magic
tech scmos
timestamp 1607758192
<< ntransistor >>
rect 11 24 13 28
rect 27 24 29 28
rect 43 24 45 28
rect 66 24 68 28
rect 71 24 73 28
rect 97 24 99 28
rect 118 24 120 28
rect 138 24 140 28
rect 143 24 145 28
rect 161 24 163 28
<< ptransistor >>
rect 11 42 13 50
rect 27 42 29 50
rect 43 42 45 50
rect 66 42 68 50
rect 71 42 73 50
rect 97 42 99 50
rect 118 42 120 50
rect 138 42 140 50
rect 143 42 145 50
rect 161 42 163 50
<< ndiffusion >>
rect 10 24 11 28
rect 13 24 14 28
rect 26 24 27 28
rect 29 24 30 28
rect 42 24 43 28
rect 45 24 46 28
rect 61 24 66 28
rect 68 24 71 28
rect 73 24 74 28
rect 95 24 97 28
rect 99 24 100 28
rect 117 24 118 28
rect 120 24 121 28
rect 133 24 138 28
rect 140 24 143 28
rect 145 24 146 28
rect 160 24 161 28
rect 163 24 164 28
<< pdiffusion >>
rect 10 42 11 50
rect 13 42 14 50
rect 26 42 27 50
rect 29 42 30 50
rect 42 42 43 50
rect 45 42 46 50
rect 61 42 66 50
rect 68 42 71 50
rect 73 42 74 50
rect 95 42 97 50
rect 99 42 100 50
rect 117 42 118 50
rect 120 42 121 50
rect 133 42 138 50
rect 140 42 143 50
rect 145 42 146 50
rect 160 42 161 50
rect 163 42 164 50
<< ndcontact >>
rect 6 24 10 28
rect 14 24 18 28
rect 22 24 26 28
rect 30 24 34 28
rect 38 24 42 28
rect 46 24 50 28
rect 57 24 61 28
rect 74 24 78 28
rect 91 24 95 28
rect 100 24 104 28
rect 113 24 117 28
rect 121 24 125 28
rect 129 24 133 28
rect 146 24 150 28
rect 156 24 160 28
rect 164 24 168 28
<< pdcontact >>
rect 6 42 10 50
rect 14 42 18 50
rect 22 42 26 50
rect 30 42 34 50
rect 38 42 42 50
rect 46 42 50 50
rect 57 42 61 50
rect 74 42 78 50
rect 91 42 95 50
rect 100 42 104 50
rect 113 42 117 50
rect 121 42 125 50
rect 129 42 133 50
rect 146 42 150 50
rect 156 42 160 50
rect 164 42 168 50
<< psubstratepcontact >>
rect -1 8 3 12
rect 17 8 22 12
rect 47 8 51 12
rect 83 8 87 12
rect 122 8 126 12
<< nsubstratencontact >>
rect -1 60 3 64
rect 17 60 22 64
rect 47 60 51 64
rect 83 60 87 64
rect 122 60 126 64
<< polysilicon >>
rect 27 57 29 60
rect 71 57 73 60
rect 97 57 99 60
rect 143 57 145 60
rect 97 53 98 57
rect 11 50 13 52
rect 27 50 29 53
rect 43 50 45 52
rect 66 50 68 52
rect 71 50 73 53
rect 97 50 99 53
rect 118 50 120 53
rect 138 50 140 52
rect 143 50 145 53
rect 161 50 163 52
rect 11 28 13 42
rect 27 40 29 42
rect 27 28 29 30
rect 43 28 45 42
rect 66 37 68 42
rect 71 40 73 42
rect 97 40 99 42
rect 62 33 68 37
rect 66 28 68 33
rect 71 28 73 30
rect 97 28 99 30
rect 118 28 120 42
rect 138 37 140 42
rect 143 40 145 42
rect 134 33 140 37
rect 138 28 140 33
rect 143 28 145 30
rect 161 28 163 42
rect 11 22 13 24
rect 27 20 29 24
rect 43 22 45 24
rect 66 22 68 24
rect 28 16 29 20
rect 71 19 73 24
rect 97 20 99 24
rect 118 22 120 24
rect 138 22 140 24
rect 27 13 29 16
rect 72 15 73 19
rect 98 16 99 20
rect 143 19 145 24
rect 161 22 163 24
rect 71 13 73 15
rect 97 12 99 16
rect 144 15 145 19
rect 143 13 145 15
<< polycontact >>
rect 27 53 31 57
rect 71 53 75 57
rect 98 53 102 57
rect 143 53 147 57
rect 7 33 11 37
rect 39 34 43 38
rect 58 33 62 37
rect 114 34 118 38
rect 130 33 134 37
rect 157 33 161 37
rect 24 16 28 20
rect 68 15 72 19
rect 93 16 98 20
rect 140 15 144 19
<< metal1 >>
rect -1 67 31 71
rect 35 67 60 71
rect 64 67 85 71
rect 89 67 149 71
rect 153 67 168 71
rect 3 60 17 64
rect 22 60 47 64
rect 51 60 83 64
rect 87 60 122 64
rect 126 60 168 64
rect 6 50 9 60
rect 38 50 41 60
rect 57 50 60 60
rect 75 53 78 57
rect 102 53 103 57
rect 113 50 116 60
rect 129 50 132 60
rect 147 53 149 57
rect 156 50 159 60
rect 2 33 7 36
rect 15 36 18 42
rect 22 36 25 42
rect 15 33 25 36
rect 15 28 18 33
rect 22 28 25 33
rect 31 38 34 42
rect 31 34 33 38
rect 37 34 39 38
rect 47 37 50 42
rect 75 39 78 42
rect 47 35 58 37
rect 31 28 34 34
rect 47 33 53 35
rect 47 28 50 33
rect 57 33 58 35
rect 76 35 78 39
rect 75 28 78 35
rect 91 38 94 42
rect 101 38 104 42
rect 101 34 110 38
rect 122 37 125 42
rect 147 38 150 42
rect 91 28 94 34
rect 101 28 104 34
rect 122 33 123 37
rect 127 33 130 36
rect 149 34 150 38
rect 122 28 125 33
rect 147 28 150 34
rect 165 28 168 42
rect 6 12 9 24
rect 38 12 41 24
rect 57 12 60 24
rect 67 15 68 19
rect 92 16 93 20
rect 113 12 116 24
rect 129 12 132 24
rect 139 15 140 19
rect 156 12 159 24
rect 3 8 17 12
rect 22 8 47 12
rect 51 8 83 12
rect 87 8 122 12
rect 126 8 168 12
rect -1 1 20 5
rect 24 1 79 5
rect 83 1 104 5
rect 108 1 135 5
rect 139 1 168 5
<< m2contact >>
rect 31 67 35 71
rect 60 67 64 71
rect 85 67 89 71
rect 149 67 153 71
rect 31 53 35 57
rect 78 53 82 57
rect 103 53 107 57
rect 149 53 153 57
rect 33 34 37 38
rect 53 31 57 35
rect 72 35 76 39
rect 91 34 95 38
rect 110 34 114 38
rect 123 33 127 37
rect 145 34 149 38
rect 153 33 157 37
rect 20 16 24 20
rect 63 15 67 19
rect 85 16 92 20
rect 135 15 139 19
rect 20 1 24 5
rect 79 1 83 5
rect 104 1 108 5
rect 135 1 139 5
<< metal2 >>
rect 32 57 35 67
rect 20 5 23 16
rect 60 15 63 67
rect 79 5 82 53
rect 85 20 88 67
rect 150 57 153 67
rect 104 5 107 53
rect 135 5 139 15
<< m3contact >>
rect 37 34 42 39
rect 52 26 57 31
rect 67 34 72 39
rect 95 34 100 39
rect 110 38 115 44
rect 140 34 145 39
rect 124 28 129 33
rect 153 28 157 33
<< metal3 >>
rect 37 40 72 45
rect 109 44 145 49
rect 36 39 43 40
rect 36 34 37 39
rect 42 34 43 39
rect 36 33 43 34
rect 66 39 73 40
rect 66 34 67 39
rect 72 34 73 39
rect 66 33 73 34
rect 94 39 101 40
rect 94 34 95 39
rect 100 34 101 39
rect 109 38 110 44
rect 115 43 145 44
rect 115 38 116 43
rect 140 40 145 43
rect 109 37 116 38
rect 139 39 146 40
rect 139 34 140 39
rect 145 34 146 39
rect 94 33 101 34
rect 123 33 130 34
rect 139 33 146 34
rect 152 33 158 34
rect 51 31 58 32
rect 51 26 52 31
rect 57 30 58 31
rect 95 30 100 33
rect 57 26 100 30
rect 123 28 124 33
rect 129 28 130 33
rect 152 28 153 33
rect 157 28 158 33
rect 123 27 158 28
rect 51 25 100 26
rect 124 23 158 27
<< labels >>
rlabel metal1 2 33 6 36 1 D
rlabel metal1 7 8 10 12 1 GND!
rlabel metal1 6 60 9 64 1 Vdd!
rlabel metal1 165 31 168 38 7 Q
rlabel metal1 -1 67 2 71 4 clk
rlabel metal1 -1 1 2 5 2 ~clk
<< end >>
