magic
tech scmos
timestamp 1608311697
<< ntransistor >>
rect 573 1706 575 1710
rect 578 1706 580 1710
rect 594 1706 596 1710
rect 610 1706 612 1710
rect 615 1706 617 1710
rect 636 1706 638 1710
rect 652 1706 654 1710
rect 668 1706 670 1710
rect 673 1706 675 1710
rect 689 1706 691 1710
rect 705 1706 707 1710
rect 710 1706 712 1710
rect 726 1706 728 1710
rect 742 1706 744 1710
rect 747 1706 749 1710
rect 768 1706 770 1710
rect 784 1706 786 1710
rect 800 1706 802 1710
rect 805 1706 807 1710
rect 821 1706 823 1710
rect 837 1706 839 1710
rect 842 1706 844 1710
rect 858 1706 860 1710
rect 874 1706 876 1710
rect 879 1706 881 1710
rect 900 1706 902 1710
rect 916 1706 918 1710
rect 932 1706 934 1710
rect 937 1706 939 1710
rect 953 1706 955 1710
rect 969 1706 971 1710
rect 974 1706 976 1710
rect 990 1706 992 1710
rect 1006 1706 1008 1710
rect 1011 1706 1013 1710
rect 1032 1706 1034 1710
rect 1048 1706 1050 1710
rect 1064 1706 1066 1710
rect 1069 1706 1071 1710
rect 1085 1706 1087 1710
rect 233 1673 235 1677
rect 238 1673 240 1677
rect 254 1673 256 1677
rect 270 1673 272 1677
rect 275 1673 277 1677
rect 296 1673 298 1677
rect 312 1673 314 1677
rect 328 1673 330 1677
rect 333 1673 335 1677
rect 349 1673 351 1677
rect 357 1636 359 1640
rect 752 1640 754 1644
rect 778 1636 780 1640
rect 783 1636 785 1640
rect 833 1640 835 1644
rect 859 1636 861 1640
rect 864 1636 866 1640
rect 806 1632 808 1636
rect 240 1627 242 1631
rect 578 1627 580 1631
rect 594 1627 596 1631
rect 610 1627 612 1631
rect 633 1627 635 1631
rect 638 1627 640 1631
rect 664 1627 666 1631
rect 685 1627 687 1631
rect 705 1627 707 1631
rect 710 1627 712 1631
rect 728 1627 730 1631
rect 887 1632 889 1636
rect 578 1581 580 1585
rect 594 1581 596 1585
rect 610 1581 612 1585
rect 633 1581 635 1585
rect 638 1581 640 1585
rect 664 1581 666 1585
rect 685 1581 687 1585
rect 705 1581 707 1585
rect 710 1581 712 1585
rect 728 1581 730 1585
rect 224 1571 226 1575
rect 240 1571 242 1575
rect 245 1571 247 1575
rect 261 1571 263 1575
rect 277 1571 279 1575
rect 298 1571 300 1575
rect 303 1571 305 1575
rect 319 1571 321 1575
rect 335 1571 337 1575
rect 340 1571 342 1575
rect 778 1580 780 1584
rect 783 1580 785 1584
rect 859 1580 861 1584
rect 864 1580 866 1584
rect 778 1504 780 1508
rect 783 1504 785 1508
rect 857 1508 859 1512
rect 883 1504 885 1508
rect 888 1504 890 1508
rect 806 1500 808 1504
rect 578 1495 580 1499
rect 594 1495 596 1499
rect 610 1495 612 1499
rect 633 1495 635 1499
rect 638 1495 640 1499
rect 664 1495 666 1499
rect 685 1495 687 1499
rect 705 1495 707 1499
rect 710 1495 712 1499
rect 728 1495 730 1499
rect 911 1500 913 1504
rect 578 1449 580 1453
rect 594 1449 596 1453
rect 610 1449 612 1453
rect 633 1449 635 1453
rect 638 1449 640 1453
rect 664 1449 666 1453
rect 685 1449 687 1453
rect 705 1449 707 1453
rect 710 1449 712 1453
rect 728 1449 730 1453
rect 778 1449 780 1453
rect 783 1449 785 1453
rect 883 1449 885 1453
rect 888 1449 890 1453
rect 778 1372 780 1376
rect 783 1372 785 1376
rect 833 1376 835 1380
rect 859 1372 861 1376
rect 864 1372 866 1376
rect 923 1376 925 1380
rect 949 1372 951 1376
rect 954 1372 956 1376
rect 806 1368 808 1372
rect 578 1363 580 1367
rect 594 1363 596 1367
rect 610 1363 612 1367
rect 633 1363 635 1367
rect 638 1363 640 1367
rect 664 1363 666 1367
rect 685 1363 687 1367
rect 705 1363 707 1367
rect 710 1363 712 1367
rect 728 1363 730 1367
rect 887 1368 889 1372
rect 977 1368 979 1372
rect 578 1317 580 1321
rect 594 1317 596 1321
rect 610 1317 612 1321
rect 633 1317 635 1321
rect 638 1317 640 1321
rect 664 1317 666 1321
rect 685 1317 687 1321
rect 705 1317 707 1321
rect 710 1317 712 1321
rect 728 1317 730 1321
rect 778 1314 780 1318
rect 783 1314 785 1318
rect 859 1314 861 1318
rect 864 1314 866 1318
rect 949 1314 951 1318
rect 954 1314 956 1318
rect 778 1240 780 1244
rect 783 1240 785 1244
rect 806 1236 808 1240
rect 578 1231 580 1235
rect 594 1231 596 1235
rect 610 1231 612 1235
rect 633 1231 635 1235
rect 638 1231 640 1235
rect 664 1231 666 1235
rect 685 1231 687 1235
rect 705 1231 707 1235
rect 710 1231 712 1235
rect 728 1231 730 1235
rect 578 1185 580 1189
rect 594 1185 596 1189
rect 610 1185 612 1189
rect 633 1185 635 1189
rect 638 1185 640 1189
rect 664 1185 666 1189
rect 685 1185 687 1189
rect 705 1185 707 1189
rect 710 1185 712 1189
rect 728 1185 730 1189
rect 812 1185 814 1189
rect 830 1185 832 1189
rect 855 1185 857 1189
rect 871 1185 873 1189
rect 894 1185 896 1189
rect 899 1185 901 1189
rect 925 1185 927 1189
rect 946 1185 948 1189
rect 966 1185 968 1189
rect 971 1185 973 1189
rect 989 1185 991 1189
rect 101 1171 103 1175
rect 106 1171 108 1175
rect 122 1171 124 1175
rect 138 1171 140 1175
rect 143 1171 145 1175
rect 164 1171 166 1175
rect 180 1171 182 1175
rect 196 1171 198 1175
rect 201 1171 203 1175
rect 217 1171 219 1175
rect 233 1171 235 1175
rect 238 1171 240 1175
rect 254 1171 256 1175
rect 270 1171 272 1175
rect 275 1171 277 1175
rect 296 1171 298 1175
rect 312 1171 314 1175
rect 328 1171 330 1175
rect 333 1171 335 1175
rect 349 1171 351 1175
rect 365 1171 367 1175
rect 370 1171 372 1175
rect 386 1171 388 1175
rect 402 1171 404 1175
rect 407 1171 409 1175
rect 428 1171 430 1175
rect 444 1171 446 1175
rect 460 1171 462 1175
rect 465 1171 467 1175
rect 481 1171 483 1175
rect 778 1178 780 1182
rect 783 1178 785 1182
rect 216 1127 218 1131
rect 240 1127 242 1131
rect 1001 1129 1005 1131
rect 236 1116 238 1120
rect 227 1102 231 1104
rect 216 1093 218 1097
rect 240 1093 242 1097
rect 872 1061 874 1065
rect 877 1061 879 1065
rect 893 1061 895 1065
rect 909 1061 911 1065
rect 914 1061 916 1065
rect 935 1061 937 1065
rect 951 1061 953 1065
rect 967 1061 969 1065
rect 972 1061 974 1065
rect 988 1061 990 1065
rect 101 1031 103 1035
rect 106 1031 108 1035
rect 122 1031 124 1035
rect 138 1031 140 1035
rect 143 1031 145 1035
rect 164 1031 166 1035
rect 180 1031 182 1035
rect 196 1031 198 1035
rect 201 1031 203 1035
rect 217 1031 219 1035
rect 233 1031 235 1035
rect 238 1031 240 1035
rect 254 1031 256 1035
rect 270 1031 272 1035
rect 275 1031 277 1035
rect 296 1031 298 1035
rect 312 1031 314 1035
rect 328 1031 330 1035
rect 333 1031 335 1035
rect 349 1031 351 1035
rect 365 1031 367 1035
rect 370 1031 372 1035
rect 386 1031 388 1035
rect 402 1031 404 1035
rect 407 1031 409 1035
rect 428 1031 430 1035
rect 444 1031 446 1035
rect 460 1031 462 1035
rect 465 1031 467 1035
rect 481 1031 483 1035
rect 1013 985 1017 987
rect 872 975 874 979
rect 877 975 879 979
rect 893 975 895 979
rect 909 975 911 979
rect 914 975 916 979
rect 935 975 937 979
rect 951 975 953 979
rect 967 975 969 979
rect 972 975 974 979
rect 988 975 990 979
rect 101 945 103 949
rect 106 945 108 949
rect 122 945 124 949
rect 138 945 140 949
rect 143 945 145 949
rect 164 945 166 949
rect 180 945 182 949
rect 196 945 198 949
rect 201 945 203 949
rect 217 945 219 949
rect 233 945 235 949
rect 238 945 240 949
rect 254 945 256 949
rect 270 945 272 949
rect 275 945 277 949
rect 296 945 298 949
rect 312 945 314 949
rect 328 945 330 949
rect 333 945 335 949
rect 349 945 351 949
rect 365 945 367 949
rect 370 945 372 949
rect 386 945 388 949
rect 402 945 404 949
rect 407 945 409 949
rect 428 945 430 949
rect 444 945 446 949
rect 460 945 462 949
rect 465 945 467 949
rect 481 945 483 949
rect 333 901 335 905
rect 357 901 359 905
rect 353 890 355 894
rect 344 876 348 878
rect 333 867 335 871
rect 357 867 359 871
rect 101 805 103 809
rect 106 805 108 809
rect 122 805 124 809
rect 138 805 140 809
rect 143 805 145 809
rect 164 805 166 809
rect 180 805 182 809
rect 196 805 198 809
rect 201 805 203 809
rect 217 805 219 809
rect 233 805 235 809
rect 238 805 240 809
rect 254 805 256 809
rect 270 805 272 809
rect 275 805 277 809
rect 296 805 298 809
rect 312 805 314 809
rect 328 805 330 809
rect 333 805 335 809
rect 349 805 351 809
rect 365 805 367 809
rect 370 805 372 809
rect 386 805 388 809
rect 402 805 404 809
rect 407 805 409 809
rect 428 805 430 809
rect 444 805 446 809
rect 460 805 462 809
rect 465 805 467 809
rect 481 805 483 809
<< ptransistor >>
rect 573 1729 575 1737
rect 578 1729 580 1737
rect 594 1729 596 1737
rect 610 1729 612 1737
rect 615 1729 617 1737
rect 636 1729 638 1737
rect 652 1729 654 1737
rect 668 1729 670 1737
rect 673 1729 675 1737
rect 689 1729 691 1737
rect 705 1729 707 1737
rect 710 1729 712 1737
rect 726 1729 728 1737
rect 742 1729 744 1737
rect 747 1729 749 1737
rect 768 1729 770 1737
rect 784 1729 786 1737
rect 800 1729 802 1737
rect 805 1729 807 1737
rect 821 1729 823 1737
rect 837 1729 839 1737
rect 842 1729 844 1737
rect 858 1729 860 1737
rect 874 1729 876 1737
rect 879 1729 881 1737
rect 900 1729 902 1737
rect 916 1729 918 1737
rect 932 1729 934 1737
rect 937 1729 939 1737
rect 953 1729 955 1737
rect 969 1729 971 1737
rect 974 1729 976 1737
rect 990 1729 992 1737
rect 1006 1729 1008 1737
rect 1011 1729 1013 1737
rect 1032 1729 1034 1737
rect 1048 1729 1050 1737
rect 1064 1729 1066 1737
rect 1069 1729 1071 1737
rect 1085 1729 1087 1737
rect 233 1696 235 1704
rect 238 1696 240 1704
rect 254 1696 256 1704
rect 270 1696 272 1704
rect 275 1696 277 1704
rect 296 1696 298 1704
rect 312 1696 314 1704
rect 328 1696 330 1704
rect 333 1696 335 1704
rect 349 1696 351 1704
rect 752 1658 754 1666
rect 578 1645 580 1653
rect 594 1645 596 1653
rect 610 1645 612 1653
rect 633 1645 635 1653
rect 638 1645 640 1653
rect 664 1645 666 1653
rect 685 1645 687 1653
rect 705 1645 707 1653
rect 710 1645 712 1653
rect 728 1645 730 1653
rect 778 1652 780 1660
rect 783 1652 785 1660
rect 806 1658 808 1666
rect 833 1658 835 1666
rect 859 1652 861 1660
rect 864 1652 866 1660
rect 887 1658 889 1666
rect 224 1594 226 1602
rect 240 1594 242 1602
rect 245 1594 247 1602
rect 261 1594 263 1602
rect 277 1594 279 1602
rect 298 1594 300 1602
rect 303 1594 305 1602
rect 319 1594 321 1602
rect 335 1594 337 1602
rect 340 1594 342 1602
rect 578 1559 580 1567
rect 594 1559 596 1567
rect 610 1559 612 1567
rect 633 1559 635 1567
rect 638 1559 640 1567
rect 664 1559 666 1567
rect 685 1559 687 1567
rect 705 1559 707 1567
rect 710 1559 712 1567
rect 728 1559 730 1567
rect 778 1560 780 1568
rect 783 1560 785 1568
rect 859 1560 861 1568
rect 864 1560 866 1568
rect 578 1513 580 1521
rect 594 1513 596 1521
rect 610 1513 612 1521
rect 633 1513 635 1521
rect 638 1513 640 1521
rect 664 1513 666 1521
rect 685 1513 687 1521
rect 705 1513 707 1521
rect 710 1513 712 1521
rect 728 1513 730 1521
rect 778 1520 780 1528
rect 783 1520 785 1528
rect 806 1526 808 1534
rect 857 1526 859 1534
rect 883 1520 885 1528
rect 888 1520 890 1528
rect 911 1526 913 1534
rect 578 1427 580 1435
rect 594 1427 596 1435
rect 610 1427 612 1435
rect 633 1427 635 1435
rect 638 1427 640 1435
rect 664 1427 666 1435
rect 685 1427 687 1435
rect 705 1427 707 1435
rect 710 1427 712 1435
rect 728 1427 730 1435
rect 778 1429 780 1437
rect 783 1429 785 1437
rect 883 1429 885 1437
rect 888 1429 890 1437
rect 578 1381 580 1389
rect 594 1381 596 1389
rect 610 1381 612 1389
rect 633 1381 635 1389
rect 638 1381 640 1389
rect 664 1381 666 1389
rect 685 1381 687 1389
rect 705 1381 707 1389
rect 710 1381 712 1389
rect 728 1381 730 1389
rect 778 1388 780 1396
rect 783 1388 785 1396
rect 806 1394 808 1402
rect 833 1394 835 1402
rect 859 1388 861 1396
rect 864 1388 866 1396
rect 887 1394 889 1402
rect 923 1394 925 1402
rect 949 1388 951 1396
rect 954 1388 956 1396
rect 977 1394 979 1402
rect 578 1295 580 1303
rect 594 1295 596 1303
rect 610 1295 612 1303
rect 633 1295 635 1303
rect 638 1295 640 1303
rect 664 1295 666 1303
rect 685 1295 687 1303
rect 705 1295 707 1303
rect 710 1295 712 1303
rect 728 1295 730 1303
rect 778 1294 780 1302
rect 783 1294 785 1302
rect 859 1294 861 1302
rect 864 1294 866 1302
rect 949 1294 951 1302
rect 954 1294 956 1302
rect 578 1249 580 1257
rect 594 1249 596 1257
rect 610 1249 612 1257
rect 633 1249 635 1257
rect 638 1249 640 1257
rect 664 1249 666 1257
rect 685 1249 687 1257
rect 705 1249 707 1257
rect 710 1249 712 1257
rect 728 1249 730 1257
rect 778 1256 780 1264
rect 783 1256 785 1264
rect 806 1262 808 1270
rect 101 1194 103 1202
rect 106 1194 108 1202
rect 122 1194 124 1202
rect 138 1194 140 1202
rect 143 1194 145 1202
rect 164 1194 166 1202
rect 180 1194 182 1202
rect 196 1194 198 1202
rect 201 1194 203 1202
rect 217 1194 219 1202
rect 233 1194 235 1202
rect 238 1194 240 1202
rect 254 1194 256 1202
rect 270 1194 272 1202
rect 275 1194 277 1202
rect 296 1194 298 1202
rect 312 1194 314 1202
rect 328 1194 330 1202
rect 333 1194 335 1202
rect 349 1194 351 1202
rect 365 1194 367 1202
rect 370 1194 372 1202
rect 386 1194 388 1202
rect 402 1194 404 1202
rect 407 1194 409 1202
rect 428 1194 430 1202
rect 444 1194 446 1202
rect 460 1194 462 1202
rect 465 1194 467 1202
rect 481 1194 483 1202
rect 578 1163 580 1171
rect 594 1163 596 1171
rect 610 1163 612 1171
rect 633 1163 635 1171
rect 638 1163 640 1171
rect 664 1163 666 1171
rect 685 1163 687 1171
rect 705 1163 707 1171
rect 710 1163 712 1171
rect 728 1163 730 1171
rect 778 1158 780 1166
rect 783 1158 785 1166
rect 812 1163 814 1171
rect 830 1163 832 1171
rect 855 1163 857 1171
rect 871 1163 873 1171
rect 894 1163 896 1171
rect 899 1163 901 1171
rect 925 1163 927 1171
rect 946 1163 948 1171
rect 966 1163 968 1171
rect 971 1163 973 1171
rect 989 1163 991 1171
rect 872 1084 874 1092
rect 877 1084 879 1092
rect 893 1084 895 1092
rect 909 1084 911 1092
rect 914 1084 916 1092
rect 935 1084 937 1092
rect 951 1084 953 1092
rect 967 1084 969 1092
rect 972 1084 974 1092
rect 988 1084 990 1092
rect 101 1054 103 1062
rect 106 1054 108 1062
rect 122 1054 124 1062
rect 138 1054 140 1062
rect 143 1054 145 1062
rect 164 1054 166 1062
rect 180 1054 182 1062
rect 196 1054 198 1062
rect 201 1054 203 1062
rect 217 1054 219 1062
rect 233 1054 235 1062
rect 238 1054 240 1062
rect 254 1054 256 1062
rect 270 1054 272 1062
rect 275 1054 277 1062
rect 296 1054 298 1062
rect 312 1054 314 1062
rect 328 1054 330 1062
rect 333 1054 335 1062
rect 349 1054 351 1062
rect 365 1054 367 1062
rect 370 1054 372 1062
rect 386 1054 388 1062
rect 402 1054 404 1062
rect 407 1054 409 1062
rect 428 1054 430 1062
rect 444 1054 446 1062
rect 460 1054 462 1062
rect 465 1054 467 1062
rect 481 1054 483 1062
rect 872 998 874 1006
rect 877 998 879 1006
rect 893 998 895 1006
rect 909 998 911 1006
rect 914 998 916 1006
rect 935 998 937 1006
rect 951 998 953 1006
rect 967 998 969 1006
rect 972 998 974 1006
rect 988 998 990 1006
rect 101 968 103 976
rect 106 968 108 976
rect 122 968 124 976
rect 138 968 140 976
rect 143 968 145 976
rect 164 968 166 976
rect 180 968 182 976
rect 196 968 198 976
rect 201 968 203 976
rect 217 968 219 976
rect 233 968 235 976
rect 238 968 240 976
rect 254 968 256 976
rect 270 968 272 976
rect 275 968 277 976
rect 296 968 298 976
rect 312 968 314 976
rect 328 968 330 976
rect 333 968 335 976
rect 349 968 351 976
rect 365 968 367 976
rect 370 968 372 976
rect 386 968 388 976
rect 402 968 404 976
rect 407 968 409 976
rect 428 968 430 976
rect 444 968 446 976
rect 460 968 462 976
rect 465 968 467 976
rect 481 968 483 976
rect 101 828 103 836
rect 106 828 108 836
rect 122 828 124 836
rect 138 828 140 836
rect 143 828 145 836
rect 164 828 166 836
rect 180 828 182 836
rect 196 828 198 836
rect 201 828 203 836
rect 217 828 219 836
rect 233 828 235 836
rect 238 828 240 836
rect 254 828 256 836
rect 270 828 272 836
rect 275 828 277 836
rect 296 828 298 836
rect 312 828 314 836
rect 328 828 330 836
rect 333 828 335 836
rect 349 828 351 836
rect 365 828 367 836
rect 370 828 372 836
rect 386 828 388 836
rect 402 828 404 836
rect 407 828 409 836
rect 428 828 430 836
rect 444 828 446 836
rect 460 828 462 836
rect 465 828 467 836
rect 481 828 483 836
<< ndiffusion >>
rect 572 1706 573 1710
rect 575 1706 578 1710
rect 580 1706 581 1710
rect 593 1706 594 1710
rect 596 1706 597 1710
rect 609 1706 610 1710
rect 612 1706 615 1710
rect 617 1706 618 1710
rect 635 1706 636 1710
rect 638 1706 639 1710
rect 651 1706 652 1710
rect 654 1706 655 1710
rect 667 1706 668 1710
rect 670 1706 673 1710
rect 675 1706 676 1710
rect 688 1706 689 1710
rect 691 1706 692 1710
rect 704 1706 705 1710
rect 707 1706 710 1710
rect 712 1706 713 1710
rect 725 1706 726 1710
rect 728 1706 729 1710
rect 741 1706 742 1710
rect 744 1706 747 1710
rect 749 1706 750 1710
rect 767 1706 768 1710
rect 770 1706 771 1710
rect 783 1706 784 1710
rect 786 1706 787 1710
rect 799 1706 800 1710
rect 802 1706 805 1710
rect 807 1706 808 1710
rect 820 1706 821 1710
rect 823 1706 824 1710
rect 836 1706 837 1710
rect 839 1706 842 1710
rect 844 1706 845 1710
rect 857 1706 858 1710
rect 860 1706 861 1710
rect 873 1706 874 1710
rect 876 1706 879 1710
rect 881 1706 882 1710
rect 899 1706 900 1710
rect 902 1706 903 1710
rect 915 1706 916 1710
rect 918 1706 919 1710
rect 931 1706 932 1710
rect 934 1706 937 1710
rect 939 1706 940 1710
rect 952 1706 953 1710
rect 955 1706 956 1710
rect 968 1706 969 1710
rect 971 1706 974 1710
rect 976 1706 977 1710
rect 989 1706 990 1710
rect 992 1706 993 1710
rect 1005 1706 1006 1710
rect 1008 1706 1011 1710
rect 1013 1706 1014 1710
rect 1031 1706 1032 1710
rect 1034 1706 1035 1710
rect 1047 1706 1048 1710
rect 1050 1706 1051 1710
rect 1063 1706 1064 1710
rect 1066 1706 1069 1710
rect 1071 1706 1072 1710
rect 1084 1706 1085 1710
rect 1087 1706 1088 1710
rect 232 1673 233 1677
rect 235 1673 238 1677
rect 240 1673 241 1677
rect 253 1673 254 1677
rect 256 1673 257 1677
rect 269 1673 270 1677
rect 272 1673 275 1677
rect 277 1673 278 1677
rect 295 1673 296 1677
rect 298 1673 299 1677
rect 311 1673 312 1677
rect 314 1673 315 1677
rect 327 1673 328 1677
rect 330 1673 333 1677
rect 335 1673 336 1677
rect 348 1673 349 1677
rect 351 1673 352 1677
rect 356 1636 357 1640
rect 359 1636 360 1640
rect 751 1640 752 1644
rect 754 1640 755 1644
rect 775 1636 778 1640
rect 780 1636 783 1640
rect 785 1636 786 1640
rect 832 1640 833 1644
rect 835 1640 836 1644
rect 856 1636 859 1640
rect 861 1636 864 1640
rect 866 1636 867 1640
rect 805 1632 806 1636
rect 808 1632 809 1636
rect 239 1627 240 1631
rect 242 1627 243 1631
rect 577 1627 578 1631
rect 580 1627 581 1631
rect 593 1627 594 1631
rect 596 1627 597 1631
rect 609 1627 610 1631
rect 612 1627 613 1631
rect 628 1627 633 1631
rect 635 1627 638 1631
rect 640 1627 641 1631
rect 662 1627 664 1631
rect 666 1627 667 1631
rect 684 1627 685 1631
rect 687 1627 688 1631
rect 700 1627 705 1631
rect 707 1627 710 1631
rect 712 1627 713 1631
rect 727 1627 728 1631
rect 730 1627 731 1631
rect 886 1632 887 1636
rect 889 1632 890 1636
rect 577 1581 578 1585
rect 580 1581 581 1585
rect 593 1581 594 1585
rect 596 1581 597 1585
rect 609 1581 610 1585
rect 612 1581 613 1585
rect 628 1581 633 1585
rect 635 1581 638 1585
rect 640 1581 641 1585
rect 662 1581 664 1585
rect 666 1581 667 1585
rect 684 1581 685 1585
rect 687 1581 688 1585
rect 700 1581 705 1585
rect 707 1581 710 1585
rect 712 1581 713 1585
rect 727 1581 728 1585
rect 730 1581 731 1585
rect 223 1571 224 1575
rect 226 1571 227 1575
rect 239 1571 240 1575
rect 242 1571 245 1575
rect 247 1571 248 1575
rect 260 1571 261 1575
rect 263 1571 264 1575
rect 276 1571 277 1575
rect 279 1571 280 1575
rect 297 1571 298 1575
rect 300 1571 303 1575
rect 305 1571 306 1575
rect 318 1571 319 1575
rect 321 1571 322 1575
rect 334 1571 335 1575
rect 337 1571 340 1575
rect 342 1571 343 1575
rect 775 1580 778 1584
rect 780 1580 783 1584
rect 785 1580 786 1584
rect 856 1580 859 1584
rect 861 1580 864 1584
rect 866 1580 867 1584
rect 775 1504 778 1508
rect 780 1504 783 1508
rect 785 1504 786 1508
rect 856 1508 857 1512
rect 859 1508 860 1512
rect 880 1504 883 1508
rect 885 1504 888 1508
rect 890 1504 891 1508
rect 805 1500 806 1504
rect 808 1500 809 1504
rect 577 1495 578 1499
rect 580 1495 581 1499
rect 593 1495 594 1499
rect 596 1495 597 1499
rect 609 1495 610 1499
rect 612 1495 613 1499
rect 628 1495 633 1499
rect 635 1495 638 1499
rect 640 1495 641 1499
rect 662 1495 664 1499
rect 666 1495 667 1499
rect 684 1495 685 1499
rect 687 1495 688 1499
rect 700 1495 705 1499
rect 707 1495 710 1499
rect 712 1495 713 1499
rect 727 1495 728 1499
rect 730 1495 731 1499
rect 910 1500 911 1504
rect 913 1500 914 1504
rect 577 1449 578 1453
rect 580 1449 581 1453
rect 593 1449 594 1453
rect 596 1449 597 1453
rect 609 1449 610 1453
rect 612 1449 613 1453
rect 628 1449 633 1453
rect 635 1449 638 1453
rect 640 1449 641 1453
rect 662 1449 664 1453
rect 666 1449 667 1453
rect 684 1449 685 1453
rect 687 1449 688 1453
rect 700 1449 705 1453
rect 707 1449 710 1453
rect 712 1449 713 1453
rect 727 1449 728 1453
rect 730 1449 731 1453
rect 775 1449 778 1453
rect 780 1449 783 1453
rect 785 1449 786 1453
rect 880 1449 883 1453
rect 885 1449 888 1453
rect 890 1449 891 1453
rect 775 1372 778 1376
rect 780 1372 783 1376
rect 785 1372 786 1376
rect 832 1376 833 1380
rect 835 1376 836 1380
rect 856 1372 859 1376
rect 861 1372 864 1376
rect 866 1372 867 1376
rect 922 1376 923 1380
rect 925 1376 926 1380
rect 946 1372 949 1376
rect 951 1372 954 1376
rect 956 1372 957 1376
rect 805 1368 806 1372
rect 808 1368 809 1372
rect 577 1363 578 1367
rect 580 1363 581 1367
rect 593 1363 594 1367
rect 596 1363 597 1367
rect 609 1363 610 1367
rect 612 1363 613 1367
rect 628 1363 633 1367
rect 635 1363 638 1367
rect 640 1363 641 1367
rect 662 1363 664 1367
rect 666 1363 667 1367
rect 684 1363 685 1367
rect 687 1363 688 1367
rect 700 1363 705 1367
rect 707 1363 710 1367
rect 712 1363 713 1367
rect 727 1363 728 1367
rect 730 1363 731 1367
rect 886 1368 887 1372
rect 889 1368 890 1372
rect 976 1368 977 1372
rect 979 1368 980 1372
rect 577 1317 578 1321
rect 580 1317 581 1321
rect 593 1317 594 1321
rect 596 1317 597 1321
rect 609 1317 610 1321
rect 612 1317 613 1321
rect 628 1317 633 1321
rect 635 1317 638 1321
rect 640 1317 641 1321
rect 662 1317 664 1321
rect 666 1317 667 1321
rect 684 1317 685 1321
rect 687 1317 688 1321
rect 700 1317 705 1321
rect 707 1317 710 1321
rect 712 1317 713 1321
rect 727 1317 728 1321
rect 730 1317 731 1321
rect 775 1314 778 1318
rect 780 1314 783 1318
rect 785 1314 786 1318
rect 856 1314 859 1318
rect 861 1314 864 1318
rect 866 1314 867 1318
rect 946 1314 949 1318
rect 951 1314 954 1318
rect 956 1314 957 1318
rect 775 1240 778 1244
rect 780 1240 783 1244
rect 785 1240 786 1244
rect 805 1236 806 1240
rect 808 1236 809 1240
rect 577 1231 578 1235
rect 580 1231 581 1235
rect 593 1231 594 1235
rect 596 1231 597 1235
rect 609 1231 610 1235
rect 612 1231 613 1235
rect 628 1231 633 1235
rect 635 1231 638 1235
rect 640 1231 641 1235
rect 662 1231 664 1235
rect 666 1231 667 1235
rect 684 1231 685 1235
rect 687 1231 688 1235
rect 700 1231 705 1235
rect 707 1231 710 1235
rect 712 1231 713 1235
rect 727 1231 728 1235
rect 730 1231 731 1235
rect 577 1185 578 1189
rect 580 1185 581 1189
rect 593 1185 594 1189
rect 596 1185 597 1189
rect 609 1185 610 1189
rect 612 1185 613 1189
rect 628 1185 633 1189
rect 635 1185 638 1189
rect 640 1185 641 1189
rect 662 1185 664 1189
rect 666 1185 667 1189
rect 684 1185 685 1189
rect 687 1185 688 1189
rect 700 1185 705 1189
rect 707 1185 710 1189
rect 712 1185 713 1189
rect 727 1185 728 1189
rect 730 1185 731 1189
rect 811 1185 812 1189
rect 814 1185 815 1189
rect 819 1185 825 1189
rect 829 1185 830 1189
rect 832 1185 833 1189
rect 854 1185 855 1189
rect 857 1185 858 1189
rect 870 1185 871 1189
rect 873 1185 874 1189
rect 889 1185 894 1189
rect 896 1185 899 1189
rect 901 1185 902 1189
rect 923 1185 925 1189
rect 927 1185 928 1189
rect 945 1185 946 1189
rect 948 1185 949 1189
rect 961 1185 966 1189
rect 968 1185 971 1189
rect 973 1185 974 1189
rect 988 1185 989 1189
rect 991 1185 992 1189
rect 100 1171 101 1175
rect 103 1171 106 1175
rect 108 1171 109 1175
rect 121 1171 122 1175
rect 124 1171 125 1175
rect 137 1171 138 1175
rect 140 1171 143 1175
rect 145 1171 146 1175
rect 163 1171 164 1175
rect 166 1171 167 1175
rect 179 1171 180 1175
rect 182 1171 183 1175
rect 195 1171 196 1175
rect 198 1171 201 1175
rect 203 1171 204 1175
rect 216 1171 217 1175
rect 219 1171 220 1175
rect 232 1171 233 1175
rect 235 1171 238 1175
rect 240 1171 241 1175
rect 253 1171 254 1175
rect 256 1171 257 1175
rect 269 1171 270 1175
rect 272 1171 275 1175
rect 277 1171 278 1175
rect 295 1171 296 1175
rect 298 1171 299 1175
rect 311 1171 312 1175
rect 314 1171 315 1175
rect 327 1171 328 1175
rect 330 1171 333 1175
rect 335 1171 336 1175
rect 348 1171 349 1175
rect 351 1171 352 1175
rect 364 1171 365 1175
rect 367 1171 370 1175
rect 372 1171 373 1175
rect 385 1171 386 1175
rect 388 1171 389 1175
rect 401 1171 402 1175
rect 404 1171 407 1175
rect 409 1171 410 1175
rect 427 1171 428 1175
rect 430 1171 431 1175
rect 443 1171 444 1175
rect 446 1171 447 1175
rect 459 1171 460 1175
rect 462 1171 465 1175
rect 467 1171 468 1175
rect 480 1171 481 1175
rect 483 1171 484 1175
rect 775 1178 778 1182
rect 780 1178 783 1182
rect 785 1178 786 1182
rect 215 1127 216 1131
rect 218 1127 219 1131
rect 239 1127 240 1131
rect 242 1127 243 1131
rect 1001 1131 1005 1132
rect 1001 1128 1005 1129
rect 235 1116 236 1120
rect 238 1116 239 1120
rect 227 1104 231 1105
rect 227 1101 231 1102
rect 215 1093 216 1097
rect 218 1093 219 1097
rect 239 1093 240 1097
rect 242 1093 243 1097
rect 871 1061 872 1065
rect 874 1061 877 1065
rect 879 1061 880 1065
rect 892 1061 893 1065
rect 895 1061 896 1065
rect 908 1061 909 1065
rect 911 1061 914 1065
rect 916 1061 917 1065
rect 934 1061 935 1065
rect 937 1061 938 1065
rect 950 1061 951 1065
rect 953 1061 954 1065
rect 966 1061 967 1065
rect 969 1061 972 1065
rect 974 1061 975 1065
rect 987 1061 988 1065
rect 990 1061 991 1065
rect 100 1031 101 1035
rect 103 1031 106 1035
rect 108 1031 109 1035
rect 121 1031 122 1035
rect 124 1031 125 1035
rect 137 1031 138 1035
rect 140 1031 143 1035
rect 145 1031 146 1035
rect 163 1031 164 1035
rect 166 1031 167 1035
rect 179 1031 180 1035
rect 182 1031 183 1035
rect 195 1031 196 1035
rect 198 1031 201 1035
rect 203 1031 204 1035
rect 216 1031 217 1035
rect 219 1031 220 1035
rect 232 1031 233 1035
rect 235 1031 238 1035
rect 240 1031 241 1035
rect 253 1031 254 1035
rect 256 1031 257 1035
rect 269 1031 270 1035
rect 272 1031 275 1035
rect 277 1031 278 1035
rect 295 1031 296 1035
rect 298 1031 299 1035
rect 311 1031 312 1035
rect 314 1031 315 1035
rect 327 1031 328 1035
rect 330 1031 333 1035
rect 335 1031 336 1035
rect 348 1031 349 1035
rect 351 1031 352 1035
rect 364 1031 365 1035
rect 367 1031 370 1035
rect 372 1031 373 1035
rect 385 1031 386 1035
rect 388 1031 389 1035
rect 401 1031 402 1035
rect 404 1031 407 1035
rect 409 1031 410 1035
rect 427 1031 428 1035
rect 430 1031 431 1035
rect 443 1031 444 1035
rect 446 1031 447 1035
rect 459 1031 460 1035
rect 462 1031 465 1035
rect 467 1031 468 1035
rect 480 1031 481 1035
rect 483 1031 484 1035
rect 1013 987 1017 988
rect 1013 984 1017 985
rect 871 975 872 979
rect 874 975 877 979
rect 879 975 880 979
rect 892 975 893 979
rect 895 975 896 979
rect 908 975 909 979
rect 911 975 914 979
rect 916 975 917 979
rect 934 975 935 979
rect 937 975 938 979
rect 950 975 951 979
rect 953 975 954 979
rect 966 975 967 979
rect 969 975 972 979
rect 974 975 975 979
rect 987 975 988 979
rect 990 975 991 979
rect 100 945 101 949
rect 103 945 106 949
rect 108 945 109 949
rect 121 945 122 949
rect 124 945 125 949
rect 137 945 138 949
rect 140 945 143 949
rect 145 945 146 949
rect 163 945 164 949
rect 166 945 167 949
rect 179 945 180 949
rect 182 945 183 949
rect 195 945 196 949
rect 198 945 201 949
rect 203 945 204 949
rect 216 945 217 949
rect 219 945 220 949
rect 232 945 233 949
rect 235 945 238 949
rect 240 945 241 949
rect 253 945 254 949
rect 256 945 257 949
rect 269 945 270 949
rect 272 945 275 949
rect 277 945 278 949
rect 295 945 296 949
rect 298 945 299 949
rect 311 945 312 949
rect 314 945 315 949
rect 327 945 328 949
rect 330 945 333 949
rect 335 945 336 949
rect 348 945 349 949
rect 351 945 352 949
rect 364 945 365 949
rect 367 945 370 949
rect 372 945 373 949
rect 385 945 386 949
rect 388 945 389 949
rect 401 945 402 949
rect 404 945 407 949
rect 409 945 410 949
rect 427 945 428 949
rect 430 945 431 949
rect 443 945 444 949
rect 446 945 447 949
rect 459 945 460 949
rect 462 945 465 949
rect 467 945 468 949
rect 480 945 481 949
rect 483 945 484 949
rect 332 901 333 905
rect 335 901 336 905
rect 356 901 357 905
rect 359 901 360 905
rect 352 890 353 894
rect 355 890 356 894
rect 344 878 348 879
rect 344 875 348 876
rect 332 867 333 871
rect 335 867 336 871
rect 356 867 357 871
rect 359 867 360 871
rect 100 805 101 809
rect 103 805 106 809
rect 108 805 109 809
rect 121 805 122 809
rect 124 805 125 809
rect 137 805 138 809
rect 140 805 143 809
rect 145 805 146 809
rect 163 805 164 809
rect 166 805 167 809
rect 179 805 180 809
rect 182 805 183 809
rect 195 805 196 809
rect 198 805 201 809
rect 203 805 204 809
rect 216 805 217 809
rect 219 805 220 809
rect 232 805 233 809
rect 235 805 238 809
rect 240 805 241 809
rect 253 805 254 809
rect 256 805 257 809
rect 269 805 270 809
rect 272 805 275 809
rect 277 805 278 809
rect 295 805 296 809
rect 298 805 299 809
rect 311 805 312 809
rect 314 805 315 809
rect 327 805 328 809
rect 330 805 333 809
rect 335 805 336 809
rect 348 805 349 809
rect 351 805 352 809
rect 364 805 365 809
rect 367 805 370 809
rect 372 805 373 809
rect 385 805 386 809
rect 388 805 389 809
rect 401 805 402 809
rect 404 805 407 809
rect 409 805 410 809
rect 427 805 428 809
rect 430 805 431 809
rect 443 805 444 809
rect 446 805 447 809
rect 459 805 460 809
rect 462 805 465 809
rect 467 805 468 809
rect 480 805 481 809
rect 483 805 484 809
<< pdiffusion >>
rect 572 1729 573 1737
rect 575 1729 578 1737
rect 580 1729 581 1737
rect 593 1729 594 1737
rect 596 1733 597 1737
rect 596 1729 601 1733
rect 609 1729 610 1737
rect 612 1729 615 1737
rect 617 1729 618 1737
rect 635 1729 636 1737
rect 638 1729 639 1737
rect 651 1729 652 1737
rect 654 1733 655 1737
rect 654 1729 659 1733
rect 667 1729 668 1737
rect 670 1729 673 1737
rect 675 1729 676 1737
rect 688 1729 689 1737
rect 691 1729 692 1737
rect 704 1729 705 1737
rect 707 1729 710 1737
rect 712 1729 713 1737
rect 725 1729 726 1737
rect 728 1733 729 1737
rect 728 1729 733 1733
rect 741 1729 742 1737
rect 744 1729 747 1737
rect 749 1729 750 1737
rect 767 1729 768 1737
rect 770 1729 771 1737
rect 783 1729 784 1737
rect 786 1733 787 1737
rect 786 1729 791 1733
rect 799 1729 800 1737
rect 802 1729 805 1737
rect 807 1729 808 1737
rect 820 1729 821 1737
rect 823 1729 824 1737
rect 836 1729 837 1737
rect 839 1729 842 1737
rect 844 1729 845 1737
rect 857 1729 858 1737
rect 860 1733 861 1737
rect 860 1729 865 1733
rect 873 1729 874 1737
rect 876 1729 879 1737
rect 881 1729 882 1737
rect 899 1729 900 1737
rect 902 1729 903 1737
rect 915 1729 916 1737
rect 918 1733 919 1737
rect 918 1729 923 1733
rect 931 1729 932 1737
rect 934 1729 937 1737
rect 939 1729 940 1737
rect 952 1729 953 1737
rect 955 1729 956 1737
rect 968 1729 969 1737
rect 971 1729 974 1737
rect 976 1729 977 1737
rect 989 1729 990 1737
rect 992 1733 993 1737
rect 992 1729 997 1733
rect 1005 1729 1006 1737
rect 1008 1729 1011 1737
rect 1013 1729 1014 1737
rect 1031 1729 1032 1737
rect 1034 1729 1035 1737
rect 1047 1729 1048 1737
rect 1050 1733 1051 1737
rect 1050 1729 1055 1733
rect 1063 1729 1064 1737
rect 1066 1729 1069 1737
rect 1071 1729 1072 1737
rect 1084 1729 1085 1737
rect 1087 1729 1088 1737
rect 232 1696 233 1704
rect 235 1696 238 1704
rect 240 1696 241 1704
rect 253 1696 254 1704
rect 256 1700 257 1704
rect 256 1696 261 1700
rect 269 1696 270 1704
rect 272 1696 275 1704
rect 277 1696 278 1704
rect 295 1696 296 1704
rect 298 1696 299 1704
rect 311 1696 312 1704
rect 314 1700 315 1704
rect 314 1696 319 1700
rect 327 1696 328 1704
rect 330 1696 333 1704
rect 335 1696 336 1704
rect 348 1696 349 1704
rect 351 1696 352 1704
rect 751 1658 752 1666
rect 754 1658 755 1666
rect 577 1645 578 1653
rect 580 1645 581 1653
rect 593 1645 594 1653
rect 596 1645 597 1653
rect 609 1645 610 1653
rect 612 1645 613 1653
rect 628 1645 633 1653
rect 635 1645 638 1653
rect 640 1645 641 1653
rect 662 1645 664 1653
rect 666 1645 667 1653
rect 684 1645 685 1653
rect 687 1645 688 1653
rect 700 1645 705 1653
rect 707 1645 710 1653
rect 712 1645 713 1653
rect 727 1645 728 1653
rect 730 1645 731 1653
rect 775 1652 778 1660
rect 780 1652 783 1660
rect 785 1652 786 1660
rect 805 1658 806 1666
rect 808 1658 809 1666
rect 832 1658 833 1666
rect 835 1658 836 1666
rect 856 1652 859 1660
rect 861 1652 864 1660
rect 866 1652 867 1660
rect 886 1658 887 1666
rect 889 1658 890 1666
rect 223 1594 224 1602
rect 226 1594 227 1602
rect 239 1594 240 1602
rect 242 1594 245 1602
rect 247 1594 248 1602
rect 260 1598 261 1602
rect 256 1594 261 1598
rect 263 1594 264 1602
rect 276 1594 277 1602
rect 279 1594 280 1602
rect 297 1594 298 1602
rect 300 1594 303 1602
rect 305 1594 306 1602
rect 318 1598 319 1602
rect 314 1594 319 1598
rect 321 1594 322 1602
rect 334 1594 335 1602
rect 337 1594 340 1602
rect 342 1594 343 1602
rect 577 1559 578 1567
rect 580 1559 581 1567
rect 593 1559 594 1567
rect 596 1559 597 1567
rect 609 1559 610 1567
rect 612 1559 613 1567
rect 628 1559 633 1567
rect 635 1559 638 1567
rect 640 1559 641 1567
rect 662 1559 664 1567
rect 666 1559 667 1567
rect 684 1559 685 1567
rect 687 1559 688 1567
rect 700 1559 705 1567
rect 707 1559 710 1567
rect 712 1559 713 1567
rect 727 1559 728 1567
rect 730 1559 731 1567
rect 775 1560 778 1568
rect 780 1560 783 1568
rect 785 1560 786 1568
rect 856 1560 859 1568
rect 861 1560 864 1568
rect 866 1560 867 1568
rect 577 1513 578 1521
rect 580 1513 581 1521
rect 593 1513 594 1521
rect 596 1513 597 1521
rect 609 1513 610 1521
rect 612 1513 613 1521
rect 628 1513 633 1521
rect 635 1513 638 1521
rect 640 1513 641 1521
rect 662 1513 664 1521
rect 666 1513 667 1521
rect 684 1513 685 1521
rect 687 1513 688 1521
rect 700 1513 705 1521
rect 707 1513 710 1521
rect 712 1513 713 1521
rect 727 1513 728 1521
rect 730 1513 731 1521
rect 775 1520 778 1528
rect 780 1520 783 1528
rect 785 1520 786 1528
rect 805 1526 806 1534
rect 808 1526 809 1534
rect 856 1526 857 1534
rect 859 1526 860 1534
rect 880 1520 883 1528
rect 885 1520 888 1528
rect 890 1520 891 1528
rect 910 1526 911 1534
rect 913 1526 914 1534
rect 577 1427 578 1435
rect 580 1427 581 1435
rect 593 1427 594 1435
rect 596 1427 597 1435
rect 609 1427 610 1435
rect 612 1427 613 1435
rect 628 1427 633 1435
rect 635 1427 638 1435
rect 640 1427 641 1435
rect 662 1427 664 1435
rect 666 1427 667 1435
rect 684 1427 685 1435
rect 687 1427 688 1435
rect 700 1427 705 1435
rect 707 1427 710 1435
rect 712 1427 713 1435
rect 727 1427 728 1435
rect 730 1427 731 1435
rect 775 1429 778 1437
rect 780 1429 783 1437
rect 785 1429 786 1437
rect 880 1429 883 1437
rect 885 1429 888 1437
rect 890 1429 891 1437
rect 577 1381 578 1389
rect 580 1381 581 1389
rect 593 1381 594 1389
rect 596 1381 597 1389
rect 609 1381 610 1389
rect 612 1381 613 1389
rect 628 1381 633 1389
rect 635 1381 638 1389
rect 640 1381 641 1389
rect 662 1381 664 1389
rect 666 1381 667 1389
rect 684 1381 685 1389
rect 687 1381 688 1389
rect 700 1381 705 1389
rect 707 1381 710 1389
rect 712 1381 713 1389
rect 727 1381 728 1389
rect 730 1381 731 1389
rect 775 1388 778 1396
rect 780 1388 783 1396
rect 785 1388 786 1396
rect 805 1394 806 1402
rect 808 1394 809 1402
rect 832 1394 833 1402
rect 835 1394 836 1402
rect 856 1388 859 1396
rect 861 1388 864 1396
rect 866 1388 867 1396
rect 886 1394 887 1402
rect 889 1394 890 1402
rect 922 1394 923 1402
rect 925 1394 926 1402
rect 946 1388 949 1396
rect 951 1388 954 1396
rect 956 1388 957 1396
rect 976 1394 977 1402
rect 979 1394 980 1402
rect 577 1295 578 1303
rect 580 1295 581 1303
rect 593 1295 594 1303
rect 596 1295 597 1303
rect 609 1295 610 1303
rect 612 1295 613 1303
rect 628 1295 633 1303
rect 635 1295 638 1303
rect 640 1295 641 1303
rect 662 1295 664 1303
rect 666 1295 667 1303
rect 684 1295 685 1303
rect 687 1295 688 1303
rect 700 1295 705 1303
rect 707 1295 710 1303
rect 712 1295 713 1303
rect 727 1295 728 1303
rect 730 1295 731 1303
rect 775 1294 778 1302
rect 780 1294 783 1302
rect 785 1294 786 1302
rect 856 1294 859 1302
rect 861 1294 864 1302
rect 866 1294 867 1302
rect 946 1294 949 1302
rect 951 1294 954 1302
rect 956 1294 957 1302
rect 577 1249 578 1257
rect 580 1249 581 1257
rect 593 1249 594 1257
rect 596 1249 597 1257
rect 609 1249 610 1257
rect 612 1249 613 1257
rect 628 1249 633 1257
rect 635 1249 638 1257
rect 640 1249 641 1257
rect 662 1249 664 1257
rect 666 1249 667 1257
rect 684 1249 685 1257
rect 687 1249 688 1257
rect 700 1249 705 1257
rect 707 1249 710 1257
rect 712 1249 713 1257
rect 727 1249 728 1257
rect 730 1249 731 1257
rect 775 1256 778 1264
rect 780 1256 783 1264
rect 785 1256 786 1264
rect 805 1262 806 1270
rect 808 1262 809 1270
rect 100 1194 101 1202
rect 103 1194 106 1202
rect 108 1194 109 1202
rect 121 1194 122 1202
rect 124 1198 125 1202
rect 124 1194 129 1198
rect 137 1194 138 1202
rect 140 1194 143 1202
rect 145 1194 146 1202
rect 163 1194 164 1202
rect 166 1194 167 1202
rect 179 1194 180 1202
rect 182 1198 183 1202
rect 182 1194 187 1198
rect 195 1194 196 1202
rect 198 1194 201 1202
rect 203 1194 204 1202
rect 216 1194 217 1202
rect 219 1194 220 1202
rect 232 1194 233 1202
rect 235 1194 238 1202
rect 240 1194 241 1202
rect 253 1194 254 1202
rect 256 1198 257 1202
rect 256 1194 261 1198
rect 269 1194 270 1202
rect 272 1194 275 1202
rect 277 1194 278 1202
rect 295 1194 296 1202
rect 298 1194 299 1202
rect 311 1194 312 1202
rect 314 1198 315 1202
rect 314 1194 319 1198
rect 327 1194 328 1202
rect 330 1194 333 1202
rect 335 1194 336 1202
rect 348 1194 349 1202
rect 351 1194 352 1202
rect 364 1194 365 1202
rect 367 1194 370 1202
rect 372 1194 373 1202
rect 385 1194 386 1202
rect 388 1198 389 1202
rect 388 1194 393 1198
rect 401 1194 402 1202
rect 404 1194 407 1202
rect 409 1194 410 1202
rect 427 1194 428 1202
rect 430 1194 431 1202
rect 443 1194 444 1202
rect 446 1198 447 1202
rect 446 1194 451 1198
rect 459 1194 460 1202
rect 462 1194 465 1202
rect 467 1194 468 1202
rect 480 1194 481 1202
rect 483 1194 484 1202
rect 577 1163 578 1171
rect 580 1163 581 1171
rect 593 1163 594 1171
rect 596 1163 597 1171
rect 609 1163 610 1171
rect 612 1163 613 1171
rect 628 1163 633 1171
rect 635 1163 638 1171
rect 640 1163 641 1171
rect 662 1163 664 1171
rect 666 1163 667 1171
rect 684 1163 685 1171
rect 687 1163 688 1171
rect 700 1163 705 1171
rect 707 1163 710 1171
rect 712 1163 713 1171
rect 727 1163 728 1171
rect 730 1163 731 1171
rect 775 1158 778 1166
rect 780 1158 783 1166
rect 785 1158 786 1166
rect 811 1163 812 1171
rect 814 1163 815 1171
rect 819 1163 825 1171
rect 829 1163 830 1171
rect 832 1163 833 1171
rect 854 1163 855 1171
rect 857 1163 858 1171
rect 870 1163 871 1171
rect 873 1163 874 1171
rect 889 1163 894 1171
rect 896 1163 899 1171
rect 901 1163 902 1171
rect 923 1163 925 1171
rect 927 1163 928 1171
rect 945 1163 946 1171
rect 948 1163 949 1171
rect 961 1163 966 1171
rect 968 1163 971 1171
rect 973 1163 974 1171
rect 988 1163 989 1171
rect 991 1163 992 1171
rect 871 1084 872 1092
rect 874 1084 877 1092
rect 879 1084 880 1092
rect 892 1084 893 1092
rect 895 1088 896 1092
rect 895 1084 900 1088
rect 908 1084 909 1092
rect 911 1084 914 1092
rect 916 1084 917 1092
rect 934 1084 935 1092
rect 937 1084 938 1092
rect 950 1084 951 1092
rect 953 1088 954 1092
rect 953 1084 958 1088
rect 966 1084 967 1092
rect 969 1084 972 1092
rect 974 1084 975 1092
rect 987 1084 988 1092
rect 990 1084 991 1092
rect 100 1054 101 1062
rect 103 1054 106 1062
rect 108 1054 109 1062
rect 121 1054 122 1062
rect 124 1058 125 1062
rect 124 1054 129 1058
rect 137 1054 138 1062
rect 140 1054 143 1062
rect 145 1054 146 1062
rect 163 1054 164 1062
rect 166 1054 167 1062
rect 179 1054 180 1062
rect 182 1058 183 1062
rect 182 1054 187 1058
rect 195 1054 196 1062
rect 198 1054 201 1062
rect 203 1054 204 1062
rect 216 1054 217 1062
rect 219 1054 220 1062
rect 232 1054 233 1062
rect 235 1054 238 1062
rect 240 1054 241 1062
rect 253 1054 254 1062
rect 256 1058 257 1062
rect 256 1054 261 1058
rect 269 1054 270 1062
rect 272 1054 275 1062
rect 277 1054 278 1062
rect 295 1054 296 1062
rect 298 1054 299 1062
rect 311 1054 312 1062
rect 314 1058 315 1062
rect 314 1054 319 1058
rect 327 1054 328 1062
rect 330 1054 333 1062
rect 335 1054 336 1062
rect 348 1054 349 1062
rect 351 1054 352 1062
rect 364 1054 365 1062
rect 367 1054 370 1062
rect 372 1054 373 1062
rect 385 1054 386 1062
rect 388 1058 389 1062
rect 388 1054 393 1058
rect 401 1054 402 1062
rect 404 1054 407 1062
rect 409 1054 410 1062
rect 427 1054 428 1062
rect 430 1054 431 1062
rect 443 1054 444 1062
rect 446 1058 447 1062
rect 446 1054 451 1058
rect 459 1054 460 1062
rect 462 1054 465 1062
rect 467 1054 468 1062
rect 480 1054 481 1062
rect 483 1054 484 1062
rect 871 998 872 1006
rect 874 998 877 1006
rect 879 998 880 1006
rect 892 998 893 1006
rect 895 1002 896 1006
rect 895 998 900 1002
rect 908 998 909 1006
rect 911 998 914 1006
rect 916 998 917 1006
rect 934 998 935 1006
rect 937 998 938 1006
rect 950 998 951 1006
rect 953 1002 954 1006
rect 953 998 958 1002
rect 966 998 967 1006
rect 969 998 972 1006
rect 974 998 975 1006
rect 987 998 988 1006
rect 990 998 991 1006
rect 100 968 101 976
rect 103 968 106 976
rect 108 968 109 976
rect 121 968 122 976
rect 124 972 125 976
rect 124 968 129 972
rect 137 968 138 976
rect 140 968 143 976
rect 145 968 146 976
rect 163 968 164 976
rect 166 968 167 976
rect 179 968 180 976
rect 182 972 183 976
rect 182 968 187 972
rect 195 968 196 976
rect 198 968 201 976
rect 203 968 204 976
rect 216 968 217 976
rect 219 968 220 976
rect 232 968 233 976
rect 235 968 238 976
rect 240 968 241 976
rect 253 968 254 976
rect 256 972 257 976
rect 256 968 261 972
rect 269 968 270 976
rect 272 968 275 976
rect 277 968 278 976
rect 295 968 296 976
rect 298 968 299 976
rect 311 968 312 976
rect 314 972 315 976
rect 314 968 319 972
rect 327 968 328 976
rect 330 968 333 976
rect 335 968 336 976
rect 348 968 349 976
rect 351 968 352 976
rect 364 968 365 976
rect 367 968 370 976
rect 372 968 373 976
rect 385 968 386 976
rect 388 972 389 976
rect 388 968 393 972
rect 401 968 402 976
rect 404 968 407 976
rect 409 968 410 976
rect 427 968 428 976
rect 430 968 431 976
rect 443 968 444 976
rect 446 972 447 976
rect 446 968 451 972
rect 459 968 460 976
rect 462 968 465 976
rect 467 968 468 976
rect 480 968 481 976
rect 483 968 484 976
rect 100 828 101 836
rect 103 828 106 836
rect 108 828 109 836
rect 121 828 122 836
rect 124 832 125 836
rect 124 828 129 832
rect 137 828 138 836
rect 140 828 143 836
rect 145 828 146 836
rect 163 828 164 836
rect 166 828 167 836
rect 179 828 180 836
rect 182 832 183 836
rect 182 828 187 832
rect 195 828 196 836
rect 198 828 201 836
rect 203 828 204 836
rect 216 828 217 836
rect 219 828 220 836
rect 232 828 233 836
rect 235 828 238 836
rect 240 828 241 836
rect 253 828 254 836
rect 256 832 257 836
rect 256 828 261 832
rect 269 828 270 836
rect 272 828 275 836
rect 277 828 278 836
rect 295 828 296 836
rect 298 828 299 836
rect 311 828 312 836
rect 314 832 315 836
rect 314 828 319 832
rect 327 828 328 836
rect 330 828 333 836
rect 335 828 336 836
rect 348 828 349 836
rect 351 828 352 836
rect 364 828 365 836
rect 367 828 370 836
rect 372 828 373 836
rect 385 828 386 836
rect 388 832 389 836
rect 388 828 393 832
rect 401 828 402 836
rect 404 828 407 836
rect 409 828 410 836
rect 427 828 428 836
rect 430 828 431 836
rect 443 828 444 836
rect 446 832 447 836
rect 446 828 451 832
rect 459 828 460 836
rect 462 828 465 836
rect 467 828 468 836
rect 480 828 481 836
rect 483 828 484 836
<< ndcontact >>
rect 568 1706 572 1710
rect 581 1706 585 1710
rect 589 1706 593 1710
rect 597 1706 601 1710
rect 605 1706 609 1710
rect 618 1706 622 1710
rect 631 1706 635 1710
rect 639 1706 643 1710
rect 647 1706 651 1710
rect 655 1706 659 1710
rect 663 1706 667 1710
rect 676 1706 680 1710
rect 684 1706 688 1710
rect 692 1706 696 1710
rect 700 1706 704 1710
rect 713 1706 717 1710
rect 721 1706 725 1710
rect 729 1706 733 1710
rect 737 1706 741 1710
rect 750 1706 754 1710
rect 763 1706 767 1710
rect 771 1706 775 1710
rect 779 1706 783 1710
rect 787 1706 791 1710
rect 795 1706 799 1710
rect 808 1706 812 1710
rect 816 1706 820 1710
rect 824 1706 828 1710
rect 832 1706 836 1710
rect 845 1706 849 1710
rect 853 1706 857 1710
rect 861 1706 865 1710
rect 869 1706 873 1710
rect 882 1706 886 1710
rect 895 1706 899 1710
rect 903 1706 907 1710
rect 911 1706 915 1710
rect 919 1706 923 1710
rect 927 1706 931 1710
rect 940 1706 944 1710
rect 948 1706 952 1710
rect 956 1706 960 1710
rect 964 1706 968 1710
rect 977 1706 981 1710
rect 985 1706 989 1710
rect 993 1706 997 1710
rect 1001 1706 1005 1710
rect 1014 1706 1018 1710
rect 1027 1706 1031 1710
rect 1035 1706 1039 1710
rect 1043 1706 1047 1710
rect 1051 1706 1055 1710
rect 1059 1706 1063 1710
rect 1072 1706 1076 1710
rect 1080 1706 1084 1710
rect 1088 1706 1092 1710
rect 228 1673 232 1677
rect 241 1673 245 1677
rect 249 1673 253 1677
rect 257 1673 261 1677
rect 265 1673 269 1677
rect 278 1673 282 1677
rect 291 1673 295 1677
rect 299 1673 303 1677
rect 307 1673 311 1677
rect 315 1673 319 1677
rect 323 1673 327 1677
rect 336 1673 340 1677
rect 344 1673 348 1677
rect 352 1673 356 1677
rect 352 1636 356 1640
rect 360 1636 364 1640
rect 747 1640 751 1644
rect 755 1640 759 1644
rect 771 1636 775 1640
rect 786 1636 790 1640
rect 828 1640 832 1644
rect 836 1640 840 1644
rect 852 1636 856 1640
rect 867 1636 871 1640
rect 801 1632 805 1636
rect 809 1632 813 1636
rect 235 1627 239 1631
rect 243 1627 247 1631
rect 573 1627 577 1631
rect 581 1627 585 1631
rect 589 1627 593 1631
rect 597 1627 601 1631
rect 605 1627 609 1631
rect 613 1627 617 1631
rect 624 1627 628 1631
rect 641 1627 645 1631
rect 658 1627 662 1631
rect 667 1627 671 1631
rect 680 1627 684 1631
rect 688 1627 692 1631
rect 696 1627 700 1631
rect 713 1627 717 1631
rect 723 1627 727 1631
rect 731 1627 735 1631
rect 882 1632 886 1636
rect 890 1632 894 1636
rect 573 1581 577 1585
rect 581 1581 585 1585
rect 589 1581 593 1585
rect 597 1581 601 1585
rect 605 1581 609 1585
rect 613 1581 617 1585
rect 624 1581 628 1585
rect 641 1581 645 1585
rect 658 1581 662 1585
rect 667 1581 671 1585
rect 680 1581 684 1585
rect 688 1581 692 1585
rect 696 1581 700 1585
rect 713 1581 717 1585
rect 723 1581 727 1585
rect 731 1581 735 1585
rect 219 1571 223 1575
rect 227 1571 231 1575
rect 235 1571 239 1575
rect 248 1571 252 1575
rect 256 1571 260 1575
rect 264 1571 268 1575
rect 272 1571 276 1575
rect 280 1571 284 1575
rect 293 1571 297 1575
rect 306 1571 310 1575
rect 314 1571 318 1575
rect 322 1571 326 1575
rect 330 1571 334 1575
rect 343 1571 347 1575
rect 771 1580 775 1584
rect 786 1580 790 1584
rect 852 1580 856 1584
rect 867 1580 871 1584
rect 771 1504 775 1508
rect 786 1504 790 1508
rect 852 1508 856 1512
rect 860 1508 864 1512
rect 876 1504 880 1508
rect 891 1504 895 1508
rect 801 1500 805 1504
rect 809 1500 813 1504
rect 573 1495 577 1499
rect 581 1495 585 1499
rect 589 1495 593 1499
rect 597 1495 601 1499
rect 605 1495 609 1499
rect 613 1495 617 1499
rect 624 1495 628 1499
rect 641 1495 645 1499
rect 658 1495 662 1499
rect 667 1495 671 1499
rect 680 1495 684 1499
rect 688 1495 692 1499
rect 696 1495 700 1499
rect 713 1495 717 1499
rect 723 1495 727 1499
rect 731 1495 735 1499
rect 906 1500 910 1504
rect 914 1500 918 1504
rect 573 1449 577 1453
rect 581 1449 585 1453
rect 589 1449 593 1453
rect 597 1449 601 1453
rect 605 1449 609 1453
rect 613 1449 617 1453
rect 624 1449 628 1453
rect 641 1449 645 1453
rect 658 1449 662 1453
rect 667 1449 671 1453
rect 680 1449 684 1453
rect 688 1449 692 1453
rect 696 1449 700 1453
rect 713 1449 717 1453
rect 723 1449 727 1453
rect 731 1449 735 1453
rect 771 1449 775 1453
rect 786 1449 790 1453
rect 876 1449 880 1453
rect 891 1449 895 1453
rect 771 1372 775 1376
rect 786 1372 790 1376
rect 828 1376 832 1380
rect 836 1376 840 1380
rect 852 1372 856 1376
rect 867 1372 871 1376
rect 918 1376 922 1380
rect 926 1376 930 1380
rect 942 1372 946 1376
rect 957 1372 961 1376
rect 801 1368 805 1372
rect 809 1368 813 1372
rect 573 1363 577 1367
rect 581 1363 585 1367
rect 589 1363 593 1367
rect 597 1363 601 1367
rect 605 1363 609 1367
rect 613 1363 617 1367
rect 624 1363 628 1367
rect 641 1363 645 1367
rect 658 1363 662 1367
rect 667 1363 671 1367
rect 680 1363 684 1367
rect 688 1363 692 1367
rect 696 1363 700 1367
rect 713 1363 717 1367
rect 723 1363 727 1367
rect 731 1363 735 1367
rect 882 1368 886 1372
rect 890 1368 894 1372
rect 972 1368 976 1372
rect 980 1368 984 1372
rect 573 1317 577 1321
rect 581 1317 585 1321
rect 589 1317 593 1321
rect 597 1317 601 1321
rect 605 1317 609 1321
rect 613 1317 617 1321
rect 624 1317 628 1321
rect 641 1317 645 1321
rect 658 1317 662 1321
rect 667 1317 671 1321
rect 680 1317 684 1321
rect 688 1317 692 1321
rect 696 1317 700 1321
rect 713 1317 717 1321
rect 723 1317 727 1321
rect 731 1317 735 1321
rect 771 1314 775 1318
rect 786 1314 790 1318
rect 852 1314 856 1318
rect 867 1314 871 1318
rect 942 1314 946 1318
rect 957 1314 961 1318
rect 771 1240 775 1244
rect 786 1240 790 1244
rect 801 1236 805 1240
rect 809 1236 813 1240
rect 573 1231 577 1235
rect 581 1231 585 1235
rect 589 1231 593 1235
rect 597 1231 601 1235
rect 605 1231 609 1235
rect 613 1231 617 1235
rect 624 1231 628 1235
rect 641 1231 645 1235
rect 658 1231 662 1235
rect 667 1231 671 1235
rect 680 1231 684 1235
rect 688 1231 692 1235
rect 696 1231 700 1235
rect 713 1231 717 1235
rect 723 1231 727 1235
rect 731 1231 735 1235
rect 573 1185 577 1189
rect 581 1185 585 1189
rect 589 1185 593 1189
rect 597 1185 601 1189
rect 605 1185 609 1189
rect 613 1185 617 1189
rect 624 1185 628 1189
rect 641 1185 645 1189
rect 658 1185 662 1189
rect 667 1185 671 1189
rect 680 1185 684 1189
rect 688 1185 692 1189
rect 696 1185 700 1189
rect 713 1185 717 1189
rect 723 1185 727 1189
rect 731 1185 735 1189
rect 807 1185 811 1189
rect 815 1185 819 1189
rect 825 1185 829 1189
rect 833 1185 837 1189
rect 842 1185 846 1189
rect 850 1185 854 1189
rect 858 1185 862 1189
rect 866 1185 870 1189
rect 874 1185 878 1189
rect 885 1185 889 1189
rect 902 1185 906 1189
rect 919 1185 923 1189
rect 928 1185 932 1189
rect 941 1185 945 1189
rect 949 1185 953 1189
rect 957 1185 961 1189
rect 974 1185 978 1189
rect 984 1185 988 1189
rect 992 1185 996 1189
rect 96 1171 100 1175
rect 109 1171 113 1175
rect 117 1171 121 1175
rect 125 1171 129 1175
rect 133 1171 137 1175
rect 146 1171 150 1175
rect 159 1171 163 1175
rect 167 1171 171 1175
rect 175 1171 179 1175
rect 183 1171 187 1175
rect 191 1171 195 1175
rect 204 1171 208 1175
rect 212 1171 216 1175
rect 220 1171 224 1175
rect 228 1171 232 1175
rect 241 1171 245 1175
rect 249 1171 253 1175
rect 257 1171 261 1175
rect 265 1171 269 1175
rect 278 1171 282 1175
rect 291 1171 295 1175
rect 299 1171 303 1175
rect 307 1171 311 1175
rect 315 1171 319 1175
rect 323 1171 327 1175
rect 336 1171 340 1175
rect 344 1171 348 1175
rect 352 1171 356 1175
rect 360 1171 364 1175
rect 373 1171 377 1175
rect 381 1171 385 1175
rect 389 1171 393 1175
rect 397 1171 401 1175
rect 410 1171 414 1175
rect 423 1171 427 1175
rect 431 1171 435 1175
rect 439 1171 443 1175
rect 447 1171 451 1175
rect 455 1171 459 1175
rect 468 1171 472 1175
rect 476 1171 480 1175
rect 484 1171 488 1175
rect 771 1178 775 1182
rect 786 1178 790 1182
rect 1001 1132 1005 1136
rect 211 1127 215 1131
rect 219 1127 223 1131
rect 235 1127 239 1131
rect 243 1127 247 1131
rect 1001 1124 1005 1128
rect 231 1116 235 1120
rect 239 1116 243 1120
rect 227 1105 231 1109
rect 227 1097 231 1101
rect 211 1093 215 1097
rect 219 1093 223 1097
rect 235 1093 239 1097
rect 243 1093 247 1097
rect 867 1061 871 1065
rect 880 1061 884 1065
rect 888 1061 892 1065
rect 896 1061 900 1065
rect 904 1061 908 1065
rect 917 1061 921 1065
rect 930 1061 934 1065
rect 938 1061 942 1065
rect 946 1061 950 1065
rect 954 1061 958 1065
rect 962 1061 966 1065
rect 975 1061 979 1065
rect 983 1061 987 1065
rect 991 1061 995 1065
rect 96 1031 100 1035
rect 109 1031 113 1035
rect 117 1031 121 1035
rect 125 1031 129 1035
rect 133 1031 137 1035
rect 146 1031 150 1035
rect 159 1031 163 1035
rect 167 1031 171 1035
rect 175 1031 179 1035
rect 183 1031 187 1035
rect 191 1031 195 1035
rect 204 1031 208 1035
rect 212 1031 216 1035
rect 220 1031 224 1035
rect 228 1031 232 1035
rect 241 1031 245 1035
rect 249 1031 253 1035
rect 257 1031 261 1035
rect 265 1031 269 1035
rect 278 1031 282 1035
rect 291 1031 295 1035
rect 299 1031 303 1035
rect 307 1031 311 1035
rect 315 1031 319 1035
rect 323 1031 327 1035
rect 336 1031 340 1035
rect 344 1031 348 1035
rect 352 1031 356 1035
rect 360 1031 364 1035
rect 373 1031 377 1035
rect 381 1031 385 1035
rect 389 1031 393 1035
rect 397 1031 401 1035
rect 410 1031 414 1035
rect 423 1031 427 1035
rect 431 1031 435 1035
rect 439 1031 443 1035
rect 447 1031 451 1035
rect 455 1031 459 1035
rect 468 1031 472 1035
rect 476 1031 480 1035
rect 484 1031 488 1035
rect 1013 988 1017 992
rect 1013 980 1017 984
rect 867 975 871 979
rect 880 975 884 979
rect 888 975 892 979
rect 896 975 900 979
rect 904 975 908 979
rect 917 975 921 979
rect 930 975 934 979
rect 938 975 942 979
rect 946 975 950 979
rect 954 975 958 979
rect 962 975 966 979
rect 975 975 979 979
rect 983 975 987 979
rect 991 975 995 979
rect 96 945 100 949
rect 109 945 113 949
rect 117 945 121 949
rect 125 945 129 949
rect 133 945 137 949
rect 146 945 150 949
rect 159 945 163 949
rect 167 945 171 949
rect 175 945 179 949
rect 183 945 187 949
rect 191 945 195 949
rect 204 945 208 949
rect 212 945 216 949
rect 220 945 224 949
rect 228 945 232 949
rect 241 945 245 949
rect 249 945 253 949
rect 257 945 261 949
rect 265 945 269 949
rect 278 945 282 949
rect 291 945 295 949
rect 299 945 303 949
rect 307 945 311 949
rect 315 945 319 949
rect 323 945 327 949
rect 336 945 340 949
rect 344 945 348 949
rect 352 945 356 949
rect 360 945 364 949
rect 373 945 377 949
rect 381 945 385 949
rect 389 945 393 949
rect 397 945 401 949
rect 410 945 414 949
rect 423 945 427 949
rect 431 945 435 949
rect 439 945 443 949
rect 447 945 451 949
rect 455 945 459 949
rect 468 945 472 949
rect 476 945 480 949
rect 484 945 488 949
rect 328 901 332 905
rect 336 901 340 905
rect 352 901 356 905
rect 360 901 364 905
rect 348 890 352 894
rect 356 890 360 894
rect 344 879 348 883
rect 344 871 348 875
rect 328 867 332 871
rect 336 867 340 871
rect 352 867 356 871
rect 360 867 364 871
rect 96 805 100 809
rect 109 805 113 809
rect 117 805 121 809
rect 125 805 129 809
rect 133 805 137 809
rect 146 805 150 809
rect 159 805 163 809
rect 167 805 171 809
rect 175 805 179 809
rect 183 805 187 809
rect 191 805 195 809
rect 204 805 208 809
rect 212 805 216 809
rect 220 805 224 809
rect 228 805 232 809
rect 241 805 245 809
rect 249 805 253 809
rect 257 805 261 809
rect 265 805 269 809
rect 278 805 282 809
rect 291 805 295 809
rect 299 805 303 809
rect 307 805 311 809
rect 315 805 319 809
rect 323 805 327 809
rect 336 805 340 809
rect 344 805 348 809
rect 352 805 356 809
rect 360 805 364 809
rect 373 805 377 809
rect 381 805 385 809
rect 389 805 393 809
rect 397 805 401 809
rect 410 805 414 809
rect 423 805 427 809
rect 431 805 435 809
rect 439 805 443 809
rect 447 805 451 809
rect 455 805 459 809
rect 468 805 472 809
rect 476 805 480 809
rect 484 805 488 809
<< pdcontact >>
rect 568 1729 572 1737
rect 581 1729 585 1737
rect 589 1729 593 1737
rect 597 1733 601 1737
rect 605 1729 609 1737
rect 618 1729 622 1737
rect 631 1729 635 1737
rect 639 1729 643 1737
rect 647 1729 651 1737
rect 655 1733 659 1737
rect 663 1729 667 1737
rect 676 1729 680 1737
rect 684 1729 688 1737
rect 692 1729 696 1737
rect 700 1729 704 1737
rect 713 1729 717 1737
rect 721 1729 725 1737
rect 729 1733 733 1737
rect 737 1729 741 1737
rect 750 1729 754 1737
rect 763 1729 767 1737
rect 771 1729 775 1737
rect 779 1729 783 1737
rect 787 1733 791 1737
rect 795 1729 799 1737
rect 808 1729 812 1737
rect 816 1729 820 1737
rect 824 1729 828 1737
rect 832 1729 836 1737
rect 845 1729 849 1737
rect 853 1729 857 1737
rect 861 1733 865 1737
rect 869 1729 873 1737
rect 882 1729 886 1737
rect 895 1729 899 1737
rect 903 1729 907 1737
rect 911 1729 915 1737
rect 919 1733 923 1737
rect 927 1729 931 1737
rect 940 1729 944 1737
rect 948 1729 952 1737
rect 956 1729 960 1737
rect 964 1729 968 1737
rect 977 1729 981 1737
rect 985 1729 989 1737
rect 993 1733 997 1737
rect 1001 1729 1005 1737
rect 1014 1729 1018 1737
rect 1027 1729 1031 1737
rect 1035 1729 1039 1737
rect 1043 1729 1047 1737
rect 1051 1733 1055 1737
rect 1059 1729 1063 1737
rect 1072 1729 1076 1737
rect 1080 1729 1084 1737
rect 1088 1729 1092 1737
rect 228 1696 232 1704
rect 241 1696 245 1704
rect 249 1696 253 1704
rect 257 1700 261 1704
rect 265 1696 269 1704
rect 278 1696 282 1704
rect 291 1696 295 1704
rect 299 1696 303 1704
rect 307 1696 311 1704
rect 315 1700 319 1704
rect 323 1696 327 1704
rect 336 1696 340 1704
rect 344 1696 348 1704
rect 352 1696 356 1704
rect 747 1658 751 1666
rect 755 1658 759 1666
rect 573 1645 577 1653
rect 581 1645 585 1653
rect 589 1645 593 1653
rect 597 1645 601 1653
rect 605 1645 609 1653
rect 613 1645 617 1653
rect 624 1645 628 1653
rect 641 1645 645 1653
rect 658 1645 662 1653
rect 667 1645 671 1653
rect 680 1645 684 1653
rect 688 1645 692 1653
rect 696 1645 700 1653
rect 713 1645 717 1653
rect 723 1645 727 1653
rect 731 1645 735 1653
rect 771 1652 775 1660
rect 786 1652 790 1660
rect 801 1658 805 1666
rect 809 1658 813 1666
rect 828 1658 832 1666
rect 836 1658 840 1666
rect 852 1652 856 1660
rect 867 1652 871 1660
rect 882 1658 886 1666
rect 890 1658 894 1666
rect 219 1594 223 1602
rect 227 1594 231 1602
rect 235 1594 239 1602
rect 248 1594 252 1602
rect 256 1598 260 1602
rect 264 1594 268 1602
rect 272 1594 276 1602
rect 280 1594 284 1602
rect 293 1594 297 1602
rect 306 1594 310 1602
rect 314 1598 318 1602
rect 322 1594 326 1602
rect 330 1594 334 1602
rect 343 1594 347 1602
rect 573 1559 577 1567
rect 581 1559 585 1567
rect 589 1559 593 1567
rect 597 1559 601 1567
rect 605 1559 609 1567
rect 613 1559 617 1567
rect 624 1559 628 1567
rect 641 1559 645 1567
rect 658 1559 662 1567
rect 667 1559 671 1567
rect 680 1559 684 1567
rect 688 1559 692 1567
rect 696 1559 700 1567
rect 713 1559 717 1567
rect 723 1559 727 1567
rect 731 1559 735 1567
rect 771 1560 775 1568
rect 786 1560 790 1568
rect 852 1560 856 1568
rect 867 1560 871 1568
rect 573 1513 577 1521
rect 581 1513 585 1521
rect 589 1513 593 1521
rect 597 1513 601 1521
rect 605 1513 609 1521
rect 613 1513 617 1521
rect 624 1513 628 1521
rect 641 1513 645 1521
rect 658 1513 662 1521
rect 667 1513 671 1521
rect 680 1513 684 1521
rect 688 1513 692 1521
rect 696 1513 700 1521
rect 713 1513 717 1521
rect 723 1513 727 1521
rect 731 1513 735 1521
rect 771 1520 775 1528
rect 786 1520 790 1528
rect 801 1526 805 1534
rect 809 1526 813 1534
rect 852 1526 856 1534
rect 860 1526 864 1534
rect 876 1520 880 1528
rect 891 1520 895 1528
rect 906 1526 910 1534
rect 914 1526 918 1534
rect 573 1427 577 1435
rect 581 1427 585 1435
rect 589 1427 593 1435
rect 597 1427 601 1435
rect 605 1427 609 1435
rect 613 1427 617 1435
rect 624 1427 628 1435
rect 641 1427 645 1435
rect 658 1427 662 1435
rect 667 1427 671 1435
rect 680 1427 684 1435
rect 688 1427 692 1435
rect 696 1427 700 1435
rect 713 1427 717 1435
rect 723 1427 727 1435
rect 731 1427 735 1435
rect 771 1429 775 1437
rect 786 1429 790 1437
rect 876 1429 880 1437
rect 891 1429 895 1437
rect 573 1381 577 1389
rect 581 1381 585 1389
rect 589 1381 593 1389
rect 597 1381 601 1389
rect 605 1381 609 1389
rect 613 1381 617 1389
rect 624 1381 628 1389
rect 641 1381 645 1389
rect 658 1381 662 1389
rect 667 1381 671 1389
rect 680 1381 684 1389
rect 688 1381 692 1389
rect 696 1381 700 1389
rect 713 1381 717 1389
rect 723 1381 727 1389
rect 731 1381 735 1389
rect 771 1388 775 1396
rect 786 1388 790 1396
rect 801 1394 805 1402
rect 809 1394 813 1402
rect 828 1394 832 1402
rect 836 1394 840 1402
rect 852 1388 856 1396
rect 867 1388 871 1396
rect 882 1394 886 1402
rect 890 1394 894 1402
rect 918 1394 922 1402
rect 926 1394 930 1402
rect 942 1388 946 1396
rect 957 1388 961 1396
rect 972 1394 976 1402
rect 980 1394 984 1402
rect 573 1295 577 1303
rect 581 1295 585 1303
rect 589 1295 593 1303
rect 597 1295 601 1303
rect 605 1295 609 1303
rect 613 1295 617 1303
rect 624 1295 628 1303
rect 641 1295 645 1303
rect 658 1295 662 1303
rect 667 1295 671 1303
rect 680 1295 684 1303
rect 688 1295 692 1303
rect 696 1295 700 1303
rect 713 1295 717 1303
rect 723 1295 727 1303
rect 731 1295 735 1303
rect 771 1294 775 1302
rect 786 1294 790 1302
rect 852 1294 856 1302
rect 867 1294 871 1302
rect 942 1294 946 1302
rect 957 1294 961 1302
rect 573 1249 577 1257
rect 581 1249 585 1257
rect 589 1249 593 1257
rect 597 1249 601 1257
rect 605 1249 609 1257
rect 613 1249 617 1257
rect 624 1249 628 1257
rect 641 1249 645 1257
rect 658 1249 662 1257
rect 667 1249 671 1257
rect 680 1249 684 1257
rect 688 1249 692 1257
rect 696 1249 700 1257
rect 713 1249 717 1257
rect 723 1249 727 1257
rect 731 1249 735 1257
rect 771 1256 775 1264
rect 786 1256 790 1264
rect 801 1262 805 1270
rect 809 1262 813 1270
rect 96 1194 100 1202
rect 109 1194 113 1202
rect 117 1194 121 1202
rect 125 1198 129 1202
rect 133 1194 137 1202
rect 146 1194 150 1202
rect 159 1194 163 1202
rect 167 1194 171 1202
rect 175 1194 179 1202
rect 183 1198 187 1202
rect 191 1194 195 1202
rect 204 1194 208 1202
rect 212 1194 216 1202
rect 220 1194 224 1202
rect 228 1194 232 1202
rect 241 1194 245 1202
rect 249 1194 253 1202
rect 257 1198 261 1202
rect 265 1194 269 1202
rect 278 1194 282 1202
rect 291 1194 295 1202
rect 299 1194 303 1202
rect 307 1194 311 1202
rect 315 1198 319 1202
rect 323 1194 327 1202
rect 336 1194 340 1202
rect 344 1194 348 1202
rect 352 1194 356 1202
rect 360 1194 364 1202
rect 373 1194 377 1202
rect 381 1194 385 1202
rect 389 1198 393 1202
rect 397 1194 401 1202
rect 410 1194 414 1202
rect 423 1194 427 1202
rect 431 1194 435 1202
rect 439 1194 443 1202
rect 447 1198 451 1202
rect 455 1194 459 1202
rect 468 1194 472 1202
rect 476 1194 480 1202
rect 484 1194 488 1202
rect 573 1163 577 1171
rect 581 1163 585 1171
rect 589 1163 593 1171
rect 597 1163 601 1171
rect 605 1163 609 1171
rect 613 1163 617 1171
rect 624 1163 628 1171
rect 641 1163 645 1171
rect 658 1163 662 1171
rect 667 1163 671 1171
rect 680 1163 684 1171
rect 688 1163 692 1171
rect 696 1163 700 1171
rect 713 1163 717 1171
rect 723 1163 727 1171
rect 731 1163 735 1171
rect 771 1158 775 1166
rect 786 1158 790 1166
rect 807 1163 811 1171
rect 815 1163 819 1171
rect 825 1163 829 1171
rect 833 1163 837 1171
rect 842 1163 846 1171
rect 850 1163 854 1171
rect 858 1163 862 1171
rect 866 1163 870 1171
rect 874 1163 878 1171
rect 885 1163 889 1171
rect 902 1163 906 1171
rect 919 1163 923 1171
rect 928 1163 932 1171
rect 941 1163 945 1171
rect 949 1163 953 1171
rect 957 1163 961 1171
rect 974 1163 978 1171
rect 984 1163 988 1171
rect 992 1163 996 1171
rect 867 1084 871 1092
rect 880 1084 884 1092
rect 888 1084 892 1092
rect 896 1088 900 1092
rect 904 1084 908 1092
rect 917 1084 921 1092
rect 930 1084 934 1092
rect 938 1084 942 1092
rect 946 1084 950 1092
rect 954 1088 958 1092
rect 962 1084 966 1092
rect 975 1084 979 1092
rect 983 1084 987 1092
rect 991 1084 995 1092
rect 96 1054 100 1062
rect 109 1054 113 1062
rect 117 1054 121 1062
rect 125 1058 129 1062
rect 133 1054 137 1062
rect 146 1054 150 1062
rect 159 1054 163 1062
rect 167 1054 171 1062
rect 175 1054 179 1062
rect 183 1058 187 1062
rect 191 1054 195 1062
rect 204 1054 208 1062
rect 212 1054 216 1062
rect 220 1054 224 1062
rect 228 1054 232 1062
rect 241 1054 245 1062
rect 249 1054 253 1062
rect 257 1058 261 1062
rect 265 1054 269 1062
rect 278 1054 282 1062
rect 291 1054 295 1062
rect 299 1054 303 1062
rect 307 1054 311 1062
rect 315 1058 319 1062
rect 323 1054 327 1062
rect 336 1054 340 1062
rect 344 1054 348 1062
rect 352 1054 356 1062
rect 360 1054 364 1062
rect 373 1054 377 1062
rect 381 1054 385 1062
rect 389 1058 393 1062
rect 397 1054 401 1062
rect 410 1054 414 1062
rect 423 1054 427 1062
rect 431 1054 435 1062
rect 439 1054 443 1062
rect 447 1058 451 1062
rect 455 1054 459 1062
rect 468 1054 472 1062
rect 476 1054 480 1062
rect 484 1054 488 1062
rect 867 998 871 1006
rect 880 998 884 1006
rect 888 998 892 1006
rect 896 1002 900 1006
rect 904 998 908 1006
rect 917 998 921 1006
rect 930 998 934 1006
rect 938 998 942 1006
rect 946 998 950 1006
rect 954 1002 958 1006
rect 962 998 966 1006
rect 975 998 979 1006
rect 983 998 987 1006
rect 991 998 995 1006
rect 96 968 100 976
rect 109 968 113 976
rect 117 968 121 976
rect 125 972 129 976
rect 133 968 137 976
rect 146 968 150 976
rect 159 968 163 976
rect 167 968 171 976
rect 175 968 179 976
rect 183 972 187 976
rect 191 968 195 976
rect 204 968 208 976
rect 212 968 216 976
rect 220 968 224 976
rect 228 968 232 976
rect 241 968 245 976
rect 249 968 253 976
rect 257 972 261 976
rect 265 968 269 976
rect 278 968 282 976
rect 291 968 295 976
rect 299 968 303 976
rect 307 968 311 976
rect 315 972 319 976
rect 323 968 327 976
rect 336 968 340 976
rect 344 968 348 976
rect 352 968 356 976
rect 360 968 364 976
rect 373 968 377 976
rect 381 968 385 976
rect 389 972 393 976
rect 397 968 401 976
rect 410 968 414 976
rect 423 968 427 976
rect 431 968 435 976
rect 439 968 443 976
rect 447 972 451 976
rect 455 968 459 976
rect 468 968 472 976
rect 476 968 480 976
rect 484 968 488 976
rect 96 828 100 836
rect 109 828 113 836
rect 117 828 121 836
rect 125 832 129 836
rect 133 828 137 836
rect 146 828 150 836
rect 159 828 163 836
rect 167 828 171 836
rect 175 828 179 836
rect 183 832 187 836
rect 191 828 195 836
rect 204 828 208 836
rect 212 828 216 836
rect 220 828 224 836
rect 228 828 232 836
rect 241 828 245 836
rect 249 828 253 836
rect 257 832 261 836
rect 265 828 269 836
rect 278 828 282 836
rect 291 828 295 836
rect 299 828 303 836
rect 307 828 311 836
rect 315 832 319 836
rect 323 828 327 836
rect 336 828 340 836
rect 344 828 348 836
rect 352 828 356 836
rect 360 828 364 836
rect 373 828 377 836
rect 381 828 385 836
rect 389 832 393 836
rect 397 828 401 836
rect 410 828 414 836
rect 423 828 427 836
rect 431 828 435 836
rect 439 828 443 836
rect 447 832 451 836
rect 455 828 459 836
rect 468 828 472 836
rect 476 828 480 836
rect 484 828 488 836
<< psubstratepcontact >>
rect 598 1690 602 1694
rect 626 1690 630 1694
rect 656 1690 660 1694
rect 730 1690 734 1694
rect 758 1690 762 1694
rect 788 1690 792 1694
rect 862 1690 866 1694
rect 890 1690 894 1694
rect 920 1690 924 1694
rect 994 1690 998 1694
rect 1022 1690 1026 1694
rect 1052 1690 1056 1694
rect 258 1657 262 1661
rect 286 1657 290 1661
rect 316 1657 320 1661
rect 579 1604 583 1608
rect 614 1604 618 1608
rect 740 1604 744 1608
rect 764 1604 768 1608
rect 818 1604 825 1608
rect 845 1604 849 1608
rect 899 1604 903 1608
rect 255 1555 259 1559
rect 285 1555 289 1559
rect 313 1555 317 1559
rect 579 1472 583 1476
rect 614 1472 618 1476
rect 740 1472 744 1476
rect 764 1472 768 1476
rect 818 1472 822 1476
rect 845 1472 849 1476
rect 869 1472 873 1476
rect 579 1340 583 1344
rect 614 1340 618 1344
rect 740 1340 744 1344
rect 764 1340 768 1344
rect 818 1340 825 1344
rect 845 1340 849 1344
rect 899 1340 903 1344
rect 935 1340 939 1344
rect 989 1340 993 1344
rect 579 1208 583 1212
rect 614 1208 618 1212
rect 740 1208 744 1212
rect 764 1208 768 1212
rect 875 1208 879 1212
rect 126 1155 130 1159
rect 154 1155 158 1159
rect 184 1155 188 1159
rect 258 1155 262 1159
rect 286 1155 290 1159
rect 316 1155 320 1159
rect 390 1155 394 1159
rect 418 1155 422 1159
rect 448 1155 452 1159
rect 897 1045 901 1049
rect 925 1045 929 1049
rect 955 1045 959 1049
rect 126 1015 130 1019
rect 154 1015 158 1019
rect 184 1015 188 1019
rect 258 1015 262 1019
rect 286 1015 290 1019
rect 316 1015 320 1019
rect 390 1015 394 1019
rect 418 1015 422 1019
rect 448 1015 452 1019
rect 897 959 901 963
rect 925 959 929 963
rect 955 959 959 963
rect 126 929 130 933
rect 154 929 158 933
rect 184 929 188 933
rect 258 929 262 933
rect 286 929 290 933
rect 316 929 320 933
rect 390 929 394 933
rect 418 929 422 933
rect 448 929 452 933
rect 126 789 130 793
rect 154 789 158 793
rect 184 789 188 793
rect 258 789 262 793
rect 286 789 290 793
rect 316 789 320 793
rect 390 789 394 793
rect 418 789 422 793
rect 448 789 452 793
<< nsubstratencontact >>
rect 598 1747 602 1751
rect 626 1747 630 1751
rect 656 1747 660 1751
rect 693 1747 697 1751
rect 730 1747 734 1751
rect 758 1747 762 1751
rect 788 1747 792 1751
rect 825 1747 829 1751
rect 862 1747 866 1751
rect 890 1747 894 1751
rect 920 1747 924 1751
rect 957 1747 961 1751
rect 994 1747 998 1751
rect 1022 1747 1026 1751
rect 1052 1747 1056 1751
rect 1089 1747 1093 1751
rect 258 1714 262 1718
rect 286 1714 290 1718
rect 316 1714 320 1718
rect 353 1714 357 1718
rect 588 1670 592 1674
rect 617 1670 621 1674
rect 642 1670 646 1674
rect 684 1670 688 1674
rect 740 1670 744 1674
rect 764 1670 768 1674
rect 818 1670 822 1674
rect 845 1670 849 1674
rect 899 1670 903 1674
rect 218 1612 222 1616
rect 255 1612 259 1616
rect 285 1612 289 1616
rect 313 1612 317 1616
rect 588 1538 592 1542
rect 617 1538 621 1542
rect 642 1538 646 1542
rect 684 1538 688 1542
rect 740 1538 744 1542
rect 764 1538 768 1542
rect 818 1538 822 1542
rect 845 1538 849 1542
rect 907 1538 911 1542
rect 588 1406 592 1410
rect 617 1406 621 1410
rect 642 1406 646 1410
rect 684 1406 688 1410
rect 740 1406 744 1410
rect 764 1406 768 1410
rect 818 1406 822 1410
rect 845 1406 849 1410
rect 899 1406 903 1410
rect 907 1406 911 1410
rect 935 1406 939 1410
rect 989 1406 993 1410
rect 588 1274 592 1278
rect 617 1274 621 1278
rect 642 1274 646 1278
rect 684 1274 688 1278
rect 740 1274 744 1278
rect 764 1274 768 1278
rect 818 1274 822 1278
rect 845 1274 849 1278
rect 935 1274 939 1278
rect 126 1212 130 1216
rect 154 1212 158 1216
rect 184 1212 188 1216
rect 221 1212 225 1216
rect 258 1212 262 1216
rect 286 1212 290 1216
rect 316 1212 320 1216
rect 353 1212 357 1216
rect 390 1212 394 1216
rect 418 1212 422 1216
rect 448 1212 452 1216
rect 485 1212 489 1216
rect 588 1142 592 1146
rect 617 1142 621 1146
rect 642 1142 646 1146
rect 684 1142 688 1146
rect 764 1142 768 1146
rect 818 1142 822 1146
rect 849 1142 853 1146
rect 878 1142 882 1146
rect 903 1142 907 1146
rect 945 1142 949 1146
rect 897 1102 901 1106
rect 925 1102 929 1106
rect 955 1102 959 1106
rect 992 1102 996 1106
rect 126 1072 130 1076
rect 154 1072 158 1076
rect 184 1072 188 1076
rect 221 1072 225 1076
rect 258 1072 262 1076
rect 286 1072 290 1076
rect 316 1072 320 1076
rect 353 1072 357 1076
rect 390 1072 394 1076
rect 418 1072 422 1076
rect 448 1072 452 1076
rect 485 1072 489 1076
rect 897 1016 901 1020
rect 925 1016 929 1020
rect 955 1016 959 1020
rect 992 1016 996 1020
rect 126 986 130 990
rect 154 986 158 990
rect 184 986 188 990
rect 221 986 225 990
rect 258 986 262 990
rect 286 986 290 990
rect 316 986 320 990
rect 353 986 357 990
rect 390 986 394 990
rect 418 986 422 990
rect 448 986 452 990
rect 485 986 489 990
rect 126 846 130 850
rect 154 846 158 850
rect 184 846 188 850
rect 221 846 225 850
rect 258 846 262 850
rect 286 846 290 850
rect 316 846 320 850
rect 353 846 357 850
rect 390 846 394 850
rect 418 846 422 850
rect 448 846 452 850
rect 485 846 489 850
<< polysilicon >>
rect 573 1737 575 1739
rect 578 1737 580 1740
rect 594 1737 596 1739
rect 610 1737 612 1739
rect 615 1737 617 1740
rect 636 1737 638 1740
rect 652 1737 654 1740
rect 668 1737 670 1739
rect 673 1737 675 1740
rect 689 1737 691 1739
rect 705 1737 707 1739
rect 710 1737 712 1740
rect 726 1737 728 1739
rect 742 1737 744 1739
rect 747 1737 749 1740
rect 768 1737 770 1740
rect 784 1737 786 1740
rect 800 1737 802 1739
rect 805 1737 807 1740
rect 821 1737 823 1739
rect 837 1737 839 1739
rect 842 1737 844 1740
rect 858 1737 860 1739
rect 874 1737 876 1739
rect 879 1737 881 1740
rect 900 1737 902 1740
rect 916 1737 918 1740
rect 932 1737 934 1739
rect 937 1737 939 1740
rect 953 1737 955 1739
rect 969 1737 971 1739
rect 974 1737 976 1740
rect 990 1737 992 1739
rect 1006 1737 1008 1739
rect 1011 1737 1013 1740
rect 1032 1737 1034 1740
rect 1048 1737 1050 1740
rect 1064 1737 1066 1739
rect 1069 1737 1071 1740
rect 1085 1737 1087 1739
rect 573 1724 575 1729
rect 578 1727 580 1729
rect 573 1710 575 1720
rect 578 1710 580 1717
rect 594 1710 596 1729
rect 610 1720 612 1729
rect 615 1727 617 1729
rect 636 1727 638 1729
rect 652 1726 654 1729
rect 610 1710 612 1713
rect 615 1710 617 1712
rect 636 1710 638 1712
rect 652 1710 654 1722
rect 668 1720 670 1729
rect 673 1727 675 1729
rect 689 1721 691 1729
rect 705 1724 707 1729
rect 710 1727 712 1729
rect 668 1710 670 1713
rect 673 1710 675 1712
rect 689 1710 691 1717
rect 705 1710 707 1720
rect 710 1710 712 1717
rect 726 1710 728 1729
rect 742 1720 744 1729
rect 747 1727 749 1729
rect 768 1727 770 1729
rect 784 1726 786 1729
rect 742 1710 744 1713
rect 747 1710 749 1712
rect 768 1710 770 1712
rect 784 1710 786 1722
rect 800 1720 802 1729
rect 805 1727 807 1729
rect 821 1721 823 1729
rect 837 1724 839 1729
rect 842 1727 844 1729
rect 800 1710 802 1713
rect 805 1710 807 1712
rect 821 1710 823 1717
rect 837 1710 839 1720
rect 842 1710 844 1717
rect 858 1710 860 1729
rect 874 1720 876 1729
rect 879 1727 881 1729
rect 900 1727 902 1729
rect 916 1726 918 1729
rect 874 1710 876 1713
rect 879 1710 881 1712
rect 900 1710 902 1712
rect 916 1710 918 1722
rect 932 1720 934 1729
rect 937 1727 939 1729
rect 953 1721 955 1729
rect 969 1724 971 1729
rect 974 1727 976 1729
rect 932 1710 934 1713
rect 937 1710 939 1712
rect 953 1710 955 1717
rect 969 1710 971 1720
rect 974 1710 976 1717
rect 990 1710 992 1729
rect 1006 1720 1008 1729
rect 1011 1727 1013 1729
rect 1032 1727 1034 1729
rect 1048 1726 1050 1729
rect 1006 1710 1008 1713
rect 1011 1710 1013 1712
rect 1032 1710 1034 1712
rect 1048 1710 1050 1722
rect 1064 1720 1066 1729
rect 1069 1727 1071 1729
rect 1085 1721 1087 1729
rect 1064 1710 1066 1713
rect 1069 1710 1071 1712
rect 1085 1710 1087 1717
rect 233 1704 235 1706
rect 238 1704 240 1707
rect 254 1704 256 1706
rect 270 1704 272 1706
rect 275 1704 277 1707
rect 296 1704 298 1707
rect 312 1704 314 1707
rect 328 1704 330 1706
rect 333 1704 335 1707
rect 349 1704 351 1706
rect 573 1704 575 1706
rect 578 1703 580 1706
rect 594 1704 596 1706
rect 610 1704 612 1706
rect 615 1701 617 1706
rect 636 1701 638 1706
rect 652 1704 654 1706
rect 668 1704 670 1706
rect 673 1701 675 1706
rect 689 1704 691 1706
rect 705 1704 707 1706
rect 710 1703 712 1706
rect 726 1704 728 1706
rect 742 1704 744 1706
rect 747 1701 749 1706
rect 768 1701 770 1706
rect 784 1704 786 1706
rect 800 1704 802 1706
rect 805 1701 807 1706
rect 821 1704 823 1706
rect 837 1704 839 1706
rect 842 1703 844 1706
rect 858 1704 860 1706
rect 874 1704 876 1706
rect 879 1701 881 1706
rect 900 1701 902 1706
rect 916 1704 918 1706
rect 932 1704 934 1706
rect 937 1701 939 1706
rect 953 1704 955 1706
rect 969 1704 971 1706
rect 974 1703 976 1706
rect 990 1704 992 1706
rect 1006 1704 1008 1706
rect 1011 1701 1013 1706
rect 1032 1701 1034 1706
rect 1048 1704 1050 1706
rect 1064 1704 1066 1706
rect 1069 1701 1071 1706
rect 1085 1704 1087 1706
rect 233 1691 235 1696
rect 238 1694 240 1696
rect 233 1677 235 1687
rect 238 1677 240 1684
rect 254 1677 256 1696
rect 270 1687 272 1696
rect 275 1694 277 1696
rect 296 1694 298 1696
rect 312 1693 314 1696
rect 270 1677 272 1680
rect 275 1677 277 1679
rect 296 1677 298 1679
rect 312 1677 314 1689
rect 328 1687 330 1696
rect 333 1694 335 1696
rect 328 1677 330 1680
rect 333 1677 335 1679
rect 349 1677 351 1696
rect 233 1671 235 1673
rect 238 1670 240 1673
rect 254 1671 256 1673
rect 270 1671 272 1673
rect 275 1668 277 1673
rect 296 1668 298 1673
rect 312 1671 314 1673
rect 328 1671 330 1673
rect 333 1668 335 1673
rect 349 1671 351 1673
rect 752 1666 754 1668
rect 594 1660 596 1663
rect 638 1660 640 1663
rect 664 1660 666 1663
rect 710 1660 712 1663
rect 664 1656 665 1660
rect 778 1660 780 1664
rect 806 1666 808 1668
rect 833 1666 835 1668
rect 783 1660 785 1663
rect 578 1653 580 1655
rect 594 1653 596 1656
rect 610 1653 612 1655
rect 633 1653 635 1655
rect 638 1653 640 1656
rect 664 1653 666 1656
rect 685 1653 687 1656
rect 705 1653 707 1655
rect 710 1653 712 1656
rect 728 1653 730 1655
rect 357 1640 359 1643
rect 357 1634 359 1636
rect 240 1631 242 1634
rect 578 1631 580 1645
rect 594 1643 596 1645
rect 594 1631 596 1633
rect 610 1631 612 1645
rect 633 1640 635 1645
rect 638 1643 640 1645
rect 664 1643 666 1645
rect 629 1636 635 1640
rect 633 1631 635 1636
rect 638 1631 640 1633
rect 664 1631 666 1633
rect 685 1631 687 1645
rect 705 1640 707 1645
rect 710 1643 712 1645
rect 701 1636 707 1640
rect 705 1631 707 1636
rect 710 1631 712 1633
rect 728 1631 730 1645
rect 752 1644 754 1658
rect 859 1660 861 1664
rect 887 1666 889 1668
rect 864 1660 866 1663
rect 778 1649 780 1652
rect 783 1650 785 1652
rect 779 1645 780 1649
rect 778 1640 780 1645
rect 783 1640 785 1642
rect 752 1638 754 1640
rect 806 1636 808 1658
rect 833 1644 835 1658
rect 859 1649 861 1652
rect 864 1650 866 1652
rect 860 1645 861 1649
rect 859 1640 861 1645
rect 864 1640 866 1642
rect 833 1638 835 1640
rect 887 1636 889 1658
rect 778 1634 780 1636
rect 783 1631 785 1636
rect 859 1634 861 1636
rect 806 1630 808 1632
rect 864 1631 866 1636
rect 887 1630 889 1632
rect 240 1625 242 1627
rect 578 1625 580 1627
rect 594 1623 596 1627
rect 610 1625 612 1627
rect 633 1625 635 1627
rect 595 1619 596 1623
rect 638 1622 640 1627
rect 664 1623 666 1627
rect 685 1625 687 1627
rect 705 1625 707 1627
rect 594 1616 596 1619
rect 639 1618 640 1622
rect 665 1619 666 1623
rect 710 1622 712 1627
rect 728 1625 730 1627
rect 638 1616 640 1618
rect 664 1615 666 1619
rect 711 1618 712 1622
rect 710 1616 712 1618
rect 224 1602 226 1604
rect 240 1602 242 1605
rect 245 1602 247 1604
rect 261 1602 263 1605
rect 277 1602 279 1605
rect 298 1602 300 1605
rect 303 1602 305 1604
rect 319 1602 321 1604
rect 335 1602 337 1605
rect 340 1602 342 1604
rect 224 1575 226 1594
rect 240 1592 242 1594
rect 245 1585 247 1594
rect 261 1591 263 1594
rect 277 1592 279 1594
rect 298 1592 300 1594
rect 240 1575 242 1577
rect 245 1575 247 1578
rect 261 1575 263 1587
rect 303 1585 305 1594
rect 277 1575 279 1577
rect 298 1575 300 1577
rect 303 1575 305 1578
rect 319 1575 321 1594
rect 335 1592 337 1594
rect 340 1589 342 1594
rect 594 1593 596 1596
rect 638 1594 640 1596
rect 595 1589 596 1593
rect 639 1590 640 1594
rect 664 1593 666 1597
rect 710 1594 712 1596
rect 578 1585 580 1587
rect 594 1585 596 1589
rect 610 1585 612 1587
rect 633 1585 635 1587
rect 638 1585 640 1590
rect 665 1589 666 1593
rect 711 1590 712 1594
rect 664 1585 666 1589
rect 685 1585 687 1587
rect 705 1585 707 1587
rect 710 1585 712 1590
rect 728 1585 730 1587
rect 335 1575 337 1582
rect 340 1575 342 1585
rect 778 1584 780 1587
rect 783 1584 785 1587
rect 859 1584 861 1587
rect 864 1584 866 1587
rect 224 1569 226 1571
rect 240 1566 242 1571
rect 245 1569 247 1571
rect 261 1569 263 1571
rect 277 1566 279 1571
rect 298 1566 300 1571
rect 303 1569 305 1571
rect 319 1569 321 1571
rect 335 1568 337 1571
rect 340 1569 342 1571
rect 578 1567 580 1581
rect 594 1579 596 1581
rect 594 1567 596 1569
rect 610 1567 612 1581
rect 633 1576 635 1581
rect 638 1579 640 1581
rect 664 1579 666 1581
rect 629 1572 635 1576
rect 633 1567 635 1572
rect 638 1567 640 1569
rect 664 1567 666 1569
rect 685 1567 687 1581
rect 705 1576 707 1581
rect 710 1579 712 1581
rect 701 1572 707 1576
rect 705 1567 707 1572
rect 710 1567 712 1569
rect 728 1567 730 1581
rect 778 1568 780 1580
rect 783 1578 785 1580
rect 783 1568 785 1570
rect 859 1568 861 1580
rect 864 1578 866 1580
rect 864 1568 866 1570
rect 578 1557 580 1559
rect 594 1556 596 1559
rect 610 1557 612 1559
rect 633 1557 635 1559
rect 638 1556 640 1559
rect 664 1556 666 1559
rect 685 1556 687 1559
rect 705 1557 707 1559
rect 710 1556 712 1559
rect 728 1557 730 1559
rect 778 1558 780 1560
rect 664 1552 665 1556
rect 783 1555 785 1560
rect 859 1558 861 1560
rect 864 1555 866 1560
rect 594 1549 596 1552
rect 638 1549 640 1552
rect 664 1549 666 1552
rect 710 1549 712 1552
rect 594 1528 596 1531
rect 638 1528 640 1531
rect 664 1528 666 1531
rect 710 1528 712 1531
rect 778 1528 780 1532
rect 806 1534 808 1536
rect 857 1534 859 1536
rect 783 1528 785 1531
rect 664 1524 665 1528
rect 578 1521 580 1523
rect 594 1521 596 1524
rect 610 1521 612 1523
rect 633 1521 635 1523
rect 638 1521 640 1524
rect 664 1521 666 1524
rect 685 1521 687 1524
rect 705 1521 707 1523
rect 710 1521 712 1524
rect 728 1521 730 1523
rect 883 1528 885 1532
rect 911 1534 913 1536
rect 888 1528 890 1531
rect 778 1517 780 1520
rect 783 1518 785 1520
rect 779 1513 780 1517
rect 578 1499 580 1513
rect 594 1511 596 1513
rect 594 1499 596 1501
rect 610 1499 612 1513
rect 633 1508 635 1513
rect 638 1511 640 1513
rect 664 1511 666 1513
rect 629 1504 635 1508
rect 633 1499 635 1504
rect 638 1499 640 1501
rect 664 1499 666 1501
rect 685 1499 687 1513
rect 705 1508 707 1513
rect 710 1511 712 1513
rect 701 1504 707 1508
rect 705 1499 707 1504
rect 710 1499 712 1501
rect 728 1499 730 1513
rect 778 1508 780 1513
rect 783 1508 785 1510
rect 806 1504 808 1526
rect 857 1512 859 1526
rect 883 1517 885 1520
rect 888 1518 890 1520
rect 884 1513 885 1517
rect 883 1508 885 1513
rect 888 1508 890 1510
rect 857 1506 859 1508
rect 911 1504 913 1526
rect 778 1502 780 1504
rect 783 1499 785 1504
rect 883 1502 885 1504
rect 806 1498 808 1500
rect 888 1499 890 1504
rect 911 1498 913 1500
rect 578 1493 580 1495
rect 594 1491 596 1495
rect 610 1493 612 1495
rect 633 1493 635 1495
rect 595 1487 596 1491
rect 638 1490 640 1495
rect 664 1491 666 1495
rect 685 1493 687 1495
rect 705 1493 707 1495
rect 594 1484 596 1487
rect 639 1486 640 1490
rect 665 1487 666 1491
rect 710 1490 712 1495
rect 728 1493 730 1495
rect 638 1484 640 1486
rect 664 1483 666 1487
rect 711 1486 712 1490
rect 710 1484 712 1486
rect 594 1461 596 1464
rect 638 1462 640 1464
rect 595 1457 596 1461
rect 639 1458 640 1462
rect 664 1461 666 1465
rect 710 1462 712 1464
rect 578 1453 580 1455
rect 594 1453 596 1457
rect 610 1453 612 1455
rect 633 1453 635 1455
rect 638 1453 640 1458
rect 665 1457 666 1461
rect 711 1458 712 1462
rect 664 1453 666 1457
rect 685 1453 687 1455
rect 705 1453 707 1455
rect 710 1453 712 1458
rect 728 1453 730 1455
rect 778 1453 780 1456
rect 783 1453 785 1456
rect 883 1453 885 1456
rect 888 1453 890 1456
rect 578 1435 580 1449
rect 594 1447 596 1449
rect 594 1435 596 1437
rect 610 1435 612 1449
rect 633 1444 635 1449
rect 638 1447 640 1449
rect 664 1447 666 1449
rect 629 1440 635 1444
rect 633 1435 635 1440
rect 638 1435 640 1437
rect 664 1435 666 1437
rect 685 1435 687 1449
rect 705 1444 707 1449
rect 710 1447 712 1449
rect 701 1440 707 1444
rect 705 1435 707 1440
rect 710 1435 712 1437
rect 728 1435 730 1449
rect 778 1437 780 1449
rect 783 1447 785 1449
rect 783 1437 785 1439
rect 883 1437 885 1449
rect 888 1447 890 1449
rect 888 1437 890 1439
rect 778 1427 780 1429
rect 578 1425 580 1427
rect 594 1424 596 1427
rect 610 1425 612 1427
rect 633 1425 635 1427
rect 638 1424 640 1427
rect 664 1424 666 1427
rect 685 1424 687 1427
rect 705 1425 707 1427
rect 710 1424 712 1427
rect 728 1425 730 1427
rect 783 1424 785 1429
rect 883 1427 885 1429
rect 888 1424 890 1429
rect 664 1420 665 1424
rect 594 1417 596 1420
rect 638 1417 640 1420
rect 664 1417 666 1420
rect 710 1417 712 1420
rect 594 1396 596 1399
rect 638 1396 640 1399
rect 664 1396 666 1399
rect 710 1396 712 1399
rect 778 1396 780 1400
rect 806 1402 808 1404
rect 833 1402 835 1404
rect 783 1396 785 1399
rect 664 1392 665 1396
rect 578 1389 580 1391
rect 594 1389 596 1392
rect 610 1389 612 1391
rect 633 1389 635 1391
rect 638 1389 640 1392
rect 664 1389 666 1392
rect 685 1389 687 1392
rect 705 1389 707 1391
rect 710 1389 712 1392
rect 728 1389 730 1391
rect 859 1396 861 1400
rect 887 1402 889 1404
rect 923 1402 925 1404
rect 864 1396 866 1399
rect 778 1385 780 1388
rect 783 1386 785 1388
rect 779 1381 780 1385
rect 578 1367 580 1381
rect 594 1379 596 1381
rect 594 1367 596 1369
rect 610 1367 612 1381
rect 633 1376 635 1381
rect 638 1379 640 1381
rect 664 1379 666 1381
rect 629 1372 635 1376
rect 633 1367 635 1372
rect 638 1367 640 1369
rect 664 1367 666 1369
rect 685 1367 687 1381
rect 705 1376 707 1381
rect 710 1379 712 1381
rect 701 1372 707 1376
rect 705 1367 707 1372
rect 710 1367 712 1369
rect 728 1367 730 1381
rect 778 1376 780 1381
rect 783 1376 785 1378
rect 806 1372 808 1394
rect 833 1380 835 1394
rect 949 1396 951 1400
rect 977 1402 979 1404
rect 954 1396 956 1399
rect 859 1385 861 1388
rect 864 1386 866 1388
rect 860 1381 861 1385
rect 859 1376 861 1381
rect 864 1376 866 1378
rect 833 1374 835 1376
rect 887 1372 889 1394
rect 923 1380 925 1394
rect 949 1385 951 1388
rect 954 1386 956 1388
rect 950 1381 951 1385
rect 949 1376 951 1381
rect 954 1376 956 1378
rect 923 1374 925 1376
rect 977 1372 979 1394
rect 778 1370 780 1372
rect 783 1367 785 1372
rect 859 1370 861 1372
rect 806 1366 808 1368
rect 864 1367 866 1372
rect 949 1370 951 1372
rect 887 1366 889 1368
rect 954 1367 956 1372
rect 977 1366 979 1368
rect 578 1361 580 1363
rect 594 1359 596 1363
rect 610 1361 612 1363
rect 633 1361 635 1363
rect 595 1355 596 1359
rect 638 1358 640 1363
rect 664 1359 666 1363
rect 685 1361 687 1363
rect 705 1361 707 1363
rect 594 1352 596 1355
rect 639 1354 640 1358
rect 665 1355 666 1359
rect 710 1358 712 1363
rect 728 1361 730 1363
rect 638 1352 640 1354
rect 664 1351 666 1355
rect 711 1354 712 1358
rect 710 1352 712 1354
rect 594 1329 596 1332
rect 638 1330 640 1332
rect 595 1325 596 1329
rect 639 1326 640 1330
rect 664 1329 666 1333
rect 710 1330 712 1332
rect 578 1321 580 1323
rect 594 1321 596 1325
rect 610 1321 612 1323
rect 633 1321 635 1323
rect 638 1321 640 1326
rect 665 1325 666 1329
rect 711 1326 712 1330
rect 664 1321 666 1325
rect 685 1321 687 1323
rect 705 1321 707 1323
rect 710 1321 712 1326
rect 728 1321 730 1323
rect 778 1318 780 1321
rect 783 1318 785 1321
rect 859 1318 861 1321
rect 864 1318 866 1321
rect 949 1318 951 1321
rect 954 1318 956 1321
rect 578 1303 580 1317
rect 594 1315 596 1317
rect 594 1303 596 1305
rect 610 1303 612 1317
rect 633 1312 635 1317
rect 638 1315 640 1317
rect 664 1315 666 1317
rect 629 1308 635 1312
rect 633 1303 635 1308
rect 638 1303 640 1305
rect 664 1303 666 1305
rect 685 1303 687 1317
rect 705 1312 707 1317
rect 710 1315 712 1317
rect 701 1308 707 1312
rect 705 1303 707 1308
rect 710 1303 712 1305
rect 728 1303 730 1317
rect 778 1302 780 1314
rect 783 1312 785 1314
rect 783 1302 785 1304
rect 859 1302 861 1314
rect 864 1312 866 1314
rect 864 1302 866 1304
rect 949 1302 951 1314
rect 954 1312 956 1314
rect 954 1302 956 1304
rect 578 1293 580 1295
rect 594 1292 596 1295
rect 610 1293 612 1295
rect 633 1293 635 1295
rect 638 1292 640 1295
rect 664 1292 666 1295
rect 685 1292 687 1295
rect 705 1293 707 1295
rect 710 1292 712 1295
rect 728 1293 730 1295
rect 778 1292 780 1294
rect 664 1288 665 1292
rect 783 1289 785 1294
rect 859 1292 861 1294
rect 864 1289 866 1294
rect 949 1292 951 1294
rect 954 1289 956 1294
rect 594 1285 596 1288
rect 638 1285 640 1288
rect 664 1285 666 1288
rect 710 1285 712 1288
rect 594 1264 596 1267
rect 638 1264 640 1267
rect 664 1264 666 1267
rect 710 1264 712 1267
rect 778 1264 780 1268
rect 806 1270 808 1272
rect 783 1264 785 1267
rect 664 1260 665 1264
rect 578 1257 580 1259
rect 594 1257 596 1260
rect 610 1257 612 1259
rect 633 1257 635 1259
rect 638 1257 640 1260
rect 664 1257 666 1260
rect 685 1257 687 1260
rect 705 1257 707 1259
rect 710 1257 712 1260
rect 728 1257 730 1259
rect 778 1253 780 1256
rect 783 1254 785 1256
rect 779 1249 780 1253
rect 578 1235 580 1249
rect 594 1247 596 1249
rect 594 1235 596 1237
rect 610 1235 612 1249
rect 633 1244 635 1249
rect 638 1247 640 1249
rect 664 1247 666 1249
rect 629 1240 635 1244
rect 633 1235 635 1240
rect 638 1235 640 1237
rect 664 1235 666 1237
rect 685 1235 687 1249
rect 705 1244 707 1249
rect 710 1247 712 1249
rect 701 1240 707 1244
rect 705 1235 707 1240
rect 710 1235 712 1237
rect 728 1235 730 1249
rect 778 1244 780 1249
rect 783 1244 785 1246
rect 806 1240 808 1262
rect 778 1238 780 1240
rect 783 1235 785 1240
rect 806 1234 808 1236
rect 578 1229 580 1231
rect 594 1227 596 1231
rect 610 1229 612 1231
rect 633 1229 635 1231
rect 595 1223 596 1227
rect 638 1226 640 1231
rect 664 1227 666 1231
rect 685 1229 687 1231
rect 705 1229 707 1231
rect 594 1220 596 1223
rect 639 1222 640 1226
rect 665 1223 666 1227
rect 710 1226 712 1231
rect 728 1229 730 1231
rect 638 1220 640 1222
rect 664 1219 666 1223
rect 711 1222 712 1226
rect 710 1220 712 1222
rect 101 1202 103 1204
rect 106 1202 108 1205
rect 122 1202 124 1204
rect 138 1202 140 1204
rect 143 1202 145 1205
rect 164 1202 166 1205
rect 180 1202 182 1205
rect 196 1202 198 1204
rect 201 1202 203 1205
rect 217 1202 219 1204
rect 233 1202 235 1204
rect 238 1202 240 1205
rect 254 1202 256 1204
rect 270 1202 272 1204
rect 275 1202 277 1205
rect 296 1202 298 1205
rect 312 1202 314 1205
rect 328 1202 330 1204
rect 333 1202 335 1205
rect 349 1202 351 1204
rect 365 1202 367 1204
rect 370 1202 372 1205
rect 386 1202 388 1204
rect 402 1202 404 1204
rect 407 1202 409 1205
rect 428 1202 430 1205
rect 444 1202 446 1205
rect 460 1202 462 1204
rect 465 1202 467 1205
rect 481 1202 483 1204
rect 594 1197 596 1200
rect 638 1198 640 1200
rect 101 1189 103 1194
rect 106 1192 108 1194
rect 101 1175 103 1185
rect 106 1175 108 1182
rect 122 1175 124 1194
rect 138 1185 140 1194
rect 143 1192 145 1194
rect 164 1192 166 1194
rect 180 1191 182 1194
rect 138 1175 140 1178
rect 143 1175 145 1177
rect 164 1175 166 1177
rect 180 1175 182 1187
rect 196 1185 198 1194
rect 201 1192 203 1194
rect 196 1175 198 1178
rect 201 1175 203 1177
rect 217 1175 219 1194
rect 233 1191 235 1194
rect 238 1192 240 1194
rect 233 1175 235 1187
rect 238 1175 240 1182
rect 254 1175 256 1194
rect 270 1185 272 1194
rect 275 1192 277 1194
rect 296 1192 298 1194
rect 312 1191 314 1194
rect 270 1175 272 1178
rect 275 1175 277 1177
rect 296 1175 298 1177
rect 312 1175 314 1187
rect 328 1185 330 1194
rect 333 1192 335 1194
rect 328 1175 330 1178
rect 333 1175 335 1177
rect 349 1175 351 1194
rect 365 1191 367 1194
rect 370 1192 372 1194
rect 365 1175 367 1187
rect 370 1175 372 1182
rect 386 1175 388 1194
rect 402 1185 404 1194
rect 407 1192 409 1194
rect 428 1192 430 1194
rect 444 1191 446 1194
rect 402 1175 404 1178
rect 407 1175 409 1177
rect 428 1175 430 1177
rect 444 1175 446 1187
rect 460 1185 462 1194
rect 465 1192 467 1194
rect 481 1186 483 1194
rect 595 1193 596 1197
rect 639 1194 640 1198
rect 664 1197 666 1201
rect 710 1198 712 1200
rect 578 1189 580 1191
rect 594 1189 596 1193
rect 610 1189 612 1191
rect 633 1189 635 1191
rect 638 1189 640 1194
rect 665 1193 666 1197
rect 711 1194 712 1198
rect 855 1197 857 1200
rect 899 1198 901 1200
rect 664 1189 666 1193
rect 685 1189 687 1191
rect 705 1189 707 1191
rect 710 1189 712 1194
rect 856 1193 857 1197
rect 900 1194 901 1198
rect 925 1197 927 1201
rect 971 1198 973 1200
rect 728 1189 730 1191
rect 812 1189 814 1192
rect 830 1189 832 1192
rect 855 1189 857 1193
rect 871 1189 873 1191
rect 894 1189 896 1191
rect 899 1189 901 1194
rect 926 1193 927 1197
rect 972 1194 973 1198
rect 925 1189 927 1193
rect 946 1189 948 1191
rect 966 1189 968 1191
rect 971 1189 973 1194
rect 989 1189 991 1191
rect 460 1175 462 1178
rect 465 1175 467 1177
rect 481 1175 483 1182
rect 578 1171 580 1185
rect 594 1183 596 1185
rect 594 1171 596 1173
rect 610 1171 612 1185
rect 633 1180 635 1185
rect 638 1183 640 1185
rect 664 1183 666 1185
rect 629 1176 635 1180
rect 633 1171 635 1176
rect 638 1171 640 1173
rect 664 1171 666 1173
rect 685 1171 687 1185
rect 705 1180 707 1185
rect 710 1183 712 1185
rect 701 1176 707 1180
rect 705 1171 707 1176
rect 710 1171 712 1173
rect 728 1171 730 1185
rect 778 1182 780 1185
rect 783 1182 785 1185
rect 812 1180 814 1185
rect 101 1169 103 1171
rect 106 1168 108 1171
rect 122 1169 124 1171
rect 138 1169 140 1171
rect 143 1166 145 1171
rect 164 1166 166 1171
rect 180 1169 182 1171
rect 196 1169 198 1171
rect 201 1166 203 1171
rect 217 1169 219 1171
rect 233 1169 235 1171
rect 238 1168 240 1171
rect 254 1169 256 1171
rect 270 1169 272 1171
rect 275 1166 277 1171
rect 296 1166 298 1171
rect 312 1169 314 1171
rect 328 1169 330 1171
rect 333 1166 335 1171
rect 349 1169 351 1171
rect 365 1169 367 1171
rect 370 1168 372 1171
rect 386 1169 388 1171
rect 402 1169 404 1171
rect 407 1166 409 1171
rect 428 1166 430 1171
rect 444 1169 446 1171
rect 460 1169 462 1171
rect 465 1166 467 1171
rect 481 1169 483 1171
rect 778 1166 780 1178
rect 783 1176 785 1178
rect 812 1171 814 1176
rect 830 1171 832 1185
rect 855 1183 857 1185
rect 855 1171 857 1173
rect 871 1171 873 1185
rect 894 1180 896 1185
rect 899 1183 901 1185
rect 925 1183 927 1185
rect 890 1176 896 1180
rect 894 1171 896 1176
rect 899 1171 901 1173
rect 925 1171 927 1173
rect 946 1171 948 1185
rect 966 1180 968 1185
rect 971 1183 973 1185
rect 962 1176 968 1180
rect 966 1171 968 1176
rect 971 1171 973 1173
rect 989 1171 991 1185
rect 783 1166 785 1168
rect 578 1161 580 1163
rect 594 1160 596 1163
rect 610 1161 612 1163
rect 633 1161 635 1163
rect 638 1160 640 1163
rect 664 1160 666 1163
rect 685 1160 687 1163
rect 705 1161 707 1163
rect 710 1160 712 1163
rect 728 1161 730 1163
rect 664 1156 665 1160
rect 812 1160 814 1163
rect 830 1160 832 1163
rect 855 1160 857 1163
rect 871 1161 873 1163
rect 894 1161 896 1163
rect 899 1160 901 1163
rect 925 1160 927 1163
rect 946 1160 948 1163
rect 966 1161 968 1163
rect 971 1160 973 1163
rect 989 1161 991 1163
rect 778 1156 780 1158
rect 594 1153 596 1156
rect 638 1153 640 1156
rect 664 1153 666 1156
rect 710 1153 712 1156
rect 783 1153 785 1158
rect 925 1156 926 1160
rect 855 1153 857 1156
rect 899 1153 901 1156
rect 925 1153 927 1156
rect 971 1153 973 1156
rect 216 1131 218 1134
rect 240 1131 242 1134
rect 998 1129 1001 1131
rect 1005 1129 1008 1131
rect 216 1125 218 1127
rect 240 1125 242 1127
rect 236 1120 238 1122
rect 236 1113 238 1116
rect 225 1102 227 1104
rect 231 1102 250 1104
rect 216 1097 218 1099
rect 240 1097 242 1099
rect 216 1090 218 1093
rect 240 1090 242 1093
rect 872 1092 874 1094
rect 877 1092 879 1095
rect 893 1092 895 1094
rect 909 1092 911 1094
rect 914 1092 916 1095
rect 935 1092 937 1095
rect 951 1092 953 1095
rect 967 1092 969 1094
rect 972 1092 974 1095
rect 988 1092 990 1094
rect 872 1079 874 1084
rect 877 1082 879 1084
rect 872 1065 874 1075
rect 877 1065 879 1072
rect 893 1065 895 1084
rect 909 1075 911 1084
rect 914 1082 916 1084
rect 935 1082 937 1084
rect 951 1081 953 1084
rect 909 1065 911 1068
rect 914 1065 916 1067
rect 935 1065 937 1067
rect 951 1065 953 1077
rect 967 1075 969 1084
rect 972 1082 974 1084
rect 967 1065 969 1068
rect 972 1065 974 1067
rect 988 1065 990 1084
rect 101 1062 103 1064
rect 106 1062 108 1065
rect 122 1062 124 1064
rect 138 1062 140 1064
rect 143 1062 145 1065
rect 164 1062 166 1065
rect 180 1062 182 1065
rect 196 1062 198 1064
rect 201 1062 203 1065
rect 217 1062 219 1064
rect 233 1062 235 1064
rect 238 1062 240 1065
rect 254 1062 256 1064
rect 270 1062 272 1064
rect 275 1062 277 1065
rect 296 1062 298 1065
rect 312 1062 314 1065
rect 328 1062 330 1064
rect 333 1062 335 1065
rect 349 1062 351 1064
rect 365 1062 367 1064
rect 370 1062 372 1065
rect 386 1062 388 1064
rect 402 1062 404 1064
rect 407 1062 409 1065
rect 428 1062 430 1065
rect 444 1062 446 1065
rect 460 1062 462 1064
rect 465 1062 467 1065
rect 481 1062 483 1064
rect 872 1059 874 1061
rect 877 1058 879 1061
rect 893 1059 895 1061
rect 909 1059 911 1061
rect 914 1056 916 1061
rect 935 1056 937 1061
rect 951 1059 953 1061
rect 967 1059 969 1061
rect 972 1056 974 1061
rect 988 1059 990 1061
rect 101 1049 103 1054
rect 106 1052 108 1054
rect 101 1035 103 1045
rect 106 1035 108 1042
rect 122 1035 124 1054
rect 138 1045 140 1054
rect 143 1052 145 1054
rect 164 1052 166 1054
rect 180 1051 182 1054
rect 138 1035 140 1038
rect 143 1035 145 1037
rect 164 1035 166 1037
rect 180 1035 182 1047
rect 196 1045 198 1054
rect 201 1052 203 1054
rect 196 1035 198 1038
rect 201 1035 203 1037
rect 217 1035 219 1054
rect 233 1051 235 1054
rect 238 1052 240 1054
rect 233 1035 235 1047
rect 238 1035 240 1042
rect 254 1035 256 1054
rect 270 1045 272 1054
rect 275 1052 277 1054
rect 296 1052 298 1054
rect 312 1051 314 1054
rect 270 1035 272 1038
rect 275 1035 277 1037
rect 296 1035 298 1037
rect 312 1035 314 1047
rect 328 1045 330 1054
rect 333 1052 335 1054
rect 328 1035 330 1038
rect 333 1035 335 1037
rect 349 1035 351 1054
rect 365 1051 367 1054
rect 370 1052 372 1054
rect 365 1035 367 1047
rect 370 1035 372 1042
rect 386 1035 388 1054
rect 402 1045 404 1054
rect 407 1052 409 1054
rect 428 1052 430 1054
rect 444 1051 446 1054
rect 402 1035 404 1038
rect 407 1035 409 1037
rect 428 1035 430 1037
rect 444 1035 446 1047
rect 460 1045 462 1054
rect 465 1052 467 1054
rect 481 1046 483 1054
rect 460 1035 462 1038
rect 465 1035 467 1037
rect 481 1035 483 1042
rect 101 1029 103 1031
rect 106 1028 108 1031
rect 122 1029 124 1031
rect 138 1029 140 1031
rect 143 1026 145 1031
rect 164 1026 166 1031
rect 180 1029 182 1031
rect 196 1029 198 1031
rect 201 1026 203 1031
rect 217 1029 219 1031
rect 233 1029 235 1031
rect 238 1028 240 1031
rect 254 1029 256 1031
rect 270 1029 272 1031
rect 275 1026 277 1031
rect 296 1026 298 1031
rect 312 1029 314 1031
rect 328 1029 330 1031
rect 333 1026 335 1031
rect 349 1029 351 1031
rect 365 1029 367 1031
rect 370 1028 372 1031
rect 386 1029 388 1031
rect 402 1029 404 1031
rect 407 1026 409 1031
rect 428 1026 430 1031
rect 444 1029 446 1031
rect 460 1029 462 1031
rect 465 1026 467 1031
rect 481 1029 483 1031
rect 872 1006 874 1008
rect 877 1006 879 1009
rect 893 1006 895 1008
rect 909 1006 911 1008
rect 914 1006 916 1009
rect 935 1006 937 1009
rect 951 1006 953 1009
rect 967 1006 969 1008
rect 972 1006 974 1009
rect 988 1006 990 1008
rect 872 993 874 998
rect 877 996 879 998
rect 872 979 874 989
rect 877 979 879 986
rect 893 979 895 998
rect 909 989 911 998
rect 914 996 916 998
rect 935 996 937 998
rect 951 995 953 998
rect 909 979 911 982
rect 914 979 916 981
rect 935 979 937 981
rect 951 979 953 991
rect 967 989 969 998
rect 972 996 974 998
rect 967 979 969 982
rect 972 979 974 981
rect 988 979 990 998
rect 1010 985 1013 987
rect 1017 985 1020 987
rect 101 976 103 978
rect 106 976 108 979
rect 122 976 124 978
rect 138 976 140 978
rect 143 976 145 979
rect 164 976 166 979
rect 180 976 182 979
rect 196 976 198 978
rect 201 976 203 979
rect 217 976 219 978
rect 233 976 235 978
rect 238 976 240 979
rect 254 976 256 978
rect 270 976 272 978
rect 275 976 277 979
rect 296 976 298 979
rect 312 976 314 979
rect 328 976 330 978
rect 333 976 335 979
rect 349 976 351 978
rect 365 976 367 978
rect 370 976 372 979
rect 386 976 388 978
rect 402 976 404 978
rect 407 976 409 979
rect 428 976 430 979
rect 444 976 446 979
rect 460 976 462 978
rect 465 976 467 979
rect 481 976 483 978
rect 872 973 874 975
rect 877 972 879 975
rect 893 973 895 975
rect 909 973 911 975
rect 914 970 916 975
rect 935 970 937 975
rect 951 973 953 975
rect 967 973 969 975
rect 972 970 974 975
rect 988 973 990 975
rect 101 963 103 968
rect 106 966 108 968
rect 101 949 103 959
rect 106 949 108 956
rect 122 949 124 968
rect 138 959 140 968
rect 143 966 145 968
rect 164 966 166 968
rect 180 965 182 968
rect 138 949 140 952
rect 143 949 145 951
rect 164 949 166 951
rect 180 949 182 961
rect 196 959 198 968
rect 201 966 203 968
rect 196 949 198 952
rect 201 949 203 951
rect 217 949 219 968
rect 233 965 235 968
rect 238 966 240 968
rect 233 949 235 961
rect 238 949 240 956
rect 254 949 256 968
rect 270 959 272 968
rect 275 966 277 968
rect 296 966 298 968
rect 312 965 314 968
rect 270 949 272 952
rect 275 949 277 951
rect 296 949 298 951
rect 312 949 314 961
rect 328 959 330 968
rect 333 966 335 968
rect 328 949 330 952
rect 333 949 335 951
rect 349 949 351 968
rect 365 965 367 968
rect 370 966 372 968
rect 365 949 367 961
rect 370 949 372 956
rect 386 949 388 968
rect 402 959 404 968
rect 407 966 409 968
rect 428 966 430 968
rect 444 965 446 968
rect 402 949 404 952
rect 407 949 409 951
rect 428 949 430 951
rect 444 949 446 961
rect 460 959 462 968
rect 465 966 467 968
rect 481 960 483 968
rect 460 949 462 952
rect 465 949 467 951
rect 481 949 483 956
rect 101 943 103 945
rect 106 942 108 945
rect 122 943 124 945
rect 138 943 140 945
rect 143 940 145 945
rect 164 940 166 945
rect 180 943 182 945
rect 196 943 198 945
rect 201 940 203 945
rect 217 943 219 945
rect 233 943 235 945
rect 238 942 240 945
rect 254 943 256 945
rect 270 943 272 945
rect 275 940 277 945
rect 296 940 298 945
rect 312 943 314 945
rect 328 943 330 945
rect 333 940 335 945
rect 349 943 351 945
rect 365 943 367 945
rect 370 942 372 945
rect 386 943 388 945
rect 402 943 404 945
rect 407 940 409 945
rect 428 940 430 945
rect 444 943 446 945
rect 460 943 462 945
rect 465 940 467 945
rect 481 943 483 945
rect 333 905 335 908
rect 357 905 359 908
rect 333 899 335 901
rect 357 899 359 901
rect 353 894 355 896
rect 353 887 355 890
rect 342 876 344 878
rect 348 876 367 878
rect 333 871 335 873
rect 357 871 359 873
rect 333 864 335 867
rect 357 864 359 867
rect 101 836 103 838
rect 106 836 108 839
rect 122 836 124 838
rect 138 836 140 838
rect 143 836 145 839
rect 164 836 166 839
rect 180 836 182 839
rect 196 836 198 838
rect 201 836 203 839
rect 217 836 219 838
rect 233 836 235 838
rect 238 836 240 839
rect 254 836 256 838
rect 270 836 272 838
rect 275 836 277 839
rect 296 836 298 839
rect 312 836 314 839
rect 328 836 330 838
rect 333 836 335 839
rect 349 836 351 838
rect 365 836 367 838
rect 370 836 372 839
rect 386 836 388 838
rect 402 836 404 838
rect 407 836 409 839
rect 428 836 430 839
rect 444 836 446 839
rect 460 836 462 838
rect 465 836 467 839
rect 481 836 483 838
rect 101 823 103 828
rect 106 826 108 828
rect 101 809 103 819
rect 106 809 108 816
rect 122 809 124 828
rect 138 819 140 828
rect 143 826 145 828
rect 164 826 166 828
rect 180 825 182 828
rect 138 809 140 812
rect 143 809 145 811
rect 164 809 166 811
rect 180 809 182 821
rect 196 819 198 828
rect 201 826 203 828
rect 196 809 198 812
rect 201 809 203 811
rect 217 809 219 828
rect 233 825 235 828
rect 238 826 240 828
rect 233 809 235 821
rect 238 809 240 816
rect 254 809 256 828
rect 270 819 272 828
rect 275 826 277 828
rect 296 826 298 828
rect 312 825 314 828
rect 270 809 272 812
rect 275 809 277 811
rect 296 809 298 811
rect 312 809 314 821
rect 328 819 330 828
rect 333 826 335 828
rect 328 809 330 812
rect 333 809 335 811
rect 349 809 351 828
rect 365 825 367 828
rect 370 826 372 828
rect 365 809 367 821
rect 370 809 372 816
rect 386 809 388 828
rect 402 819 404 828
rect 407 826 409 828
rect 428 826 430 828
rect 444 825 446 828
rect 402 809 404 812
rect 407 809 409 811
rect 428 809 430 811
rect 444 809 446 821
rect 460 819 462 828
rect 465 826 467 828
rect 481 820 483 828
rect 460 809 462 812
rect 465 809 467 811
rect 481 809 483 816
rect 101 803 103 805
rect 106 802 108 805
rect 122 803 124 805
rect 138 803 140 805
rect 143 800 145 805
rect 164 800 166 805
rect 180 803 182 805
rect 196 803 198 805
rect 201 800 203 805
rect 217 803 219 805
rect 233 803 235 805
rect 238 802 240 805
rect 254 803 256 805
rect 270 803 272 805
rect 275 800 277 805
rect 296 800 298 805
rect 312 803 314 805
rect 328 803 330 805
rect 333 800 335 805
rect 349 803 351 805
rect 365 803 367 805
rect 370 802 372 805
rect 386 803 388 805
rect 402 803 404 805
rect 407 800 409 805
rect 428 800 430 805
rect 444 803 446 805
rect 460 803 462 805
rect 465 800 467 805
rect 481 803 483 805
<< polycontact >>
rect 578 1740 582 1744
rect 615 1740 619 1744
rect 635 1740 639 1744
rect 673 1740 677 1744
rect 710 1740 714 1744
rect 747 1740 751 1744
rect 767 1740 771 1744
rect 805 1740 809 1744
rect 842 1740 846 1744
rect 879 1740 883 1744
rect 899 1740 903 1744
rect 937 1740 941 1744
rect 974 1740 978 1744
rect 1011 1740 1015 1744
rect 1031 1740 1035 1744
rect 1069 1740 1073 1744
rect 572 1720 576 1724
rect 590 1722 594 1726
rect 238 1707 242 1711
rect 275 1707 279 1711
rect 295 1707 299 1711
rect 333 1707 337 1711
rect 650 1722 654 1726
rect 608 1713 612 1720
rect 666 1713 670 1720
rect 687 1717 691 1721
rect 704 1720 708 1724
rect 722 1722 726 1726
rect 782 1722 786 1726
rect 740 1713 744 1720
rect 798 1713 802 1720
rect 819 1717 823 1721
rect 836 1720 840 1724
rect 854 1722 858 1726
rect 914 1722 918 1726
rect 872 1713 876 1720
rect 930 1713 934 1720
rect 951 1717 955 1721
rect 968 1720 972 1724
rect 986 1722 990 1726
rect 1046 1722 1050 1726
rect 1004 1713 1008 1720
rect 1062 1713 1066 1720
rect 1083 1717 1087 1721
rect 578 1699 582 1703
rect 615 1697 619 1701
rect 635 1697 639 1701
rect 671 1697 675 1701
rect 710 1699 714 1703
rect 747 1697 751 1701
rect 767 1697 771 1701
rect 803 1697 807 1701
rect 842 1699 846 1703
rect 879 1697 883 1701
rect 899 1697 903 1701
rect 935 1697 939 1701
rect 974 1699 978 1703
rect 1011 1697 1015 1701
rect 1031 1697 1035 1701
rect 1067 1697 1071 1701
rect 232 1687 236 1691
rect 250 1689 254 1693
rect 310 1689 314 1693
rect 268 1680 272 1687
rect 326 1680 330 1687
rect 345 1684 349 1688
rect 238 1666 242 1670
rect 275 1664 279 1668
rect 295 1664 299 1668
rect 331 1664 335 1668
rect 594 1656 598 1660
rect 638 1656 642 1660
rect 665 1656 669 1660
rect 710 1656 714 1660
rect 783 1663 787 1667
rect 356 1643 360 1647
rect 748 1649 752 1653
rect 239 1634 243 1638
rect 574 1636 578 1640
rect 606 1637 610 1641
rect 625 1636 629 1640
rect 681 1637 685 1641
rect 697 1636 701 1640
rect 724 1636 728 1640
rect 864 1663 868 1667
rect 775 1645 779 1649
rect 802 1641 806 1645
rect 829 1649 833 1653
rect 856 1645 860 1649
rect 883 1641 887 1645
rect 781 1627 785 1631
rect 862 1627 866 1631
rect 591 1619 595 1623
rect 635 1618 639 1622
rect 660 1619 665 1623
rect 707 1618 711 1622
rect 238 1605 242 1609
rect 276 1605 280 1609
rect 296 1605 300 1609
rect 333 1605 337 1609
rect 226 1582 230 1586
rect 261 1587 265 1591
rect 245 1578 249 1585
rect 303 1578 307 1585
rect 321 1587 325 1591
rect 591 1589 595 1593
rect 635 1590 639 1594
rect 339 1585 343 1589
rect 660 1589 665 1593
rect 707 1590 711 1594
rect 783 1587 787 1591
rect 864 1587 868 1591
rect 574 1572 578 1576
rect 240 1562 244 1566
rect 276 1562 280 1566
rect 296 1562 300 1566
rect 333 1564 337 1568
rect 606 1571 610 1575
rect 625 1572 629 1576
rect 681 1571 685 1575
rect 697 1572 701 1576
rect 724 1572 728 1576
rect 772 1571 778 1575
rect 853 1571 859 1575
rect 594 1552 598 1556
rect 638 1552 642 1556
rect 665 1552 669 1556
rect 710 1552 714 1556
rect 781 1551 785 1555
rect 862 1551 866 1555
rect 783 1531 787 1535
rect 594 1524 598 1528
rect 638 1524 642 1528
rect 665 1524 669 1528
rect 710 1524 714 1528
rect 888 1531 892 1535
rect 775 1513 779 1517
rect 574 1504 578 1508
rect 606 1505 610 1509
rect 625 1504 629 1508
rect 681 1505 685 1509
rect 697 1504 701 1508
rect 724 1504 728 1508
rect 802 1509 806 1513
rect 853 1517 857 1521
rect 880 1513 884 1517
rect 907 1509 911 1513
rect 781 1495 785 1499
rect 886 1495 890 1499
rect 591 1487 595 1491
rect 635 1486 639 1490
rect 660 1487 665 1491
rect 707 1486 711 1490
rect 591 1457 595 1461
rect 635 1458 639 1462
rect 660 1457 665 1461
rect 707 1458 711 1462
rect 783 1456 787 1460
rect 888 1456 892 1460
rect 574 1440 578 1444
rect 606 1439 610 1443
rect 625 1440 629 1444
rect 681 1439 685 1443
rect 697 1440 701 1444
rect 724 1440 728 1444
rect 772 1440 778 1444
rect 877 1440 883 1444
rect 594 1420 598 1424
rect 638 1420 642 1424
rect 665 1420 669 1424
rect 710 1420 714 1424
rect 781 1420 785 1424
rect 886 1420 890 1424
rect 783 1399 787 1403
rect 594 1392 598 1396
rect 638 1392 642 1396
rect 665 1392 669 1396
rect 710 1392 714 1396
rect 864 1399 868 1403
rect 775 1381 779 1385
rect 574 1372 578 1376
rect 606 1373 610 1377
rect 625 1372 629 1376
rect 681 1373 685 1377
rect 697 1372 701 1376
rect 724 1372 728 1376
rect 802 1377 806 1381
rect 829 1385 833 1389
rect 954 1399 958 1403
rect 856 1381 860 1385
rect 883 1377 887 1381
rect 919 1385 923 1389
rect 946 1381 950 1385
rect 973 1377 977 1381
rect 781 1363 785 1367
rect 862 1363 866 1367
rect 952 1363 956 1367
rect 591 1355 595 1359
rect 635 1354 639 1358
rect 660 1355 665 1359
rect 707 1354 711 1358
rect 591 1325 595 1329
rect 635 1326 639 1330
rect 660 1325 665 1329
rect 707 1326 711 1330
rect 783 1321 787 1325
rect 864 1321 868 1325
rect 954 1321 958 1325
rect 574 1308 578 1312
rect 606 1307 610 1311
rect 625 1308 629 1312
rect 681 1307 685 1311
rect 697 1308 701 1312
rect 724 1308 728 1312
rect 772 1305 778 1309
rect 853 1305 859 1309
rect 943 1305 949 1309
rect 594 1288 598 1292
rect 638 1288 642 1292
rect 665 1288 669 1292
rect 710 1288 714 1292
rect 781 1285 785 1289
rect 862 1285 866 1289
rect 952 1285 956 1289
rect 783 1267 787 1271
rect 594 1260 598 1264
rect 638 1260 642 1264
rect 665 1260 669 1264
rect 710 1260 714 1264
rect 775 1249 779 1253
rect 574 1240 578 1244
rect 606 1241 610 1245
rect 625 1240 629 1244
rect 681 1241 685 1245
rect 697 1240 701 1244
rect 724 1240 728 1244
rect 802 1245 806 1249
rect 781 1231 785 1235
rect 591 1223 595 1227
rect 635 1222 639 1226
rect 660 1223 665 1227
rect 707 1222 711 1226
rect 106 1205 110 1209
rect 143 1205 147 1209
rect 163 1205 167 1209
rect 201 1205 205 1209
rect 238 1205 242 1209
rect 275 1205 279 1209
rect 295 1205 299 1209
rect 333 1205 337 1209
rect 370 1205 374 1209
rect 407 1205 411 1209
rect 427 1205 431 1209
rect 465 1205 469 1209
rect 100 1185 104 1189
rect 118 1187 122 1191
rect 178 1187 182 1191
rect 136 1178 140 1185
rect 194 1178 198 1185
rect 213 1182 217 1186
rect 231 1187 235 1191
rect 250 1187 254 1191
rect 310 1187 314 1191
rect 268 1178 272 1185
rect 326 1178 330 1185
rect 345 1182 349 1186
rect 363 1187 367 1191
rect 382 1187 386 1191
rect 442 1187 446 1191
rect 400 1178 404 1185
rect 591 1193 595 1197
rect 635 1194 639 1198
rect 660 1193 665 1197
rect 707 1194 711 1198
rect 852 1193 856 1197
rect 896 1194 900 1198
rect 921 1193 926 1197
rect 968 1194 972 1198
rect 458 1178 462 1185
rect 479 1182 483 1186
rect 783 1185 787 1189
rect 574 1176 578 1180
rect 606 1175 610 1179
rect 625 1176 629 1180
rect 681 1175 685 1179
rect 697 1176 701 1180
rect 724 1176 728 1180
rect 106 1164 110 1168
rect 143 1162 147 1166
rect 163 1162 167 1166
rect 199 1162 203 1166
rect 238 1164 242 1168
rect 275 1162 279 1166
rect 295 1162 299 1166
rect 331 1162 335 1166
rect 370 1164 374 1168
rect 407 1162 411 1166
rect 427 1162 431 1166
rect 463 1162 467 1166
rect 772 1169 778 1173
rect 810 1176 814 1180
rect 867 1175 871 1179
rect 886 1176 890 1180
rect 942 1175 946 1179
rect 958 1176 962 1180
rect 985 1176 989 1180
rect 594 1156 598 1160
rect 638 1156 642 1160
rect 665 1156 669 1160
rect 710 1156 714 1160
rect 855 1156 859 1160
rect 899 1156 903 1160
rect 926 1156 930 1160
rect 971 1156 975 1160
rect 781 1149 785 1153
rect 215 1134 219 1138
rect 239 1134 243 1138
rect 994 1128 998 1132
rect 235 1109 239 1113
rect 250 1101 254 1105
rect 877 1095 881 1099
rect 914 1095 918 1099
rect 934 1095 938 1099
rect 972 1095 976 1099
rect 215 1086 219 1090
rect 239 1086 243 1090
rect 871 1075 875 1079
rect 889 1077 893 1081
rect 106 1065 110 1069
rect 143 1065 147 1069
rect 163 1065 167 1069
rect 201 1065 205 1069
rect 238 1065 242 1069
rect 275 1065 279 1069
rect 295 1065 299 1069
rect 333 1065 337 1069
rect 370 1065 374 1069
rect 407 1065 411 1069
rect 427 1065 431 1069
rect 465 1065 469 1069
rect 949 1077 953 1081
rect 907 1068 911 1075
rect 965 1068 969 1075
rect 984 1072 988 1076
rect 877 1054 881 1058
rect 100 1045 104 1049
rect 118 1047 122 1051
rect 178 1047 182 1051
rect 136 1038 140 1045
rect 194 1038 198 1045
rect 213 1042 217 1046
rect 231 1047 235 1051
rect 250 1047 254 1051
rect 310 1047 314 1051
rect 268 1038 272 1045
rect 326 1038 330 1045
rect 345 1042 349 1046
rect 363 1047 367 1051
rect 382 1047 386 1051
rect 442 1047 446 1051
rect 400 1038 404 1045
rect 914 1052 918 1056
rect 934 1052 938 1056
rect 970 1052 974 1056
rect 458 1038 462 1045
rect 479 1042 483 1046
rect 106 1024 110 1028
rect 143 1022 147 1026
rect 163 1022 167 1026
rect 199 1022 203 1026
rect 238 1024 242 1028
rect 275 1022 279 1026
rect 295 1022 299 1026
rect 331 1022 335 1026
rect 370 1024 374 1028
rect 407 1022 411 1026
rect 427 1022 431 1026
rect 463 1022 467 1026
rect 877 1009 881 1013
rect 914 1009 918 1013
rect 934 1009 938 1013
rect 972 1009 976 1013
rect 871 989 875 993
rect 889 991 893 995
rect 106 979 110 983
rect 143 979 147 983
rect 163 979 167 983
rect 201 979 205 983
rect 238 979 242 983
rect 275 979 279 983
rect 295 979 299 983
rect 333 979 337 983
rect 370 979 374 983
rect 407 979 411 983
rect 427 979 431 983
rect 465 979 469 983
rect 949 991 953 995
rect 907 982 911 989
rect 965 982 969 989
rect 984 986 988 990
rect 1006 984 1010 988
rect 877 968 881 972
rect 100 959 104 963
rect 118 961 122 965
rect 178 961 182 965
rect 136 952 140 959
rect 194 952 198 959
rect 213 956 217 960
rect 231 961 235 965
rect 250 961 254 965
rect 310 961 314 965
rect 268 952 272 959
rect 326 952 330 959
rect 345 956 349 960
rect 363 961 367 965
rect 382 961 386 965
rect 442 961 446 965
rect 400 952 404 959
rect 914 966 918 970
rect 934 966 938 970
rect 970 966 974 970
rect 458 952 462 959
rect 479 956 483 960
rect 106 938 110 942
rect 143 936 147 940
rect 163 936 167 940
rect 199 936 203 940
rect 238 938 242 942
rect 275 936 279 940
rect 295 936 299 940
rect 331 936 335 940
rect 370 938 374 942
rect 407 936 411 940
rect 427 936 431 940
rect 463 936 467 940
rect 332 908 336 912
rect 356 908 360 912
rect 352 883 356 887
rect 367 875 371 879
rect 332 860 336 864
rect 356 860 360 864
rect 106 839 110 843
rect 143 839 147 843
rect 163 839 167 843
rect 201 839 205 843
rect 238 839 242 843
rect 275 839 279 843
rect 295 839 299 843
rect 333 839 337 843
rect 370 839 374 843
rect 407 839 411 843
rect 427 839 431 843
rect 465 839 469 843
rect 100 819 104 823
rect 118 821 122 825
rect 178 821 182 825
rect 136 812 140 819
rect 194 812 198 819
rect 213 816 217 820
rect 231 821 235 825
rect 250 821 254 825
rect 310 821 314 825
rect 268 812 272 819
rect 326 812 330 819
rect 345 816 349 820
rect 363 821 367 825
rect 382 821 386 825
rect 442 821 446 825
rect 400 812 404 819
rect 458 812 462 819
rect 479 816 483 820
rect 106 798 110 802
rect 143 796 147 800
rect 163 796 167 800
rect 199 796 203 800
rect 238 798 242 802
rect 275 796 279 800
rect 295 796 299 800
rect 331 796 335 800
rect 370 798 374 802
rect 407 796 411 800
rect 427 796 431 800
rect 463 796 467 800
<< metal1 >>
rect 559 1754 574 1758
rect 578 1754 610 1758
rect 614 1754 677 1758
rect 681 1754 706 1758
rect 710 1754 742 1758
rect 746 1754 809 1758
rect 813 1754 838 1758
rect 842 1754 874 1758
rect 878 1754 941 1758
rect 945 1754 970 1758
rect 974 1754 1006 1758
rect 1010 1754 1073 1758
rect 1077 1754 1093 1758
rect 499 1747 598 1751
rect 602 1747 626 1751
rect 630 1747 656 1751
rect 660 1747 693 1751
rect 697 1747 730 1751
rect 734 1747 758 1751
rect 762 1747 788 1751
rect 792 1747 825 1751
rect 829 1747 862 1751
rect 866 1747 890 1751
rect 894 1747 920 1751
rect 924 1747 957 1751
rect 961 1747 994 1751
rect 998 1747 1022 1751
rect 1026 1747 1052 1751
rect 1056 1747 1089 1751
rect 568 1737 571 1747
rect 589 1737 592 1747
rect 605 1737 608 1747
rect 619 1740 624 1744
rect 628 1740 635 1744
rect 647 1737 650 1747
rect 663 1737 666 1747
rect 684 1737 687 1747
rect 700 1737 703 1747
rect 721 1737 724 1747
rect 737 1737 740 1747
rect 751 1740 756 1744
rect 760 1740 767 1744
rect 779 1737 782 1747
rect 795 1737 798 1747
rect 816 1737 819 1747
rect 832 1737 835 1747
rect 853 1737 856 1747
rect 869 1737 872 1747
rect 883 1740 888 1744
rect 892 1740 899 1744
rect 911 1737 914 1747
rect 927 1737 930 1747
rect 948 1737 951 1747
rect 964 1737 967 1747
rect 985 1737 988 1747
rect 1001 1737 1004 1747
rect 1015 1740 1020 1744
rect 1024 1740 1031 1744
rect 1043 1737 1046 1747
rect 1059 1737 1062 1747
rect 1080 1737 1083 1747
rect 225 1721 234 1725
rect 238 1721 270 1725
rect 274 1721 337 1725
rect 341 1721 553 1725
rect 585 1723 590 1726
rect 594 1723 618 1726
rect 643 1723 650 1726
rect 654 1723 676 1726
rect 225 1714 258 1718
rect 262 1714 286 1718
rect 290 1714 316 1718
rect 320 1714 353 1718
rect 357 1714 493 1718
rect 228 1704 231 1714
rect 249 1704 252 1714
rect 265 1704 268 1714
rect 279 1707 284 1711
rect 288 1707 295 1711
rect 307 1704 310 1714
rect 323 1704 326 1714
rect 344 1704 347 1714
rect 601 1713 608 1716
rect 612 1717 631 1720
rect 631 1710 634 1716
rect 659 1713 666 1716
rect 670 1717 687 1720
rect 717 1723 722 1726
rect 726 1723 750 1726
rect 775 1723 782 1726
rect 786 1723 808 1726
rect 733 1713 740 1716
rect 744 1717 763 1720
rect 763 1710 766 1716
rect 791 1713 798 1716
rect 802 1717 819 1720
rect 849 1723 854 1726
rect 858 1723 882 1726
rect 907 1723 914 1726
rect 918 1723 940 1726
rect 865 1713 872 1716
rect 876 1717 895 1720
rect 895 1710 898 1716
rect 923 1713 930 1716
rect 934 1717 951 1720
rect 981 1723 986 1726
rect 990 1723 1014 1726
rect 1039 1723 1046 1726
rect 1050 1723 1072 1726
rect 997 1713 1004 1716
rect 1008 1717 1027 1720
rect 223 1687 232 1691
rect 245 1690 250 1693
rect 254 1690 278 1693
rect 303 1690 310 1693
rect 314 1690 336 1693
rect 568 1694 571 1706
rect 589 1694 592 1706
rect 605 1694 608 1706
rect 619 1697 631 1700
rect 647 1694 650 1706
rect 663 1694 666 1706
rect 684 1694 687 1706
rect 700 1694 703 1706
rect 721 1694 724 1706
rect 737 1694 740 1706
rect 751 1697 763 1700
rect 779 1694 782 1706
rect 795 1694 798 1706
rect 816 1694 819 1706
rect 832 1694 835 1706
rect 853 1694 856 1706
rect 869 1694 872 1706
rect 883 1697 895 1700
rect 911 1694 914 1706
rect 927 1694 930 1706
rect 948 1694 951 1706
rect 1027 1710 1030 1716
rect 1055 1713 1062 1716
rect 1066 1717 1083 1720
rect 964 1694 967 1706
rect 985 1694 988 1706
rect 1001 1694 1004 1706
rect 1015 1697 1027 1700
rect 1043 1694 1046 1706
rect 1059 1694 1062 1706
rect 1080 1694 1083 1706
rect 511 1690 598 1694
rect 602 1690 626 1694
rect 630 1690 656 1694
rect 660 1690 730 1694
rect 734 1690 758 1694
rect 762 1690 788 1694
rect 792 1690 862 1694
rect 866 1690 890 1694
rect 894 1690 920 1694
rect 924 1690 994 1694
rect 998 1690 1022 1694
rect 1026 1690 1052 1694
rect 1056 1690 1093 1694
rect 261 1680 268 1683
rect 272 1684 291 1687
rect 291 1677 294 1683
rect 319 1680 326 1683
rect 330 1684 345 1687
rect 547 1683 574 1687
rect 578 1683 625 1687
rect 629 1683 675 1687
rect 679 1683 706 1687
rect 710 1683 757 1687
rect 761 1683 807 1687
rect 811 1683 838 1687
rect 842 1683 889 1687
rect 893 1683 939 1687
rect 943 1683 970 1687
rect 974 1683 1021 1687
rect 1025 1683 1071 1687
rect 1075 1683 1093 1687
rect 228 1661 231 1673
rect 249 1661 252 1673
rect 265 1661 268 1673
rect 279 1664 291 1667
rect 307 1661 310 1673
rect 323 1661 326 1673
rect 344 1661 347 1673
rect 499 1670 572 1674
rect 576 1670 588 1674
rect 592 1670 606 1674
rect 610 1670 617 1674
rect 621 1670 623 1674
rect 627 1670 642 1674
rect 646 1670 679 1674
rect 683 1670 684 1674
rect 688 1670 696 1674
rect 700 1670 724 1674
rect 728 1670 740 1674
rect 744 1670 764 1674
rect 768 1670 818 1674
rect 822 1670 845 1674
rect 849 1670 899 1674
rect 903 1670 922 1674
rect 535 1663 599 1667
rect 603 1663 630 1667
rect 634 1663 652 1667
rect 656 1663 717 1667
rect 721 1663 735 1667
rect 747 1666 750 1670
rect 225 1657 258 1661
rect 262 1657 286 1661
rect 290 1657 316 1661
rect 320 1657 505 1661
rect 225 1650 234 1654
rect 238 1650 285 1654
rect 289 1650 335 1654
rect 339 1650 541 1654
rect 642 1656 645 1660
rect 669 1656 670 1660
rect 714 1656 716 1660
rect 756 1653 759 1658
rect 771 1660 774 1670
rect 801 1666 804 1670
rect 828 1666 831 1670
rect 223 1634 239 1638
rect 348 1636 352 1640
rect 364 1636 368 1640
rect 372 1636 574 1640
rect 582 1639 585 1645
rect 589 1639 592 1645
rect 582 1636 592 1639
rect 582 1631 585 1636
rect 231 1627 235 1631
rect 247 1627 368 1631
rect 589 1631 592 1636
rect 598 1641 601 1645
rect 598 1637 600 1641
rect 604 1637 606 1641
rect 614 1640 617 1645
rect 642 1642 645 1645
rect 614 1638 625 1640
rect 598 1631 601 1637
rect 614 1636 620 1638
rect 614 1631 617 1636
rect 624 1636 625 1638
rect 643 1638 645 1642
rect 642 1631 645 1638
rect 745 1649 748 1652
rect 787 1649 790 1652
rect 658 1641 661 1645
rect 668 1641 671 1645
rect 668 1637 677 1641
rect 689 1640 692 1645
rect 714 1641 717 1645
rect 658 1631 661 1637
rect 668 1631 671 1637
rect 689 1636 690 1640
rect 694 1636 697 1639
rect 716 1637 717 1641
rect 732 1640 735 1645
rect 756 1644 759 1649
rect 764 1645 775 1648
rect 787 1646 795 1649
rect 689 1631 692 1636
rect 714 1631 717 1637
rect 732 1631 735 1636
rect 218 1619 234 1623
rect 238 1619 301 1623
rect 305 1619 337 1623
rect 341 1619 553 1623
rect 634 1618 635 1622
rect 659 1619 660 1623
rect 706 1618 707 1622
rect 222 1612 255 1616
rect 259 1612 285 1616
rect 289 1612 313 1616
rect 317 1612 493 1616
rect 228 1602 231 1612
rect 249 1602 252 1612
rect 265 1602 268 1612
rect 280 1605 287 1609
rect 291 1605 296 1609
rect 307 1602 310 1612
rect 323 1602 326 1612
rect 344 1602 347 1612
rect 523 1611 587 1615
rect 591 1611 646 1615
rect 650 1611 671 1615
rect 675 1611 702 1615
rect 706 1611 735 1615
rect 747 1608 750 1640
rect 764 1639 767 1645
rect 787 1640 790 1646
rect 799 1641 802 1644
rect 810 1644 813 1658
rect 837 1653 840 1658
rect 852 1660 855 1670
rect 882 1666 885 1670
rect 821 1649 822 1652
rect 826 1649 829 1652
rect 868 1649 871 1652
rect 810 1641 818 1644
rect 837 1644 840 1649
rect 810 1636 813 1641
rect 818 1637 822 1641
rect 845 1645 856 1648
rect 868 1646 876 1649
rect 762 1630 767 1635
rect 771 1608 774 1636
rect 801 1608 804 1632
rect 828 1608 831 1640
rect 845 1639 848 1645
rect 868 1640 871 1646
rect 880 1641 883 1644
rect 891 1644 894 1658
rect 891 1641 903 1644
rect 891 1636 894 1641
rect 843 1630 848 1635
rect 852 1608 855 1636
rect 882 1608 885 1632
rect 511 1604 573 1608
rect 577 1604 579 1608
rect 583 1604 587 1608
rect 591 1604 605 1608
rect 609 1604 614 1608
rect 618 1604 623 1608
rect 627 1604 646 1608
rect 650 1604 680 1608
rect 684 1604 695 1608
rect 699 1604 723 1608
rect 727 1604 740 1608
rect 744 1604 764 1608
rect 768 1604 818 1608
rect 825 1604 845 1608
rect 849 1604 899 1608
rect 239 1588 261 1591
rect 265 1588 272 1591
rect 523 1597 587 1601
rect 591 1597 646 1601
rect 650 1597 671 1601
rect 675 1597 702 1601
rect 706 1597 735 1601
rect 297 1588 321 1591
rect 325 1588 330 1591
rect 634 1590 635 1594
rect 659 1589 660 1593
rect 706 1590 707 1594
rect 343 1585 352 1589
rect 230 1582 245 1585
rect 284 1582 303 1585
rect 249 1578 256 1581
rect 281 1575 284 1581
rect 307 1578 314 1581
rect 582 1576 585 1581
rect 589 1576 592 1581
rect 572 1573 574 1576
rect 582 1573 592 1576
rect 228 1559 231 1571
rect 249 1559 252 1571
rect 265 1559 268 1571
rect 284 1562 296 1565
rect 307 1559 310 1571
rect 323 1559 326 1571
rect 344 1559 347 1571
rect 582 1567 585 1573
rect 589 1567 592 1573
rect 598 1575 601 1581
rect 614 1576 617 1581
rect 598 1571 600 1575
rect 604 1571 606 1575
rect 614 1574 620 1576
rect 624 1574 625 1576
rect 614 1572 625 1574
rect 642 1574 645 1581
rect 598 1567 601 1571
rect 614 1567 617 1572
rect 643 1570 645 1574
rect 642 1567 645 1570
rect 658 1575 661 1581
rect 668 1575 671 1581
rect 689 1576 692 1581
rect 668 1571 677 1575
rect 689 1572 690 1576
rect 694 1573 697 1576
rect 714 1575 717 1581
rect 732 1576 735 1581
rect 771 1584 774 1604
rect 852 1584 855 1604
rect 658 1567 661 1571
rect 668 1567 671 1571
rect 689 1567 692 1572
rect 716 1571 717 1575
rect 714 1567 717 1571
rect 732 1567 735 1572
rect 762 1571 767 1576
rect 771 1572 772 1575
rect 787 1574 790 1580
rect 787 1571 795 1574
rect 842 1571 847 1576
rect 851 1572 853 1575
rect 868 1574 871 1580
rect 868 1571 876 1574
rect 787 1568 790 1571
rect 868 1568 871 1571
rect 218 1555 255 1559
rect 259 1555 285 1559
rect 289 1555 313 1559
rect 317 1555 505 1559
rect 642 1552 645 1556
rect 669 1552 670 1556
rect 714 1552 716 1556
rect 218 1548 236 1552
rect 240 1548 286 1552
rect 290 1548 337 1552
rect 341 1548 541 1552
rect 587 1545 599 1549
rect 603 1545 630 1549
rect 634 1545 652 1549
rect 656 1545 717 1549
rect 721 1545 735 1549
rect 771 1542 774 1560
rect 852 1542 855 1560
rect 499 1538 572 1542
rect 576 1538 588 1542
rect 592 1538 606 1542
rect 610 1538 617 1542
rect 621 1538 623 1542
rect 627 1538 642 1542
rect 646 1538 679 1542
rect 683 1538 684 1542
rect 688 1538 696 1542
rect 700 1538 724 1542
rect 728 1538 740 1542
rect 744 1538 764 1542
rect 768 1538 818 1542
rect 822 1538 845 1542
rect 849 1538 907 1542
rect 911 1538 922 1542
rect 535 1531 583 1535
rect 587 1531 599 1535
rect 603 1531 630 1535
rect 634 1531 652 1535
rect 656 1531 717 1535
rect 721 1531 735 1535
rect 771 1528 774 1538
rect 801 1534 804 1538
rect 852 1534 855 1538
rect 642 1524 645 1528
rect 669 1524 670 1528
rect 714 1524 716 1528
rect 571 1504 574 1507
rect 582 1507 585 1513
rect 589 1507 592 1513
rect 582 1504 592 1507
rect 582 1499 585 1504
rect 589 1499 592 1504
rect 598 1509 601 1513
rect 598 1505 600 1509
rect 604 1505 606 1509
rect 614 1508 617 1513
rect 642 1510 645 1513
rect 614 1506 625 1508
rect 598 1499 601 1505
rect 614 1504 620 1506
rect 614 1499 617 1504
rect 624 1504 625 1506
rect 643 1506 645 1510
rect 642 1499 645 1506
rect 787 1517 790 1520
rect 658 1509 661 1513
rect 668 1509 671 1513
rect 668 1505 677 1509
rect 689 1508 692 1513
rect 714 1509 717 1513
rect 658 1499 661 1505
rect 668 1499 671 1505
rect 689 1504 690 1508
rect 694 1504 697 1507
rect 716 1505 717 1509
rect 732 1508 735 1513
rect 764 1513 775 1516
rect 787 1514 795 1517
rect 689 1499 692 1504
rect 714 1499 717 1505
rect 764 1507 767 1513
rect 787 1508 790 1514
rect 799 1509 802 1512
rect 810 1512 813 1526
rect 861 1521 864 1526
rect 876 1528 879 1538
rect 906 1534 909 1538
rect 845 1517 846 1520
rect 850 1517 853 1520
rect 892 1517 895 1520
rect 818 1512 823 1517
rect 861 1512 864 1517
rect 810 1509 818 1512
rect 732 1499 735 1504
rect 810 1504 813 1509
rect 869 1513 880 1516
rect 892 1514 900 1517
rect 762 1498 767 1503
rect 634 1486 635 1490
rect 659 1487 660 1491
rect 706 1486 707 1490
rect 523 1479 587 1483
rect 591 1479 646 1483
rect 650 1479 671 1483
rect 675 1479 702 1483
rect 706 1479 735 1483
rect 771 1476 774 1504
rect 801 1476 804 1500
rect 852 1476 855 1508
rect 869 1507 872 1513
rect 892 1508 895 1514
rect 904 1509 907 1512
rect 915 1512 918 1526
rect 915 1509 921 1512
rect 915 1504 918 1509
rect 867 1498 872 1503
rect 876 1476 879 1504
rect 906 1476 909 1500
rect 511 1472 573 1476
rect 577 1472 579 1476
rect 583 1472 587 1476
rect 591 1472 605 1476
rect 609 1472 614 1476
rect 618 1472 623 1476
rect 627 1472 646 1476
rect 650 1472 680 1476
rect 684 1472 695 1476
rect 699 1472 723 1476
rect 727 1472 740 1476
rect 744 1472 764 1476
rect 768 1472 818 1476
rect 822 1472 845 1476
rect 849 1472 869 1476
rect 873 1472 921 1476
rect 523 1465 587 1469
rect 591 1465 646 1469
rect 650 1465 671 1469
rect 675 1465 702 1469
rect 706 1465 735 1469
rect 634 1458 635 1462
rect 659 1457 660 1461
rect 706 1458 707 1462
rect 771 1453 774 1472
rect 876 1453 879 1472
rect 582 1444 585 1449
rect 589 1444 592 1449
rect 572 1441 574 1444
rect 582 1441 592 1444
rect 582 1435 585 1441
rect 589 1435 592 1441
rect 598 1443 601 1449
rect 614 1444 617 1449
rect 598 1439 600 1443
rect 604 1439 606 1443
rect 614 1442 620 1444
rect 624 1442 625 1444
rect 614 1440 625 1442
rect 642 1442 645 1449
rect 598 1435 601 1439
rect 614 1435 617 1440
rect 643 1438 645 1442
rect 642 1435 645 1438
rect 658 1443 661 1449
rect 668 1443 671 1449
rect 689 1444 692 1449
rect 668 1439 677 1443
rect 689 1440 690 1444
rect 694 1441 697 1444
rect 714 1443 717 1449
rect 732 1444 735 1449
rect 658 1435 661 1439
rect 668 1435 671 1439
rect 689 1435 692 1440
rect 716 1439 717 1443
rect 761 1440 766 1445
rect 770 1441 772 1444
rect 787 1443 790 1449
rect 787 1440 795 1443
rect 867 1440 872 1445
rect 876 1441 877 1444
rect 892 1443 895 1449
rect 892 1440 900 1443
rect 714 1435 717 1439
rect 732 1435 735 1440
rect 787 1437 790 1440
rect 892 1437 895 1440
rect 642 1420 645 1424
rect 669 1420 670 1424
rect 714 1420 716 1424
rect 535 1413 599 1417
rect 603 1413 630 1417
rect 634 1413 652 1417
rect 656 1413 717 1417
rect 721 1413 735 1417
rect 771 1410 774 1429
rect 876 1410 879 1429
rect 499 1406 572 1410
rect 576 1406 588 1410
rect 592 1406 606 1410
rect 610 1406 617 1410
rect 621 1406 623 1410
rect 627 1406 642 1410
rect 646 1406 679 1410
rect 683 1406 684 1410
rect 688 1406 696 1410
rect 700 1406 724 1410
rect 728 1406 740 1410
rect 744 1406 764 1410
rect 768 1406 818 1410
rect 822 1406 845 1410
rect 849 1406 899 1410
rect 903 1406 907 1410
rect 911 1406 935 1410
rect 939 1406 989 1410
rect 535 1399 599 1403
rect 603 1399 630 1403
rect 634 1399 652 1403
rect 656 1399 717 1403
rect 721 1399 735 1403
rect 771 1396 774 1406
rect 801 1402 804 1406
rect 828 1402 831 1406
rect 642 1392 645 1396
rect 669 1392 670 1396
rect 714 1392 716 1396
rect 571 1372 574 1375
rect 582 1375 585 1381
rect 589 1375 592 1381
rect 582 1372 592 1375
rect 582 1367 585 1372
rect 589 1367 592 1372
rect 598 1377 601 1381
rect 598 1373 600 1377
rect 604 1373 606 1377
rect 614 1376 617 1381
rect 642 1378 645 1381
rect 614 1374 625 1376
rect 598 1367 601 1373
rect 614 1372 620 1374
rect 614 1367 617 1372
rect 624 1372 625 1374
rect 643 1374 645 1378
rect 642 1367 645 1374
rect 787 1385 790 1388
rect 658 1377 661 1381
rect 668 1377 671 1381
rect 668 1373 677 1377
rect 689 1376 692 1381
rect 714 1377 717 1381
rect 658 1367 661 1373
rect 668 1367 671 1373
rect 689 1372 690 1376
rect 694 1372 697 1375
rect 716 1373 717 1377
rect 732 1376 735 1381
rect 764 1381 775 1384
rect 787 1382 795 1385
rect 689 1367 692 1372
rect 714 1367 717 1373
rect 764 1375 767 1381
rect 787 1376 790 1382
rect 799 1377 802 1380
rect 810 1380 813 1394
rect 837 1389 840 1394
rect 852 1396 855 1406
rect 882 1402 885 1406
rect 918 1402 921 1406
rect 821 1385 822 1388
rect 826 1385 829 1388
rect 868 1385 871 1388
rect 810 1377 818 1380
rect 837 1380 840 1385
rect 732 1367 735 1372
rect 810 1372 813 1377
rect 818 1373 822 1377
rect 845 1381 856 1384
rect 868 1382 876 1385
rect 762 1366 767 1371
rect 634 1354 635 1358
rect 659 1355 660 1359
rect 706 1354 707 1358
rect 523 1347 587 1351
rect 591 1347 646 1351
rect 650 1347 671 1351
rect 675 1347 702 1351
rect 706 1347 735 1351
rect 771 1344 774 1372
rect 801 1344 804 1368
rect 828 1344 831 1376
rect 845 1375 848 1381
rect 868 1376 871 1382
rect 880 1377 883 1380
rect 891 1380 894 1394
rect 927 1389 930 1394
rect 942 1396 945 1406
rect 972 1402 975 1406
rect 916 1385 919 1388
rect 958 1385 961 1388
rect 891 1377 900 1380
rect 927 1380 930 1385
rect 891 1372 894 1377
rect 843 1366 848 1371
rect 852 1344 855 1372
rect 934 1383 946 1384
rect 938 1381 946 1383
rect 958 1382 966 1385
rect 958 1376 961 1382
rect 970 1377 973 1380
rect 981 1380 984 1394
rect 981 1377 1001 1380
rect 882 1344 885 1368
rect 918 1344 921 1376
rect 981 1372 984 1377
rect 942 1344 945 1372
rect 972 1344 975 1368
rect 511 1340 573 1344
rect 577 1340 579 1344
rect 583 1340 587 1344
rect 591 1340 605 1344
rect 609 1340 614 1344
rect 618 1340 623 1344
rect 627 1340 646 1344
rect 650 1340 680 1344
rect 684 1340 695 1344
rect 699 1340 723 1344
rect 727 1340 740 1344
rect 744 1340 764 1344
rect 768 1340 818 1344
rect 825 1340 845 1344
rect 849 1340 899 1344
rect 903 1340 935 1344
rect 939 1340 989 1344
rect 523 1333 587 1337
rect 591 1333 646 1337
rect 650 1333 671 1337
rect 675 1333 702 1337
rect 706 1333 735 1337
rect 634 1326 635 1330
rect 659 1325 660 1329
rect 706 1326 707 1330
rect 582 1312 585 1317
rect 589 1312 592 1317
rect 572 1309 574 1312
rect 582 1309 592 1312
rect 582 1303 585 1309
rect 589 1303 592 1309
rect 598 1311 601 1317
rect 614 1312 617 1317
rect 598 1307 600 1311
rect 604 1307 606 1311
rect 614 1310 620 1312
rect 624 1310 625 1312
rect 614 1308 625 1310
rect 642 1310 645 1317
rect 598 1303 601 1307
rect 614 1303 617 1308
rect 643 1306 645 1310
rect 642 1303 645 1306
rect 658 1311 661 1317
rect 668 1311 671 1317
rect 689 1312 692 1317
rect 668 1307 677 1311
rect 689 1308 690 1312
rect 694 1309 697 1312
rect 714 1311 717 1317
rect 732 1312 735 1317
rect 771 1318 774 1340
rect 852 1318 855 1340
rect 942 1318 945 1340
rect 658 1303 661 1307
rect 668 1303 671 1307
rect 689 1303 692 1308
rect 716 1307 717 1311
rect 714 1303 717 1307
rect 732 1303 735 1308
rect 762 1305 767 1310
rect 771 1306 772 1309
rect 787 1308 790 1314
rect 787 1305 795 1308
rect 842 1305 847 1310
rect 851 1306 853 1309
rect 868 1308 871 1314
rect 868 1305 876 1308
rect 935 1306 943 1309
rect 958 1308 961 1314
rect 958 1305 966 1308
rect 787 1302 790 1305
rect 868 1302 871 1305
rect 958 1302 961 1305
rect 642 1288 645 1292
rect 669 1288 670 1292
rect 714 1288 716 1292
rect 535 1281 599 1285
rect 603 1281 630 1285
rect 634 1281 652 1285
rect 656 1281 717 1285
rect 721 1281 735 1285
rect 771 1278 774 1294
rect 852 1278 855 1294
rect 942 1278 945 1294
rect 499 1274 572 1278
rect 576 1274 588 1278
rect 592 1274 606 1278
rect 610 1274 617 1278
rect 621 1274 623 1278
rect 627 1274 642 1278
rect 646 1274 679 1278
rect 683 1274 684 1278
rect 688 1274 696 1278
rect 700 1274 724 1278
rect 728 1274 740 1278
rect 744 1274 764 1278
rect 768 1274 818 1278
rect 822 1274 845 1278
rect 849 1274 935 1278
rect 939 1274 993 1278
rect 535 1267 599 1271
rect 603 1267 630 1271
rect 634 1267 652 1271
rect 656 1267 717 1271
rect 721 1267 735 1271
rect 771 1264 774 1274
rect 801 1270 804 1274
rect 642 1260 645 1264
rect 669 1260 670 1264
rect 714 1260 716 1264
rect 571 1240 574 1243
rect 582 1243 585 1249
rect 589 1243 592 1249
rect 582 1240 592 1243
rect 582 1235 585 1240
rect 589 1235 592 1240
rect 598 1245 601 1249
rect 598 1241 600 1245
rect 604 1241 606 1245
rect 614 1244 617 1249
rect 642 1246 645 1249
rect 614 1242 625 1244
rect 598 1235 601 1241
rect 614 1240 620 1242
rect 614 1235 617 1240
rect 624 1240 625 1242
rect 643 1242 645 1246
rect 642 1235 645 1242
rect 787 1253 790 1256
rect 658 1245 661 1249
rect 668 1245 671 1249
rect 668 1241 677 1245
rect 689 1244 692 1249
rect 714 1245 717 1249
rect 658 1235 661 1241
rect 668 1235 671 1241
rect 689 1240 690 1244
rect 694 1240 697 1243
rect 716 1241 717 1245
rect 732 1244 735 1249
rect 764 1249 775 1252
rect 787 1250 795 1253
rect 689 1235 692 1240
rect 714 1235 717 1241
rect 764 1243 767 1249
rect 787 1244 790 1250
rect 799 1245 802 1248
rect 810 1248 813 1262
rect 818 1248 823 1253
rect 810 1245 818 1248
rect 732 1235 735 1240
rect 810 1240 813 1245
rect 762 1234 767 1239
rect 93 1219 102 1223
rect 106 1219 138 1223
rect 142 1219 205 1223
rect 209 1219 234 1223
rect 238 1219 270 1223
rect 274 1219 337 1223
rect 341 1219 366 1223
rect 370 1219 402 1223
rect 406 1219 469 1223
rect 473 1219 553 1223
rect 634 1222 635 1226
rect 659 1223 660 1227
rect 706 1222 707 1226
rect 93 1212 126 1216
rect 130 1212 154 1216
rect 158 1212 184 1216
rect 188 1212 221 1216
rect 225 1212 258 1216
rect 262 1212 286 1216
rect 290 1212 316 1216
rect 320 1212 353 1216
rect 357 1212 390 1216
rect 394 1212 418 1216
rect 422 1212 448 1216
rect 452 1212 485 1216
rect 489 1212 493 1216
rect 566 1215 587 1219
rect 591 1215 596 1219
rect 600 1215 646 1219
rect 650 1215 671 1219
rect 675 1215 702 1219
rect 706 1215 735 1219
rect 771 1212 774 1240
rect 801 1212 804 1236
rect 96 1202 99 1212
rect 117 1202 120 1212
rect 133 1202 136 1212
rect 147 1205 152 1209
rect 156 1205 163 1209
rect 175 1202 178 1212
rect 191 1202 194 1212
rect 212 1202 215 1212
rect 228 1202 231 1212
rect 249 1202 252 1212
rect 265 1202 268 1212
rect 279 1205 284 1209
rect 288 1205 295 1209
rect 307 1202 310 1212
rect 323 1202 326 1212
rect 344 1202 347 1212
rect 360 1202 363 1212
rect 381 1202 384 1212
rect 397 1202 400 1212
rect 411 1205 416 1209
rect 420 1205 427 1209
rect 439 1202 442 1212
rect 455 1202 458 1212
rect 476 1202 479 1212
rect 511 1208 573 1212
rect 577 1208 579 1212
rect 583 1208 587 1212
rect 591 1208 605 1212
rect 609 1208 614 1212
rect 618 1208 623 1212
rect 627 1208 646 1212
rect 650 1208 680 1212
rect 684 1208 695 1212
rect 699 1208 723 1212
rect 727 1208 740 1212
rect 744 1208 764 1212
rect 768 1208 848 1212
rect 852 1208 866 1212
rect 870 1208 875 1212
rect 879 1208 884 1212
rect 888 1208 907 1212
rect 911 1208 941 1212
rect 945 1208 956 1212
rect 960 1208 984 1212
rect 988 1208 997 1212
rect 113 1188 118 1191
rect 122 1188 146 1191
rect 171 1188 178 1191
rect 182 1188 204 1191
rect 224 1188 231 1191
rect 245 1188 250 1191
rect 254 1188 278 1191
rect 303 1188 310 1191
rect 314 1188 336 1191
rect 356 1188 363 1191
rect 377 1188 382 1191
rect 386 1188 410 1191
rect 523 1201 587 1205
rect 591 1201 596 1205
rect 600 1201 646 1205
rect 650 1201 671 1205
rect 675 1201 702 1205
rect 706 1201 735 1205
rect 435 1188 442 1191
rect 446 1188 468 1191
rect 634 1194 635 1198
rect 659 1193 660 1197
rect 706 1194 707 1198
rect 129 1178 136 1181
rect 140 1182 159 1185
rect 159 1175 162 1181
rect 187 1178 194 1181
rect 198 1182 213 1185
rect 261 1178 268 1181
rect 272 1182 291 1185
rect 291 1175 294 1181
rect 319 1178 326 1181
rect 330 1182 345 1185
rect 393 1178 400 1181
rect 404 1182 423 1185
rect 423 1175 426 1181
rect 451 1178 458 1181
rect 462 1182 479 1185
rect 582 1180 585 1185
rect 589 1180 592 1185
rect 572 1177 574 1180
rect 582 1177 592 1180
rect 582 1171 585 1177
rect 96 1159 99 1171
rect 117 1159 120 1171
rect 133 1159 136 1171
rect 147 1162 159 1165
rect 175 1159 178 1171
rect 191 1159 194 1171
rect 212 1159 215 1171
rect 228 1159 231 1171
rect 249 1159 252 1171
rect 265 1159 268 1171
rect 279 1162 291 1165
rect 307 1159 310 1171
rect 323 1159 326 1171
rect 344 1159 347 1171
rect 360 1159 363 1171
rect 381 1159 384 1171
rect 397 1159 400 1171
rect 411 1162 423 1165
rect 439 1159 442 1171
rect 455 1159 458 1171
rect 476 1159 479 1171
rect 589 1171 592 1177
rect 598 1179 601 1185
rect 614 1180 617 1185
rect 598 1175 600 1179
rect 604 1175 606 1179
rect 614 1178 620 1180
rect 624 1178 625 1180
rect 614 1176 625 1178
rect 642 1178 645 1185
rect 598 1171 601 1175
rect 614 1171 617 1176
rect 643 1174 645 1178
rect 642 1171 645 1174
rect 658 1179 661 1185
rect 668 1179 671 1185
rect 689 1180 692 1185
rect 668 1175 677 1179
rect 689 1176 690 1180
rect 694 1177 697 1180
rect 714 1179 717 1185
rect 732 1180 735 1185
rect 771 1182 774 1208
rect 807 1201 826 1205
rect 830 1201 848 1205
rect 852 1201 907 1205
rect 911 1201 932 1205
rect 936 1201 963 1205
rect 967 1201 996 1205
rect 807 1189 810 1201
rect 895 1194 896 1198
rect 920 1193 921 1197
rect 967 1194 968 1198
rect 658 1171 661 1175
rect 668 1171 671 1175
rect 689 1171 692 1176
rect 716 1175 717 1179
rect 834 1180 837 1185
rect 843 1180 846 1185
rect 850 1180 853 1185
rect 714 1171 717 1175
rect 732 1171 735 1176
rect 761 1169 766 1174
rect 770 1170 772 1173
rect 787 1172 790 1178
rect 819 1177 853 1180
rect 787 1169 795 1172
rect 787 1166 790 1169
rect 93 1155 126 1159
rect 130 1155 154 1159
rect 158 1155 184 1159
rect 188 1155 258 1159
rect 262 1155 286 1159
rect 290 1155 316 1159
rect 320 1155 390 1159
rect 394 1155 418 1159
rect 422 1155 448 1159
rect 452 1155 505 1159
rect 642 1156 645 1160
rect 669 1156 670 1160
rect 714 1156 716 1160
rect 819 1163 822 1177
rect 843 1171 846 1177
rect 850 1171 853 1177
rect 859 1179 862 1185
rect 875 1180 878 1185
rect 859 1175 861 1179
rect 865 1175 867 1179
rect 875 1178 881 1180
rect 885 1178 886 1180
rect 875 1176 886 1178
rect 903 1178 906 1185
rect 859 1171 862 1175
rect 875 1171 878 1176
rect 904 1174 906 1178
rect 903 1171 906 1174
rect 919 1179 922 1185
rect 929 1179 932 1185
rect 950 1180 953 1185
rect 929 1175 938 1179
rect 950 1176 951 1180
rect 955 1177 958 1180
rect 975 1179 978 1185
rect 993 1180 996 1185
rect 919 1171 922 1175
rect 929 1171 932 1175
rect 950 1171 953 1176
rect 977 1175 978 1179
rect 975 1171 978 1175
rect 993 1171 996 1176
rect 93 1148 102 1152
rect 106 1148 153 1152
rect 157 1148 203 1152
rect 207 1148 234 1152
rect 238 1148 285 1152
rect 289 1148 335 1152
rect 339 1148 366 1152
rect 370 1148 417 1152
rect 421 1148 467 1152
rect 471 1149 541 1152
rect 585 1149 599 1153
rect 603 1149 630 1153
rect 634 1149 652 1153
rect 656 1149 717 1153
rect 721 1149 735 1153
rect 771 1146 774 1158
rect 903 1156 906 1160
rect 930 1156 931 1160
rect 975 1156 977 1160
rect 811 1149 816 1153
rect 820 1149 860 1153
rect 864 1149 891 1153
rect 895 1149 913 1153
rect 917 1149 978 1153
rect 982 1149 996 1153
rect 100 1142 484 1145
rect 499 1142 572 1146
rect 576 1142 588 1146
rect 592 1142 606 1146
rect 610 1142 617 1146
rect 621 1142 623 1146
rect 627 1142 642 1146
rect 646 1142 679 1146
rect 683 1142 684 1146
rect 688 1142 696 1146
rect 700 1142 724 1146
rect 728 1142 764 1146
rect 768 1142 807 1146
rect 811 1142 818 1146
rect 822 1142 833 1146
rect 837 1142 849 1146
rect 853 1142 867 1146
rect 871 1142 878 1146
rect 882 1142 884 1146
rect 888 1142 903 1146
rect 907 1142 940 1146
rect 944 1142 945 1146
rect 949 1142 957 1146
rect 961 1142 985 1146
rect 989 1142 997 1146
rect 243 1135 352 1138
rect 535 1135 581 1139
rect 585 1135 815 1138
rect 1005 1136 1013 1140
rect 223 1127 227 1131
rect 231 1127 235 1131
rect 523 1128 825 1131
rect 1001 1120 1005 1124
rect 83 1116 211 1120
rect 215 1116 231 1120
rect 247 1116 1026 1120
rect 239 1109 484 1112
rect 559 1109 873 1113
rect 877 1109 909 1113
rect 913 1109 976 1113
rect 980 1109 996 1113
rect 254 1102 484 1105
rect 499 1102 859 1106
rect 863 1102 897 1106
rect 901 1102 925 1106
rect 929 1102 955 1106
rect 959 1102 992 1106
rect 223 1093 227 1097
rect 231 1093 235 1097
rect 867 1092 870 1102
rect 888 1092 891 1102
rect 904 1092 907 1102
rect 918 1095 923 1099
rect 927 1095 934 1099
rect 946 1092 949 1102
rect 962 1092 965 1102
rect 983 1092 986 1102
rect 243 1086 353 1089
rect 93 1079 102 1083
rect 106 1079 138 1083
rect 142 1079 205 1083
rect 209 1079 234 1083
rect 238 1079 270 1083
rect 274 1079 337 1083
rect 341 1079 366 1083
rect 370 1079 402 1083
rect 406 1079 469 1083
rect 473 1079 553 1083
rect 93 1072 126 1076
rect 130 1072 154 1076
rect 158 1072 184 1076
rect 188 1072 221 1076
rect 225 1072 258 1076
rect 262 1072 286 1076
rect 290 1072 316 1076
rect 320 1072 353 1076
rect 357 1072 390 1076
rect 394 1072 418 1076
rect 422 1072 448 1076
rect 452 1072 485 1076
rect 489 1072 493 1076
rect 884 1078 889 1081
rect 893 1078 917 1081
rect 942 1078 949 1081
rect 953 1078 975 1081
rect 96 1062 99 1072
rect 117 1062 120 1072
rect 133 1062 136 1072
rect 147 1065 152 1069
rect 156 1065 163 1069
rect 175 1062 178 1072
rect 191 1062 194 1072
rect 212 1062 215 1072
rect 228 1062 231 1072
rect 249 1062 252 1072
rect 265 1062 268 1072
rect 279 1065 284 1069
rect 288 1065 295 1069
rect 307 1062 310 1072
rect 323 1062 326 1072
rect 344 1062 347 1072
rect 360 1062 363 1072
rect 381 1062 384 1072
rect 397 1062 400 1072
rect 411 1065 416 1069
rect 420 1065 427 1069
rect 439 1062 442 1072
rect 455 1062 458 1072
rect 476 1062 479 1072
rect 900 1068 907 1071
rect 911 1072 930 1075
rect 113 1048 118 1051
rect 122 1048 146 1051
rect 171 1048 178 1051
rect 182 1048 204 1051
rect 224 1048 231 1051
rect 245 1048 250 1051
rect 254 1048 278 1051
rect 303 1048 310 1051
rect 314 1048 336 1051
rect 356 1048 363 1051
rect 377 1048 382 1051
rect 386 1048 410 1051
rect 435 1048 442 1051
rect 446 1048 468 1051
rect 930 1065 933 1071
rect 958 1068 965 1071
rect 969 1072 984 1075
rect 867 1049 870 1061
rect 888 1049 891 1061
rect 904 1049 907 1061
rect 918 1052 930 1055
rect 946 1049 949 1061
rect 962 1049 965 1061
rect 983 1049 986 1061
rect 129 1038 136 1041
rect 140 1042 159 1045
rect 159 1035 162 1041
rect 187 1038 194 1041
rect 198 1042 213 1045
rect 261 1038 268 1041
rect 272 1042 291 1045
rect 291 1035 294 1041
rect 319 1038 326 1041
rect 330 1042 345 1045
rect 393 1038 400 1041
rect 404 1042 423 1045
rect 423 1035 426 1041
rect 451 1038 458 1041
rect 462 1042 479 1045
rect 511 1045 897 1049
rect 901 1045 925 1049
rect 929 1045 955 1049
rect 959 1045 996 1049
rect 547 1038 873 1042
rect 877 1038 924 1042
rect 928 1038 974 1042
rect 978 1038 996 1042
rect 96 1019 99 1031
rect 117 1019 120 1031
rect 133 1019 136 1031
rect 147 1022 159 1025
rect 175 1019 178 1031
rect 191 1019 194 1031
rect 212 1019 215 1031
rect 228 1019 231 1031
rect 249 1019 252 1031
rect 265 1019 268 1031
rect 279 1022 291 1025
rect 307 1019 310 1031
rect 323 1019 326 1031
rect 344 1019 347 1031
rect 360 1019 363 1031
rect 381 1019 384 1031
rect 397 1019 400 1031
rect 411 1022 423 1025
rect 439 1019 442 1031
rect 455 1019 458 1031
rect 476 1019 479 1031
rect 870 1031 991 1034
rect 559 1023 873 1027
rect 877 1023 909 1027
rect 913 1023 976 1027
rect 980 1023 996 1027
rect 93 1015 126 1019
rect 130 1015 154 1019
rect 158 1015 184 1019
rect 188 1015 258 1019
rect 262 1015 286 1019
rect 290 1015 316 1019
rect 320 1015 390 1019
rect 394 1015 418 1019
rect 422 1015 448 1019
rect 452 1015 505 1019
rect 863 1016 897 1020
rect 901 1016 925 1020
rect 929 1016 955 1020
rect 959 1016 992 1020
rect 93 1008 102 1012
rect 106 1008 153 1012
rect 157 1008 203 1012
rect 207 1008 234 1012
rect 238 1008 285 1012
rect 289 1008 335 1012
rect 339 1008 366 1012
rect 370 1008 417 1012
rect 421 1008 467 1012
rect 471 1008 541 1012
rect 867 1006 870 1016
rect 888 1006 891 1016
rect 904 1006 907 1016
rect 918 1009 923 1013
rect 927 1009 934 1013
rect 946 1006 949 1016
rect 962 1006 965 1016
rect 983 1006 986 1016
rect 99 1001 484 1004
rect 93 993 102 997
rect 106 993 138 997
rect 142 993 205 997
rect 209 993 234 997
rect 238 993 270 997
rect 274 993 337 997
rect 341 993 366 997
rect 370 993 402 997
rect 406 993 469 997
rect 473 993 553 997
rect 93 986 126 990
rect 130 986 154 990
rect 158 986 184 990
rect 188 986 221 990
rect 225 986 258 990
rect 262 986 286 990
rect 290 986 316 990
rect 320 986 353 990
rect 357 986 390 990
rect 394 986 418 990
rect 422 986 448 990
rect 452 986 485 990
rect 489 986 493 990
rect 884 992 889 995
rect 893 992 917 995
rect 942 992 949 995
rect 953 992 975 995
rect 96 976 99 986
rect 117 976 120 986
rect 133 976 136 986
rect 147 979 152 983
rect 156 979 163 983
rect 175 976 178 986
rect 191 976 194 986
rect 212 976 215 986
rect 228 976 231 986
rect 249 976 252 986
rect 265 976 268 986
rect 279 979 284 983
rect 288 979 295 983
rect 307 976 310 986
rect 323 976 326 986
rect 344 976 347 986
rect 360 976 363 986
rect 381 976 384 986
rect 397 976 400 986
rect 411 979 416 983
rect 420 979 427 983
rect 439 976 442 986
rect 455 976 458 986
rect 476 976 479 986
rect 900 982 907 985
rect 911 986 930 989
rect 113 962 118 965
rect 122 962 146 965
rect 171 962 178 965
rect 182 962 204 965
rect 224 962 231 965
rect 245 962 250 965
rect 254 962 278 965
rect 303 962 310 965
rect 314 962 336 965
rect 356 962 363 965
rect 377 962 382 965
rect 386 962 410 965
rect 435 962 442 965
rect 446 962 468 965
rect 930 979 933 985
rect 958 982 965 985
rect 969 986 984 989
rect 995 984 1006 988
rect 867 963 870 975
rect 888 963 891 975
rect 904 963 907 975
rect 918 966 930 969
rect 946 963 949 975
rect 962 963 965 975
rect 983 963 986 975
rect 129 952 136 955
rect 140 956 159 959
rect 159 949 162 955
rect 187 952 194 955
rect 198 956 213 959
rect 261 952 268 955
rect 272 956 291 959
rect 291 949 294 955
rect 319 952 326 955
rect 330 956 345 959
rect 393 952 400 955
rect 404 956 423 959
rect 423 949 426 955
rect 451 952 458 955
rect 462 956 479 959
rect 511 959 897 963
rect 901 959 925 963
rect 929 959 955 963
rect 959 959 996 963
rect 547 952 873 956
rect 877 952 924 956
rect 928 952 974 956
rect 978 952 996 956
rect 96 933 99 945
rect 117 933 120 945
rect 133 933 136 945
rect 147 936 159 939
rect 175 933 178 945
rect 191 933 194 945
rect 212 933 215 945
rect 228 933 231 945
rect 249 933 252 945
rect 265 933 268 945
rect 279 936 291 939
rect 307 933 310 945
rect 323 933 326 945
rect 344 933 347 945
rect 360 933 363 945
rect 381 933 384 945
rect 397 933 400 945
rect 411 936 423 939
rect 439 933 442 945
rect 455 933 458 945
rect 476 933 479 945
rect 93 929 126 933
rect 130 929 154 933
rect 158 929 184 933
rect 188 929 258 933
rect 262 929 286 933
rect 290 929 316 933
rect 320 929 390 933
rect 394 929 418 933
rect 422 929 448 933
rect 452 929 505 933
rect 93 922 102 926
rect 106 922 153 926
rect 157 922 203 926
rect 207 922 234 926
rect 238 922 285 926
rect 289 922 335 926
rect 339 922 366 926
rect 370 922 417 926
rect 421 922 467 926
rect 471 922 541 926
rect 99 916 484 919
rect 224 909 328 912
rect 340 901 344 905
rect 348 901 352 905
rect 83 890 328 894
rect 332 890 348 894
rect 364 890 1013 894
rect 1017 890 1026 894
rect 356 883 484 886
rect 371 876 484 879
rect 340 867 344 871
rect 348 867 352 871
rect 224 860 328 863
rect 93 853 102 857
rect 106 853 138 857
rect 142 853 205 857
rect 209 853 234 857
rect 238 853 270 857
rect 274 853 337 857
rect 341 853 366 857
rect 370 853 402 857
rect 406 853 469 857
rect 473 853 553 857
rect 93 846 126 850
rect 130 846 154 850
rect 158 846 184 850
rect 188 846 221 850
rect 225 846 258 850
rect 262 846 286 850
rect 290 846 316 850
rect 320 846 353 850
rect 357 846 390 850
rect 394 846 418 850
rect 422 846 448 850
rect 452 846 485 850
rect 489 846 493 850
rect 96 836 99 846
rect 117 836 120 846
rect 133 836 136 846
rect 147 839 152 843
rect 156 839 163 843
rect 175 836 178 846
rect 191 836 194 846
rect 212 836 215 846
rect 228 836 231 846
rect 249 836 252 846
rect 265 836 268 846
rect 279 839 284 843
rect 288 839 295 843
rect 307 836 310 846
rect 323 836 326 846
rect 344 836 347 846
rect 360 836 363 846
rect 381 836 384 846
rect 397 836 400 846
rect 411 839 416 843
rect 420 839 427 843
rect 439 836 442 846
rect 455 836 458 846
rect 476 836 479 846
rect 113 822 118 825
rect 122 822 146 825
rect 171 822 178 825
rect 182 822 204 825
rect 224 822 231 825
rect 245 822 250 825
rect 254 822 278 825
rect 303 822 310 825
rect 314 822 336 825
rect 356 822 363 825
rect 377 822 382 825
rect 386 822 410 825
rect 435 822 442 825
rect 446 822 468 825
rect 129 812 136 815
rect 140 816 159 819
rect 159 809 162 815
rect 187 812 194 815
rect 198 816 213 819
rect 261 812 268 815
rect 272 816 291 819
rect 291 809 294 815
rect 319 812 326 815
rect 330 816 345 819
rect 393 812 400 815
rect 404 816 423 819
rect 423 809 426 815
rect 451 812 458 815
rect 462 816 479 819
rect 96 793 99 805
rect 117 793 120 805
rect 133 793 136 805
rect 147 796 159 799
rect 175 793 178 805
rect 191 793 194 805
rect 212 793 215 805
rect 228 793 231 805
rect 249 793 252 805
rect 265 793 268 805
rect 279 796 291 799
rect 307 793 310 805
rect 323 793 326 805
rect 344 793 347 805
rect 360 793 363 805
rect 381 793 384 805
rect 397 793 400 805
rect 411 796 423 799
rect 439 793 442 805
rect 455 793 458 805
rect 476 793 479 805
rect 93 789 126 793
rect 130 789 154 793
rect 158 789 184 793
rect 188 789 258 793
rect 262 789 286 793
rect 290 789 316 793
rect 320 789 390 793
rect 394 789 418 793
rect 422 789 448 793
rect 452 789 505 793
rect 93 782 102 786
rect 106 782 153 786
rect 157 782 203 786
rect 207 782 234 786
rect 238 782 285 786
rect 289 782 335 786
rect 339 782 366 786
rect 370 782 417 786
rect 421 782 467 786
rect 471 782 541 786
<< m2contact >>
rect 553 1754 559 1758
rect 574 1754 578 1758
rect 610 1754 614 1758
rect 677 1754 681 1758
rect 706 1754 710 1758
rect 742 1754 746 1758
rect 809 1754 813 1758
rect 838 1754 842 1758
rect 874 1754 878 1758
rect 941 1754 945 1758
rect 970 1754 974 1758
rect 1006 1754 1010 1758
rect 1073 1754 1077 1758
rect 493 1747 499 1751
rect 574 1740 578 1744
rect 624 1740 628 1744
rect 677 1740 681 1744
rect 706 1740 710 1744
rect 756 1740 760 1744
rect 809 1740 813 1744
rect 838 1740 842 1744
rect 888 1740 892 1744
rect 941 1740 945 1744
rect 970 1740 974 1744
rect 1020 1740 1024 1744
rect 1073 1740 1077 1744
rect 597 1729 601 1733
rect 234 1721 238 1725
rect 270 1721 274 1725
rect 337 1721 341 1725
rect 553 1721 559 1725
rect 568 1720 572 1724
rect 581 1723 585 1729
rect 618 1723 622 1729
rect 631 1725 635 1729
rect 655 1729 659 1733
rect 729 1729 733 1733
rect 639 1723 643 1729
rect 676 1723 680 1729
rect 692 1725 696 1729
rect 493 1714 499 1718
rect 234 1707 238 1711
rect 284 1707 288 1711
rect 337 1707 341 1711
rect 581 1710 585 1714
rect 597 1710 601 1716
rect 631 1716 635 1720
rect 618 1710 622 1714
rect 639 1710 643 1714
rect 655 1710 659 1716
rect 700 1720 704 1724
rect 713 1723 717 1729
rect 750 1723 754 1729
rect 763 1725 767 1729
rect 787 1729 791 1733
rect 861 1729 865 1733
rect 771 1723 775 1729
rect 808 1723 812 1729
rect 824 1725 828 1729
rect 676 1710 680 1714
rect 692 1710 696 1714
rect 713 1710 717 1714
rect 729 1710 733 1716
rect 763 1716 767 1720
rect 750 1710 754 1714
rect 771 1710 775 1714
rect 787 1710 791 1716
rect 832 1720 836 1724
rect 845 1723 849 1729
rect 882 1723 886 1729
rect 895 1725 899 1729
rect 919 1729 923 1733
rect 993 1729 997 1733
rect 903 1723 907 1729
rect 940 1723 944 1729
rect 956 1725 960 1729
rect 808 1710 812 1714
rect 824 1710 828 1714
rect 845 1710 849 1714
rect 861 1710 865 1716
rect 895 1716 899 1720
rect 882 1710 886 1714
rect 903 1710 907 1714
rect 919 1710 923 1716
rect 964 1720 968 1724
rect 977 1723 981 1729
rect 1014 1723 1018 1729
rect 1027 1725 1031 1729
rect 1051 1729 1055 1733
rect 1035 1723 1039 1729
rect 1072 1723 1076 1729
rect 1088 1725 1092 1729
rect 940 1710 944 1714
rect 956 1710 960 1714
rect 977 1710 981 1714
rect 993 1710 997 1716
rect 1027 1716 1031 1720
rect 1014 1710 1018 1714
rect 257 1696 261 1700
rect 219 1687 223 1691
rect 241 1690 245 1696
rect 278 1690 282 1696
rect 291 1692 295 1696
rect 315 1696 319 1700
rect 299 1690 303 1696
rect 336 1690 340 1696
rect 352 1690 356 1696
rect 574 1699 578 1703
rect 611 1697 615 1701
rect 631 1697 635 1701
rect 675 1697 679 1701
rect 706 1699 710 1703
rect 743 1697 747 1701
rect 763 1697 767 1701
rect 807 1697 811 1701
rect 838 1699 842 1703
rect 875 1697 879 1701
rect 895 1697 899 1701
rect 939 1697 943 1701
rect 956 1702 960 1706
rect 1035 1710 1039 1714
rect 1051 1710 1055 1716
rect 1072 1710 1076 1714
rect 1088 1710 1092 1714
rect 970 1699 974 1703
rect 1007 1697 1011 1701
rect 1027 1697 1031 1701
rect 1071 1697 1075 1701
rect 1088 1702 1092 1706
rect 505 1690 511 1694
rect 241 1677 245 1681
rect 257 1677 261 1683
rect 291 1683 295 1687
rect 278 1677 282 1681
rect 299 1677 303 1681
rect 315 1677 319 1683
rect 541 1683 547 1687
rect 574 1683 578 1687
rect 625 1683 629 1687
rect 675 1683 679 1687
rect 706 1683 710 1687
rect 757 1683 761 1687
rect 807 1683 811 1687
rect 838 1683 842 1687
rect 889 1683 893 1687
rect 939 1683 943 1687
rect 970 1683 974 1687
rect 1021 1683 1025 1687
rect 1071 1683 1075 1687
rect 336 1677 340 1681
rect 352 1677 356 1681
rect 234 1666 238 1670
rect 271 1664 275 1668
rect 291 1664 295 1668
rect 335 1664 339 1668
rect 493 1670 499 1674
rect 572 1670 576 1674
rect 606 1670 610 1674
rect 623 1670 627 1674
rect 679 1670 683 1674
rect 696 1670 700 1674
rect 724 1670 728 1674
rect 529 1663 535 1667
rect 599 1663 603 1667
rect 630 1663 634 1667
rect 652 1663 656 1667
rect 717 1663 721 1667
rect 505 1657 511 1661
rect 234 1650 238 1654
rect 285 1650 289 1654
rect 335 1650 339 1654
rect 541 1650 547 1654
rect 573 1653 577 1657
rect 598 1656 602 1660
rect 605 1653 609 1657
rect 623 1653 627 1657
rect 645 1656 649 1660
rect 670 1656 674 1660
rect 680 1653 684 1657
rect 696 1653 700 1657
rect 716 1656 720 1660
rect 723 1653 727 1657
rect 787 1663 791 1667
rect 352 1643 356 1647
rect 219 1634 223 1638
rect 344 1636 348 1640
rect 368 1636 372 1640
rect 227 1627 231 1631
rect 368 1627 372 1631
rect 600 1637 604 1641
rect 620 1634 624 1638
rect 639 1638 643 1642
rect 741 1649 745 1653
rect 756 1649 760 1653
rect 658 1637 662 1641
rect 677 1637 681 1641
rect 690 1636 694 1640
rect 712 1637 716 1641
rect 720 1636 724 1640
rect 732 1636 736 1640
rect 573 1623 577 1627
rect 605 1623 609 1627
rect 623 1623 627 1627
rect 680 1623 684 1627
rect 695 1623 699 1627
rect 723 1623 727 1627
rect 234 1619 238 1623
rect 301 1619 305 1623
rect 337 1619 341 1623
rect 553 1619 559 1623
rect 587 1619 591 1623
rect 630 1618 634 1622
rect 652 1619 659 1623
rect 702 1618 706 1622
rect 493 1612 499 1616
rect 234 1605 238 1609
rect 287 1605 291 1609
rect 337 1605 341 1609
rect 517 1611 523 1615
rect 587 1611 591 1615
rect 646 1611 650 1615
rect 671 1611 675 1615
rect 702 1611 706 1615
rect 795 1641 799 1649
rect 868 1663 872 1667
rect 822 1649 826 1653
rect 837 1649 841 1653
rect 818 1641 822 1645
rect 764 1635 768 1639
rect 777 1627 781 1631
rect 876 1641 880 1649
rect 903 1641 907 1645
rect 845 1635 849 1639
rect 858 1627 862 1631
rect 505 1604 511 1608
rect 573 1604 577 1608
rect 587 1604 591 1608
rect 605 1604 609 1608
rect 623 1604 627 1608
rect 646 1604 650 1608
rect 680 1604 684 1608
rect 695 1604 699 1608
rect 723 1604 727 1608
rect 256 1594 260 1598
rect 219 1588 223 1594
rect 235 1588 239 1594
rect 272 1588 276 1594
rect 280 1590 284 1594
rect 314 1594 318 1598
rect 517 1597 523 1601
rect 587 1597 591 1601
rect 646 1597 650 1601
rect 671 1597 675 1601
rect 702 1597 706 1601
rect 293 1588 297 1594
rect 330 1588 334 1594
rect 587 1589 591 1593
rect 630 1590 634 1594
rect 652 1589 659 1593
rect 702 1590 706 1594
rect 352 1585 356 1589
rect 573 1585 577 1589
rect 605 1585 609 1589
rect 623 1585 627 1589
rect 680 1585 684 1589
rect 695 1585 699 1589
rect 723 1585 727 1589
rect 219 1575 223 1579
rect 235 1575 239 1579
rect 280 1581 284 1585
rect 256 1575 260 1581
rect 272 1575 276 1579
rect 293 1575 297 1579
rect 314 1575 318 1581
rect 330 1575 334 1579
rect 568 1573 572 1577
rect 236 1562 240 1566
rect 280 1562 284 1566
rect 300 1562 304 1566
rect 337 1564 341 1568
rect 600 1571 604 1575
rect 620 1574 624 1578
rect 639 1570 643 1574
rect 658 1571 662 1575
rect 677 1571 681 1575
rect 690 1572 694 1576
rect 787 1587 791 1591
rect 868 1587 872 1591
rect 712 1571 716 1575
rect 720 1572 724 1576
rect 732 1572 736 1576
rect 767 1572 771 1576
rect 795 1571 799 1575
rect 847 1572 851 1576
rect 876 1571 880 1575
rect 505 1555 511 1559
rect 573 1555 577 1559
rect 598 1552 602 1556
rect 605 1555 609 1559
rect 623 1555 627 1559
rect 645 1552 649 1556
rect 670 1552 674 1556
rect 680 1555 684 1559
rect 696 1555 700 1559
rect 716 1552 720 1556
rect 723 1555 727 1559
rect 236 1548 240 1552
rect 286 1548 290 1552
rect 337 1548 341 1552
rect 541 1548 547 1552
rect 583 1545 587 1549
rect 599 1545 603 1549
rect 630 1545 634 1549
rect 652 1545 656 1549
rect 717 1545 721 1549
rect 777 1551 781 1555
rect 858 1551 862 1555
rect 493 1538 499 1542
rect 572 1538 576 1542
rect 606 1538 610 1542
rect 623 1538 627 1542
rect 679 1538 683 1542
rect 696 1538 700 1542
rect 724 1538 728 1542
rect 529 1531 535 1535
rect 583 1531 587 1535
rect 599 1531 603 1535
rect 630 1531 634 1535
rect 652 1531 656 1535
rect 717 1531 721 1535
rect 787 1531 791 1535
rect 573 1521 577 1525
rect 598 1524 602 1528
rect 605 1521 609 1525
rect 623 1521 627 1525
rect 645 1524 649 1528
rect 670 1524 674 1528
rect 680 1521 684 1525
rect 696 1521 700 1525
rect 716 1524 720 1528
rect 723 1521 727 1525
rect 567 1504 571 1508
rect 600 1505 604 1509
rect 620 1502 624 1506
rect 639 1506 643 1510
rect 658 1505 662 1509
rect 677 1505 681 1509
rect 690 1504 694 1508
rect 712 1505 716 1509
rect 720 1504 724 1508
rect 732 1504 736 1508
rect 795 1509 799 1517
rect 892 1531 896 1535
rect 846 1517 850 1521
rect 861 1517 865 1521
rect 764 1503 768 1507
rect 818 1508 822 1512
rect 573 1491 577 1495
rect 605 1491 609 1495
rect 623 1491 627 1495
rect 680 1491 684 1495
rect 695 1491 699 1495
rect 723 1491 727 1495
rect 587 1487 591 1491
rect 630 1486 634 1490
rect 652 1487 659 1491
rect 702 1486 706 1490
rect 517 1479 523 1483
rect 587 1479 591 1483
rect 646 1479 650 1483
rect 671 1479 675 1483
rect 702 1479 706 1483
rect 777 1495 781 1499
rect 900 1509 904 1517
rect 921 1509 925 1513
rect 869 1503 873 1507
rect 882 1495 886 1499
rect 505 1472 511 1476
rect 573 1472 577 1476
rect 587 1472 591 1476
rect 605 1472 609 1476
rect 623 1472 627 1476
rect 646 1472 650 1476
rect 680 1472 684 1476
rect 695 1472 699 1476
rect 723 1472 727 1476
rect 517 1465 523 1469
rect 587 1465 591 1469
rect 646 1465 650 1469
rect 671 1465 675 1469
rect 702 1465 706 1469
rect 587 1457 591 1461
rect 630 1458 634 1462
rect 652 1457 659 1461
rect 702 1458 706 1462
rect 573 1453 577 1457
rect 605 1453 609 1457
rect 623 1453 627 1457
rect 680 1453 684 1457
rect 695 1453 699 1457
rect 723 1453 727 1457
rect 787 1456 791 1460
rect 892 1456 896 1460
rect 568 1441 572 1445
rect 600 1439 604 1443
rect 620 1442 624 1446
rect 639 1438 643 1442
rect 658 1439 662 1443
rect 677 1439 681 1443
rect 690 1440 694 1444
rect 712 1439 716 1443
rect 720 1440 724 1444
rect 732 1440 736 1444
rect 766 1441 770 1445
rect 795 1440 799 1444
rect 872 1441 876 1445
rect 900 1440 904 1444
rect 573 1423 577 1427
rect 598 1420 602 1424
rect 605 1423 609 1427
rect 623 1423 627 1427
rect 645 1420 649 1424
rect 670 1420 674 1424
rect 680 1423 684 1427
rect 696 1423 700 1427
rect 716 1420 720 1424
rect 723 1423 727 1427
rect 529 1413 535 1417
rect 599 1413 603 1417
rect 630 1413 634 1417
rect 652 1413 656 1417
rect 717 1413 721 1417
rect 777 1420 781 1424
rect 882 1420 886 1424
rect 493 1406 499 1410
rect 572 1406 576 1410
rect 606 1406 610 1410
rect 623 1406 627 1410
rect 679 1406 683 1410
rect 696 1406 700 1410
rect 724 1406 728 1410
rect 529 1399 535 1403
rect 599 1399 603 1403
rect 630 1399 634 1403
rect 652 1399 656 1403
rect 717 1399 721 1403
rect 787 1399 791 1403
rect 573 1389 577 1393
rect 598 1392 602 1396
rect 605 1389 609 1393
rect 623 1389 627 1393
rect 645 1392 649 1396
rect 670 1392 674 1396
rect 680 1389 684 1393
rect 696 1389 700 1393
rect 716 1392 720 1396
rect 723 1389 727 1393
rect 567 1372 571 1376
rect 600 1373 604 1377
rect 620 1370 624 1374
rect 639 1374 643 1378
rect 658 1373 662 1377
rect 677 1373 681 1377
rect 690 1372 694 1376
rect 712 1373 716 1377
rect 720 1372 724 1376
rect 732 1372 736 1376
rect 795 1377 799 1385
rect 868 1399 872 1403
rect 822 1385 826 1389
rect 837 1385 841 1389
rect 818 1377 822 1381
rect 764 1371 768 1375
rect 573 1359 577 1363
rect 605 1359 609 1363
rect 623 1359 627 1363
rect 680 1359 684 1363
rect 695 1359 699 1363
rect 723 1359 727 1363
rect 587 1355 591 1359
rect 630 1354 634 1358
rect 652 1355 659 1359
rect 702 1354 706 1358
rect 517 1347 523 1351
rect 587 1347 591 1351
rect 646 1347 650 1351
rect 671 1347 675 1351
rect 702 1347 706 1351
rect 777 1363 781 1367
rect 876 1377 880 1385
rect 958 1399 962 1403
rect 912 1385 916 1389
rect 927 1385 931 1389
rect 900 1377 904 1381
rect 845 1371 849 1375
rect 934 1379 938 1383
rect 966 1377 970 1385
rect 858 1363 862 1367
rect 1001 1376 1005 1380
rect 948 1363 952 1367
rect 505 1340 511 1344
rect 573 1340 577 1344
rect 587 1340 591 1344
rect 605 1340 609 1344
rect 623 1340 627 1344
rect 646 1340 650 1344
rect 680 1340 684 1344
rect 695 1340 699 1344
rect 723 1340 727 1344
rect 517 1333 523 1337
rect 587 1333 591 1337
rect 646 1333 650 1337
rect 671 1333 675 1337
rect 702 1333 706 1337
rect 587 1325 591 1329
rect 630 1326 634 1330
rect 652 1325 659 1329
rect 702 1326 706 1330
rect 573 1321 577 1325
rect 605 1321 609 1325
rect 623 1321 627 1325
rect 680 1321 684 1325
rect 695 1321 699 1325
rect 723 1321 727 1325
rect 568 1309 572 1313
rect 600 1307 604 1311
rect 620 1310 624 1314
rect 639 1306 643 1310
rect 658 1307 662 1311
rect 677 1307 681 1311
rect 690 1308 694 1312
rect 787 1321 791 1325
rect 868 1321 872 1325
rect 958 1321 962 1325
rect 712 1307 716 1311
rect 720 1308 724 1312
rect 732 1308 736 1312
rect 767 1306 771 1310
rect 795 1305 799 1309
rect 847 1306 851 1310
rect 876 1305 880 1309
rect 931 1306 935 1310
rect 966 1305 970 1309
rect 573 1291 577 1295
rect 598 1288 602 1292
rect 605 1291 609 1295
rect 623 1291 627 1295
rect 645 1288 649 1292
rect 670 1288 674 1292
rect 680 1291 684 1295
rect 696 1291 700 1295
rect 716 1288 720 1292
rect 723 1291 727 1295
rect 529 1281 535 1285
rect 599 1281 603 1285
rect 630 1281 634 1285
rect 652 1281 656 1285
rect 717 1281 721 1285
rect 777 1285 781 1289
rect 858 1285 862 1289
rect 948 1285 952 1289
rect 493 1274 499 1278
rect 572 1274 576 1278
rect 606 1274 610 1278
rect 623 1274 627 1278
rect 679 1274 683 1278
rect 696 1274 700 1278
rect 724 1274 728 1278
rect 529 1267 535 1271
rect 599 1267 603 1271
rect 630 1267 634 1271
rect 652 1267 656 1271
rect 717 1267 721 1271
rect 787 1267 791 1271
rect 573 1257 577 1261
rect 598 1260 602 1264
rect 605 1257 609 1261
rect 623 1257 627 1261
rect 645 1260 649 1264
rect 670 1260 674 1264
rect 680 1257 684 1261
rect 696 1257 700 1261
rect 716 1260 720 1264
rect 723 1257 727 1261
rect 567 1240 571 1244
rect 600 1241 604 1245
rect 620 1238 624 1242
rect 639 1242 643 1246
rect 658 1241 662 1245
rect 677 1241 681 1245
rect 690 1240 694 1244
rect 712 1241 716 1245
rect 720 1240 724 1244
rect 732 1240 736 1244
rect 795 1245 799 1253
rect 764 1239 768 1243
rect 818 1244 822 1248
rect 573 1227 577 1231
rect 605 1227 609 1231
rect 623 1227 627 1231
rect 680 1227 684 1231
rect 695 1227 699 1231
rect 723 1227 727 1231
rect 587 1223 591 1227
rect 102 1219 106 1223
rect 138 1219 142 1223
rect 205 1219 209 1223
rect 234 1219 238 1223
rect 270 1219 274 1223
rect 337 1219 341 1223
rect 366 1219 370 1223
rect 402 1219 406 1223
rect 469 1219 473 1223
rect 553 1219 559 1223
rect 630 1222 634 1226
rect 652 1223 659 1227
rect 702 1222 706 1226
rect 493 1212 499 1216
rect 587 1215 591 1219
rect 596 1215 600 1219
rect 646 1215 650 1219
rect 671 1215 675 1219
rect 702 1215 706 1219
rect 777 1231 781 1235
rect 102 1205 106 1209
rect 152 1205 156 1209
rect 205 1205 209 1209
rect 234 1205 238 1209
rect 284 1205 288 1209
rect 337 1205 341 1209
rect 366 1205 370 1209
rect 416 1205 420 1209
rect 469 1205 473 1209
rect 505 1208 511 1212
rect 573 1208 577 1212
rect 587 1208 591 1212
rect 605 1208 609 1212
rect 623 1208 627 1212
rect 646 1208 650 1212
rect 680 1208 684 1212
rect 695 1208 699 1212
rect 723 1208 727 1212
rect 848 1208 852 1212
rect 866 1208 870 1212
rect 884 1208 888 1212
rect 907 1208 911 1212
rect 941 1208 945 1212
rect 956 1208 960 1212
rect 984 1208 988 1212
rect 125 1194 129 1198
rect 96 1185 100 1189
rect 109 1188 113 1194
rect 146 1188 150 1194
rect 159 1190 163 1194
rect 183 1194 187 1198
rect 257 1194 261 1198
rect 167 1188 171 1194
rect 204 1188 208 1194
rect 220 1188 224 1194
rect 241 1188 245 1194
rect 278 1188 282 1194
rect 291 1190 295 1194
rect 315 1194 319 1198
rect 389 1194 393 1198
rect 299 1188 303 1194
rect 336 1188 340 1194
rect 352 1188 356 1194
rect 373 1188 377 1194
rect 410 1188 414 1194
rect 423 1190 427 1194
rect 447 1194 451 1198
rect 517 1201 523 1205
rect 587 1201 591 1205
rect 596 1201 600 1205
rect 646 1201 650 1205
rect 671 1201 675 1205
rect 702 1201 706 1205
rect 431 1188 435 1194
rect 468 1188 472 1194
rect 484 1190 488 1194
rect 587 1193 591 1197
rect 630 1194 634 1198
rect 652 1193 659 1197
rect 702 1194 706 1198
rect 573 1189 577 1193
rect 605 1189 609 1193
rect 623 1189 627 1193
rect 680 1189 684 1193
rect 695 1189 699 1193
rect 723 1189 727 1193
rect 109 1175 113 1179
rect 125 1175 129 1181
rect 159 1181 163 1185
rect 146 1175 150 1179
rect 167 1175 171 1179
rect 183 1175 187 1181
rect 204 1175 208 1179
rect 220 1175 224 1179
rect 241 1175 245 1179
rect 257 1175 261 1181
rect 291 1181 295 1185
rect 278 1175 282 1179
rect 299 1175 303 1179
rect 315 1175 319 1181
rect 336 1175 340 1179
rect 352 1175 356 1179
rect 373 1175 377 1179
rect 389 1175 393 1181
rect 423 1181 427 1185
rect 410 1175 414 1179
rect 431 1175 435 1179
rect 447 1175 451 1181
rect 468 1175 472 1179
rect 484 1175 488 1179
rect 568 1177 572 1181
rect 102 1164 106 1168
rect 139 1162 143 1166
rect 159 1162 163 1166
rect 203 1162 207 1166
rect 234 1164 238 1168
rect 271 1162 275 1166
rect 291 1162 295 1166
rect 335 1162 339 1166
rect 366 1164 370 1168
rect 403 1162 407 1166
rect 423 1162 427 1166
rect 467 1162 471 1166
rect 600 1175 604 1179
rect 620 1178 624 1182
rect 639 1174 643 1178
rect 658 1175 662 1179
rect 677 1175 681 1179
rect 690 1176 694 1180
rect 826 1201 830 1205
rect 848 1201 852 1205
rect 907 1201 911 1205
rect 932 1201 936 1205
rect 963 1201 967 1205
rect 848 1193 852 1197
rect 891 1194 895 1198
rect 913 1193 920 1197
rect 963 1194 967 1198
rect 866 1189 870 1193
rect 884 1189 888 1193
rect 941 1189 945 1193
rect 956 1189 960 1193
rect 984 1189 988 1193
rect 787 1185 791 1189
rect 712 1175 716 1179
rect 720 1176 724 1180
rect 732 1176 736 1180
rect 766 1170 770 1174
rect 806 1176 810 1180
rect 795 1169 799 1173
rect 573 1159 577 1163
rect 505 1155 511 1159
rect 598 1156 602 1160
rect 605 1159 609 1163
rect 623 1159 627 1163
rect 645 1156 649 1160
rect 670 1156 674 1160
rect 680 1159 684 1163
rect 696 1159 700 1163
rect 716 1156 720 1160
rect 723 1159 727 1163
rect 861 1175 865 1179
rect 881 1178 885 1182
rect 900 1174 904 1178
rect 919 1175 923 1179
rect 938 1175 942 1179
rect 951 1176 955 1180
rect 973 1175 977 1179
rect 981 1176 985 1180
rect 993 1176 997 1180
rect 807 1159 811 1163
rect 833 1159 837 1163
rect 102 1148 106 1152
rect 153 1148 157 1152
rect 203 1148 207 1152
rect 234 1148 238 1152
rect 285 1148 289 1152
rect 335 1148 339 1152
rect 366 1148 370 1152
rect 417 1148 421 1152
rect 467 1148 471 1152
rect 541 1149 547 1153
rect 581 1149 585 1153
rect 599 1149 603 1153
rect 630 1149 634 1153
rect 652 1149 656 1153
rect 717 1149 721 1153
rect 859 1156 863 1160
rect 866 1159 870 1163
rect 884 1159 888 1163
rect 906 1156 910 1160
rect 931 1156 935 1160
rect 941 1159 945 1163
rect 957 1159 961 1163
rect 977 1156 981 1160
rect 984 1159 988 1163
rect 777 1149 781 1153
rect 816 1149 820 1153
rect 860 1149 864 1153
rect 891 1149 895 1153
rect 913 1149 917 1153
rect 978 1149 982 1153
rect 96 1141 100 1145
rect 484 1141 488 1145
rect 493 1142 499 1146
rect 572 1142 576 1146
rect 606 1142 610 1146
rect 623 1142 627 1146
rect 679 1142 683 1146
rect 696 1142 700 1146
rect 724 1142 728 1146
rect 807 1142 811 1146
rect 833 1142 837 1146
rect 867 1142 871 1146
rect 884 1142 888 1146
rect 940 1142 944 1146
rect 957 1142 961 1146
rect 985 1142 989 1146
rect 219 1134 224 1138
rect 352 1134 356 1138
rect 529 1135 535 1139
rect 581 1135 585 1139
rect 815 1135 819 1139
rect 1001 1136 1005 1140
rect 1013 1136 1017 1140
rect 227 1127 231 1131
rect 517 1127 523 1131
rect 825 1128 829 1132
rect 990 1128 994 1132
rect 211 1123 215 1127
rect 243 1123 247 1127
rect 211 1116 215 1120
rect 243 1116 247 1120
rect 227 1109 231 1113
rect 484 1109 488 1113
rect 553 1109 559 1113
rect 873 1109 877 1113
rect 909 1109 913 1113
rect 976 1109 980 1113
rect 484 1101 488 1105
rect 493 1102 499 1106
rect 859 1102 863 1106
rect 211 1097 215 1101
rect 243 1097 247 1101
rect 227 1093 231 1097
rect 873 1095 877 1099
rect 923 1095 927 1099
rect 976 1095 980 1099
rect 219 1086 224 1090
rect 353 1086 357 1090
rect 896 1084 900 1088
rect 102 1079 106 1083
rect 138 1079 142 1083
rect 205 1079 209 1083
rect 234 1079 238 1083
rect 270 1079 274 1083
rect 337 1079 341 1083
rect 366 1079 370 1083
rect 402 1079 406 1083
rect 469 1079 473 1083
rect 553 1079 559 1083
rect 493 1072 499 1076
rect 867 1075 871 1079
rect 880 1078 884 1084
rect 917 1078 921 1084
rect 930 1080 934 1084
rect 954 1084 958 1088
rect 938 1078 942 1084
rect 975 1078 979 1084
rect 991 1078 995 1084
rect 102 1065 106 1069
rect 152 1065 156 1069
rect 205 1065 209 1069
rect 234 1065 238 1069
rect 284 1065 288 1069
rect 337 1065 341 1069
rect 366 1065 370 1069
rect 416 1065 420 1069
rect 469 1065 473 1069
rect 880 1065 884 1069
rect 896 1065 900 1071
rect 930 1071 934 1075
rect 917 1065 921 1069
rect 125 1054 129 1058
rect 96 1045 100 1049
rect 109 1048 113 1054
rect 146 1048 150 1054
rect 159 1050 163 1054
rect 183 1054 187 1058
rect 257 1054 261 1058
rect 167 1048 171 1054
rect 204 1048 208 1054
rect 220 1048 224 1054
rect 241 1048 245 1054
rect 278 1048 282 1054
rect 291 1050 295 1054
rect 315 1054 319 1058
rect 389 1054 393 1058
rect 299 1048 303 1054
rect 336 1048 340 1054
rect 352 1048 356 1054
rect 373 1048 377 1054
rect 410 1048 414 1054
rect 423 1050 427 1054
rect 447 1054 451 1058
rect 431 1048 435 1054
rect 468 1048 472 1054
rect 484 1050 488 1054
rect 938 1065 942 1069
rect 954 1065 958 1071
rect 975 1065 979 1069
rect 991 1065 995 1069
rect 873 1054 877 1058
rect 910 1052 914 1056
rect 930 1052 934 1056
rect 974 1052 978 1056
rect 109 1035 113 1039
rect 125 1035 129 1041
rect 159 1041 163 1045
rect 146 1035 150 1039
rect 167 1035 171 1039
rect 183 1035 187 1041
rect 204 1035 208 1039
rect 220 1035 224 1039
rect 241 1035 245 1039
rect 257 1035 261 1041
rect 291 1041 295 1045
rect 278 1035 282 1039
rect 299 1035 303 1039
rect 315 1035 319 1041
rect 336 1035 340 1039
rect 352 1035 356 1039
rect 373 1035 377 1039
rect 389 1035 393 1041
rect 423 1041 427 1045
rect 410 1035 414 1039
rect 431 1035 435 1039
rect 447 1035 451 1041
rect 505 1045 511 1049
rect 468 1035 472 1039
rect 484 1035 488 1039
rect 541 1038 547 1042
rect 873 1038 877 1042
rect 924 1038 928 1042
rect 974 1038 978 1042
rect 102 1024 106 1028
rect 139 1022 143 1026
rect 159 1022 163 1026
rect 203 1022 207 1026
rect 234 1024 238 1028
rect 271 1022 275 1026
rect 291 1022 295 1026
rect 335 1022 339 1026
rect 366 1024 370 1028
rect 403 1022 407 1026
rect 423 1022 427 1026
rect 467 1022 471 1026
rect 866 1030 870 1034
rect 991 1031 995 1035
rect 553 1023 559 1027
rect 873 1023 877 1027
rect 909 1023 913 1027
rect 976 1023 980 1027
rect 505 1015 511 1019
rect 859 1016 863 1020
rect 102 1008 106 1012
rect 153 1008 157 1012
rect 203 1008 207 1012
rect 234 1008 238 1012
rect 285 1008 289 1012
rect 335 1008 339 1012
rect 366 1008 370 1012
rect 417 1008 421 1012
rect 467 1008 471 1012
rect 541 1008 547 1012
rect 873 1009 877 1013
rect 923 1009 927 1013
rect 976 1009 980 1013
rect 95 1001 99 1005
rect 484 1001 488 1005
rect 896 998 900 1002
rect 102 993 106 997
rect 138 993 142 997
rect 205 993 209 997
rect 234 993 238 997
rect 270 993 274 997
rect 337 993 341 997
rect 366 993 370 997
rect 402 993 406 997
rect 469 993 473 997
rect 553 993 559 997
rect 493 986 499 990
rect 867 989 871 993
rect 880 992 884 998
rect 917 992 921 998
rect 930 994 934 998
rect 954 998 958 1002
rect 938 992 942 998
rect 975 992 979 998
rect 991 994 995 998
rect 1013 992 1017 996
rect 102 979 106 983
rect 152 979 156 983
rect 205 979 209 983
rect 234 979 238 983
rect 284 979 288 983
rect 337 979 341 983
rect 366 979 370 983
rect 416 979 420 983
rect 469 979 473 983
rect 880 979 884 983
rect 896 979 900 985
rect 930 985 934 989
rect 917 979 921 983
rect 125 968 129 972
rect 96 959 100 963
rect 109 962 113 968
rect 146 962 150 968
rect 159 964 163 968
rect 183 968 187 972
rect 257 968 261 972
rect 167 962 171 968
rect 204 962 208 968
rect 220 962 224 968
rect 241 962 245 968
rect 278 962 282 968
rect 291 964 295 968
rect 315 968 319 972
rect 389 968 393 972
rect 299 962 303 968
rect 336 962 340 968
rect 352 962 356 968
rect 373 962 377 968
rect 410 962 414 968
rect 423 964 427 968
rect 447 968 451 972
rect 431 962 435 968
rect 468 962 472 968
rect 484 964 488 968
rect 938 979 942 983
rect 954 979 958 985
rect 975 979 979 983
rect 991 979 995 988
rect 1013 976 1017 980
rect 873 968 877 972
rect 910 966 914 970
rect 930 966 934 970
rect 974 966 978 970
rect 109 949 113 953
rect 125 949 129 955
rect 159 955 163 959
rect 146 949 150 953
rect 167 949 171 953
rect 183 949 187 955
rect 204 949 208 953
rect 220 949 224 953
rect 241 949 245 953
rect 257 949 261 955
rect 291 955 295 959
rect 278 949 282 953
rect 299 949 303 953
rect 315 949 319 955
rect 336 949 340 953
rect 352 949 356 953
rect 373 949 377 953
rect 389 949 393 955
rect 423 955 427 959
rect 410 949 414 953
rect 431 949 435 953
rect 447 949 451 955
rect 505 959 511 963
rect 468 949 472 953
rect 484 949 488 953
rect 541 952 547 956
rect 873 952 877 956
rect 924 952 928 956
rect 974 952 978 956
rect 102 938 106 942
rect 139 936 143 940
rect 159 936 163 940
rect 203 936 207 940
rect 234 938 238 942
rect 271 936 275 940
rect 291 936 295 940
rect 335 936 339 940
rect 366 938 370 942
rect 403 936 407 940
rect 423 936 427 940
rect 467 936 471 940
rect 505 929 511 933
rect 102 922 106 926
rect 153 922 157 926
rect 203 922 207 926
rect 234 922 238 926
rect 285 922 289 926
rect 335 922 339 926
rect 366 922 370 926
rect 417 922 421 926
rect 467 922 471 926
rect 541 922 547 926
rect 95 915 99 919
rect 484 915 488 919
rect 220 908 224 912
rect 328 908 332 912
rect 352 908 356 912
rect 344 901 348 905
rect 328 897 332 901
rect 360 897 364 901
rect 328 890 332 894
rect 360 890 364 894
rect 1013 890 1017 894
rect 344 883 348 887
rect 484 883 488 887
rect 484 875 488 879
rect 328 871 332 875
rect 360 871 364 875
rect 344 867 348 871
rect 220 860 224 864
rect 328 860 332 864
rect 352 860 356 864
rect 102 853 106 857
rect 138 853 142 857
rect 205 853 209 857
rect 234 853 238 857
rect 270 853 274 857
rect 337 853 341 857
rect 366 853 370 857
rect 402 853 406 857
rect 469 853 473 857
rect 553 853 559 857
rect 493 846 499 850
rect 102 839 106 843
rect 152 839 156 843
rect 205 839 209 843
rect 234 839 238 843
rect 284 839 288 843
rect 337 839 341 843
rect 366 839 370 843
rect 416 839 420 843
rect 469 839 473 843
rect 125 828 129 832
rect 96 819 100 823
rect 109 822 113 828
rect 146 822 150 828
rect 159 824 163 828
rect 183 828 187 832
rect 257 828 261 832
rect 167 822 171 828
rect 204 822 208 828
rect 220 822 224 828
rect 241 822 245 828
rect 278 822 282 828
rect 291 824 295 828
rect 315 828 319 832
rect 389 828 393 832
rect 299 822 303 828
rect 336 822 340 828
rect 352 822 356 828
rect 373 822 377 828
rect 410 822 414 828
rect 423 824 427 828
rect 447 828 451 832
rect 431 822 435 828
rect 468 822 472 828
rect 484 824 488 828
rect 109 809 113 813
rect 125 809 129 815
rect 159 815 163 819
rect 146 809 150 813
rect 167 809 171 813
rect 183 809 187 815
rect 204 809 208 813
rect 220 809 224 813
rect 241 809 245 813
rect 257 809 261 815
rect 291 815 295 819
rect 278 809 282 813
rect 299 809 303 813
rect 315 809 319 815
rect 336 809 340 813
rect 352 809 356 813
rect 373 809 377 813
rect 389 809 393 815
rect 423 815 427 819
rect 410 809 414 813
rect 431 809 435 813
rect 447 809 451 815
rect 468 809 472 813
rect 484 809 488 813
rect 102 798 106 802
rect 139 796 143 800
rect 159 796 163 800
rect 203 796 207 800
rect 234 798 238 802
rect 271 796 275 800
rect 291 796 295 800
rect 335 796 339 800
rect 366 798 370 802
rect 403 796 407 800
rect 423 796 427 800
rect 467 796 471 800
rect 505 789 511 793
rect 102 782 106 786
rect 153 782 157 786
rect 203 782 207 786
rect 234 782 238 786
rect 285 782 289 786
rect 335 782 339 786
rect 366 782 370 786
rect 417 782 421 786
rect 467 782 471 786
rect 541 782 547 786
<< metal2 >>
rect 219 1638 222 1687
rect 219 1594 222 1634
rect 227 1631 231 1774
rect 235 1711 238 1721
rect 242 1681 245 1690
rect 258 1683 261 1696
rect 271 1668 274 1721
rect 338 1711 341 1721
rect 278 1696 282 1700
rect 279 1681 282 1690
rect 234 1654 237 1666
rect 275 1664 276 1668
rect 285 1654 288 1707
rect 291 1687 294 1692
rect 300 1681 303 1690
rect 316 1683 319 1696
rect 337 1681 340 1690
rect 336 1654 339 1664
rect 219 1579 222 1588
rect 103 1209 106 1219
rect 110 1179 113 1188
rect 126 1181 129 1194
rect 139 1166 142 1219
rect 206 1209 209 1219
rect 146 1194 150 1198
rect 147 1179 150 1188
rect 102 1152 105 1164
rect 143 1162 144 1166
rect 153 1152 156 1205
rect 159 1185 162 1190
rect 168 1179 171 1188
rect 184 1181 187 1194
rect 205 1179 208 1188
rect 221 1179 224 1188
rect 204 1152 207 1162
rect 96 1049 99 1141
rect 221 1138 224 1175
rect 227 1131 231 1627
rect 344 1640 348 1774
rect 493 1751 499 1765
rect 493 1718 499 1747
rect 353 1688 356 1690
rect 353 1681 356 1684
rect 353 1647 356 1677
rect 493 1674 499 1714
rect 234 1609 237 1619
rect 235 1579 238 1588
rect 256 1581 259 1594
rect 272 1579 275 1588
rect 281 1585 284 1590
rect 236 1552 239 1562
rect 287 1552 290 1605
rect 293 1594 297 1598
rect 293 1579 296 1588
rect 301 1566 304 1619
rect 337 1609 340 1619
rect 314 1581 317 1594
rect 330 1579 333 1588
rect 299 1562 300 1566
rect 338 1552 341 1564
rect 235 1209 238 1219
rect 242 1179 245 1188
rect 258 1181 261 1194
rect 271 1166 274 1219
rect 338 1209 341 1219
rect 278 1194 282 1198
rect 279 1179 282 1188
rect 234 1152 237 1164
rect 275 1162 276 1166
rect 285 1152 288 1205
rect 291 1185 294 1190
rect 300 1179 303 1188
rect 316 1181 319 1194
rect 337 1179 340 1188
rect 336 1152 339 1162
rect 211 1120 215 1123
rect 211 1101 215 1116
rect 227 1113 231 1127
rect 243 1127 247 1131
rect 243 1120 247 1123
rect 243 1101 247 1116
rect 227 1097 231 1098
rect 243 1093 247 1097
rect 103 1069 106 1079
rect 110 1039 113 1048
rect 126 1041 129 1054
rect 139 1026 142 1079
rect 206 1069 209 1079
rect 146 1054 150 1058
rect 147 1039 150 1048
rect 102 1012 105 1024
rect 143 1022 144 1026
rect 153 1012 156 1065
rect 221 1054 224 1086
rect 159 1045 162 1050
rect 168 1039 171 1048
rect 184 1041 187 1054
rect 205 1039 208 1048
rect 221 1039 224 1048
rect 204 1012 207 1022
rect 96 963 99 1001
rect 103 983 106 993
rect 110 953 113 962
rect 126 955 129 968
rect 139 940 142 993
rect 206 983 209 993
rect 146 968 150 972
rect 147 953 150 962
rect 102 926 105 938
rect 143 936 144 940
rect 153 926 156 979
rect 159 959 162 964
rect 168 953 171 962
rect 184 955 187 968
rect 205 953 208 962
rect 221 953 224 962
rect 204 926 207 936
rect 96 823 99 915
rect 221 912 224 949
rect 103 843 106 853
rect 110 813 113 822
rect 126 815 129 828
rect 139 800 142 853
rect 206 843 209 853
rect 146 828 150 832
rect 147 813 150 822
rect 102 786 105 798
rect 143 796 144 800
rect 153 786 156 839
rect 221 828 224 860
rect 159 819 162 824
rect 168 813 171 822
rect 184 815 187 828
rect 205 813 208 822
rect 221 813 224 822
rect 204 786 207 796
rect 227 779 231 1093
rect 235 1069 238 1079
rect 242 1039 245 1048
rect 258 1041 261 1054
rect 271 1026 274 1079
rect 338 1069 341 1079
rect 278 1054 282 1058
rect 279 1039 282 1048
rect 234 1012 237 1024
rect 275 1022 276 1026
rect 285 1012 288 1065
rect 291 1045 294 1050
rect 300 1039 303 1048
rect 316 1041 319 1054
rect 337 1039 340 1048
rect 336 1012 339 1022
rect 235 983 238 993
rect 242 953 245 962
rect 258 955 261 968
rect 271 940 274 993
rect 338 983 341 993
rect 278 968 282 972
rect 279 953 282 962
rect 234 926 237 938
rect 275 936 276 940
rect 285 926 288 979
rect 291 959 294 964
rect 300 953 303 962
rect 316 955 319 968
rect 337 953 340 962
rect 336 926 339 936
rect 344 905 348 1636
rect 368 1631 372 1636
rect 493 1616 499 1670
rect 493 1542 499 1612
rect 493 1410 499 1538
rect 493 1278 499 1406
rect 367 1209 370 1219
rect 353 1179 356 1188
rect 374 1179 377 1188
rect 390 1181 393 1194
rect 353 1138 356 1175
rect 403 1166 406 1219
rect 470 1209 473 1219
rect 493 1216 499 1274
rect 410 1194 414 1198
rect 411 1179 414 1188
rect 366 1152 369 1164
rect 407 1162 408 1166
rect 417 1152 420 1205
rect 423 1185 426 1190
rect 432 1179 435 1188
rect 448 1181 451 1194
rect 469 1179 472 1188
rect 485 1179 488 1190
rect 468 1152 471 1162
rect 485 1145 488 1175
rect 485 1113 488 1141
rect 493 1146 499 1212
rect 493 1106 499 1142
rect 353 1054 356 1086
rect 367 1069 370 1079
rect 353 1039 356 1048
rect 374 1039 377 1048
rect 390 1041 393 1054
rect 403 1026 406 1079
rect 470 1069 473 1079
rect 410 1054 414 1058
rect 411 1039 414 1048
rect 366 1012 369 1024
rect 407 1022 408 1026
rect 417 1012 420 1065
rect 485 1054 488 1101
rect 423 1045 426 1050
rect 432 1039 435 1048
rect 448 1041 451 1054
rect 469 1039 472 1048
rect 485 1039 488 1050
rect 468 1012 471 1022
rect 485 1005 488 1035
rect 493 1076 499 1102
rect 367 983 370 993
rect 353 953 356 962
rect 374 953 377 962
rect 390 955 393 968
rect 353 912 356 949
rect 403 940 406 993
rect 470 983 473 993
rect 493 990 499 1072
rect 410 968 414 972
rect 411 953 414 962
rect 366 926 369 938
rect 407 936 408 940
rect 417 926 420 979
rect 423 959 426 964
rect 432 953 435 962
rect 448 955 451 968
rect 469 953 472 962
rect 485 953 488 964
rect 468 926 471 936
rect 485 919 488 949
rect 328 894 332 897
rect 328 875 332 890
rect 344 887 348 901
rect 360 901 364 905
rect 360 894 364 897
rect 360 875 364 890
rect 485 887 488 915
rect 344 871 348 872
rect 360 867 364 871
rect 235 843 238 853
rect 242 813 245 822
rect 258 815 261 828
rect 271 800 274 853
rect 338 843 341 853
rect 278 828 282 832
rect 279 813 282 822
rect 234 786 237 798
rect 275 796 276 800
rect 285 786 288 839
rect 291 819 294 824
rect 300 813 303 822
rect 316 815 319 828
rect 337 813 340 822
rect 336 786 339 796
rect 344 779 348 867
rect 353 828 356 860
rect 367 843 370 853
rect 353 813 356 822
rect 374 813 377 822
rect 390 815 393 828
rect 403 800 406 853
rect 470 843 473 853
rect 410 828 414 832
rect 411 813 414 822
rect 366 786 369 798
rect 407 796 408 800
rect 417 786 420 839
rect 485 828 488 875
rect 423 819 426 824
rect 432 813 435 822
rect 448 815 451 828
rect 469 813 472 822
rect 485 820 488 824
rect 493 850 499 986
rect 485 813 488 816
rect 468 786 471 796
rect 493 779 499 846
rect 505 1694 511 1765
rect 505 1661 511 1690
rect 505 1608 511 1657
rect 505 1559 511 1604
rect 505 1476 511 1555
rect 505 1344 511 1472
rect 505 1212 511 1340
rect 505 1159 511 1208
rect 505 1049 511 1155
rect 505 1019 511 1045
rect 505 963 511 1015
rect 505 933 511 959
rect 505 793 511 929
rect 505 779 511 789
rect 517 1615 523 1765
rect 517 1601 523 1611
rect 517 1483 523 1597
rect 517 1469 523 1479
rect 517 1351 523 1465
rect 517 1337 523 1347
rect 517 1205 523 1333
rect 517 1131 523 1201
rect 517 779 523 1127
rect 529 1667 535 1765
rect 529 1535 535 1663
rect 529 1417 535 1531
rect 529 1403 535 1413
rect 529 1285 535 1399
rect 529 1271 535 1281
rect 529 1139 535 1267
rect 529 779 535 1135
rect 541 1687 547 1765
rect 541 1654 547 1683
rect 541 1552 547 1650
rect 541 1153 547 1548
rect 541 1042 547 1149
rect 541 1012 547 1038
rect 541 956 547 1008
rect 541 926 547 952
rect 541 786 547 922
rect 541 779 547 782
rect 553 1758 559 1765
rect 553 1725 559 1754
rect 575 1744 578 1754
rect 553 1623 559 1721
rect 582 1714 585 1723
rect 598 1716 601 1729
rect 611 1701 614 1754
rect 678 1744 681 1754
rect 707 1744 710 1754
rect 618 1729 622 1733
rect 619 1714 622 1723
rect 574 1687 577 1699
rect 615 1697 616 1701
rect 625 1687 628 1740
rect 631 1720 634 1725
rect 640 1714 643 1723
rect 656 1716 659 1729
rect 677 1714 680 1723
rect 693 1723 696 1725
rect 693 1720 700 1723
rect 693 1714 696 1720
rect 714 1714 717 1723
rect 730 1716 733 1729
rect 676 1687 679 1697
rect 693 1680 696 1710
rect 743 1701 746 1754
rect 810 1744 813 1754
rect 839 1744 842 1754
rect 750 1729 754 1733
rect 751 1714 754 1723
rect 706 1687 709 1699
rect 747 1697 748 1701
rect 757 1687 760 1740
rect 763 1720 766 1725
rect 772 1714 775 1723
rect 788 1716 791 1729
rect 809 1714 812 1723
rect 825 1723 828 1725
rect 825 1720 832 1723
rect 825 1714 828 1720
rect 846 1714 849 1723
rect 862 1716 865 1729
rect 808 1687 811 1697
rect 693 1677 745 1680
rect 573 1657 576 1670
rect 599 1660 602 1663
rect 606 1657 609 1670
rect 623 1657 626 1670
rect 553 1223 559 1619
rect 573 1608 576 1623
rect 587 1615 590 1619
rect 605 1608 608 1623
rect 624 1608 627 1623
rect 630 1622 633 1663
rect 646 1615 649 1656
rect 652 1623 655 1663
rect 671 1615 674 1656
rect 680 1657 683 1670
rect 696 1657 699 1670
rect 717 1660 720 1663
rect 724 1657 727 1670
rect 742 1666 745 1677
rect 825 1674 828 1710
rect 875 1701 878 1754
rect 942 1744 945 1754
rect 971 1744 974 1754
rect 882 1729 886 1733
rect 883 1714 886 1723
rect 838 1687 841 1699
rect 879 1697 880 1701
rect 889 1687 892 1740
rect 895 1720 898 1725
rect 904 1714 907 1723
rect 920 1716 923 1729
rect 941 1714 944 1723
rect 957 1723 960 1725
rect 957 1720 964 1723
rect 957 1714 960 1720
rect 978 1714 981 1723
rect 994 1716 997 1729
rect 940 1687 943 1697
rect 957 1680 960 1702
rect 1007 1701 1010 1754
rect 1074 1744 1077 1754
rect 1014 1729 1018 1733
rect 1015 1714 1018 1723
rect 970 1687 973 1699
rect 1011 1697 1012 1701
rect 1021 1687 1024 1740
rect 1027 1720 1030 1725
rect 1036 1714 1039 1723
rect 1052 1716 1055 1729
rect 1073 1714 1076 1723
rect 1089 1723 1092 1725
rect 1089 1720 1093 1723
rect 1089 1714 1092 1720
rect 1089 1706 1092 1710
rect 1072 1687 1075 1697
rect 823 1669 828 1674
rect 885 1676 960 1680
rect 742 1663 787 1666
rect 742 1653 745 1663
rect 760 1650 780 1653
rect 777 1631 780 1650
rect 680 1608 683 1623
rect 695 1608 698 1623
rect 702 1615 706 1618
rect 723 1608 726 1623
rect 573 1589 576 1604
rect 587 1593 590 1597
rect 605 1589 608 1604
rect 624 1589 627 1604
rect 573 1542 576 1555
rect 599 1549 602 1552
rect 573 1525 576 1538
rect 583 1535 587 1545
rect 606 1542 609 1555
rect 623 1542 626 1555
rect 630 1549 633 1590
rect 646 1556 649 1597
rect 652 1549 655 1589
rect 671 1556 674 1597
rect 680 1589 683 1604
rect 695 1589 698 1604
rect 702 1594 706 1597
rect 723 1589 726 1604
rect 680 1542 683 1555
rect 599 1528 602 1531
rect 606 1525 609 1538
rect 623 1525 626 1538
rect 573 1476 576 1491
rect 587 1483 590 1487
rect 605 1476 608 1491
rect 624 1476 627 1491
rect 630 1490 633 1531
rect 646 1483 649 1524
rect 652 1491 655 1531
rect 671 1483 674 1524
rect 680 1525 683 1538
rect 696 1542 699 1555
rect 717 1549 720 1552
rect 724 1542 727 1555
rect 777 1555 780 1627
rect 788 1591 791 1663
rect 823 1666 826 1669
rect 823 1663 868 1666
rect 823 1653 826 1663
rect 696 1525 699 1538
rect 717 1528 720 1531
rect 724 1525 727 1538
rect 777 1521 780 1551
rect 788 1535 791 1587
rect 795 1575 799 1641
rect 783 1531 787 1534
rect 776 1518 780 1521
rect 777 1499 780 1518
rect 680 1476 683 1491
rect 695 1476 698 1491
rect 702 1483 706 1486
rect 723 1476 726 1491
rect 573 1457 576 1472
rect 587 1461 590 1465
rect 605 1457 608 1472
rect 624 1457 627 1472
rect 573 1410 576 1423
rect 599 1417 602 1420
rect 573 1393 576 1406
rect 606 1410 609 1423
rect 623 1410 626 1423
rect 630 1417 633 1458
rect 646 1424 649 1465
rect 652 1417 655 1457
rect 671 1424 674 1465
rect 680 1457 683 1472
rect 695 1457 698 1472
rect 702 1462 706 1465
rect 723 1457 726 1472
rect 680 1410 683 1423
rect 599 1396 602 1399
rect 606 1393 609 1406
rect 623 1393 626 1406
rect 573 1344 576 1359
rect 587 1351 590 1355
rect 605 1344 608 1359
rect 624 1344 627 1359
rect 630 1358 633 1399
rect 646 1351 649 1392
rect 652 1359 655 1399
rect 671 1351 674 1392
rect 680 1393 683 1406
rect 696 1410 699 1423
rect 717 1417 720 1420
rect 724 1410 727 1423
rect 777 1424 780 1495
rect 788 1460 791 1531
rect 696 1393 699 1406
rect 717 1396 720 1399
rect 724 1393 727 1406
rect 777 1367 780 1420
rect 788 1403 791 1456
rect 795 1444 799 1509
rect 783 1399 787 1402
rect 826 1402 829 1653
rect 841 1650 861 1653
rect 858 1631 861 1650
rect 858 1555 861 1627
rect 869 1591 872 1663
rect 876 1575 880 1641
rect 885 1542 888 1676
rect 1089 1673 1092 1702
rect 913 1670 1020 1673
rect 847 1538 888 1542
rect 847 1534 850 1538
rect 847 1531 892 1534
rect 847 1521 850 1531
rect 865 1518 885 1521
rect 847 1516 850 1517
rect 882 1499 885 1518
rect 882 1424 885 1495
rect 893 1460 896 1531
rect 900 1444 904 1509
rect 680 1344 683 1359
rect 695 1344 698 1359
rect 702 1351 706 1354
rect 723 1344 726 1359
rect 573 1325 576 1340
rect 587 1329 590 1333
rect 605 1325 608 1340
rect 624 1325 627 1340
rect 573 1278 576 1291
rect 599 1285 602 1288
rect 573 1261 576 1274
rect 606 1278 609 1291
rect 623 1278 626 1291
rect 630 1285 633 1326
rect 646 1292 649 1333
rect 652 1285 655 1325
rect 671 1292 674 1333
rect 680 1325 683 1340
rect 695 1325 698 1340
rect 702 1330 706 1333
rect 723 1325 726 1340
rect 680 1278 683 1291
rect 599 1264 602 1267
rect 606 1261 609 1274
rect 623 1261 626 1274
rect 553 1113 559 1219
rect 573 1212 576 1227
rect 587 1219 590 1223
rect 573 1193 576 1208
rect 596 1205 600 1215
rect 605 1212 608 1227
rect 624 1212 627 1227
rect 630 1226 633 1267
rect 646 1219 649 1260
rect 652 1227 655 1267
rect 671 1219 674 1260
rect 680 1261 683 1274
rect 696 1278 699 1291
rect 717 1285 720 1288
rect 724 1278 727 1291
rect 777 1289 780 1363
rect 788 1325 791 1399
rect 823 1399 868 1402
rect 823 1389 826 1399
rect 841 1386 861 1389
rect 696 1261 699 1274
rect 717 1264 720 1267
rect 724 1261 727 1274
rect 777 1235 780 1285
rect 788 1271 791 1321
rect 795 1309 799 1377
rect 858 1367 861 1386
rect 858 1289 861 1363
rect 869 1325 872 1399
rect 913 1402 916 1670
rect 1024 1670 1092 1673
rect 913 1399 958 1402
rect 913 1389 916 1399
rect 931 1386 951 1389
rect 876 1309 880 1377
rect 948 1367 951 1386
rect 948 1289 951 1363
rect 959 1325 962 1399
rect 966 1309 970 1377
rect 783 1267 787 1270
rect 680 1212 683 1227
rect 695 1212 698 1227
rect 702 1219 706 1222
rect 723 1212 726 1227
rect 587 1197 590 1201
rect 605 1193 608 1208
rect 624 1193 627 1208
rect 573 1146 576 1159
rect 599 1153 602 1156
rect 581 1139 585 1149
rect 606 1146 609 1159
rect 623 1146 626 1159
rect 630 1153 633 1194
rect 646 1160 649 1201
rect 652 1153 655 1193
rect 671 1160 674 1201
rect 680 1193 683 1208
rect 695 1193 698 1208
rect 702 1198 706 1201
rect 723 1193 726 1208
rect 680 1146 683 1159
rect 696 1146 699 1159
rect 717 1153 720 1156
rect 724 1146 727 1159
rect 777 1153 780 1231
rect 788 1189 791 1267
rect 795 1173 799 1245
rect 807 1146 811 1159
rect 816 1139 819 1149
rect 826 1132 829 1201
rect 848 1197 851 1201
rect 866 1193 869 1208
rect 885 1193 888 1208
rect 833 1146 837 1159
rect 860 1153 863 1156
rect 867 1146 870 1159
rect 884 1146 887 1159
rect 891 1153 894 1194
rect 907 1160 910 1201
rect 913 1153 916 1193
rect 932 1160 935 1201
rect 941 1193 944 1208
rect 956 1193 959 1208
rect 963 1198 967 1201
rect 984 1193 987 1208
rect 941 1146 944 1159
rect 957 1146 960 1159
rect 978 1153 981 1156
rect 985 1146 988 1159
rect 1001 1140 1005 1376
rect 994 1128 995 1131
rect 553 1083 559 1109
rect 553 1027 559 1079
rect 553 997 559 1023
rect 859 1020 863 1102
rect 874 1099 877 1109
rect 881 1069 884 1078
rect 897 1071 900 1084
rect 910 1056 913 1109
rect 977 1099 980 1109
rect 917 1084 921 1088
rect 918 1069 921 1078
rect 873 1042 876 1054
rect 914 1052 915 1056
rect 924 1042 927 1095
rect 992 1084 995 1128
rect 930 1075 933 1080
rect 939 1069 942 1078
rect 955 1071 958 1084
rect 976 1069 979 1078
rect 992 1069 995 1078
rect 975 1042 978 1052
rect 992 1035 995 1065
rect 553 857 559 993
rect 867 993 870 1030
rect 874 1013 877 1023
rect 881 983 884 992
rect 897 985 900 998
rect 910 970 913 1023
rect 977 1013 980 1023
rect 917 998 921 1002
rect 918 983 921 992
rect 873 956 876 968
rect 914 966 915 970
rect 924 956 927 1009
rect 930 989 933 994
rect 939 983 942 992
rect 955 985 958 998
rect 976 983 979 992
rect 992 993 995 994
rect 1013 996 1017 1136
rect 992 988 995 989
rect 975 956 978 966
rect 1013 894 1017 976
rect 553 779 559 853
<< m3contact >>
rect 96 1181 100 1185
rect 353 1684 357 1688
rect 352 1581 356 1585
rect 485 816 489 820
rect 564 1720 568 1724
rect 604 1637 609 1642
rect 615 1633 620 1638
rect 638 1642 643 1647
rect 662 1637 667 1642
rect 677 1641 682 1647
rect 707 1637 712 1642
rect 736 1636 741 1641
rect 691 1631 696 1636
rect 720 1631 724 1636
rect 762 1630 767 1635
rect 568 1577 573 1582
rect 604 1570 609 1575
rect 615 1574 620 1579
rect 638 1565 643 1570
rect 662 1570 667 1575
rect 691 1576 696 1581
rect 720 1576 724 1581
rect 677 1565 682 1571
rect 707 1570 712 1575
rect 736 1571 741 1576
rect 762 1571 767 1576
rect 567 1508 572 1513
rect 604 1505 609 1510
rect 615 1501 620 1506
rect 638 1510 643 1515
rect 662 1505 667 1510
rect 818 1636 823 1641
rect 677 1509 682 1515
rect 707 1505 712 1510
rect 736 1504 741 1509
rect 691 1499 696 1504
rect 720 1499 724 1504
rect 762 1498 767 1503
rect 568 1445 573 1450
rect 604 1438 609 1443
rect 615 1442 620 1447
rect 638 1433 643 1438
rect 662 1438 667 1443
rect 691 1444 696 1449
rect 720 1444 724 1449
rect 677 1433 682 1439
rect 707 1438 712 1443
rect 736 1439 741 1444
rect 761 1440 766 1445
rect 567 1376 572 1381
rect 604 1373 609 1378
rect 615 1369 620 1374
rect 638 1378 643 1383
rect 662 1373 667 1378
rect 677 1377 682 1383
rect 707 1373 712 1378
rect 736 1372 741 1377
rect 691 1367 696 1372
rect 720 1367 724 1372
rect 762 1366 767 1371
rect 818 1512 823 1517
rect 843 1630 848 1635
rect 842 1571 847 1576
rect 903 1636 908 1641
rect 867 1498 872 1503
rect 867 1440 872 1445
rect 568 1313 573 1318
rect 604 1306 609 1311
rect 615 1310 620 1315
rect 638 1301 643 1306
rect 662 1306 667 1311
rect 691 1312 696 1317
rect 720 1312 724 1317
rect 677 1301 682 1307
rect 707 1306 712 1311
rect 736 1307 741 1312
rect 762 1305 767 1310
rect 567 1244 572 1249
rect 604 1241 609 1246
rect 615 1237 620 1242
rect 638 1246 643 1251
rect 662 1241 667 1246
rect 677 1245 682 1251
rect 707 1241 712 1246
rect 736 1240 741 1245
rect 691 1235 696 1240
rect 720 1235 724 1240
rect 762 1234 767 1239
rect 818 1372 823 1377
rect 843 1366 848 1371
rect 842 1305 847 1310
rect 1020 1669 1024 1673
rect 925 1509 930 1514
rect 900 1381 905 1386
rect 934 1374 939 1379
rect 931 1301 936 1306
rect 568 1181 573 1186
rect 604 1174 609 1179
rect 615 1178 620 1183
rect 638 1169 643 1174
rect 662 1174 667 1179
rect 691 1180 696 1185
rect 720 1180 724 1185
rect 677 1169 682 1175
rect 707 1174 712 1179
rect 736 1175 741 1180
rect 761 1169 766 1174
rect 818 1248 823 1253
rect 806 1180 811 1185
rect 865 1174 870 1179
rect 876 1178 881 1183
rect 899 1169 904 1174
rect 923 1174 928 1179
rect 952 1180 957 1185
rect 981 1180 985 1185
rect 938 1169 943 1175
rect 968 1174 973 1179
rect 993 1180 998 1185
rect 867 1071 871 1075
rect 992 989 996 993
<< metal3 >>
rect 563 1724 569 1725
rect 563 1720 564 1724
rect 568 1720 569 1724
rect 563 1719 569 1720
rect 563 1689 568 1719
rect 352 1688 568 1689
rect 352 1684 353 1688
rect 357 1684 568 1688
rect 352 1683 358 1684
rect 1019 1673 1025 1674
rect 1019 1669 1020 1673
rect 1024 1669 1025 1673
rect 1019 1668 1025 1669
rect 604 1647 644 1648
rect 604 1643 638 1647
rect 603 1642 610 1643
rect 603 1637 604 1642
rect 609 1637 610 1642
rect 637 1642 638 1643
rect 643 1642 644 1647
rect 676 1647 712 1652
rect 637 1641 644 1642
rect 661 1642 668 1643
rect 603 1636 610 1637
rect 614 1638 621 1639
rect 614 1633 615 1638
rect 620 1633 621 1638
rect 661 1637 662 1642
rect 667 1637 668 1642
rect 676 1641 677 1647
rect 682 1646 712 1647
rect 682 1641 683 1646
rect 707 1643 712 1646
rect 676 1640 683 1641
rect 706 1642 713 1643
rect 706 1637 707 1642
rect 712 1637 713 1642
rect 735 1641 742 1642
rect 661 1636 668 1637
rect 690 1636 697 1637
rect 706 1636 713 1637
rect 719 1636 725 1637
rect 662 1633 667 1636
rect 614 1628 667 1633
rect 690 1631 691 1636
rect 696 1631 697 1636
rect 719 1631 720 1636
rect 724 1631 725 1636
rect 690 1630 725 1631
rect 691 1626 725 1630
rect 735 1636 736 1641
rect 741 1636 742 1641
rect 817 1641 824 1642
rect 817 1636 818 1641
rect 823 1636 824 1641
rect 902 1641 909 1642
rect 902 1636 903 1641
rect 908 1636 909 1641
rect 735 1635 742 1636
rect 761 1635 768 1636
rect 817 1635 824 1636
rect 842 1635 849 1636
rect 902 1635 909 1636
rect 735 1630 762 1635
rect 767 1630 768 1635
rect 818 1630 843 1635
rect 848 1630 849 1635
rect 735 1609 740 1630
rect 761 1629 768 1630
rect 842 1629 849 1630
rect 899 1630 908 1635
rect 568 1603 740 1609
rect 351 1585 357 1586
rect 351 1581 352 1585
rect 356 1581 489 1585
rect 568 1583 573 1603
rect 351 1580 489 1581
rect 95 1185 101 1186
rect 95 1181 96 1185
rect 100 1181 101 1185
rect 95 1180 101 1181
rect 484 821 489 1580
rect 567 1582 574 1583
rect 567 1577 568 1582
rect 573 1577 574 1582
rect 567 1576 574 1577
rect 614 1579 667 1584
rect 691 1582 725 1586
rect 603 1575 610 1576
rect 603 1570 604 1575
rect 609 1570 610 1575
rect 614 1574 615 1579
rect 620 1574 621 1579
rect 662 1576 667 1579
rect 690 1581 725 1582
rect 690 1576 691 1581
rect 696 1576 697 1581
rect 719 1576 720 1581
rect 724 1576 725 1581
rect 614 1573 621 1574
rect 661 1575 668 1576
rect 690 1575 697 1576
rect 706 1575 713 1576
rect 719 1575 725 1576
rect 735 1576 742 1577
rect 761 1576 768 1577
rect 841 1576 848 1577
rect 603 1569 610 1570
rect 637 1570 644 1571
rect 637 1569 638 1570
rect 604 1565 638 1569
rect 643 1565 644 1570
rect 661 1570 662 1575
rect 667 1570 668 1575
rect 661 1569 668 1570
rect 676 1571 683 1572
rect 604 1564 644 1565
rect 676 1565 677 1571
rect 682 1566 683 1571
rect 706 1570 707 1575
rect 712 1570 713 1575
rect 735 1571 736 1576
rect 741 1571 762 1576
rect 767 1571 768 1576
rect 735 1570 742 1571
rect 761 1570 768 1571
rect 818 1571 842 1576
rect 847 1571 848 1576
rect 706 1569 713 1570
rect 707 1566 712 1569
rect 682 1565 712 1566
rect 676 1560 712 1565
rect 736 1543 741 1570
rect 567 1537 741 1543
rect 567 1514 572 1537
rect 604 1515 644 1516
rect 566 1513 573 1514
rect 566 1508 567 1513
rect 572 1508 573 1513
rect 604 1511 638 1515
rect 566 1507 573 1508
rect 603 1510 610 1511
rect 603 1505 604 1510
rect 609 1505 610 1510
rect 637 1510 638 1511
rect 643 1510 644 1515
rect 676 1515 712 1520
rect 818 1518 823 1571
rect 841 1570 848 1571
rect 899 1542 904 1630
rect 861 1537 904 1542
rect 637 1509 644 1510
rect 661 1510 668 1511
rect 603 1504 610 1505
rect 614 1506 621 1507
rect 614 1501 615 1506
rect 620 1501 621 1506
rect 661 1505 662 1510
rect 667 1505 668 1510
rect 676 1509 677 1515
rect 682 1514 712 1515
rect 682 1509 683 1514
rect 707 1511 712 1514
rect 817 1517 824 1518
rect 817 1512 818 1517
rect 823 1512 824 1517
rect 817 1511 824 1512
rect 676 1508 683 1509
rect 706 1510 713 1511
rect 706 1505 707 1510
rect 712 1505 713 1510
rect 735 1509 742 1510
rect 661 1504 668 1505
rect 690 1504 697 1505
rect 706 1504 713 1505
rect 719 1504 725 1505
rect 662 1501 667 1504
rect 614 1496 667 1501
rect 690 1499 691 1504
rect 696 1499 697 1504
rect 719 1499 720 1504
rect 724 1499 725 1504
rect 690 1498 725 1499
rect 691 1494 725 1498
rect 735 1504 736 1509
rect 741 1504 742 1509
rect 861 1504 866 1537
rect 924 1514 931 1515
rect 924 1509 925 1514
rect 930 1509 931 1514
rect 924 1508 931 1509
rect 735 1503 742 1504
rect 761 1503 768 1504
rect 735 1498 762 1503
rect 767 1498 768 1503
rect 861 1503 873 1504
rect 861 1498 867 1503
rect 872 1498 873 1503
rect 735 1477 740 1498
rect 761 1497 768 1498
rect 866 1497 873 1498
rect 568 1471 740 1477
rect 568 1451 573 1471
rect 567 1450 574 1451
rect 567 1445 568 1450
rect 573 1445 574 1450
rect 567 1444 574 1445
rect 614 1447 667 1452
rect 691 1450 725 1454
rect 603 1443 610 1444
rect 603 1438 604 1443
rect 609 1438 610 1443
rect 614 1442 615 1447
rect 620 1442 621 1447
rect 662 1444 667 1447
rect 690 1449 725 1450
rect 690 1444 691 1449
rect 696 1444 697 1449
rect 719 1444 720 1449
rect 724 1444 725 1449
rect 760 1445 767 1446
rect 866 1445 873 1446
rect 614 1441 621 1442
rect 661 1443 668 1444
rect 690 1443 697 1444
rect 706 1443 713 1444
rect 719 1443 725 1444
rect 735 1444 761 1445
rect 603 1437 610 1438
rect 637 1438 644 1439
rect 637 1437 638 1438
rect 604 1433 638 1437
rect 643 1433 644 1438
rect 661 1438 662 1443
rect 667 1438 668 1443
rect 661 1437 668 1438
rect 676 1439 683 1440
rect 604 1432 644 1433
rect 676 1433 677 1439
rect 682 1434 683 1439
rect 706 1438 707 1443
rect 712 1438 713 1443
rect 706 1437 713 1438
rect 735 1439 736 1444
rect 741 1440 761 1444
rect 766 1440 767 1445
rect 741 1439 742 1440
rect 760 1439 767 1440
rect 862 1440 867 1445
rect 872 1440 873 1445
rect 862 1439 873 1440
rect 735 1438 742 1439
rect 707 1434 712 1437
rect 682 1433 712 1434
rect 676 1428 712 1433
rect 735 1411 740 1438
rect 567 1405 740 1411
rect 862 1411 867 1439
rect 862 1406 905 1411
rect 567 1382 572 1405
rect 604 1383 644 1384
rect 566 1381 573 1382
rect 566 1376 567 1381
rect 572 1376 573 1381
rect 604 1379 638 1383
rect 566 1375 573 1376
rect 603 1378 610 1379
rect 603 1373 604 1378
rect 609 1373 610 1378
rect 637 1378 638 1379
rect 643 1378 644 1383
rect 676 1383 712 1388
rect 900 1387 905 1406
rect 637 1377 644 1378
rect 661 1378 668 1379
rect 603 1372 610 1373
rect 614 1374 621 1375
rect 614 1369 615 1374
rect 620 1369 621 1374
rect 661 1373 662 1378
rect 667 1373 668 1378
rect 676 1377 677 1383
rect 682 1382 712 1383
rect 682 1377 683 1382
rect 707 1379 712 1382
rect 899 1386 906 1387
rect 899 1381 900 1386
rect 905 1381 906 1386
rect 899 1380 906 1381
rect 925 1379 930 1508
rect 933 1379 940 1380
rect 676 1376 683 1377
rect 706 1378 713 1379
rect 706 1373 707 1378
rect 712 1373 713 1378
rect 735 1377 742 1378
rect 661 1372 668 1373
rect 690 1372 697 1373
rect 706 1372 713 1373
rect 719 1372 725 1373
rect 662 1369 667 1372
rect 614 1364 667 1369
rect 690 1367 691 1372
rect 696 1367 697 1372
rect 719 1367 720 1372
rect 724 1367 725 1372
rect 690 1366 725 1367
rect 691 1362 725 1366
rect 735 1372 736 1377
rect 741 1372 742 1377
rect 817 1377 824 1378
rect 817 1372 818 1377
rect 823 1372 824 1377
rect 913 1374 934 1379
rect 939 1374 940 1379
rect 913 1373 925 1374
rect 933 1373 940 1374
rect 735 1371 742 1372
rect 761 1371 768 1372
rect 817 1371 824 1372
rect 842 1371 849 1372
rect 735 1366 762 1371
rect 767 1366 768 1371
rect 818 1366 843 1371
rect 848 1366 849 1371
rect 735 1345 740 1366
rect 761 1365 768 1366
rect 842 1365 849 1366
rect 913 1365 918 1373
rect 568 1339 740 1345
rect 880 1344 918 1365
rect 568 1319 573 1339
rect 567 1318 574 1319
rect 567 1313 568 1318
rect 573 1313 574 1318
rect 567 1312 574 1313
rect 614 1315 667 1320
rect 691 1318 725 1322
rect 603 1311 610 1312
rect 603 1306 604 1311
rect 609 1306 610 1311
rect 614 1310 615 1315
rect 620 1310 621 1315
rect 662 1312 667 1315
rect 690 1317 725 1318
rect 690 1312 691 1317
rect 696 1312 697 1317
rect 719 1312 720 1317
rect 724 1312 725 1317
rect 614 1309 621 1310
rect 661 1311 668 1312
rect 690 1311 697 1312
rect 706 1311 713 1312
rect 719 1311 725 1312
rect 735 1312 742 1313
rect 603 1305 610 1306
rect 637 1306 644 1307
rect 637 1305 638 1306
rect 604 1301 638 1305
rect 643 1301 644 1306
rect 661 1306 662 1311
rect 667 1306 668 1311
rect 661 1305 668 1306
rect 676 1307 683 1308
rect 604 1300 644 1301
rect 676 1301 677 1307
rect 682 1302 683 1307
rect 706 1306 707 1311
rect 712 1306 713 1311
rect 735 1307 736 1312
rect 741 1310 742 1312
rect 761 1310 768 1311
rect 841 1310 848 1311
rect 741 1307 762 1310
rect 735 1306 762 1307
rect 706 1305 713 1306
rect 736 1305 762 1306
rect 767 1305 768 1310
rect 707 1302 712 1305
rect 682 1301 712 1302
rect 676 1296 712 1301
rect 736 1279 741 1305
rect 761 1304 768 1305
rect 818 1305 842 1310
rect 847 1305 848 1310
rect 567 1273 741 1279
rect 567 1250 572 1273
rect 604 1251 644 1252
rect 566 1249 573 1250
rect 566 1244 567 1249
rect 572 1244 573 1249
rect 604 1247 638 1251
rect 566 1243 573 1244
rect 603 1246 610 1247
rect 603 1241 604 1246
rect 609 1241 610 1246
rect 637 1246 638 1247
rect 643 1246 644 1251
rect 676 1251 712 1256
rect 818 1254 823 1305
rect 841 1304 848 1305
rect 637 1245 644 1246
rect 661 1246 668 1247
rect 603 1240 610 1241
rect 614 1242 621 1243
rect 614 1237 615 1242
rect 620 1237 621 1242
rect 661 1241 662 1246
rect 667 1241 668 1246
rect 676 1245 677 1251
rect 682 1250 712 1251
rect 682 1245 683 1250
rect 707 1247 712 1250
rect 817 1253 824 1254
rect 817 1248 818 1253
rect 823 1248 824 1253
rect 817 1247 824 1248
rect 676 1244 683 1245
rect 706 1246 713 1247
rect 706 1241 707 1246
rect 712 1241 713 1246
rect 735 1245 742 1246
rect 661 1240 668 1241
rect 690 1240 697 1241
rect 706 1240 713 1241
rect 719 1240 725 1241
rect 662 1237 667 1240
rect 614 1232 667 1237
rect 690 1235 691 1240
rect 696 1235 697 1240
rect 719 1235 720 1240
rect 724 1235 725 1240
rect 690 1234 725 1235
rect 691 1230 725 1234
rect 735 1240 736 1245
rect 741 1240 742 1245
rect 735 1239 742 1240
rect 761 1239 768 1240
rect 735 1234 762 1239
rect 767 1234 768 1239
rect 880 1235 885 1344
rect 930 1306 937 1307
rect 930 1301 931 1306
rect 936 1301 937 1306
rect 930 1300 937 1301
rect 837 1234 885 1235
rect 735 1213 740 1234
rect 761 1233 768 1234
rect 568 1207 740 1213
rect 806 1229 885 1234
rect 931 1238 936 1300
rect 931 1232 998 1238
rect 568 1187 573 1207
rect 567 1186 574 1187
rect 567 1181 568 1186
rect 573 1181 574 1186
rect 567 1180 574 1181
rect 614 1183 667 1188
rect 691 1186 725 1190
rect 806 1186 811 1229
rect 603 1179 610 1180
rect 603 1174 604 1179
rect 609 1174 610 1179
rect 614 1178 615 1183
rect 620 1178 621 1183
rect 662 1180 667 1183
rect 690 1185 725 1186
rect 690 1180 691 1185
rect 696 1180 697 1185
rect 719 1180 720 1185
rect 724 1180 725 1185
rect 805 1185 812 1186
rect 614 1177 621 1178
rect 661 1179 668 1180
rect 690 1179 697 1180
rect 706 1179 713 1180
rect 719 1179 725 1180
rect 735 1180 742 1181
rect 603 1173 610 1174
rect 637 1174 644 1175
rect 637 1173 638 1174
rect 604 1169 638 1173
rect 643 1169 644 1174
rect 661 1174 662 1179
rect 667 1174 668 1179
rect 661 1173 668 1174
rect 676 1175 683 1176
rect 604 1168 644 1169
rect 676 1169 677 1175
rect 682 1170 683 1175
rect 706 1174 707 1179
rect 712 1174 713 1179
rect 735 1175 736 1180
rect 741 1175 742 1180
rect 805 1180 806 1185
rect 811 1180 812 1185
rect 875 1183 928 1188
rect 952 1186 986 1190
rect 993 1186 998 1232
rect 805 1179 812 1180
rect 864 1179 871 1180
rect 735 1174 742 1175
rect 760 1174 767 1175
rect 706 1173 713 1174
rect 707 1170 712 1173
rect 682 1169 712 1170
rect 737 1169 761 1174
rect 766 1169 767 1174
rect 864 1174 865 1179
rect 870 1174 871 1179
rect 875 1178 876 1183
rect 881 1178 882 1183
rect 923 1180 928 1183
rect 951 1185 986 1186
rect 951 1180 952 1185
rect 957 1180 958 1185
rect 980 1180 981 1185
rect 985 1180 986 1185
rect 875 1177 882 1178
rect 922 1179 929 1180
rect 951 1179 958 1180
rect 967 1179 974 1180
rect 980 1179 986 1180
rect 992 1185 999 1186
rect 992 1180 993 1185
rect 998 1180 999 1185
rect 992 1179 999 1180
rect 864 1173 871 1174
rect 898 1174 905 1175
rect 898 1173 899 1174
rect 676 1164 712 1169
rect 760 1168 767 1169
rect 865 1169 899 1173
rect 904 1169 905 1174
rect 922 1174 923 1179
rect 928 1174 929 1179
rect 922 1173 929 1174
rect 937 1175 944 1176
rect 865 1168 905 1169
rect 937 1169 938 1175
rect 943 1170 944 1175
rect 967 1174 968 1179
rect 973 1174 974 1179
rect 967 1173 974 1174
rect 968 1170 973 1173
rect 943 1169 973 1170
rect 937 1164 973 1169
rect 1020 1141 1025 1668
rect 867 1136 1025 1141
rect 867 1076 872 1136
rect 866 1075 872 1076
rect 866 1071 867 1075
rect 871 1071 872 1075
rect 866 1070 872 1071
rect 992 1008 1026 1013
rect 992 994 997 1008
rect 991 993 997 994
rect 991 989 992 993
rect 996 989 997 993
rect 991 988 997 989
rect 484 820 490 821
rect 484 816 485 820
rect 489 816 490 820
rect 484 815 490 816
rect 96 779 1026 784
<< labels >>
rlabel metal2 544 782 544 782 5 p_clk_b
rlabel metal2 556 782 556 782 5 p_clk
rlabel metal2 532 781 532 781 5 f_clk
rlabel metal2 520 782 520 782 4 f_clk_b
rlabel metal2 495 783 495 783 1 Vdd!
rlabel metal2 507 783 507 783 1 GND!
rlabel metal2 507 1763 507 1763 1 GND!
rlabel metal2 495 1763 495 1763 1 Vdd!
rlabel polysilicon 1007 1130 1007 1130 1 CB3
rlabel polysilicon 1019 986 1019 986 1 CB4
rlabel polysilicon 241 1633 241 1633 1 CB1
rlabel polysilicon 358 1641 358 1641 1 CB2
rlabel metal2 520 1762 520 1762 4 f_clk_b
rlabel metal2 532 1761 532 1761 5 f_clk
rlabel metal2 556 1762 556 1762 5 p_clk
rlabel metal2 544 1762 544 1762 5 p_clk_b
rlabel metal2 885 1674 888 1680 1 select2
rlabel metal2 825 1674 828 1681 1 select1
rlabel metal2 742 1675 745 1680 1 select0
rlabel metal2 913 1665 916 1670 1 select_out
rlabel metal1 918 1509 921 1512 7 Y
rlabel polysilicon 830 1181 832 1184 5 reset
rlabel polysilicon 353 877 353 877 1 11
rlabel polysilicon 358 865 358 865 1 10
rlabel polysilicon 334 866 334 866 1 9
rlabel polysilicon 239 1103 239 1103 1 5
rlabel polysilicon 241 1092 241 1092 1 4
rlabel polysilicon 217 1092 217 1092 1 3
rlabel polysilicon 354 889 354 889 1 8
rlabel polysilicon 358 907 358 907 1 7
rlabel polysilicon 334 907 334 907 1 6
rlabel polysilicon 237 1121 237 1121 1 2
rlabel polysilicon 241 1132 241 1132 1 1
rlabel polysilicon 217 1132 217 1132 1 0
rlabel metal2 228 1749 228 1749 1 A
rlabel metal2 346 1745 346 1745 1 B
rlabel metal1 1023 1118 1023 1118 1 C
rlabel m3contact 97 1182 97 1182 1 in
rlabel metal1 1021 892 1021 892 1 E
rlabel metal1 570 1638 570 1638 1 LB_in
rlabel metal1 995 1379 995 1379 1 LB_out
<< end >>
