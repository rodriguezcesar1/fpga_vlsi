magic
tech scmos
timestamp 1607749837
<< ntransistor >>
rect 12 24 14 28
rect 28 24 30 28
rect 47 24 49 28
rect 70 24 72 28
rect 75 24 77 28
rect 101 24 103 28
rect 129 24 131 28
rect 149 24 151 28
rect 154 24 156 28
rect 181 24 183 28
rect 197 24 199 28
rect 213 24 215 28
rect 232 24 234 28
rect 255 24 257 28
rect 260 24 262 28
rect 286 24 288 28
rect 314 24 316 28
rect 334 24 336 28
rect 339 24 341 28
rect 366 24 368 28
rect 382 24 384 28
rect 398 24 400 28
rect 417 24 419 28
rect 440 24 442 28
rect 445 24 447 28
rect 471 24 473 28
rect 499 24 501 28
rect 519 24 521 28
rect 524 24 526 28
rect 551 24 553 28
rect 567 24 569 28
rect 583 24 585 28
rect 602 24 604 28
rect 625 24 627 28
rect 630 24 632 28
rect 656 24 658 28
rect 684 24 686 28
rect 704 24 706 28
rect 709 24 711 28
rect 736 24 738 28
<< ptransistor >>
rect 12 43 14 51
rect 28 43 30 51
rect 47 44 49 52
rect 70 43 72 51
rect 75 43 77 51
rect 101 43 103 51
rect 129 44 131 52
rect 149 43 151 51
rect 154 43 156 51
rect 181 43 183 51
rect 197 43 199 51
rect 213 43 215 51
rect 232 44 234 52
rect 255 43 257 51
rect 260 43 262 51
rect 286 43 288 51
rect 314 44 316 52
rect 334 43 336 51
rect 339 43 341 51
rect 366 43 368 51
rect 382 43 384 51
rect 398 43 400 51
rect 417 44 419 52
rect 440 43 442 51
rect 445 43 447 51
rect 471 43 473 51
rect 499 44 501 52
rect 519 43 521 51
rect 524 43 526 51
rect 551 43 553 51
rect 567 43 569 51
rect 583 43 585 51
rect 602 44 604 52
rect 625 43 627 51
rect 630 43 632 51
rect 656 43 658 51
rect 684 44 686 52
rect 704 43 706 51
rect 709 43 711 51
rect 736 43 738 51
<< ndiffusion >>
rect 11 24 12 28
rect 14 24 15 28
rect 27 24 28 28
rect 30 24 31 28
rect 46 24 47 28
rect 49 24 50 28
rect 65 24 70 28
rect 72 24 75 28
rect 77 24 78 28
rect 99 24 101 28
rect 103 24 104 28
rect 128 24 129 28
rect 131 24 132 28
rect 144 24 149 28
rect 151 24 154 28
rect 156 24 157 28
rect 180 24 181 28
rect 183 24 184 28
rect 196 24 197 28
rect 199 24 200 28
rect 212 24 213 28
rect 215 24 216 28
rect 231 24 232 28
rect 234 24 235 28
rect 250 24 255 28
rect 257 24 260 28
rect 262 24 263 28
rect 284 24 286 28
rect 288 24 289 28
rect 313 24 314 28
rect 316 24 317 28
rect 329 24 334 28
rect 336 24 339 28
rect 341 24 342 28
rect 365 24 366 28
rect 368 24 369 28
rect 381 24 382 28
rect 384 24 385 28
rect 397 24 398 28
rect 400 24 401 28
rect 416 24 417 28
rect 419 24 420 28
rect 435 24 440 28
rect 442 24 445 28
rect 447 24 448 28
rect 469 24 471 28
rect 473 24 474 28
rect 498 24 499 28
rect 501 24 502 28
rect 514 24 519 28
rect 521 24 524 28
rect 526 24 527 28
rect 550 24 551 28
rect 553 24 554 28
rect 566 24 567 28
rect 569 24 570 28
rect 582 24 583 28
rect 585 24 586 28
rect 601 24 602 28
rect 604 24 605 28
rect 620 24 625 28
rect 627 24 630 28
rect 632 24 633 28
rect 654 24 656 28
rect 658 24 659 28
rect 683 24 684 28
rect 686 24 687 28
rect 699 24 704 28
rect 706 24 709 28
rect 711 24 712 28
rect 735 24 736 28
rect 738 24 739 28
<< pdiffusion >>
rect 11 43 12 51
rect 14 43 15 51
rect 27 43 28 51
rect 30 43 31 51
rect 46 44 47 52
rect 49 44 50 52
rect 65 43 70 51
rect 72 43 75 51
rect 77 43 78 51
rect 99 43 101 51
rect 103 43 104 51
rect 128 44 129 52
rect 131 44 132 52
rect 144 43 149 51
rect 151 43 154 51
rect 156 43 157 51
rect 180 43 181 51
rect 183 43 184 51
rect 196 43 197 51
rect 199 43 200 51
rect 212 43 213 51
rect 215 43 216 51
rect 231 44 232 52
rect 234 44 235 52
rect 250 43 255 51
rect 257 43 260 51
rect 262 43 263 51
rect 284 43 286 51
rect 288 43 289 51
rect 313 44 314 52
rect 316 44 317 52
rect 329 43 334 51
rect 336 43 339 51
rect 341 43 342 51
rect 365 43 366 51
rect 368 43 369 51
rect 381 43 382 51
rect 384 43 385 51
rect 397 43 398 51
rect 400 43 401 51
rect 416 44 417 52
rect 419 44 420 52
rect 435 43 440 51
rect 442 43 445 51
rect 447 43 448 51
rect 469 43 471 51
rect 473 43 474 51
rect 498 44 499 52
rect 501 44 502 52
rect 514 43 519 51
rect 521 43 524 51
rect 526 43 527 51
rect 550 43 551 51
rect 553 43 554 51
rect 566 43 567 51
rect 569 43 570 51
rect 582 43 583 51
rect 585 43 586 51
rect 601 44 602 52
rect 604 44 605 52
rect 620 43 625 51
rect 627 43 630 51
rect 632 43 633 51
rect 654 43 656 51
rect 658 43 659 51
rect 683 44 684 52
rect 686 44 687 52
rect 699 43 704 51
rect 706 43 709 51
rect 711 43 712 51
rect 735 43 736 51
rect 738 43 739 51
<< ndcontact >>
rect 7 24 11 28
rect 15 24 19 28
rect 23 24 27 28
rect 31 24 35 28
rect 42 24 46 28
rect 50 24 54 28
rect 61 24 65 28
rect 78 24 82 28
rect 95 24 99 28
rect 104 24 108 28
rect 124 24 128 28
rect 132 24 136 28
rect 140 24 144 28
rect 157 24 161 28
rect 176 24 180 28
rect 184 24 188 28
rect 192 24 196 28
rect 200 24 204 28
rect 208 24 212 28
rect 216 24 220 28
rect 227 24 231 28
rect 235 24 239 28
rect 246 24 250 28
rect 263 24 267 28
rect 280 24 284 28
rect 289 24 293 28
rect 309 24 313 28
rect 317 24 321 28
rect 325 24 329 28
rect 342 24 346 28
rect 361 24 365 28
rect 369 24 373 28
rect 377 24 381 28
rect 385 24 389 28
rect 393 24 397 28
rect 401 24 405 28
rect 412 24 416 28
rect 420 24 424 28
rect 431 24 435 28
rect 448 24 452 28
rect 465 24 469 28
rect 474 24 478 28
rect 494 24 498 28
rect 502 24 506 28
rect 510 24 514 28
rect 527 24 531 28
rect 546 24 550 28
rect 554 24 558 28
rect 562 24 566 28
rect 570 24 574 28
rect 578 24 582 28
rect 586 24 590 28
rect 597 24 601 28
rect 605 24 609 28
rect 616 24 620 28
rect 633 24 637 28
rect 650 24 654 28
rect 659 24 663 28
rect 679 24 683 28
rect 687 24 691 28
rect 695 24 699 28
rect 712 24 716 28
rect 731 24 735 28
rect 739 24 743 28
<< pdcontact >>
rect 7 43 11 51
rect 15 43 19 51
rect 23 43 27 51
rect 31 43 35 51
rect 42 44 46 52
rect 50 44 54 52
rect 61 43 65 51
rect 78 43 82 51
rect 95 43 99 51
rect 104 43 108 51
rect 124 44 128 52
rect 132 44 136 52
rect 140 43 144 51
rect 157 43 161 51
rect 176 43 180 51
rect 184 43 188 51
rect 192 43 196 51
rect 200 43 204 51
rect 208 43 212 51
rect 216 43 220 51
rect 227 44 231 52
rect 235 44 239 52
rect 246 43 250 51
rect 263 43 267 51
rect 280 43 284 51
rect 289 43 293 51
rect 309 44 313 52
rect 317 44 321 52
rect 325 43 329 51
rect 342 43 346 51
rect 361 43 365 51
rect 369 43 373 51
rect 377 43 381 51
rect 385 43 389 51
rect 393 43 397 51
rect 401 43 405 51
rect 412 44 416 52
rect 420 44 424 52
rect 431 43 435 51
rect 448 43 452 51
rect 465 43 469 51
rect 474 43 478 51
rect 494 44 498 52
rect 502 44 506 52
rect 510 43 514 51
rect 527 43 531 51
rect 546 43 550 51
rect 554 43 558 51
rect 562 43 566 51
rect 570 43 574 51
rect 578 43 582 51
rect 586 43 590 51
rect 597 44 601 52
rect 605 44 609 52
rect 616 43 620 51
rect 633 43 637 51
rect 650 43 654 51
rect 659 43 663 51
rect 679 44 683 52
rect 687 44 691 52
rect 695 43 699 51
rect 712 43 716 51
rect 731 43 735 51
rect 739 43 743 51
<< psubstratepcontact >>
rect 0 8 4 12
rect 18 8 22 12
rect 38 8 42 12
rect 51 8 55 12
rect 87 8 91 12
rect 113 8 117 12
rect 133 8 137 12
rect 185 8 189 12
rect 203 8 207 12
rect 223 8 227 12
rect 236 8 240 12
rect 272 8 276 12
rect 298 8 302 12
rect 318 8 322 12
rect 370 8 374 12
rect 388 8 392 12
rect 408 8 412 12
rect 421 8 425 12
rect 457 8 461 12
rect 483 8 487 12
rect 503 8 507 12
rect 555 8 559 12
rect 573 8 577 12
rect 593 8 597 12
rect 606 8 610 12
rect 642 8 646 12
rect 668 8 672 12
rect 688 8 692 12
<< nsubstratencontact >>
rect 0 61 4 65
rect 18 61 22 65
rect 38 61 42 65
rect 51 61 55 65
rect 87 61 91 65
rect 113 61 117 65
rect 133 61 137 65
rect 185 61 189 65
rect 203 61 207 65
rect 223 61 227 65
rect 236 61 240 65
rect 272 61 276 65
rect 298 61 302 65
rect 318 61 322 65
rect 370 61 374 65
rect 388 61 392 65
rect 408 61 412 65
rect 421 61 425 65
rect 457 61 461 65
rect 483 61 487 65
rect 503 61 507 65
rect 555 61 559 65
rect 573 61 577 65
rect 593 61 597 65
rect 606 61 610 65
rect 642 61 646 65
rect 668 61 672 65
rect 688 61 692 65
<< polysilicon >>
rect 28 58 30 61
rect 75 58 77 61
rect 101 58 103 61
rect 154 58 156 61
rect 213 58 215 61
rect 260 58 262 61
rect 286 58 288 61
rect 339 58 341 61
rect 398 58 400 61
rect 445 58 447 61
rect 471 58 473 61
rect 524 58 526 61
rect 583 58 585 61
rect 630 58 632 61
rect 656 58 658 61
rect 709 58 711 61
rect 28 54 29 58
rect 101 54 102 58
rect 213 54 214 58
rect 286 54 287 58
rect 398 54 399 58
rect 471 54 472 58
rect 583 54 584 58
rect 656 54 657 58
rect 12 51 14 53
rect 28 51 30 54
rect 47 52 49 54
rect 70 51 72 53
rect 75 51 77 54
rect 101 51 103 54
rect 129 52 131 54
rect 12 28 14 43
rect 28 41 30 43
rect 28 28 30 30
rect 47 28 49 44
rect 149 51 151 53
rect 154 51 156 54
rect 181 51 183 53
rect 197 51 199 53
rect 213 51 215 54
rect 232 52 234 54
rect 70 37 72 43
rect 75 41 77 43
rect 101 41 103 43
rect 66 33 72 37
rect 70 28 72 33
rect 75 28 77 30
rect 101 28 103 30
rect 129 28 131 44
rect 255 51 257 53
rect 260 51 262 54
rect 286 51 288 54
rect 314 52 316 54
rect 149 37 151 43
rect 154 41 156 43
rect 145 33 151 37
rect 149 28 151 33
rect 154 28 156 30
rect 181 28 183 43
rect 197 28 199 43
rect 213 41 215 43
rect 213 28 215 30
rect 232 28 234 44
rect 334 51 336 53
rect 339 51 341 54
rect 366 51 368 53
rect 382 51 384 53
rect 398 51 400 54
rect 417 52 419 54
rect 255 37 257 43
rect 260 41 262 43
rect 286 41 288 43
rect 251 33 257 37
rect 255 28 257 33
rect 260 28 262 30
rect 286 28 288 30
rect 314 28 316 44
rect 440 51 442 53
rect 445 51 447 54
rect 471 51 473 54
rect 499 52 501 54
rect 334 37 336 43
rect 339 41 341 43
rect 330 33 336 37
rect 334 28 336 33
rect 339 28 341 30
rect 366 28 368 43
rect 382 28 384 43
rect 398 41 400 43
rect 398 28 400 30
rect 417 28 419 44
rect 519 51 521 53
rect 524 51 526 54
rect 551 51 553 53
rect 567 51 569 53
rect 583 51 585 54
rect 602 52 604 54
rect 440 37 442 43
rect 445 41 447 43
rect 471 41 473 43
rect 436 33 442 37
rect 440 28 442 33
rect 445 28 447 30
rect 471 28 473 30
rect 499 28 501 44
rect 625 51 627 53
rect 630 51 632 54
rect 656 51 658 54
rect 684 52 686 54
rect 519 37 521 43
rect 524 41 526 43
rect 515 33 521 37
rect 519 28 521 33
rect 524 28 526 30
rect 551 28 553 43
rect 567 28 569 43
rect 583 41 585 43
rect 583 28 585 30
rect 602 28 604 44
rect 704 51 706 53
rect 709 51 711 54
rect 736 51 738 53
rect 625 37 627 43
rect 630 41 632 43
rect 656 41 658 43
rect 621 33 627 37
rect 625 28 627 33
rect 630 28 632 30
rect 656 28 658 30
rect 684 28 686 44
rect 704 37 706 43
rect 709 41 711 43
rect 700 33 706 37
rect 704 28 706 33
rect 709 28 711 30
rect 736 28 738 43
rect 12 22 14 24
rect 28 20 30 24
rect 47 22 49 24
rect 70 22 72 24
rect 29 16 30 20
rect 75 19 77 24
rect 101 20 103 24
rect 129 22 131 24
rect 149 22 151 24
rect 28 13 30 16
rect 76 15 77 19
rect 102 16 103 20
rect 154 19 156 24
rect 181 22 183 24
rect 197 22 199 24
rect 213 20 215 24
rect 232 22 234 24
rect 255 22 257 24
rect 75 13 77 15
rect 101 12 103 16
rect 155 15 156 19
rect 214 16 215 20
rect 260 19 262 24
rect 286 20 288 24
rect 314 22 316 24
rect 334 22 336 24
rect 154 13 156 15
rect 213 13 215 16
rect 261 15 262 19
rect 287 16 288 20
rect 339 19 341 24
rect 366 22 368 24
rect 382 22 384 24
rect 398 20 400 24
rect 417 22 419 24
rect 440 22 442 24
rect 260 13 262 15
rect 286 12 288 16
rect 340 15 341 19
rect 399 16 400 20
rect 445 19 447 24
rect 471 20 473 24
rect 499 22 501 24
rect 519 22 521 24
rect 339 13 341 15
rect 398 13 400 16
rect 446 15 447 19
rect 472 16 473 20
rect 524 19 526 24
rect 551 22 553 24
rect 567 22 569 24
rect 583 20 585 24
rect 602 22 604 24
rect 625 22 627 24
rect 445 13 447 15
rect 471 12 473 16
rect 525 15 526 19
rect 584 16 585 20
rect 630 19 632 24
rect 656 20 658 24
rect 684 22 686 24
rect 704 22 706 24
rect 524 13 526 15
rect 583 13 585 16
rect 631 15 632 19
rect 657 16 658 20
rect 709 19 711 24
rect 736 22 738 24
rect 630 13 632 15
rect 656 12 658 16
rect 710 15 711 19
rect 709 13 711 15
<< polycontact >>
rect 29 54 33 58
rect 75 54 79 58
rect 102 54 106 58
rect 154 54 158 58
rect 214 54 218 58
rect 260 54 264 58
rect 287 54 291 58
rect 339 54 343 58
rect 399 54 403 58
rect 445 54 449 58
rect 472 54 476 58
rect 524 54 528 58
rect 584 54 588 58
rect 630 54 634 58
rect 657 54 661 58
rect 709 54 713 58
rect 8 33 12 37
rect 43 34 47 38
rect 62 33 66 37
rect 125 34 129 38
rect 141 33 145 37
rect 177 33 181 37
rect 193 33 197 37
rect 228 34 232 38
rect 247 33 251 37
rect 310 34 314 38
rect 326 33 330 37
rect 362 33 366 37
rect 378 33 382 37
rect 413 34 417 38
rect 432 33 436 37
rect 495 34 499 38
rect 511 33 515 37
rect 547 33 551 37
rect 563 33 567 37
rect 598 34 602 38
rect 617 33 621 37
rect 680 34 684 38
rect 696 33 700 37
rect 732 33 736 37
rect 25 16 29 20
rect 72 15 76 19
rect 97 16 102 20
rect 151 15 155 19
rect 210 16 214 20
rect 257 15 261 19
rect 282 16 287 20
rect 336 15 340 19
rect 395 16 399 20
rect 442 15 446 19
rect 467 16 472 20
rect 521 15 525 19
rect 580 16 584 20
rect 627 15 631 19
rect 652 16 657 20
rect 706 15 710 19
<< metal1 >>
rect 0 70 34 74
rect 38 70 64 74
rect 68 70 89 74
rect 93 70 164 74
rect 168 70 219 74
rect 223 70 249 74
rect 253 70 274 74
rect 278 70 349 74
rect 353 70 404 74
rect 408 70 434 74
rect 438 70 459 74
rect 463 70 534 74
rect 538 70 589 74
rect 593 70 619 74
rect 623 70 644 74
rect 648 70 719 74
rect 723 70 743 74
rect 4 61 18 65
rect 22 61 38 65
rect 42 61 51 65
rect 55 61 87 65
rect 91 61 113 65
rect 117 61 133 65
rect 137 61 185 65
rect 189 61 203 65
rect 207 61 223 65
rect 227 61 236 65
rect 240 61 272 65
rect 276 61 298 65
rect 302 61 318 65
rect 322 61 370 65
rect 374 61 388 65
rect 392 61 408 65
rect 412 61 421 65
rect 425 61 457 65
rect 461 61 483 65
rect 487 61 503 65
rect 507 61 555 65
rect 559 61 573 65
rect 577 61 593 65
rect 597 61 606 65
rect 610 61 642 65
rect 646 61 668 65
rect 672 61 688 65
rect 692 61 743 65
rect 7 51 10 61
rect 33 54 34 58
rect 42 52 45 61
rect 3 33 8 36
rect 16 36 19 43
rect 23 36 26 43
rect 16 33 26 36
rect 16 28 19 33
rect 23 28 26 33
rect 32 38 35 43
rect 32 36 38 38
rect 42 36 43 38
rect 32 34 43 36
rect 51 37 54 44
rect 61 51 64 61
rect 79 54 82 58
rect 106 54 107 58
rect 124 52 127 61
rect 79 39 82 43
rect 51 35 62 37
rect 32 28 35 34
rect 51 33 57 35
rect 51 28 54 33
rect 61 33 62 35
rect 80 35 82 39
rect 79 28 82 35
rect 95 38 98 43
rect 105 38 108 43
rect 105 34 117 38
rect 121 34 125 38
rect 133 37 136 44
rect 140 51 143 61
rect 158 54 164 58
rect 176 51 179 61
rect 192 51 195 61
rect 218 54 219 58
rect 227 52 230 61
rect 158 38 161 43
rect 95 28 98 34
rect 105 28 108 34
rect 133 33 134 37
rect 138 33 141 36
rect 160 34 161 38
rect 133 28 136 33
rect 158 28 161 34
rect 173 33 177 37
rect 185 36 188 43
rect 185 33 193 36
rect 201 36 204 43
rect 208 36 211 43
rect 201 33 211 36
rect 185 28 188 33
rect 201 28 204 33
rect 208 28 211 33
rect 217 38 220 43
rect 217 36 223 38
rect 227 36 228 38
rect 217 34 228 36
rect 236 37 239 44
rect 246 51 249 61
rect 264 54 267 58
rect 291 54 292 58
rect 309 52 312 61
rect 264 39 267 43
rect 236 35 247 37
rect 217 28 220 34
rect 236 33 242 35
rect 236 28 239 33
rect 246 33 247 35
rect 265 35 267 39
rect 264 28 267 35
rect 280 38 283 43
rect 290 38 293 43
rect 290 34 302 38
rect 306 34 310 38
rect 318 37 321 44
rect 325 51 328 61
rect 343 54 349 58
rect 361 51 364 61
rect 377 51 380 61
rect 403 54 404 58
rect 412 52 415 61
rect 343 38 346 43
rect 280 28 283 34
rect 290 28 293 34
rect 318 33 319 37
rect 323 33 326 36
rect 345 34 346 38
rect 318 28 321 33
rect 343 28 346 34
rect 358 33 362 37
rect 370 36 373 43
rect 370 33 378 36
rect 386 36 389 43
rect 393 36 396 43
rect 386 33 396 36
rect 370 28 373 33
rect 386 28 389 33
rect 393 28 396 33
rect 402 38 405 43
rect 402 36 408 38
rect 412 36 413 38
rect 402 34 413 36
rect 421 37 424 44
rect 431 51 434 61
rect 449 54 452 58
rect 476 54 477 58
rect 494 52 497 61
rect 449 39 452 43
rect 421 35 432 37
rect 402 28 405 34
rect 421 33 427 35
rect 421 28 424 33
rect 431 33 432 35
rect 450 35 452 39
rect 449 28 452 35
rect 465 38 468 43
rect 475 38 478 43
rect 475 34 487 38
rect 491 34 495 38
rect 503 37 506 44
rect 510 51 513 61
rect 528 54 534 58
rect 546 51 549 61
rect 562 51 565 61
rect 588 54 589 58
rect 597 52 600 61
rect 528 38 531 43
rect 465 28 468 34
rect 475 28 478 34
rect 503 33 504 37
rect 508 33 511 36
rect 530 34 531 38
rect 503 28 506 33
rect 528 28 531 34
rect 543 33 547 37
rect 555 36 558 43
rect 555 33 563 36
rect 571 36 574 43
rect 578 36 581 43
rect 571 33 581 36
rect 555 28 558 33
rect 571 28 574 33
rect 578 28 581 33
rect 587 38 590 43
rect 587 36 593 38
rect 597 36 598 38
rect 587 34 598 36
rect 606 37 609 44
rect 616 51 619 61
rect 634 54 637 58
rect 661 54 662 58
rect 679 52 682 61
rect 634 39 637 43
rect 606 35 617 37
rect 587 28 590 34
rect 606 33 612 35
rect 606 28 609 33
rect 616 33 617 35
rect 635 35 637 39
rect 634 28 637 35
rect 650 38 653 43
rect 660 38 663 43
rect 660 34 672 38
rect 676 34 680 38
rect 688 37 691 44
rect 695 51 698 61
rect 713 54 719 58
rect 731 51 734 61
rect 713 38 716 43
rect 650 28 653 34
rect 660 28 663 34
rect 688 33 689 37
rect 693 33 696 36
rect 715 34 716 38
rect 688 28 691 33
rect 713 28 716 34
rect 728 33 732 37
rect 740 28 743 43
rect 7 12 10 24
rect 24 16 25 20
rect 42 12 45 24
rect 61 12 64 24
rect 71 15 72 19
rect 96 16 97 20
rect 124 12 127 24
rect 140 12 143 24
rect 150 15 151 19
rect 176 12 179 24
rect 192 12 195 24
rect 209 16 210 20
rect 227 12 230 24
rect 246 12 249 24
rect 256 15 257 19
rect 281 16 282 20
rect 309 12 312 24
rect 325 12 328 24
rect 335 15 336 19
rect 361 12 364 24
rect 377 12 380 24
rect 394 16 395 20
rect 412 12 415 24
rect 431 12 434 24
rect 441 15 442 19
rect 466 16 467 20
rect 494 12 497 24
rect 510 12 513 24
rect 520 15 521 19
rect 546 12 549 24
rect 562 12 565 24
rect 579 16 580 20
rect 597 12 600 24
rect 616 12 619 24
rect 626 15 627 19
rect 651 16 652 20
rect 679 12 682 24
rect 695 12 698 24
rect 705 15 706 19
rect 731 12 734 24
rect 4 8 18 12
rect 22 8 38 12
rect 42 8 51 12
rect 55 8 87 12
rect 91 8 113 12
rect 117 8 133 12
rect 137 8 185 12
rect 189 8 203 12
rect 207 8 223 12
rect 227 8 236 12
rect 240 8 272 12
rect 276 8 298 12
rect 302 8 318 12
rect 322 8 370 12
rect 374 8 388 12
rect 392 8 408 12
rect 412 8 421 12
rect 425 8 457 12
rect 461 8 483 12
rect 487 8 503 12
rect 507 8 555 12
rect 559 8 573 12
rect 577 8 593 12
rect 597 8 606 12
rect 610 8 642 12
rect 646 8 668 12
rect 672 8 688 12
rect 692 8 743 12
rect 0 0 20 4
rect 24 0 83 4
rect 87 0 108 4
rect 112 0 146 4
rect 150 0 205 4
rect 209 0 268 4
rect 272 0 293 4
rect 297 0 331 4
rect 335 0 390 4
rect 394 0 453 4
rect 457 0 478 4
rect 482 0 516 4
rect 520 0 575 4
rect 579 0 638 4
rect 642 0 663 4
rect 667 0 701 4
rect 705 0 743 4
<< m2contact >>
rect 34 70 38 74
rect 64 70 68 74
rect 89 70 93 74
rect 164 70 168 74
rect 219 70 223 74
rect 249 70 253 74
rect 274 70 278 74
rect 349 70 353 74
rect 404 70 408 74
rect 434 70 438 74
rect 459 70 463 74
rect 534 70 538 74
rect 589 70 593 74
rect 619 70 623 74
rect 644 70 648 74
rect 719 70 723 74
rect 34 54 38 58
rect 38 36 42 40
rect 82 54 86 58
rect 107 54 111 58
rect 57 31 61 35
rect 76 35 80 39
rect 95 34 99 38
rect 117 34 121 38
rect 164 54 168 58
rect 219 54 223 58
rect 134 33 138 37
rect 156 34 160 38
rect 169 33 173 37
rect 223 36 227 40
rect 267 54 271 58
rect 292 54 296 58
rect 242 31 246 35
rect 261 35 265 39
rect 280 34 284 38
rect 302 34 306 38
rect 349 54 353 58
rect 404 54 408 58
rect 319 33 323 37
rect 341 34 345 38
rect 354 33 358 37
rect 408 36 412 40
rect 452 54 456 58
rect 477 54 481 58
rect 427 31 431 35
rect 446 35 450 39
rect 465 34 469 38
rect 487 34 491 38
rect 534 54 538 58
rect 589 54 593 58
rect 504 33 508 37
rect 526 34 530 38
rect 539 33 543 37
rect 593 36 597 40
rect 637 54 641 58
rect 662 54 666 58
rect 612 31 616 35
rect 631 35 635 39
rect 650 34 654 38
rect 672 34 676 38
rect 719 54 723 58
rect 689 33 693 37
rect 711 34 715 38
rect 724 33 728 37
rect 20 16 24 20
rect 67 15 71 19
rect 89 16 96 20
rect 146 15 150 19
rect 205 16 209 20
rect 252 15 256 19
rect 274 16 281 20
rect 331 15 335 19
rect 390 16 394 20
rect 437 15 441 19
rect 459 16 466 20
rect 516 15 520 19
rect 575 16 579 20
rect 622 15 626 19
rect 644 16 651 20
rect 701 15 705 19
rect 20 0 24 4
rect 83 0 87 4
rect 108 0 112 4
rect 146 0 150 4
rect 205 0 209 4
rect 268 0 272 4
rect 293 0 297 4
rect 331 0 335 4
rect 390 0 394 4
rect 453 0 457 4
rect 478 0 482 4
rect 516 0 520 4
rect 575 0 579 4
rect 638 0 642 4
rect 663 0 667 4
rect 701 0 705 4
<< metal2 >>
rect 34 58 38 70
rect 20 4 24 16
rect 64 15 67 70
rect 83 4 86 54
rect 89 20 92 70
rect 164 58 168 70
rect 219 58 223 70
rect 108 4 111 54
rect 146 4 150 15
rect 205 4 209 16
rect 249 15 252 70
rect 268 4 271 54
rect 274 20 277 70
rect 349 58 353 70
rect 404 58 408 70
rect 293 4 296 54
rect 331 4 335 15
rect 390 4 394 16
rect 434 15 437 70
rect 453 4 456 54
rect 459 20 462 70
rect 534 58 538 70
rect 589 58 593 70
rect 478 4 481 54
rect 516 4 520 15
rect 575 4 579 16
rect 619 15 622 70
rect 638 4 641 54
rect 644 20 647 70
rect 719 58 723 70
rect 663 4 666 54
rect 701 4 705 15
<< m3contact >>
rect 42 35 47 40
rect 56 26 61 31
rect 71 34 76 39
rect 99 34 104 39
rect 117 38 122 43
rect 151 34 156 39
rect 227 35 232 40
rect 135 28 140 33
rect 168 28 173 33
rect 241 26 246 31
rect 256 34 261 39
rect 284 34 289 39
rect 302 38 307 43
rect 336 34 341 39
rect 412 35 417 40
rect 320 28 325 33
rect 353 28 358 33
rect 426 26 431 31
rect 441 34 446 39
rect 469 34 474 39
rect 487 38 492 43
rect 521 34 526 39
rect 597 35 602 40
rect 505 28 510 33
rect 538 28 543 33
rect 611 26 616 31
rect 626 34 631 39
rect 654 34 659 39
rect 672 38 677 43
rect 706 34 711 39
rect 690 28 695 33
rect 723 28 728 33
<< metal3 >>
rect 117 45 156 50
rect 302 45 341 50
rect 487 45 526 50
rect 672 45 711 50
rect 42 41 76 45
rect 117 44 126 45
rect 134 44 156 45
rect 41 40 76 41
rect 116 43 123 44
rect 41 35 42 40
rect 47 35 48 40
rect 41 34 48 35
rect 70 39 77 40
rect 70 34 71 39
rect 76 34 77 39
rect 70 33 77 34
rect 98 39 105 40
rect 98 34 99 39
rect 104 34 105 39
rect 116 38 117 43
rect 122 38 123 43
rect 151 40 156 44
rect 227 41 261 45
rect 302 44 311 45
rect 319 44 341 45
rect 226 40 261 41
rect 301 43 308 44
rect 116 37 123 38
rect 150 39 157 40
rect 150 34 151 39
rect 156 34 157 39
rect 226 35 227 40
rect 232 35 233 40
rect 226 34 233 35
rect 255 39 262 40
rect 255 34 256 39
rect 261 34 262 39
rect 98 33 105 34
rect 134 33 141 34
rect 150 33 157 34
rect 167 33 174 34
rect 255 33 262 34
rect 283 39 290 40
rect 283 34 284 39
rect 289 34 290 39
rect 301 38 302 43
rect 307 38 308 43
rect 336 40 341 44
rect 412 41 446 45
rect 487 44 496 45
rect 504 44 526 45
rect 411 40 446 41
rect 486 43 493 44
rect 301 37 308 38
rect 335 39 342 40
rect 335 34 336 39
rect 341 34 342 39
rect 411 35 412 40
rect 417 35 418 40
rect 411 34 418 35
rect 440 39 447 40
rect 440 34 441 39
rect 446 34 447 39
rect 283 33 290 34
rect 319 33 326 34
rect 335 33 342 34
rect 352 33 359 34
rect 440 33 447 34
rect 468 39 475 40
rect 468 34 469 39
rect 474 34 475 39
rect 486 38 487 43
rect 492 38 493 43
rect 521 40 526 44
rect 597 41 631 45
rect 672 44 681 45
rect 689 44 711 45
rect 596 40 631 41
rect 671 43 678 44
rect 486 37 493 38
rect 520 39 527 40
rect 520 34 521 39
rect 526 34 527 39
rect 596 35 597 40
rect 602 35 603 40
rect 596 34 603 35
rect 625 39 632 40
rect 625 34 626 39
rect 631 34 632 39
rect 468 33 475 34
rect 504 33 511 34
rect 520 33 527 34
rect 537 33 544 34
rect 625 33 632 34
rect 653 39 660 40
rect 653 34 654 39
rect 659 34 660 39
rect 671 38 672 43
rect 677 38 678 43
rect 706 40 711 44
rect 671 37 678 38
rect 705 39 712 40
rect 705 34 706 39
rect 711 34 712 39
rect 653 33 660 34
rect 689 33 696 34
rect 705 33 712 34
rect 722 33 729 34
rect 55 31 62 32
rect 55 26 56 31
rect 61 30 62 31
rect 99 30 104 33
rect 61 26 104 30
rect 134 28 135 33
rect 140 28 141 33
rect 167 28 168 33
rect 173 28 174 33
rect 134 27 174 28
rect 55 25 104 26
rect 135 23 174 27
rect 240 31 247 32
rect 240 26 241 31
rect 246 30 247 31
rect 284 30 289 33
rect 246 26 289 30
rect 319 28 320 33
rect 325 28 326 33
rect 352 28 353 33
rect 358 28 359 33
rect 319 27 359 28
rect 240 25 289 26
rect 320 23 359 27
rect 425 31 432 32
rect 425 26 426 31
rect 431 30 432 31
rect 469 30 474 33
rect 431 26 474 30
rect 504 28 505 33
rect 510 28 511 33
rect 537 28 538 33
rect 543 28 544 33
rect 504 27 544 28
rect 425 25 474 26
rect 505 23 544 27
rect 610 31 617 32
rect 610 26 611 31
rect 616 30 617 31
rect 654 30 659 33
rect 616 26 659 30
rect 689 28 690 33
rect 695 28 696 33
rect 722 28 723 33
rect 728 28 729 33
rect 689 27 729 28
rect 610 25 659 26
rect 690 23 729 27
<< labels >>
rlabel metal1 3 33 7 36 1 D
rlabel metal1 0 70 3 74 4 clk
rlabel metal1 0 0 3 4 2 ~clk
rlabel metal1 7 61 10 65 1 Vdd!
rlabel metal1 8 8 11 12 1 GND!
rlabel metal1 95 36 98 39 1 test2
rlabel metal1 105 34 108 37 1 test1
rlabel metal1 193 8 196 12 1 GND!
rlabel metal1 192 61 195 65 1 Vdd!
rlabel metal1 185 0 188 4 2 ~clk
rlabel metal1 185 70 188 74 4 clk
rlabel metal1 185 32 188 36 1 q0
rlabel metal1 555 70 558 74 4 clk
rlabel metal1 555 0 558 4 2 ~clk
rlabel metal1 562 61 565 65 1 Vdd!
rlabel metal1 563 8 566 12 1 GND!
rlabel metal1 378 8 381 12 1 GND!
rlabel metal1 377 61 380 65 1 Vdd!
rlabel metal1 370 0 373 4 2 ~clk
rlabel metal1 370 70 373 74 4 clk
rlabel metal1 370 32 373 37 1 q1
rlabel metal1 555 32 558 36 1 q2
rlabel metal1 740 32 743 36 7 q3
<< end >>
