magic
tech scmos
timestamp 1608269925
<< ntransistor >>
rect 2763 4183 2765 4187
rect 2789 4179 2791 4183
rect 2794 4179 2796 4183
rect 2817 4175 2819 4179
rect 2718 4156 2720 4166
rect 2789 4149 2791 4153
rect 2794 4149 2796 4153
<< ptransistor >>
rect 2718 4186 2720 4206
rect 2763 4201 2765 4209
rect 2789 4195 2791 4203
rect 2794 4195 2796 4203
rect 2817 4201 2819 4209
rect 2789 4129 2791 4137
rect 2794 4129 2796 4137
<< ndiffusion >>
rect 2762 4183 2763 4187
rect 2765 4183 2766 4187
rect 2786 4179 2789 4183
rect 2791 4179 2794 4183
rect 2796 4179 2797 4183
rect 2816 4175 2817 4179
rect 2819 4175 2820 4179
rect 2717 4156 2718 4166
rect 2720 4156 2721 4166
rect 2786 4149 2789 4153
rect 2791 4149 2794 4153
rect 2796 4149 2797 4153
<< pdiffusion >>
rect 2717 4186 2718 4206
rect 2720 4186 2721 4206
rect 2762 4201 2763 4209
rect 2765 4201 2766 4209
rect 2786 4195 2789 4203
rect 2791 4195 2794 4203
rect 2796 4195 2797 4203
rect 2816 4201 2817 4209
rect 2819 4201 2820 4209
rect 2786 4129 2789 4137
rect 2791 4129 2794 4137
rect 2796 4129 2797 4137
<< ndcontact >>
rect 2758 4183 2762 4187
rect 2766 4183 2770 4187
rect 2782 4179 2786 4183
rect 2797 4179 2801 4183
rect 2812 4175 2816 4179
rect 2820 4175 2824 4179
rect 2693 4156 2717 4166
rect 2721 4156 2745 4166
rect 2782 4149 2786 4153
rect 2797 4149 2801 4153
<< pdcontact >>
rect 2693 4186 2717 4206
rect 2721 4186 2745 4206
rect 2758 4201 2762 4209
rect 2766 4201 2770 4209
rect 2782 4195 2786 4203
rect 2797 4195 2801 4203
rect 2812 4201 2816 4209
rect 2820 4201 2824 4209
rect 2782 4129 2786 4137
rect 2797 4129 2801 4137
<< psubstratepcontact >>
rect 2751 4163 2755 4167
rect 2775 4163 2779 4167
rect 2829 4163 2833 4167
<< nsubstratencontact >>
rect 2751 4213 2755 4217
rect 2775 4213 2779 4217
rect 2829 4213 2833 4217
rect 2775 4113 2779 4117
<< polysilicon >>
rect 2763 4209 2765 4211
rect 2718 4206 2720 4209
rect 2789 4203 2791 4207
rect 2817 4209 2819 4211
rect 2794 4203 2796 4206
rect 2763 4187 2765 4201
rect 2789 4192 2791 4195
rect 2794 4193 2796 4195
rect 2790 4188 2791 4192
rect 2718 4178 2720 4186
rect 2789 4183 2791 4188
rect 2794 4183 2796 4185
rect 2763 4181 2765 4183
rect 2817 4179 2819 4201
rect 2789 4177 2791 4179
rect 2794 4174 2796 4179
rect 2718 4166 2720 4174
rect 2817 4173 2819 4175
rect 2718 4154 2720 4156
rect 2789 4153 2791 4156
rect 2794 4153 2796 4156
rect 2789 4137 2791 4149
rect 2794 4147 2796 4149
rect 2794 4137 2796 4139
rect 2789 4127 2791 4129
rect 2794 4124 2796 4129
<< polycontact >>
rect 2794 4206 2798 4210
rect 2759 4192 2763 4196
rect 2786 4188 2790 4192
rect 2813 4184 2817 4188
rect 2716 4174 2720 4178
rect 2792 4170 2796 4174
rect 2794 4156 2798 4160
rect 2783 4140 2789 4144
rect 2792 4120 2796 4124
<< metal1 >>
rect 1376 4845 1460 4930
rect 1679 4820 1757 4909
rect 1986 4825 2064 4914
rect 2303 4825 2381 4914
rect 2614 4827 2692 4916
rect 2918 4817 2996 4906
rect 3232 4825 3310 4914
rect 3522 4810 3634 4924
rect 1718 4300 1731 4326
rect 2027 4300 2040 4326
rect 2336 4300 2349 4354
rect 2645 4316 2658 4338
rect 2954 4300 2967 4338
rect 3263 4300 3276 4338
rect 2686 4213 2751 4217
rect 2755 4213 2775 4217
rect 2779 4213 2829 4217
rect 2693 4206 2696 4213
rect 2758 4209 2761 4213
rect 2767 4196 2770 4201
rect 2782 4203 2785 4213
rect 2812 4209 2815 4213
rect 2751 4192 2752 4195
rect 2756 4192 2759 4195
rect 2798 4192 2801 4195
rect 2767 4187 2770 4192
rect 2778 4188 2786 4191
rect 2798 4189 2806 4192
rect 2658 4174 2716 4178
rect 2742 4166 2745 4186
rect 2798 4183 2801 4189
rect 2810 4184 2813 4187
rect 2821 4187 2824 4201
rect 2821 4184 2833 4187
rect 2758 4167 2761 4183
rect 2821 4179 2824 4184
rect 2782 4167 2785 4179
rect 2812 4167 2815 4175
rect 2755 4163 2775 4167
rect 2779 4163 2829 4167
rect 2693 4149 2696 4156
rect 2782 4153 2785 4163
rect 2684 4145 2748 4149
rect 2778 4141 2783 4144
rect 2798 4143 2801 4149
rect 2798 4140 2806 4143
rect 2798 4137 2801 4140
rect 2782 4117 2785 4129
rect 2751 4113 2775 4117
rect 2779 4113 2833 4117
<< m2contact >>
rect 2645 4312 2658 4316
rect 2798 4206 2802 4210
rect 2752 4192 2756 4196
rect 2767 4192 2771 4196
rect 2645 4174 2658 4178
rect 2806 4184 2810 4192
rect 2788 4170 2792 4174
rect 2798 4156 2802 4160
rect 2806 4140 2810 4144
rect 2788 4120 2792 4124
<< metal2 >>
rect 2080 4448 2088 4450
rect 2080 4443 2081 4448
rect 2086 4443 2088 4448
rect 2080 4330 2088 4443
rect 2080 4323 2093 4330
rect 2087 4300 2093 4323
rect 2171 4326 2172 4330
rect 2171 4300 2175 4326
rect 2645 4178 2658 4312
rect 2753 4206 2798 4209
rect 2753 4196 2756 4206
rect 2771 4193 2791 4196
rect 2788 4174 2791 4193
rect 2788 4124 2791 4170
rect 2799 4160 2802 4206
rect 2806 4144 2810 4184
<< m3contact >>
rect 2081 4443 2086 4448
rect 2172 4326 2176 4330
<< metal3 >>
rect 2080 4448 2088 4450
rect 2080 4443 2081 4448
rect 2086 4443 2088 4448
rect 2080 4442 2088 4443
rect 2171 4330 2177 4331
rect 2171 4326 2172 4330
rect 2176 4326 2177 4330
rect 2171 4325 2177 4326
use OutPad  OutPad_0
timestamp 1012172318
transform 1 0 2565 0 1 5183
box 17 -26 326 657
use BlankPad  t0
timestamp 1006127261
transform 1 0 960 0 1 4368
box -11 -51 298 632
use GNDPad  t1
timestamp 1509371954
transform 1 0 1258 0 1 4352
box 0 -35 309 648
use InPad  t2
timestamp 1509371954
transform 1 0 1599 0 1 4683
box -32 -366 277 317
use InPad  t3
timestamp 1509371954
transform 1 0 1908 0 1 4683
box -32 -366 277 317
use InPad  t4
timestamp 1509371954
transform 1 0 2217 0 1 4683
box -32 -366 277 317
use InPad  InPad_0
timestamp 1509371954
transform 1 0 2526 0 1 4683
box -32 -366 277 317
use InPad  InPad_1
timestamp 1509371954
transform 1 0 2835 0 1 4683
box -32 -366 277 317
use OutPad  t7
timestamp 1012172318
transform 1 0 3095 0 1 4343
box 17 -26 326 657
use VddPad  t8
timestamp 1509371954
transform 1 0 3421 0 1 4352
box 0 -35 309 648
use BlankPad  t9
timestamp 1006127261
transform 1 0 3741 0 1 4368
box -11 -51 298 632
use Corner  crt
timestamp 1012241868
transform 0 1 4369 -1 0 4825
box -143 -333 774 618
use Corner  clt
timestamp 1012241868
transform 1 0 175 0 1 4369
box -143 -333 774 618
use BlankPad  l9
timestamp 1006127261
transform 0 -1 632 1 0 3740
box -11 -51 298 632
use BlankPad  l8
timestamp 1006127261
transform 0 -1 632 1 0 3431
box -11 -51 298 632
use BlankPad  l7
timestamp 1006127261
transform 0 -1 632 1 0 3122
box -11 -51 298 632
use BlankPad  l6
timestamp 1006127261
transform 0 -1 632 1 0 2813
box -11 -51 298 632
use BlankPad  l5
timestamp 1006127261
transform 0 -1 632 1 0 2504
box -11 -51 298 632
use BlankPad  l4
timestamp 1006127261
transform 0 -1 632 1 0 2195
box -11 -51 298 632
use BlankPad  l3
timestamp 1006127261
transform 0 -1 632 1 0 1886
box -11 -51 298 632
use BlankPad  l2
timestamp 1006127261
transform 0 -1 632 1 0 1577
box -11 -51 298 632
use BlankPad  l1
timestamp 1006127261
transform 0 -1 632 1 0 1268
box -11 -51 298 632
use BlankPad  r9
timestamp 1006127261
transform 0 1 4368 -1 0 4040
box -11 -51 298 632
use BlankPad  r8
timestamp 1006127261
transform 0 1 4368 -1 0 3731
box -11 -51 298 632
use BlankPad  r7
timestamp 1006127261
transform 0 1 4368 -1 0 3422
box -11 -51 298 632
use BlankPad  r6
timestamp 1006127261
transform 0 1 4368 -1 0 3113
box -11 -51 298 632
use BlankPad  r5
timestamp 1006127261
transform 0 1 4368 -1 0 2804
box -11 -51 298 632
use BlankPad  r4
timestamp 1006127261
transform 0 1 4368 -1 0 2495
box -11 -51 298 632
use BlankPad  r3
timestamp 1006127261
transform 0 1 4368 -1 0 2186
box -11 -51 298 632
use BlankPad  r2
timestamp 1006127261
transform 0 1 4368 -1 0 1877
box -11 -51 298 632
use BlankPad  r1
timestamp 1006127261
transform 0 1 4368 -1 0 1568
box -11 -51 298 632
use BlankPad  r0
timestamp 1006127261
transform 0 1 4368 -1 0 1259
box -11 -51 298 632
use BlankPad  l0
timestamp 1006127261
transform 0 -1 632 1 0 959
box -11 -51 298 632
use Corner  clb
timestamp 1012241868
transform 0 -1 631 1 0 175
box -143 -333 774 618
use BlankPad  b0
timestamp 1006127261
transform -1 0 1260 0 -1 632
box -11 -51 298 632
use BlankPad  b1
timestamp 1006127261
transform -1 0 1569 0 -1 632
box -11 -51 298 632
use BlankPad  b2
timestamp 1006127261
transform -1 0 1878 0 -1 632
box -11 -51 298 632
use BlankPad  b3
timestamp 1006127261
transform -1 0 2187 0 -1 632
box -11 -51 298 632
use BlankPad  b4
timestamp 1006127261
transform -1 0 2496 0 -1 632
box -11 -51 298 632
use BlankPad  b5
timestamp 1006127261
transform -1 0 2805 0 -1 632
box -11 -51 298 632
use BlankPad  b6
timestamp 1006127261
transform -1 0 3114 0 -1 632
box -11 -51 298 632
use BlankPad  b7
timestamp 1006127261
transform -1 0 3423 0 -1 632
box -11 -51 298 632
use BlankPad  b8
timestamp 1006127261
transform -1 0 3732 0 -1 632
box -11 -51 298 632
use Corner  crb
timestamp 1012241868
transform -1 0 4825 0 -1 631
box -143 -333 774 618
use BlankPad  b9
timestamp 1006127261
transform -1 0 4041 0 -1 632
box -11 -51 298 632
<< labels >>
rlabel space 2500 2500 2500 2500 2 Core
rlabel metal1 1716 4857 1720 4857 1 p0
rlabel metal1 2031 4873 2031 4873 1 p1
rlabel metal1 2340 4865 2340 4865 1 p2
rlabel metal1 3267 4862 3267 4862 1 p5
rlabel metal1 1417 4883 1419 4884 1 p6
rlabel metal1 3571 4861 3572 4861 1 p7
rlabel metal1 2637 4868 2637 4868 1 p3
rlabel metal1 2951 4862 2951 4862 1 p4
rlabel metal1 2830 4184 2833 4187 7 y0
rlabel metal1 2779 4113 2783 4117 1 Vdd!
rlabel metal1 2780 4163 2783 4167 1 GND!
rlabel metal1 2778 4141 2782 4144 3 a1
rlabel metal1 2779 4213 2783 4217 1 Vdd!
rlabel metal1 2778 4188 2782 4191 3 a0
rlabel metal1 2751 4192 2752 4195 3 select0
<< end >>
