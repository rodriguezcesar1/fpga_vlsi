magic
tech scmos
timestamp 1608329531
<< ntransistor >>
rect 2770 4006 2772 4010
rect 2775 4006 2777 4010
rect 2791 4006 2793 4010
rect 2807 4006 2809 4010
rect 2812 4006 2814 4010
rect 2833 4006 2835 4010
rect 2849 4006 2851 4010
rect 2865 4006 2867 4010
rect 2870 4006 2872 4010
rect 2886 4006 2888 4010
rect 2902 4006 2904 4010
rect 2907 4006 2909 4010
rect 2923 4006 2925 4010
rect 2939 4006 2941 4010
rect 2944 4006 2946 4010
rect 2965 4006 2967 4010
rect 2981 4006 2983 4010
rect 2997 4006 2999 4010
rect 3002 4006 3004 4010
rect 3018 4006 3020 4010
rect 3034 4006 3036 4010
rect 3039 4006 3041 4010
rect 3055 4006 3057 4010
rect 3071 4006 3073 4010
rect 3076 4006 3078 4010
rect 3097 4006 3099 4010
rect 3113 4006 3115 4010
rect 3129 4006 3131 4010
rect 3134 4006 3136 4010
rect 3150 4006 3152 4010
rect 3166 4006 3168 4010
rect 3171 4006 3173 4010
rect 3187 4006 3189 4010
rect 3203 4006 3205 4010
rect 3208 4006 3210 4010
rect 3229 4006 3231 4010
rect 3245 4006 3247 4010
rect 3261 4006 3263 4010
rect 3266 4006 3268 4010
rect 3282 4006 3284 4010
rect 3715 4006 3717 4010
rect 3720 4006 3722 4010
rect 3736 4006 3738 4010
rect 3752 4006 3754 4010
rect 3757 4006 3759 4010
rect 3778 4006 3780 4010
rect 3794 4006 3796 4010
rect 3810 4006 3812 4010
rect 3815 4006 3817 4010
rect 3831 4006 3833 4010
rect 3847 4006 3849 4010
rect 3852 4006 3854 4010
rect 3868 4006 3870 4010
rect 3884 4006 3886 4010
rect 3889 4006 3891 4010
rect 3910 4006 3912 4010
rect 3926 4006 3928 4010
rect 3942 4006 3944 4010
rect 3947 4006 3949 4010
rect 3963 4006 3965 4010
rect 3979 4006 3981 4010
rect 3984 4006 3986 4010
rect 4000 4006 4002 4010
rect 4016 4006 4018 4010
rect 4021 4006 4023 4010
rect 4042 4006 4044 4010
rect 4058 4006 4060 4010
rect 4074 4006 4076 4010
rect 4079 4006 4081 4010
rect 4095 4006 4097 4010
rect 4111 4006 4113 4010
rect 4116 4006 4118 4010
rect 4132 4006 4134 4010
rect 4148 4006 4150 4010
rect 4153 4006 4155 4010
rect 4174 4006 4176 4010
rect 4190 4006 4192 4010
rect 4206 4006 4208 4010
rect 4211 4006 4213 4010
rect 4227 4006 4229 4010
rect 2418 3973 2420 3977
rect 2423 3973 2425 3977
rect 2439 3973 2441 3977
rect 2455 3973 2457 3977
rect 2460 3973 2462 3977
rect 2481 3973 2483 3977
rect 2497 3973 2499 3977
rect 2513 3973 2515 3977
rect 2518 3973 2520 3977
rect 2534 3973 2536 3977
rect 3363 3973 3365 3977
rect 3368 3973 3370 3977
rect 3384 3973 3386 3977
rect 3400 3973 3402 3977
rect 3405 3973 3407 3977
rect 3426 3973 3428 3977
rect 3442 3973 3444 3977
rect 3458 3973 3460 3977
rect 3463 3973 3465 3977
rect 3479 3973 3481 3977
rect 2542 3936 2544 3940
rect 2949 3940 2951 3944
rect 2975 3936 2977 3940
rect 2980 3936 2982 3940
rect 3030 3940 3032 3944
rect 3056 3936 3058 3940
rect 3061 3936 3063 3940
rect 3003 3932 3005 3936
rect 2425 3927 2427 3931
rect 2775 3927 2777 3931
rect 2791 3927 2793 3931
rect 2807 3927 2809 3931
rect 2830 3927 2832 3931
rect 2835 3927 2837 3931
rect 2861 3927 2863 3931
rect 2882 3927 2884 3931
rect 2902 3927 2904 3931
rect 2907 3927 2909 3931
rect 2925 3927 2927 3931
rect 3084 3932 3086 3936
rect 3487 3936 3489 3940
rect 3894 3940 3896 3944
rect 3920 3936 3922 3940
rect 3925 3936 3927 3940
rect 3975 3940 3977 3944
rect 4001 3936 4003 3940
rect 4006 3936 4008 3940
rect 3948 3932 3950 3936
rect 3370 3927 3372 3931
rect 3720 3927 3722 3931
rect 3736 3927 3738 3931
rect 3752 3927 3754 3931
rect 3775 3927 3777 3931
rect 3780 3927 3782 3931
rect 3806 3927 3808 3931
rect 3827 3927 3829 3931
rect 3847 3927 3849 3931
rect 3852 3927 3854 3931
rect 3870 3927 3872 3931
rect 4029 3932 4031 3936
rect 2775 3881 2777 3885
rect 2791 3881 2793 3885
rect 2807 3881 2809 3885
rect 2830 3881 2832 3885
rect 2835 3881 2837 3885
rect 2861 3881 2863 3885
rect 2882 3881 2884 3885
rect 2902 3881 2904 3885
rect 2907 3881 2909 3885
rect 2925 3881 2927 3885
rect 2409 3871 2411 3875
rect 2425 3871 2427 3875
rect 2430 3871 2432 3875
rect 2446 3871 2448 3875
rect 2462 3871 2464 3875
rect 2483 3871 2485 3875
rect 2488 3871 2490 3875
rect 2504 3871 2506 3875
rect 2520 3871 2522 3875
rect 2525 3871 2527 3875
rect 2975 3880 2977 3884
rect 2980 3880 2982 3884
rect 3056 3880 3058 3884
rect 3061 3880 3063 3884
rect 3720 3881 3722 3885
rect 3736 3881 3738 3885
rect 3752 3881 3754 3885
rect 3775 3881 3777 3885
rect 3780 3881 3782 3885
rect 3806 3881 3808 3885
rect 3827 3881 3829 3885
rect 3847 3881 3849 3885
rect 3852 3881 3854 3885
rect 3870 3881 3872 3885
rect 3354 3871 3356 3875
rect 3370 3871 3372 3875
rect 3375 3871 3377 3875
rect 3391 3871 3393 3875
rect 3407 3871 3409 3875
rect 3428 3871 3430 3875
rect 3433 3871 3435 3875
rect 3449 3871 3451 3875
rect 3465 3871 3467 3875
rect 3470 3871 3472 3875
rect 3920 3880 3922 3884
rect 3925 3880 3927 3884
rect 4001 3880 4003 3884
rect 4006 3880 4008 3884
rect 2975 3804 2977 3808
rect 2980 3804 2982 3808
rect 3054 3808 3056 3812
rect 3080 3804 3082 3808
rect 3085 3804 3087 3808
rect 3003 3800 3005 3804
rect 2775 3795 2777 3799
rect 2791 3795 2793 3799
rect 2807 3795 2809 3799
rect 2830 3795 2832 3799
rect 2835 3795 2837 3799
rect 2861 3795 2863 3799
rect 2882 3795 2884 3799
rect 2902 3795 2904 3799
rect 2907 3795 2909 3799
rect 2925 3795 2927 3799
rect 3108 3800 3110 3804
rect 3285 3779 3287 3783
rect 3311 3775 3313 3779
rect 3316 3775 3318 3779
rect 3339 3771 3341 3775
rect 3920 3804 3922 3808
rect 3925 3804 3927 3808
rect 3999 3808 4001 3812
rect 4025 3804 4027 3808
rect 4030 3804 4032 3808
rect 3948 3800 3950 3804
rect 3720 3795 3722 3799
rect 3736 3795 3738 3799
rect 3752 3795 3754 3799
rect 3775 3795 3777 3799
rect 3780 3795 3782 3799
rect 3806 3795 3808 3799
rect 3827 3795 3829 3799
rect 3847 3795 3849 3799
rect 3852 3795 3854 3799
rect 3870 3795 3872 3799
rect 4053 3800 4055 3804
rect 2775 3749 2777 3753
rect 2791 3749 2793 3753
rect 2807 3749 2809 3753
rect 2830 3749 2832 3753
rect 2835 3749 2837 3753
rect 2861 3749 2863 3753
rect 2882 3749 2884 3753
rect 2902 3749 2904 3753
rect 2907 3749 2909 3753
rect 2925 3749 2927 3753
rect 2975 3749 2977 3753
rect 2980 3749 2982 3753
rect 3080 3749 3082 3753
rect 3085 3749 3087 3753
rect 3471 3740 3473 3752
rect 3524 3740 3526 3752
rect 3720 3749 3722 3753
rect 3736 3749 3738 3753
rect 3752 3749 3754 3753
rect 3775 3749 3777 3753
rect 3780 3749 3782 3753
rect 3806 3749 3808 3753
rect 3827 3749 3829 3753
rect 3847 3749 3849 3753
rect 3852 3749 3854 3753
rect 3870 3749 3872 3753
rect 3920 3749 3922 3753
rect 3925 3749 3927 3753
rect 4025 3749 4027 3753
rect 4030 3749 4032 3753
rect 3311 3715 3313 3719
rect 3316 3715 3318 3719
rect 2975 3672 2977 3676
rect 2980 3672 2982 3676
rect 3030 3676 3032 3680
rect 3056 3672 3058 3676
rect 3061 3672 3063 3676
rect 3120 3676 3122 3680
rect 3146 3672 3148 3676
rect 3151 3672 3153 3676
rect 3003 3668 3005 3672
rect 2775 3663 2777 3667
rect 2791 3663 2793 3667
rect 2807 3663 2809 3667
rect 2830 3663 2832 3667
rect 2835 3663 2837 3667
rect 2861 3663 2863 3667
rect 2882 3663 2884 3667
rect 2902 3663 2904 3667
rect 2907 3663 2909 3667
rect 2925 3663 2927 3667
rect 3084 3668 3086 3672
rect 3174 3668 3176 3672
rect 3263 3649 3265 3653
rect 3285 3649 3287 3653
rect 3311 3645 3313 3649
rect 3316 3645 3318 3649
rect 3339 3641 3341 3645
rect 3920 3672 3922 3676
rect 3925 3672 3927 3676
rect 3975 3676 3977 3680
rect 4001 3672 4003 3676
rect 4006 3672 4008 3676
rect 4065 3676 4067 3680
rect 4091 3672 4093 3676
rect 4096 3672 4098 3676
rect 3948 3668 3950 3672
rect 3720 3663 3722 3667
rect 3736 3663 3738 3667
rect 3752 3663 3754 3667
rect 3775 3663 3777 3667
rect 3780 3663 3782 3667
rect 3806 3663 3808 3667
rect 3827 3663 3829 3667
rect 3847 3663 3849 3667
rect 3852 3663 3854 3667
rect 3870 3663 3872 3667
rect 4029 3668 4031 3672
rect 4119 3668 4121 3672
rect 2775 3617 2777 3621
rect 2791 3617 2793 3621
rect 2807 3617 2809 3621
rect 2830 3617 2832 3621
rect 2835 3617 2837 3621
rect 2861 3617 2863 3621
rect 2882 3617 2884 3621
rect 2902 3617 2904 3621
rect 2907 3617 2909 3621
rect 2925 3617 2927 3621
rect 2975 3614 2977 3618
rect 2980 3614 2982 3618
rect 3056 3614 3058 3618
rect 3061 3614 3063 3618
rect 3146 3614 3148 3618
rect 3151 3614 3153 3618
rect 3377 3610 3379 3622
rect 3430 3610 3432 3622
rect 3720 3617 3722 3621
rect 3736 3617 3738 3621
rect 3752 3617 3754 3621
rect 3775 3617 3777 3621
rect 3780 3617 3782 3621
rect 3806 3617 3808 3621
rect 3827 3617 3829 3621
rect 3847 3617 3849 3621
rect 3852 3617 3854 3621
rect 3870 3617 3872 3621
rect 3920 3614 3922 3618
rect 3925 3614 3927 3618
rect 4001 3614 4003 3618
rect 4006 3614 4008 3618
rect 4091 3614 4093 3618
rect 4096 3614 4098 3618
rect 3311 3585 3313 3589
rect 3316 3585 3318 3589
rect 2975 3540 2977 3544
rect 2980 3540 2982 3544
rect 3003 3536 3005 3540
rect 2775 3531 2777 3535
rect 2791 3531 2793 3535
rect 2807 3531 2809 3535
rect 2830 3531 2832 3535
rect 2835 3531 2837 3535
rect 2861 3531 2863 3535
rect 2882 3531 2884 3535
rect 2902 3531 2904 3535
rect 2907 3531 2909 3535
rect 2925 3531 2927 3535
rect 3920 3540 3922 3544
rect 3925 3540 3927 3544
rect 3948 3536 3950 3540
rect 3720 3531 3722 3535
rect 3736 3531 3738 3535
rect 3752 3531 3754 3535
rect 3775 3531 3777 3535
rect 3780 3531 3782 3535
rect 3806 3531 3808 3535
rect 3827 3531 3829 3535
rect 3847 3531 3849 3535
rect 3852 3531 3854 3535
rect 3870 3531 3872 3535
rect 2775 3485 2777 3489
rect 2791 3485 2793 3489
rect 2807 3485 2809 3489
rect 2830 3485 2832 3489
rect 2835 3485 2837 3489
rect 2861 3485 2863 3489
rect 2882 3485 2884 3489
rect 2902 3485 2904 3489
rect 2907 3485 2909 3489
rect 2925 3485 2927 3489
rect 3009 3485 3011 3489
rect 3027 3485 3029 3489
rect 3052 3485 3054 3489
rect 3068 3485 3070 3489
rect 3091 3485 3093 3489
rect 3096 3485 3098 3489
rect 3122 3485 3124 3489
rect 3143 3485 3145 3489
rect 3163 3485 3165 3489
rect 3168 3485 3170 3489
rect 3186 3485 3188 3489
rect 2286 3471 2288 3475
rect 2291 3471 2293 3475
rect 2307 3471 2309 3475
rect 2323 3471 2325 3475
rect 2328 3471 2330 3475
rect 2349 3471 2351 3475
rect 2365 3471 2367 3475
rect 2381 3471 2383 3475
rect 2386 3471 2388 3475
rect 2402 3471 2404 3475
rect 2418 3471 2420 3475
rect 2423 3471 2425 3475
rect 2439 3471 2441 3475
rect 2455 3471 2457 3475
rect 2460 3471 2462 3475
rect 2481 3471 2483 3475
rect 2497 3471 2499 3475
rect 2513 3471 2515 3475
rect 2518 3471 2520 3475
rect 2534 3471 2536 3475
rect 2550 3471 2552 3475
rect 2555 3471 2557 3475
rect 2571 3471 2573 3475
rect 2587 3471 2589 3475
rect 2592 3471 2594 3475
rect 2613 3471 2615 3475
rect 2629 3471 2631 3475
rect 2645 3471 2647 3475
rect 2650 3471 2652 3475
rect 2666 3471 2668 3475
rect 2975 3478 2977 3482
rect 2980 3478 2982 3482
rect 3720 3485 3722 3489
rect 3736 3485 3738 3489
rect 3752 3485 3754 3489
rect 3775 3485 3777 3489
rect 3780 3485 3782 3489
rect 3806 3485 3808 3489
rect 3827 3485 3829 3489
rect 3847 3485 3849 3489
rect 3852 3485 3854 3489
rect 3870 3485 3872 3489
rect 3954 3485 3956 3489
rect 3972 3485 3974 3489
rect 3997 3485 3999 3489
rect 4013 3485 4015 3489
rect 4036 3485 4038 3489
rect 4041 3485 4043 3489
rect 4067 3485 4069 3489
rect 4088 3485 4090 3489
rect 4108 3485 4110 3489
rect 4113 3485 4115 3489
rect 4131 3485 4133 3489
rect 3231 3471 3233 3475
rect 3236 3471 3238 3475
rect 3252 3471 3254 3475
rect 3268 3471 3270 3475
rect 3273 3471 3275 3475
rect 3294 3471 3296 3475
rect 3310 3471 3312 3475
rect 3326 3471 3328 3475
rect 3331 3471 3333 3475
rect 3347 3471 3349 3475
rect 3363 3471 3365 3475
rect 3368 3471 3370 3475
rect 3384 3471 3386 3475
rect 3400 3471 3402 3475
rect 3405 3471 3407 3475
rect 3426 3471 3428 3475
rect 3442 3471 3444 3475
rect 3458 3471 3460 3475
rect 3463 3471 3465 3475
rect 3479 3471 3481 3475
rect 3495 3471 3497 3475
rect 3500 3471 3502 3475
rect 3516 3471 3518 3475
rect 3532 3471 3534 3475
rect 3537 3471 3539 3475
rect 3558 3471 3560 3475
rect 3574 3471 3576 3475
rect 3590 3471 3592 3475
rect 3595 3471 3597 3475
rect 3611 3471 3613 3475
rect 3920 3478 3922 3482
rect 3925 3478 3927 3482
rect 2401 3427 2403 3431
rect 2425 3427 2427 3431
rect 3198 3429 3202 3431
rect 3346 3427 3348 3431
rect 3370 3427 3372 3431
rect 4143 3429 4147 3431
rect 2421 3414 2423 3418
rect 3366 3414 3368 3418
rect 2412 3400 2416 3402
rect 3357 3400 3361 3402
rect 2401 3391 2403 3395
rect 2425 3391 2427 3395
rect 3346 3391 3348 3395
rect 3370 3391 3372 3395
rect 3069 3359 3071 3363
rect 3074 3359 3076 3363
rect 3090 3359 3092 3363
rect 3106 3359 3108 3363
rect 3111 3359 3113 3363
rect 3132 3359 3134 3363
rect 3148 3359 3150 3363
rect 3164 3359 3166 3363
rect 3169 3359 3171 3363
rect 3185 3359 3187 3363
rect 4014 3359 4016 3363
rect 4019 3359 4021 3363
rect 4035 3359 4037 3363
rect 4051 3359 4053 3363
rect 4056 3359 4058 3363
rect 4077 3359 4079 3363
rect 4093 3359 4095 3363
rect 4109 3359 4111 3363
rect 4114 3359 4116 3363
rect 4130 3359 4132 3363
rect 2286 3329 2288 3333
rect 2291 3329 2293 3333
rect 2307 3329 2309 3333
rect 2323 3329 2325 3333
rect 2328 3329 2330 3333
rect 2349 3329 2351 3333
rect 2365 3329 2367 3333
rect 2381 3329 2383 3333
rect 2386 3329 2388 3333
rect 2402 3329 2404 3333
rect 2418 3329 2420 3333
rect 2423 3329 2425 3333
rect 2439 3329 2441 3333
rect 2455 3329 2457 3333
rect 2460 3329 2462 3333
rect 2481 3329 2483 3333
rect 2497 3329 2499 3333
rect 2513 3329 2515 3333
rect 2518 3329 2520 3333
rect 2534 3329 2536 3333
rect 2550 3329 2552 3333
rect 2555 3329 2557 3333
rect 2571 3329 2573 3333
rect 2587 3329 2589 3333
rect 2592 3329 2594 3333
rect 2613 3329 2615 3333
rect 2629 3329 2631 3333
rect 2645 3329 2647 3333
rect 2650 3329 2652 3333
rect 2666 3329 2668 3333
rect 3231 3329 3233 3333
rect 3236 3329 3238 3333
rect 3252 3329 3254 3333
rect 3268 3329 3270 3333
rect 3273 3329 3275 3333
rect 3294 3329 3296 3333
rect 3310 3329 3312 3333
rect 3326 3329 3328 3333
rect 3331 3329 3333 3333
rect 3347 3329 3349 3333
rect 3363 3329 3365 3333
rect 3368 3329 3370 3333
rect 3384 3329 3386 3333
rect 3400 3329 3402 3333
rect 3405 3329 3407 3333
rect 3426 3329 3428 3333
rect 3442 3329 3444 3333
rect 3458 3329 3460 3333
rect 3463 3329 3465 3333
rect 3479 3329 3481 3333
rect 3495 3329 3497 3333
rect 3500 3329 3502 3333
rect 3516 3329 3518 3333
rect 3532 3329 3534 3333
rect 3537 3329 3539 3333
rect 3558 3329 3560 3333
rect 3574 3329 3576 3333
rect 3590 3329 3592 3333
rect 3595 3329 3597 3333
rect 3611 3329 3613 3333
rect 3210 3283 3214 3285
rect 4155 3283 4159 3285
rect 3069 3273 3071 3277
rect 3074 3273 3076 3277
rect 3090 3273 3092 3277
rect 3106 3273 3108 3277
rect 3111 3273 3113 3277
rect 3132 3273 3134 3277
rect 3148 3273 3150 3277
rect 3164 3273 3166 3277
rect 3169 3273 3171 3277
rect 3185 3273 3187 3277
rect 4014 3273 4016 3277
rect 4019 3273 4021 3277
rect 4035 3273 4037 3277
rect 4051 3273 4053 3277
rect 4056 3273 4058 3277
rect 4077 3273 4079 3277
rect 4093 3273 4095 3277
rect 4109 3273 4111 3277
rect 4114 3273 4116 3277
rect 4130 3273 4132 3277
rect 2286 3243 2288 3247
rect 2291 3243 2293 3247
rect 2307 3243 2309 3247
rect 2323 3243 2325 3247
rect 2328 3243 2330 3247
rect 2349 3243 2351 3247
rect 2365 3243 2367 3247
rect 2381 3243 2383 3247
rect 2386 3243 2388 3247
rect 2402 3243 2404 3247
rect 2418 3243 2420 3247
rect 2423 3243 2425 3247
rect 2439 3243 2441 3247
rect 2455 3243 2457 3247
rect 2460 3243 2462 3247
rect 2481 3243 2483 3247
rect 2497 3243 2499 3247
rect 2513 3243 2515 3247
rect 2518 3243 2520 3247
rect 2534 3243 2536 3247
rect 2550 3243 2552 3247
rect 2555 3243 2557 3247
rect 2571 3243 2573 3247
rect 2587 3243 2589 3247
rect 2592 3243 2594 3247
rect 2613 3243 2615 3247
rect 2629 3243 2631 3247
rect 2645 3243 2647 3247
rect 2650 3243 2652 3247
rect 2666 3243 2668 3247
rect 3231 3243 3233 3247
rect 3236 3243 3238 3247
rect 3252 3243 3254 3247
rect 3268 3243 3270 3247
rect 3273 3243 3275 3247
rect 3294 3243 3296 3247
rect 3310 3243 3312 3247
rect 3326 3243 3328 3247
rect 3331 3243 3333 3247
rect 3347 3243 3349 3247
rect 3363 3243 3365 3247
rect 3368 3243 3370 3247
rect 3384 3243 3386 3247
rect 3400 3243 3402 3247
rect 3405 3243 3407 3247
rect 3426 3243 3428 3247
rect 3442 3243 3444 3247
rect 3458 3243 3460 3247
rect 3463 3243 3465 3247
rect 3479 3243 3481 3247
rect 3495 3243 3497 3247
rect 3500 3243 3502 3247
rect 3516 3243 3518 3247
rect 3532 3243 3534 3247
rect 3537 3243 3539 3247
rect 3558 3243 3560 3247
rect 3574 3243 3576 3247
rect 3590 3243 3592 3247
rect 3595 3243 3597 3247
rect 3611 3243 3613 3247
rect 2518 3199 2520 3203
rect 2542 3199 2544 3203
rect 3463 3199 3465 3203
rect 3487 3199 3489 3203
rect 2538 3188 2540 3192
rect 3483 3188 3485 3192
rect 2529 3174 2533 3176
rect 3474 3174 3478 3176
rect 2518 3165 2520 3169
rect 2542 3165 2544 3169
rect 3463 3165 3465 3169
rect 3487 3165 3489 3169
rect 2286 3103 2288 3107
rect 2291 3103 2293 3107
rect 2307 3103 2309 3107
rect 2323 3103 2325 3107
rect 2328 3103 2330 3107
rect 2349 3103 2351 3107
rect 2365 3103 2367 3107
rect 2381 3103 2383 3107
rect 2386 3103 2388 3107
rect 2402 3103 2404 3107
rect 2418 3103 2420 3107
rect 2423 3103 2425 3107
rect 2439 3103 2441 3107
rect 2455 3103 2457 3107
rect 2460 3103 2462 3107
rect 2481 3103 2483 3107
rect 2497 3103 2499 3107
rect 2513 3103 2515 3107
rect 2518 3103 2520 3107
rect 2534 3103 2536 3107
rect 2550 3103 2552 3107
rect 2555 3103 2557 3107
rect 2571 3103 2573 3107
rect 2587 3103 2589 3107
rect 2592 3103 2594 3107
rect 2613 3103 2615 3107
rect 2629 3103 2631 3107
rect 2645 3103 2647 3107
rect 2650 3103 2652 3107
rect 2666 3103 2668 3107
rect 3231 3103 3233 3107
rect 3236 3103 3238 3107
rect 3252 3103 3254 3107
rect 3268 3103 3270 3107
rect 3273 3103 3275 3107
rect 3294 3103 3296 3107
rect 3310 3103 3312 3107
rect 3326 3103 3328 3107
rect 3331 3103 3333 3107
rect 3347 3103 3349 3107
rect 3363 3103 3365 3107
rect 3368 3103 3370 3107
rect 3384 3103 3386 3107
rect 3400 3103 3402 3107
rect 3405 3103 3407 3107
rect 3426 3103 3428 3107
rect 3442 3103 3444 3107
rect 3458 3103 3460 3107
rect 3463 3103 3465 3107
rect 3479 3103 3481 3107
rect 3495 3103 3497 3107
rect 3500 3103 3502 3107
rect 3516 3103 3518 3107
rect 3532 3103 3534 3107
rect 3537 3103 3539 3107
rect 3558 3103 3560 3107
rect 3574 3103 3576 3107
rect 3590 3103 3592 3107
rect 3595 3103 3597 3107
rect 3611 3103 3613 3107
rect 2770 3024 2772 3028
rect 2775 3024 2777 3028
rect 2791 3024 2793 3028
rect 2807 3024 2809 3028
rect 2812 3024 2814 3028
rect 2833 3024 2835 3028
rect 2849 3024 2851 3028
rect 2865 3024 2867 3028
rect 2870 3024 2872 3028
rect 2886 3024 2888 3028
rect 2902 3024 2904 3028
rect 2907 3024 2909 3028
rect 2923 3024 2925 3028
rect 2939 3024 2941 3028
rect 2944 3024 2946 3028
rect 2965 3024 2967 3028
rect 2981 3024 2983 3028
rect 2997 3024 2999 3028
rect 3002 3024 3004 3028
rect 3018 3024 3020 3028
rect 3034 3024 3036 3028
rect 3039 3024 3041 3028
rect 3055 3024 3057 3028
rect 3071 3024 3073 3028
rect 3076 3024 3078 3028
rect 3097 3024 3099 3028
rect 3113 3024 3115 3028
rect 3129 3024 3131 3028
rect 3134 3024 3136 3028
rect 3150 3024 3152 3028
rect 3166 3024 3168 3028
rect 3171 3024 3173 3028
rect 3187 3024 3189 3028
rect 3203 3024 3205 3028
rect 3208 3024 3210 3028
rect 3229 3024 3231 3028
rect 3245 3024 3247 3028
rect 3261 3024 3263 3028
rect 3266 3024 3268 3028
rect 3282 3024 3284 3028
rect 3715 3024 3717 3028
rect 3720 3024 3722 3028
rect 3736 3024 3738 3028
rect 3752 3024 3754 3028
rect 3757 3024 3759 3028
rect 3778 3024 3780 3028
rect 3794 3024 3796 3028
rect 3810 3024 3812 3028
rect 3815 3024 3817 3028
rect 3831 3024 3833 3028
rect 3847 3024 3849 3028
rect 3852 3024 3854 3028
rect 3868 3024 3870 3028
rect 3884 3024 3886 3028
rect 3889 3024 3891 3028
rect 3910 3024 3912 3028
rect 3926 3024 3928 3028
rect 3942 3024 3944 3028
rect 3947 3024 3949 3028
rect 3963 3024 3965 3028
rect 3979 3024 3981 3028
rect 3984 3024 3986 3028
rect 4000 3024 4002 3028
rect 4016 3024 4018 3028
rect 4021 3024 4023 3028
rect 4042 3024 4044 3028
rect 4058 3024 4060 3028
rect 4074 3024 4076 3028
rect 4079 3024 4081 3028
rect 4095 3024 4097 3028
rect 4111 3024 4113 3028
rect 4116 3024 4118 3028
rect 4132 3024 4134 3028
rect 4148 3024 4150 3028
rect 4153 3024 4155 3028
rect 4174 3024 4176 3028
rect 4190 3024 4192 3028
rect 4206 3024 4208 3028
rect 4211 3024 4213 3028
rect 4227 3024 4229 3028
rect 2418 2991 2420 2995
rect 2423 2991 2425 2995
rect 2439 2991 2441 2995
rect 2455 2991 2457 2995
rect 2460 2991 2462 2995
rect 2481 2991 2483 2995
rect 2497 2991 2499 2995
rect 2513 2991 2515 2995
rect 2518 2991 2520 2995
rect 2534 2991 2536 2995
rect 3363 2991 3365 2995
rect 3368 2991 3370 2995
rect 3384 2991 3386 2995
rect 3400 2991 3402 2995
rect 3405 2991 3407 2995
rect 3426 2991 3428 2995
rect 3442 2991 3444 2995
rect 3458 2991 3460 2995
rect 3463 2991 3465 2995
rect 3479 2991 3481 2995
rect 2542 2954 2544 2958
rect 2949 2958 2951 2962
rect 2975 2954 2977 2958
rect 2980 2954 2982 2958
rect 3030 2958 3032 2962
rect 3056 2954 3058 2958
rect 3061 2954 3063 2958
rect 3003 2950 3005 2954
rect 2425 2945 2427 2949
rect 2775 2945 2777 2949
rect 2791 2945 2793 2949
rect 2807 2945 2809 2949
rect 2830 2945 2832 2949
rect 2835 2945 2837 2949
rect 2861 2945 2863 2949
rect 2882 2945 2884 2949
rect 2902 2945 2904 2949
rect 2907 2945 2909 2949
rect 2925 2945 2927 2949
rect 3084 2950 3086 2954
rect 3487 2954 3489 2958
rect 3894 2958 3896 2962
rect 3920 2954 3922 2958
rect 3925 2954 3927 2958
rect 3975 2958 3977 2962
rect 4001 2954 4003 2958
rect 4006 2954 4008 2958
rect 3948 2950 3950 2954
rect 3370 2945 3372 2949
rect 3720 2945 3722 2949
rect 3736 2945 3738 2949
rect 3752 2945 3754 2949
rect 3775 2945 3777 2949
rect 3780 2945 3782 2949
rect 3806 2945 3808 2949
rect 3827 2945 3829 2949
rect 3847 2945 3849 2949
rect 3852 2945 3854 2949
rect 3870 2945 3872 2949
rect 4029 2950 4031 2954
rect 2775 2899 2777 2903
rect 2791 2899 2793 2903
rect 2807 2899 2809 2903
rect 2830 2899 2832 2903
rect 2835 2899 2837 2903
rect 2861 2899 2863 2903
rect 2882 2899 2884 2903
rect 2902 2899 2904 2903
rect 2907 2899 2909 2903
rect 2925 2899 2927 2903
rect 2409 2889 2411 2893
rect 2425 2889 2427 2893
rect 2430 2889 2432 2893
rect 2446 2889 2448 2893
rect 2462 2889 2464 2893
rect 2483 2889 2485 2893
rect 2488 2889 2490 2893
rect 2504 2889 2506 2893
rect 2520 2889 2522 2893
rect 2525 2889 2527 2893
rect 2975 2898 2977 2902
rect 2980 2898 2982 2902
rect 3056 2898 3058 2902
rect 3061 2898 3063 2902
rect 3720 2899 3722 2903
rect 3736 2899 3738 2903
rect 3752 2899 3754 2903
rect 3775 2899 3777 2903
rect 3780 2899 3782 2903
rect 3806 2899 3808 2903
rect 3827 2899 3829 2903
rect 3847 2899 3849 2903
rect 3852 2899 3854 2903
rect 3870 2899 3872 2903
rect 3354 2889 3356 2893
rect 3370 2889 3372 2893
rect 3375 2889 3377 2893
rect 3391 2889 3393 2893
rect 3407 2889 3409 2893
rect 3428 2889 3430 2893
rect 3433 2889 3435 2893
rect 3449 2889 3451 2893
rect 3465 2889 3467 2893
rect 3470 2889 3472 2893
rect 3920 2898 3922 2902
rect 3925 2898 3927 2902
rect 4001 2898 4003 2902
rect 4006 2898 4008 2902
rect 2975 2822 2977 2826
rect 2980 2822 2982 2826
rect 3054 2826 3056 2830
rect 3080 2822 3082 2826
rect 3085 2822 3087 2826
rect 3003 2818 3005 2822
rect 2775 2813 2777 2817
rect 2791 2813 2793 2817
rect 2807 2813 2809 2817
rect 2830 2813 2832 2817
rect 2835 2813 2837 2817
rect 2861 2813 2863 2817
rect 2882 2813 2884 2817
rect 2902 2813 2904 2817
rect 2907 2813 2909 2817
rect 2925 2813 2927 2817
rect 3108 2818 3110 2822
rect 3920 2822 3922 2826
rect 3925 2822 3927 2826
rect 3999 2826 4001 2830
rect 4025 2822 4027 2826
rect 4030 2822 4032 2826
rect 3948 2818 3950 2822
rect 3720 2813 3722 2817
rect 3736 2813 3738 2817
rect 3752 2813 3754 2817
rect 3775 2813 3777 2817
rect 3780 2813 3782 2817
rect 3806 2813 3808 2817
rect 3827 2813 3829 2817
rect 3847 2813 3849 2817
rect 3852 2813 3854 2817
rect 3870 2813 3872 2817
rect 4053 2818 4055 2822
rect 2775 2767 2777 2771
rect 2791 2767 2793 2771
rect 2807 2767 2809 2771
rect 2830 2767 2832 2771
rect 2835 2767 2837 2771
rect 2861 2767 2863 2771
rect 2882 2767 2884 2771
rect 2902 2767 2904 2771
rect 2907 2767 2909 2771
rect 2925 2767 2927 2771
rect 2975 2767 2977 2771
rect 2980 2767 2982 2771
rect 3080 2767 3082 2771
rect 3085 2767 3087 2771
rect 3720 2767 3722 2771
rect 3736 2767 3738 2771
rect 3752 2767 3754 2771
rect 3775 2767 3777 2771
rect 3780 2767 3782 2771
rect 3806 2767 3808 2771
rect 3827 2767 3829 2771
rect 3847 2767 3849 2771
rect 3852 2767 3854 2771
rect 3870 2767 3872 2771
rect 3920 2767 3922 2771
rect 3925 2767 3927 2771
rect 4025 2767 4027 2771
rect 4030 2767 4032 2771
rect 2975 2690 2977 2694
rect 2980 2690 2982 2694
rect 3030 2694 3032 2698
rect 3056 2690 3058 2694
rect 3061 2690 3063 2694
rect 3120 2694 3122 2698
rect 3146 2690 3148 2694
rect 3151 2690 3153 2694
rect 3003 2686 3005 2690
rect 2775 2681 2777 2685
rect 2791 2681 2793 2685
rect 2807 2681 2809 2685
rect 2830 2681 2832 2685
rect 2835 2681 2837 2685
rect 2861 2681 2863 2685
rect 2882 2681 2884 2685
rect 2902 2681 2904 2685
rect 2907 2681 2909 2685
rect 2925 2681 2927 2685
rect 3084 2686 3086 2690
rect 3174 2686 3176 2690
rect 3920 2690 3922 2694
rect 3925 2690 3927 2694
rect 3975 2694 3977 2698
rect 4001 2690 4003 2694
rect 4006 2690 4008 2694
rect 4065 2694 4067 2698
rect 4091 2690 4093 2694
rect 4096 2690 4098 2694
rect 3948 2686 3950 2690
rect 3720 2681 3722 2685
rect 3736 2681 3738 2685
rect 3752 2681 3754 2685
rect 3775 2681 3777 2685
rect 3780 2681 3782 2685
rect 3806 2681 3808 2685
rect 3827 2681 3829 2685
rect 3847 2681 3849 2685
rect 3852 2681 3854 2685
rect 3870 2681 3872 2685
rect 4029 2686 4031 2690
rect 4119 2686 4121 2690
rect 2775 2635 2777 2639
rect 2791 2635 2793 2639
rect 2807 2635 2809 2639
rect 2830 2635 2832 2639
rect 2835 2635 2837 2639
rect 2861 2635 2863 2639
rect 2882 2635 2884 2639
rect 2902 2635 2904 2639
rect 2907 2635 2909 2639
rect 2925 2635 2927 2639
rect 2975 2632 2977 2636
rect 2980 2632 2982 2636
rect 3056 2632 3058 2636
rect 3061 2632 3063 2636
rect 3146 2632 3148 2636
rect 3151 2632 3153 2636
rect 3720 2635 3722 2639
rect 3736 2635 3738 2639
rect 3752 2635 3754 2639
rect 3775 2635 3777 2639
rect 3780 2635 3782 2639
rect 3806 2635 3808 2639
rect 3827 2635 3829 2639
rect 3847 2635 3849 2639
rect 3852 2635 3854 2639
rect 3870 2635 3872 2639
rect 3920 2632 3922 2636
rect 3925 2632 3927 2636
rect 4001 2632 4003 2636
rect 4006 2632 4008 2636
rect 4091 2632 4093 2636
rect 4096 2632 4098 2636
rect 2975 2558 2977 2562
rect 2980 2558 2982 2562
rect 3003 2554 3005 2558
rect 2775 2549 2777 2553
rect 2791 2549 2793 2553
rect 2807 2549 2809 2553
rect 2830 2549 2832 2553
rect 2835 2549 2837 2553
rect 2861 2549 2863 2553
rect 2882 2549 2884 2553
rect 2902 2549 2904 2553
rect 2907 2549 2909 2553
rect 2925 2549 2927 2553
rect 3920 2558 3922 2562
rect 3925 2558 3927 2562
rect 3948 2554 3950 2558
rect 3720 2549 3722 2553
rect 3736 2549 3738 2553
rect 3752 2549 3754 2553
rect 3775 2549 3777 2553
rect 3780 2549 3782 2553
rect 3806 2549 3808 2553
rect 3827 2549 3829 2553
rect 3847 2549 3849 2553
rect 3852 2549 3854 2553
rect 3870 2549 3872 2553
rect 2775 2503 2777 2507
rect 2791 2503 2793 2507
rect 2807 2503 2809 2507
rect 2830 2503 2832 2507
rect 2835 2503 2837 2507
rect 2861 2503 2863 2507
rect 2882 2503 2884 2507
rect 2902 2503 2904 2507
rect 2907 2503 2909 2507
rect 2925 2503 2927 2507
rect 3009 2503 3011 2507
rect 3027 2503 3029 2507
rect 3052 2503 3054 2507
rect 3068 2503 3070 2507
rect 3091 2503 3093 2507
rect 3096 2503 3098 2507
rect 3122 2503 3124 2507
rect 3143 2503 3145 2507
rect 3163 2503 3165 2507
rect 3168 2503 3170 2507
rect 3186 2503 3188 2507
rect 2286 2489 2288 2493
rect 2291 2489 2293 2493
rect 2307 2489 2309 2493
rect 2323 2489 2325 2493
rect 2328 2489 2330 2493
rect 2349 2489 2351 2493
rect 2365 2489 2367 2493
rect 2381 2489 2383 2493
rect 2386 2489 2388 2493
rect 2402 2489 2404 2493
rect 2418 2489 2420 2493
rect 2423 2489 2425 2493
rect 2439 2489 2441 2493
rect 2455 2489 2457 2493
rect 2460 2489 2462 2493
rect 2481 2489 2483 2493
rect 2497 2489 2499 2493
rect 2513 2489 2515 2493
rect 2518 2489 2520 2493
rect 2534 2489 2536 2493
rect 2550 2489 2552 2493
rect 2555 2489 2557 2493
rect 2571 2489 2573 2493
rect 2587 2489 2589 2493
rect 2592 2489 2594 2493
rect 2613 2489 2615 2493
rect 2629 2489 2631 2493
rect 2645 2489 2647 2493
rect 2650 2489 2652 2493
rect 2666 2489 2668 2493
rect 2975 2496 2977 2500
rect 2980 2496 2982 2500
rect 3720 2503 3722 2507
rect 3736 2503 3738 2507
rect 3752 2503 3754 2507
rect 3775 2503 3777 2507
rect 3780 2503 3782 2507
rect 3806 2503 3808 2507
rect 3827 2503 3829 2507
rect 3847 2503 3849 2507
rect 3852 2503 3854 2507
rect 3870 2503 3872 2507
rect 3954 2503 3956 2507
rect 3972 2503 3974 2507
rect 3997 2503 3999 2507
rect 4013 2503 4015 2507
rect 4036 2503 4038 2507
rect 4041 2503 4043 2507
rect 4067 2503 4069 2507
rect 4088 2503 4090 2507
rect 4108 2503 4110 2507
rect 4113 2503 4115 2507
rect 4131 2503 4133 2507
rect 3231 2489 3233 2493
rect 3236 2489 3238 2493
rect 3252 2489 3254 2493
rect 3268 2489 3270 2493
rect 3273 2489 3275 2493
rect 3294 2489 3296 2493
rect 3310 2489 3312 2493
rect 3326 2489 3328 2493
rect 3331 2489 3333 2493
rect 3347 2489 3349 2493
rect 3363 2489 3365 2493
rect 3368 2489 3370 2493
rect 3384 2489 3386 2493
rect 3400 2489 3402 2493
rect 3405 2489 3407 2493
rect 3426 2489 3428 2493
rect 3442 2489 3444 2493
rect 3458 2489 3460 2493
rect 3463 2489 3465 2493
rect 3479 2489 3481 2493
rect 3495 2489 3497 2493
rect 3500 2489 3502 2493
rect 3516 2489 3518 2493
rect 3532 2489 3534 2493
rect 3537 2489 3539 2493
rect 3558 2489 3560 2493
rect 3574 2489 3576 2493
rect 3590 2489 3592 2493
rect 3595 2489 3597 2493
rect 3611 2489 3613 2493
rect 3920 2496 3922 2500
rect 3925 2496 3927 2500
rect 2401 2445 2403 2449
rect 2425 2445 2427 2449
rect 3198 2447 3202 2449
rect 3346 2445 3348 2449
rect 3370 2445 3372 2449
rect 4143 2447 4147 2449
rect 2421 2432 2423 2436
rect 3366 2432 3368 2436
rect 2412 2418 2416 2420
rect 3357 2418 3361 2420
rect 2401 2409 2403 2413
rect 2425 2409 2427 2413
rect 3346 2409 3348 2413
rect 3370 2409 3372 2413
rect 3069 2377 3071 2381
rect 3074 2377 3076 2381
rect 3090 2377 3092 2381
rect 3106 2377 3108 2381
rect 3111 2377 3113 2381
rect 3132 2377 3134 2381
rect 3148 2377 3150 2381
rect 3164 2377 3166 2381
rect 3169 2377 3171 2381
rect 3185 2377 3187 2381
rect 4014 2377 4016 2381
rect 4019 2377 4021 2381
rect 4035 2377 4037 2381
rect 4051 2377 4053 2381
rect 4056 2377 4058 2381
rect 4077 2377 4079 2381
rect 4093 2377 4095 2381
rect 4109 2377 4111 2381
rect 4114 2377 4116 2381
rect 4130 2377 4132 2381
rect 2286 2347 2288 2351
rect 2291 2347 2293 2351
rect 2307 2347 2309 2351
rect 2323 2347 2325 2351
rect 2328 2347 2330 2351
rect 2349 2347 2351 2351
rect 2365 2347 2367 2351
rect 2381 2347 2383 2351
rect 2386 2347 2388 2351
rect 2402 2347 2404 2351
rect 2418 2347 2420 2351
rect 2423 2347 2425 2351
rect 2439 2347 2441 2351
rect 2455 2347 2457 2351
rect 2460 2347 2462 2351
rect 2481 2347 2483 2351
rect 2497 2347 2499 2351
rect 2513 2347 2515 2351
rect 2518 2347 2520 2351
rect 2534 2347 2536 2351
rect 2550 2347 2552 2351
rect 2555 2347 2557 2351
rect 2571 2347 2573 2351
rect 2587 2347 2589 2351
rect 2592 2347 2594 2351
rect 2613 2347 2615 2351
rect 2629 2347 2631 2351
rect 2645 2347 2647 2351
rect 2650 2347 2652 2351
rect 2666 2347 2668 2351
rect 3231 2347 3233 2351
rect 3236 2347 3238 2351
rect 3252 2347 3254 2351
rect 3268 2347 3270 2351
rect 3273 2347 3275 2351
rect 3294 2347 3296 2351
rect 3310 2347 3312 2351
rect 3326 2347 3328 2351
rect 3331 2347 3333 2351
rect 3347 2347 3349 2351
rect 3363 2347 3365 2351
rect 3368 2347 3370 2351
rect 3384 2347 3386 2351
rect 3400 2347 3402 2351
rect 3405 2347 3407 2351
rect 3426 2347 3428 2351
rect 3442 2347 3444 2351
rect 3458 2347 3460 2351
rect 3463 2347 3465 2351
rect 3479 2347 3481 2351
rect 3495 2347 3497 2351
rect 3500 2347 3502 2351
rect 3516 2347 3518 2351
rect 3532 2347 3534 2351
rect 3537 2347 3539 2351
rect 3558 2347 3560 2351
rect 3574 2347 3576 2351
rect 3590 2347 3592 2351
rect 3595 2347 3597 2351
rect 3611 2347 3613 2351
rect 3210 2301 3214 2303
rect 4155 2301 4159 2303
rect 3069 2291 3071 2295
rect 3074 2291 3076 2295
rect 3090 2291 3092 2295
rect 3106 2291 3108 2295
rect 3111 2291 3113 2295
rect 3132 2291 3134 2295
rect 3148 2291 3150 2295
rect 3164 2291 3166 2295
rect 3169 2291 3171 2295
rect 3185 2291 3187 2295
rect 4014 2291 4016 2295
rect 4019 2291 4021 2295
rect 4035 2291 4037 2295
rect 4051 2291 4053 2295
rect 4056 2291 4058 2295
rect 4077 2291 4079 2295
rect 4093 2291 4095 2295
rect 4109 2291 4111 2295
rect 4114 2291 4116 2295
rect 4130 2291 4132 2295
rect 2286 2261 2288 2265
rect 2291 2261 2293 2265
rect 2307 2261 2309 2265
rect 2323 2261 2325 2265
rect 2328 2261 2330 2265
rect 2349 2261 2351 2265
rect 2365 2261 2367 2265
rect 2381 2261 2383 2265
rect 2386 2261 2388 2265
rect 2402 2261 2404 2265
rect 2418 2261 2420 2265
rect 2423 2261 2425 2265
rect 2439 2261 2441 2265
rect 2455 2261 2457 2265
rect 2460 2261 2462 2265
rect 2481 2261 2483 2265
rect 2497 2261 2499 2265
rect 2513 2261 2515 2265
rect 2518 2261 2520 2265
rect 2534 2261 2536 2265
rect 2550 2261 2552 2265
rect 2555 2261 2557 2265
rect 2571 2261 2573 2265
rect 2587 2261 2589 2265
rect 2592 2261 2594 2265
rect 2613 2261 2615 2265
rect 2629 2261 2631 2265
rect 2645 2261 2647 2265
rect 2650 2261 2652 2265
rect 2666 2261 2668 2265
rect 3231 2261 3233 2265
rect 3236 2261 3238 2265
rect 3252 2261 3254 2265
rect 3268 2261 3270 2265
rect 3273 2261 3275 2265
rect 3294 2261 3296 2265
rect 3310 2261 3312 2265
rect 3326 2261 3328 2265
rect 3331 2261 3333 2265
rect 3347 2261 3349 2265
rect 3363 2261 3365 2265
rect 3368 2261 3370 2265
rect 3384 2261 3386 2265
rect 3400 2261 3402 2265
rect 3405 2261 3407 2265
rect 3426 2261 3428 2265
rect 3442 2261 3444 2265
rect 3458 2261 3460 2265
rect 3463 2261 3465 2265
rect 3479 2261 3481 2265
rect 3495 2261 3497 2265
rect 3500 2261 3502 2265
rect 3516 2261 3518 2265
rect 3532 2261 3534 2265
rect 3537 2261 3539 2265
rect 3558 2261 3560 2265
rect 3574 2261 3576 2265
rect 3590 2261 3592 2265
rect 3595 2261 3597 2265
rect 3611 2261 3613 2265
rect 2518 2217 2520 2221
rect 2542 2217 2544 2221
rect 3463 2217 3465 2221
rect 3487 2217 3489 2221
rect 2538 2206 2540 2210
rect 3483 2206 3485 2210
rect 2529 2192 2533 2194
rect 3474 2192 3478 2194
rect 2518 2183 2520 2187
rect 2542 2183 2544 2187
rect 3463 2183 3465 2187
rect 3487 2183 3489 2187
rect 2286 2121 2288 2125
rect 2291 2121 2293 2125
rect 2307 2121 2309 2125
rect 2323 2121 2325 2125
rect 2328 2121 2330 2125
rect 2349 2121 2351 2125
rect 2365 2121 2367 2125
rect 2381 2121 2383 2125
rect 2386 2121 2388 2125
rect 2402 2121 2404 2125
rect 2418 2121 2420 2125
rect 2423 2121 2425 2125
rect 2439 2121 2441 2125
rect 2455 2121 2457 2125
rect 2460 2121 2462 2125
rect 2481 2121 2483 2125
rect 2497 2121 2499 2125
rect 2513 2121 2515 2125
rect 2518 2121 2520 2125
rect 2534 2121 2536 2125
rect 2550 2121 2552 2125
rect 2555 2121 2557 2125
rect 2571 2121 2573 2125
rect 2587 2121 2589 2125
rect 2592 2121 2594 2125
rect 2613 2121 2615 2125
rect 2629 2121 2631 2125
rect 2645 2121 2647 2125
rect 2650 2121 2652 2125
rect 2666 2121 2668 2125
rect 3231 2121 3233 2125
rect 3236 2121 3238 2125
rect 3252 2121 3254 2125
rect 3268 2121 3270 2125
rect 3273 2121 3275 2125
rect 3294 2121 3296 2125
rect 3310 2121 3312 2125
rect 3326 2121 3328 2125
rect 3331 2121 3333 2125
rect 3347 2121 3349 2125
rect 3363 2121 3365 2125
rect 3368 2121 3370 2125
rect 3384 2121 3386 2125
rect 3400 2121 3402 2125
rect 3405 2121 3407 2125
rect 3426 2121 3428 2125
rect 3442 2121 3444 2125
rect 3458 2121 3460 2125
rect 3463 2121 3465 2125
rect 3479 2121 3481 2125
rect 3495 2121 3497 2125
rect 3500 2121 3502 2125
rect 3516 2121 3518 2125
rect 3532 2121 3534 2125
rect 3537 2121 3539 2125
rect 3558 2121 3560 2125
rect 3574 2121 3576 2125
rect 3590 2121 3592 2125
rect 3595 2121 3597 2125
rect 3611 2121 3613 2125
<< ptransistor >>
rect 2770 4029 2772 4037
rect 2775 4029 2777 4037
rect 2791 4029 2793 4037
rect 2807 4029 2809 4037
rect 2812 4029 2814 4037
rect 2833 4029 2835 4037
rect 2849 4029 2851 4037
rect 2865 4029 2867 4037
rect 2870 4029 2872 4037
rect 2886 4029 2888 4037
rect 2902 4029 2904 4037
rect 2907 4029 2909 4037
rect 2923 4029 2925 4037
rect 2939 4029 2941 4037
rect 2944 4029 2946 4037
rect 2965 4029 2967 4037
rect 2981 4029 2983 4037
rect 2997 4029 2999 4037
rect 3002 4029 3004 4037
rect 3018 4029 3020 4037
rect 3034 4029 3036 4037
rect 3039 4029 3041 4037
rect 3055 4029 3057 4037
rect 3071 4029 3073 4037
rect 3076 4029 3078 4037
rect 3097 4029 3099 4037
rect 3113 4029 3115 4037
rect 3129 4029 3131 4037
rect 3134 4029 3136 4037
rect 3150 4029 3152 4037
rect 3166 4029 3168 4037
rect 3171 4029 3173 4037
rect 3187 4029 3189 4037
rect 3203 4029 3205 4037
rect 3208 4029 3210 4037
rect 3229 4029 3231 4037
rect 3245 4029 3247 4037
rect 3261 4029 3263 4037
rect 3266 4029 3268 4037
rect 3282 4029 3284 4037
rect 3715 4029 3717 4037
rect 3720 4029 3722 4037
rect 3736 4029 3738 4037
rect 3752 4029 3754 4037
rect 3757 4029 3759 4037
rect 3778 4029 3780 4037
rect 3794 4029 3796 4037
rect 3810 4029 3812 4037
rect 3815 4029 3817 4037
rect 3831 4029 3833 4037
rect 3847 4029 3849 4037
rect 3852 4029 3854 4037
rect 3868 4029 3870 4037
rect 3884 4029 3886 4037
rect 3889 4029 3891 4037
rect 3910 4029 3912 4037
rect 3926 4029 3928 4037
rect 3942 4029 3944 4037
rect 3947 4029 3949 4037
rect 3963 4029 3965 4037
rect 3979 4029 3981 4037
rect 3984 4029 3986 4037
rect 4000 4029 4002 4037
rect 4016 4029 4018 4037
rect 4021 4029 4023 4037
rect 4042 4029 4044 4037
rect 4058 4029 4060 4037
rect 4074 4029 4076 4037
rect 4079 4029 4081 4037
rect 4095 4029 4097 4037
rect 4111 4029 4113 4037
rect 4116 4029 4118 4037
rect 4132 4029 4134 4037
rect 4148 4029 4150 4037
rect 4153 4029 4155 4037
rect 4174 4029 4176 4037
rect 4190 4029 4192 4037
rect 4206 4029 4208 4037
rect 4211 4029 4213 4037
rect 4227 4029 4229 4037
rect 2418 3996 2420 4004
rect 2423 3996 2425 4004
rect 2439 3996 2441 4004
rect 2455 3996 2457 4004
rect 2460 3996 2462 4004
rect 2481 3996 2483 4004
rect 2497 3996 2499 4004
rect 2513 3996 2515 4004
rect 2518 3996 2520 4004
rect 2534 3996 2536 4004
rect 3363 3996 3365 4004
rect 3368 3996 3370 4004
rect 3384 3996 3386 4004
rect 3400 3996 3402 4004
rect 3405 3996 3407 4004
rect 3426 3996 3428 4004
rect 3442 3996 3444 4004
rect 3458 3996 3460 4004
rect 3463 3996 3465 4004
rect 3479 3996 3481 4004
rect 2949 3958 2951 3966
rect 2775 3945 2777 3953
rect 2791 3945 2793 3953
rect 2807 3945 2809 3953
rect 2830 3945 2832 3953
rect 2835 3945 2837 3953
rect 2861 3945 2863 3953
rect 2882 3945 2884 3953
rect 2902 3945 2904 3953
rect 2907 3945 2909 3953
rect 2925 3945 2927 3953
rect 2975 3952 2977 3960
rect 2980 3952 2982 3960
rect 3003 3958 3005 3966
rect 3030 3958 3032 3966
rect 3056 3952 3058 3960
rect 3061 3952 3063 3960
rect 3084 3958 3086 3966
rect 3894 3958 3896 3966
rect 3720 3945 3722 3953
rect 3736 3945 3738 3953
rect 3752 3945 3754 3953
rect 3775 3945 3777 3953
rect 3780 3945 3782 3953
rect 3806 3945 3808 3953
rect 3827 3945 3829 3953
rect 3847 3945 3849 3953
rect 3852 3945 3854 3953
rect 3870 3945 3872 3953
rect 3920 3952 3922 3960
rect 3925 3952 3927 3960
rect 3948 3958 3950 3966
rect 3975 3958 3977 3966
rect 4001 3952 4003 3960
rect 4006 3952 4008 3960
rect 4029 3958 4031 3966
rect 2409 3894 2411 3902
rect 2425 3894 2427 3902
rect 2430 3894 2432 3902
rect 2446 3894 2448 3902
rect 2462 3894 2464 3902
rect 2483 3894 2485 3902
rect 2488 3894 2490 3902
rect 2504 3894 2506 3902
rect 2520 3894 2522 3902
rect 2525 3894 2527 3902
rect 3354 3894 3356 3902
rect 3370 3894 3372 3902
rect 3375 3894 3377 3902
rect 3391 3894 3393 3902
rect 3407 3894 3409 3902
rect 3428 3894 3430 3902
rect 3433 3894 3435 3902
rect 3449 3894 3451 3902
rect 3465 3894 3467 3902
rect 3470 3894 3472 3902
rect 2775 3859 2777 3867
rect 2791 3859 2793 3867
rect 2807 3859 2809 3867
rect 2830 3859 2832 3867
rect 2835 3859 2837 3867
rect 2861 3859 2863 3867
rect 2882 3859 2884 3867
rect 2902 3859 2904 3867
rect 2907 3859 2909 3867
rect 2925 3859 2927 3867
rect 2975 3860 2977 3868
rect 2980 3860 2982 3868
rect 3056 3860 3058 3868
rect 3061 3860 3063 3868
rect 3720 3859 3722 3867
rect 3736 3859 3738 3867
rect 3752 3859 3754 3867
rect 3775 3859 3777 3867
rect 3780 3859 3782 3867
rect 3806 3859 3808 3867
rect 3827 3859 3829 3867
rect 3847 3859 3849 3867
rect 3852 3859 3854 3867
rect 3870 3859 3872 3867
rect 3920 3860 3922 3868
rect 3925 3860 3927 3868
rect 4001 3860 4003 3868
rect 4006 3860 4008 3868
rect 2775 3813 2777 3821
rect 2791 3813 2793 3821
rect 2807 3813 2809 3821
rect 2830 3813 2832 3821
rect 2835 3813 2837 3821
rect 2861 3813 2863 3821
rect 2882 3813 2884 3821
rect 2902 3813 2904 3821
rect 2907 3813 2909 3821
rect 2925 3813 2927 3821
rect 2975 3820 2977 3828
rect 2980 3820 2982 3828
rect 3003 3826 3005 3834
rect 3054 3826 3056 3834
rect 3080 3820 3082 3828
rect 3085 3820 3087 3828
rect 3108 3826 3110 3834
rect 3720 3813 3722 3821
rect 3736 3813 3738 3821
rect 3752 3813 3754 3821
rect 3775 3813 3777 3821
rect 3780 3813 3782 3821
rect 3806 3813 3808 3821
rect 3827 3813 3829 3821
rect 3847 3813 3849 3821
rect 3852 3813 3854 3821
rect 3870 3813 3872 3821
rect 3920 3820 3922 3828
rect 3925 3820 3927 3828
rect 3948 3826 3950 3834
rect 3999 3826 4001 3834
rect 3285 3797 3287 3805
rect 3311 3791 3313 3799
rect 3316 3791 3318 3799
rect 3339 3797 3341 3805
rect 3471 3772 3473 3802
rect 3524 3772 3526 3802
rect 4025 3820 4027 3828
rect 4030 3820 4032 3828
rect 4053 3826 4055 3834
rect 2775 3727 2777 3735
rect 2791 3727 2793 3735
rect 2807 3727 2809 3735
rect 2830 3727 2832 3735
rect 2835 3727 2837 3735
rect 2861 3727 2863 3735
rect 2882 3727 2884 3735
rect 2902 3727 2904 3735
rect 2907 3727 2909 3735
rect 2925 3727 2927 3735
rect 2975 3729 2977 3737
rect 2980 3729 2982 3737
rect 3080 3729 3082 3737
rect 3085 3729 3087 3737
rect 3720 3727 3722 3735
rect 3736 3727 3738 3735
rect 3752 3727 3754 3735
rect 3775 3727 3777 3735
rect 3780 3727 3782 3735
rect 3806 3727 3808 3735
rect 3827 3727 3829 3735
rect 3847 3727 3849 3735
rect 3852 3727 3854 3735
rect 3870 3727 3872 3735
rect 3920 3729 3922 3737
rect 3925 3729 3927 3737
rect 4025 3729 4027 3737
rect 4030 3729 4032 3737
rect 2775 3681 2777 3689
rect 2791 3681 2793 3689
rect 2807 3681 2809 3689
rect 2830 3681 2832 3689
rect 2835 3681 2837 3689
rect 2861 3681 2863 3689
rect 2882 3681 2884 3689
rect 2902 3681 2904 3689
rect 2907 3681 2909 3689
rect 2925 3681 2927 3689
rect 2975 3688 2977 3696
rect 2980 3688 2982 3696
rect 3003 3694 3005 3702
rect 3030 3694 3032 3702
rect 3056 3688 3058 3696
rect 3061 3688 3063 3696
rect 3084 3694 3086 3702
rect 3120 3694 3122 3702
rect 3146 3688 3148 3696
rect 3151 3688 3153 3696
rect 3174 3694 3176 3702
rect 3311 3695 3313 3703
rect 3316 3695 3318 3703
rect 3720 3681 3722 3689
rect 3736 3681 3738 3689
rect 3752 3681 3754 3689
rect 3775 3681 3777 3689
rect 3780 3681 3782 3689
rect 3806 3681 3808 3689
rect 3827 3681 3829 3689
rect 3847 3681 3849 3689
rect 3852 3681 3854 3689
rect 3870 3681 3872 3689
rect 3920 3688 3922 3696
rect 3925 3688 3927 3696
rect 3948 3694 3950 3702
rect 3975 3694 3977 3702
rect 3263 3667 3265 3675
rect 3285 3667 3287 3675
rect 3311 3661 3313 3669
rect 3316 3661 3318 3669
rect 3339 3667 3341 3675
rect 3377 3642 3379 3672
rect 3430 3642 3432 3672
rect 4001 3688 4003 3696
rect 4006 3688 4008 3696
rect 4029 3694 4031 3702
rect 4065 3694 4067 3702
rect 4091 3688 4093 3696
rect 4096 3688 4098 3696
rect 4119 3694 4121 3702
rect 2775 3595 2777 3603
rect 2791 3595 2793 3603
rect 2807 3595 2809 3603
rect 2830 3595 2832 3603
rect 2835 3595 2837 3603
rect 2861 3595 2863 3603
rect 2882 3595 2884 3603
rect 2902 3595 2904 3603
rect 2907 3595 2909 3603
rect 2925 3595 2927 3603
rect 2975 3594 2977 3602
rect 2980 3594 2982 3602
rect 3056 3594 3058 3602
rect 3061 3594 3063 3602
rect 3146 3594 3148 3602
rect 3151 3594 3153 3602
rect 3720 3595 3722 3603
rect 3736 3595 3738 3603
rect 3752 3595 3754 3603
rect 3775 3595 3777 3603
rect 3780 3595 3782 3603
rect 3806 3595 3808 3603
rect 3827 3595 3829 3603
rect 3847 3595 3849 3603
rect 3852 3595 3854 3603
rect 3870 3595 3872 3603
rect 3920 3594 3922 3602
rect 3925 3594 3927 3602
rect 4001 3594 4003 3602
rect 4006 3594 4008 3602
rect 4091 3594 4093 3602
rect 4096 3594 4098 3602
rect 2775 3549 2777 3557
rect 2791 3549 2793 3557
rect 2807 3549 2809 3557
rect 2830 3549 2832 3557
rect 2835 3549 2837 3557
rect 2861 3549 2863 3557
rect 2882 3549 2884 3557
rect 2902 3549 2904 3557
rect 2907 3549 2909 3557
rect 2925 3549 2927 3557
rect 2975 3556 2977 3564
rect 2980 3556 2982 3564
rect 3003 3562 3005 3570
rect 3311 3565 3313 3573
rect 3316 3565 3318 3573
rect 3720 3549 3722 3557
rect 3736 3549 3738 3557
rect 3752 3549 3754 3557
rect 3775 3549 3777 3557
rect 3780 3549 3782 3557
rect 3806 3549 3808 3557
rect 3827 3549 3829 3557
rect 3847 3549 3849 3557
rect 3852 3549 3854 3557
rect 3870 3549 3872 3557
rect 3920 3556 3922 3564
rect 3925 3556 3927 3564
rect 3948 3562 3950 3570
rect 2286 3494 2288 3502
rect 2291 3494 2293 3502
rect 2307 3494 2309 3502
rect 2323 3494 2325 3502
rect 2328 3494 2330 3502
rect 2349 3494 2351 3502
rect 2365 3494 2367 3502
rect 2381 3494 2383 3502
rect 2386 3494 2388 3502
rect 2402 3494 2404 3502
rect 2418 3494 2420 3502
rect 2423 3494 2425 3502
rect 2439 3494 2441 3502
rect 2455 3494 2457 3502
rect 2460 3494 2462 3502
rect 2481 3494 2483 3502
rect 2497 3494 2499 3502
rect 2513 3494 2515 3502
rect 2518 3494 2520 3502
rect 2534 3494 2536 3502
rect 2550 3494 2552 3502
rect 2555 3494 2557 3502
rect 2571 3494 2573 3502
rect 2587 3494 2589 3502
rect 2592 3494 2594 3502
rect 2613 3494 2615 3502
rect 2629 3494 2631 3502
rect 2645 3494 2647 3502
rect 2650 3494 2652 3502
rect 2666 3494 2668 3502
rect 3231 3494 3233 3502
rect 3236 3494 3238 3502
rect 3252 3494 3254 3502
rect 3268 3494 3270 3502
rect 3273 3494 3275 3502
rect 3294 3494 3296 3502
rect 3310 3494 3312 3502
rect 3326 3494 3328 3502
rect 3331 3494 3333 3502
rect 3347 3494 3349 3502
rect 3363 3494 3365 3502
rect 3368 3494 3370 3502
rect 3384 3494 3386 3502
rect 3400 3494 3402 3502
rect 3405 3494 3407 3502
rect 3426 3494 3428 3502
rect 3442 3494 3444 3502
rect 3458 3494 3460 3502
rect 3463 3494 3465 3502
rect 3479 3494 3481 3502
rect 3495 3494 3497 3502
rect 3500 3494 3502 3502
rect 3516 3494 3518 3502
rect 3532 3494 3534 3502
rect 3537 3494 3539 3502
rect 3558 3494 3560 3502
rect 3574 3494 3576 3502
rect 3590 3494 3592 3502
rect 3595 3494 3597 3502
rect 3611 3494 3613 3502
rect 2775 3463 2777 3471
rect 2791 3463 2793 3471
rect 2807 3463 2809 3471
rect 2830 3463 2832 3471
rect 2835 3463 2837 3471
rect 2861 3463 2863 3471
rect 2882 3463 2884 3471
rect 2902 3463 2904 3471
rect 2907 3463 2909 3471
rect 2925 3463 2927 3471
rect 2975 3458 2977 3466
rect 2980 3458 2982 3466
rect 3009 3463 3011 3471
rect 3027 3463 3029 3471
rect 3052 3463 3054 3471
rect 3068 3463 3070 3471
rect 3091 3463 3093 3471
rect 3096 3463 3098 3471
rect 3122 3463 3124 3471
rect 3143 3463 3145 3471
rect 3163 3463 3165 3471
rect 3168 3463 3170 3471
rect 3186 3463 3188 3471
rect 3720 3463 3722 3471
rect 3736 3463 3738 3471
rect 3752 3463 3754 3471
rect 3775 3463 3777 3471
rect 3780 3463 3782 3471
rect 3806 3463 3808 3471
rect 3827 3463 3829 3471
rect 3847 3463 3849 3471
rect 3852 3463 3854 3471
rect 3870 3463 3872 3471
rect 3920 3458 3922 3466
rect 3925 3458 3927 3466
rect 3954 3463 3956 3471
rect 3972 3463 3974 3471
rect 3997 3463 3999 3471
rect 4013 3463 4015 3471
rect 4036 3463 4038 3471
rect 4041 3463 4043 3471
rect 4067 3463 4069 3471
rect 4088 3463 4090 3471
rect 4108 3463 4110 3471
rect 4113 3463 4115 3471
rect 4131 3463 4133 3471
rect 3069 3382 3071 3390
rect 3074 3382 3076 3390
rect 3090 3382 3092 3390
rect 3106 3382 3108 3390
rect 3111 3382 3113 3390
rect 3132 3382 3134 3390
rect 3148 3382 3150 3390
rect 3164 3382 3166 3390
rect 3169 3382 3171 3390
rect 3185 3382 3187 3390
rect 4014 3382 4016 3390
rect 4019 3382 4021 3390
rect 4035 3382 4037 3390
rect 4051 3382 4053 3390
rect 4056 3382 4058 3390
rect 4077 3382 4079 3390
rect 4093 3382 4095 3390
rect 4109 3382 4111 3390
rect 4114 3382 4116 3390
rect 4130 3382 4132 3390
rect 2286 3352 2288 3360
rect 2291 3352 2293 3360
rect 2307 3352 2309 3360
rect 2323 3352 2325 3360
rect 2328 3352 2330 3360
rect 2349 3352 2351 3360
rect 2365 3352 2367 3360
rect 2381 3352 2383 3360
rect 2386 3352 2388 3360
rect 2402 3352 2404 3360
rect 2418 3352 2420 3360
rect 2423 3352 2425 3360
rect 2439 3352 2441 3360
rect 2455 3352 2457 3360
rect 2460 3352 2462 3360
rect 2481 3352 2483 3360
rect 2497 3352 2499 3360
rect 2513 3352 2515 3360
rect 2518 3352 2520 3360
rect 2534 3352 2536 3360
rect 2550 3352 2552 3360
rect 2555 3352 2557 3360
rect 2571 3352 2573 3360
rect 2587 3352 2589 3360
rect 2592 3352 2594 3360
rect 2613 3352 2615 3360
rect 2629 3352 2631 3360
rect 2645 3352 2647 3360
rect 2650 3352 2652 3360
rect 2666 3352 2668 3360
rect 3231 3352 3233 3360
rect 3236 3352 3238 3360
rect 3252 3352 3254 3360
rect 3268 3352 3270 3360
rect 3273 3352 3275 3360
rect 3294 3352 3296 3360
rect 3310 3352 3312 3360
rect 3326 3352 3328 3360
rect 3331 3352 3333 3360
rect 3347 3352 3349 3360
rect 3363 3352 3365 3360
rect 3368 3352 3370 3360
rect 3384 3352 3386 3360
rect 3400 3352 3402 3360
rect 3405 3352 3407 3360
rect 3426 3352 3428 3360
rect 3442 3352 3444 3360
rect 3458 3352 3460 3360
rect 3463 3352 3465 3360
rect 3479 3352 3481 3360
rect 3495 3352 3497 3360
rect 3500 3352 3502 3360
rect 3516 3352 3518 3360
rect 3532 3352 3534 3360
rect 3537 3352 3539 3360
rect 3558 3352 3560 3360
rect 3574 3352 3576 3360
rect 3590 3352 3592 3360
rect 3595 3352 3597 3360
rect 3611 3352 3613 3360
rect 3069 3296 3071 3304
rect 3074 3296 3076 3304
rect 3090 3296 3092 3304
rect 3106 3296 3108 3304
rect 3111 3296 3113 3304
rect 3132 3296 3134 3304
rect 3148 3296 3150 3304
rect 3164 3296 3166 3304
rect 3169 3296 3171 3304
rect 3185 3296 3187 3304
rect 4014 3296 4016 3304
rect 4019 3296 4021 3304
rect 4035 3296 4037 3304
rect 4051 3296 4053 3304
rect 4056 3296 4058 3304
rect 4077 3296 4079 3304
rect 4093 3296 4095 3304
rect 4109 3296 4111 3304
rect 4114 3296 4116 3304
rect 4130 3296 4132 3304
rect 2286 3266 2288 3274
rect 2291 3266 2293 3274
rect 2307 3266 2309 3274
rect 2323 3266 2325 3274
rect 2328 3266 2330 3274
rect 2349 3266 2351 3274
rect 2365 3266 2367 3274
rect 2381 3266 2383 3274
rect 2386 3266 2388 3274
rect 2402 3266 2404 3274
rect 2418 3266 2420 3274
rect 2423 3266 2425 3274
rect 2439 3266 2441 3274
rect 2455 3266 2457 3274
rect 2460 3266 2462 3274
rect 2481 3266 2483 3274
rect 2497 3266 2499 3274
rect 2513 3266 2515 3274
rect 2518 3266 2520 3274
rect 2534 3266 2536 3274
rect 2550 3266 2552 3274
rect 2555 3266 2557 3274
rect 2571 3266 2573 3274
rect 2587 3266 2589 3274
rect 2592 3266 2594 3274
rect 2613 3266 2615 3274
rect 2629 3266 2631 3274
rect 2645 3266 2647 3274
rect 2650 3266 2652 3274
rect 2666 3266 2668 3274
rect 3231 3266 3233 3274
rect 3236 3266 3238 3274
rect 3252 3266 3254 3274
rect 3268 3266 3270 3274
rect 3273 3266 3275 3274
rect 3294 3266 3296 3274
rect 3310 3266 3312 3274
rect 3326 3266 3328 3274
rect 3331 3266 3333 3274
rect 3347 3266 3349 3274
rect 3363 3266 3365 3274
rect 3368 3266 3370 3274
rect 3384 3266 3386 3274
rect 3400 3266 3402 3274
rect 3405 3266 3407 3274
rect 3426 3266 3428 3274
rect 3442 3266 3444 3274
rect 3458 3266 3460 3274
rect 3463 3266 3465 3274
rect 3479 3266 3481 3274
rect 3495 3266 3497 3274
rect 3500 3266 3502 3274
rect 3516 3266 3518 3274
rect 3532 3266 3534 3274
rect 3537 3266 3539 3274
rect 3558 3266 3560 3274
rect 3574 3266 3576 3274
rect 3590 3266 3592 3274
rect 3595 3266 3597 3274
rect 3611 3266 3613 3274
rect 2286 3126 2288 3134
rect 2291 3126 2293 3134
rect 2307 3126 2309 3134
rect 2323 3126 2325 3134
rect 2328 3126 2330 3134
rect 2349 3126 2351 3134
rect 2365 3126 2367 3134
rect 2381 3126 2383 3134
rect 2386 3126 2388 3134
rect 2402 3126 2404 3134
rect 2418 3126 2420 3134
rect 2423 3126 2425 3134
rect 2439 3126 2441 3134
rect 2455 3126 2457 3134
rect 2460 3126 2462 3134
rect 2481 3126 2483 3134
rect 2497 3126 2499 3134
rect 2513 3126 2515 3134
rect 2518 3126 2520 3134
rect 2534 3126 2536 3134
rect 2550 3126 2552 3134
rect 2555 3126 2557 3134
rect 2571 3126 2573 3134
rect 2587 3126 2589 3134
rect 2592 3126 2594 3134
rect 2613 3126 2615 3134
rect 2629 3126 2631 3134
rect 2645 3126 2647 3134
rect 2650 3126 2652 3134
rect 2666 3126 2668 3134
rect 3231 3126 3233 3134
rect 3236 3126 3238 3134
rect 3252 3126 3254 3134
rect 3268 3126 3270 3134
rect 3273 3126 3275 3134
rect 3294 3126 3296 3134
rect 3310 3126 3312 3134
rect 3326 3126 3328 3134
rect 3331 3126 3333 3134
rect 3347 3126 3349 3134
rect 3363 3126 3365 3134
rect 3368 3126 3370 3134
rect 3384 3126 3386 3134
rect 3400 3126 3402 3134
rect 3405 3126 3407 3134
rect 3426 3126 3428 3134
rect 3442 3126 3444 3134
rect 3458 3126 3460 3134
rect 3463 3126 3465 3134
rect 3479 3126 3481 3134
rect 3495 3126 3497 3134
rect 3500 3126 3502 3134
rect 3516 3126 3518 3134
rect 3532 3126 3534 3134
rect 3537 3126 3539 3134
rect 3558 3126 3560 3134
rect 3574 3126 3576 3134
rect 3590 3126 3592 3134
rect 3595 3126 3597 3134
rect 3611 3126 3613 3134
rect 2770 3047 2772 3055
rect 2775 3047 2777 3055
rect 2791 3047 2793 3055
rect 2807 3047 2809 3055
rect 2812 3047 2814 3055
rect 2833 3047 2835 3055
rect 2849 3047 2851 3055
rect 2865 3047 2867 3055
rect 2870 3047 2872 3055
rect 2886 3047 2888 3055
rect 2902 3047 2904 3055
rect 2907 3047 2909 3055
rect 2923 3047 2925 3055
rect 2939 3047 2941 3055
rect 2944 3047 2946 3055
rect 2965 3047 2967 3055
rect 2981 3047 2983 3055
rect 2997 3047 2999 3055
rect 3002 3047 3004 3055
rect 3018 3047 3020 3055
rect 3034 3047 3036 3055
rect 3039 3047 3041 3055
rect 3055 3047 3057 3055
rect 3071 3047 3073 3055
rect 3076 3047 3078 3055
rect 3097 3047 3099 3055
rect 3113 3047 3115 3055
rect 3129 3047 3131 3055
rect 3134 3047 3136 3055
rect 3150 3047 3152 3055
rect 3166 3047 3168 3055
rect 3171 3047 3173 3055
rect 3187 3047 3189 3055
rect 3203 3047 3205 3055
rect 3208 3047 3210 3055
rect 3229 3047 3231 3055
rect 3245 3047 3247 3055
rect 3261 3047 3263 3055
rect 3266 3047 3268 3055
rect 3282 3047 3284 3055
rect 3715 3047 3717 3055
rect 3720 3047 3722 3055
rect 3736 3047 3738 3055
rect 3752 3047 3754 3055
rect 3757 3047 3759 3055
rect 3778 3047 3780 3055
rect 3794 3047 3796 3055
rect 3810 3047 3812 3055
rect 3815 3047 3817 3055
rect 3831 3047 3833 3055
rect 3847 3047 3849 3055
rect 3852 3047 3854 3055
rect 3868 3047 3870 3055
rect 3884 3047 3886 3055
rect 3889 3047 3891 3055
rect 3910 3047 3912 3055
rect 3926 3047 3928 3055
rect 3942 3047 3944 3055
rect 3947 3047 3949 3055
rect 3963 3047 3965 3055
rect 3979 3047 3981 3055
rect 3984 3047 3986 3055
rect 4000 3047 4002 3055
rect 4016 3047 4018 3055
rect 4021 3047 4023 3055
rect 4042 3047 4044 3055
rect 4058 3047 4060 3055
rect 4074 3047 4076 3055
rect 4079 3047 4081 3055
rect 4095 3047 4097 3055
rect 4111 3047 4113 3055
rect 4116 3047 4118 3055
rect 4132 3047 4134 3055
rect 4148 3047 4150 3055
rect 4153 3047 4155 3055
rect 4174 3047 4176 3055
rect 4190 3047 4192 3055
rect 4206 3047 4208 3055
rect 4211 3047 4213 3055
rect 4227 3047 4229 3055
rect 2418 3014 2420 3022
rect 2423 3014 2425 3022
rect 2439 3014 2441 3022
rect 2455 3014 2457 3022
rect 2460 3014 2462 3022
rect 2481 3014 2483 3022
rect 2497 3014 2499 3022
rect 2513 3014 2515 3022
rect 2518 3014 2520 3022
rect 2534 3014 2536 3022
rect 3363 3014 3365 3022
rect 3368 3014 3370 3022
rect 3384 3014 3386 3022
rect 3400 3014 3402 3022
rect 3405 3014 3407 3022
rect 3426 3014 3428 3022
rect 3442 3014 3444 3022
rect 3458 3014 3460 3022
rect 3463 3014 3465 3022
rect 3479 3014 3481 3022
rect 2949 2976 2951 2984
rect 2775 2963 2777 2971
rect 2791 2963 2793 2971
rect 2807 2963 2809 2971
rect 2830 2963 2832 2971
rect 2835 2963 2837 2971
rect 2861 2963 2863 2971
rect 2882 2963 2884 2971
rect 2902 2963 2904 2971
rect 2907 2963 2909 2971
rect 2925 2963 2927 2971
rect 2975 2970 2977 2978
rect 2980 2970 2982 2978
rect 3003 2976 3005 2984
rect 3030 2976 3032 2984
rect 3056 2970 3058 2978
rect 3061 2970 3063 2978
rect 3084 2976 3086 2984
rect 3894 2976 3896 2984
rect 3720 2963 3722 2971
rect 3736 2963 3738 2971
rect 3752 2963 3754 2971
rect 3775 2963 3777 2971
rect 3780 2963 3782 2971
rect 3806 2963 3808 2971
rect 3827 2963 3829 2971
rect 3847 2963 3849 2971
rect 3852 2963 3854 2971
rect 3870 2963 3872 2971
rect 3920 2970 3922 2978
rect 3925 2970 3927 2978
rect 3948 2976 3950 2984
rect 3975 2976 3977 2984
rect 4001 2970 4003 2978
rect 4006 2970 4008 2978
rect 4029 2976 4031 2984
rect 2409 2912 2411 2920
rect 2425 2912 2427 2920
rect 2430 2912 2432 2920
rect 2446 2912 2448 2920
rect 2462 2912 2464 2920
rect 2483 2912 2485 2920
rect 2488 2912 2490 2920
rect 2504 2912 2506 2920
rect 2520 2912 2522 2920
rect 2525 2912 2527 2920
rect 3354 2912 3356 2920
rect 3370 2912 3372 2920
rect 3375 2912 3377 2920
rect 3391 2912 3393 2920
rect 3407 2912 3409 2920
rect 3428 2912 3430 2920
rect 3433 2912 3435 2920
rect 3449 2912 3451 2920
rect 3465 2912 3467 2920
rect 3470 2912 3472 2920
rect 2775 2877 2777 2885
rect 2791 2877 2793 2885
rect 2807 2877 2809 2885
rect 2830 2877 2832 2885
rect 2835 2877 2837 2885
rect 2861 2877 2863 2885
rect 2882 2877 2884 2885
rect 2902 2877 2904 2885
rect 2907 2877 2909 2885
rect 2925 2877 2927 2885
rect 2975 2878 2977 2886
rect 2980 2878 2982 2886
rect 3056 2878 3058 2886
rect 3061 2878 3063 2886
rect 3720 2877 3722 2885
rect 3736 2877 3738 2885
rect 3752 2877 3754 2885
rect 3775 2877 3777 2885
rect 3780 2877 3782 2885
rect 3806 2877 3808 2885
rect 3827 2877 3829 2885
rect 3847 2877 3849 2885
rect 3852 2877 3854 2885
rect 3870 2877 3872 2885
rect 3920 2878 3922 2886
rect 3925 2878 3927 2886
rect 4001 2878 4003 2886
rect 4006 2878 4008 2886
rect 2775 2831 2777 2839
rect 2791 2831 2793 2839
rect 2807 2831 2809 2839
rect 2830 2831 2832 2839
rect 2835 2831 2837 2839
rect 2861 2831 2863 2839
rect 2882 2831 2884 2839
rect 2902 2831 2904 2839
rect 2907 2831 2909 2839
rect 2925 2831 2927 2839
rect 2975 2838 2977 2846
rect 2980 2838 2982 2846
rect 3003 2844 3005 2852
rect 3054 2844 3056 2852
rect 3080 2838 3082 2846
rect 3085 2838 3087 2846
rect 3108 2844 3110 2852
rect 3720 2831 3722 2839
rect 3736 2831 3738 2839
rect 3752 2831 3754 2839
rect 3775 2831 3777 2839
rect 3780 2831 3782 2839
rect 3806 2831 3808 2839
rect 3827 2831 3829 2839
rect 3847 2831 3849 2839
rect 3852 2831 3854 2839
rect 3870 2831 3872 2839
rect 3920 2838 3922 2846
rect 3925 2838 3927 2846
rect 3948 2844 3950 2852
rect 3999 2844 4001 2852
rect 4025 2838 4027 2846
rect 4030 2838 4032 2846
rect 4053 2844 4055 2852
rect 2775 2745 2777 2753
rect 2791 2745 2793 2753
rect 2807 2745 2809 2753
rect 2830 2745 2832 2753
rect 2835 2745 2837 2753
rect 2861 2745 2863 2753
rect 2882 2745 2884 2753
rect 2902 2745 2904 2753
rect 2907 2745 2909 2753
rect 2925 2745 2927 2753
rect 2975 2747 2977 2755
rect 2980 2747 2982 2755
rect 3080 2747 3082 2755
rect 3085 2747 3087 2755
rect 3720 2745 3722 2753
rect 3736 2745 3738 2753
rect 3752 2745 3754 2753
rect 3775 2745 3777 2753
rect 3780 2745 3782 2753
rect 3806 2745 3808 2753
rect 3827 2745 3829 2753
rect 3847 2745 3849 2753
rect 3852 2745 3854 2753
rect 3870 2745 3872 2753
rect 3920 2747 3922 2755
rect 3925 2747 3927 2755
rect 4025 2747 4027 2755
rect 4030 2747 4032 2755
rect 2775 2699 2777 2707
rect 2791 2699 2793 2707
rect 2807 2699 2809 2707
rect 2830 2699 2832 2707
rect 2835 2699 2837 2707
rect 2861 2699 2863 2707
rect 2882 2699 2884 2707
rect 2902 2699 2904 2707
rect 2907 2699 2909 2707
rect 2925 2699 2927 2707
rect 2975 2706 2977 2714
rect 2980 2706 2982 2714
rect 3003 2712 3005 2720
rect 3030 2712 3032 2720
rect 3056 2706 3058 2714
rect 3061 2706 3063 2714
rect 3084 2712 3086 2720
rect 3120 2712 3122 2720
rect 3146 2706 3148 2714
rect 3151 2706 3153 2714
rect 3174 2712 3176 2720
rect 3720 2699 3722 2707
rect 3736 2699 3738 2707
rect 3752 2699 3754 2707
rect 3775 2699 3777 2707
rect 3780 2699 3782 2707
rect 3806 2699 3808 2707
rect 3827 2699 3829 2707
rect 3847 2699 3849 2707
rect 3852 2699 3854 2707
rect 3870 2699 3872 2707
rect 3920 2706 3922 2714
rect 3925 2706 3927 2714
rect 3948 2712 3950 2720
rect 3975 2712 3977 2720
rect 4001 2706 4003 2714
rect 4006 2706 4008 2714
rect 4029 2712 4031 2720
rect 4065 2712 4067 2720
rect 4091 2706 4093 2714
rect 4096 2706 4098 2714
rect 4119 2712 4121 2720
rect 2775 2613 2777 2621
rect 2791 2613 2793 2621
rect 2807 2613 2809 2621
rect 2830 2613 2832 2621
rect 2835 2613 2837 2621
rect 2861 2613 2863 2621
rect 2882 2613 2884 2621
rect 2902 2613 2904 2621
rect 2907 2613 2909 2621
rect 2925 2613 2927 2621
rect 2975 2612 2977 2620
rect 2980 2612 2982 2620
rect 3056 2612 3058 2620
rect 3061 2612 3063 2620
rect 3146 2612 3148 2620
rect 3151 2612 3153 2620
rect 3720 2613 3722 2621
rect 3736 2613 3738 2621
rect 3752 2613 3754 2621
rect 3775 2613 3777 2621
rect 3780 2613 3782 2621
rect 3806 2613 3808 2621
rect 3827 2613 3829 2621
rect 3847 2613 3849 2621
rect 3852 2613 3854 2621
rect 3870 2613 3872 2621
rect 3920 2612 3922 2620
rect 3925 2612 3927 2620
rect 4001 2612 4003 2620
rect 4006 2612 4008 2620
rect 4091 2612 4093 2620
rect 4096 2612 4098 2620
rect 2775 2567 2777 2575
rect 2791 2567 2793 2575
rect 2807 2567 2809 2575
rect 2830 2567 2832 2575
rect 2835 2567 2837 2575
rect 2861 2567 2863 2575
rect 2882 2567 2884 2575
rect 2902 2567 2904 2575
rect 2907 2567 2909 2575
rect 2925 2567 2927 2575
rect 2975 2574 2977 2582
rect 2980 2574 2982 2582
rect 3003 2580 3005 2588
rect 3720 2567 3722 2575
rect 3736 2567 3738 2575
rect 3752 2567 3754 2575
rect 3775 2567 3777 2575
rect 3780 2567 3782 2575
rect 3806 2567 3808 2575
rect 3827 2567 3829 2575
rect 3847 2567 3849 2575
rect 3852 2567 3854 2575
rect 3870 2567 3872 2575
rect 3920 2574 3922 2582
rect 3925 2574 3927 2582
rect 3948 2580 3950 2588
rect 2286 2512 2288 2520
rect 2291 2512 2293 2520
rect 2307 2512 2309 2520
rect 2323 2512 2325 2520
rect 2328 2512 2330 2520
rect 2349 2512 2351 2520
rect 2365 2512 2367 2520
rect 2381 2512 2383 2520
rect 2386 2512 2388 2520
rect 2402 2512 2404 2520
rect 2418 2512 2420 2520
rect 2423 2512 2425 2520
rect 2439 2512 2441 2520
rect 2455 2512 2457 2520
rect 2460 2512 2462 2520
rect 2481 2512 2483 2520
rect 2497 2512 2499 2520
rect 2513 2512 2515 2520
rect 2518 2512 2520 2520
rect 2534 2512 2536 2520
rect 2550 2512 2552 2520
rect 2555 2512 2557 2520
rect 2571 2512 2573 2520
rect 2587 2512 2589 2520
rect 2592 2512 2594 2520
rect 2613 2512 2615 2520
rect 2629 2512 2631 2520
rect 2645 2512 2647 2520
rect 2650 2512 2652 2520
rect 2666 2512 2668 2520
rect 3231 2512 3233 2520
rect 3236 2512 3238 2520
rect 3252 2512 3254 2520
rect 3268 2512 3270 2520
rect 3273 2512 3275 2520
rect 3294 2512 3296 2520
rect 3310 2512 3312 2520
rect 3326 2512 3328 2520
rect 3331 2512 3333 2520
rect 3347 2512 3349 2520
rect 3363 2512 3365 2520
rect 3368 2512 3370 2520
rect 3384 2512 3386 2520
rect 3400 2512 3402 2520
rect 3405 2512 3407 2520
rect 3426 2512 3428 2520
rect 3442 2512 3444 2520
rect 3458 2512 3460 2520
rect 3463 2512 3465 2520
rect 3479 2512 3481 2520
rect 3495 2512 3497 2520
rect 3500 2512 3502 2520
rect 3516 2512 3518 2520
rect 3532 2512 3534 2520
rect 3537 2512 3539 2520
rect 3558 2512 3560 2520
rect 3574 2512 3576 2520
rect 3590 2512 3592 2520
rect 3595 2512 3597 2520
rect 3611 2512 3613 2520
rect 2775 2481 2777 2489
rect 2791 2481 2793 2489
rect 2807 2481 2809 2489
rect 2830 2481 2832 2489
rect 2835 2481 2837 2489
rect 2861 2481 2863 2489
rect 2882 2481 2884 2489
rect 2902 2481 2904 2489
rect 2907 2481 2909 2489
rect 2925 2481 2927 2489
rect 2975 2476 2977 2484
rect 2980 2476 2982 2484
rect 3009 2481 3011 2489
rect 3027 2481 3029 2489
rect 3052 2481 3054 2489
rect 3068 2481 3070 2489
rect 3091 2481 3093 2489
rect 3096 2481 3098 2489
rect 3122 2481 3124 2489
rect 3143 2481 3145 2489
rect 3163 2481 3165 2489
rect 3168 2481 3170 2489
rect 3186 2481 3188 2489
rect 3720 2481 3722 2489
rect 3736 2481 3738 2489
rect 3752 2481 3754 2489
rect 3775 2481 3777 2489
rect 3780 2481 3782 2489
rect 3806 2481 3808 2489
rect 3827 2481 3829 2489
rect 3847 2481 3849 2489
rect 3852 2481 3854 2489
rect 3870 2481 3872 2489
rect 3920 2476 3922 2484
rect 3925 2476 3927 2484
rect 3954 2481 3956 2489
rect 3972 2481 3974 2489
rect 3997 2481 3999 2489
rect 4013 2481 4015 2489
rect 4036 2481 4038 2489
rect 4041 2481 4043 2489
rect 4067 2481 4069 2489
rect 4088 2481 4090 2489
rect 4108 2481 4110 2489
rect 4113 2481 4115 2489
rect 4131 2481 4133 2489
rect 3069 2400 3071 2408
rect 3074 2400 3076 2408
rect 3090 2400 3092 2408
rect 3106 2400 3108 2408
rect 3111 2400 3113 2408
rect 3132 2400 3134 2408
rect 3148 2400 3150 2408
rect 3164 2400 3166 2408
rect 3169 2400 3171 2408
rect 3185 2400 3187 2408
rect 4014 2400 4016 2408
rect 4019 2400 4021 2408
rect 4035 2400 4037 2408
rect 4051 2400 4053 2408
rect 4056 2400 4058 2408
rect 4077 2400 4079 2408
rect 4093 2400 4095 2408
rect 4109 2400 4111 2408
rect 4114 2400 4116 2408
rect 4130 2400 4132 2408
rect 2286 2370 2288 2378
rect 2291 2370 2293 2378
rect 2307 2370 2309 2378
rect 2323 2370 2325 2378
rect 2328 2370 2330 2378
rect 2349 2370 2351 2378
rect 2365 2370 2367 2378
rect 2381 2370 2383 2378
rect 2386 2370 2388 2378
rect 2402 2370 2404 2378
rect 2418 2370 2420 2378
rect 2423 2370 2425 2378
rect 2439 2370 2441 2378
rect 2455 2370 2457 2378
rect 2460 2370 2462 2378
rect 2481 2370 2483 2378
rect 2497 2370 2499 2378
rect 2513 2370 2515 2378
rect 2518 2370 2520 2378
rect 2534 2370 2536 2378
rect 2550 2370 2552 2378
rect 2555 2370 2557 2378
rect 2571 2370 2573 2378
rect 2587 2370 2589 2378
rect 2592 2370 2594 2378
rect 2613 2370 2615 2378
rect 2629 2370 2631 2378
rect 2645 2370 2647 2378
rect 2650 2370 2652 2378
rect 2666 2370 2668 2378
rect 3231 2370 3233 2378
rect 3236 2370 3238 2378
rect 3252 2370 3254 2378
rect 3268 2370 3270 2378
rect 3273 2370 3275 2378
rect 3294 2370 3296 2378
rect 3310 2370 3312 2378
rect 3326 2370 3328 2378
rect 3331 2370 3333 2378
rect 3347 2370 3349 2378
rect 3363 2370 3365 2378
rect 3368 2370 3370 2378
rect 3384 2370 3386 2378
rect 3400 2370 3402 2378
rect 3405 2370 3407 2378
rect 3426 2370 3428 2378
rect 3442 2370 3444 2378
rect 3458 2370 3460 2378
rect 3463 2370 3465 2378
rect 3479 2370 3481 2378
rect 3495 2370 3497 2378
rect 3500 2370 3502 2378
rect 3516 2370 3518 2378
rect 3532 2370 3534 2378
rect 3537 2370 3539 2378
rect 3558 2370 3560 2378
rect 3574 2370 3576 2378
rect 3590 2370 3592 2378
rect 3595 2370 3597 2378
rect 3611 2370 3613 2378
rect 3069 2314 3071 2322
rect 3074 2314 3076 2322
rect 3090 2314 3092 2322
rect 3106 2314 3108 2322
rect 3111 2314 3113 2322
rect 3132 2314 3134 2322
rect 3148 2314 3150 2322
rect 3164 2314 3166 2322
rect 3169 2314 3171 2322
rect 3185 2314 3187 2322
rect 4014 2314 4016 2322
rect 4019 2314 4021 2322
rect 4035 2314 4037 2322
rect 4051 2314 4053 2322
rect 4056 2314 4058 2322
rect 4077 2314 4079 2322
rect 4093 2314 4095 2322
rect 4109 2314 4111 2322
rect 4114 2314 4116 2322
rect 4130 2314 4132 2322
rect 2286 2284 2288 2292
rect 2291 2284 2293 2292
rect 2307 2284 2309 2292
rect 2323 2284 2325 2292
rect 2328 2284 2330 2292
rect 2349 2284 2351 2292
rect 2365 2284 2367 2292
rect 2381 2284 2383 2292
rect 2386 2284 2388 2292
rect 2402 2284 2404 2292
rect 2418 2284 2420 2292
rect 2423 2284 2425 2292
rect 2439 2284 2441 2292
rect 2455 2284 2457 2292
rect 2460 2284 2462 2292
rect 2481 2284 2483 2292
rect 2497 2284 2499 2292
rect 2513 2284 2515 2292
rect 2518 2284 2520 2292
rect 2534 2284 2536 2292
rect 2550 2284 2552 2292
rect 2555 2284 2557 2292
rect 2571 2284 2573 2292
rect 2587 2284 2589 2292
rect 2592 2284 2594 2292
rect 2613 2284 2615 2292
rect 2629 2284 2631 2292
rect 2645 2284 2647 2292
rect 2650 2284 2652 2292
rect 2666 2284 2668 2292
rect 3231 2284 3233 2292
rect 3236 2284 3238 2292
rect 3252 2284 3254 2292
rect 3268 2284 3270 2292
rect 3273 2284 3275 2292
rect 3294 2284 3296 2292
rect 3310 2284 3312 2292
rect 3326 2284 3328 2292
rect 3331 2284 3333 2292
rect 3347 2284 3349 2292
rect 3363 2284 3365 2292
rect 3368 2284 3370 2292
rect 3384 2284 3386 2292
rect 3400 2284 3402 2292
rect 3405 2284 3407 2292
rect 3426 2284 3428 2292
rect 3442 2284 3444 2292
rect 3458 2284 3460 2292
rect 3463 2284 3465 2292
rect 3479 2284 3481 2292
rect 3495 2284 3497 2292
rect 3500 2284 3502 2292
rect 3516 2284 3518 2292
rect 3532 2284 3534 2292
rect 3537 2284 3539 2292
rect 3558 2284 3560 2292
rect 3574 2284 3576 2292
rect 3590 2284 3592 2292
rect 3595 2284 3597 2292
rect 3611 2284 3613 2292
rect 2286 2144 2288 2152
rect 2291 2144 2293 2152
rect 2307 2144 2309 2152
rect 2323 2144 2325 2152
rect 2328 2144 2330 2152
rect 2349 2144 2351 2152
rect 2365 2144 2367 2152
rect 2381 2144 2383 2152
rect 2386 2144 2388 2152
rect 2402 2144 2404 2152
rect 2418 2144 2420 2152
rect 2423 2144 2425 2152
rect 2439 2144 2441 2152
rect 2455 2144 2457 2152
rect 2460 2144 2462 2152
rect 2481 2144 2483 2152
rect 2497 2144 2499 2152
rect 2513 2144 2515 2152
rect 2518 2144 2520 2152
rect 2534 2144 2536 2152
rect 2550 2144 2552 2152
rect 2555 2144 2557 2152
rect 2571 2144 2573 2152
rect 2587 2144 2589 2152
rect 2592 2144 2594 2152
rect 2613 2144 2615 2152
rect 2629 2144 2631 2152
rect 2645 2144 2647 2152
rect 2650 2144 2652 2152
rect 2666 2144 2668 2152
rect 3231 2144 3233 2152
rect 3236 2144 3238 2152
rect 3252 2144 3254 2152
rect 3268 2144 3270 2152
rect 3273 2144 3275 2152
rect 3294 2144 3296 2152
rect 3310 2144 3312 2152
rect 3326 2144 3328 2152
rect 3331 2144 3333 2152
rect 3347 2144 3349 2152
rect 3363 2144 3365 2152
rect 3368 2144 3370 2152
rect 3384 2144 3386 2152
rect 3400 2144 3402 2152
rect 3405 2144 3407 2152
rect 3426 2144 3428 2152
rect 3442 2144 3444 2152
rect 3458 2144 3460 2152
rect 3463 2144 3465 2152
rect 3479 2144 3481 2152
rect 3495 2144 3497 2152
rect 3500 2144 3502 2152
rect 3516 2144 3518 2152
rect 3532 2144 3534 2152
rect 3537 2144 3539 2152
rect 3558 2144 3560 2152
rect 3574 2144 3576 2152
rect 3590 2144 3592 2152
rect 3595 2144 3597 2152
rect 3611 2144 3613 2152
<< ndiffusion >>
rect 2769 4006 2770 4010
rect 2772 4006 2775 4010
rect 2777 4006 2778 4010
rect 2790 4006 2791 4010
rect 2793 4006 2794 4010
rect 2806 4006 2807 4010
rect 2809 4006 2812 4010
rect 2814 4006 2815 4010
rect 2832 4006 2833 4010
rect 2835 4006 2836 4010
rect 2848 4006 2849 4010
rect 2851 4006 2852 4010
rect 2864 4006 2865 4010
rect 2867 4006 2870 4010
rect 2872 4006 2873 4010
rect 2885 4006 2886 4010
rect 2888 4006 2889 4010
rect 2901 4006 2902 4010
rect 2904 4006 2907 4010
rect 2909 4006 2910 4010
rect 2922 4006 2923 4010
rect 2925 4006 2926 4010
rect 2938 4006 2939 4010
rect 2941 4006 2944 4010
rect 2946 4006 2947 4010
rect 2964 4006 2965 4010
rect 2967 4006 2968 4010
rect 2980 4006 2981 4010
rect 2983 4006 2984 4010
rect 2996 4006 2997 4010
rect 2999 4006 3002 4010
rect 3004 4006 3005 4010
rect 3017 4006 3018 4010
rect 3020 4006 3021 4010
rect 3033 4006 3034 4010
rect 3036 4006 3039 4010
rect 3041 4006 3042 4010
rect 3054 4006 3055 4010
rect 3057 4006 3058 4010
rect 3070 4006 3071 4010
rect 3073 4006 3076 4010
rect 3078 4006 3079 4010
rect 3096 4006 3097 4010
rect 3099 4006 3100 4010
rect 3112 4006 3113 4010
rect 3115 4006 3116 4010
rect 3128 4006 3129 4010
rect 3131 4006 3134 4010
rect 3136 4006 3137 4010
rect 3149 4006 3150 4010
rect 3152 4006 3153 4010
rect 3165 4006 3166 4010
rect 3168 4006 3171 4010
rect 3173 4006 3174 4010
rect 3186 4006 3187 4010
rect 3189 4006 3190 4010
rect 3202 4006 3203 4010
rect 3205 4006 3208 4010
rect 3210 4006 3211 4010
rect 3228 4006 3229 4010
rect 3231 4006 3232 4010
rect 3244 4006 3245 4010
rect 3247 4006 3248 4010
rect 3260 4006 3261 4010
rect 3263 4006 3266 4010
rect 3268 4006 3269 4010
rect 3281 4006 3282 4010
rect 3284 4006 3285 4010
rect 3714 4006 3715 4010
rect 3717 4006 3720 4010
rect 3722 4006 3723 4010
rect 3735 4006 3736 4010
rect 3738 4006 3739 4010
rect 3751 4006 3752 4010
rect 3754 4006 3757 4010
rect 3759 4006 3760 4010
rect 3777 4006 3778 4010
rect 3780 4006 3781 4010
rect 3793 4006 3794 4010
rect 3796 4006 3797 4010
rect 3809 4006 3810 4010
rect 3812 4006 3815 4010
rect 3817 4006 3818 4010
rect 3830 4006 3831 4010
rect 3833 4006 3834 4010
rect 3846 4006 3847 4010
rect 3849 4006 3852 4010
rect 3854 4006 3855 4010
rect 3867 4006 3868 4010
rect 3870 4006 3871 4010
rect 3883 4006 3884 4010
rect 3886 4006 3889 4010
rect 3891 4006 3892 4010
rect 3909 4006 3910 4010
rect 3912 4006 3913 4010
rect 3925 4006 3926 4010
rect 3928 4006 3929 4010
rect 3941 4006 3942 4010
rect 3944 4006 3947 4010
rect 3949 4006 3950 4010
rect 3962 4006 3963 4010
rect 3965 4006 3966 4010
rect 3978 4006 3979 4010
rect 3981 4006 3984 4010
rect 3986 4006 3987 4010
rect 3999 4006 4000 4010
rect 4002 4006 4003 4010
rect 4015 4006 4016 4010
rect 4018 4006 4021 4010
rect 4023 4006 4024 4010
rect 4041 4006 4042 4010
rect 4044 4006 4045 4010
rect 4057 4006 4058 4010
rect 4060 4006 4061 4010
rect 4073 4006 4074 4010
rect 4076 4006 4079 4010
rect 4081 4006 4082 4010
rect 4094 4006 4095 4010
rect 4097 4006 4098 4010
rect 4110 4006 4111 4010
rect 4113 4006 4116 4010
rect 4118 4006 4119 4010
rect 4131 4006 4132 4010
rect 4134 4006 4135 4010
rect 4147 4006 4148 4010
rect 4150 4006 4153 4010
rect 4155 4006 4156 4010
rect 4173 4006 4174 4010
rect 4176 4006 4177 4010
rect 4189 4006 4190 4010
rect 4192 4006 4193 4010
rect 4205 4006 4206 4010
rect 4208 4006 4211 4010
rect 4213 4006 4214 4010
rect 4226 4006 4227 4010
rect 4229 4006 4230 4010
rect 2417 3973 2418 3977
rect 2420 3973 2423 3977
rect 2425 3973 2426 3977
rect 2438 3973 2439 3977
rect 2441 3973 2442 3977
rect 2454 3973 2455 3977
rect 2457 3973 2460 3977
rect 2462 3973 2463 3977
rect 2480 3973 2481 3977
rect 2483 3973 2484 3977
rect 2496 3973 2497 3977
rect 2499 3973 2500 3977
rect 2512 3973 2513 3977
rect 2515 3973 2518 3977
rect 2520 3973 2521 3977
rect 2533 3973 2534 3977
rect 2536 3973 2537 3977
rect 3362 3973 3363 3977
rect 3365 3973 3368 3977
rect 3370 3973 3371 3977
rect 3383 3973 3384 3977
rect 3386 3973 3387 3977
rect 3399 3973 3400 3977
rect 3402 3973 3405 3977
rect 3407 3973 3408 3977
rect 3425 3973 3426 3977
rect 3428 3973 3429 3977
rect 3441 3973 3442 3977
rect 3444 3973 3445 3977
rect 3457 3973 3458 3977
rect 3460 3973 3463 3977
rect 3465 3973 3466 3977
rect 3478 3973 3479 3977
rect 3481 3973 3482 3977
rect 2541 3936 2542 3940
rect 2544 3936 2545 3940
rect 2948 3940 2949 3944
rect 2951 3940 2952 3944
rect 2972 3936 2975 3940
rect 2977 3936 2980 3940
rect 2982 3936 2983 3940
rect 3029 3940 3030 3944
rect 3032 3940 3033 3944
rect 3053 3936 3056 3940
rect 3058 3936 3061 3940
rect 3063 3936 3064 3940
rect 3002 3932 3003 3936
rect 3005 3932 3006 3936
rect 2424 3927 2425 3931
rect 2427 3927 2428 3931
rect 2774 3927 2775 3931
rect 2777 3927 2778 3931
rect 2790 3927 2791 3931
rect 2793 3927 2794 3931
rect 2806 3927 2807 3931
rect 2809 3927 2810 3931
rect 2825 3927 2830 3931
rect 2832 3927 2835 3931
rect 2837 3927 2838 3931
rect 2859 3927 2861 3931
rect 2863 3927 2864 3931
rect 2881 3927 2882 3931
rect 2884 3927 2885 3931
rect 2897 3927 2902 3931
rect 2904 3927 2907 3931
rect 2909 3927 2910 3931
rect 2924 3927 2925 3931
rect 2927 3927 2928 3931
rect 3083 3932 3084 3936
rect 3086 3932 3087 3936
rect 3486 3936 3487 3940
rect 3489 3936 3490 3940
rect 3893 3940 3894 3944
rect 3896 3940 3897 3944
rect 3917 3936 3920 3940
rect 3922 3936 3925 3940
rect 3927 3936 3928 3940
rect 3974 3940 3975 3944
rect 3977 3940 3978 3944
rect 3998 3936 4001 3940
rect 4003 3936 4006 3940
rect 4008 3936 4009 3940
rect 3947 3932 3948 3936
rect 3950 3932 3951 3936
rect 3369 3927 3370 3931
rect 3372 3927 3373 3931
rect 3719 3927 3720 3931
rect 3722 3927 3723 3931
rect 3735 3927 3736 3931
rect 3738 3927 3739 3931
rect 3751 3927 3752 3931
rect 3754 3927 3755 3931
rect 3770 3927 3775 3931
rect 3777 3927 3780 3931
rect 3782 3927 3783 3931
rect 3804 3927 3806 3931
rect 3808 3927 3809 3931
rect 3826 3927 3827 3931
rect 3829 3927 3830 3931
rect 3842 3927 3847 3931
rect 3849 3927 3852 3931
rect 3854 3927 3855 3931
rect 3869 3927 3870 3931
rect 3872 3927 3873 3931
rect 4028 3932 4029 3936
rect 4031 3932 4032 3936
rect 2774 3881 2775 3885
rect 2777 3881 2778 3885
rect 2790 3881 2791 3885
rect 2793 3881 2794 3885
rect 2806 3881 2807 3885
rect 2809 3881 2810 3885
rect 2825 3881 2830 3885
rect 2832 3881 2835 3885
rect 2837 3881 2838 3885
rect 2859 3881 2861 3885
rect 2863 3881 2864 3885
rect 2881 3881 2882 3885
rect 2884 3881 2885 3885
rect 2897 3881 2902 3885
rect 2904 3881 2907 3885
rect 2909 3881 2910 3885
rect 2924 3881 2925 3885
rect 2927 3881 2928 3885
rect 2408 3871 2409 3875
rect 2411 3871 2412 3875
rect 2424 3871 2425 3875
rect 2427 3871 2430 3875
rect 2432 3871 2433 3875
rect 2445 3871 2446 3875
rect 2448 3871 2449 3875
rect 2461 3871 2462 3875
rect 2464 3871 2465 3875
rect 2482 3871 2483 3875
rect 2485 3871 2488 3875
rect 2490 3871 2491 3875
rect 2503 3871 2504 3875
rect 2506 3871 2507 3875
rect 2519 3871 2520 3875
rect 2522 3871 2525 3875
rect 2527 3871 2528 3875
rect 2972 3880 2975 3884
rect 2977 3880 2980 3884
rect 2982 3880 2983 3884
rect 3053 3880 3056 3884
rect 3058 3880 3061 3884
rect 3063 3880 3064 3884
rect 3719 3881 3720 3885
rect 3722 3881 3723 3885
rect 3735 3881 3736 3885
rect 3738 3881 3739 3885
rect 3751 3881 3752 3885
rect 3754 3881 3755 3885
rect 3770 3881 3775 3885
rect 3777 3881 3780 3885
rect 3782 3881 3783 3885
rect 3804 3881 3806 3885
rect 3808 3881 3809 3885
rect 3826 3881 3827 3885
rect 3829 3881 3830 3885
rect 3842 3881 3847 3885
rect 3849 3881 3852 3885
rect 3854 3881 3855 3885
rect 3869 3881 3870 3885
rect 3872 3881 3873 3885
rect 3353 3871 3354 3875
rect 3356 3871 3357 3875
rect 3369 3871 3370 3875
rect 3372 3871 3375 3875
rect 3377 3871 3378 3875
rect 3390 3871 3391 3875
rect 3393 3871 3394 3875
rect 3406 3871 3407 3875
rect 3409 3871 3410 3875
rect 3427 3871 3428 3875
rect 3430 3871 3433 3875
rect 3435 3871 3436 3875
rect 3448 3871 3449 3875
rect 3451 3871 3452 3875
rect 3464 3871 3465 3875
rect 3467 3871 3470 3875
rect 3472 3871 3473 3875
rect 3917 3880 3920 3884
rect 3922 3880 3925 3884
rect 3927 3880 3928 3884
rect 3998 3880 4001 3884
rect 4003 3880 4006 3884
rect 4008 3880 4009 3884
rect 2972 3804 2975 3808
rect 2977 3804 2980 3808
rect 2982 3804 2983 3808
rect 3053 3808 3054 3812
rect 3056 3808 3057 3812
rect 3077 3804 3080 3808
rect 3082 3804 3085 3808
rect 3087 3804 3088 3808
rect 3002 3800 3003 3804
rect 3005 3800 3006 3804
rect 2774 3795 2775 3799
rect 2777 3795 2778 3799
rect 2790 3795 2791 3799
rect 2793 3795 2794 3799
rect 2806 3795 2807 3799
rect 2809 3795 2810 3799
rect 2825 3795 2830 3799
rect 2832 3795 2835 3799
rect 2837 3795 2838 3799
rect 2859 3795 2861 3799
rect 2863 3795 2864 3799
rect 2881 3795 2882 3799
rect 2884 3795 2885 3799
rect 2897 3795 2902 3799
rect 2904 3795 2907 3799
rect 2909 3795 2910 3799
rect 2924 3795 2925 3799
rect 2927 3795 2928 3799
rect 3107 3800 3108 3804
rect 3110 3800 3111 3804
rect 3284 3779 3285 3783
rect 3287 3779 3288 3783
rect 3308 3775 3311 3779
rect 3313 3775 3316 3779
rect 3318 3775 3319 3779
rect 3338 3771 3339 3775
rect 3341 3771 3342 3775
rect 3917 3804 3920 3808
rect 3922 3804 3925 3808
rect 3927 3804 3928 3808
rect 3998 3808 3999 3812
rect 4001 3808 4002 3812
rect 4022 3804 4025 3808
rect 4027 3804 4030 3808
rect 4032 3804 4033 3808
rect 3947 3800 3948 3804
rect 3950 3800 3951 3804
rect 3719 3795 3720 3799
rect 3722 3795 3723 3799
rect 3735 3795 3736 3799
rect 3738 3795 3739 3799
rect 3751 3795 3752 3799
rect 3754 3795 3755 3799
rect 3770 3795 3775 3799
rect 3777 3795 3780 3799
rect 3782 3795 3783 3799
rect 3804 3795 3806 3799
rect 3808 3795 3809 3799
rect 3826 3795 3827 3799
rect 3829 3795 3830 3799
rect 3842 3795 3847 3799
rect 3849 3795 3852 3799
rect 3854 3795 3855 3799
rect 3869 3795 3870 3799
rect 3872 3795 3873 3799
rect 4052 3800 4053 3804
rect 4055 3800 4056 3804
rect 2774 3749 2775 3753
rect 2777 3749 2778 3753
rect 2790 3749 2791 3753
rect 2793 3749 2794 3753
rect 2806 3749 2807 3753
rect 2809 3749 2810 3753
rect 2825 3749 2830 3753
rect 2832 3749 2835 3753
rect 2837 3749 2838 3753
rect 2859 3749 2861 3753
rect 2863 3749 2864 3753
rect 2881 3749 2882 3753
rect 2884 3749 2885 3753
rect 2897 3749 2902 3753
rect 2904 3749 2907 3753
rect 2909 3749 2910 3753
rect 2924 3749 2925 3753
rect 2927 3749 2928 3753
rect 2972 3749 2975 3753
rect 2977 3749 2980 3753
rect 2982 3749 2983 3753
rect 3077 3749 3080 3753
rect 3082 3749 3085 3753
rect 3087 3749 3088 3753
rect 3470 3740 3471 3752
rect 3473 3740 3474 3752
rect 3523 3740 3524 3752
rect 3526 3740 3527 3752
rect 3719 3749 3720 3753
rect 3722 3749 3723 3753
rect 3735 3749 3736 3753
rect 3738 3749 3739 3753
rect 3751 3749 3752 3753
rect 3754 3749 3755 3753
rect 3770 3749 3775 3753
rect 3777 3749 3780 3753
rect 3782 3749 3783 3753
rect 3804 3749 3806 3753
rect 3808 3749 3809 3753
rect 3826 3749 3827 3753
rect 3829 3749 3830 3753
rect 3842 3749 3847 3753
rect 3849 3749 3852 3753
rect 3854 3749 3855 3753
rect 3869 3749 3870 3753
rect 3872 3749 3873 3753
rect 3917 3749 3920 3753
rect 3922 3749 3925 3753
rect 3927 3749 3928 3753
rect 4022 3749 4025 3753
rect 4027 3749 4030 3753
rect 4032 3749 4033 3753
rect 3308 3715 3311 3719
rect 3313 3715 3316 3719
rect 3318 3715 3319 3719
rect 2972 3672 2975 3676
rect 2977 3672 2980 3676
rect 2982 3672 2983 3676
rect 3029 3676 3030 3680
rect 3032 3676 3033 3680
rect 3053 3672 3056 3676
rect 3058 3672 3061 3676
rect 3063 3672 3064 3676
rect 3119 3676 3120 3680
rect 3122 3676 3123 3680
rect 3143 3672 3146 3676
rect 3148 3672 3151 3676
rect 3153 3672 3154 3676
rect 3002 3668 3003 3672
rect 3005 3668 3006 3672
rect 2774 3663 2775 3667
rect 2777 3663 2778 3667
rect 2790 3663 2791 3667
rect 2793 3663 2794 3667
rect 2806 3663 2807 3667
rect 2809 3663 2810 3667
rect 2825 3663 2830 3667
rect 2832 3663 2835 3667
rect 2837 3663 2838 3667
rect 2859 3663 2861 3667
rect 2863 3663 2864 3667
rect 2881 3663 2882 3667
rect 2884 3663 2885 3667
rect 2897 3663 2902 3667
rect 2904 3663 2907 3667
rect 2909 3663 2910 3667
rect 2924 3663 2925 3667
rect 2927 3663 2928 3667
rect 3083 3668 3084 3672
rect 3086 3668 3087 3672
rect 3173 3668 3174 3672
rect 3176 3668 3177 3672
rect 3262 3649 3263 3653
rect 3265 3649 3266 3653
rect 3284 3649 3285 3653
rect 3287 3649 3288 3653
rect 3308 3645 3311 3649
rect 3313 3645 3316 3649
rect 3318 3645 3319 3649
rect 3338 3641 3339 3645
rect 3341 3641 3342 3645
rect 3917 3672 3920 3676
rect 3922 3672 3925 3676
rect 3927 3672 3928 3676
rect 3974 3676 3975 3680
rect 3977 3676 3978 3680
rect 3998 3672 4001 3676
rect 4003 3672 4006 3676
rect 4008 3672 4009 3676
rect 4064 3676 4065 3680
rect 4067 3676 4068 3680
rect 4088 3672 4091 3676
rect 4093 3672 4096 3676
rect 4098 3672 4099 3676
rect 3947 3668 3948 3672
rect 3950 3668 3951 3672
rect 3719 3663 3720 3667
rect 3722 3663 3723 3667
rect 3735 3663 3736 3667
rect 3738 3663 3739 3667
rect 3751 3663 3752 3667
rect 3754 3663 3755 3667
rect 3770 3663 3775 3667
rect 3777 3663 3780 3667
rect 3782 3663 3783 3667
rect 3804 3663 3806 3667
rect 3808 3663 3809 3667
rect 3826 3663 3827 3667
rect 3829 3663 3830 3667
rect 3842 3663 3847 3667
rect 3849 3663 3852 3667
rect 3854 3663 3855 3667
rect 3869 3663 3870 3667
rect 3872 3663 3873 3667
rect 4028 3668 4029 3672
rect 4031 3668 4032 3672
rect 4118 3668 4119 3672
rect 4121 3668 4122 3672
rect 2774 3617 2775 3621
rect 2777 3617 2778 3621
rect 2790 3617 2791 3621
rect 2793 3617 2794 3621
rect 2806 3617 2807 3621
rect 2809 3617 2810 3621
rect 2825 3617 2830 3621
rect 2832 3617 2835 3621
rect 2837 3617 2838 3621
rect 2859 3617 2861 3621
rect 2863 3617 2864 3621
rect 2881 3617 2882 3621
rect 2884 3617 2885 3621
rect 2897 3617 2902 3621
rect 2904 3617 2907 3621
rect 2909 3617 2910 3621
rect 2924 3617 2925 3621
rect 2927 3617 2928 3621
rect 2972 3614 2975 3618
rect 2977 3614 2980 3618
rect 2982 3614 2983 3618
rect 3053 3614 3056 3618
rect 3058 3614 3061 3618
rect 3063 3614 3064 3618
rect 3143 3614 3146 3618
rect 3148 3614 3151 3618
rect 3153 3614 3154 3618
rect 3376 3610 3377 3622
rect 3379 3610 3380 3622
rect 3429 3610 3430 3622
rect 3432 3610 3433 3622
rect 3719 3617 3720 3621
rect 3722 3617 3723 3621
rect 3735 3617 3736 3621
rect 3738 3617 3739 3621
rect 3751 3617 3752 3621
rect 3754 3617 3755 3621
rect 3770 3617 3775 3621
rect 3777 3617 3780 3621
rect 3782 3617 3783 3621
rect 3804 3617 3806 3621
rect 3808 3617 3809 3621
rect 3826 3617 3827 3621
rect 3829 3617 3830 3621
rect 3842 3617 3847 3621
rect 3849 3617 3852 3621
rect 3854 3617 3855 3621
rect 3869 3617 3870 3621
rect 3872 3617 3873 3621
rect 3917 3614 3920 3618
rect 3922 3614 3925 3618
rect 3927 3614 3928 3618
rect 3998 3614 4001 3618
rect 4003 3614 4006 3618
rect 4008 3614 4009 3618
rect 4088 3614 4091 3618
rect 4093 3614 4096 3618
rect 4098 3614 4099 3618
rect 3308 3585 3311 3589
rect 3313 3585 3316 3589
rect 3318 3585 3319 3589
rect 2972 3540 2975 3544
rect 2977 3540 2980 3544
rect 2982 3540 2983 3544
rect 3002 3536 3003 3540
rect 3005 3536 3006 3540
rect 2774 3531 2775 3535
rect 2777 3531 2778 3535
rect 2790 3531 2791 3535
rect 2793 3531 2794 3535
rect 2806 3531 2807 3535
rect 2809 3531 2810 3535
rect 2825 3531 2830 3535
rect 2832 3531 2835 3535
rect 2837 3531 2838 3535
rect 2859 3531 2861 3535
rect 2863 3531 2864 3535
rect 2881 3531 2882 3535
rect 2884 3531 2885 3535
rect 2897 3531 2902 3535
rect 2904 3531 2907 3535
rect 2909 3531 2910 3535
rect 2924 3531 2925 3535
rect 2927 3531 2928 3535
rect 3917 3540 3920 3544
rect 3922 3540 3925 3544
rect 3927 3540 3928 3544
rect 3947 3536 3948 3540
rect 3950 3536 3951 3540
rect 3719 3531 3720 3535
rect 3722 3531 3723 3535
rect 3735 3531 3736 3535
rect 3738 3531 3739 3535
rect 3751 3531 3752 3535
rect 3754 3531 3755 3535
rect 3770 3531 3775 3535
rect 3777 3531 3780 3535
rect 3782 3531 3783 3535
rect 3804 3531 3806 3535
rect 3808 3531 3809 3535
rect 3826 3531 3827 3535
rect 3829 3531 3830 3535
rect 3842 3531 3847 3535
rect 3849 3531 3852 3535
rect 3854 3531 3855 3535
rect 3869 3531 3870 3535
rect 3872 3531 3873 3535
rect 2774 3485 2775 3489
rect 2777 3485 2778 3489
rect 2790 3485 2791 3489
rect 2793 3485 2794 3489
rect 2806 3485 2807 3489
rect 2809 3485 2810 3489
rect 2825 3485 2830 3489
rect 2832 3485 2835 3489
rect 2837 3485 2838 3489
rect 2859 3485 2861 3489
rect 2863 3485 2864 3489
rect 2881 3485 2882 3489
rect 2884 3485 2885 3489
rect 2897 3485 2902 3489
rect 2904 3485 2907 3489
rect 2909 3485 2910 3489
rect 2924 3485 2925 3489
rect 2927 3485 2928 3489
rect 3008 3485 3009 3489
rect 3011 3485 3012 3489
rect 3016 3485 3022 3489
rect 3026 3485 3027 3489
rect 3029 3485 3030 3489
rect 3051 3485 3052 3489
rect 3054 3485 3055 3489
rect 3067 3485 3068 3489
rect 3070 3485 3071 3489
rect 3086 3485 3091 3489
rect 3093 3485 3096 3489
rect 3098 3485 3099 3489
rect 3120 3485 3122 3489
rect 3124 3485 3125 3489
rect 3142 3485 3143 3489
rect 3145 3485 3146 3489
rect 3158 3485 3163 3489
rect 3165 3485 3168 3489
rect 3170 3485 3171 3489
rect 3185 3485 3186 3489
rect 3188 3485 3189 3489
rect 2285 3471 2286 3475
rect 2288 3471 2291 3475
rect 2293 3471 2294 3475
rect 2306 3471 2307 3475
rect 2309 3471 2310 3475
rect 2322 3471 2323 3475
rect 2325 3471 2328 3475
rect 2330 3471 2331 3475
rect 2348 3471 2349 3475
rect 2351 3471 2352 3475
rect 2364 3471 2365 3475
rect 2367 3471 2368 3475
rect 2380 3471 2381 3475
rect 2383 3471 2386 3475
rect 2388 3471 2389 3475
rect 2401 3471 2402 3475
rect 2404 3471 2405 3475
rect 2417 3471 2418 3475
rect 2420 3471 2423 3475
rect 2425 3471 2426 3475
rect 2438 3471 2439 3475
rect 2441 3471 2442 3475
rect 2454 3471 2455 3475
rect 2457 3471 2460 3475
rect 2462 3471 2463 3475
rect 2480 3471 2481 3475
rect 2483 3471 2484 3475
rect 2496 3471 2497 3475
rect 2499 3471 2500 3475
rect 2512 3471 2513 3475
rect 2515 3471 2518 3475
rect 2520 3471 2521 3475
rect 2533 3471 2534 3475
rect 2536 3471 2537 3475
rect 2549 3471 2550 3475
rect 2552 3471 2555 3475
rect 2557 3471 2558 3475
rect 2570 3471 2571 3475
rect 2573 3471 2574 3475
rect 2586 3471 2587 3475
rect 2589 3471 2592 3475
rect 2594 3471 2595 3475
rect 2612 3471 2613 3475
rect 2615 3471 2616 3475
rect 2628 3471 2629 3475
rect 2631 3471 2632 3475
rect 2644 3471 2645 3475
rect 2647 3471 2650 3475
rect 2652 3471 2653 3475
rect 2665 3471 2666 3475
rect 2668 3471 2669 3475
rect 2972 3478 2975 3482
rect 2977 3478 2980 3482
rect 2982 3478 2983 3482
rect 3719 3485 3720 3489
rect 3722 3485 3723 3489
rect 3735 3485 3736 3489
rect 3738 3485 3739 3489
rect 3751 3485 3752 3489
rect 3754 3485 3755 3489
rect 3770 3485 3775 3489
rect 3777 3485 3780 3489
rect 3782 3485 3783 3489
rect 3804 3485 3806 3489
rect 3808 3485 3809 3489
rect 3826 3485 3827 3489
rect 3829 3485 3830 3489
rect 3842 3485 3847 3489
rect 3849 3485 3852 3489
rect 3854 3485 3855 3489
rect 3869 3485 3870 3489
rect 3872 3485 3873 3489
rect 3953 3485 3954 3489
rect 3956 3485 3957 3489
rect 3961 3485 3967 3489
rect 3971 3485 3972 3489
rect 3974 3485 3975 3489
rect 3996 3485 3997 3489
rect 3999 3485 4000 3489
rect 4012 3485 4013 3489
rect 4015 3485 4016 3489
rect 4031 3485 4036 3489
rect 4038 3485 4041 3489
rect 4043 3485 4044 3489
rect 4065 3485 4067 3489
rect 4069 3485 4070 3489
rect 4087 3485 4088 3489
rect 4090 3485 4091 3489
rect 4103 3485 4108 3489
rect 4110 3485 4113 3489
rect 4115 3485 4116 3489
rect 4130 3485 4131 3489
rect 4133 3485 4134 3489
rect 3230 3471 3231 3475
rect 3233 3471 3236 3475
rect 3238 3471 3239 3475
rect 3251 3471 3252 3475
rect 3254 3471 3255 3475
rect 3267 3471 3268 3475
rect 3270 3471 3273 3475
rect 3275 3471 3276 3475
rect 3293 3471 3294 3475
rect 3296 3471 3297 3475
rect 3309 3471 3310 3475
rect 3312 3471 3313 3475
rect 3325 3471 3326 3475
rect 3328 3471 3331 3475
rect 3333 3471 3334 3475
rect 3346 3471 3347 3475
rect 3349 3471 3350 3475
rect 3362 3471 3363 3475
rect 3365 3471 3368 3475
rect 3370 3471 3371 3475
rect 3383 3471 3384 3475
rect 3386 3471 3387 3475
rect 3399 3471 3400 3475
rect 3402 3471 3405 3475
rect 3407 3471 3408 3475
rect 3425 3471 3426 3475
rect 3428 3471 3429 3475
rect 3441 3471 3442 3475
rect 3444 3471 3445 3475
rect 3457 3471 3458 3475
rect 3460 3471 3463 3475
rect 3465 3471 3466 3475
rect 3478 3471 3479 3475
rect 3481 3471 3482 3475
rect 3494 3471 3495 3475
rect 3497 3471 3500 3475
rect 3502 3471 3503 3475
rect 3515 3471 3516 3475
rect 3518 3471 3519 3475
rect 3531 3471 3532 3475
rect 3534 3471 3537 3475
rect 3539 3471 3540 3475
rect 3557 3471 3558 3475
rect 3560 3471 3561 3475
rect 3573 3471 3574 3475
rect 3576 3471 3577 3475
rect 3589 3471 3590 3475
rect 3592 3471 3595 3475
rect 3597 3471 3598 3475
rect 3610 3471 3611 3475
rect 3613 3471 3614 3475
rect 3917 3478 3920 3482
rect 3922 3478 3925 3482
rect 3927 3478 3928 3482
rect 2400 3427 2401 3431
rect 2403 3427 2404 3431
rect 2424 3427 2425 3431
rect 2427 3427 2428 3431
rect 3198 3431 3202 3432
rect 3198 3428 3202 3429
rect 3345 3427 3346 3431
rect 3348 3427 3349 3431
rect 3369 3427 3370 3431
rect 3372 3427 3373 3431
rect 4143 3431 4147 3432
rect 4143 3428 4147 3429
rect 2420 3414 2421 3418
rect 2423 3414 2424 3418
rect 3365 3414 3366 3418
rect 3368 3414 3369 3418
rect 2412 3402 2416 3403
rect 2412 3399 2416 3400
rect 3357 3402 3361 3403
rect 3357 3399 3361 3400
rect 2400 3391 2401 3395
rect 2403 3391 2404 3395
rect 2424 3391 2425 3395
rect 2427 3391 2428 3395
rect 3345 3391 3346 3395
rect 3348 3391 3349 3395
rect 3369 3391 3370 3395
rect 3372 3391 3373 3395
rect 3068 3359 3069 3363
rect 3071 3359 3074 3363
rect 3076 3359 3077 3363
rect 3089 3359 3090 3363
rect 3092 3359 3093 3363
rect 3105 3359 3106 3363
rect 3108 3359 3111 3363
rect 3113 3359 3114 3363
rect 3131 3359 3132 3363
rect 3134 3359 3135 3363
rect 3147 3359 3148 3363
rect 3150 3359 3151 3363
rect 3163 3359 3164 3363
rect 3166 3359 3169 3363
rect 3171 3359 3172 3363
rect 3184 3359 3185 3363
rect 3187 3359 3188 3363
rect 4013 3359 4014 3363
rect 4016 3359 4019 3363
rect 4021 3359 4022 3363
rect 4034 3359 4035 3363
rect 4037 3359 4038 3363
rect 4050 3359 4051 3363
rect 4053 3359 4056 3363
rect 4058 3359 4059 3363
rect 4076 3359 4077 3363
rect 4079 3359 4080 3363
rect 4092 3359 4093 3363
rect 4095 3359 4096 3363
rect 4108 3359 4109 3363
rect 4111 3359 4114 3363
rect 4116 3359 4117 3363
rect 4129 3359 4130 3363
rect 4132 3359 4133 3363
rect 2285 3329 2286 3333
rect 2288 3329 2291 3333
rect 2293 3329 2294 3333
rect 2306 3329 2307 3333
rect 2309 3329 2310 3333
rect 2322 3329 2323 3333
rect 2325 3329 2328 3333
rect 2330 3329 2331 3333
rect 2348 3329 2349 3333
rect 2351 3329 2352 3333
rect 2364 3329 2365 3333
rect 2367 3329 2368 3333
rect 2380 3329 2381 3333
rect 2383 3329 2386 3333
rect 2388 3329 2389 3333
rect 2401 3329 2402 3333
rect 2404 3329 2405 3333
rect 2417 3329 2418 3333
rect 2420 3329 2423 3333
rect 2425 3329 2426 3333
rect 2438 3329 2439 3333
rect 2441 3329 2442 3333
rect 2454 3329 2455 3333
rect 2457 3329 2460 3333
rect 2462 3329 2463 3333
rect 2480 3329 2481 3333
rect 2483 3329 2484 3333
rect 2496 3329 2497 3333
rect 2499 3329 2500 3333
rect 2512 3329 2513 3333
rect 2515 3329 2518 3333
rect 2520 3329 2521 3333
rect 2533 3329 2534 3333
rect 2536 3329 2537 3333
rect 2549 3329 2550 3333
rect 2552 3329 2555 3333
rect 2557 3329 2558 3333
rect 2570 3329 2571 3333
rect 2573 3329 2574 3333
rect 2586 3329 2587 3333
rect 2589 3329 2592 3333
rect 2594 3329 2595 3333
rect 2612 3329 2613 3333
rect 2615 3329 2616 3333
rect 2628 3329 2629 3333
rect 2631 3329 2632 3333
rect 2644 3329 2645 3333
rect 2647 3329 2650 3333
rect 2652 3329 2653 3333
rect 2665 3329 2666 3333
rect 2668 3329 2669 3333
rect 3230 3329 3231 3333
rect 3233 3329 3236 3333
rect 3238 3329 3239 3333
rect 3251 3329 3252 3333
rect 3254 3329 3255 3333
rect 3267 3329 3268 3333
rect 3270 3329 3273 3333
rect 3275 3329 3276 3333
rect 3293 3329 3294 3333
rect 3296 3329 3297 3333
rect 3309 3329 3310 3333
rect 3312 3329 3313 3333
rect 3325 3329 3326 3333
rect 3328 3329 3331 3333
rect 3333 3329 3334 3333
rect 3346 3329 3347 3333
rect 3349 3329 3350 3333
rect 3362 3329 3363 3333
rect 3365 3329 3368 3333
rect 3370 3329 3371 3333
rect 3383 3329 3384 3333
rect 3386 3329 3387 3333
rect 3399 3329 3400 3333
rect 3402 3329 3405 3333
rect 3407 3329 3408 3333
rect 3425 3329 3426 3333
rect 3428 3329 3429 3333
rect 3441 3329 3442 3333
rect 3444 3329 3445 3333
rect 3457 3329 3458 3333
rect 3460 3329 3463 3333
rect 3465 3329 3466 3333
rect 3478 3329 3479 3333
rect 3481 3329 3482 3333
rect 3494 3329 3495 3333
rect 3497 3329 3500 3333
rect 3502 3329 3503 3333
rect 3515 3329 3516 3333
rect 3518 3329 3519 3333
rect 3531 3329 3532 3333
rect 3534 3329 3537 3333
rect 3539 3329 3540 3333
rect 3557 3329 3558 3333
rect 3560 3329 3561 3333
rect 3573 3329 3574 3333
rect 3576 3329 3577 3333
rect 3589 3329 3590 3333
rect 3592 3329 3595 3333
rect 3597 3329 3598 3333
rect 3610 3329 3611 3333
rect 3613 3329 3614 3333
rect 3210 3285 3214 3286
rect 3210 3282 3214 3283
rect 4155 3285 4159 3286
rect 4155 3282 4159 3283
rect 3068 3273 3069 3277
rect 3071 3273 3074 3277
rect 3076 3273 3077 3277
rect 3089 3273 3090 3277
rect 3092 3273 3093 3277
rect 3105 3273 3106 3277
rect 3108 3273 3111 3277
rect 3113 3273 3114 3277
rect 3131 3273 3132 3277
rect 3134 3273 3135 3277
rect 3147 3273 3148 3277
rect 3150 3273 3151 3277
rect 3163 3273 3164 3277
rect 3166 3273 3169 3277
rect 3171 3273 3172 3277
rect 3184 3273 3185 3277
rect 3187 3273 3188 3277
rect 4013 3273 4014 3277
rect 4016 3273 4019 3277
rect 4021 3273 4022 3277
rect 4034 3273 4035 3277
rect 4037 3273 4038 3277
rect 4050 3273 4051 3277
rect 4053 3273 4056 3277
rect 4058 3273 4059 3277
rect 4076 3273 4077 3277
rect 4079 3273 4080 3277
rect 4092 3273 4093 3277
rect 4095 3273 4096 3277
rect 4108 3273 4109 3277
rect 4111 3273 4114 3277
rect 4116 3273 4117 3277
rect 4129 3273 4130 3277
rect 4132 3273 4133 3277
rect 2285 3243 2286 3247
rect 2288 3243 2291 3247
rect 2293 3243 2294 3247
rect 2306 3243 2307 3247
rect 2309 3243 2310 3247
rect 2322 3243 2323 3247
rect 2325 3243 2328 3247
rect 2330 3243 2331 3247
rect 2348 3243 2349 3247
rect 2351 3243 2352 3247
rect 2364 3243 2365 3247
rect 2367 3243 2368 3247
rect 2380 3243 2381 3247
rect 2383 3243 2386 3247
rect 2388 3243 2389 3247
rect 2401 3243 2402 3247
rect 2404 3243 2405 3247
rect 2417 3243 2418 3247
rect 2420 3243 2423 3247
rect 2425 3243 2426 3247
rect 2438 3243 2439 3247
rect 2441 3243 2442 3247
rect 2454 3243 2455 3247
rect 2457 3243 2460 3247
rect 2462 3243 2463 3247
rect 2480 3243 2481 3247
rect 2483 3243 2484 3247
rect 2496 3243 2497 3247
rect 2499 3243 2500 3247
rect 2512 3243 2513 3247
rect 2515 3243 2518 3247
rect 2520 3243 2521 3247
rect 2533 3243 2534 3247
rect 2536 3243 2537 3247
rect 2549 3243 2550 3247
rect 2552 3243 2555 3247
rect 2557 3243 2558 3247
rect 2570 3243 2571 3247
rect 2573 3243 2574 3247
rect 2586 3243 2587 3247
rect 2589 3243 2592 3247
rect 2594 3243 2595 3247
rect 2612 3243 2613 3247
rect 2615 3243 2616 3247
rect 2628 3243 2629 3247
rect 2631 3243 2632 3247
rect 2644 3243 2645 3247
rect 2647 3243 2650 3247
rect 2652 3243 2653 3247
rect 2665 3243 2666 3247
rect 2668 3243 2669 3247
rect 3230 3243 3231 3247
rect 3233 3243 3236 3247
rect 3238 3243 3239 3247
rect 3251 3243 3252 3247
rect 3254 3243 3255 3247
rect 3267 3243 3268 3247
rect 3270 3243 3273 3247
rect 3275 3243 3276 3247
rect 3293 3243 3294 3247
rect 3296 3243 3297 3247
rect 3309 3243 3310 3247
rect 3312 3243 3313 3247
rect 3325 3243 3326 3247
rect 3328 3243 3331 3247
rect 3333 3243 3334 3247
rect 3346 3243 3347 3247
rect 3349 3243 3350 3247
rect 3362 3243 3363 3247
rect 3365 3243 3368 3247
rect 3370 3243 3371 3247
rect 3383 3243 3384 3247
rect 3386 3243 3387 3247
rect 3399 3243 3400 3247
rect 3402 3243 3405 3247
rect 3407 3243 3408 3247
rect 3425 3243 3426 3247
rect 3428 3243 3429 3247
rect 3441 3243 3442 3247
rect 3444 3243 3445 3247
rect 3457 3243 3458 3247
rect 3460 3243 3463 3247
rect 3465 3243 3466 3247
rect 3478 3243 3479 3247
rect 3481 3243 3482 3247
rect 3494 3243 3495 3247
rect 3497 3243 3500 3247
rect 3502 3243 3503 3247
rect 3515 3243 3516 3247
rect 3518 3243 3519 3247
rect 3531 3243 3532 3247
rect 3534 3243 3537 3247
rect 3539 3243 3540 3247
rect 3557 3243 3558 3247
rect 3560 3243 3561 3247
rect 3573 3243 3574 3247
rect 3576 3243 3577 3247
rect 3589 3243 3590 3247
rect 3592 3243 3595 3247
rect 3597 3243 3598 3247
rect 3610 3243 3611 3247
rect 3613 3243 3614 3247
rect 2517 3199 2518 3203
rect 2520 3199 2521 3203
rect 2541 3199 2542 3203
rect 2544 3199 2545 3203
rect 3462 3199 3463 3203
rect 3465 3199 3466 3203
rect 3486 3199 3487 3203
rect 3489 3199 3490 3203
rect 2537 3188 2538 3192
rect 2540 3188 2541 3192
rect 3482 3188 3483 3192
rect 3485 3188 3486 3192
rect 2529 3176 2533 3177
rect 2529 3173 2533 3174
rect 3474 3176 3478 3177
rect 3474 3173 3478 3174
rect 2517 3165 2518 3169
rect 2520 3165 2521 3169
rect 2541 3165 2542 3169
rect 2544 3165 2545 3169
rect 3462 3165 3463 3169
rect 3465 3165 3466 3169
rect 3486 3165 3487 3169
rect 3489 3165 3490 3169
rect 2285 3103 2286 3107
rect 2288 3103 2291 3107
rect 2293 3103 2294 3107
rect 2306 3103 2307 3107
rect 2309 3103 2310 3107
rect 2322 3103 2323 3107
rect 2325 3103 2328 3107
rect 2330 3103 2331 3107
rect 2348 3103 2349 3107
rect 2351 3103 2352 3107
rect 2364 3103 2365 3107
rect 2367 3103 2368 3107
rect 2380 3103 2381 3107
rect 2383 3103 2386 3107
rect 2388 3103 2389 3107
rect 2401 3103 2402 3107
rect 2404 3103 2405 3107
rect 2417 3103 2418 3107
rect 2420 3103 2423 3107
rect 2425 3103 2426 3107
rect 2438 3103 2439 3107
rect 2441 3103 2442 3107
rect 2454 3103 2455 3107
rect 2457 3103 2460 3107
rect 2462 3103 2463 3107
rect 2480 3103 2481 3107
rect 2483 3103 2484 3107
rect 2496 3103 2497 3107
rect 2499 3103 2500 3107
rect 2512 3103 2513 3107
rect 2515 3103 2518 3107
rect 2520 3103 2521 3107
rect 2533 3103 2534 3107
rect 2536 3103 2537 3107
rect 2549 3103 2550 3107
rect 2552 3103 2555 3107
rect 2557 3103 2558 3107
rect 2570 3103 2571 3107
rect 2573 3103 2574 3107
rect 2586 3103 2587 3107
rect 2589 3103 2592 3107
rect 2594 3103 2595 3107
rect 2612 3103 2613 3107
rect 2615 3103 2616 3107
rect 2628 3103 2629 3107
rect 2631 3103 2632 3107
rect 2644 3103 2645 3107
rect 2647 3103 2650 3107
rect 2652 3103 2653 3107
rect 2665 3103 2666 3107
rect 2668 3103 2669 3107
rect 3230 3103 3231 3107
rect 3233 3103 3236 3107
rect 3238 3103 3239 3107
rect 3251 3103 3252 3107
rect 3254 3103 3255 3107
rect 3267 3103 3268 3107
rect 3270 3103 3273 3107
rect 3275 3103 3276 3107
rect 3293 3103 3294 3107
rect 3296 3103 3297 3107
rect 3309 3103 3310 3107
rect 3312 3103 3313 3107
rect 3325 3103 3326 3107
rect 3328 3103 3331 3107
rect 3333 3103 3334 3107
rect 3346 3103 3347 3107
rect 3349 3103 3350 3107
rect 3362 3103 3363 3107
rect 3365 3103 3368 3107
rect 3370 3103 3371 3107
rect 3383 3103 3384 3107
rect 3386 3103 3387 3107
rect 3399 3103 3400 3107
rect 3402 3103 3405 3107
rect 3407 3103 3408 3107
rect 3425 3103 3426 3107
rect 3428 3103 3429 3107
rect 3441 3103 3442 3107
rect 3444 3103 3445 3107
rect 3457 3103 3458 3107
rect 3460 3103 3463 3107
rect 3465 3103 3466 3107
rect 3478 3103 3479 3107
rect 3481 3103 3482 3107
rect 3494 3103 3495 3107
rect 3497 3103 3500 3107
rect 3502 3103 3503 3107
rect 3515 3103 3516 3107
rect 3518 3103 3519 3107
rect 3531 3103 3532 3107
rect 3534 3103 3537 3107
rect 3539 3103 3540 3107
rect 3557 3103 3558 3107
rect 3560 3103 3561 3107
rect 3573 3103 3574 3107
rect 3576 3103 3577 3107
rect 3589 3103 3590 3107
rect 3592 3103 3595 3107
rect 3597 3103 3598 3107
rect 3610 3103 3611 3107
rect 3613 3103 3614 3107
rect 2769 3024 2770 3028
rect 2772 3024 2775 3028
rect 2777 3024 2778 3028
rect 2790 3024 2791 3028
rect 2793 3024 2794 3028
rect 2806 3024 2807 3028
rect 2809 3024 2812 3028
rect 2814 3024 2815 3028
rect 2832 3024 2833 3028
rect 2835 3024 2836 3028
rect 2848 3024 2849 3028
rect 2851 3024 2852 3028
rect 2864 3024 2865 3028
rect 2867 3024 2870 3028
rect 2872 3024 2873 3028
rect 2885 3024 2886 3028
rect 2888 3024 2889 3028
rect 2901 3024 2902 3028
rect 2904 3024 2907 3028
rect 2909 3024 2910 3028
rect 2922 3024 2923 3028
rect 2925 3024 2926 3028
rect 2938 3024 2939 3028
rect 2941 3024 2944 3028
rect 2946 3024 2947 3028
rect 2964 3024 2965 3028
rect 2967 3024 2968 3028
rect 2980 3024 2981 3028
rect 2983 3024 2984 3028
rect 2996 3024 2997 3028
rect 2999 3024 3002 3028
rect 3004 3024 3005 3028
rect 3017 3024 3018 3028
rect 3020 3024 3021 3028
rect 3033 3024 3034 3028
rect 3036 3024 3039 3028
rect 3041 3024 3042 3028
rect 3054 3024 3055 3028
rect 3057 3024 3058 3028
rect 3070 3024 3071 3028
rect 3073 3024 3076 3028
rect 3078 3024 3079 3028
rect 3096 3024 3097 3028
rect 3099 3024 3100 3028
rect 3112 3024 3113 3028
rect 3115 3024 3116 3028
rect 3128 3024 3129 3028
rect 3131 3024 3134 3028
rect 3136 3024 3137 3028
rect 3149 3024 3150 3028
rect 3152 3024 3153 3028
rect 3165 3024 3166 3028
rect 3168 3024 3171 3028
rect 3173 3024 3174 3028
rect 3186 3024 3187 3028
rect 3189 3024 3190 3028
rect 3202 3024 3203 3028
rect 3205 3024 3208 3028
rect 3210 3024 3211 3028
rect 3228 3024 3229 3028
rect 3231 3024 3232 3028
rect 3244 3024 3245 3028
rect 3247 3024 3248 3028
rect 3260 3024 3261 3028
rect 3263 3024 3266 3028
rect 3268 3024 3269 3028
rect 3281 3024 3282 3028
rect 3284 3024 3285 3028
rect 3714 3024 3715 3028
rect 3717 3024 3720 3028
rect 3722 3024 3723 3028
rect 3735 3024 3736 3028
rect 3738 3024 3739 3028
rect 3751 3024 3752 3028
rect 3754 3024 3757 3028
rect 3759 3024 3760 3028
rect 3777 3024 3778 3028
rect 3780 3024 3781 3028
rect 3793 3024 3794 3028
rect 3796 3024 3797 3028
rect 3809 3024 3810 3028
rect 3812 3024 3815 3028
rect 3817 3024 3818 3028
rect 3830 3024 3831 3028
rect 3833 3024 3834 3028
rect 3846 3024 3847 3028
rect 3849 3024 3852 3028
rect 3854 3024 3855 3028
rect 3867 3024 3868 3028
rect 3870 3024 3871 3028
rect 3883 3024 3884 3028
rect 3886 3024 3889 3028
rect 3891 3024 3892 3028
rect 3909 3024 3910 3028
rect 3912 3024 3913 3028
rect 3925 3024 3926 3028
rect 3928 3024 3929 3028
rect 3941 3024 3942 3028
rect 3944 3024 3947 3028
rect 3949 3024 3950 3028
rect 3962 3024 3963 3028
rect 3965 3024 3966 3028
rect 3978 3024 3979 3028
rect 3981 3024 3984 3028
rect 3986 3024 3987 3028
rect 3999 3024 4000 3028
rect 4002 3024 4003 3028
rect 4015 3024 4016 3028
rect 4018 3024 4021 3028
rect 4023 3024 4024 3028
rect 4041 3024 4042 3028
rect 4044 3024 4045 3028
rect 4057 3024 4058 3028
rect 4060 3024 4061 3028
rect 4073 3024 4074 3028
rect 4076 3024 4079 3028
rect 4081 3024 4082 3028
rect 4094 3024 4095 3028
rect 4097 3024 4098 3028
rect 4110 3024 4111 3028
rect 4113 3024 4116 3028
rect 4118 3024 4119 3028
rect 4131 3024 4132 3028
rect 4134 3024 4135 3028
rect 4147 3024 4148 3028
rect 4150 3024 4153 3028
rect 4155 3024 4156 3028
rect 4173 3024 4174 3028
rect 4176 3024 4177 3028
rect 4189 3024 4190 3028
rect 4192 3024 4193 3028
rect 4205 3024 4206 3028
rect 4208 3024 4211 3028
rect 4213 3024 4214 3028
rect 4226 3024 4227 3028
rect 4229 3024 4230 3028
rect 2417 2991 2418 2995
rect 2420 2991 2423 2995
rect 2425 2991 2426 2995
rect 2438 2991 2439 2995
rect 2441 2991 2442 2995
rect 2454 2991 2455 2995
rect 2457 2991 2460 2995
rect 2462 2991 2463 2995
rect 2480 2991 2481 2995
rect 2483 2991 2484 2995
rect 2496 2991 2497 2995
rect 2499 2991 2500 2995
rect 2512 2991 2513 2995
rect 2515 2991 2518 2995
rect 2520 2991 2521 2995
rect 2533 2991 2534 2995
rect 2536 2991 2537 2995
rect 3362 2991 3363 2995
rect 3365 2991 3368 2995
rect 3370 2991 3371 2995
rect 3383 2991 3384 2995
rect 3386 2991 3387 2995
rect 3399 2991 3400 2995
rect 3402 2991 3405 2995
rect 3407 2991 3408 2995
rect 3425 2991 3426 2995
rect 3428 2991 3429 2995
rect 3441 2991 3442 2995
rect 3444 2991 3445 2995
rect 3457 2991 3458 2995
rect 3460 2991 3463 2995
rect 3465 2991 3466 2995
rect 3478 2991 3479 2995
rect 3481 2991 3482 2995
rect 2541 2954 2542 2958
rect 2544 2954 2545 2958
rect 2948 2958 2949 2962
rect 2951 2958 2952 2962
rect 2972 2954 2975 2958
rect 2977 2954 2980 2958
rect 2982 2954 2983 2958
rect 3029 2958 3030 2962
rect 3032 2958 3033 2962
rect 3053 2954 3056 2958
rect 3058 2954 3061 2958
rect 3063 2954 3064 2958
rect 3002 2950 3003 2954
rect 3005 2950 3006 2954
rect 2424 2945 2425 2949
rect 2427 2945 2428 2949
rect 2774 2945 2775 2949
rect 2777 2945 2778 2949
rect 2790 2945 2791 2949
rect 2793 2945 2794 2949
rect 2806 2945 2807 2949
rect 2809 2945 2810 2949
rect 2825 2945 2830 2949
rect 2832 2945 2835 2949
rect 2837 2945 2838 2949
rect 2859 2945 2861 2949
rect 2863 2945 2864 2949
rect 2881 2945 2882 2949
rect 2884 2945 2885 2949
rect 2897 2945 2902 2949
rect 2904 2945 2907 2949
rect 2909 2945 2910 2949
rect 2924 2945 2925 2949
rect 2927 2945 2928 2949
rect 3083 2950 3084 2954
rect 3086 2950 3087 2954
rect 3486 2954 3487 2958
rect 3489 2954 3490 2958
rect 3893 2958 3894 2962
rect 3896 2958 3897 2962
rect 3917 2954 3920 2958
rect 3922 2954 3925 2958
rect 3927 2954 3928 2958
rect 3974 2958 3975 2962
rect 3977 2958 3978 2962
rect 3998 2954 4001 2958
rect 4003 2954 4006 2958
rect 4008 2954 4009 2958
rect 3947 2950 3948 2954
rect 3950 2950 3951 2954
rect 3369 2945 3370 2949
rect 3372 2945 3373 2949
rect 3719 2945 3720 2949
rect 3722 2945 3723 2949
rect 3735 2945 3736 2949
rect 3738 2945 3739 2949
rect 3751 2945 3752 2949
rect 3754 2945 3755 2949
rect 3770 2945 3775 2949
rect 3777 2945 3780 2949
rect 3782 2945 3783 2949
rect 3804 2945 3806 2949
rect 3808 2945 3809 2949
rect 3826 2945 3827 2949
rect 3829 2945 3830 2949
rect 3842 2945 3847 2949
rect 3849 2945 3852 2949
rect 3854 2945 3855 2949
rect 3869 2945 3870 2949
rect 3872 2945 3873 2949
rect 4028 2950 4029 2954
rect 4031 2950 4032 2954
rect 2774 2899 2775 2903
rect 2777 2899 2778 2903
rect 2790 2899 2791 2903
rect 2793 2899 2794 2903
rect 2806 2899 2807 2903
rect 2809 2899 2810 2903
rect 2825 2899 2830 2903
rect 2832 2899 2835 2903
rect 2837 2899 2838 2903
rect 2859 2899 2861 2903
rect 2863 2899 2864 2903
rect 2881 2899 2882 2903
rect 2884 2899 2885 2903
rect 2897 2899 2902 2903
rect 2904 2899 2907 2903
rect 2909 2899 2910 2903
rect 2924 2899 2925 2903
rect 2927 2899 2928 2903
rect 2408 2889 2409 2893
rect 2411 2889 2412 2893
rect 2424 2889 2425 2893
rect 2427 2889 2430 2893
rect 2432 2889 2433 2893
rect 2445 2889 2446 2893
rect 2448 2889 2449 2893
rect 2461 2889 2462 2893
rect 2464 2889 2465 2893
rect 2482 2889 2483 2893
rect 2485 2889 2488 2893
rect 2490 2889 2491 2893
rect 2503 2889 2504 2893
rect 2506 2889 2507 2893
rect 2519 2889 2520 2893
rect 2522 2889 2525 2893
rect 2527 2889 2528 2893
rect 2972 2898 2975 2902
rect 2977 2898 2980 2902
rect 2982 2898 2983 2902
rect 3053 2898 3056 2902
rect 3058 2898 3061 2902
rect 3063 2898 3064 2902
rect 3719 2899 3720 2903
rect 3722 2899 3723 2903
rect 3735 2899 3736 2903
rect 3738 2899 3739 2903
rect 3751 2899 3752 2903
rect 3754 2899 3755 2903
rect 3770 2899 3775 2903
rect 3777 2899 3780 2903
rect 3782 2899 3783 2903
rect 3804 2899 3806 2903
rect 3808 2899 3809 2903
rect 3826 2899 3827 2903
rect 3829 2899 3830 2903
rect 3842 2899 3847 2903
rect 3849 2899 3852 2903
rect 3854 2899 3855 2903
rect 3869 2899 3870 2903
rect 3872 2899 3873 2903
rect 3353 2889 3354 2893
rect 3356 2889 3357 2893
rect 3369 2889 3370 2893
rect 3372 2889 3375 2893
rect 3377 2889 3378 2893
rect 3390 2889 3391 2893
rect 3393 2889 3394 2893
rect 3406 2889 3407 2893
rect 3409 2889 3410 2893
rect 3427 2889 3428 2893
rect 3430 2889 3433 2893
rect 3435 2889 3436 2893
rect 3448 2889 3449 2893
rect 3451 2889 3452 2893
rect 3464 2889 3465 2893
rect 3467 2889 3470 2893
rect 3472 2889 3473 2893
rect 3917 2898 3920 2902
rect 3922 2898 3925 2902
rect 3927 2898 3928 2902
rect 3998 2898 4001 2902
rect 4003 2898 4006 2902
rect 4008 2898 4009 2902
rect 2972 2822 2975 2826
rect 2977 2822 2980 2826
rect 2982 2822 2983 2826
rect 3053 2826 3054 2830
rect 3056 2826 3057 2830
rect 3077 2822 3080 2826
rect 3082 2822 3085 2826
rect 3087 2822 3088 2826
rect 3002 2818 3003 2822
rect 3005 2818 3006 2822
rect 2774 2813 2775 2817
rect 2777 2813 2778 2817
rect 2790 2813 2791 2817
rect 2793 2813 2794 2817
rect 2806 2813 2807 2817
rect 2809 2813 2810 2817
rect 2825 2813 2830 2817
rect 2832 2813 2835 2817
rect 2837 2813 2838 2817
rect 2859 2813 2861 2817
rect 2863 2813 2864 2817
rect 2881 2813 2882 2817
rect 2884 2813 2885 2817
rect 2897 2813 2902 2817
rect 2904 2813 2907 2817
rect 2909 2813 2910 2817
rect 2924 2813 2925 2817
rect 2927 2813 2928 2817
rect 3107 2818 3108 2822
rect 3110 2818 3111 2822
rect 3917 2822 3920 2826
rect 3922 2822 3925 2826
rect 3927 2822 3928 2826
rect 3998 2826 3999 2830
rect 4001 2826 4002 2830
rect 4022 2822 4025 2826
rect 4027 2822 4030 2826
rect 4032 2822 4033 2826
rect 3947 2818 3948 2822
rect 3950 2818 3951 2822
rect 3719 2813 3720 2817
rect 3722 2813 3723 2817
rect 3735 2813 3736 2817
rect 3738 2813 3739 2817
rect 3751 2813 3752 2817
rect 3754 2813 3755 2817
rect 3770 2813 3775 2817
rect 3777 2813 3780 2817
rect 3782 2813 3783 2817
rect 3804 2813 3806 2817
rect 3808 2813 3809 2817
rect 3826 2813 3827 2817
rect 3829 2813 3830 2817
rect 3842 2813 3847 2817
rect 3849 2813 3852 2817
rect 3854 2813 3855 2817
rect 3869 2813 3870 2817
rect 3872 2813 3873 2817
rect 4052 2818 4053 2822
rect 4055 2818 4056 2822
rect 2774 2767 2775 2771
rect 2777 2767 2778 2771
rect 2790 2767 2791 2771
rect 2793 2767 2794 2771
rect 2806 2767 2807 2771
rect 2809 2767 2810 2771
rect 2825 2767 2830 2771
rect 2832 2767 2835 2771
rect 2837 2767 2838 2771
rect 2859 2767 2861 2771
rect 2863 2767 2864 2771
rect 2881 2767 2882 2771
rect 2884 2767 2885 2771
rect 2897 2767 2902 2771
rect 2904 2767 2907 2771
rect 2909 2767 2910 2771
rect 2924 2767 2925 2771
rect 2927 2767 2928 2771
rect 2972 2767 2975 2771
rect 2977 2767 2980 2771
rect 2982 2767 2983 2771
rect 3077 2767 3080 2771
rect 3082 2767 3085 2771
rect 3087 2767 3088 2771
rect 3719 2767 3720 2771
rect 3722 2767 3723 2771
rect 3735 2767 3736 2771
rect 3738 2767 3739 2771
rect 3751 2767 3752 2771
rect 3754 2767 3755 2771
rect 3770 2767 3775 2771
rect 3777 2767 3780 2771
rect 3782 2767 3783 2771
rect 3804 2767 3806 2771
rect 3808 2767 3809 2771
rect 3826 2767 3827 2771
rect 3829 2767 3830 2771
rect 3842 2767 3847 2771
rect 3849 2767 3852 2771
rect 3854 2767 3855 2771
rect 3869 2767 3870 2771
rect 3872 2767 3873 2771
rect 3917 2767 3920 2771
rect 3922 2767 3925 2771
rect 3927 2767 3928 2771
rect 4022 2767 4025 2771
rect 4027 2767 4030 2771
rect 4032 2767 4033 2771
rect 2972 2690 2975 2694
rect 2977 2690 2980 2694
rect 2982 2690 2983 2694
rect 3029 2694 3030 2698
rect 3032 2694 3033 2698
rect 3053 2690 3056 2694
rect 3058 2690 3061 2694
rect 3063 2690 3064 2694
rect 3119 2694 3120 2698
rect 3122 2694 3123 2698
rect 3143 2690 3146 2694
rect 3148 2690 3151 2694
rect 3153 2690 3154 2694
rect 3002 2686 3003 2690
rect 3005 2686 3006 2690
rect 2774 2681 2775 2685
rect 2777 2681 2778 2685
rect 2790 2681 2791 2685
rect 2793 2681 2794 2685
rect 2806 2681 2807 2685
rect 2809 2681 2810 2685
rect 2825 2681 2830 2685
rect 2832 2681 2835 2685
rect 2837 2681 2838 2685
rect 2859 2681 2861 2685
rect 2863 2681 2864 2685
rect 2881 2681 2882 2685
rect 2884 2681 2885 2685
rect 2897 2681 2902 2685
rect 2904 2681 2907 2685
rect 2909 2681 2910 2685
rect 2924 2681 2925 2685
rect 2927 2681 2928 2685
rect 3083 2686 3084 2690
rect 3086 2686 3087 2690
rect 3173 2686 3174 2690
rect 3176 2686 3177 2690
rect 3917 2690 3920 2694
rect 3922 2690 3925 2694
rect 3927 2690 3928 2694
rect 3974 2694 3975 2698
rect 3977 2694 3978 2698
rect 3998 2690 4001 2694
rect 4003 2690 4006 2694
rect 4008 2690 4009 2694
rect 4064 2694 4065 2698
rect 4067 2694 4068 2698
rect 4088 2690 4091 2694
rect 4093 2690 4096 2694
rect 4098 2690 4099 2694
rect 3947 2686 3948 2690
rect 3950 2686 3951 2690
rect 3719 2681 3720 2685
rect 3722 2681 3723 2685
rect 3735 2681 3736 2685
rect 3738 2681 3739 2685
rect 3751 2681 3752 2685
rect 3754 2681 3755 2685
rect 3770 2681 3775 2685
rect 3777 2681 3780 2685
rect 3782 2681 3783 2685
rect 3804 2681 3806 2685
rect 3808 2681 3809 2685
rect 3826 2681 3827 2685
rect 3829 2681 3830 2685
rect 3842 2681 3847 2685
rect 3849 2681 3852 2685
rect 3854 2681 3855 2685
rect 3869 2681 3870 2685
rect 3872 2681 3873 2685
rect 4028 2686 4029 2690
rect 4031 2686 4032 2690
rect 4118 2686 4119 2690
rect 4121 2686 4122 2690
rect 2774 2635 2775 2639
rect 2777 2635 2778 2639
rect 2790 2635 2791 2639
rect 2793 2635 2794 2639
rect 2806 2635 2807 2639
rect 2809 2635 2810 2639
rect 2825 2635 2830 2639
rect 2832 2635 2835 2639
rect 2837 2635 2838 2639
rect 2859 2635 2861 2639
rect 2863 2635 2864 2639
rect 2881 2635 2882 2639
rect 2884 2635 2885 2639
rect 2897 2635 2902 2639
rect 2904 2635 2907 2639
rect 2909 2635 2910 2639
rect 2924 2635 2925 2639
rect 2927 2635 2928 2639
rect 2972 2632 2975 2636
rect 2977 2632 2980 2636
rect 2982 2632 2983 2636
rect 3053 2632 3056 2636
rect 3058 2632 3061 2636
rect 3063 2632 3064 2636
rect 3143 2632 3146 2636
rect 3148 2632 3151 2636
rect 3153 2632 3154 2636
rect 3719 2635 3720 2639
rect 3722 2635 3723 2639
rect 3735 2635 3736 2639
rect 3738 2635 3739 2639
rect 3751 2635 3752 2639
rect 3754 2635 3755 2639
rect 3770 2635 3775 2639
rect 3777 2635 3780 2639
rect 3782 2635 3783 2639
rect 3804 2635 3806 2639
rect 3808 2635 3809 2639
rect 3826 2635 3827 2639
rect 3829 2635 3830 2639
rect 3842 2635 3847 2639
rect 3849 2635 3852 2639
rect 3854 2635 3855 2639
rect 3869 2635 3870 2639
rect 3872 2635 3873 2639
rect 3917 2632 3920 2636
rect 3922 2632 3925 2636
rect 3927 2632 3928 2636
rect 3998 2632 4001 2636
rect 4003 2632 4006 2636
rect 4008 2632 4009 2636
rect 4088 2632 4091 2636
rect 4093 2632 4096 2636
rect 4098 2632 4099 2636
rect 2972 2558 2975 2562
rect 2977 2558 2980 2562
rect 2982 2558 2983 2562
rect 3002 2554 3003 2558
rect 3005 2554 3006 2558
rect 2774 2549 2775 2553
rect 2777 2549 2778 2553
rect 2790 2549 2791 2553
rect 2793 2549 2794 2553
rect 2806 2549 2807 2553
rect 2809 2549 2810 2553
rect 2825 2549 2830 2553
rect 2832 2549 2835 2553
rect 2837 2549 2838 2553
rect 2859 2549 2861 2553
rect 2863 2549 2864 2553
rect 2881 2549 2882 2553
rect 2884 2549 2885 2553
rect 2897 2549 2902 2553
rect 2904 2549 2907 2553
rect 2909 2549 2910 2553
rect 2924 2549 2925 2553
rect 2927 2549 2928 2553
rect 3917 2558 3920 2562
rect 3922 2558 3925 2562
rect 3927 2558 3928 2562
rect 3947 2554 3948 2558
rect 3950 2554 3951 2558
rect 3719 2549 3720 2553
rect 3722 2549 3723 2553
rect 3735 2549 3736 2553
rect 3738 2549 3739 2553
rect 3751 2549 3752 2553
rect 3754 2549 3755 2553
rect 3770 2549 3775 2553
rect 3777 2549 3780 2553
rect 3782 2549 3783 2553
rect 3804 2549 3806 2553
rect 3808 2549 3809 2553
rect 3826 2549 3827 2553
rect 3829 2549 3830 2553
rect 3842 2549 3847 2553
rect 3849 2549 3852 2553
rect 3854 2549 3855 2553
rect 3869 2549 3870 2553
rect 3872 2549 3873 2553
rect 2774 2503 2775 2507
rect 2777 2503 2778 2507
rect 2790 2503 2791 2507
rect 2793 2503 2794 2507
rect 2806 2503 2807 2507
rect 2809 2503 2810 2507
rect 2825 2503 2830 2507
rect 2832 2503 2835 2507
rect 2837 2503 2838 2507
rect 2859 2503 2861 2507
rect 2863 2503 2864 2507
rect 2881 2503 2882 2507
rect 2884 2503 2885 2507
rect 2897 2503 2902 2507
rect 2904 2503 2907 2507
rect 2909 2503 2910 2507
rect 2924 2503 2925 2507
rect 2927 2503 2928 2507
rect 3008 2503 3009 2507
rect 3011 2503 3012 2507
rect 3016 2503 3022 2507
rect 3026 2503 3027 2507
rect 3029 2503 3030 2507
rect 3051 2503 3052 2507
rect 3054 2503 3055 2507
rect 3067 2503 3068 2507
rect 3070 2503 3071 2507
rect 3086 2503 3091 2507
rect 3093 2503 3096 2507
rect 3098 2503 3099 2507
rect 3120 2503 3122 2507
rect 3124 2503 3125 2507
rect 3142 2503 3143 2507
rect 3145 2503 3146 2507
rect 3158 2503 3163 2507
rect 3165 2503 3168 2507
rect 3170 2503 3171 2507
rect 3185 2503 3186 2507
rect 3188 2503 3189 2507
rect 2285 2489 2286 2493
rect 2288 2489 2291 2493
rect 2293 2489 2294 2493
rect 2306 2489 2307 2493
rect 2309 2489 2310 2493
rect 2322 2489 2323 2493
rect 2325 2489 2328 2493
rect 2330 2489 2331 2493
rect 2348 2489 2349 2493
rect 2351 2489 2352 2493
rect 2364 2489 2365 2493
rect 2367 2489 2368 2493
rect 2380 2489 2381 2493
rect 2383 2489 2386 2493
rect 2388 2489 2389 2493
rect 2401 2489 2402 2493
rect 2404 2489 2405 2493
rect 2417 2489 2418 2493
rect 2420 2489 2423 2493
rect 2425 2489 2426 2493
rect 2438 2489 2439 2493
rect 2441 2489 2442 2493
rect 2454 2489 2455 2493
rect 2457 2489 2460 2493
rect 2462 2489 2463 2493
rect 2480 2489 2481 2493
rect 2483 2489 2484 2493
rect 2496 2489 2497 2493
rect 2499 2489 2500 2493
rect 2512 2489 2513 2493
rect 2515 2489 2518 2493
rect 2520 2489 2521 2493
rect 2533 2489 2534 2493
rect 2536 2489 2537 2493
rect 2549 2489 2550 2493
rect 2552 2489 2555 2493
rect 2557 2489 2558 2493
rect 2570 2489 2571 2493
rect 2573 2489 2574 2493
rect 2586 2489 2587 2493
rect 2589 2489 2592 2493
rect 2594 2489 2595 2493
rect 2612 2489 2613 2493
rect 2615 2489 2616 2493
rect 2628 2489 2629 2493
rect 2631 2489 2632 2493
rect 2644 2489 2645 2493
rect 2647 2489 2650 2493
rect 2652 2489 2653 2493
rect 2665 2489 2666 2493
rect 2668 2489 2669 2493
rect 2972 2496 2975 2500
rect 2977 2496 2980 2500
rect 2982 2496 2983 2500
rect 3719 2503 3720 2507
rect 3722 2503 3723 2507
rect 3735 2503 3736 2507
rect 3738 2503 3739 2507
rect 3751 2503 3752 2507
rect 3754 2503 3755 2507
rect 3770 2503 3775 2507
rect 3777 2503 3780 2507
rect 3782 2503 3783 2507
rect 3804 2503 3806 2507
rect 3808 2503 3809 2507
rect 3826 2503 3827 2507
rect 3829 2503 3830 2507
rect 3842 2503 3847 2507
rect 3849 2503 3852 2507
rect 3854 2503 3855 2507
rect 3869 2503 3870 2507
rect 3872 2503 3873 2507
rect 3953 2503 3954 2507
rect 3956 2503 3957 2507
rect 3961 2503 3967 2507
rect 3971 2503 3972 2507
rect 3974 2503 3975 2507
rect 3996 2503 3997 2507
rect 3999 2503 4000 2507
rect 4012 2503 4013 2507
rect 4015 2503 4016 2507
rect 4031 2503 4036 2507
rect 4038 2503 4041 2507
rect 4043 2503 4044 2507
rect 4065 2503 4067 2507
rect 4069 2503 4070 2507
rect 4087 2503 4088 2507
rect 4090 2503 4091 2507
rect 4103 2503 4108 2507
rect 4110 2503 4113 2507
rect 4115 2503 4116 2507
rect 4130 2503 4131 2507
rect 4133 2503 4134 2507
rect 3230 2489 3231 2493
rect 3233 2489 3236 2493
rect 3238 2489 3239 2493
rect 3251 2489 3252 2493
rect 3254 2489 3255 2493
rect 3267 2489 3268 2493
rect 3270 2489 3273 2493
rect 3275 2489 3276 2493
rect 3293 2489 3294 2493
rect 3296 2489 3297 2493
rect 3309 2489 3310 2493
rect 3312 2489 3313 2493
rect 3325 2489 3326 2493
rect 3328 2489 3331 2493
rect 3333 2489 3334 2493
rect 3346 2489 3347 2493
rect 3349 2489 3350 2493
rect 3362 2489 3363 2493
rect 3365 2489 3368 2493
rect 3370 2489 3371 2493
rect 3383 2489 3384 2493
rect 3386 2489 3387 2493
rect 3399 2489 3400 2493
rect 3402 2489 3405 2493
rect 3407 2489 3408 2493
rect 3425 2489 3426 2493
rect 3428 2489 3429 2493
rect 3441 2489 3442 2493
rect 3444 2489 3445 2493
rect 3457 2489 3458 2493
rect 3460 2489 3463 2493
rect 3465 2489 3466 2493
rect 3478 2489 3479 2493
rect 3481 2489 3482 2493
rect 3494 2489 3495 2493
rect 3497 2489 3500 2493
rect 3502 2489 3503 2493
rect 3515 2489 3516 2493
rect 3518 2489 3519 2493
rect 3531 2489 3532 2493
rect 3534 2489 3537 2493
rect 3539 2489 3540 2493
rect 3557 2489 3558 2493
rect 3560 2489 3561 2493
rect 3573 2489 3574 2493
rect 3576 2489 3577 2493
rect 3589 2489 3590 2493
rect 3592 2489 3595 2493
rect 3597 2489 3598 2493
rect 3610 2489 3611 2493
rect 3613 2489 3614 2493
rect 3917 2496 3920 2500
rect 3922 2496 3925 2500
rect 3927 2496 3928 2500
rect 2400 2445 2401 2449
rect 2403 2445 2404 2449
rect 2424 2445 2425 2449
rect 2427 2445 2428 2449
rect 3198 2449 3202 2450
rect 3198 2446 3202 2447
rect 3345 2445 3346 2449
rect 3348 2445 3349 2449
rect 3369 2445 3370 2449
rect 3372 2445 3373 2449
rect 4143 2449 4147 2450
rect 4143 2446 4147 2447
rect 2420 2432 2421 2436
rect 2423 2432 2424 2436
rect 3365 2432 3366 2436
rect 3368 2432 3369 2436
rect 2412 2420 2416 2421
rect 2412 2417 2416 2418
rect 3357 2420 3361 2421
rect 3357 2417 3361 2418
rect 2400 2409 2401 2413
rect 2403 2409 2404 2413
rect 2424 2409 2425 2413
rect 2427 2409 2428 2413
rect 3345 2409 3346 2413
rect 3348 2409 3349 2413
rect 3369 2409 3370 2413
rect 3372 2409 3373 2413
rect 3068 2377 3069 2381
rect 3071 2377 3074 2381
rect 3076 2377 3077 2381
rect 3089 2377 3090 2381
rect 3092 2377 3093 2381
rect 3105 2377 3106 2381
rect 3108 2377 3111 2381
rect 3113 2377 3114 2381
rect 3131 2377 3132 2381
rect 3134 2377 3135 2381
rect 3147 2377 3148 2381
rect 3150 2377 3151 2381
rect 3163 2377 3164 2381
rect 3166 2377 3169 2381
rect 3171 2377 3172 2381
rect 3184 2377 3185 2381
rect 3187 2377 3188 2381
rect 4013 2377 4014 2381
rect 4016 2377 4019 2381
rect 4021 2377 4022 2381
rect 4034 2377 4035 2381
rect 4037 2377 4038 2381
rect 4050 2377 4051 2381
rect 4053 2377 4056 2381
rect 4058 2377 4059 2381
rect 4076 2377 4077 2381
rect 4079 2377 4080 2381
rect 4092 2377 4093 2381
rect 4095 2377 4096 2381
rect 4108 2377 4109 2381
rect 4111 2377 4114 2381
rect 4116 2377 4117 2381
rect 4129 2377 4130 2381
rect 4132 2377 4133 2381
rect 2285 2347 2286 2351
rect 2288 2347 2291 2351
rect 2293 2347 2294 2351
rect 2306 2347 2307 2351
rect 2309 2347 2310 2351
rect 2322 2347 2323 2351
rect 2325 2347 2328 2351
rect 2330 2347 2331 2351
rect 2348 2347 2349 2351
rect 2351 2347 2352 2351
rect 2364 2347 2365 2351
rect 2367 2347 2368 2351
rect 2380 2347 2381 2351
rect 2383 2347 2386 2351
rect 2388 2347 2389 2351
rect 2401 2347 2402 2351
rect 2404 2347 2405 2351
rect 2417 2347 2418 2351
rect 2420 2347 2423 2351
rect 2425 2347 2426 2351
rect 2438 2347 2439 2351
rect 2441 2347 2442 2351
rect 2454 2347 2455 2351
rect 2457 2347 2460 2351
rect 2462 2347 2463 2351
rect 2480 2347 2481 2351
rect 2483 2347 2484 2351
rect 2496 2347 2497 2351
rect 2499 2347 2500 2351
rect 2512 2347 2513 2351
rect 2515 2347 2518 2351
rect 2520 2347 2521 2351
rect 2533 2347 2534 2351
rect 2536 2347 2537 2351
rect 2549 2347 2550 2351
rect 2552 2347 2555 2351
rect 2557 2347 2558 2351
rect 2570 2347 2571 2351
rect 2573 2347 2574 2351
rect 2586 2347 2587 2351
rect 2589 2347 2592 2351
rect 2594 2347 2595 2351
rect 2612 2347 2613 2351
rect 2615 2347 2616 2351
rect 2628 2347 2629 2351
rect 2631 2347 2632 2351
rect 2644 2347 2645 2351
rect 2647 2347 2650 2351
rect 2652 2347 2653 2351
rect 2665 2347 2666 2351
rect 2668 2347 2669 2351
rect 3230 2347 3231 2351
rect 3233 2347 3236 2351
rect 3238 2347 3239 2351
rect 3251 2347 3252 2351
rect 3254 2347 3255 2351
rect 3267 2347 3268 2351
rect 3270 2347 3273 2351
rect 3275 2347 3276 2351
rect 3293 2347 3294 2351
rect 3296 2347 3297 2351
rect 3309 2347 3310 2351
rect 3312 2347 3313 2351
rect 3325 2347 3326 2351
rect 3328 2347 3331 2351
rect 3333 2347 3334 2351
rect 3346 2347 3347 2351
rect 3349 2347 3350 2351
rect 3362 2347 3363 2351
rect 3365 2347 3368 2351
rect 3370 2347 3371 2351
rect 3383 2347 3384 2351
rect 3386 2347 3387 2351
rect 3399 2347 3400 2351
rect 3402 2347 3405 2351
rect 3407 2347 3408 2351
rect 3425 2347 3426 2351
rect 3428 2347 3429 2351
rect 3441 2347 3442 2351
rect 3444 2347 3445 2351
rect 3457 2347 3458 2351
rect 3460 2347 3463 2351
rect 3465 2347 3466 2351
rect 3478 2347 3479 2351
rect 3481 2347 3482 2351
rect 3494 2347 3495 2351
rect 3497 2347 3500 2351
rect 3502 2347 3503 2351
rect 3515 2347 3516 2351
rect 3518 2347 3519 2351
rect 3531 2347 3532 2351
rect 3534 2347 3537 2351
rect 3539 2347 3540 2351
rect 3557 2347 3558 2351
rect 3560 2347 3561 2351
rect 3573 2347 3574 2351
rect 3576 2347 3577 2351
rect 3589 2347 3590 2351
rect 3592 2347 3595 2351
rect 3597 2347 3598 2351
rect 3610 2347 3611 2351
rect 3613 2347 3614 2351
rect 3210 2303 3214 2304
rect 3210 2300 3214 2301
rect 4155 2303 4159 2304
rect 4155 2300 4159 2301
rect 3068 2291 3069 2295
rect 3071 2291 3074 2295
rect 3076 2291 3077 2295
rect 3089 2291 3090 2295
rect 3092 2291 3093 2295
rect 3105 2291 3106 2295
rect 3108 2291 3111 2295
rect 3113 2291 3114 2295
rect 3131 2291 3132 2295
rect 3134 2291 3135 2295
rect 3147 2291 3148 2295
rect 3150 2291 3151 2295
rect 3163 2291 3164 2295
rect 3166 2291 3169 2295
rect 3171 2291 3172 2295
rect 3184 2291 3185 2295
rect 3187 2291 3188 2295
rect 4013 2291 4014 2295
rect 4016 2291 4019 2295
rect 4021 2291 4022 2295
rect 4034 2291 4035 2295
rect 4037 2291 4038 2295
rect 4050 2291 4051 2295
rect 4053 2291 4056 2295
rect 4058 2291 4059 2295
rect 4076 2291 4077 2295
rect 4079 2291 4080 2295
rect 4092 2291 4093 2295
rect 4095 2291 4096 2295
rect 4108 2291 4109 2295
rect 4111 2291 4114 2295
rect 4116 2291 4117 2295
rect 4129 2291 4130 2295
rect 4132 2291 4133 2295
rect 2285 2261 2286 2265
rect 2288 2261 2291 2265
rect 2293 2261 2294 2265
rect 2306 2261 2307 2265
rect 2309 2261 2310 2265
rect 2322 2261 2323 2265
rect 2325 2261 2328 2265
rect 2330 2261 2331 2265
rect 2348 2261 2349 2265
rect 2351 2261 2352 2265
rect 2364 2261 2365 2265
rect 2367 2261 2368 2265
rect 2380 2261 2381 2265
rect 2383 2261 2386 2265
rect 2388 2261 2389 2265
rect 2401 2261 2402 2265
rect 2404 2261 2405 2265
rect 2417 2261 2418 2265
rect 2420 2261 2423 2265
rect 2425 2261 2426 2265
rect 2438 2261 2439 2265
rect 2441 2261 2442 2265
rect 2454 2261 2455 2265
rect 2457 2261 2460 2265
rect 2462 2261 2463 2265
rect 2480 2261 2481 2265
rect 2483 2261 2484 2265
rect 2496 2261 2497 2265
rect 2499 2261 2500 2265
rect 2512 2261 2513 2265
rect 2515 2261 2518 2265
rect 2520 2261 2521 2265
rect 2533 2261 2534 2265
rect 2536 2261 2537 2265
rect 2549 2261 2550 2265
rect 2552 2261 2555 2265
rect 2557 2261 2558 2265
rect 2570 2261 2571 2265
rect 2573 2261 2574 2265
rect 2586 2261 2587 2265
rect 2589 2261 2592 2265
rect 2594 2261 2595 2265
rect 2612 2261 2613 2265
rect 2615 2261 2616 2265
rect 2628 2261 2629 2265
rect 2631 2261 2632 2265
rect 2644 2261 2645 2265
rect 2647 2261 2650 2265
rect 2652 2261 2653 2265
rect 2665 2261 2666 2265
rect 2668 2261 2669 2265
rect 3230 2261 3231 2265
rect 3233 2261 3236 2265
rect 3238 2261 3239 2265
rect 3251 2261 3252 2265
rect 3254 2261 3255 2265
rect 3267 2261 3268 2265
rect 3270 2261 3273 2265
rect 3275 2261 3276 2265
rect 3293 2261 3294 2265
rect 3296 2261 3297 2265
rect 3309 2261 3310 2265
rect 3312 2261 3313 2265
rect 3325 2261 3326 2265
rect 3328 2261 3331 2265
rect 3333 2261 3334 2265
rect 3346 2261 3347 2265
rect 3349 2261 3350 2265
rect 3362 2261 3363 2265
rect 3365 2261 3368 2265
rect 3370 2261 3371 2265
rect 3383 2261 3384 2265
rect 3386 2261 3387 2265
rect 3399 2261 3400 2265
rect 3402 2261 3405 2265
rect 3407 2261 3408 2265
rect 3425 2261 3426 2265
rect 3428 2261 3429 2265
rect 3441 2261 3442 2265
rect 3444 2261 3445 2265
rect 3457 2261 3458 2265
rect 3460 2261 3463 2265
rect 3465 2261 3466 2265
rect 3478 2261 3479 2265
rect 3481 2261 3482 2265
rect 3494 2261 3495 2265
rect 3497 2261 3500 2265
rect 3502 2261 3503 2265
rect 3515 2261 3516 2265
rect 3518 2261 3519 2265
rect 3531 2261 3532 2265
rect 3534 2261 3537 2265
rect 3539 2261 3540 2265
rect 3557 2261 3558 2265
rect 3560 2261 3561 2265
rect 3573 2261 3574 2265
rect 3576 2261 3577 2265
rect 3589 2261 3590 2265
rect 3592 2261 3595 2265
rect 3597 2261 3598 2265
rect 3610 2261 3611 2265
rect 3613 2261 3614 2265
rect 2517 2217 2518 2221
rect 2520 2217 2521 2221
rect 2541 2217 2542 2221
rect 2544 2217 2545 2221
rect 3462 2217 3463 2221
rect 3465 2217 3466 2221
rect 3486 2217 3487 2221
rect 3489 2217 3490 2221
rect 2537 2206 2538 2210
rect 2540 2206 2541 2210
rect 3482 2206 3483 2210
rect 3485 2206 3486 2210
rect 2529 2194 2533 2195
rect 2529 2191 2533 2192
rect 3474 2194 3478 2195
rect 3474 2191 3478 2192
rect 2517 2183 2518 2187
rect 2520 2183 2521 2187
rect 2541 2183 2542 2187
rect 2544 2183 2545 2187
rect 3462 2183 3463 2187
rect 3465 2183 3466 2187
rect 3486 2183 3487 2187
rect 3489 2183 3490 2187
rect 2285 2121 2286 2125
rect 2288 2121 2291 2125
rect 2293 2121 2294 2125
rect 2306 2121 2307 2125
rect 2309 2121 2310 2125
rect 2322 2121 2323 2125
rect 2325 2121 2328 2125
rect 2330 2121 2331 2125
rect 2348 2121 2349 2125
rect 2351 2121 2352 2125
rect 2364 2121 2365 2125
rect 2367 2121 2368 2125
rect 2380 2121 2381 2125
rect 2383 2121 2386 2125
rect 2388 2121 2389 2125
rect 2401 2121 2402 2125
rect 2404 2121 2405 2125
rect 2417 2121 2418 2125
rect 2420 2121 2423 2125
rect 2425 2121 2426 2125
rect 2438 2121 2439 2125
rect 2441 2121 2442 2125
rect 2454 2121 2455 2125
rect 2457 2121 2460 2125
rect 2462 2121 2463 2125
rect 2480 2121 2481 2125
rect 2483 2121 2484 2125
rect 2496 2121 2497 2125
rect 2499 2121 2500 2125
rect 2512 2121 2513 2125
rect 2515 2121 2518 2125
rect 2520 2121 2521 2125
rect 2533 2121 2534 2125
rect 2536 2121 2537 2125
rect 2549 2121 2550 2125
rect 2552 2121 2555 2125
rect 2557 2121 2558 2125
rect 2570 2121 2571 2125
rect 2573 2121 2574 2125
rect 2586 2121 2587 2125
rect 2589 2121 2592 2125
rect 2594 2121 2595 2125
rect 2612 2121 2613 2125
rect 2615 2121 2616 2125
rect 2628 2121 2629 2125
rect 2631 2121 2632 2125
rect 2644 2121 2645 2125
rect 2647 2121 2650 2125
rect 2652 2121 2653 2125
rect 2665 2121 2666 2125
rect 2668 2121 2669 2125
rect 3230 2121 3231 2125
rect 3233 2121 3236 2125
rect 3238 2121 3239 2125
rect 3251 2121 3252 2125
rect 3254 2121 3255 2125
rect 3267 2121 3268 2125
rect 3270 2121 3273 2125
rect 3275 2121 3276 2125
rect 3293 2121 3294 2125
rect 3296 2121 3297 2125
rect 3309 2121 3310 2125
rect 3312 2121 3313 2125
rect 3325 2121 3326 2125
rect 3328 2121 3331 2125
rect 3333 2121 3334 2125
rect 3346 2121 3347 2125
rect 3349 2121 3350 2125
rect 3362 2121 3363 2125
rect 3365 2121 3368 2125
rect 3370 2121 3371 2125
rect 3383 2121 3384 2125
rect 3386 2121 3387 2125
rect 3399 2121 3400 2125
rect 3402 2121 3405 2125
rect 3407 2121 3408 2125
rect 3425 2121 3426 2125
rect 3428 2121 3429 2125
rect 3441 2121 3442 2125
rect 3444 2121 3445 2125
rect 3457 2121 3458 2125
rect 3460 2121 3463 2125
rect 3465 2121 3466 2125
rect 3478 2121 3479 2125
rect 3481 2121 3482 2125
rect 3494 2121 3495 2125
rect 3497 2121 3500 2125
rect 3502 2121 3503 2125
rect 3515 2121 3516 2125
rect 3518 2121 3519 2125
rect 3531 2121 3532 2125
rect 3534 2121 3537 2125
rect 3539 2121 3540 2125
rect 3557 2121 3558 2125
rect 3560 2121 3561 2125
rect 3573 2121 3574 2125
rect 3576 2121 3577 2125
rect 3589 2121 3590 2125
rect 3592 2121 3595 2125
rect 3597 2121 3598 2125
rect 3610 2121 3611 2125
rect 3613 2121 3614 2125
<< pdiffusion >>
rect 2769 4029 2770 4037
rect 2772 4029 2775 4037
rect 2777 4029 2778 4037
rect 2790 4029 2791 4037
rect 2793 4033 2794 4037
rect 2793 4029 2798 4033
rect 2806 4029 2807 4037
rect 2809 4029 2812 4037
rect 2814 4029 2815 4037
rect 2832 4029 2833 4037
rect 2835 4029 2836 4037
rect 2848 4029 2849 4037
rect 2851 4033 2852 4037
rect 2851 4029 2856 4033
rect 2864 4029 2865 4037
rect 2867 4029 2870 4037
rect 2872 4029 2873 4037
rect 2885 4029 2886 4037
rect 2888 4029 2889 4037
rect 2901 4029 2902 4037
rect 2904 4029 2907 4037
rect 2909 4029 2910 4037
rect 2922 4029 2923 4037
rect 2925 4033 2926 4037
rect 2925 4029 2930 4033
rect 2938 4029 2939 4037
rect 2941 4029 2944 4037
rect 2946 4029 2947 4037
rect 2964 4029 2965 4037
rect 2967 4029 2968 4037
rect 2980 4029 2981 4037
rect 2983 4033 2984 4037
rect 2983 4029 2988 4033
rect 2996 4029 2997 4037
rect 2999 4029 3002 4037
rect 3004 4029 3005 4037
rect 3017 4029 3018 4037
rect 3020 4029 3021 4037
rect 3033 4029 3034 4037
rect 3036 4029 3039 4037
rect 3041 4029 3042 4037
rect 3054 4029 3055 4037
rect 3057 4033 3058 4037
rect 3057 4029 3062 4033
rect 3070 4029 3071 4037
rect 3073 4029 3076 4037
rect 3078 4029 3079 4037
rect 3096 4029 3097 4037
rect 3099 4029 3100 4037
rect 3112 4029 3113 4037
rect 3115 4033 3116 4037
rect 3115 4029 3120 4033
rect 3128 4029 3129 4037
rect 3131 4029 3134 4037
rect 3136 4029 3137 4037
rect 3149 4029 3150 4037
rect 3152 4029 3153 4037
rect 3165 4029 3166 4037
rect 3168 4029 3171 4037
rect 3173 4029 3174 4037
rect 3186 4029 3187 4037
rect 3189 4033 3190 4037
rect 3189 4029 3194 4033
rect 3202 4029 3203 4037
rect 3205 4029 3208 4037
rect 3210 4029 3211 4037
rect 3228 4029 3229 4037
rect 3231 4029 3232 4037
rect 3244 4029 3245 4037
rect 3247 4033 3248 4037
rect 3247 4029 3252 4033
rect 3260 4029 3261 4037
rect 3263 4029 3266 4037
rect 3268 4029 3269 4037
rect 3281 4029 3282 4037
rect 3284 4029 3285 4037
rect 3714 4029 3715 4037
rect 3717 4029 3720 4037
rect 3722 4029 3723 4037
rect 3735 4029 3736 4037
rect 3738 4033 3739 4037
rect 3738 4029 3743 4033
rect 3751 4029 3752 4037
rect 3754 4029 3757 4037
rect 3759 4029 3760 4037
rect 3777 4029 3778 4037
rect 3780 4029 3781 4037
rect 3793 4029 3794 4037
rect 3796 4033 3797 4037
rect 3796 4029 3801 4033
rect 3809 4029 3810 4037
rect 3812 4029 3815 4037
rect 3817 4029 3818 4037
rect 3830 4029 3831 4037
rect 3833 4029 3834 4037
rect 3846 4029 3847 4037
rect 3849 4029 3852 4037
rect 3854 4029 3855 4037
rect 3867 4029 3868 4037
rect 3870 4033 3871 4037
rect 3870 4029 3875 4033
rect 3883 4029 3884 4037
rect 3886 4029 3889 4037
rect 3891 4029 3892 4037
rect 3909 4029 3910 4037
rect 3912 4029 3913 4037
rect 3925 4029 3926 4037
rect 3928 4033 3929 4037
rect 3928 4029 3933 4033
rect 3941 4029 3942 4037
rect 3944 4029 3947 4037
rect 3949 4029 3950 4037
rect 3962 4029 3963 4037
rect 3965 4029 3966 4037
rect 3978 4029 3979 4037
rect 3981 4029 3984 4037
rect 3986 4029 3987 4037
rect 3999 4029 4000 4037
rect 4002 4033 4003 4037
rect 4002 4029 4007 4033
rect 4015 4029 4016 4037
rect 4018 4029 4021 4037
rect 4023 4029 4024 4037
rect 4041 4029 4042 4037
rect 4044 4029 4045 4037
rect 4057 4029 4058 4037
rect 4060 4033 4061 4037
rect 4060 4029 4065 4033
rect 4073 4029 4074 4037
rect 4076 4029 4079 4037
rect 4081 4029 4082 4037
rect 4094 4029 4095 4037
rect 4097 4029 4098 4037
rect 4110 4029 4111 4037
rect 4113 4029 4116 4037
rect 4118 4029 4119 4037
rect 4131 4029 4132 4037
rect 4134 4033 4135 4037
rect 4134 4029 4139 4033
rect 4147 4029 4148 4037
rect 4150 4029 4153 4037
rect 4155 4029 4156 4037
rect 4173 4029 4174 4037
rect 4176 4029 4177 4037
rect 4189 4029 4190 4037
rect 4192 4033 4193 4037
rect 4192 4029 4197 4033
rect 4205 4029 4206 4037
rect 4208 4029 4211 4037
rect 4213 4029 4214 4037
rect 4226 4029 4227 4037
rect 4229 4029 4230 4037
rect 2417 3996 2418 4004
rect 2420 3996 2423 4004
rect 2425 3996 2426 4004
rect 2438 3996 2439 4004
rect 2441 4000 2442 4004
rect 2441 3996 2446 4000
rect 2454 3996 2455 4004
rect 2457 3996 2460 4004
rect 2462 3996 2463 4004
rect 2480 3996 2481 4004
rect 2483 3996 2484 4004
rect 2496 3996 2497 4004
rect 2499 4000 2500 4004
rect 2499 3996 2504 4000
rect 2512 3996 2513 4004
rect 2515 3996 2518 4004
rect 2520 3996 2521 4004
rect 2533 3996 2534 4004
rect 2536 3996 2537 4004
rect 3362 3996 3363 4004
rect 3365 3996 3368 4004
rect 3370 3996 3371 4004
rect 3383 3996 3384 4004
rect 3386 4000 3387 4004
rect 3386 3996 3391 4000
rect 3399 3996 3400 4004
rect 3402 3996 3405 4004
rect 3407 3996 3408 4004
rect 3425 3996 3426 4004
rect 3428 3996 3429 4004
rect 3441 3996 3442 4004
rect 3444 4000 3445 4004
rect 3444 3996 3449 4000
rect 3457 3996 3458 4004
rect 3460 3996 3463 4004
rect 3465 3996 3466 4004
rect 3478 3996 3479 4004
rect 3481 3996 3482 4004
rect 2948 3958 2949 3966
rect 2951 3958 2952 3966
rect 2774 3945 2775 3953
rect 2777 3945 2778 3953
rect 2790 3945 2791 3953
rect 2793 3945 2794 3953
rect 2806 3945 2807 3953
rect 2809 3945 2810 3953
rect 2825 3945 2830 3953
rect 2832 3945 2835 3953
rect 2837 3945 2838 3953
rect 2859 3945 2861 3953
rect 2863 3945 2864 3953
rect 2881 3945 2882 3953
rect 2884 3945 2885 3953
rect 2897 3945 2902 3953
rect 2904 3945 2907 3953
rect 2909 3945 2910 3953
rect 2924 3945 2925 3953
rect 2927 3945 2928 3953
rect 2972 3952 2975 3960
rect 2977 3952 2980 3960
rect 2982 3952 2983 3960
rect 3002 3958 3003 3966
rect 3005 3958 3006 3966
rect 3029 3958 3030 3966
rect 3032 3958 3033 3966
rect 3053 3952 3056 3960
rect 3058 3952 3061 3960
rect 3063 3952 3064 3960
rect 3083 3958 3084 3966
rect 3086 3958 3087 3966
rect 3893 3958 3894 3966
rect 3896 3958 3897 3966
rect 3719 3945 3720 3953
rect 3722 3945 3723 3953
rect 3735 3945 3736 3953
rect 3738 3945 3739 3953
rect 3751 3945 3752 3953
rect 3754 3945 3755 3953
rect 3770 3945 3775 3953
rect 3777 3945 3780 3953
rect 3782 3945 3783 3953
rect 3804 3945 3806 3953
rect 3808 3945 3809 3953
rect 3826 3945 3827 3953
rect 3829 3945 3830 3953
rect 3842 3945 3847 3953
rect 3849 3945 3852 3953
rect 3854 3945 3855 3953
rect 3869 3945 3870 3953
rect 3872 3945 3873 3953
rect 3917 3952 3920 3960
rect 3922 3952 3925 3960
rect 3927 3952 3928 3960
rect 3947 3958 3948 3966
rect 3950 3958 3951 3966
rect 3974 3958 3975 3966
rect 3977 3958 3978 3966
rect 3998 3952 4001 3960
rect 4003 3952 4006 3960
rect 4008 3952 4009 3960
rect 4028 3958 4029 3966
rect 4031 3958 4032 3966
rect 2408 3894 2409 3902
rect 2411 3894 2412 3902
rect 2424 3894 2425 3902
rect 2427 3894 2430 3902
rect 2432 3894 2433 3902
rect 2445 3898 2446 3902
rect 2441 3894 2446 3898
rect 2448 3894 2449 3902
rect 2461 3894 2462 3902
rect 2464 3894 2465 3902
rect 2482 3894 2483 3902
rect 2485 3894 2488 3902
rect 2490 3894 2491 3902
rect 2503 3898 2504 3902
rect 2499 3894 2504 3898
rect 2506 3894 2507 3902
rect 2519 3894 2520 3902
rect 2522 3894 2525 3902
rect 2527 3894 2528 3902
rect 3353 3894 3354 3902
rect 3356 3894 3357 3902
rect 3369 3894 3370 3902
rect 3372 3894 3375 3902
rect 3377 3894 3378 3902
rect 3390 3898 3391 3902
rect 3386 3894 3391 3898
rect 3393 3894 3394 3902
rect 3406 3894 3407 3902
rect 3409 3894 3410 3902
rect 3427 3894 3428 3902
rect 3430 3894 3433 3902
rect 3435 3894 3436 3902
rect 3448 3898 3449 3902
rect 3444 3894 3449 3898
rect 3451 3894 3452 3902
rect 3464 3894 3465 3902
rect 3467 3894 3470 3902
rect 3472 3894 3473 3902
rect 2774 3859 2775 3867
rect 2777 3859 2778 3867
rect 2790 3859 2791 3867
rect 2793 3859 2794 3867
rect 2806 3859 2807 3867
rect 2809 3859 2810 3867
rect 2825 3859 2830 3867
rect 2832 3859 2835 3867
rect 2837 3859 2838 3867
rect 2859 3859 2861 3867
rect 2863 3859 2864 3867
rect 2881 3859 2882 3867
rect 2884 3859 2885 3867
rect 2897 3859 2902 3867
rect 2904 3859 2907 3867
rect 2909 3859 2910 3867
rect 2924 3859 2925 3867
rect 2927 3859 2928 3867
rect 2972 3860 2975 3868
rect 2977 3860 2980 3868
rect 2982 3860 2983 3868
rect 3053 3860 3056 3868
rect 3058 3860 3061 3868
rect 3063 3860 3064 3868
rect 3719 3859 3720 3867
rect 3722 3859 3723 3867
rect 3735 3859 3736 3867
rect 3738 3859 3739 3867
rect 3751 3859 3752 3867
rect 3754 3859 3755 3867
rect 3770 3859 3775 3867
rect 3777 3859 3780 3867
rect 3782 3859 3783 3867
rect 3804 3859 3806 3867
rect 3808 3859 3809 3867
rect 3826 3859 3827 3867
rect 3829 3859 3830 3867
rect 3842 3859 3847 3867
rect 3849 3859 3852 3867
rect 3854 3859 3855 3867
rect 3869 3859 3870 3867
rect 3872 3859 3873 3867
rect 3917 3860 3920 3868
rect 3922 3860 3925 3868
rect 3927 3860 3928 3868
rect 3998 3860 4001 3868
rect 4003 3860 4006 3868
rect 4008 3860 4009 3868
rect 2774 3813 2775 3821
rect 2777 3813 2778 3821
rect 2790 3813 2791 3821
rect 2793 3813 2794 3821
rect 2806 3813 2807 3821
rect 2809 3813 2810 3821
rect 2825 3813 2830 3821
rect 2832 3813 2835 3821
rect 2837 3813 2838 3821
rect 2859 3813 2861 3821
rect 2863 3813 2864 3821
rect 2881 3813 2882 3821
rect 2884 3813 2885 3821
rect 2897 3813 2902 3821
rect 2904 3813 2907 3821
rect 2909 3813 2910 3821
rect 2924 3813 2925 3821
rect 2927 3813 2928 3821
rect 2972 3820 2975 3828
rect 2977 3820 2980 3828
rect 2982 3820 2983 3828
rect 3002 3826 3003 3834
rect 3005 3826 3006 3834
rect 3053 3826 3054 3834
rect 3056 3826 3057 3834
rect 3077 3820 3080 3828
rect 3082 3820 3085 3828
rect 3087 3820 3088 3828
rect 3107 3826 3108 3834
rect 3110 3826 3111 3834
rect 3719 3813 3720 3821
rect 3722 3813 3723 3821
rect 3735 3813 3736 3821
rect 3738 3813 3739 3821
rect 3751 3813 3752 3821
rect 3754 3813 3755 3821
rect 3770 3813 3775 3821
rect 3777 3813 3780 3821
rect 3782 3813 3783 3821
rect 3804 3813 3806 3821
rect 3808 3813 3809 3821
rect 3826 3813 3827 3821
rect 3829 3813 3830 3821
rect 3842 3813 3847 3821
rect 3849 3813 3852 3821
rect 3854 3813 3855 3821
rect 3869 3813 3870 3821
rect 3872 3813 3873 3821
rect 3917 3820 3920 3828
rect 3922 3820 3925 3828
rect 3927 3820 3928 3828
rect 3947 3826 3948 3834
rect 3950 3826 3951 3834
rect 3998 3826 3999 3834
rect 4001 3826 4002 3834
rect 3284 3797 3285 3805
rect 3287 3797 3288 3805
rect 3308 3791 3311 3799
rect 3313 3791 3316 3799
rect 3318 3791 3319 3799
rect 3338 3797 3339 3805
rect 3341 3797 3342 3805
rect 3470 3772 3471 3802
rect 3473 3772 3474 3802
rect 3523 3772 3524 3802
rect 3526 3772 3527 3802
rect 4022 3820 4025 3828
rect 4027 3820 4030 3828
rect 4032 3820 4033 3828
rect 4052 3826 4053 3834
rect 4055 3826 4056 3834
rect 2774 3727 2775 3735
rect 2777 3727 2778 3735
rect 2790 3727 2791 3735
rect 2793 3727 2794 3735
rect 2806 3727 2807 3735
rect 2809 3727 2810 3735
rect 2825 3727 2830 3735
rect 2832 3727 2835 3735
rect 2837 3727 2838 3735
rect 2859 3727 2861 3735
rect 2863 3727 2864 3735
rect 2881 3727 2882 3735
rect 2884 3727 2885 3735
rect 2897 3727 2902 3735
rect 2904 3727 2907 3735
rect 2909 3727 2910 3735
rect 2924 3727 2925 3735
rect 2927 3727 2928 3735
rect 2972 3729 2975 3737
rect 2977 3729 2980 3737
rect 2982 3729 2983 3737
rect 3077 3729 3080 3737
rect 3082 3729 3085 3737
rect 3087 3729 3088 3737
rect 3719 3727 3720 3735
rect 3722 3727 3723 3735
rect 3735 3727 3736 3735
rect 3738 3727 3739 3735
rect 3751 3727 3752 3735
rect 3754 3727 3755 3735
rect 3770 3727 3775 3735
rect 3777 3727 3780 3735
rect 3782 3727 3783 3735
rect 3804 3727 3806 3735
rect 3808 3727 3809 3735
rect 3826 3727 3827 3735
rect 3829 3727 3830 3735
rect 3842 3727 3847 3735
rect 3849 3727 3852 3735
rect 3854 3727 3855 3735
rect 3869 3727 3870 3735
rect 3872 3727 3873 3735
rect 3917 3729 3920 3737
rect 3922 3729 3925 3737
rect 3927 3729 3928 3737
rect 4022 3729 4025 3737
rect 4027 3729 4030 3737
rect 4032 3729 4033 3737
rect 2774 3681 2775 3689
rect 2777 3681 2778 3689
rect 2790 3681 2791 3689
rect 2793 3681 2794 3689
rect 2806 3681 2807 3689
rect 2809 3681 2810 3689
rect 2825 3681 2830 3689
rect 2832 3681 2835 3689
rect 2837 3681 2838 3689
rect 2859 3681 2861 3689
rect 2863 3681 2864 3689
rect 2881 3681 2882 3689
rect 2884 3681 2885 3689
rect 2897 3681 2902 3689
rect 2904 3681 2907 3689
rect 2909 3681 2910 3689
rect 2924 3681 2925 3689
rect 2927 3681 2928 3689
rect 2972 3688 2975 3696
rect 2977 3688 2980 3696
rect 2982 3688 2983 3696
rect 3002 3694 3003 3702
rect 3005 3694 3006 3702
rect 3029 3694 3030 3702
rect 3032 3694 3033 3702
rect 3053 3688 3056 3696
rect 3058 3688 3061 3696
rect 3063 3688 3064 3696
rect 3083 3694 3084 3702
rect 3086 3694 3087 3702
rect 3119 3694 3120 3702
rect 3122 3694 3123 3702
rect 3143 3688 3146 3696
rect 3148 3688 3151 3696
rect 3153 3688 3154 3696
rect 3173 3694 3174 3702
rect 3176 3694 3177 3702
rect 3308 3695 3311 3703
rect 3313 3695 3316 3703
rect 3318 3695 3319 3703
rect 3719 3681 3720 3689
rect 3722 3681 3723 3689
rect 3735 3681 3736 3689
rect 3738 3681 3739 3689
rect 3751 3681 3752 3689
rect 3754 3681 3755 3689
rect 3770 3681 3775 3689
rect 3777 3681 3780 3689
rect 3782 3681 3783 3689
rect 3804 3681 3806 3689
rect 3808 3681 3809 3689
rect 3826 3681 3827 3689
rect 3829 3681 3830 3689
rect 3842 3681 3847 3689
rect 3849 3681 3852 3689
rect 3854 3681 3855 3689
rect 3869 3681 3870 3689
rect 3872 3681 3873 3689
rect 3917 3688 3920 3696
rect 3922 3688 3925 3696
rect 3927 3688 3928 3696
rect 3947 3694 3948 3702
rect 3950 3694 3951 3702
rect 3974 3694 3975 3702
rect 3977 3694 3978 3702
rect 3262 3667 3263 3675
rect 3265 3667 3266 3675
rect 3284 3667 3285 3675
rect 3287 3667 3288 3675
rect 3308 3661 3311 3669
rect 3313 3661 3316 3669
rect 3318 3661 3319 3669
rect 3338 3667 3339 3675
rect 3341 3667 3342 3675
rect 3376 3642 3377 3672
rect 3379 3642 3380 3672
rect 3429 3642 3430 3672
rect 3432 3642 3433 3672
rect 3998 3688 4001 3696
rect 4003 3688 4006 3696
rect 4008 3688 4009 3696
rect 4028 3694 4029 3702
rect 4031 3694 4032 3702
rect 4064 3694 4065 3702
rect 4067 3694 4068 3702
rect 4088 3688 4091 3696
rect 4093 3688 4096 3696
rect 4098 3688 4099 3696
rect 4118 3694 4119 3702
rect 4121 3694 4122 3702
rect 2774 3595 2775 3603
rect 2777 3595 2778 3603
rect 2790 3595 2791 3603
rect 2793 3595 2794 3603
rect 2806 3595 2807 3603
rect 2809 3595 2810 3603
rect 2825 3595 2830 3603
rect 2832 3595 2835 3603
rect 2837 3595 2838 3603
rect 2859 3595 2861 3603
rect 2863 3595 2864 3603
rect 2881 3595 2882 3603
rect 2884 3595 2885 3603
rect 2897 3595 2902 3603
rect 2904 3595 2907 3603
rect 2909 3595 2910 3603
rect 2924 3595 2925 3603
rect 2927 3595 2928 3603
rect 2972 3594 2975 3602
rect 2977 3594 2980 3602
rect 2982 3594 2983 3602
rect 3053 3594 3056 3602
rect 3058 3594 3061 3602
rect 3063 3594 3064 3602
rect 3143 3594 3146 3602
rect 3148 3594 3151 3602
rect 3153 3594 3154 3602
rect 3719 3595 3720 3603
rect 3722 3595 3723 3603
rect 3735 3595 3736 3603
rect 3738 3595 3739 3603
rect 3751 3595 3752 3603
rect 3754 3595 3755 3603
rect 3770 3595 3775 3603
rect 3777 3595 3780 3603
rect 3782 3595 3783 3603
rect 3804 3595 3806 3603
rect 3808 3595 3809 3603
rect 3826 3595 3827 3603
rect 3829 3595 3830 3603
rect 3842 3595 3847 3603
rect 3849 3595 3852 3603
rect 3854 3595 3855 3603
rect 3869 3595 3870 3603
rect 3872 3595 3873 3603
rect 3917 3594 3920 3602
rect 3922 3594 3925 3602
rect 3927 3594 3928 3602
rect 3998 3594 4001 3602
rect 4003 3594 4006 3602
rect 4008 3594 4009 3602
rect 4088 3594 4091 3602
rect 4093 3594 4096 3602
rect 4098 3594 4099 3602
rect 2774 3549 2775 3557
rect 2777 3549 2778 3557
rect 2790 3549 2791 3557
rect 2793 3549 2794 3557
rect 2806 3549 2807 3557
rect 2809 3549 2810 3557
rect 2825 3549 2830 3557
rect 2832 3549 2835 3557
rect 2837 3549 2838 3557
rect 2859 3549 2861 3557
rect 2863 3549 2864 3557
rect 2881 3549 2882 3557
rect 2884 3549 2885 3557
rect 2897 3549 2902 3557
rect 2904 3549 2907 3557
rect 2909 3549 2910 3557
rect 2924 3549 2925 3557
rect 2927 3549 2928 3557
rect 2972 3556 2975 3564
rect 2977 3556 2980 3564
rect 2982 3556 2983 3564
rect 3002 3562 3003 3570
rect 3005 3562 3006 3570
rect 3308 3565 3311 3573
rect 3313 3565 3316 3573
rect 3318 3565 3319 3573
rect 3719 3549 3720 3557
rect 3722 3549 3723 3557
rect 3735 3549 3736 3557
rect 3738 3549 3739 3557
rect 3751 3549 3752 3557
rect 3754 3549 3755 3557
rect 3770 3549 3775 3557
rect 3777 3549 3780 3557
rect 3782 3549 3783 3557
rect 3804 3549 3806 3557
rect 3808 3549 3809 3557
rect 3826 3549 3827 3557
rect 3829 3549 3830 3557
rect 3842 3549 3847 3557
rect 3849 3549 3852 3557
rect 3854 3549 3855 3557
rect 3869 3549 3870 3557
rect 3872 3549 3873 3557
rect 3917 3556 3920 3564
rect 3922 3556 3925 3564
rect 3927 3556 3928 3564
rect 3947 3562 3948 3570
rect 3950 3562 3951 3570
rect 2285 3494 2286 3502
rect 2288 3494 2291 3502
rect 2293 3494 2294 3502
rect 2306 3494 2307 3502
rect 2309 3498 2310 3502
rect 2309 3494 2314 3498
rect 2322 3494 2323 3502
rect 2325 3494 2328 3502
rect 2330 3494 2331 3502
rect 2348 3494 2349 3502
rect 2351 3494 2352 3502
rect 2364 3494 2365 3502
rect 2367 3498 2368 3502
rect 2367 3494 2372 3498
rect 2380 3494 2381 3502
rect 2383 3494 2386 3502
rect 2388 3494 2389 3502
rect 2401 3494 2402 3502
rect 2404 3494 2405 3502
rect 2417 3494 2418 3502
rect 2420 3494 2423 3502
rect 2425 3494 2426 3502
rect 2438 3494 2439 3502
rect 2441 3498 2442 3502
rect 2441 3494 2446 3498
rect 2454 3494 2455 3502
rect 2457 3494 2460 3502
rect 2462 3494 2463 3502
rect 2480 3494 2481 3502
rect 2483 3494 2484 3502
rect 2496 3494 2497 3502
rect 2499 3498 2500 3502
rect 2499 3494 2504 3498
rect 2512 3494 2513 3502
rect 2515 3494 2518 3502
rect 2520 3494 2521 3502
rect 2533 3494 2534 3502
rect 2536 3494 2537 3502
rect 2549 3494 2550 3502
rect 2552 3494 2555 3502
rect 2557 3494 2558 3502
rect 2570 3494 2571 3502
rect 2573 3498 2574 3502
rect 2573 3494 2578 3498
rect 2586 3494 2587 3502
rect 2589 3494 2592 3502
rect 2594 3494 2595 3502
rect 2612 3494 2613 3502
rect 2615 3494 2616 3502
rect 2628 3494 2629 3502
rect 2631 3498 2632 3502
rect 2631 3494 2636 3498
rect 2644 3494 2645 3502
rect 2647 3494 2650 3502
rect 2652 3494 2653 3502
rect 2665 3494 2666 3502
rect 2668 3494 2669 3502
rect 3230 3494 3231 3502
rect 3233 3494 3236 3502
rect 3238 3494 3239 3502
rect 3251 3494 3252 3502
rect 3254 3498 3255 3502
rect 3254 3494 3259 3498
rect 3267 3494 3268 3502
rect 3270 3494 3273 3502
rect 3275 3494 3276 3502
rect 3293 3494 3294 3502
rect 3296 3494 3297 3502
rect 3309 3494 3310 3502
rect 3312 3498 3313 3502
rect 3312 3494 3317 3498
rect 3325 3494 3326 3502
rect 3328 3494 3331 3502
rect 3333 3494 3334 3502
rect 3346 3494 3347 3502
rect 3349 3494 3350 3502
rect 3362 3494 3363 3502
rect 3365 3494 3368 3502
rect 3370 3494 3371 3502
rect 3383 3494 3384 3502
rect 3386 3498 3387 3502
rect 3386 3494 3391 3498
rect 3399 3494 3400 3502
rect 3402 3494 3405 3502
rect 3407 3494 3408 3502
rect 3425 3494 3426 3502
rect 3428 3494 3429 3502
rect 3441 3494 3442 3502
rect 3444 3498 3445 3502
rect 3444 3494 3449 3498
rect 3457 3494 3458 3502
rect 3460 3494 3463 3502
rect 3465 3494 3466 3502
rect 3478 3494 3479 3502
rect 3481 3494 3482 3502
rect 3494 3494 3495 3502
rect 3497 3494 3500 3502
rect 3502 3494 3503 3502
rect 3515 3494 3516 3502
rect 3518 3498 3519 3502
rect 3518 3494 3523 3498
rect 3531 3494 3532 3502
rect 3534 3494 3537 3502
rect 3539 3494 3540 3502
rect 3557 3494 3558 3502
rect 3560 3494 3561 3502
rect 3573 3494 3574 3502
rect 3576 3498 3577 3502
rect 3576 3494 3581 3498
rect 3589 3494 3590 3502
rect 3592 3494 3595 3502
rect 3597 3494 3598 3502
rect 3610 3494 3611 3502
rect 3613 3494 3614 3502
rect 2774 3463 2775 3471
rect 2777 3463 2778 3471
rect 2790 3463 2791 3471
rect 2793 3463 2794 3471
rect 2806 3463 2807 3471
rect 2809 3463 2810 3471
rect 2825 3463 2830 3471
rect 2832 3463 2835 3471
rect 2837 3463 2838 3471
rect 2859 3463 2861 3471
rect 2863 3463 2864 3471
rect 2881 3463 2882 3471
rect 2884 3463 2885 3471
rect 2897 3463 2902 3471
rect 2904 3463 2907 3471
rect 2909 3463 2910 3471
rect 2924 3463 2925 3471
rect 2927 3463 2928 3471
rect 2972 3458 2975 3466
rect 2977 3458 2980 3466
rect 2982 3458 2983 3466
rect 3008 3463 3009 3471
rect 3011 3463 3012 3471
rect 3016 3463 3022 3471
rect 3026 3463 3027 3471
rect 3029 3463 3030 3471
rect 3051 3463 3052 3471
rect 3054 3463 3055 3471
rect 3067 3463 3068 3471
rect 3070 3463 3071 3471
rect 3086 3463 3091 3471
rect 3093 3463 3096 3471
rect 3098 3463 3099 3471
rect 3120 3463 3122 3471
rect 3124 3463 3125 3471
rect 3142 3463 3143 3471
rect 3145 3463 3146 3471
rect 3158 3463 3163 3471
rect 3165 3463 3168 3471
rect 3170 3463 3171 3471
rect 3185 3463 3186 3471
rect 3188 3463 3189 3471
rect 3719 3463 3720 3471
rect 3722 3463 3723 3471
rect 3735 3463 3736 3471
rect 3738 3463 3739 3471
rect 3751 3463 3752 3471
rect 3754 3463 3755 3471
rect 3770 3463 3775 3471
rect 3777 3463 3780 3471
rect 3782 3463 3783 3471
rect 3804 3463 3806 3471
rect 3808 3463 3809 3471
rect 3826 3463 3827 3471
rect 3829 3463 3830 3471
rect 3842 3463 3847 3471
rect 3849 3463 3852 3471
rect 3854 3463 3855 3471
rect 3869 3463 3870 3471
rect 3872 3463 3873 3471
rect 3917 3458 3920 3466
rect 3922 3458 3925 3466
rect 3927 3458 3928 3466
rect 3953 3463 3954 3471
rect 3956 3463 3957 3471
rect 3961 3463 3967 3471
rect 3971 3463 3972 3471
rect 3974 3463 3975 3471
rect 3996 3463 3997 3471
rect 3999 3463 4000 3471
rect 4012 3463 4013 3471
rect 4015 3463 4016 3471
rect 4031 3463 4036 3471
rect 4038 3463 4041 3471
rect 4043 3463 4044 3471
rect 4065 3463 4067 3471
rect 4069 3463 4070 3471
rect 4087 3463 4088 3471
rect 4090 3463 4091 3471
rect 4103 3463 4108 3471
rect 4110 3463 4113 3471
rect 4115 3463 4116 3471
rect 4130 3463 4131 3471
rect 4133 3463 4134 3471
rect 3068 3382 3069 3390
rect 3071 3382 3074 3390
rect 3076 3382 3077 3390
rect 3089 3382 3090 3390
rect 3092 3386 3093 3390
rect 3092 3382 3097 3386
rect 3105 3382 3106 3390
rect 3108 3382 3111 3390
rect 3113 3382 3114 3390
rect 3131 3382 3132 3390
rect 3134 3382 3135 3390
rect 3147 3382 3148 3390
rect 3150 3386 3151 3390
rect 3150 3382 3155 3386
rect 3163 3382 3164 3390
rect 3166 3382 3169 3390
rect 3171 3382 3172 3390
rect 3184 3382 3185 3390
rect 3187 3382 3188 3390
rect 4013 3382 4014 3390
rect 4016 3382 4019 3390
rect 4021 3382 4022 3390
rect 4034 3382 4035 3390
rect 4037 3386 4038 3390
rect 4037 3382 4042 3386
rect 4050 3382 4051 3390
rect 4053 3382 4056 3390
rect 4058 3382 4059 3390
rect 4076 3382 4077 3390
rect 4079 3382 4080 3390
rect 4092 3382 4093 3390
rect 4095 3386 4096 3390
rect 4095 3382 4100 3386
rect 4108 3382 4109 3390
rect 4111 3382 4114 3390
rect 4116 3382 4117 3390
rect 4129 3382 4130 3390
rect 4132 3382 4133 3390
rect 2285 3352 2286 3360
rect 2288 3352 2291 3360
rect 2293 3352 2294 3360
rect 2306 3352 2307 3360
rect 2309 3356 2310 3360
rect 2309 3352 2314 3356
rect 2322 3352 2323 3360
rect 2325 3352 2328 3360
rect 2330 3352 2331 3360
rect 2348 3352 2349 3360
rect 2351 3352 2352 3360
rect 2364 3352 2365 3360
rect 2367 3356 2368 3360
rect 2367 3352 2372 3356
rect 2380 3352 2381 3360
rect 2383 3352 2386 3360
rect 2388 3352 2389 3360
rect 2401 3352 2402 3360
rect 2404 3352 2405 3360
rect 2417 3352 2418 3360
rect 2420 3352 2423 3360
rect 2425 3352 2426 3360
rect 2438 3352 2439 3360
rect 2441 3356 2442 3360
rect 2441 3352 2446 3356
rect 2454 3352 2455 3360
rect 2457 3352 2460 3360
rect 2462 3352 2463 3360
rect 2480 3352 2481 3360
rect 2483 3352 2484 3360
rect 2496 3352 2497 3360
rect 2499 3356 2500 3360
rect 2499 3352 2504 3356
rect 2512 3352 2513 3360
rect 2515 3352 2518 3360
rect 2520 3352 2521 3360
rect 2533 3352 2534 3360
rect 2536 3352 2537 3360
rect 2549 3352 2550 3360
rect 2552 3352 2555 3360
rect 2557 3352 2558 3360
rect 2570 3352 2571 3360
rect 2573 3356 2574 3360
rect 2573 3352 2578 3356
rect 2586 3352 2587 3360
rect 2589 3352 2592 3360
rect 2594 3352 2595 3360
rect 2612 3352 2613 3360
rect 2615 3352 2616 3360
rect 2628 3352 2629 3360
rect 2631 3356 2632 3360
rect 2631 3352 2636 3356
rect 2644 3352 2645 3360
rect 2647 3352 2650 3360
rect 2652 3352 2653 3360
rect 2665 3352 2666 3360
rect 2668 3352 2669 3360
rect 3230 3352 3231 3360
rect 3233 3352 3236 3360
rect 3238 3352 3239 3360
rect 3251 3352 3252 3360
rect 3254 3356 3255 3360
rect 3254 3352 3259 3356
rect 3267 3352 3268 3360
rect 3270 3352 3273 3360
rect 3275 3352 3276 3360
rect 3293 3352 3294 3360
rect 3296 3352 3297 3360
rect 3309 3352 3310 3360
rect 3312 3356 3313 3360
rect 3312 3352 3317 3356
rect 3325 3352 3326 3360
rect 3328 3352 3331 3360
rect 3333 3352 3334 3360
rect 3346 3352 3347 3360
rect 3349 3352 3350 3360
rect 3362 3352 3363 3360
rect 3365 3352 3368 3360
rect 3370 3352 3371 3360
rect 3383 3352 3384 3360
rect 3386 3356 3387 3360
rect 3386 3352 3391 3356
rect 3399 3352 3400 3360
rect 3402 3352 3405 3360
rect 3407 3352 3408 3360
rect 3425 3352 3426 3360
rect 3428 3352 3429 3360
rect 3441 3352 3442 3360
rect 3444 3356 3445 3360
rect 3444 3352 3449 3356
rect 3457 3352 3458 3360
rect 3460 3352 3463 3360
rect 3465 3352 3466 3360
rect 3478 3352 3479 3360
rect 3481 3352 3482 3360
rect 3494 3352 3495 3360
rect 3497 3352 3500 3360
rect 3502 3352 3503 3360
rect 3515 3352 3516 3360
rect 3518 3356 3519 3360
rect 3518 3352 3523 3356
rect 3531 3352 3532 3360
rect 3534 3352 3537 3360
rect 3539 3352 3540 3360
rect 3557 3352 3558 3360
rect 3560 3352 3561 3360
rect 3573 3352 3574 3360
rect 3576 3356 3577 3360
rect 3576 3352 3581 3356
rect 3589 3352 3590 3360
rect 3592 3352 3595 3360
rect 3597 3352 3598 3360
rect 3610 3352 3611 3360
rect 3613 3352 3614 3360
rect 3068 3296 3069 3304
rect 3071 3296 3074 3304
rect 3076 3296 3077 3304
rect 3089 3296 3090 3304
rect 3092 3300 3093 3304
rect 3092 3296 3097 3300
rect 3105 3296 3106 3304
rect 3108 3296 3111 3304
rect 3113 3296 3114 3304
rect 3131 3296 3132 3304
rect 3134 3296 3135 3304
rect 3147 3296 3148 3304
rect 3150 3300 3151 3304
rect 3150 3296 3155 3300
rect 3163 3296 3164 3304
rect 3166 3296 3169 3304
rect 3171 3296 3172 3304
rect 3184 3296 3185 3304
rect 3187 3296 3188 3304
rect 4013 3296 4014 3304
rect 4016 3296 4019 3304
rect 4021 3296 4022 3304
rect 4034 3296 4035 3304
rect 4037 3300 4038 3304
rect 4037 3296 4042 3300
rect 4050 3296 4051 3304
rect 4053 3296 4056 3304
rect 4058 3296 4059 3304
rect 4076 3296 4077 3304
rect 4079 3296 4080 3304
rect 4092 3296 4093 3304
rect 4095 3300 4096 3304
rect 4095 3296 4100 3300
rect 4108 3296 4109 3304
rect 4111 3296 4114 3304
rect 4116 3296 4117 3304
rect 4129 3296 4130 3304
rect 4132 3296 4133 3304
rect 2285 3266 2286 3274
rect 2288 3266 2291 3274
rect 2293 3266 2294 3274
rect 2306 3266 2307 3274
rect 2309 3270 2310 3274
rect 2309 3266 2314 3270
rect 2322 3266 2323 3274
rect 2325 3266 2328 3274
rect 2330 3266 2331 3274
rect 2348 3266 2349 3274
rect 2351 3266 2352 3274
rect 2364 3266 2365 3274
rect 2367 3270 2368 3274
rect 2367 3266 2372 3270
rect 2380 3266 2381 3274
rect 2383 3266 2386 3274
rect 2388 3266 2389 3274
rect 2401 3266 2402 3274
rect 2404 3266 2405 3274
rect 2417 3266 2418 3274
rect 2420 3266 2423 3274
rect 2425 3266 2426 3274
rect 2438 3266 2439 3274
rect 2441 3270 2442 3274
rect 2441 3266 2446 3270
rect 2454 3266 2455 3274
rect 2457 3266 2460 3274
rect 2462 3266 2463 3274
rect 2480 3266 2481 3274
rect 2483 3266 2484 3274
rect 2496 3266 2497 3274
rect 2499 3270 2500 3274
rect 2499 3266 2504 3270
rect 2512 3266 2513 3274
rect 2515 3266 2518 3274
rect 2520 3266 2521 3274
rect 2533 3266 2534 3274
rect 2536 3266 2537 3274
rect 2549 3266 2550 3274
rect 2552 3266 2555 3274
rect 2557 3266 2558 3274
rect 2570 3266 2571 3274
rect 2573 3270 2574 3274
rect 2573 3266 2578 3270
rect 2586 3266 2587 3274
rect 2589 3266 2592 3274
rect 2594 3266 2595 3274
rect 2612 3266 2613 3274
rect 2615 3266 2616 3274
rect 2628 3266 2629 3274
rect 2631 3270 2632 3274
rect 2631 3266 2636 3270
rect 2644 3266 2645 3274
rect 2647 3266 2650 3274
rect 2652 3266 2653 3274
rect 2665 3266 2666 3274
rect 2668 3266 2669 3274
rect 3230 3266 3231 3274
rect 3233 3266 3236 3274
rect 3238 3266 3239 3274
rect 3251 3266 3252 3274
rect 3254 3270 3255 3274
rect 3254 3266 3259 3270
rect 3267 3266 3268 3274
rect 3270 3266 3273 3274
rect 3275 3266 3276 3274
rect 3293 3266 3294 3274
rect 3296 3266 3297 3274
rect 3309 3266 3310 3274
rect 3312 3270 3313 3274
rect 3312 3266 3317 3270
rect 3325 3266 3326 3274
rect 3328 3266 3331 3274
rect 3333 3266 3334 3274
rect 3346 3266 3347 3274
rect 3349 3266 3350 3274
rect 3362 3266 3363 3274
rect 3365 3266 3368 3274
rect 3370 3266 3371 3274
rect 3383 3266 3384 3274
rect 3386 3270 3387 3274
rect 3386 3266 3391 3270
rect 3399 3266 3400 3274
rect 3402 3266 3405 3274
rect 3407 3266 3408 3274
rect 3425 3266 3426 3274
rect 3428 3266 3429 3274
rect 3441 3266 3442 3274
rect 3444 3270 3445 3274
rect 3444 3266 3449 3270
rect 3457 3266 3458 3274
rect 3460 3266 3463 3274
rect 3465 3266 3466 3274
rect 3478 3266 3479 3274
rect 3481 3266 3482 3274
rect 3494 3266 3495 3274
rect 3497 3266 3500 3274
rect 3502 3266 3503 3274
rect 3515 3266 3516 3274
rect 3518 3270 3519 3274
rect 3518 3266 3523 3270
rect 3531 3266 3532 3274
rect 3534 3266 3537 3274
rect 3539 3266 3540 3274
rect 3557 3266 3558 3274
rect 3560 3266 3561 3274
rect 3573 3266 3574 3274
rect 3576 3270 3577 3274
rect 3576 3266 3581 3270
rect 3589 3266 3590 3274
rect 3592 3266 3595 3274
rect 3597 3266 3598 3274
rect 3610 3266 3611 3274
rect 3613 3266 3614 3274
rect 2285 3126 2286 3134
rect 2288 3126 2291 3134
rect 2293 3126 2294 3134
rect 2306 3126 2307 3134
rect 2309 3130 2310 3134
rect 2309 3126 2314 3130
rect 2322 3126 2323 3134
rect 2325 3126 2328 3134
rect 2330 3126 2331 3134
rect 2348 3126 2349 3134
rect 2351 3126 2352 3134
rect 2364 3126 2365 3134
rect 2367 3130 2368 3134
rect 2367 3126 2372 3130
rect 2380 3126 2381 3134
rect 2383 3126 2386 3134
rect 2388 3126 2389 3134
rect 2401 3126 2402 3134
rect 2404 3126 2405 3134
rect 2417 3126 2418 3134
rect 2420 3126 2423 3134
rect 2425 3126 2426 3134
rect 2438 3126 2439 3134
rect 2441 3130 2442 3134
rect 2441 3126 2446 3130
rect 2454 3126 2455 3134
rect 2457 3126 2460 3134
rect 2462 3126 2463 3134
rect 2480 3126 2481 3134
rect 2483 3126 2484 3134
rect 2496 3126 2497 3134
rect 2499 3130 2500 3134
rect 2499 3126 2504 3130
rect 2512 3126 2513 3134
rect 2515 3126 2518 3134
rect 2520 3126 2521 3134
rect 2533 3126 2534 3134
rect 2536 3126 2537 3134
rect 2549 3126 2550 3134
rect 2552 3126 2555 3134
rect 2557 3126 2558 3134
rect 2570 3126 2571 3134
rect 2573 3130 2574 3134
rect 2573 3126 2578 3130
rect 2586 3126 2587 3134
rect 2589 3126 2592 3134
rect 2594 3126 2595 3134
rect 2612 3126 2613 3134
rect 2615 3126 2616 3134
rect 2628 3126 2629 3134
rect 2631 3130 2632 3134
rect 2631 3126 2636 3130
rect 2644 3126 2645 3134
rect 2647 3126 2650 3134
rect 2652 3126 2653 3134
rect 2665 3126 2666 3134
rect 2668 3126 2669 3134
rect 3230 3126 3231 3134
rect 3233 3126 3236 3134
rect 3238 3126 3239 3134
rect 3251 3126 3252 3134
rect 3254 3130 3255 3134
rect 3254 3126 3259 3130
rect 3267 3126 3268 3134
rect 3270 3126 3273 3134
rect 3275 3126 3276 3134
rect 3293 3126 3294 3134
rect 3296 3126 3297 3134
rect 3309 3126 3310 3134
rect 3312 3130 3313 3134
rect 3312 3126 3317 3130
rect 3325 3126 3326 3134
rect 3328 3126 3331 3134
rect 3333 3126 3334 3134
rect 3346 3126 3347 3134
rect 3349 3126 3350 3134
rect 3362 3126 3363 3134
rect 3365 3126 3368 3134
rect 3370 3126 3371 3134
rect 3383 3126 3384 3134
rect 3386 3130 3387 3134
rect 3386 3126 3391 3130
rect 3399 3126 3400 3134
rect 3402 3126 3405 3134
rect 3407 3126 3408 3134
rect 3425 3126 3426 3134
rect 3428 3126 3429 3134
rect 3441 3126 3442 3134
rect 3444 3130 3445 3134
rect 3444 3126 3449 3130
rect 3457 3126 3458 3134
rect 3460 3126 3463 3134
rect 3465 3126 3466 3134
rect 3478 3126 3479 3134
rect 3481 3126 3482 3134
rect 3494 3126 3495 3134
rect 3497 3126 3500 3134
rect 3502 3126 3503 3134
rect 3515 3126 3516 3134
rect 3518 3130 3519 3134
rect 3518 3126 3523 3130
rect 3531 3126 3532 3134
rect 3534 3126 3537 3134
rect 3539 3126 3540 3134
rect 3557 3126 3558 3134
rect 3560 3126 3561 3134
rect 3573 3126 3574 3134
rect 3576 3130 3577 3134
rect 3576 3126 3581 3130
rect 3589 3126 3590 3134
rect 3592 3126 3595 3134
rect 3597 3126 3598 3134
rect 3610 3126 3611 3134
rect 3613 3126 3614 3134
rect 2769 3047 2770 3055
rect 2772 3047 2775 3055
rect 2777 3047 2778 3055
rect 2790 3047 2791 3055
rect 2793 3051 2794 3055
rect 2793 3047 2798 3051
rect 2806 3047 2807 3055
rect 2809 3047 2812 3055
rect 2814 3047 2815 3055
rect 2832 3047 2833 3055
rect 2835 3047 2836 3055
rect 2848 3047 2849 3055
rect 2851 3051 2852 3055
rect 2851 3047 2856 3051
rect 2864 3047 2865 3055
rect 2867 3047 2870 3055
rect 2872 3047 2873 3055
rect 2885 3047 2886 3055
rect 2888 3047 2889 3055
rect 2901 3047 2902 3055
rect 2904 3047 2907 3055
rect 2909 3047 2910 3055
rect 2922 3047 2923 3055
rect 2925 3051 2926 3055
rect 2925 3047 2930 3051
rect 2938 3047 2939 3055
rect 2941 3047 2944 3055
rect 2946 3047 2947 3055
rect 2964 3047 2965 3055
rect 2967 3047 2968 3055
rect 2980 3047 2981 3055
rect 2983 3051 2984 3055
rect 2983 3047 2988 3051
rect 2996 3047 2997 3055
rect 2999 3047 3002 3055
rect 3004 3047 3005 3055
rect 3017 3047 3018 3055
rect 3020 3047 3021 3055
rect 3033 3047 3034 3055
rect 3036 3047 3039 3055
rect 3041 3047 3042 3055
rect 3054 3047 3055 3055
rect 3057 3051 3058 3055
rect 3057 3047 3062 3051
rect 3070 3047 3071 3055
rect 3073 3047 3076 3055
rect 3078 3047 3079 3055
rect 3096 3047 3097 3055
rect 3099 3047 3100 3055
rect 3112 3047 3113 3055
rect 3115 3051 3116 3055
rect 3115 3047 3120 3051
rect 3128 3047 3129 3055
rect 3131 3047 3134 3055
rect 3136 3047 3137 3055
rect 3149 3047 3150 3055
rect 3152 3047 3153 3055
rect 3165 3047 3166 3055
rect 3168 3047 3171 3055
rect 3173 3047 3174 3055
rect 3186 3047 3187 3055
rect 3189 3051 3190 3055
rect 3189 3047 3194 3051
rect 3202 3047 3203 3055
rect 3205 3047 3208 3055
rect 3210 3047 3211 3055
rect 3228 3047 3229 3055
rect 3231 3047 3232 3055
rect 3244 3047 3245 3055
rect 3247 3051 3248 3055
rect 3247 3047 3252 3051
rect 3260 3047 3261 3055
rect 3263 3047 3266 3055
rect 3268 3047 3269 3055
rect 3281 3047 3282 3055
rect 3284 3047 3285 3055
rect 3714 3047 3715 3055
rect 3717 3047 3720 3055
rect 3722 3047 3723 3055
rect 3735 3047 3736 3055
rect 3738 3051 3739 3055
rect 3738 3047 3743 3051
rect 3751 3047 3752 3055
rect 3754 3047 3757 3055
rect 3759 3047 3760 3055
rect 3777 3047 3778 3055
rect 3780 3047 3781 3055
rect 3793 3047 3794 3055
rect 3796 3051 3797 3055
rect 3796 3047 3801 3051
rect 3809 3047 3810 3055
rect 3812 3047 3815 3055
rect 3817 3047 3818 3055
rect 3830 3047 3831 3055
rect 3833 3047 3834 3055
rect 3846 3047 3847 3055
rect 3849 3047 3852 3055
rect 3854 3047 3855 3055
rect 3867 3047 3868 3055
rect 3870 3051 3871 3055
rect 3870 3047 3875 3051
rect 3883 3047 3884 3055
rect 3886 3047 3889 3055
rect 3891 3047 3892 3055
rect 3909 3047 3910 3055
rect 3912 3047 3913 3055
rect 3925 3047 3926 3055
rect 3928 3051 3929 3055
rect 3928 3047 3933 3051
rect 3941 3047 3942 3055
rect 3944 3047 3947 3055
rect 3949 3047 3950 3055
rect 3962 3047 3963 3055
rect 3965 3047 3966 3055
rect 3978 3047 3979 3055
rect 3981 3047 3984 3055
rect 3986 3047 3987 3055
rect 3999 3047 4000 3055
rect 4002 3051 4003 3055
rect 4002 3047 4007 3051
rect 4015 3047 4016 3055
rect 4018 3047 4021 3055
rect 4023 3047 4024 3055
rect 4041 3047 4042 3055
rect 4044 3047 4045 3055
rect 4057 3047 4058 3055
rect 4060 3051 4061 3055
rect 4060 3047 4065 3051
rect 4073 3047 4074 3055
rect 4076 3047 4079 3055
rect 4081 3047 4082 3055
rect 4094 3047 4095 3055
rect 4097 3047 4098 3055
rect 4110 3047 4111 3055
rect 4113 3047 4116 3055
rect 4118 3047 4119 3055
rect 4131 3047 4132 3055
rect 4134 3051 4135 3055
rect 4134 3047 4139 3051
rect 4147 3047 4148 3055
rect 4150 3047 4153 3055
rect 4155 3047 4156 3055
rect 4173 3047 4174 3055
rect 4176 3047 4177 3055
rect 4189 3047 4190 3055
rect 4192 3051 4193 3055
rect 4192 3047 4197 3051
rect 4205 3047 4206 3055
rect 4208 3047 4211 3055
rect 4213 3047 4214 3055
rect 4226 3047 4227 3055
rect 4229 3047 4230 3055
rect 2417 3014 2418 3022
rect 2420 3014 2423 3022
rect 2425 3014 2426 3022
rect 2438 3014 2439 3022
rect 2441 3018 2442 3022
rect 2441 3014 2446 3018
rect 2454 3014 2455 3022
rect 2457 3014 2460 3022
rect 2462 3014 2463 3022
rect 2480 3014 2481 3022
rect 2483 3014 2484 3022
rect 2496 3014 2497 3022
rect 2499 3018 2500 3022
rect 2499 3014 2504 3018
rect 2512 3014 2513 3022
rect 2515 3014 2518 3022
rect 2520 3014 2521 3022
rect 2533 3014 2534 3022
rect 2536 3014 2537 3022
rect 3362 3014 3363 3022
rect 3365 3014 3368 3022
rect 3370 3014 3371 3022
rect 3383 3014 3384 3022
rect 3386 3018 3387 3022
rect 3386 3014 3391 3018
rect 3399 3014 3400 3022
rect 3402 3014 3405 3022
rect 3407 3014 3408 3022
rect 3425 3014 3426 3022
rect 3428 3014 3429 3022
rect 3441 3014 3442 3022
rect 3444 3018 3445 3022
rect 3444 3014 3449 3018
rect 3457 3014 3458 3022
rect 3460 3014 3463 3022
rect 3465 3014 3466 3022
rect 3478 3014 3479 3022
rect 3481 3014 3482 3022
rect 2948 2976 2949 2984
rect 2951 2976 2952 2984
rect 2774 2963 2775 2971
rect 2777 2963 2778 2971
rect 2790 2963 2791 2971
rect 2793 2963 2794 2971
rect 2806 2963 2807 2971
rect 2809 2963 2810 2971
rect 2825 2963 2830 2971
rect 2832 2963 2835 2971
rect 2837 2963 2838 2971
rect 2859 2963 2861 2971
rect 2863 2963 2864 2971
rect 2881 2963 2882 2971
rect 2884 2963 2885 2971
rect 2897 2963 2902 2971
rect 2904 2963 2907 2971
rect 2909 2963 2910 2971
rect 2924 2963 2925 2971
rect 2927 2963 2928 2971
rect 2972 2970 2975 2978
rect 2977 2970 2980 2978
rect 2982 2970 2983 2978
rect 3002 2976 3003 2984
rect 3005 2976 3006 2984
rect 3029 2976 3030 2984
rect 3032 2976 3033 2984
rect 3053 2970 3056 2978
rect 3058 2970 3061 2978
rect 3063 2970 3064 2978
rect 3083 2976 3084 2984
rect 3086 2976 3087 2984
rect 3893 2976 3894 2984
rect 3896 2976 3897 2984
rect 3719 2963 3720 2971
rect 3722 2963 3723 2971
rect 3735 2963 3736 2971
rect 3738 2963 3739 2971
rect 3751 2963 3752 2971
rect 3754 2963 3755 2971
rect 3770 2963 3775 2971
rect 3777 2963 3780 2971
rect 3782 2963 3783 2971
rect 3804 2963 3806 2971
rect 3808 2963 3809 2971
rect 3826 2963 3827 2971
rect 3829 2963 3830 2971
rect 3842 2963 3847 2971
rect 3849 2963 3852 2971
rect 3854 2963 3855 2971
rect 3869 2963 3870 2971
rect 3872 2963 3873 2971
rect 3917 2970 3920 2978
rect 3922 2970 3925 2978
rect 3927 2970 3928 2978
rect 3947 2976 3948 2984
rect 3950 2976 3951 2984
rect 3974 2976 3975 2984
rect 3977 2976 3978 2984
rect 3998 2970 4001 2978
rect 4003 2970 4006 2978
rect 4008 2970 4009 2978
rect 4028 2976 4029 2984
rect 4031 2976 4032 2984
rect 2408 2912 2409 2920
rect 2411 2912 2412 2920
rect 2424 2912 2425 2920
rect 2427 2912 2430 2920
rect 2432 2912 2433 2920
rect 2445 2916 2446 2920
rect 2441 2912 2446 2916
rect 2448 2912 2449 2920
rect 2461 2912 2462 2920
rect 2464 2912 2465 2920
rect 2482 2912 2483 2920
rect 2485 2912 2488 2920
rect 2490 2912 2491 2920
rect 2503 2916 2504 2920
rect 2499 2912 2504 2916
rect 2506 2912 2507 2920
rect 2519 2912 2520 2920
rect 2522 2912 2525 2920
rect 2527 2912 2528 2920
rect 3353 2912 3354 2920
rect 3356 2912 3357 2920
rect 3369 2912 3370 2920
rect 3372 2912 3375 2920
rect 3377 2912 3378 2920
rect 3390 2916 3391 2920
rect 3386 2912 3391 2916
rect 3393 2912 3394 2920
rect 3406 2912 3407 2920
rect 3409 2912 3410 2920
rect 3427 2912 3428 2920
rect 3430 2912 3433 2920
rect 3435 2912 3436 2920
rect 3448 2916 3449 2920
rect 3444 2912 3449 2916
rect 3451 2912 3452 2920
rect 3464 2912 3465 2920
rect 3467 2912 3470 2920
rect 3472 2912 3473 2920
rect 2774 2877 2775 2885
rect 2777 2877 2778 2885
rect 2790 2877 2791 2885
rect 2793 2877 2794 2885
rect 2806 2877 2807 2885
rect 2809 2877 2810 2885
rect 2825 2877 2830 2885
rect 2832 2877 2835 2885
rect 2837 2877 2838 2885
rect 2859 2877 2861 2885
rect 2863 2877 2864 2885
rect 2881 2877 2882 2885
rect 2884 2877 2885 2885
rect 2897 2877 2902 2885
rect 2904 2877 2907 2885
rect 2909 2877 2910 2885
rect 2924 2877 2925 2885
rect 2927 2877 2928 2885
rect 2972 2878 2975 2886
rect 2977 2878 2980 2886
rect 2982 2878 2983 2886
rect 3053 2878 3056 2886
rect 3058 2878 3061 2886
rect 3063 2878 3064 2886
rect 3719 2877 3720 2885
rect 3722 2877 3723 2885
rect 3735 2877 3736 2885
rect 3738 2877 3739 2885
rect 3751 2877 3752 2885
rect 3754 2877 3755 2885
rect 3770 2877 3775 2885
rect 3777 2877 3780 2885
rect 3782 2877 3783 2885
rect 3804 2877 3806 2885
rect 3808 2877 3809 2885
rect 3826 2877 3827 2885
rect 3829 2877 3830 2885
rect 3842 2877 3847 2885
rect 3849 2877 3852 2885
rect 3854 2877 3855 2885
rect 3869 2877 3870 2885
rect 3872 2877 3873 2885
rect 3917 2878 3920 2886
rect 3922 2878 3925 2886
rect 3927 2878 3928 2886
rect 3998 2878 4001 2886
rect 4003 2878 4006 2886
rect 4008 2878 4009 2886
rect 2774 2831 2775 2839
rect 2777 2831 2778 2839
rect 2790 2831 2791 2839
rect 2793 2831 2794 2839
rect 2806 2831 2807 2839
rect 2809 2831 2810 2839
rect 2825 2831 2830 2839
rect 2832 2831 2835 2839
rect 2837 2831 2838 2839
rect 2859 2831 2861 2839
rect 2863 2831 2864 2839
rect 2881 2831 2882 2839
rect 2884 2831 2885 2839
rect 2897 2831 2902 2839
rect 2904 2831 2907 2839
rect 2909 2831 2910 2839
rect 2924 2831 2925 2839
rect 2927 2831 2928 2839
rect 2972 2838 2975 2846
rect 2977 2838 2980 2846
rect 2982 2838 2983 2846
rect 3002 2844 3003 2852
rect 3005 2844 3006 2852
rect 3053 2844 3054 2852
rect 3056 2844 3057 2852
rect 3077 2838 3080 2846
rect 3082 2838 3085 2846
rect 3087 2838 3088 2846
rect 3107 2844 3108 2852
rect 3110 2844 3111 2852
rect 3719 2831 3720 2839
rect 3722 2831 3723 2839
rect 3735 2831 3736 2839
rect 3738 2831 3739 2839
rect 3751 2831 3752 2839
rect 3754 2831 3755 2839
rect 3770 2831 3775 2839
rect 3777 2831 3780 2839
rect 3782 2831 3783 2839
rect 3804 2831 3806 2839
rect 3808 2831 3809 2839
rect 3826 2831 3827 2839
rect 3829 2831 3830 2839
rect 3842 2831 3847 2839
rect 3849 2831 3852 2839
rect 3854 2831 3855 2839
rect 3869 2831 3870 2839
rect 3872 2831 3873 2839
rect 3917 2838 3920 2846
rect 3922 2838 3925 2846
rect 3927 2838 3928 2846
rect 3947 2844 3948 2852
rect 3950 2844 3951 2852
rect 3998 2844 3999 2852
rect 4001 2844 4002 2852
rect 4022 2838 4025 2846
rect 4027 2838 4030 2846
rect 4032 2838 4033 2846
rect 4052 2844 4053 2852
rect 4055 2844 4056 2852
rect 2774 2745 2775 2753
rect 2777 2745 2778 2753
rect 2790 2745 2791 2753
rect 2793 2745 2794 2753
rect 2806 2745 2807 2753
rect 2809 2745 2810 2753
rect 2825 2745 2830 2753
rect 2832 2745 2835 2753
rect 2837 2745 2838 2753
rect 2859 2745 2861 2753
rect 2863 2745 2864 2753
rect 2881 2745 2882 2753
rect 2884 2745 2885 2753
rect 2897 2745 2902 2753
rect 2904 2745 2907 2753
rect 2909 2745 2910 2753
rect 2924 2745 2925 2753
rect 2927 2745 2928 2753
rect 2972 2747 2975 2755
rect 2977 2747 2980 2755
rect 2982 2747 2983 2755
rect 3077 2747 3080 2755
rect 3082 2747 3085 2755
rect 3087 2747 3088 2755
rect 3719 2745 3720 2753
rect 3722 2745 3723 2753
rect 3735 2745 3736 2753
rect 3738 2745 3739 2753
rect 3751 2745 3752 2753
rect 3754 2745 3755 2753
rect 3770 2745 3775 2753
rect 3777 2745 3780 2753
rect 3782 2745 3783 2753
rect 3804 2745 3806 2753
rect 3808 2745 3809 2753
rect 3826 2745 3827 2753
rect 3829 2745 3830 2753
rect 3842 2745 3847 2753
rect 3849 2745 3852 2753
rect 3854 2745 3855 2753
rect 3869 2745 3870 2753
rect 3872 2745 3873 2753
rect 3917 2747 3920 2755
rect 3922 2747 3925 2755
rect 3927 2747 3928 2755
rect 4022 2747 4025 2755
rect 4027 2747 4030 2755
rect 4032 2747 4033 2755
rect 2774 2699 2775 2707
rect 2777 2699 2778 2707
rect 2790 2699 2791 2707
rect 2793 2699 2794 2707
rect 2806 2699 2807 2707
rect 2809 2699 2810 2707
rect 2825 2699 2830 2707
rect 2832 2699 2835 2707
rect 2837 2699 2838 2707
rect 2859 2699 2861 2707
rect 2863 2699 2864 2707
rect 2881 2699 2882 2707
rect 2884 2699 2885 2707
rect 2897 2699 2902 2707
rect 2904 2699 2907 2707
rect 2909 2699 2910 2707
rect 2924 2699 2925 2707
rect 2927 2699 2928 2707
rect 2972 2706 2975 2714
rect 2977 2706 2980 2714
rect 2982 2706 2983 2714
rect 3002 2712 3003 2720
rect 3005 2712 3006 2720
rect 3029 2712 3030 2720
rect 3032 2712 3033 2720
rect 3053 2706 3056 2714
rect 3058 2706 3061 2714
rect 3063 2706 3064 2714
rect 3083 2712 3084 2720
rect 3086 2712 3087 2720
rect 3119 2712 3120 2720
rect 3122 2712 3123 2720
rect 3143 2706 3146 2714
rect 3148 2706 3151 2714
rect 3153 2706 3154 2714
rect 3173 2712 3174 2720
rect 3176 2712 3177 2720
rect 3719 2699 3720 2707
rect 3722 2699 3723 2707
rect 3735 2699 3736 2707
rect 3738 2699 3739 2707
rect 3751 2699 3752 2707
rect 3754 2699 3755 2707
rect 3770 2699 3775 2707
rect 3777 2699 3780 2707
rect 3782 2699 3783 2707
rect 3804 2699 3806 2707
rect 3808 2699 3809 2707
rect 3826 2699 3827 2707
rect 3829 2699 3830 2707
rect 3842 2699 3847 2707
rect 3849 2699 3852 2707
rect 3854 2699 3855 2707
rect 3869 2699 3870 2707
rect 3872 2699 3873 2707
rect 3917 2706 3920 2714
rect 3922 2706 3925 2714
rect 3927 2706 3928 2714
rect 3947 2712 3948 2720
rect 3950 2712 3951 2720
rect 3974 2712 3975 2720
rect 3977 2712 3978 2720
rect 3998 2706 4001 2714
rect 4003 2706 4006 2714
rect 4008 2706 4009 2714
rect 4028 2712 4029 2720
rect 4031 2712 4032 2720
rect 4064 2712 4065 2720
rect 4067 2712 4068 2720
rect 4088 2706 4091 2714
rect 4093 2706 4096 2714
rect 4098 2706 4099 2714
rect 4118 2712 4119 2720
rect 4121 2712 4122 2720
rect 2774 2613 2775 2621
rect 2777 2613 2778 2621
rect 2790 2613 2791 2621
rect 2793 2613 2794 2621
rect 2806 2613 2807 2621
rect 2809 2613 2810 2621
rect 2825 2613 2830 2621
rect 2832 2613 2835 2621
rect 2837 2613 2838 2621
rect 2859 2613 2861 2621
rect 2863 2613 2864 2621
rect 2881 2613 2882 2621
rect 2884 2613 2885 2621
rect 2897 2613 2902 2621
rect 2904 2613 2907 2621
rect 2909 2613 2910 2621
rect 2924 2613 2925 2621
rect 2927 2613 2928 2621
rect 2972 2612 2975 2620
rect 2977 2612 2980 2620
rect 2982 2612 2983 2620
rect 3053 2612 3056 2620
rect 3058 2612 3061 2620
rect 3063 2612 3064 2620
rect 3143 2612 3146 2620
rect 3148 2612 3151 2620
rect 3153 2612 3154 2620
rect 3719 2613 3720 2621
rect 3722 2613 3723 2621
rect 3735 2613 3736 2621
rect 3738 2613 3739 2621
rect 3751 2613 3752 2621
rect 3754 2613 3755 2621
rect 3770 2613 3775 2621
rect 3777 2613 3780 2621
rect 3782 2613 3783 2621
rect 3804 2613 3806 2621
rect 3808 2613 3809 2621
rect 3826 2613 3827 2621
rect 3829 2613 3830 2621
rect 3842 2613 3847 2621
rect 3849 2613 3852 2621
rect 3854 2613 3855 2621
rect 3869 2613 3870 2621
rect 3872 2613 3873 2621
rect 3917 2612 3920 2620
rect 3922 2612 3925 2620
rect 3927 2612 3928 2620
rect 3998 2612 4001 2620
rect 4003 2612 4006 2620
rect 4008 2612 4009 2620
rect 4088 2612 4091 2620
rect 4093 2612 4096 2620
rect 4098 2612 4099 2620
rect 2774 2567 2775 2575
rect 2777 2567 2778 2575
rect 2790 2567 2791 2575
rect 2793 2567 2794 2575
rect 2806 2567 2807 2575
rect 2809 2567 2810 2575
rect 2825 2567 2830 2575
rect 2832 2567 2835 2575
rect 2837 2567 2838 2575
rect 2859 2567 2861 2575
rect 2863 2567 2864 2575
rect 2881 2567 2882 2575
rect 2884 2567 2885 2575
rect 2897 2567 2902 2575
rect 2904 2567 2907 2575
rect 2909 2567 2910 2575
rect 2924 2567 2925 2575
rect 2927 2567 2928 2575
rect 2972 2574 2975 2582
rect 2977 2574 2980 2582
rect 2982 2574 2983 2582
rect 3002 2580 3003 2588
rect 3005 2580 3006 2588
rect 3719 2567 3720 2575
rect 3722 2567 3723 2575
rect 3735 2567 3736 2575
rect 3738 2567 3739 2575
rect 3751 2567 3752 2575
rect 3754 2567 3755 2575
rect 3770 2567 3775 2575
rect 3777 2567 3780 2575
rect 3782 2567 3783 2575
rect 3804 2567 3806 2575
rect 3808 2567 3809 2575
rect 3826 2567 3827 2575
rect 3829 2567 3830 2575
rect 3842 2567 3847 2575
rect 3849 2567 3852 2575
rect 3854 2567 3855 2575
rect 3869 2567 3870 2575
rect 3872 2567 3873 2575
rect 3917 2574 3920 2582
rect 3922 2574 3925 2582
rect 3927 2574 3928 2582
rect 3947 2580 3948 2588
rect 3950 2580 3951 2588
rect 2285 2512 2286 2520
rect 2288 2512 2291 2520
rect 2293 2512 2294 2520
rect 2306 2512 2307 2520
rect 2309 2516 2310 2520
rect 2309 2512 2314 2516
rect 2322 2512 2323 2520
rect 2325 2512 2328 2520
rect 2330 2512 2331 2520
rect 2348 2512 2349 2520
rect 2351 2512 2352 2520
rect 2364 2512 2365 2520
rect 2367 2516 2368 2520
rect 2367 2512 2372 2516
rect 2380 2512 2381 2520
rect 2383 2512 2386 2520
rect 2388 2512 2389 2520
rect 2401 2512 2402 2520
rect 2404 2512 2405 2520
rect 2417 2512 2418 2520
rect 2420 2512 2423 2520
rect 2425 2512 2426 2520
rect 2438 2512 2439 2520
rect 2441 2516 2442 2520
rect 2441 2512 2446 2516
rect 2454 2512 2455 2520
rect 2457 2512 2460 2520
rect 2462 2512 2463 2520
rect 2480 2512 2481 2520
rect 2483 2512 2484 2520
rect 2496 2512 2497 2520
rect 2499 2516 2500 2520
rect 2499 2512 2504 2516
rect 2512 2512 2513 2520
rect 2515 2512 2518 2520
rect 2520 2512 2521 2520
rect 2533 2512 2534 2520
rect 2536 2512 2537 2520
rect 2549 2512 2550 2520
rect 2552 2512 2555 2520
rect 2557 2512 2558 2520
rect 2570 2512 2571 2520
rect 2573 2516 2574 2520
rect 2573 2512 2578 2516
rect 2586 2512 2587 2520
rect 2589 2512 2592 2520
rect 2594 2512 2595 2520
rect 2612 2512 2613 2520
rect 2615 2512 2616 2520
rect 2628 2512 2629 2520
rect 2631 2516 2632 2520
rect 2631 2512 2636 2516
rect 2644 2512 2645 2520
rect 2647 2512 2650 2520
rect 2652 2512 2653 2520
rect 2665 2512 2666 2520
rect 2668 2512 2669 2520
rect 3230 2512 3231 2520
rect 3233 2512 3236 2520
rect 3238 2512 3239 2520
rect 3251 2512 3252 2520
rect 3254 2516 3255 2520
rect 3254 2512 3259 2516
rect 3267 2512 3268 2520
rect 3270 2512 3273 2520
rect 3275 2512 3276 2520
rect 3293 2512 3294 2520
rect 3296 2512 3297 2520
rect 3309 2512 3310 2520
rect 3312 2516 3313 2520
rect 3312 2512 3317 2516
rect 3325 2512 3326 2520
rect 3328 2512 3331 2520
rect 3333 2512 3334 2520
rect 3346 2512 3347 2520
rect 3349 2512 3350 2520
rect 3362 2512 3363 2520
rect 3365 2512 3368 2520
rect 3370 2512 3371 2520
rect 3383 2512 3384 2520
rect 3386 2516 3387 2520
rect 3386 2512 3391 2516
rect 3399 2512 3400 2520
rect 3402 2512 3405 2520
rect 3407 2512 3408 2520
rect 3425 2512 3426 2520
rect 3428 2512 3429 2520
rect 3441 2512 3442 2520
rect 3444 2516 3445 2520
rect 3444 2512 3449 2516
rect 3457 2512 3458 2520
rect 3460 2512 3463 2520
rect 3465 2512 3466 2520
rect 3478 2512 3479 2520
rect 3481 2512 3482 2520
rect 3494 2512 3495 2520
rect 3497 2512 3500 2520
rect 3502 2512 3503 2520
rect 3515 2512 3516 2520
rect 3518 2516 3519 2520
rect 3518 2512 3523 2516
rect 3531 2512 3532 2520
rect 3534 2512 3537 2520
rect 3539 2512 3540 2520
rect 3557 2512 3558 2520
rect 3560 2512 3561 2520
rect 3573 2512 3574 2520
rect 3576 2516 3577 2520
rect 3576 2512 3581 2516
rect 3589 2512 3590 2520
rect 3592 2512 3595 2520
rect 3597 2512 3598 2520
rect 3610 2512 3611 2520
rect 3613 2512 3614 2520
rect 2774 2481 2775 2489
rect 2777 2481 2778 2489
rect 2790 2481 2791 2489
rect 2793 2481 2794 2489
rect 2806 2481 2807 2489
rect 2809 2481 2810 2489
rect 2825 2481 2830 2489
rect 2832 2481 2835 2489
rect 2837 2481 2838 2489
rect 2859 2481 2861 2489
rect 2863 2481 2864 2489
rect 2881 2481 2882 2489
rect 2884 2481 2885 2489
rect 2897 2481 2902 2489
rect 2904 2481 2907 2489
rect 2909 2481 2910 2489
rect 2924 2481 2925 2489
rect 2927 2481 2928 2489
rect 2972 2476 2975 2484
rect 2977 2476 2980 2484
rect 2982 2476 2983 2484
rect 3008 2481 3009 2489
rect 3011 2481 3012 2489
rect 3016 2481 3022 2489
rect 3026 2481 3027 2489
rect 3029 2481 3030 2489
rect 3051 2481 3052 2489
rect 3054 2481 3055 2489
rect 3067 2481 3068 2489
rect 3070 2481 3071 2489
rect 3086 2481 3091 2489
rect 3093 2481 3096 2489
rect 3098 2481 3099 2489
rect 3120 2481 3122 2489
rect 3124 2481 3125 2489
rect 3142 2481 3143 2489
rect 3145 2481 3146 2489
rect 3158 2481 3163 2489
rect 3165 2481 3168 2489
rect 3170 2481 3171 2489
rect 3185 2481 3186 2489
rect 3188 2481 3189 2489
rect 3719 2481 3720 2489
rect 3722 2481 3723 2489
rect 3735 2481 3736 2489
rect 3738 2481 3739 2489
rect 3751 2481 3752 2489
rect 3754 2481 3755 2489
rect 3770 2481 3775 2489
rect 3777 2481 3780 2489
rect 3782 2481 3783 2489
rect 3804 2481 3806 2489
rect 3808 2481 3809 2489
rect 3826 2481 3827 2489
rect 3829 2481 3830 2489
rect 3842 2481 3847 2489
rect 3849 2481 3852 2489
rect 3854 2481 3855 2489
rect 3869 2481 3870 2489
rect 3872 2481 3873 2489
rect 3917 2476 3920 2484
rect 3922 2476 3925 2484
rect 3927 2476 3928 2484
rect 3953 2481 3954 2489
rect 3956 2481 3957 2489
rect 3961 2481 3967 2489
rect 3971 2481 3972 2489
rect 3974 2481 3975 2489
rect 3996 2481 3997 2489
rect 3999 2481 4000 2489
rect 4012 2481 4013 2489
rect 4015 2481 4016 2489
rect 4031 2481 4036 2489
rect 4038 2481 4041 2489
rect 4043 2481 4044 2489
rect 4065 2481 4067 2489
rect 4069 2481 4070 2489
rect 4087 2481 4088 2489
rect 4090 2481 4091 2489
rect 4103 2481 4108 2489
rect 4110 2481 4113 2489
rect 4115 2481 4116 2489
rect 4130 2481 4131 2489
rect 4133 2481 4134 2489
rect 3068 2400 3069 2408
rect 3071 2400 3074 2408
rect 3076 2400 3077 2408
rect 3089 2400 3090 2408
rect 3092 2404 3093 2408
rect 3092 2400 3097 2404
rect 3105 2400 3106 2408
rect 3108 2400 3111 2408
rect 3113 2400 3114 2408
rect 3131 2400 3132 2408
rect 3134 2400 3135 2408
rect 3147 2400 3148 2408
rect 3150 2404 3151 2408
rect 3150 2400 3155 2404
rect 3163 2400 3164 2408
rect 3166 2400 3169 2408
rect 3171 2400 3172 2408
rect 3184 2400 3185 2408
rect 3187 2400 3188 2408
rect 4013 2400 4014 2408
rect 4016 2400 4019 2408
rect 4021 2400 4022 2408
rect 4034 2400 4035 2408
rect 4037 2404 4038 2408
rect 4037 2400 4042 2404
rect 4050 2400 4051 2408
rect 4053 2400 4056 2408
rect 4058 2400 4059 2408
rect 4076 2400 4077 2408
rect 4079 2400 4080 2408
rect 4092 2400 4093 2408
rect 4095 2404 4096 2408
rect 4095 2400 4100 2404
rect 4108 2400 4109 2408
rect 4111 2400 4114 2408
rect 4116 2400 4117 2408
rect 4129 2400 4130 2408
rect 4132 2400 4133 2408
rect 2285 2370 2286 2378
rect 2288 2370 2291 2378
rect 2293 2370 2294 2378
rect 2306 2370 2307 2378
rect 2309 2374 2310 2378
rect 2309 2370 2314 2374
rect 2322 2370 2323 2378
rect 2325 2370 2328 2378
rect 2330 2370 2331 2378
rect 2348 2370 2349 2378
rect 2351 2370 2352 2378
rect 2364 2370 2365 2378
rect 2367 2374 2368 2378
rect 2367 2370 2372 2374
rect 2380 2370 2381 2378
rect 2383 2370 2386 2378
rect 2388 2370 2389 2378
rect 2401 2370 2402 2378
rect 2404 2370 2405 2378
rect 2417 2370 2418 2378
rect 2420 2370 2423 2378
rect 2425 2370 2426 2378
rect 2438 2370 2439 2378
rect 2441 2374 2442 2378
rect 2441 2370 2446 2374
rect 2454 2370 2455 2378
rect 2457 2370 2460 2378
rect 2462 2370 2463 2378
rect 2480 2370 2481 2378
rect 2483 2370 2484 2378
rect 2496 2370 2497 2378
rect 2499 2374 2500 2378
rect 2499 2370 2504 2374
rect 2512 2370 2513 2378
rect 2515 2370 2518 2378
rect 2520 2370 2521 2378
rect 2533 2370 2534 2378
rect 2536 2370 2537 2378
rect 2549 2370 2550 2378
rect 2552 2370 2555 2378
rect 2557 2370 2558 2378
rect 2570 2370 2571 2378
rect 2573 2374 2574 2378
rect 2573 2370 2578 2374
rect 2586 2370 2587 2378
rect 2589 2370 2592 2378
rect 2594 2370 2595 2378
rect 2612 2370 2613 2378
rect 2615 2370 2616 2378
rect 2628 2370 2629 2378
rect 2631 2374 2632 2378
rect 2631 2370 2636 2374
rect 2644 2370 2645 2378
rect 2647 2370 2650 2378
rect 2652 2370 2653 2378
rect 2665 2370 2666 2378
rect 2668 2370 2669 2378
rect 3230 2370 3231 2378
rect 3233 2370 3236 2378
rect 3238 2370 3239 2378
rect 3251 2370 3252 2378
rect 3254 2374 3255 2378
rect 3254 2370 3259 2374
rect 3267 2370 3268 2378
rect 3270 2370 3273 2378
rect 3275 2370 3276 2378
rect 3293 2370 3294 2378
rect 3296 2370 3297 2378
rect 3309 2370 3310 2378
rect 3312 2374 3313 2378
rect 3312 2370 3317 2374
rect 3325 2370 3326 2378
rect 3328 2370 3331 2378
rect 3333 2370 3334 2378
rect 3346 2370 3347 2378
rect 3349 2370 3350 2378
rect 3362 2370 3363 2378
rect 3365 2370 3368 2378
rect 3370 2370 3371 2378
rect 3383 2370 3384 2378
rect 3386 2374 3387 2378
rect 3386 2370 3391 2374
rect 3399 2370 3400 2378
rect 3402 2370 3405 2378
rect 3407 2370 3408 2378
rect 3425 2370 3426 2378
rect 3428 2370 3429 2378
rect 3441 2370 3442 2378
rect 3444 2374 3445 2378
rect 3444 2370 3449 2374
rect 3457 2370 3458 2378
rect 3460 2370 3463 2378
rect 3465 2370 3466 2378
rect 3478 2370 3479 2378
rect 3481 2370 3482 2378
rect 3494 2370 3495 2378
rect 3497 2370 3500 2378
rect 3502 2370 3503 2378
rect 3515 2370 3516 2378
rect 3518 2374 3519 2378
rect 3518 2370 3523 2374
rect 3531 2370 3532 2378
rect 3534 2370 3537 2378
rect 3539 2370 3540 2378
rect 3557 2370 3558 2378
rect 3560 2370 3561 2378
rect 3573 2370 3574 2378
rect 3576 2374 3577 2378
rect 3576 2370 3581 2374
rect 3589 2370 3590 2378
rect 3592 2370 3595 2378
rect 3597 2370 3598 2378
rect 3610 2370 3611 2378
rect 3613 2370 3614 2378
rect 3068 2314 3069 2322
rect 3071 2314 3074 2322
rect 3076 2314 3077 2322
rect 3089 2314 3090 2322
rect 3092 2318 3093 2322
rect 3092 2314 3097 2318
rect 3105 2314 3106 2322
rect 3108 2314 3111 2322
rect 3113 2314 3114 2322
rect 3131 2314 3132 2322
rect 3134 2314 3135 2322
rect 3147 2314 3148 2322
rect 3150 2318 3151 2322
rect 3150 2314 3155 2318
rect 3163 2314 3164 2322
rect 3166 2314 3169 2322
rect 3171 2314 3172 2322
rect 3184 2314 3185 2322
rect 3187 2314 3188 2322
rect 4013 2314 4014 2322
rect 4016 2314 4019 2322
rect 4021 2314 4022 2322
rect 4034 2314 4035 2322
rect 4037 2318 4038 2322
rect 4037 2314 4042 2318
rect 4050 2314 4051 2322
rect 4053 2314 4056 2322
rect 4058 2314 4059 2322
rect 4076 2314 4077 2322
rect 4079 2314 4080 2322
rect 4092 2314 4093 2322
rect 4095 2318 4096 2322
rect 4095 2314 4100 2318
rect 4108 2314 4109 2322
rect 4111 2314 4114 2322
rect 4116 2314 4117 2322
rect 4129 2314 4130 2322
rect 4132 2314 4133 2322
rect 2285 2284 2286 2292
rect 2288 2284 2291 2292
rect 2293 2284 2294 2292
rect 2306 2284 2307 2292
rect 2309 2288 2310 2292
rect 2309 2284 2314 2288
rect 2322 2284 2323 2292
rect 2325 2284 2328 2292
rect 2330 2284 2331 2292
rect 2348 2284 2349 2292
rect 2351 2284 2352 2292
rect 2364 2284 2365 2292
rect 2367 2288 2368 2292
rect 2367 2284 2372 2288
rect 2380 2284 2381 2292
rect 2383 2284 2386 2292
rect 2388 2284 2389 2292
rect 2401 2284 2402 2292
rect 2404 2284 2405 2292
rect 2417 2284 2418 2292
rect 2420 2284 2423 2292
rect 2425 2284 2426 2292
rect 2438 2284 2439 2292
rect 2441 2288 2442 2292
rect 2441 2284 2446 2288
rect 2454 2284 2455 2292
rect 2457 2284 2460 2292
rect 2462 2284 2463 2292
rect 2480 2284 2481 2292
rect 2483 2284 2484 2292
rect 2496 2284 2497 2292
rect 2499 2288 2500 2292
rect 2499 2284 2504 2288
rect 2512 2284 2513 2292
rect 2515 2284 2518 2292
rect 2520 2284 2521 2292
rect 2533 2284 2534 2292
rect 2536 2284 2537 2292
rect 2549 2284 2550 2292
rect 2552 2284 2555 2292
rect 2557 2284 2558 2292
rect 2570 2284 2571 2292
rect 2573 2288 2574 2292
rect 2573 2284 2578 2288
rect 2586 2284 2587 2292
rect 2589 2284 2592 2292
rect 2594 2284 2595 2292
rect 2612 2284 2613 2292
rect 2615 2284 2616 2292
rect 2628 2284 2629 2292
rect 2631 2288 2632 2292
rect 2631 2284 2636 2288
rect 2644 2284 2645 2292
rect 2647 2284 2650 2292
rect 2652 2284 2653 2292
rect 2665 2284 2666 2292
rect 2668 2284 2669 2292
rect 3230 2284 3231 2292
rect 3233 2284 3236 2292
rect 3238 2284 3239 2292
rect 3251 2284 3252 2292
rect 3254 2288 3255 2292
rect 3254 2284 3259 2288
rect 3267 2284 3268 2292
rect 3270 2284 3273 2292
rect 3275 2284 3276 2292
rect 3293 2284 3294 2292
rect 3296 2284 3297 2292
rect 3309 2284 3310 2292
rect 3312 2288 3313 2292
rect 3312 2284 3317 2288
rect 3325 2284 3326 2292
rect 3328 2284 3331 2292
rect 3333 2284 3334 2292
rect 3346 2284 3347 2292
rect 3349 2284 3350 2292
rect 3362 2284 3363 2292
rect 3365 2284 3368 2292
rect 3370 2284 3371 2292
rect 3383 2284 3384 2292
rect 3386 2288 3387 2292
rect 3386 2284 3391 2288
rect 3399 2284 3400 2292
rect 3402 2284 3405 2292
rect 3407 2284 3408 2292
rect 3425 2284 3426 2292
rect 3428 2284 3429 2292
rect 3441 2284 3442 2292
rect 3444 2288 3445 2292
rect 3444 2284 3449 2288
rect 3457 2284 3458 2292
rect 3460 2284 3463 2292
rect 3465 2284 3466 2292
rect 3478 2284 3479 2292
rect 3481 2284 3482 2292
rect 3494 2284 3495 2292
rect 3497 2284 3500 2292
rect 3502 2284 3503 2292
rect 3515 2284 3516 2292
rect 3518 2288 3519 2292
rect 3518 2284 3523 2288
rect 3531 2284 3532 2292
rect 3534 2284 3537 2292
rect 3539 2284 3540 2292
rect 3557 2284 3558 2292
rect 3560 2284 3561 2292
rect 3573 2284 3574 2292
rect 3576 2288 3577 2292
rect 3576 2284 3581 2288
rect 3589 2284 3590 2292
rect 3592 2284 3595 2292
rect 3597 2284 3598 2292
rect 3610 2284 3611 2292
rect 3613 2284 3614 2292
rect 2285 2144 2286 2152
rect 2288 2144 2291 2152
rect 2293 2144 2294 2152
rect 2306 2144 2307 2152
rect 2309 2148 2310 2152
rect 2309 2144 2314 2148
rect 2322 2144 2323 2152
rect 2325 2144 2328 2152
rect 2330 2144 2331 2152
rect 2348 2144 2349 2152
rect 2351 2144 2352 2152
rect 2364 2144 2365 2152
rect 2367 2148 2368 2152
rect 2367 2144 2372 2148
rect 2380 2144 2381 2152
rect 2383 2144 2386 2152
rect 2388 2144 2389 2152
rect 2401 2144 2402 2152
rect 2404 2144 2405 2152
rect 2417 2144 2418 2152
rect 2420 2144 2423 2152
rect 2425 2144 2426 2152
rect 2438 2144 2439 2152
rect 2441 2148 2442 2152
rect 2441 2144 2446 2148
rect 2454 2144 2455 2152
rect 2457 2144 2460 2152
rect 2462 2144 2463 2152
rect 2480 2144 2481 2152
rect 2483 2144 2484 2152
rect 2496 2144 2497 2152
rect 2499 2148 2500 2152
rect 2499 2144 2504 2148
rect 2512 2144 2513 2152
rect 2515 2144 2518 2152
rect 2520 2144 2521 2152
rect 2533 2144 2534 2152
rect 2536 2144 2537 2152
rect 2549 2144 2550 2152
rect 2552 2144 2555 2152
rect 2557 2144 2558 2152
rect 2570 2144 2571 2152
rect 2573 2148 2574 2152
rect 2573 2144 2578 2148
rect 2586 2144 2587 2152
rect 2589 2144 2592 2152
rect 2594 2144 2595 2152
rect 2612 2144 2613 2152
rect 2615 2144 2616 2152
rect 2628 2144 2629 2152
rect 2631 2148 2632 2152
rect 2631 2144 2636 2148
rect 2644 2144 2645 2152
rect 2647 2144 2650 2152
rect 2652 2144 2653 2152
rect 2665 2144 2666 2152
rect 2668 2144 2669 2152
rect 3230 2144 3231 2152
rect 3233 2144 3236 2152
rect 3238 2144 3239 2152
rect 3251 2144 3252 2152
rect 3254 2148 3255 2152
rect 3254 2144 3259 2148
rect 3267 2144 3268 2152
rect 3270 2144 3273 2152
rect 3275 2144 3276 2152
rect 3293 2144 3294 2152
rect 3296 2144 3297 2152
rect 3309 2144 3310 2152
rect 3312 2148 3313 2152
rect 3312 2144 3317 2148
rect 3325 2144 3326 2152
rect 3328 2144 3331 2152
rect 3333 2144 3334 2152
rect 3346 2144 3347 2152
rect 3349 2144 3350 2152
rect 3362 2144 3363 2152
rect 3365 2144 3368 2152
rect 3370 2144 3371 2152
rect 3383 2144 3384 2152
rect 3386 2148 3387 2152
rect 3386 2144 3391 2148
rect 3399 2144 3400 2152
rect 3402 2144 3405 2152
rect 3407 2144 3408 2152
rect 3425 2144 3426 2152
rect 3428 2144 3429 2152
rect 3441 2144 3442 2152
rect 3444 2148 3445 2152
rect 3444 2144 3449 2148
rect 3457 2144 3458 2152
rect 3460 2144 3463 2152
rect 3465 2144 3466 2152
rect 3478 2144 3479 2152
rect 3481 2144 3482 2152
rect 3494 2144 3495 2152
rect 3497 2144 3500 2152
rect 3502 2144 3503 2152
rect 3515 2144 3516 2152
rect 3518 2148 3519 2152
rect 3518 2144 3523 2148
rect 3531 2144 3532 2152
rect 3534 2144 3537 2152
rect 3539 2144 3540 2152
rect 3557 2144 3558 2152
rect 3560 2144 3561 2152
rect 3573 2144 3574 2152
rect 3576 2148 3577 2152
rect 3576 2144 3581 2148
rect 3589 2144 3590 2152
rect 3592 2144 3595 2152
rect 3597 2144 3598 2152
rect 3610 2144 3611 2152
rect 3613 2144 3614 2152
<< ndcontact >>
rect 2765 4006 2769 4010
rect 2778 4006 2782 4010
rect 2786 4006 2790 4010
rect 2794 4006 2798 4010
rect 2802 4006 2806 4010
rect 2815 4006 2819 4010
rect 2828 4006 2832 4010
rect 2836 4006 2840 4010
rect 2844 4006 2848 4010
rect 2852 4006 2856 4010
rect 2860 4006 2864 4010
rect 2873 4006 2877 4010
rect 2881 4006 2885 4010
rect 2889 4006 2893 4010
rect 2897 4006 2901 4010
rect 2910 4006 2914 4010
rect 2918 4006 2922 4010
rect 2926 4006 2930 4010
rect 2934 4006 2938 4010
rect 2947 4006 2951 4010
rect 2960 4006 2964 4010
rect 2968 4006 2972 4010
rect 2976 4006 2980 4010
rect 2984 4006 2988 4010
rect 2992 4006 2996 4010
rect 3005 4006 3009 4010
rect 3013 4006 3017 4010
rect 3021 4006 3025 4010
rect 3029 4006 3033 4010
rect 3042 4006 3046 4010
rect 3050 4006 3054 4010
rect 3058 4006 3062 4010
rect 3066 4006 3070 4010
rect 3079 4006 3083 4010
rect 3092 4006 3096 4010
rect 3100 4006 3104 4010
rect 3108 4006 3112 4010
rect 3116 4006 3120 4010
rect 3124 4006 3128 4010
rect 3137 4006 3141 4010
rect 3145 4006 3149 4010
rect 3153 4006 3157 4010
rect 3161 4006 3165 4010
rect 3174 4006 3178 4010
rect 3182 4006 3186 4010
rect 3190 4006 3194 4010
rect 3198 4006 3202 4010
rect 3211 4006 3215 4010
rect 3224 4006 3228 4010
rect 3232 4006 3236 4010
rect 3240 4006 3244 4010
rect 3248 4006 3252 4010
rect 3256 4006 3260 4010
rect 3269 4006 3273 4010
rect 3277 4006 3281 4010
rect 3285 4006 3289 4010
rect 3710 4006 3714 4010
rect 3723 4006 3727 4010
rect 3731 4006 3735 4010
rect 3739 4006 3743 4010
rect 3747 4006 3751 4010
rect 3760 4006 3764 4010
rect 3773 4006 3777 4010
rect 3781 4006 3785 4010
rect 3789 4006 3793 4010
rect 3797 4006 3801 4010
rect 3805 4006 3809 4010
rect 3818 4006 3822 4010
rect 3826 4006 3830 4010
rect 3834 4006 3838 4010
rect 3842 4006 3846 4010
rect 3855 4006 3859 4010
rect 3863 4006 3867 4010
rect 3871 4006 3875 4010
rect 3879 4006 3883 4010
rect 3892 4006 3896 4010
rect 3905 4006 3909 4010
rect 3913 4006 3917 4010
rect 3921 4006 3925 4010
rect 3929 4006 3933 4010
rect 3937 4006 3941 4010
rect 3950 4006 3954 4010
rect 3958 4006 3962 4010
rect 3966 4006 3970 4010
rect 3974 4006 3978 4010
rect 3987 4006 3991 4010
rect 3995 4006 3999 4010
rect 4003 4006 4007 4010
rect 4011 4006 4015 4010
rect 4024 4006 4028 4010
rect 4037 4006 4041 4010
rect 4045 4006 4049 4010
rect 4053 4006 4057 4010
rect 4061 4006 4065 4010
rect 4069 4006 4073 4010
rect 4082 4006 4086 4010
rect 4090 4006 4094 4010
rect 4098 4006 4102 4010
rect 4106 4006 4110 4010
rect 4119 4006 4123 4010
rect 4127 4006 4131 4010
rect 4135 4006 4139 4010
rect 4143 4006 4147 4010
rect 4156 4006 4160 4010
rect 4169 4006 4173 4010
rect 4177 4006 4181 4010
rect 4185 4006 4189 4010
rect 4193 4006 4197 4010
rect 4201 4006 4205 4010
rect 4214 4006 4218 4010
rect 4222 4006 4226 4010
rect 4230 4006 4234 4010
rect 2413 3973 2417 3977
rect 2426 3973 2430 3977
rect 2434 3973 2438 3977
rect 2442 3973 2446 3977
rect 2450 3973 2454 3977
rect 2463 3973 2467 3977
rect 2476 3973 2480 3977
rect 2484 3973 2488 3977
rect 2492 3973 2496 3977
rect 2500 3973 2504 3977
rect 2508 3973 2512 3977
rect 2521 3973 2525 3977
rect 2529 3973 2533 3977
rect 2537 3973 2541 3977
rect 3358 3973 3362 3977
rect 3371 3973 3375 3977
rect 3379 3973 3383 3977
rect 3387 3973 3391 3977
rect 3395 3973 3399 3977
rect 3408 3973 3412 3977
rect 3421 3973 3425 3977
rect 3429 3973 3433 3977
rect 3437 3973 3441 3977
rect 3445 3973 3449 3977
rect 3453 3973 3457 3977
rect 3466 3973 3470 3977
rect 3474 3973 3478 3977
rect 3482 3973 3486 3977
rect 2537 3936 2541 3940
rect 2545 3936 2549 3940
rect 2944 3940 2948 3944
rect 2952 3940 2956 3944
rect 2968 3936 2972 3940
rect 2983 3936 2987 3940
rect 3025 3940 3029 3944
rect 3033 3940 3037 3944
rect 3049 3936 3053 3940
rect 3064 3936 3068 3940
rect 2998 3932 3002 3936
rect 3006 3932 3010 3936
rect 2420 3927 2424 3931
rect 2428 3927 2432 3931
rect 2770 3927 2774 3931
rect 2778 3927 2782 3931
rect 2786 3927 2790 3931
rect 2794 3927 2798 3931
rect 2802 3927 2806 3931
rect 2810 3927 2814 3931
rect 2821 3927 2825 3931
rect 2838 3927 2842 3931
rect 2855 3927 2859 3931
rect 2864 3927 2868 3931
rect 2877 3927 2881 3931
rect 2885 3927 2889 3931
rect 2893 3927 2897 3931
rect 2910 3927 2914 3931
rect 2920 3927 2924 3931
rect 2928 3927 2932 3931
rect 3079 3932 3083 3936
rect 3087 3932 3091 3936
rect 3482 3936 3486 3940
rect 3490 3936 3494 3940
rect 3889 3940 3893 3944
rect 3897 3940 3901 3944
rect 3913 3936 3917 3940
rect 3928 3936 3932 3940
rect 3970 3940 3974 3944
rect 3978 3940 3982 3944
rect 3994 3936 3998 3940
rect 4009 3936 4013 3940
rect 3943 3932 3947 3936
rect 3951 3932 3955 3936
rect 3365 3927 3369 3931
rect 3373 3927 3377 3931
rect 3715 3927 3719 3931
rect 3723 3927 3727 3931
rect 3731 3927 3735 3931
rect 3739 3927 3743 3931
rect 3747 3927 3751 3931
rect 3755 3927 3759 3931
rect 3766 3927 3770 3931
rect 3783 3927 3787 3931
rect 3800 3927 3804 3931
rect 3809 3927 3813 3931
rect 3822 3927 3826 3931
rect 3830 3927 3834 3931
rect 3838 3927 3842 3931
rect 3855 3927 3859 3931
rect 3865 3927 3869 3931
rect 3873 3927 3877 3931
rect 4024 3932 4028 3936
rect 4032 3932 4036 3936
rect 2770 3881 2774 3885
rect 2778 3881 2782 3885
rect 2786 3881 2790 3885
rect 2794 3881 2798 3885
rect 2802 3881 2806 3885
rect 2810 3881 2814 3885
rect 2821 3881 2825 3885
rect 2838 3881 2842 3885
rect 2855 3881 2859 3885
rect 2864 3881 2868 3885
rect 2877 3881 2881 3885
rect 2885 3881 2889 3885
rect 2893 3881 2897 3885
rect 2910 3881 2914 3885
rect 2920 3881 2924 3885
rect 2928 3881 2932 3885
rect 2404 3871 2408 3875
rect 2412 3871 2416 3875
rect 2420 3871 2424 3875
rect 2433 3871 2437 3875
rect 2441 3871 2445 3875
rect 2449 3871 2453 3875
rect 2457 3871 2461 3875
rect 2465 3871 2469 3875
rect 2478 3871 2482 3875
rect 2491 3871 2495 3875
rect 2499 3871 2503 3875
rect 2507 3871 2511 3875
rect 2515 3871 2519 3875
rect 2528 3871 2532 3875
rect 2968 3880 2972 3884
rect 2983 3880 2987 3884
rect 3049 3880 3053 3884
rect 3064 3880 3068 3884
rect 3715 3881 3719 3885
rect 3723 3881 3727 3885
rect 3731 3881 3735 3885
rect 3739 3881 3743 3885
rect 3747 3881 3751 3885
rect 3755 3881 3759 3885
rect 3766 3881 3770 3885
rect 3783 3881 3787 3885
rect 3800 3881 3804 3885
rect 3809 3881 3813 3885
rect 3822 3881 3826 3885
rect 3830 3881 3834 3885
rect 3838 3881 3842 3885
rect 3855 3881 3859 3885
rect 3865 3881 3869 3885
rect 3873 3881 3877 3885
rect 3349 3871 3353 3875
rect 3357 3871 3361 3875
rect 3365 3871 3369 3875
rect 3378 3871 3382 3875
rect 3386 3871 3390 3875
rect 3394 3871 3398 3875
rect 3402 3871 3406 3875
rect 3410 3871 3414 3875
rect 3423 3871 3427 3875
rect 3436 3871 3440 3875
rect 3444 3871 3448 3875
rect 3452 3871 3456 3875
rect 3460 3871 3464 3875
rect 3473 3871 3477 3875
rect 3913 3880 3917 3884
rect 3928 3880 3932 3884
rect 3994 3880 3998 3884
rect 4009 3880 4013 3884
rect 2968 3804 2972 3808
rect 2983 3804 2987 3808
rect 3049 3808 3053 3812
rect 3057 3808 3061 3812
rect 3073 3804 3077 3808
rect 3088 3804 3092 3808
rect 2998 3800 3002 3804
rect 3006 3800 3010 3804
rect 2770 3795 2774 3799
rect 2778 3795 2782 3799
rect 2786 3795 2790 3799
rect 2794 3795 2798 3799
rect 2802 3795 2806 3799
rect 2810 3795 2814 3799
rect 2821 3795 2825 3799
rect 2838 3795 2842 3799
rect 2855 3795 2859 3799
rect 2864 3795 2868 3799
rect 2877 3795 2881 3799
rect 2885 3795 2889 3799
rect 2893 3795 2897 3799
rect 2910 3795 2914 3799
rect 2920 3795 2924 3799
rect 2928 3795 2932 3799
rect 3103 3800 3107 3804
rect 3111 3800 3115 3804
rect 3280 3779 3284 3783
rect 3288 3779 3292 3783
rect 3304 3775 3308 3779
rect 3319 3775 3323 3779
rect 3334 3771 3338 3775
rect 3342 3771 3346 3775
rect 3913 3804 3917 3808
rect 3928 3804 3932 3808
rect 3994 3808 3998 3812
rect 4002 3808 4006 3812
rect 4018 3804 4022 3808
rect 4033 3804 4037 3808
rect 3943 3800 3947 3804
rect 3951 3800 3955 3804
rect 3715 3795 3719 3799
rect 3723 3795 3727 3799
rect 3731 3795 3735 3799
rect 3739 3795 3743 3799
rect 3747 3795 3751 3799
rect 3755 3795 3759 3799
rect 3766 3795 3770 3799
rect 3783 3795 3787 3799
rect 3800 3795 3804 3799
rect 3809 3795 3813 3799
rect 3822 3795 3826 3799
rect 3830 3795 3834 3799
rect 3838 3795 3842 3799
rect 3855 3795 3859 3799
rect 3865 3795 3869 3799
rect 3873 3795 3877 3799
rect 4048 3800 4052 3804
rect 4056 3800 4060 3804
rect 2770 3749 2774 3753
rect 2778 3749 2782 3753
rect 2786 3749 2790 3753
rect 2794 3749 2798 3753
rect 2802 3749 2806 3753
rect 2810 3749 2814 3753
rect 2821 3749 2825 3753
rect 2838 3749 2842 3753
rect 2855 3749 2859 3753
rect 2864 3749 2868 3753
rect 2877 3749 2881 3753
rect 2885 3749 2889 3753
rect 2893 3749 2897 3753
rect 2910 3749 2914 3753
rect 2920 3749 2924 3753
rect 2928 3749 2932 3753
rect 2968 3749 2972 3753
rect 2983 3749 2987 3753
rect 3073 3749 3077 3753
rect 3088 3749 3092 3753
rect 3454 3740 3470 3752
rect 3474 3740 3490 3752
rect 3507 3740 3523 3752
rect 3527 3740 3543 3752
rect 3715 3749 3719 3753
rect 3723 3749 3727 3753
rect 3731 3749 3735 3753
rect 3739 3749 3743 3753
rect 3747 3749 3751 3753
rect 3755 3749 3759 3753
rect 3766 3749 3770 3753
rect 3783 3749 3787 3753
rect 3800 3749 3804 3753
rect 3809 3749 3813 3753
rect 3822 3749 3826 3753
rect 3830 3749 3834 3753
rect 3838 3749 3842 3753
rect 3855 3749 3859 3753
rect 3865 3749 3869 3753
rect 3873 3749 3877 3753
rect 3913 3749 3917 3753
rect 3928 3749 3932 3753
rect 4018 3749 4022 3753
rect 4033 3749 4037 3753
rect 3304 3715 3308 3719
rect 3319 3715 3323 3719
rect 2968 3672 2972 3676
rect 2983 3672 2987 3676
rect 3025 3676 3029 3680
rect 3033 3676 3037 3680
rect 3049 3672 3053 3676
rect 3064 3672 3068 3676
rect 3115 3676 3119 3680
rect 3123 3676 3127 3680
rect 3139 3672 3143 3676
rect 3154 3672 3158 3676
rect 2998 3668 3002 3672
rect 3006 3668 3010 3672
rect 2770 3663 2774 3667
rect 2778 3663 2782 3667
rect 2786 3663 2790 3667
rect 2794 3663 2798 3667
rect 2802 3663 2806 3667
rect 2810 3663 2814 3667
rect 2821 3663 2825 3667
rect 2838 3663 2842 3667
rect 2855 3663 2859 3667
rect 2864 3663 2868 3667
rect 2877 3663 2881 3667
rect 2885 3663 2889 3667
rect 2893 3663 2897 3667
rect 2910 3663 2914 3667
rect 2920 3663 2924 3667
rect 2928 3663 2932 3667
rect 3079 3668 3083 3672
rect 3087 3668 3091 3672
rect 3169 3668 3173 3672
rect 3177 3668 3181 3672
rect 3258 3649 3262 3653
rect 3266 3649 3270 3653
rect 3280 3649 3284 3653
rect 3288 3649 3292 3653
rect 3304 3645 3308 3649
rect 3319 3645 3323 3649
rect 3334 3641 3338 3645
rect 3342 3641 3346 3645
rect 3913 3672 3917 3676
rect 3928 3672 3932 3676
rect 3970 3676 3974 3680
rect 3978 3676 3982 3680
rect 3994 3672 3998 3676
rect 4009 3672 4013 3676
rect 4060 3676 4064 3680
rect 4068 3676 4072 3680
rect 4084 3672 4088 3676
rect 4099 3672 4103 3676
rect 3943 3668 3947 3672
rect 3951 3668 3955 3672
rect 3715 3663 3719 3667
rect 3723 3663 3727 3667
rect 3731 3663 3735 3667
rect 3739 3663 3743 3667
rect 3747 3663 3751 3667
rect 3755 3663 3759 3667
rect 3766 3663 3770 3667
rect 3783 3663 3787 3667
rect 3800 3663 3804 3667
rect 3809 3663 3813 3667
rect 3822 3663 3826 3667
rect 3830 3663 3834 3667
rect 3838 3663 3842 3667
rect 3855 3663 3859 3667
rect 3865 3663 3869 3667
rect 3873 3663 3877 3667
rect 4024 3668 4028 3672
rect 4032 3668 4036 3672
rect 4114 3668 4118 3672
rect 4122 3668 4126 3672
rect 2770 3617 2774 3621
rect 2778 3617 2782 3621
rect 2786 3617 2790 3621
rect 2794 3617 2798 3621
rect 2802 3617 2806 3621
rect 2810 3617 2814 3621
rect 2821 3617 2825 3621
rect 2838 3617 2842 3621
rect 2855 3617 2859 3621
rect 2864 3617 2868 3621
rect 2877 3617 2881 3621
rect 2885 3617 2889 3621
rect 2893 3617 2897 3621
rect 2910 3617 2914 3621
rect 2920 3617 2924 3621
rect 2928 3617 2932 3621
rect 2968 3614 2972 3618
rect 2983 3614 2987 3618
rect 3049 3614 3053 3618
rect 3064 3614 3068 3618
rect 3139 3614 3143 3618
rect 3154 3614 3158 3618
rect 3360 3610 3376 3622
rect 3380 3610 3396 3622
rect 3413 3610 3429 3622
rect 3433 3610 3449 3622
rect 3715 3617 3719 3621
rect 3723 3617 3727 3621
rect 3731 3617 3735 3621
rect 3739 3617 3743 3621
rect 3747 3617 3751 3621
rect 3755 3617 3759 3621
rect 3766 3617 3770 3621
rect 3783 3617 3787 3621
rect 3800 3617 3804 3621
rect 3809 3617 3813 3621
rect 3822 3617 3826 3621
rect 3830 3617 3834 3621
rect 3838 3617 3842 3621
rect 3855 3617 3859 3621
rect 3865 3617 3869 3621
rect 3873 3617 3877 3621
rect 3913 3614 3917 3618
rect 3928 3614 3932 3618
rect 3994 3614 3998 3618
rect 4009 3614 4013 3618
rect 4084 3614 4088 3618
rect 4099 3614 4103 3618
rect 3304 3585 3308 3589
rect 3319 3585 3323 3589
rect 2968 3540 2972 3544
rect 2983 3540 2987 3544
rect 2998 3536 3002 3540
rect 3006 3536 3010 3540
rect 2770 3531 2774 3535
rect 2778 3531 2782 3535
rect 2786 3531 2790 3535
rect 2794 3531 2798 3535
rect 2802 3531 2806 3535
rect 2810 3531 2814 3535
rect 2821 3531 2825 3535
rect 2838 3531 2842 3535
rect 2855 3531 2859 3535
rect 2864 3531 2868 3535
rect 2877 3531 2881 3535
rect 2885 3531 2889 3535
rect 2893 3531 2897 3535
rect 2910 3531 2914 3535
rect 2920 3531 2924 3535
rect 2928 3531 2932 3535
rect 3913 3540 3917 3544
rect 3928 3540 3932 3544
rect 3943 3536 3947 3540
rect 3951 3536 3955 3540
rect 3715 3531 3719 3535
rect 3723 3531 3727 3535
rect 3731 3531 3735 3535
rect 3739 3531 3743 3535
rect 3747 3531 3751 3535
rect 3755 3531 3759 3535
rect 3766 3531 3770 3535
rect 3783 3531 3787 3535
rect 3800 3531 3804 3535
rect 3809 3531 3813 3535
rect 3822 3531 3826 3535
rect 3830 3531 3834 3535
rect 3838 3531 3842 3535
rect 3855 3531 3859 3535
rect 3865 3531 3869 3535
rect 3873 3531 3877 3535
rect 2770 3485 2774 3489
rect 2778 3485 2782 3489
rect 2786 3485 2790 3489
rect 2794 3485 2798 3489
rect 2802 3485 2806 3489
rect 2810 3485 2814 3489
rect 2821 3485 2825 3489
rect 2838 3485 2842 3489
rect 2855 3485 2859 3489
rect 2864 3485 2868 3489
rect 2877 3485 2881 3489
rect 2885 3485 2889 3489
rect 2893 3485 2897 3489
rect 2910 3485 2914 3489
rect 2920 3485 2924 3489
rect 2928 3485 2932 3489
rect 3004 3485 3008 3489
rect 3012 3485 3016 3489
rect 3022 3485 3026 3489
rect 3030 3485 3034 3489
rect 3039 3485 3043 3489
rect 3047 3485 3051 3489
rect 3055 3485 3059 3489
rect 3063 3485 3067 3489
rect 3071 3485 3075 3489
rect 3082 3485 3086 3489
rect 3099 3485 3103 3489
rect 3116 3485 3120 3489
rect 3125 3485 3129 3489
rect 3138 3485 3142 3489
rect 3146 3485 3150 3489
rect 3154 3485 3158 3489
rect 3171 3485 3175 3489
rect 3181 3485 3185 3489
rect 3189 3485 3193 3489
rect 2281 3471 2285 3475
rect 2294 3471 2298 3475
rect 2302 3471 2306 3475
rect 2310 3471 2314 3475
rect 2318 3471 2322 3475
rect 2331 3471 2335 3475
rect 2344 3471 2348 3475
rect 2352 3471 2356 3475
rect 2360 3471 2364 3475
rect 2368 3471 2372 3475
rect 2376 3471 2380 3475
rect 2389 3471 2393 3475
rect 2397 3471 2401 3475
rect 2405 3471 2409 3475
rect 2413 3471 2417 3475
rect 2426 3471 2430 3475
rect 2434 3471 2438 3475
rect 2442 3471 2446 3475
rect 2450 3471 2454 3475
rect 2463 3471 2467 3475
rect 2476 3471 2480 3475
rect 2484 3471 2488 3475
rect 2492 3471 2496 3475
rect 2500 3471 2504 3475
rect 2508 3471 2512 3475
rect 2521 3471 2525 3475
rect 2529 3471 2533 3475
rect 2537 3471 2541 3475
rect 2545 3471 2549 3475
rect 2558 3471 2562 3475
rect 2566 3471 2570 3475
rect 2574 3471 2578 3475
rect 2582 3471 2586 3475
rect 2595 3471 2599 3475
rect 2608 3471 2612 3475
rect 2616 3471 2620 3475
rect 2624 3471 2628 3475
rect 2632 3471 2636 3475
rect 2640 3471 2644 3475
rect 2653 3471 2657 3475
rect 2661 3471 2665 3475
rect 2669 3471 2673 3475
rect 2968 3478 2972 3482
rect 2983 3478 2987 3482
rect 3715 3485 3719 3489
rect 3723 3485 3727 3489
rect 3731 3485 3735 3489
rect 3739 3485 3743 3489
rect 3747 3485 3751 3489
rect 3755 3485 3759 3489
rect 3766 3485 3770 3489
rect 3783 3485 3787 3489
rect 3800 3485 3804 3489
rect 3809 3485 3813 3489
rect 3822 3485 3826 3489
rect 3830 3485 3834 3489
rect 3838 3485 3842 3489
rect 3855 3485 3859 3489
rect 3865 3485 3869 3489
rect 3873 3485 3877 3489
rect 3949 3485 3953 3489
rect 3957 3485 3961 3489
rect 3967 3485 3971 3489
rect 3975 3485 3979 3489
rect 3984 3485 3988 3489
rect 3992 3485 3996 3489
rect 4000 3485 4004 3489
rect 4008 3485 4012 3489
rect 4016 3485 4020 3489
rect 4027 3485 4031 3489
rect 4044 3485 4048 3489
rect 4061 3485 4065 3489
rect 4070 3485 4074 3489
rect 4083 3485 4087 3489
rect 4091 3485 4095 3489
rect 4099 3485 4103 3489
rect 4116 3485 4120 3489
rect 4126 3485 4130 3489
rect 4134 3485 4138 3489
rect 3226 3471 3230 3475
rect 3239 3471 3243 3475
rect 3247 3471 3251 3475
rect 3255 3471 3259 3475
rect 3263 3471 3267 3475
rect 3276 3471 3280 3475
rect 3289 3471 3293 3475
rect 3297 3471 3301 3475
rect 3305 3471 3309 3475
rect 3313 3471 3317 3475
rect 3321 3471 3325 3475
rect 3334 3471 3338 3475
rect 3342 3471 3346 3475
rect 3350 3471 3354 3475
rect 3358 3471 3362 3475
rect 3371 3471 3375 3475
rect 3379 3471 3383 3475
rect 3387 3471 3391 3475
rect 3395 3471 3399 3475
rect 3408 3471 3412 3475
rect 3421 3471 3425 3475
rect 3429 3471 3433 3475
rect 3437 3471 3441 3475
rect 3445 3471 3449 3475
rect 3453 3471 3457 3475
rect 3466 3471 3470 3475
rect 3474 3471 3478 3475
rect 3482 3471 3486 3475
rect 3490 3471 3494 3475
rect 3503 3471 3507 3475
rect 3511 3471 3515 3475
rect 3519 3471 3523 3475
rect 3527 3471 3531 3475
rect 3540 3471 3544 3475
rect 3553 3471 3557 3475
rect 3561 3471 3565 3475
rect 3569 3471 3573 3475
rect 3577 3471 3581 3475
rect 3585 3471 3589 3475
rect 3598 3471 3602 3475
rect 3606 3471 3610 3475
rect 3614 3471 3618 3475
rect 3913 3478 3917 3482
rect 3928 3478 3932 3482
rect 2396 3427 2400 3431
rect 2404 3427 2408 3431
rect 2420 3427 2424 3431
rect 2428 3427 2432 3431
rect 3198 3432 3202 3436
rect 3198 3423 3202 3428
rect 3341 3427 3345 3431
rect 3349 3427 3353 3431
rect 3365 3427 3369 3431
rect 3373 3427 3377 3431
rect 4143 3432 4147 3436
rect 4143 3423 4147 3428
rect 2416 3414 2420 3418
rect 2424 3414 2428 3418
rect 3361 3414 3365 3418
rect 3369 3414 3373 3418
rect 2412 3403 2416 3407
rect 3357 3403 3361 3407
rect 2412 3395 2416 3399
rect 2396 3391 2400 3395
rect 2404 3391 2408 3395
rect 2420 3391 2424 3395
rect 2428 3391 2432 3395
rect 3357 3395 3361 3399
rect 3341 3391 3345 3395
rect 3349 3391 3353 3395
rect 3365 3391 3369 3395
rect 3373 3391 3377 3395
rect 3064 3359 3068 3363
rect 3077 3359 3081 3363
rect 3085 3359 3089 3363
rect 3093 3359 3097 3363
rect 3101 3359 3105 3363
rect 3114 3359 3118 3363
rect 3127 3359 3131 3363
rect 3135 3359 3139 3363
rect 3143 3359 3147 3363
rect 3151 3359 3155 3363
rect 3159 3359 3163 3363
rect 3172 3359 3176 3363
rect 3180 3359 3184 3363
rect 3188 3359 3192 3363
rect 4009 3359 4013 3363
rect 4022 3359 4026 3363
rect 4030 3359 4034 3363
rect 4038 3359 4042 3363
rect 4046 3359 4050 3363
rect 4059 3359 4063 3363
rect 4072 3359 4076 3363
rect 4080 3359 4084 3363
rect 4088 3359 4092 3363
rect 4096 3359 4100 3363
rect 4104 3359 4108 3363
rect 4117 3359 4121 3363
rect 4125 3359 4129 3363
rect 4133 3359 4137 3363
rect 2281 3329 2285 3333
rect 2294 3329 2298 3333
rect 2302 3329 2306 3333
rect 2310 3329 2314 3333
rect 2318 3329 2322 3333
rect 2331 3329 2335 3333
rect 2344 3329 2348 3333
rect 2352 3329 2356 3333
rect 2360 3329 2364 3333
rect 2368 3329 2372 3333
rect 2376 3329 2380 3333
rect 2389 3329 2393 3333
rect 2397 3329 2401 3333
rect 2405 3329 2409 3333
rect 2413 3329 2417 3333
rect 2426 3329 2430 3333
rect 2434 3329 2438 3333
rect 2442 3329 2446 3333
rect 2450 3329 2454 3333
rect 2463 3329 2467 3333
rect 2476 3329 2480 3333
rect 2484 3329 2488 3333
rect 2492 3329 2496 3333
rect 2500 3329 2504 3333
rect 2508 3329 2512 3333
rect 2521 3329 2525 3333
rect 2529 3329 2533 3333
rect 2537 3329 2541 3333
rect 2545 3329 2549 3333
rect 2558 3329 2562 3333
rect 2566 3329 2570 3333
rect 2574 3329 2578 3333
rect 2582 3329 2586 3333
rect 2595 3329 2599 3333
rect 2608 3329 2612 3333
rect 2616 3329 2620 3333
rect 2624 3329 2628 3333
rect 2632 3329 2636 3333
rect 2640 3329 2644 3333
rect 2653 3329 2657 3333
rect 2661 3329 2665 3333
rect 2669 3329 2673 3333
rect 3226 3329 3230 3333
rect 3239 3329 3243 3333
rect 3247 3329 3251 3333
rect 3255 3329 3259 3333
rect 3263 3329 3267 3333
rect 3276 3329 3280 3333
rect 3289 3329 3293 3333
rect 3297 3329 3301 3333
rect 3305 3329 3309 3333
rect 3313 3329 3317 3333
rect 3321 3329 3325 3333
rect 3334 3329 3338 3333
rect 3342 3329 3346 3333
rect 3350 3329 3354 3333
rect 3358 3329 3362 3333
rect 3371 3329 3375 3333
rect 3379 3329 3383 3333
rect 3387 3329 3391 3333
rect 3395 3329 3399 3333
rect 3408 3329 3412 3333
rect 3421 3329 3425 3333
rect 3429 3329 3433 3333
rect 3437 3329 3441 3333
rect 3445 3329 3449 3333
rect 3453 3329 3457 3333
rect 3466 3329 3470 3333
rect 3474 3329 3478 3333
rect 3482 3329 3486 3333
rect 3490 3329 3494 3333
rect 3503 3329 3507 3333
rect 3511 3329 3515 3333
rect 3519 3329 3523 3333
rect 3527 3329 3531 3333
rect 3540 3329 3544 3333
rect 3553 3329 3557 3333
rect 3561 3329 3565 3333
rect 3569 3329 3573 3333
rect 3577 3329 3581 3333
rect 3585 3329 3589 3333
rect 3598 3329 3602 3333
rect 3606 3329 3610 3333
rect 3614 3329 3618 3333
rect 3210 3286 3214 3290
rect 3210 3278 3214 3282
rect 4155 3286 4159 3290
rect 4155 3278 4159 3282
rect 3064 3273 3068 3277
rect 3077 3273 3081 3277
rect 3085 3273 3089 3277
rect 3093 3273 3097 3277
rect 3101 3273 3105 3277
rect 3114 3273 3118 3277
rect 3127 3273 3131 3277
rect 3135 3273 3139 3277
rect 3143 3273 3147 3277
rect 3151 3273 3155 3277
rect 3159 3273 3163 3277
rect 3172 3273 3176 3277
rect 3180 3273 3184 3277
rect 3188 3273 3192 3277
rect 4009 3273 4013 3277
rect 4022 3273 4026 3277
rect 4030 3273 4034 3277
rect 4038 3273 4042 3277
rect 4046 3273 4050 3277
rect 4059 3273 4063 3277
rect 4072 3273 4076 3277
rect 4080 3273 4084 3277
rect 4088 3273 4092 3277
rect 4096 3273 4100 3277
rect 4104 3273 4108 3277
rect 4117 3273 4121 3277
rect 4125 3273 4129 3277
rect 4133 3273 4137 3277
rect 2281 3243 2285 3247
rect 2294 3243 2298 3247
rect 2302 3243 2306 3247
rect 2310 3243 2314 3247
rect 2318 3243 2322 3247
rect 2331 3243 2335 3247
rect 2344 3243 2348 3247
rect 2352 3243 2356 3247
rect 2360 3243 2364 3247
rect 2368 3243 2372 3247
rect 2376 3243 2380 3247
rect 2389 3243 2393 3247
rect 2397 3243 2401 3247
rect 2405 3243 2409 3247
rect 2413 3243 2417 3247
rect 2426 3243 2430 3247
rect 2434 3243 2438 3247
rect 2442 3243 2446 3247
rect 2450 3243 2454 3247
rect 2463 3243 2467 3247
rect 2476 3243 2480 3247
rect 2484 3243 2488 3247
rect 2492 3243 2496 3247
rect 2500 3243 2504 3247
rect 2508 3243 2512 3247
rect 2521 3243 2525 3247
rect 2529 3243 2533 3247
rect 2537 3243 2541 3247
rect 2545 3243 2549 3247
rect 2558 3243 2562 3247
rect 2566 3243 2570 3247
rect 2574 3243 2578 3247
rect 2582 3243 2586 3247
rect 2595 3243 2599 3247
rect 2608 3243 2612 3247
rect 2616 3243 2620 3247
rect 2624 3243 2628 3247
rect 2632 3243 2636 3247
rect 2640 3243 2644 3247
rect 2653 3243 2657 3247
rect 2661 3243 2665 3247
rect 2669 3243 2673 3247
rect 3226 3243 3230 3247
rect 3239 3243 3243 3247
rect 3247 3243 3251 3247
rect 3255 3243 3259 3247
rect 3263 3243 3267 3247
rect 3276 3243 3280 3247
rect 3289 3243 3293 3247
rect 3297 3243 3301 3247
rect 3305 3243 3309 3247
rect 3313 3243 3317 3247
rect 3321 3243 3325 3247
rect 3334 3243 3338 3247
rect 3342 3243 3346 3247
rect 3350 3243 3354 3247
rect 3358 3243 3362 3247
rect 3371 3243 3375 3247
rect 3379 3243 3383 3247
rect 3387 3243 3391 3247
rect 3395 3243 3399 3247
rect 3408 3243 3412 3247
rect 3421 3243 3425 3247
rect 3429 3243 3433 3247
rect 3437 3243 3441 3247
rect 3445 3243 3449 3247
rect 3453 3243 3457 3247
rect 3466 3243 3470 3247
rect 3474 3243 3478 3247
rect 3482 3243 3486 3247
rect 3490 3243 3494 3247
rect 3503 3243 3507 3247
rect 3511 3243 3515 3247
rect 3519 3243 3523 3247
rect 3527 3243 3531 3247
rect 3540 3243 3544 3247
rect 3553 3243 3557 3247
rect 3561 3243 3565 3247
rect 3569 3243 3573 3247
rect 3577 3243 3581 3247
rect 3585 3243 3589 3247
rect 3598 3243 3602 3247
rect 3606 3243 3610 3247
rect 3614 3243 3618 3247
rect 2513 3199 2517 3203
rect 2521 3199 2525 3203
rect 2537 3199 2541 3203
rect 2545 3199 2549 3203
rect 3458 3199 3462 3203
rect 3466 3199 3470 3203
rect 3482 3199 3486 3203
rect 3490 3199 3494 3203
rect 2533 3188 2537 3192
rect 2541 3188 2545 3192
rect 3478 3188 3482 3192
rect 3486 3188 3490 3192
rect 2529 3177 2533 3181
rect 3474 3177 3478 3181
rect 2529 3169 2533 3173
rect 3474 3169 3478 3173
rect 2513 3165 2517 3169
rect 2521 3165 2525 3169
rect 2537 3165 2541 3169
rect 2545 3165 2549 3169
rect 3458 3165 3462 3169
rect 3466 3165 3470 3169
rect 3482 3165 3486 3169
rect 3490 3165 3494 3169
rect 2281 3103 2285 3107
rect 2294 3103 2298 3107
rect 2302 3103 2306 3107
rect 2310 3103 2314 3107
rect 2318 3103 2322 3107
rect 2331 3103 2335 3107
rect 2344 3103 2348 3107
rect 2352 3103 2356 3107
rect 2360 3103 2364 3107
rect 2368 3103 2372 3107
rect 2376 3103 2380 3107
rect 2389 3103 2393 3107
rect 2397 3103 2401 3107
rect 2405 3103 2409 3107
rect 2413 3103 2417 3107
rect 2426 3103 2430 3107
rect 2434 3103 2438 3107
rect 2442 3103 2446 3107
rect 2450 3103 2454 3107
rect 2463 3103 2467 3107
rect 2476 3103 2480 3107
rect 2484 3103 2488 3107
rect 2492 3103 2496 3107
rect 2500 3103 2504 3107
rect 2508 3103 2512 3107
rect 2521 3103 2525 3107
rect 2529 3103 2533 3107
rect 2537 3103 2541 3107
rect 2545 3103 2549 3107
rect 2558 3103 2562 3107
rect 2566 3103 2570 3107
rect 2574 3103 2578 3107
rect 2582 3103 2586 3107
rect 2595 3103 2599 3107
rect 2608 3103 2612 3107
rect 2616 3103 2620 3107
rect 2624 3103 2628 3107
rect 2632 3103 2636 3107
rect 2640 3103 2644 3107
rect 2653 3103 2657 3107
rect 2661 3103 2665 3107
rect 2669 3103 2673 3107
rect 3226 3103 3230 3107
rect 3239 3103 3243 3107
rect 3247 3103 3251 3107
rect 3255 3103 3259 3107
rect 3263 3103 3267 3107
rect 3276 3103 3280 3107
rect 3289 3103 3293 3107
rect 3297 3103 3301 3107
rect 3305 3103 3309 3107
rect 3313 3103 3317 3107
rect 3321 3103 3325 3107
rect 3334 3103 3338 3107
rect 3342 3103 3346 3107
rect 3350 3103 3354 3107
rect 3358 3103 3362 3107
rect 3371 3103 3375 3107
rect 3379 3103 3383 3107
rect 3387 3103 3391 3107
rect 3395 3103 3399 3107
rect 3408 3103 3412 3107
rect 3421 3103 3425 3107
rect 3429 3103 3433 3107
rect 3437 3103 3441 3107
rect 3445 3103 3449 3107
rect 3453 3103 3457 3107
rect 3466 3103 3470 3107
rect 3474 3103 3478 3107
rect 3482 3103 3486 3107
rect 3490 3103 3494 3107
rect 3503 3103 3507 3107
rect 3511 3103 3515 3107
rect 3519 3103 3523 3107
rect 3527 3103 3531 3107
rect 3540 3103 3544 3107
rect 3553 3103 3557 3107
rect 3561 3103 3565 3107
rect 3569 3103 3573 3107
rect 3577 3103 3581 3107
rect 3585 3103 3589 3107
rect 3598 3103 3602 3107
rect 3606 3103 3610 3107
rect 3614 3103 3618 3107
rect 2765 3024 2769 3028
rect 2778 3024 2782 3028
rect 2786 3024 2790 3028
rect 2794 3024 2798 3028
rect 2802 3024 2806 3028
rect 2815 3024 2819 3028
rect 2828 3024 2832 3028
rect 2836 3024 2840 3028
rect 2844 3024 2848 3028
rect 2852 3024 2856 3028
rect 2860 3024 2864 3028
rect 2873 3024 2877 3028
rect 2881 3024 2885 3028
rect 2889 3024 2893 3028
rect 2897 3024 2901 3028
rect 2910 3024 2914 3028
rect 2918 3024 2922 3028
rect 2926 3024 2930 3028
rect 2934 3024 2938 3028
rect 2947 3024 2951 3028
rect 2960 3024 2964 3028
rect 2968 3024 2972 3028
rect 2976 3024 2980 3028
rect 2984 3024 2988 3028
rect 2992 3024 2996 3028
rect 3005 3024 3009 3028
rect 3013 3024 3017 3028
rect 3021 3024 3025 3028
rect 3029 3024 3033 3028
rect 3042 3024 3046 3028
rect 3050 3024 3054 3028
rect 3058 3024 3062 3028
rect 3066 3024 3070 3028
rect 3079 3024 3083 3028
rect 3092 3024 3096 3028
rect 3100 3024 3104 3028
rect 3108 3024 3112 3028
rect 3116 3024 3120 3028
rect 3124 3024 3128 3028
rect 3137 3024 3141 3028
rect 3145 3024 3149 3028
rect 3153 3024 3157 3028
rect 3161 3024 3165 3028
rect 3174 3024 3178 3028
rect 3182 3024 3186 3028
rect 3190 3024 3194 3028
rect 3198 3024 3202 3028
rect 3211 3024 3215 3028
rect 3224 3024 3228 3028
rect 3232 3024 3236 3028
rect 3240 3024 3244 3028
rect 3248 3024 3252 3028
rect 3256 3024 3260 3028
rect 3269 3024 3273 3028
rect 3277 3024 3281 3028
rect 3285 3024 3289 3028
rect 3710 3024 3714 3028
rect 3723 3024 3727 3028
rect 3731 3024 3735 3028
rect 3739 3024 3743 3028
rect 3747 3024 3751 3028
rect 3760 3024 3764 3028
rect 3773 3024 3777 3028
rect 3781 3024 3785 3028
rect 3789 3024 3793 3028
rect 3797 3024 3801 3028
rect 3805 3024 3809 3028
rect 3818 3024 3822 3028
rect 3826 3024 3830 3028
rect 3834 3024 3838 3028
rect 3842 3024 3846 3028
rect 3855 3024 3859 3028
rect 3863 3024 3867 3028
rect 3871 3024 3875 3028
rect 3879 3024 3883 3028
rect 3892 3024 3896 3028
rect 3905 3024 3909 3028
rect 3913 3024 3917 3028
rect 3921 3024 3925 3028
rect 3929 3024 3933 3028
rect 3937 3024 3941 3028
rect 3950 3024 3954 3028
rect 3958 3024 3962 3028
rect 3966 3024 3970 3028
rect 3974 3024 3978 3028
rect 3987 3024 3991 3028
rect 3995 3024 3999 3028
rect 4003 3024 4007 3028
rect 4011 3024 4015 3028
rect 4024 3024 4028 3028
rect 4037 3024 4041 3028
rect 4045 3024 4049 3028
rect 4053 3024 4057 3028
rect 4061 3024 4065 3028
rect 4069 3024 4073 3028
rect 4082 3024 4086 3028
rect 4090 3024 4094 3028
rect 4098 3024 4102 3028
rect 4106 3024 4110 3028
rect 4119 3024 4123 3028
rect 4127 3024 4131 3028
rect 4135 3024 4139 3028
rect 4143 3024 4147 3028
rect 4156 3024 4160 3028
rect 4169 3024 4173 3028
rect 4177 3024 4181 3028
rect 4185 3024 4189 3028
rect 4193 3024 4197 3028
rect 4201 3024 4205 3028
rect 4214 3024 4218 3028
rect 4222 3024 4226 3028
rect 4230 3024 4234 3028
rect 2413 2991 2417 2995
rect 2426 2991 2430 2995
rect 2434 2991 2438 2995
rect 2442 2991 2446 2995
rect 2450 2991 2454 2995
rect 2463 2991 2467 2995
rect 2476 2991 2480 2995
rect 2484 2991 2488 2995
rect 2492 2991 2496 2995
rect 2500 2991 2504 2995
rect 2508 2991 2512 2995
rect 2521 2991 2525 2995
rect 2529 2991 2533 2995
rect 2537 2991 2541 2995
rect 3358 2991 3362 2995
rect 3371 2991 3375 2995
rect 3379 2991 3383 2995
rect 3387 2991 3391 2995
rect 3395 2991 3399 2995
rect 3408 2991 3412 2995
rect 3421 2991 3425 2995
rect 3429 2991 3433 2995
rect 3437 2991 3441 2995
rect 3445 2991 3449 2995
rect 3453 2991 3457 2995
rect 3466 2991 3470 2995
rect 3474 2991 3478 2995
rect 3482 2991 3486 2995
rect 2537 2954 2541 2958
rect 2545 2954 2549 2958
rect 2944 2958 2948 2962
rect 2952 2958 2956 2962
rect 2968 2954 2972 2958
rect 2983 2954 2987 2958
rect 3025 2958 3029 2962
rect 3033 2958 3037 2962
rect 3049 2954 3053 2958
rect 3064 2954 3068 2958
rect 2998 2950 3002 2954
rect 3006 2950 3010 2954
rect 2420 2945 2424 2949
rect 2428 2945 2432 2949
rect 2770 2945 2774 2949
rect 2778 2945 2782 2949
rect 2786 2945 2790 2949
rect 2794 2945 2798 2949
rect 2802 2945 2806 2949
rect 2810 2945 2814 2949
rect 2821 2945 2825 2949
rect 2838 2945 2842 2949
rect 2855 2945 2859 2949
rect 2864 2945 2868 2949
rect 2877 2945 2881 2949
rect 2885 2945 2889 2949
rect 2893 2945 2897 2949
rect 2910 2945 2914 2949
rect 2920 2945 2924 2949
rect 2928 2945 2932 2949
rect 3079 2950 3083 2954
rect 3087 2950 3091 2954
rect 3482 2954 3486 2958
rect 3490 2954 3494 2958
rect 3889 2958 3893 2962
rect 3897 2958 3901 2962
rect 3913 2954 3917 2958
rect 3928 2954 3932 2958
rect 3970 2958 3974 2962
rect 3978 2958 3982 2962
rect 3994 2954 3998 2958
rect 4009 2954 4013 2958
rect 3943 2950 3947 2954
rect 3951 2950 3955 2954
rect 3365 2945 3369 2949
rect 3373 2945 3377 2949
rect 3715 2945 3719 2949
rect 3723 2945 3727 2949
rect 3731 2945 3735 2949
rect 3739 2945 3743 2949
rect 3747 2945 3751 2949
rect 3755 2945 3759 2949
rect 3766 2945 3770 2949
rect 3783 2945 3787 2949
rect 3800 2945 3804 2949
rect 3809 2945 3813 2949
rect 3822 2945 3826 2949
rect 3830 2945 3834 2949
rect 3838 2945 3842 2949
rect 3855 2945 3859 2949
rect 3865 2945 3869 2949
rect 3873 2945 3877 2949
rect 4024 2950 4028 2954
rect 4032 2950 4036 2954
rect 2770 2899 2774 2903
rect 2778 2899 2782 2903
rect 2786 2899 2790 2903
rect 2794 2899 2798 2903
rect 2802 2899 2806 2903
rect 2810 2899 2814 2903
rect 2821 2899 2825 2903
rect 2838 2899 2842 2903
rect 2855 2899 2859 2903
rect 2864 2899 2868 2903
rect 2877 2899 2881 2903
rect 2885 2899 2889 2903
rect 2893 2899 2897 2903
rect 2910 2899 2914 2903
rect 2920 2899 2924 2903
rect 2928 2899 2932 2903
rect 2404 2889 2408 2893
rect 2412 2889 2416 2893
rect 2420 2889 2424 2893
rect 2433 2889 2437 2893
rect 2441 2889 2445 2893
rect 2449 2889 2453 2893
rect 2457 2889 2461 2893
rect 2465 2889 2469 2893
rect 2478 2889 2482 2893
rect 2491 2889 2495 2893
rect 2499 2889 2503 2893
rect 2507 2889 2511 2893
rect 2515 2889 2519 2893
rect 2528 2889 2532 2893
rect 2968 2898 2972 2902
rect 2983 2898 2987 2902
rect 3049 2898 3053 2902
rect 3064 2898 3068 2902
rect 3715 2899 3719 2903
rect 3723 2899 3727 2903
rect 3731 2899 3735 2903
rect 3739 2899 3743 2903
rect 3747 2899 3751 2903
rect 3755 2899 3759 2903
rect 3766 2899 3770 2903
rect 3783 2899 3787 2903
rect 3800 2899 3804 2903
rect 3809 2899 3813 2903
rect 3822 2899 3826 2903
rect 3830 2899 3834 2903
rect 3838 2899 3842 2903
rect 3855 2899 3859 2903
rect 3865 2899 3869 2903
rect 3873 2899 3877 2903
rect 3349 2889 3353 2893
rect 3357 2889 3361 2893
rect 3365 2889 3369 2893
rect 3378 2889 3382 2893
rect 3386 2889 3390 2893
rect 3394 2889 3398 2893
rect 3402 2889 3406 2893
rect 3410 2889 3414 2893
rect 3423 2889 3427 2893
rect 3436 2889 3440 2893
rect 3444 2889 3448 2893
rect 3452 2889 3456 2893
rect 3460 2889 3464 2893
rect 3473 2889 3477 2893
rect 3913 2898 3917 2902
rect 3928 2898 3932 2902
rect 3994 2898 3998 2902
rect 4009 2898 4013 2902
rect 2968 2822 2972 2826
rect 2983 2822 2987 2826
rect 3049 2826 3053 2830
rect 3057 2826 3061 2830
rect 3073 2822 3077 2826
rect 3088 2822 3092 2826
rect 2998 2818 3002 2822
rect 3006 2818 3010 2822
rect 2770 2813 2774 2817
rect 2778 2813 2782 2817
rect 2786 2813 2790 2817
rect 2794 2813 2798 2817
rect 2802 2813 2806 2817
rect 2810 2813 2814 2817
rect 2821 2813 2825 2817
rect 2838 2813 2842 2817
rect 2855 2813 2859 2817
rect 2864 2813 2868 2817
rect 2877 2813 2881 2817
rect 2885 2813 2889 2817
rect 2893 2813 2897 2817
rect 2910 2813 2914 2817
rect 2920 2813 2924 2817
rect 2928 2813 2932 2817
rect 3103 2818 3107 2822
rect 3111 2818 3115 2822
rect 3913 2822 3917 2826
rect 3928 2822 3932 2826
rect 3994 2826 3998 2830
rect 4002 2826 4006 2830
rect 4018 2822 4022 2826
rect 4033 2822 4037 2826
rect 3943 2818 3947 2822
rect 3951 2818 3955 2822
rect 3715 2813 3719 2817
rect 3723 2813 3727 2817
rect 3731 2813 3735 2817
rect 3739 2813 3743 2817
rect 3747 2813 3751 2817
rect 3755 2813 3759 2817
rect 3766 2813 3770 2817
rect 3783 2813 3787 2817
rect 3800 2813 3804 2817
rect 3809 2813 3813 2817
rect 3822 2813 3826 2817
rect 3830 2813 3834 2817
rect 3838 2813 3842 2817
rect 3855 2813 3859 2817
rect 3865 2813 3869 2817
rect 3873 2813 3877 2817
rect 4048 2818 4052 2822
rect 4056 2818 4060 2822
rect 2770 2767 2774 2771
rect 2778 2767 2782 2771
rect 2786 2767 2790 2771
rect 2794 2767 2798 2771
rect 2802 2767 2806 2771
rect 2810 2767 2814 2771
rect 2821 2767 2825 2771
rect 2838 2767 2842 2771
rect 2855 2767 2859 2771
rect 2864 2767 2868 2771
rect 2877 2767 2881 2771
rect 2885 2767 2889 2771
rect 2893 2767 2897 2771
rect 2910 2767 2914 2771
rect 2920 2767 2924 2771
rect 2928 2767 2932 2771
rect 2968 2767 2972 2771
rect 2983 2767 2987 2771
rect 3073 2767 3077 2771
rect 3088 2767 3092 2771
rect 3715 2767 3719 2771
rect 3723 2767 3727 2771
rect 3731 2767 3735 2771
rect 3739 2767 3743 2771
rect 3747 2767 3751 2771
rect 3755 2767 3759 2771
rect 3766 2767 3770 2771
rect 3783 2767 3787 2771
rect 3800 2767 3804 2771
rect 3809 2767 3813 2771
rect 3822 2767 3826 2771
rect 3830 2767 3834 2771
rect 3838 2767 3842 2771
rect 3855 2767 3859 2771
rect 3865 2767 3869 2771
rect 3873 2767 3877 2771
rect 3913 2767 3917 2771
rect 3928 2767 3932 2771
rect 4018 2767 4022 2771
rect 4033 2767 4037 2771
rect 2968 2690 2972 2694
rect 2983 2690 2987 2694
rect 3025 2694 3029 2698
rect 3033 2694 3037 2698
rect 3049 2690 3053 2694
rect 3064 2690 3068 2694
rect 3115 2694 3119 2698
rect 3123 2694 3127 2698
rect 3139 2690 3143 2694
rect 3154 2690 3158 2694
rect 2998 2686 3002 2690
rect 3006 2686 3010 2690
rect 2770 2681 2774 2685
rect 2778 2681 2782 2685
rect 2786 2681 2790 2685
rect 2794 2681 2798 2685
rect 2802 2681 2806 2685
rect 2810 2681 2814 2685
rect 2821 2681 2825 2685
rect 2838 2681 2842 2685
rect 2855 2681 2859 2685
rect 2864 2681 2868 2685
rect 2877 2681 2881 2685
rect 2885 2681 2889 2685
rect 2893 2681 2897 2685
rect 2910 2681 2914 2685
rect 2920 2681 2924 2685
rect 2928 2681 2932 2685
rect 3079 2686 3083 2690
rect 3087 2686 3091 2690
rect 3169 2686 3173 2690
rect 3177 2686 3181 2690
rect 3913 2690 3917 2694
rect 3928 2690 3932 2694
rect 3970 2694 3974 2698
rect 3978 2694 3982 2698
rect 3994 2690 3998 2694
rect 4009 2690 4013 2694
rect 4060 2694 4064 2698
rect 4068 2694 4072 2698
rect 4084 2690 4088 2694
rect 4099 2690 4103 2694
rect 3943 2686 3947 2690
rect 3951 2686 3955 2690
rect 3715 2681 3719 2685
rect 3723 2681 3727 2685
rect 3731 2681 3735 2685
rect 3739 2681 3743 2685
rect 3747 2681 3751 2685
rect 3755 2681 3759 2685
rect 3766 2681 3770 2685
rect 3783 2681 3787 2685
rect 3800 2681 3804 2685
rect 3809 2681 3813 2685
rect 3822 2681 3826 2685
rect 3830 2681 3834 2685
rect 3838 2681 3842 2685
rect 3855 2681 3859 2685
rect 3865 2681 3869 2685
rect 3873 2681 3877 2685
rect 4024 2686 4028 2690
rect 4032 2686 4036 2690
rect 4114 2686 4118 2690
rect 4122 2686 4126 2690
rect 2770 2635 2774 2639
rect 2778 2635 2782 2639
rect 2786 2635 2790 2639
rect 2794 2635 2798 2639
rect 2802 2635 2806 2639
rect 2810 2635 2814 2639
rect 2821 2635 2825 2639
rect 2838 2635 2842 2639
rect 2855 2635 2859 2639
rect 2864 2635 2868 2639
rect 2877 2635 2881 2639
rect 2885 2635 2889 2639
rect 2893 2635 2897 2639
rect 2910 2635 2914 2639
rect 2920 2635 2924 2639
rect 2928 2635 2932 2639
rect 2968 2632 2972 2636
rect 2983 2632 2987 2636
rect 3049 2632 3053 2636
rect 3064 2632 3068 2636
rect 3139 2632 3143 2636
rect 3154 2632 3158 2636
rect 3715 2635 3719 2639
rect 3723 2635 3727 2639
rect 3731 2635 3735 2639
rect 3739 2635 3743 2639
rect 3747 2635 3751 2639
rect 3755 2635 3759 2639
rect 3766 2635 3770 2639
rect 3783 2635 3787 2639
rect 3800 2635 3804 2639
rect 3809 2635 3813 2639
rect 3822 2635 3826 2639
rect 3830 2635 3834 2639
rect 3838 2635 3842 2639
rect 3855 2635 3859 2639
rect 3865 2635 3869 2639
rect 3873 2635 3877 2639
rect 3913 2632 3917 2636
rect 3928 2632 3932 2636
rect 3994 2632 3998 2636
rect 4009 2632 4013 2636
rect 4084 2632 4088 2636
rect 4099 2632 4103 2636
rect 2968 2558 2972 2562
rect 2983 2558 2987 2562
rect 2998 2554 3002 2558
rect 3006 2554 3010 2558
rect 2770 2549 2774 2553
rect 2778 2549 2782 2553
rect 2786 2549 2790 2553
rect 2794 2549 2798 2553
rect 2802 2549 2806 2553
rect 2810 2549 2814 2553
rect 2821 2549 2825 2553
rect 2838 2549 2842 2553
rect 2855 2549 2859 2553
rect 2864 2549 2868 2553
rect 2877 2549 2881 2553
rect 2885 2549 2889 2553
rect 2893 2549 2897 2553
rect 2910 2549 2914 2553
rect 2920 2549 2924 2553
rect 2928 2549 2932 2553
rect 3913 2558 3917 2562
rect 3928 2558 3932 2562
rect 3943 2554 3947 2558
rect 3951 2554 3955 2558
rect 3715 2549 3719 2553
rect 3723 2549 3727 2553
rect 3731 2549 3735 2553
rect 3739 2549 3743 2553
rect 3747 2549 3751 2553
rect 3755 2549 3759 2553
rect 3766 2549 3770 2553
rect 3783 2549 3787 2553
rect 3800 2549 3804 2553
rect 3809 2549 3813 2553
rect 3822 2549 3826 2553
rect 3830 2549 3834 2553
rect 3838 2549 3842 2553
rect 3855 2549 3859 2553
rect 3865 2549 3869 2553
rect 3873 2549 3877 2553
rect 2770 2503 2774 2507
rect 2778 2503 2782 2507
rect 2786 2503 2790 2507
rect 2794 2503 2798 2507
rect 2802 2503 2806 2507
rect 2810 2503 2814 2507
rect 2821 2503 2825 2507
rect 2838 2503 2842 2507
rect 2855 2503 2859 2507
rect 2864 2503 2868 2507
rect 2877 2503 2881 2507
rect 2885 2503 2889 2507
rect 2893 2503 2897 2507
rect 2910 2503 2914 2507
rect 2920 2503 2924 2507
rect 2928 2503 2932 2507
rect 3004 2503 3008 2507
rect 3012 2503 3016 2507
rect 3022 2503 3026 2507
rect 3030 2503 3034 2507
rect 3039 2503 3043 2507
rect 3047 2503 3051 2507
rect 3055 2503 3059 2507
rect 3063 2503 3067 2507
rect 3071 2503 3075 2507
rect 3082 2503 3086 2507
rect 3099 2503 3103 2507
rect 3116 2503 3120 2507
rect 3125 2503 3129 2507
rect 3138 2503 3142 2507
rect 3146 2503 3150 2507
rect 3154 2503 3158 2507
rect 3171 2503 3175 2507
rect 3181 2503 3185 2507
rect 3189 2503 3193 2507
rect 2281 2489 2285 2493
rect 2294 2489 2298 2493
rect 2302 2489 2306 2493
rect 2310 2489 2314 2493
rect 2318 2489 2322 2493
rect 2331 2489 2335 2493
rect 2344 2489 2348 2493
rect 2352 2489 2356 2493
rect 2360 2489 2364 2493
rect 2368 2489 2372 2493
rect 2376 2489 2380 2493
rect 2389 2489 2393 2493
rect 2397 2489 2401 2493
rect 2405 2489 2409 2493
rect 2413 2489 2417 2493
rect 2426 2489 2430 2493
rect 2434 2489 2438 2493
rect 2442 2489 2446 2493
rect 2450 2489 2454 2493
rect 2463 2489 2467 2493
rect 2476 2489 2480 2493
rect 2484 2489 2488 2493
rect 2492 2489 2496 2493
rect 2500 2489 2504 2493
rect 2508 2489 2512 2493
rect 2521 2489 2525 2493
rect 2529 2489 2533 2493
rect 2537 2489 2541 2493
rect 2545 2489 2549 2493
rect 2558 2489 2562 2493
rect 2566 2489 2570 2493
rect 2574 2489 2578 2493
rect 2582 2489 2586 2493
rect 2595 2489 2599 2493
rect 2608 2489 2612 2493
rect 2616 2489 2620 2493
rect 2624 2489 2628 2493
rect 2632 2489 2636 2493
rect 2640 2489 2644 2493
rect 2653 2489 2657 2493
rect 2661 2489 2665 2493
rect 2669 2489 2673 2493
rect 2968 2496 2972 2500
rect 2983 2496 2987 2500
rect 3715 2503 3719 2507
rect 3723 2503 3727 2507
rect 3731 2503 3735 2507
rect 3739 2503 3743 2507
rect 3747 2503 3751 2507
rect 3755 2503 3759 2507
rect 3766 2503 3770 2507
rect 3783 2503 3787 2507
rect 3800 2503 3804 2507
rect 3809 2503 3813 2507
rect 3822 2503 3826 2507
rect 3830 2503 3834 2507
rect 3838 2503 3842 2507
rect 3855 2503 3859 2507
rect 3865 2503 3869 2507
rect 3873 2503 3877 2507
rect 3949 2503 3953 2507
rect 3957 2503 3961 2507
rect 3967 2503 3971 2507
rect 3975 2503 3979 2507
rect 3984 2503 3988 2507
rect 3992 2503 3996 2507
rect 4000 2503 4004 2507
rect 4008 2503 4012 2507
rect 4016 2503 4020 2507
rect 4027 2503 4031 2507
rect 4044 2503 4048 2507
rect 4061 2503 4065 2507
rect 4070 2503 4074 2507
rect 4083 2503 4087 2507
rect 4091 2503 4095 2507
rect 4099 2503 4103 2507
rect 4116 2503 4120 2507
rect 4126 2503 4130 2507
rect 4134 2503 4138 2507
rect 3226 2489 3230 2493
rect 3239 2489 3243 2493
rect 3247 2489 3251 2493
rect 3255 2489 3259 2493
rect 3263 2489 3267 2493
rect 3276 2489 3280 2493
rect 3289 2489 3293 2493
rect 3297 2489 3301 2493
rect 3305 2489 3309 2493
rect 3313 2489 3317 2493
rect 3321 2489 3325 2493
rect 3334 2489 3338 2493
rect 3342 2489 3346 2493
rect 3350 2489 3354 2493
rect 3358 2489 3362 2493
rect 3371 2489 3375 2493
rect 3379 2489 3383 2493
rect 3387 2489 3391 2493
rect 3395 2489 3399 2493
rect 3408 2489 3412 2493
rect 3421 2489 3425 2493
rect 3429 2489 3433 2493
rect 3437 2489 3441 2493
rect 3445 2489 3449 2493
rect 3453 2489 3457 2493
rect 3466 2489 3470 2493
rect 3474 2489 3478 2493
rect 3482 2489 3486 2493
rect 3490 2489 3494 2493
rect 3503 2489 3507 2493
rect 3511 2489 3515 2493
rect 3519 2489 3523 2493
rect 3527 2489 3531 2493
rect 3540 2489 3544 2493
rect 3553 2489 3557 2493
rect 3561 2489 3565 2493
rect 3569 2489 3573 2493
rect 3577 2489 3581 2493
rect 3585 2489 3589 2493
rect 3598 2489 3602 2493
rect 3606 2489 3610 2493
rect 3614 2489 3618 2493
rect 3913 2496 3917 2500
rect 3928 2496 3932 2500
rect 2396 2445 2400 2449
rect 2404 2445 2408 2449
rect 2420 2445 2424 2449
rect 2428 2445 2432 2449
rect 3198 2450 3202 2454
rect 3198 2442 3202 2446
rect 3341 2445 3345 2449
rect 3349 2445 3353 2449
rect 3365 2445 3369 2449
rect 3373 2445 3377 2449
rect 4143 2450 4147 2454
rect 4143 2442 4147 2446
rect 2416 2432 2420 2436
rect 2424 2432 2428 2436
rect 3361 2432 3365 2436
rect 3369 2432 3373 2436
rect 2412 2421 2416 2425
rect 3357 2421 3361 2425
rect 2412 2413 2416 2417
rect 2396 2409 2400 2413
rect 2404 2409 2408 2413
rect 2420 2409 2424 2413
rect 2428 2409 2432 2413
rect 3357 2413 3361 2417
rect 3341 2409 3345 2413
rect 3349 2409 3353 2413
rect 3365 2409 3369 2413
rect 3373 2409 3377 2413
rect 3064 2377 3068 2381
rect 3077 2377 3081 2381
rect 3085 2377 3089 2381
rect 3093 2377 3097 2381
rect 3101 2377 3105 2381
rect 3114 2377 3118 2381
rect 3127 2377 3131 2381
rect 3135 2377 3139 2381
rect 3143 2377 3147 2381
rect 3151 2377 3155 2381
rect 3159 2377 3163 2381
rect 3172 2377 3176 2381
rect 3180 2377 3184 2381
rect 3188 2377 3192 2381
rect 4009 2377 4013 2381
rect 4022 2377 4026 2381
rect 4030 2377 4034 2381
rect 4038 2377 4042 2381
rect 4046 2377 4050 2381
rect 4059 2377 4063 2381
rect 4072 2377 4076 2381
rect 4080 2377 4084 2381
rect 4088 2377 4092 2381
rect 4096 2377 4100 2381
rect 4104 2377 4108 2381
rect 4117 2377 4121 2381
rect 4125 2377 4129 2381
rect 4133 2377 4137 2381
rect 2281 2347 2285 2351
rect 2294 2347 2298 2351
rect 2302 2347 2306 2351
rect 2310 2347 2314 2351
rect 2318 2347 2322 2351
rect 2331 2347 2335 2351
rect 2344 2347 2348 2351
rect 2352 2347 2356 2351
rect 2360 2347 2364 2351
rect 2368 2347 2372 2351
rect 2376 2347 2380 2351
rect 2389 2347 2393 2351
rect 2397 2347 2401 2351
rect 2405 2347 2409 2351
rect 2413 2347 2417 2351
rect 2426 2347 2430 2351
rect 2434 2347 2438 2351
rect 2442 2347 2446 2351
rect 2450 2347 2454 2351
rect 2463 2347 2467 2351
rect 2476 2347 2480 2351
rect 2484 2347 2488 2351
rect 2492 2347 2496 2351
rect 2500 2347 2504 2351
rect 2508 2347 2512 2351
rect 2521 2347 2525 2351
rect 2529 2347 2533 2351
rect 2537 2347 2541 2351
rect 2545 2347 2549 2351
rect 2558 2347 2562 2351
rect 2566 2347 2570 2351
rect 2574 2347 2578 2351
rect 2582 2347 2586 2351
rect 2595 2347 2599 2351
rect 2608 2347 2612 2351
rect 2616 2347 2620 2351
rect 2624 2347 2628 2351
rect 2632 2347 2636 2351
rect 2640 2347 2644 2351
rect 2653 2347 2657 2351
rect 2661 2347 2665 2351
rect 2669 2347 2673 2351
rect 3226 2347 3230 2351
rect 3239 2347 3243 2351
rect 3247 2347 3251 2351
rect 3255 2347 3259 2351
rect 3263 2347 3267 2351
rect 3276 2347 3280 2351
rect 3289 2347 3293 2351
rect 3297 2347 3301 2351
rect 3305 2347 3309 2351
rect 3313 2347 3317 2351
rect 3321 2347 3325 2351
rect 3334 2347 3338 2351
rect 3342 2347 3346 2351
rect 3350 2347 3354 2351
rect 3358 2347 3362 2351
rect 3371 2347 3375 2351
rect 3379 2347 3383 2351
rect 3387 2347 3391 2351
rect 3395 2347 3399 2351
rect 3408 2347 3412 2351
rect 3421 2347 3425 2351
rect 3429 2347 3433 2351
rect 3437 2347 3441 2351
rect 3445 2347 3449 2351
rect 3453 2347 3457 2351
rect 3466 2347 3470 2351
rect 3474 2347 3478 2351
rect 3482 2347 3486 2351
rect 3490 2347 3494 2351
rect 3503 2347 3507 2351
rect 3511 2347 3515 2351
rect 3519 2347 3523 2351
rect 3527 2347 3531 2351
rect 3540 2347 3544 2351
rect 3553 2347 3557 2351
rect 3561 2347 3565 2351
rect 3569 2347 3573 2351
rect 3577 2347 3581 2351
rect 3585 2347 3589 2351
rect 3598 2347 3602 2351
rect 3606 2347 3610 2351
rect 3614 2347 3618 2351
rect 3210 2304 3214 2308
rect 3210 2296 3214 2300
rect 4155 2304 4159 2308
rect 4155 2296 4159 2300
rect 3064 2291 3068 2295
rect 3077 2291 3081 2295
rect 3085 2291 3089 2295
rect 3093 2291 3097 2295
rect 3101 2291 3105 2295
rect 3114 2291 3118 2295
rect 3127 2291 3131 2295
rect 3135 2291 3139 2295
rect 3143 2291 3147 2295
rect 3151 2291 3155 2295
rect 3159 2291 3163 2295
rect 3172 2291 3176 2295
rect 3180 2291 3184 2295
rect 3188 2291 3192 2295
rect 4009 2291 4013 2295
rect 4022 2291 4026 2295
rect 4030 2291 4034 2295
rect 4038 2291 4042 2295
rect 4046 2291 4050 2295
rect 4059 2291 4063 2295
rect 4072 2291 4076 2295
rect 4080 2291 4084 2295
rect 4088 2291 4092 2295
rect 4096 2291 4100 2295
rect 4104 2291 4108 2295
rect 4117 2291 4121 2295
rect 4125 2291 4129 2295
rect 4133 2291 4137 2295
rect 2281 2261 2285 2265
rect 2294 2261 2298 2265
rect 2302 2261 2306 2265
rect 2310 2261 2314 2265
rect 2318 2261 2322 2265
rect 2331 2261 2335 2265
rect 2344 2261 2348 2265
rect 2352 2261 2356 2265
rect 2360 2261 2364 2265
rect 2368 2261 2372 2265
rect 2376 2261 2380 2265
rect 2389 2261 2393 2265
rect 2397 2261 2401 2265
rect 2405 2261 2409 2265
rect 2413 2261 2417 2265
rect 2426 2261 2430 2265
rect 2434 2261 2438 2265
rect 2442 2261 2446 2265
rect 2450 2261 2454 2265
rect 2463 2261 2467 2265
rect 2476 2261 2480 2265
rect 2484 2261 2488 2265
rect 2492 2261 2496 2265
rect 2500 2261 2504 2265
rect 2508 2261 2512 2265
rect 2521 2261 2525 2265
rect 2529 2261 2533 2265
rect 2537 2261 2541 2265
rect 2545 2261 2549 2265
rect 2558 2261 2562 2265
rect 2566 2261 2570 2265
rect 2574 2261 2578 2265
rect 2582 2261 2586 2265
rect 2595 2261 2599 2265
rect 2608 2261 2612 2265
rect 2616 2261 2620 2265
rect 2624 2261 2628 2265
rect 2632 2261 2636 2265
rect 2640 2261 2644 2265
rect 2653 2261 2657 2265
rect 2661 2261 2665 2265
rect 2669 2261 2673 2265
rect 3226 2261 3230 2265
rect 3239 2261 3243 2265
rect 3247 2261 3251 2265
rect 3255 2261 3259 2265
rect 3263 2261 3267 2265
rect 3276 2261 3280 2265
rect 3289 2261 3293 2265
rect 3297 2261 3301 2265
rect 3305 2261 3309 2265
rect 3313 2261 3317 2265
rect 3321 2261 3325 2265
rect 3334 2261 3338 2265
rect 3342 2261 3346 2265
rect 3350 2261 3354 2265
rect 3358 2261 3362 2265
rect 3371 2261 3375 2265
rect 3379 2261 3383 2265
rect 3387 2261 3391 2265
rect 3395 2261 3399 2265
rect 3408 2261 3412 2265
rect 3421 2261 3425 2265
rect 3429 2261 3433 2265
rect 3437 2261 3441 2265
rect 3445 2261 3449 2265
rect 3453 2261 3457 2265
rect 3466 2261 3470 2265
rect 3474 2261 3478 2265
rect 3482 2261 3486 2265
rect 3490 2261 3494 2265
rect 3503 2261 3507 2265
rect 3511 2261 3515 2265
rect 3519 2261 3523 2265
rect 3527 2261 3531 2265
rect 3540 2261 3544 2265
rect 3553 2261 3557 2265
rect 3561 2261 3565 2265
rect 3569 2261 3573 2265
rect 3577 2261 3581 2265
rect 3585 2261 3589 2265
rect 3598 2261 3602 2265
rect 3606 2261 3610 2265
rect 3614 2261 3618 2265
rect 2513 2217 2517 2221
rect 2521 2217 2525 2221
rect 2537 2217 2541 2221
rect 2545 2217 2549 2221
rect 3458 2217 3462 2221
rect 3466 2217 3470 2221
rect 3482 2217 3486 2221
rect 3490 2217 3494 2221
rect 2533 2206 2537 2210
rect 2541 2206 2545 2210
rect 3478 2206 3482 2210
rect 3486 2206 3490 2210
rect 2529 2195 2533 2199
rect 3474 2195 3478 2199
rect 2529 2187 2533 2191
rect 3474 2187 3478 2191
rect 2513 2183 2517 2187
rect 2521 2183 2525 2187
rect 2537 2183 2541 2187
rect 2545 2183 2549 2187
rect 3458 2183 3462 2187
rect 3466 2183 3470 2187
rect 3482 2183 3486 2187
rect 3490 2183 3494 2187
rect 2281 2121 2285 2125
rect 2294 2121 2298 2125
rect 2302 2121 2306 2125
rect 2310 2121 2314 2125
rect 2318 2121 2322 2125
rect 2331 2121 2335 2125
rect 2344 2121 2348 2125
rect 2352 2121 2356 2125
rect 2360 2121 2364 2125
rect 2368 2121 2372 2125
rect 2376 2121 2380 2125
rect 2389 2121 2393 2125
rect 2397 2121 2401 2125
rect 2405 2121 2409 2125
rect 2413 2121 2417 2125
rect 2426 2121 2430 2125
rect 2434 2121 2438 2125
rect 2442 2121 2446 2125
rect 2450 2121 2454 2125
rect 2463 2121 2467 2125
rect 2476 2121 2480 2125
rect 2484 2121 2488 2125
rect 2492 2121 2496 2125
rect 2500 2121 2504 2125
rect 2508 2121 2512 2125
rect 2521 2121 2525 2125
rect 2529 2121 2533 2125
rect 2537 2121 2541 2125
rect 2545 2121 2549 2125
rect 2558 2121 2562 2125
rect 2566 2121 2570 2125
rect 2574 2121 2578 2125
rect 2582 2121 2586 2125
rect 2595 2121 2599 2125
rect 2608 2121 2612 2125
rect 2616 2121 2620 2125
rect 2624 2121 2628 2125
rect 2632 2121 2636 2125
rect 2640 2121 2644 2125
rect 2653 2121 2657 2125
rect 2661 2121 2665 2125
rect 2669 2121 2673 2125
rect 3226 2121 3230 2125
rect 3239 2121 3243 2125
rect 3247 2121 3251 2125
rect 3255 2121 3259 2125
rect 3263 2121 3267 2125
rect 3276 2121 3280 2125
rect 3289 2121 3293 2125
rect 3297 2121 3301 2125
rect 3305 2121 3309 2125
rect 3313 2121 3317 2125
rect 3321 2121 3325 2125
rect 3334 2121 3338 2125
rect 3342 2121 3346 2125
rect 3350 2121 3354 2125
rect 3358 2121 3362 2125
rect 3371 2121 3375 2125
rect 3379 2121 3383 2125
rect 3387 2121 3391 2125
rect 3395 2121 3399 2125
rect 3408 2121 3412 2125
rect 3421 2121 3425 2125
rect 3429 2121 3433 2125
rect 3437 2121 3441 2125
rect 3445 2121 3449 2125
rect 3453 2121 3457 2125
rect 3466 2121 3470 2125
rect 3474 2121 3478 2125
rect 3482 2121 3486 2125
rect 3490 2121 3494 2125
rect 3503 2121 3507 2125
rect 3511 2121 3515 2125
rect 3519 2121 3523 2125
rect 3527 2121 3531 2125
rect 3540 2121 3544 2125
rect 3553 2121 3557 2125
rect 3561 2121 3565 2125
rect 3569 2121 3573 2125
rect 3577 2121 3581 2125
rect 3585 2121 3589 2125
rect 3598 2121 3602 2125
rect 3606 2121 3610 2125
rect 3614 2121 3618 2125
<< pdcontact >>
rect 2765 4029 2769 4037
rect 2778 4029 2782 4037
rect 2786 4029 2790 4037
rect 2794 4033 2798 4037
rect 2802 4029 2806 4037
rect 2815 4029 2819 4037
rect 2828 4029 2832 4037
rect 2836 4029 2840 4037
rect 2844 4029 2848 4037
rect 2852 4033 2856 4037
rect 2860 4029 2864 4037
rect 2873 4029 2877 4037
rect 2881 4029 2885 4037
rect 2889 4029 2893 4037
rect 2897 4029 2901 4037
rect 2910 4029 2914 4037
rect 2918 4029 2922 4037
rect 2926 4033 2930 4037
rect 2934 4029 2938 4037
rect 2947 4029 2951 4037
rect 2960 4029 2964 4037
rect 2968 4029 2972 4037
rect 2976 4029 2980 4037
rect 2984 4033 2988 4037
rect 2992 4029 2996 4037
rect 3005 4029 3009 4037
rect 3013 4029 3017 4037
rect 3021 4029 3025 4037
rect 3029 4029 3033 4037
rect 3042 4029 3046 4037
rect 3050 4029 3054 4037
rect 3058 4033 3062 4037
rect 3066 4029 3070 4037
rect 3079 4029 3083 4037
rect 3092 4029 3096 4037
rect 3100 4029 3104 4037
rect 3108 4029 3112 4037
rect 3116 4033 3120 4037
rect 3124 4029 3128 4037
rect 3137 4029 3141 4037
rect 3145 4029 3149 4037
rect 3153 4029 3157 4037
rect 3161 4029 3165 4037
rect 3174 4029 3178 4037
rect 3182 4029 3186 4037
rect 3190 4033 3194 4037
rect 3198 4029 3202 4037
rect 3211 4029 3215 4037
rect 3224 4029 3228 4037
rect 3232 4029 3236 4037
rect 3240 4029 3244 4037
rect 3248 4033 3252 4037
rect 3256 4029 3260 4037
rect 3269 4029 3273 4037
rect 3277 4029 3281 4037
rect 3285 4029 3289 4037
rect 3710 4029 3714 4037
rect 3723 4029 3727 4037
rect 3731 4029 3735 4037
rect 3739 4033 3743 4037
rect 3747 4029 3751 4037
rect 3760 4029 3764 4037
rect 3773 4029 3777 4037
rect 3781 4029 3785 4037
rect 3789 4029 3793 4037
rect 3797 4033 3801 4037
rect 3805 4029 3809 4037
rect 3818 4029 3822 4037
rect 3826 4029 3830 4037
rect 3834 4029 3838 4037
rect 3842 4029 3846 4037
rect 3855 4029 3859 4037
rect 3863 4029 3867 4037
rect 3871 4033 3875 4037
rect 3879 4029 3883 4037
rect 3892 4029 3896 4037
rect 3905 4029 3909 4037
rect 3913 4029 3917 4037
rect 3921 4029 3925 4037
rect 3929 4033 3933 4037
rect 3937 4029 3941 4037
rect 3950 4029 3954 4037
rect 3958 4029 3962 4037
rect 3966 4029 3970 4037
rect 3974 4029 3978 4037
rect 3987 4029 3991 4037
rect 3995 4029 3999 4037
rect 4003 4033 4007 4037
rect 4011 4029 4015 4037
rect 4024 4029 4028 4037
rect 4037 4029 4041 4037
rect 4045 4029 4049 4037
rect 4053 4029 4057 4037
rect 4061 4033 4065 4037
rect 4069 4029 4073 4037
rect 4082 4029 4086 4037
rect 4090 4029 4094 4037
rect 4098 4029 4102 4037
rect 4106 4029 4110 4037
rect 4119 4029 4123 4037
rect 4127 4029 4131 4037
rect 4135 4033 4139 4037
rect 4143 4029 4147 4037
rect 4156 4029 4160 4037
rect 4169 4029 4173 4037
rect 4177 4029 4181 4037
rect 4185 4029 4189 4037
rect 4193 4033 4197 4037
rect 4201 4029 4205 4037
rect 4214 4029 4218 4037
rect 4222 4029 4226 4037
rect 4230 4029 4234 4037
rect 2413 3996 2417 4004
rect 2426 3996 2430 4004
rect 2434 3996 2438 4004
rect 2442 4000 2446 4004
rect 2450 3996 2454 4004
rect 2463 3996 2467 4004
rect 2476 3996 2480 4004
rect 2484 3996 2488 4004
rect 2492 3996 2496 4004
rect 2500 4000 2504 4004
rect 2508 3996 2512 4004
rect 2521 3996 2525 4004
rect 2529 3996 2533 4004
rect 2537 3996 2541 4004
rect 3358 3996 3362 4004
rect 3371 3996 3375 4004
rect 3379 3996 3383 4004
rect 3387 4000 3391 4004
rect 3395 3996 3399 4004
rect 3408 3996 3412 4004
rect 3421 3996 3425 4004
rect 3429 3996 3433 4004
rect 3437 3996 3441 4004
rect 3445 4000 3449 4004
rect 3453 3996 3457 4004
rect 3466 3996 3470 4004
rect 3474 3996 3478 4004
rect 3482 3996 3486 4004
rect 2944 3958 2948 3966
rect 2952 3958 2956 3966
rect 2770 3945 2774 3953
rect 2778 3945 2782 3953
rect 2786 3945 2790 3953
rect 2794 3945 2798 3953
rect 2802 3945 2806 3953
rect 2810 3945 2814 3953
rect 2821 3945 2825 3953
rect 2838 3945 2842 3953
rect 2855 3945 2859 3953
rect 2864 3945 2868 3953
rect 2877 3945 2881 3953
rect 2885 3945 2889 3953
rect 2893 3945 2897 3953
rect 2910 3945 2914 3953
rect 2920 3945 2924 3953
rect 2928 3945 2932 3953
rect 2968 3952 2972 3960
rect 2983 3952 2987 3960
rect 2998 3958 3002 3966
rect 3006 3958 3010 3966
rect 3025 3958 3029 3966
rect 3033 3958 3037 3966
rect 3049 3952 3053 3960
rect 3064 3952 3068 3960
rect 3079 3958 3083 3966
rect 3087 3958 3091 3966
rect 3889 3958 3893 3966
rect 3897 3958 3901 3966
rect 3715 3945 3719 3953
rect 3723 3945 3727 3953
rect 3731 3945 3735 3953
rect 3739 3945 3743 3953
rect 3747 3945 3751 3953
rect 3755 3945 3759 3953
rect 3766 3945 3770 3953
rect 3783 3945 3787 3953
rect 3800 3945 3804 3953
rect 3809 3945 3813 3953
rect 3822 3945 3826 3953
rect 3830 3945 3834 3953
rect 3838 3945 3842 3953
rect 3855 3945 3859 3953
rect 3865 3945 3869 3953
rect 3873 3945 3877 3953
rect 3913 3952 3917 3960
rect 3928 3952 3932 3960
rect 3943 3958 3947 3966
rect 3951 3958 3955 3966
rect 3970 3958 3974 3966
rect 3978 3958 3982 3966
rect 3994 3952 3998 3960
rect 4009 3952 4013 3960
rect 4024 3958 4028 3966
rect 4032 3958 4036 3966
rect 2404 3894 2408 3902
rect 2412 3894 2416 3902
rect 2420 3894 2424 3902
rect 2433 3894 2437 3902
rect 2441 3898 2445 3902
rect 2449 3894 2453 3902
rect 2457 3894 2461 3902
rect 2465 3894 2469 3902
rect 2478 3894 2482 3902
rect 2491 3894 2495 3902
rect 2499 3898 2503 3902
rect 2507 3894 2511 3902
rect 2515 3894 2519 3902
rect 2528 3894 2532 3902
rect 3349 3894 3353 3902
rect 3357 3894 3361 3902
rect 3365 3894 3369 3902
rect 3378 3894 3382 3902
rect 3386 3898 3390 3902
rect 3394 3894 3398 3902
rect 3402 3894 3406 3902
rect 3410 3894 3414 3902
rect 3423 3894 3427 3902
rect 3436 3894 3440 3902
rect 3444 3898 3448 3902
rect 3452 3894 3456 3902
rect 3460 3894 3464 3902
rect 3473 3894 3477 3902
rect 2770 3859 2774 3867
rect 2778 3859 2782 3867
rect 2786 3859 2790 3867
rect 2794 3859 2798 3867
rect 2802 3859 2806 3867
rect 2810 3859 2814 3867
rect 2821 3859 2825 3867
rect 2838 3859 2842 3867
rect 2855 3859 2859 3867
rect 2864 3859 2868 3867
rect 2877 3859 2881 3867
rect 2885 3859 2889 3867
rect 2893 3859 2897 3867
rect 2910 3859 2914 3867
rect 2920 3859 2924 3867
rect 2928 3859 2932 3867
rect 2968 3860 2972 3868
rect 2983 3860 2987 3868
rect 3049 3860 3053 3868
rect 3064 3860 3068 3868
rect 3715 3859 3719 3867
rect 3723 3859 3727 3867
rect 3731 3859 3735 3867
rect 3739 3859 3743 3867
rect 3747 3859 3751 3867
rect 3755 3859 3759 3867
rect 3766 3859 3770 3867
rect 3783 3859 3787 3867
rect 3800 3859 3804 3867
rect 3809 3859 3813 3867
rect 3822 3859 3826 3867
rect 3830 3859 3834 3867
rect 3838 3859 3842 3867
rect 3855 3859 3859 3867
rect 3865 3859 3869 3867
rect 3873 3859 3877 3867
rect 3913 3860 3917 3868
rect 3928 3860 3932 3868
rect 3994 3860 3998 3868
rect 4009 3860 4013 3868
rect 2770 3813 2774 3821
rect 2778 3813 2782 3821
rect 2786 3813 2790 3821
rect 2794 3813 2798 3821
rect 2802 3813 2806 3821
rect 2810 3813 2814 3821
rect 2821 3813 2825 3821
rect 2838 3813 2842 3821
rect 2855 3813 2859 3821
rect 2864 3813 2868 3821
rect 2877 3813 2881 3821
rect 2885 3813 2889 3821
rect 2893 3813 2897 3821
rect 2910 3813 2914 3821
rect 2920 3813 2924 3821
rect 2928 3813 2932 3821
rect 2968 3820 2972 3828
rect 2983 3820 2987 3828
rect 2998 3826 3002 3834
rect 3006 3826 3010 3834
rect 3049 3826 3053 3834
rect 3057 3826 3061 3834
rect 3073 3820 3077 3828
rect 3088 3820 3092 3828
rect 3103 3826 3107 3834
rect 3111 3826 3115 3834
rect 3715 3813 3719 3821
rect 3723 3813 3727 3821
rect 3731 3813 3735 3821
rect 3739 3813 3743 3821
rect 3747 3813 3751 3821
rect 3755 3813 3759 3821
rect 3766 3813 3770 3821
rect 3783 3813 3787 3821
rect 3800 3813 3804 3821
rect 3809 3813 3813 3821
rect 3822 3813 3826 3821
rect 3830 3813 3834 3821
rect 3838 3813 3842 3821
rect 3855 3813 3859 3821
rect 3865 3813 3869 3821
rect 3873 3813 3877 3821
rect 3913 3820 3917 3828
rect 3928 3820 3932 3828
rect 3943 3826 3947 3834
rect 3951 3826 3955 3834
rect 3994 3826 3998 3834
rect 4002 3826 4006 3834
rect 3280 3797 3284 3805
rect 3288 3797 3292 3805
rect 3304 3791 3308 3799
rect 3319 3791 3323 3799
rect 3334 3797 3338 3805
rect 3342 3797 3346 3805
rect 3454 3772 3470 3802
rect 3474 3772 3490 3802
rect 3507 3772 3523 3802
rect 3527 3772 3543 3802
rect 4018 3820 4022 3828
rect 4033 3820 4037 3828
rect 4048 3826 4052 3834
rect 4056 3826 4060 3834
rect 2770 3727 2774 3735
rect 2778 3727 2782 3735
rect 2786 3727 2790 3735
rect 2794 3727 2798 3735
rect 2802 3727 2806 3735
rect 2810 3727 2814 3735
rect 2821 3727 2825 3735
rect 2838 3727 2842 3735
rect 2855 3727 2859 3735
rect 2864 3727 2868 3735
rect 2877 3727 2881 3735
rect 2885 3727 2889 3735
rect 2893 3727 2897 3735
rect 2910 3727 2914 3735
rect 2920 3727 2924 3735
rect 2928 3727 2932 3735
rect 2968 3729 2972 3737
rect 2983 3729 2987 3737
rect 3073 3729 3077 3737
rect 3088 3729 3092 3737
rect 3715 3727 3719 3735
rect 3723 3727 3727 3735
rect 3731 3727 3735 3735
rect 3739 3727 3743 3735
rect 3747 3727 3751 3735
rect 3755 3727 3759 3735
rect 3766 3727 3770 3735
rect 3783 3727 3787 3735
rect 3800 3727 3804 3735
rect 3809 3727 3813 3735
rect 3822 3727 3826 3735
rect 3830 3727 3834 3735
rect 3838 3727 3842 3735
rect 3855 3727 3859 3735
rect 3865 3727 3869 3735
rect 3873 3727 3877 3735
rect 3913 3729 3917 3737
rect 3928 3729 3932 3737
rect 4018 3729 4022 3737
rect 4033 3729 4037 3737
rect 2770 3681 2774 3689
rect 2778 3681 2782 3689
rect 2786 3681 2790 3689
rect 2794 3681 2798 3689
rect 2802 3681 2806 3689
rect 2810 3681 2814 3689
rect 2821 3681 2825 3689
rect 2838 3681 2842 3689
rect 2855 3681 2859 3689
rect 2864 3681 2868 3689
rect 2877 3681 2881 3689
rect 2885 3681 2889 3689
rect 2893 3681 2897 3689
rect 2910 3681 2914 3689
rect 2920 3681 2924 3689
rect 2928 3681 2932 3689
rect 2968 3688 2972 3696
rect 2983 3688 2987 3696
rect 2998 3694 3002 3702
rect 3006 3694 3010 3702
rect 3025 3694 3029 3702
rect 3033 3694 3037 3702
rect 3049 3688 3053 3696
rect 3064 3688 3068 3696
rect 3079 3694 3083 3702
rect 3087 3694 3091 3702
rect 3115 3694 3119 3702
rect 3123 3694 3127 3702
rect 3139 3688 3143 3696
rect 3154 3688 3158 3696
rect 3169 3694 3173 3702
rect 3177 3694 3181 3702
rect 3304 3695 3308 3703
rect 3319 3695 3323 3703
rect 3715 3681 3719 3689
rect 3723 3681 3727 3689
rect 3731 3681 3735 3689
rect 3739 3681 3743 3689
rect 3747 3681 3751 3689
rect 3755 3681 3759 3689
rect 3766 3681 3770 3689
rect 3783 3681 3787 3689
rect 3800 3681 3804 3689
rect 3809 3681 3813 3689
rect 3822 3681 3826 3689
rect 3830 3681 3834 3689
rect 3838 3681 3842 3689
rect 3855 3681 3859 3689
rect 3865 3681 3869 3689
rect 3873 3681 3877 3689
rect 3913 3688 3917 3696
rect 3928 3688 3932 3696
rect 3943 3694 3947 3702
rect 3951 3694 3955 3702
rect 3970 3694 3974 3702
rect 3978 3694 3982 3702
rect 3258 3667 3262 3675
rect 3266 3667 3270 3675
rect 3280 3667 3284 3675
rect 3288 3667 3292 3675
rect 3304 3661 3308 3669
rect 3319 3661 3323 3669
rect 3334 3667 3338 3675
rect 3342 3667 3346 3675
rect 3360 3642 3376 3672
rect 3380 3642 3396 3672
rect 3413 3642 3429 3672
rect 3433 3642 3449 3672
rect 3994 3688 3998 3696
rect 4009 3688 4013 3696
rect 4024 3694 4028 3702
rect 4032 3694 4036 3702
rect 4060 3694 4064 3702
rect 4068 3694 4072 3702
rect 4084 3688 4088 3696
rect 4099 3688 4103 3696
rect 4114 3694 4118 3702
rect 4122 3694 4126 3702
rect 2770 3595 2774 3603
rect 2778 3595 2782 3603
rect 2786 3595 2790 3603
rect 2794 3595 2798 3603
rect 2802 3595 2806 3603
rect 2810 3595 2814 3603
rect 2821 3595 2825 3603
rect 2838 3595 2842 3603
rect 2855 3595 2859 3603
rect 2864 3595 2868 3603
rect 2877 3595 2881 3603
rect 2885 3595 2889 3603
rect 2893 3595 2897 3603
rect 2910 3595 2914 3603
rect 2920 3595 2924 3603
rect 2928 3595 2932 3603
rect 2968 3594 2972 3602
rect 2983 3594 2987 3602
rect 3049 3594 3053 3602
rect 3064 3594 3068 3602
rect 3139 3594 3143 3602
rect 3154 3594 3158 3602
rect 3715 3595 3719 3603
rect 3723 3595 3727 3603
rect 3731 3595 3735 3603
rect 3739 3595 3743 3603
rect 3747 3595 3751 3603
rect 3755 3595 3759 3603
rect 3766 3595 3770 3603
rect 3783 3595 3787 3603
rect 3800 3595 3804 3603
rect 3809 3595 3813 3603
rect 3822 3595 3826 3603
rect 3830 3595 3834 3603
rect 3838 3595 3842 3603
rect 3855 3595 3859 3603
rect 3865 3595 3869 3603
rect 3873 3595 3877 3603
rect 3913 3594 3917 3602
rect 3928 3594 3932 3602
rect 3994 3594 3998 3602
rect 4009 3594 4013 3602
rect 4084 3594 4088 3602
rect 4099 3594 4103 3602
rect 2770 3549 2774 3557
rect 2778 3549 2782 3557
rect 2786 3549 2790 3557
rect 2794 3549 2798 3557
rect 2802 3549 2806 3557
rect 2810 3549 2814 3557
rect 2821 3549 2825 3557
rect 2838 3549 2842 3557
rect 2855 3549 2859 3557
rect 2864 3549 2868 3557
rect 2877 3549 2881 3557
rect 2885 3549 2889 3557
rect 2893 3549 2897 3557
rect 2910 3549 2914 3557
rect 2920 3549 2924 3557
rect 2928 3549 2932 3557
rect 2968 3556 2972 3564
rect 2983 3556 2987 3564
rect 2998 3562 3002 3570
rect 3006 3562 3010 3570
rect 3304 3565 3308 3573
rect 3319 3565 3323 3573
rect 3715 3549 3719 3557
rect 3723 3549 3727 3557
rect 3731 3549 3735 3557
rect 3739 3549 3743 3557
rect 3747 3549 3751 3557
rect 3755 3549 3759 3557
rect 3766 3549 3770 3557
rect 3783 3549 3787 3557
rect 3800 3549 3804 3557
rect 3809 3549 3813 3557
rect 3822 3549 3826 3557
rect 3830 3549 3834 3557
rect 3838 3549 3842 3557
rect 3855 3549 3859 3557
rect 3865 3549 3869 3557
rect 3873 3549 3877 3557
rect 3913 3556 3917 3564
rect 3928 3556 3932 3564
rect 3943 3562 3947 3570
rect 3951 3562 3955 3570
rect 2281 3494 2285 3502
rect 2294 3494 2298 3502
rect 2302 3494 2306 3502
rect 2310 3498 2314 3502
rect 2318 3494 2322 3502
rect 2331 3494 2335 3502
rect 2344 3494 2348 3502
rect 2352 3494 2356 3502
rect 2360 3494 2364 3502
rect 2368 3498 2372 3502
rect 2376 3494 2380 3502
rect 2389 3494 2393 3502
rect 2397 3494 2401 3502
rect 2405 3494 2409 3502
rect 2413 3494 2417 3502
rect 2426 3494 2430 3502
rect 2434 3494 2438 3502
rect 2442 3498 2446 3502
rect 2450 3494 2454 3502
rect 2463 3494 2467 3502
rect 2476 3494 2480 3502
rect 2484 3494 2488 3502
rect 2492 3494 2496 3502
rect 2500 3498 2504 3502
rect 2508 3494 2512 3502
rect 2521 3494 2525 3502
rect 2529 3494 2533 3502
rect 2537 3494 2541 3502
rect 2545 3494 2549 3502
rect 2558 3494 2562 3502
rect 2566 3494 2570 3502
rect 2574 3498 2578 3502
rect 2582 3494 2586 3502
rect 2595 3494 2599 3502
rect 2608 3494 2612 3502
rect 2616 3494 2620 3502
rect 2624 3494 2628 3502
rect 2632 3498 2636 3502
rect 2640 3494 2644 3502
rect 2653 3494 2657 3502
rect 2661 3494 2665 3502
rect 2669 3494 2673 3502
rect 3226 3494 3230 3502
rect 3239 3494 3243 3502
rect 3247 3494 3251 3502
rect 3255 3498 3259 3502
rect 3263 3494 3267 3502
rect 3276 3494 3280 3502
rect 3289 3494 3293 3502
rect 3297 3494 3301 3502
rect 3305 3494 3309 3502
rect 3313 3498 3317 3502
rect 3321 3494 3325 3502
rect 3334 3494 3338 3502
rect 3342 3494 3346 3502
rect 3350 3494 3354 3502
rect 3358 3494 3362 3502
rect 3371 3494 3375 3502
rect 3379 3494 3383 3502
rect 3387 3498 3391 3502
rect 3395 3494 3399 3502
rect 3408 3494 3412 3502
rect 3421 3494 3425 3502
rect 3429 3494 3433 3502
rect 3437 3494 3441 3502
rect 3445 3498 3449 3502
rect 3453 3494 3457 3502
rect 3466 3494 3470 3502
rect 3474 3494 3478 3502
rect 3482 3494 3486 3502
rect 3490 3494 3494 3502
rect 3503 3494 3507 3502
rect 3511 3494 3515 3502
rect 3519 3498 3523 3502
rect 3527 3494 3531 3502
rect 3540 3494 3544 3502
rect 3553 3494 3557 3502
rect 3561 3494 3565 3502
rect 3569 3494 3573 3502
rect 3577 3498 3581 3502
rect 3585 3494 3589 3502
rect 3598 3494 3602 3502
rect 3606 3494 3610 3502
rect 3614 3494 3618 3502
rect 2770 3463 2774 3471
rect 2778 3463 2782 3471
rect 2786 3463 2790 3471
rect 2794 3463 2798 3471
rect 2802 3463 2806 3471
rect 2810 3463 2814 3471
rect 2821 3463 2825 3471
rect 2838 3463 2842 3471
rect 2855 3463 2859 3471
rect 2864 3463 2868 3471
rect 2877 3463 2881 3471
rect 2885 3463 2889 3471
rect 2893 3463 2897 3471
rect 2910 3463 2914 3471
rect 2920 3463 2924 3471
rect 2928 3463 2932 3471
rect 2968 3458 2972 3466
rect 2983 3458 2987 3466
rect 3004 3463 3008 3471
rect 3012 3463 3016 3471
rect 3022 3463 3026 3471
rect 3030 3463 3034 3471
rect 3039 3463 3043 3471
rect 3047 3463 3051 3471
rect 3055 3463 3059 3471
rect 3063 3463 3067 3471
rect 3071 3463 3075 3471
rect 3082 3463 3086 3471
rect 3099 3463 3103 3471
rect 3116 3463 3120 3471
rect 3125 3463 3129 3471
rect 3138 3463 3142 3471
rect 3146 3463 3150 3471
rect 3154 3463 3158 3471
rect 3171 3463 3175 3471
rect 3181 3463 3185 3471
rect 3189 3463 3193 3471
rect 3715 3463 3719 3471
rect 3723 3463 3727 3471
rect 3731 3463 3735 3471
rect 3739 3463 3743 3471
rect 3747 3463 3751 3471
rect 3755 3463 3759 3471
rect 3766 3463 3770 3471
rect 3783 3463 3787 3471
rect 3800 3463 3804 3471
rect 3809 3463 3813 3471
rect 3822 3463 3826 3471
rect 3830 3463 3834 3471
rect 3838 3463 3842 3471
rect 3855 3463 3859 3471
rect 3865 3463 3869 3471
rect 3873 3463 3877 3471
rect 3913 3458 3917 3466
rect 3928 3458 3932 3466
rect 3949 3463 3953 3471
rect 3957 3463 3961 3471
rect 3967 3463 3971 3471
rect 3975 3463 3979 3471
rect 3984 3463 3988 3471
rect 3992 3463 3996 3471
rect 4000 3463 4004 3471
rect 4008 3463 4012 3471
rect 4016 3463 4020 3471
rect 4027 3463 4031 3471
rect 4044 3463 4048 3471
rect 4061 3463 4065 3471
rect 4070 3463 4074 3471
rect 4083 3463 4087 3471
rect 4091 3463 4095 3471
rect 4099 3463 4103 3471
rect 4116 3463 4120 3471
rect 4126 3463 4130 3471
rect 4134 3463 4138 3471
rect 3064 3382 3068 3390
rect 3077 3382 3081 3390
rect 3085 3382 3089 3390
rect 3093 3386 3097 3390
rect 3101 3382 3105 3390
rect 3114 3382 3118 3390
rect 3127 3382 3131 3390
rect 3135 3382 3139 3390
rect 3143 3382 3147 3390
rect 3151 3386 3155 3390
rect 3159 3382 3163 3390
rect 3172 3382 3176 3390
rect 3180 3382 3184 3390
rect 3188 3382 3192 3390
rect 4009 3382 4013 3390
rect 4022 3382 4026 3390
rect 4030 3382 4034 3390
rect 4038 3386 4042 3390
rect 4046 3382 4050 3390
rect 4059 3382 4063 3390
rect 4072 3382 4076 3390
rect 4080 3382 4084 3390
rect 4088 3382 4092 3390
rect 4096 3386 4100 3390
rect 4104 3382 4108 3390
rect 4117 3382 4121 3390
rect 4125 3382 4129 3390
rect 4133 3382 4137 3390
rect 2281 3352 2285 3360
rect 2294 3352 2298 3360
rect 2302 3352 2306 3360
rect 2310 3356 2314 3360
rect 2318 3352 2322 3360
rect 2331 3352 2335 3360
rect 2344 3352 2348 3360
rect 2352 3352 2356 3360
rect 2360 3352 2364 3360
rect 2368 3356 2372 3360
rect 2376 3352 2380 3360
rect 2389 3352 2393 3360
rect 2397 3352 2401 3360
rect 2405 3352 2409 3360
rect 2413 3352 2417 3360
rect 2426 3352 2430 3360
rect 2434 3352 2438 3360
rect 2442 3356 2446 3360
rect 2450 3352 2454 3360
rect 2463 3352 2467 3360
rect 2476 3352 2480 3360
rect 2484 3352 2488 3360
rect 2492 3352 2496 3360
rect 2500 3356 2504 3360
rect 2508 3352 2512 3360
rect 2521 3352 2525 3360
rect 2529 3352 2533 3360
rect 2537 3352 2541 3360
rect 2545 3352 2549 3360
rect 2558 3352 2562 3360
rect 2566 3352 2570 3360
rect 2574 3356 2578 3360
rect 2582 3352 2586 3360
rect 2595 3352 2599 3360
rect 2608 3352 2612 3360
rect 2616 3352 2620 3360
rect 2624 3352 2628 3360
rect 2632 3356 2636 3360
rect 2640 3352 2644 3360
rect 2653 3352 2657 3360
rect 2661 3352 2665 3360
rect 2669 3352 2673 3360
rect 3226 3352 3230 3360
rect 3239 3352 3243 3360
rect 3247 3352 3251 3360
rect 3255 3356 3259 3360
rect 3263 3352 3267 3360
rect 3276 3352 3280 3360
rect 3289 3352 3293 3360
rect 3297 3352 3301 3360
rect 3305 3352 3309 3360
rect 3313 3356 3317 3360
rect 3321 3352 3325 3360
rect 3334 3352 3338 3360
rect 3342 3352 3346 3360
rect 3350 3352 3354 3360
rect 3358 3352 3362 3360
rect 3371 3352 3375 3360
rect 3379 3352 3383 3360
rect 3387 3356 3391 3360
rect 3395 3352 3399 3360
rect 3408 3352 3412 3360
rect 3421 3352 3425 3360
rect 3429 3352 3433 3360
rect 3437 3352 3441 3360
rect 3445 3356 3449 3360
rect 3453 3352 3457 3360
rect 3466 3352 3470 3360
rect 3474 3352 3478 3360
rect 3482 3352 3486 3360
rect 3490 3352 3494 3360
rect 3503 3352 3507 3360
rect 3511 3352 3515 3360
rect 3519 3356 3523 3360
rect 3527 3352 3531 3360
rect 3540 3352 3544 3360
rect 3553 3352 3557 3360
rect 3561 3352 3565 3360
rect 3569 3352 3573 3360
rect 3577 3356 3581 3360
rect 3585 3352 3589 3360
rect 3598 3352 3602 3360
rect 3606 3352 3610 3360
rect 3614 3352 3618 3360
rect 3064 3296 3068 3304
rect 3077 3296 3081 3304
rect 3085 3296 3089 3304
rect 3093 3300 3097 3304
rect 3101 3296 3105 3304
rect 3114 3296 3118 3304
rect 3127 3296 3131 3304
rect 3135 3296 3139 3304
rect 3143 3296 3147 3304
rect 3151 3300 3155 3304
rect 3159 3296 3163 3304
rect 3172 3296 3176 3304
rect 3180 3296 3184 3304
rect 3188 3296 3192 3304
rect 4009 3296 4013 3304
rect 4022 3296 4026 3304
rect 4030 3296 4034 3304
rect 4038 3300 4042 3304
rect 4046 3296 4050 3304
rect 4059 3296 4063 3304
rect 4072 3296 4076 3304
rect 4080 3296 4084 3304
rect 4088 3296 4092 3304
rect 4096 3300 4100 3304
rect 4104 3296 4108 3304
rect 4117 3296 4121 3304
rect 4125 3296 4129 3304
rect 4133 3296 4137 3304
rect 2281 3266 2285 3274
rect 2294 3266 2298 3274
rect 2302 3266 2306 3274
rect 2310 3270 2314 3274
rect 2318 3266 2322 3274
rect 2331 3266 2335 3274
rect 2344 3266 2348 3274
rect 2352 3266 2356 3274
rect 2360 3266 2364 3274
rect 2368 3270 2372 3274
rect 2376 3266 2380 3274
rect 2389 3266 2393 3274
rect 2397 3266 2401 3274
rect 2405 3266 2409 3274
rect 2413 3266 2417 3274
rect 2426 3266 2430 3274
rect 2434 3266 2438 3274
rect 2442 3270 2446 3274
rect 2450 3266 2454 3274
rect 2463 3266 2467 3274
rect 2476 3266 2480 3274
rect 2484 3266 2488 3274
rect 2492 3266 2496 3274
rect 2500 3270 2504 3274
rect 2508 3266 2512 3274
rect 2521 3266 2525 3274
rect 2529 3266 2533 3274
rect 2537 3266 2541 3274
rect 2545 3266 2549 3274
rect 2558 3266 2562 3274
rect 2566 3266 2570 3274
rect 2574 3270 2578 3274
rect 2582 3266 2586 3274
rect 2595 3266 2599 3274
rect 2608 3266 2612 3274
rect 2616 3266 2620 3274
rect 2624 3266 2628 3274
rect 2632 3270 2636 3274
rect 2640 3266 2644 3274
rect 2653 3266 2657 3274
rect 2661 3266 2665 3274
rect 2669 3266 2673 3274
rect 3226 3266 3230 3274
rect 3239 3266 3243 3274
rect 3247 3266 3251 3274
rect 3255 3270 3259 3274
rect 3263 3266 3267 3274
rect 3276 3266 3280 3274
rect 3289 3266 3293 3274
rect 3297 3266 3301 3274
rect 3305 3266 3309 3274
rect 3313 3270 3317 3274
rect 3321 3266 3325 3274
rect 3334 3266 3338 3274
rect 3342 3266 3346 3274
rect 3350 3266 3354 3274
rect 3358 3266 3362 3274
rect 3371 3266 3375 3274
rect 3379 3266 3383 3274
rect 3387 3270 3391 3274
rect 3395 3266 3399 3274
rect 3408 3266 3412 3274
rect 3421 3266 3425 3274
rect 3429 3266 3433 3274
rect 3437 3266 3441 3274
rect 3445 3270 3449 3274
rect 3453 3266 3457 3274
rect 3466 3266 3470 3274
rect 3474 3266 3478 3274
rect 3482 3266 3486 3274
rect 3490 3266 3494 3274
rect 3503 3266 3507 3274
rect 3511 3266 3515 3274
rect 3519 3270 3523 3274
rect 3527 3266 3531 3274
rect 3540 3266 3544 3274
rect 3553 3266 3557 3274
rect 3561 3266 3565 3274
rect 3569 3266 3573 3274
rect 3577 3270 3581 3274
rect 3585 3266 3589 3274
rect 3598 3266 3602 3274
rect 3606 3266 3610 3274
rect 3614 3266 3618 3274
rect 2281 3126 2285 3134
rect 2294 3126 2298 3134
rect 2302 3126 2306 3134
rect 2310 3130 2314 3134
rect 2318 3126 2322 3134
rect 2331 3126 2335 3134
rect 2344 3126 2348 3134
rect 2352 3126 2356 3134
rect 2360 3126 2364 3134
rect 2368 3130 2372 3134
rect 2376 3126 2380 3134
rect 2389 3126 2393 3134
rect 2397 3126 2401 3134
rect 2405 3126 2409 3134
rect 2413 3126 2417 3134
rect 2426 3126 2430 3134
rect 2434 3126 2438 3134
rect 2442 3130 2446 3134
rect 2450 3126 2454 3134
rect 2463 3126 2467 3134
rect 2476 3126 2480 3134
rect 2484 3126 2488 3134
rect 2492 3126 2496 3134
rect 2500 3130 2504 3134
rect 2508 3126 2512 3134
rect 2521 3126 2525 3134
rect 2529 3126 2533 3134
rect 2537 3126 2541 3134
rect 2545 3126 2549 3134
rect 2558 3126 2562 3134
rect 2566 3126 2570 3134
rect 2574 3130 2578 3134
rect 2582 3126 2586 3134
rect 2595 3126 2599 3134
rect 2608 3126 2612 3134
rect 2616 3126 2620 3134
rect 2624 3126 2628 3134
rect 2632 3130 2636 3134
rect 2640 3126 2644 3134
rect 2653 3126 2657 3134
rect 2661 3126 2665 3134
rect 2669 3126 2673 3134
rect 3226 3126 3230 3134
rect 3239 3126 3243 3134
rect 3247 3126 3251 3134
rect 3255 3130 3259 3134
rect 3263 3126 3267 3134
rect 3276 3126 3280 3134
rect 3289 3126 3293 3134
rect 3297 3126 3301 3134
rect 3305 3126 3309 3134
rect 3313 3130 3317 3134
rect 3321 3126 3325 3134
rect 3334 3126 3338 3134
rect 3342 3126 3346 3134
rect 3350 3126 3354 3134
rect 3358 3126 3362 3134
rect 3371 3126 3375 3134
rect 3379 3126 3383 3134
rect 3387 3130 3391 3134
rect 3395 3126 3399 3134
rect 3408 3126 3412 3134
rect 3421 3126 3425 3134
rect 3429 3126 3433 3134
rect 3437 3126 3441 3134
rect 3445 3130 3449 3134
rect 3453 3126 3457 3134
rect 3466 3126 3470 3134
rect 3474 3126 3478 3134
rect 3482 3126 3486 3134
rect 3490 3126 3494 3134
rect 3503 3126 3507 3134
rect 3511 3126 3515 3134
rect 3519 3130 3523 3134
rect 3527 3126 3531 3134
rect 3540 3126 3544 3134
rect 3553 3126 3557 3134
rect 3561 3126 3565 3134
rect 3569 3126 3573 3134
rect 3577 3130 3581 3134
rect 3585 3126 3589 3134
rect 3598 3126 3602 3134
rect 3606 3126 3610 3134
rect 3614 3126 3618 3134
rect 2765 3047 2769 3055
rect 2778 3047 2782 3055
rect 2786 3047 2790 3055
rect 2794 3051 2798 3055
rect 2802 3047 2806 3055
rect 2815 3047 2819 3055
rect 2828 3047 2832 3055
rect 2836 3047 2840 3055
rect 2844 3047 2848 3055
rect 2852 3051 2856 3055
rect 2860 3047 2864 3055
rect 2873 3047 2877 3055
rect 2881 3047 2885 3055
rect 2889 3047 2893 3055
rect 2897 3047 2901 3055
rect 2910 3047 2914 3055
rect 2918 3047 2922 3055
rect 2926 3051 2930 3055
rect 2934 3047 2938 3055
rect 2947 3047 2951 3055
rect 2960 3047 2964 3055
rect 2968 3047 2972 3055
rect 2976 3047 2980 3055
rect 2984 3051 2988 3055
rect 2992 3047 2996 3055
rect 3005 3047 3009 3055
rect 3013 3047 3017 3055
rect 3021 3047 3025 3055
rect 3029 3047 3033 3055
rect 3042 3047 3046 3055
rect 3050 3047 3054 3055
rect 3058 3051 3062 3055
rect 3066 3047 3070 3055
rect 3079 3047 3083 3055
rect 3092 3047 3096 3055
rect 3100 3047 3104 3055
rect 3108 3047 3112 3055
rect 3116 3051 3120 3055
rect 3124 3047 3128 3055
rect 3137 3047 3141 3055
rect 3145 3047 3149 3055
rect 3153 3047 3157 3055
rect 3161 3047 3165 3055
rect 3174 3047 3178 3055
rect 3182 3047 3186 3055
rect 3190 3051 3194 3055
rect 3198 3047 3202 3055
rect 3211 3047 3215 3055
rect 3224 3047 3228 3055
rect 3232 3047 3236 3055
rect 3240 3047 3244 3055
rect 3248 3051 3252 3055
rect 3256 3047 3260 3055
rect 3269 3047 3273 3055
rect 3277 3047 3281 3055
rect 3285 3047 3289 3055
rect 3710 3047 3714 3055
rect 3723 3047 3727 3055
rect 3731 3047 3735 3055
rect 3739 3051 3743 3055
rect 3747 3047 3751 3055
rect 3760 3047 3764 3055
rect 3773 3047 3777 3055
rect 3781 3047 3785 3055
rect 3789 3047 3793 3055
rect 3797 3051 3801 3055
rect 3805 3047 3809 3055
rect 3818 3047 3822 3055
rect 3826 3047 3830 3055
rect 3834 3047 3838 3055
rect 3842 3047 3846 3055
rect 3855 3047 3859 3055
rect 3863 3047 3867 3055
rect 3871 3051 3875 3055
rect 3879 3047 3883 3055
rect 3892 3047 3896 3055
rect 3905 3047 3909 3055
rect 3913 3047 3917 3055
rect 3921 3047 3925 3055
rect 3929 3051 3933 3055
rect 3937 3047 3941 3055
rect 3950 3047 3954 3055
rect 3958 3047 3962 3055
rect 3966 3047 3970 3055
rect 3974 3047 3978 3055
rect 3987 3047 3991 3055
rect 3995 3047 3999 3055
rect 4003 3051 4007 3055
rect 4011 3047 4015 3055
rect 4024 3047 4028 3055
rect 4037 3047 4041 3055
rect 4045 3047 4049 3055
rect 4053 3047 4057 3055
rect 4061 3051 4065 3055
rect 4069 3047 4073 3055
rect 4082 3047 4086 3055
rect 4090 3047 4094 3055
rect 4098 3047 4102 3055
rect 4106 3047 4110 3055
rect 4119 3047 4123 3055
rect 4127 3047 4131 3055
rect 4135 3051 4139 3055
rect 4143 3047 4147 3055
rect 4156 3047 4160 3055
rect 4169 3047 4173 3055
rect 4177 3047 4181 3055
rect 4185 3047 4189 3055
rect 4193 3051 4197 3055
rect 4201 3047 4205 3055
rect 4214 3047 4218 3055
rect 4222 3047 4226 3055
rect 4230 3047 4234 3055
rect 2413 3014 2417 3022
rect 2426 3014 2430 3022
rect 2434 3014 2438 3022
rect 2442 3018 2446 3022
rect 2450 3014 2454 3022
rect 2463 3014 2467 3022
rect 2476 3014 2480 3022
rect 2484 3014 2488 3022
rect 2492 3014 2496 3022
rect 2500 3018 2504 3022
rect 2508 3014 2512 3022
rect 2521 3014 2525 3022
rect 2529 3014 2533 3022
rect 2537 3014 2541 3022
rect 3358 3014 3362 3022
rect 3371 3014 3375 3022
rect 3379 3014 3383 3022
rect 3387 3018 3391 3022
rect 3395 3014 3399 3022
rect 3408 3014 3412 3022
rect 3421 3014 3425 3022
rect 3429 3014 3433 3022
rect 3437 3014 3441 3022
rect 3445 3018 3449 3022
rect 3453 3014 3457 3022
rect 3466 3014 3470 3022
rect 3474 3014 3478 3022
rect 3482 3014 3486 3022
rect 2944 2976 2948 2984
rect 2952 2976 2956 2984
rect 2770 2963 2774 2971
rect 2778 2963 2782 2971
rect 2786 2963 2790 2971
rect 2794 2963 2798 2971
rect 2802 2963 2806 2971
rect 2810 2963 2814 2971
rect 2821 2963 2825 2971
rect 2838 2963 2842 2971
rect 2855 2963 2859 2971
rect 2864 2963 2868 2971
rect 2877 2963 2881 2971
rect 2885 2963 2889 2971
rect 2893 2963 2897 2971
rect 2910 2963 2914 2971
rect 2920 2963 2924 2971
rect 2928 2963 2932 2971
rect 2968 2970 2972 2978
rect 2983 2970 2987 2978
rect 2998 2976 3002 2984
rect 3006 2976 3010 2984
rect 3025 2976 3029 2984
rect 3033 2976 3037 2984
rect 3049 2970 3053 2978
rect 3064 2970 3068 2978
rect 3079 2976 3083 2984
rect 3087 2976 3091 2984
rect 3889 2976 3893 2984
rect 3897 2976 3901 2984
rect 3715 2963 3719 2971
rect 3723 2963 3727 2971
rect 3731 2963 3735 2971
rect 3739 2963 3743 2971
rect 3747 2963 3751 2971
rect 3755 2963 3759 2971
rect 3766 2963 3770 2971
rect 3783 2963 3787 2971
rect 3800 2963 3804 2971
rect 3809 2963 3813 2971
rect 3822 2963 3826 2971
rect 3830 2963 3834 2971
rect 3838 2963 3842 2971
rect 3855 2963 3859 2971
rect 3865 2963 3869 2971
rect 3873 2963 3877 2971
rect 3913 2970 3917 2978
rect 3928 2970 3932 2978
rect 3943 2976 3947 2984
rect 3951 2976 3955 2984
rect 3970 2976 3974 2984
rect 3978 2976 3982 2984
rect 3994 2970 3998 2978
rect 4009 2970 4013 2978
rect 4024 2976 4028 2984
rect 4032 2976 4036 2984
rect 2404 2912 2408 2920
rect 2412 2912 2416 2920
rect 2420 2912 2424 2920
rect 2433 2912 2437 2920
rect 2441 2916 2445 2920
rect 2449 2912 2453 2920
rect 2457 2912 2461 2920
rect 2465 2912 2469 2920
rect 2478 2912 2482 2920
rect 2491 2912 2495 2920
rect 2499 2916 2503 2920
rect 2507 2912 2511 2920
rect 2515 2912 2519 2920
rect 2528 2912 2532 2920
rect 3349 2912 3353 2920
rect 3357 2912 3361 2920
rect 3365 2912 3369 2920
rect 3378 2912 3382 2920
rect 3386 2916 3390 2920
rect 3394 2912 3398 2920
rect 3402 2912 3406 2920
rect 3410 2912 3414 2920
rect 3423 2912 3427 2920
rect 3436 2912 3440 2920
rect 3444 2916 3448 2920
rect 3452 2912 3456 2920
rect 3460 2912 3464 2920
rect 3473 2912 3477 2920
rect 2770 2877 2774 2885
rect 2778 2877 2782 2885
rect 2786 2877 2790 2885
rect 2794 2877 2798 2885
rect 2802 2877 2806 2885
rect 2810 2877 2814 2885
rect 2821 2877 2825 2885
rect 2838 2877 2842 2885
rect 2855 2877 2859 2885
rect 2864 2877 2868 2885
rect 2877 2877 2881 2885
rect 2885 2877 2889 2885
rect 2893 2877 2897 2885
rect 2910 2877 2914 2885
rect 2920 2877 2924 2885
rect 2928 2877 2932 2885
rect 2968 2878 2972 2886
rect 2983 2878 2987 2886
rect 3049 2878 3053 2886
rect 3064 2878 3068 2886
rect 3715 2877 3719 2885
rect 3723 2877 3727 2885
rect 3731 2877 3735 2885
rect 3739 2877 3743 2885
rect 3747 2877 3751 2885
rect 3755 2877 3759 2885
rect 3766 2877 3770 2885
rect 3783 2877 3787 2885
rect 3800 2877 3804 2885
rect 3809 2877 3813 2885
rect 3822 2877 3826 2885
rect 3830 2877 3834 2885
rect 3838 2877 3842 2885
rect 3855 2877 3859 2885
rect 3865 2877 3869 2885
rect 3873 2877 3877 2885
rect 3913 2878 3917 2886
rect 3928 2878 3932 2886
rect 3994 2878 3998 2886
rect 4009 2878 4013 2886
rect 2770 2831 2774 2839
rect 2778 2831 2782 2839
rect 2786 2831 2790 2839
rect 2794 2831 2798 2839
rect 2802 2831 2806 2839
rect 2810 2831 2814 2839
rect 2821 2831 2825 2839
rect 2838 2831 2842 2839
rect 2855 2831 2859 2839
rect 2864 2831 2868 2839
rect 2877 2831 2881 2839
rect 2885 2831 2889 2839
rect 2893 2831 2897 2839
rect 2910 2831 2914 2839
rect 2920 2831 2924 2839
rect 2928 2831 2932 2839
rect 2968 2838 2972 2846
rect 2983 2838 2987 2846
rect 2998 2844 3002 2852
rect 3006 2844 3010 2852
rect 3049 2844 3053 2852
rect 3057 2844 3061 2852
rect 3073 2838 3077 2846
rect 3088 2838 3092 2846
rect 3103 2844 3107 2852
rect 3111 2844 3115 2852
rect 3715 2831 3719 2839
rect 3723 2831 3727 2839
rect 3731 2831 3735 2839
rect 3739 2831 3743 2839
rect 3747 2831 3751 2839
rect 3755 2831 3759 2839
rect 3766 2831 3770 2839
rect 3783 2831 3787 2839
rect 3800 2831 3804 2839
rect 3809 2831 3813 2839
rect 3822 2831 3826 2839
rect 3830 2831 3834 2839
rect 3838 2831 3842 2839
rect 3855 2831 3859 2839
rect 3865 2831 3869 2839
rect 3873 2831 3877 2839
rect 3913 2838 3917 2846
rect 3928 2838 3932 2846
rect 3943 2844 3947 2852
rect 3951 2844 3955 2852
rect 3994 2844 3998 2852
rect 4002 2844 4006 2852
rect 4018 2838 4022 2846
rect 4033 2838 4037 2846
rect 4048 2844 4052 2852
rect 4056 2844 4060 2852
rect 2770 2745 2774 2753
rect 2778 2745 2782 2753
rect 2786 2745 2790 2753
rect 2794 2745 2798 2753
rect 2802 2745 2806 2753
rect 2810 2745 2814 2753
rect 2821 2745 2825 2753
rect 2838 2745 2842 2753
rect 2855 2745 2859 2753
rect 2864 2745 2868 2753
rect 2877 2745 2881 2753
rect 2885 2745 2889 2753
rect 2893 2745 2897 2753
rect 2910 2745 2914 2753
rect 2920 2745 2924 2753
rect 2928 2745 2932 2753
rect 2968 2747 2972 2755
rect 2983 2747 2987 2755
rect 3073 2747 3077 2755
rect 3088 2747 3092 2755
rect 3715 2745 3719 2753
rect 3723 2745 3727 2753
rect 3731 2745 3735 2753
rect 3739 2745 3743 2753
rect 3747 2745 3751 2753
rect 3755 2745 3759 2753
rect 3766 2745 3770 2753
rect 3783 2745 3787 2753
rect 3800 2745 3804 2753
rect 3809 2745 3813 2753
rect 3822 2745 3826 2753
rect 3830 2745 3834 2753
rect 3838 2745 3842 2753
rect 3855 2745 3859 2753
rect 3865 2745 3869 2753
rect 3873 2745 3877 2753
rect 3913 2747 3917 2755
rect 3928 2747 3932 2755
rect 4018 2747 4022 2755
rect 4033 2747 4037 2755
rect 2770 2699 2774 2707
rect 2778 2699 2782 2707
rect 2786 2699 2790 2707
rect 2794 2699 2798 2707
rect 2802 2699 2806 2707
rect 2810 2699 2814 2707
rect 2821 2699 2825 2707
rect 2838 2699 2842 2707
rect 2855 2699 2859 2707
rect 2864 2699 2868 2707
rect 2877 2699 2881 2707
rect 2885 2699 2889 2707
rect 2893 2699 2897 2707
rect 2910 2699 2914 2707
rect 2920 2699 2924 2707
rect 2928 2699 2932 2707
rect 2968 2706 2972 2714
rect 2983 2706 2987 2714
rect 2998 2712 3002 2720
rect 3006 2712 3010 2720
rect 3025 2712 3029 2720
rect 3033 2712 3037 2720
rect 3049 2706 3053 2714
rect 3064 2706 3068 2714
rect 3079 2712 3083 2720
rect 3087 2712 3091 2720
rect 3115 2712 3119 2720
rect 3123 2712 3127 2720
rect 3139 2706 3143 2714
rect 3154 2706 3158 2714
rect 3169 2712 3173 2720
rect 3177 2712 3181 2720
rect 3715 2699 3719 2707
rect 3723 2699 3727 2707
rect 3731 2699 3735 2707
rect 3739 2699 3743 2707
rect 3747 2699 3751 2707
rect 3755 2699 3759 2707
rect 3766 2699 3770 2707
rect 3783 2699 3787 2707
rect 3800 2699 3804 2707
rect 3809 2699 3813 2707
rect 3822 2699 3826 2707
rect 3830 2699 3834 2707
rect 3838 2699 3842 2707
rect 3855 2699 3859 2707
rect 3865 2699 3869 2707
rect 3873 2699 3877 2707
rect 3913 2706 3917 2714
rect 3928 2706 3932 2714
rect 3943 2712 3947 2720
rect 3951 2712 3955 2720
rect 3970 2712 3974 2720
rect 3978 2712 3982 2720
rect 3994 2706 3998 2714
rect 4009 2706 4013 2714
rect 4024 2712 4028 2720
rect 4032 2712 4036 2720
rect 4060 2712 4064 2720
rect 4068 2712 4072 2720
rect 4084 2706 4088 2714
rect 4099 2706 4103 2714
rect 4114 2712 4118 2720
rect 4122 2712 4126 2720
rect 2770 2613 2774 2621
rect 2778 2613 2782 2621
rect 2786 2613 2790 2621
rect 2794 2613 2798 2621
rect 2802 2613 2806 2621
rect 2810 2613 2814 2621
rect 2821 2613 2825 2621
rect 2838 2613 2842 2621
rect 2855 2613 2859 2621
rect 2864 2613 2868 2621
rect 2877 2613 2881 2621
rect 2885 2613 2889 2621
rect 2893 2613 2897 2621
rect 2910 2613 2914 2621
rect 2920 2613 2924 2621
rect 2928 2613 2932 2621
rect 2968 2612 2972 2620
rect 2983 2612 2987 2620
rect 3049 2612 3053 2620
rect 3064 2612 3068 2620
rect 3139 2612 3143 2620
rect 3154 2612 3158 2620
rect 3715 2613 3719 2621
rect 3723 2613 3727 2621
rect 3731 2613 3735 2621
rect 3739 2613 3743 2621
rect 3747 2613 3751 2621
rect 3755 2613 3759 2621
rect 3766 2613 3770 2621
rect 3783 2613 3787 2621
rect 3800 2613 3804 2621
rect 3809 2613 3813 2621
rect 3822 2613 3826 2621
rect 3830 2613 3834 2621
rect 3838 2613 3842 2621
rect 3855 2613 3859 2621
rect 3865 2613 3869 2621
rect 3873 2613 3877 2621
rect 3913 2612 3917 2620
rect 3928 2612 3932 2620
rect 3994 2612 3998 2620
rect 4009 2612 4013 2620
rect 4084 2612 4088 2620
rect 4099 2612 4103 2620
rect 2770 2567 2774 2575
rect 2778 2567 2782 2575
rect 2786 2567 2790 2575
rect 2794 2567 2798 2575
rect 2802 2567 2806 2575
rect 2810 2567 2814 2575
rect 2821 2567 2825 2575
rect 2838 2567 2842 2575
rect 2855 2567 2859 2575
rect 2864 2567 2868 2575
rect 2877 2567 2881 2575
rect 2885 2567 2889 2575
rect 2893 2567 2897 2575
rect 2910 2567 2914 2575
rect 2920 2567 2924 2575
rect 2928 2567 2932 2575
rect 2968 2574 2972 2582
rect 2983 2574 2987 2582
rect 2998 2580 3002 2588
rect 3006 2580 3010 2588
rect 3715 2567 3719 2575
rect 3723 2567 3727 2575
rect 3731 2567 3735 2575
rect 3739 2567 3743 2575
rect 3747 2567 3751 2575
rect 3755 2567 3759 2575
rect 3766 2567 3770 2575
rect 3783 2567 3787 2575
rect 3800 2567 3804 2575
rect 3809 2567 3813 2575
rect 3822 2567 3826 2575
rect 3830 2567 3834 2575
rect 3838 2567 3842 2575
rect 3855 2567 3859 2575
rect 3865 2567 3869 2575
rect 3873 2567 3877 2575
rect 3913 2574 3917 2582
rect 3928 2574 3932 2582
rect 3943 2580 3947 2588
rect 3951 2580 3955 2588
rect 2281 2512 2285 2520
rect 2294 2512 2298 2520
rect 2302 2512 2306 2520
rect 2310 2516 2314 2520
rect 2318 2512 2322 2520
rect 2331 2512 2335 2520
rect 2344 2512 2348 2520
rect 2352 2512 2356 2520
rect 2360 2512 2364 2520
rect 2368 2516 2372 2520
rect 2376 2512 2380 2520
rect 2389 2512 2393 2520
rect 2397 2512 2401 2520
rect 2405 2512 2409 2520
rect 2413 2512 2417 2520
rect 2426 2512 2430 2520
rect 2434 2512 2438 2520
rect 2442 2516 2446 2520
rect 2450 2512 2454 2520
rect 2463 2512 2467 2520
rect 2476 2512 2480 2520
rect 2484 2512 2488 2520
rect 2492 2512 2496 2520
rect 2500 2516 2504 2520
rect 2508 2512 2512 2520
rect 2521 2512 2525 2520
rect 2529 2512 2533 2520
rect 2537 2512 2541 2520
rect 2545 2512 2549 2520
rect 2558 2512 2562 2520
rect 2566 2512 2570 2520
rect 2574 2516 2578 2520
rect 2582 2512 2586 2520
rect 2595 2512 2599 2520
rect 2608 2512 2612 2520
rect 2616 2512 2620 2520
rect 2624 2512 2628 2520
rect 2632 2516 2636 2520
rect 2640 2512 2644 2520
rect 2653 2512 2657 2520
rect 2661 2512 2665 2520
rect 2669 2512 2673 2520
rect 3226 2512 3230 2520
rect 3239 2512 3243 2520
rect 3247 2512 3251 2520
rect 3255 2516 3259 2520
rect 3263 2512 3267 2520
rect 3276 2512 3280 2520
rect 3289 2512 3293 2520
rect 3297 2512 3301 2520
rect 3305 2512 3309 2520
rect 3313 2516 3317 2520
rect 3321 2512 3325 2520
rect 3334 2512 3338 2520
rect 3342 2512 3346 2520
rect 3350 2512 3354 2520
rect 3358 2512 3362 2520
rect 3371 2512 3375 2520
rect 3379 2512 3383 2520
rect 3387 2516 3391 2520
rect 3395 2512 3399 2520
rect 3408 2512 3412 2520
rect 3421 2512 3425 2520
rect 3429 2512 3433 2520
rect 3437 2512 3441 2520
rect 3445 2516 3449 2520
rect 3453 2512 3457 2520
rect 3466 2512 3470 2520
rect 3474 2512 3478 2520
rect 3482 2512 3486 2520
rect 3490 2512 3494 2520
rect 3503 2512 3507 2520
rect 3511 2512 3515 2520
rect 3519 2516 3523 2520
rect 3527 2512 3531 2520
rect 3540 2512 3544 2520
rect 3553 2512 3557 2520
rect 3561 2512 3565 2520
rect 3569 2512 3573 2520
rect 3577 2516 3581 2520
rect 3585 2512 3589 2520
rect 3598 2512 3602 2520
rect 3606 2512 3610 2520
rect 3614 2512 3618 2520
rect 2770 2481 2774 2489
rect 2778 2481 2782 2489
rect 2786 2481 2790 2489
rect 2794 2481 2798 2489
rect 2802 2481 2806 2489
rect 2810 2481 2814 2489
rect 2821 2481 2825 2489
rect 2838 2481 2842 2489
rect 2855 2481 2859 2489
rect 2864 2481 2868 2489
rect 2877 2481 2881 2489
rect 2885 2481 2889 2489
rect 2893 2481 2897 2489
rect 2910 2481 2914 2489
rect 2920 2481 2924 2489
rect 2928 2481 2932 2489
rect 2968 2476 2972 2484
rect 2983 2476 2987 2484
rect 3004 2481 3008 2489
rect 3012 2481 3016 2489
rect 3022 2481 3026 2489
rect 3030 2481 3034 2489
rect 3039 2481 3043 2489
rect 3047 2481 3051 2489
rect 3055 2481 3059 2489
rect 3063 2481 3067 2489
rect 3071 2481 3075 2489
rect 3082 2481 3086 2489
rect 3099 2481 3103 2489
rect 3116 2481 3120 2489
rect 3125 2481 3129 2489
rect 3138 2481 3142 2489
rect 3146 2481 3150 2489
rect 3154 2481 3158 2489
rect 3171 2481 3175 2489
rect 3181 2481 3185 2489
rect 3189 2481 3193 2489
rect 3715 2481 3719 2489
rect 3723 2481 3727 2489
rect 3731 2481 3735 2489
rect 3739 2481 3743 2489
rect 3747 2481 3751 2489
rect 3755 2481 3759 2489
rect 3766 2481 3770 2489
rect 3783 2481 3787 2489
rect 3800 2481 3804 2489
rect 3809 2481 3813 2489
rect 3822 2481 3826 2489
rect 3830 2481 3834 2489
rect 3838 2481 3842 2489
rect 3855 2481 3859 2489
rect 3865 2481 3869 2489
rect 3873 2481 3877 2489
rect 3913 2476 3917 2484
rect 3928 2476 3932 2484
rect 3949 2481 3953 2489
rect 3957 2481 3961 2489
rect 3967 2481 3971 2489
rect 3975 2481 3979 2489
rect 3984 2481 3988 2489
rect 3992 2481 3996 2489
rect 4000 2481 4004 2489
rect 4008 2481 4012 2489
rect 4016 2481 4020 2489
rect 4027 2481 4031 2489
rect 4044 2481 4048 2489
rect 4061 2481 4065 2489
rect 4070 2481 4074 2489
rect 4083 2481 4087 2489
rect 4091 2481 4095 2489
rect 4099 2481 4103 2489
rect 4116 2481 4120 2489
rect 4126 2481 4130 2489
rect 4134 2481 4138 2489
rect 3064 2400 3068 2408
rect 3077 2400 3081 2408
rect 3085 2400 3089 2408
rect 3093 2404 3097 2408
rect 3101 2400 3105 2408
rect 3114 2400 3118 2408
rect 3127 2400 3131 2408
rect 3135 2400 3139 2408
rect 3143 2400 3147 2408
rect 3151 2404 3155 2408
rect 3159 2400 3163 2408
rect 3172 2400 3176 2408
rect 3180 2400 3184 2408
rect 3188 2400 3192 2408
rect 4009 2400 4013 2408
rect 4022 2400 4026 2408
rect 4030 2400 4034 2408
rect 4038 2404 4042 2408
rect 4046 2400 4050 2408
rect 4059 2400 4063 2408
rect 4072 2400 4076 2408
rect 4080 2400 4084 2408
rect 4088 2400 4092 2408
rect 4096 2404 4100 2408
rect 4104 2400 4108 2408
rect 4117 2400 4121 2408
rect 4125 2400 4129 2408
rect 4133 2400 4137 2408
rect 2281 2370 2285 2378
rect 2294 2370 2298 2378
rect 2302 2370 2306 2378
rect 2310 2374 2314 2378
rect 2318 2370 2322 2378
rect 2331 2370 2335 2378
rect 2344 2370 2348 2378
rect 2352 2370 2356 2378
rect 2360 2370 2364 2378
rect 2368 2374 2372 2378
rect 2376 2370 2380 2378
rect 2389 2370 2393 2378
rect 2397 2370 2401 2378
rect 2405 2370 2409 2378
rect 2413 2370 2417 2378
rect 2426 2370 2430 2378
rect 2434 2370 2438 2378
rect 2442 2374 2446 2378
rect 2450 2370 2454 2378
rect 2463 2370 2467 2378
rect 2476 2370 2480 2378
rect 2484 2370 2488 2378
rect 2492 2370 2496 2378
rect 2500 2374 2504 2378
rect 2508 2370 2512 2378
rect 2521 2370 2525 2378
rect 2529 2370 2533 2378
rect 2537 2370 2541 2378
rect 2545 2370 2549 2378
rect 2558 2370 2562 2378
rect 2566 2370 2570 2378
rect 2574 2374 2578 2378
rect 2582 2370 2586 2378
rect 2595 2370 2599 2378
rect 2608 2370 2612 2378
rect 2616 2370 2620 2378
rect 2624 2370 2628 2378
rect 2632 2374 2636 2378
rect 2640 2370 2644 2378
rect 2653 2370 2657 2378
rect 2661 2370 2665 2378
rect 2669 2370 2673 2378
rect 3226 2370 3230 2378
rect 3239 2370 3243 2378
rect 3247 2370 3251 2378
rect 3255 2374 3259 2378
rect 3263 2370 3267 2378
rect 3276 2370 3280 2378
rect 3289 2370 3293 2378
rect 3297 2370 3301 2378
rect 3305 2370 3309 2378
rect 3313 2374 3317 2378
rect 3321 2370 3325 2378
rect 3334 2370 3338 2378
rect 3342 2370 3346 2378
rect 3350 2370 3354 2378
rect 3358 2370 3362 2378
rect 3371 2370 3375 2378
rect 3379 2370 3383 2378
rect 3387 2374 3391 2378
rect 3395 2370 3399 2378
rect 3408 2370 3412 2378
rect 3421 2370 3425 2378
rect 3429 2370 3433 2378
rect 3437 2370 3441 2378
rect 3445 2374 3449 2378
rect 3453 2370 3457 2378
rect 3466 2370 3470 2378
rect 3474 2370 3478 2378
rect 3482 2370 3486 2378
rect 3490 2370 3494 2378
rect 3503 2370 3507 2378
rect 3511 2370 3515 2378
rect 3519 2374 3523 2378
rect 3527 2370 3531 2378
rect 3540 2370 3544 2378
rect 3553 2370 3557 2378
rect 3561 2370 3565 2378
rect 3569 2370 3573 2378
rect 3577 2374 3581 2378
rect 3585 2370 3589 2378
rect 3598 2370 3602 2378
rect 3606 2370 3610 2378
rect 3614 2370 3618 2378
rect 3064 2314 3068 2322
rect 3077 2314 3081 2322
rect 3085 2314 3089 2322
rect 3093 2318 3097 2322
rect 3101 2314 3105 2322
rect 3114 2314 3118 2322
rect 3127 2314 3131 2322
rect 3135 2314 3139 2322
rect 3143 2314 3147 2322
rect 3151 2318 3155 2322
rect 3159 2314 3163 2322
rect 3172 2314 3176 2322
rect 3180 2314 3184 2322
rect 3188 2314 3192 2322
rect 4009 2314 4013 2322
rect 4022 2314 4026 2322
rect 4030 2314 4034 2322
rect 4038 2318 4042 2322
rect 4046 2314 4050 2322
rect 4059 2314 4063 2322
rect 4072 2314 4076 2322
rect 4080 2314 4084 2322
rect 4088 2314 4092 2322
rect 4096 2318 4100 2322
rect 4104 2314 4108 2322
rect 4117 2314 4121 2322
rect 4125 2314 4129 2322
rect 4133 2314 4137 2322
rect 2281 2284 2285 2292
rect 2294 2284 2298 2292
rect 2302 2284 2306 2292
rect 2310 2288 2314 2292
rect 2318 2284 2322 2292
rect 2331 2284 2335 2292
rect 2344 2284 2348 2292
rect 2352 2284 2356 2292
rect 2360 2284 2364 2292
rect 2368 2288 2372 2292
rect 2376 2284 2380 2292
rect 2389 2284 2393 2292
rect 2397 2284 2401 2292
rect 2405 2284 2409 2292
rect 2413 2284 2417 2292
rect 2426 2284 2430 2292
rect 2434 2284 2438 2292
rect 2442 2288 2446 2292
rect 2450 2284 2454 2292
rect 2463 2284 2467 2292
rect 2476 2284 2480 2292
rect 2484 2284 2488 2292
rect 2492 2284 2496 2292
rect 2500 2288 2504 2292
rect 2508 2284 2512 2292
rect 2521 2284 2525 2292
rect 2529 2284 2533 2292
rect 2537 2284 2541 2292
rect 2545 2284 2549 2292
rect 2558 2284 2562 2292
rect 2566 2284 2570 2292
rect 2574 2288 2578 2292
rect 2582 2284 2586 2292
rect 2595 2284 2599 2292
rect 2608 2284 2612 2292
rect 2616 2284 2620 2292
rect 2624 2284 2628 2292
rect 2632 2288 2636 2292
rect 2640 2284 2644 2292
rect 2653 2284 2657 2292
rect 2661 2284 2665 2292
rect 2669 2284 2673 2292
rect 3226 2284 3230 2292
rect 3239 2284 3243 2292
rect 3247 2284 3251 2292
rect 3255 2288 3259 2292
rect 3263 2284 3267 2292
rect 3276 2284 3280 2292
rect 3289 2284 3293 2292
rect 3297 2284 3301 2292
rect 3305 2284 3309 2292
rect 3313 2288 3317 2292
rect 3321 2284 3325 2292
rect 3334 2284 3338 2292
rect 3342 2284 3346 2292
rect 3350 2284 3354 2292
rect 3358 2284 3362 2292
rect 3371 2284 3375 2292
rect 3379 2284 3383 2292
rect 3387 2288 3391 2292
rect 3395 2284 3399 2292
rect 3408 2284 3412 2292
rect 3421 2284 3425 2292
rect 3429 2284 3433 2292
rect 3437 2284 3441 2292
rect 3445 2288 3449 2292
rect 3453 2284 3457 2292
rect 3466 2284 3470 2292
rect 3474 2284 3478 2292
rect 3482 2284 3486 2292
rect 3490 2284 3494 2292
rect 3503 2284 3507 2292
rect 3511 2284 3515 2292
rect 3519 2288 3523 2292
rect 3527 2284 3531 2292
rect 3540 2284 3544 2292
rect 3553 2284 3557 2292
rect 3561 2284 3565 2292
rect 3569 2284 3573 2292
rect 3577 2288 3581 2292
rect 3585 2284 3589 2292
rect 3598 2284 3602 2292
rect 3606 2284 3610 2292
rect 3614 2284 3618 2292
rect 2281 2144 2285 2152
rect 2294 2144 2298 2152
rect 2302 2144 2306 2152
rect 2310 2148 2314 2152
rect 2318 2144 2322 2152
rect 2331 2144 2335 2152
rect 2344 2144 2348 2152
rect 2352 2144 2356 2152
rect 2360 2144 2364 2152
rect 2368 2148 2372 2152
rect 2376 2144 2380 2152
rect 2389 2144 2393 2152
rect 2397 2144 2401 2152
rect 2405 2144 2409 2152
rect 2413 2144 2417 2152
rect 2426 2144 2430 2152
rect 2434 2144 2438 2152
rect 2442 2148 2446 2152
rect 2450 2144 2454 2152
rect 2463 2144 2467 2152
rect 2476 2144 2480 2152
rect 2484 2144 2488 2152
rect 2492 2144 2496 2152
rect 2500 2148 2504 2152
rect 2508 2144 2512 2152
rect 2521 2144 2525 2152
rect 2529 2144 2533 2152
rect 2537 2144 2541 2152
rect 2545 2144 2549 2152
rect 2558 2144 2562 2152
rect 2566 2144 2570 2152
rect 2574 2148 2578 2152
rect 2582 2144 2586 2152
rect 2595 2144 2599 2152
rect 2608 2144 2612 2152
rect 2616 2144 2620 2152
rect 2624 2144 2628 2152
rect 2632 2148 2636 2152
rect 2640 2144 2644 2152
rect 2653 2144 2657 2152
rect 2661 2144 2665 2152
rect 2669 2144 2673 2152
rect 3226 2144 3230 2152
rect 3239 2144 3243 2152
rect 3247 2144 3251 2152
rect 3255 2148 3259 2152
rect 3263 2144 3267 2152
rect 3276 2144 3280 2152
rect 3289 2144 3293 2152
rect 3297 2144 3301 2152
rect 3305 2144 3309 2152
rect 3313 2148 3317 2152
rect 3321 2144 3325 2152
rect 3334 2144 3338 2152
rect 3342 2144 3346 2152
rect 3350 2144 3354 2152
rect 3358 2144 3362 2152
rect 3371 2144 3375 2152
rect 3379 2144 3383 2152
rect 3387 2148 3391 2152
rect 3395 2144 3399 2152
rect 3408 2144 3412 2152
rect 3421 2144 3425 2152
rect 3429 2144 3433 2152
rect 3437 2144 3441 2152
rect 3445 2148 3449 2152
rect 3453 2144 3457 2152
rect 3466 2144 3470 2152
rect 3474 2144 3478 2152
rect 3482 2144 3486 2152
rect 3490 2144 3494 2152
rect 3503 2144 3507 2152
rect 3511 2144 3515 2152
rect 3519 2148 3523 2152
rect 3527 2144 3531 2152
rect 3540 2144 3544 2152
rect 3553 2144 3557 2152
rect 3561 2144 3565 2152
rect 3569 2144 3573 2152
rect 3577 2148 3581 2152
rect 3585 2144 3589 2152
rect 3598 2144 3602 2152
rect 3606 2144 3610 2152
rect 3614 2144 3618 2152
<< psubstratepcontact >>
rect 2795 3990 2799 3994
rect 2823 3990 2827 3994
rect 2853 3990 2857 3994
rect 2927 3990 2931 3994
rect 2955 3990 2959 3994
rect 2985 3990 2989 3994
rect 3059 3990 3063 3994
rect 3087 3990 3091 3994
rect 3117 3990 3121 3994
rect 3191 3990 3195 3994
rect 3219 3990 3223 3994
rect 3249 3990 3253 3994
rect 3740 3990 3744 3994
rect 3768 3990 3772 3994
rect 3798 3990 3802 3994
rect 3872 3990 3876 3994
rect 3900 3990 3904 3994
rect 3930 3990 3934 3994
rect 4004 3990 4008 3994
rect 4032 3990 4036 3994
rect 4062 3990 4066 3994
rect 4136 3990 4140 3994
rect 4164 3990 4168 3994
rect 4194 3990 4198 3994
rect 2443 3957 2447 3961
rect 2471 3957 2475 3961
rect 2501 3957 2505 3961
rect 3388 3957 3392 3961
rect 3416 3957 3420 3961
rect 3446 3957 3450 3961
rect 2776 3904 2780 3908
rect 2811 3904 2815 3908
rect 2937 3904 2941 3908
rect 2961 3904 2965 3908
rect 3015 3904 3022 3908
rect 3042 3904 3046 3908
rect 3096 3904 3100 3908
rect 3721 3904 3725 3908
rect 3756 3904 3760 3908
rect 3882 3904 3886 3908
rect 3906 3904 3910 3908
rect 3960 3904 3967 3908
rect 3987 3904 3991 3908
rect 4041 3904 4045 3908
rect 2440 3855 2444 3859
rect 2470 3855 2474 3859
rect 2498 3855 2502 3859
rect 3385 3855 3389 3859
rect 3415 3855 3419 3859
rect 3443 3855 3447 3859
rect 2776 3772 2780 3776
rect 2811 3772 2815 3776
rect 2937 3772 2941 3776
rect 2961 3772 2965 3776
rect 3015 3772 3019 3776
rect 3042 3772 3046 3776
rect 3066 3772 3070 3776
rect 3721 3772 3725 3776
rect 3756 3772 3760 3776
rect 3882 3772 3886 3776
rect 3906 3772 3910 3776
rect 3960 3772 3964 3776
rect 3987 3772 3991 3776
rect 4011 3772 4015 3776
rect 3273 3729 3277 3733
rect 3297 3729 3301 3733
rect 3351 3729 3355 3733
rect 3494 3729 3498 3733
rect 2776 3640 2780 3644
rect 2811 3640 2815 3644
rect 2937 3640 2941 3644
rect 2961 3640 2965 3644
rect 3015 3640 3022 3644
rect 3042 3640 3046 3644
rect 3096 3640 3100 3644
rect 3132 3640 3136 3644
rect 3186 3640 3190 3644
rect 3721 3640 3725 3644
rect 3756 3640 3760 3644
rect 3882 3640 3886 3644
rect 3906 3640 3910 3644
rect 3960 3640 3967 3644
rect 3987 3640 3991 3644
rect 4041 3640 4045 3644
rect 4077 3640 4081 3644
rect 4131 3640 4135 3644
rect 3251 3599 3255 3603
rect 3273 3599 3277 3603
rect 3297 3599 3301 3603
rect 3351 3599 3355 3603
rect 3400 3599 3404 3603
rect 2776 3508 2780 3512
rect 2811 3508 2815 3512
rect 2937 3508 2941 3512
rect 2961 3508 2965 3512
rect 3072 3508 3076 3512
rect 3721 3508 3725 3512
rect 3756 3508 3760 3512
rect 3882 3508 3886 3512
rect 3906 3508 3910 3512
rect 4017 3508 4021 3512
rect 2311 3455 2315 3459
rect 2339 3455 2343 3459
rect 2369 3455 2373 3459
rect 2443 3455 2447 3459
rect 2471 3455 2475 3459
rect 2501 3455 2505 3459
rect 2575 3455 2579 3459
rect 2603 3455 2607 3459
rect 2633 3455 2637 3459
rect 3256 3455 3260 3459
rect 3284 3455 3288 3459
rect 3314 3455 3318 3459
rect 3388 3455 3392 3459
rect 3416 3455 3420 3459
rect 3446 3455 3450 3459
rect 3520 3455 3524 3459
rect 3548 3455 3552 3459
rect 3578 3455 3582 3459
rect 3094 3343 3098 3347
rect 3122 3343 3126 3347
rect 3152 3343 3156 3347
rect 4039 3343 4043 3347
rect 4067 3343 4071 3347
rect 4097 3343 4101 3347
rect 2311 3313 2315 3317
rect 2339 3313 2343 3317
rect 2369 3313 2373 3317
rect 2443 3313 2447 3317
rect 2471 3313 2475 3317
rect 2501 3313 2505 3317
rect 2575 3313 2579 3317
rect 2603 3313 2607 3317
rect 2633 3313 2637 3317
rect 3256 3313 3260 3317
rect 3284 3313 3288 3317
rect 3314 3313 3318 3317
rect 3388 3313 3392 3317
rect 3416 3313 3420 3317
rect 3446 3313 3450 3317
rect 3520 3313 3524 3317
rect 3548 3313 3552 3317
rect 3578 3313 3582 3317
rect 3094 3257 3098 3261
rect 3122 3257 3126 3261
rect 3152 3257 3156 3261
rect 4039 3257 4043 3261
rect 4067 3257 4071 3261
rect 4097 3257 4101 3261
rect 2311 3227 2315 3231
rect 2339 3227 2343 3231
rect 2369 3227 2373 3231
rect 2443 3227 2447 3231
rect 2471 3227 2475 3231
rect 2501 3227 2505 3231
rect 2575 3227 2579 3231
rect 2603 3227 2607 3231
rect 2633 3227 2637 3231
rect 3256 3227 3260 3231
rect 3284 3227 3288 3231
rect 3314 3227 3318 3231
rect 3388 3227 3392 3231
rect 3416 3227 3420 3231
rect 3446 3227 3450 3231
rect 3520 3227 3524 3231
rect 3548 3227 3552 3231
rect 3578 3227 3582 3231
rect 2311 3087 2315 3091
rect 2339 3087 2343 3091
rect 2369 3087 2373 3091
rect 2443 3087 2447 3091
rect 2471 3087 2475 3091
rect 2501 3087 2505 3091
rect 2575 3087 2579 3091
rect 2603 3087 2607 3091
rect 2633 3087 2637 3091
rect 3256 3087 3260 3091
rect 3284 3087 3288 3091
rect 3314 3087 3318 3091
rect 3388 3087 3392 3091
rect 3416 3087 3420 3091
rect 3446 3087 3450 3091
rect 3520 3087 3524 3091
rect 3548 3087 3552 3091
rect 3578 3087 3582 3091
rect 2795 3008 2799 3012
rect 2823 3008 2827 3012
rect 2853 3008 2857 3012
rect 2927 3008 2931 3012
rect 2955 3008 2959 3012
rect 2985 3008 2989 3012
rect 3059 3008 3063 3012
rect 3087 3008 3091 3012
rect 3117 3008 3121 3012
rect 3191 3008 3195 3012
rect 3219 3008 3223 3012
rect 3249 3008 3253 3012
rect 3740 3008 3744 3012
rect 3768 3008 3772 3012
rect 3798 3008 3802 3012
rect 3872 3008 3876 3012
rect 3900 3008 3904 3012
rect 3930 3008 3934 3012
rect 4004 3008 4008 3012
rect 4032 3008 4036 3012
rect 4062 3008 4066 3012
rect 4136 3008 4140 3012
rect 4164 3008 4168 3012
rect 4194 3008 4198 3012
rect 2443 2975 2447 2979
rect 2471 2975 2475 2979
rect 2501 2975 2505 2979
rect 3388 2975 3392 2979
rect 3416 2975 3420 2979
rect 3446 2975 3450 2979
rect 2776 2922 2780 2926
rect 2811 2922 2815 2926
rect 2937 2922 2941 2926
rect 2961 2922 2965 2926
rect 3015 2922 3022 2926
rect 3042 2922 3046 2926
rect 3096 2922 3100 2926
rect 3721 2922 3725 2926
rect 3756 2922 3760 2926
rect 3882 2922 3886 2926
rect 3906 2922 3910 2926
rect 3960 2922 3967 2926
rect 3987 2922 3991 2926
rect 4041 2922 4045 2926
rect 2440 2873 2444 2877
rect 2470 2873 2474 2877
rect 2498 2873 2502 2877
rect 3385 2873 3389 2877
rect 3415 2873 3419 2877
rect 3443 2873 3447 2877
rect 2776 2790 2780 2794
rect 2811 2790 2815 2794
rect 2937 2790 2941 2794
rect 2961 2790 2965 2794
rect 3015 2790 3019 2794
rect 3042 2790 3046 2794
rect 3066 2790 3070 2794
rect 3721 2790 3725 2794
rect 3756 2790 3760 2794
rect 3882 2790 3886 2794
rect 3906 2790 3910 2794
rect 3960 2790 3964 2794
rect 3987 2790 3991 2794
rect 4011 2790 4015 2794
rect 2776 2658 2780 2662
rect 2811 2658 2815 2662
rect 2937 2658 2941 2662
rect 2961 2658 2965 2662
rect 3015 2658 3022 2662
rect 3042 2658 3046 2662
rect 3096 2658 3100 2662
rect 3132 2658 3136 2662
rect 3186 2658 3190 2662
rect 3721 2658 3725 2662
rect 3756 2658 3760 2662
rect 3882 2658 3886 2662
rect 3906 2658 3910 2662
rect 3960 2658 3967 2662
rect 3987 2658 3991 2662
rect 4041 2658 4045 2662
rect 4077 2658 4081 2662
rect 4131 2658 4135 2662
rect 2776 2526 2780 2530
rect 2811 2526 2815 2530
rect 2937 2526 2941 2530
rect 2961 2526 2965 2530
rect 3072 2526 3076 2530
rect 3721 2526 3725 2530
rect 3756 2526 3760 2530
rect 3882 2526 3886 2530
rect 3906 2526 3910 2530
rect 4017 2526 4021 2530
rect 2311 2473 2315 2477
rect 2339 2473 2343 2477
rect 2369 2473 2373 2477
rect 2443 2473 2447 2477
rect 2471 2473 2475 2477
rect 2501 2473 2505 2477
rect 2575 2473 2579 2477
rect 2603 2473 2607 2477
rect 2633 2473 2637 2477
rect 3256 2473 3260 2477
rect 3284 2473 3288 2477
rect 3314 2473 3318 2477
rect 3388 2473 3392 2477
rect 3416 2473 3420 2477
rect 3446 2473 3450 2477
rect 3520 2473 3524 2477
rect 3548 2473 3552 2477
rect 3578 2473 3582 2477
rect 3094 2361 3098 2365
rect 3122 2361 3126 2365
rect 3152 2361 3156 2365
rect 4039 2361 4043 2365
rect 4067 2361 4071 2365
rect 4097 2361 4101 2365
rect 2311 2331 2315 2335
rect 2339 2331 2343 2335
rect 2369 2331 2373 2335
rect 2443 2331 2447 2335
rect 2471 2331 2475 2335
rect 2501 2331 2505 2335
rect 2575 2331 2579 2335
rect 2603 2331 2607 2335
rect 2633 2331 2637 2335
rect 3256 2331 3260 2335
rect 3284 2331 3288 2335
rect 3314 2331 3318 2335
rect 3388 2331 3392 2335
rect 3416 2331 3420 2335
rect 3446 2331 3450 2335
rect 3520 2331 3524 2335
rect 3548 2331 3552 2335
rect 3578 2331 3582 2335
rect 3094 2275 3098 2279
rect 3122 2275 3126 2279
rect 3152 2275 3156 2279
rect 4039 2275 4043 2279
rect 4067 2275 4071 2279
rect 4097 2275 4101 2279
rect 2311 2245 2315 2249
rect 2339 2245 2343 2249
rect 2369 2245 2373 2249
rect 2443 2245 2447 2249
rect 2471 2245 2475 2249
rect 2501 2245 2505 2249
rect 2575 2245 2579 2249
rect 2603 2245 2607 2249
rect 2633 2245 2637 2249
rect 3256 2245 3260 2249
rect 3284 2245 3288 2249
rect 3314 2245 3318 2249
rect 3388 2245 3392 2249
rect 3416 2245 3420 2249
rect 3446 2245 3450 2249
rect 3520 2245 3524 2249
rect 3548 2245 3552 2249
rect 3578 2245 3582 2249
rect 2311 2105 2315 2109
rect 2339 2105 2343 2109
rect 2369 2105 2373 2109
rect 2443 2105 2447 2109
rect 2471 2105 2475 2109
rect 2501 2105 2505 2109
rect 2575 2105 2579 2109
rect 2603 2105 2607 2109
rect 2633 2105 2637 2109
rect 3256 2105 3260 2109
rect 3284 2105 3288 2109
rect 3314 2105 3318 2109
rect 3388 2105 3392 2109
rect 3416 2105 3420 2109
rect 3446 2105 3450 2109
rect 3520 2105 3524 2109
rect 3548 2105 3552 2109
rect 3578 2105 3582 2109
<< nsubstratencontact >>
rect 2795 4047 2799 4051
rect 2823 4047 2827 4051
rect 2853 4047 2857 4051
rect 2890 4047 2894 4051
rect 2927 4047 2931 4051
rect 2955 4047 2959 4051
rect 2985 4047 2989 4051
rect 3022 4047 3026 4051
rect 3059 4047 3063 4051
rect 3087 4047 3091 4051
rect 3117 4047 3121 4051
rect 3154 4047 3158 4051
rect 3191 4047 3195 4051
rect 3219 4047 3223 4051
rect 3249 4047 3253 4051
rect 3286 4047 3290 4051
rect 3740 4047 3744 4051
rect 3768 4047 3772 4051
rect 3798 4047 3802 4051
rect 3835 4047 3839 4051
rect 3872 4047 3876 4051
rect 3900 4047 3904 4051
rect 3930 4047 3934 4051
rect 3967 4047 3971 4051
rect 4004 4047 4008 4051
rect 4032 4047 4036 4051
rect 4062 4047 4066 4051
rect 4099 4047 4103 4051
rect 4136 4047 4140 4051
rect 4164 4047 4168 4051
rect 4194 4047 4198 4051
rect 4231 4047 4235 4051
rect 2443 4014 2447 4018
rect 2471 4014 2475 4018
rect 2501 4014 2505 4018
rect 2538 4014 2542 4018
rect 3388 4014 3392 4018
rect 3416 4014 3420 4018
rect 3446 4014 3450 4018
rect 3483 4014 3487 4018
rect 2785 3970 2789 3974
rect 2814 3970 2818 3974
rect 2839 3970 2843 3974
rect 2881 3970 2885 3974
rect 2937 3970 2941 3974
rect 2961 3970 2965 3974
rect 3015 3970 3019 3974
rect 3042 3970 3046 3974
rect 3096 3970 3100 3974
rect 3730 3970 3734 3974
rect 3759 3970 3763 3974
rect 3784 3970 3788 3974
rect 3826 3970 3830 3974
rect 3882 3970 3886 3974
rect 3906 3970 3910 3974
rect 3960 3970 3964 3974
rect 3987 3970 3991 3974
rect 4041 3970 4045 3974
rect 2403 3912 2407 3916
rect 2440 3912 2444 3916
rect 2470 3912 2474 3916
rect 2498 3912 2502 3916
rect 3348 3912 3352 3916
rect 3385 3912 3389 3916
rect 3415 3912 3419 3916
rect 3443 3912 3447 3916
rect 2785 3838 2789 3842
rect 2814 3838 2818 3842
rect 2839 3838 2843 3842
rect 2881 3838 2885 3842
rect 2937 3838 2941 3842
rect 2961 3838 2965 3842
rect 3015 3838 3019 3842
rect 3042 3838 3046 3842
rect 3104 3838 3108 3842
rect 3730 3838 3734 3842
rect 3759 3838 3763 3842
rect 3784 3838 3788 3842
rect 3826 3838 3830 3842
rect 3882 3838 3886 3842
rect 3906 3838 3910 3842
rect 3960 3838 3964 3842
rect 3987 3838 3991 3842
rect 4049 3838 4053 3842
rect 3273 3809 3277 3813
rect 3297 3809 3301 3813
rect 3351 3809 3355 3813
rect 3494 3809 3498 3813
rect 2785 3706 2789 3710
rect 2814 3706 2818 3710
rect 2839 3706 2843 3710
rect 2881 3706 2885 3710
rect 2937 3706 2941 3710
rect 2961 3706 2965 3710
rect 3015 3706 3019 3710
rect 3042 3706 3046 3710
rect 3096 3706 3100 3710
rect 3104 3706 3108 3710
rect 3132 3706 3136 3710
rect 3186 3706 3190 3710
rect 3730 3706 3734 3710
rect 3759 3706 3763 3710
rect 3784 3706 3788 3710
rect 3826 3706 3830 3710
rect 3882 3706 3886 3710
rect 3906 3706 3910 3710
rect 3960 3706 3964 3710
rect 3987 3706 3991 3710
rect 4041 3706 4045 3710
rect 4049 3706 4053 3710
rect 4077 3706 4081 3710
rect 4131 3706 4135 3710
rect 3251 3679 3255 3683
rect 3273 3679 3277 3683
rect 3297 3679 3301 3683
rect 3351 3679 3355 3683
rect 3400 3679 3404 3683
rect 2785 3574 2789 3578
rect 2814 3574 2818 3578
rect 2839 3574 2843 3578
rect 2881 3574 2885 3578
rect 2937 3574 2941 3578
rect 2961 3574 2965 3578
rect 3015 3574 3019 3578
rect 3042 3574 3046 3578
rect 3132 3574 3136 3578
rect 3730 3574 3734 3578
rect 3759 3574 3763 3578
rect 3784 3574 3788 3578
rect 3826 3574 3830 3578
rect 3882 3574 3886 3578
rect 3906 3574 3910 3578
rect 3960 3574 3964 3578
rect 3987 3574 3991 3578
rect 4077 3574 4081 3578
rect 3297 3549 3301 3553
rect 2311 3512 2315 3516
rect 2339 3512 2343 3516
rect 2369 3512 2373 3516
rect 2406 3512 2410 3516
rect 2443 3512 2447 3516
rect 2471 3512 2475 3516
rect 2501 3512 2505 3516
rect 2538 3512 2542 3516
rect 2575 3512 2579 3516
rect 2603 3512 2607 3516
rect 2633 3512 2637 3516
rect 2670 3512 2674 3516
rect 3256 3512 3260 3516
rect 3284 3512 3288 3516
rect 3314 3512 3318 3516
rect 3351 3512 3355 3516
rect 3388 3512 3392 3516
rect 3416 3512 3420 3516
rect 3446 3512 3450 3516
rect 3483 3512 3487 3516
rect 3520 3512 3524 3516
rect 3548 3512 3552 3516
rect 3578 3512 3582 3516
rect 3615 3512 3619 3516
rect 2785 3442 2789 3446
rect 2814 3442 2818 3446
rect 2839 3442 2843 3446
rect 2881 3442 2885 3446
rect 2961 3442 2965 3446
rect 3015 3442 3019 3446
rect 3046 3442 3050 3446
rect 3075 3442 3079 3446
rect 3100 3442 3104 3446
rect 3142 3442 3146 3446
rect 3730 3442 3734 3446
rect 3759 3442 3763 3446
rect 3784 3442 3788 3446
rect 3826 3442 3830 3446
rect 3906 3442 3910 3446
rect 3960 3442 3964 3446
rect 3991 3442 3995 3446
rect 4020 3442 4024 3446
rect 4045 3442 4049 3446
rect 4087 3442 4091 3446
rect 3094 3400 3098 3404
rect 3122 3400 3126 3404
rect 3152 3400 3156 3404
rect 3189 3400 3193 3404
rect 4039 3400 4043 3404
rect 4067 3400 4071 3404
rect 4097 3400 4101 3404
rect 4134 3400 4138 3404
rect 2311 3370 2315 3374
rect 2339 3370 2343 3374
rect 2369 3370 2373 3374
rect 2406 3370 2410 3374
rect 2443 3370 2447 3374
rect 2471 3370 2475 3374
rect 2501 3370 2505 3374
rect 2538 3370 2542 3374
rect 2575 3370 2579 3374
rect 2603 3370 2607 3374
rect 2633 3370 2637 3374
rect 2670 3370 2674 3374
rect 3256 3370 3260 3374
rect 3284 3370 3288 3374
rect 3314 3370 3318 3374
rect 3351 3370 3355 3374
rect 3388 3370 3392 3374
rect 3416 3370 3420 3374
rect 3446 3370 3450 3374
rect 3483 3370 3487 3374
rect 3520 3370 3524 3374
rect 3548 3370 3552 3374
rect 3578 3370 3582 3374
rect 3615 3370 3619 3374
rect 3094 3314 3098 3318
rect 3122 3314 3126 3318
rect 3152 3314 3156 3318
rect 3189 3314 3193 3318
rect 4039 3314 4043 3318
rect 4067 3314 4071 3318
rect 4097 3314 4101 3318
rect 4134 3314 4138 3318
rect 2311 3284 2315 3288
rect 2339 3284 2343 3288
rect 2369 3284 2373 3288
rect 2406 3284 2410 3288
rect 2443 3284 2447 3288
rect 2471 3284 2475 3288
rect 2501 3284 2505 3288
rect 2538 3284 2542 3288
rect 2575 3284 2579 3288
rect 2603 3284 2607 3288
rect 2633 3284 2637 3288
rect 2670 3284 2674 3288
rect 3256 3284 3260 3288
rect 3284 3284 3288 3288
rect 3314 3284 3318 3288
rect 3351 3284 3355 3288
rect 3388 3284 3392 3288
rect 3416 3284 3420 3288
rect 3446 3284 3450 3288
rect 3483 3284 3487 3288
rect 3520 3284 3524 3288
rect 3548 3284 3552 3288
rect 3578 3284 3582 3288
rect 3615 3284 3619 3288
rect 2311 3144 2315 3148
rect 2339 3144 2343 3148
rect 2369 3144 2373 3148
rect 2406 3144 2410 3148
rect 2443 3144 2447 3148
rect 2471 3144 2475 3148
rect 2501 3144 2505 3148
rect 2538 3144 2542 3148
rect 2575 3144 2579 3148
rect 2603 3144 2607 3148
rect 2633 3144 2637 3148
rect 2670 3144 2674 3148
rect 3256 3144 3260 3148
rect 3284 3144 3288 3148
rect 3314 3144 3318 3148
rect 3351 3144 3355 3148
rect 3388 3144 3392 3148
rect 3416 3144 3420 3148
rect 3446 3144 3450 3148
rect 3483 3144 3487 3148
rect 3520 3144 3524 3148
rect 3548 3144 3552 3148
rect 3578 3144 3582 3148
rect 3615 3144 3619 3148
rect 2795 3065 2799 3069
rect 2823 3065 2827 3069
rect 2853 3065 2857 3069
rect 2890 3065 2894 3069
rect 2927 3065 2931 3069
rect 2955 3065 2959 3069
rect 2985 3065 2989 3069
rect 3022 3065 3026 3069
rect 3059 3065 3063 3069
rect 3087 3065 3091 3069
rect 3117 3065 3121 3069
rect 3154 3065 3158 3069
rect 3191 3065 3195 3069
rect 3219 3065 3223 3069
rect 3249 3065 3253 3069
rect 3286 3065 3290 3069
rect 3740 3065 3744 3069
rect 3768 3065 3772 3069
rect 3798 3065 3802 3069
rect 3835 3065 3839 3069
rect 3872 3065 3876 3069
rect 3900 3065 3904 3069
rect 3930 3065 3934 3069
rect 3967 3065 3971 3069
rect 4004 3065 4008 3069
rect 4032 3065 4036 3069
rect 4062 3065 4066 3069
rect 4099 3065 4103 3069
rect 4136 3065 4140 3069
rect 4164 3065 4168 3069
rect 4194 3065 4198 3069
rect 4231 3065 4235 3069
rect 2443 3032 2447 3036
rect 2471 3032 2475 3036
rect 2501 3032 2505 3036
rect 2538 3032 2542 3036
rect 3388 3032 3392 3036
rect 3416 3032 3420 3036
rect 3446 3032 3450 3036
rect 3483 3032 3487 3036
rect 2785 2988 2789 2992
rect 2814 2988 2818 2992
rect 2839 2988 2843 2992
rect 2881 2988 2885 2992
rect 2937 2988 2941 2992
rect 2961 2988 2965 2992
rect 3015 2988 3019 2992
rect 3042 2988 3046 2992
rect 3096 2988 3100 2992
rect 3730 2988 3734 2992
rect 3759 2988 3763 2992
rect 3784 2988 3788 2992
rect 3826 2988 3830 2992
rect 3882 2988 3886 2992
rect 3906 2988 3910 2992
rect 3960 2988 3964 2992
rect 3987 2988 3991 2992
rect 4041 2988 4045 2992
rect 2403 2930 2407 2934
rect 2440 2930 2444 2934
rect 2470 2930 2474 2934
rect 2498 2930 2502 2934
rect 3348 2930 3352 2934
rect 3385 2930 3389 2934
rect 3415 2930 3419 2934
rect 3443 2930 3447 2934
rect 2785 2856 2789 2860
rect 2814 2856 2818 2860
rect 2839 2856 2843 2860
rect 2881 2856 2885 2860
rect 2937 2856 2941 2860
rect 2961 2856 2965 2860
rect 3015 2856 3019 2860
rect 3042 2856 3046 2860
rect 3104 2856 3108 2860
rect 3730 2856 3734 2860
rect 3759 2856 3763 2860
rect 3784 2856 3788 2860
rect 3826 2856 3830 2860
rect 3882 2856 3886 2860
rect 3906 2856 3910 2860
rect 3960 2856 3964 2860
rect 3987 2856 3991 2860
rect 4049 2856 4053 2860
rect 2785 2724 2789 2728
rect 2814 2724 2818 2728
rect 2839 2724 2843 2728
rect 2881 2724 2885 2728
rect 2937 2724 2941 2728
rect 2961 2724 2965 2728
rect 3015 2724 3019 2728
rect 3042 2724 3046 2728
rect 3096 2724 3100 2728
rect 3104 2724 3108 2728
rect 3132 2724 3136 2728
rect 3186 2724 3190 2728
rect 3730 2724 3734 2728
rect 3759 2724 3763 2728
rect 3784 2724 3788 2728
rect 3826 2724 3830 2728
rect 3882 2724 3886 2728
rect 3906 2724 3910 2728
rect 3960 2724 3964 2728
rect 3987 2724 3991 2728
rect 4041 2724 4045 2728
rect 4049 2724 4053 2728
rect 4077 2724 4081 2728
rect 4131 2724 4135 2728
rect 2785 2592 2789 2596
rect 2814 2592 2818 2596
rect 2839 2592 2843 2596
rect 2881 2592 2885 2596
rect 2937 2592 2941 2596
rect 2961 2592 2965 2596
rect 3015 2592 3019 2596
rect 3042 2592 3046 2596
rect 3132 2592 3136 2596
rect 3730 2592 3734 2596
rect 3759 2592 3763 2596
rect 3784 2592 3788 2596
rect 3826 2592 3830 2596
rect 3882 2592 3886 2596
rect 3906 2592 3910 2596
rect 3960 2592 3964 2596
rect 3987 2592 3991 2596
rect 4077 2592 4081 2596
rect 2311 2530 2315 2534
rect 2339 2530 2343 2534
rect 2369 2530 2373 2534
rect 2406 2530 2410 2534
rect 2443 2530 2447 2534
rect 2471 2530 2475 2534
rect 2501 2530 2505 2534
rect 2538 2530 2542 2534
rect 2575 2530 2579 2534
rect 2603 2530 2607 2534
rect 2633 2530 2637 2534
rect 2670 2530 2674 2534
rect 3256 2530 3260 2534
rect 3284 2530 3288 2534
rect 3314 2530 3318 2534
rect 3351 2530 3355 2534
rect 3388 2530 3392 2534
rect 3416 2530 3420 2534
rect 3446 2530 3450 2534
rect 3483 2530 3487 2534
rect 3520 2530 3524 2534
rect 3548 2530 3552 2534
rect 3578 2530 3582 2534
rect 3615 2530 3619 2534
rect 2785 2460 2789 2464
rect 2814 2460 2818 2464
rect 2839 2460 2843 2464
rect 2881 2460 2885 2464
rect 2961 2460 2965 2464
rect 3015 2460 3019 2464
rect 3046 2460 3050 2464
rect 3075 2460 3079 2464
rect 3100 2460 3104 2464
rect 3142 2460 3146 2464
rect 3730 2460 3734 2464
rect 3759 2460 3763 2464
rect 3784 2460 3788 2464
rect 3826 2460 3830 2464
rect 3906 2460 3910 2464
rect 3960 2460 3964 2464
rect 3991 2460 3995 2464
rect 4020 2460 4024 2464
rect 4045 2460 4049 2464
rect 4087 2460 4091 2464
rect 3094 2418 3098 2422
rect 3122 2418 3126 2422
rect 3152 2418 3156 2422
rect 3189 2418 3193 2422
rect 4039 2418 4043 2422
rect 4067 2418 4071 2422
rect 4097 2418 4101 2422
rect 4134 2418 4138 2422
rect 2311 2388 2315 2392
rect 2339 2388 2343 2392
rect 2369 2388 2373 2392
rect 2406 2388 2410 2392
rect 2443 2388 2447 2392
rect 2471 2388 2475 2392
rect 2501 2388 2505 2392
rect 2538 2388 2542 2392
rect 2575 2388 2579 2392
rect 2603 2388 2607 2392
rect 2633 2388 2637 2392
rect 2670 2388 2674 2392
rect 3256 2388 3260 2392
rect 3284 2388 3288 2392
rect 3314 2388 3318 2392
rect 3351 2388 3355 2392
rect 3388 2388 3392 2392
rect 3416 2388 3420 2392
rect 3446 2388 3450 2392
rect 3483 2388 3487 2392
rect 3520 2388 3524 2392
rect 3548 2388 3552 2392
rect 3578 2388 3582 2392
rect 3615 2388 3619 2392
rect 3094 2332 3098 2336
rect 3122 2332 3126 2336
rect 3152 2332 3156 2336
rect 3189 2332 3193 2336
rect 4039 2332 4043 2336
rect 4067 2332 4071 2336
rect 4097 2332 4101 2336
rect 4134 2332 4138 2336
rect 2311 2302 2315 2306
rect 2339 2302 2343 2306
rect 2369 2302 2373 2306
rect 2406 2302 2410 2306
rect 2443 2302 2447 2306
rect 2471 2302 2475 2306
rect 2501 2302 2505 2306
rect 2538 2302 2542 2306
rect 2575 2302 2579 2306
rect 2603 2302 2607 2306
rect 2633 2302 2637 2306
rect 2670 2302 2674 2306
rect 3256 2302 3260 2306
rect 3284 2302 3288 2306
rect 3314 2302 3318 2306
rect 3351 2302 3355 2306
rect 3388 2302 3392 2306
rect 3416 2302 3420 2306
rect 3446 2302 3450 2306
rect 3483 2302 3487 2306
rect 3520 2302 3524 2306
rect 3548 2302 3552 2306
rect 3578 2302 3582 2306
rect 3615 2302 3619 2306
rect 2311 2162 2315 2166
rect 2339 2162 2343 2166
rect 2369 2162 2373 2166
rect 2406 2162 2410 2166
rect 2443 2162 2447 2166
rect 2471 2162 2475 2166
rect 2501 2162 2505 2166
rect 2538 2162 2542 2166
rect 2575 2162 2579 2166
rect 2603 2162 2607 2166
rect 2633 2162 2637 2166
rect 2670 2162 2674 2166
rect 3256 2162 3260 2166
rect 3284 2162 3288 2166
rect 3314 2162 3318 2166
rect 3351 2162 3355 2166
rect 3388 2162 3392 2166
rect 3416 2162 3420 2166
rect 3446 2162 3450 2166
rect 3483 2162 3487 2166
rect 3520 2162 3524 2166
rect 3548 2162 3552 2166
rect 3578 2162 3582 2166
rect 3615 2162 3619 2166
<< polysilicon >>
rect 2770 4037 2772 4039
rect 2775 4037 2777 4040
rect 2791 4037 2793 4039
rect 2807 4037 2809 4039
rect 2812 4037 2814 4040
rect 2833 4037 2835 4040
rect 2849 4037 2851 4040
rect 2865 4037 2867 4039
rect 2870 4037 2872 4040
rect 2886 4037 2888 4039
rect 2902 4037 2904 4039
rect 2907 4037 2909 4040
rect 2923 4037 2925 4039
rect 2939 4037 2941 4039
rect 2944 4037 2946 4040
rect 2965 4037 2967 4040
rect 2981 4037 2983 4040
rect 2997 4037 2999 4039
rect 3002 4037 3004 4040
rect 3018 4037 3020 4039
rect 3034 4037 3036 4039
rect 3039 4037 3041 4040
rect 3055 4037 3057 4039
rect 3071 4037 3073 4039
rect 3076 4037 3078 4040
rect 3097 4037 3099 4040
rect 3113 4037 3115 4040
rect 3129 4037 3131 4039
rect 3134 4037 3136 4040
rect 3150 4037 3152 4039
rect 3166 4037 3168 4039
rect 3171 4037 3173 4040
rect 3187 4037 3189 4039
rect 3203 4037 3205 4039
rect 3208 4037 3210 4040
rect 3229 4037 3231 4040
rect 3245 4037 3247 4040
rect 3261 4037 3263 4039
rect 3266 4037 3268 4040
rect 3282 4037 3284 4039
rect 3715 4037 3717 4039
rect 3720 4037 3722 4040
rect 3736 4037 3738 4039
rect 3752 4037 3754 4039
rect 3757 4037 3759 4040
rect 3778 4037 3780 4040
rect 3794 4037 3796 4040
rect 3810 4037 3812 4039
rect 3815 4037 3817 4040
rect 3831 4037 3833 4039
rect 3847 4037 3849 4039
rect 3852 4037 3854 4040
rect 3868 4037 3870 4039
rect 3884 4037 3886 4039
rect 3889 4037 3891 4040
rect 3910 4037 3912 4040
rect 3926 4037 3928 4040
rect 3942 4037 3944 4039
rect 3947 4037 3949 4040
rect 3963 4037 3965 4039
rect 3979 4037 3981 4039
rect 3984 4037 3986 4040
rect 4000 4037 4002 4039
rect 4016 4037 4018 4039
rect 4021 4037 4023 4040
rect 4042 4037 4044 4040
rect 4058 4037 4060 4040
rect 4074 4037 4076 4039
rect 4079 4037 4081 4040
rect 4095 4037 4097 4039
rect 4111 4037 4113 4039
rect 4116 4037 4118 4040
rect 4132 4037 4134 4039
rect 4148 4037 4150 4039
rect 4153 4037 4155 4040
rect 4174 4037 4176 4040
rect 4190 4037 4192 4040
rect 4206 4037 4208 4039
rect 4211 4037 4213 4040
rect 4227 4037 4229 4039
rect 2770 4024 2772 4029
rect 2775 4027 2777 4029
rect 2770 4010 2772 4020
rect 2775 4010 2777 4017
rect 2791 4010 2793 4029
rect 2807 4020 2809 4029
rect 2812 4027 2814 4029
rect 2833 4027 2835 4029
rect 2849 4026 2851 4029
rect 2807 4010 2809 4013
rect 2812 4010 2814 4012
rect 2833 4010 2835 4012
rect 2849 4010 2851 4022
rect 2865 4020 2867 4029
rect 2870 4027 2872 4029
rect 2886 4021 2888 4029
rect 2902 4024 2904 4029
rect 2907 4027 2909 4029
rect 2865 4010 2867 4013
rect 2870 4010 2872 4012
rect 2886 4010 2888 4017
rect 2902 4010 2904 4020
rect 2907 4010 2909 4017
rect 2923 4010 2925 4029
rect 2939 4020 2941 4029
rect 2944 4027 2946 4029
rect 2965 4027 2967 4029
rect 2981 4026 2983 4029
rect 2939 4010 2941 4013
rect 2944 4010 2946 4012
rect 2965 4010 2967 4012
rect 2981 4010 2983 4022
rect 2997 4020 2999 4029
rect 3002 4027 3004 4029
rect 3018 4021 3020 4029
rect 3034 4024 3036 4029
rect 3039 4027 3041 4029
rect 2997 4010 2999 4013
rect 3002 4010 3004 4012
rect 3018 4010 3020 4017
rect 3034 4010 3036 4020
rect 3039 4010 3041 4017
rect 3055 4010 3057 4029
rect 3071 4020 3073 4029
rect 3076 4027 3078 4029
rect 3097 4027 3099 4029
rect 3113 4026 3115 4029
rect 3071 4010 3073 4013
rect 3076 4010 3078 4012
rect 3097 4010 3099 4012
rect 3113 4010 3115 4022
rect 3129 4020 3131 4029
rect 3134 4027 3136 4029
rect 3150 4021 3152 4029
rect 3166 4024 3168 4029
rect 3171 4027 3173 4029
rect 3129 4010 3131 4013
rect 3134 4010 3136 4012
rect 3150 4010 3152 4017
rect 3166 4010 3168 4020
rect 3171 4010 3173 4017
rect 3187 4010 3189 4029
rect 3203 4020 3205 4029
rect 3208 4027 3210 4029
rect 3229 4027 3231 4029
rect 3245 4026 3247 4029
rect 3203 4010 3205 4013
rect 3208 4010 3210 4012
rect 3229 4010 3231 4012
rect 3245 4010 3247 4022
rect 3261 4020 3263 4029
rect 3266 4027 3268 4029
rect 3282 4021 3284 4029
rect 3715 4024 3717 4029
rect 3720 4027 3722 4029
rect 3261 4010 3263 4013
rect 3266 4010 3268 4012
rect 3282 4010 3284 4017
rect 2418 4004 2420 4006
rect 2423 4004 2425 4007
rect 2439 4004 2441 4006
rect 2455 4004 2457 4006
rect 2460 4004 2462 4007
rect 2481 4004 2483 4007
rect 2497 4004 2499 4007
rect 2513 4004 2515 4006
rect 2518 4004 2520 4007
rect 3715 4010 3717 4020
rect 3720 4010 3722 4017
rect 3736 4010 3738 4029
rect 3752 4020 3754 4029
rect 3757 4027 3759 4029
rect 3778 4027 3780 4029
rect 3794 4026 3796 4029
rect 3752 4010 3754 4013
rect 3757 4010 3759 4012
rect 3778 4010 3780 4012
rect 3794 4010 3796 4022
rect 3810 4020 3812 4029
rect 3815 4027 3817 4029
rect 3831 4021 3833 4029
rect 3847 4024 3849 4029
rect 3852 4027 3854 4029
rect 3810 4010 3812 4013
rect 3815 4010 3817 4012
rect 3831 4010 3833 4017
rect 3847 4010 3849 4020
rect 3852 4010 3854 4017
rect 3868 4010 3870 4029
rect 3884 4020 3886 4029
rect 3889 4027 3891 4029
rect 3910 4027 3912 4029
rect 3926 4026 3928 4029
rect 3884 4010 3886 4013
rect 3889 4010 3891 4012
rect 3910 4010 3912 4012
rect 3926 4010 3928 4022
rect 3942 4020 3944 4029
rect 3947 4027 3949 4029
rect 3963 4021 3965 4029
rect 3979 4024 3981 4029
rect 3984 4027 3986 4029
rect 3942 4010 3944 4013
rect 3947 4010 3949 4012
rect 3963 4010 3965 4017
rect 3979 4010 3981 4020
rect 3984 4010 3986 4017
rect 4000 4010 4002 4029
rect 4016 4020 4018 4029
rect 4021 4027 4023 4029
rect 4042 4027 4044 4029
rect 4058 4026 4060 4029
rect 4016 4010 4018 4013
rect 4021 4010 4023 4012
rect 4042 4010 4044 4012
rect 4058 4010 4060 4022
rect 4074 4020 4076 4029
rect 4079 4027 4081 4029
rect 4095 4021 4097 4029
rect 4111 4024 4113 4029
rect 4116 4027 4118 4029
rect 4074 4010 4076 4013
rect 4079 4010 4081 4012
rect 4095 4010 4097 4017
rect 4111 4010 4113 4020
rect 4116 4010 4118 4017
rect 4132 4010 4134 4029
rect 4148 4020 4150 4029
rect 4153 4027 4155 4029
rect 4174 4027 4176 4029
rect 4190 4026 4192 4029
rect 4148 4010 4150 4013
rect 4153 4010 4155 4012
rect 4174 4010 4176 4012
rect 4190 4010 4192 4022
rect 4206 4020 4208 4029
rect 4211 4027 4213 4029
rect 4227 4021 4229 4029
rect 4206 4010 4208 4013
rect 4211 4010 4213 4012
rect 4227 4010 4229 4017
rect 2534 4004 2536 4006
rect 2770 4004 2772 4006
rect 2775 4003 2777 4006
rect 2791 4004 2793 4006
rect 2807 4004 2809 4006
rect 2812 4001 2814 4006
rect 2833 4001 2835 4006
rect 2849 4004 2851 4006
rect 2865 4004 2867 4006
rect 2870 4001 2872 4006
rect 2886 4004 2888 4006
rect 2902 4004 2904 4006
rect 2907 4003 2909 4006
rect 2923 4004 2925 4006
rect 2939 4004 2941 4006
rect 2944 4001 2946 4006
rect 2965 4001 2967 4006
rect 2981 4004 2983 4006
rect 2997 4004 2999 4006
rect 3002 4001 3004 4006
rect 3018 4004 3020 4006
rect 3034 4004 3036 4006
rect 3039 4003 3041 4006
rect 3055 4004 3057 4006
rect 3071 4004 3073 4006
rect 3076 4001 3078 4006
rect 3097 4001 3099 4006
rect 3113 4004 3115 4006
rect 3129 4004 3131 4006
rect 3134 4001 3136 4006
rect 3150 4004 3152 4006
rect 3166 4004 3168 4006
rect 3171 4003 3173 4006
rect 3187 4004 3189 4006
rect 3203 4004 3205 4006
rect 3208 4001 3210 4006
rect 3229 4001 3231 4006
rect 3245 4004 3247 4006
rect 3261 4004 3263 4006
rect 3266 4001 3268 4006
rect 3282 4004 3284 4006
rect 3363 4004 3365 4006
rect 3368 4004 3370 4007
rect 3384 4004 3386 4006
rect 3400 4004 3402 4006
rect 3405 4004 3407 4007
rect 3426 4004 3428 4007
rect 3442 4004 3444 4007
rect 3458 4004 3460 4006
rect 3463 4004 3465 4007
rect 3479 4004 3481 4006
rect 3715 4004 3717 4006
rect 3720 4003 3722 4006
rect 3736 4004 3738 4006
rect 3752 4004 3754 4006
rect 3757 4001 3759 4006
rect 3778 4001 3780 4006
rect 3794 4004 3796 4006
rect 3810 4004 3812 4006
rect 3815 4001 3817 4006
rect 3831 4004 3833 4006
rect 3847 4004 3849 4006
rect 3852 4003 3854 4006
rect 3868 4004 3870 4006
rect 3884 4004 3886 4006
rect 3889 4001 3891 4006
rect 3910 4001 3912 4006
rect 3926 4004 3928 4006
rect 3942 4004 3944 4006
rect 3947 4001 3949 4006
rect 3963 4004 3965 4006
rect 3979 4004 3981 4006
rect 3984 4003 3986 4006
rect 4000 4004 4002 4006
rect 4016 4004 4018 4006
rect 4021 4001 4023 4006
rect 4042 4001 4044 4006
rect 4058 4004 4060 4006
rect 4074 4004 4076 4006
rect 4079 4001 4081 4006
rect 4095 4004 4097 4006
rect 4111 4004 4113 4006
rect 4116 4003 4118 4006
rect 4132 4004 4134 4006
rect 4148 4004 4150 4006
rect 4153 4001 4155 4006
rect 4174 4001 4176 4006
rect 4190 4004 4192 4006
rect 4206 4004 4208 4006
rect 4211 4001 4213 4006
rect 4227 4004 4229 4006
rect 2418 3991 2420 3996
rect 2423 3994 2425 3996
rect 2418 3977 2420 3987
rect 2423 3977 2425 3984
rect 2439 3977 2441 3996
rect 2455 3987 2457 3996
rect 2460 3994 2462 3996
rect 2481 3994 2483 3996
rect 2497 3993 2499 3996
rect 2455 3977 2457 3980
rect 2460 3977 2462 3979
rect 2481 3977 2483 3979
rect 2497 3977 2499 3989
rect 2513 3987 2515 3996
rect 2518 3994 2520 3996
rect 2513 3977 2515 3980
rect 2518 3977 2520 3979
rect 2534 3977 2536 3996
rect 3363 3991 3365 3996
rect 3368 3994 3370 3996
rect 3363 3977 3365 3987
rect 3368 3977 3370 3984
rect 3384 3977 3386 3996
rect 3400 3987 3402 3996
rect 3405 3994 3407 3996
rect 3426 3994 3428 3996
rect 3442 3993 3444 3996
rect 3400 3977 3402 3980
rect 3405 3977 3407 3979
rect 3426 3977 3428 3979
rect 3442 3977 3444 3989
rect 3458 3987 3460 3996
rect 3463 3994 3465 3996
rect 3458 3977 3460 3980
rect 3463 3977 3465 3979
rect 3479 3977 3481 3996
rect 2418 3971 2420 3973
rect 2423 3970 2425 3973
rect 2439 3971 2441 3973
rect 2455 3971 2457 3973
rect 2460 3968 2462 3973
rect 2481 3968 2483 3973
rect 2497 3971 2499 3973
rect 2513 3971 2515 3973
rect 2518 3968 2520 3973
rect 2534 3971 2536 3973
rect 3363 3971 3365 3973
rect 3368 3970 3370 3973
rect 3384 3971 3386 3973
rect 3400 3971 3402 3973
rect 2949 3966 2951 3968
rect 2791 3960 2793 3963
rect 2835 3960 2837 3963
rect 2861 3960 2863 3963
rect 2907 3960 2909 3963
rect 2861 3956 2862 3960
rect 2975 3960 2977 3964
rect 3003 3966 3005 3968
rect 3030 3966 3032 3968
rect 2980 3960 2982 3963
rect 2775 3953 2777 3955
rect 2791 3953 2793 3956
rect 2807 3953 2809 3955
rect 2830 3953 2832 3955
rect 2835 3953 2837 3956
rect 2861 3953 2863 3956
rect 2882 3953 2884 3956
rect 2902 3953 2904 3955
rect 2907 3953 2909 3956
rect 2925 3953 2927 3955
rect 2542 3940 2544 3943
rect 2542 3934 2544 3936
rect 2425 3931 2427 3934
rect 2775 3931 2777 3945
rect 2791 3943 2793 3945
rect 2791 3931 2793 3933
rect 2807 3931 2809 3945
rect 2830 3940 2832 3945
rect 2835 3943 2837 3945
rect 2861 3943 2863 3945
rect 2826 3936 2832 3940
rect 2830 3931 2832 3936
rect 2835 3931 2837 3933
rect 2861 3931 2863 3933
rect 2882 3931 2884 3945
rect 2902 3940 2904 3945
rect 2907 3943 2909 3945
rect 2898 3936 2904 3940
rect 2902 3931 2904 3936
rect 2907 3931 2909 3933
rect 2925 3931 2927 3945
rect 2949 3944 2951 3958
rect 3056 3960 3058 3964
rect 3084 3966 3086 3968
rect 3405 3968 3407 3973
rect 3426 3968 3428 3973
rect 3442 3971 3444 3973
rect 3458 3971 3460 3973
rect 3463 3968 3465 3973
rect 3479 3971 3481 3973
rect 3061 3960 3063 3963
rect 2975 3949 2977 3952
rect 2980 3950 2982 3952
rect 2976 3945 2977 3949
rect 2975 3940 2977 3945
rect 2980 3940 2982 3942
rect 2949 3938 2951 3940
rect 3003 3936 3005 3958
rect 3030 3944 3032 3958
rect 3894 3966 3896 3968
rect 3056 3949 3058 3952
rect 3061 3950 3063 3952
rect 3057 3945 3058 3949
rect 3056 3940 3058 3945
rect 3061 3940 3063 3942
rect 3030 3938 3032 3940
rect 3084 3936 3086 3958
rect 3736 3960 3738 3963
rect 3780 3960 3782 3963
rect 3806 3960 3808 3963
rect 3852 3960 3854 3963
rect 3806 3956 3807 3960
rect 3920 3960 3922 3964
rect 3948 3966 3950 3968
rect 3975 3966 3977 3968
rect 3925 3960 3927 3963
rect 3720 3953 3722 3955
rect 3736 3953 3738 3956
rect 3752 3953 3754 3955
rect 3775 3953 3777 3955
rect 3780 3953 3782 3956
rect 3806 3953 3808 3956
rect 3827 3953 3829 3956
rect 3847 3953 3849 3955
rect 3852 3953 3854 3956
rect 3870 3953 3872 3955
rect 3487 3940 3489 3943
rect 2975 3934 2977 3936
rect 2980 3931 2982 3936
rect 3056 3934 3058 3936
rect 3003 3930 3005 3932
rect 3061 3931 3063 3936
rect 3487 3934 3489 3936
rect 3084 3930 3086 3932
rect 3370 3931 3372 3934
rect 3720 3931 3722 3945
rect 3736 3943 3738 3945
rect 3736 3931 3738 3933
rect 3752 3931 3754 3945
rect 3775 3940 3777 3945
rect 3780 3943 3782 3945
rect 3806 3943 3808 3945
rect 3771 3936 3777 3940
rect 3775 3931 3777 3936
rect 3780 3931 3782 3933
rect 3806 3931 3808 3933
rect 3827 3931 3829 3945
rect 3847 3940 3849 3945
rect 3852 3943 3854 3945
rect 3843 3936 3849 3940
rect 3847 3931 3849 3936
rect 3852 3931 3854 3933
rect 3870 3931 3872 3945
rect 3894 3944 3896 3958
rect 4001 3960 4003 3964
rect 4029 3966 4031 3968
rect 4006 3960 4008 3963
rect 3920 3949 3922 3952
rect 3925 3950 3927 3952
rect 3921 3945 3922 3949
rect 3920 3940 3922 3945
rect 3925 3940 3927 3942
rect 3894 3938 3896 3940
rect 3948 3936 3950 3958
rect 3975 3944 3977 3958
rect 4001 3949 4003 3952
rect 4006 3950 4008 3952
rect 4002 3945 4003 3949
rect 4001 3940 4003 3945
rect 4006 3940 4008 3942
rect 3975 3938 3977 3940
rect 4029 3936 4031 3958
rect 3920 3934 3922 3936
rect 3925 3931 3927 3936
rect 4001 3934 4003 3936
rect 3948 3930 3950 3932
rect 4006 3931 4008 3936
rect 4029 3930 4031 3932
rect 2425 3925 2427 3927
rect 2775 3925 2777 3927
rect 2791 3923 2793 3927
rect 2807 3925 2809 3927
rect 2830 3925 2832 3927
rect 2792 3919 2793 3923
rect 2835 3922 2837 3927
rect 2861 3923 2863 3927
rect 2882 3925 2884 3927
rect 2902 3925 2904 3927
rect 2791 3916 2793 3919
rect 2836 3918 2837 3922
rect 2862 3919 2863 3923
rect 2907 3922 2909 3927
rect 2925 3925 2927 3927
rect 3370 3925 3372 3927
rect 3720 3925 3722 3927
rect 3736 3923 3738 3927
rect 3752 3925 3754 3927
rect 3775 3925 3777 3927
rect 2835 3916 2837 3918
rect 2861 3915 2863 3919
rect 2908 3918 2909 3922
rect 3737 3919 3738 3923
rect 3780 3922 3782 3927
rect 3806 3923 3808 3927
rect 3827 3925 3829 3927
rect 3847 3925 3849 3927
rect 2907 3916 2909 3918
rect 3736 3916 3738 3919
rect 3781 3918 3782 3922
rect 3807 3919 3808 3923
rect 3852 3922 3854 3927
rect 3870 3925 3872 3927
rect 3780 3916 3782 3918
rect 3806 3915 3808 3919
rect 3853 3918 3854 3922
rect 3852 3916 3854 3918
rect 2409 3902 2411 3904
rect 2425 3902 2427 3905
rect 2430 3902 2432 3904
rect 2446 3902 2448 3905
rect 2462 3902 2464 3905
rect 2483 3902 2485 3905
rect 2488 3902 2490 3904
rect 2504 3902 2506 3904
rect 2520 3902 2522 3905
rect 2525 3902 2527 3904
rect 3354 3902 3356 3904
rect 3370 3902 3372 3905
rect 3375 3902 3377 3904
rect 3391 3902 3393 3905
rect 3407 3902 3409 3905
rect 3428 3902 3430 3905
rect 3433 3902 3435 3904
rect 3449 3902 3451 3904
rect 3465 3902 3467 3905
rect 3470 3902 3472 3904
rect 2409 3875 2411 3894
rect 2425 3892 2427 3894
rect 2430 3885 2432 3894
rect 2446 3891 2448 3894
rect 2462 3892 2464 3894
rect 2483 3892 2485 3894
rect 2425 3875 2427 3877
rect 2430 3875 2432 3878
rect 2446 3875 2448 3887
rect 2488 3885 2490 3894
rect 2462 3875 2464 3877
rect 2483 3875 2485 3877
rect 2488 3875 2490 3878
rect 2504 3875 2506 3894
rect 2520 3892 2522 3894
rect 2525 3889 2527 3894
rect 2791 3893 2793 3896
rect 2835 3894 2837 3896
rect 2792 3889 2793 3893
rect 2836 3890 2837 3894
rect 2861 3893 2863 3897
rect 2907 3894 2909 3896
rect 2775 3885 2777 3887
rect 2791 3885 2793 3889
rect 2807 3885 2809 3887
rect 2830 3885 2832 3887
rect 2835 3885 2837 3890
rect 2862 3889 2863 3893
rect 2908 3890 2909 3894
rect 2861 3885 2863 3889
rect 2882 3885 2884 3887
rect 2902 3885 2904 3887
rect 2907 3885 2909 3890
rect 2925 3885 2927 3887
rect 2520 3875 2522 3882
rect 2525 3875 2527 3885
rect 2975 3884 2977 3887
rect 2980 3884 2982 3887
rect 3056 3884 3058 3887
rect 3061 3884 3063 3887
rect 2409 3869 2411 3871
rect 2425 3866 2427 3871
rect 2430 3869 2432 3871
rect 2446 3869 2448 3871
rect 2462 3866 2464 3871
rect 2483 3866 2485 3871
rect 2488 3869 2490 3871
rect 2504 3869 2506 3871
rect 2520 3868 2522 3871
rect 2525 3869 2527 3871
rect 2775 3867 2777 3881
rect 2791 3879 2793 3881
rect 2791 3867 2793 3869
rect 2807 3867 2809 3881
rect 2830 3876 2832 3881
rect 2835 3879 2837 3881
rect 2861 3879 2863 3881
rect 2826 3872 2832 3876
rect 2830 3867 2832 3872
rect 2835 3867 2837 3869
rect 2861 3867 2863 3869
rect 2882 3867 2884 3881
rect 2902 3876 2904 3881
rect 2907 3879 2909 3881
rect 2898 3872 2904 3876
rect 2902 3867 2904 3872
rect 2907 3867 2909 3869
rect 2925 3867 2927 3881
rect 2975 3868 2977 3880
rect 2980 3878 2982 3880
rect 2980 3868 2982 3870
rect 3056 3868 3058 3880
rect 3061 3878 3063 3880
rect 3354 3875 3356 3894
rect 3370 3892 3372 3894
rect 3375 3885 3377 3894
rect 3391 3891 3393 3894
rect 3407 3892 3409 3894
rect 3428 3892 3430 3894
rect 3370 3875 3372 3877
rect 3375 3875 3377 3878
rect 3391 3875 3393 3887
rect 3433 3885 3435 3894
rect 3407 3875 3409 3877
rect 3428 3875 3430 3877
rect 3433 3875 3435 3878
rect 3449 3875 3451 3894
rect 3465 3892 3467 3894
rect 3470 3889 3472 3894
rect 3736 3893 3738 3896
rect 3780 3894 3782 3896
rect 3737 3889 3738 3893
rect 3781 3890 3782 3894
rect 3806 3893 3808 3897
rect 3852 3894 3854 3896
rect 3720 3885 3722 3887
rect 3736 3885 3738 3889
rect 3752 3885 3754 3887
rect 3775 3885 3777 3887
rect 3780 3885 3782 3890
rect 3807 3889 3808 3893
rect 3853 3890 3854 3894
rect 3806 3885 3808 3889
rect 3827 3885 3829 3887
rect 3847 3885 3849 3887
rect 3852 3885 3854 3890
rect 3870 3885 3872 3887
rect 3465 3875 3467 3882
rect 3470 3875 3472 3885
rect 3920 3884 3922 3887
rect 3925 3884 3927 3887
rect 4001 3884 4003 3887
rect 4006 3884 4008 3887
rect 3061 3868 3063 3870
rect 3354 3869 3356 3871
rect 3370 3866 3372 3871
rect 3375 3869 3377 3871
rect 3391 3869 3393 3871
rect 3407 3866 3409 3871
rect 3428 3866 3430 3871
rect 3433 3869 3435 3871
rect 3449 3869 3451 3871
rect 3465 3868 3467 3871
rect 3470 3869 3472 3871
rect 3720 3867 3722 3881
rect 3736 3879 3738 3881
rect 3736 3867 3738 3869
rect 3752 3867 3754 3881
rect 3775 3876 3777 3881
rect 3780 3879 3782 3881
rect 3806 3879 3808 3881
rect 3771 3872 3777 3876
rect 3775 3867 3777 3872
rect 3780 3867 3782 3869
rect 3806 3867 3808 3869
rect 3827 3867 3829 3881
rect 3847 3876 3849 3881
rect 3852 3879 3854 3881
rect 3843 3872 3849 3876
rect 3847 3867 3849 3872
rect 3852 3867 3854 3869
rect 3870 3867 3872 3881
rect 3920 3868 3922 3880
rect 3925 3878 3927 3880
rect 3925 3868 3927 3870
rect 4001 3868 4003 3880
rect 4006 3878 4008 3880
rect 4006 3868 4008 3870
rect 2775 3857 2777 3859
rect 2791 3856 2793 3859
rect 2807 3857 2809 3859
rect 2830 3857 2832 3859
rect 2835 3856 2837 3859
rect 2861 3856 2863 3859
rect 2882 3856 2884 3859
rect 2902 3857 2904 3859
rect 2907 3856 2909 3859
rect 2925 3857 2927 3859
rect 2975 3858 2977 3860
rect 2861 3852 2862 3856
rect 2980 3855 2982 3860
rect 3056 3858 3058 3860
rect 3061 3855 3063 3860
rect 3720 3857 3722 3859
rect 3736 3856 3738 3859
rect 3752 3857 3754 3859
rect 3775 3857 3777 3859
rect 3780 3856 3782 3859
rect 3806 3856 3808 3859
rect 3827 3856 3829 3859
rect 3847 3857 3849 3859
rect 3852 3856 3854 3859
rect 3870 3857 3872 3859
rect 3920 3858 3922 3860
rect 2791 3849 2793 3852
rect 2835 3849 2837 3852
rect 2861 3849 2863 3852
rect 2907 3849 2909 3852
rect 3806 3852 3807 3856
rect 3925 3855 3927 3860
rect 4001 3858 4003 3860
rect 4006 3855 4008 3860
rect 3736 3849 3738 3852
rect 3780 3849 3782 3852
rect 3806 3849 3808 3852
rect 3852 3849 3854 3852
rect 2791 3828 2793 3831
rect 2835 3828 2837 3831
rect 2861 3828 2863 3831
rect 2907 3828 2909 3831
rect 2975 3828 2977 3832
rect 3003 3834 3005 3836
rect 3054 3834 3056 3836
rect 2980 3828 2982 3831
rect 2861 3824 2862 3828
rect 2775 3821 2777 3823
rect 2791 3821 2793 3824
rect 2807 3821 2809 3823
rect 2830 3821 2832 3823
rect 2835 3821 2837 3824
rect 2861 3821 2863 3824
rect 2882 3821 2884 3824
rect 2902 3821 2904 3823
rect 2907 3821 2909 3824
rect 2925 3821 2927 3823
rect 3080 3828 3082 3832
rect 3108 3834 3110 3836
rect 3085 3828 3087 3831
rect 2975 3817 2977 3820
rect 2980 3818 2982 3820
rect 2976 3813 2977 3817
rect 2775 3799 2777 3813
rect 2791 3811 2793 3813
rect 2791 3799 2793 3801
rect 2807 3799 2809 3813
rect 2830 3808 2832 3813
rect 2835 3811 2837 3813
rect 2861 3811 2863 3813
rect 2826 3804 2832 3808
rect 2830 3799 2832 3804
rect 2835 3799 2837 3801
rect 2861 3799 2863 3801
rect 2882 3799 2884 3813
rect 2902 3808 2904 3813
rect 2907 3811 2909 3813
rect 2898 3804 2904 3808
rect 2902 3799 2904 3804
rect 2907 3799 2909 3801
rect 2925 3799 2927 3813
rect 2975 3808 2977 3813
rect 2980 3808 2982 3810
rect 3003 3804 3005 3826
rect 3054 3812 3056 3826
rect 3736 3828 3738 3831
rect 3780 3828 3782 3831
rect 3806 3828 3808 3831
rect 3852 3828 3854 3831
rect 3920 3828 3922 3832
rect 3948 3834 3950 3836
rect 3999 3834 4001 3836
rect 3925 3828 3927 3831
rect 3080 3817 3082 3820
rect 3085 3818 3087 3820
rect 3081 3813 3082 3817
rect 3080 3808 3082 3813
rect 3085 3808 3087 3810
rect 3054 3806 3056 3808
rect 3108 3804 3110 3826
rect 3806 3824 3807 3828
rect 3720 3821 3722 3823
rect 3736 3821 3738 3824
rect 3752 3821 3754 3823
rect 3775 3821 3777 3823
rect 3780 3821 3782 3824
rect 3806 3821 3808 3824
rect 3827 3821 3829 3824
rect 3847 3821 3849 3823
rect 3852 3821 3854 3824
rect 3870 3821 3872 3823
rect 4025 3828 4027 3832
rect 4053 3834 4055 3836
rect 4030 3828 4032 3831
rect 3920 3817 3922 3820
rect 3925 3818 3927 3820
rect 3921 3813 3922 3817
rect 3285 3805 3287 3807
rect 2975 3802 2977 3804
rect 2980 3799 2982 3804
rect 3080 3802 3082 3804
rect 3003 3798 3005 3800
rect 3085 3799 3087 3804
rect 3108 3798 3110 3800
rect 3311 3799 3313 3803
rect 3339 3805 3341 3807
rect 3316 3799 3318 3802
rect 2775 3793 2777 3795
rect 2791 3791 2793 3795
rect 2807 3793 2809 3795
rect 2830 3793 2832 3795
rect 2792 3787 2793 3791
rect 2835 3790 2837 3795
rect 2861 3791 2863 3795
rect 2882 3793 2884 3795
rect 2902 3793 2904 3795
rect 2791 3784 2793 3787
rect 2836 3786 2837 3790
rect 2862 3787 2863 3791
rect 2907 3790 2909 3795
rect 2925 3793 2927 3795
rect 2835 3784 2837 3786
rect 2861 3783 2863 3787
rect 2908 3786 2909 3790
rect 2907 3784 2909 3786
rect 3285 3783 3287 3797
rect 3471 3802 3473 3805
rect 3524 3802 3526 3805
rect 3311 3788 3313 3791
rect 3316 3789 3318 3791
rect 3312 3784 3313 3788
rect 3311 3779 3313 3784
rect 3316 3779 3318 3781
rect 3285 3777 3287 3779
rect 3339 3775 3341 3797
rect 3311 3773 3313 3775
rect 3316 3770 3318 3775
rect 3720 3799 3722 3813
rect 3736 3811 3738 3813
rect 3736 3799 3738 3801
rect 3752 3799 3754 3813
rect 3775 3808 3777 3813
rect 3780 3811 3782 3813
rect 3806 3811 3808 3813
rect 3771 3804 3777 3808
rect 3775 3799 3777 3804
rect 3780 3799 3782 3801
rect 3806 3799 3808 3801
rect 3827 3799 3829 3813
rect 3847 3808 3849 3813
rect 3852 3811 3854 3813
rect 3843 3804 3849 3808
rect 3847 3799 3849 3804
rect 3852 3799 3854 3801
rect 3870 3799 3872 3813
rect 3920 3808 3922 3813
rect 3925 3808 3927 3810
rect 3948 3804 3950 3826
rect 3999 3812 4001 3826
rect 4025 3817 4027 3820
rect 4030 3818 4032 3820
rect 4026 3813 4027 3817
rect 4025 3808 4027 3813
rect 4030 3808 4032 3810
rect 3999 3806 4001 3808
rect 4053 3804 4055 3826
rect 3920 3802 3922 3804
rect 3925 3799 3927 3804
rect 4025 3802 4027 3804
rect 3948 3798 3950 3800
rect 4030 3799 4032 3804
rect 4053 3798 4055 3800
rect 3720 3793 3722 3795
rect 3736 3791 3738 3795
rect 3752 3793 3754 3795
rect 3775 3793 3777 3795
rect 3737 3787 3738 3791
rect 3780 3790 3782 3795
rect 3806 3791 3808 3795
rect 3827 3793 3829 3795
rect 3847 3793 3849 3795
rect 3736 3784 3738 3787
rect 3781 3786 3782 3790
rect 3807 3787 3808 3791
rect 3852 3790 3854 3795
rect 3870 3793 3872 3795
rect 3780 3784 3782 3786
rect 3806 3783 3808 3787
rect 3853 3786 3854 3790
rect 3852 3784 3854 3786
rect 3339 3769 3341 3771
rect 2791 3761 2793 3764
rect 2835 3762 2837 3764
rect 2792 3757 2793 3761
rect 2836 3758 2837 3762
rect 2861 3761 2863 3765
rect 3471 3764 3473 3772
rect 3524 3764 3526 3772
rect 2907 3762 2909 3764
rect 2775 3753 2777 3755
rect 2791 3753 2793 3757
rect 2807 3753 2809 3755
rect 2830 3753 2832 3755
rect 2835 3753 2837 3758
rect 2862 3757 2863 3761
rect 2908 3758 2909 3762
rect 3736 3761 3738 3764
rect 3780 3762 3782 3764
rect 2861 3753 2863 3757
rect 2882 3753 2884 3755
rect 2902 3753 2904 3755
rect 2907 3753 2909 3758
rect 2925 3753 2927 3755
rect 2975 3753 2977 3756
rect 2980 3753 2982 3756
rect 3080 3753 3082 3756
rect 3085 3753 3087 3756
rect 3471 3752 3473 3760
rect 3524 3752 3526 3760
rect 3737 3757 3738 3761
rect 3781 3758 3782 3762
rect 3806 3761 3808 3765
rect 3852 3762 3854 3764
rect 3720 3753 3722 3755
rect 3736 3753 3738 3757
rect 3752 3753 3754 3755
rect 3775 3753 3777 3755
rect 3780 3753 3782 3758
rect 3807 3757 3808 3761
rect 3853 3758 3854 3762
rect 3806 3753 3808 3757
rect 3827 3753 3829 3755
rect 3847 3753 3849 3755
rect 3852 3753 3854 3758
rect 3870 3753 3872 3755
rect 3920 3753 3922 3756
rect 3925 3753 3927 3756
rect 4025 3753 4027 3756
rect 4030 3753 4032 3756
rect 2775 3735 2777 3749
rect 2791 3747 2793 3749
rect 2791 3735 2793 3737
rect 2807 3735 2809 3749
rect 2830 3744 2832 3749
rect 2835 3747 2837 3749
rect 2861 3747 2863 3749
rect 2826 3740 2832 3744
rect 2830 3735 2832 3740
rect 2835 3735 2837 3737
rect 2861 3735 2863 3737
rect 2882 3735 2884 3749
rect 2902 3744 2904 3749
rect 2907 3747 2909 3749
rect 2898 3740 2904 3744
rect 2902 3735 2904 3740
rect 2907 3735 2909 3737
rect 2925 3735 2927 3749
rect 2975 3737 2977 3749
rect 2980 3747 2982 3749
rect 2980 3737 2982 3739
rect 3080 3737 3082 3749
rect 3085 3747 3087 3749
rect 3085 3737 3087 3739
rect 3471 3738 3473 3740
rect 3524 3738 3526 3740
rect 3720 3735 3722 3749
rect 3736 3747 3738 3749
rect 3736 3735 3738 3737
rect 3752 3735 3754 3749
rect 3775 3744 3777 3749
rect 3780 3747 3782 3749
rect 3806 3747 3808 3749
rect 3771 3740 3777 3744
rect 3775 3735 3777 3740
rect 3780 3735 3782 3737
rect 3806 3735 3808 3737
rect 3827 3735 3829 3749
rect 3847 3744 3849 3749
rect 3852 3747 3854 3749
rect 3843 3740 3849 3744
rect 3847 3735 3849 3740
rect 3852 3735 3854 3737
rect 3870 3735 3872 3749
rect 3920 3737 3922 3749
rect 3925 3747 3927 3749
rect 3925 3737 3927 3739
rect 4025 3737 4027 3749
rect 4030 3747 4032 3749
rect 4030 3737 4032 3739
rect 2975 3727 2977 3729
rect 2775 3725 2777 3727
rect 2791 3724 2793 3727
rect 2807 3725 2809 3727
rect 2830 3725 2832 3727
rect 2835 3724 2837 3727
rect 2861 3724 2863 3727
rect 2882 3724 2884 3727
rect 2902 3725 2904 3727
rect 2907 3724 2909 3727
rect 2925 3725 2927 3727
rect 2980 3724 2982 3729
rect 3080 3727 3082 3729
rect 3085 3724 3087 3729
rect 3920 3727 3922 3729
rect 2861 3720 2862 3724
rect 3720 3725 3722 3727
rect 3736 3724 3738 3727
rect 3752 3725 3754 3727
rect 3775 3725 3777 3727
rect 3780 3724 3782 3727
rect 3806 3724 3808 3727
rect 3827 3724 3829 3727
rect 3847 3725 3849 3727
rect 3852 3724 3854 3727
rect 3870 3725 3872 3727
rect 3925 3724 3927 3729
rect 4025 3727 4027 3729
rect 4030 3724 4032 3729
rect 2791 3717 2793 3720
rect 2835 3717 2837 3720
rect 2861 3717 2863 3720
rect 2907 3717 2909 3720
rect 3311 3719 3313 3722
rect 3316 3719 3318 3722
rect 3806 3720 3807 3724
rect 3736 3717 3738 3720
rect 3780 3717 3782 3720
rect 3806 3717 3808 3720
rect 3852 3717 3854 3720
rect 2791 3696 2793 3699
rect 2835 3696 2837 3699
rect 2861 3696 2863 3699
rect 2907 3696 2909 3699
rect 2975 3696 2977 3700
rect 3003 3702 3005 3704
rect 3030 3702 3032 3704
rect 2980 3696 2982 3699
rect 2861 3692 2862 3696
rect 2775 3689 2777 3691
rect 2791 3689 2793 3692
rect 2807 3689 2809 3691
rect 2830 3689 2832 3691
rect 2835 3689 2837 3692
rect 2861 3689 2863 3692
rect 2882 3689 2884 3692
rect 2902 3689 2904 3691
rect 2907 3689 2909 3692
rect 2925 3689 2927 3691
rect 3056 3696 3058 3700
rect 3084 3702 3086 3704
rect 3120 3702 3122 3704
rect 3061 3696 3063 3699
rect 2975 3685 2977 3688
rect 2980 3686 2982 3688
rect 2976 3681 2977 3685
rect 2775 3667 2777 3681
rect 2791 3679 2793 3681
rect 2791 3667 2793 3669
rect 2807 3667 2809 3681
rect 2830 3676 2832 3681
rect 2835 3679 2837 3681
rect 2861 3679 2863 3681
rect 2826 3672 2832 3676
rect 2830 3667 2832 3672
rect 2835 3667 2837 3669
rect 2861 3667 2863 3669
rect 2882 3667 2884 3681
rect 2902 3676 2904 3681
rect 2907 3679 2909 3681
rect 2898 3672 2904 3676
rect 2902 3667 2904 3672
rect 2907 3667 2909 3669
rect 2925 3667 2927 3681
rect 2975 3676 2977 3681
rect 2980 3676 2982 3678
rect 3003 3672 3005 3694
rect 3030 3680 3032 3694
rect 3146 3696 3148 3700
rect 3174 3702 3176 3704
rect 3311 3703 3313 3715
rect 3316 3713 3318 3715
rect 3316 3703 3318 3705
rect 3151 3696 3153 3699
rect 3056 3685 3058 3688
rect 3061 3686 3063 3688
rect 3057 3681 3058 3685
rect 3056 3676 3058 3681
rect 3061 3676 3063 3678
rect 3030 3674 3032 3676
rect 3084 3672 3086 3694
rect 3120 3680 3122 3694
rect 3736 3696 3738 3699
rect 3780 3696 3782 3699
rect 3806 3696 3808 3699
rect 3852 3696 3854 3699
rect 3920 3696 3922 3700
rect 3948 3702 3950 3704
rect 3975 3702 3977 3704
rect 3925 3696 3927 3699
rect 3146 3685 3148 3688
rect 3151 3686 3153 3688
rect 3147 3681 3148 3685
rect 3146 3676 3148 3681
rect 3151 3676 3153 3678
rect 3120 3674 3122 3676
rect 3174 3672 3176 3694
rect 3311 3693 3313 3695
rect 3316 3690 3318 3695
rect 3806 3692 3807 3696
rect 3720 3689 3722 3691
rect 3736 3689 3738 3692
rect 3752 3689 3754 3691
rect 3775 3689 3777 3691
rect 3780 3689 3782 3692
rect 3806 3689 3808 3692
rect 3827 3689 3829 3692
rect 3847 3689 3849 3691
rect 3852 3689 3854 3692
rect 3870 3689 3872 3691
rect 4001 3696 4003 3700
rect 4029 3702 4031 3704
rect 4065 3702 4067 3704
rect 4006 3696 4008 3699
rect 3920 3685 3922 3688
rect 3925 3686 3927 3688
rect 3921 3681 3922 3685
rect 3263 3675 3265 3677
rect 3285 3675 3287 3677
rect 2975 3670 2977 3672
rect 2980 3667 2982 3672
rect 3056 3670 3058 3672
rect 3003 3666 3005 3668
rect 3061 3667 3063 3672
rect 3146 3670 3148 3672
rect 3084 3666 3086 3668
rect 3151 3667 3153 3672
rect 3174 3666 3176 3668
rect 3311 3669 3313 3673
rect 3339 3675 3341 3677
rect 3316 3669 3318 3672
rect 2775 3661 2777 3663
rect 2791 3659 2793 3663
rect 2807 3661 2809 3663
rect 2830 3661 2832 3663
rect 2792 3655 2793 3659
rect 2835 3658 2837 3663
rect 2861 3659 2863 3663
rect 2882 3661 2884 3663
rect 2902 3661 2904 3663
rect 2791 3652 2793 3655
rect 2836 3654 2837 3658
rect 2862 3655 2863 3659
rect 2907 3658 2909 3663
rect 2925 3661 2927 3663
rect 2835 3652 2837 3654
rect 2861 3651 2863 3655
rect 2908 3654 2909 3658
rect 2907 3652 2909 3654
rect 3263 3653 3265 3667
rect 3285 3653 3287 3667
rect 3377 3672 3379 3675
rect 3430 3672 3432 3675
rect 3311 3658 3313 3661
rect 3316 3659 3318 3661
rect 3312 3654 3313 3658
rect 3311 3649 3313 3654
rect 3316 3649 3318 3651
rect 3263 3647 3265 3649
rect 3285 3647 3287 3649
rect 3339 3645 3341 3667
rect 3311 3643 3313 3645
rect 3316 3640 3318 3645
rect 3720 3667 3722 3681
rect 3736 3679 3738 3681
rect 3736 3667 3738 3669
rect 3752 3667 3754 3681
rect 3775 3676 3777 3681
rect 3780 3679 3782 3681
rect 3806 3679 3808 3681
rect 3771 3672 3777 3676
rect 3775 3667 3777 3672
rect 3780 3667 3782 3669
rect 3806 3667 3808 3669
rect 3827 3667 3829 3681
rect 3847 3676 3849 3681
rect 3852 3679 3854 3681
rect 3843 3672 3849 3676
rect 3847 3667 3849 3672
rect 3852 3667 3854 3669
rect 3870 3667 3872 3681
rect 3920 3676 3922 3681
rect 3925 3676 3927 3678
rect 3948 3672 3950 3694
rect 3975 3680 3977 3694
rect 4091 3696 4093 3700
rect 4119 3702 4121 3704
rect 4096 3696 4098 3699
rect 4001 3685 4003 3688
rect 4006 3686 4008 3688
rect 4002 3681 4003 3685
rect 4001 3676 4003 3681
rect 4006 3676 4008 3678
rect 3975 3674 3977 3676
rect 4029 3672 4031 3694
rect 4065 3680 4067 3694
rect 4091 3685 4093 3688
rect 4096 3686 4098 3688
rect 4092 3681 4093 3685
rect 4091 3676 4093 3681
rect 4096 3676 4098 3678
rect 4065 3674 4067 3676
rect 4119 3672 4121 3694
rect 3920 3670 3922 3672
rect 3925 3667 3927 3672
rect 4001 3670 4003 3672
rect 3948 3666 3950 3668
rect 4006 3667 4008 3672
rect 4091 3670 4093 3672
rect 4029 3666 4031 3668
rect 4096 3667 4098 3672
rect 4119 3666 4121 3668
rect 3720 3661 3722 3663
rect 3736 3659 3738 3663
rect 3752 3661 3754 3663
rect 3775 3661 3777 3663
rect 3737 3655 3738 3659
rect 3780 3658 3782 3663
rect 3806 3659 3808 3663
rect 3827 3661 3829 3663
rect 3847 3661 3849 3663
rect 3736 3652 3738 3655
rect 3781 3654 3782 3658
rect 3807 3655 3808 3659
rect 3852 3658 3854 3663
rect 3870 3661 3872 3663
rect 3780 3652 3782 3654
rect 3806 3651 3808 3655
rect 3853 3654 3854 3658
rect 3852 3652 3854 3654
rect 3339 3639 3341 3641
rect 3377 3634 3379 3642
rect 3430 3634 3432 3642
rect 2791 3629 2793 3632
rect 2835 3630 2837 3632
rect 2792 3625 2793 3629
rect 2836 3626 2837 3630
rect 2861 3629 2863 3633
rect 2907 3630 2909 3632
rect 2775 3621 2777 3623
rect 2791 3621 2793 3625
rect 2807 3621 2809 3623
rect 2830 3621 2832 3623
rect 2835 3621 2837 3626
rect 2862 3625 2863 3629
rect 2908 3626 2909 3630
rect 2861 3621 2863 3625
rect 2882 3621 2884 3623
rect 2902 3621 2904 3623
rect 2907 3621 2909 3626
rect 2925 3621 2927 3623
rect 3377 3622 3379 3630
rect 3430 3622 3432 3630
rect 3736 3629 3738 3632
rect 3780 3630 3782 3632
rect 3737 3625 3738 3629
rect 3781 3626 3782 3630
rect 3806 3629 3808 3633
rect 3852 3630 3854 3632
rect 2975 3618 2977 3621
rect 2980 3618 2982 3621
rect 3056 3618 3058 3621
rect 3061 3618 3063 3621
rect 3146 3618 3148 3621
rect 3151 3618 3153 3621
rect 2775 3603 2777 3617
rect 2791 3615 2793 3617
rect 2791 3603 2793 3605
rect 2807 3603 2809 3617
rect 2830 3612 2832 3617
rect 2835 3615 2837 3617
rect 2861 3615 2863 3617
rect 2826 3608 2832 3612
rect 2830 3603 2832 3608
rect 2835 3603 2837 3605
rect 2861 3603 2863 3605
rect 2882 3603 2884 3617
rect 2902 3612 2904 3617
rect 2907 3615 2909 3617
rect 2898 3608 2904 3612
rect 2902 3603 2904 3608
rect 2907 3603 2909 3605
rect 2925 3603 2927 3617
rect 2975 3602 2977 3614
rect 2980 3612 2982 3614
rect 2980 3602 2982 3604
rect 3056 3602 3058 3614
rect 3061 3612 3063 3614
rect 3061 3602 3063 3604
rect 3146 3602 3148 3614
rect 3151 3612 3153 3614
rect 3720 3621 3722 3623
rect 3736 3621 3738 3625
rect 3752 3621 3754 3623
rect 3775 3621 3777 3623
rect 3780 3621 3782 3626
rect 3807 3625 3808 3629
rect 3853 3626 3854 3630
rect 3806 3621 3808 3625
rect 3827 3621 3829 3623
rect 3847 3621 3849 3623
rect 3852 3621 3854 3626
rect 3870 3621 3872 3623
rect 3920 3618 3922 3621
rect 3925 3618 3927 3621
rect 4001 3618 4003 3621
rect 4006 3618 4008 3621
rect 4091 3618 4093 3621
rect 4096 3618 4098 3621
rect 3377 3608 3379 3610
rect 3430 3608 3432 3610
rect 3151 3602 3153 3604
rect 3720 3603 3722 3617
rect 3736 3615 3738 3617
rect 3736 3603 3738 3605
rect 3752 3603 3754 3617
rect 3775 3612 3777 3617
rect 3780 3615 3782 3617
rect 3806 3615 3808 3617
rect 3771 3608 3777 3612
rect 3775 3603 3777 3608
rect 3780 3603 3782 3605
rect 3806 3603 3808 3605
rect 3827 3603 3829 3617
rect 3847 3612 3849 3617
rect 3852 3615 3854 3617
rect 3843 3608 3849 3612
rect 3847 3603 3849 3608
rect 3852 3603 3854 3605
rect 3870 3603 3872 3617
rect 2775 3593 2777 3595
rect 2791 3592 2793 3595
rect 2807 3593 2809 3595
rect 2830 3593 2832 3595
rect 2835 3592 2837 3595
rect 2861 3592 2863 3595
rect 2882 3592 2884 3595
rect 2902 3593 2904 3595
rect 2907 3592 2909 3595
rect 2925 3593 2927 3595
rect 2975 3592 2977 3594
rect 2861 3588 2862 3592
rect 2980 3589 2982 3594
rect 3056 3592 3058 3594
rect 3061 3589 3063 3594
rect 3146 3592 3148 3594
rect 3151 3589 3153 3594
rect 3920 3602 3922 3614
rect 3925 3612 3927 3614
rect 3925 3602 3927 3604
rect 4001 3602 4003 3614
rect 4006 3612 4008 3614
rect 4006 3602 4008 3604
rect 4091 3602 4093 3614
rect 4096 3612 4098 3614
rect 4096 3602 4098 3604
rect 3720 3593 3722 3595
rect 3736 3592 3738 3595
rect 3752 3593 3754 3595
rect 3775 3593 3777 3595
rect 3780 3592 3782 3595
rect 3806 3592 3808 3595
rect 3827 3592 3829 3595
rect 3847 3593 3849 3595
rect 3852 3592 3854 3595
rect 3870 3593 3872 3595
rect 3920 3592 3922 3594
rect 3311 3589 3313 3592
rect 3316 3589 3318 3592
rect 2791 3585 2793 3588
rect 2835 3585 2837 3588
rect 2861 3585 2863 3588
rect 2907 3585 2909 3588
rect 3806 3588 3807 3592
rect 3925 3589 3927 3594
rect 4001 3592 4003 3594
rect 4006 3589 4008 3594
rect 4091 3592 4093 3594
rect 4096 3589 4098 3594
rect 3736 3585 3738 3588
rect 3780 3585 3782 3588
rect 3806 3585 3808 3588
rect 3852 3585 3854 3588
rect 3311 3573 3313 3585
rect 3316 3583 3318 3585
rect 3316 3573 3318 3575
rect 2791 3564 2793 3567
rect 2835 3564 2837 3567
rect 2861 3564 2863 3567
rect 2907 3564 2909 3567
rect 2975 3564 2977 3568
rect 3003 3570 3005 3572
rect 2980 3564 2982 3567
rect 2861 3560 2862 3564
rect 2775 3557 2777 3559
rect 2791 3557 2793 3560
rect 2807 3557 2809 3559
rect 2830 3557 2832 3559
rect 2835 3557 2837 3560
rect 2861 3557 2863 3560
rect 2882 3557 2884 3560
rect 2902 3557 2904 3559
rect 2907 3557 2909 3560
rect 2925 3557 2927 3559
rect 3311 3563 3313 3565
rect 2975 3553 2977 3556
rect 2980 3554 2982 3556
rect 2976 3549 2977 3553
rect 2775 3535 2777 3549
rect 2791 3547 2793 3549
rect 2791 3535 2793 3537
rect 2807 3535 2809 3549
rect 2830 3544 2832 3549
rect 2835 3547 2837 3549
rect 2861 3547 2863 3549
rect 2826 3540 2832 3544
rect 2830 3535 2832 3540
rect 2835 3535 2837 3537
rect 2861 3535 2863 3537
rect 2882 3535 2884 3549
rect 2902 3544 2904 3549
rect 2907 3547 2909 3549
rect 2898 3540 2904 3544
rect 2902 3535 2904 3540
rect 2907 3535 2909 3537
rect 2925 3535 2927 3549
rect 2975 3544 2977 3549
rect 2980 3544 2982 3546
rect 3003 3540 3005 3562
rect 3316 3560 3318 3565
rect 3736 3564 3738 3567
rect 3780 3564 3782 3567
rect 3806 3564 3808 3567
rect 3852 3564 3854 3567
rect 3920 3564 3922 3568
rect 3948 3570 3950 3572
rect 3925 3564 3927 3567
rect 3806 3560 3807 3564
rect 3720 3557 3722 3559
rect 3736 3557 3738 3560
rect 3752 3557 3754 3559
rect 3775 3557 3777 3559
rect 3780 3557 3782 3560
rect 3806 3557 3808 3560
rect 3827 3557 3829 3560
rect 3847 3557 3849 3559
rect 3852 3557 3854 3560
rect 3870 3557 3872 3559
rect 3920 3553 3922 3556
rect 3925 3554 3927 3556
rect 3921 3549 3922 3553
rect 2975 3538 2977 3540
rect 2980 3535 2982 3540
rect 3003 3534 3005 3536
rect 3720 3535 3722 3549
rect 3736 3547 3738 3549
rect 3736 3535 3738 3537
rect 3752 3535 3754 3549
rect 3775 3544 3777 3549
rect 3780 3547 3782 3549
rect 3806 3547 3808 3549
rect 3771 3540 3777 3544
rect 3775 3535 3777 3540
rect 3780 3535 3782 3537
rect 3806 3535 3808 3537
rect 3827 3535 3829 3549
rect 3847 3544 3849 3549
rect 3852 3547 3854 3549
rect 3843 3540 3849 3544
rect 3847 3535 3849 3540
rect 3852 3535 3854 3537
rect 3870 3535 3872 3549
rect 3920 3544 3922 3549
rect 3925 3544 3927 3546
rect 3948 3540 3950 3562
rect 3920 3538 3922 3540
rect 3925 3535 3927 3540
rect 3948 3534 3950 3536
rect 2775 3529 2777 3531
rect 2791 3527 2793 3531
rect 2807 3529 2809 3531
rect 2830 3529 2832 3531
rect 2792 3523 2793 3527
rect 2835 3526 2837 3531
rect 2861 3527 2863 3531
rect 2882 3529 2884 3531
rect 2902 3529 2904 3531
rect 2791 3520 2793 3523
rect 2836 3522 2837 3526
rect 2862 3523 2863 3527
rect 2907 3526 2909 3531
rect 2925 3529 2927 3531
rect 3720 3529 3722 3531
rect 3736 3527 3738 3531
rect 3752 3529 3754 3531
rect 3775 3529 3777 3531
rect 2835 3520 2837 3522
rect 2861 3519 2863 3523
rect 2908 3522 2909 3526
rect 3737 3523 3738 3527
rect 3780 3526 3782 3531
rect 3806 3527 3808 3531
rect 3827 3529 3829 3531
rect 3847 3529 3849 3531
rect 2907 3520 2909 3522
rect 3736 3520 3738 3523
rect 3781 3522 3782 3526
rect 3807 3523 3808 3527
rect 3852 3526 3854 3531
rect 3870 3529 3872 3531
rect 3780 3520 3782 3522
rect 3806 3519 3808 3523
rect 3853 3522 3854 3526
rect 3852 3520 3854 3522
rect 2286 3502 2288 3504
rect 2291 3502 2293 3505
rect 2307 3502 2309 3504
rect 2323 3502 2325 3504
rect 2328 3502 2330 3505
rect 2349 3502 2351 3505
rect 2365 3502 2367 3505
rect 2381 3502 2383 3504
rect 2386 3502 2388 3505
rect 2402 3502 2404 3504
rect 2418 3502 2420 3504
rect 2423 3502 2425 3505
rect 2439 3502 2441 3504
rect 2455 3502 2457 3504
rect 2460 3502 2462 3505
rect 2481 3502 2483 3505
rect 2497 3502 2499 3505
rect 2513 3502 2515 3504
rect 2518 3502 2520 3505
rect 2534 3502 2536 3504
rect 2550 3502 2552 3504
rect 2555 3502 2557 3505
rect 2571 3502 2573 3504
rect 2587 3502 2589 3504
rect 2592 3502 2594 3505
rect 2613 3502 2615 3505
rect 2629 3502 2631 3505
rect 2645 3502 2647 3504
rect 2650 3502 2652 3505
rect 2666 3502 2668 3504
rect 3231 3502 3233 3504
rect 3236 3502 3238 3505
rect 3252 3502 3254 3504
rect 3268 3502 3270 3504
rect 3273 3502 3275 3505
rect 3294 3502 3296 3505
rect 3310 3502 3312 3505
rect 3326 3502 3328 3504
rect 3331 3502 3333 3505
rect 3347 3502 3349 3504
rect 3363 3502 3365 3504
rect 3368 3502 3370 3505
rect 3384 3502 3386 3504
rect 3400 3502 3402 3504
rect 3405 3502 3407 3505
rect 3426 3502 3428 3505
rect 3442 3502 3444 3505
rect 3458 3502 3460 3504
rect 3463 3502 3465 3505
rect 3479 3502 3481 3504
rect 3495 3502 3497 3504
rect 3500 3502 3502 3505
rect 3516 3502 3518 3504
rect 3532 3502 3534 3504
rect 3537 3502 3539 3505
rect 3558 3502 3560 3505
rect 3574 3502 3576 3505
rect 3590 3502 3592 3504
rect 3595 3502 3597 3505
rect 3611 3502 3613 3504
rect 2791 3497 2793 3500
rect 2835 3498 2837 3500
rect 2286 3489 2288 3494
rect 2291 3492 2293 3494
rect 2286 3475 2288 3485
rect 2291 3475 2293 3482
rect 2307 3475 2309 3494
rect 2323 3485 2325 3494
rect 2328 3492 2330 3494
rect 2349 3492 2351 3494
rect 2365 3491 2367 3494
rect 2323 3475 2325 3478
rect 2328 3475 2330 3477
rect 2349 3475 2351 3477
rect 2365 3475 2367 3487
rect 2381 3485 2383 3494
rect 2386 3492 2388 3494
rect 2381 3475 2383 3478
rect 2386 3475 2388 3477
rect 2402 3475 2404 3494
rect 2418 3491 2420 3494
rect 2423 3492 2425 3494
rect 2418 3475 2420 3487
rect 2423 3475 2425 3482
rect 2439 3475 2441 3494
rect 2455 3485 2457 3494
rect 2460 3492 2462 3494
rect 2481 3492 2483 3494
rect 2497 3491 2499 3494
rect 2455 3475 2457 3478
rect 2460 3475 2462 3477
rect 2481 3475 2483 3477
rect 2497 3475 2499 3487
rect 2513 3485 2515 3494
rect 2518 3492 2520 3494
rect 2513 3475 2515 3478
rect 2518 3475 2520 3477
rect 2534 3475 2536 3494
rect 2550 3491 2552 3494
rect 2555 3492 2557 3494
rect 2550 3475 2552 3487
rect 2555 3475 2557 3482
rect 2571 3475 2573 3494
rect 2587 3485 2589 3494
rect 2592 3492 2594 3494
rect 2613 3492 2615 3494
rect 2629 3491 2631 3494
rect 2587 3475 2589 3478
rect 2592 3475 2594 3477
rect 2613 3475 2615 3477
rect 2629 3475 2631 3487
rect 2645 3485 2647 3494
rect 2650 3492 2652 3494
rect 2666 3486 2668 3494
rect 2792 3493 2793 3497
rect 2836 3494 2837 3498
rect 2861 3497 2863 3501
rect 2907 3498 2909 3500
rect 2775 3489 2777 3491
rect 2791 3489 2793 3493
rect 2807 3489 2809 3491
rect 2830 3489 2832 3491
rect 2835 3489 2837 3494
rect 2862 3493 2863 3497
rect 2908 3494 2909 3498
rect 3052 3497 3054 3500
rect 3096 3498 3098 3500
rect 2861 3489 2863 3493
rect 2882 3489 2884 3491
rect 2902 3489 2904 3491
rect 2907 3489 2909 3494
rect 3053 3493 3054 3497
rect 3097 3494 3098 3498
rect 3122 3497 3124 3501
rect 3168 3498 3170 3500
rect 2925 3489 2927 3491
rect 3009 3489 3011 3492
rect 3027 3489 3029 3492
rect 3052 3489 3054 3493
rect 3068 3489 3070 3491
rect 3091 3489 3093 3491
rect 3096 3489 3098 3494
rect 3123 3493 3124 3497
rect 3169 3494 3170 3498
rect 3736 3497 3738 3500
rect 3780 3498 3782 3500
rect 3122 3489 3124 3493
rect 3143 3489 3145 3491
rect 3163 3489 3165 3491
rect 3168 3489 3170 3494
rect 3186 3489 3188 3491
rect 3231 3489 3233 3494
rect 3236 3492 3238 3494
rect 2645 3475 2647 3478
rect 2650 3475 2652 3477
rect 2666 3475 2668 3482
rect 2775 3471 2777 3485
rect 2791 3483 2793 3485
rect 2791 3471 2793 3473
rect 2807 3471 2809 3485
rect 2830 3480 2832 3485
rect 2835 3483 2837 3485
rect 2861 3483 2863 3485
rect 2826 3476 2832 3480
rect 2830 3471 2832 3476
rect 2835 3471 2837 3473
rect 2861 3471 2863 3473
rect 2882 3471 2884 3485
rect 2902 3480 2904 3485
rect 2907 3483 2909 3485
rect 2898 3476 2904 3480
rect 2902 3471 2904 3476
rect 2907 3471 2909 3473
rect 2925 3471 2927 3485
rect 2975 3482 2977 3485
rect 2980 3482 2982 3485
rect 3009 3480 3011 3485
rect 2286 3469 2288 3471
rect 2291 3468 2293 3471
rect 2307 3469 2309 3471
rect 2323 3469 2325 3471
rect 2328 3466 2330 3471
rect 2349 3466 2351 3471
rect 2365 3469 2367 3471
rect 2381 3469 2383 3471
rect 2386 3466 2388 3471
rect 2402 3469 2404 3471
rect 2418 3469 2420 3471
rect 2423 3468 2425 3471
rect 2439 3469 2441 3471
rect 2455 3469 2457 3471
rect 2460 3466 2462 3471
rect 2481 3466 2483 3471
rect 2497 3469 2499 3471
rect 2513 3469 2515 3471
rect 2518 3466 2520 3471
rect 2534 3469 2536 3471
rect 2550 3469 2552 3471
rect 2555 3468 2557 3471
rect 2571 3469 2573 3471
rect 2587 3469 2589 3471
rect 2592 3466 2594 3471
rect 2613 3466 2615 3471
rect 2629 3469 2631 3471
rect 2645 3469 2647 3471
rect 2650 3466 2652 3471
rect 2666 3469 2668 3471
rect 2975 3466 2977 3478
rect 2980 3476 2982 3478
rect 3009 3471 3011 3476
rect 3027 3471 3029 3485
rect 3052 3483 3054 3485
rect 3052 3471 3054 3473
rect 3068 3471 3070 3485
rect 3091 3480 3093 3485
rect 3096 3483 3098 3485
rect 3122 3483 3124 3485
rect 3087 3476 3093 3480
rect 3091 3471 3093 3476
rect 3096 3471 3098 3473
rect 3122 3471 3124 3473
rect 3143 3471 3145 3485
rect 3163 3480 3165 3485
rect 3168 3483 3170 3485
rect 3159 3476 3165 3480
rect 3163 3471 3165 3476
rect 3168 3471 3170 3473
rect 3186 3471 3188 3485
rect 3231 3475 3233 3485
rect 3236 3475 3238 3482
rect 3252 3475 3254 3494
rect 3268 3485 3270 3494
rect 3273 3492 3275 3494
rect 3294 3492 3296 3494
rect 3310 3491 3312 3494
rect 3268 3475 3270 3478
rect 3273 3475 3275 3477
rect 3294 3475 3296 3477
rect 3310 3475 3312 3487
rect 3326 3485 3328 3494
rect 3331 3492 3333 3494
rect 3326 3475 3328 3478
rect 3331 3475 3333 3477
rect 3347 3475 3349 3494
rect 3363 3491 3365 3494
rect 3368 3492 3370 3494
rect 3363 3475 3365 3487
rect 3368 3475 3370 3482
rect 3384 3475 3386 3494
rect 3400 3485 3402 3494
rect 3405 3492 3407 3494
rect 3426 3492 3428 3494
rect 3442 3491 3444 3494
rect 3400 3475 3402 3478
rect 3405 3475 3407 3477
rect 3426 3475 3428 3477
rect 3442 3475 3444 3487
rect 3458 3485 3460 3494
rect 3463 3492 3465 3494
rect 3458 3475 3460 3478
rect 3463 3475 3465 3477
rect 3479 3475 3481 3494
rect 3495 3491 3497 3494
rect 3500 3492 3502 3494
rect 3495 3475 3497 3487
rect 3500 3475 3502 3482
rect 3516 3475 3518 3494
rect 3532 3485 3534 3494
rect 3537 3492 3539 3494
rect 3558 3492 3560 3494
rect 3574 3491 3576 3494
rect 3532 3475 3534 3478
rect 3537 3475 3539 3477
rect 3558 3475 3560 3477
rect 3574 3475 3576 3487
rect 3590 3485 3592 3494
rect 3595 3492 3597 3494
rect 3611 3486 3613 3494
rect 3737 3493 3738 3497
rect 3781 3494 3782 3498
rect 3806 3497 3808 3501
rect 3852 3498 3854 3500
rect 3720 3489 3722 3491
rect 3736 3489 3738 3493
rect 3752 3489 3754 3491
rect 3775 3489 3777 3491
rect 3780 3489 3782 3494
rect 3807 3493 3808 3497
rect 3853 3494 3854 3498
rect 3997 3497 3999 3500
rect 4041 3498 4043 3500
rect 3806 3489 3808 3493
rect 3827 3489 3829 3491
rect 3847 3489 3849 3491
rect 3852 3489 3854 3494
rect 3998 3493 3999 3497
rect 4042 3494 4043 3498
rect 4067 3497 4069 3501
rect 4113 3498 4115 3500
rect 3870 3489 3872 3491
rect 3954 3489 3956 3492
rect 3972 3489 3974 3492
rect 3997 3489 3999 3493
rect 4013 3489 4015 3491
rect 4036 3489 4038 3491
rect 4041 3489 4043 3494
rect 4068 3493 4069 3497
rect 4114 3494 4115 3498
rect 4067 3489 4069 3493
rect 4088 3489 4090 3491
rect 4108 3489 4110 3491
rect 4113 3489 4115 3494
rect 4131 3489 4133 3491
rect 3590 3475 3592 3478
rect 3595 3475 3597 3477
rect 3611 3475 3613 3482
rect 3720 3471 3722 3485
rect 3736 3483 3738 3485
rect 3736 3471 3738 3473
rect 3752 3471 3754 3485
rect 3775 3480 3777 3485
rect 3780 3483 3782 3485
rect 3806 3483 3808 3485
rect 3771 3476 3777 3480
rect 3775 3471 3777 3476
rect 3780 3471 3782 3473
rect 3806 3471 3808 3473
rect 3827 3471 3829 3485
rect 3847 3480 3849 3485
rect 3852 3483 3854 3485
rect 3843 3476 3849 3480
rect 3847 3471 3849 3476
rect 3852 3471 3854 3473
rect 3870 3471 3872 3485
rect 3920 3482 3922 3485
rect 3925 3482 3927 3485
rect 3954 3480 3956 3485
rect 2980 3466 2982 3468
rect 2775 3461 2777 3463
rect 2791 3460 2793 3463
rect 2807 3461 2809 3463
rect 2830 3461 2832 3463
rect 2835 3460 2837 3463
rect 2861 3460 2863 3463
rect 2882 3460 2884 3463
rect 2902 3461 2904 3463
rect 2907 3460 2909 3463
rect 2925 3461 2927 3463
rect 2861 3456 2862 3460
rect 3231 3469 3233 3471
rect 3236 3468 3238 3471
rect 3252 3469 3254 3471
rect 3268 3469 3270 3471
rect 3273 3466 3275 3471
rect 3294 3466 3296 3471
rect 3310 3469 3312 3471
rect 3326 3469 3328 3471
rect 3331 3466 3333 3471
rect 3347 3469 3349 3471
rect 3363 3469 3365 3471
rect 3009 3460 3011 3463
rect 2975 3456 2977 3458
rect 2791 3453 2793 3456
rect 2835 3453 2837 3456
rect 2861 3453 2863 3456
rect 2907 3453 2909 3456
rect 2980 3453 2982 3458
rect 2401 3431 2403 3434
rect 2425 3431 2427 3434
rect 2401 3424 2403 3427
rect 2425 3424 2427 3427
rect 3027 3421 3029 3463
rect 3052 3460 3054 3463
rect 3068 3461 3070 3463
rect 3091 3461 3093 3463
rect 3096 3460 3098 3463
rect 3122 3460 3124 3463
rect 3143 3460 3145 3463
rect 3163 3461 3165 3463
rect 3168 3460 3170 3463
rect 3186 3461 3188 3463
rect 3368 3468 3370 3471
rect 3384 3469 3386 3471
rect 3400 3469 3402 3471
rect 3405 3466 3407 3471
rect 3426 3466 3428 3471
rect 3442 3469 3444 3471
rect 3458 3469 3460 3471
rect 3463 3466 3465 3471
rect 3479 3469 3481 3471
rect 3495 3469 3497 3471
rect 3500 3468 3502 3471
rect 3516 3469 3518 3471
rect 3532 3469 3534 3471
rect 3537 3466 3539 3471
rect 3558 3466 3560 3471
rect 3574 3469 3576 3471
rect 3590 3469 3592 3471
rect 3595 3466 3597 3471
rect 3611 3469 3613 3471
rect 3920 3466 3922 3478
rect 3925 3476 3927 3478
rect 3954 3471 3956 3476
rect 3972 3471 3974 3485
rect 3997 3483 3999 3485
rect 3997 3471 3999 3473
rect 4013 3471 4015 3485
rect 4036 3480 4038 3485
rect 4041 3483 4043 3485
rect 4067 3483 4069 3485
rect 4032 3476 4038 3480
rect 4036 3471 4038 3476
rect 4041 3471 4043 3473
rect 4067 3471 4069 3473
rect 4088 3471 4090 3485
rect 4108 3480 4110 3485
rect 4113 3483 4115 3485
rect 4104 3476 4110 3480
rect 4108 3471 4110 3476
rect 4113 3471 4115 3473
rect 4131 3471 4133 3485
rect 3925 3466 3927 3468
rect 3720 3461 3722 3463
rect 3736 3460 3738 3463
rect 3752 3461 3754 3463
rect 3775 3461 3777 3463
rect 3780 3460 3782 3463
rect 3806 3460 3808 3463
rect 3827 3460 3829 3463
rect 3847 3461 3849 3463
rect 3852 3460 3854 3463
rect 3870 3461 3872 3463
rect 3122 3456 3123 3460
rect 3052 3453 3054 3456
rect 3096 3453 3098 3456
rect 3122 3453 3124 3456
rect 3168 3453 3170 3456
rect 3806 3456 3807 3460
rect 3954 3460 3956 3463
rect 3920 3456 3922 3458
rect 3736 3453 3738 3456
rect 3780 3453 3782 3456
rect 3806 3453 3808 3456
rect 3852 3453 3854 3456
rect 3925 3453 3927 3458
rect 3346 3431 3348 3434
rect 3370 3431 3372 3434
rect 3195 3429 3198 3431
rect 3202 3429 3205 3431
rect 3346 3424 3348 3427
rect 3370 3424 3372 3427
rect 3972 3425 3974 3463
rect 3997 3460 3999 3463
rect 4013 3461 4015 3463
rect 4036 3461 4038 3463
rect 4041 3460 4043 3463
rect 4067 3460 4069 3463
rect 4088 3460 4090 3463
rect 4108 3461 4110 3463
rect 4113 3460 4115 3463
rect 4131 3461 4133 3463
rect 4067 3456 4068 3460
rect 3997 3453 3999 3456
rect 4041 3453 4043 3456
rect 4067 3453 4069 3456
rect 4113 3453 4115 3456
rect 4140 3429 4143 3431
rect 4147 3429 4150 3431
rect 2421 3418 2423 3420
rect 3366 3418 3368 3420
rect 2421 3411 2423 3414
rect 3366 3411 3368 3414
rect 2410 3400 2412 3402
rect 2416 3400 2435 3402
rect 3355 3400 3357 3402
rect 3361 3400 3380 3402
rect 2401 3395 2403 3397
rect 2425 3395 2427 3397
rect 3346 3395 3348 3397
rect 3370 3395 3372 3397
rect 2401 3388 2403 3391
rect 2425 3388 2427 3391
rect 3069 3390 3071 3392
rect 3074 3390 3076 3393
rect 3090 3390 3092 3392
rect 3106 3390 3108 3392
rect 3111 3390 3113 3393
rect 3132 3390 3134 3393
rect 3148 3390 3150 3393
rect 3164 3390 3166 3392
rect 3169 3390 3171 3393
rect 3185 3390 3187 3392
rect 3346 3388 3348 3391
rect 3370 3388 3372 3391
rect 4014 3390 4016 3392
rect 4019 3390 4021 3393
rect 4035 3390 4037 3392
rect 4051 3390 4053 3392
rect 4056 3390 4058 3393
rect 4077 3390 4079 3393
rect 4093 3390 4095 3393
rect 4109 3390 4111 3392
rect 4114 3390 4116 3393
rect 4130 3390 4132 3392
rect 3069 3377 3071 3382
rect 3074 3380 3076 3382
rect 3069 3363 3071 3373
rect 3074 3363 3076 3370
rect 3090 3363 3092 3382
rect 3106 3373 3108 3382
rect 3111 3380 3113 3382
rect 3132 3380 3134 3382
rect 3148 3379 3150 3382
rect 3106 3363 3108 3366
rect 3111 3363 3113 3365
rect 3132 3363 3134 3365
rect 3148 3363 3150 3375
rect 3164 3373 3166 3382
rect 3169 3380 3171 3382
rect 3164 3363 3166 3366
rect 3169 3363 3171 3365
rect 3185 3363 3187 3382
rect 4014 3377 4016 3382
rect 4019 3380 4021 3382
rect 4014 3363 4016 3373
rect 4019 3363 4021 3370
rect 4035 3363 4037 3382
rect 4051 3373 4053 3382
rect 4056 3380 4058 3382
rect 4077 3380 4079 3382
rect 4093 3379 4095 3382
rect 4051 3363 4053 3366
rect 4056 3363 4058 3365
rect 4077 3363 4079 3365
rect 4093 3363 4095 3375
rect 4109 3373 4111 3382
rect 4114 3380 4116 3382
rect 4109 3363 4111 3366
rect 4114 3363 4116 3365
rect 4130 3363 4132 3382
rect 2286 3360 2288 3362
rect 2291 3360 2293 3363
rect 2307 3360 2309 3362
rect 2323 3360 2325 3362
rect 2328 3360 2330 3363
rect 2349 3360 2351 3363
rect 2365 3360 2367 3363
rect 2381 3360 2383 3362
rect 2386 3360 2388 3363
rect 2402 3360 2404 3362
rect 2418 3360 2420 3362
rect 2423 3360 2425 3363
rect 2439 3360 2441 3362
rect 2455 3360 2457 3362
rect 2460 3360 2462 3363
rect 2481 3360 2483 3363
rect 2497 3360 2499 3363
rect 2513 3360 2515 3362
rect 2518 3360 2520 3363
rect 2534 3360 2536 3362
rect 2550 3360 2552 3362
rect 2555 3360 2557 3363
rect 2571 3360 2573 3362
rect 2587 3360 2589 3362
rect 2592 3360 2594 3363
rect 2613 3360 2615 3363
rect 2629 3360 2631 3363
rect 2645 3360 2647 3362
rect 2650 3360 2652 3363
rect 2666 3360 2668 3362
rect 3231 3360 3233 3362
rect 3236 3360 3238 3363
rect 3252 3360 3254 3362
rect 3268 3360 3270 3362
rect 3273 3360 3275 3363
rect 3294 3360 3296 3363
rect 3310 3360 3312 3363
rect 3326 3360 3328 3362
rect 3331 3360 3333 3363
rect 3347 3360 3349 3362
rect 3363 3360 3365 3362
rect 3368 3360 3370 3363
rect 3384 3360 3386 3362
rect 3400 3360 3402 3362
rect 3405 3360 3407 3363
rect 3426 3360 3428 3363
rect 3442 3360 3444 3363
rect 3458 3360 3460 3362
rect 3463 3360 3465 3363
rect 3479 3360 3481 3362
rect 3495 3360 3497 3362
rect 3500 3360 3502 3363
rect 3516 3360 3518 3362
rect 3532 3360 3534 3362
rect 3537 3360 3539 3363
rect 3558 3360 3560 3363
rect 3574 3360 3576 3363
rect 3590 3360 3592 3362
rect 3595 3360 3597 3363
rect 3611 3360 3613 3362
rect 3069 3357 3071 3359
rect 3074 3356 3076 3359
rect 3090 3357 3092 3359
rect 3106 3357 3108 3359
rect 3111 3354 3113 3359
rect 3132 3354 3134 3359
rect 3148 3357 3150 3359
rect 3164 3357 3166 3359
rect 3169 3354 3171 3359
rect 3185 3357 3187 3359
rect 2286 3347 2288 3352
rect 2291 3350 2293 3352
rect 2286 3333 2288 3343
rect 2291 3333 2293 3340
rect 2307 3333 2309 3352
rect 2323 3343 2325 3352
rect 2328 3350 2330 3352
rect 2349 3350 2351 3352
rect 2365 3349 2367 3352
rect 2323 3333 2325 3336
rect 2328 3333 2330 3335
rect 2349 3333 2351 3335
rect 2365 3333 2367 3345
rect 2381 3343 2383 3352
rect 2386 3350 2388 3352
rect 2381 3333 2383 3336
rect 2386 3333 2388 3335
rect 2402 3333 2404 3352
rect 2418 3349 2420 3352
rect 2423 3350 2425 3352
rect 2418 3333 2420 3345
rect 2423 3333 2425 3340
rect 2439 3333 2441 3352
rect 2455 3343 2457 3352
rect 2460 3350 2462 3352
rect 2481 3350 2483 3352
rect 2497 3349 2499 3352
rect 2455 3333 2457 3336
rect 2460 3333 2462 3335
rect 2481 3333 2483 3335
rect 2497 3333 2499 3345
rect 2513 3343 2515 3352
rect 2518 3350 2520 3352
rect 2513 3333 2515 3336
rect 2518 3333 2520 3335
rect 2534 3333 2536 3352
rect 2550 3349 2552 3352
rect 2555 3350 2557 3352
rect 2550 3333 2552 3345
rect 2555 3333 2557 3340
rect 2571 3333 2573 3352
rect 2587 3343 2589 3352
rect 2592 3350 2594 3352
rect 2613 3350 2615 3352
rect 2629 3349 2631 3352
rect 2587 3333 2589 3336
rect 2592 3333 2594 3335
rect 2613 3333 2615 3335
rect 2629 3333 2631 3345
rect 2645 3343 2647 3352
rect 2650 3350 2652 3352
rect 2666 3344 2668 3352
rect 4014 3357 4016 3359
rect 4019 3356 4021 3359
rect 4035 3357 4037 3359
rect 4051 3357 4053 3359
rect 4056 3354 4058 3359
rect 4077 3354 4079 3359
rect 4093 3357 4095 3359
rect 4109 3357 4111 3359
rect 4114 3354 4116 3359
rect 4130 3357 4132 3359
rect 3231 3347 3233 3352
rect 3236 3350 3238 3352
rect 2645 3333 2647 3336
rect 2650 3333 2652 3335
rect 2666 3333 2668 3340
rect 3231 3333 3233 3343
rect 3236 3333 3238 3340
rect 3252 3333 3254 3352
rect 3268 3343 3270 3352
rect 3273 3350 3275 3352
rect 3294 3350 3296 3352
rect 3310 3349 3312 3352
rect 3268 3333 3270 3336
rect 3273 3333 3275 3335
rect 3294 3333 3296 3335
rect 3310 3333 3312 3345
rect 3326 3343 3328 3352
rect 3331 3350 3333 3352
rect 3326 3333 3328 3336
rect 3331 3333 3333 3335
rect 3347 3333 3349 3352
rect 3363 3349 3365 3352
rect 3368 3350 3370 3352
rect 3363 3333 3365 3345
rect 3368 3333 3370 3340
rect 3384 3333 3386 3352
rect 3400 3343 3402 3352
rect 3405 3350 3407 3352
rect 3426 3350 3428 3352
rect 3442 3349 3444 3352
rect 3400 3333 3402 3336
rect 3405 3333 3407 3335
rect 3426 3333 3428 3335
rect 3442 3333 3444 3345
rect 3458 3343 3460 3352
rect 3463 3350 3465 3352
rect 3458 3333 3460 3336
rect 3463 3333 3465 3335
rect 3479 3333 3481 3352
rect 3495 3349 3497 3352
rect 3500 3350 3502 3352
rect 3495 3333 3497 3345
rect 3500 3333 3502 3340
rect 3516 3333 3518 3352
rect 3532 3343 3534 3352
rect 3537 3350 3539 3352
rect 3558 3350 3560 3352
rect 3574 3349 3576 3352
rect 3532 3333 3534 3336
rect 3537 3333 3539 3335
rect 3558 3333 3560 3335
rect 3574 3333 3576 3345
rect 3590 3343 3592 3352
rect 3595 3350 3597 3352
rect 3611 3344 3613 3352
rect 3590 3333 3592 3336
rect 3595 3333 3597 3335
rect 3611 3333 3613 3340
rect 2286 3327 2288 3329
rect 2291 3326 2293 3329
rect 2307 3327 2309 3329
rect 2323 3327 2325 3329
rect 2328 3324 2330 3329
rect 2349 3324 2351 3329
rect 2365 3327 2367 3329
rect 2381 3327 2383 3329
rect 2386 3324 2388 3329
rect 2402 3327 2404 3329
rect 2418 3327 2420 3329
rect 2423 3326 2425 3329
rect 2439 3327 2441 3329
rect 2455 3327 2457 3329
rect 2460 3324 2462 3329
rect 2481 3324 2483 3329
rect 2497 3327 2499 3329
rect 2513 3327 2515 3329
rect 2518 3324 2520 3329
rect 2534 3327 2536 3329
rect 2550 3327 2552 3329
rect 2555 3326 2557 3329
rect 2571 3327 2573 3329
rect 2587 3327 2589 3329
rect 2592 3324 2594 3329
rect 2613 3324 2615 3329
rect 2629 3327 2631 3329
rect 2645 3327 2647 3329
rect 2650 3324 2652 3329
rect 2666 3327 2668 3329
rect 3231 3327 3233 3329
rect 3236 3326 3238 3329
rect 3252 3327 3254 3329
rect 3268 3327 3270 3329
rect 3273 3324 3275 3329
rect 3294 3324 3296 3329
rect 3310 3327 3312 3329
rect 3326 3327 3328 3329
rect 3331 3324 3333 3329
rect 3347 3327 3349 3329
rect 3363 3327 3365 3329
rect 3368 3326 3370 3329
rect 3384 3327 3386 3329
rect 3400 3327 3402 3329
rect 3405 3324 3407 3329
rect 3426 3324 3428 3329
rect 3442 3327 3444 3329
rect 3458 3327 3460 3329
rect 3463 3324 3465 3329
rect 3479 3327 3481 3329
rect 3495 3327 3497 3329
rect 3500 3326 3502 3329
rect 3516 3327 3518 3329
rect 3532 3327 3534 3329
rect 3537 3324 3539 3329
rect 3558 3324 3560 3329
rect 3574 3327 3576 3329
rect 3590 3327 3592 3329
rect 3595 3324 3597 3329
rect 3611 3327 3613 3329
rect 3069 3304 3071 3306
rect 3074 3304 3076 3307
rect 3090 3304 3092 3306
rect 3106 3304 3108 3306
rect 3111 3304 3113 3307
rect 3132 3304 3134 3307
rect 3148 3304 3150 3307
rect 3164 3304 3166 3306
rect 3169 3304 3171 3307
rect 3185 3304 3187 3306
rect 4014 3304 4016 3306
rect 4019 3304 4021 3307
rect 4035 3304 4037 3306
rect 4051 3304 4053 3306
rect 4056 3304 4058 3307
rect 4077 3304 4079 3307
rect 4093 3304 4095 3307
rect 4109 3304 4111 3306
rect 4114 3304 4116 3307
rect 4130 3304 4132 3306
rect 3069 3291 3071 3296
rect 3074 3294 3076 3296
rect 3069 3277 3071 3287
rect 3074 3277 3076 3284
rect 3090 3277 3092 3296
rect 3106 3287 3108 3296
rect 3111 3294 3113 3296
rect 3132 3294 3134 3296
rect 3148 3293 3150 3296
rect 3106 3277 3108 3280
rect 3111 3277 3113 3279
rect 3132 3277 3134 3279
rect 3148 3277 3150 3289
rect 3164 3287 3166 3296
rect 3169 3294 3171 3296
rect 3164 3277 3166 3280
rect 3169 3277 3171 3279
rect 3185 3277 3187 3296
rect 4014 3291 4016 3296
rect 4019 3294 4021 3296
rect 3207 3283 3210 3285
rect 3214 3283 3217 3285
rect 4014 3277 4016 3287
rect 4019 3277 4021 3284
rect 4035 3277 4037 3296
rect 4051 3287 4053 3296
rect 4056 3294 4058 3296
rect 4077 3294 4079 3296
rect 4093 3293 4095 3296
rect 4051 3277 4053 3280
rect 4056 3277 4058 3279
rect 4077 3277 4079 3279
rect 4093 3277 4095 3289
rect 4109 3287 4111 3296
rect 4114 3294 4116 3296
rect 4109 3277 4111 3280
rect 4114 3277 4116 3279
rect 4130 3277 4132 3296
rect 4152 3283 4155 3285
rect 4159 3283 4162 3285
rect 2286 3274 2288 3276
rect 2291 3274 2293 3277
rect 2307 3274 2309 3276
rect 2323 3274 2325 3276
rect 2328 3274 2330 3277
rect 2349 3274 2351 3277
rect 2365 3274 2367 3277
rect 2381 3274 2383 3276
rect 2386 3274 2388 3277
rect 2402 3274 2404 3276
rect 2418 3274 2420 3276
rect 2423 3274 2425 3277
rect 2439 3274 2441 3276
rect 2455 3274 2457 3276
rect 2460 3274 2462 3277
rect 2481 3274 2483 3277
rect 2497 3274 2499 3277
rect 2513 3274 2515 3276
rect 2518 3274 2520 3277
rect 2534 3274 2536 3276
rect 2550 3274 2552 3276
rect 2555 3274 2557 3277
rect 2571 3274 2573 3276
rect 2587 3274 2589 3276
rect 2592 3274 2594 3277
rect 2613 3274 2615 3277
rect 2629 3274 2631 3277
rect 2645 3274 2647 3276
rect 2650 3274 2652 3277
rect 2666 3274 2668 3276
rect 3231 3274 3233 3276
rect 3236 3274 3238 3277
rect 3252 3274 3254 3276
rect 3268 3274 3270 3276
rect 3273 3274 3275 3277
rect 3294 3274 3296 3277
rect 3310 3274 3312 3277
rect 3326 3274 3328 3276
rect 3331 3274 3333 3277
rect 3347 3274 3349 3276
rect 3363 3274 3365 3276
rect 3368 3274 3370 3277
rect 3384 3274 3386 3276
rect 3400 3274 3402 3276
rect 3405 3274 3407 3277
rect 3426 3274 3428 3277
rect 3442 3274 3444 3277
rect 3458 3274 3460 3276
rect 3463 3274 3465 3277
rect 3479 3274 3481 3276
rect 3495 3274 3497 3276
rect 3500 3274 3502 3277
rect 3516 3274 3518 3276
rect 3532 3274 3534 3276
rect 3537 3274 3539 3277
rect 3558 3274 3560 3277
rect 3574 3274 3576 3277
rect 3590 3274 3592 3276
rect 3595 3274 3597 3277
rect 3611 3274 3613 3276
rect 3069 3271 3071 3273
rect 3074 3270 3076 3273
rect 3090 3271 3092 3273
rect 3106 3271 3108 3273
rect 3111 3268 3113 3273
rect 3132 3268 3134 3273
rect 3148 3271 3150 3273
rect 3164 3271 3166 3273
rect 3169 3268 3171 3273
rect 3185 3271 3187 3273
rect 2286 3261 2288 3266
rect 2291 3264 2293 3266
rect 2286 3247 2288 3257
rect 2291 3247 2293 3254
rect 2307 3247 2309 3266
rect 2323 3257 2325 3266
rect 2328 3264 2330 3266
rect 2349 3264 2351 3266
rect 2365 3263 2367 3266
rect 2323 3247 2325 3250
rect 2328 3247 2330 3249
rect 2349 3247 2351 3249
rect 2365 3247 2367 3259
rect 2381 3257 2383 3266
rect 2386 3264 2388 3266
rect 2381 3247 2383 3250
rect 2386 3247 2388 3249
rect 2402 3247 2404 3266
rect 2418 3263 2420 3266
rect 2423 3264 2425 3266
rect 2418 3247 2420 3259
rect 2423 3247 2425 3254
rect 2439 3247 2441 3266
rect 2455 3257 2457 3266
rect 2460 3264 2462 3266
rect 2481 3264 2483 3266
rect 2497 3263 2499 3266
rect 2455 3247 2457 3250
rect 2460 3247 2462 3249
rect 2481 3247 2483 3249
rect 2497 3247 2499 3259
rect 2513 3257 2515 3266
rect 2518 3264 2520 3266
rect 2513 3247 2515 3250
rect 2518 3247 2520 3249
rect 2534 3247 2536 3266
rect 2550 3263 2552 3266
rect 2555 3264 2557 3266
rect 2550 3247 2552 3259
rect 2555 3247 2557 3254
rect 2571 3247 2573 3266
rect 2587 3257 2589 3266
rect 2592 3264 2594 3266
rect 2613 3264 2615 3266
rect 2629 3263 2631 3266
rect 2587 3247 2589 3250
rect 2592 3247 2594 3249
rect 2613 3247 2615 3249
rect 2629 3247 2631 3259
rect 2645 3257 2647 3266
rect 2650 3264 2652 3266
rect 2666 3258 2668 3266
rect 4014 3271 4016 3273
rect 4019 3270 4021 3273
rect 4035 3271 4037 3273
rect 4051 3271 4053 3273
rect 4056 3268 4058 3273
rect 4077 3268 4079 3273
rect 4093 3271 4095 3273
rect 4109 3271 4111 3273
rect 4114 3268 4116 3273
rect 4130 3271 4132 3273
rect 3231 3261 3233 3266
rect 3236 3264 3238 3266
rect 2645 3247 2647 3250
rect 2650 3247 2652 3249
rect 2666 3247 2668 3254
rect 3231 3247 3233 3257
rect 3236 3247 3238 3254
rect 3252 3247 3254 3266
rect 3268 3257 3270 3266
rect 3273 3264 3275 3266
rect 3294 3264 3296 3266
rect 3310 3263 3312 3266
rect 3268 3247 3270 3250
rect 3273 3247 3275 3249
rect 3294 3247 3296 3249
rect 3310 3247 3312 3259
rect 3326 3257 3328 3266
rect 3331 3264 3333 3266
rect 3326 3247 3328 3250
rect 3331 3247 3333 3249
rect 3347 3247 3349 3266
rect 3363 3263 3365 3266
rect 3368 3264 3370 3266
rect 3363 3247 3365 3259
rect 3368 3247 3370 3254
rect 3384 3247 3386 3266
rect 3400 3257 3402 3266
rect 3405 3264 3407 3266
rect 3426 3264 3428 3266
rect 3442 3263 3444 3266
rect 3400 3247 3402 3250
rect 3405 3247 3407 3249
rect 3426 3247 3428 3249
rect 3442 3247 3444 3259
rect 3458 3257 3460 3266
rect 3463 3264 3465 3266
rect 3458 3247 3460 3250
rect 3463 3247 3465 3249
rect 3479 3247 3481 3266
rect 3495 3263 3497 3266
rect 3500 3264 3502 3266
rect 3495 3247 3497 3259
rect 3500 3247 3502 3254
rect 3516 3247 3518 3266
rect 3532 3257 3534 3266
rect 3537 3264 3539 3266
rect 3558 3264 3560 3266
rect 3574 3263 3576 3266
rect 3532 3247 3534 3250
rect 3537 3247 3539 3249
rect 3558 3247 3560 3249
rect 3574 3247 3576 3259
rect 3590 3257 3592 3266
rect 3595 3264 3597 3266
rect 3611 3258 3613 3266
rect 3590 3247 3592 3250
rect 3595 3247 3597 3249
rect 3611 3247 3613 3254
rect 2286 3241 2288 3243
rect 2291 3240 2293 3243
rect 2307 3241 2309 3243
rect 2323 3241 2325 3243
rect 2328 3238 2330 3243
rect 2349 3238 2351 3243
rect 2365 3241 2367 3243
rect 2381 3241 2383 3243
rect 2386 3238 2388 3243
rect 2402 3241 2404 3243
rect 2418 3241 2420 3243
rect 2423 3240 2425 3243
rect 2439 3241 2441 3243
rect 2455 3241 2457 3243
rect 2460 3238 2462 3243
rect 2481 3238 2483 3243
rect 2497 3241 2499 3243
rect 2513 3241 2515 3243
rect 2518 3238 2520 3243
rect 2534 3241 2536 3243
rect 2550 3241 2552 3243
rect 2555 3240 2557 3243
rect 2571 3241 2573 3243
rect 2587 3241 2589 3243
rect 2592 3238 2594 3243
rect 2613 3238 2615 3243
rect 2629 3241 2631 3243
rect 2645 3241 2647 3243
rect 2650 3238 2652 3243
rect 2666 3241 2668 3243
rect 3231 3241 3233 3243
rect 3236 3240 3238 3243
rect 3252 3241 3254 3243
rect 3268 3241 3270 3243
rect 3273 3238 3275 3243
rect 3294 3238 3296 3243
rect 3310 3241 3312 3243
rect 3326 3241 3328 3243
rect 3331 3238 3333 3243
rect 3347 3241 3349 3243
rect 3363 3241 3365 3243
rect 3368 3240 3370 3243
rect 3384 3241 3386 3243
rect 3400 3241 3402 3243
rect 3405 3238 3407 3243
rect 3426 3238 3428 3243
rect 3442 3241 3444 3243
rect 3458 3241 3460 3243
rect 3463 3238 3465 3243
rect 3479 3241 3481 3243
rect 3495 3241 3497 3243
rect 3500 3240 3502 3243
rect 3516 3241 3518 3243
rect 3532 3241 3534 3243
rect 3537 3238 3539 3243
rect 3558 3238 3560 3243
rect 3574 3241 3576 3243
rect 3590 3241 3592 3243
rect 3595 3238 3597 3243
rect 3611 3241 3613 3243
rect 2518 3203 2520 3206
rect 2542 3203 2544 3206
rect 3463 3203 3465 3206
rect 3487 3203 3489 3206
rect 2518 3197 2520 3199
rect 2542 3197 2544 3199
rect 3463 3197 3465 3199
rect 3487 3197 3489 3199
rect 2538 3192 2540 3194
rect 3483 3192 3485 3194
rect 2538 3185 2540 3188
rect 3483 3185 3485 3188
rect 2527 3174 2529 3176
rect 2533 3174 2552 3176
rect 3472 3174 3474 3176
rect 3478 3174 3497 3176
rect 2518 3169 2520 3171
rect 2542 3169 2544 3171
rect 3463 3169 3465 3171
rect 3487 3169 3489 3171
rect 2518 3162 2520 3165
rect 2542 3162 2544 3165
rect 3463 3162 3465 3165
rect 3487 3162 3489 3165
rect 2286 3134 2288 3136
rect 2291 3134 2293 3137
rect 2307 3134 2309 3136
rect 2323 3134 2325 3136
rect 2328 3134 2330 3137
rect 2349 3134 2351 3137
rect 2365 3134 2367 3137
rect 2381 3134 2383 3136
rect 2386 3134 2388 3137
rect 2402 3134 2404 3136
rect 2418 3134 2420 3136
rect 2423 3134 2425 3137
rect 2439 3134 2441 3136
rect 2455 3134 2457 3136
rect 2460 3134 2462 3137
rect 2481 3134 2483 3137
rect 2497 3134 2499 3137
rect 2513 3134 2515 3136
rect 2518 3134 2520 3137
rect 2534 3134 2536 3136
rect 2550 3134 2552 3136
rect 2555 3134 2557 3137
rect 2571 3134 2573 3136
rect 2587 3134 2589 3136
rect 2592 3134 2594 3137
rect 2613 3134 2615 3137
rect 2629 3134 2631 3137
rect 2645 3134 2647 3136
rect 2650 3134 2652 3137
rect 2666 3134 2668 3136
rect 3231 3134 3233 3136
rect 3236 3134 3238 3137
rect 3252 3134 3254 3136
rect 3268 3134 3270 3136
rect 3273 3134 3275 3137
rect 3294 3134 3296 3137
rect 3310 3134 3312 3137
rect 3326 3134 3328 3136
rect 3331 3134 3333 3137
rect 3347 3134 3349 3136
rect 3363 3134 3365 3136
rect 3368 3134 3370 3137
rect 3384 3134 3386 3136
rect 3400 3134 3402 3136
rect 3405 3134 3407 3137
rect 3426 3134 3428 3137
rect 3442 3134 3444 3137
rect 3458 3134 3460 3136
rect 3463 3134 3465 3137
rect 3479 3134 3481 3136
rect 3495 3134 3497 3136
rect 3500 3134 3502 3137
rect 3516 3134 3518 3136
rect 3532 3134 3534 3136
rect 3537 3134 3539 3137
rect 3558 3134 3560 3137
rect 3574 3134 3576 3137
rect 3590 3134 3592 3136
rect 3595 3134 3597 3137
rect 3611 3134 3613 3136
rect 2286 3121 2288 3126
rect 2291 3124 2293 3126
rect 2286 3107 2288 3117
rect 2291 3107 2293 3114
rect 2307 3107 2309 3126
rect 2323 3117 2325 3126
rect 2328 3124 2330 3126
rect 2349 3124 2351 3126
rect 2365 3123 2367 3126
rect 2323 3107 2325 3110
rect 2328 3107 2330 3109
rect 2349 3107 2351 3109
rect 2365 3107 2367 3119
rect 2381 3117 2383 3126
rect 2386 3124 2388 3126
rect 2381 3107 2383 3110
rect 2386 3107 2388 3109
rect 2402 3107 2404 3126
rect 2418 3123 2420 3126
rect 2423 3124 2425 3126
rect 2418 3107 2420 3119
rect 2423 3107 2425 3114
rect 2439 3107 2441 3126
rect 2455 3117 2457 3126
rect 2460 3124 2462 3126
rect 2481 3124 2483 3126
rect 2497 3123 2499 3126
rect 2455 3107 2457 3110
rect 2460 3107 2462 3109
rect 2481 3107 2483 3109
rect 2497 3107 2499 3119
rect 2513 3117 2515 3126
rect 2518 3124 2520 3126
rect 2513 3107 2515 3110
rect 2518 3107 2520 3109
rect 2534 3107 2536 3126
rect 2550 3123 2552 3126
rect 2555 3124 2557 3126
rect 2550 3107 2552 3119
rect 2555 3107 2557 3114
rect 2571 3107 2573 3126
rect 2587 3117 2589 3126
rect 2592 3124 2594 3126
rect 2613 3124 2615 3126
rect 2629 3123 2631 3126
rect 2587 3107 2589 3110
rect 2592 3107 2594 3109
rect 2613 3107 2615 3109
rect 2629 3107 2631 3119
rect 2645 3117 2647 3126
rect 2650 3124 2652 3126
rect 2666 3118 2668 3126
rect 3231 3121 3233 3126
rect 3236 3124 3238 3126
rect 2645 3107 2647 3110
rect 2650 3107 2652 3109
rect 2666 3107 2668 3114
rect 3231 3107 3233 3117
rect 3236 3107 3238 3114
rect 3252 3107 3254 3126
rect 3268 3117 3270 3126
rect 3273 3124 3275 3126
rect 3294 3124 3296 3126
rect 3310 3123 3312 3126
rect 3268 3107 3270 3110
rect 3273 3107 3275 3109
rect 3294 3107 3296 3109
rect 3310 3107 3312 3119
rect 3326 3117 3328 3126
rect 3331 3124 3333 3126
rect 3326 3107 3328 3110
rect 3331 3107 3333 3109
rect 3347 3107 3349 3126
rect 3363 3123 3365 3126
rect 3368 3124 3370 3126
rect 3363 3107 3365 3119
rect 3368 3107 3370 3114
rect 3384 3107 3386 3126
rect 3400 3117 3402 3126
rect 3405 3124 3407 3126
rect 3426 3124 3428 3126
rect 3442 3123 3444 3126
rect 3400 3107 3402 3110
rect 3405 3107 3407 3109
rect 3426 3107 3428 3109
rect 3442 3107 3444 3119
rect 3458 3117 3460 3126
rect 3463 3124 3465 3126
rect 3458 3107 3460 3110
rect 3463 3107 3465 3109
rect 3479 3107 3481 3126
rect 3495 3123 3497 3126
rect 3500 3124 3502 3126
rect 3495 3107 3497 3119
rect 3500 3107 3502 3114
rect 3516 3107 3518 3126
rect 3532 3117 3534 3126
rect 3537 3124 3539 3126
rect 3558 3124 3560 3126
rect 3574 3123 3576 3126
rect 3532 3107 3534 3110
rect 3537 3107 3539 3109
rect 3558 3107 3560 3109
rect 3574 3107 3576 3119
rect 3590 3117 3592 3126
rect 3595 3124 3597 3126
rect 3611 3118 3613 3126
rect 3590 3107 3592 3110
rect 3595 3107 3597 3109
rect 3611 3107 3613 3114
rect 2286 3101 2288 3103
rect 2291 3100 2293 3103
rect 2307 3101 2309 3103
rect 2323 3101 2325 3103
rect 2328 3098 2330 3103
rect 2349 3098 2351 3103
rect 2365 3101 2367 3103
rect 2381 3101 2383 3103
rect 2386 3098 2388 3103
rect 2402 3101 2404 3103
rect 2418 3101 2420 3103
rect 2423 3100 2425 3103
rect 2439 3101 2441 3103
rect 2455 3101 2457 3103
rect 2460 3098 2462 3103
rect 2481 3098 2483 3103
rect 2497 3101 2499 3103
rect 2513 3101 2515 3103
rect 2518 3098 2520 3103
rect 2534 3101 2536 3103
rect 2550 3101 2552 3103
rect 2555 3100 2557 3103
rect 2571 3101 2573 3103
rect 2587 3101 2589 3103
rect 2592 3098 2594 3103
rect 2613 3098 2615 3103
rect 2629 3101 2631 3103
rect 2645 3101 2647 3103
rect 2650 3098 2652 3103
rect 2666 3101 2668 3103
rect 3231 3101 3233 3103
rect 3236 3100 3238 3103
rect 3252 3101 3254 3103
rect 3268 3101 3270 3103
rect 3273 3098 3275 3103
rect 3294 3098 3296 3103
rect 3310 3101 3312 3103
rect 3326 3101 3328 3103
rect 3331 3098 3333 3103
rect 3347 3101 3349 3103
rect 3363 3101 3365 3103
rect 3368 3100 3370 3103
rect 3384 3101 3386 3103
rect 3400 3101 3402 3103
rect 3405 3098 3407 3103
rect 3426 3098 3428 3103
rect 3442 3101 3444 3103
rect 3458 3101 3460 3103
rect 3463 3098 3465 3103
rect 3479 3101 3481 3103
rect 3495 3101 3497 3103
rect 3500 3100 3502 3103
rect 3516 3101 3518 3103
rect 3532 3101 3534 3103
rect 3537 3098 3539 3103
rect 3558 3098 3560 3103
rect 3574 3101 3576 3103
rect 3590 3101 3592 3103
rect 3595 3098 3597 3103
rect 3611 3101 3613 3103
rect 2770 3055 2772 3057
rect 2775 3055 2777 3058
rect 2791 3055 2793 3057
rect 2807 3055 2809 3057
rect 2812 3055 2814 3058
rect 2833 3055 2835 3058
rect 2849 3055 2851 3058
rect 2865 3055 2867 3057
rect 2870 3055 2872 3058
rect 2886 3055 2888 3057
rect 2902 3055 2904 3057
rect 2907 3055 2909 3058
rect 2923 3055 2925 3057
rect 2939 3055 2941 3057
rect 2944 3055 2946 3058
rect 2965 3055 2967 3058
rect 2981 3055 2983 3058
rect 2997 3055 2999 3057
rect 3002 3055 3004 3058
rect 3018 3055 3020 3057
rect 3034 3055 3036 3057
rect 3039 3055 3041 3058
rect 3055 3055 3057 3057
rect 3071 3055 3073 3057
rect 3076 3055 3078 3058
rect 3097 3055 3099 3058
rect 3113 3055 3115 3058
rect 3129 3055 3131 3057
rect 3134 3055 3136 3058
rect 3150 3055 3152 3057
rect 3166 3055 3168 3057
rect 3171 3055 3173 3058
rect 3187 3055 3189 3057
rect 3203 3055 3205 3057
rect 3208 3055 3210 3058
rect 3229 3055 3231 3058
rect 3245 3055 3247 3058
rect 3261 3055 3263 3057
rect 3266 3055 3268 3058
rect 3282 3055 3284 3057
rect 3715 3055 3717 3057
rect 3720 3055 3722 3058
rect 3736 3055 3738 3057
rect 3752 3055 3754 3057
rect 3757 3055 3759 3058
rect 3778 3055 3780 3058
rect 3794 3055 3796 3058
rect 3810 3055 3812 3057
rect 3815 3055 3817 3058
rect 3831 3055 3833 3057
rect 3847 3055 3849 3057
rect 3852 3055 3854 3058
rect 3868 3055 3870 3057
rect 3884 3055 3886 3057
rect 3889 3055 3891 3058
rect 3910 3055 3912 3058
rect 3926 3055 3928 3058
rect 3942 3055 3944 3057
rect 3947 3055 3949 3058
rect 3963 3055 3965 3057
rect 3979 3055 3981 3057
rect 3984 3055 3986 3058
rect 4000 3055 4002 3057
rect 4016 3055 4018 3057
rect 4021 3055 4023 3058
rect 4042 3055 4044 3058
rect 4058 3055 4060 3058
rect 4074 3055 4076 3057
rect 4079 3055 4081 3058
rect 4095 3055 4097 3057
rect 4111 3055 4113 3057
rect 4116 3055 4118 3058
rect 4132 3055 4134 3057
rect 4148 3055 4150 3057
rect 4153 3055 4155 3058
rect 4174 3055 4176 3058
rect 4190 3055 4192 3058
rect 4206 3055 4208 3057
rect 4211 3055 4213 3058
rect 4227 3055 4229 3057
rect 2770 3042 2772 3047
rect 2775 3045 2777 3047
rect 2770 3028 2772 3038
rect 2775 3028 2777 3035
rect 2791 3028 2793 3047
rect 2807 3038 2809 3047
rect 2812 3045 2814 3047
rect 2833 3045 2835 3047
rect 2849 3044 2851 3047
rect 2807 3028 2809 3031
rect 2812 3028 2814 3030
rect 2833 3028 2835 3030
rect 2849 3028 2851 3040
rect 2865 3038 2867 3047
rect 2870 3045 2872 3047
rect 2886 3039 2888 3047
rect 2902 3042 2904 3047
rect 2907 3045 2909 3047
rect 2865 3028 2867 3031
rect 2870 3028 2872 3030
rect 2886 3028 2888 3035
rect 2902 3028 2904 3038
rect 2907 3028 2909 3035
rect 2923 3028 2925 3047
rect 2939 3038 2941 3047
rect 2944 3045 2946 3047
rect 2965 3045 2967 3047
rect 2981 3044 2983 3047
rect 2939 3028 2941 3031
rect 2944 3028 2946 3030
rect 2965 3028 2967 3030
rect 2981 3028 2983 3040
rect 2997 3038 2999 3047
rect 3002 3045 3004 3047
rect 3018 3039 3020 3047
rect 3034 3042 3036 3047
rect 3039 3045 3041 3047
rect 2997 3028 2999 3031
rect 3002 3028 3004 3030
rect 3018 3028 3020 3035
rect 3034 3028 3036 3038
rect 3039 3028 3041 3035
rect 3055 3028 3057 3047
rect 3071 3038 3073 3047
rect 3076 3045 3078 3047
rect 3097 3045 3099 3047
rect 3113 3044 3115 3047
rect 3071 3028 3073 3031
rect 3076 3028 3078 3030
rect 3097 3028 3099 3030
rect 3113 3028 3115 3040
rect 3129 3038 3131 3047
rect 3134 3045 3136 3047
rect 3150 3039 3152 3047
rect 3166 3042 3168 3047
rect 3171 3045 3173 3047
rect 3129 3028 3131 3031
rect 3134 3028 3136 3030
rect 3150 3028 3152 3035
rect 3166 3028 3168 3038
rect 3171 3028 3173 3035
rect 3187 3028 3189 3047
rect 3203 3038 3205 3047
rect 3208 3045 3210 3047
rect 3229 3045 3231 3047
rect 3245 3044 3247 3047
rect 3203 3028 3205 3031
rect 3208 3028 3210 3030
rect 3229 3028 3231 3030
rect 3245 3028 3247 3040
rect 3261 3038 3263 3047
rect 3266 3045 3268 3047
rect 3282 3039 3284 3047
rect 3715 3042 3717 3047
rect 3720 3045 3722 3047
rect 3261 3028 3263 3031
rect 3266 3028 3268 3030
rect 3282 3028 3284 3035
rect 2418 3022 2420 3024
rect 2423 3022 2425 3025
rect 2439 3022 2441 3024
rect 2455 3022 2457 3024
rect 2460 3022 2462 3025
rect 2481 3022 2483 3025
rect 2497 3022 2499 3025
rect 2513 3022 2515 3024
rect 2518 3022 2520 3025
rect 3715 3028 3717 3038
rect 3720 3028 3722 3035
rect 3736 3028 3738 3047
rect 3752 3038 3754 3047
rect 3757 3045 3759 3047
rect 3778 3045 3780 3047
rect 3794 3044 3796 3047
rect 3752 3028 3754 3031
rect 3757 3028 3759 3030
rect 3778 3028 3780 3030
rect 3794 3028 3796 3040
rect 3810 3038 3812 3047
rect 3815 3045 3817 3047
rect 3831 3039 3833 3047
rect 3847 3042 3849 3047
rect 3852 3045 3854 3047
rect 3810 3028 3812 3031
rect 3815 3028 3817 3030
rect 3831 3028 3833 3035
rect 3847 3028 3849 3038
rect 3852 3028 3854 3035
rect 3868 3028 3870 3047
rect 3884 3038 3886 3047
rect 3889 3045 3891 3047
rect 3910 3045 3912 3047
rect 3926 3044 3928 3047
rect 3884 3028 3886 3031
rect 3889 3028 3891 3030
rect 3910 3028 3912 3030
rect 3926 3028 3928 3040
rect 3942 3038 3944 3047
rect 3947 3045 3949 3047
rect 3963 3039 3965 3047
rect 3979 3042 3981 3047
rect 3984 3045 3986 3047
rect 3942 3028 3944 3031
rect 3947 3028 3949 3030
rect 3963 3028 3965 3035
rect 3979 3028 3981 3038
rect 3984 3028 3986 3035
rect 4000 3028 4002 3047
rect 4016 3038 4018 3047
rect 4021 3045 4023 3047
rect 4042 3045 4044 3047
rect 4058 3044 4060 3047
rect 4016 3028 4018 3031
rect 4021 3028 4023 3030
rect 4042 3028 4044 3030
rect 4058 3028 4060 3040
rect 4074 3038 4076 3047
rect 4079 3045 4081 3047
rect 4095 3039 4097 3047
rect 4111 3042 4113 3047
rect 4116 3045 4118 3047
rect 4074 3028 4076 3031
rect 4079 3028 4081 3030
rect 4095 3028 4097 3035
rect 4111 3028 4113 3038
rect 4116 3028 4118 3035
rect 4132 3028 4134 3047
rect 4148 3038 4150 3047
rect 4153 3045 4155 3047
rect 4174 3045 4176 3047
rect 4190 3044 4192 3047
rect 4148 3028 4150 3031
rect 4153 3028 4155 3030
rect 4174 3028 4176 3030
rect 4190 3028 4192 3040
rect 4206 3038 4208 3047
rect 4211 3045 4213 3047
rect 4227 3039 4229 3047
rect 4206 3028 4208 3031
rect 4211 3028 4213 3030
rect 4227 3028 4229 3035
rect 2534 3022 2536 3024
rect 2770 3022 2772 3024
rect 2775 3021 2777 3024
rect 2791 3022 2793 3024
rect 2807 3022 2809 3024
rect 2812 3019 2814 3024
rect 2833 3019 2835 3024
rect 2849 3022 2851 3024
rect 2865 3022 2867 3024
rect 2870 3019 2872 3024
rect 2886 3022 2888 3024
rect 2902 3022 2904 3024
rect 2907 3021 2909 3024
rect 2923 3022 2925 3024
rect 2939 3022 2941 3024
rect 2944 3019 2946 3024
rect 2965 3019 2967 3024
rect 2981 3022 2983 3024
rect 2997 3022 2999 3024
rect 3002 3019 3004 3024
rect 3018 3022 3020 3024
rect 3034 3022 3036 3024
rect 3039 3021 3041 3024
rect 3055 3022 3057 3024
rect 3071 3022 3073 3024
rect 3076 3019 3078 3024
rect 3097 3019 3099 3024
rect 3113 3022 3115 3024
rect 3129 3022 3131 3024
rect 3134 3019 3136 3024
rect 3150 3022 3152 3024
rect 3166 3022 3168 3024
rect 3171 3021 3173 3024
rect 3187 3022 3189 3024
rect 3203 3022 3205 3024
rect 3208 3019 3210 3024
rect 3229 3019 3231 3024
rect 3245 3022 3247 3024
rect 3261 3022 3263 3024
rect 3266 3019 3268 3024
rect 3282 3022 3284 3024
rect 3363 3022 3365 3024
rect 3368 3022 3370 3025
rect 3384 3022 3386 3024
rect 3400 3022 3402 3024
rect 3405 3022 3407 3025
rect 3426 3022 3428 3025
rect 3442 3022 3444 3025
rect 3458 3022 3460 3024
rect 3463 3022 3465 3025
rect 3479 3022 3481 3024
rect 3715 3022 3717 3024
rect 3720 3021 3722 3024
rect 3736 3022 3738 3024
rect 3752 3022 3754 3024
rect 3757 3019 3759 3024
rect 3778 3019 3780 3024
rect 3794 3022 3796 3024
rect 3810 3022 3812 3024
rect 3815 3019 3817 3024
rect 3831 3022 3833 3024
rect 3847 3022 3849 3024
rect 3852 3021 3854 3024
rect 3868 3022 3870 3024
rect 3884 3022 3886 3024
rect 3889 3019 3891 3024
rect 3910 3019 3912 3024
rect 3926 3022 3928 3024
rect 3942 3022 3944 3024
rect 3947 3019 3949 3024
rect 3963 3022 3965 3024
rect 3979 3022 3981 3024
rect 3984 3021 3986 3024
rect 4000 3022 4002 3024
rect 4016 3022 4018 3024
rect 4021 3019 4023 3024
rect 4042 3019 4044 3024
rect 4058 3022 4060 3024
rect 4074 3022 4076 3024
rect 4079 3019 4081 3024
rect 4095 3022 4097 3024
rect 4111 3022 4113 3024
rect 4116 3021 4118 3024
rect 4132 3022 4134 3024
rect 4148 3022 4150 3024
rect 4153 3019 4155 3024
rect 4174 3019 4176 3024
rect 4190 3022 4192 3024
rect 4206 3022 4208 3024
rect 4211 3019 4213 3024
rect 4227 3022 4229 3024
rect 2418 3009 2420 3014
rect 2423 3012 2425 3014
rect 2418 2995 2420 3005
rect 2423 2995 2425 3002
rect 2439 2995 2441 3014
rect 2455 3005 2457 3014
rect 2460 3012 2462 3014
rect 2481 3012 2483 3014
rect 2497 3011 2499 3014
rect 2455 2995 2457 2998
rect 2460 2995 2462 2997
rect 2481 2995 2483 2997
rect 2497 2995 2499 3007
rect 2513 3005 2515 3014
rect 2518 3012 2520 3014
rect 2513 2995 2515 2998
rect 2518 2995 2520 2997
rect 2534 2995 2536 3014
rect 3363 3009 3365 3014
rect 3368 3012 3370 3014
rect 3363 2995 3365 3005
rect 3368 2995 3370 3002
rect 3384 2995 3386 3014
rect 3400 3005 3402 3014
rect 3405 3012 3407 3014
rect 3426 3012 3428 3014
rect 3442 3011 3444 3014
rect 3400 2995 3402 2998
rect 3405 2995 3407 2997
rect 3426 2995 3428 2997
rect 3442 2995 3444 3007
rect 3458 3005 3460 3014
rect 3463 3012 3465 3014
rect 3458 2995 3460 2998
rect 3463 2995 3465 2997
rect 3479 2995 3481 3014
rect 2418 2989 2420 2991
rect 2423 2988 2425 2991
rect 2439 2989 2441 2991
rect 2455 2989 2457 2991
rect 2460 2986 2462 2991
rect 2481 2986 2483 2991
rect 2497 2989 2499 2991
rect 2513 2989 2515 2991
rect 2518 2986 2520 2991
rect 2534 2989 2536 2991
rect 3363 2989 3365 2991
rect 3368 2988 3370 2991
rect 3384 2989 3386 2991
rect 3400 2989 3402 2991
rect 2949 2984 2951 2986
rect 2791 2978 2793 2981
rect 2835 2978 2837 2981
rect 2861 2978 2863 2981
rect 2907 2978 2909 2981
rect 2861 2974 2862 2978
rect 2975 2978 2977 2982
rect 3003 2984 3005 2986
rect 3030 2984 3032 2986
rect 2980 2978 2982 2981
rect 2775 2971 2777 2973
rect 2791 2971 2793 2974
rect 2807 2971 2809 2973
rect 2830 2971 2832 2973
rect 2835 2971 2837 2974
rect 2861 2971 2863 2974
rect 2882 2971 2884 2974
rect 2902 2971 2904 2973
rect 2907 2971 2909 2974
rect 2925 2971 2927 2973
rect 2542 2958 2544 2961
rect 2542 2952 2544 2954
rect 2425 2949 2427 2952
rect 2775 2949 2777 2963
rect 2791 2961 2793 2963
rect 2791 2949 2793 2951
rect 2807 2949 2809 2963
rect 2830 2958 2832 2963
rect 2835 2961 2837 2963
rect 2861 2961 2863 2963
rect 2826 2954 2832 2958
rect 2830 2949 2832 2954
rect 2835 2949 2837 2951
rect 2861 2949 2863 2951
rect 2882 2949 2884 2963
rect 2902 2958 2904 2963
rect 2907 2961 2909 2963
rect 2898 2954 2904 2958
rect 2902 2949 2904 2954
rect 2907 2949 2909 2951
rect 2925 2949 2927 2963
rect 2949 2962 2951 2976
rect 3056 2978 3058 2982
rect 3084 2984 3086 2986
rect 3405 2986 3407 2991
rect 3426 2986 3428 2991
rect 3442 2989 3444 2991
rect 3458 2989 3460 2991
rect 3463 2986 3465 2991
rect 3479 2989 3481 2991
rect 3061 2978 3063 2981
rect 2975 2967 2977 2970
rect 2980 2968 2982 2970
rect 2976 2963 2977 2967
rect 2975 2958 2977 2963
rect 2980 2958 2982 2960
rect 2949 2956 2951 2958
rect 3003 2954 3005 2976
rect 3030 2962 3032 2976
rect 3894 2984 3896 2986
rect 3056 2967 3058 2970
rect 3061 2968 3063 2970
rect 3057 2963 3058 2967
rect 3056 2958 3058 2963
rect 3061 2958 3063 2960
rect 3030 2956 3032 2958
rect 3084 2954 3086 2976
rect 3736 2978 3738 2981
rect 3780 2978 3782 2981
rect 3806 2978 3808 2981
rect 3852 2978 3854 2981
rect 3806 2974 3807 2978
rect 3920 2978 3922 2982
rect 3948 2984 3950 2986
rect 3975 2984 3977 2986
rect 3925 2978 3927 2981
rect 3720 2971 3722 2973
rect 3736 2971 3738 2974
rect 3752 2971 3754 2973
rect 3775 2971 3777 2973
rect 3780 2971 3782 2974
rect 3806 2971 3808 2974
rect 3827 2971 3829 2974
rect 3847 2971 3849 2973
rect 3852 2971 3854 2974
rect 3870 2971 3872 2973
rect 3487 2958 3489 2961
rect 2975 2952 2977 2954
rect 2980 2949 2982 2954
rect 3056 2952 3058 2954
rect 3003 2948 3005 2950
rect 3061 2949 3063 2954
rect 3487 2952 3489 2954
rect 3084 2948 3086 2950
rect 3370 2949 3372 2952
rect 3720 2949 3722 2963
rect 3736 2961 3738 2963
rect 3736 2949 3738 2951
rect 3752 2949 3754 2963
rect 3775 2958 3777 2963
rect 3780 2961 3782 2963
rect 3806 2961 3808 2963
rect 3771 2954 3777 2958
rect 3775 2949 3777 2954
rect 3780 2949 3782 2951
rect 3806 2949 3808 2951
rect 3827 2949 3829 2963
rect 3847 2958 3849 2963
rect 3852 2961 3854 2963
rect 3843 2954 3849 2958
rect 3847 2949 3849 2954
rect 3852 2949 3854 2951
rect 3870 2949 3872 2963
rect 3894 2962 3896 2976
rect 4001 2978 4003 2982
rect 4029 2984 4031 2986
rect 4006 2978 4008 2981
rect 3920 2967 3922 2970
rect 3925 2968 3927 2970
rect 3921 2963 3922 2967
rect 3920 2958 3922 2963
rect 3925 2958 3927 2960
rect 3894 2956 3896 2958
rect 3948 2954 3950 2976
rect 3975 2962 3977 2976
rect 4001 2967 4003 2970
rect 4006 2968 4008 2970
rect 4002 2963 4003 2967
rect 4001 2958 4003 2963
rect 4006 2958 4008 2960
rect 3975 2956 3977 2958
rect 4029 2954 4031 2976
rect 3920 2952 3922 2954
rect 3925 2949 3927 2954
rect 4001 2952 4003 2954
rect 3948 2948 3950 2950
rect 4006 2949 4008 2954
rect 4029 2948 4031 2950
rect 2425 2943 2427 2945
rect 2775 2943 2777 2945
rect 2791 2941 2793 2945
rect 2807 2943 2809 2945
rect 2830 2943 2832 2945
rect 2792 2937 2793 2941
rect 2835 2940 2837 2945
rect 2861 2941 2863 2945
rect 2882 2943 2884 2945
rect 2902 2943 2904 2945
rect 2791 2934 2793 2937
rect 2836 2936 2837 2940
rect 2862 2937 2863 2941
rect 2907 2940 2909 2945
rect 2925 2943 2927 2945
rect 3370 2943 3372 2945
rect 3720 2943 3722 2945
rect 3736 2941 3738 2945
rect 3752 2943 3754 2945
rect 3775 2943 3777 2945
rect 2835 2934 2837 2936
rect 2861 2933 2863 2937
rect 2908 2936 2909 2940
rect 3737 2937 3738 2941
rect 3780 2940 3782 2945
rect 3806 2941 3808 2945
rect 3827 2943 3829 2945
rect 3847 2943 3849 2945
rect 2907 2934 2909 2936
rect 3736 2934 3738 2937
rect 3781 2936 3782 2940
rect 3807 2937 3808 2941
rect 3852 2940 3854 2945
rect 3870 2943 3872 2945
rect 3780 2934 3782 2936
rect 3806 2933 3808 2937
rect 3853 2936 3854 2940
rect 3852 2934 3854 2936
rect 2409 2920 2411 2922
rect 2425 2920 2427 2923
rect 2430 2920 2432 2922
rect 2446 2920 2448 2923
rect 2462 2920 2464 2923
rect 2483 2920 2485 2923
rect 2488 2920 2490 2922
rect 2504 2920 2506 2922
rect 2520 2920 2522 2923
rect 2525 2920 2527 2922
rect 3354 2920 3356 2922
rect 3370 2920 3372 2923
rect 3375 2920 3377 2922
rect 3391 2920 3393 2923
rect 3407 2920 3409 2923
rect 3428 2920 3430 2923
rect 3433 2920 3435 2922
rect 3449 2920 3451 2922
rect 3465 2920 3467 2923
rect 3470 2920 3472 2922
rect 2409 2893 2411 2912
rect 2425 2910 2427 2912
rect 2430 2903 2432 2912
rect 2446 2909 2448 2912
rect 2462 2910 2464 2912
rect 2483 2910 2485 2912
rect 2425 2893 2427 2895
rect 2430 2893 2432 2896
rect 2446 2893 2448 2905
rect 2488 2903 2490 2912
rect 2462 2893 2464 2895
rect 2483 2893 2485 2895
rect 2488 2893 2490 2896
rect 2504 2893 2506 2912
rect 2520 2910 2522 2912
rect 2525 2907 2527 2912
rect 2791 2911 2793 2914
rect 2835 2912 2837 2914
rect 2792 2907 2793 2911
rect 2836 2908 2837 2912
rect 2861 2911 2863 2915
rect 2907 2912 2909 2914
rect 2775 2903 2777 2905
rect 2791 2903 2793 2907
rect 2807 2903 2809 2905
rect 2830 2903 2832 2905
rect 2835 2903 2837 2908
rect 2862 2907 2863 2911
rect 2908 2908 2909 2912
rect 2861 2903 2863 2907
rect 2882 2903 2884 2905
rect 2902 2903 2904 2905
rect 2907 2903 2909 2908
rect 2925 2903 2927 2905
rect 2520 2893 2522 2900
rect 2525 2893 2527 2903
rect 2975 2902 2977 2905
rect 2980 2902 2982 2905
rect 3056 2902 3058 2905
rect 3061 2902 3063 2905
rect 2409 2887 2411 2889
rect 2425 2884 2427 2889
rect 2430 2887 2432 2889
rect 2446 2887 2448 2889
rect 2462 2884 2464 2889
rect 2483 2884 2485 2889
rect 2488 2887 2490 2889
rect 2504 2887 2506 2889
rect 2520 2886 2522 2889
rect 2525 2887 2527 2889
rect 2775 2885 2777 2899
rect 2791 2897 2793 2899
rect 2791 2885 2793 2887
rect 2807 2885 2809 2899
rect 2830 2894 2832 2899
rect 2835 2897 2837 2899
rect 2861 2897 2863 2899
rect 2826 2890 2832 2894
rect 2830 2885 2832 2890
rect 2835 2885 2837 2887
rect 2861 2885 2863 2887
rect 2882 2885 2884 2899
rect 2902 2894 2904 2899
rect 2907 2897 2909 2899
rect 2898 2890 2904 2894
rect 2902 2885 2904 2890
rect 2907 2885 2909 2887
rect 2925 2885 2927 2899
rect 2975 2886 2977 2898
rect 2980 2896 2982 2898
rect 2980 2886 2982 2888
rect 3056 2886 3058 2898
rect 3061 2896 3063 2898
rect 3354 2893 3356 2912
rect 3370 2910 3372 2912
rect 3375 2903 3377 2912
rect 3391 2909 3393 2912
rect 3407 2910 3409 2912
rect 3428 2910 3430 2912
rect 3370 2893 3372 2895
rect 3375 2893 3377 2896
rect 3391 2893 3393 2905
rect 3433 2903 3435 2912
rect 3407 2893 3409 2895
rect 3428 2893 3430 2895
rect 3433 2893 3435 2896
rect 3449 2893 3451 2912
rect 3465 2910 3467 2912
rect 3470 2907 3472 2912
rect 3736 2911 3738 2914
rect 3780 2912 3782 2914
rect 3737 2907 3738 2911
rect 3781 2908 3782 2912
rect 3806 2911 3808 2915
rect 3852 2912 3854 2914
rect 3720 2903 3722 2905
rect 3736 2903 3738 2907
rect 3752 2903 3754 2905
rect 3775 2903 3777 2905
rect 3780 2903 3782 2908
rect 3807 2907 3808 2911
rect 3853 2908 3854 2912
rect 3806 2903 3808 2907
rect 3827 2903 3829 2905
rect 3847 2903 3849 2905
rect 3852 2903 3854 2908
rect 3870 2903 3872 2905
rect 3465 2893 3467 2900
rect 3470 2893 3472 2903
rect 3920 2902 3922 2905
rect 3925 2902 3927 2905
rect 4001 2902 4003 2905
rect 4006 2902 4008 2905
rect 3061 2886 3063 2888
rect 3354 2887 3356 2889
rect 3370 2884 3372 2889
rect 3375 2887 3377 2889
rect 3391 2887 3393 2889
rect 3407 2884 3409 2889
rect 3428 2884 3430 2889
rect 3433 2887 3435 2889
rect 3449 2887 3451 2889
rect 3465 2886 3467 2889
rect 3470 2887 3472 2889
rect 3720 2885 3722 2899
rect 3736 2897 3738 2899
rect 3736 2885 3738 2887
rect 3752 2885 3754 2899
rect 3775 2894 3777 2899
rect 3780 2897 3782 2899
rect 3806 2897 3808 2899
rect 3771 2890 3777 2894
rect 3775 2885 3777 2890
rect 3780 2885 3782 2887
rect 3806 2885 3808 2887
rect 3827 2885 3829 2899
rect 3847 2894 3849 2899
rect 3852 2897 3854 2899
rect 3843 2890 3849 2894
rect 3847 2885 3849 2890
rect 3852 2885 3854 2887
rect 3870 2885 3872 2899
rect 3920 2886 3922 2898
rect 3925 2896 3927 2898
rect 3925 2886 3927 2888
rect 4001 2886 4003 2898
rect 4006 2896 4008 2898
rect 4006 2886 4008 2888
rect 2775 2875 2777 2877
rect 2791 2874 2793 2877
rect 2807 2875 2809 2877
rect 2830 2875 2832 2877
rect 2835 2874 2837 2877
rect 2861 2874 2863 2877
rect 2882 2874 2884 2877
rect 2902 2875 2904 2877
rect 2907 2874 2909 2877
rect 2925 2875 2927 2877
rect 2975 2876 2977 2878
rect 2861 2870 2862 2874
rect 2980 2873 2982 2878
rect 3056 2876 3058 2878
rect 3061 2873 3063 2878
rect 3720 2875 3722 2877
rect 3736 2874 3738 2877
rect 3752 2875 3754 2877
rect 3775 2875 3777 2877
rect 3780 2874 3782 2877
rect 3806 2874 3808 2877
rect 3827 2874 3829 2877
rect 3847 2875 3849 2877
rect 3852 2874 3854 2877
rect 3870 2875 3872 2877
rect 3920 2876 3922 2878
rect 2791 2867 2793 2870
rect 2835 2867 2837 2870
rect 2861 2867 2863 2870
rect 2907 2867 2909 2870
rect 3806 2870 3807 2874
rect 3925 2873 3927 2878
rect 4001 2876 4003 2878
rect 4006 2873 4008 2878
rect 3736 2867 3738 2870
rect 3780 2867 3782 2870
rect 3806 2867 3808 2870
rect 3852 2867 3854 2870
rect 2791 2846 2793 2849
rect 2835 2846 2837 2849
rect 2861 2846 2863 2849
rect 2907 2846 2909 2849
rect 2975 2846 2977 2850
rect 3003 2852 3005 2854
rect 3054 2852 3056 2854
rect 2980 2846 2982 2849
rect 2861 2842 2862 2846
rect 2775 2839 2777 2841
rect 2791 2839 2793 2842
rect 2807 2839 2809 2841
rect 2830 2839 2832 2841
rect 2835 2839 2837 2842
rect 2861 2839 2863 2842
rect 2882 2839 2884 2842
rect 2902 2839 2904 2841
rect 2907 2839 2909 2842
rect 2925 2839 2927 2841
rect 3080 2846 3082 2850
rect 3108 2852 3110 2854
rect 3085 2846 3087 2849
rect 2975 2835 2977 2838
rect 2980 2836 2982 2838
rect 2976 2831 2977 2835
rect 2775 2817 2777 2831
rect 2791 2829 2793 2831
rect 2791 2817 2793 2819
rect 2807 2817 2809 2831
rect 2830 2826 2832 2831
rect 2835 2829 2837 2831
rect 2861 2829 2863 2831
rect 2826 2822 2832 2826
rect 2830 2817 2832 2822
rect 2835 2817 2837 2819
rect 2861 2817 2863 2819
rect 2882 2817 2884 2831
rect 2902 2826 2904 2831
rect 2907 2829 2909 2831
rect 2898 2822 2904 2826
rect 2902 2817 2904 2822
rect 2907 2817 2909 2819
rect 2925 2817 2927 2831
rect 2975 2826 2977 2831
rect 2980 2826 2982 2828
rect 3003 2822 3005 2844
rect 3054 2830 3056 2844
rect 3736 2846 3738 2849
rect 3780 2846 3782 2849
rect 3806 2846 3808 2849
rect 3852 2846 3854 2849
rect 3920 2846 3922 2850
rect 3948 2852 3950 2854
rect 3999 2852 4001 2854
rect 3925 2846 3927 2849
rect 3080 2835 3082 2838
rect 3085 2836 3087 2838
rect 3081 2831 3082 2835
rect 3080 2826 3082 2831
rect 3085 2826 3087 2828
rect 3054 2824 3056 2826
rect 3108 2822 3110 2844
rect 3806 2842 3807 2846
rect 3720 2839 3722 2841
rect 3736 2839 3738 2842
rect 3752 2839 3754 2841
rect 3775 2839 3777 2841
rect 3780 2839 3782 2842
rect 3806 2839 3808 2842
rect 3827 2839 3829 2842
rect 3847 2839 3849 2841
rect 3852 2839 3854 2842
rect 3870 2839 3872 2841
rect 4025 2846 4027 2850
rect 4053 2852 4055 2854
rect 4030 2846 4032 2849
rect 3920 2835 3922 2838
rect 3925 2836 3927 2838
rect 3921 2831 3922 2835
rect 2975 2820 2977 2822
rect 2980 2817 2982 2822
rect 3080 2820 3082 2822
rect 3003 2816 3005 2818
rect 3085 2817 3087 2822
rect 3108 2816 3110 2818
rect 3720 2817 3722 2831
rect 3736 2829 3738 2831
rect 3736 2817 3738 2819
rect 3752 2817 3754 2831
rect 3775 2826 3777 2831
rect 3780 2829 3782 2831
rect 3806 2829 3808 2831
rect 3771 2822 3777 2826
rect 3775 2817 3777 2822
rect 3780 2817 3782 2819
rect 3806 2817 3808 2819
rect 3827 2817 3829 2831
rect 3847 2826 3849 2831
rect 3852 2829 3854 2831
rect 3843 2822 3849 2826
rect 3847 2817 3849 2822
rect 3852 2817 3854 2819
rect 3870 2817 3872 2831
rect 3920 2826 3922 2831
rect 3925 2826 3927 2828
rect 3948 2822 3950 2844
rect 3999 2830 4001 2844
rect 4025 2835 4027 2838
rect 4030 2836 4032 2838
rect 4026 2831 4027 2835
rect 4025 2826 4027 2831
rect 4030 2826 4032 2828
rect 3999 2824 4001 2826
rect 4053 2822 4055 2844
rect 3920 2820 3922 2822
rect 3925 2817 3927 2822
rect 4025 2820 4027 2822
rect 3948 2816 3950 2818
rect 4030 2817 4032 2822
rect 4053 2816 4055 2818
rect 2775 2811 2777 2813
rect 2791 2809 2793 2813
rect 2807 2811 2809 2813
rect 2830 2811 2832 2813
rect 2792 2805 2793 2809
rect 2835 2808 2837 2813
rect 2861 2809 2863 2813
rect 2882 2811 2884 2813
rect 2902 2811 2904 2813
rect 2791 2802 2793 2805
rect 2836 2804 2837 2808
rect 2862 2805 2863 2809
rect 2907 2808 2909 2813
rect 2925 2811 2927 2813
rect 3720 2811 3722 2813
rect 3736 2809 3738 2813
rect 3752 2811 3754 2813
rect 3775 2811 3777 2813
rect 2835 2802 2837 2804
rect 2861 2801 2863 2805
rect 2908 2804 2909 2808
rect 3737 2805 3738 2809
rect 3780 2808 3782 2813
rect 3806 2809 3808 2813
rect 3827 2811 3829 2813
rect 3847 2811 3849 2813
rect 2907 2802 2909 2804
rect 3736 2802 3738 2805
rect 3781 2804 3782 2808
rect 3807 2805 3808 2809
rect 3852 2808 3854 2813
rect 3870 2811 3872 2813
rect 3780 2802 3782 2804
rect 3806 2801 3808 2805
rect 3853 2804 3854 2808
rect 3852 2802 3854 2804
rect 2791 2779 2793 2782
rect 2835 2780 2837 2782
rect 2792 2775 2793 2779
rect 2836 2776 2837 2780
rect 2861 2779 2863 2783
rect 2907 2780 2909 2782
rect 2775 2771 2777 2773
rect 2791 2771 2793 2775
rect 2807 2771 2809 2773
rect 2830 2771 2832 2773
rect 2835 2771 2837 2776
rect 2862 2775 2863 2779
rect 2908 2776 2909 2780
rect 3736 2779 3738 2782
rect 3780 2780 3782 2782
rect 2861 2771 2863 2775
rect 2882 2771 2884 2773
rect 2902 2771 2904 2773
rect 2907 2771 2909 2776
rect 3737 2775 3738 2779
rect 3781 2776 3782 2780
rect 3806 2779 3808 2783
rect 3852 2780 3854 2782
rect 2925 2771 2927 2773
rect 2975 2771 2977 2774
rect 2980 2771 2982 2774
rect 3080 2771 3082 2774
rect 3085 2771 3087 2774
rect 3720 2771 3722 2773
rect 3736 2771 3738 2775
rect 3752 2771 3754 2773
rect 3775 2771 3777 2773
rect 3780 2771 3782 2776
rect 3807 2775 3808 2779
rect 3853 2776 3854 2780
rect 3806 2771 3808 2775
rect 3827 2771 3829 2773
rect 3847 2771 3849 2773
rect 3852 2771 3854 2776
rect 3870 2771 3872 2773
rect 3920 2771 3922 2774
rect 3925 2771 3927 2774
rect 4025 2771 4027 2774
rect 4030 2771 4032 2774
rect 2775 2753 2777 2767
rect 2791 2765 2793 2767
rect 2791 2753 2793 2755
rect 2807 2753 2809 2767
rect 2830 2762 2832 2767
rect 2835 2765 2837 2767
rect 2861 2765 2863 2767
rect 2826 2758 2832 2762
rect 2830 2753 2832 2758
rect 2835 2753 2837 2755
rect 2861 2753 2863 2755
rect 2882 2753 2884 2767
rect 2902 2762 2904 2767
rect 2907 2765 2909 2767
rect 2898 2758 2904 2762
rect 2902 2753 2904 2758
rect 2907 2753 2909 2755
rect 2925 2753 2927 2767
rect 2975 2755 2977 2767
rect 2980 2765 2982 2767
rect 2980 2755 2982 2757
rect 3080 2755 3082 2767
rect 3085 2765 3087 2767
rect 3085 2755 3087 2757
rect 3720 2753 3722 2767
rect 3736 2765 3738 2767
rect 3736 2753 3738 2755
rect 3752 2753 3754 2767
rect 3775 2762 3777 2767
rect 3780 2765 3782 2767
rect 3806 2765 3808 2767
rect 3771 2758 3777 2762
rect 3775 2753 3777 2758
rect 3780 2753 3782 2755
rect 3806 2753 3808 2755
rect 3827 2753 3829 2767
rect 3847 2762 3849 2767
rect 3852 2765 3854 2767
rect 3843 2758 3849 2762
rect 3847 2753 3849 2758
rect 3852 2753 3854 2755
rect 3870 2753 3872 2767
rect 3920 2755 3922 2767
rect 3925 2765 3927 2767
rect 3925 2755 3927 2757
rect 4025 2755 4027 2767
rect 4030 2765 4032 2767
rect 4030 2755 4032 2757
rect 2975 2745 2977 2747
rect 2775 2743 2777 2745
rect 2791 2742 2793 2745
rect 2807 2743 2809 2745
rect 2830 2743 2832 2745
rect 2835 2742 2837 2745
rect 2861 2742 2863 2745
rect 2882 2742 2884 2745
rect 2902 2743 2904 2745
rect 2907 2742 2909 2745
rect 2925 2743 2927 2745
rect 2980 2742 2982 2747
rect 3080 2745 3082 2747
rect 3085 2742 3087 2747
rect 3920 2745 3922 2747
rect 3720 2743 3722 2745
rect 2861 2738 2862 2742
rect 3736 2742 3738 2745
rect 3752 2743 3754 2745
rect 3775 2743 3777 2745
rect 3780 2742 3782 2745
rect 3806 2742 3808 2745
rect 3827 2742 3829 2745
rect 3847 2743 3849 2745
rect 3852 2742 3854 2745
rect 3870 2743 3872 2745
rect 3925 2742 3927 2747
rect 4025 2745 4027 2747
rect 4030 2742 4032 2747
rect 3806 2738 3807 2742
rect 2791 2735 2793 2738
rect 2835 2735 2837 2738
rect 2861 2735 2863 2738
rect 2907 2735 2909 2738
rect 3736 2735 3738 2738
rect 3780 2735 3782 2738
rect 3806 2735 3808 2738
rect 3852 2735 3854 2738
rect 2791 2714 2793 2717
rect 2835 2714 2837 2717
rect 2861 2714 2863 2717
rect 2907 2714 2909 2717
rect 2975 2714 2977 2718
rect 3003 2720 3005 2722
rect 3030 2720 3032 2722
rect 2980 2714 2982 2717
rect 2861 2710 2862 2714
rect 2775 2707 2777 2709
rect 2791 2707 2793 2710
rect 2807 2707 2809 2709
rect 2830 2707 2832 2709
rect 2835 2707 2837 2710
rect 2861 2707 2863 2710
rect 2882 2707 2884 2710
rect 2902 2707 2904 2709
rect 2907 2707 2909 2710
rect 2925 2707 2927 2709
rect 3056 2714 3058 2718
rect 3084 2720 3086 2722
rect 3120 2720 3122 2722
rect 3061 2714 3063 2717
rect 2975 2703 2977 2706
rect 2980 2704 2982 2706
rect 2976 2699 2977 2703
rect 2775 2685 2777 2699
rect 2791 2697 2793 2699
rect 2791 2685 2793 2687
rect 2807 2685 2809 2699
rect 2830 2694 2832 2699
rect 2835 2697 2837 2699
rect 2861 2697 2863 2699
rect 2826 2690 2832 2694
rect 2830 2685 2832 2690
rect 2835 2685 2837 2687
rect 2861 2685 2863 2687
rect 2882 2685 2884 2699
rect 2902 2694 2904 2699
rect 2907 2697 2909 2699
rect 2898 2690 2904 2694
rect 2902 2685 2904 2690
rect 2907 2685 2909 2687
rect 2925 2685 2927 2699
rect 2975 2694 2977 2699
rect 2980 2694 2982 2696
rect 3003 2690 3005 2712
rect 3030 2698 3032 2712
rect 3146 2714 3148 2718
rect 3174 2720 3176 2722
rect 3151 2714 3153 2717
rect 3056 2703 3058 2706
rect 3061 2704 3063 2706
rect 3057 2699 3058 2703
rect 3056 2694 3058 2699
rect 3061 2694 3063 2696
rect 3030 2692 3032 2694
rect 3084 2690 3086 2712
rect 3120 2698 3122 2712
rect 3736 2714 3738 2717
rect 3780 2714 3782 2717
rect 3806 2714 3808 2717
rect 3852 2714 3854 2717
rect 3920 2714 3922 2718
rect 3948 2720 3950 2722
rect 3975 2720 3977 2722
rect 3925 2714 3927 2717
rect 3146 2703 3148 2706
rect 3151 2704 3153 2706
rect 3147 2699 3148 2703
rect 3146 2694 3148 2699
rect 3151 2694 3153 2696
rect 3120 2692 3122 2694
rect 3174 2690 3176 2712
rect 3806 2710 3807 2714
rect 3720 2707 3722 2709
rect 3736 2707 3738 2710
rect 3752 2707 3754 2709
rect 3775 2707 3777 2709
rect 3780 2707 3782 2710
rect 3806 2707 3808 2710
rect 3827 2707 3829 2710
rect 3847 2707 3849 2709
rect 3852 2707 3854 2710
rect 3870 2707 3872 2709
rect 4001 2714 4003 2718
rect 4029 2720 4031 2722
rect 4065 2720 4067 2722
rect 4006 2714 4008 2717
rect 3920 2703 3922 2706
rect 3925 2704 3927 2706
rect 3921 2699 3922 2703
rect 2975 2688 2977 2690
rect 2980 2685 2982 2690
rect 3056 2688 3058 2690
rect 3003 2684 3005 2686
rect 3061 2685 3063 2690
rect 3146 2688 3148 2690
rect 3084 2684 3086 2686
rect 3151 2685 3153 2690
rect 3174 2684 3176 2686
rect 3720 2685 3722 2699
rect 3736 2697 3738 2699
rect 3736 2685 3738 2687
rect 3752 2685 3754 2699
rect 3775 2694 3777 2699
rect 3780 2697 3782 2699
rect 3806 2697 3808 2699
rect 3771 2690 3777 2694
rect 3775 2685 3777 2690
rect 3780 2685 3782 2687
rect 3806 2685 3808 2687
rect 3827 2685 3829 2699
rect 3847 2694 3849 2699
rect 3852 2697 3854 2699
rect 3843 2690 3849 2694
rect 3847 2685 3849 2690
rect 3852 2685 3854 2687
rect 3870 2685 3872 2699
rect 3920 2694 3922 2699
rect 3925 2694 3927 2696
rect 3948 2690 3950 2712
rect 3975 2698 3977 2712
rect 4091 2714 4093 2718
rect 4119 2720 4121 2722
rect 4096 2714 4098 2717
rect 4001 2703 4003 2706
rect 4006 2704 4008 2706
rect 4002 2699 4003 2703
rect 4001 2694 4003 2699
rect 4006 2694 4008 2696
rect 3975 2692 3977 2694
rect 4029 2690 4031 2712
rect 4065 2698 4067 2712
rect 4091 2703 4093 2706
rect 4096 2704 4098 2706
rect 4092 2699 4093 2703
rect 4091 2694 4093 2699
rect 4096 2694 4098 2696
rect 4065 2692 4067 2694
rect 4119 2690 4121 2712
rect 3920 2688 3922 2690
rect 3925 2685 3927 2690
rect 4001 2688 4003 2690
rect 3948 2684 3950 2686
rect 4006 2685 4008 2690
rect 4091 2688 4093 2690
rect 4029 2684 4031 2686
rect 4096 2685 4098 2690
rect 4119 2684 4121 2686
rect 2775 2679 2777 2681
rect 2791 2677 2793 2681
rect 2807 2679 2809 2681
rect 2830 2679 2832 2681
rect 2792 2673 2793 2677
rect 2835 2676 2837 2681
rect 2861 2677 2863 2681
rect 2882 2679 2884 2681
rect 2902 2679 2904 2681
rect 2791 2670 2793 2673
rect 2836 2672 2837 2676
rect 2862 2673 2863 2677
rect 2907 2676 2909 2681
rect 2925 2679 2927 2681
rect 3720 2679 3722 2681
rect 3736 2677 3738 2681
rect 3752 2679 3754 2681
rect 3775 2679 3777 2681
rect 2835 2670 2837 2672
rect 2861 2669 2863 2673
rect 2908 2672 2909 2676
rect 3737 2673 3738 2677
rect 3780 2676 3782 2681
rect 3806 2677 3808 2681
rect 3827 2679 3829 2681
rect 3847 2679 3849 2681
rect 2907 2670 2909 2672
rect 3736 2670 3738 2673
rect 3781 2672 3782 2676
rect 3807 2673 3808 2677
rect 3852 2676 3854 2681
rect 3870 2679 3872 2681
rect 3780 2670 3782 2672
rect 3806 2669 3808 2673
rect 3853 2672 3854 2676
rect 3852 2670 3854 2672
rect 2791 2647 2793 2650
rect 2835 2648 2837 2650
rect 2792 2643 2793 2647
rect 2836 2644 2837 2648
rect 2861 2647 2863 2651
rect 2907 2648 2909 2650
rect 2775 2639 2777 2641
rect 2791 2639 2793 2643
rect 2807 2639 2809 2641
rect 2830 2639 2832 2641
rect 2835 2639 2837 2644
rect 2862 2643 2863 2647
rect 2908 2644 2909 2648
rect 3736 2647 3738 2650
rect 3780 2648 3782 2650
rect 2861 2639 2863 2643
rect 2882 2639 2884 2641
rect 2902 2639 2904 2641
rect 2907 2639 2909 2644
rect 3737 2643 3738 2647
rect 3781 2644 3782 2648
rect 3806 2647 3808 2651
rect 3852 2648 3854 2650
rect 2925 2639 2927 2641
rect 3720 2639 3722 2641
rect 3736 2639 3738 2643
rect 3752 2639 3754 2641
rect 3775 2639 3777 2641
rect 3780 2639 3782 2644
rect 3807 2643 3808 2647
rect 3853 2644 3854 2648
rect 3806 2639 3808 2643
rect 3827 2639 3829 2641
rect 3847 2639 3849 2641
rect 3852 2639 3854 2644
rect 3870 2639 3872 2641
rect 2975 2636 2977 2639
rect 2980 2636 2982 2639
rect 3056 2636 3058 2639
rect 3061 2636 3063 2639
rect 3146 2636 3148 2639
rect 3151 2636 3153 2639
rect 2775 2621 2777 2635
rect 2791 2633 2793 2635
rect 2791 2621 2793 2623
rect 2807 2621 2809 2635
rect 2830 2630 2832 2635
rect 2835 2633 2837 2635
rect 2861 2633 2863 2635
rect 2826 2626 2832 2630
rect 2830 2621 2832 2626
rect 2835 2621 2837 2623
rect 2861 2621 2863 2623
rect 2882 2621 2884 2635
rect 2902 2630 2904 2635
rect 2907 2633 2909 2635
rect 2898 2626 2904 2630
rect 2902 2621 2904 2626
rect 2907 2621 2909 2623
rect 2925 2621 2927 2635
rect 3920 2636 3922 2639
rect 3925 2636 3927 2639
rect 4001 2636 4003 2639
rect 4006 2636 4008 2639
rect 4091 2636 4093 2639
rect 4096 2636 4098 2639
rect 2975 2620 2977 2632
rect 2980 2630 2982 2632
rect 2980 2620 2982 2622
rect 3056 2620 3058 2632
rect 3061 2630 3063 2632
rect 3061 2620 3063 2622
rect 3146 2620 3148 2632
rect 3151 2630 3153 2632
rect 3151 2620 3153 2622
rect 3720 2621 3722 2635
rect 3736 2633 3738 2635
rect 3736 2621 3738 2623
rect 3752 2621 3754 2635
rect 3775 2630 3777 2635
rect 3780 2633 3782 2635
rect 3806 2633 3808 2635
rect 3771 2626 3777 2630
rect 3775 2621 3777 2626
rect 3780 2621 3782 2623
rect 3806 2621 3808 2623
rect 3827 2621 3829 2635
rect 3847 2630 3849 2635
rect 3852 2633 3854 2635
rect 3843 2626 3849 2630
rect 3847 2621 3849 2626
rect 3852 2621 3854 2623
rect 3870 2621 3872 2635
rect 2775 2611 2777 2613
rect 2791 2610 2793 2613
rect 2807 2611 2809 2613
rect 2830 2611 2832 2613
rect 2835 2610 2837 2613
rect 2861 2610 2863 2613
rect 2882 2610 2884 2613
rect 2902 2611 2904 2613
rect 2907 2610 2909 2613
rect 2925 2611 2927 2613
rect 3920 2620 3922 2632
rect 3925 2630 3927 2632
rect 3925 2620 3927 2622
rect 4001 2620 4003 2632
rect 4006 2630 4008 2632
rect 4006 2620 4008 2622
rect 4091 2620 4093 2632
rect 4096 2630 4098 2632
rect 4096 2620 4098 2622
rect 2975 2610 2977 2612
rect 2861 2606 2862 2610
rect 2980 2607 2982 2612
rect 3056 2610 3058 2612
rect 3061 2607 3063 2612
rect 3146 2610 3148 2612
rect 3151 2607 3153 2612
rect 3720 2611 3722 2613
rect 2791 2603 2793 2606
rect 2835 2603 2837 2606
rect 2861 2603 2863 2606
rect 2907 2603 2909 2606
rect 3736 2610 3738 2613
rect 3752 2611 3754 2613
rect 3775 2611 3777 2613
rect 3780 2610 3782 2613
rect 3806 2610 3808 2613
rect 3827 2610 3829 2613
rect 3847 2611 3849 2613
rect 3852 2610 3854 2613
rect 3870 2611 3872 2613
rect 3920 2610 3922 2612
rect 3806 2606 3807 2610
rect 3925 2607 3927 2612
rect 4001 2610 4003 2612
rect 4006 2607 4008 2612
rect 4091 2610 4093 2612
rect 4096 2607 4098 2612
rect 3736 2603 3738 2606
rect 3780 2603 3782 2606
rect 3806 2603 3808 2606
rect 3852 2603 3854 2606
rect 2791 2582 2793 2585
rect 2835 2582 2837 2585
rect 2861 2582 2863 2585
rect 2907 2582 2909 2585
rect 2975 2582 2977 2586
rect 3003 2588 3005 2590
rect 2980 2582 2982 2585
rect 2861 2578 2862 2582
rect 2775 2575 2777 2577
rect 2791 2575 2793 2578
rect 2807 2575 2809 2577
rect 2830 2575 2832 2577
rect 2835 2575 2837 2578
rect 2861 2575 2863 2578
rect 2882 2575 2884 2578
rect 2902 2575 2904 2577
rect 2907 2575 2909 2578
rect 2925 2575 2927 2577
rect 3736 2582 3738 2585
rect 3780 2582 3782 2585
rect 3806 2582 3808 2585
rect 3852 2582 3854 2585
rect 3920 2582 3922 2586
rect 3948 2588 3950 2590
rect 3925 2582 3927 2585
rect 2975 2571 2977 2574
rect 2980 2572 2982 2574
rect 2976 2567 2977 2571
rect 2775 2553 2777 2567
rect 2791 2565 2793 2567
rect 2791 2553 2793 2555
rect 2807 2553 2809 2567
rect 2830 2562 2832 2567
rect 2835 2565 2837 2567
rect 2861 2565 2863 2567
rect 2826 2558 2832 2562
rect 2830 2553 2832 2558
rect 2835 2553 2837 2555
rect 2861 2553 2863 2555
rect 2882 2553 2884 2567
rect 2902 2562 2904 2567
rect 2907 2565 2909 2567
rect 2898 2558 2904 2562
rect 2902 2553 2904 2558
rect 2907 2553 2909 2555
rect 2925 2553 2927 2567
rect 2975 2562 2977 2567
rect 2980 2562 2982 2564
rect 3003 2558 3005 2580
rect 3806 2578 3807 2582
rect 3720 2575 3722 2577
rect 3736 2575 3738 2578
rect 3752 2575 3754 2577
rect 3775 2575 3777 2577
rect 3780 2575 3782 2578
rect 3806 2575 3808 2578
rect 3827 2575 3829 2578
rect 3847 2575 3849 2577
rect 3852 2575 3854 2578
rect 3870 2575 3872 2577
rect 3920 2571 3922 2574
rect 3925 2572 3927 2574
rect 3921 2567 3922 2571
rect 2975 2556 2977 2558
rect 2980 2553 2982 2558
rect 3003 2552 3005 2554
rect 3720 2553 3722 2567
rect 3736 2565 3738 2567
rect 3736 2553 3738 2555
rect 3752 2553 3754 2567
rect 3775 2562 3777 2567
rect 3780 2565 3782 2567
rect 3806 2565 3808 2567
rect 3771 2558 3777 2562
rect 3775 2553 3777 2558
rect 3780 2553 3782 2555
rect 3806 2553 3808 2555
rect 3827 2553 3829 2567
rect 3847 2562 3849 2567
rect 3852 2565 3854 2567
rect 3843 2558 3849 2562
rect 3847 2553 3849 2558
rect 3852 2553 3854 2555
rect 3870 2553 3872 2567
rect 3920 2562 3922 2567
rect 3925 2562 3927 2564
rect 3948 2558 3950 2580
rect 3920 2556 3922 2558
rect 3925 2553 3927 2558
rect 3948 2552 3950 2554
rect 2775 2547 2777 2549
rect 2791 2545 2793 2549
rect 2807 2547 2809 2549
rect 2830 2547 2832 2549
rect 2792 2541 2793 2545
rect 2835 2544 2837 2549
rect 2861 2545 2863 2549
rect 2882 2547 2884 2549
rect 2902 2547 2904 2549
rect 2791 2538 2793 2541
rect 2836 2540 2837 2544
rect 2862 2541 2863 2545
rect 2907 2544 2909 2549
rect 2925 2547 2927 2549
rect 3720 2547 3722 2549
rect 3736 2545 3738 2549
rect 3752 2547 3754 2549
rect 3775 2547 3777 2549
rect 2835 2538 2837 2540
rect 2861 2537 2863 2541
rect 2908 2540 2909 2544
rect 3737 2541 3738 2545
rect 3780 2544 3782 2549
rect 3806 2545 3808 2549
rect 3827 2547 3829 2549
rect 3847 2547 3849 2549
rect 2907 2538 2909 2540
rect 3736 2538 3738 2541
rect 3781 2540 3782 2544
rect 3807 2541 3808 2545
rect 3852 2544 3854 2549
rect 3870 2547 3872 2549
rect 3780 2538 3782 2540
rect 3806 2537 3808 2541
rect 3853 2540 3854 2544
rect 3852 2538 3854 2540
rect 2286 2520 2288 2522
rect 2291 2520 2293 2523
rect 2307 2520 2309 2522
rect 2323 2520 2325 2522
rect 2328 2520 2330 2523
rect 2349 2520 2351 2523
rect 2365 2520 2367 2523
rect 2381 2520 2383 2522
rect 2386 2520 2388 2523
rect 2402 2520 2404 2522
rect 2418 2520 2420 2522
rect 2423 2520 2425 2523
rect 2439 2520 2441 2522
rect 2455 2520 2457 2522
rect 2460 2520 2462 2523
rect 2481 2520 2483 2523
rect 2497 2520 2499 2523
rect 2513 2520 2515 2522
rect 2518 2520 2520 2523
rect 2534 2520 2536 2522
rect 2550 2520 2552 2522
rect 2555 2520 2557 2523
rect 2571 2520 2573 2522
rect 2587 2520 2589 2522
rect 2592 2520 2594 2523
rect 2613 2520 2615 2523
rect 2629 2520 2631 2523
rect 2645 2520 2647 2522
rect 2650 2520 2652 2523
rect 2666 2520 2668 2522
rect 3231 2520 3233 2522
rect 3236 2520 3238 2523
rect 3252 2520 3254 2522
rect 3268 2520 3270 2522
rect 3273 2520 3275 2523
rect 3294 2520 3296 2523
rect 3310 2520 3312 2523
rect 3326 2520 3328 2522
rect 3331 2520 3333 2523
rect 3347 2520 3349 2522
rect 3363 2520 3365 2522
rect 3368 2520 3370 2523
rect 3384 2520 3386 2522
rect 3400 2520 3402 2522
rect 3405 2520 3407 2523
rect 3426 2520 3428 2523
rect 3442 2520 3444 2523
rect 3458 2520 3460 2522
rect 3463 2520 3465 2523
rect 3479 2520 3481 2522
rect 3495 2520 3497 2522
rect 3500 2520 3502 2523
rect 3516 2520 3518 2522
rect 3532 2520 3534 2522
rect 3537 2520 3539 2523
rect 3558 2520 3560 2523
rect 3574 2520 3576 2523
rect 3590 2520 3592 2522
rect 3595 2520 3597 2523
rect 3611 2520 3613 2522
rect 2791 2515 2793 2518
rect 2835 2516 2837 2518
rect 2286 2507 2288 2512
rect 2291 2510 2293 2512
rect 2286 2493 2288 2503
rect 2291 2493 2293 2500
rect 2307 2493 2309 2512
rect 2323 2503 2325 2512
rect 2328 2510 2330 2512
rect 2349 2510 2351 2512
rect 2365 2509 2367 2512
rect 2323 2493 2325 2496
rect 2328 2493 2330 2495
rect 2349 2493 2351 2495
rect 2365 2493 2367 2505
rect 2381 2503 2383 2512
rect 2386 2510 2388 2512
rect 2381 2493 2383 2496
rect 2386 2493 2388 2495
rect 2402 2493 2404 2512
rect 2418 2509 2420 2512
rect 2423 2510 2425 2512
rect 2418 2493 2420 2505
rect 2423 2493 2425 2500
rect 2439 2493 2441 2512
rect 2455 2503 2457 2512
rect 2460 2510 2462 2512
rect 2481 2510 2483 2512
rect 2497 2509 2499 2512
rect 2455 2493 2457 2496
rect 2460 2493 2462 2495
rect 2481 2493 2483 2495
rect 2497 2493 2499 2505
rect 2513 2503 2515 2512
rect 2518 2510 2520 2512
rect 2513 2493 2515 2496
rect 2518 2493 2520 2495
rect 2534 2493 2536 2512
rect 2550 2509 2552 2512
rect 2555 2510 2557 2512
rect 2550 2493 2552 2505
rect 2555 2493 2557 2500
rect 2571 2493 2573 2512
rect 2587 2503 2589 2512
rect 2592 2510 2594 2512
rect 2613 2510 2615 2512
rect 2629 2509 2631 2512
rect 2587 2493 2589 2496
rect 2592 2493 2594 2495
rect 2613 2493 2615 2495
rect 2629 2493 2631 2505
rect 2645 2503 2647 2512
rect 2650 2510 2652 2512
rect 2666 2504 2668 2512
rect 2792 2511 2793 2515
rect 2836 2512 2837 2516
rect 2861 2515 2863 2519
rect 2907 2516 2909 2518
rect 2775 2507 2777 2509
rect 2791 2507 2793 2511
rect 2807 2507 2809 2509
rect 2830 2507 2832 2509
rect 2835 2507 2837 2512
rect 2862 2511 2863 2515
rect 2908 2512 2909 2516
rect 3052 2515 3054 2518
rect 3096 2516 3098 2518
rect 2861 2507 2863 2511
rect 2882 2507 2884 2509
rect 2902 2507 2904 2509
rect 2907 2507 2909 2512
rect 3053 2511 3054 2515
rect 3097 2512 3098 2516
rect 3122 2515 3124 2519
rect 3168 2516 3170 2518
rect 2925 2507 2927 2509
rect 3009 2507 3011 2510
rect 3027 2507 3029 2510
rect 3052 2507 3054 2511
rect 3068 2507 3070 2509
rect 3091 2507 3093 2509
rect 3096 2507 3098 2512
rect 3123 2511 3124 2515
rect 3169 2512 3170 2516
rect 3736 2515 3738 2518
rect 3780 2516 3782 2518
rect 3122 2507 3124 2511
rect 3143 2507 3145 2509
rect 3163 2507 3165 2509
rect 3168 2507 3170 2512
rect 3186 2507 3188 2509
rect 3231 2507 3233 2512
rect 3236 2510 3238 2512
rect 2645 2493 2647 2496
rect 2650 2493 2652 2495
rect 2666 2493 2668 2500
rect 2775 2489 2777 2503
rect 2791 2501 2793 2503
rect 2791 2489 2793 2491
rect 2807 2489 2809 2503
rect 2830 2498 2832 2503
rect 2835 2501 2837 2503
rect 2861 2501 2863 2503
rect 2826 2494 2832 2498
rect 2830 2489 2832 2494
rect 2835 2489 2837 2491
rect 2861 2489 2863 2491
rect 2882 2489 2884 2503
rect 2902 2498 2904 2503
rect 2907 2501 2909 2503
rect 2898 2494 2904 2498
rect 2902 2489 2904 2494
rect 2907 2489 2909 2491
rect 2925 2489 2927 2503
rect 2975 2500 2977 2503
rect 2980 2500 2982 2503
rect 3009 2498 3011 2503
rect 2286 2487 2288 2489
rect 2291 2486 2293 2489
rect 2307 2487 2309 2489
rect 2323 2487 2325 2489
rect 2328 2484 2330 2489
rect 2349 2484 2351 2489
rect 2365 2487 2367 2489
rect 2381 2487 2383 2489
rect 2386 2484 2388 2489
rect 2402 2487 2404 2489
rect 2418 2487 2420 2489
rect 2423 2486 2425 2489
rect 2439 2487 2441 2489
rect 2455 2487 2457 2489
rect 2460 2484 2462 2489
rect 2481 2484 2483 2489
rect 2497 2487 2499 2489
rect 2513 2487 2515 2489
rect 2518 2484 2520 2489
rect 2534 2487 2536 2489
rect 2550 2487 2552 2489
rect 2555 2486 2557 2489
rect 2571 2487 2573 2489
rect 2587 2487 2589 2489
rect 2592 2484 2594 2489
rect 2613 2484 2615 2489
rect 2629 2487 2631 2489
rect 2645 2487 2647 2489
rect 2650 2484 2652 2489
rect 2666 2487 2668 2489
rect 2975 2484 2977 2496
rect 2980 2494 2982 2496
rect 3009 2489 3011 2494
rect 3027 2489 3029 2503
rect 3052 2501 3054 2503
rect 3052 2489 3054 2491
rect 3068 2489 3070 2503
rect 3091 2498 3093 2503
rect 3096 2501 3098 2503
rect 3122 2501 3124 2503
rect 3087 2494 3093 2498
rect 3091 2489 3093 2494
rect 3096 2489 3098 2491
rect 3122 2489 3124 2491
rect 3143 2489 3145 2503
rect 3163 2498 3165 2503
rect 3168 2501 3170 2503
rect 3159 2494 3165 2498
rect 3163 2489 3165 2494
rect 3168 2489 3170 2491
rect 3186 2489 3188 2503
rect 3231 2493 3233 2503
rect 3236 2493 3238 2500
rect 3252 2493 3254 2512
rect 3268 2503 3270 2512
rect 3273 2510 3275 2512
rect 3294 2510 3296 2512
rect 3310 2509 3312 2512
rect 3268 2493 3270 2496
rect 3273 2493 3275 2495
rect 3294 2493 3296 2495
rect 3310 2493 3312 2505
rect 3326 2503 3328 2512
rect 3331 2510 3333 2512
rect 3326 2493 3328 2496
rect 3331 2493 3333 2495
rect 3347 2493 3349 2512
rect 3363 2509 3365 2512
rect 3368 2510 3370 2512
rect 3363 2493 3365 2505
rect 3368 2493 3370 2500
rect 3384 2493 3386 2512
rect 3400 2503 3402 2512
rect 3405 2510 3407 2512
rect 3426 2510 3428 2512
rect 3442 2509 3444 2512
rect 3400 2493 3402 2496
rect 3405 2493 3407 2495
rect 3426 2493 3428 2495
rect 3442 2493 3444 2505
rect 3458 2503 3460 2512
rect 3463 2510 3465 2512
rect 3458 2493 3460 2496
rect 3463 2493 3465 2495
rect 3479 2493 3481 2512
rect 3495 2509 3497 2512
rect 3500 2510 3502 2512
rect 3495 2493 3497 2505
rect 3500 2493 3502 2500
rect 3516 2493 3518 2512
rect 3532 2503 3534 2512
rect 3537 2510 3539 2512
rect 3558 2510 3560 2512
rect 3574 2509 3576 2512
rect 3532 2493 3534 2496
rect 3537 2493 3539 2495
rect 3558 2493 3560 2495
rect 3574 2493 3576 2505
rect 3590 2503 3592 2512
rect 3595 2510 3597 2512
rect 3611 2504 3613 2512
rect 3737 2511 3738 2515
rect 3781 2512 3782 2516
rect 3806 2515 3808 2519
rect 3852 2516 3854 2518
rect 3720 2507 3722 2509
rect 3736 2507 3738 2511
rect 3752 2507 3754 2509
rect 3775 2507 3777 2509
rect 3780 2507 3782 2512
rect 3807 2511 3808 2515
rect 3853 2512 3854 2516
rect 3997 2515 3999 2518
rect 4041 2516 4043 2518
rect 3806 2507 3808 2511
rect 3827 2507 3829 2509
rect 3847 2507 3849 2509
rect 3852 2507 3854 2512
rect 3998 2511 3999 2515
rect 4042 2512 4043 2516
rect 4067 2515 4069 2519
rect 4113 2516 4115 2518
rect 3870 2507 3872 2509
rect 3954 2507 3956 2510
rect 3972 2507 3974 2510
rect 3997 2507 3999 2511
rect 4013 2507 4015 2509
rect 4036 2507 4038 2509
rect 4041 2507 4043 2512
rect 4068 2511 4069 2515
rect 4114 2512 4115 2516
rect 4067 2507 4069 2511
rect 4088 2507 4090 2509
rect 4108 2507 4110 2509
rect 4113 2507 4115 2512
rect 4131 2507 4133 2509
rect 3590 2493 3592 2496
rect 3595 2493 3597 2495
rect 3611 2493 3613 2500
rect 3720 2489 3722 2503
rect 3736 2501 3738 2503
rect 3736 2489 3738 2491
rect 3752 2489 3754 2503
rect 3775 2498 3777 2503
rect 3780 2501 3782 2503
rect 3806 2501 3808 2503
rect 3771 2494 3777 2498
rect 3775 2489 3777 2494
rect 3780 2489 3782 2491
rect 3806 2489 3808 2491
rect 3827 2489 3829 2503
rect 3847 2498 3849 2503
rect 3852 2501 3854 2503
rect 3843 2494 3849 2498
rect 3847 2489 3849 2494
rect 3852 2489 3854 2491
rect 3870 2489 3872 2503
rect 3920 2500 3922 2503
rect 3925 2500 3927 2503
rect 3954 2498 3956 2503
rect 2980 2484 2982 2486
rect 2775 2479 2777 2481
rect 2791 2478 2793 2481
rect 2807 2479 2809 2481
rect 2830 2479 2832 2481
rect 2835 2478 2837 2481
rect 2861 2478 2863 2481
rect 2882 2478 2884 2481
rect 2902 2479 2904 2481
rect 2907 2478 2909 2481
rect 2925 2479 2927 2481
rect 2861 2474 2862 2478
rect 3231 2487 3233 2489
rect 3236 2486 3238 2489
rect 3252 2487 3254 2489
rect 3268 2487 3270 2489
rect 3273 2484 3275 2489
rect 3294 2484 3296 2489
rect 3310 2487 3312 2489
rect 3326 2487 3328 2489
rect 3331 2484 3333 2489
rect 3347 2487 3349 2489
rect 3363 2487 3365 2489
rect 3009 2478 3011 2481
rect 2975 2474 2977 2476
rect 2791 2471 2793 2474
rect 2835 2471 2837 2474
rect 2861 2471 2863 2474
rect 2907 2471 2909 2474
rect 2980 2471 2982 2476
rect 2401 2449 2403 2452
rect 2425 2449 2427 2452
rect 2401 2443 2403 2445
rect 2425 2443 2427 2445
rect 3027 2439 3029 2481
rect 3052 2478 3054 2481
rect 3068 2479 3070 2481
rect 3091 2479 3093 2481
rect 3096 2478 3098 2481
rect 3122 2478 3124 2481
rect 3143 2478 3145 2481
rect 3163 2479 3165 2481
rect 3168 2478 3170 2481
rect 3186 2479 3188 2481
rect 3368 2486 3370 2489
rect 3384 2487 3386 2489
rect 3400 2487 3402 2489
rect 3405 2484 3407 2489
rect 3426 2484 3428 2489
rect 3442 2487 3444 2489
rect 3458 2487 3460 2489
rect 3463 2484 3465 2489
rect 3479 2487 3481 2489
rect 3495 2487 3497 2489
rect 3500 2486 3502 2489
rect 3516 2487 3518 2489
rect 3532 2487 3534 2489
rect 3537 2484 3539 2489
rect 3558 2484 3560 2489
rect 3574 2487 3576 2489
rect 3590 2487 3592 2489
rect 3595 2484 3597 2489
rect 3611 2487 3613 2489
rect 3920 2484 3922 2496
rect 3925 2494 3927 2496
rect 3954 2489 3956 2494
rect 3972 2489 3974 2503
rect 3997 2501 3999 2503
rect 3997 2489 3999 2491
rect 4013 2489 4015 2503
rect 4036 2498 4038 2503
rect 4041 2501 4043 2503
rect 4067 2501 4069 2503
rect 4032 2494 4038 2498
rect 4036 2489 4038 2494
rect 4041 2489 4043 2491
rect 4067 2489 4069 2491
rect 4088 2489 4090 2503
rect 4108 2498 4110 2503
rect 4113 2501 4115 2503
rect 4104 2494 4110 2498
rect 4108 2489 4110 2494
rect 4113 2489 4115 2491
rect 4131 2489 4133 2503
rect 3925 2484 3927 2486
rect 3720 2479 3722 2481
rect 3736 2478 3738 2481
rect 3752 2479 3754 2481
rect 3775 2479 3777 2481
rect 3780 2478 3782 2481
rect 3806 2478 3808 2481
rect 3827 2478 3829 2481
rect 3847 2479 3849 2481
rect 3852 2478 3854 2481
rect 3870 2479 3872 2481
rect 3122 2474 3123 2478
rect 3052 2471 3054 2474
rect 3096 2471 3098 2474
rect 3122 2471 3124 2474
rect 3168 2471 3170 2474
rect 3806 2474 3807 2478
rect 3954 2478 3956 2481
rect 3920 2474 3922 2476
rect 3736 2471 3738 2474
rect 3780 2471 3782 2474
rect 3806 2471 3808 2474
rect 3852 2471 3854 2474
rect 3925 2471 3927 2476
rect 3346 2449 3348 2452
rect 3370 2449 3372 2452
rect 3195 2447 3198 2449
rect 3202 2447 3205 2449
rect 3346 2443 3348 2445
rect 3370 2443 3372 2445
rect 3972 2443 3974 2481
rect 3997 2478 3999 2481
rect 4013 2479 4015 2481
rect 4036 2479 4038 2481
rect 4041 2478 4043 2481
rect 4067 2478 4069 2481
rect 4088 2478 4090 2481
rect 4108 2479 4110 2481
rect 4113 2478 4115 2481
rect 4131 2479 4133 2481
rect 4067 2474 4068 2478
rect 3997 2471 3999 2474
rect 4041 2471 4043 2474
rect 4067 2471 4069 2474
rect 4113 2471 4115 2474
rect 4140 2447 4143 2449
rect 4147 2447 4150 2449
rect 2421 2436 2423 2438
rect 3366 2436 3368 2438
rect 2421 2429 2423 2432
rect 3366 2429 3368 2432
rect 2410 2418 2412 2420
rect 2416 2418 2435 2420
rect 3355 2418 3357 2420
rect 3361 2418 3380 2420
rect 2401 2413 2403 2415
rect 2425 2413 2427 2415
rect 3346 2413 3348 2415
rect 3370 2413 3372 2415
rect 2401 2406 2403 2409
rect 2425 2406 2427 2409
rect 3069 2408 3071 2410
rect 3074 2408 3076 2411
rect 3090 2408 3092 2410
rect 3106 2408 3108 2410
rect 3111 2408 3113 2411
rect 3132 2408 3134 2411
rect 3148 2408 3150 2411
rect 3164 2408 3166 2410
rect 3169 2408 3171 2411
rect 3185 2408 3187 2410
rect 3346 2406 3348 2409
rect 3370 2406 3372 2409
rect 4014 2408 4016 2410
rect 4019 2408 4021 2411
rect 4035 2408 4037 2410
rect 4051 2408 4053 2410
rect 4056 2408 4058 2411
rect 4077 2408 4079 2411
rect 4093 2408 4095 2411
rect 4109 2408 4111 2410
rect 4114 2408 4116 2411
rect 4130 2408 4132 2410
rect 3069 2395 3071 2400
rect 3074 2398 3076 2400
rect 3069 2381 3071 2391
rect 3074 2381 3076 2388
rect 3090 2381 3092 2400
rect 3106 2391 3108 2400
rect 3111 2398 3113 2400
rect 3132 2398 3134 2400
rect 3148 2397 3150 2400
rect 3106 2381 3108 2384
rect 3111 2381 3113 2383
rect 3132 2381 3134 2383
rect 3148 2381 3150 2393
rect 3164 2391 3166 2400
rect 3169 2398 3171 2400
rect 3164 2381 3166 2384
rect 3169 2381 3171 2383
rect 3185 2381 3187 2400
rect 4014 2395 4016 2400
rect 4019 2398 4021 2400
rect 4014 2381 4016 2391
rect 4019 2381 4021 2388
rect 4035 2381 4037 2400
rect 4051 2391 4053 2400
rect 4056 2398 4058 2400
rect 4077 2398 4079 2400
rect 4093 2397 4095 2400
rect 4051 2381 4053 2384
rect 4056 2381 4058 2383
rect 4077 2381 4079 2383
rect 4093 2381 4095 2393
rect 4109 2391 4111 2400
rect 4114 2398 4116 2400
rect 4109 2381 4111 2384
rect 4114 2381 4116 2383
rect 4130 2381 4132 2400
rect 2286 2378 2288 2380
rect 2291 2378 2293 2381
rect 2307 2378 2309 2380
rect 2323 2378 2325 2380
rect 2328 2378 2330 2381
rect 2349 2378 2351 2381
rect 2365 2378 2367 2381
rect 2381 2378 2383 2380
rect 2386 2378 2388 2381
rect 2402 2378 2404 2380
rect 2418 2378 2420 2380
rect 2423 2378 2425 2381
rect 2439 2378 2441 2380
rect 2455 2378 2457 2380
rect 2460 2378 2462 2381
rect 2481 2378 2483 2381
rect 2497 2378 2499 2381
rect 2513 2378 2515 2380
rect 2518 2378 2520 2381
rect 2534 2378 2536 2380
rect 2550 2378 2552 2380
rect 2555 2378 2557 2381
rect 2571 2378 2573 2380
rect 2587 2378 2589 2380
rect 2592 2378 2594 2381
rect 2613 2378 2615 2381
rect 2629 2378 2631 2381
rect 2645 2378 2647 2380
rect 2650 2378 2652 2381
rect 2666 2378 2668 2380
rect 3231 2378 3233 2380
rect 3236 2378 3238 2381
rect 3252 2378 3254 2380
rect 3268 2378 3270 2380
rect 3273 2378 3275 2381
rect 3294 2378 3296 2381
rect 3310 2378 3312 2381
rect 3326 2378 3328 2380
rect 3331 2378 3333 2381
rect 3347 2378 3349 2380
rect 3363 2378 3365 2380
rect 3368 2378 3370 2381
rect 3384 2378 3386 2380
rect 3400 2378 3402 2380
rect 3405 2378 3407 2381
rect 3426 2378 3428 2381
rect 3442 2378 3444 2381
rect 3458 2378 3460 2380
rect 3463 2378 3465 2381
rect 3479 2378 3481 2380
rect 3495 2378 3497 2380
rect 3500 2378 3502 2381
rect 3516 2378 3518 2380
rect 3532 2378 3534 2380
rect 3537 2378 3539 2381
rect 3558 2378 3560 2381
rect 3574 2378 3576 2381
rect 3590 2378 3592 2380
rect 3595 2378 3597 2381
rect 3611 2378 3613 2380
rect 3069 2375 3071 2377
rect 3074 2374 3076 2377
rect 3090 2375 3092 2377
rect 3106 2375 3108 2377
rect 3111 2372 3113 2377
rect 3132 2372 3134 2377
rect 3148 2375 3150 2377
rect 3164 2375 3166 2377
rect 3169 2372 3171 2377
rect 3185 2375 3187 2377
rect 2286 2365 2288 2370
rect 2291 2368 2293 2370
rect 2286 2351 2288 2361
rect 2291 2351 2293 2358
rect 2307 2351 2309 2370
rect 2323 2361 2325 2370
rect 2328 2368 2330 2370
rect 2349 2368 2351 2370
rect 2365 2367 2367 2370
rect 2323 2351 2325 2354
rect 2328 2351 2330 2353
rect 2349 2351 2351 2353
rect 2365 2351 2367 2363
rect 2381 2361 2383 2370
rect 2386 2368 2388 2370
rect 2381 2351 2383 2354
rect 2386 2351 2388 2353
rect 2402 2351 2404 2370
rect 2418 2367 2420 2370
rect 2423 2368 2425 2370
rect 2418 2351 2420 2363
rect 2423 2351 2425 2358
rect 2439 2351 2441 2370
rect 2455 2361 2457 2370
rect 2460 2368 2462 2370
rect 2481 2368 2483 2370
rect 2497 2367 2499 2370
rect 2455 2351 2457 2354
rect 2460 2351 2462 2353
rect 2481 2351 2483 2353
rect 2497 2351 2499 2363
rect 2513 2361 2515 2370
rect 2518 2368 2520 2370
rect 2513 2351 2515 2354
rect 2518 2351 2520 2353
rect 2534 2351 2536 2370
rect 2550 2367 2552 2370
rect 2555 2368 2557 2370
rect 2550 2351 2552 2363
rect 2555 2351 2557 2358
rect 2571 2351 2573 2370
rect 2587 2361 2589 2370
rect 2592 2368 2594 2370
rect 2613 2368 2615 2370
rect 2629 2367 2631 2370
rect 2587 2351 2589 2354
rect 2592 2351 2594 2353
rect 2613 2351 2615 2353
rect 2629 2351 2631 2363
rect 2645 2361 2647 2370
rect 2650 2368 2652 2370
rect 2666 2362 2668 2370
rect 4014 2375 4016 2377
rect 4019 2374 4021 2377
rect 4035 2375 4037 2377
rect 4051 2375 4053 2377
rect 4056 2372 4058 2377
rect 4077 2372 4079 2377
rect 4093 2375 4095 2377
rect 4109 2375 4111 2377
rect 4114 2372 4116 2377
rect 4130 2375 4132 2377
rect 3231 2365 3233 2370
rect 3236 2368 3238 2370
rect 2645 2351 2647 2354
rect 2650 2351 2652 2353
rect 2666 2351 2668 2358
rect 3231 2351 3233 2361
rect 3236 2351 3238 2358
rect 3252 2351 3254 2370
rect 3268 2361 3270 2370
rect 3273 2368 3275 2370
rect 3294 2368 3296 2370
rect 3310 2367 3312 2370
rect 3268 2351 3270 2354
rect 3273 2351 3275 2353
rect 3294 2351 3296 2353
rect 3310 2351 3312 2363
rect 3326 2361 3328 2370
rect 3331 2368 3333 2370
rect 3326 2351 3328 2354
rect 3331 2351 3333 2353
rect 3347 2351 3349 2370
rect 3363 2367 3365 2370
rect 3368 2368 3370 2370
rect 3363 2351 3365 2363
rect 3368 2351 3370 2358
rect 3384 2351 3386 2370
rect 3400 2361 3402 2370
rect 3405 2368 3407 2370
rect 3426 2368 3428 2370
rect 3442 2367 3444 2370
rect 3400 2351 3402 2354
rect 3405 2351 3407 2353
rect 3426 2351 3428 2353
rect 3442 2351 3444 2363
rect 3458 2361 3460 2370
rect 3463 2368 3465 2370
rect 3458 2351 3460 2354
rect 3463 2351 3465 2353
rect 3479 2351 3481 2370
rect 3495 2367 3497 2370
rect 3500 2368 3502 2370
rect 3495 2351 3497 2363
rect 3500 2351 3502 2358
rect 3516 2351 3518 2370
rect 3532 2361 3534 2370
rect 3537 2368 3539 2370
rect 3558 2368 3560 2370
rect 3574 2367 3576 2370
rect 3532 2351 3534 2354
rect 3537 2351 3539 2353
rect 3558 2351 3560 2353
rect 3574 2351 3576 2363
rect 3590 2361 3592 2370
rect 3595 2368 3597 2370
rect 3611 2362 3613 2370
rect 3590 2351 3592 2354
rect 3595 2351 3597 2353
rect 3611 2351 3613 2358
rect 2286 2345 2288 2347
rect 2291 2344 2293 2347
rect 2307 2345 2309 2347
rect 2323 2345 2325 2347
rect 2328 2342 2330 2347
rect 2349 2342 2351 2347
rect 2365 2345 2367 2347
rect 2381 2345 2383 2347
rect 2386 2342 2388 2347
rect 2402 2345 2404 2347
rect 2418 2345 2420 2347
rect 2423 2344 2425 2347
rect 2439 2345 2441 2347
rect 2455 2345 2457 2347
rect 2460 2342 2462 2347
rect 2481 2342 2483 2347
rect 2497 2345 2499 2347
rect 2513 2345 2515 2347
rect 2518 2342 2520 2347
rect 2534 2345 2536 2347
rect 2550 2345 2552 2347
rect 2555 2344 2557 2347
rect 2571 2345 2573 2347
rect 2587 2345 2589 2347
rect 2592 2342 2594 2347
rect 2613 2342 2615 2347
rect 2629 2345 2631 2347
rect 2645 2345 2647 2347
rect 2650 2342 2652 2347
rect 2666 2345 2668 2347
rect 3231 2345 3233 2347
rect 3236 2344 3238 2347
rect 3252 2345 3254 2347
rect 3268 2345 3270 2347
rect 3273 2342 3275 2347
rect 3294 2342 3296 2347
rect 3310 2345 3312 2347
rect 3326 2345 3328 2347
rect 3331 2342 3333 2347
rect 3347 2345 3349 2347
rect 3363 2345 3365 2347
rect 3368 2344 3370 2347
rect 3384 2345 3386 2347
rect 3400 2345 3402 2347
rect 3405 2342 3407 2347
rect 3426 2342 3428 2347
rect 3442 2345 3444 2347
rect 3458 2345 3460 2347
rect 3463 2342 3465 2347
rect 3479 2345 3481 2347
rect 3495 2345 3497 2347
rect 3500 2344 3502 2347
rect 3516 2345 3518 2347
rect 3532 2345 3534 2347
rect 3537 2342 3539 2347
rect 3558 2342 3560 2347
rect 3574 2345 3576 2347
rect 3590 2345 3592 2347
rect 3595 2342 3597 2347
rect 3611 2345 3613 2347
rect 3069 2322 3071 2324
rect 3074 2322 3076 2325
rect 3090 2322 3092 2324
rect 3106 2322 3108 2324
rect 3111 2322 3113 2325
rect 3132 2322 3134 2325
rect 3148 2322 3150 2325
rect 3164 2322 3166 2324
rect 3169 2322 3171 2325
rect 3185 2322 3187 2324
rect 4014 2322 4016 2324
rect 4019 2322 4021 2325
rect 4035 2322 4037 2324
rect 4051 2322 4053 2324
rect 4056 2322 4058 2325
rect 4077 2322 4079 2325
rect 4093 2322 4095 2325
rect 4109 2322 4111 2324
rect 4114 2322 4116 2325
rect 4130 2322 4132 2324
rect 3069 2309 3071 2314
rect 3074 2312 3076 2314
rect 3069 2295 3071 2305
rect 3074 2295 3076 2302
rect 3090 2295 3092 2314
rect 3106 2305 3108 2314
rect 3111 2312 3113 2314
rect 3132 2312 3134 2314
rect 3148 2311 3150 2314
rect 3106 2295 3108 2298
rect 3111 2295 3113 2297
rect 3132 2295 3134 2297
rect 3148 2295 3150 2307
rect 3164 2305 3166 2314
rect 3169 2312 3171 2314
rect 3164 2295 3166 2298
rect 3169 2295 3171 2297
rect 3185 2295 3187 2314
rect 4014 2309 4016 2314
rect 4019 2312 4021 2314
rect 3207 2301 3210 2303
rect 3214 2301 3217 2303
rect 4014 2295 4016 2305
rect 4019 2295 4021 2302
rect 4035 2295 4037 2314
rect 4051 2305 4053 2314
rect 4056 2312 4058 2314
rect 4077 2312 4079 2314
rect 4093 2311 4095 2314
rect 4051 2295 4053 2298
rect 4056 2295 4058 2297
rect 4077 2295 4079 2297
rect 4093 2295 4095 2307
rect 4109 2305 4111 2314
rect 4114 2312 4116 2314
rect 4109 2295 4111 2298
rect 4114 2295 4116 2297
rect 4130 2295 4132 2314
rect 4152 2301 4155 2303
rect 4159 2301 4162 2303
rect 2286 2292 2288 2294
rect 2291 2292 2293 2295
rect 2307 2292 2309 2294
rect 2323 2292 2325 2294
rect 2328 2292 2330 2295
rect 2349 2292 2351 2295
rect 2365 2292 2367 2295
rect 2381 2292 2383 2294
rect 2386 2292 2388 2295
rect 2402 2292 2404 2294
rect 2418 2292 2420 2294
rect 2423 2292 2425 2295
rect 2439 2292 2441 2294
rect 2455 2292 2457 2294
rect 2460 2292 2462 2295
rect 2481 2292 2483 2295
rect 2497 2292 2499 2295
rect 2513 2292 2515 2294
rect 2518 2292 2520 2295
rect 2534 2292 2536 2294
rect 2550 2292 2552 2294
rect 2555 2292 2557 2295
rect 2571 2292 2573 2294
rect 2587 2292 2589 2294
rect 2592 2292 2594 2295
rect 2613 2292 2615 2295
rect 2629 2292 2631 2295
rect 2645 2292 2647 2294
rect 2650 2292 2652 2295
rect 2666 2292 2668 2294
rect 3231 2292 3233 2294
rect 3236 2292 3238 2295
rect 3252 2292 3254 2294
rect 3268 2292 3270 2294
rect 3273 2292 3275 2295
rect 3294 2292 3296 2295
rect 3310 2292 3312 2295
rect 3326 2292 3328 2294
rect 3331 2292 3333 2295
rect 3347 2292 3349 2294
rect 3363 2292 3365 2294
rect 3368 2292 3370 2295
rect 3384 2292 3386 2294
rect 3400 2292 3402 2294
rect 3405 2292 3407 2295
rect 3426 2292 3428 2295
rect 3442 2292 3444 2295
rect 3458 2292 3460 2294
rect 3463 2292 3465 2295
rect 3479 2292 3481 2294
rect 3495 2292 3497 2294
rect 3500 2292 3502 2295
rect 3516 2292 3518 2294
rect 3532 2292 3534 2294
rect 3537 2292 3539 2295
rect 3558 2292 3560 2295
rect 3574 2292 3576 2295
rect 3590 2292 3592 2294
rect 3595 2292 3597 2295
rect 3611 2292 3613 2294
rect 3069 2289 3071 2291
rect 3074 2288 3076 2291
rect 3090 2289 3092 2291
rect 3106 2289 3108 2291
rect 3111 2286 3113 2291
rect 3132 2286 3134 2291
rect 3148 2289 3150 2291
rect 3164 2289 3166 2291
rect 3169 2286 3171 2291
rect 3185 2289 3187 2291
rect 2286 2279 2288 2284
rect 2291 2282 2293 2284
rect 2286 2265 2288 2275
rect 2291 2265 2293 2272
rect 2307 2265 2309 2284
rect 2323 2275 2325 2284
rect 2328 2282 2330 2284
rect 2349 2282 2351 2284
rect 2365 2281 2367 2284
rect 2323 2265 2325 2268
rect 2328 2265 2330 2267
rect 2349 2265 2351 2267
rect 2365 2265 2367 2277
rect 2381 2275 2383 2284
rect 2386 2282 2388 2284
rect 2381 2265 2383 2268
rect 2386 2265 2388 2267
rect 2402 2265 2404 2284
rect 2418 2281 2420 2284
rect 2423 2282 2425 2284
rect 2418 2265 2420 2277
rect 2423 2265 2425 2272
rect 2439 2265 2441 2284
rect 2455 2275 2457 2284
rect 2460 2282 2462 2284
rect 2481 2282 2483 2284
rect 2497 2281 2499 2284
rect 2455 2265 2457 2268
rect 2460 2265 2462 2267
rect 2481 2265 2483 2267
rect 2497 2265 2499 2277
rect 2513 2275 2515 2284
rect 2518 2282 2520 2284
rect 2513 2265 2515 2268
rect 2518 2265 2520 2267
rect 2534 2265 2536 2284
rect 2550 2281 2552 2284
rect 2555 2282 2557 2284
rect 2550 2265 2552 2277
rect 2555 2265 2557 2272
rect 2571 2265 2573 2284
rect 2587 2275 2589 2284
rect 2592 2282 2594 2284
rect 2613 2282 2615 2284
rect 2629 2281 2631 2284
rect 2587 2265 2589 2268
rect 2592 2265 2594 2267
rect 2613 2265 2615 2267
rect 2629 2265 2631 2277
rect 2645 2275 2647 2284
rect 2650 2282 2652 2284
rect 2666 2276 2668 2284
rect 4014 2289 4016 2291
rect 4019 2288 4021 2291
rect 4035 2289 4037 2291
rect 4051 2289 4053 2291
rect 4056 2286 4058 2291
rect 4077 2286 4079 2291
rect 4093 2289 4095 2291
rect 4109 2289 4111 2291
rect 4114 2286 4116 2291
rect 4130 2289 4132 2291
rect 3231 2279 3233 2284
rect 3236 2282 3238 2284
rect 2645 2265 2647 2268
rect 2650 2265 2652 2267
rect 2666 2265 2668 2272
rect 3231 2265 3233 2275
rect 3236 2265 3238 2272
rect 3252 2265 3254 2284
rect 3268 2275 3270 2284
rect 3273 2282 3275 2284
rect 3294 2282 3296 2284
rect 3310 2281 3312 2284
rect 3268 2265 3270 2268
rect 3273 2265 3275 2267
rect 3294 2265 3296 2267
rect 3310 2265 3312 2277
rect 3326 2275 3328 2284
rect 3331 2282 3333 2284
rect 3326 2265 3328 2268
rect 3331 2265 3333 2267
rect 3347 2265 3349 2284
rect 3363 2281 3365 2284
rect 3368 2282 3370 2284
rect 3363 2265 3365 2277
rect 3368 2265 3370 2272
rect 3384 2265 3386 2284
rect 3400 2275 3402 2284
rect 3405 2282 3407 2284
rect 3426 2282 3428 2284
rect 3442 2281 3444 2284
rect 3400 2265 3402 2268
rect 3405 2265 3407 2267
rect 3426 2265 3428 2267
rect 3442 2265 3444 2277
rect 3458 2275 3460 2284
rect 3463 2282 3465 2284
rect 3458 2265 3460 2268
rect 3463 2265 3465 2267
rect 3479 2265 3481 2284
rect 3495 2281 3497 2284
rect 3500 2282 3502 2284
rect 3495 2265 3497 2277
rect 3500 2265 3502 2272
rect 3516 2265 3518 2284
rect 3532 2275 3534 2284
rect 3537 2282 3539 2284
rect 3558 2282 3560 2284
rect 3574 2281 3576 2284
rect 3532 2265 3534 2268
rect 3537 2265 3539 2267
rect 3558 2265 3560 2267
rect 3574 2265 3576 2277
rect 3590 2275 3592 2284
rect 3595 2282 3597 2284
rect 3611 2276 3613 2284
rect 3590 2265 3592 2268
rect 3595 2265 3597 2267
rect 3611 2265 3613 2272
rect 2286 2259 2288 2261
rect 2291 2258 2293 2261
rect 2307 2259 2309 2261
rect 2323 2259 2325 2261
rect 2328 2256 2330 2261
rect 2349 2256 2351 2261
rect 2365 2259 2367 2261
rect 2381 2259 2383 2261
rect 2386 2256 2388 2261
rect 2402 2259 2404 2261
rect 2418 2259 2420 2261
rect 2423 2258 2425 2261
rect 2439 2259 2441 2261
rect 2455 2259 2457 2261
rect 2460 2256 2462 2261
rect 2481 2256 2483 2261
rect 2497 2259 2499 2261
rect 2513 2259 2515 2261
rect 2518 2256 2520 2261
rect 2534 2259 2536 2261
rect 2550 2259 2552 2261
rect 2555 2258 2557 2261
rect 2571 2259 2573 2261
rect 2587 2259 2589 2261
rect 2592 2256 2594 2261
rect 2613 2256 2615 2261
rect 2629 2259 2631 2261
rect 2645 2259 2647 2261
rect 2650 2256 2652 2261
rect 2666 2259 2668 2261
rect 3231 2259 3233 2261
rect 3236 2258 3238 2261
rect 3252 2259 3254 2261
rect 3268 2259 3270 2261
rect 3273 2256 3275 2261
rect 3294 2256 3296 2261
rect 3310 2259 3312 2261
rect 3326 2259 3328 2261
rect 3331 2256 3333 2261
rect 3347 2259 3349 2261
rect 3363 2259 3365 2261
rect 3368 2258 3370 2261
rect 3384 2259 3386 2261
rect 3400 2259 3402 2261
rect 3405 2256 3407 2261
rect 3426 2256 3428 2261
rect 3442 2259 3444 2261
rect 3458 2259 3460 2261
rect 3463 2256 3465 2261
rect 3479 2259 3481 2261
rect 3495 2259 3497 2261
rect 3500 2258 3502 2261
rect 3516 2259 3518 2261
rect 3532 2259 3534 2261
rect 3537 2256 3539 2261
rect 3558 2256 3560 2261
rect 3574 2259 3576 2261
rect 3590 2259 3592 2261
rect 3595 2256 3597 2261
rect 3611 2259 3613 2261
rect 2518 2221 2520 2224
rect 2542 2221 2544 2224
rect 3463 2221 3465 2224
rect 3487 2221 3489 2224
rect 2518 2215 2520 2217
rect 2542 2215 2544 2217
rect 3463 2215 3465 2217
rect 3487 2215 3489 2217
rect 2538 2210 2540 2212
rect 3483 2210 3485 2212
rect 2538 2203 2540 2206
rect 3483 2203 3485 2206
rect 2527 2192 2529 2194
rect 2533 2192 2552 2194
rect 3472 2192 3474 2194
rect 3478 2192 3497 2194
rect 2518 2187 2520 2189
rect 2542 2187 2544 2189
rect 3463 2187 3465 2189
rect 3487 2187 3489 2189
rect 2518 2180 2520 2183
rect 2542 2180 2544 2183
rect 3463 2180 3465 2183
rect 3487 2180 3489 2183
rect 2286 2152 2288 2154
rect 2291 2152 2293 2155
rect 2307 2152 2309 2154
rect 2323 2152 2325 2154
rect 2328 2152 2330 2155
rect 2349 2152 2351 2155
rect 2365 2152 2367 2155
rect 2381 2152 2383 2154
rect 2386 2152 2388 2155
rect 2402 2152 2404 2154
rect 2418 2152 2420 2154
rect 2423 2152 2425 2155
rect 2439 2152 2441 2154
rect 2455 2152 2457 2154
rect 2460 2152 2462 2155
rect 2481 2152 2483 2155
rect 2497 2152 2499 2155
rect 2513 2152 2515 2154
rect 2518 2152 2520 2155
rect 2534 2152 2536 2154
rect 2550 2152 2552 2154
rect 2555 2152 2557 2155
rect 2571 2152 2573 2154
rect 2587 2152 2589 2154
rect 2592 2152 2594 2155
rect 2613 2152 2615 2155
rect 2629 2152 2631 2155
rect 2645 2152 2647 2154
rect 2650 2152 2652 2155
rect 2666 2152 2668 2154
rect 3231 2152 3233 2154
rect 3236 2152 3238 2155
rect 3252 2152 3254 2154
rect 3268 2152 3270 2154
rect 3273 2152 3275 2155
rect 3294 2152 3296 2155
rect 3310 2152 3312 2155
rect 3326 2152 3328 2154
rect 3331 2152 3333 2155
rect 3347 2152 3349 2154
rect 3363 2152 3365 2154
rect 3368 2152 3370 2155
rect 3384 2152 3386 2154
rect 3400 2152 3402 2154
rect 3405 2152 3407 2155
rect 3426 2152 3428 2155
rect 3442 2152 3444 2155
rect 3458 2152 3460 2154
rect 3463 2152 3465 2155
rect 3479 2152 3481 2154
rect 3495 2152 3497 2154
rect 3500 2152 3502 2155
rect 3516 2152 3518 2154
rect 3532 2152 3534 2154
rect 3537 2152 3539 2155
rect 3558 2152 3560 2155
rect 3574 2152 3576 2155
rect 3590 2152 3592 2154
rect 3595 2152 3597 2155
rect 3611 2152 3613 2154
rect 2286 2139 2288 2144
rect 2291 2142 2293 2144
rect 2286 2125 2288 2135
rect 2291 2125 2293 2132
rect 2307 2125 2309 2144
rect 2323 2135 2325 2144
rect 2328 2142 2330 2144
rect 2349 2142 2351 2144
rect 2365 2141 2367 2144
rect 2323 2125 2325 2128
rect 2328 2125 2330 2127
rect 2349 2125 2351 2127
rect 2365 2125 2367 2137
rect 2381 2135 2383 2144
rect 2386 2142 2388 2144
rect 2381 2125 2383 2128
rect 2386 2125 2388 2127
rect 2402 2125 2404 2144
rect 2418 2141 2420 2144
rect 2423 2142 2425 2144
rect 2418 2125 2420 2137
rect 2423 2125 2425 2132
rect 2439 2125 2441 2144
rect 2455 2135 2457 2144
rect 2460 2142 2462 2144
rect 2481 2142 2483 2144
rect 2497 2141 2499 2144
rect 2455 2125 2457 2128
rect 2460 2125 2462 2127
rect 2481 2125 2483 2127
rect 2497 2125 2499 2137
rect 2513 2135 2515 2144
rect 2518 2142 2520 2144
rect 2513 2125 2515 2128
rect 2518 2125 2520 2127
rect 2534 2125 2536 2144
rect 2550 2141 2552 2144
rect 2555 2142 2557 2144
rect 2550 2125 2552 2137
rect 2555 2125 2557 2132
rect 2571 2125 2573 2144
rect 2587 2135 2589 2144
rect 2592 2142 2594 2144
rect 2613 2142 2615 2144
rect 2629 2141 2631 2144
rect 2587 2125 2589 2128
rect 2592 2125 2594 2127
rect 2613 2125 2615 2127
rect 2629 2125 2631 2137
rect 2645 2135 2647 2144
rect 2650 2142 2652 2144
rect 2666 2136 2668 2144
rect 3231 2139 3233 2144
rect 3236 2142 3238 2144
rect 2645 2125 2647 2128
rect 2650 2125 2652 2127
rect 2666 2125 2668 2132
rect 3231 2125 3233 2135
rect 3236 2125 3238 2132
rect 3252 2125 3254 2144
rect 3268 2135 3270 2144
rect 3273 2142 3275 2144
rect 3294 2142 3296 2144
rect 3310 2141 3312 2144
rect 3268 2125 3270 2128
rect 3273 2125 3275 2127
rect 3294 2125 3296 2127
rect 3310 2125 3312 2137
rect 3326 2135 3328 2144
rect 3331 2142 3333 2144
rect 3326 2125 3328 2128
rect 3331 2125 3333 2127
rect 3347 2125 3349 2144
rect 3363 2141 3365 2144
rect 3368 2142 3370 2144
rect 3363 2125 3365 2137
rect 3368 2125 3370 2132
rect 3384 2125 3386 2144
rect 3400 2135 3402 2144
rect 3405 2142 3407 2144
rect 3426 2142 3428 2144
rect 3442 2141 3444 2144
rect 3400 2125 3402 2128
rect 3405 2125 3407 2127
rect 3426 2125 3428 2127
rect 3442 2125 3444 2137
rect 3458 2135 3460 2144
rect 3463 2142 3465 2144
rect 3458 2125 3460 2128
rect 3463 2125 3465 2127
rect 3479 2125 3481 2144
rect 3495 2141 3497 2144
rect 3500 2142 3502 2144
rect 3495 2125 3497 2137
rect 3500 2125 3502 2132
rect 3516 2125 3518 2144
rect 3532 2135 3534 2144
rect 3537 2142 3539 2144
rect 3558 2142 3560 2144
rect 3574 2141 3576 2144
rect 3532 2125 3534 2128
rect 3537 2125 3539 2127
rect 3558 2125 3560 2127
rect 3574 2125 3576 2137
rect 3590 2135 3592 2144
rect 3595 2142 3597 2144
rect 3611 2136 3613 2144
rect 3590 2125 3592 2128
rect 3595 2125 3597 2127
rect 3611 2125 3613 2132
rect 2286 2119 2288 2121
rect 2291 2118 2293 2121
rect 2307 2119 2309 2121
rect 2323 2119 2325 2121
rect 2328 2116 2330 2121
rect 2349 2116 2351 2121
rect 2365 2119 2367 2121
rect 2381 2119 2383 2121
rect 2386 2116 2388 2121
rect 2402 2119 2404 2121
rect 2418 2119 2420 2121
rect 2423 2118 2425 2121
rect 2439 2119 2441 2121
rect 2455 2119 2457 2121
rect 2460 2116 2462 2121
rect 2481 2116 2483 2121
rect 2497 2119 2499 2121
rect 2513 2119 2515 2121
rect 2518 2116 2520 2121
rect 2534 2119 2536 2121
rect 2550 2119 2552 2121
rect 2555 2118 2557 2121
rect 2571 2119 2573 2121
rect 2587 2119 2589 2121
rect 2592 2116 2594 2121
rect 2613 2116 2615 2121
rect 2629 2119 2631 2121
rect 2645 2119 2647 2121
rect 2650 2116 2652 2121
rect 2666 2119 2668 2121
rect 3231 2119 3233 2121
rect 3236 2118 3238 2121
rect 3252 2119 3254 2121
rect 3268 2119 3270 2121
rect 3273 2116 3275 2121
rect 3294 2116 3296 2121
rect 3310 2119 3312 2121
rect 3326 2119 3328 2121
rect 3331 2116 3333 2121
rect 3347 2119 3349 2121
rect 3363 2119 3365 2121
rect 3368 2118 3370 2121
rect 3384 2119 3386 2121
rect 3400 2119 3402 2121
rect 3405 2116 3407 2121
rect 3426 2116 3428 2121
rect 3442 2119 3444 2121
rect 3458 2119 3460 2121
rect 3463 2116 3465 2121
rect 3479 2119 3481 2121
rect 3495 2119 3497 2121
rect 3500 2118 3502 2121
rect 3516 2119 3518 2121
rect 3532 2119 3534 2121
rect 3537 2116 3539 2121
rect 3558 2116 3560 2121
rect 3574 2119 3576 2121
rect 3590 2119 3592 2121
rect 3595 2116 3597 2121
rect 3611 2119 3613 2121
<< polycontact >>
rect 2775 4040 2779 4044
rect 2812 4040 2816 4044
rect 2832 4040 2836 4044
rect 2870 4040 2874 4044
rect 2907 4040 2911 4044
rect 2944 4040 2948 4044
rect 2964 4040 2968 4044
rect 3002 4040 3006 4044
rect 3039 4040 3043 4044
rect 3076 4040 3080 4044
rect 3096 4040 3100 4044
rect 3134 4040 3138 4044
rect 3171 4040 3175 4044
rect 3208 4040 3212 4044
rect 3228 4040 3232 4044
rect 3266 4040 3270 4044
rect 3720 4040 3724 4044
rect 3757 4040 3761 4044
rect 3777 4040 3781 4044
rect 3815 4040 3819 4044
rect 3852 4040 3856 4044
rect 3889 4040 3893 4044
rect 3909 4040 3913 4044
rect 3947 4040 3951 4044
rect 3984 4040 3988 4044
rect 4021 4040 4025 4044
rect 4041 4040 4045 4044
rect 4079 4040 4083 4044
rect 4116 4040 4120 4044
rect 4153 4040 4157 4044
rect 4173 4040 4177 4044
rect 4211 4040 4215 4044
rect 2769 4020 2773 4024
rect 2787 4022 2791 4026
rect 2423 4007 2427 4011
rect 2460 4007 2464 4011
rect 2480 4007 2484 4011
rect 2518 4007 2522 4011
rect 2847 4022 2851 4026
rect 2805 4013 2809 4020
rect 2863 4013 2867 4020
rect 2884 4017 2888 4021
rect 2901 4020 2905 4024
rect 2919 4022 2923 4026
rect 2979 4022 2983 4026
rect 2937 4013 2941 4020
rect 2995 4013 2999 4020
rect 3016 4017 3020 4021
rect 3033 4020 3037 4024
rect 3051 4022 3055 4026
rect 3111 4022 3115 4026
rect 3069 4013 3073 4020
rect 3127 4013 3131 4020
rect 3148 4017 3152 4021
rect 3165 4020 3169 4024
rect 3183 4022 3187 4026
rect 3243 4022 3247 4026
rect 3201 4013 3205 4020
rect 3259 4013 3263 4020
rect 3280 4017 3284 4021
rect 3714 4020 3718 4024
rect 3732 4022 3736 4026
rect 3368 4007 3372 4011
rect 3405 4007 3409 4011
rect 3425 4007 3429 4011
rect 3463 4007 3467 4011
rect 3792 4022 3796 4026
rect 3750 4013 3754 4020
rect 3808 4013 3812 4020
rect 3829 4017 3833 4021
rect 3846 4020 3850 4024
rect 3864 4022 3868 4026
rect 3924 4022 3928 4026
rect 3882 4013 3886 4020
rect 3940 4013 3944 4020
rect 3961 4017 3965 4021
rect 3978 4020 3982 4024
rect 3996 4022 4000 4026
rect 4056 4022 4060 4026
rect 4014 4013 4018 4020
rect 4072 4013 4076 4020
rect 4093 4017 4097 4021
rect 4110 4020 4114 4024
rect 4128 4022 4132 4026
rect 4188 4022 4192 4026
rect 4146 4013 4150 4020
rect 4204 4013 4208 4020
rect 4225 4017 4229 4021
rect 2775 3999 2779 4003
rect 2812 3997 2816 4001
rect 2832 3997 2836 4001
rect 2868 3997 2872 4001
rect 2907 3999 2911 4003
rect 2944 3997 2948 4001
rect 2964 3997 2968 4001
rect 3000 3997 3004 4001
rect 3039 3999 3043 4003
rect 3076 3997 3080 4001
rect 3096 3997 3100 4001
rect 3132 3997 3136 4001
rect 3171 3999 3175 4003
rect 3208 3997 3212 4001
rect 3228 3997 3232 4001
rect 3264 3997 3268 4001
rect 3720 3999 3724 4003
rect 3757 3997 3761 4001
rect 3777 3997 3781 4001
rect 3813 3997 3817 4001
rect 3852 3999 3856 4003
rect 3889 3997 3893 4001
rect 3909 3997 3913 4001
rect 3945 3997 3949 4001
rect 3984 3999 3988 4003
rect 4021 3997 4025 4001
rect 4041 3997 4045 4001
rect 4077 3997 4081 4001
rect 4116 3999 4120 4003
rect 4153 3997 4157 4001
rect 4173 3997 4177 4001
rect 4209 3997 4213 4001
rect 2417 3987 2421 3991
rect 2435 3989 2439 3993
rect 2495 3989 2499 3993
rect 2453 3980 2457 3987
rect 2511 3980 2515 3987
rect 2530 3984 2534 3988
rect 3362 3987 3366 3991
rect 3380 3989 3384 3993
rect 3440 3989 3444 3993
rect 3398 3980 3402 3987
rect 3456 3980 3460 3987
rect 3475 3984 3479 3988
rect 2423 3966 2427 3970
rect 2460 3964 2464 3968
rect 2480 3964 2484 3968
rect 2516 3964 2520 3968
rect 2791 3956 2795 3960
rect 2835 3956 2839 3960
rect 2862 3956 2866 3960
rect 2907 3956 2911 3960
rect 2980 3963 2984 3967
rect 2541 3943 2545 3947
rect 2945 3949 2949 3953
rect 2424 3934 2428 3938
rect 2771 3936 2775 3940
rect 2803 3937 2807 3941
rect 2822 3936 2826 3940
rect 2878 3937 2882 3941
rect 2894 3936 2898 3940
rect 2921 3936 2925 3940
rect 3061 3963 3065 3967
rect 3368 3966 3372 3970
rect 2972 3945 2976 3949
rect 2999 3941 3003 3945
rect 3026 3949 3030 3953
rect 3405 3964 3409 3968
rect 3425 3964 3429 3968
rect 3461 3964 3465 3968
rect 3053 3945 3057 3949
rect 3080 3941 3084 3945
rect 3736 3956 3740 3960
rect 3780 3956 3784 3960
rect 3807 3956 3811 3960
rect 3852 3956 3856 3960
rect 3925 3963 3929 3967
rect 3486 3943 3490 3947
rect 3890 3949 3894 3953
rect 2978 3927 2982 3931
rect 3369 3934 3373 3938
rect 3716 3936 3720 3940
rect 3059 3927 3063 3931
rect 3748 3937 3752 3941
rect 3767 3936 3771 3940
rect 3823 3937 3827 3941
rect 3839 3936 3843 3940
rect 3866 3936 3870 3940
rect 4006 3963 4010 3967
rect 3917 3945 3921 3949
rect 3944 3941 3948 3945
rect 3971 3949 3975 3953
rect 3998 3945 4002 3949
rect 4025 3941 4029 3945
rect 3923 3927 3927 3931
rect 4004 3927 4008 3931
rect 2788 3919 2792 3923
rect 2832 3918 2836 3922
rect 2857 3919 2862 3923
rect 2904 3918 2908 3922
rect 3733 3919 3737 3923
rect 3777 3918 3781 3922
rect 3802 3919 3807 3923
rect 3849 3918 3853 3922
rect 2423 3905 2427 3909
rect 2461 3905 2465 3909
rect 2481 3905 2485 3909
rect 2518 3905 2522 3909
rect 3368 3905 3372 3909
rect 3406 3905 3410 3909
rect 3426 3905 3430 3909
rect 3463 3905 3467 3909
rect 2411 3882 2415 3886
rect 2446 3887 2450 3891
rect 2430 3878 2434 3885
rect 2488 3878 2492 3885
rect 2506 3887 2510 3891
rect 2788 3889 2792 3893
rect 2832 3890 2836 3894
rect 2524 3885 2528 3889
rect 2857 3889 2862 3893
rect 2904 3890 2908 3894
rect 2980 3887 2984 3891
rect 3061 3887 3065 3891
rect 2771 3872 2775 3876
rect 2425 3862 2429 3866
rect 2461 3862 2465 3866
rect 2481 3862 2485 3866
rect 2518 3864 2522 3868
rect 2803 3871 2807 3875
rect 2822 3872 2826 3876
rect 2878 3871 2882 3875
rect 2894 3872 2898 3876
rect 2921 3872 2925 3876
rect 2969 3871 2975 3875
rect 3050 3871 3056 3875
rect 3356 3882 3360 3886
rect 3391 3887 3395 3891
rect 3375 3878 3379 3885
rect 3433 3878 3437 3885
rect 3451 3887 3455 3891
rect 3733 3889 3737 3893
rect 3777 3890 3781 3894
rect 3469 3885 3473 3889
rect 3802 3889 3807 3893
rect 3849 3890 3853 3894
rect 3925 3887 3929 3891
rect 4006 3887 4010 3891
rect 3716 3872 3720 3876
rect 3370 3862 3374 3866
rect 3406 3862 3410 3866
rect 3426 3862 3430 3866
rect 3463 3864 3467 3868
rect 3748 3871 3752 3875
rect 3767 3872 3771 3876
rect 3823 3871 3827 3875
rect 3839 3872 3843 3876
rect 3866 3872 3870 3876
rect 3914 3871 3920 3875
rect 3995 3871 4001 3875
rect 2791 3852 2795 3856
rect 2835 3852 2839 3856
rect 2862 3852 2866 3856
rect 2907 3852 2911 3856
rect 2978 3851 2982 3855
rect 3059 3851 3063 3855
rect 3736 3852 3740 3856
rect 3780 3852 3784 3856
rect 3807 3852 3811 3856
rect 3852 3852 3856 3856
rect 3923 3851 3927 3855
rect 4004 3851 4008 3855
rect 2980 3831 2984 3835
rect 2791 3824 2795 3828
rect 2835 3824 2839 3828
rect 2862 3824 2866 3828
rect 2907 3824 2911 3828
rect 3085 3831 3089 3835
rect 2972 3813 2976 3817
rect 2771 3804 2775 3808
rect 2803 3805 2807 3809
rect 2822 3804 2826 3808
rect 2878 3805 2882 3809
rect 2894 3804 2898 3808
rect 2921 3804 2925 3808
rect 2999 3809 3003 3813
rect 3050 3817 3054 3821
rect 3925 3831 3929 3835
rect 3077 3813 3081 3817
rect 3104 3809 3108 3813
rect 3736 3824 3740 3828
rect 3780 3824 3784 3828
rect 3807 3824 3811 3828
rect 3852 3824 3856 3828
rect 4030 3831 4034 3835
rect 3917 3813 3921 3817
rect 2978 3795 2982 3799
rect 3083 3795 3087 3799
rect 3316 3802 3320 3806
rect 2788 3787 2792 3791
rect 2832 3786 2836 3790
rect 2857 3787 2862 3791
rect 2904 3786 2908 3790
rect 3281 3788 3285 3792
rect 3716 3804 3720 3808
rect 3308 3784 3312 3788
rect 3335 3780 3339 3784
rect 3748 3805 3752 3809
rect 3767 3804 3771 3808
rect 3823 3805 3827 3809
rect 3839 3804 3843 3808
rect 3866 3804 3870 3808
rect 3944 3809 3948 3813
rect 3995 3817 3999 3821
rect 4022 3813 4026 3817
rect 4049 3809 4053 3813
rect 3923 3795 3927 3799
rect 4028 3795 4032 3799
rect 3733 3787 3737 3791
rect 3777 3786 3781 3790
rect 3802 3787 3807 3791
rect 3849 3786 3853 3790
rect 3314 3766 3318 3770
rect 2788 3757 2792 3761
rect 2832 3758 2836 3762
rect 2857 3757 2862 3761
rect 2904 3758 2908 3762
rect 3469 3760 3473 3764
rect 3522 3760 3526 3764
rect 2980 3756 2984 3760
rect 3085 3756 3089 3760
rect 3733 3757 3737 3761
rect 3777 3758 3781 3762
rect 3802 3757 3807 3761
rect 3849 3758 3853 3762
rect 3925 3756 3929 3760
rect 4030 3756 4034 3760
rect 2771 3740 2775 3744
rect 2803 3739 2807 3743
rect 2822 3740 2826 3744
rect 2878 3739 2882 3743
rect 2894 3740 2898 3744
rect 2921 3740 2925 3744
rect 2969 3740 2975 3744
rect 3074 3740 3080 3744
rect 3716 3740 3720 3744
rect 3748 3739 3752 3743
rect 3767 3740 3771 3744
rect 3823 3739 3827 3743
rect 3839 3740 3843 3744
rect 3866 3740 3870 3744
rect 3914 3740 3920 3744
rect 4019 3740 4025 3744
rect 2791 3720 2795 3724
rect 2835 3720 2839 3724
rect 2862 3720 2866 3724
rect 2907 3720 2911 3724
rect 2978 3720 2982 3724
rect 3083 3720 3087 3724
rect 3316 3722 3320 3726
rect 3736 3720 3740 3724
rect 3780 3720 3784 3724
rect 3807 3720 3811 3724
rect 3852 3720 3856 3724
rect 3923 3720 3927 3724
rect 4028 3720 4032 3724
rect 3305 3706 3311 3710
rect 2980 3699 2984 3703
rect 2791 3692 2795 3696
rect 2835 3692 2839 3696
rect 2862 3692 2866 3696
rect 2907 3692 2911 3696
rect 3061 3699 3065 3703
rect 2972 3681 2976 3685
rect 2771 3672 2775 3676
rect 2803 3673 2807 3677
rect 2822 3672 2826 3676
rect 2878 3673 2882 3677
rect 2894 3672 2898 3676
rect 2921 3672 2925 3676
rect 2999 3677 3003 3681
rect 3026 3685 3030 3689
rect 3151 3699 3155 3703
rect 3053 3681 3057 3685
rect 3080 3677 3084 3681
rect 3116 3685 3120 3689
rect 3925 3699 3929 3703
rect 3143 3681 3147 3685
rect 3170 3677 3174 3681
rect 3736 3692 3740 3696
rect 3780 3692 3784 3696
rect 3807 3692 3811 3696
rect 3852 3692 3856 3696
rect 3314 3686 3318 3690
rect 4006 3699 4010 3703
rect 3917 3681 3921 3685
rect 2978 3663 2982 3667
rect 3059 3663 3063 3667
rect 3149 3663 3153 3667
rect 3316 3672 3320 3676
rect 2788 3655 2792 3659
rect 2832 3654 2836 3658
rect 2857 3655 2862 3659
rect 3259 3658 3263 3662
rect 2904 3654 2908 3658
rect 3281 3658 3285 3662
rect 3716 3672 3720 3676
rect 3308 3654 3312 3658
rect 3335 3650 3339 3654
rect 3748 3673 3752 3677
rect 3767 3672 3771 3676
rect 3823 3673 3827 3677
rect 3839 3672 3843 3676
rect 3866 3672 3870 3676
rect 3944 3677 3948 3681
rect 3971 3685 3975 3689
rect 4096 3699 4100 3703
rect 3998 3681 4002 3685
rect 4025 3677 4029 3681
rect 4061 3685 4065 3689
rect 4088 3681 4092 3685
rect 4115 3677 4119 3681
rect 3923 3663 3927 3667
rect 4004 3663 4008 3667
rect 4094 3663 4098 3667
rect 3733 3655 3737 3659
rect 3777 3654 3781 3658
rect 3802 3655 3807 3659
rect 3849 3654 3853 3658
rect 3314 3636 3318 3640
rect 2788 3625 2792 3629
rect 2832 3626 2836 3630
rect 3375 3630 3379 3634
rect 3428 3630 3432 3634
rect 2857 3625 2862 3629
rect 2904 3626 2908 3630
rect 2980 3621 2984 3625
rect 3061 3621 3065 3625
rect 3151 3621 3155 3625
rect 3733 3625 3737 3629
rect 3777 3626 3781 3630
rect 2771 3608 2775 3612
rect 2803 3607 2807 3611
rect 2822 3608 2826 3612
rect 2878 3607 2882 3611
rect 2894 3608 2898 3612
rect 2921 3608 2925 3612
rect 2969 3605 2975 3609
rect 3050 3605 3056 3609
rect 3140 3605 3146 3609
rect 3802 3625 3807 3629
rect 3849 3626 3853 3630
rect 3925 3621 3929 3625
rect 4006 3621 4010 3625
rect 4096 3621 4100 3625
rect 3716 3608 3720 3612
rect 3748 3607 3752 3611
rect 3767 3608 3771 3612
rect 3823 3607 3827 3611
rect 3839 3608 3843 3612
rect 3866 3608 3870 3612
rect 3914 3605 3920 3609
rect 2791 3588 2795 3592
rect 2835 3588 2839 3592
rect 2862 3588 2866 3592
rect 2907 3588 2911 3592
rect 3316 3592 3320 3596
rect 3995 3605 4001 3609
rect 4085 3605 4091 3609
rect 2978 3585 2982 3589
rect 3059 3585 3063 3589
rect 3149 3585 3153 3589
rect 3736 3588 3740 3592
rect 3780 3588 3784 3592
rect 3807 3588 3811 3592
rect 3852 3588 3856 3592
rect 3923 3585 3927 3589
rect 4004 3585 4008 3589
rect 4094 3585 4098 3589
rect 3305 3576 3311 3580
rect 2980 3567 2984 3571
rect 2791 3560 2795 3564
rect 2835 3560 2839 3564
rect 2862 3560 2866 3564
rect 2907 3560 2911 3564
rect 2972 3549 2976 3553
rect 2771 3540 2775 3544
rect 2803 3541 2807 3545
rect 2822 3540 2826 3544
rect 2878 3541 2882 3545
rect 2894 3540 2898 3544
rect 2921 3540 2925 3544
rect 2999 3545 3003 3549
rect 3314 3556 3318 3560
rect 3925 3567 3929 3571
rect 3736 3560 3740 3564
rect 3780 3560 3784 3564
rect 3807 3560 3811 3564
rect 3852 3560 3856 3564
rect 3917 3549 3921 3553
rect 3716 3540 3720 3544
rect 2978 3531 2982 3535
rect 3748 3541 3752 3545
rect 3767 3540 3771 3544
rect 3823 3541 3827 3545
rect 3839 3540 3843 3544
rect 3866 3540 3870 3544
rect 3944 3545 3948 3549
rect 3923 3531 3927 3535
rect 2788 3523 2792 3527
rect 2832 3522 2836 3526
rect 2857 3523 2862 3527
rect 2904 3522 2908 3526
rect 3733 3523 3737 3527
rect 3777 3522 3781 3526
rect 3802 3523 3807 3527
rect 3849 3522 3853 3526
rect 2291 3505 2295 3509
rect 2328 3505 2332 3509
rect 2348 3505 2352 3509
rect 2386 3505 2390 3509
rect 2423 3505 2427 3509
rect 2460 3505 2464 3509
rect 2480 3505 2484 3509
rect 2518 3505 2522 3509
rect 2555 3505 2559 3509
rect 2592 3505 2596 3509
rect 2612 3505 2616 3509
rect 2650 3505 2654 3509
rect 3236 3505 3240 3509
rect 3273 3505 3277 3509
rect 3293 3505 3297 3509
rect 3331 3505 3335 3509
rect 3368 3505 3372 3509
rect 3405 3505 3409 3509
rect 3425 3505 3429 3509
rect 3463 3505 3467 3509
rect 3500 3505 3504 3509
rect 3537 3505 3541 3509
rect 3557 3505 3561 3509
rect 3595 3505 3599 3509
rect 2285 3485 2289 3489
rect 2303 3487 2307 3491
rect 2363 3487 2367 3491
rect 2321 3478 2325 3485
rect 2379 3478 2383 3485
rect 2398 3482 2402 3486
rect 2416 3487 2420 3491
rect 2435 3487 2439 3491
rect 2495 3487 2499 3491
rect 2453 3478 2457 3485
rect 2511 3478 2515 3485
rect 2530 3482 2534 3486
rect 2548 3487 2552 3491
rect 2567 3487 2571 3491
rect 2627 3487 2631 3491
rect 2585 3478 2589 3485
rect 2788 3493 2792 3497
rect 2832 3494 2836 3498
rect 2857 3493 2862 3497
rect 2904 3494 2908 3498
rect 3049 3493 3053 3497
rect 3093 3494 3097 3498
rect 3118 3493 3123 3497
rect 3165 3494 3169 3498
rect 2643 3478 2647 3485
rect 2664 3482 2668 3486
rect 2980 3485 2984 3489
rect 3230 3485 3234 3489
rect 3248 3487 3252 3491
rect 2771 3476 2775 3480
rect 2803 3475 2807 3479
rect 2822 3476 2826 3480
rect 2878 3475 2882 3479
rect 2894 3476 2898 3480
rect 2921 3476 2925 3480
rect 2291 3464 2295 3468
rect 2328 3462 2332 3466
rect 2348 3462 2352 3466
rect 2384 3462 2388 3466
rect 2423 3464 2427 3468
rect 2460 3462 2464 3466
rect 2480 3462 2484 3466
rect 2516 3462 2520 3466
rect 2555 3464 2559 3468
rect 2592 3462 2596 3466
rect 2612 3462 2616 3466
rect 2648 3462 2652 3466
rect 2969 3469 2975 3473
rect 3007 3476 3011 3480
rect 3064 3475 3068 3479
rect 3083 3476 3087 3480
rect 3139 3475 3143 3479
rect 3155 3476 3159 3480
rect 3182 3476 3186 3480
rect 3308 3487 3312 3491
rect 3266 3478 3270 3485
rect 3324 3478 3328 3485
rect 3343 3482 3347 3486
rect 3361 3487 3365 3491
rect 3380 3487 3384 3491
rect 3440 3487 3444 3491
rect 3398 3478 3402 3485
rect 3456 3478 3460 3485
rect 3475 3482 3479 3486
rect 3493 3487 3497 3491
rect 3512 3487 3516 3491
rect 3572 3487 3576 3491
rect 3530 3478 3534 3485
rect 3733 3493 3737 3497
rect 3777 3494 3781 3498
rect 3802 3493 3807 3497
rect 3849 3494 3853 3498
rect 3994 3493 3998 3497
rect 4038 3494 4042 3498
rect 4063 3493 4068 3497
rect 4110 3494 4114 3498
rect 3588 3478 3592 3485
rect 3609 3482 3613 3486
rect 3925 3485 3929 3489
rect 3716 3476 3720 3480
rect 3748 3475 3752 3479
rect 3767 3476 3771 3480
rect 3823 3475 3827 3479
rect 3839 3476 3843 3480
rect 3866 3476 3870 3480
rect 2791 3456 2795 3460
rect 2835 3456 2839 3460
rect 2862 3456 2866 3460
rect 2907 3456 2911 3460
rect 3236 3464 3240 3468
rect 2978 3449 2982 3453
rect 2400 3434 2404 3438
rect 2424 3434 2428 3438
rect 3273 3462 3277 3466
rect 3293 3462 3297 3466
rect 3329 3462 3333 3466
rect 3368 3464 3372 3468
rect 3405 3462 3409 3466
rect 3425 3462 3429 3466
rect 3461 3462 3465 3466
rect 3500 3464 3504 3468
rect 3537 3462 3541 3466
rect 3557 3462 3561 3466
rect 3593 3462 3597 3466
rect 3914 3469 3920 3473
rect 3952 3476 3956 3480
rect 4009 3475 4013 3479
rect 4028 3476 4032 3480
rect 4084 3475 4088 3479
rect 4100 3476 4104 3480
rect 4127 3476 4131 3480
rect 3052 3456 3056 3460
rect 3096 3456 3100 3460
rect 3123 3456 3127 3460
rect 3168 3456 3172 3460
rect 3736 3456 3740 3460
rect 3780 3456 3784 3460
rect 3807 3456 3811 3460
rect 3852 3456 3856 3460
rect 3923 3449 3927 3453
rect 3345 3434 3349 3438
rect 3369 3434 3373 3438
rect 3191 3428 3195 3432
rect 3029 3421 3033 3425
rect 3997 3456 4001 3460
rect 4041 3456 4045 3460
rect 4068 3456 4072 3460
rect 4113 3456 4117 3460
rect 4136 3428 4140 3432
rect 3972 3421 3976 3425
rect 2420 3407 2424 3411
rect 3365 3407 3369 3411
rect 2435 3399 2439 3403
rect 3380 3399 3384 3403
rect 3074 3393 3078 3397
rect 3111 3393 3115 3397
rect 3131 3393 3135 3397
rect 3169 3393 3173 3397
rect 4019 3393 4023 3397
rect 4056 3393 4060 3397
rect 4076 3393 4080 3397
rect 4114 3393 4118 3397
rect 2400 3384 2404 3388
rect 2424 3384 2428 3388
rect 3345 3384 3349 3388
rect 3369 3384 3373 3388
rect 3068 3373 3072 3377
rect 3086 3375 3090 3379
rect 2291 3363 2295 3367
rect 2328 3363 2332 3367
rect 2348 3363 2352 3367
rect 2386 3363 2390 3367
rect 2423 3363 2427 3367
rect 2460 3363 2464 3367
rect 2480 3363 2484 3367
rect 2518 3363 2522 3367
rect 2555 3363 2559 3367
rect 2592 3363 2596 3367
rect 2612 3363 2616 3367
rect 2650 3363 2654 3367
rect 3146 3375 3150 3379
rect 3104 3366 3108 3373
rect 3162 3366 3166 3373
rect 3181 3370 3185 3374
rect 4013 3373 4017 3377
rect 4031 3375 4035 3379
rect 3236 3363 3240 3367
rect 3273 3363 3277 3367
rect 3293 3363 3297 3367
rect 3331 3363 3335 3367
rect 3368 3363 3372 3367
rect 3405 3363 3409 3367
rect 3425 3363 3429 3367
rect 3463 3363 3467 3367
rect 3500 3363 3504 3367
rect 3537 3363 3541 3367
rect 3557 3363 3561 3367
rect 3595 3363 3599 3367
rect 4091 3375 4095 3379
rect 4049 3366 4053 3373
rect 4107 3366 4111 3373
rect 4126 3370 4130 3374
rect 3074 3352 3078 3356
rect 2285 3343 2289 3347
rect 2303 3345 2307 3349
rect 2363 3345 2367 3349
rect 2321 3336 2325 3343
rect 2379 3336 2383 3343
rect 2398 3340 2402 3344
rect 2416 3345 2420 3349
rect 2435 3345 2439 3349
rect 2495 3345 2499 3349
rect 2453 3336 2457 3343
rect 2511 3336 2515 3343
rect 2530 3340 2534 3344
rect 2548 3345 2552 3349
rect 2567 3345 2571 3349
rect 2627 3345 2631 3349
rect 2585 3336 2589 3343
rect 3111 3350 3115 3354
rect 3131 3350 3135 3354
rect 3167 3350 3171 3354
rect 4019 3352 4023 3356
rect 2643 3336 2647 3343
rect 2664 3340 2668 3344
rect 3230 3343 3234 3347
rect 3248 3345 3252 3349
rect 3308 3345 3312 3349
rect 3266 3336 3270 3343
rect 3324 3336 3328 3343
rect 3343 3340 3347 3344
rect 3361 3345 3365 3349
rect 3380 3345 3384 3349
rect 3440 3345 3444 3349
rect 3398 3336 3402 3343
rect 3456 3336 3460 3343
rect 3475 3340 3479 3344
rect 3493 3345 3497 3349
rect 3512 3345 3516 3349
rect 3572 3345 3576 3349
rect 3530 3336 3534 3343
rect 4056 3350 4060 3354
rect 4076 3350 4080 3354
rect 4112 3350 4116 3354
rect 3588 3336 3592 3343
rect 3609 3340 3613 3344
rect 2291 3322 2295 3326
rect 2328 3320 2332 3324
rect 2348 3320 2352 3324
rect 2384 3320 2388 3324
rect 2423 3322 2427 3326
rect 2460 3320 2464 3324
rect 2480 3320 2484 3324
rect 2516 3320 2520 3324
rect 2555 3322 2559 3326
rect 2592 3320 2596 3324
rect 2612 3320 2616 3324
rect 2648 3320 2652 3324
rect 3236 3322 3240 3326
rect 3273 3320 3277 3324
rect 3293 3320 3297 3324
rect 3329 3320 3333 3324
rect 3368 3322 3372 3326
rect 3405 3320 3409 3324
rect 3425 3320 3429 3324
rect 3461 3320 3465 3324
rect 3500 3322 3504 3326
rect 3537 3320 3541 3324
rect 3557 3320 3561 3324
rect 3593 3320 3597 3324
rect 3074 3307 3078 3311
rect 3111 3307 3115 3311
rect 3131 3307 3135 3311
rect 3169 3307 3173 3311
rect 4019 3307 4023 3311
rect 4056 3307 4060 3311
rect 4076 3307 4080 3311
rect 4114 3307 4118 3311
rect 3068 3287 3072 3291
rect 3086 3289 3090 3293
rect 2291 3277 2295 3281
rect 2328 3277 2332 3281
rect 2348 3277 2352 3281
rect 2386 3277 2390 3281
rect 2423 3277 2427 3281
rect 2460 3277 2464 3281
rect 2480 3277 2484 3281
rect 2518 3277 2522 3281
rect 2555 3277 2559 3281
rect 2592 3277 2596 3281
rect 2612 3277 2616 3281
rect 2650 3277 2654 3281
rect 3146 3289 3150 3293
rect 3104 3280 3108 3287
rect 3162 3280 3166 3287
rect 3181 3284 3185 3288
rect 3203 3282 3207 3286
rect 4013 3287 4017 3291
rect 4031 3289 4035 3293
rect 3236 3277 3240 3281
rect 3273 3277 3277 3281
rect 3293 3277 3297 3281
rect 3331 3277 3335 3281
rect 3368 3277 3372 3281
rect 3405 3277 3409 3281
rect 3425 3277 3429 3281
rect 3463 3277 3467 3281
rect 3500 3277 3504 3281
rect 3537 3277 3541 3281
rect 3557 3277 3561 3281
rect 3595 3277 3599 3281
rect 4091 3289 4095 3293
rect 4049 3280 4053 3287
rect 4107 3280 4111 3287
rect 4126 3284 4130 3288
rect 4148 3282 4152 3286
rect 3074 3266 3078 3270
rect 2285 3257 2289 3261
rect 2303 3259 2307 3263
rect 2363 3259 2367 3263
rect 2321 3250 2325 3257
rect 2379 3250 2383 3257
rect 2398 3254 2402 3258
rect 2416 3259 2420 3263
rect 2435 3259 2439 3263
rect 2495 3259 2499 3263
rect 2453 3250 2457 3257
rect 2511 3250 2515 3257
rect 2530 3254 2534 3258
rect 2548 3259 2552 3263
rect 2567 3259 2571 3263
rect 2627 3259 2631 3263
rect 2585 3250 2589 3257
rect 3111 3264 3115 3268
rect 3131 3264 3135 3268
rect 3167 3264 3171 3268
rect 4019 3266 4023 3270
rect 2643 3250 2647 3257
rect 2664 3254 2668 3258
rect 3230 3257 3234 3261
rect 3248 3259 3252 3263
rect 3308 3259 3312 3263
rect 3266 3250 3270 3257
rect 3324 3250 3328 3257
rect 3343 3254 3347 3258
rect 3361 3259 3365 3263
rect 3380 3259 3384 3263
rect 3440 3259 3444 3263
rect 3398 3250 3402 3257
rect 3456 3250 3460 3257
rect 3475 3254 3479 3258
rect 3493 3259 3497 3263
rect 3512 3259 3516 3263
rect 3572 3259 3576 3263
rect 3530 3250 3534 3257
rect 4056 3264 4060 3268
rect 4076 3264 4080 3268
rect 4112 3264 4116 3268
rect 3588 3250 3592 3257
rect 3609 3254 3613 3258
rect 2291 3236 2295 3240
rect 2328 3234 2332 3238
rect 2348 3234 2352 3238
rect 2384 3234 2388 3238
rect 2423 3236 2427 3240
rect 2460 3234 2464 3238
rect 2480 3234 2484 3238
rect 2516 3234 2520 3238
rect 2555 3236 2559 3240
rect 2592 3234 2596 3238
rect 2612 3234 2616 3238
rect 2648 3234 2652 3238
rect 3236 3236 3240 3240
rect 3273 3234 3277 3238
rect 3293 3234 3297 3238
rect 3329 3234 3333 3238
rect 3368 3236 3372 3240
rect 3405 3234 3409 3238
rect 3425 3234 3429 3238
rect 3461 3234 3465 3238
rect 3500 3236 3504 3240
rect 3537 3234 3541 3238
rect 3557 3234 3561 3238
rect 3593 3234 3597 3238
rect 2517 3206 2521 3210
rect 2541 3206 2545 3210
rect 3462 3206 3466 3210
rect 3486 3206 3490 3210
rect 2537 3181 2541 3185
rect 3482 3181 3486 3185
rect 2552 3173 2556 3177
rect 3497 3173 3501 3177
rect 2517 3158 2521 3162
rect 2541 3158 2545 3162
rect 3462 3158 3466 3162
rect 3486 3158 3490 3162
rect 2291 3137 2295 3141
rect 2328 3137 2332 3141
rect 2348 3137 2352 3141
rect 2386 3137 2390 3141
rect 2423 3137 2427 3141
rect 2460 3137 2464 3141
rect 2480 3137 2484 3141
rect 2518 3137 2522 3141
rect 2555 3137 2559 3141
rect 2592 3137 2596 3141
rect 2612 3137 2616 3141
rect 2650 3137 2654 3141
rect 3236 3137 3240 3141
rect 3273 3137 3277 3141
rect 3293 3137 3297 3141
rect 3331 3137 3335 3141
rect 3368 3137 3372 3141
rect 3405 3137 3409 3141
rect 3425 3137 3429 3141
rect 3463 3137 3467 3141
rect 3500 3137 3504 3141
rect 3537 3137 3541 3141
rect 3557 3137 3561 3141
rect 3595 3137 3599 3141
rect 2285 3117 2289 3121
rect 2303 3119 2307 3123
rect 2363 3119 2367 3123
rect 2321 3110 2325 3117
rect 2379 3110 2383 3117
rect 2398 3114 2402 3118
rect 2416 3119 2420 3123
rect 2435 3119 2439 3123
rect 2495 3119 2499 3123
rect 2453 3110 2457 3117
rect 2511 3110 2515 3117
rect 2530 3114 2534 3118
rect 2548 3119 2552 3123
rect 2567 3119 2571 3123
rect 2627 3119 2631 3123
rect 2585 3110 2589 3117
rect 2643 3110 2647 3117
rect 2664 3114 2668 3118
rect 3230 3117 3234 3121
rect 3248 3119 3252 3123
rect 3308 3119 3312 3123
rect 3266 3110 3270 3117
rect 3324 3110 3328 3117
rect 3343 3114 3347 3118
rect 3361 3119 3365 3123
rect 3380 3119 3384 3123
rect 3440 3119 3444 3123
rect 3398 3110 3402 3117
rect 3456 3110 3460 3117
rect 3475 3114 3479 3118
rect 3493 3119 3497 3123
rect 3512 3119 3516 3123
rect 3572 3119 3576 3123
rect 3530 3110 3534 3117
rect 3588 3110 3592 3117
rect 3609 3114 3613 3118
rect 2291 3096 2295 3100
rect 2328 3094 2332 3098
rect 2348 3094 2352 3098
rect 2384 3094 2388 3098
rect 2423 3096 2427 3100
rect 2460 3094 2464 3098
rect 2480 3094 2484 3098
rect 2516 3094 2520 3098
rect 2555 3096 2559 3100
rect 2592 3094 2596 3098
rect 2612 3094 2616 3098
rect 2648 3094 2652 3098
rect 3236 3096 3240 3100
rect 3273 3094 3277 3098
rect 3293 3094 3297 3098
rect 3329 3094 3333 3098
rect 3368 3096 3372 3100
rect 3405 3094 3409 3098
rect 3425 3094 3429 3098
rect 3461 3094 3465 3098
rect 3500 3096 3504 3100
rect 3537 3094 3541 3098
rect 3557 3094 3561 3098
rect 3593 3094 3597 3098
rect 2775 3058 2779 3062
rect 2812 3058 2816 3062
rect 2832 3058 2836 3062
rect 2870 3058 2874 3062
rect 2907 3058 2911 3062
rect 2944 3058 2948 3062
rect 2964 3058 2968 3062
rect 3002 3058 3006 3062
rect 3039 3058 3043 3062
rect 3076 3058 3080 3062
rect 3096 3058 3100 3062
rect 3134 3058 3138 3062
rect 3171 3058 3175 3062
rect 3208 3058 3212 3062
rect 3228 3058 3232 3062
rect 3266 3058 3270 3062
rect 3720 3058 3724 3062
rect 3757 3058 3761 3062
rect 3777 3058 3781 3062
rect 3815 3058 3819 3062
rect 3852 3058 3856 3062
rect 3889 3058 3893 3062
rect 3909 3058 3913 3062
rect 3947 3058 3951 3062
rect 3984 3058 3988 3062
rect 4021 3058 4025 3062
rect 4041 3058 4045 3062
rect 4079 3058 4083 3062
rect 4116 3058 4120 3062
rect 4153 3058 4157 3062
rect 4173 3058 4177 3062
rect 4211 3058 4215 3062
rect 2769 3038 2773 3042
rect 2787 3040 2791 3044
rect 2423 3025 2427 3029
rect 2460 3025 2464 3029
rect 2480 3025 2484 3029
rect 2518 3025 2522 3029
rect 2847 3040 2851 3044
rect 2805 3031 2809 3038
rect 2863 3031 2867 3038
rect 2884 3035 2888 3039
rect 2901 3038 2905 3042
rect 2919 3040 2923 3044
rect 2979 3040 2983 3044
rect 2937 3031 2941 3038
rect 2995 3031 2999 3038
rect 3016 3035 3020 3039
rect 3033 3038 3037 3042
rect 3051 3040 3055 3044
rect 3111 3040 3115 3044
rect 3069 3031 3073 3038
rect 3127 3031 3131 3038
rect 3148 3035 3152 3039
rect 3165 3038 3169 3042
rect 3183 3040 3187 3044
rect 3243 3040 3247 3044
rect 3201 3031 3205 3038
rect 3259 3031 3263 3038
rect 3280 3035 3284 3039
rect 3714 3038 3718 3042
rect 3732 3040 3736 3044
rect 3368 3025 3372 3029
rect 3405 3025 3409 3029
rect 3425 3025 3429 3029
rect 3463 3025 3467 3029
rect 3792 3040 3796 3044
rect 3750 3031 3754 3038
rect 3808 3031 3812 3038
rect 3829 3035 3833 3039
rect 3846 3038 3850 3042
rect 3864 3040 3868 3044
rect 3924 3040 3928 3044
rect 3882 3031 3886 3038
rect 3940 3031 3944 3038
rect 3961 3035 3965 3039
rect 3978 3038 3982 3042
rect 3996 3040 4000 3044
rect 4056 3040 4060 3044
rect 4014 3031 4018 3038
rect 4072 3031 4076 3038
rect 4093 3035 4097 3039
rect 4110 3038 4114 3042
rect 4128 3040 4132 3044
rect 4188 3040 4192 3044
rect 4146 3031 4150 3038
rect 4204 3031 4208 3038
rect 4225 3035 4229 3039
rect 2775 3017 2779 3021
rect 2812 3015 2816 3019
rect 2832 3015 2836 3019
rect 2868 3015 2872 3019
rect 2907 3017 2911 3021
rect 2944 3015 2948 3019
rect 2964 3015 2968 3019
rect 3000 3015 3004 3019
rect 3039 3017 3043 3021
rect 3076 3015 3080 3019
rect 3096 3015 3100 3019
rect 3132 3015 3136 3019
rect 3171 3017 3175 3021
rect 3208 3015 3212 3019
rect 3228 3015 3232 3019
rect 3264 3015 3268 3019
rect 3720 3017 3724 3021
rect 3757 3015 3761 3019
rect 3777 3015 3781 3019
rect 3813 3015 3817 3019
rect 3852 3017 3856 3021
rect 3889 3015 3893 3019
rect 3909 3015 3913 3019
rect 3945 3015 3949 3019
rect 3984 3017 3988 3021
rect 4021 3015 4025 3019
rect 4041 3015 4045 3019
rect 4077 3015 4081 3019
rect 4116 3017 4120 3021
rect 4153 3015 4157 3019
rect 4173 3015 4177 3019
rect 4209 3015 4213 3019
rect 2417 3005 2421 3009
rect 2435 3007 2439 3011
rect 2495 3007 2499 3011
rect 2453 2998 2457 3005
rect 2511 2998 2515 3005
rect 2530 3002 2534 3006
rect 3362 3005 3366 3009
rect 3380 3007 3384 3011
rect 3440 3007 3444 3011
rect 3398 2998 3402 3005
rect 3456 2998 3460 3005
rect 3475 3002 3479 3006
rect 2423 2984 2427 2988
rect 2460 2982 2464 2986
rect 2480 2982 2484 2986
rect 2516 2982 2520 2986
rect 2791 2974 2795 2978
rect 2835 2974 2839 2978
rect 2862 2974 2866 2978
rect 2907 2974 2911 2978
rect 2980 2981 2984 2985
rect 2541 2961 2545 2965
rect 2945 2967 2949 2971
rect 2424 2952 2428 2956
rect 2771 2954 2775 2958
rect 2803 2955 2807 2959
rect 2822 2954 2826 2958
rect 2878 2955 2882 2959
rect 2894 2954 2898 2958
rect 2921 2954 2925 2958
rect 3061 2981 3065 2985
rect 3368 2984 3372 2988
rect 2972 2963 2976 2967
rect 2999 2959 3003 2963
rect 3026 2967 3030 2971
rect 3405 2982 3409 2986
rect 3425 2982 3429 2986
rect 3461 2982 3465 2986
rect 3053 2963 3057 2967
rect 3080 2959 3084 2963
rect 3736 2974 3740 2978
rect 3780 2974 3784 2978
rect 3807 2974 3811 2978
rect 3852 2974 3856 2978
rect 3925 2981 3929 2985
rect 3486 2961 3490 2965
rect 3890 2967 3894 2971
rect 2978 2945 2982 2949
rect 3369 2952 3373 2956
rect 3716 2954 3720 2958
rect 3059 2945 3063 2949
rect 3748 2955 3752 2959
rect 3767 2954 3771 2958
rect 3823 2955 3827 2959
rect 3839 2954 3843 2958
rect 3866 2954 3870 2958
rect 4006 2981 4010 2985
rect 3917 2963 3921 2967
rect 3944 2959 3948 2963
rect 3971 2967 3975 2971
rect 3998 2963 4002 2967
rect 4025 2959 4029 2963
rect 3923 2945 3927 2949
rect 4004 2945 4008 2949
rect 2788 2937 2792 2941
rect 2832 2936 2836 2940
rect 2857 2937 2862 2941
rect 2904 2936 2908 2940
rect 3733 2937 3737 2941
rect 3777 2936 3781 2940
rect 3802 2937 3807 2941
rect 3849 2936 3853 2940
rect 2423 2923 2427 2927
rect 2461 2923 2465 2927
rect 2481 2923 2485 2927
rect 2518 2923 2522 2927
rect 3368 2923 3372 2927
rect 3406 2923 3410 2927
rect 3426 2923 3430 2927
rect 3463 2923 3467 2927
rect 2411 2900 2415 2904
rect 2446 2905 2450 2909
rect 2430 2896 2434 2903
rect 2488 2896 2492 2903
rect 2506 2905 2510 2909
rect 2788 2907 2792 2911
rect 2832 2908 2836 2912
rect 2524 2903 2528 2907
rect 2857 2907 2862 2911
rect 2904 2908 2908 2912
rect 2980 2905 2984 2909
rect 3061 2905 3065 2909
rect 2771 2890 2775 2894
rect 2425 2880 2429 2884
rect 2461 2880 2465 2884
rect 2481 2880 2485 2884
rect 2518 2882 2522 2886
rect 2803 2889 2807 2893
rect 2822 2890 2826 2894
rect 2878 2889 2882 2893
rect 2894 2890 2898 2894
rect 2921 2890 2925 2894
rect 2969 2889 2975 2893
rect 3050 2889 3056 2893
rect 3356 2900 3360 2904
rect 3391 2905 3395 2909
rect 3375 2896 3379 2903
rect 3433 2896 3437 2903
rect 3451 2905 3455 2909
rect 3733 2907 3737 2911
rect 3777 2908 3781 2912
rect 3469 2903 3473 2907
rect 3802 2907 3807 2911
rect 3849 2908 3853 2912
rect 3925 2905 3929 2909
rect 4006 2905 4010 2909
rect 3716 2890 3720 2894
rect 3370 2880 3374 2884
rect 3406 2880 3410 2884
rect 3426 2880 3430 2884
rect 3463 2882 3467 2886
rect 3748 2889 3752 2893
rect 3767 2890 3771 2894
rect 3823 2889 3827 2893
rect 3839 2890 3843 2894
rect 3866 2890 3870 2894
rect 3914 2889 3920 2893
rect 3995 2889 4001 2893
rect 2791 2870 2795 2874
rect 2835 2870 2839 2874
rect 2862 2870 2866 2874
rect 2907 2870 2911 2874
rect 2978 2869 2982 2873
rect 3059 2869 3063 2873
rect 3736 2870 3740 2874
rect 3780 2870 3784 2874
rect 3807 2870 3811 2874
rect 3852 2870 3856 2874
rect 3923 2869 3927 2873
rect 4004 2869 4008 2873
rect 2980 2849 2984 2853
rect 2791 2842 2795 2846
rect 2835 2842 2839 2846
rect 2862 2842 2866 2846
rect 2907 2842 2911 2846
rect 3085 2849 3089 2853
rect 2972 2831 2976 2835
rect 2771 2822 2775 2826
rect 2803 2823 2807 2827
rect 2822 2822 2826 2826
rect 2878 2823 2882 2827
rect 2894 2822 2898 2826
rect 2921 2822 2925 2826
rect 2999 2827 3003 2831
rect 3050 2835 3054 2839
rect 3925 2849 3929 2853
rect 3077 2831 3081 2835
rect 3104 2827 3108 2831
rect 3736 2842 3740 2846
rect 3780 2842 3784 2846
rect 3807 2842 3811 2846
rect 3852 2842 3856 2846
rect 4030 2849 4034 2853
rect 3917 2831 3921 2835
rect 3716 2822 3720 2826
rect 2978 2813 2982 2817
rect 3083 2813 3087 2817
rect 3748 2823 3752 2827
rect 3767 2822 3771 2826
rect 3823 2823 3827 2827
rect 3839 2822 3843 2826
rect 3866 2822 3870 2826
rect 3944 2827 3948 2831
rect 3995 2835 3999 2839
rect 4022 2831 4026 2835
rect 4049 2827 4053 2831
rect 3923 2813 3927 2817
rect 4028 2813 4032 2817
rect 2788 2805 2792 2809
rect 2832 2804 2836 2808
rect 2857 2805 2862 2809
rect 2904 2804 2908 2808
rect 3733 2805 3737 2809
rect 3777 2804 3781 2808
rect 3802 2805 3807 2809
rect 3849 2804 3853 2808
rect 2788 2775 2792 2779
rect 2832 2776 2836 2780
rect 2857 2775 2862 2779
rect 2904 2776 2908 2780
rect 2980 2774 2984 2778
rect 3085 2774 3089 2778
rect 3733 2775 3737 2779
rect 3777 2776 3781 2780
rect 3802 2775 3807 2779
rect 3849 2776 3853 2780
rect 3925 2774 3929 2778
rect 4030 2774 4034 2778
rect 2771 2758 2775 2762
rect 2803 2757 2807 2761
rect 2822 2758 2826 2762
rect 2878 2757 2882 2761
rect 2894 2758 2898 2762
rect 2921 2758 2925 2762
rect 2969 2758 2975 2762
rect 3074 2758 3080 2762
rect 3716 2758 3720 2762
rect 3748 2757 3752 2761
rect 3767 2758 3771 2762
rect 3823 2757 3827 2761
rect 3839 2758 3843 2762
rect 3866 2758 3870 2762
rect 3914 2758 3920 2762
rect 4019 2758 4025 2762
rect 2791 2738 2795 2742
rect 2835 2738 2839 2742
rect 2862 2738 2866 2742
rect 2907 2738 2911 2742
rect 2978 2738 2982 2742
rect 3083 2738 3087 2742
rect 3736 2738 3740 2742
rect 3780 2738 3784 2742
rect 3807 2738 3811 2742
rect 3852 2738 3856 2742
rect 3923 2738 3927 2742
rect 4028 2738 4032 2742
rect 2980 2717 2984 2721
rect 2791 2710 2795 2714
rect 2835 2710 2839 2714
rect 2862 2710 2866 2714
rect 2907 2710 2911 2714
rect 3061 2717 3065 2721
rect 2972 2699 2976 2703
rect 2771 2690 2775 2694
rect 2803 2691 2807 2695
rect 2822 2690 2826 2694
rect 2878 2691 2882 2695
rect 2894 2690 2898 2694
rect 2921 2690 2925 2694
rect 2999 2695 3003 2699
rect 3026 2703 3030 2707
rect 3151 2717 3155 2721
rect 3053 2699 3057 2703
rect 3080 2695 3084 2699
rect 3116 2703 3120 2707
rect 3925 2717 3929 2721
rect 3143 2699 3147 2703
rect 3170 2695 3174 2699
rect 3736 2710 3740 2714
rect 3780 2710 3784 2714
rect 3807 2710 3811 2714
rect 3852 2710 3856 2714
rect 4006 2717 4010 2721
rect 3917 2699 3921 2703
rect 3716 2690 3720 2694
rect 2978 2681 2982 2685
rect 3059 2681 3063 2685
rect 3149 2681 3153 2685
rect 3748 2691 3752 2695
rect 3767 2690 3771 2694
rect 3823 2691 3827 2695
rect 3839 2690 3843 2694
rect 3866 2690 3870 2694
rect 3944 2695 3948 2699
rect 3971 2703 3975 2707
rect 4096 2717 4100 2721
rect 3998 2699 4002 2703
rect 4025 2695 4029 2699
rect 4061 2703 4065 2707
rect 4088 2699 4092 2703
rect 4115 2695 4119 2699
rect 3923 2681 3927 2685
rect 4004 2681 4008 2685
rect 4094 2681 4098 2685
rect 2788 2673 2792 2677
rect 2832 2672 2836 2676
rect 2857 2673 2862 2677
rect 2904 2672 2908 2676
rect 3733 2673 3737 2677
rect 3777 2672 3781 2676
rect 3802 2673 3807 2677
rect 3849 2672 3853 2676
rect 2788 2643 2792 2647
rect 2832 2644 2836 2648
rect 2857 2643 2862 2647
rect 2904 2644 2908 2648
rect 3733 2643 3737 2647
rect 3777 2644 3781 2648
rect 2980 2639 2984 2643
rect 3061 2639 3065 2643
rect 3151 2639 3155 2643
rect 3802 2643 3807 2647
rect 3849 2644 3853 2648
rect 3925 2639 3929 2643
rect 4006 2639 4010 2643
rect 4096 2639 4100 2643
rect 2771 2626 2775 2630
rect 2803 2625 2807 2629
rect 2822 2626 2826 2630
rect 2878 2625 2882 2629
rect 2894 2626 2898 2630
rect 2921 2626 2925 2630
rect 2969 2623 2975 2627
rect 3050 2623 3056 2627
rect 3140 2623 3146 2627
rect 3716 2626 3720 2630
rect 3748 2625 3752 2629
rect 3767 2626 3771 2630
rect 3823 2625 3827 2629
rect 3839 2626 3843 2630
rect 3866 2626 3870 2630
rect 3914 2623 3920 2627
rect 3995 2623 4001 2627
rect 4085 2623 4091 2627
rect 2791 2606 2795 2610
rect 2835 2606 2839 2610
rect 2862 2606 2866 2610
rect 2907 2606 2911 2610
rect 2978 2603 2982 2607
rect 3059 2603 3063 2607
rect 3149 2603 3153 2607
rect 3736 2606 3740 2610
rect 3780 2606 3784 2610
rect 3807 2606 3811 2610
rect 3852 2606 3856 2610
rect 3923 2603 3927 2607
rect 4004 2603 4008 2607
rect 4094 2603 4098 2607
rect 2980 2585 2984 2589
rect 2791 2578 2795 2582
rect 2835 2578 2839 2582
rect 2862 2578 2866 2582
rect 2907 2578 2911 2582
rect 3925 2585 3929 2589
rect 2972 2567 2976 2571
rect 2771 2558 2775 2562
rect 2803 2559 2807 2563
rect 2822 2558 2826 2562
rect 2878 2559 2882 2563
rect 2894 2558 2898 2562
rect 2921 2558 2925 2562
rect 2999 2563 3003 2567
rect 3736 2578 3740 2582
rect 3780 2578 3784 2582
rect 3807 2578 3811 2582
rect 3852 2578 3856 2582
rect 3917 2567 3921 2571
rect 3716 2558 3720 2562
rect 2978 2549 2982 2553
rect 3748 2559 3752 2563
rect 3767 2558 3771 2562
rect 3823 2559 3827 2563
rect 3839 2558 3843 2562
rect 3866 2558 3870 2562
rect 3944 2563 3948 2567
rect 3923 2549 3927 2553
rect 2788 2541 2792 2545
rect 2832 2540 2836 2544
rect 2857 2541 2862 2545
rect 2904 2540 2908 2544
rect 3733 2541 3737 2545
rect 3777 2540 3781 2544
rect 3802 2541 3807 2545
rect 3849 2540 3853 2544
rect 2291 2523 2295 2527
rect 2328 2523 2332 2527
rect 2348 2523 2352 2527
rect 2386 2523 2390 2527
rect 2423 2523 2427 2527
rect 2460 2523 2464 2527
rect 2480 2523 2484 2527
rect 2518 2523 2522 2527
rect 2555 2523 2559 2527
rect 2592 2523 2596 2527
rect 2612 2523 2616 2527
rect 2650 2523 2654 2527
rect 3236 2523 3240 2527
rect 3273 2523 3277 2527
rect 3293 2523 3297 2527
rect 3331 2523 3335 2527
rect 3368 2523 3372 2527
rect 3405 2523 3409 2527
rect 3425 2523 3429 2527
rect 3463 2523 3467 2527
rect 3500 2523 3504 2527
rect 3537 2523 3541 2527
rect 3557 2523 3561 2527
rect 3595 2523 3599 2527
rect 2285 2503 2289 2507
rect 2303 2505 2307 2509
rect 2363 2505 2367 2509
rect 2321 2496 2325 2503
rect 2379 2496 2383 2503
rect 2398 2500 2402 2504
rect 2416 2505 2420 2509
rect 2435 2505 2439 2509
rect 2495 2505 2499 2509
rect 2453 2496 2457 2503
rect 2511 2496 2515 2503
rect 2530 2500 2534 2504
rect 2548 2505 2552 2509
rect 2567 2505 2571 2509
rect 2627 2505 2631 2509
rect 2585 2496 2589 2503
rect 2788 2511 2792 2515
rect 2832 2512 2836 2516
rect 2857 2511 2862 2515
rect 2904 2512 2908 2516
rect 3049 2511 3053 2515
rect 3093 2512 3097 2516
rect 3118 2511 3123 2515
rect 3165 2512 3169 2516
rect 2643 2496 2647 2503
rect 2664 2500 2668 2504
rect 2980 2503 2984 2507
rect 3230 2503 3234 2507
rect 3248 2505 3252 2509
rect 2771 2494 2775 2498
rect 2803 2493 2807 2497
rect 2822 2494 2826 2498
rect 2878 2493 2882 2497
rect 2894 2494 2898 2498
rect 2921 2494 2925 2498
rect 2291 2482 2295 2486
rect 2328 2480 2332 2484
rect 2348 2480 2352 2484
rect 2384 2480 2388 2484
rect 2423 2482 2427 2486
rect 2460 2480 2464 2484
rect 2480 2480 2484 2484
rect 2516 2480 2520 2484
rect 2555 2482 2559 2486
rect 2592 2480 2596 2484
rect 2612 2480 2616 2484
rect 2648 2480 2652 2484
rect 2969 2487 2975 2491
rect 3007 2494 3011 2498
rect 3064 2493 3068 2497
rect 3083 2494 3087 2498
rect 3139 2493 3143 2497
rect 3155 2494 3159 2498
rect 3182 2494 3186 2498
rect 3308 2505 3312 2509
rect 3266 2496 3270 2503
rect 3324 2496 3328 2503
rect 3343 2500 3347 2504
rect 3361 2505 3365 2509
rect 3380 2505 3384 2509
rect 3440 2505 3444 2509
rect 3398 2496 3402 2503
rect 3456 2496 3460 2503
rect 3475 2500 3479 2504
rect 3493 2505 3497 2509
rect 3512 2505 3516 2509
rect 3572 2505 3576 2509
rect 3530 2496 3534 2503
rect 3733 2511 3737 2515
rect 3777 2512 3781 2516
rect 3802 2511 3807 2515
rect 3849 2512 3853 2516
rect 3994 2511 3998 2515
rect 4038 2512 4042 2516
rect 4063 2511 4068 2515
rect 4110 2512 4114 2516
rect 3588 2496 3592 2503
rect 3609 2500 3613 2504
rect 3925 2503 3929 2507
rect 3716 2494 3720 2498
rect 3748 2493 3752 2497
rect 3767 2494 3771 2498
rect 3823 2493 3827 2497
rect 3839 2494 3843 2498
rect 3866 2494 3870 2498
rect 2791 2474 2795 2478
rect 2835 2474 2839 2478
rect 2862 2474 2866 2478
rect 2907 2474 2911 2478
rect 3236 2482 3240 2486
rect 2978 2467 2982 2471
rect 2400 2452 2404 2456
rect 2424 2452 2428 2456
rect 3273 2480 3277 2484
rect 3293 2480 3297 2484
rect 3329 2480 3333 2484
rect 3368 2482 3372 2486
rect 3405 2480 3409 2484
rect 3425 2480 3429 2484
rect 3461 2480 3465 2484
rect 3500 2482 3504 2486
rect 3537 2480 3541 2484
rect 3557 2480 3561 2484
rect 3593 2480 3597 2484
rect 3914 2487 3920 2491
rect 3952 2494 3956 2498
rect 4009 2493 4013 2497
rect 4028 2494 4032 2498
rect 4084 2493 4088 2497
rect 4100 2494 4104 2498
rect 4127 2494 4131 2498
rect 3052 2474 3056 2478
rect 3096 2474 3100 2478
rect 3123 2474 3127 2478
rect 3168 2474 3172 2478
rect 3736 2474 3740 2478
rect 3780 2474 3784 2478
rect 3807 2474 3811 2478
rect 3852 2474 3856 2478
rect 3923 2467 3927 2471
rect 3345 2452 3349 2456
rect 3369 2452 3373 2456
rect 3191 2446 3195 2450
rect 3029 2439 3033 2443
rect 3997 2474 4001 2478
rect 4041 2474 4045 2478
rect 4068 2474 4072 2478
rect 4113 2474 4117 2478
rect 4136 2446 4140 2450
rect 3972 2439 3976 2443
rect 2420 2425 2424 2429
rect 3365 2425 3369 2429
rect 2435 2417 2439 2421
rect 3380 2417 3384 2421
rect 3074 2411 3078 2415
rect 3111 2411 3115 2415
rect 3131 2411 3135 2415
rect 3169 2411 3173 2415
rect 4019 2411 4023 2415
rect 4056 2411 4060 2415
rect 4076 2411 4080 2415
rect 4114 2411 4118 2415
rect 2400 2402 2404 2406
rect 2424 2402 2428 2406
rect 3345 2402 3349 2406
rect 3369 2402 3373 2406
rect 3068 2391 3072 2395
rect 3086 2393 3090 2397
rect 2291 2381 2295 2385
rect 2328 2381 2332 2385
rect 2348 2381 2352 2385
rect 2386 2381 2390 2385
rect 2423 2381 2427 2385
rect 2460 2381 2464 2385
rect 2480 2381 2484 2385
rect 2518 2381 2522 2385
rect 2555 2381 2559 2385
rect 2592 2381 2596 2385
rect 2612 2381 2616 2385
rect 2650 2381 2654 2385
rect 3146 2393 3150 2397
rect 3104 2384 3108 2391
rect 3162 2384 3166 2391
rect 3181 2388 3185 2392
rect 4013 2391 4017 2395
rect 4031 2393 4035 2397
rect 3236 2381 3240 2385
rect 3273 2381 3277 2385
rect 3293 2381 3297 2385
rect 3331 2381 3335 2385
rect 3368 2381 3372 2385
rect 3405 2381 3409 2385
rect 3425 2381 3429 2385
rect 3463 2381 3467 2385
rect 3500 2381 3504 2385
rect 3537 2381 3541 2385
rect 3557 2381 3561 2385
rect 3595 2381 3599 2385
rect 4091 2393 4095 2397
rect 4049 2384 4053 2391
rect 4107 2384 4111 2391
rect 4126 2388 4130 2392
rect 3074 2370 3078 2374
rect 2285 2361 2289 2365
rect 2303 2363 2307 2367
rect 2363 2363 2367 2367
rect 2321 2354 2325 2361
rect 2379 2354 2383 2361
rect 2398 2358 2402 2362
rect 2416 2363 2420 2367
rect 2435 2363 2439 2367
rect 2495 2363 2499 2367
rect 2453 2354 2457 2361
rect 2511 2354 2515 2361
rect 2530 2358 2534 2362
rect 2548 2363 2552 2367
rect 2567 2363 2571 2367
rect 2627 2363 2631 2367
rect 2585 2354 2589 2361
rect 3111 2368 3115 2372
rect 3131 2368 3135 2372
rect 3167 2368 3171 2372
rect 4019 2370 4023 2374
rect 2643 2354 2647 2361
rect 2664 2358 2668 2362
rect 3230 2361 3234 2365
rect 3248 2363 3252 2367
rect 3308 2363 3312 2367
rect 3266 2354 3270 2361
rect 3324 2354 3328 2361
rect 3343 2358 3347 2362
rect 3361 2363 3365 2367
rect 3380 2363 3384 2367
rect 3440 2363 3444 2367
rect 3398 2354 3402 2361
rect 3456 2354 3460 2361
rect 3475 2358 3479 2362
rect 3493 2363 3497 2367
rect 3512 2363 3516 2367
rect 3572 2363 3576 2367
rect 3530 2354 3534 2361
rect 4056 2368 4060 2372
rect 4076 2368 4080 2372
rect 4112 2368 4116 2372
rect 3588 2354 3592 2361
rect 3609 2358 3613 2362
rect 2291 2340 2295 2344
rect 2328 2338 2332 2342
rect 2348 2338 2352 2342
rect 2384 2338 2388 2342
rect 2423 2340 2427 2344
rect 2460 2338 2464 2342
rect 2480 2338 2484 2342
rect 2516 2338 2520 2342
rect 2555 2340 2559 2344
rect 2592 2338 2596 2342
rect 2612 2338 2616 2342
rect 2648 2338 2652 2342
rect 3236 2340 3240 2344
rect 3273 2338 3277 2342
rect 3293 2338 3297 2342
rect 3329 2338 3333 2342
rect 3368 2340 3372 2344
rect 3405 2338 3409 2342
rect 3425 2338 3429 2342
rect 3461 2338 3465 2342
rect 3500 2340 3504 2344
rect 3537 2338 3541 2342
rect 3557 2338 3561 2342
rect 3593 2338 3597 2342
rect 3074 2325 3078 2329
rect 3111 2325 3115 2329
rect 3131 2325 3135 2329
rect 3169 2325 3173 2329
rect 4019 2325 4023 2329
rect 4056 2325 4060 2329
rect 4076 2325 4080 2329
rect 4114 2325 4118 2329
rect 3068 2305 3072 2309
rect 3086 2307 3090 2311
rect 2291 2295 2295 2299
rect 2328 2295 2332 2299
rect 2348 2295 2352 2299
rect 2386 2295 2390 2299
rect 2423 2295 2427 2299
rect 2460 2295 2464 2299
rect 2480 2295 2484 2299
rect 2518 2295 2522 2299
rect 2555 2295 2559 2299
rect 2592 2295 2596 2299
rect 2612 2295 2616 2299
rect 2650 2295 2654 2299
rect 3146 2307 3150 2311
rect 3104 2298 3108 2305
rect 3162 2298 3166 2305
rect 3181 2302 3185 2306
rect 3203 2300 3207 2304
rect 4013 2305 4017 2309
rect 4031 2307 4035 2311
rect 3236 2295 3240 2299
rect 3273 2295 3277 2299
rect 3293 2295 3297 2299
rect 3331 2295 3335 2299
rect 3368 2295 3372 2299
rect 3405 2295 3409 2299
rect 3425 2295 3429 2299
rect 3463 2295 3467 2299
rect 3500 2295 3504 2299
rect 3537 2295 3541 2299
rect 3557 2295 3561 2299
rect 3595 2295 3599 2299
rect 4091 2307 4095 2311
rect 4049 2298 4053 2305
rect 4107 2298 4111 2305
rect 4126 2302 4130 2306
rect 4148 2300 4152 2304
rect 3074 2284 3078 2288
rect 2285 2275 2289 2279
rect 2303 2277 2307 2281
rect 2363 2277 2367 2281
rect 2321 2268 2325 2275
rect 2379 2268 2383 2275
rect 2398 2272 2402 2276
rect 2416 2277 2420 2281
rect 2435 2277 2439 2281
rect 2495 2277 2499 2281
rect 2453 2268 2457 2275
rect 2511 2268 2515 2275
rect 2530 2272 2534 2276
rect 2548 2277 2552 2281
rect 2567 2277 2571 2281
rect 2627 2277 2631 2281
rect 2585 2268 2589 2275
rect 3111 2282 3115 2286
rect 3131 2282 3135 2286
rect 3167 2282 3171 2286
rect 4019 2284 4023 2288
rect 2643 2268 2647 2275
rect 2664 2272 2668 2276
rect 3230 2275 3234 2279
rect 3248 2277 3252 2281
rect 3308 2277 3312 2281
rect 3266 2268 3270 2275
rect 3324 2268 3328 2275
rect 3343 2272 3347 2276
rect 3361 2277 3365 2281
rect 3380 2277 3384 2281
rect 3440 2277 3444 2281
rect 3398 2268 3402 2275
rect 3456 2268 3460 2275
rect 3475 2272 3479 2276
rect 3493 2277 3497 2281
rect 3512 2277 3516 2281
rect 3572 2277 3576 2281
rect 3530 2268 3534 2275
rect 4056 2282 4060 2286
rect 4076 2282 4080 2286
rect 4112 2282 4116 2286
rect 3588 2268 3592 2275
rect 3609 2272 3613 2276
rect 2291 2254 2295 2258
rect 2328 2252 2332 2256
rect 2348 2252 2352 2256
rect 2384 2252 2388 2256
rect 2423 2254 2427 2258
rect 2460 2252 2464 2256
rect 2480 2252 2484 2256
rect 2516 2252 2520 2256
rect 2555 2254 2559 2258
rect 2592 2252 2596 2256
rect 2612 2252 2616 2256
rect 2648 2252 2652 2256
rect 3236 2254 3240 2258
rect 3273 2252 3277 2256
rect 3293 2252 3297 2256
rect 3329 2252 3333 2256
rect 3368 2254 3372 2258
rect 3405 2252 3409 2256
rect 3425 2252 3429 2256
rect 3461 2252 3465 2256
rect 3500 2254 3504 2258
rect 3537 2252 3541 2256
rect 3557 2252 3561 2256
rect 3593 2252 3597 2256
rect 2517 2224 2521 2228
rect 2541 2224 2545 2228
rect 3462 2224 3466 2228
rect 3486 2224 3490 2228
rect 2537 2199 2541 2203
rect 3482 2199 3486 2203
rect 2552 2191 2556 2195
rect 3497 2191 3501 2195
rect 2517 2176 2521 2180
rect 2541 2176 2545 2180
rect 3462 2176 3466 2180
rect 3486 2176 3490 2180
rect 2291 2155 2295 2159
rect 2328 2155 2332 2159
rect 2348 2155 2352 2159
rect 2386 2155 2390 2159
rect 2423 2155 2427 2159
rect 2460 2155 2464 2159
rect 2480 2155 2484 2159
rect 2518 2155 2522 2159
rect 2555 2155 2559 2159
rect 2592 2155 2596 2159
rect 2612 2155 2616 2159
rect 2650 2155 2654 2159
rect 3236 2155 3240 2159
rect 3273 2155 3277 2159
rect 3293 2155 3297 2159
rect 3331 2155 3335 2159
rect 3368 2155 3372 2159
rect 3405 2155 3409 2159
rect 3425 2155 3429 2159
rect 3463 2155 3467 2159
rect 3500 2155 3504 2159
rect 3537 2155 3541 2159
rect 3557 2155 3561 2159
rect 3595 2155 3599 2159
rect 2285 2135 2289 2139
rect 2303 2137 2307 2141
rect 2363 2137 2367 2141
rect 2321 2128 2325 2135
rect 2379 2128 2383 2135
rect 2398 2132 2402 2136
rect 2416 2137 2420 2141
rect 2435 2137 2439 2141
rect 2495 2137 2499 2141
rect 2453 2128 2457 2135
rect 2511 2128 2515 2135
rect 2530 2132 2534 2136
rect 2548 2137 2552 2141
rect 2567 2137 2571 2141
rect 2627 2137 2631 2141
rect 2585 2128 2589 2135
rect 2643 2128 2647 2135
rect 2664 2132 2668 2136
rect 3230 2135 3234 2139
rect 3248 2137 3252 2141
rect 3308 2137 3312 2141
rect 3266 2128 3270 2135
rect 3324 2128 3328 2135
rect 3343 2132 3347 2136
rect 3361 2137 3365 2141
rect 3380 2137 3384 2141
rect 3440 2137 3444 2141
rect 3398 2128 3402 2135
rect 3456 2128 3460 2135
rect 3475 2132 3479 2136
rect 3493 2137 3497 2141
rect 3512 2137 3516 2141
rect 3572 2137 3576 2141
rect 3530 2128 3534 2135
rect 3588 2128 3592 2135
rect 3609 2132 3613 2136
rect 2291 2114 2295 2118
rect 2328 2112 2332 2116
rect 2348 2112 2352 2116
rect 2384 2112 2388 2116
rect 2423 2114 2427 2118
rect 2460 2112 2464 2116
rect 2480 2112 2484 2116
rect 2516 2112 2520 2116
rect 2555 2114 2559 2118
rect 2592 2112 2596 2116
rect 2612 2112 2616 2116
rect 2648 2112 2652 2116
rect 3236 2114 3240 2118
rect 3273 2112 3277 2116
rect 3293 2112 3297 2116
rect 3329 2112 3333 2116
rect 3368 2114 3372 2118
rect 3405 2112 3409 2116
rect 3425 2112 3429 2116
rect 3461 2112 3465 2116
rect 3500 2114 3504 2118
rect 3537 2112 3541 2116
rect 3557 2112 3561 2116
rect 3593 2112 3597 2116
<< metal1 >>
rect 1376 4845 1460 4930
rect 1679 4820 1757 4909
rect 1986 4825 2064 4914
rect 2303 4825 2381 4914
rect 2614 4827 2692 4916
rect 2918 4817 2996 4906
rect 3232 4825 3310 4914
rect 3522 4810 3634 4924
rect 1718 4300 1731 4326
rect 2027 4304 2040 4326
rect 2336 4304 2349 4354
rect 2645 4316 2658 4338
rect 2954 4318 2967 4338
rect 3263 4318 3276 4338
rect 2645 4312 2935 4316
rect 3548 4316 3604 4336
rect 2645 4311 2911 4312
rect 2349 4282 2411 4304
rect 3881 4281 3894 4328
rect 2048 4256 2315 4278
rect 2328 4256 2390 4278
rect 2048 4254 2330 4256
rect 2744 4204 3683 4208
rect 2732 4196 3671 4200
rect 2720 4189 3659 4193
rect 2708 4182 3647 4186
rect 2696 4174 3241 4178
rect 3296 4174 3635 4178
rect 3641 4174 3702 4178
rect 3606 4170 3623 4171
rect 2684 4166 3549 4170
rect 3604 4167 3623 4170
rect 3629 4167 3702 4171
rect 3604 4166 3612 4167
rect 3882 4163 3894 4281
rect 2756 4159 3695 4163
rect 3701 4159 3894 4163
rect 2967 4151 3337 4155
rect 2940 4141 3325 4145
rect 2744 4054 2771 4058
rect 2775 4054 2807 4058
rect 2811 4054 2874 4058
rect 2878 4054 2903 4058
rect 2907 4054 2939 4058
rect 2943 4054 3006 4058
rect 3010 4054 3035 4058
rect 3039 4054 3071 4058
rect 3075 4054 3138 4058
rect 3142 4054 3167 4058
rect 3171 4054 3203 4058
rect 3207 4054 3270 4058
rect 3274 4054 3290 4058
rect 3689 4054 3716 4058
rect 3720 4054 3752 4058
rect 3756 4054 3819 4058
rect 3823 4054 3848 4058
rect 3852 4054 3884 4058
rect 3888 4054 3951 4058
rect 3955 4054 3980 4058
rect 3984 4054 4016 4058
rect 4020 4054 4083 4058
rect 4087 4054 4112 4058
rect 4116 4054 4148 4058
rect 4152 4054 4215 4058
rect 4219 4054 4235 4058
rect 2684 4047 2795 4051
rect 2799 4047 2823 4051
rect 2827 4047 2853 4051
rect 2857 4047 2890 4051
rect 2894 4047 2927 4051
rect 2931 4047 2955 4051
rect 2959 4047 2985 4051
rect 2989 4047 3022 4051
rect 3026 4047 3059 4051
rect 3063 4047 3087 4051
rect 3091 4047 3117 4051
rect 3121 4047 3154 4051
rect 3158 4047 3191 4051
rect 3195 4047 3219 4051
rect 3223 4047 3249 4051
rect 3253 4047 3286 4051
rect 3629 4047 3740 4051
rect 3744 4047 3768 4051
rect 3772 4047 3798 4051
rect 3802 4047 3835 4051
rect 3839 4047 3872 4051
rect 3876 4047 3900 4051
rect 3904 4047 3930 4051
rect 3934 4047 3967 4051
rect 3971 4047 4004 4051
rect 4008 4047 4032 4051
rect 4036 4047 4062 4051
rect 4066 4047 4099 4051
rect 4103 4047 4136 4051
rect 4140 4047 4164 4051
rect 4168 4047 4194 4051
rect 4198 4047 4231 4051
rect 2765 4037 2768 4047
rect 2786 4037 2789 4047
rect 2802 4037 2805 4047
rect 2816 4040 2821 4044
rect 2825 4040 2832 4044
rect 2844 4037 2847 4047
rect 2860 4037 2863 4047
rect 2881 4037 2884 4047
rect 2897 4037 2900 4047
rect 2918 4037 2921 4047
rect 2934 4037 2937 4047
rect 2948 4040 2953 4044
rect 2957 4040 2964 4044
rect 2976 4037 2979 4047
rect 2992 4037 2995 4047
rect 3013 4037 3016 4047
rect 3029 4037 3032 4047
rect 3050 4037 3053 4047
rect 3066 4037 3069 4047
rect 3080 4040 3085 4044
rect 3089 4040 3096 4044
rect 3108 4037 3111 4047
rect 3124 4037 3127 4047
rect 3145 4037 3148 4047
rect 3161 4037 3164 4047
rect 3182 4037 3185 4047
rect 3198 4037 3201 4047
rect 3212 4040 3217 4044
rect 3221 4040 3228 4044
rect 3240 4037 3243 4047
rect 3256 4037 3259 4047
rect 3277 4037 3280 4047
rect 3710 4037 3713 4047
rect 3731 4037 3734 4047
rect 3747 4037 3750 4047
rect 3761 4040 3766 4044
rect 3770 4040 3777 4044
rect 3789 4037 3792 4047
rect 3805 4037 3808 4047
rect 3826 4037 3829 4047
rect 3842 4037 3845 4047
rect 3863 4037 3866 4047
rect 3879 4037 3882 4047
rect 3893 4040 3898 4044
rect 3902 4040 3909 4044
rect 3921 4037 3924 4047
rect 3937 4037 3940 4047
rect 3958 4037 3961 4047
rect 3974 4037 3977 4047
rect 3995 4037 3998 4047
rect 4011 4037 4014 4047
rect 4025 4040 4030 4044
rect 4034 4040 4041 4044
rect 4053 4037 4056 4047
rect 4069 4037 4072 4047
rect 4090 4037 4093 4047
rect 4106 4037 4109 4047
rect 4127 4037 4130 4047
rect 4143 4037 4146 4047
rect 4157 4040 4162 4044
rect 4166 4040 4173 4044
rect 4185 4037 4188 4047
rect 4201 4037 4204 4047
rect 4222 4037 4225 4047
rect 2410 4021 2419 4025
rect 2423 4021 2455 4025
rect 2459 4021 2522 4025
rect 2526 4021 2738 4025
rect 2782 4023 2787 4026
rect 2791 4023 2815 4026
rect 2840 4023 2847 4026
rect 2851 4023 2873 4026
rect 2410 4014 2443 4018
rect 2447 4014 2471 4018
rect 2475 4014 2501 4018
rect 2505 4014 2538 4018
rect 2542 4014 2678 4018
rect 2413 4004 2416 4014
rect 2434 4004 2437 4014
rect 2450 4004 2453 4014
rect 2464 4007 2469 4011
rect 2473 4007 2480 4011
rect 2492 4004 2495 4014
rect 2508 4004 2511 4014
rect 2529 4004 2532 4014
rect 2798 4013 2805 4016
rect 2809 4017 2828 4020
rect 2828 4010 2831 4016
rect 2856 4013 2863 4016
rect 2867 4017 2884 4020
rect 2914 4023 2919 4026
rect 2923 4023 2947 4026
rect 2972 4023 2979 4026
rect 2983 4023 3005 4026
rect 2930 4013 2937 4016
rect 2941 4017 2960 4020
rect 2960 4010 2963 4016
rect 2988 4013 2995 4016
rect 2999 4017 3016 4020
rect 3046 4023 3051 4026
rect 3055 4023 3079 4026
rect 3104 4023 3111 4026
rect 3115 4023 3137 4026
rect 3062 4013 3069 4016
rect 3073 4017 3092 4020
rect 3092 4010 3095 4016
rect 3120 4013 3127 4016
rect 3131 4017 3148 4020
rect 3178 4023 3183 4026
rect 3187 4023 3211 4026
rect 3236 4023 3243 4026
rect 3247 4023 3269 4026
rect 3355 4021 3364 4025
rect 3368 4021 3400 4025
rect 3404 4021 3467 4025
rect 3471 4021 3683 4025
rect 3194 4013 3201 4016
rect 3205 4017 3224 4020
rect 2408 3987 2417 3991
rect 2430 3990 2435 3993
rect 2439 3990 2463 3993
rect 2488 3990 2495 3993
rect 2499 3990 2521 3993
rect 2765 3994 2768 4006
rect 2786 3994 2789 4006
rect 2802 3994 2805 4006
rect 2816 3997 2828 4000
rect 2844 3994 2847 4006
rect 2860 3994 2863 4006
rect 2881 3994 2884 4006
rect 2897 3994 2900 4006
rect 2918 3994 2921 4006
rect 2934 3994 2937 4006
rect 2948 3997 2960 4000
rect 2976 3994 2979 4006
rect 2992 3994 2995 4006
rect 3013 3994 3016 4006
rect 3029 3994 3032 4006
rect 3050 3994 3053 4006
rect 3066 3994 3069 4006
rect 3080 3997 3092 4000
rect 3108 3994 3111 4006
rect 3124 3994 3127 4006
rect 3145 3994 3148 4006
rect 3224 4010 3227 4016
rect 3252 4013 3259 4016
rect 3263 4017 3280 4020
rect 3727 4023 3732 4026
rect 3736 4023 3760 4026
rect 3785 4023 3792 4026
rect 3796 4023 3818 4026
rect 3355 4014 3388 4018
rect 3392 4014 3416 4018
rect 3420 4014 3446 4018
rect 3450 4014 3483 4018
rect 3487 4014 3623 4018
rect 3161 3994 3164 4006
rect 3182 3994 3185 4006
rect 3198 3994 3201 4006
rect 3212 3997 3224 4000
rect 3240 3994 3243 4006
rect 3256 3994 3259 4006
rect 3277 3994 3280 4006
rect 3358 4004 3361 4014
rect 3379 4004 3382 4014
rect 3395 4004 3398 4014
rect 3409 4007 3414 4011
rect 3418 4007 3425 4011
rect 3437 4004 3440 4014
rect 3453 4004 3456 4014
rect 3474 4004 3477 4014
rect 3743 4013 3750 4016
rect 3754 4017 3773 4020
rect 3773 4010 3776 4016
rect 3801 4013 3808 4016
rect 3812 4017 3829 4020
rect 3859 4023 3864 4026
rect 3868 4023 3892 4026
rect 3917 4023 3924 4026
rect 3928 4023 3950 4026
rect 3875 4013 3882 4016
rect 3886 4017 3905 4020
rect 3905 4010 3908 4016
rect 3933 4013 3940 4016
rect 3944 4017 3961 4020
rect 3991 4023 3996 4026
rect 4000 4023 4024 4026
rect 4049 4023 4056 4026
rect 4060 4023 4082 4026
rect 4007 4013 4014 4016
rect 4018 4017 4037 4020
rect 4037 4010 4040 4016
rect 4065 4013 4072 4016
rect 4076 4017 4093 4020
rect 4123 4023 4128 4026
rect 4132 4023 4156 4026
rect 4181 4023 4188 4026
rect 4192 4023 4214 4026
rect 4139 4013 4146 4016
rect 4150 4017 4169 4020
rect 2696 3990 2795 3994
rect 2799 3990 2823 3994
rect 2827 3990 2853 3994
rect 2857 3990 2927 3994
rect 2931 3990 2955 3994
rect 2959 3990 2985 3994
rect 2989 3990 3059 3994
rect 3063 3990 3087 3994
rect 3091 3990 3117 3994
rect 3121 3990 3191 3994
rect 3195 3990 3219 3994
rect 3223 3990 3249 3994
rect 3253 3990 3290 3994
rect 2446 3980 2453 3983
rect 2457 3984 2476 3987
rect 2476 3977 2479 3983
rect 2504 3980 2511 3983
rect 2515 3984 2530 3987
rect 3353 3987 3362 3991
rect 3375 3990 3380 3993
rect 3384 3990 3408 3993
rect 3433 3990 3440 3993
rect 3444 3990 3466 3993
rect 3710 3994 3713 4006
rect 3731 3994 3734 4006
rect 3747 3994 3750 4006
rect 3761 3997 3773 4000
rect 3789 3994 3792 4006
rect 3805 3994 3808 4006
rect 3826 3994 3829 4006
rect 3842 3994 3845 4006
rect 3863 3994 3866 4006
rect 3879 3994 3882 4006
rect 3893 3997 3905 4000
rect 3921 3994 3924 4006
rect 3937 3994 3940 4006
rect 3958 3994 3961 4006
rect 3974 3994 3977 4006
rect 3995 3994 3998 4006
rect 4011 3994 4014 4006
rect 4025 3997 4037 4000
rect 4053 3994 4056 4006
rect 4069 3994 4072 4006
rect 4090 3994 4093 4006
rect 4169 4010 4172 4016
rect 4197 4013 4204 4016
rect 4208 4017 4225 4020
rect 4106 3994 4109 4006
rect 4127 3994 4130 4006
rect 4143 3994 4146 4006
rect 4157 3997 4169 4000
rect 4185 3994 4188 4006
rect 4201 3994 4204 4006
rect 4222 3994 4225 4006
rect 3641 3990 3740 3994
rect 3744 3990 3768 3994
rect 3772 3990 3798 3994
rect 3802 3990 3872 3994
rect 3876 3990 3900 3994
rect 3904 3990 3930 3994
rect 3934 3990 4004 3994
rect 4008 3990 4032 3994
rect 4036 3990 4062 3994
rect 4066 3990 4136 3994
rect 4140 3990 4164 3994
rect 4168 3990 4194 3994
rect 4198 3990 4235 3994
rect 2732 3983 2771 3987
rect 2775 3983 2822 3987
rect 2826 3983 2872 3987
rect 2876 3983 2903 3987
rect 2907 3983 2954 3987
rect 2958 3983 3004 3987
rect 3008 3983 3035 3987
rect 3039 3983 3086 3987
rect 3090 3983 3136 3987
rect 3140 3983 3167 3987
rect 3171 3983 3218 3987
rect 3222 3983 3268 3987
rect 3272 3983 3290 3987
rect 3391 3980 3398 3983
rect 3402 3984 3421 3987
rect 2413 3961 2416 3973
rect 2434 3961 2437 3973
rect 2450 3961 2453 3973
rect 2464 3964 2476 3967
rect 2492 3961 2495 3973
rect 2508 3961 2511 3973
rect 2529 3961 2532 3973
rect 2684 3970 2769 3974
rect 2773 3970 2785 3974
rect 2789 3970 2803 3974
rect 2807 3970 2814 3974
rect 2818 3970 2820 3974
rect 2824 3970 2839 3974
rect 2843 3970 2876 3974
rect 2880 3970 2881 3974
rect 2885 3970 2893 3974
rect 2897 3970 2921 3974
rect 2925 3970 2937 3974
rect 2941 3970 2961 3974
rect 2965 3970 3015 3974
rect 3019 3970 3042 3974
rect 3046 3970 3096 3974
rect 3100 3970 3119 3974
rect 3421 3977 3424 3983
rect 3449 3980 3456 3983
rect 3460 3984 3475 3987
rect 3677 3983 3716 3987
rect 3720 3983 3767 3987
rect 3771 3983 3817 3987
rect 3821 3983 3848 3987
rect 3852 3983 3899 3987
rect 3903 3983 3949 3987
rect 3953 3983 3980 3987
rect 3984 3983 4031 3987
rect 4035 3983 4081 3987
rect 4085 3983 4112 3987
rect 4116 3983 4163 3987
rect 4167 3983 4213 3987
rect 4217 3983 4235 3987
rect 2720 3963 2796 3967
rect 2800 3963 2827 3967
rect 2831 3963 2849 3967
rect 2853 3963 2914 3967
rect 2918 3963 2932 3967
rect 2944 3966 2947 3970
rect 2410 3957 2443 3961
rect 2447 3957 2471 3961
rect 2475 3957 2501 3961
rect 2505 3957 2690 3961
rect 2410 3950 2419 3954
rect 2423 3950 2470 3954
rect 2474 3950 2520 3954
rect 2524 3950 2726 3954
rect 2839 3956 2842 3960
rect 2866 3956 2867 3960
rect 2911 3956 2913 3960
rect 2953 3953 2956 3958
rect 2968 3960 2971 3970
rect 2998 3966 3001 3970
rect 3025 3966 3028 3970
rect 2408 3934 2424 3938
rect 2533 3936 2537 3940
rect 2549 3936 2553 3940
rect 2557 3936 2771 3940
rect 2779 3939 2782 3945
rect 2786 3939 2789 3945
rect 2779 3936 2789 3939
rect 2779 3931 2782 3936
rect 2416 3927 2420 3931
rect 2432 3927 2553 3931
rect 2786 3931 2789 3936
rect 2795 3941 2798 3945
rect 2795 3937 2797 3941
rect 2801 3937 2803 3941
rect 2811 3940 2814 3945
rect 2839 3942 2842 3945
rect 2811 3938 2822 3940
rect 2795 3931 2798 3937
rect 2811 3936 2817 3938
rect 2811 3931 2814 3936
rect 2821 3936 2822 3938
rect 2840 3938 2842 3942
rect 2839 3931 2842 3938
rect 2942 3949 2945 3952
rect 2984 3949 2987 3952
rect 2855 3941 2858 3945
rect 2865 3941 2868 3945
rect 2865 3937 2874 3941
rect 2886 3940 2889 3945
rect 2911 3941 2914 3945
rect 2855 3931 2858 3937
rect 2865 3931 2868 3937
rect 2886 3936 2887 3940
rect 2891 3936 2894 3939
rect 2913 3937 2914 3941
rect 2929 3940 2932 3945
rect 2953 3944 2956 3949
rect 2961 3945 2972 3948
rect 2984 3946 2992 3949
rect 2886 3931 2889 3936
rect 2911 3931 2914 3937
rect 2929 3931 2932 3936
rect 2403 3919 2419 3923
rect 2423 3919 2486 3923
rect 2490 3919 2522 3923
rect 2526 3919 2738 3923
rect 2831 3918 2832 3922
rect 2856 3919 2857 3923
rect 2903 3918 2904 3922
rect 2407 3912 2440 3916
rect 2444 3912 2470 3916
rect 2474 3912 2498 3916
rect 2502 3912 2678 3916
rect 2413 3902 2416 3912
rect 2434 3902 2437 3912
rect 2450 3902 2453 3912
rect 2465 3905 2472 3909
rect 2476 3905 2481 3909
rect 2492 3902 2495 3912
rect 2508 3902 2511 3912
rect 2529 3902 2532 3912
rect 2708 3911 2784 3915
rect 2788 3911 2843 3915
rect 2847 3911 2868 3915
rect 2872 3911 2899 3915
rect 2903 3911 2932 3915
rect 2944 3908 2947 3940
rect 2961 3939 2964 3945
rect 2984 3940 2987 3946
rect 2996 3941 2999 3944
rect 3007 3944 3010 3958
rect 3034 3953 3037 3958
rect 3049 3960 3052 3970
rect 3079 3966 3082 3970
rect 3018 3949 3019 3952
rect 3023 3949 3026 3952
rect 3065 3949 3068 3952
rect 3007 3941 3015 3944
rect 3034 3944 3037 3949
rect 3007 3936 3010 3941
rect 3015 3937 3019 3941
rect 3042 3945 3053 3948
rect 3065 3946 3073 3949
rect 2959 3930 2964 3935
rect 2968 3908 2971 3936
rect 2998 3908 3001 3932
rect 3025 3908 3028 3940
rect 3042 3939 3045 3945
rect 3065 3940 3068 3946
rect 3077 3941 3080 3944
rect 3088 3944 3091 3958
rect 3242 3957 3325 3965
rect 3358 3961 3361 3973
rect 3379 3961 3382 3973
rect 3395 3961 3398 3973
rect 3409 3964 3421 3967
rect 3437 3961 3440 3973
rect 3453 3961 3456 3973
rect 3474 3961 3477 3973
rect 3629 3970 3714 3974
rect 3718 3970 3730 3974
rect 3734 3970 3748 3974
rect 3752 3970 3759 3974
rect 3763 3970 3765 3974
rect 3769 3970 3784 3974
rect 3788 3970 3821 3974
rect 3825 3970 3826 3974
rect 3830 3970 3838 3974
rect 3842 3970 3866 3974
rect 3870 3970 3882 3974
rect 3886 3970 3906 3974
rect 3910 3970 3960 3974
rect 3964 3970 3987 3974
rect 3991 3970 4041 3974
rect 4045 3970 4064 3974
rect 3665 3963 3741 3967
rect 3745 3963 3772 3967
rect 3776 3963 3794 3967
rect 3798 3963 3859 3967
rect 3863 3963 3877 3967
rect 3889 3966 3892 3970
rect 3355 3957 3388 3961
rect 3392 3957 3416 3961
rect 3420 3957 3446 3961
rect 3450 3957 3635 3961
rect 3279 3948 3337 3952
rect 3355 3950 3364 3954
rect 3368 3950 3415 3954
rect 3419 3950 3465 3954
rect 3469 3950 3671 3954
rect 3784 3956 3787 3960
rect 3811 3956 3812 3960
rect 3856 3956 3858 3960
rect 3898 3953 3901 3958
rect 3913 3960 3916 3970
rect 3943 3966 3946 3970
rect 3970 3966 3973 3970
rect 3088 3941 3100 3944
rect 3088 3936 3091 3941
rect 3040 3930 3045 3935
rect 3049 3908 3052 3936
rect 3353 3934 3369 3938
rect 3478 3936 3482 3940
rect 3494 3936 3498 3940
rect 3502 3936 3707 3940
rect 3711 3936 3716 3940
rect 3724 3939 3727 3945
rect 3731 3939 3734 3945
rect 3724 3936 3734 3939
rect 3079 3908 3082 3932
rect 3724 3931 3727 3936
rect 3361 3927 3365 3931
rect 3377 3927 3498 3931
rect 3731 3931 3734 3936
rect 3740 3941 3743 3945
rect 3740 3937 3742 3941
rect 3746 3937 3748 3941
rect 3756 3940 3759 3945
rect 3784 3942 3787 3945
rect 3756 3938 3767 3940
rect 3740 3931 3743 3937
rect 3756 3936 3762 3938
rect 3756 3931 3759 3936
rect 3766 3936 3767 3938
rect 3785 3938 3787 3942
rect 3784 3931 3787 3938
rect 3887 3949 3890 3952
rect 3929 3949 3932 3952
rect 3800 3941 3803 3945
rect 3810 3941 3813 3945
rect 3810 3937 3819 3941
rect 3831 3940 3834 3945
rect 3856 3941 3859 3945
rect 3800 3931 3803 3937
rect 3810 3931 3813 3937
rect 3831 3936 3832 3940
rect 3836 3936 3839 3939
rect 3858 3937 3859 3941
rect 3874 3940 3877 3945
rect 3898 3944 3901 3949
rect 3906 3945 3917 3948
rect 3929 3946 3937 3949
rect 3831 3931 3834 3936
rect 3856 3931 3859 3937
rect 3874 3931 3877 3936
rect 3348 3919 3364 3923
rect 3368 3919 3431 3923
rect 3435 3919 3467 3923
rect 3471 3919 3683 3923
rect 3776 3918 3777 3922
rect 3801 3919 3802 3923
rect 3848 3918 3849 3922
rect 3352 3912 3385 3916
rect 3389 3912 3415 3916
rect 3419 3912 3443 3916
rect 3447 3912 3623 3916
rect 2696 3904 2770 3908
rect 2774 3904 2776 3908
rect 2780 3904 2784 3908
rect 2788 3904 2802 3908
rect 2806 3904 2811 3908
rect 2815 3904 2820 3908
rect 2824 3904 2843 3908
rect 2847 3904 2877 3908
rect 2881 3904 2892 3908
rect 2896 3904 2920 3908
rect 2924 3904 2937 3908
rect 2941 3904 2961 3908
rect 2965 3904 3015 3908
rect 3022 3904 3042 3908
rect 3046 3904 3096 3908
rect 2424 3888 2446 3891
rect 2450 3888 2457 3891
rect 2708 3897 2784 3901
rect 2788 3897 2843 3901
rect 2847 3897 2868 3901
rect 2872 3897 2899 3901
rect 2903 3897 2932 3901
rect 2482 3888 2506 3891
rect 2510 3888 2515 3891
rect 2831 3890 2832 3894
rect 2856 3889 2857 3893
rect 2903 3890 2904 3894
rect 2528 3885 2537 3889
rect 2415 3882 2430 3885
rect 2469 3882 2488 3885
rect 2434 3878 2441 3881
rect 2466 3875 2469 3881
rect 2492 3878 2499 3881
rect 2779 3876 2782 3881
rect 2786 3876 2789 3881
rect 2769 3873 2771 3876
rect 2779 3873 2789 3876
rect 2413 3859 2416 3871
rect 2434 3859 2437 3871
rect 2450 3859 2453 3871
rect 2469 3862 2481 3865
rect 2492 3859 2495 3871
rect 2508 3859 2511 3871
rect 2529 3859 2532 3871
rect 2779 3867 2782 3873
rect 2786 3867 2789 3873
rect 2795 3875 2798 3881
rect 2811 3876 2814 3881
rect 2795 3871 2797 3875
rect 2801 3871 2803 3875
rect 2811 3874 2817 3876
rect 2821 3874 2822 3876
rect 2811 3872 2822 3874
rect 2839 3874 2842 3881
rect 2795 3867 2798 3871
rect 2811 3867 2814 3872
rect 2840 3870 2842 3874
rect 2839 3867 2842 3870
rect 2855 3875 2858 3881
rect 2865 3875 2868 3881
rect 2886 3876 2889 3881
rect 2865 3871 2874 3875
rect 2886 3872 2887 3876
rect 2891 3873 2894 3876
rect 2911 3875 2914 3881
rect 2929 3876 2932 3881
rect 2968 3884 2971 3904
rect 3049 3884 3052 3904
rect 3358 3902 3361 3912
rect 3379 3902 3382 3912
rect 3395 3902 3398 3912
rect 3410 3905 3417 3909
rect 3421 3905 3426 3909
rect 3437 3902 3440 3912
rect 3453 3902 3456 3912
rect 3474 3902 3477 3912
rect 3653 3911 3729 3915
rect 3733 3911 3788 3915
rect 3792 3911 3813 3915
rect 3817 3911 3844 3915
rect 3848 3911 3877 3915
rect 3889 3908 3892 3940
rect 3906 3939 3909 3945
rect 3929 3940 3932 3946
rect 3941 3941 3944 3944
rect 3952 3944 3955 3958
rect 3979 3953 3982 3958
rect 3994 3960 3997 3970
rect 4024 3966 4027 3970
rect 3963 3949 3964 3952
rect 3968 3949 3971 3952
rect 4010 3949 4013 3952
rect 3952 3941 3960 3944
rect 3979 3944 3982 3949
rect 3952 3936 3955 3941
rect 3960 3937 3964 3941
rect 3987 3945 3998 3948
rect 4010 3946 4018 3949
rect 3904 3930 3909 3935
rect 3913 3908 3916 3936
rect 3943 3908 3946 3932
rect 3970 3908 3973 3940
rect 3987 3939 3990 3945
rect 4010 3940 4013 3946
rect 4022 3941 4025 3944
rect 4033 3944 4036 3958
rect 4033 3941 4045 3944
rect 4033 3936 4036 3941
rect 3985 3930 3990 3935
rect 3994 3908 3997 3936
rect 4024 3908 4027 3932
rect 3641 3904 3715 3908
rect 3719 3904 3721 3908
rect 3725 3904 3729 3908
rect 3733 3904 3747 3908
rect 3751 3904 3756 3908
rect 3760 3904 3765 3908
rect 3769 3904 3788 3908
rect 3792 3904 3822 3908
rect 3826 3904 3837 3908
rect 3841 3904 3865 3908
rect 3869 3904 3882 3908
rect 3886 3904 3906 3908
rect 3910 3904 3960 3908
rect 3967 3904 3987 3908
rect 3991 3904 4041 3908
rect 3369 3888 3391 3891
rect 3395 3888 3402 3891
rect 3653 3897 3729 3901
rect 3733 3897 3788 3901
rect 3792 3897 3813 3901
rect 3817 3897 3844 3901
rect 3848 3897 3877 3901
rect 3427 3888 3451 3891
rect 3455 3888 3460 3891
rect 3776 3890 3777 3894
rect 3801 3889 3802 3893
rect 3848 3890 3849 3894
rect 3473 3885 3482 3889
rect 3360 3882 3375 3885
rect 2855 3867 2858 3871
rect 2865 3867 2868 3871
rect 2886 3867 2889 3872
rect 2913 3871 2914 3875
rect 2911 3867 2914 3871
rect 2929 3867 2932 3872
rect 2959 3871 2964 3876
rect 2968 3872 2969 3875
rect 2984 3874 2987 3880
rect 2984 3871 2992 3874
rect 3039 3871 3044 3876
rect 3048 3872 3050 3875
rect 3065 3874 3068 3880
rect 3414 3882 3433 3885
rect 3379 3878 3386 3881
rect 3411 3875 3414 3881
rect 3065 3871 3073 3874
rect 3437 3878 3444 3881
rect 3724 3876 3727 3881
rect 3731 3876 3734 3881
rect 3714 3873 3716 3876
rect 3724 3873 3734 3876
rect 2984 3868 2987 3871
rect 3065 3868 3068 3871
rect 2403 3855 2440 3859
rect 2444 3855 2470 3859
rect 2474 3855 2498 3859
rect 2502 3855 2690 3859
rect 2839 3852 2842 3856
rect 2866 3852 2867 3856
rect 2911 3852 2913 3856
rect 2403 3848 2421 3852
rect 2425 3848 2471 3852
rect 2475 3848 2522 3852
rect 2526 3848 2726 3852
rect 2784 3845 2796 3849
rect 2800 3845 2827 3849
rect 2831 3845 2849 3849
rect 2853 3845 2914 3849
rect 2918 3845 2932 3849
rect 2968 3842 2971 3860
rect 3049 3842 3052 3860
rect 3358 3859 3361 3871
rect 3379 3859 3382 3871
rect 3395 3859 3398 3871
rect 3414 3862 3426 3865
rect 3437 3859 3440 3871
rect 3453 3859 3456 3871
rect 3474 3859 3477 3871
rect 3724 3867 3727 3873
rect 3731 3867 3734 3873
rect 3740 3875 3743 3881
rect 3756 3876 3759 3881
rect 3740 3871 3742 3875
rect 3746 3871 3748 3875
rect 3756 3874 3762 3876
rect 3766 3874 3767 3876
rect 3756 3872 3767 3874
rect 3784 3874 3787 3881
rect 3740 3867 3743 3871
rect 3756 3867 3759 3872
rect 3785 3870 3787 3874
rect 3784 3867 3787 3870
rect 3800 3875 3803 3881
rect 3810 3875 3813 3881
rect 3831 3876 3834 3881
rect 3810 3871 3819 3875
rect 3831 3872 3832 3876
rect 3836 3873 3839 3876
rect 3856 3875 3859 3881
rect 3874 3876 3877 3881
rect 3913 3884 3916 3904
rect 3994 3884 3997 3904
rect 3800 3867 3803 3871
rect 3810 3867 3813 3871
rect 3831 3867 3834 3872
rect 3858 3871 3859 3875
rect 3856 3867 3859 3871
rect 3874 3867 3877 3872
rect 3904 3871 3909 3876
rect 3913 3872 3914 3875
rect 3929 3874 3932 3880
rect 3929 3871 3937 3874
rect 3984 3871 3989 3876
rect 3993 3872 3995 3875
rect 4010 3874 4013 3880
rect 4010 3871 4018 3874
rect 3929 3868 3932 3871
rect 4010 3868 4013 3871
rect 3348 3855 3385 3859
rect 3389 3855 3415 3859
rect 3419 3855 3443 3859
rect 3447 3855 3635 3859
rect 3784 3852 3787 3856
rect 3811 3852 3812 3856
rect 3856 3852 3858 3856
rect 3348 3848 3366 3852
rect 3370 3848 3416 3852
rect 3420 3848 3467 3852
rect 3471 3848 3671 3852
rect 3729 3845 3741 3849
rect 3745 3845 3772 3849
rect 3776 3845 3794 3849
rect 3798 3845 3859 3849
rect 3863 3845 3877 3849
rect 3913 3842 3916 3860
rect 3994 3842 3997 3860
rect 2684 3838 2769 3842
rect 2773 3838 2785 3842
rect 2789 3838 2803 3842
rect 2807 3838 2814 3842
rect 2818 3838 2820 3842
rect 2824 3838 2839 3842
rect 2843 3838 2876 3842
rect 2880 3838 2881 3842
rect 2885 3838 2893 3842
rect 2897 3838 2921 3842
rect 2925 3838 2937 3842
rect 2941 3838 2961 3842
rect 2965 3838 3015 3842
rect 3019 3838 3042 3842
rect 3046 3838 3104 3842
rect 3108 3838 3119 3842
rect 3629 3838 3714 3842
rect 3718 3838 3730 3842
rect 3734 3838 3748 3842
rect 3752 3838 3759 3842
rect 3763 3838 3765 3842
rect 3769 3838 3784 3842
rect 3788 3838 3821 3842
rect 3825 3838 3826 3842
rect 3830 3838 3838 3842
rect 3842 3838 3866 3842
rect 3870 3838 3882 3842
rect 3886 3838 3906 3842
rect 3910 3838 3960 3842
rect 3964 3838 3987 3842
rect 3991 3838 4049 3842
rect 4053 3838 4064 3842
rect 2720 3831 2780 3835
rect 2784 3831 2796 3835
rect 2800 3831 2827 3835
rect 2831 3831 2849 3835
rect 2853 3831 2914 3835
rect 2918 3831 2932 3835
rect 2968 3828 2971 3838
rect 2998 3834 3001 3838
rect 3049 3834 3052 3838
rect 2839 3824 2842 3828
rect 2866 3824 2867 3828
rect 2911 3824 2913 3828
rect 2768 3804 2771 3807
rect 2779 3807 2782 3813
rect 2786 3807 2789 3813
rect 2779 3804 2789 3807
rect 2779 3799 2782 3804
rect 2786 3799 2789 3804
rect 2795 3809 2798 3813
rect 2795 3805 2797 3809
rect 2801 3805 2803 3809
rect 2811 3808 2814 3813
rect 2839 3810 2842 3813
rect 2811 3806 2822 3808
rect 2795 3799 2798 3805
rect 2811 3804 2817 3806
rect 2811 3799 2814 3804
rect 2821 3804 2822 3806
rect 2840 3806 2842 3810
rect 2839 3799 2842 3806
rect 2984 3817 2987 3820
rect 2855 3809 2858 3813
rect 2865 3809 2868 3813
rect 2865 3805 2874 3809
rect 2886 3808 2889 3813
rect 2911 3809 2914 3813
rect 2855 3799 2858 3805
rect 2865 3799 2868 3805
rect 2886 3804 2887 3808
rect 2891 3804 2894 3807
rect 2913 3805 2914 3809
rect 2929 3808 2932 3813
rect 2961 3813 2972 3816
rect 2984 3814 2992 3817
rect 2886 3799 2889 3804
rect 2911 3799 2914 3805
rect 2961 3807 2964 3813
rect 2984 3808 2987 3814
rect 2996 3809 2999 3812
rect 3007 3812 3010 3826
rect 3058 3821 3061 3826
rect 3073 3828 3076 3838
rect 3103 3834 3106 3838
rect 3042 3817 3043 3820
rect 3047 3817 3050 3820
rect 3279 3827 3535 3832
rect 3665 3831 3725 3835
rect 3729 3831 3741 3835
rect 3745 3831 3772 3835
rect 3776 3831 3794 3835
rect 3798 3831 3859 3835
rect 3863 3831 3877 3835
rect 3913 3828 3916 3838
rect 3943 3834 3946 3838
rect 3994 3834 3997 3838
rect 3089 3817 3092 3820
rect 3015 3812 3020 3817
rect 3058 3812 3061 3817
rect 3007 3809 3015 3812
rect 2929 3799 2932 3804
rect 3007 3804 3010 3809
rect 3066 3813 3077 3816
rect 3089 3814 3097 3817
rect 2959 3798 2964 3803
rect 2831 3786 2832 3790
rect 2856 3787 2857 3791
rect 2903 3786 2904 3790
rect 2708 3779 2784 3783
rect 2788 3779 2843 3783
rect 2847 3779 2868 3783
rect 2872 3779 2899 3783
rect 2903 3779 2932 3783
rect 2968 3776 2971 3804
rect 2998 3776 3001 3800
rect 3049 3776 3052 3808
rect 3066 3807 3069 3813
rect 3089 3808 3092 3814
rect 3101 3809 3104 3812
rect 3112 3812 3115 3826
rect 3784 3824 3787 3828
rect 3811 3824 3812 3828
rect 3856 3824 3858 3828
rect 3112 3809 3118 3812
rect 3277 3809 3297 3813
rect 3301 3809 3351 3813
rect 3355 3809 3494 3813
rect 3498 3809 3582 3813
rect 3112 3804 3115 3809
rect 3064 3798 3069 3803
rect 3073 3776 3076 3804
rect 3280 3805 3283 3809
rect 3103 3776 3106 3800
rect 3289 3792 3292 3797
rect 3304 3799 3307 3809
rect 3334 3805 3337 3809
rect 3273 3788 3274 3791
rect 3278 3788 3281 3791
rect 3320 3788 3323 3791
rect 3289 3783 3292 3788
rect 3297 3784 3308 3787
rect 3320 3785 3328 3788
rect 3320 3779 3323 3785
rect 3332 3780 3335 3783
rect 3343 3783 3346 3797
rect 3454 3802 3457 3809
rect 3507 3802 3510 3809
rect 3713 3804 3716 3807
rect 3724 3807 3727 3813
rect 3731 3807 3734 3813
rect 3724 3804 3734 3807
rect 3343 3780 3355 3783
rect 2696 3772 2770 3776
rect 2774 3772 2776 3776
rect 2780 3772 2784 3776
rect 2788 3772 2802 3776
rect 2806 3772 2811 3776
rect 2815 3772 2820 3776
rect 2824 3772 2843 3776
rect 2847 3772 2877 3776
rect 2881 3772 2892 3776
rect 2896 3772 2920 3776
rect 2924 3772 2937 3776
rect 2941 3772 2961 3776
rect 2965 3772 3015 3776
rect 3019 3772 3042 3776
rect 3046 3772 3066 3776
rect 3070 3772 3118 3776
rect 2708 3765 2784 3769
rect 2788 3765 2843 3769
rect 2847 3765 2868 3769
rect 2872 3765 2899 3769
rect 2903 3765 2932 3769
rect 2831 3758 2832 3762
rect 2856 3757 2857 3761
rect 2903 3758 2904 3762
rect 2968 3753 2971 3772
rect 3073 3753 3076 3772
rect 2779 3744 2782 3749
rect 2786 3744 2789 3749
rect 2769 3741 2771 3744
rect 2779 3741 2789 3744
rect 2779 3735 2782 3741
rect 2786 3735 2789 3741
rect 2795 3743 2798 3749
rect 2811 3744 2814 3749
rect 2795 3739 2797 3743
rect 2801 3739 2803 3743
rect 2811 3742 2817 3744
rect 2821 3742 2822 3744
rect 2811 3740 2822 3742
rect 2839 3742 2842 3749
rect 2795 3735 2798 3739
rect 2811 3735 2814 3740
rect 2840 3738 2842 3742
rect 2839 3735 2842 3738
rect 2855 3743 2858 3749
rect 2865 3743 2868 3749
rect 2886 3744 2889 3749
rect 2865 3739 2874 3743
rect 2886 3740 2887 3744
rect 2891 3741 2894 3744
rect 2911 3743 2914 3749
rect 2929 3744 2932 3749
rect 2855 3735 2858 3739
rect 2865 3735 2868 3739
rect 2886 3735 2889 3740
rect 2913 3739 2914 3743
rect 2958 3740 2963 3745
rect 2967 3741 2969 3744
rect 2984 3743 2987 3749
rect 2984 3740 2992 3743
rect 3064 3740 3069 3745
rect 3073 3741 3074 3744
rect 3089 3743 3092 3749
rect 3089 3740 3097 3743
rect 2911 3735 2914 3739
rect 2929 3735 2932 3740
rect 2984 3737 2987 3740
rect 3089 3737 3092 3740
rect 3280 3733 3283 3779
rect 3343 3775 3346 3780
rect 3304 3733 3307 3775
rect 3334 3733 3337 3771
rect 3352 3765 3355 3780
rect 3724 3799 3727 3804
rect 3731 3799 3734 3804
rect 3740 3809 3743 3813
rect 3740 3805 3742 3809
rect 3746 3805 3748 3809
rect 3756 3808 3759 3813
rect 3784 3810 3787 3813
rect 3756 3806 3767 3808
rect 3740 3799 3743 3805
rect 3756 3804 3762 3806
rect 3756 3799 3759 3804
rect 3766 3804 3767 3806
rect 3785 3806 3787 3810
rect 3784 3799 3787 3806
rect 3929 3817 3932 3820
rect 3800 3809 3803 3813
rect 3810 3809 3813 3813
rect 3810 3805 3819 3809
rect 3831 3808 3834 3813
rect 3856 3809 3859 3813
rect 3800 3799 3803 3805
rect 3810 3799 3813 3805
rect 3831 3804 3832 3808
rect 3836 3804 3839 3807
rect 3858 3805 3859 3809
rect 3874 3808 3877 3813
rect 3906 3813 3917 3816
rect 3929 3814 3937 3817
rect 3831 3799 3834 3804
rect 3856 3799 3859 3805
rect 3906 3807 3909 3813
rect 3929 3808 3932 3814
rect 3941 3809 3944 3812
rect 3952 3812 3955 3826
rect 4003 3821 4006 3826
rect 4018 3828 4021 3838
rect 4048 3834 4051 3838
rect 3987 3817 3988 3820
rect 3992 3817 3995 3820
rect 4034 3817 4037 3820
rect 3960 3812 3965 3817
rect 4003 3812 4006 3817
rect 3952 3809 3960 3812
rect 3874 3799 3877 3804
rect 3952 3804 3955 3809
rect 4011 3813 4022 3816
rect 4034 3814 4042 3817
rect 3904 3798 3909 3803
rect 3776 3786 3777 3790
rect 3801 3787 3802 3791
rect 3848 3786 3849 3790
rect 3653 3779 3729 3783
rect 3733 3779 3788 3783
rect 3792 3779 3813 3783
rect 3817 3779 3844 3783
rect 3848 3779 3877 3783
rect 3913 3776 3916 3804
rect 3943 3776 3946 3800
rect 3994 3776 3997 3808
rect 4011 3807 4014 3813
rect 4034 3808 4037 3814
rect 4046 3809 4049 3812
rect 4057 3812 4060 3826
rect 4057 3809 4063 3812
rect 4057 3804 4060 3809
rect 4009 3798 4014 3803
rect 4018 3776 4021 3804
rect 4048 3776 4051 3800
rect 3641 3772 3715 3776
rect 3719 3772 3721 3776
rect 3725 3772 3729 3776
rect 3733 3772 3747 3776
rect 3751 3772 3756 3776
rect 3760 3772 3765 3776
rect 3769 3772 3788 3776
rect 3792 3772 3822 3776
rect 3826 3772 3837 3776
rect 3841 3772 3865 3776
rect 3869 3772 3882 3776
rect 3886 3772 3906 3776
rect 3910 3772 3960 3776
rect 3964 3772 3987 3776
rect 3991 3772 4011 3776
rect 4015 3772 4063 3776
rect 3352 3760 3469 3765
rect 3487 3764 3490 3772
rect 3487 3760 3507 3764
rect 3511 3760 3522 3764
rect 3487 3752 3490 3760
rect 3540 3756 3543 3772
rect 3653 3765 3729 3769
rect 3733 3765 3788 3769
rect 3792 3765 3813 3769
rect 3817 3765 3844 3769
rect 3848 3765 3877 3769
rect 3776 3758 3777 3762
rect 3801 3757 3802 3761
rect 3848 3758 3849 3762
rect 3544 3752 3659 3756
rect 3913 3753 3916 3772
rect 4018 3753 4021 3772
rect 3586 3740 3623 3744
rect 3724 3744 3727 3749
rect 3731 3744 3734 3749
rect 3714 3741 3716 3744
rect 3724 3741 3734 3744
rect 3454 3733 3457 3740
rect 3507 3733 3510 3740
rect 3574 3733 3635 3737
rect 3724 3735 3727 3741
rect 3277 3729 3297 3733
rect 3301 3729 3351 3733
rect 3355 3729 3494 3733
rect 3498 3729 3574 3733
rect 2839 3720 2842 3724
rect 2866 3720 2867 3724
rect 2911 3720 2913 3724
rect 2720 3713 2796 3717
rect 2800 3713 2827 3717
rect 2831 3713 2849 3717
rect 2853 3713 2914 3717
rect 2918 3713 2932 3717
rect 2968 3710 2971 3729
rect 3073 3710 3076 3729
rect 3304 3719 3307 3729
rect 3594 3724 3695 3728
rect 3731 3735 3734 3741
rect 3740 3743 3743 3749
rect 3756 3744 3759 3749
rect 3740 3739 3742 3743
rect 3746 3739 3748 3743
rect 3756 3742 3762 3744
rect 3766 3742 3767 3744
rect 3756 3740 3767 3742
rect 3784 3742 3787 3749
rect 3740 3735 3743 3739
rect 3756 3735 3759 3740
rect 3785 3738 3787 3742
rect 3784 3735 3787 3738
rect 3800 3743 3803 3749
rect 3810 3743 3813 3749
rect 3831 3744 3834 3749
rect 3810 3739 3819 3743
rect 3831 3740 3832 3744
rect 3836 3741 3839 3744
rect 3856 3743 3859 3749
rect 3874 3744 3877 3749
rect 3800 3735 3803 3739
rect 3810 3735 3813 3739
rect 3831 3735 3834 3740
rect 3858 3739 3859 3743
rect 3903 3740 3908 3745
rect 3912 3741 3914 3744
rect 3929 3743 3932 3749
rect 3929 3740 3937 3743
rect 4009 3740 4014 3745
rect 4018 3741 4019 3744
rect 4034 3743 4037 3749
rect 4034 3740 4042 3743
rect 3856 3735 3859 3739
rect 3874 3735 3877 3740
rect 3929 3737 3932 3740
rect 4034 3737 4037 3740
rect 3784 3720 3787 3724
rect 3811 3720 3812 3724
rect 3856 3720 3858 3724
rect 3512 3715 3647 3719
rect 2684 3706 2769 3710
rect 2773 3706 2785 3710
rect 2789 3706 2803 3710
rect 2807 3706 2814 3710
rect 2818 3706 2820 3710
rect 2824 3706 2839 3710
rect 2843 3706 2876 3710
rect 2880 3706 2881 3710
rect 2885 3706 2893 3710
rect 2897 3706 2921 3710
rect 2925 3706 2937 3710
rect 2941 3706 2961 3710
rect 2965 3706 3015 3710
rect 3019 3706 3042 3710
rect 3046 3706 3096 3710
rect 3100 3706 3104 3710
rect 3108 3706 3132 3710
rect 3136 3706 3186 3710
rect 3244 3707 3305 3710
rect 3320 3709 3323 3715
rect 3665 3713 3741 3717
rect 3745 3713 3772 3717
rect 3776 3713 3794 3717
rect 3798 3713 3859 3717
rect 3863 3713 3877 3717
rect 3913 3710 3916 3729
rect 4018 3710 4021 3729
rect 3320 3706 3328 3709
rect 3629 3706 3714 3710
rect 3718 3706 3730 3710
rect 3734 3706 3748 3710
rect 3752 3706 3759 3710
rect 3763 3706 3765 3710
rect 3769 3706 3784 3710
rect 3788 3706 3821 3710
rect 3825 3706 3826 3710
rect 3830 3706 3838 3710
rect 3842 3706 3866 3710
rect 3870 3706 3882 3710
rect 3886 3706 3906 3710
rect 3910 3706 3960 3710
rect 3964 3706 3987 3710
rect 3991 3706 4041 3710
rect 4045 3706 4049 3710
rect 4053 3706 4077 3710
rect 4081 3706 4131 3710
rect 2720 3699 2796 3703
rect 2800 3699 2827 3703
rect 2831 3699 2849 3703
rect 2853 3699 2914 3703
rect 2918 3699 2932 3703
rect 2968 3696 2971 3706
rect 2998 3702 3001 3706
rect 3025 3702 3028 3706
rect 2839 3692 2842 3696
rect 2866 3692 2867 3696
rect 2911 3692 2913 3696
rect 2768 3672 2771 3675
rect 2779 3675 2782 3681
rect 2786 3675 2789 3681
rect 2779 3672 2789 3675
rect 2779 3667 2782 3672
rect 2786 3667 2789 3672
rect 2795 3677 2798 3681
rect 2795 3673 2797 3677
rect 2801 3673 2803 3677
rect 2811 3676 2814 3681
rect 2839 3678 2842 3681
rect 2811 3674 2822 3676
rect 2795 3667 2798 3673
rect 2811 3672 2817 3674
rect 2811 3667 2814 3672
rect 2821 3672 2822 3674
rect 2840 3674 2842 3678
rect 2839 3667 2842 3674
rect 2984 3685 2987 3688
rect 2855 3677 2858 3681
rect 2865 3677 2868 3681
rect 2865 3673 2874 3677
rect 2886 3676 2889 3681
rect 2911 3677 2914 3681
rect 2855 3667 2858 3673
rect 2865 3667 2868 3673
rect 2886 3672 2887 3676
rect 2891 3672 2894 3675
rect 2913 3673 2914 3677
rect 2929 3676 2932 3681
rect 2961 3681 2972 3684
rect 2984 3682 2992 3685
rect 2886 3667 2889 3672
rect 2911 3667 2914 3673
rect 2961 3675 2964 3681
rect 2984 3676 2987 3682
rect 2996 3677 2999 3680
rect 3007 3680 3010 3694
rect 3034 3689 3037 3694
rect 3049 3696 3052 3706
rect 3079 3702 3082 3706
rect 3115 3702 3118 3706
rect 3018 3685 3019 3688
rect 3023 3685 3026 3688
rect 3065 3685 3068 3688
rect 3007 3677 3015 3680
rect 3034 3680 3037 3685
rect 2929 3667 2932 3672
rect 3007 3672 3010 3677
rect 3015 3673 3019 3677
rect 3042 3681 3053 3684
rect 3065 3682 3073 3685
rect 2959 3666 2964 3671
rect 2831 3654 2832 3658
rect 2856 3655 2857 3659
rect 2903 3654 2904 3658
rect 2708 3647 2784 3651
rect 2788 3647 2843 3651
rect 2847 3647 2868 3651
rect 2872 3647 2899 3651
rect 2903 3647 2932 3651
rect 2968 3644 2971 3672
rect 2998 3644 3001 3668
rect 3025 3644 3028 3676
rect 3042 3675 3045 3681
rect 3065 3676 3068 3682
rect 3077 3677 3080 3680
rect 3088 3680 3091 3694
rect 3124 3689 3127 3694
rect 3139 3696 3142 3706
rect 3169 3702 3172 3706
rect 3320 3703 3323 3706
rect 3113 3685 3116 3688
rect 3155 3685 3158 3688
rect 3088 3677 3097 3680
rect 3124 3680 3127 3685
rect 3088 3672 3091 3677
rect 3040 3666 3045 3671
rect 3049 3644 3052 3672
rect 3131 3683 3143 3684
rect 3135 3681 3143 3683
rect 3155 3682 3163 3685
rect 3155 3676 3158 3682
rect 3167 3677 3170 3680
rect 3178 3680 3181 3694
rect 3665 3699 3741 3703
rect 3745 3699 3772 3703
rect 3776 3699 3794 3703
rect 3798 3699 3859 3703
rect 3863 3699 3877 3703
rect 3913 3696 3916 3706
rect 3943 3702 3946 3706
rect 3970 3702 3973 3706
rect 3304 3683 3307 3695
rect 3784 3692 3787 3696
rect 3811 3692 3812 3696
rect 3856 3692 3858 3696
rect 3178 3677 3198 3680
rect 3079 3644 3082 3668
rect 3115 3644 3118 3676
rect 3178 3672 3181 3677
rect 3255 3679 3273 3683
rect 3277 3679 3297 3683
rect 3301 3679 3351 3683
rect 3355 3679 3400 3683
rect 3404 3679 3582 3683
rect 3139 3644 3142 3672
rect 3258 3675 3261 3679
rect 3280 3675 3283 3679
rect 3169 3644 3172 3668
rect 3267 3662 3270 3667
rect 3289 3662 3292 3667
rect 3304 3669 3307 3679
rect 3334 3675 3337 3679
rect 3251 3658 3252 3661
rect 3256 3658 3259 3661
rect 3271 3658 3274 3662
rect 3278 3658 3281 3661
rect 3320 3658 3323 3661
rect 3267 3653 3270 3658
rect 3289 3653 3292 3658
rect 3297 3654 3308 3657
rect 3320 3655 3328 3658
rect 3320 3649 3323 3655
rect 3332 3650 3335 3653
rect 3343 3653 3346 3667
rect 3360 3672 3363 3679
rect 3413 3672 3416 3679
rect 3713 3672 3716 3675
rect 3724 3675 3727 3681
rect 3731 3675 3734 3681
rect 3724 3672 3734 3675
rect 3343 3650 3355 3653
rect 2696 3640 2770 3644
rect 2774 3640 2776 3644
rect 2780 3640 2784 3644
rect 2788 3640 2802 3644
rect 2806 3640 2811 3644
rect 2815 3640 2820 3644
rect 2824 3640 2843 3644
rect 2847 3640 2877 3644
rect 2881 3640 2892 3644
rect 2896 3640 2920 3644
rect 2924 3640 2937 3644
rect 2941 3640 2961 3644
rect 2965 3640 3015 3644
rect 3022 3640 3042 3644
rect 3046 3640 3096 3644
rect 3100 3640 3132 3644
rect 3136 3640 3186 3644
rect 2708 3633 2784 3637
rect 2788 3633 2843 3637
rect 2847 3633 2868 3637
rect 2872 3633 2899 3637
rect 2903 3633 2932 3637
rect 2831 3626 2832 3630
rect 2856 3625 2857 3629
rect 2903 3626 2904 3630
rect 2779 3612 2782 3617
rect 2786 3612 2789 3617
rect 2769 3609 2771 3612
rect 2779 3609 2789 3612
rect 2779 3603 2782 3609
rect 2786 3603 2789 3609
rect 2795 3611 2798 3617
rect 2811 3612 2814 3617
rect 2795 3607 2797 3611
rect 2801 3607 2803 3611
rect 2811 3610 2817 3612
rect 2821 3610 2822 3612
rect 2811 3608 2822 3610
rect 2839 3610 2842 3617
rect 2795 3603 2798 3607
rect 2811 3603 2814 3608
rect 2840 3606 2842 3610
rect 2839 3603 2842 3606
rect 2855 3611 2858 3617
rect 2865 3611 2868 3617
rect 2886 3612 2889 3617
rect 2865 3607 2874 3611
rect 2886 3608 2887 3612
rect 2891 3609 2894 3612
rect 2911 3611 2914 3617
rect 2929 3612 2932 3617
rect 2968 3618 2971 3640
rect 3049 3618 3052 3640
rect 3139 3618 3142 3640
rect 2855 3603 2858 3607
rect 2865 3603 2868 3607
rect 2886 3603 2889 3608
rect 2913 3607 2914 3611
rect 2911 3603 2914 3607
rect 2929 3603 2932 3608
rect 2959 3605 2964 3610
rect 2968 3606 2969 3609
rect 2984 3608 2987 3614
rect 2984 3605 2992 3608
rect 3039 3605 3044 3610
rect 3048 3606 3050 3609
rect 3065 3608 3068 3614
rect 3065 3605 3073 3608
rect 3132 3606 3140 3609
rect 3155 3608 3158 3614
rect 3155 3605 3163 3608
rect 2984 3602 2987 3605
rect 3065 3602 3068 3605
rect 3155 3602 3158 3605
rect 3258 3603 3261 3649
rect 3280 3603 3283 3649
rect 3343 3645 3346 3650
rect 3304 3603 3307 3645
rect 3334 3603 3337 3641
rect 3352 3635 3355 3650
rect 3724 3667 3727 3672
rect 3731 3667 3734 3672
rect 3740 3677 3743 3681
rect 3740 3673 3742 3677
rect 3746 3673 3748 3677
rect 3756 3676 3759 3681
rect 3784 3678 3787 3681
rect 3756 3674 3767 3676
rect 3740 3667 3743 3673
rect 3756 3672 3762 3674
rect 3756 3667 3759 3672
rect 3766 3672 3767 3674
rect 3785 3674 3787 3678
rect 3784 3667 3787 3674
rect 3929 3685 3932 3688
rect 3800 3677 3803 3681
rect 3810 3677 3813 3681
rect 3810 3673 3819 3677
rect 3831 3676 3834 3681
rect 3856 3677 3859 3681
rect 3800 3667 3803 3673
rect 3810 3667 3813 3673
rect 3831 3672 3832 3676
rect 3836 3672 3839 3675
rect 3858 3673 3859 3677
rect 3874 3676 3877 3681
rect 3906 3681 3917 3684
rect 3929 3682 3937 3685
rect 3831 3667 3834 3672
rect 3856 3667 3859 3673
rect 3906 3675 3909 3681
rect 3929 3676 3932 3682
rect 3941 3677 3944 3680
rect 3952 3680 3955 3694
rect 3979 3689 3982 3694
rect 3994 3696 3997 3706
rect 4024 3702 4027 3706
rect 4060 3702 4063 3706
rect 3963 3685 3964 3688
rect 3968 3685 3971 3688
rect 4010 3685 4013 3688
rect 3952 3677 3960 3680
rect 3979 3680 3982 3685
rect 3874 3667 3877 3672
rect 3952 3672 3955 3677
rect 3960 3673 3964 3677
rect 3987 3681 3998 3684
rect 4010 3682 4018 3685
rect 3904 3666 3909 3671
rect 3776 3654 3777 3658
rect 3801 3655 3802 3659
rect 3848 3654 3849 3658
rect 3653 3647 3729 3651
rect 3733 3647 3788 3651
rect 3792 3647 3813 3651
rect 3817 3647 3844 3651
rect 3848 3647 3877 3651
rect 3913 3644 3916 3672
rect 3943 3644 3946 3668
rect 3970 3644 3973 3676
rect 3987 3675 3990 3681
rect 4010 3676 4013 3682
rect 4022 3677 4025 3680
rect 4033 3680 4036 3694
rect 4069 3689 4072 3694
rect 4084 3696 4087 3706
rect 4114 3702 4117 3706
rect 4058 3685 4061 3688
rect 4100 3685 4103 3688
rect 4033 3677 4042 3680
rect 4069 3680 4072 3685
rect 4033 3672 4036 3677
rect 3985 3666 3990 3671
rect 3994 3644 3997 3672
rect 4076 3683 4088 3684
rect 4080 3681 4088 3683
rect 4100 3682 4108 3685
rect 4100 3676 4103 3682
rect 4112 3677 4115 3680
rect 4123 3680 4126 3694
rect 4123 3677 4143 3680
rect 4024 3644 4027 3668
rect 4060 3644 4063 3676
rect 4123 3672 4126 3677
rect 4084 3644 4087 3672
rect 4114 3644 4117 3668
rect 3352 3630 3375 3635
rect 3393 3634 3396 3642
rect 3393 3630 3402 3634
rect 3406 3630 3428 3634
rect 3393 3622 3396 3630
rect 3446 3626 3449 3642
rect 3641 3640 3715 3644
rect 3719 3640 3721 3644
rect 3725 3640 3729 3644
rect 3733 3640 3747 3644
rect 3751 3640 3756 3644
rect 3760 3640 3765 3644
rect 3769 3640 3788 3644
rect 3792 3640 3822 3644
rect 3826 3640 3837 3644
rect 3841 3640 3865 3644
rect 3869 3640 3882 3644
rect 3886 3640 3906 3644
rect 3910 3640 3960 3644
rect 3967 3640 3987 3644
rect 3991 3640 4041 3644
rect 4045 3640 4077 3644
rect 4081 3640 4131 3644
rect 3653 3633 3729 3637
rect 3733 3633 3788 3637
rect 3792 3633 3813 3637
rect 3817 3633 3844 3637
rect 3848 3633 3877 3637
rect 3776 3626 3777 3630
rect 3801 3625 3802 3629
rect 3848 3626 3849 3630
rect 3450 3622 3683 3623
rect 3449 3619 3683 3622
rect 3360 3603 3363 3610
rect 3413 3603 3416 3610
rect 3724 3612 3727 3617
rect 3731 3612 3734 3617
rect 3714 3609 3716 3612
rect 3724 3609 3734 3612
rect 3724 3603 3727 3609
rect 2839 3588 2842 3592
rect 2866 3588 2867 3592
rect 2911 3588 2913 3592
rect 3255 3599 3273 3603
rect 3277 3599 3297 3603
rect 3301 3599 3351 3603
rect 3355 3599 3400 3603
rect 3404 3599 3574 3603
rect 2720 3581 2796 3585
rect 2800 3581 2827 3585
rect 2831 3581 2849 3585
rect 2853 3581 2914 3585
rect 2918 3581 2932 3585
rect 2968 3578 2971 3594
rect 3049 3578 3052 3594
rect 3139 3578 3142 3594
rect 3304 3589 3307 3599
rect 3731 3603 3734 3609
rect 3740 3611 3743 3617
rect 3756 3612 3759 3617
rect 3740 3607 3742 3611
rect 3746 3607 3748 3611
rect 3756 3610 3762 3612
rect 3766 3610 3767 3612
rect 3756 3608 3767 3610
rect 3784 3610 3787 3617
rect 3740 3603 3743 3607
rect 3756 3603 3759 3608
rect 3785 3606 3787 3610
rect 3784 3603 3787 3606
rect 3800 3611 3803 3617
rect 3810 3611 3813 3617
rect 3831 3612 3834 3617
rect 3810 3607 3819 3611
rect 3831 3608 3832 3612
rect 3836 3609 3839 3612
rect 3856 3611 3859 3617
rect 3874 3612 3877 3617
rect 3913 3618 3916 3640
rect 3994 3618 3997 3640
rect 4084 3618 4087 3640
rect 3800 3603 3803 3607
rect 3810 3603 3813 3607
rect 3831 3603 3834 3608
rect 3858 3607 3859 3611
rect 3856 3603 3859 3607
rect 3874 3603 3877 3608
rect 3904 3605 3909 3610
rect 3913 3606 3914 3609
rect 3929 3608 3932 3614
rect 3929 3605 3937 3608
rect 3984 3605 3989 3610
rect 3993 3606 3995 3609
rect 4010 3608 4013 3614
rect 4010 3605 4018 3608
rect 4077 3606 4085 3609
rect 4100 3608 4103 3614
rect 4100 3605 4108 3608
rect 3929 3602 3932 3605
rect 4010 3602 4013 3605
rect 4100 3602 4103 3605
rect 3406 3589 3671 3593
rect 3784 3588 3787 3592
rect 3811 3588 3812 3592
rect 3856 3588 3858 3592
rect 2684 3574 2769 3578
rect 2773 3574 2785 3578
rect 2789 3574 2803 3578
rect 2807 3574 2814 3578
rect 2818 3574 2820 3578
rect 2824 3574 2839 3578
rect 2843 3574 2876 3578
rect 2880 3574 2881 3578
rect 2885 3574 2893 3578
rect 2897 3574 2921 3578
rect 2925 3574 2937 3578
rect 2941 3574 2961 3578
rect 2965 3574 3015 3578
rect 3019 3574 3042 3578
rect 3046 3574 3132 3578
rect 3136 3574 3190 3578
rect 3246 3577 3305 3580
rect 3320 3579 3323 3585
rect 3665 3581 3741 3585
rect 3745 3581 3772 3585
rect 3776 3581 3794 3585
rect 3798 3581 3859 3585
rect 3863 3581 3877 3585
rect 3320 3576 3328 3579
rect 3913 3578 3916 3594
rect 3994 3578 3997 3594
rect 4084 3578 4087 3594
rect 2720 3567 2796 3571
rect 2800 3567 2827 3571
rect 2831 3567 2849 3571
rect 2853 3567 2914 3571
rect 2918 3567 2932 3571
rect 2968 3564 2971 3574
rect 2998 3570 3001 3574
rect 3320 3573 3323 3576
rect 3629 3574 3714 3578
rect 3718 3574 3730 3578
rect 3734 3574 3748 3578
rect 3752 3574 3759 3578
rect 3763 3574 3765 3578
rect 3769 3574 3784 3578
rect 3788 3574 3821 3578
rect 3825 3574 3826 3578
rect 3830 3574 3838 3578
rect 3842 3574 3866 3578
rect 3870 3574 3882 3578
rect 3886 3574 3906 3578
rect 3910 3574 3960 3578
rect 3964 3574 3987 3578
rect 3991 3574 4077 3578
rect 4081 3574 4135 3578
rect 2839 3560 2842 3564
rect 2866 3560 2867 3564
rect 2911 3560 2913 3564
rect 2768 3540 2771 3543
rect 2779 3543 2782 3549
rect 2786 3543 2789 3549
rect 2779 3540 2789 3543
rect 2779 3535 2782 3540
rect 2786 3535 2789 3540
rect 2795 3545 2798 3549
rect 2795 3541 2797 3545
rect 2801 3541 2803 3545
rect 2811 3544 2814 3549
rect 2839 3546 2842 3549
rect 2811 3542 2822 3544
rect 2795 3535 2798 3541
rect 2811 3540 2817 3542
rect 2811 3535 2814 3540
rect 2821 3540 2822 3542
rect 2840 3542 2842 3546
rect 2839 3535 2842 3542
rect 2984 3553 2987 3556
rect 2855 3545 2858 3549
rect 2865 3545 2868 3549
rect 2865 3541 2874 3545
rect 2886 3544 2889 3549
rect 2911 3545 2914 3549
rect 2855 3535 2858 3541
rect 2865 3535 2868 3541
rect 2886 3540 2887 3544
rect 2891 3540 2894 3543
rect 2913 3541 2914 3545
rect 2929 3544 2932 3549
rect 2961 3549 2972 3552
rect 2984 3550 2992 3553
rect 2886 3535 2889 3540
rect 2911 3535 2914 3541
rect 2961 3543 2964 3549
rect 2984 3544 2987 3550
rect 2996 3545 2999 3548
rect 3007 3548 3010 3562
rect 3665 3567 3741 3571
rect 3745 3567 3772 3571
rect 3776 3567 3794 3571
rect 3798 3567 3859 3571
rect 3863 3567 3877 3571
rect 3304 3553 3307 3565
rect 3913 3564 3916 3574
rect 3943 3570 3946 3574
rect 3784 3560 3787 3564
rect 3811 3560 3812 3564
rect 3856 3560 3858 3564
rect 3015 3548 3020 3553
rect 3273 3549 3297 3553
rect 3301 3549 3582 3553
rect 3007 3545 3015 3548
rect 2929 3535 2932 3540
rect 3007 3540 3010 3545
rect 3713 3540 3716 3543
rect 3724 3543 3727 3549
rect 3731 3543 3734 3549
rect 3724 3540 3734 3543
rect 2959 3534 2964 3539
rect 2269 3526 2390 3530
rect 2278 3519 2287 3523
rect 2291 3519 2323 3523
rect 2327 3519 2390 3523
rect 2394 3519 2419 3523
rect 2423 3519 2455 3523
rect 2459 3519 2522 3523
rect 2526 3519 2551 3523
rect 2555 3519 2587 3523
rect 2591 3519 2654 3523
rect 2658 3519 2738 3523
rect 2831 3522 2832 3526
rect 2856 3523 2857 3527
rect 2903 3522 2904 3526
rect 2278 3512 2311 3516
rect 2315 3512 2339 3516
rect 2343 3512 2369 3516
rect 2373 3512 2406 3516
rect 2410 3512 2443 3516
rect 2447 3512 2471 3516
rect 2475 3512 2501 3516
rect 2505 3512 2538 3516
rect 2542 3512 2575 3516
rect 2579 3512 2603 3516
rect 2607 3512 2633 3516
rect 2637 3512 2670 3516
rect 2674 3512 2678 3516
rect 2763 3515 2784 3519
rect 2788 3515 2793 3519
rect 2797 3515 2843 3519
rect 2847 3515 2868 3519
rect 2872 3515 2899 3519
rect 2903 3515 2932 3519
rect 2968 3512 2971 3540
rect 2998 3512 3001 3536
rect 3724 3535 3727 3540
rect 3731 3535 3734 3540
rect 3740 3545 3743 3549
rect 3740 3541 3742 3545
rect 3746 3541 3748 3545
rect 3756 3544 3759 3549
rect 3784 3546 3787 3549
rect 3756 3542 3767 3544
rect 3740 3535 3743 3541
rect 3756 3540 3762 3542
rect 3756 3535 3759 3540
rect 3766 3540 3767 3542
rect 3785 3542 3787 3546
rect 3784 3535 3787 3542
rect 3929 3553 3932 3556
rect 3800 3545 3803 3549
rect 3810 3545 3813 3549
rect 3810 3541 3819 3545
rect 3831 3544 3834 3549
rect 3856 3545 3859 3549
rect 3800 3535 3803 3541
rect 3810 3535 3813 3541
rect 3831 3540 3832 3544
rect 3836 3540 3839 3543
rect 3858 3541 3859 3545
rect 3874 3544 3877 3549
rect 3906 3549 3917 3552
rect 3929 3550 3937 3553
rect 3831 3535 3834 3540
rect 3856 3535 3859 3541
rect 3906 3543 3909 3549
rect 3929 3544 3932 3550
rect 3941 3545 3944 3548
rect 3952 3548 3955 3562
rect 3960 3548 3965 3553
rect 3952 3545 3960 3548
rect 3874 3535 3877 3540
rect 3952 3540 3955 3545
rect 3904 3534 3909 3539
rect 3223 3519 3232 3523
rect 3236 3519 3268 3523
rect 3272 3519 3335 3523
rect 3339 3519 3364 3523
rect 3368 3519 3400 3523
rect 3404 3519 3467 3523
rect 3471 3519 3496 3523
rect 3500 3519 3532 3523
rect 3536 3519 3599 3523
rect 3603 3519 3683 3523
rect 3776 3522 3777 3526
rect 3801 3523 3802 3527
rect 3848 3522 3849 3526
rect 3223 3512 3256 3516
rect 3260 3512 3284 3516
rect 3288 3512 3314 3516
rect 3318 3512 3351 3516
rect 3355 3512 3388 3516
rect 3392 3512 3416 3516
rect 3420 3512 3446 3516
rect 3450 3512 3483 3516
rect 3487 3512 3520 3516
rect 3524 3512 3548 3516
rect 3552 3512 3578 3516
rect 3582 3512 3615 3516
rect 3619 3512 3623 3516
rect 3708 3515 3729 3519
rect 3733 3515 3738 3519
rect 3742 3515 3788 3519
rect 3792 3515 3813 3519
rect 3817 3515 3844 3519
rect 3848 3515 3877 3519
rect 3913 3512 3916 3540
rect 3943 3512 3946 3536
rect 2281 3502 2284 3512
rect 2302 3502 2305 3512
rect 2318 3502 2321 3512
rect 2332 3505 2337 3509
rect 2341 3505 2348 3509
rect 2360 3502 2363 3512
rect 2376 3502 2379 3512
rect 2397 3502 2400 3512
rect 2413 3502 2416 3512
rect 2434 3502 2437 3512
rect 2450 3502 2453 3512
rect 2464 3505 2469 3509
rect 2473 3505 2480 3509
rect 2492 3502 2495 3512
rect 2508 3502 2511 3512
rect 2529 3502 2532 3512
rect 2545 3502 2548 3512
rect 2566 3502 2569 3512
rect 2582 3502 2585 3512
rect 2596 3505 2601 3509
rect 2605 3505 2612 3509
rect 2624 3502 2627 3512
rect 2640 3502 2643 3512
rect 2661 3502 2664 3512
rect 2696 3508 2770 3512
rect 2774 3508 2776 3512
rect 2780 3508 2784 3512
rect 2788 3508 2802 3512
rect 2806 3508 2811 3512
rect 2815 3508 2820 3512
rect 2824 3508 2843 3512
rect 2847 3508 2877 3512
rect 2881 3508 2892 3512
rect 2896 3508 2920 3512
rect 2924 3508 2937 3512
rect 2941 3508 2961 3512
rect 2965 3508 3045 3512
rect 3049 3508 3063 3512
rect 3067 3508 3072 3512
rect 3076 3508 3081 3512
rect 3085 3508 3104 3512
rect 3108 3508 3138 3512
rect 3142 3508 3153 3512
rect 3157 3508 3181 3512
rect 3185 3508 3194 3512
rect 2298 3488 2303 3491
rect 2307 3488 2331 3491
rect 2356 3488 2363 3491
rect 2367 3488 2389 3491
rect 2409 3488 2416 3491
rect 2430 3488 2435 3491
rect 2439 3488 2463 3491
rect 2488 3488 2495 3491
rect 2499 3488 2521 3491
rect 2541 3488 2548 3491
rect 2562 3488 2567 3491
rect 2571 3488 2595 3491
rect 2708 3501 2784 3505
rect 2788 3501 2793 3505
rect 2797 3501 2843 3505
rect 2847 3501 2868 3505
rect 2872 3501 2899 3505
rect 2903 3501 2932 3505
rect 2620 3488 2627 3491
rect 2631 3488 2653 3491
rect 2831 3494 2832 3498
rect 2856 3493 2857 3497
rect 2903 3494 2904 3498
rect 2314 3478 2321 3481
rect 2325 3482 2344 3485
rect 2344 3475 2347 3481
rect 2372 3478 2379 3481
rect 2383 3482 2398 3485
rect 2446 3478 2453 3481
rect 2457 3482 2476 3485
rect 2476 3475 2479 3481
rect 2504 3478 2511 3481
rect 2515 3482 2530 3485
rect 2578 3478 2585 3481
rect 2589 3482 2608 3485
rect 2608 3475 2611 3481
rect 2636 3478 2643 3481
rect 2647 3482 2664 3485
rect 2779 3480 2782 3485
rect 2786 3480 2789 3485
rect 2769 3477 2771 3480
rect 2779 3477 2789 3480
rect 2779 3471 2782 3477
rect 2281 3459 2284 3471
rect 2302 3459 2305 3471
rect 2318 3459 2321 3471
rect 2332 3462 2344 3465
rect 2360 3459 2363 3471
rect 2376 3459 2379 3471
rect 2397 3459 2400 3471
rect 2413 3459 2416 3471
rect 2434 3459 2437 3471
rect 2450 3459 2453 3471
rect 2464 3462 2476 3465
rect 2492 3459 2495 3471
rect 2508 3459 2511 3471
rect 2529 3459 2532 3471
rect 2545 3459 2548 3471
rect 2566 3459 2569 3471
rect 2582 3459 2585 3471
rect 2596 3462 2608 3465
rect 2624 3459 2627 3471
rect 2640 3459 2643 3471
rect 2661 3459 2664 3471
rect 2786 3471 2789 3477
rect 2795 3479 2798 3485
rect 2811 3480 2814 3485
rect 2795 3475 2797 3479
rect 2801 3475 2803 3479
rect 2811 3478 2817 3480
rect 2821 3478 2822 3480
rect 2811 3476 2822 3478
rect 2839 3478 2842 3485
rect 2795 3471 2798 3475
rect 2811 3471 2814 3476
rect 2840 3474 2842 3478
rect 2839 3471 2842 3474
rect 2855 3479 2858 3485
rect 2865 3479 2868 3485
rect 2886 3480 2889 3485
rect 2865 3475 2874 3479
rect 2886 3476 2887 3480
rect 2891 3477 2894 3480
rect 2911 3479 2914 3485
rect 2929 3480 2932 3485
rect 2968 3482 2971 3508
rect 3004 3501 3023 3505
rect 3027 3501 3045 3505
rect 3049 3501 3104 3505
rect 3108 3501 3129 3505
rect 3133 3501 3160 3505
rect 3164 3501 3193 3505
rect 3226 3502 3229 3512
rect 3247 3502 3250 3512
rect 3263 3502 3266 3512
rect 3277 3505 3282 3509
rect 3286 3505 3293 3509
rect 3305 3502 3308 3512
rect 3321 3502 3324 3512
rect 3342 3502 3345 3512
rect 3358 3502 3361 3512
rect 3379 3502 3382 3512
rect 3395 3502 3398 3512
rect 3409 3505 3414 3509
rect 3418 3505 3425 3509
rect 3437 3502 3440 3512
rect 3453 3502 3456 3512
rect 3474 3502 3477 3512
rect 3490 3502 3493 3512
rect 3511 3502 3514 3512
rect 3527 3502 3530 3512
rect 3541 3505 3546 3509
rect 3550 3505 3557 3509
rect 3569 3502 3572 3512
rect 3585 3502 3588 3512
rect 3606 3502 3609 3512
rect 3641 3508 3715 3512
rect 3719 3508 3721 3512
rect 3725 3508 3729 3512
rect 3733 3508 3747 3512
rect 3751 3508 3756 3512
rect 3760 3508 3765 3512
rect 3769 3508 3788 3512
rect 3792 3508 3822 3512
rect 3826 3508 3837 3512
rect 3841 3508 3865 3512
rect 3869 3508 3882 3512
rect 3886 3508 3906 3512
rect 3910 3508 3990 3512
rect 3994 3508 4008 3512
rect 4012 3508 4017 3512
rect 4021 3508 4026 3512
rect 4030 3508 4049 3512
rect 4053 3508 4083 3512
rect 4087 3508 4098 3512
rect 4102 3508 4126 3512
rect 4130 3508 4139 3512
rect 3004 3489 3007 3501
rect 3092 3494 3093 3498
rect 3117 3493 3118 3497
rect 3164 3494 3165 3498
rect 2855 3471 2858 3475
rect 2865 3471 2868 3475
rect 2886 3471 2889 3476
rect 2913 3475 2914 3479
rect 3031 3480 3034 3485
rect 3040 3480 3043 3485
rect 3047 3480 3050 3485
rect 2911 3471 2914 3475
rect 2929 3471 2932 3476
rect 2958 3469 2963 3474
rect 2967 3470 2969 3473
rect 2984 3472 2987 3478
rect 3016 3477 3050 3480
rect 2984 3469 2992 3472
rect 2984 3466 2987 3469
rect 2278 3455 2311 3459
rect 2315 3455 2339 3459
rect 2343 3455 2369 3459
rect 2373 3455 2443 3459
rect 2447 3455 2471 3459
rect 2475 3455 2501 3459
rect 2505 3455 2575 3459
rect 2579 3455 2603 3459
rect 2607 3455 2633 3459
rect 2637 3455 2690 3459
rect 2839 3456 2842 3460
rect 2866 3456 2867 3460
rect 2911 3456 2913 3460
rect 3016 3463 3019 3477
rect 3040 3471 3043 3477
rect 3047 3471 3050 3477
rect 3056 3479 3059 3485
rect 3072 3480 3075 3485
rect 3056 3475 3058 3479
rect 3062 3475 3064 3479
rect 3072 3478 3078 3480
rect 3082 3478 3083 3480
rect 3072 3476 3083 3478
rect 3100 3478 3103 3485
rect 3056 3471 3059 3475
rect 3072 3471 3075 3476
rect 3101 3474 3103 3478
rect 3100 3471 3103 3474
rect 3243 3488 3248 3491
rect 3252 3488 3276 3491
rect 3301 3488 3308 3491
rect 3312 3488 3334 3491
rect 3354 3488 3361 3491
rect 3375 3488 3380 3491
rect 3384 3488 3408 3491
rect 3433 3488 3440 3491
rect 3444 3488 3466 3491
rect 3486 3488 3493 3491
rect 3507 3488 3512 3491
rect 3516 3488 3540 3491
rect 3653 3501 3729 3505
rect 3733 3501 3738 3505
rect 3742 3501 3788 3505
rect 3792 3501 3813 3505
rect 3817 3501 3844 3505
rect 3848 3501 3877 3505
rect 3565 3488 3572 3491
rect 3576 3488 3598 3491
rect 3776 3494 3777 3498
rect 3801 3493 3802 3497
rect 3848 3494 3849 3498
rect 3116 3479 3119 3485
rect 3126 3479 3129 3485
rect 3147 3480 3150 3485
rect 3126 3475 3135 3479
rect 3147 3476 3148 3480
rect 3152 3477 3155 3480
rect 3172 3479 3175 3485
rect 3190 3480 3193 3485
rect 3116 3471 3119 3475
rect 3126 3471 3129 3475
rect 3147 3471 3150 3476
rect 3174 3475 3175 3479
rect 3172 3471 3175 3475
rect 3190 3471 3193 3476
rect 3259 3478 3266 3481
rect 3270 3482 3289 3485
rect 3289 3475 3292 3481
rect 3317 3478 3324 3481
rect 3328 3482 3343 3485
rect 3391 3478 3398 3481
rect 3402 3482 3421 3485
rect 3421 3475 3424 3481
rect 3449 3478 3456 3481
rect 3460 3482 3475 3485
rect 3523 3478 3530 3481
rect 3534 3482 3553 3485
rect 3553 3475 3556 3481
rect 3581 3478 3588 3481
rect 3592 3482 3609 3485
rect 3724 3480 3727 3485
rect 3731 3480 3734 3485
rect 3714 3477 3716 3480
rect 3724 3477 3734 3480
rect 3724 3471 3727 3477
rect 2278 3448 2287 3452
rect 2291 3448 2338 3452
rect 2342 3448 2388 3452
rect 2392 3448 2419 3452
rect 2423 3448 2470 3452
rect 2474 3448 2520 3452
rect 2524 3448 2551 3452
rect 2555 3448 2602 3452
rect 2606 3448 2652 3452
rect 2656 3449 2726 3452
rect 2782 3449 2796 3453
rect 2800 3449 2827 3453
rect 2831 3449 2849 3453
rect 2853 3449 2914 3453
rect 2918 3449 2932 3453
rect 2968 3446 2971 3458
rect 3100 3456 3103 3460
rect 3127 3456 3128 3460
rect 3172 3456 3174 3460
rect 3226 3459 3229 3471
rect 3247 3459 3250 3471
rect 3263 3459 3266 3471
rect 3277 3462 3289 3465
rect 3305 3459 3308 3471
rect 3321 3459 3324 3471
rect 3342 3459 3345 3471
rect 3358 3459 3361 3471
rect 3379 3459 3382 3471
rect 3395 3459 3398 3471
rect 3409 3462 3421 3465
rect 3437 3459 3440 3471
rect 3453 3459 3456 3471
rect 3474 3459 3477 3471
rect 3490 3459 3493 3471
rect 3511 3459 3514 3471
rect 3527 3459 3530 3471
rect 3541 3462 3553 3465
rect 3569 3459 3572 3471
rect 3585 3459 3588 3471
rect 3606 3459 3609 3471
rect 3731 3471 3734 3477
rect 3740 3479 3743 3485
rect 3756 3480 3759 3485
rect 3740 3475 3742 3479
rect 3746 3475 3748 3479
rect 3756 3478 3762 3480
rect 3766 3478 3767 3480
rect 3756 3476 3767 3478
rect 3784 3478 3787 3485
rect 3740 3471 3743 3475
rect 3756 3471 3759 3476
rect 3785 3474 3787 3478
rect 3784 3471 3787 3474
rect 3800 3479 3803 3485
rect 3810 3479 3813 3485
rect 3831 3480 3834 3485
rect 3810 3475 3819 3479
rect 3831 3476 3832 3480
rect 3836 3477 3839 3480
rect 3856 3479 3859 3485
rect 3874 3480 3877 3485
rect 3913 3482 3916 3508
rect 3949 3501 3968 3505
rect 3972 3501 3990 3505
rect 3994 3501 4049 3505
rect 4053 3501 4074 3505
rect 4078 3501 4105 3505
rect 4109 3501 4138 3505
rect 3949 3489 3952 3501
rect 4037 3494 4038 3498
rect 4062 3493 4063 3497
rect 4109 3494 4110 3498
rect 3800 3471 3803 3475
rect 3810 3471 3813 3475
rect 3831 3471 3834 3476
rect 3858 3475 3859 3479
rect 3976 3480 3979 3485
rect 3985 3480 3988 3485
rect 3992 3480 3995 3485
rect 3856 3471 3859 3475
rect 3874 3471 3877 3476
rect 3903 3469 3908 3474
rect 3912 3470 3914 3473
rect 3929 3472 3932 3478
rect 3961 3477 3995 3480
rect 3929 3469 3937 3472
rect 3929 3466 3932 3469
rect 3223 3455 3256 3459
rect 3260 3455 3284 3459
rect 3288 3455 3314 3459
rect 3318 3455 3388 3459
rect 3392 3455 3416 3459
rect 3420 3455 3446 3459
rect 3450 3455 3520 3459
rect 3524 3455 3548 3459
rect 3552 3455 3578 3459
rect 3582 3455 3635 3459
rect 3784 3456 3787 3460
rect 3811 3456 3812 3460
rect 3856 3456 3858 3460
rect 3961 3463 3964 3477
rect 3985 3471 3988 3477
rect 3992 3471 3995 3477
rect 4001 3479 4004 3485
rect 4017 3480 4020 3485
rect 4001 3475 4003 3479
rect 4007 3475 4009 3479
rect 4017 3478 4023 3480
rect 4027 3478 4028 3480
rect 4017 3476 4028 3478
rect 4045 3478 4048 3485
rect 4001 3471 4004 3475
rect 4017 3471 4020 3476
rect 4046 3474 4048 3478
rect 4045 3471 4048 3474
rect 4061 3479 4064 3485
rect 4071 3479 4074 3485
rect 4092 3480 4095 3485
rect 4071 3475 4080 3479
rect 4092 3476 4093 3480
rect 4097 3477 4100 3480
rect 4117 3479 4120 3485
rect 4135 3480 4138 3485
rect 4061 3471 4064 3475
rect 4071 3471 4074 3475
rect 4092 3471 4095 3476
rect 4119 3475 4120 3479
rect 4117 3471 4120 3475
rect 4135 3471 4138 3476
rect 3008 3449 3013 3453
rect 3017 3449 3057 3453
rect 3061 3449 3088 3453
rect 3092 3449 3110 3453
rect 3114 3449 3175 3453
rect 3179 3449 3193 3453
rect 3223 3448 3232 3452
rect 3236 3448 3283 3452
rect 3287 3448 3333 3452
rect 3337 3448 3364 3452
rect 3368 3448 3415 3452
rect 3419 3448 3465 3452
rect 3469 3448 3496 3452
rect 3500 3448 3547 3452
rect 3551 3448 3597 3452
rect 3601 3449 3671 3452
rect 3727 3449 3741 3453
rect 3745 3449 3772 3453
rect 3776 3449 3794 3453
rect 3798 3449 3859 3453
rect 3863 3449 3877 3453
rect 3913 3446 3916 3458
rect 4045 3456 4048 3460
rect 4072 3456 4073 3460
rect 4117 3456 4119 3460
rect 3953 3449 3958 3453
rect 3962 3449 4002 3453
rect 4006 3449 4033 3453
rect 4037 3449 4055 3453
rect 4059 3449 4120 3453
rect 4124 3449 4138 3453
rect 2285 3442 2669 3445
rect 2684 3442 2769 3446
rect 2773 3442 2785 3446
rect 2789 3442 2803 3446
rect 2807 3442 2814 3446
rect 2818 3442 2820 3446
rect 2824 3442 2839 3446
rect 2843 3442 2876 3446
rect 2880 3442 2881 3446
rect 2885 3442 2893 3446
rect 2897 3442 2921 3446
rect 2925 3442 2961 3446
rect 2965 3442 3004 3446
rect 3008 3442 3015 3446
rect 3019 3442 3030 3446
rect 3034 3442 3046 3446
rect 3050 3442 3064 3446
rect 3068 3442 3075 3446
rect 3079 3442 3081 3446
rect 3085 3442 3100 3446
rect 3104 3442 3137 3446
rect 3141 3442 3142 3446
rect 3146 3442 3154 3446
rect 3158 3442 3182 3446
rect 3186 3442 3194 3446
rect 3230 3442 3614 3445
rect 3629 3442 3714 3446
rect 3718 3442 3730 3446
rect 3734 3442 3748 3446
rect 3752 3442 3759 3446
rect 3763 3442 3765 3446
rect 3769 3442 3784 3446
rect 3788 3442 3821 3446
rect 3825 3442 3826 3446
rect 3830 3442 3838 3446
rect 3842 3442 3866 3446
rect 3870 3442 3906 3446
rect 3910 3442 3949 3446
rect 3953 3442 3960 3446
rect 3964 3442 3975 3446
rect 3979 3442 3991 3446
rect 3995 3442 4009 3446
rect 4013 3442 4020 3446
rect 4024 3442 4026 3446
rect 4030 3442 4045 3446
rect 4049 3442 4082 3446
rect 4086 3442 4087 3446
rect 4091 3442 4099 3446
rect 4103 3442 4127 3446
rect 4131 3442 4139 3446
rect 2428 3435 2537 3438
rect 2720 3435 2778 3439
rect 2782 3435 3012 3438
rect 3202 3436 3210 3440
rect 3373 3435 3482 3438
rect 3665 3435 3723 3439
rect 3727 3435 3957 3438
rect 4147 3436 4155 3440
rect 2408 3427 2412 3431
rect 2416 3427 2420 3431
rect 2708 3428 3022 3431
rect 2396 3426 2400 3427
rect 2428 3426 2432 3427
rect 2756 3421 3029 3424
rect 3198 3418 3202 3423
rect 3353 3427 3357 3431
rect 3361 3427 3365 3431
rect 3653 3428 3967 3431
rect 3341 3426 3345 3427
rect 3373 3426 3377 3427
rect 3701 3421 3972 3425
rect 4143 3418 4147 3423
rect 2269 3414 2396 3418
rect 2400 3414 2416 3418
rect 2432 3414 3341 3418
rect 3345 3414 3361 3418
rect 3377 3414 4235 3418
rect 2424 3407 2669 3410
rect 2744 3407 3070 3411
rect 3074 3407 3106 3411
rect 3110 3407 3173 3411
rect 3177 3407 3193 3411
rect 3369 3407 3614 3410
rect 3689 3407 4015 3411
rect 4019 3407 4051 3411
rect 4055 3407 4118 3411
rect 4122 3407 4138 3411
rect 2439 3400 2669 3403
rect 2684 3400 3056 3404
rect 3060 3400 3094 3404
rect 3098 3400 3122 3404
rect 3126 3400 3152 3404
rect 3156 3400 3189 3404
rect 2408 3391 2412 3395
rect 2416 3391 2420 3395
rect 3064 3390 3067 3400
rect 3085 3390 3088 3400
rect 3101 3390 3104 3400
rect 3115 3393 3120 3397
rect 3124 3393 3131 3397
rect 3143 3390 3146 3400
rect 3159 3390 3162 3400
rect 3180 3390 3183 3400
rect 3384 3400 3614 3403
rect 3629 3400 4001 3404
rect 4005 3400 4039 3404
rect 4043 3400 4067 3404
rect 4071 3400 4097 3404
rect 4101 3400 4134 3404
rect 3353 3391 3357 3395
rect 3361 3391 3365 3395
rect 4009 3390 4012 3400
rect 4030 3390 4033 3400
rect 4046 3390 4049 3400
rect 4060 3393 4065 3397
rect 4069 3393 4076 3397
rect 4088 3390 4091 3400
rect 4104 3390 4107 3400
rect 4125 3390 4128 3400
rect 2428 3384 2538 3387
rect 2278 3377 2287 3381
rect 2291 3377 2323 3381
rect 2327 3377 2390 3381
rect 2394 3377 2419 3381
rect 2423 3377 2455 3381
rect 2459 3377 2522 3381
rect 2526 3377 2551 3381
rect 2555 3377 2587 3381
rect 2591 3377 2654 3381
rect 2658 3377 2738 3381
rect 2278 3370 2311 3374
rect 2315 3370 2339 3374
rect 2343 3370 2369 3374
rect 2373 3370 2406 3374
rect 2410 3370 2443 3374
rect 2447 3370 2471 3374
rect 2475 3370 2501 3374
rect 2505 3370 2538 3374
rect 2542 3370 2575 3374
rect 2579 3370 2603 3374
rect 2607 3370 2633 3374
rect 2637 3370 2670 3374
rect 2674 3370 2678 3374
rect 3081 3376 3086 3379
rect 3090 3376 3114 3379
rect 3373 3384 3483 3387
rect 3139 3376 3146 3379
rect 3150 3376 3172 3379
rect 3223 3377 3232 3381
rect 3236 3377 3268 3381
rect 3272 3377 3335 3381
rect 3339 3377 3364 3381
rect 3368 3377 3400 3381
rect 3404 3377 3467 3381
rect 3471 3377 3496 3381
rect 3500 3377 3532 3381
rect 3536 3377 3599 3381
rect 3603 3377 3683 3381
rect 2281 3360 2284 3370
rect 2302 3360 2305 3370
rect 2318 3360 2321 3370
rect 2332 3363 2337 3367
rect 2341 3363 2348 3367
rect 2360 3360 2363 3370
rect 2376 3360 2379 3370
rect 2397 3360 2400 3370
rect 2413 3360 2416 3370
rect 2434 3360 2437 3370
rect 2450 3360 2453 3370
rect 2464 3363 2469 3367
rect 2473 3363 2480 3367
rect 2492 3360 2495 3370
rect 2508 3360 2511 3370
rect 2529 3360 2532 3370
rect 2545 3360 2548 3370
rect 2566 3360 2569 3370
rect 2582 3360 2585 3370
rect 2596 3363 2601 3367
rect 2605 3363 2612 3367
rect 2624 3360 2627 3370
rect 2640 3360 2643 3370
rect 2661 3360 2664 3370
rect 3097 3366 3104 3369
rect 3108 3370 3127 3373
rect 2298 3346 2303 3349
rect 2307 3346 2331 3349
rect 2356 3346 2363 3349
rect 2367 3346 2389 3349
rect 2409 3346 2416 3349
rect 2430 3346 2435 3349
rect 2439 3346 2463 3349
rect 2488 3346 2495 3349
rect 2499 3346 2521 3349
rect 2541 3346 2548 3349
rect 2562 3346 2567 3349
rect 2571 3346 2595 3349
rect 2620 3346 2627 3349
rect 2631 3346 2653 3349
rect 3127 3363 3130 3369
rect 3155 3366 3162 3369
rect 3166 3370 3181 3373
rect 3223 3370 3256 3374
rect 3260 3370 3284 3374
rect 3288 3370 3314 3374
rect 3318 3370 3351 3374
rect 3355 3370 3388 3374
rect 3392 3370 3416 3374
rect 3420 3370 3446 3374
rect 3450 3370 3483 3374
rect 3487 3370 3520 3374
rect 3524 3370 3548 3374
rect 3552 3370 3578 3374
rect 3582 3370 3615 3374
rect 3619 3370 3623 3374
rect 4026 3376 4031 3379
rect 4035 3376 4059 3379
rect 4084 3376 4091 3379
rect 4095 3376 4117 3379
rect 3226 3360 3229 3370
rect 3247 3360 3250 3370
rect 3263 3360 3266 3370
rect 3277 3363 3282 3367
rect 3286 3363 3293 3367
rect 3305 3360 3308 3370
rect 3321 3360 3324 3370
rect 3342 3360 3345 3370
rect 3358 3360 3361 3370
rect 3379 3360 3382 3370
rect 3395 3360 3398 3370
rect 3409 3363 3414 3367
rect 3418 3363 3425 3367
rect 3437 3360 3440 3370
rect 3453 3360 3456 3370
rect 3474 3360 3477 3370
rect 3490 3360 3493 3370
rect 3511 3360 3514 3370
rect 3527 3360 3530 3370
rect 3541 3363 3546 3367
rect 3550 3363 3557 3367
rect 3569 3360 3572 3370
rect 3585 3360 3588 3370
rect 3606 3360 3609 3370
rect 4042 3366 4049 3369
rect 4053 3370 4072 3373
rect 3064 3347 3067 3359
rect 3085 3347 3088 3359
rect 3101 3347 3104 3359
rect 3115 3350 3127 3353
rect 3143 3347 3146 3359
rect 3159 3347 3162 3359
rect 3180 3347 3183 3359
rect 2314 3336 2321 3339
rect 2325 3340 2344 3343
rect 2344 3333 2347 3339
rect 2372 3336 2379 3339
rect 2383 3340 2398 3343
rect 2446 3336 2453 3339
rect 2457 3340 2476 3343
rect 2476 3333 2479 3339
rect 2504 3336 2511 3339
rect 2515 3340 2530 3343
rect 2578 3336 2585 3339
rect 2589 3340 2608 3343
rect 2608 3333 2611 3339
rect 2636 3336 2643 3339
rect 2647 3340 2664 3343
rect 2696 3343 3094 3347
rect 3098 3343 3122 3347
rect 3126 3343 3152 3347
rect 3156 3343 3193 3347
rect 3243 3346 3248 3349
rect 3252 3346 3276 3349
rect 3301 3346 3308 3349
rect 3312 3346 3334 3349
rect 3354 3346 3361 3349
rect 3375 3346 3380 3349
rect 3384 3346 3408 3349
rect 3433 3346 3440 3349
rect 3444 3346 3466 3349
rect 3486 3346 3493 3349
rect 3507 3346 3512 3349
rect 3516 3346 3540 3349
rect 3565 3346 3572 3349
rect 3576 3346 3598 3349
rect 4072 3363 4075 3369
rect 4100 3366 4107 3369
rect 4111 3370 4126 3373
rect 4009 3347 4012 3359
rect 4030 3347 4033 3359
rect 4046 3347 4049 3359
rect 4060 3350 4072 3353
rect 4088 3347 4091 3359
rect 4104 3347 4107 3359
rect 4125 3347 4128 3359
rect 2732 3336 3070 3340
rect 3074 3336 3121 3340
rect 3125 3336 3171 3340
rect 3175 3336 3193 3340
rect 3259 3336 3266 3339
rect 3270 3340 3289 3343
rect 2281 3317 2284 3329
rect 2302 3317 2305 3329
rect 2318 3317 2321 3329
rect 2332 3320 2344 3323
rect 2360 3317 2363 3329
rect 2376 3317 2379 3329
rect 2397 3317 2400 3329
rect 2413 3317 2416 3329
rect 2434 3317 2437 3329
rect 2450 3317 2453 3329
rect 2464 3320 2476 3323
rect 2492 3317 2495 3329
rect 2508 3317 2511 3329
rect 2529 3317 2532 3329
rect 2545 3317 2548 3329
rect 2566 3317 2569 3329
rect 2582 3317 2585 3329
rect 2596 3320 2608 3323
rect 2624 3317 2627 3329
rect 2640 3317 2643 3329
rect 2661 3317 2664 3329
rect 3067 3329 3188 3332
rect 3289 3333 3292 3339
rect 3317 3336 3324 3339
rect 3328 3340 3343 3343
rect 3391 3336 3398 3339
rect 3402 3340 3421 3343
rect 3421 3333 3424 3339
rect 3449 3336 3456 3339
rect 3460 3340 3475 3343
rect 3523 3336 3530 3339
rect 3534 3340 3553 3343
rect 3553 3333 3556 3339
rect 3581 3336 3588 3339
rect 3592 3340 3609 3343
rect 3641 3343 4039 3347
rect 4043 3343 4067 3347
rect 4071 3343 4097 3347
rect 4101 3343 4138 3347
rect 3677 3336 4015 3340
rect 4019 3336 4066 3340
rect 4070 3336 4116 3340
rect 4120 3336 4138 3340
rect 2744 3321 3070 3325
rect 3074 3321 3106 3325
rect 3110 3321 3173 3325
rect 3177 3321 3193 3325
rect 2278 3313 2311 3317
rect 2315 3313 2339 3317
rect 2343 3313 2369 3317
rect 2373 3313 2443 3317
rect 2447 3313 2471 3317
rect 2475 3313 2501 3317
rect 2505 3313 2575 3317
rect 2579 3313 2603 3317
rect 2607 3313 2633 3317
rect 2637 3313 2690 3317
rect 3060 3314 3094 3318
rect 3098 3314 3122 3318
rect 3126 3314 3152 3318
rect 3156 3314 3189 3318
rect 3226 3317 3229 3329
rect 3247 3317 3250 3329
rect 3263 3317 3266 3329
rect 3277 3320 3289 3323
rect 3305 3317 3308 3329
rect 3321 3317 3324 3329
rect 3342 3317 3345 3329
rect 3358 3317 3361 3329
rect 3379 3317 3382 3329
rect 3395 3317 3398 3329
rect 3409 3320 3421 3323
rect 3437 3317 3440 3329
rect 3453 3317 3456 3329
rect 3474 3317 3477 3329
rect 3490 3317 3493 3329
rect 3511 3317 3514 3329
rect 3527 3317 3530 3329
rect 3541 3320 3553 3323
rect 3569 3317 3572 3329
rect 3585 3317 3588 3329
rect 3606 3317 3609 3329
rect 4012 3329 4133 3332
rect 3689 3321 4015 3325
rect 4019 3321 4051 3325
rect 4055 3321 4118 3325
rect 4122 3321 4138 3325
rect 2278 3306 2287 3310
rect 2291 3306 2338 3310
rect 2342 3306 2388 3310
rect 2392 3306 2419 3310
rect 2423 3306 2470 3310
rect 2474 3306 2520 3310
rect 2524 3306 2551 3310
rect 2555 3306 2602 3310
rect 2606 3306 2652 3310
rect 2656 3306 2726 3310
rect 3064 3304 3067 3314
rect 3085 3304 3088 3314
rect 3101 3304 3104 3314
rect 3115 3307 3120 3311
rect 3124 3307 3131 3311
rect 3143 3304 3146 3314
rect 3159 3304 3162 3314
rect 3180 3304 3183 3314
rect 3223 3313 3256 3317
rect 3260 3313 3284 3317
rect 3288 3313 3314 3317
rect 3318 3313 3388 3317
rect 3392 3313 3416 3317
rect 3420 3313 3446 3317
rect 3450 3313 3520 3317
rect 3524 3313 3548 3317
rect 3552 3313 3578 3317
rect 3582 3313 3635 3317
rect 4005 3314 4039 3318
rect 4043 3314 4067 3318
rect 4071 3314 4097 3318
rect 4101 3314 4134 3318
rect 3223 3306 3232 3310
rect 3236 3306 3283 3310
rect 3287 3306 3333 3310
rect 3337 3306 3364 3310
rect 3368 3306 3415 3310
rect 3419 3306 3465 3310
rect 3469 3306 3496 3310
rect 3500 3306 3547 3310
rect 3551 3306 3597 3310
rect 3601 3306 3671 3310
rect 4009 3304 4012 3314
rect 4030 3304 4033 3314
rect 4046 3304 4049 3314
rect 4060 3307 4065 3311
rect 4069 3307 4076 3311
rect 4088 3304 4091 3314
rect 4104 3304 4107 3314
rect 4125 3304 4128 3314
rect 2284 3299 2669 3302
rect 2278 3291 2287 3295
rect 2291 3291 2323 3295
rect 2327 3291 2390 3295
rect 2394 3291 2419 3295
rect 2423 3291 2455 3295
rect 2459 3291 2522 3295
rect 2526 3291 2551 3295
rect 2555 3291 2587 3295
rect 2591 3291 2654 3295
rect 2658 3291 2738 3295
rect 2278 3284 2311 3288
rect 2315 3284 2339 3288
rect 2343 3284 2369 3288
rect 2373 3284 2406 3288
rect 2410 3284 2443 3288
rect 2447 3284 2471 3288
rect 2475 3284 2501 3288
rect 2505 3284 2538 3288
rect 2542 3284 2575 3288
rect 2579 3284 2603 3288
rect 2607 3284 2633 3288
rect 2637 3284 2670 3288
rect 2674 3284 2678 3288
rect 3081 3290 3086 3293
rect 3090 3290 3114 3293
rect 3229 3299 3614 3302
rect 3139 3290 3146 3293
rect 3150 3290 3172 3293
rect 3223 3291 3232 3295
rect 3236 3291 3268 3295
rect 3272 3291 3335 3295
rect 3339 3291 3364 3295
rect 3368 3291 3400 3295
rect 3404 3291 3467 3295
rect 3471 3291 3496 3295
rect 3500 3291 3532 3295
rect 3536 3291 3599 3295
rect 3603 3291 3683 3295
rect 2281 3274 2284 3284
rect 2302 3274 2305 3284
rect 2318 3274 2321 3284
rect 2332 3277 2337 3281
rect 2341 3277 2348 3281
rect 2360 3274 2363 3284
rect 2376 3274 2379 3284
rect 2397 3274 2400 3284
rect 2413 3274 2416 3284
rect 2434 3274 2437 3284
rect 2450 3274 2453 3284
rect 2464 3277 2469 3281
rect 2473 3277 2480 3281
rect 2492 3274 2495 3284
rect 2508 3274 2511 3284
rect 2529 3274 2532 3284
rect 2545 3274 2548 3284
rect 2566 3274 2569 3284
rect 2582 3274 2585 3284
rect 2596 3277 2601 3281
rect 2605 3277 2612 3281
rect 2624 3274 2627 3284
rect 2640 3274 2643 3284
rect 2661 3274 2664 3284
rect 3097 3280 3104 3283
rect 3108 3284 3127 3287
rect 2298 3260 2303 3263
rect 2307 3260 2331 3263
rect 2356 3260 2363 3263
rect 2367 3260 2389 3263
rect 2409 3260 2416 3263
rect 2430 3260 2435 3263
rect 2439 3260 2463 3263
rect 2488 3260 2495 3263
rect 2499 3260 2521 3263
rect 2541 3260 2548 3263
rect 2562 3260 2567 3263
rect 2571 3260 2595 3263
rect 2620 3260 2627 3263
rect 2631 3260 2653 3263
rect 3127 3277 3130 3283
rect 3155 3280 3162 3283
rect 3166 3284 3181 3287
rect 3192 3282 3203 3286
rect 3223 3284 3256 3288
rect 3260 3284 3284 3288
rect 3288 3284 3314 3288
rect 3318 3284 3351 3288
rect 3355 3284 3388 3288
rect 3392 3284 3416 3288
rect 3420 3284 3446 3288
rect 3450 3284 3483 3288
rect 3487 3284 3520 3288
rect 3524 3284 3548 3288
rect 3552 3284 3578 3288
rect 3582 3284 3615 3288
rect 3619 3284 3623 3288
rect 4026 3290 4031 3293
rect 4035 3290 4059 3293
rect 4084 3290 4091 3293
rect 4095 3290 4117 3293
rect 3226 3274 3229 3284
rect 3247 3274 3250 3284
rect 3263 3274 3266 3284
rect 3277 3277 3282 3281
rect 3286 3277 3293 3281
rect 3305 3274 3308 3284
rect 3321 3274 3324 3284
rect 3342 3274 3345 3284
rect 3358 3274 3361 3284
rect 3379 3274 3382 3284
rect 3395 3274 3398 3284
rect 3409 3277 3414 3281
rect 3418 3277 3425 3281
rect 3437 3274 3440 3284
rect 3453 3274 3456 3284
rect 3474 3274 3477 3284
rect 3490 3274 3493 3284
rect 3511 3274 3514 3284
rect 3527 3274 3530 3284
rect 3541 3277 3546 3281
rect 3550 3277 3557 3281
rect 3569 3274 3572 3284
rect 3585 3274 3588 3284
rect 3606 3274 3609 3284
rect 4042 3280 4049 3283
rect 4053 3284 4072 3287
rect 3064 3261 3067 3273
rect 3085 3261 3088 3273
rect 3101 3261 3104 3273
rect 3115 3264 3127 3267
rect 3143 3261 3146 3273
rect 3159 3261 3162 3273
rect 3180 3261 3183 3273
rect 2314 3250 2321 3253
rect 2325 3254 2344 3257
rect 2344 3247 2347 3253
rect 2372 3250 2379 3253
rect 2383 3254 2398 3257
rect 2446 3250 2453 3253
rect 2457 3254 2476 3257
rect 2476 3247 2479 3253
rect 2504 3250 2511 3253
rect 2515 3254 2530 3257
rect 2578 3250 2585 3253
rect 2589 3254 2608 3257
rect 2608 3247 2611 3253
rect 2636 3250 2643 3253
rect 2647 3254 2664 3257
rect 2696 3257 3094 3261
rect 3098 3257 3122 3261
rect 3126 3257 3152 3261
rect 3156 3257 3193 3261
rect 3243 3260 3248 3263
rect 3252 3260 3276 3263
rect 3301 3260 3308 3263
rect 3312 3260 3334 3263
rect 3354 3260 3361 3263
rect 3375 3260 3380 3263
rect 3384 3260 3408 3263
rect 3433 3260 3440 3263
rect 3444 3260 3466 3263
rect 3486 3260 3493 3263
rect 3507 3260 3512 3263
rect 3516 3260 3540 3263
rect 3565 3260 3572 3263
rect 3576 3260 3598 3263
rect 4072 3277 4075 3283
rect 4100 3280 4107 3283
rect 4111 3284 4126 3287
rect 4137 3282 4148 3286
rect 4009 3261 4012 3273
rect 4030 3261 4033 3273
rect 4046 3261 4049 3273
rect 4060 3264 4072 3267
rect 4088 3261 4091 3273
rect 4104 3261 4107 3273
rect 4125 3261 4128 3273
rect 2732 3250 3070 3254
rect 3074 3250 3121 3254
rect 3125 3250 3171 3254
rect 3175 3250 3193 3254
rect 3259 3250 3266 3253
rect 3270 3254 3289 3257
rect 3289 3247 3292 3253
rect 3317 3250 3324 3253
rect 3328 3254 3343 3257
rect 3391 3250 3398 3253
rect 3402 3254 3421 3257
rect 3421 3247 3424 3253
rect 3449 3250 3456 3253
rect 3460 3254 3475 3257
rect 3523 3250 3530 3253
rect 3534 3254 3553 3257
rect 3553 3247 3556 3253
rect 3581 3250 3588 3253
rect 3592 3254 3609 3257
rect 3641 3257 4039 3261
rect 4043 3257 4067 3261
rect 4071 3257 4097 3261
rect 4101 3257 4138 3261
rect 3677 3250 4015 3254
rect 4019 3250 4066 3254
rect 4070 3250 4116 3254
rect 4120 3250 4138 3254
rect 2281 3231 2284 3243
rect 2302 3231 2305 3243
rect 2318 3231 2321 3243
rect 2332 3234 2344 3237
rect 2360 3231 2363 3243
rect 2376 3231 2379 3243
rect 2397 3231 2400 3243
rect 2413 3231 2416 3243
rect 2434 3231 2437 3243
rect 2450 3231 2453 3243
rect 2464 3234 2476 3237
rect 2492 3231 2495 3243
rect 2508 3231 2511 3243
rect 2529 3231 2532 3243
rect 2545 3231 2548 3243
rect 2566 3231 2569 3243
rect 2582 3231 2585 3243
rect 2596 3234 2608 3237
rect 2624 3231 2627 3243
rect 2640 3231 2643 3243
rect 2661 3231 2664 3243
rect 3226 3231 3229 3243
rect 3247 3231 3250 3243
rect 3263 3231 3266 3243
rect 3277 3234 3289 3237
rect 3305 3231 3308 3243
rect 3321 3231 3324 3243
rect 3342 3231 3345 3243
rect 3358 3231 3361 3243
rect 3379 3231 3382 3243
rect 3395 3231 3398 3243
rect 3409 3234 3421 3237
rect 3437 3231 3440 3243
rect 3453 3231 3456 3243
rect 3474 3231 3477 3243
rect 3490 3231 3493 3243
rect 3511 3231 3514 3243
rect 3527 3231 3530 3243
rect 3541 3234 3553 3237
rect 3569 3231 3572 3243
rect 3585 3231 3588 3243
rect 3606 3231 3609 3243
rect 2278 3227 2311 3231
rect 2315 3227 2339 3231
rect 2343 3227 2369 3231
rect 2373 3227 2443 3231
rect 2447 3227 2471 3231
rect 2475 3227 2501 3231
rect 2505 3227 2575 3231
rect 2579 3227 2603 3231
rect 2607 3227 2633 3231
rect 2637 3227 2690 3231
rect 3223 3227 3256 3231
rect 3260 3227 3284 3231
rect 3288 3227 3314 3231
rect 3318 3227 3388 3231
rect 3392 3227 3416 3231
rect 3420 3227 3446 3231
rect 3450 3227 3520 3231
rect 3524 3227 3548 3231
rect 3552 3227 3578 3231
rect 3582 3227 3635 3231
rect 2278 3220 2287 3224
rect 2291 3220 2338 3224
rect 2342 3220 2388 3224
rect 2392 3220 2419 3224
rect 2423 3220 2470 3224
rect 2474 3220 2520 3224
rect 2524 3220 2551 3224
rect 2555 3220 2602 3224
rect 2606 3220 2652 3224
rect 2656 3220 2726 3224
rect 3223 3220 3232 3224
rect 3236 3220 3283 3224
rect 3287 3220 3333 3224
rect 3337 3220 3364 3224
rect 3368 3220 3415 3224
rect 3419 3220 3465 3224
rect 3469 3220 3496 3224
rect 3500 3220 3547 3224
rect 3551 3220 3597 3224
rect 3601 3220 3671 3224
rect 2284 3214 2669 3217
rect 3229 3214 3614 3217
rect 2409 3207 2513 3210
rect 3354 3207 3458 3210
rect 2525 3199 2529 3203
rect 2533 3199 2537 3203
rect 3470 3199 3474 3203
rect 3478 3199 3482 3203
rect 2268 3188 2513 3192
rect 2517 3188 2533 3192
rect 2549 3188 3210 3192
rect 3214 3188 3458 3192
rect 3462 3188 3478 3192
rect 3494 3188 4155 3192
rect 4159 3188 4237 3192
rect 2541 3181 2669 3184
rect 3486 3181 3614 3184
rect 2556 3174 2669 3177
rect 3501 3174 3614 3177
rect 2525 3165 2529 3169
rect 2533 3165 2537 3169
rect 3470 3165 3474 3169
rect 3478 3165 3482 3169
rect 2409 3158 2513 3161
rect 3354 3158 3458 3161
rect 2278 3151 2287 3155
rect 2291 3151 2323 3155
rect 2327 3151 2390 3155
rect 2394 3151 2419 3155
rect 2423 3151 2455 3155
rect 2459 3151 2522 3155
rect 2526 3151 2551 3155
rect 2555 3151 2587 3155
rect 2591 3151 2654 3155
rect 2658 3151 2738 3155
rect 3223 3151 3232 3155
rect 3236 3151 3268 3155
rect 3272 3151 3335 3155
rect 3339 3151 3364 3155
rect 3368 3151 3400 3155
rect 3404 3151 3467 3155
rect 3471 3151 3496 3155
rect 3500 3151 3532 3155
rect 3536 3151 3599 3155
rect 3603 3151 3683 3155
rect 2278 3144 2311 3148
rect 2315 3144 2339 3148
rect 2343 3144 2369 3148
rect 2373 3144 2406 3148
rect 2410 3144 2443 3148
rect 2447 3144 2471 3148
rect 2475 3144 2501 3148
rect 2505 3144 2538 3148
rect 2542 3144 2575 3148
rect 2579 3144 2603 3148
rect 2607 3144 2633 3148
rect 2637 3144 2670 3148
rect 2674 3144 2678 3148
rect 3223 3144 3256 3148
rect 3260 3144 3284 3148
rect 3288 3144 3314 3148
rect 3318 3144 3351 3148
rect 3355 3144 3388 3148
rect 3392 3144 3416 3148
rect 3420 3144 3446 3148
rect 3450 3144 3483 3148
rect 3487 3144 3520 3148
rect 3524 3144 3548 3148
rect 3552 3144 3578 3148
rect 3582 3144 3615 3148
rect 3619 3144 3623 3148
rect 2281 3134 2284 3144
rect 2302 3134 2305 3144
rect 2318 3134 2321 3144
rect 2332 3137 2337 3141
rect 2341 3137 2348 3141
rect 2360 3134 2363 3144
rect 2376 3134 2379 3144
rect 2397 3134 2400 3144
rect 2413 3134 2416 3144
rect 2434 3134 2437 3144
rect 2450 3134 2453 3144
rect 2464 3137 2469 3141
rect 2473 3137 2480 3141
rect 2492 3134 2495 3144
rect 2508 3134 2511 3144
rect 2529 3134 2532 3144
rect 2545 3134 2548 3144
rect 2566 3134 2569 3144
rect 2582 3134 2585 3144
rect 2596 3137 2601 3141
rect 2605 3137 2612 3141
rect 2624 3134 2627 3144
rect 2640 3134 2643 3144
rect 2661 3134 2664 3144
rect 3226 3134 3229 3144
rect 3247 3134 3250 3144
rect 3263 3134 3266 3144
rect 3277 3137 3282 3141
rect 3286 3137 3293 3141
rect 3305 3134 3308 3144
rect 3321 3134 3324 3144
rect 3342 3134 3345 3144
rect 3358 3134 3361 3144
rect 3379 3134 3382 3144
rect 3395 3134 3398 3144
rect 3409 3137 3414 3141
rect 3418 3137 3425 3141
rect 3437 3134 3440 3144
rect 3453 3134 3456 3144
rect 3474 3134 3477 3144
rect 3490 3134 3493 3144
rect 3511 3134 3514 3144
rect 3527 3134 3530 3144
rect 3541 3137 3546 3141
rect 3550 3137 3557 3141
rect 3569 3134 3572 3144
rect 3585 3134 3588 3144
rect 3606 3134 3609 3144
rect 2298 3120 2303 3123
rect 2307 3120 2331 3123
rect 2356 3120 2363 3123
rect 2367 3120 2389 3123
rect 2409 3120 2416 3123
rect 2430 3120 2435 3123
rect 2439 3120 2463 3123
rect 2488 3120 2495 3123
rect 2499 3120 2521 3123
rect 2541 3120 2548 3123
rect 2562 3120 2567 3123
rect 2571 3120 2595 3123
rect 2620 3120 2627 3123
rect 2631 3120 2653 3123
rect 2314 3110 2321 3113
rect 2325 3114 2344 3117
rect 2344 3107 2347 3113
rect 2372 3110 2379 3113
rect 2383 3114 2398 3117
rect 2446 3110 2453 3113
rect 2457 3114 2476 3117
rect 2476 3107 2479 3113
rect 2504 3110 2511 3113
rect 2515 3114 2530 3117
rect 2578 3110 2585 3113
rect 2589 3114 2608 3117
rect 2608 3107 2611 3113
rect 2636 3110 2643 3113
rect 2647 3114 2664 3117
rect 3243 3120 3248 3123
rect 3252 3120 3276 3123
rect 3301 3120 3308 3123
rect 3312 3120 3334 3123
rect 3354 3120 3361 3123
rect 3375 3120 3380 3123
rect 3384 3120 3408 3123
rect 3433 3120 3440 3123
rect 3444 3120 3466 3123
rect 3486 3120 3493 3123
rect 3507 3120 3512 3123
rect 3516 3120 3540 3123
rect 3565 3120 3572 3123
rect 3576 3120 3598 3123
rect 3259 3110 3266 3113
rect 3270 3114 3289 3117
rect 3289 3107 3292 3113
rect 3317 3110 3324 3113
rect 3328 3114 3343 3117
rect 3391 3110 3398 3113
rect 3402 3114 3421 3117
rect 3421 3107 3424 3113
rect 3449 3110 3456 3113
rect 3460 3114 3475 3117
rect 3523 3110 3530 3113
rect 3534 3114 3553 3117
rect 3553 3107 3556 3113
rect 3581 3110 3588 3113
rect 3592 3114 3609 3117
rect 2281 3091 2284 3103
rect 2302 3091 2305 3103
rect 2318 3091 2321 3103
rect 2332 3094 2344 3097
rect 2360 3091 2363 3103
rect 2376 3091 2379 3103
rect 2397 3091 2400 3103
rect 2413 3091 2416 3103
rect 2434 3091 2437 3103
rect 2450 3091 2453 3103
rect 2464 3094 2476 3097
rect 2492 3091 2495 3103
rect 2508 3091 2511 3103
rect 2529 3091 2532 3103
rect 2545 3091 2548 3103
rect 2566 3091 2569 3103
rect 2582 3091 2585 3103
rect 2596 3094 2608 3097
rect 2624 3091 2627 3103
rect 2640 3091 2643 3103
rect 2661 3091 2664 3103
rect 3226 3091 3229 3103
rect 3247 3091 3250 3103
rect 3263 3091 3266 3103
rect 3277 3094 3289 3097
rect 3305 3091 3308 3103
rect 3321 3091 3324 3103
rect 3342 3091 3345 3103
rect 3358 3091 3361 3103
rect 3379 3091 3382 3103
rect 3395 3091 3398 3103
rect 3409 3094 3421 3097
rect 3437 3091 3440 3103
rect 3453 3091 3456 3103
rect 3474 3091 3477 3103
rect 3490 3091 3493 3103
rect 3511 3091 3514 3103
rect 3527 3091 3530 3103
rect 3541 3094 3553 3097
rect 3569 3091 3572 3103
rect 3585 3091 3588 3103
rect 3606 3091 3609 3103
rect 2278 3087 2311 3091
rect 2315 3087 2339 3091
rect 2343 3087 2369 3091
rect 2373 3087 2443 3091
rect 2447 3087 2471 3091
rect 2475 3087 2501 3091
rect 2505 3087 2575 3091
rect 2579 3087 2603 3091
rect 2607 3087 2633 3091
rect 2637 3087 2690 3091
rect 3223 3087 3256 3091
rect 3260 3087 3284 3091
rect 3288 3087 3314 3091
rect 3318 3087 3388 3091
rect 3392 3087 3416 3091
rect 3420 3087 3446 3091
rect 3450 3087 3520 3091
rect 3524 3087 3548 3091
rect 3552 3087 3578 3091
rect 3582 3087 3635 3091
rect 2278 3080 2287 3084
rect 2291 3080 2338 3084
rect 2342 3080 2388 3084
rect 2392 3080 2419 3084
rect 2423 3080 2470 3084
rect 2474 3080 2520 3084
rect 2524 3080 2551 3084
rect 2555 3080 2602 3084
rect 2606 3080 2652 3084
rect 2656 3080 2726 3084
rect 3223 3080 3232 3084
rect 3236 3080 3283 3084
rect 3287 3080 3333 3084
rect 3337 3080 3364 3084
rect 3368 3080 3415 3084
rect 3419 3080 3465 3084
rect 3469 3080 3496 3084
rect 3500 3080 3547 3084
rect 3551 3080 3597 3084
rect 3601 3080 3671 3084
rect 2744 3072 2771 3076
rect 2775 3072 2807 3076
rect 2811 3072 2874 3076
rect 2878 3072 2903 3076
rect 2907 3072 2939 3076
rect 2943 3072 3006 3076
rect 3010 3072 3035 3076
rect 3039 3072 3071 3076
rect 3075 3072 3138 3076
rect 3142 3072 3167 3076
rect 3171 3072 3203 3076
rect 3207 3072 3270 3076
rect 3274 3072 3290 3076
rect 3689 3072 3716 3076
rect 3720 3072 3752 3076
rect 3756 3072 3819 3076
rect 3823 3072 3848 3076
rect 3852 3072 3884 3076
rect 3888 3072 3951 3076
rect 3955 3072 3980 3076
rect 3984 3072 4016 3076
rect 4020 3072 4083 3076
rect 4087 3072 4112 3076
rect 4116 3072 4148 3076
rect 4152 3072 4215 3076
rect 4219 3072 4235 3076
rect 2684 3065 2795 3069
rect 2799 3065 2823 3069
rect 2827 3065 2853 3069
rect 2857 3065 2890 3069
rect 2894 3065 2927 3069
rect 2931 3065 2955 3069
rect 2959 3065 2985 3069
rect 2989 3065 3022 3069
rect 3026 3065 3059 3069
rect 3063 3065 3087 3069
rect 3091 3065 3117 3069
rect 3121 3065 3154 3069
rect 3158 3065 3191 3069
rect 3195 3065 3219 3069
rect 3223 3065 3249 3069
rect 3253 3065 3286 3069
rect 3629 3065 3740 3069
rect 3744 3065 3768 3069
rect 3772 3065 3798 3069
rect 3802 3065 3835 3069
rect 3839 3065 3872 3069
rect 3876 3065 3900 3069
rect 3904 3065 3930 3069
rect 3934 3065 3967 3069
rect 3971 3065 4004 3069
rect 4008 3065 4032 3069
rect 4036 3065 4062 3069
rect 4066 3065 4099 3069
rect 4103 3065 4136 3069
rect 4140 3065 4164 3069
rect 4168 3065 4194 3069
rect 4198 3065 4231 3069
rect 2765 3055 2768 3065
rect 2786 3055 2789 3065
rect 2802 3055 2805 3065
rect 2816 3058 2821 3062
rect 2825 3058 2832 3062
rect 2844 3055 2847 3065
rect 2860 3055 2863 3065
rect 2881 3055 2884 3065
rect 2897 3055 2900 3065
rect 2918 3055 2921 3065
rect 2934 3055 2937 3065
rect 2948 3058 2953 3062
rect 2957 3058 2964 3062
rect 2976 3055 2979 3065
rect 2992 3055 2995 3065
rect 3013 3055 3016 3065
rect 3029 3055 3032 3065
rect 3050 3055 3053 3065
rect 3066 3055 3069 3065
rect 3080 3058 3085 3062
rect 3089 3058 3096 3062
rect 3108 3055 3111 3065
rect 3124 3055 3127 3065
rect 3145 3055 3148 3065
rect 3161 3055 3164 3065
rect 3182 3055 3185 3065
rect 3198 3055 3201 3065
rect 3212 3058 3217 3062
rect 3221 3058 3228 3062
rect 3240 3055 3243 3065
rect 3256 3055 3259 3065
rect 3277 3055 3280 3065
rect 3710 3055 3713 3065
rect 3731 3055 3734 3065
rect 3747 3055 3750 3065
rect 3761 3058 3766 3062
rect 3770 3058 3777 3062
rect 3789 3055 3792 3065
rect 3805 3055 3808 3065
rect 3826 3055 3829 3065
rect 3842 3055 3845 3065
rect 3863 3055 3866 3065
rect 3879 3055 3882 3065
rect 3893 3058 3898 3062
rect 3902 3058 3909 3062
rect 3921 3055 3924 3065
rect 3937 3055 3940 3065
rect 3958 3055 3961 3065
rect 3974 3055 3977 3065
rect 3995 3055 3998 3065
rect 4011 3055 4014 3065
rect 4025 3058 4030 3062
rect 4034 3058 4041 3062
rect 4053 3055 4056 3065
rect 4069 3055 4072 3065
rect 4090 3055 4093 3065
rect 4106 3055 4109 3065
rect 4127 3055 4130 3065
rect 4143 3055 4146 3065
rect 4157 3058 4162 3062
rect 4166 3058 4173 3062
rect 4185 3055 4188 3065
rect 4201 3055 4204 3065
rect 4222 3055 4225 3065
rect 2410 3039 2419 3043
rect 2423 3039 2455 3043
rect 2459 3039 2522 3043
rect 2526 3039 2738 3043
rect 2782 3041 2787 3044
rect 2791 3041 2815 3044
rect 2840 3041 2847 3044
rect 2851 3041 2873 3044
rect 2410 3032 2443 3036
rect 2447 3032 2471 3036
rect 2475 3032 2501 3036
rect 2505 3032 2538 3036
rect 2542 3032 2678 3036
rect 2413 3022 2416 3032
rect 2434 3022 2437 3032
rect 2450 3022 2453 3032
rect 2464 3025 2469 3029
rect 2473 3025 2480 3029
rect 2492 3022 2495 3032
rect 2508 3022 2511 3032
rect 2529 3022 2532 3032
rect 2798 3031 2805 3034
rect 2809 3035 2828 3038
rect 2828 3028 2831 3034
rect 2856 3031 2863 3034
rect 2867 3035 2884 3038
rect 2914 3041 2919 3044
rect 2923 3041 2947 3044
rect 2972 3041 2979 3044
rect 2983 3041 3005 3044
rect 2930 3031 2937 3034
rect 2941 3035 2960 3038
rect 2960 3028 2963 3034
rect 2988 3031 2995 3034
rect 2999 3035 3016 3038
rect 3046 3041 3051 3044
rect 3055 3041 3079 3044
rect 3104 3041 3111 3044
rect 3115 3041 3137 3044
rect 3062 3031 3069 3034
rect 3073 3035 3092 3038
rect 3092 3028 3095 3034
rect 3120 3031 3127 3034
rect 3131 3035 3148 3038
rect 3178 3041 3183 3044
rect 3187 3041 3211 3044
rect 3236 3041 3243 3044
rect 3247 3041 3269 3044
rect 3355 3039 3364 3043
rect 3368 3039 3400 3043
rect 3404 3039 3467 3043
rect 3471 3039 3683 3043
rect 3194 3031 3201 3034
rect 3205 3035 3224 3038
rect 2408 3005 2417 3009
rect 2430 3008 2435 3011
rect 2439 3008 2463 3011
rect 2488 3008 2495 3011
rect 2499 3008 2521 3011
rect 2765 3012 2768 3024
rect 2786 3012 2789 3024
rect 2802 3012 2805 3024
rect 2816 3015 2828 3018
rect 2844 3012 2847 3024
rect 2860 3012 2863 3024
rect 2881 3012 2884 3024
rect 2897 3012 2900 3024
rect 2918 3012 2921 3024
rect 2934 3012 2937 3024
rect 2948 3015 2960 3018
rect 2976 3012 2979 3024
rect 2992 3012 2995 3024
rect 3013 3012 3016 3024
rect 3029 3012 3032 3024
rect 3050 3012 3053 3024
rect 3066 3012 3069 3024
rect 3080 3015 3092 3018
rect 3108 3012 3111 3024
rect 3124 3012 3127 3024
rect 3145 3012 3148 3024
rect 3224 3028 3227 3034
rect 3252 3031 3259 3034
rect 3263 3035 3280 3038
rect 3727 3041 3732 3044
rect 3736 3041 3760 3044
rect 3785 3041 3792 3044
rect 3796 3041 3818 3044
rect 3355 3032 3388 3036
rect 3392 3032 3416 3036
rect 3420 3032 3446 3036
rect 3450 3032 3483 3036
rect 3487 3032 3623 3036
rect 3161 3012 3164 3024
rect 3182 3012 3185 3024
rect 3198 3012 3201 3024
rect 3212 3015 3224 3018
rect 3240 3012 3243 3024
rect 3256 3012 3259 3024
rect 3277 3012 3280 3024
rect 3358 3022 3361 3032
rect 3379 3022 3382 3032
rect 3395 3022 3398 3032
rect 3409 3025 3414 3029
rect 3418 3025 3425 3029
rect 3437 3022 3440 3032
rect 3453 3022 3456 3032
rect 3474 3022 3477 3032
rect 3743 3031 3750 3034
rect 3754 3035 3773 3038
rect 3773 3028 3776 3034
rect 3801 3031 3808 3034
rect 3812 3035 3829 3038
rect 3859 3041 3864 3044
rect 3868 3041 3892 3044
rect 3917 3041 3924 3044
rect 3928 3041 3950 3044
rect 3875 3031 3882 3034
rect 3886 3035 3905 3038
rect 3905 3028 3908 3034
rect 3933 3031 3940 3034
rect 3944 3035 3961 3038
rect 3991 3041 3996 3044
rect 4000 3041 4024 3044
rect 4049 3041 4056 3044
rect 4060 3041 4082 3044
rect 4007 3031 4014 3034
rect 4018 3035 4037 3038
rect 4037 3028 4040 3034
rect 4065 3031 4072 3034
rect 4076 3035 4093 3038
rect 4123 3041 4128 3044
rect 4132 3041 4156 3044
rect 4181 3041 4188 3044
rect 4192 3041 4214 3044
rect 4139 3031 4146 3034
rect 4150 3035 4169 3038
rect 2696 3008 2795 3012
rect 2799 3008 2823 3012
rect 2827 3008 2853 3012
rect 2857 3008 2927 3012
rect 2931 3008 2955 3012
rect 2959 3008 2985 3012
rect 2989 3008 3059 3012
rect 3063 3008 3087 3012
rect 3091 3008 3117 3012
rect 3121 3008 3191 3012
rect 3195 3008 3219 3012
rect 3223 3008 3249 3012
rect 3253 3008 3290 3012
rect 2446 2998 2453 3001
rect 2457 3002 2476 3005
rect 2476 2995 2479 3001
rect 2504 2998 2511 3001
rect 2515 3002 2530 3005
rect 3353 3005 3362 3009
rect 3375 3008 3380 3011
rect 3384 3008 3408 3011
rect 3433 3008 3440 3011
rect 3444 3008 3466 3011
rect 3710 3012 3713 3024
rect 3731 3012 3734 3024
rect 3747 3012 3750 3024
rect 3761 3015 3773 3018
rect 3789 3012 3792 3024
rect 3805 3012 3808 3024
rect 3826 3012 3829 3024
rect 3842 3012 3845 3024
rect 3863 3012 3866 3024
rect 3879 3012 3882 3024
rect 3893 3015 3905 3018
rect 3921 3012 3924 3024
rect 3937 3012 3940 3024
rect 3958 3012 3961 3024
rect 3974 3012 3977 3024
rect 3995 3012 3998 3024
rect 4011 3012 4014 3024
rect 4025 3015 4037 3018
rect 4053 3012 4056 3024
rect 4069 3012 4072 3024
rect 4090 3012 4093 3024
rect 4169 3028 4172 3034
rect 4197 3031 4204 3034
rect 4208 3035 4225 3038
rect 4106 3012 4109 3024
rect 4127 3012 4130 3024
rect 4143 3012 4146 3024
rect 4157 3015 4169 3018
rect 4185 3012 4188 3024
rect 4201 3012 4204 3024
rect 4222 3012 4225 3024
rect 3641 3008 3740 3012
rect 3744 3008 3768 3012
rect 3772 3008 3798 3012
rect 3802 3008 3872 3012
rect 3876 3008 3900 3012
rect 3904 3008 3930 3012
rect 3934 3008 4004 3012
rect 4008 3008 4032 3012
rect 4036 3008 4062 3012
rect 4066 3008 4136 3012
rect 4140 3008 4164 3012
rect 4168 3008 4194 3012
rect 4198 3008 4235 3012
rect 2732 3001 2771 3005
rect 2775 3001 2822 3005
rect 2826 3001 2872 3005
rect 2876 3001 2903 3005
rect 2907 3001 2954 3005
rect 2958 3001 3004 3005
rect 3008 3001 3035 3005
rect 3039 3001 3086 3005
rect 3090 3001 3136 3005
rect 3140 3001 3167 3005
rect 3171 3001 3218 3005
rect 3222 3001 3268 3005
rect 3272 3001 3290 3005
rect 3391 2998 3398 3001
rect 3402 3002 3421 3005
rect 2413 2979 2416 2991
rect 2434 2979 2437 2991
rect 2450 2979 2453 2991
rect 2464 2982 2476 2985
rect 2492 2979 2495 2991
rect 2508 2979 2511 2991
rect 2529 2979 2532 2991
rect 2684 2988 2769 2992
rect 2773 2988 2785 2992
rect 2789 2988 2803 2992
rect 2807 2988 2814 2992
rect 2818 2988 2820 2992
rect 2824 2988 2839 2992
rect 2843 2988 2876 2992
rect 2880 2988 2881 2992
rect 2885 2988 2893 2992
rect 2897 2988 2921 2992
rect 2925 2988 2937 2992
rect 2941 2988 2961 2992
rect 2965 2988 3015 2992
rect 3019 2988 3042 2992
rect 3046 2988 3096 2992
rect 3100 2988 3119 2992
rect 3421 2995 3424 3001
rect 3449 2998 3456 3001
rect 3460 3002 3475 3005
rect 3677 3001 3716 3005
rect 3720 3001 3767 3005
rect 3771 3001 3817 3005
rect 3821 3001 3848 3005
rect 3852 3001 3899 3005
rect 3903 3001 3949 3005
rect 3953 3001 3980 3005
rect 3984 3001 4031 3005
rect 4035 3001 4081 3005
rect 4085 3001 4112 3005
rect 4116 3001 4163 3005
rect 4167 3001 4213 3005
rect 4217 3001 4235 3005
rect 2720 2981 2796 2985
rect 2800 2981 2827 2985
rect 2831 2981 2849 2985
rect 2853 2981 2914 2985
rect 2918 2981 2932 2985
rect 2944 2984 2947 2988
rect 2410 2975 2443 2979
rect 2447 2975 2471 2979
rect 2475 2975 2501 2979
rect 2505 2975 2690 2979
rect 2410 2968 2419 2972
rect 2423 2968 2470 2972
rect 2474 2968 2520 2972
rect 2524 2968 2726 2972
rect 2839 2974 2842 2978
rect 2866 2974 2867 2978
rect 2911 2974 2913 2978
rect 2953 2971 2956 2976
rect 2968 2978 2971 2988
rect 2998 2984 3001 2988
rect 3025 2984 3028 2988
rect 2408 2952 2424 2956
rect 2533 2954 2537 2958
rect 2549 2954 2553 2958
rect 2557 2954 2763 2958
rect 2767 2954 2771 2958
rect 2779 2957 2782 2963
rect 2786 2957 2789 2963
rect 2779 2954 2789 2957
rect 2779 2949 2782 2954
rect 2416 2945 2420 2949
rect 2432 2945 2553 2949
rect 2786 2949 2789 2954
rect 2795 2959 2798 2963
rect 2795 2955 2797 2959
rect 2801 2955 2803 2959
rect 2811 2958 2814 2963
rect 2839 2960 2842 2963
rect 2811 2956 2822 2958
rect 2795 2949 2798 2955
rect 2811 2954 2817 2956
rect 2811 2949 2814 2954
rect 2821 2954 2822 2956
rect 2840 2956 2842 2960
rect 2839 2949 2842 2956
rect 2942 2967 2945 2970
rect 2984 2967 2987 2970
rect 2855 2959 2858 2963
rect 2865 2959 2868 2963
rect 2865 2955 2874 2959
rect 2886 2958 2889 2963
rect 2911 2959 2914 2963
rect 2855 2949 2858 2955
rect 2865 2949 2868 2955
rect 2886 2954 2887 2958
rect 2891 2954 2894 2957
rect 2913 2955 2914 2959
rect 2929 2958 2932 2963
rect 2953 2962 2956 2967
rect 2961 2963 2972 2966
rect 2984 2964 2992 2967
rect 2886 2949 2889 2954
rect 2911 2949 2914 2955
rect 2929 2949 2932 2954
rect 2403 2937 2419 2941
rect 2423 2937 2486 2941
rect 2490 2937 2522 2941
rect 2526 2937 2738 2941
rect 2831 2936 2832 2940
rect 2856 2937 2857 2941
rect 2903 2936 2904 2940
rect 2407 2930 2440 2934
rect 2444 2930 2470 2934
rect 2474 2930 2498 2934
rect 2502 2930 2678 2934
rect 2413 2920 2416 2930
rect 2434 2920 2437 2930
rect 2450 2920 2453 2930
rect 2465 2923 2472 2927
rect 2476 2923 2481 2927
rect 2492 2920 2495 2930
rect 2508 2920 2511 2930
rect 2529 2920 2532 2930
rect 2708 2929 2784 2933
rect 2788 2929 2843 2933
rect 2847 2929 2868 2933
rect 2872 2929 2899 2933
rect 2903 2929 2932 2933
rect 2944 2926 2947 2958
rect 2961 2957 2964 2963
rect 2984 2958 2987 2964
rect 2996 2959 2999 2962
rect 3007 2962 3010 2976
rect 3034 2971 3037 2976
rect 3049 2978 3052 2988
rect 3079 2984 3082 2988
rect 3018 2967 3019 2970
rect 3023 2967 3026 2970
rect 3358 2979 3361 2991
rect 3379 2979 3382 2991
rect 3395 2979 3398 2991
rect 3409 2982 3421 2985
rect 3437 2979 3440 2991
rect 3453 2979 3456 2991
rect 3474 2979 3477 2991
rect 3629 2988 3714 2992
rect 3718 2988 3730 2992
rect 3734 2988 3748 2992
rect 3752 2988 3759 2992
rect 3763 2988 3765 2992
rect 3769 2988 3784 2992
rect 3788 2988 3821 2992
rect 3825 2988 3826 2992
rect 3830 2988 3838 2992
rect 3842 2988 3866 2992
rect 3870 2988 3882 2992
rect 3886 2988 3906 2992
rect 3910 2988 3960 2992
rect 3964 2988 3987 2992
rect 3991 2988 4041 2992
rect 4045 2988 4064 2992
rect 3665 2981 3741 2985
rect 3745 2981 3772 2985
rect 3776 2981 3794 2985
rect 3798 2981 3859 2985
rect 3863 2981 3877 2985
rect 3889 2984 3892 2988
rect 3065 2967 3068 2970
rect 3007 2959 3015 2962
rect 3034 2962 3037 2967
rect 3007 2954 3010 2959
rect 3015 2955 3019 2959
rect 3042 2963 3053 2966
rect 3065 2964 3073 2967
rect 2959 2948 2964 2953
rect 2968 2926 2971 2954
rect 2998 2926 3001 2950
rect 3025 2926 3028 2958
rect 3042 2957 3045 2963
rect 3065 2958 3068 2964
rect 3077 2959 3080 2962
rect 3088 2962 3091 2976
rect 3355 2975 3388 2979
rect 3392 2975 3416 2979
rect 3420 2975 3446 2979
rect 3450 2975 3635 2979
rect 3355 2968 3364 2972
rect 3368 2968 3415 2972
rect 3419 2968 3465 2972
rect 3469 2968 3671 2972
rect 3784 2974 3787 2978
rect 3811 2974 3812 2978
rect 3856 2974 3858 2978
rect 3898 2971 3901 2976
rect 3913 2978 3916 2988
rect 3943 2984 3946 2988
rect 3970 2984 3973 2988
rect 3088 2959 3100 2962
rect 3088 2954 3091 2959
rect 3040 2948 3045 2953
rect 3049 2926 3052 2954
rect 3353 2952 3369 2956
rect 3478 2954 3482 2958
rect 3494 2954 3498 2958
rect 3502 2954 3708 2958
rect 3712 2954 3716 2958
rect 3724 2957 3727 2963
rect 3731 2957 3734 2963
rect 3724 2954 3734 2957
rect 3079 2926 3082 2950
rect 3724 2949 3727 2954
rect 3361 2945 3365 2949
rect 3377 2945 3498 2949
rect 3731 2949 3734 2954
rect 3740 2959 3743 2963
rect 3740 2955 3742 2959
rect 3746 2955 3748 2959
rect 3756 2958 3759 2963
rect 3784 2960 3787 2963
rect 3756 2956 3767 2958
rect 3740 2949 3743 2955
rect 3756 2954 3762 2956
rect 3756 2949 3759 2954
rect 3766 2954 3767 2956
rect 3785 2956 3787 2960
rect 3784 2949 3787 2956
rect 3887 2967 3890 2970
rect 3929 2967 3932 2970
rect 3800 2959 3803 2963
rect 3810 2959 3813 2963
rect 3810 2955 3819 2959
rect 3831 2958 3834 2963
rect 3856 2959 3859 2963
rect 3800 2949 3803 2955
rect 3810 2949 3813 2955
rect 3831 2954 3832 2958
rect 3836 2954 3839 2957
rect 3858 2955 3859 2959
rect 3874 2958 3877 2963
rect 3898 2962 3901 2967
rect 3906 2963 3917 2966
rect 3929 2964 3937 2967
rect 3831 2949 3834 2954
rect 3856 2949 3859 2955
rect 3874 2949 3877 2954
rect 3348 2937 3364 2941
rect 3368 2937 3431 2941
rect 3435 2937 3467 2941
rect 3471 2937 3683 2941
rect 3776 2936 3777 2940
rect 3801 2937 3802 2941
rect 3848 2936 3849 2940
rect 3352 2930 3385 2934
rect 3389 2930 3415 2934
rect 3419 2930 3443 2934
rect 3447 2930 3623 2934
rect 2696 2922 2770 2926
rect 2774 2922 2776 2926
rect 2780 2922 2784 2926
rect 2788 2922 2802 2926
rect 2806 2922 2811 2926
rect 2815 2922 2820 2926
rect 2824 2922 2843 2926
rect 2847 2922 2877 2926
rect 2881 2922 2892 2926
rect 2896 2922 2920 2926
rect 2924 2922 2937 2926
rect 2941 2922 2961 2926
rect 2965 2922 3015 2926
rect 3022 2922 3042 2926
rect 3046 2922 3096 2926
rect 2424 2906 2446 2909
rect 2450 2906 2457 2909
rect 2708 2915 2784 2919
rect 2788 2915 2843 2919
rect 2847 2915 2868 2919
rect 2872 2915 2899 2919
rect 2903 2915 2932 2919
rect 2482 2906 2506 2909
rect 2510 2906 2515 2909
rect 2831 2908 2832 2912
rect 2856 2907 2857 2911
rect 2903 2908 2904 2912
rect 2528 2903 2537 2907
rect 2415 2900 2430 2903
rect 2469 2900 2488 2903
rect 2434 2896 2441 2899
rect 2466 2893 2469 2899
rect 2492 2896 2499 2899
rect 2779 2894 2782 2899
rect 2786 2894 2789 2899
rect 2769 2891 2771 2894
rect 2779 2891 2789 2894
rect 2413 2877 2416 2889
rect 2434 2877 2437 2889
rect 2450 2877 2453 2889
rect 2469 2880 2481 2883
rect 2492 2877 2495 2889
rect 2508 2877 2511 2889
rect 2529 2877 2532 2889
rect 2779 2885 2782 2891
rect 2786 2885 2789 2891
rect 2795 2893 2798 2899
rect 2811 2894 2814 2899
rect 2795 2889 2797 2893
rect 2801 2889 2803 2893
rect 2811 2892 2817 2894
rect 2821 2892 2822 2894
rect 2811 2890 2822 2892
rect 2839 2892 2842 2899
rect 2795 2885 2798 2889
rect 2811 2885 2814 2890
rect 2840 2888 2842 2892
rect 2839 2885 2842 2888
rect 2855 2893 2858 2899
rect 2865 2893 2868 2899
rect 2886 2894 2889 2899
rect 2865 2889 2874 2893
rect 2886 2890 2887 2894
rect 2891 2891 2894 2894
rect 2911 2893 2914 2899
rect 2929 2894 2932 2899
rect 2968 2902 2971 2922
rect 3049 2902 3052 2922
rect 3358 2920 3361 2930
rect 3379 2920 3382 2930
rect 3395 2920 3398 2930
rect 3410 2923 3417 2927
rect 3421 2923 3426 2927
rect 3437 2920 3440 2930
rect 3453 2920 3456 2930
rect 3474 2920 3477 2930
rect 3653 2929 3729 2933
rect 3733 2929 3788 2933
rect 3792 2929 3813 2933
rect 3817 2929 3844 2933
rect 3848 2929 3877 2933
rect 3889 2926 3892 2958
rect 3906 2957 3909 2963
rect 3929 2958 3932 2964
rect 3941 2959 3944 2962
rect 3952 2962 3955 2976
rect 3979 2971 3982 2976
rect 3994 2978 3997 2988
rect 4024 2984 4027 2988
rect 3963 2967 3964 2970
rect 3968 2967 3971 2970
rect 4010 2967 4013 2970
rect 3952 2959 3960 2962
rect 3979 2962 3982 2967
rect 3952 2954 3955 2959
rect 3960 2955 3964 2959
rect 3987 2963 3998 2966
rect 4010 2964 4018 2967
rect 3904 2948 3909 2953
rect 3913 2926 3916 2954
rect 3943 2926 3946 2950
rect 3970 2926 3973 2958
rect 3987 2957 3990 2963
rect 4010 2958 4013 2964
rect 4022 2959 4025 2962
rect 4033 2962 4036 2976
rect 4033 2959 4045 2962
rect 4033 2954 4036 2959
rect 3985 2948 3990 2953
rect 3994 2926 3997 2954
rect 4024 2926 4027 2950
rect 3641 2922 3715 2926
rect 3719 2922 3721 2926
rect 3725 2922 3729 2926
rect 3733 2922 3747 2926
rect 3751 2922 3756 2926
rect 3760 2922 3765 2926
rect 3769 2922 3788 2926
rect 3792 2922 3822 2926
rect 3826 2922 3837 2926
rect 3841 2922 3865 2926
rect 3869 2922 3882 2926
rect 3886 2922 3906 2926
rect 3910 2922 3960 2926
rect 3967 2922 3987 2926
rect 3991 2922 4041 2926
rect 3369 2906 3391 2909
rect 3395 2906 3402 2909
rect 3653 2915 3729 2919
rect 3733 2915 3788 2919
rect 3792 2915 3813 2919
rect 3817 2915 3844 2919
rect 3848 2915 3877 2919
rect 3427 2906 3451 2909
rect 3455 2906 3460 2909
rect 3776 2908 3777 2912
rect 3801 2907 3802 2911
rect 3848 2908 3849 2912
rect 3473 2903 3482 2907
rect 3360 2900 3375 2903
rect 2855 2885 2858 2889
rect 2865 2885 2868 2889
rect 2886 2885 2889 2890
rect 2913 2889 2914 2893
rect 2911 2885 2914 2889
rect 2929 2885 2932 2890
rect 2959 2889 2964 2894
rect 2968 2890 2969 2893
rect 2984 2892 2987 2898
rect 2984 2889 2992 2892
rect 3039 2889 3044 2894
rect 3048 2890 3050 2893
rect 3065 2892 3068 2898
rect 3414 2900 3433 2903
rect 3379 2896 3386 2899
rect 3411 2893 3414 2899
rect 3065 2889 3073 2892
rect 3437 2896 3444 2899
rect 3724 2894 3727 2899
rect 3731 2894 3734 2899
rect 3714 2891 3716 2894
rect 3724 2891 3734 2894
rect 2984 2886 2987 2889
rect 3065 2886 3068 2889
rect 2403 2873 2440 2877
rect 2444 2873 2470 2877
rect 2474 2873 2498 2877
rect 2502 2873 2690 2877
rect 2839 2870 2842 2874
rect 2866 2870 2867 2874
rect 2911 2870 2913 2874
rect 2403 2866 2421 2870
rect 2425 2866 2471 2870
rect 2475 2866 2522 2870
rect 2526 2866 2726 2870
rect 2784 2863 2796 2867
rect 2800 2863 2827 2867
rect 2831 2863 2849 2867
rect 2853 2863 2914 2867
rect 2918 2863 2932 2867
rect 2968 2860 2971 2878
rect 3049 2860 3052 2878
rect 3358 2877 3361 2889
rect 3379 2877 3382 2889
rect 3395 2877 3398 2889
rect 3414 2880 3426 2883
rect 3437 2877 3440 2889
rect 3453 2877 3456 2889
rect 3474 2877 3477 2889
rect 3724 2885 3727 2891
rect 3731 2885 3734 2891
rect 3740 2893 3743 2899
rect 3756 2894 3759 2899
rect 3740 2889 3742 2893
rect 3746 2889 3748 2893
rect 3756 2892 3762 2894
rect 3766 2892 3767 2894
rect 3756 2890 3767 2892
rect 3784 2892 3787 2899
rect 3740 2885 3743 2889
rect 3756 2885 3759 2890
rect 3785 2888 3787 2892
rect 3784 2885 3787 2888
rect 3800 2893 3803 2899
rect 3810 2893 3813 2899
rect 3831 2894 3834 2899
rect 3810 2889 3819 2893
rect 3831 2890 3832 2894
rect 3836 2891 3839 2894
rect 3856 2893 3859 2899
rect 3874 2894 3877 2899
rect 3913 2902 3916 2922
rect 3994 2902 3997 2922
rect 3800 2885 3803 2889
rect 3810 2885 3813 2889
rect 3831 2885 3834 2890
rect 3858 2889 3859 2893
rect 3856 2885 3859 2889
rect 3874 2885 3877 2890
rect 3904 2889 3909 2894
rect 3913 2890 3914 2893
rect 3929 2892 3932 2898
rect 3929 2889 3937 2892
rect 3984 2889 3989 2894
rect 3993 2890 3995 2893
rect 4010 2892 4013 2898
rect 4010 2889 4018 2892
rect 3929 2886 3932 2889
rect 4010 2886 4013 2889
rect 3348 2873 3385 2877
rect 3389 2873 3415 2877
rect 3419 2873 3443 2877
rect 3447 2873 3635 2877
rect 3784 2870 3787 2874
rect 3811 2870 3812 2874
rect 3856 2870 3858 2874
rect 3348 2866 3366 2870
rect 3370 2866 3416 2870
rect 3420 2866 3467 2870
rect 3471 2866 3671 2870
rect 3729 2863 3741 2867
rect 3745 2863 3772 2867
rect 3776 2863 3794 2867
rect 3798 2863 3859 2867
rect 3863 2863 3877 2867
rect 3913 2860 3916 2878
rect 3994 2860 3997 2878
rect 2684 2856 2769 2860
rect 2773 2856 2785 2860
rect 2789 2856 2803 2860
rect 2807 2856 2814 2860
rect 2818 2856 2820 2860
rect 2824 2856 2839 2860
rect 2843 2856 2876 2860
rect 2880 2856 2881 2860
rect 2885 2856 2893 2860
rect 2897 2856 2921 2860
rect 2925 2856 2937 2860
rect 2941 2856 2961 2860
rect 2965 2856 3015 2860
rect 3019 2856 3042 2860
rect 3046 2856 3104 2860
rect 3108 2856 3119 2860
rect 3629 2856 3714 2860
rect 3718 2856 3730 2860
rect 3734 2856 3748 2860
rect 3752 2856 3759 2860
rect 3763 2856 3765 2860
rect 3769 2856 3784 2860
rect 3788 2856 3821 2860
rect 3825 2856 3826 2860
rect 3830 2856 3838 2860
rect 3842 2856 3866 2860
rect 3870 2856 3882 2860
rect 3886 2856 3906 2860
rect 3910 2856 3960 2860
rect 3964 2856 3987 2860
rect 3991 2856 4049 2860
rect 4053 2856 4064 2860
rect 2720 2849 2780 2853
rect 2784 2849 2796 2853
rect 2800 2849 2827 2853
rect 2831 2849 2849 2853
rect 2853 2849 2914 2853
rect 2918 2849 2932 2853
rect 2968 2846 2971 2856
rect 2998 2852 3001 2856
rect 3049 2852 3052 2856
rect 2839 2842 2842 2846
rect 2866 2842 2867 2846
rect 2911 2842 2913 2846
rect 2768 2822 2771 2825
rect 2779 2825 2782 2831
rect 2786 2825 2789 2831
rect 2779 2822 2789 2825
rect 2779 2817 2782 2822
rect 2786 2817 2789 2822
rect 2795 2827 2798 2831
rect 2795 2823 2797 2827
rect 2801 2823 2803 2827
rect 2811 2826 2814 2831
rect 2839 2828 2842 2831
rect 2811 2824 2822 2826
rect 2795 2817 2798 2823
rect 2811 2822 2817 2824
rect 2811 2817 2814 2822
rect 2821 2822 2822 2824
rect 2840 2824 2842 2828
rect 2839 2817 2842 2824
rect 2984 2835 2987 2838
rect 2855 2827 2858 2831
rect 2865 2827 2868 2831
rect 2865 2823 2874 2827
rect 2886 2826 2889 2831
rect 2911 2827 2914 2831
rect 2855 2817 2858 2823
rect 2865 2817 2868 2823
rect 2886 2822 2887 2826
rect 2891 2822 2894 2825
rect 2913 2823 2914 2827
rect 2929 2826 2932 2831
rect 2961 2831 2972 2834
rect 2984 2832 2992 2835
rect 2886 2817 2889 2822
rect 2911 2817 2914 2823
rect 2961 2825 2964 2831
rect 2984 2826 2987 2832
rect 2996 2827 2999 2830
rect 3007 2830 3010 2844
rect 3058 2839 3061 2844
rect 3073 2846 3076 2856
rect 3103 2852 3106 2856
rect 3042 2835 3043 2838
rect 3047 2835 3050 2838
rect 3665 2849 3725 2853
rect 3729 2849 3741 2853
rect 3745 2849 3772 2853
rect 3776 2849 3794 2853
rect 3798 2849 3859 2853
rect 3863 2849 3877 2853
rect 3913 2846 3916 2856
rect 3943 2852 3946 2856
rect 3994 2852 3997 2856
rect 3089 2835 3092 2838
rect 3015 2830 3020 2835
rect 3058 2830 3061 2835
rect 3007 2827 3015 2830
rect 2929 2817 2932 2822
rect 3007 2822 3010 2827
rect 3066 2831 3077 2834
rect 3089 2832 3097 2835
rect 2959 2816 2964 2821
rect 2831 2804 2832 2808
rect 2856 2805 2857 2809
rect 2903 2804 2904 2808
rect 2708 2797 2784 2801
rect 2788 2797 2843 2801
rect 2847 2797 2868 2801
rect 2872 2797 2899 2801
rect 2903 2797 2932 2801
rect 2968 2794 2971 2822
rect 2998 2794 3001 2818
rect 3049 2794 3052 2826
rect 3066 2825 3069 2831
rect 3089 2826 3092 2832
rect 3101 2827 3104 2830
rect 3112 2830 3115 2844
rect 3784 2842 3787 2846
rect 3811 2842 3812 2846
rect 3856 2842 3858 2846
rect 3112 2827 3118 2830
rect 3112 2822 3115 2827
rect 3713 2822 3716 2825
rect 3724 2825 3727 2831
rect 3731 2825 3734 2831
rect 3724 2822 3734 2825
rect 3064 2816 3069 2821
rect 3073 2794 3076 2822
rect 3103 2794 3106 2818
rect 3724 2817 3727 2822
rect 3731 2817 3734 2822
rect 3740 2827 3743 2831
rect 3740 2823 3742 2827
rect 3746 2823 3748 2827
rect 3756 2826 3759 2831
rect 3784 2828 3787 2831
rect 3756 2824 3767 2826
rect 3740 2817 3743 2823
rect 3756 2822 3762 2824
rect 3756 2817 3759 2822
rect 3766 2822 3767 2824
rect 3785 2824 3787 2828
rect 3784 2817 3787 2824
rect 3929 2835 3932 2838
rect 3800 2827 3803 2831
rect 3810 2827 3813 2831
rect 3810 2823 3819 2827
rect 3831 2826 3834 2831
rect 3856 2827 3859 2831
rect 3800 2817 3803 2823
rect 3810 2817 3813 2823
rect 3831 2822 3832 2826
rect 3836 2822 3839 2825
rect 3858 2823 3859 2827
rect 3874 2826 3877 2831
rect 3906 2831 3917 2834
rect 3929 2832 3937 2835
rect 3831 2817 3834 2822
rect 3856 2817 3859 2823
rect 3906 2825 3909 2831
rect 3929 2826 3932 2832
rect 3941 2827 3944 2830
rect 3952 2830 3955 2844
rect 4003 2839 4006 2844
rect 4018 2846 4021 2856
rect 4048 2852 4051 2856
rect 3987 2835 3988 2838
rect 3992 2835 3995 2838
rect 4034 2835 4037 2838
rect 3960 2830 3965 2835
rect 4003 2830 4006 2835
rect 3952 2827 3960 2830
rect 3874 2817 3877 2822
rect 3952 2822 3955 2827
rect 4011 2831 4022 2834
rect 4034 2832 4042 2835
rect 3904 2816 3909 2821
rect 3776 2804 3777 2808
rect 3801 2805 3802 2809
rect 3848 2804 3849 2808
rect 3653 2797 3729 2801
rect 3733 2797 3788 2801
rect 3792 2797 3813 2801
rect 3817 2797 3844 2801
rect 3848 2797 3877 2801
rect 3913 2794 3916 2822
rect 3943 2794 3946 2818
rect 3994 2794 3997 2826
rect 4011 2825 4014 2831
rect 4034 2826 4037 2832
rect 4046 2827 4049 2830
rect 4057 2830 4060 2844
rect 4057 2827 4063 2830
rect 4057 2822 4060 2827
rect 4009 2816 4014 2821
rect 4018 2794 4021 2822
rect 4048 2794 4051 2818
rect 2696 2790 2770 2794
rect 2774 2790 2776 2794
rect 2780 2790 2784 2794
rect 2788 2790 2802 2794
rect 2806 2790 2811 2794
rect 2815 2790 2820 2794
rect 2824 2790 2843 2794
rect 2847 2790 2877 2794
rect 2881 2790 2892 2794
rect 2896 2790 2920 2794
rect 2924 2790 2937 2794
rect 2941 2790 2961 2794
rect 2965 2790 3015 2794
rect 3019 2790 3042 2794
rect 3046 2790 3066 2794
rect 3070 2790 3118 2794
rect 3641 2790 3715 2794
rect 3719 2790 3721 2794
rect 3725 2790 3729 2794
rect 3733 2790 3747 2794
rect 3751 2790 3756 2794
rect 3760 2790 3765 2794
rect 3769 2790 3788 2794
rect 3792 2790 3822 2794
rect 3826 2790 3837 2794
rect 3841 2790 3865 2794
rect 3869 2790 3882 2794
rect 3886 2790 3906 2794
rect 3910 2790 3960 2794
rect 3964 2790 3987 2794
rect 3991 2790 4011 2794
rect 4015 2790 4063 2794
rect 2708 2783 2784 2787
rect 2788 2783 2843 2787
rect 2847 2783 2868 2787
rect 2872 2783 2899 2787
rect 2903 2783 2932 2787
rect 2831 2776 2832 2780
rect 2856 2775 2857 2779
rect 2903 2776 2904 2780
rect 2968 2771 2971 2790
rect 3073 2771 3076 2790
rect 3653 2783 3729 2787
rect 3733 2783 3788 2787
rect 3792 2783 3813 2787
rect 3817 2783 3844 2787
rect 3848 2783 3877 2787
rect 3776 2776 3777 2780
rect 3801 2775 3802 2779
rect 3848 2776 3849 2780
rect 3913 2771 3916 2790
rect 4018 2771 4021 2790
rect 2779 2762 2782 2767
rect 2786 2762 2789 2767
rect 2769 2759 2771 2762
rect 2779 2759 2789 2762
rect 2779 2753 2782 2759
rect 2786 2753 2789 2759
rect 2795 2761 2798 2767
rect 2811 2762 2814 2767
rect 2795 2757 2797 2761
rect 2801 2757 2803 2761
rect 2811 2760 2817 2762
rect 2821 2760 2822 2762
rect 2811 2758 2822 2760
rect 2839 2760 2842 2767
rect 2795 2753 2798 2757
rect 2811 2753 2814 2758
rect 2840 2756 2842 2760
rect 2839 2753 2842 2756
rect 2855 2761 2858 2767
rect 2865 2761 2868 2767
rect 2886 2762 2889 2767
rect 2865 2757 2874 2761
rect 2886 2758 2887 2762
rect 2891 2759 2894 2762
rect 2911 2761 2914 2767
rect 2929 2762 2932 2767
rect 2855 2753 2858 2757
rect 2865 2753 2868 2757
rect 2886 2753 2889 2758
rect 2913 2757 2914 2761
rect 2958 2758 2963 2763
rect 2967 2759 2969 2762
rect 2984 2761 2987 2767
rect 2984 2758 2992 2761
rect 3064 2758 3069 2763
rect 3073 2759 3074 2762
rect 3089 2761 3092 2767
rect 3089 2758 3097 2761
rect 3724 2762 3727 2767
rect 3731 2762 3734 2767
rect 3714 2759 3716 2762
rect 3724 2759 3734 2762
rect 2911 2753 2914 2757
rect 2929 2753 2932 2758
rect 2984 2755 2987 2758
rect 3089 2755 3092 2758
rect 3724 2753 3727 2759
rect 2839 2738 2842 2742
rect 2866 2738 2867 2742
rect 2911 2738 2913 2742
rect 2720 2731 2796 2735
rect 2800 2731 2827 2735
rect 2831 2731 2849 2735
rect 2853 2731 2914 2735
rect 2918 2731 2932 2735
rect 2968 2728 2971 2747
rect 3073 2728 3076 2747
rect 3731 2753 3734 2759
rect 3740 2761 3743 2767
rect 3756 2762 3759 2767
rect 3740 2757 3742 2761
rect 3746 2757 3748 2761
rect 3756 2760 3762 2762
rect 3766 2760 3767 2762
rect 3756 2758 3767 2760
rect 3784 2760 3787 2767
rect 3740 2753 3743 2757
rect 3756 2753 3759 2758
rect 3785 2756 3787 2760
rect 3784 2753 3787 2756
rect 3800 2761 3803 2767
rect 3810 2761 3813 2767
rect 3831 2762 3834 2767
rect 3810 2757 3819 2761
rect 3831 2758 3832 2762
rect 3836 2759 3839 2762
rect 3856 2761 3859 2767
rect 3874 2762 3877 2767
rect 3800 2753 3803 2757
rect 3810 2753 3813 2757
rect 3831 2753 3834 2758
rect 3858 2757 3859 2761
rect 3903 2758 3908 2763
rect 3912 2759 3914 2762
rect 3929 2761 3932 2767
rect 3929 2758 3937 2761
rect 4009 2758 4014 2763
rect 4018 2759 4019 2762
rect 4034 2761 4037 2767
rect 4034 2758 4042 2761
rect 3856 2753 3859 2757
rect 3874 2753 3877 2758
rect 3929 2755 3932 2758
rect 4034 2755 4037 2758
rect 3784 2738 3787 2742
rect 3811 2738 3812 2742
rect 3856 2738 3858 2742
rect 3665 2731 3741 2735
rect 3745 2731 3772 2735
rect 3776 2731 3794 2735
rect 3798 2731 3859 2735
rect 3863 2731 3877 2735
rect 3913 2728 3916 2747
rect 4018 2728 4021 2747
rect 2684 2724 2769 2728
rect 2773 2724 2785 2728
rect 2789 2724 2803 2728
rect 2807 2724 2814 2728
rect 2818 2724 2820 2728
rect 2824 2724 2839 2728
rect 2843 2724 2876 2728
rect 2880 2724 2881 2728
rect 2885 2724 2893 2728
rect 2897 2724 2921 2728
rect 2925 2724 2937 2728
rect 2941 2724 2961 2728
rect 2965 2724 3015 2728
rect 3019 2724 3042 2728
rect 3046 2724 3096 2728
rect 3100 2724 3104 2728
rect 3108 2724 3132 2728
rect 3136 2724 3186 2728
rect 3629 2724 3714 2728
rect 3718 2724 3730 2728
rect 3734 2724 3748 2728
rect 3752 2724 3759 2728
rect 3763 2724 3765 2728
rect 3769 2724 3784 2728
rect 3788 2724 3821 2728
rect 3825 2724 3826 2728
rect 3830 2724 3838 2728
rect 3842 2724 3866 2728
rect 3870 2724 3882 2728
rect 3886 2724 3906 2728
rect 3910 2724 3960 2728
rect 3964 2724 3987 2728
rect 3991 2724 4041 2728
rect 4045 2724 4049 2728
rect 4053 2724 4077 2728
rect 4081 2724 4131 2728
rect 2720 2717 2796 2721
rect 2800 2717 2827 2721
rect 2831 2717 2849 2721
rect 2853 2717 2914 2721
rect 2918 2717 2932 2721
rect 2968 2714 2971 2724
rect 2998 2720 3001 2724
rect 3025 2720 3028 2724
rect 2839 2710 2842 2714
rect 2866 2710 2867 2714
rect 2911 2710 2913 2714
rect 2768 2690 2771 2693
rect 2779 2693 2782 2699
rect 2786 2693 2789 2699
rect 2779 2690 2789 2693
rect 2779 2685 2782 2690
rect 2786 2685 2789 2690
rect 2795 2695 2798 2699
rect 2795 2691 2797 2695
rect 2801 2691 2803 2695
rect 2811 2694 2814 2699
rect 2839 2696 2842 2699
rect 2811 2692 2822 2694
rect 2795 2685 2798 2691
rect 2811 2690 2817 2692
rect 2811 2685 2814 2690
rect 2821 2690 2822 2692
rect 2840 2692 2842 2696
rect 2839 2685 2842 2692
rect 2984 2703 2987 2706
rect 2855 2695 2858 2699
rect 2865 2695 2868 2699
rect 2865 2691 2874 2695
rect 2886 2694 2889 2699
rect 2911 2695 2914 2699
rect 2855 2685 2858 2691
rect 2865 2685 2868 2691
rect 2886 2690 2887 2694
rect 2891 2690 2894 2693
rect 2913 2691 2914 2695
rect 2929 2694 2932 2699
rect 2961 2699 2972 2702
rect 2984 2700 2992 2703
rect 2886 2685 2889 2690
rect 2911 2685 2914 2691
rect 2961 2693 2964 2699
rect 2984 2694 2987 2700
rect 2996 2695 2999 2698
rect 3007 2698 3010 2712
rect 3034 2707 3037 2712
rect 3049 2714 3052 2724
rect 3079 2720 3082 2724
rect 3115 2720 3118 2724
rect 3018 2703 3019 2706
rect 3023 2703 3026 2706
rect 3065 2703 3068 2706
rect 3007 2695 3015 2698
rect 3034 2698 3037 2703
rect 2929 2685 2932 2690
rect 3007 2690 3010 2695
rect 3015 2691 3019 2695
rect 3042 2699 3053 2702
rect 3065 2700 3073 2703
rect 2959 2684 2964 2689
rect 2831 2672 2832 2676
rect 2856 2673 2857 2677
rect 2903 2672 2904 2676
rect 2708 2665 2784 2669
rect 2788 2665 2843 2669
rect 2847 2665 2868 2669
rect 2872 2665 2899 2669
rect 2903 2665 2932 2669
rect 2968 2662 2971 2690
rect 2998 2662 3001 2686
rect 3025 2662 3028 2694
rect 3042 2693 3045 2699
rect 3065 2694 3068 2700
rect 3077 2695 3080 2698
rect 3088 2698 3091 2712
rect 3124 2707 3127 2712
rect 3139 2714 3142 2724
rect 3169 2720 3172 2724
rect 3113 2703 3116 2706
rect 3665 2717 3741 2721
rect 3745 2717 3772 2721
rect 3776 2717 3794 2721
rect 3798 2717 3859 2721
rect 3863 2717 3877 2721
rect 3913 2714 3916 2724
rect 3943 2720 3946 2724
rect 3970 2720 3973 2724
rect 3155 2703 3158 2706
rect 3088 2695 3097 2698
rect 3124 2698 3127 2703
rect 3088 2690 3091 2695
rect 3040 2684 3045 2689
rect 3049 2662 3052 2690
rect 3131 2701 3143 2702
rect 3135 2699 3143 2701
rect 3155 2700 3163 2703
rect 3155 2694 3158 2700
rect 3167 2695 3170 2698
rect 3178 2698 3181 2712
rect 3784 2710 3787 2714
rect 3811 2710 3812 2714
rect 3856 2710 3858 2714
rect 3178 2695 3198 2698
rect 3079 2662 3082 2686
rect 3115 2662 3118 2694
rect 3178 2690 3181 2695
rect 3713 2690 3716 2693
rect 3724 2693 3727 2699
rect 3731 2693 3734 2699
rect 3724 2690 3734 2693
rect 3139 2662 3142 2690
rect 3169 2662 3172 2686
rect 3724 2685 3727 2690
rect 3731 2685 3734 2690
rect 3740 2695 3743 2699
rect 3740 2691 3742 2695
rect 3746 2691 3748 2695
rect 3756 2694 3759 2699
rect 3784 2696 3787 2699
rect 3756 2692 3767 2694
rect 3740 2685 3743 2691
rect 3756 2690 3762 2692
rect 3756 2685 3759 2690
rect 3766 2690 3767 2692
rect 3785 2692 3787 2696
rect 3784 2685 3787 2692
rect 3929 2703 3932 2706
rect 3800 2695 3803 2699
rect 3810 2695 3813 2699
rect 3810 2691 3819 2695
rect 3831 2694 3834 2699
rect 3856 2695 3859 2699
rect 3800 2685 3803 2691
rect 3810 2685 3813 2691
rect 3831 2690 3832 2694
rect 3836 2690 3839 2693
rect 3858 2691 3859 2695
rect 3874 2694 3877 2699
rect 3906 2699 3917 2702
rect 3929 2700 3937 2703
rect 3831 2685 3834 2690
rect 3856 2685 3859 2691
rect 3906 2693 3909 2699
rect 3929 2694 3932 2700
rect 3941 2695 3944 2698
rect 3952 2698 3955 2712
rect 3979 2707 3982 2712
rect 3994 2714 3997 2724
rect 4024 2720 4027 2724
rect 4060 2720 4063 2724
rect 3963 2703 3964 2706
rect 3968 2703 3971 2706
rect 4010 2703 4013 2706
rect 3952 2695 3960 2698
rect 3979 2698 3982 2703
rect 3874 2685 3877 2690
rect 3952 2690 3955 2695
rect 3960 2691 3964 2695
rect 3987 2699 3998 2702
rect 4010 2700 4018 2703
rect 3904 2684 3909 2689
rect 3776 2672 3777 2676
rect 3801 2673 3802 2677
rect 3848 2672 3849 2676
rect 3653 2665 3729 2669
rect 3733 2665 3788 2669
rect 3792 2665 3813 2669
rect 3817 2665 3844 2669
rect 3848 2665 3877 2669
rect 3913 2662 3916 2690
rect 3943 2662 3946 2686
rect 3970 2662 3973 2694
rect 3987 2693 3990 2699
rect 4010 2694 4013 2700
rect 4022 2695 4025 2698
rect 4033 2698 4036 2712
rect 4069 2707 4072 2712
rect 4084 2714 4087 2724
rect 4114 2720 4117 2724
rect 4058 2703 4061 2706
rect 4100 2703 4103 2706
rect 4033 2695 4042 2698
rect 4069 2698 4072 2703
rect 4033 2690 4036 2695
rect 3985 2684 3990 2689
rect 3994 2662 3997 2690
rect 4076 2701 4088 2702
rect 4080 2699 4088 2701
rect 4100 2700 4108 2703
rect 4100 2694 4103 2700
rect 4112 2695 4115 2698
rect 4123 2698 4126 2712
rect 4242 2698 4291 2699
rect 4123 2695 4143 2698
rect 4024 2662 4027 2686
rect 4060 2662 4063 2694
rect 4123 2690 4126 2695
rect 4147 2694 4291 2698
rect 4084 2662 4087 2690
rect 4114 2662 4117 2686
rect 2696 2658 2770 2662
rect 2774 2658 2776 2662
rect 2780 2658 2784 2662
rect 2788 2658 2802 2662
rect 2806 2658 2811 2662
rect 2815 2658 2820 2662
rect 2824 2658 2843 2662
rect 2847 2658 2877 2662
rect 2881 2658 2892 2662
rect 2896 2658 2920 2662
rect 2924 2658 2937 2662
rect 2941 2658 2961 2662
rect 2965 2658 3015 2662
rect 3022 2658 3042 2662
rect 3046 2658 3096 2662
rect 3100 2658 3132 2662
rect 3136 2658 3186 2662
rect 3641 2658 3715 2662
rect 3719 2658 3721 2662
rect 3725 2658 3729 2662
rect 3733 2658 3747 2662
rect 3751 2658 3756 2662
rect 3760 2658 3765 2662
rect 3769 2658 3788 2662
rect 3792 2658 3822 2662
rect 3826 2658 3837 2662
rect 3841 2658 3865 2662
rect 3869 2658 3882 2662
rect 3886 2658 3906 2662
rect 3910 2658 3960 2662
rect 3967 2658 3987 2662
rect 3991 2658 4041 2662
rect 4045 2658 4077 2662
rect 4081 2658 4131 2662
rect 2708 2651 2784 2655
rect 2788 2651 2843 2655
rect 2847 2651 2868 2655
rect 2872 2651 2899 2655
rect 2903 2651 2932 2655
rect 2831 2644 2832 2648
rect 2856 2643 2857 2647
rect 2903 2644 2904 2648
rect 2779 2630 2782 2635
rect 2786 2630 2789 2635
rect 2769 2627 2771 2630
rect 2779 2627 2789 2630
rect 2779 2621 2782 2627
rect 2786 2621 2789 2627
rect 2795 2629 2798 2635
rect 2811 2630 2814 2635
rect 2795 2625 2797 2629
rect 2801 2625 2803 2629
rect 2811 2628 2817 2630
rect 2821 2628 2822 2630
rect 2811 2626 2822 2628
rect 2839 2628 2842 2635
rect 2795 2621 2798 2625
rect 2811 2621 2814 2626
rect 2840 2624 2842 2628
rect 2839 2621 2842 2624
rect 2855 2629 2858 2635
rect 2865 2629 2868 2635
rect 2886 2630 2889 2635
rect 2865 2625 2874 2629
rect 2886 2626 2887 2630
rect 2891 2627 2894 2630
rect 2911 2629 2914 2635
rect 2929 2630 2932 2635
rect 2968 2636 2971 2658
rect 3049 2636 3052 2658
rect 3139 2636 3142 2658
rect 3653 2651 3729 2655
rect 3733 2651 3788 2655
rect 3792 2651 3813 2655
rect 3817 2651 3844 2655
rect 3848 2651 3877 2655
rect 3776 2644 3777 2648
rect 3801 2643 3802 2647
rect 3848 2644 3849 2648
rect 2855 2621 2858 2625
rect 2865 2621 2868 2625
rect 2886 2621 2889 2626
rect 2913 2625 2914 2629
rect 2911 2621 2914 2625
rect 2929 2621 2932 2626
rect 2959 2623 2964 2628
rect 2968 2624 2969 2627
rect 2984 2626 2987 2632
rect 2984 2623 2992 2626
rect 3039 2623 3044 2628
rect 3048 2624 3050 2627
rect 3065 2626 3068 2632
rect 3065 2623 3073 2626
rect 3132 2624 3140 2627
rect 3155 2626 3158 2632
rect 3724 2630 3727 2635
rect 3731 2630 3734 2635
rect 3714 2627 3716 2630
rect 3155 2623 3163 2626
rect 3724 2627 3734 2630
rect 2984 2620 2987 2623
rect 3065 2620 3068 2623
rect 3155 2620 3158 2623
rect 3724 2621 3727 2627
rect 2839 2606 2842 2610
rect 2866 2606 2867 2610
rect 2911 2606 2913 2610
rect 3731 2621 3734 2627
rect 3740 2629 3743 2635
rect 3756 2630 3759 2635
rect 3740 2625 3742 2629
rect 3746 2625 3748 2629
rect 3756 2628 3762 2630
rect 3766 2628 3767 2630
rect 3756 2626 3767 2628
rect 3784 2628 3787 2635
rect 3740 2621 3743 2625
rect 3756 2621 3759 2626
rect 3785 2624 3787 2628
rect 3784 2621 3787 2624
rect 3800 2629 3803 2635
rect 3810 2629 3813 2635
rect 3831 2630 3834 2635
rect 3810 2625 3819 2629
rect 3831 2626 3832 2630
rect 3836 2627 3839 2630
rect 3856 2629 3859 2635
rect 3874 2630 3877 2635
rect 3913 2636 3916 2658
rect 3994 2636 3997 2658
rect 4084 2636 4087 2658
rect 4300 2657 4341 2670
rect 3800 2621 3803 2625
rect 3810 2621 3813 2625
rect 3831 2621 3834 2626
rect 3858 2625 3859 2629
rect 3856 2621 3859 2625
rect 3874 2621 3877 2626
rect 3904 2623 3909 2628
rect 3913 2624 3914 2627
rect 3929 2626 3932 2632
rect 3929 2623 3937 2626
rect 3984 2623 3989 2628
rect 3993 2624 3995 2627
rect 4010 2626 4013 2632
rect 4010 2623 4018 2626
rect 4077 2624 4085 2627
rect 4100 2626 4103 2632
rect 4100 2623 4108 2626
rect 3929 2620 3932 2623
rect 4010 2620 4013 2623
rect 4100 2620 4103 2623
rect 2720 2599 2796 2603
rect 2800 2599 2827 2603
rect 2831 2599 2849 2603
rect 2853 2599 2914 2603
rect 2918 2599 2932 2603
rect 2968 2596 2971 2612
rect 3049 2596 3052 2612
rect 3139 2596 3142 2612
rect 3784 2606 3787 2610
rect 3811 2606 3812 2610
rect 3856 2606 3858 2610
rect 3665 2599 3741 2603
rect 3745 2599 3772 2603
rect 3776 2599 3794 2603
rect 3798 2599 3859 2603
rect 3863 2599 3877 2603
rect 3913 2596 3916 2612
rect 3994 2596 3997 2612
rect 4084 2596 4087 2612
rect 2684 2592 2769 2596
rect 2773 2592 2785 2596
rect 2789 2592 2803 2596
rect 2807 2592 2814 2596
rect 2818 2592 2820 2596
rect 2824 2592 2839 2596
rect 2843 2592 2876 2596
rect 2880 2592 2881 2596
rect 2885 2592 2893 2596
rect 2897 2592 2921 2596
rect 2925 2592 2937 2596
rect 2941 2592 2961 2596
rect 2965 2592 3015 2596
rect 3019 2592 3042 2596
rect 3046 2592 3132 2596
rect 3136 2592 3190 2596
rect 3629 2592 3714 2596
rect 3718 2592 3730 2596
rect 3734 2592 3748 2596
rect 3752 2592 3759 2596
rect 3763 2592 3765 2596
rect 3769 2592 3784 2596
rect 3788 2592 3821 2596
rect 3825 2592 3826 2596
rect 3830 2592 3838 2596
rect 3842 2592 3866 2596
rect 3870 2592 3882 2596
rect 3886 2592 3906 2596
rect 3910 2592 3960 2596
rect 3964 2592 3987 2596
rect 3991 2592 4077 2596
rect 4081 2592 4135 2596
rect 2720 2585 2796 2589
rect 2800 2585 2827 2589
rect 2831 2585 2849 2589
rect 2853 2585 2914 2589
rect 2918 2585 2932 2589
rect 2968 2582 2971 2592
rect 2998 2588 3001 2592
rect 2839 2578 2842 2582
rect 2866 2578 2867 2582
rect 2911 2578 2913 2582
rect 2768 2558 2771 2561
rect 2779 2561 2782 2567
rect 2786 2561 2789 2567
rect 2779 2558 2789 2561
rect 2779 2553 2782 2558
rect 2786 2553 2789 2558
rect 2795 2563 2798 2567
rect 2795 2559 2797 2563
rect 2801 2559 2803 2563
rect 2811 2562 2814 2567
rect 2839 2564 2842 2567
rect 2811 2560 2822 2562
rect 2795 2553 2798 2559
rect 2811 2558 2817 2560
rect 2811 2553 2814 2558
rect 2821 2558 2822 2560
rect 2840 2560 2842 2564
rect 2839 2553 2842 2560
rect 3665 2585 3741 2589
rect 3745 2585 3772 2589
rect 3776 2585 3794 2589
rect 3798 2585 3859 2589
rect 3863 2585 3877 2589
rect 3913 2582 3916 2592
rect 3943 2588 3946 2592
rect 2984 2571 2987 2574
rect 2855 2563 2858 2567
rect 2865 2563 2868 2567
rect 2865 2559 2874 2563
rect 2886 2562 2889 2567
rect 2911 2563 2914 2567
rect 2855 2553 2858 2559
rect 2865 2553 2868 2559
rect 2886 2558 2887 2562
rect 2891 2558 2894 2561
rect 2913 2559 2914 2563
rect 2929 2562 2932 2567
rect 2961 2567 2972 2570
rect 2984 2568 2992 2571
rect 2886 2553 2889 2558
rect 2911 2553 2914 2559
rect 2961 2561 2964 2567
rect 2984 2562 2987 2568
rect 2996 2563 2999 2566
rect 3007 2566 3010 2580
rect 3784 2578 3787 2582
rect 3811 2578 3812 2582
rect 3856 2578 3858 2582
rect 3015 2566 3020 2571
rect 3007 2563 3015 2566
rect 2929 2553 2932 2558
rect 3007 2558 3010 2563
rect 3713 2558 3716 2561
rect 3724 2561 3727 2567
rect 3731 2561 3734 2567
rect 3724 2558 3734 2561
rect 2959 2552 2964 2557
rect 2278 2537 2287 2541
rect 2291 2537 2323 2541
rect 2327 2537 2390 2541
rect 2394 2537 2419 2541
rect 2423 2537 2455 2541
rect 2459 2537 2522 2541
rect 2526 2537 2551 2541
rect 2555 2537 2587 2541
rect 2591 2537 2654 2541
rect 2658 2537 2738 2541
rect 2831 2540 2832 2544
rect 2856 2541 2857 2545
rect 2903 2540 2904 2544
rect 2278 2530 2311 2534
rect 2315 2530 2339 2534
rect 2343 2530 2369 2534
rect 2373 2530 2406 2534
rect 2410 2530 2443 2534
rect 2447 2530 2471 2534
rect 2475 2530 2501 2534
rect 2505 2530 2538 2534
rect 2542 2530 2575 2534
rect 2579 2530 2603 2534
rect 2607 2530 2633 2534
rect 2637 2530 2670 2534
rect 2674 2530 2678 2534
rect 2763 2533 2784 2537
rect 2788 2533 2793 2537
rect 2797 2533 2843 2537
rect 2847 2533 2868 2537
rect 2872 2533 2899 2537
rect 2903 2533 2932 2537
rect 2968 2530 2971 2558
rect 2998 2530 3001 2554
rect 3724 2553 3727 2558
rect 3731 2553 3734 2558
rect 3740 2563 3743 2567
rect 3740 2559 3742 2563
rect 3746 2559 3748 2563
rect 3756 2562 3759 2567
rect 3784 2564 3787 2567
rect 3756 2560 3767 2562
rect 3740 2553 3743 2559
rect 3756 2558 3762 2560
rect 3756 2553 3759 2558
rect 3766 2558 3767 2560
rect 3785 2560 3787 2564
rect 3784 2553 3787 2560
rect 3929 2571 3932 2574
rect 3800 2563 3803 2567
rect 3810 2563 3813 2567
rect 3810 2559 3819 2563
rect 3831 2562 3834 2567
rect 3856 2563 3859 2567
rect 3800 2553 3803 2559
rect 3810 2553 3813 2559
rect 3831 2558 3832 2562
rect 3836 2558 3839 2561
rect 3858 2559 3859 2563
rect 3874 2562 3877 2567
rect 3906 2567 3917 2570
rect 3929 2568 3937 2571
rect 3831 2553 3834 2558
rect 3856 2553 3859 2559
rect 3906 2561 3909 2567
rect 3929 2562 3932 2568
rect 3941 2563 3944 2566
rect 3952 2566 3955 2580
rect 3960 2566 3965 2571
rect 3952 2563 3960 2566
rect 3874 2553 3877 2558
rect 3952 2558 3955 2563
rect 3904 2552 3909 2557
rect 3223 2537 3232 2541
rect 3236 2537 3268 2541
rect 3272 2537 3335 2541
rect 3339 2537 3364 2541
rect 3368 2537 3400 2541
rect 3404 2537 3467 2541
rect 3471 2537 3496 2541
rect 3500 2537 3532 2541
rect 3536 2537 3599 2541
rect 3603 2537 3683 2541
rect 3776 2540 3777 2544
rect 3801 2541 3802 2545
rect 3848 2540 3849 2544
rect 3223 2530 3256 2534
rect 3260 2530 3284 2534
rect 3288 2530 3314 2534
rect 3318 2530 3351 2534
rect 3355 2530 3388 2534
rect 3392 2530 3416 2534
rect 3420 2530 3446 2534
rect 3450 2530 3483 2534
rect 3487 2530 3520 2534
rect 3524 2530 3548 2534
rect 3552 2530 3578 2534
rect 3582 2530 3615 2534
rect 3619 2530 3623 2534
rect 3708 2533 3729 2537
rect 3733 2533 3738 2537
rect 3742 2533 3788 2537
rect 3792 2533 3813 2537
rect 3817 2533 3844 2537
rect 3848 2533 3877 2537
rect 3913 2530 3916 2558
rect 3943 2530 3946 2554
rect 2281 2520 2284 2530
rect 2302 2520 2305 2530
rect 2318 2520 2321 2530
rect 2332 2523 2337 2527
rect 2341 2523 2348 2527
rect 2360 2520 2363 2530
rect 2376 2520 2379 2530
rect 2397 2520 2400 2530
rect 2413 2520 2416 2530
rect 2434 2520 2437 2530
rect 2450 2520 2453 2530
rect 2464 2523 2469 2527
rect 2473 2523 2480 2527
rect 2492 2520 2495 2530
rect 2508 2520 2511 2530
rect 2529 2520 2532 2530
rect 2545 2520 2548 2530
rect 2566 2520 2569 2530
rect 2582 2520 2585 2530
rect 2596 2523 2601 2527
rect 2605 2523 2612 2527
rect 2624 2520 2627 2530
rect 2640 2520 2643 2530
rect 2661 2520 2664 2530
rect 2696 2526 2770 2530
rect 2774 2526 2776 2530
rect 2780 2526 2784 2530
rect 2788 2526 2802 2530
rect 2806 2526 2811 2530
rect 2815 2526 2820 2530
rect 2824 2526 2843 2530
rect 2847 2526 2877 2530
rect 2881 2526 2892 2530
rect 2896 2526 2920 2530
rect 2924 2526 2937 2530
rect 2941 2526 2961 2530
rect 2965 2526 3045 2530
rect 3049 2526 3063 2530
rect 3067 2526 3072 2530
rect 3076 2526 3081 2530
rect 3085 2526 3104 2530
rect 3108 2526 3138 2530
rect 3142 2526 3153 2530
rect 3157 2526 3181 2530
rect 3185 2526 3194 2530
rect 2298 2506 2303 2509
rect 2307 2506 2331 2509
rect 2356 2506 2363 2509
rect 2367 2506 2389 2509
rect 2409 2506 2416 2509
rect 2430 2506 2435 2509
rect 2439 2506 2463 2509
rect 2488 2506 2495 2509
rect 2499 2506 2521 2509
rect 2541 2506 2548 2509
rect 2562 2506 2567 2509
rect 2571 2506 2595 2509
rect 2708 2519 2784 2523
rect 2788 2519 2793 2523
rect 2797 2519 2843 2523
rect 2847 2519 2868 2523
rect 2872 2519 2899 2523
rect 2903 2519 2932 2523
rect 2620 2506 2627 2509
rect 2631 2506 2653 2509
rect 2831 2512 2832 2516
rect 2856 2511 2857 2515
rect 2903 2512 2904 2516
rect 2314 2496 2321 2499
rect 2325 2500 2344 2503
rect 2344 2493 2347 2499
rect 2372 2496 2379 2499
rect 2383 2500 2398 2503
rect 2446 2496 2453 2499
rect 2457 2500 2476 2503
rect 2476 2493 2479 2499
rect 2504 2496 2511 2499
rect 2515 2500 2530 2503
rect 2578 2496 2585 2499
rect 2589 2500 2608 2503
rect 2608 2493 2611 2499
rect 2636 2496 2643 2499
rect 2647 2500 2664 2503
rect 2779 2498 2782 2503
rect 2786 2498 2789 2503
rect 2769 2495 2771 2498
rect 2779 2495 2789 2498
rect 2779 2489 2782 2495
rect 2281 2477 2284 2489
rect 2302 2477 2305 2489
rect 2318 2477 2321 2489
rect 2332 2480 2344 2483
rect 2360 2477 2363 2489
rect 2376 2477 2379 2489
rect 2397 2477 2400 2489
rect 2413 2477 2416 2489
rect 2434 2477 2437 2489
rect 2450 2477 2453 2489
rect 2464 2480 2476 2483
rect 2492 2477 2495 2489
rect 2508 2477 2511 2489
rect 2529 2477 2532 2489
rect 2545 2477 2548 2489
rect 2566 2477 2569 2489
rect 2582 2477 2585 2489
rect 2596 2480 2608 2483
rect 2624 2477 2627 2489
rect 2640 2477 2643 2489
rect 2661 2477 2664 2489
rect 2786 2489 2789 2495
rect 2795 2497 2798 2503
rect 2811 2498 2814 2503
rect 2795 2493 2797 2497
rect 2801 2493 2803 2497
rect 2811 2496 2817 2498
rect 2821 2496 2822 2498
rect 2811 2494 2822 2496
rect 2839 2496 2842 2503
rect 2795 2489 2798 2493
rect 2811 2489 2814 2494
rect 2840 2492 2842 2496
rect 2839 2489 2842 2492
rect 2855 2497 2858 2503
rect 2865 2497 2868 2503
rect 2886 2498 2889 2503
rect 2865 2493 2874 2497
rect 2886 2494 2887 2498
rect 2891 2495 2894 2498
rect 2911 2497 2914 2503
rect 2929 2498 2932 2503
rect 2968 2500 2971 2526
rect 3004 2519 3023 2523
rect 3027 2519 3045 2523
rect 3049 2519 3104 2523
rect 3108 2519 3129 2523
rect 3133 2519 3160 2523
rect 3164 2519 3193 2523
rect 3226 2520 3229 2530
rect 3247 2520 3250 2530
rect 3263 2520 3266 2530
rect 3277 2523 3282 2527
rect 3286 2523 3293 2527
rect 3305 2520 3308 2530
rect 3321 2520 3324 2530
rect 3342 2520 3345 2530
rect 3358 2520 3361 2530
rect 3379 2520 3382 2530
rect 3395 2520 3398 2530
rect 3409 2523 3414 2527
rect 3418 2523 3425 2527
rect 3437 2520 3440 2530
rect 3453 2520 3456 2530
rect 3474 2520 3477 2530
rect 3490 2520 3493 2530
rect 3511 2520 3514 2530
rect 3527 2520 3530 2530
rect 3541 2523 3546 2527
rect 3550 2523 3557 2527
rect 3569 2520 3572 2530
rect 3585 2520 3588 2530
rect 3606 2520 3609 2530
rect 3641 2526 3715 2530
rect 3719 2526 3721 2530
rect 3725 2526 3729 2530
rect 3733 2526 3747 2530
rect 3751 2526 3756 2530
rect 3760 2526 3765 2530
rect 3769 2526 3788 2530
rect 3792 2526 3822 2530
rect 3826 2526 3837 2530
rect 3841 2526 3865 2530
rect 3869 2526 3882 2530
rect 3886 2526 3906 2530
rect 3910 2526 3990 2530
rect 3994 2526 4008 2530
rect 4012 2526 4017 2530
rect 4021 2526 4026 2530
rect 4030 2526 4049 2530
rect 4053 2526 4083 2530
rect 4087 2526 4098 2530
rect 4102 2526 4126 2530
rect 4130 2526 4139 2530
rect 3004 2507 3007 2519
rect 3092 2512 3093 2516
rect 3117 2511 3118 2515
rect 3164 2512 3165 2516
rect 2855 2489 2858 2493
rect 2865 2489 2868 2493
rect 2886 2489 2889 2494
rect 2913 2493 2914 2497
rect 3031 2498 3034 2503
rect 3040 2498 3043 2503
rect 3047 2498 3050 2503
rect 2911 2489 2914 2493
rect 2929 2489 2932 2494
rect 2958 2487 2963 2492
rect 2967 2488 2969 2491
rect 2984 2490 2987 2496
rect 3016 2495 3050 2498
rect 2984 2487 2992 2490
rect 2984 2484 2987 2487
rect 2278 2473 2311 2477
rect 2315 2473 2339 2477
rect 2343 2473 2369 2477
rect 2373 2473 2443 2477
rect 2447 2473 2471 2477
rect 2475 2473 2501 2477
rect 2505 2473 2575 2477
rect 2579 2473 2603 2477
rect 2607 2473 2633 2477
rect 2637 2473 2690 2477
rect 2839 2474 2842 2478
rect 2866 2474 2867 2478
rect 2911 2474 2913 2478
rect 3016 2481 3019 2495
rect 3040 2489 3043 2495
rect 3047 2489 3050 2495
rect 3056 2497 3059 2503
rect 3072 2498 3075 2503
rect 3056 2493 3058 2497
rect 3062 2493 3064 2497
rect 3072 2496 3078 2498
rect 3082 2496 3083 2498
rect 3072 2494 3083 2496
rect 3100 2496 3103 2503
rect 3056 2489 3059 2493
rect 3072 2489 3075 2494
rect 3101 2492 3103 2496
rect 3100 2489 3103 2492
rect 3243 2506 3248 2509
rect 3252 2506 3276 2509
rect 3301 2506 3308 2509
rect 3312 2506 3334 2509
rect 3354 2506 3361 2509
rect 3375 2506 3380 2509
rect 3384 2506 3408 2509
rect 3433 2506 3440 2509
rect 3444 2506 3466 2509
rect 3486 2506 3493 2509
rect 3507 2506 3512 2509
rect 3516 2506 3540 2509
rect 3653 2519 3729 2523
rect 3733 2519 3738 2523
rect 3742 2519 3788 2523
rect 3792 2519 3813 2523
rect 3817 2519 3844 2523
rect 3848 2519 3877 2523
rect 3565 2506 3572 2509
rect 3576 2506 3598 2509
rect 3776 2512 3777 2516
rect 3801 2511 3802 2515
rect 3848 2512 3849 2516
rect 3116 2497 3119 2503
rect 3126 2497 3129 2503
rect 3147 2498 3150 2503
rect 3126 2493 3135 2497
rect 3147 2494 3148 2498
rect 3152 2495 3155 2498
rect 3172 2497 3175 2503
rect 3190 2498 3193 2503
rect 3116 2489 3119 2493
rect 3126 2489 3129 2493
rect 3147 2489 3150 2494
rect 3174 2493 3175 2497
rect 3172 2489 3175 2493
rect 3190 2489 3193 2494
rect 3259 2496 3266 2499
rect 3270 2500 3289 2503
rect 3289 2493 3292 2499
rect 3317 2496 3324 2499
rect 3328 2500 3343 2503
rect 3391 2496 3398 2499
rect 3402 2500 3421 2503
rect 3421 2493 3424 2499
rect 3449 2496 3456 2499
rect 3460 2500 3475 2503
rect 3523 2496 3530 2499
rect 3534 2500 3553 2503
rect 3553 2493 3556 2499
rect 3581 2496 3588 2499
rect 3592 2500 3609 2503
rect 3724 2498 3727 2503
rect 3731 2498 3734 2503
rect 3714 2495 3716 2498
rect 3724 2495 3734 2498
rect 3724 2489 3727 2495
rect 2278 2466 2287 2470
rect 2291 2466 2338 2470
rect 2342 2466 2388 2470
rect 2392 2466 2419 2470
rect 2423 2466 2470 2470
rect 2474 2466 2520 2470
rect 2524 2466 2551 2470
rect 2555 2466 2602 2470
rect 2606 2466 2652 2470
rect 2656 2467 2726 2470
rect 2782 2467 2796 2471
rect 2800 2467 2827 2471
rect 2831 2467 2849 2471
rect 2853 2467 2914 2471
rect 2918 2467 2932 2471
rect 2968 2464 2971 2476
rect 3100 2474 3103 2478
rect 3127 2474 3128 2478
rect 3172 2474 3174 2478
rect 3226 2477 3229 2489
rect 3247 2477 3250 2489
rect 3263 2477 3266 2489
rect 3277 2480 3289 2483
rect 3305 2477 3308 2489
rect 3321 2477 3324 2489
rect 3342 2477 3345 2489
rect 3358 2477 3361 2489
rect 3379 2477 3382 2489
rect 3395 2477 3398 2489
rect 3409 2480 3421 2483
rect 3437 2477 3440 2489
rect 3453 2477 3456 2489
rect 3474 2477 3477 2489
rect 3490 2477 3493 2489
rect 3511 2477 3514 2489
rect 3527 2477 3530 2489
rect 3541 2480 3553 2483
rect 3569 2477 3572 2489
rect 3585 2477 3588 2489
rect 3606 2477 3609 2489
rect 3731 2489 3734 2495
rect 3740 2497 3743 2503
rect 3756 2498 3759 2503
rect 3740 2493 3742 2497
rect 3746 2493 3748 2497
rect 3756 2496 3762 2498
rect 3766 2496 3767 2498
rect 3756 2494 3767 2496
rect 3784 2496 3787 2503
rect 3740 2489 3743 2493
rect 3756 2489 3759 2494
rect 3785 2492 3787 2496
rect 3784 2489 3787 2492
rect 3800 2497 3803 2503
rect 3810 2497 3813 2503
rect 3831 2498 3834 2503
rect 3810 2493 3819 2497
rect 3831 2494 3832 2498
rect 3836 2495 3839 2498
rect 3856 2497 3859 2503
rect 3874 2498 3877 2503
rect 3913 2500 3916 2526
rect 3949 2519 3968 2523
rect 3972 2519 3990 2523
rect 3994 2519 4049 2523
rect 4053 2519 4074 2523
rect 4078 2519 4105 2523
rect 4109 2519 4138 2523
rect 3949 2507 3952 2519
rect 4037 2512 4038 2516
rect 4062 2511 4063 2515
rect 4109 2512 4110 2516
rect 3800 2489 3803 2493
rect 3810 2489 3813 2493
rect 3831 2489 3834 2494
rect 3858 2493 3859 2497
rect 3976 2498 3979 2503
rect 3985 2498 3988 2503
rect 3992 2498 3995 2503
rect 3856 2489 3859 2493
rect 3874 2489 3877 2494
rect 3903 2487 3908 2492
rect 3912 2488 3914 2491
rect 3929 2490 3932 2496
rect 3961 2495 3995 2498
rect 3929 2487 3937 2490
rect 3929 2484 3932 2487
rect 3223 2473 3256 2477
rect 3260 2473 3284 2477
rect 3288 2473 3314 2477
rect 3318 2473 3388 2477
rect 3392 2473 3416 2477
rect 3420 2473 3446 2477
rect 3450 2473 3520 2477
rect 3524 2473 3548 2477
rect 3552 2473 3578 2477
rect 3582 2473 3635 2477
rect 3784 2474 3787 2478
rect 3811 2474 3812 2478
rect 3856 2474 3858 2478
rect 3961 2481 3964 2495
rect 3985 2489 3988 2495
rect 3992 2489 3995 2495
rect 4001 2497 4004 2503
rect 4017 2498 4020 2503
rect 4001 2493 4003 2497
rect 4007 2493 4009 2497
rect 4017 2496 4023 2498
rect 4027 2496 4028 2498
rect 4017 2494 4028 2496
rect 4045 2496 4048 2503
rect 4001 2489 4004 2493
rect 4017 2489 4020 2494
rect 4046 2492 4048 2496
rect 4045 2489 4048 2492
rect 4061 2497 4064 2503
rect 4071 2497 4074 2503
rect 4092 2498 4095 2503
rect 4071 2493 4080 2497
rect 4092 2494 4093 2498
rect 4097 2495 4100 2498
rect 4117 2497 4120 2503
rect 4135 2498 4138 2503
rect 4061 2489 4064 2493
rect 4071 2489 4074 2493
rect 4092 2489 4095 2494
rect 4119 2493 4120 2497
rect 4117 2489 4120 2493
rect 4135 2489 4138 2494
rect 3008 2467 3013 2471
rect 3017 2467 3057 2471
rect 3061 2467 3088 2471
rect 3092 2467 3110 2471
rect 3114 2467 3175 2471
rect 3179 2467 3193 2471
rect 3223 2466 3232 2470
rect 3236 2466 3283 2470
rect 3287 2466 3333 2470
rect 3337 2466 3364 2470
rect 3368 2466 3415 2470
rect 3419 2466 3465 2470
rect 3469 2466 3496 2470
rect 3500 2466 3547 2470
rect 3551 2466 3597 2470
rect 3601 2467 3671 2470
rect 3727 2467 3741 2471
rect 3745 2467 3772 2471
rect 3776 2467 3794 2471
rect 3798 2467 3859 2471
rect 3863 2467 3877 2471
rect 3913 2464 3916 2476
rect 4045 2474 4048 2478
rect 4072 2474 4073 2478
rect 4117 2474 4119 2478
rect 3953 2467 3958 2471
rect 3962 2467 4002 2471
rect 4006 2467 4033 2471
rect 4037 2467 4055 2471
rect 4059 2467 4120 2471
rect 4124 2467 4138 2471
rect 2285 2460 2669 2463
rect 2684 2460 2769 2464
rect 2773 2460 2785 2464
rect 2789 2460 2803 2464
rect 2807 2460 2814 2464
rect 2818 2460 2820 2464
rect 2824 2460 2839 2464
rect 2843 2460 2876 2464
rect 2880 2460 2881 2464
rect 2885 2460 2893 2464
rect 2897 2460 2921 2464
rect 2925 2460 2961 2464
rect 2965 2460 3004 2464
rect 3008 2460 3015 2464
rect 3019 2460 3030 2464
rect 3034 2460 3046 2464
rect 3050 2460 3064 2464
rect 3068 2460 3075 2464
rect 3079 2460 3081 2464
rect 3085 2460 3100 2464
rect 3104 2460 3137 2464
rect 3141 2460 3142 2464
rect 3146 2460 3154 2464
rect 3158 2460 3182 2464
rect 3186 2460 3194 2464
rect 3230 2460 3614 2463
rect 3629 2460 3714 2464
rect 3718 2460 3730 2464
rect 3734 2460 3748 2464
rect 3752 2460 3759 2464
rect 3763 2460 3765 2464
rect 3769 2460 3784 2464
rect 3788 2460 3821 2464
rect 3825 2460 3826 2464
rect 3830 2460 3838 2464
rect 3842 2460 3866 2464
rect 3870 2460 3906 2464
rect 3910 2460 3949 2464
rect 3953 2460 3960 2464
rect 3964 2460 3975 2464
rect 3979 2460 3991 2464
rect 3995 2460 4009 2464
rect 4013 2460 4020 2464
rect 4024 2460 4026 2464
rect 4030 2460 4045 2464
rect 4049 2460 4082 2464
rect 4086 2460 4087 2464
rect 4091 2460 4099 2464
rect 4103 2460 4127 2464
rect 4131 2460 4139 2464
rect 2428 2453 2537 2456
rect 2720 2453 2778 2457
rect 2782 2453 3012 2456
rect 3202 2454 3210 2458
rect 3373 2453 3482 2456
rect 3665 2453 3723 2457
rect 3727 2453 3957 2456
rect 4147 2454 4155 2458
rect 2408 2445 2412 2449
rect 2416 2445 2420 2449
rect 2708 2446 3022 2449
rect 2756 2439 3029 2443
rect 3198 2436 3202 2442
rect 3353 2445 3357 2449
rect 3361 2445 3365 2449
rect 3653 2446 3967 2449
rect 3701 2439 3972 2443
rect 4143 2436 4147 2442
rect 2264 2432 2396 2436
rect 2400 2432 2416 2436
rect 2432 2432 3341 2436
rect 3345 2432 3361 2436
rect 3377 2432 4235 2436
rect 2424 2425 2669 2428
rect 2744 2425 3070 2429
rect 3074 2425 3106 2429
rect 3110 2425 3173 2429
rect 3177 2425 3193 2429
rect 3369 2425 3614 2428
rect 3689 2425 4015 2429
rect 4019 2425 4051 2429
rect 4055 2425 4118 2429
rect 4122 2425 4138 2429
rect 2439 2418 2669 2421
rect 2684 2418 3056 2422
rect 3060 2418 3094 2422
rect 3098 2418 3122 2422
rect 3126 2418 3152 2422
rect 3156 2418 3189 2422
rect 2408 2409 2412 2413
rect 2416 2409 2420 2413
rect 3064 2408 3067 2418
rect 3085 2408 3088 2418
rect 3101 2408 3104 2418
rect 3115 2411 3120 2415
rect 3124 2411 3131 2415
rect 3143 2408 3146 2418
rect 3159 2408 3162 2418
rect 3180 2408 3183 2418
rect 3384 2418 3614 2421
rect 3629 2418 4001 2422
rect 4005 2418 4039 2422
rect 4043 2418 4067 2422
rect 4071 2418 4097 2422
rect 4101 2418 4134 2422
rect 3353 2409 3357 2413
rect 3361 2409 3365 2413
rect 4009 2408 4012 2418
rect 4030 2408 4033 2418
rect 4046 2408 4049 2418
rect 4060 2411 4065 2415
rect 4069 2411 4076 2415
rect 4088 2408 4091 2418
rect 4104 2408 4107 2418
rect 4125 2408 4128 2418
rect 2428 2402 2538 2405
rect 2278 2395 2287 2399
rect 2291 2395 2323 2399
rect 2327 2395 2390 2399
rect 2394 2395 2419 2399
rect 2423 2395 2455 2399
rect 2459 2395 2522 2399
rect 2526 2395 2551 2399
rect 2555 2395 2587 2399
rect 2591 2395 2654 2399
rect 2658 2395 2738 2399
rect 2278 2388 2311 2392
rect 2315 2388 2339 2392
rect 2343 2388 2369 2392
rect 2373 2388 2406 2392
rect 2410 2388 2443 2392
rect 2447 2388 2471 2392
rect 2475 2388 2501 2392
rect 2505 2388 2538 2392
rect 2542 2388 2575 2392
rect 2579 2388 2603 2392
rect 2607 2388 2633 2392
rect 2637 2388 2670 2392
rect 2674 2388 2678 2392
rect 3081 2394 3086 2397
rect 3090 2394 3114 2397
rect 3373 2402 3483 2405
rect 3139 2394 3146 2397
rect 3150 2394 3172 2397
rect 3223 2395 3232 2399
rect 3236 2395 3268 2399
rect 3272 2395 3335 2399
rect 3339 2395 3364 2399
rect 3368 2395 3400 2399
rect 3404 2395 3467 2399
rect 3471 2395 3496 2399
rect 3500 2395 3532 2399
rect 3536 2395 3599 2399
rect 3603 2395 3683 2399
rect 2281 2378 2284 2388
rect 2302 2378 2305 2388
rect 2318 2378 2321 2388
rect 2332 2381 2337 2385
rect 2341 2381 2348 2385
rect 2360 2378 2363 2388
rect 2376 2378 2379 2388
rect 2397 2378 2400 2388
rect 2413 2378 2416 2388
rect 2434 2378 2437 2388
rect 2450 2378 2453 2388
rect 2464 2381 2469 2385
rect 2473 2381 2480 2385
rect 2492 2378 2495 2388
rect 2508 2378 2511 2388
rect 2529 2378 2532 2388
rect 2545 2378 2548 2388
rect 2566 2378 2569 2388
rect 2582 2378 2585 2388
rect 2596 2381 2601 2385
rect 2605 2381 2612 2385
rect 2624 2378 2627 2388
rect 2640 2378 2643 2388
rect 2661 2378 2664 2388
rect 3097 2384 3104 2387
rect 3108 2388 3127 2391
rect 2298 2364 2303 2367
rect 2307 2364 2331 2367
rect 2356 2364 2363 2367
rect 2367 2364 2389 2367
rect 2409 2364 2416 2367
rect 2430 2364 2435 2367
rect 2439 2364 2463 2367
rect 2488 2364 2495 2367
rect 2499 2364 2521 2367
rect 2541 2364 2548 2367
rect 2562 2364 2567 2367
rect 2571 2364 2595 2367
rect 2620 2364 2627 2367
rect 2631 2364 2653 2367
rect 3127 2381 3130 2387
rect 3155 2384 3162 2387
rect 3166 2388 3181 2391
rect 3223 2388 3256 2392
rect 3260 2388 3284 2392
rect 3288 2388 3314 2392
rect 3318 2388 3351 2392
rect 3355 2388 3388 2392
rect 3392 2388 3416 2392
rect 3420 2388 3446 2392
rect 3450 2388 3483 2392
rect 3487 2388 3520 2392
rect 3524 2388 3548 2392
rect 3552 2388 3578 2392
rect 3582 2388 3615 2392
rect 3619 2388 3623 2392
rect 4026 2394 4031 2397
rect 4035 2394 4059 2397
rect 4084 2394 4091 2397
rect 4095 2394 4117 2397
rect 3226 2378 3229 2388
rect 3247 2378 3250 2388
rect 3263 2378 3266 2388
rect 3277 2381 3282 2385
rect 3286 2381 3293 2385
rect 3305 2378 3308 2388
rect 3321 2378 3324 2388
rect 3342 2378 3345 2388
rect 3358 2378 3361 2388
rect 3379 2378 3382 2388
rect 3395 2378 3398 2388
rect 3409 2381 3414 2385
rect 3418 2381 3425 2385
rect 3437 2378 3440 2388
rect 3453 2378 3456 2388
rect 3474 2378 3477 2388
rect 3490 2378 3493 2388
rect 3511 2378 3514 2388
rect 3527 2378 3530 2388
rect 3541 2381 3546 2385
rect 3550 2381 3557 2385
rect 3569 2378 3572 2388
rect 3585 2378 3588 2388
rect 3606 2378 3609 2388
rect 4042 2384 4049 2387
rect 4053 2388 4072 2391
rect 3064 2365 3067 2377
rect 3085 2365 3088 2377
rect 3101 2365 3104 2377
rect 3115 2368 3127 2371
rect 3143 2365 3146 2377
rect 3159 2365 3162 2377
rect 3180 2365 3183 2377
rect 2314 2354 2321 2357
rect 2325 2358 2344 2361
rect 2344 2351 2347 2357
rect 2372 2354 2379 2357
rect 2383 2358 2398 2361
rect 2446 2354 2453 2357
rect 2457 2358 2476 2361
rect 2476 2351 2479 2357
rect 2504 2354 2511 2357
rect 2515 2358 2530 2361
rect 2578 2354 2585 2357
rect 2589 2358 2608 2361
rect 2608 2351 2611 2357
rect 2636 2354 2643 2357
rect 2647 2358 2664 2361
rect 2696 2361 3094 2365
rect 3098 2361 3122 2365
rect 3126 2361 3152 2365
rect 3156 2361 3193 2365
rect 3243 2364 3248 2367
rect 3252 2364 3276 2367
rect 3301 2364 3308 2367
rect 3312 2364 3334 2367
rect 3354 2364 3361 2367
rect 3375 2364 3380 2367
rect 3384 2364 3408 2367
rect 3433 2364 3440 2367
rect 3444 2364 3466 2367
rect 3486 2364 3493 2367
rect 3507 2364 3512 2367
rect 3516 2364 3540 2367
rect 3565 2364 3572 2367
rect 3576 2364 3598 2367
rect 4072 2381 4075 2387
rect 4100 2384 4107 2387
rect 4111 2388 4126 2391
rect 4009 2365 4012 2377
rect 4030 2365 4033 2377
rect 4046 2365 4049 2377
rect 4060 2368 4072 2371
rect 4088 2365 4091 2377
rect 4104 2365 4107 2377
rect 4125 2365 4128 2377
rect 2732 2354 3070 2358
rect 3074 2354 3121 2358
rect 3125 2354 3171 2358
rect 3175 2354 3193 2358
rect 3259 2354 3266 2357
rect 3270 2358 3289 2361
rect 2281 2335 2284 2347
rect 2302 2335 2305 2347
rect 2318 2335 2321 2347
rect 2332 2338 2344 2341
rect 2360 2335 2363 2347
rect 2376 2335 2379 2347
rect 2397 2335 2400 2347
rect 2413 2335 2416 2347
rect 2434 2335 2437 2347
rect 2450 2335 2453 2347
rect 2464 2338 2476 2341
rect 2492 2335 2495 2347
rect 2508 2335 2511 2347
rect 2529 2335 2532 2347
rect 2545 2335 2548 2347
rect 2566 2335 2569 2347
rect 2582 2335 2585 2347
rect 2596 2338 2608 2341
rect 2624 2335 2627 2347
rect 2640 2335 2643 2347
rect 2661 2335 2664 2347
rect 3067 2347 3188 2350
rect 3289 2351 3292 2357
rect 3317 2354 3324 2357
rect 3328 2358 3343 2361
rect 3391 2354 3398 2357
rect 3402 2358 3421 2361
rect 3421 2351 3424 2357
rect 3449 2354 3456 2357
rect 3460 2358 3475 2361
rect 3523 2354 3530 2357
rect 3534 2358 3553 2361
rect 3553 2351 3556 2357
rect 3581 2354 3588 2357
rect 3592 2358 3609 2361
rect 3641 2361 4039 2365
rect 4043 2361 4067 2365
rect 4071 2361 4097 2365
rect 4101 2361 4138 2365
rect 3677 2354 4015 2358
rect 4019 2354 4066 2358
rect 4070 2354 4116 2358
rect 4120 2354 4138 2358
rect 2744 2339 3070 2343
rect 3074 2339 3106 2343
rect 3110 2339 3173 2343
rect 3177 2339 3193 2343
rect 2278 2331 2311 2335
rect 2315 2331 2339 2335
rect 2343 2331 2369 2335
rect 2373 2331 2443 2335
rect 2447 2331 2471 2335
rect 2475 2331 2501 2335
rect 2505 2331 2575 2335
rect 2579 2331 2603 2335
rect 2607 2331 2633 2335
rect 2637 2331 2690 2335
rect 3060 2332 3094 2336
rect 3098 2332 3122 2336
rect 3126 2332 3152 2336
rect 3156 2332 3189 2336
rect 3226 2335 3229 2347
rect 3247 2335 3250 2347
rect 3263 2335 3266 2347
rect 3277 2338 3289 2341
rect 3305 2335 3308 2347
rect 3321 2335 3324 2347
rect 3342 2335 3345 2347
rect 3358 2335 3361 2347
rect 3379 2335 3382 2347
rect 3395 2335 3398 2347
rect 3409 2338 3421 2341
rect 3437 2335 3440 2347
rect 3453 2335 3456 2347
rect 3474 2335 3477 2347
rect 3490 2335 3493 2347
rect 3511 2335 3514 2347
rect 3527 2335 3530 2347
rect 3541 2338 3553 2341
rect 3569 2335 3572 2347
rect 3585 2335 3588 2347
rect 3606 2335 3609 2347
rect 4012 2347 4133 2350
rect 3689 2339 4015 2343
rect 4019 2339 4051 2343
rect 4055 2339 4118 2343
rect 4122 2339 4138 2343
rect 4298 2342 4324 2355
rect 2278 2324 2287 2328
rect 2291 2324 2338 2328
rect 2342 2324 2388 2328
rect 2392 2324 2419 2328
rect 2423 2324 2470 2328
rect 2474 2324 2520 2328
rect 2524 2324 2551 2328
rect 2555 2324 2602 2328
rect 2606 2324 2652 2328
rect 2656 2324 2726 2328
rect 3064 2322 3067 2332
rect 3085 2322 3088 2332
rect 3101 2322 3104 2332
rect 3115 2325 3120 2329
rect 3124 2325 3131 2329
rect 3143 2322 3146 2332
rect 3159 2322 3162 2332
rect 3180 2322 3183 2332
rect 3223 2331 3256 2335
rect 3260 2331 3284 2335
rect 3288 2331 3314 2335
rect 3318 2331 3388 2335
rect 3392 2331 3416 2335
rect 3420 2331 3446 2335
rect 3450 2331 3520 2335
rect 3524 2331 3548 2335
rect 3552 2331 3578 2335
rect 3582 2331 3635 2335
rect 4005 2332 4039 2336
rect 4043 2332 4067 2336
rect 4071 2332 4097 2336
rect 4101 2332 4134 2336
rect 3223 2324 3232 2328
rect 3236 2324 3283 2328
rect 3287 2324 3333 2328
rect 3337 2324 3364 2328
rect 3368 2324 3415 2328
rect 3419 2324 3465 2328
rect 3469 2324 3496 2328
rect 3500 2324 3547 2328
rect 3551 2324 3597 2328
rect 3601 2324 3671 2328
rect 4009 2322 4012 2332
rect 4030 2322 4033 2332
rect 4046 2322 4049 2332
rect 4060 2325 4065 2329
rect 4069 2325 4076 2329
rect 4088 2322 4091 2332
rect 4104 2322 4107 2332
rect 4125 2322 4128 2332
rect 2284 2317 2669 2320
rect 2278 2309 2287 2313
rect 2291 2309 2323 2313
rect 2327 2309 2390 2313
rect 2394 2309 2419 2313
rect 2423 2309 2455 2313
rect 2459 2309 2522 2313
rect 2526 2309 2551 2313
rect 2555 2309 2587 2313
rect 2591 2309 2654 2313
rect 2658 2309 2738 2313
rect 2278 2302 2311 2306
rect 2315 2302 2339 2306
rect 2343 2302 2369 2306
rect 2373 2302 2406 2306
rect 2410 2302 2443 2306
rect 2447 2302 2471 2306
rect 2475 2302 2501 2306
rect 2505 2302 2538 2306
rect 2542 2302 2575 2306
rect 2579 2302 2603 2306
rect 2607 2302 2633 2306
rect 2637 2302 2670 2306
rect 2674 2302 2678 2306
rect 3081 2308 3086 2311
rect 3090 2308 3114 2311
rect 3229 2317 3614 2320
rect 3139 2308 3146 2311
rect 3150 2308 3172 2311
rect 3223 2309 3232 2313
rect 3236 2309 3268 2313
rect 3272 2309 3335 2313
rect 3339 2309 3364 2313
rect 3368 2309 3400 2313
rect 3404 2309 3467 2313
rect 3471 2309 3496 2313
rect 3500 2309 3532 2313
rect 3536 2309 3599 2313
rect 3603 2309 3683 2313
rect 2281 2292 2284 2302
rect 2302 2292 2305 2302
rect 2318 2292 2321 2302
rect 2332 2295 2337 2299
rect 2341 2295 2348 2299
rect 2360 2292 2363 2302
rect 2376 2292 2379 2302
rect 2397 2292 2400 2302
rect 2413 2292 2416 2302
rect 2434 2292 2437 2302
rect 2450 2292 2453 2302
rect 2464 2295 2469 2299
rect 2473 2295 2480 2299
rect 2492 2292 2495 2302
rect 2508 2292 2511 2302
rect 2529 2292 2532 2302
rect 2545 2292 2548 2302
rect 2566 2292 2569 2302
rect 2582 2292 2585 2302
rect 2596 2295 2601 2299
rect 2605 2295 2612 2299
rect 2624 2292 2627 2302
rect 2640 2292 2643 2302
rect 2661 2292 2664 2302
rect 3097 2298 3104 2301
rect 3108 2302 3127 2305
rect 2298 2278 2303 2281
rect 2307 2278 2331 2281
rect 2356 2278 2363 2281
rect 2367 2278 2389 2281
rect 2409 2278 2416 2281
rect 2430 2278 2435 2281
rect 2439 2278 2463 2281
rect 2488 2278 2495 2281
rect 2499 2278 2521 2281
rect 2541 2278 2548 2281
rect 2562 2278 2567 2281
rect 2571 2278 2595 2281
rect 2620 2278 2627 2281
rect 2631 2278 2653 2281
rect 3127 2295 3130 2301
rect 3155 2298 3162 2301
rect 3166 2302 3181 2305
rect 3192 2300 3203 2304
rect 3223 2302 3256 2306
rect 3260 2302 3284 2306
rect 3288 2302 3314 2306
rect 3318 2302 3351 2306
rect 3355 2302 3388 2306
rect 3392 2302 3416 2306
rect 3420 2302 3446 2306
rect 3450 2302 3483 2306
rect 3487 2302 3520 2306
rect 3524 2302 3548 2306
rect 3552 2302 3578 2306
rect 3582 2302 3615 2306
rect 3619 2302 3623 2306
rect 4026 2308 4031 2311
rect 4035 2308 4059 2311
rect 4084 2308 4091 2311
rect 4095 2308 4117 2311
rect 3226 2292 3229 2302
rect 3247 2292 3250 2302
rect 3263 2292 3266 2302
rect 3277 2295 3282 2299
rect 3286 2295 3293 2299
rect 3305 2292 3308 2302
rect 3321 2292 3324 2302
rect 3342 2292 3345 2302
rect 3358 2292 3361 2302
rect 3379 2292 3382 2302
rect 3395 2292 3398 2302
rect 3409 2295 3414 2299
rect 3418 2295 3425 2299
rect 3437 2292 3440 2302
rect 3453 2292 3456 2302
rect 3474 2292 3477 2302
rect 3490 2292 3493 2302
rect 3511 2292 3514 2302
rect 3527 2292 3530 2302
rect 3541 2295 3546 2299
rect 3550 2295 3557 2299
rect 3569 2292 3572 2302
rect 3585 2292 3588 2302
rect 3606 2292 3609 2302
rect 4042 2298 4049 2301
rect 4053 2302 4072 2305
rect 3064 2279 3067 2291
rect 3085 2279 3088 2291
rect 3101 2279 3104 2291
rect 3115 2282 3127 2285
rect 3143 2279 3146 2291
rect 3159 2279 3162 2291
rect 3180 2279 3183 2291
rect 2314 2268 2321 2271
rect 2325 2272 2344 2275
rect 2344 2265 2347 2271
rect 2372 2268 2379 2271
rect 2383 2272 2398 2275
rect 2446 2268 2453 2271
rect 2457 2272 2476 2275
rect 2476 2265 2479 2271
rect 2504 2268 2511 2271
rect 2515 2272 2530 2275
rect 2578 2268 2585 2271
rect 2589 2272 2608 2275
rect 2608 2265 2611 2271
rect 2636 2268 2643 2271
rect 2647 2272 2664 2275
rect 2696 2275 3094 2279
rect 3098 2275 3122 2279
rect 3126 2275 3152 2279
rect 3156 2275 3193 2279
rect 3243 2278 3248 2281
rect 3252 2278 3276 2281
rect 3301 2278 3308 2281
rect 3312 2278 3334 2281
rect 3354 2278 3361 2281
rect 3375 2278 3380 2281
rect 3384 2278 3408 2281
rect 3433 2278 3440 2281
rect 3444 2278 3466 2281
rect 3486 2278 3493 2281
rect 3507 2278 3512 2281
rect 3516 2278 3540 2281
rect 3565 2278 3572 2281
rect 3576 2278 3598 2281
rect 4072 2295 4075 2301
rect 4100 2298 4107 2301
rect 4111 2302 4126 2305
rect 4137 2300 4148 2304
rect 4009 2279 4012 2291
rect 4030 2279 4033 2291
rect 4046 2279 4049 2291
rect 4060 2282 4072 2285
rect 4088 2279 4091 2291
rect 4104 2279 4107 2291
rect 4125 2279 4128 2291
rect 2732 2268 3070 2272
rect 3074 2268 3121 2272
rect 3125 2268 3171 2272
rect 3175 2268 3193 2272
rect 3259 2268 3266 2271
rect 3270 2272 3289 2275
rect 3289 2265 3292 2271
rect 3317 2268 3324 2271
rect 3328 2272 3343 2275
rect 3391 2268 3398 2271
rect 3402 2272 3421 2275
rect 3421 2265 3424 2271
rect 3449 2268 3456 2271
rect 3460 2272 3475 2275
rect 3523 2268 3530 2271
rect 3534 2272 3553 2275
rect 3553 2265 3556 2271
rect 3581 2268 3588 2271
rect 3592 2272 3609 2275
rect 3641 2275 4039 2279
rect 4043 2275 4067 2279
rect 4071 2275 4097 2279
rect 4101 2275 4138 2279
rect 3677 2268 4015 2272
rect 4019 2268 4066 2272
rect 4070 2268 4116 2272
rect 4120 2268 4138 2272
rect 2281 2249 2284 2261
rect 2302 2249 2305 2261
rect 2318 2249 2321 2261
rect 2332 2252 2344 2255
rect 2360 2249 2363 2261
rect 2376 2249 2379 2261
rect 2397 2249 2400 2261
rect 2413 2249 2416 2261
rect 2434 2249 2437 2261
rect 2450 2249 2453 2261
rect 2464 2252 2476 2255
rect 2492 2249 2495 2261
rect 2508 2249 2511 2261
rect 2529 2249 2532 2261
rect 2545 2249 2548 2261
rect 2566 2249 2569 2261
rect 2582 2249 2585 2261
rect 2596 2252 2608 2255
rect 2624 2249 2627 2261
rect 2640 2249 2643 2261
rect 2661 2249 2664 2261
rect 3226 2249 3229 2261
rect 3247 2249 3250 2261
rect 3263 2249 3266 2261
rect 3277 2252 3289 2255
rect 3305 2249 3308 2261
rect 3321 2249 3324 2261
rect 3342 2249 3345 2261
rect 3358 2249 3361 2261
rect 3379 2249 3382 2261
rect 3395 2249 3398 2261
rect 3409 2252 3421 2255
rect 3437 2249 3440 2261
rect 3453 2249 3456 2261
rect 3474 2249 3477 2261
rect 3490 2249 3493 2261
rect 3511 2249 3514 2261
rect 3527 2249 3530 2261
rect 3541 2252 3553 2255
rect 3569 2249 3572 2261
rect 3585 2249 3588 2261
rect 3606 2249 3609 2261
rect 2278 2245 2311 2249
rect 2315 2245 2339 2249
rect 2343 2245 2369 2249
rect 2373 2245 2443 2249
rect 2447 2245 2471 2249
rect 2475 2245 2501 2249
rect 2505 2245 2575 2249
rect 2579 2245 2603 2249
rect 2607 2245 2633 2249
rect 2637 2245 2690 2249
rect 3223 2245 3256 2249
rect 3260 2245 3284 2249
rect 3288 2245 3314 2249
rect 3318 2245 3388 2249
rect 3392 2245 3416 2249
rect 3420 2245 3446 2249
rect 3450 2245 3520 2249
rect 3524 2245 3548 2249
rect 3552 2245 3578 2249
rect 3582 2245 3635 2249
rect 2278 2238 2287 2242
rect 2291 2238 2338 2242
rect 2342 2238 2388 2242
rect 2392 2238 2419 2242
rect 2423 2238 2470 2242
rect 2474 2238 2520 2242
rect 2524 2238 2551 2242
rect 2555 2238 2602 2242
rect 2606 2238 2652 2242
rect 2656 2238 2726 2242
rect 3223 2238 3232 2242
rect 3236 2238 3283 2242
rect 3287 2238 3333 2242
rect 3337 2238 3364 2242
rect 3368 2238 3415 2242
rect 3419 2238 3465 2242
rect 3469 2238 3496 2242
rect 3500 2238 3547 2242
rect 3551 2238 3597 2242
rect 3601 2238 3671 2242
rect 2284 2232 2669 2235
rect 3229 2232 3614 2235
rect 2409 2225 2513 2228
rect 3354 2225 3458 2228
rect 2525 2217 2529 2221
rect 2533 2217 2537 2221
rect 3470 2217 3474 2221
rect 3478 2217 3482 2221
rect 2261 2206 2513 2210
rect 2517 2206 2533 2210
rect 2549 2206 3210 2210
rect 3214 2206 3458 2210
rect 3462 2206 3478 2210
rect 3494 2206 4155 2210
rect 4159 2206 4242 2210
rect 2541 2199 2669 2202
rect 3486 2199 3614 2202
rect 2556 2192 2669 2195
rect 3501 2192 3614 2195
rect 2525 2183 2529 2187
rect 2533 2183 2537 2187
rect 3470 2183 3474 2187
rect 3478 2183 3482 2187
rect 2409 2176 2513 2179
rect 3354 2176 3458 2179
rect 2278 2169 2287 2173
rect 2291 2169 2323 2173
rect 2327 2169 2390 2173
rect 2394 2169 2419 2173
rect 2423 2169 2455 2173
rect 2459 2169 2522 2173
rect 2526 2169 2551 2173
rect 2555 2169 2587 2173
rect 2591 2169 2654 2173
rect 2658 2169 2738 2173
rect 3223 2169 3232 2173
rect 3236 2169 3268 2173
rect 3272 2169 3335 2173
rect 3339 2169 3364 2173
rect 3368 2169 3400 2173
rect 3404 2169 3467 2173
rect 3471 2169 3496 2173
rect 3500 2169 3532 2173
rect 3536 2169 3599 2173
rect 3603 2169 3683 2173
rect 2278 2162 2311 2166
rect 2315 2162 2339 2166
rect 2343 2162 2369 2166
rect 2373 2162 2406 2166
rect 2410 2162 2443 2166
rect 2447 2162 2471 2166
rect 2475 2162 2501 2166
rect 2505 2162 2538 2166
rect 2542 2162 2575 2166
rect 2579 2162 2603 2166
rect 2607 2162 2633 2166
rect 2637 2162 2670 2166
rect 2674 2162 2678 2166
rect 3223 2162 3256 2166
rect 3260 2162 3284 2166
rect 3288 2162 3314 2166
rect 3318 2162 3351 2166
rect 3355 2162 3388 2166
rect 3392 2162 3416 2166
rect 3420 2162 3446 2166
rect 3450 2162 3483 2166
rect 3487 2162 3520 2166
rect 3524 2162 3548 2166
rect 3552 2162 3578 2166
rect 3582 2162 3615 2166
rect 3619 2162 3623 2166
rect 2281 2152 2284 2162
rect 2302 2152 2305 2162
rect 2318 2152 2321 2162
rect 2332 2155 2337 2159
rect 2341 2155 2348 2159
rect 2360 2152 2363 2162
rect 2376 2152 2379 2162
rect 2397 2152 2400 2162
rect 2413 2152 2416 2162
rect 2434 2152 2437 2162
rect 2450 2152 2453 2162
rect 2464 2155 2469 2159
rect 2473 2155 2480 2159
rect 2492 2152 2495 2162
rect 2508 2152 2511 2162
rect 2529 2152 2532 2162
rect 2545 2152 2548 2162
rect 2566 2152 2569 2162
rect 2582 2152 2585 2162
rect 2596 2155 2601 2159
rect 2605 2155 2612 2159
rect 2624 2152 2627 2162
rect 2640 2152 2643 2162
rect 2661 2152 2664 2162
rect 3226 2152 3229 2162
rect 3247 2152 3250 2162
rect 3263 2152 3266 2162
rect 3277 2155 3282 2159
rect 3286 2155 3293 2159
rect 3305 2152 3308 2162
rect 3321 2152 3324 2162
rect 3342 2152 3345 2162
rect 3358 2152 3361 2162
rect 3379 2152 3382 2162
rect 3395 2152 3398 2162
rect 3409 2155 3414 2159
rect 3418 2155 3425 2159
rect 3437 2152 3440 2162
rect 3453 2152 3456 2162
rect 3474 2152 3477 2162
rect 3490 2152 3493 2162
rect 3511 2152 3514 2162
rect 3527 2152 3530 2162
rect 3541 2155 3546 2159
rect 3550 2155 3557 2159
rect 3569 2152 3572 2162
rect 3585 2152 3588 2162
rect 3606 2152 3609 2162
rect 2298 2138 2303 2141
rect 2307 2138 2331 2141
rect 2356 2138 2363 2141
rect 2367 2138 2389 2141
rect 2409 2138 2416 2141
rect 2430 2138 2435 2141
rect 2439 2138 2463 2141
rect 2488 2138 2495 2141
rect 2499 2138 2521 2141
rect 2541 2138 2548 2141
rect 2562 2138 2567 2141
rect 2571 2138 2595 2141
rect 2620 2138 2627 2141
rect 2631 2138 2653 2141
rect 2314 2128 2321 2131
rect 2325 2132 2344 2135
rect 2344 2125 2347 2131
rect 2372 2128 2379 2131
rect 2383 2132 2398 2135
rect 2446 2128 2453 2131
rect 2457 2132 2476 2135
rect 2476 2125 2479 2131
rect 2504 2128 2511 2131
rect 2515 2132 2530 2135
rect 2578 2128 2585 2131
rect 2589 2132 2608 2135
rect 2608 2125 2611 2131
rect 2636 2128 2643 2131
rect 2647 2132 2664 2135
rect 3243 2138 3248 2141
rect 3252 2138 3276 2141
rect 3301 2138 3308 2141
rect 3312 2138 3334 2141
rect 3354 2138 3361 2141
rect 3375 2138 3380 2141
rect 3384 2138 3408 2141
rect 3433 2138 3440 2141
rect 3444 2138 3466 2141
rect 3486 2138 3493 2141
rect 3507 2138 3512 2141
rect 3516 2138 3540 2141
rect 3565 2138 3572 2141
rect 3576 2138 3598 2141
rect 3259 2128 3266 2131
rect 3270 2132 3289 2135
rect 3289 2125 3292 2131
rect 3317 2128 3324 2131
rect 3328 2132 3343 2135
rect 3391 2128 3398 2131
rect 3402 2132 3421 2135
rect 3421 2125 3424 2131
rect 3449 2128 3456 2131
rect 3460 2132 3475 2135
rect 3523 2128 3530 2131
rect 3534 2132 3553 2135
rect 3553 2125 3556 2131
rect 3581 2128 3588 2131
rect 3592 2132 3609 2135
rect 2281 2109 2284 2121
rect 2302 2109 2305 2121
rect 2318 2109 2321 2121
rect 2332 2112 2344 2115
rect 2360 2109 2363 2121
rect 2376 2109 2379 2121
rect 2397 2109 2400 2121
rect 2413 2109 2416 2121
rect 2434 2109 2437 2121
rect 2450 2109 2453 2121
rect 2464 2112 2476 2115
rect 2492 2109 2495 2121
rect 2508 2109 2511 2121
rect 2529 2109 2532 2121
rect 2545 2109 2548 2121
rect 2566 2109 2569 2121
rect 2582 2109 2585 2121
rect 2596 2112 2608 2115
rect 2624 2109 2627 2121
rect 2640 2109 2643 2121
rect 2661 2109 2664 2121
rect 3226 2109 3229 2121
rect 3247 2109 3250 2121
rect 3263 2109 3266 2121
rect 3277 2112 3289 2115
rect 3305 2109 3308 2121
rect 3321 2109 3324 2121
rect 3342 2109 3345 2121
rect 3358 2109 3361 2121
rect 3379 2109 3382 2121
rect 3395 2109 3398 2121
rect 3409 2112 3421 2115
rect 3437 2109 3440 2121
rect 3453 2109 3456 2121
rect 3474 2109 3477 2121
rect 3490 2109 3493 2121
rect 3511 2109 3514 2121
rect 3527 2109 3530 2121
rect 3541 2112 3553 2115
rect 3569 2109 3572 2121
rect 3585 2109 3588 2121
rect 3606 2109 3609 2121
rect 2278 2105 2311 2109
rect 2315 2105 2339 2109
rect 2343 2105 2369 2109
rect 2373 2105 2443 2109
rect 2447 2105 2471 2109
rect 2475 2105 2501 2109
rect 2505 2105 2575 2109
rect 2579 2105 2603 2109
rect 2607 2105 2633 2109
rect 2637 2105 2690 2109
rect 3223 2105 3256 2109
rect 3260 2105 3284 2109
rect 3288 2105 3314 2109
rect 3318 2105 3388 2109
rect 3392 2105 3416 2109
rect 3420 2105 3446 2109
rect 3450 2105 3520 2109
rect 3524 2105 3548 2109
rect 3552 2105 3578 2109
rect 3582 2105 3635 2109
rect 2278 2098 2287 2102
rect 2291 2098 2338 2102
rect 2342 2098 2388 2102
rect 2392 2098 2419 2102
rect 2423 2098 2470 2102
rect 2474 2098 2520 2102
rect 2524 2098 2551 2102
rect 2555 2098 2602 2102
rect 2606 2098 2652 2102
rect 2656 2098 2726 2102
rect 3223 2098 3232 2102
rect 3236 2098 3283 2102
rect 3287 2098 3333 2102
rect 3337 2098 3364 2102
rect 3368 2098 3415 2102
rect 3419 2098 3465 2102
rect 3469 2098 3496 2102
rect 3500 2098 3547 2102
rect 3551 2098 3597 2102
rect 3601 2098 3671 2102
<< m2contact >>
rect 2027 4300 2040 4304
rect 2935 4312 2940 4316
rect 2954 4314 2967 4318
rect 3241 4313 3293 4317
rect 3548 4311 3604 4316
rect 2336 4282 2349 4304
rect 2411 4282 2416 4304
rect 2027 4254 2048 4279
rect 2315 4256 2328 4278
rect 2390 4256 2395 4278
rect 2738 4204 2744 4208
rect 3683 4204 3689 4208
rect 2726 4196 2732 4200
rect 3671 4196 3677 4200
rect 2714 4189 2720 4193
rect 3659 4189 3665 4193
rect 2702 4182 2708 4186
rect 3647 4182 3653 4186
rect 2690 4173 2696 4178
rect 3241 4174 3296 4178
rect 3635 4174 3641 4178
rect 2678 4166 2684 4170
rect 3549 4166 3604 4170
rect 3623 4167 3629 4171
rect 2750 4159 2756 4163
rect 3695 4159 3701 4163
rect 2954 4151 2967 4155
rect 3337 4151 3341 4155
rect 2935 4141 2940 4145
rect 3325 4141 3330 4145
rect 3671 4119 3677 4123
rect 3659 4111 3665 4115
rect 3647 4103 3653 4107
rect 3635 4095 3641 4099
rect 3623 4087 3629 4091
rect 2738 4054 2744 4058
rect 2771 4054 2775 4058
rect 2807 4054 2811 4058
rect 2874 4054 2878 4058
rect 2903 4054 2907 4058
rect 2939 4054 2943 4058
rect 3006 4054 3010 4058
rect 3035 4054 3039 4058
rect 3071 4054 3075 4058
rect 3138 4054 3142 4058
rect 3167 4054 3171 4058
rect 3203 4054 3207 4058
rect 3270 4054 3274 4058
rect 3683 4054 3689 4058
rect 3716 4054 3720 4058
rect 3752 4054 3756 4058
rect 3819 4054 3823 4058
rect 3848 4054 3852 4058
rect 3884 4054 3888 4058
rect 3951 4054 3955 4058
rect 3980 4054 3984 4058
rect 4016 4054 4020 4058
rect 4083 4054 4087 4058
rect 4112 4054 4116 4058
rect 4148 4054 4152 4058
rect 4215 4054 4219 4058
rect 2678 4047 2684 4051
rect 3623 4047 3629 4051
rect 2771 4040 2775 4044
rect 2821 4040 2825 4044
rect 2874 4040 2878 4044
rect 2903 4040 2907 4044
rect 2953 4040 2957 4044
rect 3006 4040 3010 4044
rect 3035 4040 3039 4044
rect 3085 4040 3089 4044
rect 3138 4040 3142 4044
rect 3167 4040 3171 4044
rect 3217 4040 3221 4044
rect 3270 4040 3274 4044
rect 3716 4040 3720 4044
rect 3766 4040 3770 4044
rect 3819 4040 3823 4044
rect 3848 4040 3852 4044
rect 3898 4040 3902 4044
rect 3951 4040 3955 4044
rect 3980 4040 3984 4044
rect 4030 4040 4034 4044
rect 4083 4040 4087 4044
rect 4112 4040 4116 4044
rect 4162 4040 4166 4044
rect 4215 4040 4219 4044
rect 2794 4029 2798 4033
rect 2419 4021 2423 4025
rect 2455 4021 2459 4025
rect 2522 4021 2526 4025
rect 2738 4021 2744 4025
rect 2765 4020 2769 4024
rect 2778 4023 2782 4029
rect 2815 4023 2819 4029
rect 2828 4025 2832 4029
rect 2852 4029 2856 4033
rect 2926 4029 2930 4033
rect 2836 4023 2840 4029
rect 2873 4023 2877 4029
rect 2889 4025 2893 4029
rect 2678 4014 2684 4018
rect 2419 4007 2423 4011
rect 2469 4007 2473 4011
rect 2522 4007 2526 4011
rect 2778 4010 2782 4014
rect 2794 4010 2798 4016
rect 2828 4016 2832 4020
rect 2815 4010 2819 4014
rect 2836 4010 2840 4014
rect 2852 4010 2856 4016
rect 2897 4020 2901 4024
rect 2910 4023 2914 4029
rect 2947 4023 2951 4029
rect 2960 4025 2964 4029
rect 2984 4029 2988 4033
rect 3058 4029 3062 4033
rect 2968 4023 2972 4029
rect 3005 4023 3009 4029
rect 3021 4025 3025 4029
rect 2873 4010 2877 4014
rect 2889 4010 2893 4014
rect 2910 4010 2914 4014
rect 2926 4010 2930 4016
rect 2960 4016 2964 4020
rect 2947 4010 2951 4014
rect 2968 4010 2972 4014
rect 2984 4010 2988 4016
rect 3029 4020 3033 4024
rect 3042 4023 3046 4029
rect 3079 4023 3083 4029
rect 3092 4025 3096 4029
rect 3116 4029 3120 4033
rect 3190 4029 3194 4033
rect 3100 4023 3104 4029
rect 3137 4023 3141 4029
rect 3153 4025 3157 4029
rect 3005 4010 3009 4014
rect 3021 4010 3025 4014
rect 3042 4010 3046 4014
rect 3058 4010 3062 4016
rect 3092 4016 3096 4020
rect 3079 4010 3083 4014
rect 3100 4010 3104 4014
rect 3116 4010 3120 4016
rect 3161 4020 3165 4024
rect 3174 4023 3178 4029
rect 3211 4023 3215 4029
rect 3224 4025 3228 4029
rect 3248 4029 3252 4033
rect 3739 4029 3743 4033
rect 3232 4023 3236 4029
rect 3269 4023 3273 4029
rect 3285 4025 3289 4029
rect 3364 4021 3368 4025
rect 3400 4021 3404 4025
rect 3467 4021 3471 4025
rect 3683 4021 3689 4025
rect 3137 4010 3141 4014
rect 3153 4010 3157 4014
rect 3174 4010 3178 4014
rect 3190 4010 3194 4016
rect 3224 4016 3228 4020
rect 3211 4010 3215 4014
rect 2442 3996 2446 4000
rect 2404 3987 2408 3991
rect 2426 3990 2430 3996
rect 2463 3990 2467 3996
rect 2476 3992 2480 3996
rect 2500 3996 2504 4000
rect 2484 3990 2488 3996
rect 2521 3990 2525 3996
rect 2537 3990 2541 3996
rect 2771 3999 2775 4003
rect 2808 3997 2812 4001
rect 2828 3997 2832 4001
rect 2872 3997 2876 4001
rect 2903 3999 2907 4003
rect 2940 3997 2944 4001
rect 2960 3997 2964 4001
rect 3004 3997 3008 4001
rect 3035 3999 3039 4003
rect 3072 3997 3076 4001
rect 3092 3997 3096 4001
rect 3136 3997 3140 4001
rect 3153 4002 3157 4006
rect 3232 4010 3236 4014
rect 3248 4010 3252 4016
rect 3710 4020 3714 4024
rect 3723 4023 3727 4029
rect 3760 4023 3764 4029
rect 3773 4025 3777 4029
rect 3797 4029 3801 4033
rect 3871 4029 3875 4033
rect 3781 4023 3785 4029
rect 3818 4023 3822 4029
rect 3834 4025 3838 4029
rect 3623 4014 3629 4018
rect 3269 4010 3273 4014
rect 3285 4010 3289 4014
rect 3167 3999 3171 4003
rect 3204 3997 3208 4001
rect 3224 3997 3228 4001
rect 3268 3997 3272 4001
rect 3285 4002 3289 4006
rect 3364 4007 3368 4011
rect 3414 4007 3418 4011
rect 3467 4007 3471 4011
rect 3723 4010 3727 4014
rect 3739 4010 3743 4016
rect 3773 4016 3777 4020
rect 3760 4010 3764 4014
rect 3781 4010 3785 4014
rect 3797 4010 3801 4016
rect 3842 4020 3846 4024
rect 3855 4023 3859 4029
rect 3892 4023 3896 4029
rect 3905 4025 3909 4029
rect 3929 4029 3933 4033
rect 4003 4029 4007 4033
rect 3913 4023 3917 4029
rect 3950 4023 3954 4029
rect 3966 4025 3970 4029
rect 3818 4010 3822 4014
rect 3834 4010 3838 4014
rect 3855 4010 3859 4014
rect 3871 4010 3875 4016
rect 3905 4016 3909 4020
rect 3892 4010 3896 4014
rect 3913 4010 3917 4014
rect 3929 4010 3933 4016
rect 3974 4020 3978 4024
rect 3987 4023 3991 4029
rect 4024 4023 4028 4029
rect 4037 4025 4041 4029
rect 4061 4029 4065 4033
rect 4135 4029 4139 4033
rect 4045 4023 4049 4029
rect 4082 4023 4086 4029
rect 4098 4025 4102 4029
rect 3950 4010 3954 4014
rect 3966 4010 3970 4014
rect 3987 4010 3991 4014
rect 4003 4010 4007 4016
rect 4037 4016 4041 4020
rect 4024 4010 4028 4014
rect 4045 4010 4049 4014
rect 4061 4010 4065 4016
rect 4106 4020 4110 4024
rect 4119 4023 4123 4029
rect 4156 4023 4160 4029
rect 4169 4025 4173 4029
rect 4193 4029 4197 4033
rect 4177 4023 4181 4029
rect 4214 4023 4218 4029
rect 4230 4025 4234 4029
rect 4082 4010 4086 4014
rect 4098 4010 4102 4014
rect 4119 4010 4123 4014
rect 4135 4010 4139 4016
rect 4169 4016 4173 4020
rect 4156 4010 4160 4014
rect 3387 3996 3391 4000
rect 2690 3990 2696 3994
rect 2426 3977 2430 3981
rect 2442 3977 2446 3983
rect 2476 3983 2480 3987
rect 2463 3977 2467 3981
rect 2484 3977 2488 3981
rect 2500 3977 2504 3983
rect 3349 3987 3353 3991
rect 3371 3990 3375 3996
rect 3408 3990 3412 3996
rect 3421 3992 3425 3996
rect 3445 3996 3449 4000
rect 3429 3990 3433 3996
rect 3466 3990 3470 3996
rect 3482 3990 3486 3996
rect 3716 3999 3720 4003
rect 3753 3997 3757 4001
rect 3773 3997 3777 4001
rect 3817 3997 3821 4001
rect 3848 3999 3852 4003
rect 3885 3997 3889 4001
rect 3905 3997 3909 4001
rect 3949 3997 3953 4001
rect 3980 3999 3984 4003
rect 4017 3997 4021 4001
rect 4037 3997 4041 4001
rect 4081 3997 4085 4001
rect 4098 4002 4102 4006
rect 4177 4010 4181 4014
rect 4193 4010 4197 4016
rect 4214 4010 4218 4014
rect 4230 4010 4234 4014
rect 4112 3999 4116 4003
rect 4149 3997 4153 4001
rect 4169 3997 4173 4001
rect 4213 3997 4217 4001
rect 4230 4002 4234 4006
rect 3635 3990 3641 3994
rect 2726 3983 2732 3987
rect 2771 3983 2775 3987
rect 2822 3983 2826 3987
rect 2872 3983 2876 3987
rect 2903 3983 2907 3987
rect 2954 3983 2958 3987
rect 3004 3983 3008 3987
rect 3035 3983 3039 3987
rect 3086 3983 3090 3987
rect 3136 3983 3140 3987
rect 3167 3983 3171 3987
rect 3218 3983 3222 3987
rect 3268 3983 3272 3987
rect 2521 3977 2525 3981
rect 2537 3977 2541 3981
rect 3371 3977 3375 3981
rect 3387 3977 3391 3983
rect 3421 3983 3425 3987
rect 3408 3977 3412 3981
rect 2419 3966 2423 3970
rect 2456 3964 2460 3968
rect 2476 3964 2480 3968
rect 2520 3964 2524 3968
rect 2678 3970 2684 3974
rect 2769 3970 2773 3974
rect 2803 3970 2807 3974
rect 2820 3970 2824 3974
rect 2876 3970 2880 3974
rect 2893 3970 2897 3974
rect 2921 3970 2925 3974
rect 3429 3977 3433 3981
rect 3445 3977 3449 3983
rect 3671 3983 3677 3987
rect 3716 3983 3720 3987
rect 3767 3983 3771 3987
rect 3817 3983 3821 3987
rect 3848 3983 3852 3987
rect 3899 3983 3903 3987
rect 3949 3983 3953 3987
rect 3980 3983 3984 3987
rect 4031 3983 4035 3987
rect 4081 3983 4085 3987
rect 4112 3983 4116 3987
rect 4163 3983 4167 3987
rect 4213 3983 4217 3987
rect 3466 3977 3470 3981
rect 3482 3977 3486 3981
rect 2714 3963 2720 3967
rect 2796 3963 2800 3967
rect 2827 3963 2831 3967
rect 2849 3963 2853 3967
rect 2914 3963 2918 3967
rect 2690 3957 2696 3961
rect 2419 3950 2423 3954
rect 2470 3950 2474 3954
rect 2520 3950 2524 3954
rect 2726 3950 2732 3954
rect 2770 3953 2774 3957
rect 2795 3956 2799 3960
rect 2802 3953 2806 3957
rect 2820 3953 2824 3957
rect 2842 3956 2846 3960
rect 2867 3956 2871 3960
rect 2877 3953 2881 3957
rect 2893 3953 2897 3957
rect 2913 3956 2917 3960
rect 2920 3953 2924 3957
rect 2984 3963 2988 3967
rect 2537 3943 2541 3947
rect 2404 3934 2408 3938
rect 2529 3936 2533 3940
rect 2553 3936 2557 3940
rect 2412 3927 2416 3931
rect 2553 3927 2557 3931
rect 2797 3937 2801 3941
rect 2817 3934 2821 3938
rect 2836 3938 2840 3942
rect 2938 3949 2942 3953
rect 2953 3949 2957 3953
rect 2855 3937 2859 3941
rect 2874 3937 2878 3941
rect 2887 3936 2891 3940
rect 2909 3937 2913 3941
rect 2917 3936 2921 3940
rect 2929 3936 2933 3940
rect 2770 3923 2774 3927
rect 2802 3923 2806 3927
rect 2820 3923 2824 3927
rect 2877 3923 2881 3927
rect 2892 3923 2896 3927
rect 2920 3923 2924 3927
rect 2419 3919 2423 3923
rect 2486 3919 2490 3923
rect 2522 3919 2526 3923
rect 2738 3919 2744 3923
rect 2784 3919 2788 3923
rect 2827 3918 2831 3922
rect 2849 3919 2856 3923
rect 2899 3918 2903 3922
rect 2678 3912 2684 3916
rect 2419 3905 2423 3909
rect 2472 3905 2476 3909
rect 2522 3905 2526 3909
rect 2702 3911 2708 3915
rect 2784 3911 2788 3915
rect 2843 3911 2847 3915
rect 2868 3911 2872 3915
rect 2899 3911 2903 3915
rect 2992 3941 2996 3949
rect 3065 3963 3069 3967
rect 3019 3949 3023 3953
rect 3034 3949 3038 3953
rect 3015 3941 3019 3945
rect 2961 3935 2965 3939
rect 2974 3927 2978 3931
rect 3073 3941 3077 3949
rect 3229 3957 3242 3965
rect 3325 3957 3330 3965
rect 3364 3966 3368 3970
rect 3401 3964 3405 3968
rect 3421 3964 3425 3968
rect 3465 3964 3469 3968
rect 3623 3970 3629 3974
rect 3714 3970 3718 3974
rect 3748 3970 3752 3974
rect 3765 3970 3769 3974
rect 3821 3970 3825 3974
rect 3838 3970 3842 3974
rect 3866 3970 3870 3974
rect 3659 3963 3665 3967
rect 3741 3963 3745 3967
rect 3772 3963 3776 3967
rect 3794 3963 3798 3967
rect 3859 3963 3863 3967
rect 3635 3957 3641 3961
rect 3275 3948 3279 3952
rect 3337 3948 3341 3952
rect 3364 3950 3368 3954
rect 3415 3950 3419 3954
rect 3465 3950 3469 3954
rect 3671 3950 3677 3954
rect 3715 3953 3719 3957
rect 3740 3956 3744 3960
rect 3747 3953 3751 3957
rect 3765 3953 3769 3957
rect 3787 3956 3791 3960
rect 3812 3956 3816 3960
rect 3822 3953 3826 3957
rect 3838 3953 3842 3957
rect 3858 3956 3862 3960
rect 3865 3953 3869 3957
rect 3929 3963 3933 3967
rect 3100 3941 3104 3945
rect 3482 3943 3486 3947
rect 3042 3935 3046 3939
rect 3349 3934 3353 3938
rect 3474 3936 3478 3940
rect 3498 3936 3502 3940
rect 3707 3936 3711 3940
rect 3055 3927 3059 3931
rect 3357 3927 3361 3931
rect 3498 3927 3502 3931
rect 3742 3937 3746 3941
rect 3762 3934 3766 3938
rect 3781 3938 3785 3942
rect 3883 3949 3887 3953
rect 3898 3949 3902 3953
rect 3800 3937 3804 3941
rect 3819 3937 3823 3941
rect 3832 3936 3836 3940
rect 3854 3937 3858 3941
rect 3862 3936 3866 3940
rect 3874 3936 3878 3940
rect 3715 3923 3719 3927
rect 3747 3923 3751 3927
rect 3765 3923 3769 3927
rect 3822 3923 3826 3927
rect 3837 3923 3841 3927
rect 3865 3923 3869 3927
rect 3364 3919 3368 3923
rect 3431 3919 3435 3923
rect 3467 3919 3471 3923
rect 3683 3919 3689 3923
rect 3729 3919 3733 3923
rect 3772 3918 3776 3922
rect 3794 3919 3801 3923
rect 3844 3918 3848 3922
rect 3623 3912 3629 3916
rect 2690 3904 2696 3908
rect 2770 3904 2774 3908
rect 2784 3904 2788 3908
rect 2802 3904 2806 3908
rect 2820 3904 2824 3908
rect 2843 3904 2847 3908
rect 2877 3904 2881 3908
rect 2892 3904 2896 3908
rect 2920 3904 2924 3908
rect 2441 3894 2445 3898
rect 2404 3888 2408 3894
rect 2420 3888 2424 3894
rect 2457 3888 2461 3894
rect 2465 3890 2469 3894
rect 2499 3894 2503 3898
rect 2702 3897 2708 3901
rect 2784 3897 2788 3901
rect 2843 3897 2847 3901
rect 2868 3897 2872 3901
rect 2899 3897 2903 3901
rect 2478 3888 2482 3894
rect 2515 3888 2519 3894
rect 2784 3889 2788 3893
rect 2827 3890 2831 3894
rect 2849 3889 2856 3893
rect 2899 3890 2903 3894
rect 2537 3885 2541 3889
rect 2770 3885 2774 3889
rect 2802 3885 2806 3889
rect 2820 3885 2824 3889
rect 2877 3885 2881 3889
rect 2892 3885 2896 3889
rect 2920 3885 2924 3889
rect 2404 3875 2408 3879
rect 2420 3875 2424 3879
rect 2465 3881 2469 3885
rect 2441 3875 2445 3881
rect 2457 3875 2461 3879
rect 2478 3875 2482 3879
rect 2499 3875 2503 3881
rect 2515 3875 2519 3879
rect 2765 3873 2769 3877
rect 2421 3862 2425 3866
rect 2465 3862 2469 3866
rect 2485 3862 2489 3866
rect 2522 3864 2526 3868
rect 2797 3871 2801 3875
rect 2817 3874 2821 3878
rect 2836 3870 2840 3874
rect 2855 3871 2859 3875
rect 2874 3871 2878 3875
rect 2887 3872 2891 3876
rect 2984 3887 2988 3891
rect 3364 3905 3368 3909
rect 3417 3905 3421 3909
rect 3467 3905 3471 3909
rect 3647 3911 3653 3915
rect 3729 3911 3733 3915
rect 3788 3911 3792 3915
rect 3813 3911 3817 3915
rect 3844 3911 3848 3915
rect 3937 3941 3941 3949
rect 4010 3963 4014 3967
rect 3964 3949 3968 3953
rect 3979 3949 3983 3953
rect 3960 3941 3964 3945
rect 3906 3935 3910 3939
rect 3919 3927 3923 3931
rect 4018 3941 4022 3949
rect 4045 3941 4049 3945
rect 3987 3935 3991 3939
rect 4000 3927 4004 3931
rect 3635 3904 3641 3908
rect 3715 3904 3719 3908
rect 3729 3904 3733 3908
rect 3747 3904 3751 3908
rect 3765 3904 3769 3908
rect 3788 3904 3792 3908
rect 3822 3904 3826 3908
rect 3837 3904 3841 3908
rect 3865 3904 3869 3908
rect 3386 3894 3390 3898
rect 3065 3887 3069 3891
rect 3349 3888 3353 3894
rect 3365 3888 3369 3894
rect 3402 3888 3406 3894
rect 3410 3890 3414 3894
rect 3444 3894 3448 3898
rect 3647 3897 3653 3901
rect 3729 3897 3733 3901
rect 3788 3897 3792 3901
rect 3813 3897 3817 3901
rect 3844 3897 3848 3901
rect 3423 3888 3427 3894
rect 3460 3888 3464 3894
rect 3729 3889 3733 3893
rect 3772 3890 3776 3894
rect 3794 3889 3801 3893
rect 3844 3890 3848 3894
rect 3482 3885 3486 3889
rect 3715 3885 3719 3889
rect 3747 3885 3751 3889
rect 3765 3885 3769 3889
rect 3822 3885 3826 3889
rect 3837 3885 3841 3889
rect 3865 3885 3869 3889
rect 2909 3871 2913 3875
rect 2917 3872 2921 3876
rect 2929 3872 2933 3876
rect 2964 3872 2968 3876
rect 2992 3871 2996 3875
rect 3044 3872 3048 3876
rect 3349 3875 3353 3879
rect 3365 3875 3369 3879
rect 3410 3881 3414 3885
rect 3386 3875 3390 3881
rect 3402 3875 3406 3879
rect 3073 3871 3077 3875
rect 3423 3875 3427 3879
rect 3444 3875 3448 3881
rect 3460 3875 3464 3879
rect 3710 3873 3714 3877
rect 2690 3855 2696 3859
rect 2770 3855 2774 3859
rect 2795 3852 2799 3856
rect 2802 3855 2806 3859
rect 2820 3855 2824 3859
rect 2842 3852 2846 3856
rect 2867 3852 2871 3856
rect 2877 3855 2881 3859
rect 2893 3855 2897 3859
rect 2913 3852 2917 3856
rect 2920 3855 2924 3859
rect 2421 3848 2425 3852
rect 2471 3848 2475 3852
rect 2522 3848 2526 3852
rect 2726 3848 2732 3852
rect 2780 3845 2784 3849
rect 2796 3845 2800 3849
rect 2827 3845 2831 3849
rect 2849 3845 2853 3849
rect 2914 3845 2918 3849
rect 2974 3851 2978 3855
rect 3366 3862 3370 3866
rect 3410 3862 3414 3866
rect 3430 3862 3434 3866
rect 3467 3864 3471 3868
rect 3742 3871 3746 3875
rect 3762 3874 3766 3878
rect 3781 3870 3785 3874
rect 3800 3871 3804 3875
rect 3819 3871 3823 3875
rect 3832 3872 3836 3876
rect 3929 3887 3933 3891
rect 4010 3887 4014 3891
rect 3854 3871 3858 3875
rect 3862 3872 3866 3876
rect 3874 3872 3878 3876
rect 3909 3872 3913 3876
rect 3937 3871 3941 3875
rect 3989 3872 3993 3876
rect 4018 3871 4022 3875
rect 3635 3855 3641 3859
rect 3715 3855 3719 3859
rect 3055 3851 3059 3855
rect 3740 3852 3744 3856
rect 3747 3855 3751 3859
rect 3765 3855 3769 3859
rect 3787 3852 3791 3856
rect 3812 3852 3816 3856
rect 3822 3855 3826 3859
rect 3838 3855 3842 3859
rect 3858 3852 3862 3856
rect 3865 3855 3869 3859
rect 3366 3848 3370 3852
rect 3416 3848 3420 3852
rect 3467 3848 3471 3852
rect 3671 3848 3677 3852
rect 3725 3845 3729 3849
rect 3741 3845 3745 3849
rect 3772 3845 3776 3849
rect 3794 3845 3798 3849
rect 3859 3845 3863 3849
rect 3919 3851 3923 3855
rect 4000 3851 4004 3855
rect 2678 3838 2684 3842
rect 2769 3838 2773 3842
rect 2803 3838 2807 3842
rect 2820 3838 2824 3842
rect 2876 3838 2880 3842
rect 2893 3838 2897 3842
rect 2921 3838 2925 3842
rect 3623 3838 3629 3842
rect 3714 3838 3718 3842
rect 3748 3838 3752 3842
rect 3765 3838 3769 3842
rect 3821 3838 3825 3842
rect 3838 3838 3842 3842
rect 3866 3838 3870 3842
rect 2714 3831 2720 3835
rect 2780 3831 2784 3835
rect 2796 3831 2800 3835
rect 2827 3831 2831 3835
rect 2849 3831 2853 3835
rect 2914 3831 2918 3835
rect 2984 3831 2988 3835
rect 2770 3821 2774 3825
rect 2795 3824 2799 3828
rect 2802 3821 2806 3825
rect 2820 3821 2824 3825
rect 2842 3824 2846 3828
rect 2867 3824 2871 3828
rect 2877 3821 2881 3825
rect 2893 3821 2897 3825
rect 2913 3824 2917 3828
rect 2920 3821 2924 3825
rect 2764 3804 2768 3808
rect 2797 3805 2801 3809
rect 2817 3802 2821 3806
rect 2836 3806 2840 3810
rect 2855 3805 2859 3809
rect 2874 3805 2878 3809
rect 2887 3804 2891 3808
rect 2909 3805 2913 3809
rect 2917 3804 2921 3808
rect 2929 3804 2933 3808
rect 2992 3809 2996 3817
rect 3089 3831 3093 3835
rect 3043 3817 3047 3821
rect 3058 3817 3062 3821
rect 3275 3827 3279 3831
rect 3659 3831 3665 3835
rect 3725 3831 3729 3835
rect 3741 3831 3745 3835
rect 3772 3831 3776 3835
rect 3794 3831 3798 3835
rect 3859 3831 3863 3835
rect 3929 3831 3933 3835
rect 2961 3803 2965 3807
rect 3015 3808 3019 3812
rect 2770 3791 2774 3795
rect 2802 3791 2806 3795
rect 2820 3791 2824 3795
rect 2877 3791 2881 3795
rect 2892 3791 2896 3795
rect 2920 3791 2924 3795
rect 2784 3787 2788 3791
rect 2827 3786 2831 3790
rect 2849 3787 2856 3791
rect 2899 3786 2903 3790
rect 2702 3779 2708 3783
rect 2784 3779 2788 3783
rect 2843 3779 2847 3783
rect 2868 3779 2872 3783
rect 2899 3779 2903 3783
rect 2974 3795 2978 3799
rect 3097 3809 3101 3817
rect 3715 3821 3719 3825
rect 3740 3824 3744 3828
rect 3747 3821 3751 3825
rect 3765 3821 3769 3825
rect 3787 3824 3791 3828
rect 3812 3824 3816 3828
rect 3822 3821 3826 3825
rect 3838 3821 3842 3825
rect 3858 3824 3862 3828
rect 3865 3821 3869 3825
rect 3118 3809 3122 3813
rect 3582 3809 3586 3813
rect 3066 3803 3070 3807
rect 3079 3795 3083 3799
rect 3320 3802 3324 3806
rect 3274 3788 3278 3792
rect 3289 3788 3293 3792
rect 3297 3780 3301 3784
rect 3328 3780 3332 3788
rect 3709 3804 3713 3808
rect 2690 3772 2696 3776
rect 2770 3772 2774 3776
rect 2784 3772 2788 3776
rect 2802 3772 2806 3776
rect 2820 3772 2824 3776
rect 2843 3772 2847 3776
rect 2877 3772 2881 3776
rect 2892 3772 2896 3776
rect 2920 3772 2924 3776
rect 2702 3765 2708 3769
rect 2784 3765 2788 3769
rect 2843 3765 2847 3769
rect 2868 3765 2872 3769
rect 2899 3765 2903 3769
rect 2784 3757 2788 3761
rect 2827 3758 2831 3762
rect 2849 3757 2856 3761
rect 2899 3758 2903 3762
rect 2770 3753 2774 3757
rect 2802 3753 2806 3757
rect 2820 3753 2824 3757
rect 2877 3753 2881 3757
rect 2892 3753 2896 3757
rect 2920 3753 2924 3757
rect 2984 3756 2988 3760
rect 3089 3756 3093 3760
rect 2765 3741 2769 3745
rect 2797 3739 2801 3743
rect 2817 3742 2821 3746
rect 2836 3738 2840 3742
rect 2855 3739 2859 3743
rect 2874 3739 2878 3743
rect 2887 3740 2891 3744
rect 2909 3739 2913 3743
rect 2917 3740 2921 3744
rect 2929 3740 2933 3744
rect 2963 3741 2967 3745
rect 2992 3740 2996 3744
rect 3069 3741 3073 3745
rect 3097 3740 3101 3744
rect 3310 3766 3314 3770
rect 3742 3805 3746 3809
rect 3762 3802 3766 3806
rect 3781 3806 3785 3810
rect 3800 3805 3804 3809
rect 3819 3805 3823 3809
rect 3832 3804 3836 3808
rect 3854 3805 3858 3809
rect 3862 3804 3866 3808
rect 3874 3804 3878 3808
rect 3937 3809 3941 3817
rect 4034 3831 4038 3835
rect 3988 3817 3992 3821
rect 4003 3817 4007 3821
rect 3906 3803 3910 3807
rect 3960 3808 3964 3812
rect 3715 3791 3719 3795
rect 3747 3791 3751 3795
rect 3765 3791 3769 3795
rect 3822 3791 3826 3795
rect 3837 3791 3841 3795
rect 3865 3791 3869 3795
rect 3729 3787 3733 3791
rect 3772 3786 3776 3790
rect 3794 3787 3801 3791
rect 3844 3786 3848 3790
rect 3647 3779 3653 3783
rect 3729 3779 3733 3783
rect 3788 3779 3792 3783
rect 3813 3779 3817 3783
rect 3844 3779 3848 3783
rect 3919 3795 3923 3799
rect 4042 3809 4046 3817
rect 4063 3809 4067 3813
rect 4011 3803 4015 3807
rect 4024 3795 4028 3799
rect 3635 3772 3641 3776
rect 3715 3772 3719 3776
rect 3729 3772 3733 3776
rect 3747 3772 3751 3776
rect 3765 3772 3769 3776
rect 3788 3772 3792 3776
rect 3822 3772 3826 3776
rect 3837 3772 3841 3776
rect 3865 3772 3869 3776
rect 3507 3760 3511 3764
rect 3647 3765 3653 3769
rect 3729 3765 3733 3769
rect 3788 3765 3792 3769
rect 3813 3765 3817 3769
rect 3844 3765 3848 3769
rect 3729 3757 3733 3761
rect 3772 3758 3776 3762
rect 3794 3757 3801 3761
rect 3844 3758 3848 3762
rect 3540 3752 3544 3756
rect 3659 3752 3665 3756
rect 3715 3753 3719 3757
rect 3747 3753 3751 3757
rect 3765 3753 3769 3757
rect 3822 3753 3826 3757
rect 3837 3753 3841 3757
rect 3865 3753 3869 3757
rect 3929 3756 3933 3760
rect 4034 3756 4038 3760
rect 3582 3740 3586 3744
rect 3623 3740 3629 3744
rect 3710 3741 3714 3745
rect 3635 3733 3641 3737
rect 3574 3729 3579 3733
rect 2770 3723 2774 3727
rect 2795 3720 2799 3724
rect 2802 3723 2806 3727
rect 2820 3723 2824 3727
rect 2842 3720 2846 3724
rect 2867 3720 2871 3724
rect 2877 3723 2881 3727
rect 2893 3723 2897 3727
rect 2913 3720 2917 3724
rect 2920 3723 2924 3727
rect 2714 3713 2720 3717
rect 2796 3713 2800 3717
rect 2827 3713 2831 3717
rect 2849 3713 2853 3717
rect 2914 3713 2918 3717
rect 2974 3720 2978 3724
rect 3079 3720 3083 3724
rect 3320 3722 3324 3726
rect 3590 3724 3594 3728
rect 3695 3724 3701 3728
rect 3742 3739 3746 3743
rect 3762 3742 3766 3746
rect 3781 3738 3785 3742
rect 3800 3739 3804 3743
rect 3819 3739 3823 3743
rect 3832 3740 3836 3744
rect 3854 3739 3858 3743
rect 3862 3740 3866 3744
rect 3874 3740 3878 3744
rect 3908 3741 3912 3745
rect 3937 3740 3941 3744
rect 4014 3741 4018 3745
rect 4042 3740 4046 3744
rect 3715 3723 3719 3727
rect 3740 3720 3744 3724
rect 3747 3723 3751 3727
rect 3765 3723 3769 3727
rect 3787 3720 3791 3724
rect 3812 3720 3816 3724
rect 3822 3723 3826 3727
rect 3838 3723 3842 3727
rect 3858 3720 3862 3724
rect 3865 3723 3869 3727
rect 3507 3715 3512 3719
rect 3647 3715 3653 3719
rect 2678 3706 2684 3710
rect 2769 3706 2773 3710
rect 2803 3706 2807 3710
rect 2820 3706 2824 3710
rect 2876 3706 2880 3710
rect 2893 3706 2897 3710
rect 2921 3706 2925 3710
rect 3240 3707 3244 3711
rect 3659 3713 3665 3717
rect 3741 3713 3745 3717
rect 3772 3713 3776 3717
rect 3794 3713 3798 3717
rect 3859 3713 3863 3717
rect 3919 3720 3923 3724
rect 4024 3720 4028 3724
rect 3328 3706 3332 3710
rect 3623 3706 3629 3710
rect 3714 3706 3718 3710
rect 3748 3706 3752 3710
rect 3765 3706 3769 3710
rect 3821 3706 3825 3710
rect 3838 3706 3842 3710
rect 3866 3706 3870 3710
rect 2714 3699 2720 3703
rect 2796 3699 2800 3703
rect 2827 3699 2831 3703
rect 2849 3699 2853 3703
rect 2914 3699 2918 3703
rect 2984 3699 2988 3703
rect 2770 3689 2774 3693
rect 2795 3692 2799 3696
rect 2802 3689 2806 3693
rect 2820 3689 2824 3693
rect 2842 3692 2846 3696
rect 2867 3692 2871 3696
rect 2877 3689 2881 3693
rect 2893 3689 2897 3693
rect 2913 3692 2917 3696
rect 2920 3689 2924 3693
rect 2764 3672 2768 3676
rect 2797 3673 2801 3677
rect 2817 3670 2821 3674
rect 2836 3674 2840 3678
rect 2855 3673 2859 3677
rect 2874 3673 2878 3677
rect 2887 3672 2891 3676
rect 2909 3673 2913 3677
rect 2917 3672 2921 3676
rect 2929 3672 2933 3676
rect 2992 3677 2996 3685
rect 3065 3699 3069 3703
rect 3019 3685 3023 3689
rect 3034 3685 3038 3689
rect 3015 3677 3019 3681
rect 2961 3671 2965 3675
rect 2770 3659 2774 3663
rect 2802 3659 2806 3663
rect 2820 3659 2824 3663
rect 2877 3659 2881 3663
rect 2892 3659 2896 3663
rect 2920 3659 2924 3663
rect 2784 3655 2788 3659
rect 2827 3654 2831 3658
rect 2849 3655 2856 3659
rect 2899 3654 2903 3658
rect 2702 3647 2708 3651
rect 2784 3647 2788 3651
rect 2843 3647 2847 3651
rect 2868 3647 2872 3651
rect 2899 3647 2903 3651
rect 2974 3663 2978 3667
rect 3073 3677 3077 3685
rect 3155 3699 3159 3703
rect 3109 3685 3113 3689
rect 3124 3685 3128 3689
rect 3097 3677 3101 3681
rect 3042 3671 3046 3675
rect 3131 3679 3135 3683
rect 3163 3677 3167 3685
rect 3659 3699 3665 3703
rect 3741 3699 3745 3703
rect 3772 3699 3776 3703
rect 3794 3699 3798 3703
rect 3859 3699 3863 3703
rect 3929 3699 3933 3703
rect 3310 3686 3314 3690
rect 3715 3689 3719 3693
rect 3740 3692 3744 3696
rect 3747 3689 3751 3693
rect 3765 3689 3769 3693
rect 3787 3692 3791 3696
rect 3812 3692 3816 3696
rect 3822 3689 3826 3693
rect 3838 3689 3842 3693
rect 3858 3692 3862 3696
rect 3865 3689 3869 3693
rect 3055 3663 3059 3667
rect 3198 3676 3202 3680
rect 3582 3679 3586 3683
rect 3145 3663 3149 3667
rect 3320 3672 3324 3676
rect 3252 3658 3256 3662
rect 3267 3658 3271 3662
rect 3274 3658 3278 3662
rect 3289 3658 3293 3662
rect 3297 3650 3301 3654
rect 3328 3650 3332 3658
rect 3709 3672 3713 3676
rect 2690 3640 2696 3644
rect 2770 3640 2774 3644
rect 2784 3640 2788 3644
rect 2802 3640 2806 3644
rect 2820 3640 2824 3644
rect 2843 3640 2847 3644
rect 2877 3640 2881 3644
rect 2892 3640 2896 3644
rect 2920 3640 2924 3644
rect 2702 3633 2708 3637
rect 2784 3633 2788 3637
rect 2843 3633 2847 3637
rect 2868 3633 2872 3637
rect 2899 3633 2903 3637
rect 2784 3625 2788 3629
rect 2827 3626 2831 3630
rect 2849 3625 2856 3629
rect 2899 3626 2903 3630
rect 2770 3621 2774 3625
rect 2802 3621 2806 3625
rect 2820 3621 2824 3625
rect 2877 3621 2881 3625
rect 2892 3621 2896 3625
rect 2920 3621 2924 3625
rect 2765 3609 2769 3613
rect 2797 3607 2801 3611
rect 2817 3610 2821 3614
rect 2836 3606 2840 3610
rect 2855 3607 2859 3611
rect 2874 3607 2878 3611
rect 2887 3608 2891 3612
rect 2984 3621 2988 3625
rect 3065 3621 3069 3625
rect 3155 3621 3159 3625
rect 2909 3607 2913 3611
rect 2917 3608 2921 3612
rect 2929 3608 2933 3612
rect 2964 3606 2968 3610
rect 2992 3605 2996 3609
rect 3044 3606 3048 3610
rect 3073 3605 3077 3609
rect 3128 3606 3132 3610
rect 3163 3605 3167 3609
rect 3310 3636 3314 3640
rect 3742 3673 3746 3677
rect 3762 3670 3766 3674
rect 3781 3674 3785 3678
rect 3800 3673 3804 3677
rect 3819 3673 3823 3677
rect 3832 3672 3836 3676
rect 3854 3673 3858 3677
rect 3862 3672 3866 3676
rect 3874 3672 3878 3676
rect 3937 3677 3941 3685
rect 4010 3699 4014 3703
rect 3964 3685 3968 3689
rect 3979 3685 3983 3689
rect 3960 3677 3964 3681
rect 3906 3671 3910 3675
rect 3715 3659 3719 3663
rect 3747 3659 3751 3663
rect 3765 3659 3769 3663
rect 3822 3659 3826 3663
rect 3837 3659 3841 3663
rect 3865 3659 3869 3663
rect 3729 3655 3733 3659
rect 3772 3654 3776 3658
rect 3794 3655 3801 3659
rect 3844 3654 3848 3658
rect 3647 3647 3653 3651
rect 3729 3647 3733 3651
rect 3788 3647 3792 3651
rect 3813 3647 3817 3651
rect 3844 3647 3848 3651
rect 3919 3663 3923 3667
rect 4018 3677 4022 3685
rect 4100 3699 4104 3703
rect 4054 3685 4058 3689
rect 4069 3685 4073 3689
rect 4042 3677 4046 3681
rect 3987 3671 3991 3675
rect 4076 3679 4080 3683
rect 4108 3677 4112 3685
rect 4000 3663 4004 3667
rect 4143 3676 4147 3680
rect 4090 3663 4094 3667
rect 3402 3630 3406 3634
rect 3635 3640 3641 3644
rect 3715 3640 3719 3644
rect 3729 3640 3733 3644
rect 3747 3640 3751 3644
rect 3765 3640 3769 3644
rect 3788 3640 3792 3644
rect 3822 3640 3826 3644
rect 3837 3640 3841 3644
rect 3865 3640 3869 3644
rect 3647 3633 3653 3637
rect 3729 3633 3733 3637
rect 3788 3633 3792 3637
rect 3813 3633 3817 3637
rect 3844 3633 3848 3637
rect 3446 3622 3450 3626
rect 3729 3625 3733 3629
rect 3772 3626 3776 3630
rect 3794 3625 3801 3629
rect 3844 3626 3848 3630
rect 3683 3619 3689 3623
rect 3715 3621 3719 3625
rect 3747 3621 3751 3625
rect 3765 3621 3769 3625
rect 3822 3621 3826 3625
rect 3837 3621 3841 3625
rect 3865 3621 3869 3625
rect 3710 3609 3714 3613
rect 2770 3591 2774 3595
rect 2795 3588 2799 3592
rect 2802 3591 2806 3595
rect 2820 3591 2824 3595
rect 2842 3588 2846 3592
rect 2867 3588 2871 3592
rect 2877 3591 2881 3595
rect 2893 3591 2897 3595
rect 2913 3588 2917 3592
rect 2920 3591 2924 3595
rect 3574 3599 3579 3603
rect 2714 3581 2720 3585
rect 2796 3581 2800 3585
rect 2827 3581 2831 3585
rect 2849 3581 2853 3585
rect 2914 3581 2918 3585
rect 2974 3585 2978 3589
rect 3055 3585 3059 3589
rect 3320 3592 3324 3596
rect 3742 3607 3746 3611
rect 3762 3610 3766 3614
rect 3781 3606 3785 3610
rect 3800 3607 3804 3611
rect 3819 3607 3823 3611
rect 3832 3608 3836 3612
rect 3929 3621 3933 3625
rect 4010 3621 4014 3625
rect 4100 3621 4104 3625
rect 3854 3607 3858 3611
rect 3862 3608 3866 3612
rect 3874 3608 3878 3612
rect 3909 3606 3913 3610
rect 3937 3605 3941 3609
rect 3989 3606 3993 3610
rect 4018 3605 4022 3609
rect 4073 3606 4077 3610
rect 4108 3605 4112 3609
rect 3402 3589 3406 3593
rect 3671 3589 3677 3593
rect 3715 3591 3719 3595
rect 3145 3585 3149 3589
rect 3740 3588 3744 3592
rect 3747 3591 3751 3595
rect 3765 3591 3769 3595
rect 3787 3588 3791 3592
rect 3812 3588 3816 3592
rect 3822 3591 3826 3595
rect 3838 3591 3842 3595
rect 3858 3588 3862 3592
rect 3865 3591 3869 3595
rect 2678 3574 2684 3578
rect 2769 3574 2773 3578
rect 2803 3574 2807 3578
rect 2820 3574 2824 3578
rect 2876 3574 2880 3578
rect 2893 3574 2897 3578
rect 2921 3574 2925 3578
rect 3242 3577 3246 3581
rect 3659 3581 3665 3585
rect 3741 3581 3745 3585
rect 3772 3581 3776 3585
rect 3794 3581 3798 3585
rect 3859 3581 3863 3585
rect 3328 3576 3332 3580
rect 3919 3585 3923 3589
rect 4000 3585 4004 3589
rect 4090 3585 4094 3589
rect 2714 3567 2720 3571
rect 2796 3567 2800 3571
rect 2827 3567 2831 3571
rect 2849 3567 2853 3571
rect 2914 3567 2918 3571
rect 2984 3567 2988 3571
rect 3623 3574 3629 3578
rect 3714 3574 3718 3578
rect 3748 3574 3752 3578
rect 3765 3574 3769 3578
rect 3821 3574 3825 3578
rect 3838 3574 3842 3578
rect 3866 3574 3870 3578
rect 2770 3557 2774 3561
rect 2795 3560 2799 3564
rect 2802 3557 2806 3561
rect 2820 3557 2824 3561
rect 2842 3560 2846 3564
rect 2867 3560 2871 3564
rect 2877 3557 2881 3561
rect 2893 3557 2897 3561
rect 2913 3560 2917 3564
rect 2920 3557 2924 3561
rect 2764 3540 2768 3544
rect 2797 3541 2801 3545
rect 2817 3538 2821 3542
rect 2836 3542 2840 3546
rect 2855 3541 2859 3545
rect 2874 3541 2878 3545
rect 2887 3540 2891 3544
rect 2909 3541 2913 3545
rect 2917 3540 2921 3544
rect 2929 3540 2933 3544
rect 2992 3545 2996 3553
rect 3659 3567 3665 3571
rect 3741 3567 3745 3571
rect 3772 3567 3776 3571
rect 3794 3567 3798 3571
rect 3859 3567 3863 3571
rect 3929 3567 3933 3571
rect 3310 3556 3314 3560
rect 3715 3557 3719 3561
rect 3740 3560 3744 3564
rect 3747 3557 3751 3561
rect 3765 3557 3769 3561
rect 3787 3560 3791 3564
rect 3812 3560 3816 3564
rect 3822 3557 3826 3561
rect 3838 3557 3842 3561
rect 3858 3560 3862 3564
rect 3865 3557 3869 3561
rect 3582 3549 3586 3553
rect 2961 3539 2965 3543
rect 3015 3544 3019 3548
rect 3709 3540 3713 3544
rect 2265 3526 2269 3530
rect 2390 3526 2394 3530
rect 2770 3527 2774 3531
rect 2802 3527 2806 3531
rect 2820 3527 2824 3531
rect 2877 3527 2881 3531
rect 2892 3527 2896 3531
rect 2920 3527 2924 3531
rect 2784 3523 2788 3527
rect 2287 3519 2291 3523
rect 2323 3519 2327 3523
rect 2390 3519 2394 3523
rect 2419 3519 2423 3523
rect 2455 3519 2459 3523
rect 2522 3519 2526 3523
rect 2551 3519 2555 3523
rect 2587 3519 2591 3523
rect 2654 3519 2658 3523
rect 2738 3519 2744 3523
rect 2827 3522 2831 3526
rect 2849 3523 2856 3527
rect 2899 3522 2903 3526
rect 2678 3512 2684 3516
rect 2784 3515 2788 3519
rect 2793 3515 2797 3519
rect 2843 3515 2847 3519
rect 2868 3515 2872 3519
rect 2899 3515 2903 3519
rect 2974 3531 2978 3535
rect 3742 3541 3746 3545
rect 3762 3538 3766 3542
rect 3781 3542 3785 3546
rect 3800 3541 3804 3545
rect 3819 3541 3823 3545
rect 3832 3540 3836 3544
rect 3854 3541 3858 3545
rect 3862 3540 3866 3544
rect 3874 3540 3878 3544
rect 3937 3545 3941 3553
rect 3906 3539 3910 3543
rect 3960 3544 3964 3548
rect 3715 3527 3719 3531
rect 3747 3527 3751 3531
rect 3765 3527 3769 3531
rect 3822 3527 3826 3531
rect 3837 3527 3841 3531
rect 3865 3527 3869 3531
rect 3729 3523 3733 3527
rect 3232 3519 3236 3523
rect 3268 3519 3272 3523
rect 3335 3519 3339 3523
rect 3364 3519 3368 3523
rect 3400 3519 3404 3523
rect 3467 3519 3471 3523
rect 3496 3519 3500 3523
rect 3532 3519 3536 3523
rect 3599 3519 3603 3523
rect 3683 3519 3689 3523
rect 3772 3522 3776 3526
rect 3794 3523 3801 3527
rect 3844 3522 3848 3526
rect 3623 3512 3629 3516
rect 3729 3515 3733 3519
rect 3738 3515 3742 3519
rect 3788 3515 3792 3519
rect 3813 3515 3817 3519
rect 3844 3515 3848 3519
rect 3919 3531 3923 3535
rect 2287 3505 2291 3509
rect 2337 3505 2341 3509
rect 2390 3505 2394 3509
rect 2419 3505 2423 3509
rect 2469 3505 2473 3509
rect 2522 3505 2526 3509
rect 2551 3505 2555 3509
rect 2601 3505 2605 3509
rect 2654 3505 2658 3509
rect 2690 3508 2696 3512
rect 2770 3508 2774 3512
rect 2784 3508 2788 3512
rect 2802 3508 2806 3512
rect 2820 3508 2824 3512
rect 2843 3508 2847 3512
rect 2877 3508 2881 3512
rect 2892 3508 2896 3512
rect 2920 3508 2924 3512
rect 3045 3508 3049 3512
rect 3063 3508 3067 3512
rect 3081 3508 3085 3512
rect 3104 3508 3108 3512
rect 3138 3508 3142 3512
rect 3153 3508 3157 3512
rect 3181 3508 3185 3512
rect 2310 3494 2314 3498
rect 2281 3485 2285 3489
rect 2294 3488 2298 3494
rect 2331 3488 2335 3494
rect 2344 3490 2348 3494
rect 2368 3494 2372 3498
rect 2442 3494 2446 3498
rect 2352 3488 2356 3494
rect 2389 3488 2393 3494
rect 2405 3488 2409 3494
rect 2426 3488 2430 3494
rect 2463 3488 2467 3494
rect 2476 3490 2480 3494
rect 2500 3494 2504 3498
rect 2574 3494 2578 3498
rect 2484 3488 2488 3494
rect 2521 3488 2525 3494
rect 2537 3488 2541 3494
rect 2558 3488 2562 3494
rect 2595 3488 2599 3494
rect 2608 3490 2612 3494
rect 2632 3494 2636 3498
rect 2702 3501 2708 3505
rect 2784 3501 2788 3505
rect 2793 3501 2797 3505
rect 2843 3501 2847 3505
rect 2868 3501 2872 3505
rect 2899 3501 2903 3505
rect 2616 3488 2620 3494
rect 2653 3488 2657 3494
rect 2669 3490 2673 3494
rect 2784 3493 2788 3497
rect 2827 3494 2831 3498
rect 2849 3493 2856 3497
rect 2899 3494 2903 3498
rect 2770 3489 2774 3493
rect 2802 3489 2806 3493
rect 2820 3489 2824 3493
rect 2877 3489 2881 3493
rect 2892 3489 2896 3493
rect 2920 3489 2924 3493
rect 2294 3475 2298 3479
rect 2310 3475 2314 3481
rect 2344 3481 2348 3485
rect 2331 3475 2335 3479
rect 2352 3475 2356 3479
rect 2368 3475 2372 3481
rect 2389 3475 2393 3479
rect 2405 3475 2409 3479
rect 2426 3475 2430 3479
rect 2442 3475 2446 3481
rect 2476 3481 2480 3485
rect 2463 3475 2467 3479
rect 2484 3475 2488 3479
rect 2500 3475 2504 3481
rect 2521 3475 2525 3479
rect 2537 3475 2541 3479
rect 2558 3475 2562 3479
rect 2574 3475 2578 3481
rect 2608 3481 2612 3485
rect 2595 3475 2599 3479
rect 2616 3475 2620 3479
rect 2632 3475 2636 3481
rect 2653 3475 2657 3479
rect 2669 3475 2673 3479
rect 2765 3477 2769 3481
rect 2287 3464 2291 3468
rect 2324 3462 2328 3466
rect 2344 3462 2348 3466
rect 2388 3462 2392 3466
rect 2419 3464 2423 3468
rect 2456 3462 2460 3466
rect 2476 3462 2480 3466
rect 2520 3462 2524 3466
rect 2551 3464 2555 3468
rect 2588 3462 2592 3466
rect 2608 3462 2612 3466
rect 2652 3462 2656 3466
rect 2797 3475 2801 3479
rect 2817 3478 2821 3482
rect 2836 3474 2840 3478
rect 2855 3475 2859 3479
rect 2874 3475 2878 3479
rect 2887 3476 2891 3480
rect 3023 3501 3027 3505
rect 3045 3501 3049 3505
rect 3104 3501 3108 3505
rect 3129 3501 3133 3505
rect 3160 3501 3164 3505
rect 3232 3505 3236 3509
rect 3282 3505 3286 3509
rect 3335 3505 3339 3509
rect 3364 3505 3368 3509
rect 3414 3505 3418 3509
rect 3467 3505 3471 3509
rect 3496 3505 3500 3509
rect 3546 3505 3550 3509
rect 3599 3505 3603 3509
rect 3635 3508 3641 3512
rect 3715 3508 3719 3512
rect 3729 3508 3733 3512
rect 3747 3508 3751 3512
rect 3765 3508 3769 3512
rect 3788 3508 3792 3512
rect 3822 3508 3826 3512
rect 3837 3508 3841 3512
rect 3865 3508 3869 3512
rect 3990 3508 3994 3512
rect 4008 3508 4012 3512
rect 4026 3508 4030 3512
rect 4049 3508 4053 3512
rect 4083 3508 4087 3512
rect 4098 3508 4102 3512
rect 4126 3508 4130 3512
rect 3045 3493 3049 3497
rect 3088 3494 3092 3498
rect 3110 3493 3117 3497
rect 3160 3494 3164 3498
rect 3255 3494 3259 3498
rect 3063 3489 3067 3493
rect 3081 3489 3085 3493
rect 3138 3489 3142 3493
rect 3153 3489 3157 3493
rect 3181 3489 3185 3493
rect 2984 3485 2988 3489
rect 2909 3475 2913 3479
rect 2917 3476 2921 3480
rect 2929 3476 2933 3480
rect 2963 3470 2967 3474
rect 3003 3476 3007 3480
rect 2992 3469 2996 3473
rect 2770 3459 2774 3463
rect 2690 3455 2696 3459
rect 2795 3456 2799 3460
rect 2802 3459 2806 3463
rect 2820 3459 2824 3463
rect 2842 3456 2846 3460
rect 2867 3456 2871 3460
rect 2877 3459 2881 3463
rect 2893 3459 2897 3463
rect 2913 3456 2917 3460
rect 2920 3459 2924 3463
rect 3058 3475 3062 3479
rect 3078 3478 3082 3482
rect 3097 3474 3101 3478
rect 3226 3485 3230 3489
rect 3239 3488 3243 3494
rect 3276 3488 3280 3494
rect 3289 3490 3293 3494
rect 3313 3494 3317 3498
rect 3387 3494 3391 3498
rect 3297 3488 3301 3494
rect 3334 3488 3338 3494
rect 3350 3488 3354 3494
rect 3371 3488 3375 3494
rect 3408 3488 3412 3494
rect 3421 3490 3425 3494
rect 3445 3494 3449 3498
rect 3519 3494 3523 3498
rect 3429 3488 3433 3494
rect 3466 3488 3470 3494
rect 3482 3488 3486 3494
rect 3503 3488 3507 3494
rect 3540 3488 3544 3494
rect 3553 3490 3557 3494
rect 3577 3494 3581 3498
rect 3647 3501 3653 3505
rect 3729 3501 3733 3505
rect 3738 3501 3742 3505
rect 3788 3501 3792 3505
rect 3813 3501 3817 3505
rect 3844 3501 3848 3505
rect 3561 3488 3565 3494
rect 3598 3488 3602 3494
rect 3614 3490 3618 3494
rect 3729 3493 3733 3497
rect 3772 3494 3776 3498
rect 3794 3493 3801 3497
rect 3844 3494 3848 3498
rect 3715 3489 3719 3493
rect 3747 3489 3751 3493
rect 3765 3489 3769 3493
rect 3822 3489 3826 3493
rect 3837 3489 3841 3493
rect 3865 3489 3869 3493
rect 3116 3475 3120 3479
rect 3135 3475 3139 3479
rect 3148 3476 3152 3480
rect 3170 3475 3174 3479
rect 3178 3476 3182 3480
rect 3190 3476 3194 3480
rect 3239 3475 3243 3479
rect 3255 3475 3259 3481
rect 3289 3481 3293 3485
rect 3276 3475 3280 3479
rect 3297 3475 3301 3479
rect 3313 3475 3317 3481
rect 3334 3475 3338 3479
rect 3350 3475 3354 3479
rect 3371 3475 3375 3479
rect 3387 3475 3391 3481
rect 3421 3481 3425 3485
rect 3408 3475 3412 3479
rect 3429 3475 3433 3479
rect 3445 3475 3449 3481
rect 3466 3475 3470 3479
rect 3482 3475 3486 3479
rect 3503 3475 3507 3479
rect 3519 3475 3523 3481
rect 3553 3481 3557 3485
rect 3540 3475 3544 3479
rect 3561 3475 3565 3479
rect 3577 3475 3581 3481
rect 3598 3475 3602 3479
rect 3614 3475 3618 3479
rect 3710 3477 3714 3481
rect 3004 3459 3008 3463
rect 3030 3459 3034 3463
rect 2287 3448 2291 3452
rect 2338 3448 2342 3452
rect 2388 3448 2392 3452
rect 2419 3448 2423 3452
rect 2470 3448 2474 3452
rect 2520 3448 2524 3452
rect 2551 3448 2555 3452
rect 2602 3448 2606 3452
rect 2652 3448 2656 3452
rect 2726 3449 2732 3453
rect 2778 3449 2782 3453
rect 2796 3449 2800 3453
rect 2827 3449 2831 3453
rect 2849 3449 2853 3453
rect 2914 3449 2918 3453
rect 3056 3456 3060 3460
rect 3063 3459 3067 3463
rect 3081 3459 3085 3463
rect 3103 3456 3107 3460
rect 3128 3456 3132 3460
rect 3138 3459 3142 3463
rect 3154 3459 3158 3463
rect 3174 3456 3178 3460
rect 3181 3459 3185 3463
rect 3232 3464 3236 3468
rect 3269 3462 3273 3466
rect 3289 3462 3293 3466
rect 3333 3462 3337 3466
rect 3364 3464 3368 3468
rect 3401 3462 3405 3466
rect 3421 3462 3425 3466
rect 3465 3462 3469 3466
rect 3496 3464 3500 3468
rect 3533 3462 3537 3466
rect 3553 3462 3557 3466
rect 3597 3462 3601 3466
rect 3742 3475 3746 3479
rect 3762 3478 3766 3482
rect 3781 3474 3785 3478
rect 3800 3475 3804 3479
rect 3819 3475 3823 3479
rect 3832 3476 3836 3480
rect 3968 3501 3972 3505
rect 3990 3501 3994 3505
rect 4049 3501 4053 3505
rect 4074 3501 4078 3505
rect 4105 3501 4109 3505
rect 3990 3493 3994 3497
rect 4033 3494 4037 3498
rect 4055 3493 4062 3497
rect 4105 3494 4109 3498
rect 4008 3489 4012 3493
rect 4026 3489 4030 3493
rect 4083 3489 4087 3493
rect 4098 3489 4102 3493
rect 4126 3489 4130 3493
rect 3929 3485 3933 3489
rect 3854 3475 3858 3479
rect 3862 3476 3866 3480
rect 3874 3476 3878 3480
rect 3908 3470 3912 3474
rect 3948 3476 3952 3480
rect 3937 3469 3941 3473
rect 3715 3459 3719 3463
rect 3635 3455 3641 3459
rect 3740 3456 3744 3460
rect 3747 3459 3751 3463
rect 3765 3459 3769 3463
rect 3787 3456 3791 3460
rect 3812 3456 3816 3460
rect 3822 3459 3826 3463
rect 3838 3459 3842 3463
rect 3858 3456 3862 3460
rect 3865 3459 3869 3463
rect 4003 3475 4007 3479
rect 4023 3478 4027 3482
rect 4042 3474 4046 3478
rect 4061 3475 4065 3479
rect 4080 3475 4084 3479
rect 4093 3476 4097 3480
rect 4115 3475 4119 3479
rect 4123 3476 4127 3480
rect 4135 3476 4139 3480
rect 3949 3459 3953 3463
rect 3975 3459 3979 3463
rect 2974 3449 2978 3453
rect 3013 3449 3017 3453
rect 3057 3449 3061 3453
rect 3088 3449 3092 3453
rect 3110 3449 3114 3453
rect 3175 3449 3179 3453
rect 3232 3448 3236 3452
rect 3283 3448 3287 3452
rect 3333 3448 3337 3452
rect 3364 3448 3368 3452
rect 3415 3448 3419 3452
rect 3465 3448 3469 3452
rect 3496 3448 3500 3452
rect 3547 3448 3551 3452
rect 3597 3448 3601 3452
rect 3671 3449 3677 3453
rect 3723 3449 3727 3453
rect 3741 3449 3745 3453
rect 3772 3449 3776 3453
rect 3794 3449 3798 3453
rect 3859 3449 3863 3453
rect 4001 3456 4005 3460
rect 4008 3459 4012 3463
rect 4026 3459 4030 3463
rect 4048 3456 4052 3460
rect 4073 3456 4077 3460
rect 4083 3459 4087 3463
rect 4099 3459 4103 3463
rect 4119 3456 4123 3460
rect 4126 3459 4130 3463
rect 3919 3449 3923 3453
rect 3958 3449 3962 3453
rect 4002 3449 4006 3453
rect 4033 3449 4037 3453
rect 4055 3449 4059 3453
rect 4120 3449 4124 3453
rect 2281 3441 2285 3445
rect 2669 3441 2673 3445
rect 2678 3442 2684 3446
rect 2769 3442 2773 3446
rect 2803 3442 2807 3446
rect 2820 3442 2824 3446
rect 2876 3442 2880 3446
rect 2893 3442 2897 3446
rect 2921 3442 2925 3446
rect 3004 3442 3008 3446
rect 3030 3442 3034 3446
rect 3064 3442 3068 3446
rect 3081 3442 3085 3446
rect 3137 3442 3141 3446
rect 3154 3442 3158 3446
rect 3182 3442 3186 3446
rect 3226 3441 3230 3445
rect 3614 3441 3618 3445
rect 3623 3442 3629 3446
rect 3714 3442 3718 3446
rect 3748 3442 3752 3446
rect 3765 3442 3769 3446
rect 3821 3442 3825 3446
rect 3838 3442 3842 3446
rect 3866 3442 3870 3446
rect 3949 3442 3953 3446
rect 3975 3442 3979 3446
rect 4009 3442 4013 3446
rect 4026 3442 4030 3446
rect 4082 3442 4086 3446
rect 4099 3442 4103 3446
rect 4127 3442 4131 3446
rect 2404 3434 2409 3438
rect 2537 3434 2541 3438
rect 2714 3435 2720 3439
rect 2778 3435 2782 3439
rect 3012 3435 3016 3439
rect 3198 3436 3202 3440
rect 3210 3436 3214 3440
rect 3349 3434 3354 3438
rect 3482 3434 3486 3438
rect 3659 3435 3665 3439
rect 3723 3435 3727 3439
rect 3957 3435 3961 3439
rect 4143 3436 4147 3440
rect 4155 3436 4159 3440
rect 2412 3427 2416 3431
rect 2702 3427 2708 3431
rect 3022 3428 3026 3432
rect 3187 3428 3191 3432
rect 2396 3422 2400 3426
rect 2428 3422 2432 3426
rect 2750 3421 2756 3425
rect 3357 3427 3361 3431
rect 3647 3427 3653 3431
rect 3967 3428 3971 3432
rect 4132 3428 4136 3432
rect 3341 3422 3345 3426
rect 3373 3422 3377 3426
rect 3695 3421 3701 3425
rect 2265 3414 2269 3418
rect 2396 3414 2400 3418
rect 2428 3414 2432 3418
rect 3341 3414 3345 3418
rect 3373 3414 3377 3418
rect 2412 3407 2416 3411
rect 2669 3407 2673 3411
rect 2738 3407 2744 3411
rect 3070 3407 3074 3411
rect 3106 3407 3110 3411
rect 3173 3407 3177 3411
rect 3357 3407 3361 3411
rect 3614 3407 3618 3411
rect 3683 3407 3689 3411
rect 4015 3407 4019 3411
rect 4051 3407 4055 3411
rect 4118 3407 4122 3411
rect 2669 3399 2673 3403
rect 2678 3400 2684 3404
rect 3056 3400 3060 3404
rect 2396 3395 2400 3399
rect 2428 3395 2432 3399
rect 2412 3391 2416 3395
rect 3070 3393 3074 3397
rect 3120 3393 3124 3397
rect 3173 3393 3177 3397
rect 3614 3399 3618 3403
rect 3623 3400 3629 3404
rect 4001 3400 4005 3404
rect 3341 3395 3345 3399
rect 3373 3395 3377 3399
rect 3357 3391 3361 3395
rect 4015 3393 4019 3397
rect 4065 3393 4069 3397
rect 4118 3393 4122 3397
rect 2404 3384 2409 3388
rect 2538 3384 2542 3388
rect 3093 3382 3097 3386
rect 2287 3377 2291 3381
rect 2323 3377 2327 3381
rect 2390 3377 2394 3381
rect 2419 3377 2423 3381
rect 2455 3377 2459 3381
rect 2522 3377 2526 3381
rect 2551 3377 2555 3381
rect 2587 3377 2591 3381
rect 2654 3377 2658 3381
rect 2738 3377 2744 3381
rect 2678 3370 2684 3374
rect 3064 3373 3068 3377
rect 3077 3376 3081 3382
rect 3114 3376 3118 3382
rect 3127 3378 3131 3382
rect 3151 3382 3155 3386
rect 3349 3384 3354 3388
rect 3483 3384 3487 3388
rect 4038 3382 4042 3386
rect 3135 3376 3139 3382
rect 3172 3376 3176 3382
rect 3188 3376 3192 3382
rect 3232 3377 3236 3381
rect 3268 3377 3272 3381
rect 3335 3377 3339 3381
rect 3364 3377 3368 3381
rect 3400 3377 3404 3381
rect 3467 3377 3471 3381
rect 3496 3377 3500 3381
rect 3532 3377 3536 3381
rect 3599 3377 3603 3381
rect 3683 3377 3689 3381
rect 2287 3363 2291 3367
rect 2337 3363 2341 3367
rect 2390 3363 2394 3367
rect 2419 3363 2423 3367
rect 2469 3363 2473 3367
rect 2522 3363 2526 3367
rect 2551 3363 2555 3367
rect 2601 3363 2605 3367
rect 2654 3363 2658 3367
rect 3077 3363 3081 3367
rect 3093 3363 3097 3369
rect 3127 3369 3131 3373
rect 3114 3363 3118 3367
rect 2310 3352 2314 3356
rect 2281 3343 2285 3347
rect 2294 3346 2298 3352
rect 2331 3346 2335 3352
rect 2344 3348 2348 3352
rect 2368 3352 2372 3356
rect 2442 3352 2446 3356
rect 2352 3346 2356 3352
rect 2389 3346 2393 3352
rect 2405 3346 2409 3352
rect 2426 3346 2430 3352
rect 2463 3346 2467 3352
rect 2476 3348 2480 3352
rect 2500 3352 2504 3356
rect 2574 3352 2578 3356
rect 2484 3346 2488 3352
rect 2521 3346 2525 3352
rect 2537 3346 2541 3352
rect 2558 3346 2562 3352
rect 2595 3346 2599 3352
rect 2608 3348 2612 3352
rect 2632 3352 2636 3356
rect 2616 3346 2620 3352
rect 2653 3346 2657 3352
rect 2669 3348 2673 3352
rect 3135 3363 3139 3367
rect 3151 3363 3155 3369
rect 3623 3370 3629 3374
rect 4009 3373 4013 3377
rect 4022 3376 4026 3382
rect 4059 3376 4063 3382
rect 4072 3378 4076 3382
rect 4096 3382 4100 3386
rect 4080 3376 4084 3382
rect 4117 3376 4121 3382
rect 4133 3376 4137 3382
rect 3172 3363 3176 3367
rect 3188 3363 3192 3367
rect 3232 3363 3236 3367
rect 3282 3363 3286 3367
rect 3335 3363 3339 3367
rect 3364 3363 3368 3367
rect 3414 3363 3418 3367
rect 3467 3363 3471 3367
rect 3496 3363 3500 3367
rect 3546 3363 3550 3367
rect 3599 3363 3603 3367
rect 4022 3363 4026 3367
rect 4038 3363 4042 3369
rect 4072 3369 4076 3373
rect 4059 3363 4063 3367
rect 3070 3352 3074 3356
rect 3107 3350 3111 3354
rect 3127 3350 3131 3354
rect 3171 3350 3175 3354
rect 3255 3352 3259 3356
rect 2294 3333 2298 3337
rect 2310 3333 2314 3339
rect 2344 3339 2348 3343
rect 2331 3333 2335 3337
rect 2352 3333 2356 3337
rect 2368 3333 2372 3339
rect 2389 3333 2393 3337
rect 2405 3333 2409 3337
rect 2426 3333 2430 3337
rect 2442 3333 2446 3339
rect 2476 3339 2480 3343
rect 2463 3333 2467 3337
rect 2484 3333 2488 3337
rect 2500 3333 2504 3339
rect 2521 3333 2525 3337
rect 2537 3333 2541 3337
rect 2558 3333 2562 3337
rect 2574 3333 2578 3339
rect 2608 3339 2612 3343
rect 2595 3333 2599 3337
rect 2616 3333 2620 3337
rect 2632 3333 2636 3339
rect 2690 3343 2696 3347
rect 3226 3343 3230 3347
rect 3239 3346 3243 3352
rect 3276 3346 3280 3352
rect 3289 3348 3293 3352
rect 3313 3352 3317 3356
rect 3387 3352 3391 3356
rect 3297 3346 3301 3352
rect 3334 3346 3338 3352
rect 3350 3346 3354 3352
rect 3371 3346 3375 3352
rect 3408 3346 3412 3352
rect 3421 3348 3425 3352
rect 3445 3352 3449 3356
rect 3519 3352 3523 3356
rect 3429 3346 3433 3352
rect 3466 3346 3470 3352
rect 3482 3346 3486 3352
rect 3503 3346 3507 3352
rect 3540 3346 3544 3352
rect 3553 3348 3557 3352
rect 3577 3352 3581 3356
rect 3561 3346 3565 3352
rect 3598 3346 3602 3352
rect 3614 3348 3618 3352
rect 4080 3363 4084 3367
rect 4096 3363 4100 3369
rect 4117 3363 4121 3367
rect 4133 3363 4137 3367
rect 4015 3352 4019 3356
rect 4052 3350 4056 3354
rect 4072 3350 4076 3354
rect 4116 3350 4120 3354
rect 2653 3333 2657 3337
rect 2669 3333 2673 3337
rect 2726 3336 2732 3340
rect 3070 3336 3074 3340
rect 3121 3336 3125 3340
rect 3171 3336 3175 3340
rect 3239 3333 3243 3337
rect 3255 3333 3259 3339
rect 3289 3339 3293 3343
rect 3276 3333 3280 3337
rect 2287 3322 2291 3326
rect 2324 3320 2328 3324
rect 2344 3320 2348 3324
rect 2388 3320 2392 3324
rect 2419 3322 2423 3326
rect 2456 3320 2460 3324
rect 2476 3320 2480 3324
rect 2520 3320 2524 3324
rect 2551 3322 2555 3326
rect 2588 3320 2592 3324
rect 2608 3320 2612 3324
rect 2652 3320 2656 3324
rect 3063 3328 3067 3332
rect 3188 3329 3192 3333
rect 3297 3333 3301 3337
rect 3313 3333 3317 3339
rect 3334 3333 3338 3337
rect 3350 3333 3354 3337
rect 3371 3333 3375 3337
rect 3387 3333 3391 3339
rect 3421 3339 3425 3343
rect 3408 3333 3412 3337
rect 3429 3333 3433 3337
rect 3445 3333 3449 3339
rect 3466 3333 3470 3337
rect 3482 3333 3486 3337
rect 3503 3333 3507 3337
rect 3519 3333 3523 3339
rect 3553 3339 3557 3343
rect 3540 3333 3544 3337
rect 3561 3333 3565 3337
rect 3577 3333 3581 3339
rect 3635 3343 3641 3347
rect 3598 3333 3602 3337
rect 3614 3333 3618 3337
rect 3671 3336 3677 3340
rect 4015 3336 4019 3340
rect 4066 3336 4070 3340
rect 4116 3336 4120 3340
rect 2738 3321 2744 3325
rect 3070 3321 3074 3325
rect 3106 3321 3110 3325
rect 3173 3321 3177 3325
rect 2690 3313 2696 3317
rect 3056 3314 3060 3318
rect 3232 3322 3236 3326
rect 3269 3320 3273 3324
rect 3289 3320 3293 3324
rect 3333 3320 3337 3324
rect 3364 3322 3368 3326
rect 3401 3320 3405 3324
rect 3421 3320 3425 3324
rect 3465 3320 3469 3324
rect 3496 3322 3500 3326
rect 3533 3320 3537 3324
rect 3553 3320 3557 3324
rect 3597 3320 3601 3324
rect 4008 3328 4012 3332
rect 4133 3329 4137 3333
rect 3683 3321 3689 3325
rect 4015 3321 4019 3325
rect 4051 3321 4055 3325
rect 4118 3321 4122 3325
rect 2287 3306 2291 3310
rect 2338 3306 2342 3310
rect 2388 3306 2392 3310
rect 2419 3306 2423 3310
rect 2470 3306 2474 3310
rect 2520 3306 2524 3310
rect 2551 3306 2555 3310
rect 2602 3306 2606 3310
rect 2652 3306 2656 3310
rect 2726 3306 2732 3310
rect 3070 3307 3074 3311
rect 3120 3307 3124 3311
rect 3173 3307 3177 3311
rect 3635 3313 3641 3317
rect 4001 3314 4005 3318
rect 3232 3306 3236 3310
rect 3283 3306 3287 3310
rect 3333 3306 3337 3310
rect 3364 3306 3368 3310
rect 3415 3306 3419 3310
rect 3465 3306 3469 3310
rect 3496 3306 3500 3310
rect 3547 3306 3551 3310
rect 3597 3306 3601 3310
rect 3671 3306 3677 3310
rect 4015 3307 4019 3311
rect 4065 3307 4069 3311
rect 4118 3307 4122 3311
rect 2280 3299 2284 3303
rect 2669 3299 2673 3303
rect 3093 3296 3097 3300
rect 2287 3291 2291 3295
rect 2323 3291 2327 3295
rect 2390 3291 2394 3295
rect 2419 3291 2423 3295
rect 2455 3291 2459 3295
rect 2522 3291 2526 3295
rect 2551 3291 2555 3295
rect 2587 3291 2591 3295
rect 2654 3291 2658 3295
rect 2738 3291 2744 3295
rect 2678 3284 2684 3288
rect 3064 3287 3068 3291
rect 3077 3290 3081 3296
rect 3114 3290 3118 3296
rect 3127 3292 3131 3296
rect 3151 3296 3155 3300
rect 3225 3299 3229 3303
rect 3614 3299 3618 3303
rect 4038 3296 4042 3300
rect 3135 3290 3139 3296
rect 3172 3290 3176 3296
rect 3188 3292 3192 3296
rect 3210 3290 3214 3294
rect 3232 3291 3236 3295
rect 3268 3291 3272 3295
rect 3335 3291 3339 3295
rect 3364 3291 3368 3295
rect 3400 3291 3404 3295
rect 3467 3291 3471 3295
rect 3496 3291 3500 3295
rect 3532 3291 3536 3295
rect 3599 3291 3603 3295
rect 3683 3291 3689 3295
rect 2287 3277 2291 3281
rect 2337 3277 2341 3281
rect 2390 3277 2394 3281
rect 2419 3277 2423 3281
rect 2469 3277 2473 3281
rect 2522 3277 2526 3281
rect 2551 3277 2555 3281
rect 2601 3277 2605 3281
rect 2654 3277 2658 3281
rect 3077 3277 3081 3281
rect 3093 3277 3097 3283
rect 3127 3283 3131 3287
rect 3114 3277 3118 3281
rect 2310 3266 2314 3270
rect 2281 3257 2285 3261
rect 2294 3260 2298 3266
rect 2331 3260 2335 3266
rect 2344 3262 2348 3266
rect 2368 3266 2372 3270
rect 2442 3266 2446 3270
rect 2352 3260 2356 3266
rect 2389 3260 2393 3266
rect 2405 3260 2409 3266
rect 2426 3260 2430 3266
rect 2463 3260 2467 3266
rect 2476 3262 2480 3266
rect 2500 3266 2504 3270
rect 2574 3266 2578 3270
rect 2484 3260 2488 3266
rect 2521 3260 2525 3266
rect 2537 3260 2541 3266
rect 2558 3260 2562 3266
rect 2595 3260 2599 3266
rect 2608 3262 2612 3266
rect 2632 3266 2636 3270
rect 2616 3260 2620 3266
rect 2653 3260 2657 3266
rect 2669 3262 2673 3266
rect 3135 3277 3139 3281
rect 3151 3277 3155 3283
rect 3172 3277 3176 3281
rect 3188 3277 3192 3286
rect 3623 3284 3629 3288
rect 4009 3287 4013 3291
rect 4022 3290 4026 3296
rect 4059 3290 4063 3296
rect 4072 3292 4076 3296
rect 4096 3296 4100 3300
rect 4080 3290 4084 3296
rect 4117 3290 4121 3296
rect 4133 3292 4137 3296
rect 4155 3290 4159 3294
rect 3210 3274 3214 3278
rect 3232 3277 3236 3281
rect 3282 3277 3286 3281
rect 3335 3277 3339 3281
rect 3364 3277 3368 3281
rect 3414 3277 3418 3281
rect 3467 3277 3471 3281
rect 3496 3277 3500 3281
rect 3546 3277 3550 3281
rect 3599 3277 3603 3281
rect 4022 3277 4026 3281
rect 4038 3277 4042 3283
rect 4072 3283 4076 3287
rect 4059 3277 4063 3281
rect 3070 3266 3074 3270
rect 3107 3264 3111 3268
rect 3127 3264 3131 3268
rect 3171 3264 3175 3268
rect 3255 3266 3259 3270
rect 2294 3247 2298 3251
rect 2310 3247 2314 3253
rect 2344 3253 2348 3257
rect 2331 3247 2335 3251
rect 2352 3247 2356 3251
rect 2368 3247 2372 3253
rect 2389 3247 2393 3251
rect 2405 3247 2409 3251
rect 2426 3247 2430 3251
rect 2442 3247 2446 3253
rect 2476 3253 2480 3257
rect 2463 3247 2467 3251
rect 2484 3247 2488 3251
rect 2500 3247 2504 3253
rect 2521 3247 2525 3251
rect 2537 3247 2541 3251
rect 2558 3247 2562 3251
rect 2574 3247 2578 3253
rect 2608 3253 2612 3257
rect 2595 3247 2599 3251
rect 2616 3247 2620 3251
rect 2632 3247 2636 3253
rect 2690 3257 2696 3261
rect 3226 3257 3230 3261
rect 3239 3260 3243 3266
rect 3276 3260 3280 3266
rect 3289 3262 3293 3266
rect 3313 3266 3317 3270
rect 3387 3266 3391 3270
rect 3297 3260 3301 3266
rect 3334 3260 3338 3266
rect 3350 3260 3354 3266
rect 3371 3260 3375 3266
rect 3408 3260 3412 3266
rect 3421 3262 3425 3266
rect 3445 3266 3449 3270
rect 3519 3266 3523 3270
rect 3429 3260 3433 3266
rect 3466 3260 3470 3266
rect 3482 3260 3486 3266
rect 3503 3260 3507 3266
rect 3540 3260 3544 3266
rect 3553 3262 3557 3266
rect 3577 3266 3581 3270
rect 3561 3260 3565 3266
rect 3598 3260 3602 3266
rect 3614 3262 3618 3266
rect 4080 3277 4084 3281
rect 4096 3277 4100 3283
rect 4117 3277 4121 3281
rect 4133 3277 4137 3286
rect 4155 3274 4159 3278
rect 4015 3266 4019 3270
rect 4052 3264 4056 3268
rect 4072 3264 4076 3268
rect 4116 3264 4120 3268
rect 2653 3247 2657 3251
rect 2669 3247 2673 3251
rect 2726 3250 2732 3254
rect 3070 3250 3074 3254
rect 3121 3250 3125 3254
rect 3171 3250 3175 3254
rect 3239 3247 3243 3251
rect 3255 3247 3259 3253
rect 3289 3253 3293 3257
rect 3276 3247 3280 3251
rect 3297 3247 3301 3251
rect 3313 3247 3317 3253
rect 3334 3247 3338 3251
rect 3350 3247 3354 3251
rect 3371 3247 3375 3251
rect 3387 3247 3391 3253
rect 3421 3253 3425 3257
rect 3408 3247 3412 3251
rect 3429 3247 3433 3251
rect 3445 3247 3449 3253
rect 3466 3247 3470 3251
rect 3482 3247 3486 3251
rect 3503 3247 3507 3251
rect 3519 3247 3523 3253
rect 3553 3253 3557 3257
rect 3540 3247 3544 3251
rect 3561 3247 3565 3251
rect 3577 3247 3581 3253
rect 3635 3257 3641 3261
rect 3598 3247 3602 3251
rect 3614 3247 3618 3251
rect 3671 3250 3677 3254
rect 4015 3250 4019 3254
rect 4066 3250 4070 3254
rect 4116 3250 4120 3254
rect 2287 3236 2291 3240
rect 2324 3234 2328 3238
rect 2344 3234 2348 3238
rect 2388 3234 2392 3238
rect 2419 3236 2423 3240
rect 2456 3234 2460 3238
rect 2476 3234 2480 3238
rect 2520 3234 2524 3238
rect 2551 3236 2555 3240
rect 2588 3234 2592 3238
rect 2608 3234 2612 3238
rect 2652 3234 2656 3238
rect 3232 3236 3236 3240
rect 3269 3234 3273 3238
rect 3289 3234 3293 3238
rect 3333 3234 3337 3238
rect 3364 3236 3368 3240
rect 3401 3234 3405 3238
rect 3421 3234 3425 3238
rect 3465 3234 3469 3238
rect 3496 3236 3500 3240
rect 3533 3234 3537 3238
rect 3553 3234 3557 3238
rect 3597 3234 3601 3238
rect 2690 3227 2696 3231
rect 3635 3227 3641 3231
rect 2287 3220 2291 3224
rect 2338 3220 2342 3224
rect 2388 3220 2392 3224
rect 2419 3220 2423 3224
rect 2470 3220 2474 3224
rect 2520 3220 2524 3224
rect 2551 3220 2555 3224
rect 2602 3220 2606 3224
rect 2652 3220 2656 3224
rect 2726 3220 2732 3224
rect 3232 3220 3236 3224
rect 3283 3220 3287 3224
rect 3333 3220 3337 3224
rect 3364 3220 3368 3224
rect 3415 3220 3419 3224
rect 3465 3220 3469 3224
rect 3496 3220 3500 3224
rect 3547 3220 3551 3224
rect 3597 3220 3601 3224
rect 3671 3220 3677 3224
rect 2280 3213 2284 3217
rect 2669 3213 2673 3217
rect 3225 3213 3229 3217
rect 3614 3213 3618 3217
rect 2405 3206 2409 3210
rect 2513 3206 2517 3210
rect 2537 3206 2541 3210
rect 3350 3206 3354 3210
rect 3458 3206 3462 3210
rect 3482 3206 3486 3210
rect 2529 3199 2533 3203
rect 2513 3195 2517 3199
rect 2545 3195 2549 3199
rect 3474 3199 3478 3203
rect 3458 3195 3462 3199
rect 3490 3195 3494 3199
rect 2513 3188 2517 3192
rect 2545 3188 2549 3192
rect 3210 3188 3214 3192
rect 3458 3188 3462 3192
rect 3490 3188 3494 3192
rect 4155 3188 4159 3192
rect 2529 3181 2533 3185
rect 2669 3181 2673 3185
rect 3474 3181 3478 3185
rect 3614 3181 3618 3185
rect 2669 3173 2673 3177
rect 3614 3173 3618 3177
rect 2513 3169 2517 3173
rect 2545 3169 2549 3173
rect 2529 3165 2533 3169
rect 3458 3169 3462 3173
rect 3490 3169 3494 3173
rect 3474 3165 3478 3169
rect 2405 3158 2409 3162
rect 2513 3158 2517 3162
rect 2537 3158 2541 3162
rect 3350 3158 3354 3162
rect 3458 3158 3462 3162
rect 3482 3158 3486 3162
rect 2287 3151 2291 3155
rect 2323 3151 2327 3155
rect 2390 3151 2394 3155
rect 2419 3151 2423 3155
rect 2455 3151 2459 3155
rect 2522 3151 2526 3155
rect 2551 3151 2555 3155
rect 2587 3151 2591 3155
rect 2654 3151 2658 3155
rect 2738 3151 2744 3155
rect 3232 3151 3236 3155
rect 3268 3151 3272 3155
rect 3335 3151 3339 3155
rect 3364 3151 3368 3155
rect 3400 3151 3404 3155
rect 3467 3151 3471 3155
rect 3496 3151 3500 3155
rect 3532 3151 3536 3155
rect 3599 3151 3603 3155
rect 3683 3151 3689 3155
rect 2678 3144 2684 3148
rect 3623 3144 3629 3148
rect 2287 3137 2291 3141
rect 2337 3137 2341 3141
rect 2390 3137 2394 3141
rect 2419 3137 2423 3141
rect 2469 3137 2473 3141
rect 2522 3137 2526 3141
rect 2551 3137 2555 3141
rect 2601 3137 2605 3141
rect 2654 3137 2658 3141
rect 3232 3137 3236 3141
rect 3282 3137 3286 3141
rect 3335 3137 3339 3141
rect 3364 3137 3368 3141
rect 3414 3137 3418 3141
rect 3467 3137 3471 3141
rect 3496 3137 3500 3141
rect 3546 3137 3550 3141
rect 3599 3137 3603 3141
rect 2310 3126 2314 3130
rect 2281 3117 2285 3121
rect 2294 3120 2298 3126
rect 2331 3120 2335 3126
rect 2344 3122 2348 3126
rect 2368 3126 2372 3130
rect 2442 3126 2446 3130
rect 2352 3120 2356 3126
rect 2389 3120 2393 3126
rect 2405 3120 2409 3126
rect 2426 3120 2430 3126
rect 2463 3120 2467 3126
rect 2476 3122 2480 3126
rect 2500 3126 2504 3130
rect 2574 3126 2578 3130
rect 2484 3120 2488 3126
rect 2521 3120 2525 3126
rect 2537 3120 2541 3126
rect 2558 3120 2562 3126
rect 2595 3120 2599 3126
rect 2608 3122 2612 3126
rect 2632 3126 2636 3130
rect 3255 3126 3259 3130
rect 2616 3120 2620 3126
rect 2653 3120 2657 3126
rect 2669 3122 2673 3126
rect 2294 3107 2298 3111
rect 2310 3107 2314 3113
rect 2344 3113 2348 3117
rect 2331 3107 2335 3111
rect 2352 3107 2356 3111
rect 2368 3107 2372 3113
rect 2389 3107 2393 3111
rect 2405 3107 2409 3111
rect 2426 3107 2430 3111
rect 2442 3107 2446 3113
rect 2476 3113 2480 3117
rect 2463 3107 2467 3111
rect 2484 3107 2488 3111
rect 2500 3107 2504 3113
rect 2521 3107 2525 3111
rect 2537 3107 2541 3111
rect 2558 3107 2562 3111
rect 2574 3107 2578 3113
rect 2608 3113 2612 3117
rect 2595 3107 2599 3111
rect 2616 3107 2620 3111
rect 2632 3107 2636 3113
rect 3226 3117 3230 3121
rect 3239 3120 3243 3126
rect 3276 3120 3280 3126
rect 3289 3122 3293 3126
rect 3313 3126 3317 3130
rect 3387 3126 3391 3130
rect 3297 3120 3301 3126
rect 3334 3120 3338 3126
rect 3350 3120 3354 3126
rect 3371 3120 3375 3126
rect 3408 3120 3412 3126
rect 3421 3122 3425 3126
rect 3445 3126 3449 3130
rect 3519 3126 3523 3130
rect 3429 3120 3433 3126
rect 3466 3120 3470 3126
rect 3482 3120 3486 3126
rect 3503 3120 3507 3126
rect 3540 3120 3544 3126
rect 3553 3122 3557 3126
rect 3577 3126 3581 3130
rect 3561 3120 3565 3126
rect 3598 3120 3602 3126
rect 3614 3122 3618 3126
rect 2653 3107 2657 3111
rect 2669 3107 2673 3111
rect 3239 3107 3243 3111
rect 3255 3107 3259 3113
rect 3289 3113 3293 3117
rect 3276 3107 3280 3111
rect 3297 3107 3301 3111
rect 3313 3107 3317 3113
rect 3334 3107 3338 3111
rect 3350 3107 3354 3111
rect 3371 3107 3375 3111
rect 3387 3107 3391 3113
rect 3421 3113 3425 3117
rect 3408 3107 3412 3111
rect 3429 3107 3433 3111
rect 3445 3107 3449 3113
rect 3466 3107 3470 3111
rect 3482 3107 3486 3111
rect 3503 3107 3507 3111
rect 3519 3107 3523 3113
rect 3553 3113 3557 3117
rect 3540 3107 3544 3111
rect 3561 3107 3565 3111
rect 3577 3107 3581 3113
rect 3598 3107 3602 3111
rect 3614 3107 3618 3111
rect 2287 3096 2291 3100
rect 2324 3094 2328 3098
rect 2344 3094 2348 3098
rect 2388 3094 2392 3098
rect 2419 3096 2423 3100
rect 2456 3094 2460 3098
rect 2476 3094 2480 3098
rect 2520 3094 2524 3098
rect 2551 3096 2555 3100
rect 2588 3094 2592 3098
rect 2608 3094 2612 3098
rect 2652 3094 2656 3098
rect 3232 3096 3236 3100
rect 3269 3094 3273 3098
rect 3289 3094 3293 3098
rect 3333 3094 3337 3098
rect 3364 3096 3368 3100
rect 3401 3094 3405 3098
rect 3421 3094 3425 3098
rect 3465 3094 3469 3098
rect 3496 3096 3500 3100
rect 3533 3094 3537 3098
rect 3553 3094 3557 3098
rect 3597 3094 3601 3098
rect 2690 3087 2696 3091
rect 3635 3087 3641 3091
rect 2287 3080 2291 3084
rect 2338 3080 2342 3084
rect 2388 3080 2392 3084
rect 2419 3080 2423 3084
rect 2470 3080 2474 3084
rect 2520 3080 2524 3084
rect 2551 3080 2555 3084
rect 2602 3080 2606 3084
rect 2652 3080 2656 3084
rect 2726 3080 2732 3084
rect 3232 3080 3236 3084
rect 3283 3080 3287 3084
rect 3333 3080 3337 3084
rect 3364 3080 3368 3084
rect 3415 3080 3419 3084
rect 3465 3080 3469 3084
rect 3496 3080 3500 3084
rect 3547 3080 3551 3084
rect 3597 3080 3601 3084
rect 3671 3080 3677 3084
rect 2738 3072 2744 3076
rect 2771 3072 2775 3076
rect 2807 3072 2811 3076
rect 2874 3072 2878 3076
rect 2903 3072 2907 3076
rect 2939 3072 2943 3076
rect 3006 3072 3010 3076
rect 3035 3072 3039 3076
rect 3071 3072 3075 3076
rect 3138 3072 3142 3076
rect 3167 3072 3171 3076
rect 3203 3072 3207 3076
rect 3270 3072 3274 3076
rect 3683 3072 3689 3076
rect 3716 3072 3720 3076
rect 3752 3072 3756 3076
rect 3819 3072 3823 3076
rect 3848 3072 3852 3076
rect 3884 3072 3888 3076
rect 3951 3072 3955 3076
rect 3980 3072 3984 3076
rect 4016 3072 4020 3076
rect 4083 3072 4087 3076
rect 4112 3072 4116 3076
rect 4148 3072 4152 3076
rect 4215 3072 4219 3076
rect 2678 3065 2684 3069
rect 3623 3065 3629 3069
rect 2771 3058 2775 3062
rect 2821 3058 2825 3062
rect 2874 3058 2878 3062
rect 2903 3058 2907 3062
rect 2953 3058 2957 3062
rect 3006 3058 3010 3062
rect 3035 3058 3039 3062
rect 3085 3058 3089 3062
rect 3138 3058 3142 3062
rect 3167 3058 3171 3062
rect 3217 3058 3221 3062
rect 3270 3058 3274 3062
rect 3716 3058 3720 3062
rect 3766 3058 3770 3062
rect 3819 3058 3823 3062
rect 3848 3058 3852 3062
rect 3898 3058 3902 3062
rect 3951 3058 3955 3062
rect 3980 3058 3984 3062
rect 4030 3058 4034 3062
rect 4083 3058 4087 3062
rect 4112 3058 4116 3062
rect 4162 3058 4166 3062
rect 4215 3058 4219 3062
rect 2794 3047 2798 3051
rect 2419 3039 2423 3043
rect 2455 3039 2459 3043
rect 2522 3039 2526 3043
rect 2738 3039 2744 3043
rect 2765 3038 2769 3042
rect 2778 3041 2782 3047
rect 2815 3041 2819 3047
rect 2828 3043 2832 3047
rect 2852 3047 2856 3051
rect 2926 3047 2930 3051
rect 2836 3041 2840 3047
rect 2873 3041 2877 3047
rect 2889 3043 2893 3047
rect 2678 3032 2684 3036
rect 2419 3025 2423 3029
rect 2469 3025 2473 3029
rect 2522 3025 2526 3029
rect 2778 3028 2782 3032
rect 2794 3028 2798 3034
rect 2828 3034 2832 3038
rect 2815 3028 2819 3032
rect 2836 3028 2840 3032
rect 2852 3028 2856 3034
rect 2897 3038 2901 3042
rect 2910 3041 2914 3047
rect 2947 3041 2951 3047
rect 2960 3043 2964 3047
rect 2984 3047 2988 3051
rect 3058 3047 3062 3051
rect 2968 3041 2972 3047
rect 3005 3041 3009 3047
rect 3021 3043 3025 3047
rect 2873 3028 2877 3032
rect 2889 3028 2893 3032
rect 2910 3028 2914 3032
rect 2926 3028 2930 3034
rect 2960 3034 2964 3038
rect 2947 3028 2951 3032
rect 2968 3028 2972 3032
rect 2984 3028 2988 3034
rect 3029 3038 3033 3042
rect 3042 3041 3046 3047
rect 3079 3041 3083 3047
rect 3092 3043 3096 3047
rect 3116 3047 3120 3051
rect 3190 3047 3194 3051
rect 3100 3041 3104 3047
rect 3137 3041 3141 3047
rect 3153 3043 3157 3047
rect 3005 3028 3009 3032
rect 3021 3028 3025 3032
rect 3042 3028 3046 3032
rect 3058 3028 3062 3034
rect 3092 3034 3096 3038
rect 3079 3028 3083 3032
rect 3100 3028 3104 3032
rect 3116 3028 3120 3034
rect 3161 3038 3165 3042
rect 3174 3041 3178 3047
rect 3211 3041 3215 3047
rect 3224 3043 3228 3047
rect 3248 3047 3252 3051
rect 3739 3047 3743 3051
rect 3232 3041 3236 3047
rect 3269 3041 3273 3047
rect 3285 3043 3289 3047
rect 3364 3039 3368 3043
rect 3400 3039 3404 3043
rect 3467 3039 3471 3043
rect 3683 3039 3689 3043
rect 3137 3028 3141 3032
rect 3153 3028 3157 3032
rect 3174 3028 3178 3032
rect 3190 3028 3194 3034
rect 3224 3034 3228 3038
rect 3211 3028 3215 3032
rect 2442 3014 2446 3018
rect 2404 3005 2408 3009
rect 2426 3008 2430 3014
rect 2463 3008 2467 3014
rect 2476 3010 2480 3014
rect 2500 3014 2504 3018
rect 2484 3008 2488 3014
rect 2521 3008 2525 3014
rect 2537 3008 2541 3014
rect 2771 3017 2775 3021
rect 2808 3015 2812 3019
rect 2828 3015 2832 3019
rect 2872 3015 2876 3019
rect 2903 3017 2907 3021
rect 2940 3015 2944 3019
rect 2960 3015 2964 3019
rect 3004 3015 3008 3019
rect 3035 3017 3039 3021
rect 3072 3015 3076 3019
rect 3092 3015 3096 3019
rect 3136 3015 3140 3019
rect 3153 3020 3157 3024
rect 3232 3028 3236 3032
rect 3248 3028 3252 3034
rect 3710 3038 3714 3042
rect 3723 3041 3727 3047
rect 3760 3041 3764 3047
rect 3773 3043 3777 3047
rect 3797 3047 3801 3051
rect 3871 3047 3875 3051
rect 3781 3041 3785 3047
rect 3818 3041 3822 3047
rect 3834 3043 3838 3047
rect 3623 3032 3629 3036
rect 3269 3028 3273 3032
rect 3285 3028 3289 3032
rect 3167 3017 3171 3021
rect 3204 3015 3208 3019
rect 3224 3015 3228 3019
rect 3268 3015 3272 3019
rect 3285 3020 3289 3024
rect 3364 3025 3368 3029
rect 3414 3025 3418 3029
rect 3467 3025 3471 3029
rect 3723 3028 3727 3032
rect 3739 3028 3743 3034
rect 3773 3034 3777 3038
rect 3760 3028 3764 3032
rect 3781 3028 3785 3032
rect 3797 3028 3801 3034
rect 3842 3038 3846 3042
rect 3855 3041 3859 3047
rect 3892 3041 3896 3047
rect 3905 3043 3909 3047
rect 3929 3047 3933 3051
rect 4003 3047 4007 3051
rect 3913 3041 3917 3047
rect 3950 3041 3954 3047
rect 3966 3043 3970 3047
rect 3818 3028 3822 3032
rect 3834 3028 3838 3032
rect 3855 3028 3859 3032
rect 3871 3028 3875 3034
rect 3905 3034 3909 3038
rect 3892 3028 3896 3032
rect 3913 3028 3917 3032
rect 3929 3028 3933 3034
rect 3974 3038 3978 3042
rect 3987 3041 3991 3047
rect 4024 3041 4028 3047
rect 4037 3043 4041 3047
rect 4061 3047 4065 3051
rect 4135 3047 4139 3051
rect 4045 3041 4049 3047
rect 4082 3041 4086 3047
rect 4098 3043 4102 3047
rect 3950 3028 3954 3032
rect 3966 3028 3970 3032
rect 3987 3028 3991 3032
rect 4003 3028 4007 3034
rect 4037 3034 4041 3038
rect 4024 3028 4028 3032
rect 4045 3028 4049 3032
rect 4061 3028 4065 3034
rect 4106 3038 4110 3042
rect 4119 3041 4123 3047
rect 4156 3041 4160 3047
rect 4169 3043 4173 3047
rect 4193 3047 4197 3051
rect 4177 3041 4181 3047
rect 4214 3041 4218 3047
rect 4230 3043 4234 3047
rect 4082 3028 4086 3032
rect 4098 3028 4102 3032
rect 4119 3028 4123 3032
rect 4135 3028 4139 3034
rect 4169 3034 4173 3038
rect 4156 3028 4160 3032
rect 3387 3014 3391 3018
rect 2690 3008 2696 3012
rect 2426 2995 2430 2999
rect 2442 2995 2446 3001
rect 2476 3001 2480 3005
rect 2463 2995 2467 2999
rect 2484 2995 2488 2999
rect 2500 2995 2504 3001
rect 3349 3005 3353 3009
rect 3371 3008 3375 3014
rect 3408 3008 3412 3014
rect 3421 3010 3425 3014
rect 3445 3014 3449 3018
rect 3429 3008 3433 3014
rect 3466 3008 3470 3014
rect 3482 3008 3486 3014
rect 3716 3017 3720 3021
rect 3753 3015 3757 3019
rect 3773 3015 3777 3019
rect 3817 3015 3821 3019
rect 3848 3017 3852 3021
rect 3885 3015 3889 3019
rect 3905 3015 3909 3019
rect 3949 3015 3953 3019
rect 3980 3017 3984 3021
rect 4017 3015 4021 3019
rect 4037 3015 4041 3019
rect 4081 3015 4085 3019
rect 4098 3020 4102 3024
rect 4177 3028 4181 3032
rect 4193 3028 4197 3034
rect 4214 3028 4218 3032
rect 4230 3028 4234 3032
rect 4112 3017 4116 3021
rect 4149 3015 4153 3019
rect 4169 3015 4173 3019
rect 4213 3015 4217 3019
rect 4230 3020 4234 3024
rect 3635 3008 3641 3012
rect 2726 3001 2732 3005
rect 2771 3001 2775 3005
rect 2822 3001 2826 3005
rect 2872 3001 2876 3005
rect 2903 3001 2907 3005
rect 2954 3001 2958 3005
rect 3004 3001 3008 3005
rect 3035 3001 3039 3005
rect 3086 3001 3090 3005
rect 3136 3001 3140 3005
rect 3167 3001 3171 3005
rect 3218 3001 3222 3005
rect 3268 3001 3272 3005
rect 2521 2995 2525 2999
rect 2537 2995 2541 2999
rect 3371 2995 3375 2999
rect 3387 2995 3391 3001
rect 3421 3001 3425 3005
rect 3408 2995 3412 2999
rect 2419 2984 2423 2988
rect 2456 2982 2460 2986
rect 2476 2982 2480 2986
rect 2520 2982 2524 2986
rect 2678 2988 2684 2992
rect 2769 2988 2773 2992
rect 2803 2988 2807 2992
rect 2820 2988 2824 2992
rect 2876 2988 2880 2992
rect 2893 2988 2897 2992
rect 2921 2988 2925 2992
rect 3429 2995 3433 2999
rect 3445 2995 3449 3001
rect 3671 3001 3677 3005
rect 3716 3001 3720 3005
rect 3767 3001 3771 3005
rect 3817 3001 3821 3005
rect 3848 3001 3852 3005
rect 3899 3001 3903 3005
rect 3949 3001 3953 3005
rect 3980 3001 3984 3005
rect 4031 3001 4035 3005
rect 4081 3001 4085 3005
rect 4112 3001 4116 3005
rect 4163 3001 4167 3005
rect 4213 3001 4217 3005
rect 3466 2995 3470 2999
rect 3482 2995 3486 2999
rect 2714 2981 2720 2985
rect 2796 2981 2800 2985
rect 2827 2981 2831 2985
rect 2849 2981 2853 2985
rect 2914 2981 2918 2985
rect 2690 2975 2696 2979
rect 2419 2968 2423 2972
rect 2470 2968 2474 2972
rect 2520 2968 2524 2972
rect 2726 2968 2732 2972
rect 2770 2971 2774 2975
rect 2795 2974 2799 2978
rect 2802 2971 2806 2975
rect 2820 2971 2824 2975
rect 2842 2974 2846 2978
rect 2867 2974 2871 2978
rect 2877 2971 2881 2975
rect 2893 2971 2897 2975
rect 2913 2974 2917 2978
rect 2920 2971 2924 2975
rect 2984 2981 2988 2985
rect 2537 2961 2541 2965
rect 2404 2952 2408 2956
rect 2529 2954 2533 2958
rect 2553 2954 2557 2958
rect 2763 2954 2767 2958
rect 2412 2945 2416 2949
rect 2553 2945 2557 2949
rect 2797 2955 2801 2959
rect 2817 2952 2821 2956
rect 2836 2956 2840 2960
rect 2938 2967 2942 2971
rect 2953 2967 2957 2971
rect 2855 2955 2859 2959
rect 2874 2955 2878 2959
rect 2887 2954 2891 2958
rect 2909 2955 2913 2959
rect 2917 2954 2921 2958
rect 2929 2954 2933 2958
rect 2770 2941 2774 2945
rect 2802 2941 2806 2945
rect 2820 2941 2824 2945
rect 2877 2941 2881 2945
rect 2892 2941 2896 2945
rect 2920 2941 2924 2945
rect 2419 2937 2423 2941
rect 2486 2937 2490 2941
rect 2522 2937 2526 2941
rect 2738 2937 2744 2941
rect 2784 2937 2788 2941
rect 2827 2936 2831 2940
rect 2849 2937 2856 2941
rect 2899 2936 2903 2940
rect 2678 2930 2684 2934
rect 2419 2923 2423 2927
rect 2472 2923 2476 2927
rect 2522 2923 2526 2927
rect 2702 2929 2708 2933
rect 2784 2929 2788 2933
rect 2843 2929 2847 2933
rect 2868 2929 2872 2933
rect 2899 2929 2903 2933
rect 2992 2959 2996 2967
rect 3065 2981 3069 2985
rect 3019 2967 3023 2971
rect 3034 2967 3038 2971
rect 3364 2984 3368 2988
rect 3401 2982 3405 2986
rect 3421 2982 3425 2986
rect 3465 2982 3469 2986
rect 3623 2988 3629 2992
rect 3714 2988 3718 2992
rect 3748 2988 3752 2992
rect 3765 2988 3769 2992
rect 3821 2988 3825 2992
rect 3838 2988 3842 2992
rect 3866 2988 3870 2992
rect 3659 2981 3665 2985
rect 3741 2981 3745 2985
rect 3772 2981 3776 2985
rect 3794 2981 3798 2985
rect 3859 2981 3863 2985
rect 3015 2959 3019 2963
rect 2961 2953 2965 2957
rect 2974 2945 2978 2949
rect 3073 2959 3077 2967
rect 3635 2975 3641 2979
rect 3364 2968 3368 2972
rect 3415 2968 3419 2972
rect 3465 2968 3469 2972
rect 3671 2968 3677 2972
rect 3715 2971 3719 2975
rect 3740 2974 3744 2978
rect 3747 2971 3751 2975
rect 3765 2971 3769 2975
rect 3787 2974 3791 2978
rect 3812 2974 3816 2978
rect 3822 2971 3826 2975
rect 3838 2971 3842 2975
rect 3858 2974 3862 2978
rect 3865 2971 3869 2975
rect 3929 2981 3933 2985
rect 3100 2959 3104 2963
rect 3482 2961 3486 2965
rect 3042 2953 3046 2957
rect 3349 2952 3353 2956
rect 3474 2954 3478 2958
rect 3498 2954 3502 2958
rect 3708 2954 3712 2958
rect 3055 2945 3059 2949
rect 3357 2945 3361 2949
rect 3498 2945 3502 2949
rect 3742 2955 3746 2959
rect 3762 2952 3766 2956
rect 3781 2956 3785 2960
rect 3883 2967 3887 2971
rect 3898 2967 3902 2971
rect 3800 2955 3804 2959
rect 3819 2955 3823 2959
rect 3832 2954 3836 2958
rect 3854 2955 3858 2959
rect 3862 2954 3866 2958
rect 3874 2954 3878 2958
rect 3715 2941 3719 2945
rect 3747 2941 3751 2945
rect 3765 2941 3769 2945
rect 3822 2941 3826 2945
rect 3837 2941 3841 2945
rect 3865 2941 3869 2945
rect 3364 2937 3368 2941
rect 3431 2937 3435 2941
rect 3467 2937 3471 2941
rect 3683 2937 3689 2941
rect 3729 2937 3733 2941
rect 3772 2936 3776 2940
rect 3794 2937 3801 2941
rect 3844 2936 3848 2940
rect 3623 2930 3629 2934
rect 2690 2922 2696 2926
rect 2770 2922 2774 2926
rect 2784 2922 2788 2926
rect 2802 2922 2806 2926
rect 2820 2922 2824 2926
rect 2843 2922 2847 2926
rect 2877 2922 2881 2926
rect 2892 2922 2896 2926
rect 2920 2922 2924 2926
rect 2441 2912 2445 2916
rect 2404 2906 2408 2912
rect 2420 2906 2424 2912
rect 2457 2906 2461 2912
rect 2465 2908 2469 2912
rect 2499 2912 2503 2916
rect 2702 2915 2708 2919
rect 2784 2915 2788 2919
rect 2843 2915 2847 2919
rect 2868 2915 2872 2919
rect 2899 2915 2903 2919
rect 2478 2906 2482 2912
rect 2515 2906 2519 2912
rect 2784 2907 2788 2911
rect 2827 2908 2831 2912
rect 2849 2907 2856 2911
rect 2899 2908 2903 2912
rect 2537 2903 2541 2907
rect 2770 2903 2774 2907
rect 2802 2903 2806 2907
rect 2820 2903 2824 2907
rect 2877 2903 2881 2907
rect 2892 2903 2896 2907
rect 2920 2903 2924 2907
rect 2404 2893 2408 2897
rect 2420 2893 2424 2897
rect 2465 2899 2469 2903
rect 2441 2893 2445 2899
rect 2457 2893 2461 2897
rect 2478 2893 2482 2897
rect 2499 2893 2503 2899
rect 2515 2893 2519 2897
rect 2765 2891 2769 2895
rect 2421 2880 2425 2884
rect 2465 2880 2469 2884
rect 2485 2880 2489 2884
rect 2522 2882 2526 2886
rect 2797 2889 2801 2893
rect 2817 2892 2821 2896
rect 2836 2888 2840 2892
rect 2855 2889 2859 2893
rect 2874 2889 2878 2893
rect 2887 2890 2891 2894
rect 2984 2905 2988 2909
rect 3364 2923 3368 2927
rect 3417 2923 3421 2927
rect 3467 2923 3471 2927
rect 3647 2929 3653 2933
rect 3729 2929 3733 2933
rect 3788 2929 3792 2933
rect 3813 2929 3817 2933
rect 3844 2929 3848 2933
rect 3937 2959 3941 2967
rect 4010 2981 4014 2985
rect 3964 2967 3968 2971
rect 3979 2967 3983 2971
rect 3960 2959 3964 2963
rect 3906 2953 3910 2957
rect 3919 2945 3923 2949
rect 4018 2959 4022 2967
rect 4045 2959 4049 2963
rect 3987 2953 3991 2957
rect 4000 2945 4004 2949
rect 3635 2922 3641 2926
rect 3715 2922 3719 2926
rect 3729 2922 3733 2926
rect 3747 2922 3751 2926
rect 3765 2922 3769 2926
rect 3788 2922 3792 2926
rect 3822 2922 3826 2926
rect 3837 2922 3841 2926
rect 3865 2922 3869 2926
rect 3386 2912 3390 2916
rect 3065 2905 3069 2909
rect 3349 2906 3353 2912
rect 3365 2906 3369 2912
rect 3402 2906 3406 2912
rect 3410 2908 3414 2912
rect 3444 2912 3448 2916
rect 3647 2915 3653 2919
rect 3729 2915 3733 2919
rect 3788 2915 3792 2919
rect 3813 2915 3817 2919
rect 3844 2915 3848 2919
rect 3423 2906 3427 2912
rect 3460 2906 3464 2912
rect 3729 2907 3733 2911
rect 3772 2908 3776 2912
rect 3794 2907 3801 2911
rect 3844 2908 3848 2912
rect 3482 2903 3486 2907
rect 3715 2903 3719 2907
rect 3747 2903 3751 2907
rect 3765 2903 3769 2907
rect 3822 2903 3826 2907
rect 3837 2903 3841 2907
rect 3865 2903 3869 2907
rect 2909 2889 2913 2893
rect 2917 2890 2921 2894
rect 2929 2890 2933 2894
rect 2964 2890 2968 2894
rect 2992 2889 2996 2893
rect 3044 2890 3048 2894
rect 3349 2893 3353 2897
rect 3365 2893 3369 2897
rect 3410 2899 3414 2903
rect 3386 2893 3390 2899
rect 3402 2893 3406 2897
rect 3073 2889 3077 2893
rect 3423 2893 3427 2897
rect 3444 2893 3448 2899
rect 3460 2893 3464 2897
rect 3710 2891 3714 2895
rect 2690 2873 2696 2877
rect 2770 2873 2774 2877
rect 2795 2870 2799 2874
rect 2802 2873 2806 2877
rect 2820 2873 2824 2877
rect 2842 2870 2846 2874
rect 2867 2870 2871 2874
rect 2877 2873 2881 2877
rect 2893 2873 2897 2877
rect 2913 2870 2917 2874
rect 2920 2873 2924 2877
rect 2421 2866 2425 2870
rect 2471 2866 2475 2870
rect 2522 2866 2526 2870
rect 2726 2866 2732 2870
rect 2780 2863 2784 2867
rect 2796 2863 2800 2867
rect 2827 2863 2831 2867
rect 2849 2863 2853 2867
rect 2914 2863 2918 2867
rect 2974 2869 2978 2873
rect 3366 2880 3370 2884
rect 3410 2880 3414 2884
rect 3430 2880 3434 2884
rect 3467 2882 3471 2886
rect 3742 2889 3746 2893
rect 3762 2892 3766 2896
rect 3781 2888 3785 2892
rect 3800 2889 3804 2893
rect 3819 2889 3823 2893
rect 3832 2890 3836 2894
rect 3929 2905 3933 2909
rect 4010 2905 4014 2909
rect 3854 2889 3858 2893
rect 3862 2890 3866 2894
rect 3874 2890 3878 2894
rect 3909 2890 3913 2894
rect 3937 2889 3941 2893
rect 3989 2890 3993 2894
rect 4018 2889 4022 2893
rect 3635 2873 3641 2877
rect 3715 2873 3719 2877
rect 3055 2869 3059 2873
rect 3740 2870 3744 2874
rect 3747 2873 3751 2877
rect 3765 2873 3769 2877
rect 3787 2870 3791 2874
rect 3812 2870 3816 2874
rect 3822 2873 3826 2877
rect 3838 2873 3842 2877
rect 3858 2870 3862 2874
rect 3865 2873 3869 2877
rect 3366 2866 3370 2870
rect 3416 2866 3420 2870
rect 3467 2866 3471 2870
rect 3671 2866 3677 2870
rect 3725 2863 3729 2867
rect 3741 2863 3745 2867
rect 3772 2863 3776 2867
rect 3794 2863 3798 2867
rect 3859 2863 3863 2867
rect 3919 2869 3923 2873
rect 4000 2869 4004 2873
rect 2678 2856 2684 2860
rect 2769 2856 2773 2860
rect 2803 2856 2807 2860
rect 2820 2856 2824 2860
rect 2876 2856 2880 2860
rect 2893 2856 2897 2860
rect 2921 2856 2925 2860
rect 3623 2856 3629 2860
rect 3714 2856 3718 2860
rect 3748 2856 3752 2860
rect 3765 2856 3769 2860
rect 3821 2856 3825 2860
rect 3838 2856 3842 2860
rect 3866 2856 3870 2860
rect 2714 2849 2720 2853
rect 2780 2849 2784 2853
rect 2796 2849 2800 2853
rect 2827 2849 2831 2853
rect 2849 2849 2853 2853
rect 2914 2849 2918 2853
rect 2984 2849 2988 2853
rect 2770 2839 2774 2843
rect 2795 2842 2799 2846
rect 2802 2839 2806 2843
rect 2820 2839 2824 2843
rect 2842 2842 2846 2846
rect 2867 2842 2871 2846
rect 2877 2839 2881 2843
rect 2893 2839 2897 2843
rect 2913 2842 2917 2846
rect 2920 2839 2924 2843
rect 2764 2822 2768 2826
rect 2797 2823 2801 2827
rect 2817 2820 2821 2824
rect 2836 2824 2840 2828
rect 2855 2823 2859 2827
rect 2874 2823 2878 2827
rect 2887 2822 2891 2826
rect 2909 2823 2913 2827
rect 2917 2822 2921 2826
rect 2929 2822 2933 2826
rect 2992 2827 2996 2835
rect 3089 2849 3093 2853
rect 3043 2835 3047 2839
rect 3058 2835 3062 2839
rect 3659 2849 3665 2853
rect 3725 2849 3729 2853
rect 3741 2849 3745 2853
rect 3772 2849 3776 2853
rect 3794 2849 3798 2853
rect 3859 2849 3863 2853
rect 3929 2849 3933 2853
rect 2961 2821 2965 2825
rect 3015 2826 3019 2830
rect 2770 2809 2774 2813
rect 2802 2809 2806 2813
rect 2820 2809 2824 2813
rect 2877 2809 2881 2813
rect 2892 2809 2896 2813
rect 2920 2809 2924 2813
rect 2784 2805 2788 2809
rect 2827 2804 2831 2808
rect 2849 2805 2856 2809
rect 2899 2804 2903 2808
rect 2702 2797 2708 2801
rect 2784 2797 2788 2801
rect 2843 2797 2847 2801
rect 2868 2797 2872 2801
rect 2899 2797 2903 2801
rect 2974 2813 2978 2817
rect 3097 2827 3101 2835
rect 3715 2839 3719 2843
rect 3740 2842 3744 2846
rect 3747 2839 3751 2843
rect 3765 2839 3769 2843
rect 3787 2842 3791 2846
rect 3812 2842 3816 2846
rect 3822 2839 3826 2843
rect 3838 2839 3842 2843
rect 3858 2842 3862 2846
rect 3865 2839 3869 2843
rect 3118 2827 3122 2831
rect 3066 2821 3070 2825
rect 3709 2822 3713 2826
rect 3079 2813 3083 2817
rect 3742 2823 3746 2827
rect 3762 2820 3766 2824
rect 3781 2824 3785 2828
rect 3800 2823 3804 2827
rect 3819 2823 3823 2827
rect 3832 2822 3836 2826
rect 3854 2823 3858 2827
rect 3862 2822 3866 2826
rect 3874 2822 3878 2826
rect 3937 2827 3941 2835
rect 4034 2849 4038 2853
rect 3988 2835 3992 2839
rect 4003 2835 4007 2839
rect 3906 2821 3910 2825
rect 3960 2826 3964 2830
rect 3715 2809 3719 2813
rect 3747 2809 3751 2813
rect 3765 2809 3769 2813
rect 3822 2809 3826 2813
rect 3837 2809 3841 2813
rect 3865 2809 3869 2813
rect 3729 2805 3733 2809
rect 3772 2804 3776 2808
rect 3794 2805 3801 2809
rect 3844 2804 3848 2808
rect 3647 2797 3653 2801
rect 3729 2797 3733 2801
rect 3788 2797 3792 2801
rect 3813 2797 3817 2801
rect 3844 2797 3848 2801
rect 3919 2813 3923 2817
rect 4042 2827 4046 2835
rect 4063 2827 4067 2831
rect 4011 2821 4015 2825
rect 4024 2813 4028 2817
rect 2690 2790 2696 2794
rect 2770 2790 2774 2794
rect 2784 2790 2788 2794
rect 2802 2790 2806 2794
rect 2820 2790 2824 2794
rect 2843 2790 2847 2794
rect 2877 2790 2881 2794
rect 2892 2790 2896 2794
rect 2920 2790 2924 2794
rect 3635 2790 3641 2794
rect 3715 2790 3719 2794
rect 3729 2790 3733 2794
rect 3747 2790 3751 2794
rect 3765 2790 3769 2794
rect 3788 2790 3792 2794
rect 3822 2790 3826 2794
rect 3837 2790 3841 2794
rect 3865 2790 3869 2794
rect 2702 2783 2708 2787
rect 2784 2783 2788 2787
rect 2843 2783 2847 2787
rect 2868 2783 2872 2787
rect 2899 2783 2903 2787
rect 2784 2775 2788 2779
rect 2827 2776 2831 2780
rect 2849 2775 2856 2779
rect 2899 2776 2903 2780
rect 2770 2771 2774 2775
rect 2802 2771 2806 2775
rect 2820 2771 2824 2775
rect 2877 2771 2881 2775
rect 2892 2771 2896 2775
rect 2920 2771 2924 2775
rect 2984 2774 2988 2778
rect 3647 2783 3653 2787
rect 3729 2783 3733 2787
rect 3788 2783 3792 2787
rect 3813 2783 3817 2787
rect 3844 2783 3848 2787
rect 3089 2774 3093 2778
rect 3729 2775 3733 2779
rect 3772 2776 3776 2780
rect 3794 2775 3801 2779
rect 3844 2776 3848 2780
rect 3715 2771 3719 2775
rect 3747 2771 3751 2775
rect 3765 2771 3769 2775
rect 3822 2771 3826 2775
rect 3837 2771 3841 2775
rect 3865 2771 3869 2775
rect 3929 2774 3933 2778
rect 4034 2774 4038 2778
rect 2765 2759 2769 2763
rect 2797 2757 2801 2761
rect 2817 2760 2821 2764
rect 2836 2756 2840 2760
rect 2855 2757 2859 2761
rect 2874 2757 2878 2761
rect 2887 2758 2891 2762
rect 2909 2757 2913 2761
rect 2917 2758 2921 2762
rect 2929 2758 2933 2762
rect 2963 2759 2967 2763
rect 2992 2758 2996 2762
rect 3069 2759 3073 2763
rect 3097 2758 3101 2762
rect 3710 2759 3714 2763
rect 2770 2741 2774 2745
rect 2795 2738 2799 2742
rect 2802 2741 2806 2745
rect 2820 2741 2824 2745
rect 2842 2738 2846 2742
rect 2867 2738 2871 2742
rect 2877 2741 2881 2745
rect 2893 2741 2897 2745
rect 2913 2738 2917 2742
rect 2920 2741 2924 2745
rect 2714 2731 2720 2735
rect 2796 2731 2800 2735
rect 2827 2731 2831 2735
rect 2849 2731 2853 2735
rect 2914 2731 2918 2735
rect 2974 2738 2978 2742
rect 3742 2757 3746 2761
rect 3762 2760 3766 2764
rect 3781 2756 3785 2760
rect 3800 2757 3804 2761
rect 3819 2757 3823 2761
rect 3832 2758 3836 2762
rect 3854 2757 3858 2761
rect 3862 2758 3866 2762
rect 3874 2758 3878 2762
rect 3908 2759 3912 2763
rect 3937 2758 3941 2762
rect 4014 2759 4018 2763
rect 4042 2758 4046 2762
rect 3079 2738 3083 2742
rect 3715 2741 3719 2745
rect 3740 2738 3744 2742
rect 3747 2741 3751 2745
rect 3765 2741 3769 2745
rect 3787 2738 3791 2742
rect 3812 2738 3816 2742
rect 3822 2741 3826 2745
rect 3838 2741 3842 2745
rect 3858 2738 3862 2742
rect 3865 2741 3869 2745
rect 3659 2731 3665 2735
rect 3741 2731 3745 2735
rect 3772 2731 3776 2735
rect 3794 2731 3798 2735
rect 3859 2731 3863 2735
rect 3919 2738 3923 2742
rect 4024 2738 4028 2742
rect 2678 2724 2684 2728
rect 2769 2724 2773 2728
rect 2803 2724 2807 2728
rect 2820 2724 2824 2728
rect 2876 2724 2880 2728
rect 2893 2724 2897 2728
rect 2921 2724 2925 2728
rect 3623 2724 3629 2728
rect 3714 2724 3718 2728
rect 3748 2724 3752 2728
rect 3765 2724 3769 2728
rect 3821 2724 3825 2728
rect 3838 2724 3842 2728
rect 3866 2724 3870 2728
rect 2714 2717 2720 2721
rect 2796 2717 2800 2721
rect 2827 2717 2831 2721
rect 2849 2717 2853 2721
rect 2914 2717 2918 2721
rect 2984 2717 2988 2721
rect 2770 2707 2774 2711
rect 2795 2710 2799 2714
rect 2802 2707 2806 2711
rect 2820 2707 2824 2711
rect 2842 2710 2846 2714
rect 2867 2710 2871 2714
rect 2877 2707 2881 2711
rect 2893 2707 2897 2711
rect 2913 2710 2917 2714
rect 2920 2707 2924 2711
rect 2764 2690 2768 2694
rect 2797 2691 2801 2695
rect 2817 2688 2821 2692
rect 2836 2692 2840 2696
rect 2855 2691 2859 2695
rect 2874 2691 2878 2695
rect 2887 2690 2891 2694
rect 2909 2691 2913 2695
rect 2917 2690 2921 2694
rect 2929 2690 2933 2694
rect 2992 2695 2996 2703
rect 3065 2717 3069 2721
rect 3019 2703 3023 2707
rect 3034 2703 3038 2707
rect 3015 2695 3019 2699
rect 2961 2689 2965 2693
rect 2770 2677 2774 2681
rect 2802 2677 2806 2681
rect 2820 2677 2824 2681
rect 2877 2677 2881 2681
rect 2892 2677 2896 2681
rect 2920 2677 2924 2681
rect 2784 2673 2788 2677
rect 2827 2672 2831 2676
rect 2849 2673 2856 2677
rect 2899 2672 2903 2676
rect 2702 2665 2708 2669
rect 2784 2665 2788 2669
rect 2843 2665 2847 2669
rect 2868 2665 2872 2669
rect 2899 2665 2903 2669
rect 2974 2681 2978 2685
rect 3073 2695 3077 2703
rect 3155 2717 3159 2721
rect 3109 2703 3113 2707
rect 3124 2703 3128 2707
rect 3659 2717 3665 2721
rect 3741 2717 3745 2721
rect 3772 2717 3776 2721
rect 3794 2717 3798 2721
rect 3859 2717 3863 2721
rect 3929 2717 3933 2721
rect 3097 2695 3101 2699
rect 3042 2689 3046 2693
rect 3131 2697 3135 2701
rect 3163 2695 3167 2703
rect 3715 2707 3719 2711
rect 3740 2710 3744 2714
rect 3747 2707 3751 2711
rect 3765 2707 3769 2711
rect 3787 2710 3791 2714
rect 3812 2710 3816 2714
rect 3822 2707 3826 2711
rect 3838 2707 3842 2711
rect 3858 2710 3862 2714
rect 3865 2707 3869 2711
rect 3055 2681 3059 2685
rect 3198 2694 3202 2698
rect 3709 2690 3713 2694
rect 3145 2681 3149 2685
rect 3742 2691 3746 2695
rect 3762 2688 3766 2692
rect 3781 2692 3785 2696
rect 3800 2691 3804 2695
rect 3819 2691 3823 2695
rect 3832 2690 3836 2694
rect 3854 2691 3858 2695
rect 3862 2690 3866 2694
rect 3874 2690 3878 2694
rect 3937 2695 3941 2703
rect 4010 2717 4014 2721
rect 3964 2703 3968 2707
rect 3979 2703 3983 2707
rect 3960 2695 3964 2699
rect 3906 2689 3910 2693
rect 3715 2677 3719 2681
rect 3747 2677 3751 2681
rect 3765 2677 3769 2681
rect 3822 2677 3826 2681
rect 3837 2677 3841 2681
rect 3865 2677 3869 2681
rect 3729 2673 3733 2677
rect 3772 2672 3776 2676
rect 3794 2673 3801 2677
rect 3844 2672 3848 2676
rect 3647 2665 3653 2669
rect 3729 2665 3733 2669
rect 3788 2665 3792 2669
rect 3813 2665 3817 2669
rect 3844 2665 3848 2669
rect 3919 2681 3923 2685
rect 4018 2695 4022 2703
rect 4100 2717 4104 2721
rect 4054 2703 4058 2707
rect 4069 2703 4073 2707
rect 4042 2695 4046 2699
rect 3987 2689 3991 2693
rect 4076 2697 4080 2701
rect 4108 2695 4112 2703
rect 4000 2681 4004 2685
rect 4143 2694 4147 2698
rect 4291 2694 4300 2699
rect 4090 2681 4094 2685
rect 2690 2658 2696 2662
rect 2770 2658 2774 2662
rect 2784 2658 2788 2662
rect 2802 2658 2806 2662
rect 2820 2658 2824 2662
rect 2843 2658 2847 2662
rect 2877 2658 2881 2662
rect 2892 2658 2896 2662
rect 2920 2658 2924 2662
rect 3635 2658 3641 2662
rect 3715 2658 3719 2662
rect 3729 2658 3733 2662
rect 3747 2658 3751 2662
rect 3765 2658 3769 2662
rect 3788 2658 3792 2662
rect 3822 2658 3826 2662
rect 3837 2658 3841 2662
rect 3865 2658 3869 2662
rect 2702 2651 2708 2655
rect 2784 2651 2788 2655
rect 2843 2651 2847 2655
rect 2868 2651 2872 2655
rect 2899 2651 2903 2655
rect 2784 2643 2788 2647
rect 2827 2644 2831 2648
rect 2849 2643 2856 2647
rect 2899 2644 2903 2648
rect 2770 2639 2774 2643
rect 2802 2639 2806 2643
rect 2820 2639 2824 2643
rect 2877 2639 2881 2643
rect 2892 2639 2896 2643
rect 2920 2639 2924 2643
rect 2765 2627 2769 2631
rect 2797 2625 2801 2629
rect 2817 2628 2821 2632
rect 2836 2624 2840 2628
rect 2855 2625 2859 2629
rect 2874 2625 2878 2629
rect 2887 2626 2891 2630
rect 2984 2639 2988 2643
rect 3065 2639 3069 2643
rect 3647 2651 3653 2655
rect 3729 2651 3733 2655
rect 3788 2651 3792 2655
rect 3813 2651 3817 2655
rect 3844 2651 3848 2655
rect 3729 2643 3733 2647
rect 3772 2644 3776 2648
rect 3794 2643 3801 2647
rect 3844 2644 3848 2648
rect 3155 2639 3159 2643
rect 3715 2639 3719 2643
rect 3747 2639 3751 2643
rect 3765 2639 3769 2643
rect 3822 2639 3826 2643
rect 3837 2639 3841 2643
rect 3865 2639 3869 2643
rect 2909 2625 2913 2629
rect 2917 2626 2921 2630
rect 2929 2626 2933 2630
rect 2964 2624 2968 2628
rect 2992 2623 2996 2627
rect 3044 2624 3048 2628
rect 3073 2623 3077 2627
rect 3128 2624 3132 2628
rect 3710 2627 3714 2631
rect 3163 2623 3167 2627
rect 2770 2609 2774 2613
rect 2795 2606 2799 2610
rect 2802 2609 2806 2613
rect 2820 2609 2824 2613
rect 2842 2606 2846 2610
rect 2867 2606 2871 2610
rect 2877 2609 2881 2613
rect 2893 2609 2897 2613
rect 2913 2606 2917 2610
rect 2920 2609 2924 2613
rect 3742 2625 3746 2629
rect 3762 2628 3766 2632
rect 3781 2624 3785 2628
rect 3800 2625 3804 2629
rect 3819 2625 3823 2629
rect 3832 2626 3836 2630
rect 3929 2639 3933 2643
rect 4010 2639 4014 2643
rect 4291 2657 4300 2670
rect 4100 2639 4104 2643
rect 3854 2625 3858 2629
rect 3862 2626 3866 2630
rect 3874 2626 3878 2630
rect 3909 2624 3913 2628
rect 3937 2623 3941 2627
rect 3989 2624 3993 2628
rect 4018 2623 4022 2627
rect 4073 2624 4077 2628
rect 4108 2623 4112 2627
rect 2714 2599 2720 2603
rect 2796 2599 2800 2603
rect 2827 2599 2831 2603
rect 2849 2599 2853 2603
rect 2914 2599 2918 2603
rect 2974 2603 2978 2607
rect 3055 2603 3059 2607
rect 3715 2609 3719 2613
rect 3145 2603 3149 2607
rect 3740 2606 3744 2610
rect 3747 2609 3751 2613
rect 3765 2609 3769 2613
rect 3787 2606 3791 2610
rect 3812 2606 3816 2610
rect 3822 2609 3826 2613
rect 3838 2609 3842 2613
rect 3858 2606 3862 2610
rect 3865 2609 3869 2613
rect 3659 2599 3665 2603
rect 3741 2599 3745 2603
rect 3772 2599 3776 2603
rect 3794 2599 3798 2603
rect 3859 2599 3863 2603
rect 3919 2603 3923 2607
rect 4000 2603 4004 2607
rect 4090 2603 4094 2607
rect 2678 2592 2684 2596
rect 2769 2592 2773 2596
rect 2803 2592 2807 2596
rect 2820 2592 2824 2596
rect 2876 2592 2880 2596
rect 2893 2592 2897 2596
rect 2921 2592 2925 2596
rect 3623 2592 3629 2596
rect 3714 2592 3718 2596
rect 3748 2592 3752 2596
rect 3765 2592 3769 2596
rect 3821 2592 3825 2596
rect 3838 2592 3842 2596
rect 3866 2592 3870 2596
rect 2714 2585 2720 2589
rect 2796 2585 2800 2589
rect 2827 2585 2831 2589
rect 2849 2585 2853 2589
rect 2914 2585 2918 2589
rect 2984 2585 2988 2589
rect 2770 2575 2774 2579
rect 2795 2578 2799 2582
rect 2802 2575 2806 2579
rect 2820 2575 2824 2579
rect 2842 2578 2846 2582
rect 2867 2578 2871 2582
rect 2877 2575 2881 2579
rect 2893 2575 2897 2579
rect 2913 2578 2917 2582
rect 2920 2575 2924 2579
rect 2764 2558 2768 2562
rect 2797 2559 2801 2563
rect 2817 2556 2821 2560
rect 2836 2560 2840 2564
rect 3659 2585 3665 2589
rect 3741 2585 3745 2589
rect 3772 2585 3776 2589
rect 3794 2585 3798 2589
rect 3859 2585 3863 2589
rect 3929 2585 3933 2589
rect 2855 2559 2859 2563
rect 2874 2559 2878 2563
rect 2887 2558 2891 2562
rect 2909 2559 2913 2563
rect 2917 2558 2921 2562
rect 2929 2558 2933 2562
rect 2992 2563 2996 2571
rect 3715 2575 3719 2579
rect 3740 2578 3744 2582
rect 3747 2575 3751 2579
rect 3765 2575 3769 2579
rect 3787 2578 3791 2582
rect 3812 2578 3816 2582
rect 3822 2575 3826 2579
rect 3838 2575 3842 2579
rect 3858 2578 3862 2582
rect 3865 2575 3869 2579
rect 2961 2557 2965 2561
rect 3015 2562 3019 2566
rect 3709 2558 3713 2562
rect 2770 2545 2774 2549
rect 2802 2545 2806 2549
rect 2820 2545 2824 2549
rect 2877 2545 2881 2549
rect 2892 2545 2896 2549
rect 2920 2545 2924 2549
rect 2784 2541 2788 2545
rect 2287 2537 2291 2541
rect 2323 2537 2327 2541
rect 2390 2537 2394 2541
rect 2419 2537 2423 2541
rect 2455 2537 2459 2541
rect 2522 2537 2526 2541
rect 2551 2537 2555 2541
rect 2587 2537 2591 2541
rect 2654 2537 2658 2541
rect 2738 2537 2744 2541
rect 2827 2540 2831 2544
rect 2849 2541 2856 2545
rect 2899 2540 2903 2544
rect 2678 2530 2684 2534
rect 2784 2533 2788 2537
rect 2793 2533 2797 2537
rect 2843 2533 2847 2537
rect 2868 2533 2872 2537
rect 2899 2533 2903 2537
rect 2974 2549 2978 2553
rect 3742 2559 3746 2563
rect 3762 2556 3766 2560
rect 3781 2560 3785 2564
rect 3800 2559 3804 2563
rect 3819 2559 3823 2563
rect 3832 2558 3836 2562
rect 3854 2559 3858 2563
rect 3862 2558 3866 2562
rect 3874 2558 3878 2562
rect 3937 2563 3941 2571
rect 3906 2557 3910 2561
rect 3960 2562 3964 2566
rect 3715 2545 3719 2549
rect 3747 2545 3751 2549
rect 3765 2545 3769 2549
rect 3822 2545 3826 2549
rect 3837 2545 3841 2549
rect 3865 2545 3869 2549
rect 3729 2541 3733 2545
rect 3232 2537 3236 2541
rect 3268 2537 3272 2541
rect 3335 2537 3339 2541
rect 3364 2537 3368 2541
rect 3400 2537 3404 2541
rect 3467 2537 3471 2541
rect 3496 2537 3500 2541
rect 3532 2537 3536 2541
rect 3599 2537 3603 2541
rect 3683 2537 3689 2541
rect 3772 2540 3776 2544
rect 3794 2541 3801 2545
rect 3844 2540 3848 2544
rect 3623 2530 3629 2534
rect 3729 2533 3733 2537
rect 3738 2533 3742 2537
rect 3788 2533 3792 2537
rect 3813 2533 3817 2537
rect 3844 2533 3848 2537
rect 3919 2549 3923 2553
rect 2287 2523 2291 2527
rect 2337 2523 2341 2527
rect 2390 2523 2394 2527
rect 2419 2523 2423 2527
rect 2469 2523 2473 2527
rect 2522 2523 2526 2527
rect 2551 2523 2555 2527
rect 2601 2523 2605 2527
rect 2654 2523 2658 2527
rect 2690 2526 2696 2530
rect 2770 2526 2774 2530
rect 2784 2526 2788 2530
rect 2802 2526 2806 2530
rect 2820 2526 2824 2530
rect 2843 2526 2847 2530
rect 2877 2526 2881 2530
rect 2892 2526 2896 2530
rect 2920 2526 2924 2530
rect 3045 2526 3049 2530
rect 3063 2526 3067 2530
rect 3081 2526 3085 2530
rect 3104 2526 3108 2530
rect 3138 2526 3142 2530
rect 3153 2526 3157 2530
rect 3181 2526 3185 2530
rect 2310 2512 2314 2516
rect 2281 2503 2285 2507
rect 2294 2506 2298 2512
rect 2331 2506 2335 2512
rect 2344 2508 2348 2512
rect 2368 2512 2372 2516
rect 2442 2512 2446 2516
rect 2352 2506 2356 2512
rect 2389 2506 2393 2512
rect 2405 2506 2409 2512
rect 2426 2506 2430 2512
rect 2463 2506 2467 2512
rect 2476 2508 2480 2512
rect 2500 2512 2504 2516
rect 2574 2512 2578 2516
rect 2484 2506 2488 2512
rect 2521 2506 2525 2512
rect 2537 2506 2541 2512
rect 2558 2506 2562 2512
rect 2595 2506 2599 2512
rect 2608 2508 2612 2512
rect 2632 2512 2636 2516
rect 2702 2519 2708 2523
rect 2784 2519 2788 2523
rect 2793 2519 2797 2523
rect 2843 2519 2847 2523
rect 2868 2519 2872 2523
rect 2899 2519 2903 2523
rect 2616 2506 2620 2512
rect 2653 2506 2657 2512
rect 2669 2508 2673 2512
rect 2784 2511 2788 2515
rect 2827 2512 2831 2516
rect 2849 2511 2856 2515
rect 2899 2512 2903 2516
rect 2770 2507 2774 2511
rect 2802 2507 2806 2511
rect 2820 2507 2824 2511
rect 2877 2507 2881 2511
rect 2892 2507 2896 2511
rect 2920 2507 2924 2511
rect 2294 2493 2298 2497
rect 2310 2493 2314 2499
rect 2344 2499 2348 2503
rect 2331 2493 2335 2497
rect 2352 2493 2356 2497
rect 2368 2493 2372 2499
rect 2389 2493 2393 2497
rect 2405 2493 2409 2497
rect 2426 2493 2430 2497
rect 2442 2493 2446 2499
rect 2476 2499 2480 2503
rect 2463 2493 2467 2497
rect 2484 2493 2488 2497
rect 2500 2493 2504 2499
rect 2521 2493 2525 2497
rect 2537 2493 2541 2497
rect 2558 2493 2562 2497
rect 2574 2493 2578 2499
rect 2608 2499 2612 2503
rect 2595 2493 2599 2497
rect 2616 2493 2620 2497
rect 2632 2493 2636 2499
rect 2653 2493 2657 2497
rect 2669 2493 2673 2497
rect 2765 2495 2769 2499
rect 2287 2482 2291 2486
rect 2324 2480 2328 2484
rect 2344 2480 2348 2484
rect 2388 2480 2392 2484
rect 2419 2482 2423 2486
rect 2456 2480 2460 2484
rect 2476 2480 2480 2484
rect 2520 2480 2524 2484
rect 2551 2482 2555 2486
rect 2588 2480 2592 2484
rect 2608 2480 2612 2484
rect 2652 2480 2656 2484
rect 2797 2493 2801 2497
rect 2817 2496 2821 2500
rect 2836 2492 2840 2496
rect 2855 2493 2859 2497
rect 2874 2493 2878 2497
rect 2887 2494 2891 2498
rect 3023 2519 3027 2523
rect 3045 2519 3049 2523
rect 3104 2519 3108 2523
rect 3129 2519 3133 2523
rect 3160 2519 3164 2523
rect 3232 2523 3236 2527
rect 3282 2523 3286 2527
rect 3335 2523 3339 2527
rect 3364 2523 3368 2527
rect 3414 2523 3418 2527
rect 3467 2523 3471 2527
rect 3496 2523 3500 2527
rect 3546 2523 3550 2527
rect 3599 2523 3603 2527
rect 3635 2526 3641 2530
rect 3715 2526 3719 2530
rect 3729 2526 3733 2530
rect 3747 2526 3751 2530
rect 3765 2526 3769 2530
rect 3788 2526 3792 2530
rect 3822 2526 3826 2530
rect 3837 2526 3841 2530
rect 3865 2526 3869 2530
rect 3990 2526 3994 2530
rect 4008 2526 4012 2530
rect 4026 2526 4030 2530
rect 4049 2526 4053 2530
rect 4083 2526 4087 2530
rect 4098 2526 4102 2530
rect 4126 2526 4130 2530
rect 3045 2511 3049 2515
rect 3088 2512 3092 2516
rect 3110 2511 3117 2515
rect 3160 2512 3164 2516
rect 3255 2512 3259 2516
rect 3063 2507 3067 2511
rect 3081 2507 3085 2511
rect 3138 2507 3142 2511
rect 3153 2507 3157 2511
rect 3181 2507 3185 2511
rect 2984 2503 2988 2507
rect 2909 2493 2913 2497
rect 2917 2494 2921 2498
rect 2929 2494 2933 2498
rect 2963 2488 2967 2492
rect 3003 2494 3007 2498
rect 2992 2487 2996 2491
rect 2770 2477 2774 2481
rect 2690 2473 2696 2477
rect 2795 2474 2799 2478
rect 2802 2477 2806 2481
rect 2820 2477 2824 2481
rect 2842 2474 2846 2478
rect 2867 2474 2871 2478
rect 2877 2477 2881 2481
rect 2893 2477 2897 2481
rect 2913 2474 2917 2478
rect 2920 2477 2924 2481
rect 3058 2493 3062 2497
rect 3078 2496 3082 2500
rect 3097 2492 3101 2496
rect 3226 2503 3230 2507
rect 3239 2506 3243 2512
rect 3276 2506 3280 2512
rect 3289 2508 3293 2512
rect 3313 2512 3317 2516
rect 3387 2512 3391 2516
rect 3297 2506 3301 2512
rect 3334 2506 3338 2512
rect 3350 2506 3354 2512
rect 3371 2506 3375 2512
rect 3408 2506 3412 2512
rect 3421 2508 3425 2512
rect 3445 2512 3449 2516
rect 3519 2512 3523 2516
rect 3429 2506 3433 2512
rect 3466 2506 3470 2512
rect 3482 2506 3486 2512
rect 3503 2506 3507 2512
rect 3540 2506 3544 2512
rect 3553 2508 3557 2512
rect 3577 2512 3581 2516
rect 3647 2519 3653 2523
rect 3729 2519 3733 2523
rect 3738 2519 3742 2523
rect 3788 2519 3792 2523
rect 3813 2519 3817 2523
rect 3844 2519 3848 2523
rect 3561 2506 3565 2512
rect 3598 2506 3602 2512
rect 3614 2508 3618 2512
rect 3729 2511 3733 2515
rect 3772 2512 3776 2516
rect 3794 2511 3801 2515
rect 3844 2512 3848 2516
rect 3715 2507 3719 2511
rect 3747 2507 3751 2511
rect 3765 2507 3769 2511
rect 3822 2507 3826 2511
rect 3837 2507 3841 2511
rect 3865 2507 3869 2511
rect 3116 2493 3120 2497
rect 3135 2493 3139 2497
rect 3148 2494 3152 2498
rect 3170 2493 3174 2497
rect 3178 2494 3182 2498
rect 3190 2494 3194 2498
rect 3239 2493 3243 2497
rect 3255 2493 3259 2499
rect 3289 2499 3293 2503
rect 3276 2493 3280 2497
rect 3297 2493 3301 2497
rect 3313 2493 3317 2499
rect 3334 2493 3338 2497
rect 3350 2493 3354 2497
rect 3371 2493 3375 2497
rect 3387 2493 3391 2499
rect 3421 2499 3425 2503
rect 3408 2493 3412 2497
rect 3429 2493 3433 2497
rect 3445 2493 3449 2499
rect 3466 2493 3470 2497
rect 3482 2493 3486 2497
rect 3503 2493 3507 2497
rect 3519 2493 3523 2499
rect 3553 2499 3557 2503
rect 3540 2493 3544 2497
rect 3561 2493 3565 2497
rect 3577 2493 3581 2499
rect 3598 2493 3602 2497
rect 3614 2493 3618 2497
rect 3710 2495 3714 2499
rect 3004 2477 3008 2481
rect 3030 2477 3034 2481
rect 2287 2466 2291 2470
rect 2338 2466 2342 2470
rect 2388 2466 2392 2470
rect 2419 2466 2423 2470
rect 2470 2466 2474 2470
rect 2520 2466 2524 2470
rect 2551 2466 2555 2470
rect 2602 2466 2606 2470
rect 2652 2466 2656 2470
rect 2726 2467 2732 2471
rect 2778 2467 2782 2471
rect 2796 2467 2800 2471
rect 2827 2467 2831 2471
rect 2849 2467 2853 2471
rect 2914 2467 2918 2471
rect 3056 2474 3060 2478
rect 3063 2477 3067 2481
rect 3081 2477 3085 2481
rect 3103 2474 3107 2478
rect 3128 2474 3132 2478
rect 3138 2477 3142 2481
rect 3154 2477 3158 2481
rect 3174 2474 3178 2478
rect 3181 2477 3185 2481
rect 3232 2482 3236 2486
rect 3269 2480 3273 2484
rect 3289 2480 3293 2484
rect 3333 2480 3337 2484
rect 3364 2482 3368 2486
rect 3401 2480 3405 2484
rect 3421 2480 3425 2484
rect 3465 2480 3469 2484
rect 3496 2482 3500 2486
rect 3533 2480 3537 2484
rect 3553 2480 3557 2484
rect 3597 2480 3601 2484
rect 3742 2493 3746 2497
rect 3762 2496 3766 2500
rect 3781 2492 3785 2496
rect 3800 2493 3804 2497
rect 3819 2493 3823 2497
rect 3832 2494 3836 2498
rect 3968 2519 3972 2523
rect 3990 2519 3994 2523
rect 4049 2519 4053 2523
rect 4074 2519 4078 2523
rect 4105 2519 4109 2523
rect 3990 2511 3994 2515
rect 4033 2512 4037 2516
rect 4055 2511 4062 2515
rect 4105 2512 4109 2516
rect 4008 2507 4012 2511
rect 4026 2507 4030 2511
rect 4083 2507 4087 2511
rect 4098 2507 4102 2511
rect 4126 2507 4130 2511
rect 3929 2503 3933 2507
rect 3854 2493 3858 2497
rect 3862 2494 3866 2498
rect 3874 2494 3878 2498
rect 3908 2488 3912 2492
rect 3948 2494 3952 2498
rect 3937 2487 3941 2491
rect 3715 2477 3719 2481
rect 3635 2473 3641 2477
rect 3740 2474 3744 2478
rect 3747 2477 3751 2481
rect 3765 2477 3769 2481
rect 3787 2474 3791 2478
rect 3812 2474 3816 2478
rect 3822 2477 3826 2481
rect 3838 2477 3842 2481
rect 3858 2474 3862 2478
rect 3865 2477 3869 2481
rect 4003 2493 4007 2497
rect 4023 2496 4027 2500
rect 4042 2492 4046 2496
rect 4061 2493 4065 2497
rect 4080 2493 4084 2497
rect 4093 2494 4097 2498
rect 4115 2493 4119 2497
rect 4123 2494 4127 2498
rect 4135 2494 4139 2498
rect 3949 2477 3953 2481
rect 3975 2477 3979 2481
rect 2974 2467 2978 2471
rect 3013 2467 3017 2471
rect 3057 2467 3061 2471
rect 3088 2467 3092 2471
rect 3110 2467 3114 2471
rect 3175 2467 3179 2471
rect 3232 2466 3236 2470
rect 3283 2466 3287 2470
rect 3333 2466 3337 2470
rect 3364 2466 3368 2470
rect 3415 2466 3419 2470
rect 3465 2466 3469 2470
rect 3496 2466 3500 2470
rect 3547 2466 3551 2470
rect 3597 2466 3601 2470
rect 3671 2467 3677 2471
rect 3723 2467 3727 2471
rect 3741 2467 3745 2471
rect 3772 2467 3776 2471
rect 3794 2467 3798 2471
rect 3859 2467 3863 2471
rect 4001 2474 4005 2478
rect 4008 2477 4012 2481
rect 4026 2477 4030 2481
rect 4048 2474 4052 2478
rect 4073 2474 4077 2478
rect 4083 2477 4087 2481
rect 4099 2477 4103 2481
rect 4119 2474 4123 2478
rect 4126 2477 4130 2481
rect 3919 2467 3923 2471
rect 3958 2467 3962 2471
rect 4002 2467 4006 2471
rect 4033 2467 4037 2471
rect 4055 2467 4059 2471
rect 4120 2467 4124 2471
rect 2281 2459 2285 2463
rect 2669 2459 2673 2463
rect 2678 2460 2684 2464
rect 2769 2460 2773 2464
rect 2803 2460 2807 2464
rect 2820 2460 2824 2464
rect 2876 2460 2880 2464
rect 2893 2460 2897 2464
rect 2921 2460 2925 2464
rect 3004 2460 3008 2464
rect 3030 2460 3034 2464
rect 3064 2460 3068 2464
rect 3081 2460 3085 2464
rect 3137 2460 3141 2464
rect 3154 2460 3158 2464
rect 3182 2460 3186 2464
rect 3226 2459 3230 2463
rect 3614 2459 3618 2463
rect 3623 2460 3629 2464
rect 3714 2460 3718 2464
rect 3748 2460 3752 2464
rect 3765 2460 3769 2464
rect 3821 2460 3825 2464
rect 3838 2460 3842 2464
rect 3866 2460 3870 2464
rect 3949 2460 3953 2464
rect 3975 2460 3979 2464
rect 4009 2460 4013 2464
rect 4026 2460 4030 2464
rect 4082 2460 4086 2464
rect 4099 2460 4103 2464
rect 4127 2460 4131 2464
rect 2404 2452 2409 2456
rect 2537 2452 2541 2456
rect 2714 2453 2720 2457
rect 2778 2453 2782 2457
rect 3012 2453 3016 2457
rect 3198 2454 3202 2458
rect 3210 2454 3214 2458
rect 3349 2452 3354 2456
rect 3482 2452 3486 2456
rect 3659 2453 3665 2457
rect 3723 2453 3727 2457
rect 3957 2453 3961 2457
rect 4143 2454 4147 2458
rect 4155 2454 4159 2458
rect 2412 2445 2416 2449
rect 2702 2445 2708 2449
rect 3022 2446 3026 2450
rect 3187 2446 3191 2450
rect 2396 2441 2400 2445
rect 2428 2441 2432 2445
rect 2750 2439 2756 2443
rect 3357 2445 3361 2449
rect 3647 2445 3653 2449
rect 3967 2446 3971 2450
rect 4132 2446 4136 2450
rect 3341 2441 3345 2445
rect 3373 2441 3377 2445
rect 3695 2439 3701 2443
rect 2396 2432 2400 2436
rect 2428 2432 2432 2436
rect 3341 2432 3345 2436
rect 3373 2432 3377 2436
rect 2412 2425 2416 2429
rect 2669 2425 2673 2429
rect 2738 2425 2744 2429
rect 3070 2425 3074 2429
rect 3106 2425 3110 2429
rect 3173 2425 3177 2429
rect 3357 2425 3361 2429
rect 3614 2425 3618 2429
rect 3683 2425 3689 2429
rect 4015 2425 4019 2429
rect 4051 2425 4055 2429
rect 4118 2425 4122 2429
rect 2669 2417 2673 2421
rect 2678 2418 2684 2422
rect 3056 2418 3060 2422
rect 2396 2413 2400 2417
rect 2428 2413 2432 2417
rect 2412 2409 2416 2413
rect 3070 2411 3074 2415
rect 3120 2411 3124 2415
rect 3173 2411 3177 2415
rect 3614 2417 3618 2421
rect 3623 2418 3629 2422
rect 4001 2418 4005 2422
rect 3341 2413 3345 2417
rect 3373 2413 3377 2417
rect 3357 2409 3361 2413
rect 4015 2411 4019 2415
rect 4065 2411 4069 2415
rect 4118 2411 4122 2415
rect 2404 2402 2409 2406
rect 2538 2402 2542 2406
rect 3093 2400 3097 2404
rect 2287 2395 2291 2399
rect 2323 2395 2327 2399
rect 2390 2395 2394 2399
rect 2419 2395 2423 2399
rect 2455 2395 2459 2399
rect 2522 2395 2526 2399
rect 2551 2395 2555 2399
rect 2587 2395 2591 2399
rect 2654 2395 2658 2399
rect 2738 2395 2744 2399
rect 2678 2388 2684 2392
rect 3064 2391 3068 2395
rect 3077 2394 3081 2400
rect 3114 2394 3118 2400
rect 3127 2396 3131 2400
rect 3151 2400 3155 2404
rect 3349 2402 3354 2406
rect 3483 2402 3487 2406
rect 4038 2400 4042 2404
rect 3135 2394 3139 2400
rect 3172 2394 3176 2400
rect 3188 2394 3192 2400
rect 3232 2395 3236 2399
rect 3268 2395 3272 2399
rect 3335 2395 3339 2399
rect 3364 2395 3368 2399
rect 3400 2395 3404 2399
rect 3467 2395 3471 2399
rect 3496 2395 3500 2399
rect 3532 2395 3536 2399
rect 3599 2395 3603 2399
rect 3683 2395 3689 2399
rect 2287 2381 2291 2385
rect 2337 2381 2341 2385
rect 2390 2381 2394 2385
rect 2419 2381 2423 2385
rect 2469 2381 2473 2385
rect 2522 2381 2526 2385
rect 2551 2381 2555 2385
rect 2601 2381 2605 2385
rect 2654 2381 2658 2385
rect 3077 2381 3081 2385
rect 3093 2381 3097 2387
rect 3127 2387 3131 2391
rect 3114 2381 3118 2385
rect 2310 2370 2314 2374
rect 2281 2361 2285 2365
rect 2294 2364 2298 2370
rect 2331 2364 2335 2370
rect 2344 2366 2348 2370
rect 2368 2370 2372 2374
rect 2442 2370 2446 2374
rect 2352 2364 2356 2370
rect 2389 2364 2393 2370
rect 2405 2364 2409 2370
rect 2426 2364 2430 2370
rect 2463 2364 2467 2370
rect 2476 2366 2480 2370
rect 2500 2370 2504 2374
rect 2574 2370 2578 2374
rect 2484 2364 2488 2370
rect 2521 2364 2525 2370
rect 2537 2364 2541 2370
rect 2558 2364 2562 2370
rect 2595 2364 2599 2370
rect 2608 2366 2612 2370
rect 2632 2370 2636 2374
rect 2616 2364 2620 2370
rect 2653 2364 2657 2370
rect 2669 2366 2673 2370
rect 3135 2381 3139 2385
rect 3151 2381 3155 2387
rect 3623 2388 3629 2392
rect 4009 2391 4013 2395
rect 4022 2394 4026 2400
rect 4059 2394 4063 2400
rect 4072 2396 4076 2400
rect 4096 2400 4100 2404
rect 4080 2394 4084 2400
rect 4117 2394 4121 2400
rect 4133 2394 4137 2400
rect 3172 2381 3176 2385
rect 3188 2381 3192 2385
rect 3232 2381 3236 2385
rect 3282 2381 3286 2385
rect 3335 2381 3339 2385
rect 3364 2381 3368 2385
rect 3414 2381 3418 2385
rect 3467 2381 3471 2385
rect 3496 2381 3500 2385
rect 3546 2381 3550 2385
rect 3599 2381 3603 2385
rect 4022 2381 4026 2385
rect 4038 2381 4042 2387
rect 4072 2387 4076 2391
rect 4059 2381 4063 2385
rect 3070 2370 3074 2374
rect 3107 2368 3111 2372
rect 3127 2368 3131 2372
rect 3171 2368 3175 2372
rect 3255 2370 3259 2374
rect 2294 2351 2298 2355
rect 2310 2351 2314 2357
rect 2344 2357 2348 2361
rect 2331 2351 2335 2355
rect 2352 2351 2356 2355
rect 2368 2351 2372 2357
rect 2389 2351 2393 2355
rect 2405 2351 2409 2355
rect 2426 2351 2430 2355
rect 2442 2351 2446 2357
rect 2476 2357 2480 2361
rect 2463 2351 2467 2355
rect 2484 2351 2488 2355
rect 2500 2351 2504 2357
rect 2521 2351 2525 2355
rect 2537 2351 2541 2355
rect 2558 2351 2562 2355
rect 2574 2351 2578 2357
rect 2608 2357 2612 2361
rect 2595 2351 2599 2355
rect 2616 2351 2620 2355
rect 2632 2351 2636 2357
rect 2690 2361 2696 2365
rect 3226 2361 3230 2365
rect 3239 2364 3243 2370
rect 3276 2364 3280 2370
rect 3289 2366 3293 2370
rect 3313 2370 3317 2374
rect 3387 2370 3391 2374
rect 3297 2364 3301 2370
rect 3334 2364 3338 2370
rect 3350 2364 3354 2370
rect 3371 2364 3375 2370
rect 3408 2364 3412 2370
rect 3421 2366 3425 2370
rect 3445 2370 3449 2374
rect 3519 2370 3523 2374
rect 3429 2364 3433 2370
rect 3466 2364 3470 2370
rect 3482 2364 3486 2370
rect 3503 2364 3507 2370
rect 3540 2364 3544 2370
rect 3553 2366 3557 2370
rect 3577 2370 3581 2374
rect 3561 2364 3565 2370
rect 3598 2364 3602 2370
rect 3614 2366 3618 2370
rect 4080 2381 4084 2385
rect 4096 2381 4100 2387
rect 4117 2381 4121 2385
rect 4133 2381 4137 2385
rect 4015 2370 4019 2374
rect 4052 2368 4056 2372
rect 4072 2368 4076 2372
rect 4116 2368 4120 2372
rect 2653 2351 2657 2355
rect 2669 2351 2673 2355
rect 2726 2354 2732 2358
rect 3070 2354 3074 2358
rect 3121 2354 3125 2358
rect 3171 2354 3175 2358
rect 3239 2351 3243 2355
rect 3255 2351 3259 2357
rect 3289 2357 3293 2361
rect 3276 2351 3280 2355
rect 2287 2340 2291 2344
rect 2324 2338 2328 2342
rect 2344 2338 2348 2342
rect 2388 2338 2392 2342
rect 2419 2340 2423 2344
rect 2456 2338 2460 2342
rect 2476 2338 2480 2342
rect 2520 2338 2524 2342
rect 2551 2340 2555 2344
rect 2588 2338 2592 2342
rect 2608 2338 2612 2342
rect 2652 2338 2656 2342
rect 3063 2346 3067 2350
rect 3188 2347 3192 2351
rect 3297 2351 3301 2355
rect 3313 2351 3317 2357
rect 3334 2351 3338 2355
rect 3350 2351 3354 2355
rect 3371 2351 3375 2355
rect 3387 2351 3391 2357
rect 3421 2357 3425 2361
rect 3408 2351 3412 2355
rect 3429 2351 3433 2355
rect 3445 2351 3449 2357
rect 3466 2351 3470 2355
rect 3482 2351 3486 2355
rect 3503 2351 3507 2355
rect 3519 2351 3523 2357
rect 3553 2357 3557 2361
rect 3540 2351 3544 2355
rect 3561 2351 3565 2355
rect 3577 2351 3581 2357
rect 3635 2361 3641 2365
rect 3598 2351 3602 2355
rect 3614 2351 3618 2355
rect 3671 2354 3677 2358
rect 4015 2354 4019 2358
rect 4066 2354 4070 2358
rect 4116 2354 4120 2358
rect 2738 2339 2744 2343
rect 3070 2339 3074 2343
rect 3106 2339 3110 2343
rect 3173 2339 3177 2343
rect 2690 2331 2696 2335
rect 3056 2332 3060 2336
rect 3232 2340 3236 2344
rect 3269 2338 3273 2342
rect 3289 2338 3293 2342
rect 3333 2338 3337 2342
rect 3364 2340 3368 2344
rect 3401 2338 3405 2342
rect 3421 2338 3425 2342
rect 3465 2338 3469 2342
rect 3496 2340 3500 2344
rect 3533 2338 3537 2342
rect 3553 2338 3557 2342
rect 3597 2338 3601 2342
rect 4008 2346 4012 2350
rect 4133 2347 4137 2351
rect 3683 2339 3689 2343
rect 4015 2339 4019 2343
rect 4051 2339 4055 2343
rect 4118 2339 4122 2343
rect 2287 2324 2291 2328
rect 2338 2324 2342 2328
rect 2388 2324 2392 2328
rect 2419 2324 2423 2328
rect 2470 2324 2474 2328
rect 2520 2324 2524 2328
rect 2551 2324 2555 2328
rect 2602 2324 2606 2328
rect 2652 2324 2656 2328
rect 2726 2324 2732 2328
rect 3070 2325 3074 2329
rect 3120 2325 3124 2329
rect 3173 2325 3177 2329
rect 3635 2331 3641 2335
rect 4001 2332 4005 2336
rect 3232 2324 3236 2328
rect 3283 2324 3287 2328
rect 3333 2324 3337 2328
rect 3364 2324 3368 2328
rect 3415 2324 3419 2328
rect 3465 2324 3469 2328
rect 3496 2324 3500 2328
rect 3547 2324 3551 2328
rect 3597 2324 3601 2328
rect 3671 2324 3677 2328
rect 4015 2325 4019 2329
rect 4065 2325 4069 2329
rect 4118 2325 4122 2329
rect 2280 2317 2284 2321
rect 2669 2317 2673 2321
rect 3093 2314 3097 2318
rect 2287 2309 2291 2313
rect 2323 2309 2327 2313
rect 2390 2309 2394 2313
rect 2419 2309 2423 2313
rect 2455 2309 2459 2313
rect 2522 2309 2526 2313
rect 2551 2309 2555 2313
rect 2587 2309 2591 2313
rect 2654 2309 2658 2313
rect 2738 2309 2744 2313
rect 2678 2302 2684 2306
rect 3064 2305 3068 2309
rect 3077 2308 3081 2314
rect 3114 2308 3118 2314
rect 3127 2310 3131 2314
rect 3151 2314 3155 2318
rect 3225 2317 3229 2321
rect 3614 2317 3618 2321
rect 4038 2314 4042 2318
rect 3135 2308 3139 2314
rect 3172 2308 3176 2314
rect 3188 2310 3192 2314
rect 3210 2308 3214 2312
rect 3232 2309 3236 2313
rect 3268 2309 3272 2313
rect 3335 2309 3339 2313
rect 3364 2309 3368 2313
rect 3400 2309 3404 2313
rect 3467 2309 3471 2313
rect 3496 2309 3500 2313
rect 3532 2309 3536 2313
rect 3599 2309 3603 2313
rect 3683 2309 3689 2313
rect 2287 2295 2291 2299
rect 2337 2295 2341 2299
rect 2390 2295 2394 2299
rect 2419 2295 2423 2299
rect 2469 2295 2473 2299
rect 2522 2295 2526 2299
rect 2551 2295 2555 2299
rect 2601 2295 2605 2299
rect 2654 2295 2658 2299
rect 3077 2295 3081 2299
rect 3093 2295 3097 2301
rect 3127 2301 3131 2305
rect 3114 2295 3118 2299
rect 2310 2284 2314 2288
rect 2281 2275 2285 2279
rect 2294 2278 2298 2284
rect 2331 2278 2335 2284
rect 2344 2280 2348 2284
rect 2368 2284 2372 2288
rect 2442 2284 2446 2288
rect 2352 2278 2356 2284
rect 2389 2278 2393 2284
rect 2405 2278 2409 2284
rect 2426 2278 2430 2284
rect 2463 2278 2467 2284
rect 2476 2280 2480 2284
rect 2500 2284 2504 2288
rect 2574 2284 2578 2288
rect 2484 2278 2488 2284
rect 2521 2278 2525 2284
rect 2537 2278 2541 2284
rect 2558 2278 2562 2284
rect 2595 2278 2599 2284
rect 2608 2280 2612 2284
rect 2632 2284 2636 2288
rect 2616 2278 2620 2284
rect 2653 2278 2657 2284
rect 2669 2280 2673 2284
rect 3135 2295 3139 2299
rect 3151 2295 3155 2301
rect 3172 2295 3176 2299
rect 3188 2295 3192 2304
rect 3623 2302 3629 2306
rect 4009 2305 4013 2309
rect 4022 2308 4026 2314
rect 4059 2308 4063 2314
rect 4072 2310 4076 2314
rect 4096 2314 4100 2318
rect 4080 2308 4084 2314
rect 4117 2308 4121 2314
rect 4133 2310 4137 2314
rect 4155 2308 4159 2312
rect 3210 2292 3214 2296
rect 3232 2295 3236 2299
rect 3282 2295 3286 2299
rect 3335 2295 3339 2299
rect 3364 2295 3368 2299
rect 3414 2295 3418 2299
rect 3467 2295 3471 2299
rect 3496 2295 3500 2299
rect 3546 2295 3550 2299
rect 3599 2295 3603 2299
rect 4022 2295 4026 2299
rect 4038 2295 4042 2301
rect 4072 2301 4076 2305
rect 4059 2295 4063 2299
rect 3070 2284 3074 2288
rect 3107 2282 3111 2286
rect 3127 2282 3131 2286
rect 3171 2282 3175 2286
rect 3255 2284 3259 2288
rect 2294 2265 2298 2269
rect 2310 2265 2314 2271
rect 2344 2271 2348 2275
rect 2331 2265 2335 2269
rect 2352 2265 2356 2269
rect 2368 2265 2372 2271
rect 2389 2265 2393 2269
rect 2405 2265 2409 2269
rect 2426 2265 2430 2269
rect 2442 2265 2446 2271
rect 2476 2271 2480 2275
rect 2463 2265 2467 2269
rect 2484 2265 2488 2269
rect 2500 2265 2504 2271
rect 2521 2265 2525 2269
rect 2537 2265 2541 2269
rect 2558 2265 2562 2269
rect 2574 2265 2578 2271
rect 2608 2271 2612 2275
rect 2595 2265 2599 2269
rect 2616 2265 2620 2269
rect 2632 2265 2636 2271
rect 2690 2275 2696 2279
rect 3226 2275 3230 2279
rect 3239 2278 3243 2284
rect 3276 2278 3280 2284
rect 3289 2280 3293 2284
rect 3313 2284 3317 2288
rect 3387 2284 3391 2288
rect 3297 2278 3301 2284
rect 3334 2278 3338 2284
rect 3350 2278 3354 2284
rect 3371 2278 3375 2284
rect 3408 2278 3412 2284
rect 3421 2280 3425 2284
rect 3445 2284 3449 2288
rect 3519 2284 3523 2288
rect 3429 2278 3433 2284
rect 3466 2278 3470 2284
rect 3482 2278 3486 2284
rect 3503 2278 3507 2284
rect 3540 2278 3544 2284
rect 3553 2280 3557 2284
rect 3577 2284 3581 2288
rect 3561 2278 3565 2284
rect 3598 2278 3602 2284
rect 3614 2280 3618 2284
rect 4080 2295 4084 2299
rect 4096 2295 4100 2301
rect 4117 2295 4121 2299
rect 4133 2295 4137 2304
rect 4155 2292 4159 2296
rect 4015 2284 4019 2288
rect 4052 2282 4056 2286
rect 4072 2282 4076 2286
rect 4116 2282 4120 2286
rect 2653 2265 2657 2269
rect 2669 2265 2673 2269
rect 2726 2268 2732 2272
rect 3070 2268 3074 2272
rect 3121 2268 3125 2272
rect 3171 2268 3175 2272
rect 3239 2265 3243 2269
rect 3255 2265 3259 2271
rect 3289 2271 3293 2275
rect 3276 2265 3280 2269
rect 3297 2265 3301 2269
rect 3313 2265 3317 2271
rect 3334 2265 3338 2269
rect 3350 2265 3354 2269
rect 3371 2265 3375 2269
rect 3387 2265 3391 2271
rect 3421 2271 3425 2275
rect 3408 2265 3412 2269
rect 3429 2265 3433 2269
rect 3445 2265 3449 2271
rect 3466 2265 3470 2269
rect 3482 2265 3486 2269
rect 3503 2265 3507 2269
rect 3519 2265 3523 2271
rect 3553 2271 3557 2275
rect 3540 2265 3544 2269
rect 3561 2265 3565 2269
rect 3577 2265 3581 2271
rect 3635 2275 3641 2279
rect 3598 2265 3602 2269
rect 3614 2265 3618 2269
rect 3671 2268 3677 2272
rect 4015 2268 4019 2272
rect 4066 2268 4070 2272
rect 4116 2268 4120 2272
rect 2287 2254 2291 2258
rect 2324 2252 2328 2256
rect 2344 2252 2348 2256
rect 2388 2252 2392 2256
rect 2419 2254 2423 2258
rect 2456 2252 2460 2256
rect 2476 2252 2480 2256
rect 2520 2252 2524 2256
rect 2551 2254 2555 2258
rect 2588 2252 2592 2256
rect 2608 2252 2612 2256
rect 2652 2252 2656 2256
rect 3232 2254 3236 2258
rect 3269 2252 3273 2256
rect 3289 2252 3293 2256
rect 3333 2252 3337 2256
rect 3364 2254 3368 2258
rect 3401 2252 3405 2256
rect 3421 2252 3425 2256
rect 3465 2252 3469 2256
rect 3496 2254 3500 2258
rect 3533 2252 3537 2256
rect 3553 2252 3557 2256
rect 3597 2252 3601 2256
rect 2690 2245 2696 2249
rect 3635 2245 3641 2249
rect 2287 2238 2291 2242
rect 2338 2238 2342 2242
rect 2388 2238 2392 2242
rect 2419 2238 2423 2242
rect 2470 2238 2474 2242
rect 2520 2238 2524 2242
rect 2551 2238 2555 2242
rect 2602 2238 2606 2242
rect 2652 2238 2656 2242
rect 2726 2238 2732 2242
rect 3232 2238 3236 2242
rect 3283 2238 3287 2242
rect 3333 2238 3337 2242
rect 3364 2238 3368 2242
rect 3415 2238 3419 2242
rect 3465 2238 3469 2242
rect 3496 2238 3500 2242
rect 3547 2238 3551 2242
rect 3597 2238 3601 2242
rect 3671 2238 3677 2242
rect 2280 2231 2284 2235
rect 2669 2231 2673 2235
rect 3225 2231 3229 2235
rect 3614 2231 3618 2235
rect 2405 2224 2409 2228
rect 2513 2224 2517 2228
rect 2537 2224 2541 2228
rect 3350 2224 3354 2228
rect 3458 2224 3462 2228
rect 3482 2224 3486 2228
rect 2529 2217 2533 2221
rect 2513 2213 2517 2217
rect 2545 2213 2549 2217
rect 3474 2217 3478 2221
rect 3458 2213 3462 2217
rect 3490 2213 3494 2217
rect 2513 2206 2517 2210
rect 2545 2206 2549 2210
rect 3210 2206 3214 2210
rect 3458 2206 3462 2210
rect 3490 2206 3494 2210
rect 4155 2206 4159 2210
rect 2529 2199 2533 2203
rect 2669 2199 2673 2203
rect 3474 2199 3478 2203
rect 3614 2199 3618 2203
rect 2669 2191 2673 2195
rect 3614 2191 3618 2195
rect 2513 2187 2517 2191
rect 2545 2187 2549 2191
rect 2529 2183 2533 2187
rect 3458 2187 3462 2191
rect 3490 2187 3494 2191
rect 3474 2183 3478 2187
rect 2405 2176 2409 2180
rect 2513 2176 2517 2180
rect 2537 2176 2541 2180
rect 3350 2176 3354 2180
rect 3458 2176 3462 2180
rect 3482 2176 3486 2180
rect 2287 2169 2291 2173
rect 2323 2169 2327 2173
rect 2390 2169 2394 2173
rect 2419 2169 2423 2173
rect 2455 2169 2459 2173
rect 2522 2169 2526 2173
rect 2551 2169 2555 2173
rect 2587 2169 2591 2173
rect 2654 2169 2658 2173
rect 2738 2169 2744 2173
rect 3232 2169 3236 2173
rect 3268 2169 3272 2173
rect 3335 2169 3339 2173
rect 3364 2169 3368 2173
rect 3400 2169 3404 2173
rect 3467 2169 3471 2173
rect 3496 2169 3500 2173
rect 3532 2169 3536 2173
rect 3599 2169 3603 2173
rect 3683 2169 3689 2173
rect 2678 2162 2684 2166
rect 3623 2162 3629 2166
rect 2287 2155 2291 2159
rect 2337 2155 2341 2159
rect 2390 2155 2394 2159
rect 2419 2155 2423 2159
rect 2469 2155 2473 2159
rect 2522 2155 2526 2159
rect 2551 2155 2555 2159
rect 2601 2155 2605 2159
rect 2654 2155 2658 2159
rect 3232 2155 3236 2159
rect 3282 2155 3286 2159
rect 3335 2155 3339 2159
rect 3364 2155 3368 2159
rect 3414 2155 3418 2159
rect 3467 2155 3471 2159
rect 3496 2155 3500 2159
rect 3546 2155 3550 2159
rect 3599 2155 3603 2159
rect 2310 2144 2314 2148
rect 2281 2135 2285 2139
rect 2294 2138 2298 2144
rect 2331 2138 2335 2144
rect 2344 2140 2348 2144
rect 2368 2144 2372 2148
rect 2442 2144 2446 2148
rect 2352 2138 2356 2144
rect 2389 2138 2393 2144
rect 2405 2138 2409 2144
rect 2426 2138 2430 2144
rect 2463 2138 2467 2144
rect 2476 2140 2480 2144
rect 2500 2144 2504 2148
rect 2574 2144 2578 2148
rect 2484 2138 2488 2144
rect 2521 2138 2525 2144
rect 2537 2138 2541 2144
rect 2558 2138 2562 2144
rect 2595 2138 2599 2144
rect 2608 2140 2612 2144
rect 2632 2144 2636 2148
rect 3255 2144 3259 2148
rect 2616 2138 2620 2144
rect 2653 2138 2657 2144
rect 2669 2140 2673 2144
rect 2294 2125 2298 2129
rect 2310 2125 2314 2131
rect 2344 2131 2348 2135
rect 2331 2125 2335 2129
rect 2352 2125 2356 2129
rect 2368 2125 2372 2131
rect 2389 2125 2393 2129
rect 2405 2125 2409 2129
rect 2426 2125 2430 2129
rect 2442 2125 2446 2131
rect 2476 2131 2480 2135
rect 2463 2125 2467 2129
rect 2484 2125 2488 2129
rect 2500 2125 2504 2131
rect 2521 2125 2525 2129
rect 2537 2125 2541 2129
rect 2558 2125 2562 2129
rect 2574 2125 2578 2131
rect 2608 2131 2612 2135
rect 2595 2125 2599 2129
rect 2616 2125 2620 2129
rect 2632 2125 2636 2131
rect 3226 2135 3230 2139
rect 3239 2138 3243 2144
rect 3276 2138 3280 2144
rect 3289 2140 3293 2144
rect 3313 2144 3317 2148
rect 3387 2144 3391 2148
rect 3297 2138 3301 2144
rect 3334 2138 3338 2144
rect 3350 2138 3354 2144
rect 3371 2138 3375 2144
rect 3408 2138 3412 2144
rect 3421 2140 3425 2144
rect 3445 2144 3449 2148
rect 3519 2144 3523 2148
rect 3429 2138 3433 2144
rect 3466 2138 3470 2144
rect 3482 2138 3486 2144
rect 3503 2138 3507 2144
rect 3540 2138 3544 2144
rect 3553 2140 3557 2144
rect 3577 2144 3581 2148
rect 3561 2138 3565 2144
rect 3598 2138 3602 2144
rect 3614 2140 3618 2144
rect 2653 2125 2657 2129
rect 2669 2125 2673 2129
rect 3239 2125 3243 2129
rect 3255 2125 3259 2131
rect 3289 2131 3293 2135
rect 3276 2125 3280 2129
rect 3297 2125 3301 2129
rect 3313 2125 3317 2131
rect 3334 2125 3338 2129
rect 3350 2125 3354 2129
rect 3371 2125 3375 2129
rect 3387 2125 3391 2131
rect 3421 2131 3425 2135
rect 3408 2125 3412 2129
rect 3429 2125 3433 2129
rect 3445 2125 3449 2131
rect 3466 2125 3470 2129
rect 3482 2125 3486 2129
rect 3503 2125 3507 2129
rect 3519 2125 3523 2131
rect 3553 2131 3557 2135
rect 3540 2125 3544 2129
rect 3561 2125 3565 2129
rect 3577 2125 3581 2131
rect 3598 2125 3602 2129
rect 3614 2125 3618 2129
rect 2287 2114 2291 2118
rect 2324 2112 2328 2116
rect 2344 2112 2348 2116
rect 2388 2112 2392 2116
rect 2419 2114 2423 2118
rect 2456 2112 2460 2116
rect 2476 2112 2480 2116
rect 2520 2112 2524 2116
rect 2551 2114 2555 2118
rect 2588 2112 2592 2116
rect 2608 2112 2612 2116
rect 2652 2112 2656 2116
rect 3232 2114 3236 2118
rect 3269 2112 3273 2116
rect 3289 2112 3293 2116
rect 3333 2112 3337 2116
rect 3364 2114 3368 2118
rect 3401 2112 3405 2116
rect 3421 2112 3425 2116
rect 3465 2112 3469 2116
rect 3496 2114 3500 2118
rect 3533 2112 3537 2116
rect 3553 2112 3557 2116
rect 3597 2112 3601 2116
rect 2690 2105 2696 2109
rect 3635 2105 3641 2109
rect 2287 2098 2291 2102
rect 2338 2098 2342 2102
rect 2388 2098 2392 2102
rect 2419 2098 2423 2102
rect 2470 2098 2474 2102
rect 2520 2098 2524 2102
rect 2551 2098 2555 2102
rect 2602 2098 2606 2102
rect 2652 2098 2656 2102
rect 2726 2098 2732 2102
rect 3232 2098 3236 2102
rect 3283 2098 3287 2102
rect 3333 2098 3337 2102
rect 3364 2098 3368 2102
rect 3415 2098 3419 2102
rect 3465 2098 3469 2102
rect 3496 2098 3500 2102
rect 3547 2098 3551 2102
rect 3597 2098 3601 2102
rect 3671 2098 3677 2102
<< metal2 >>
rect 2080 4448 2088 4450
rect 2080 4443 2081 4448
rect 2086 4443 2088 4448
rect 2080 4330 2088 4443
rect 2080 4323 2093 4330
rect 2087 4300 2093 4323
rect 2171 4326 2172 4330
rect 2171 4300 2175 4326
rect 2027 4279 2040 4300
rect 2390 4255 2395 4256
rect 2390 3530 2394 4255
rect 2411 4093 2416 4282
rect 2702 4186 2708 4208
rect 2678 4137 2684 4166
rect 2690 4137 2696 4173
rect 2702 4137 2708 4182
rect 2714 4193 2720 4208
rect 2714 4137 2720 4189
rect 2726 4200 2732 4208
rect 2726 4137 2732 4196
rect 2738 4137 2744 4204
rect 2750 4137 2756 4159
rect 2935 4145 2940 4312
rect 2954 4155 2967 4314
rect 3293 4313 3296 4315
rect 3241 4178 3296 4313
rect 3548 4176 3604 4311
rect 3241 4173 3296 4174
rect 3549 4170 3604 4176
rect 2404 3938 2407 3987
rect 2404 3894 2407 3934
rect 2412 3931 2416 4093
rect 2420 4011 2423 4021
rect 2427 3981 2430 3990
rect 2443 3983 2446 3996
rect 2456 3968 2459 4021
rect 2523 4011 2526 4021
rect 2463 3996 2467 4000
rect 2464 3981 2467 3990
rect 2419 3954 2422 3966
rect 2460 3964 2461 3968
rect 2470 3954 2473 4007
rect 2476 3987 2479 3992
rect 2485 3981 2488 3990
rect 2501 3983 2504 3996
rect 2522 3981 2525 3990
rect 2521 3954 2524 3964
rect 2404 3879 2407 3888
rect 2265 3418 2269 3526
rect 2288 3509 2291 3519
rect 2295 3479 2298 3488
rect 2311 3481 2314 3494
rect 2324 3466 2327 3519
rect 2391 3509 2394 3519
rect 2331 3494 2335 3498
rect 2332 3479 2335 3488
rect 2287 3452 2290 3464
rect 2328 3462 2329 3466
rect 2338 3452 2341 3505
rect 2344 3485 2347 3490
rect 2353 3479 2356 3488
rect 2369 3481 2372 3494
rect 2390 3479 2393 3488
rect 2406 3479 2409 3488
rect 2389 3452 2392 3462
rect 2281 3347 2284 3441
rect 2406 3438 2409 3475
rect 2412 3431 2416 3927
rect 2529 3940 2533 4074
rect 2678 4051 2684 4098
rect 2678 4018 2684 4047
rect 2538 3988 2541 3990
rect 2538 3981 2541 3984
rect 2538 3947 2541 3977
rect 2678 3974 2684 4014
rect 2419 3909 2422 3919
rect 2420 3879 2423 3888
rect 2441 3881 2444 3894
rect 2457 3879 2460 3888
rect 2466 3885 2469 3890
rect 2421 3852 2424 3862
rect 2472 3852 2475 3905
rect 2478 3894 2482 3898
rect 2478 3879 2481 3888
rect 2486 3866 2489 3919
rect 2522 3909 2525 3919
rect 2499 3881 2502 3894
rect 2515 3879 2518 3888
rect 2484 3862 2485 3866
rect 2523 3852 2526 3864
rect 2420 3509 2423 3519
rect 2427 3479 2430 3488
rect 2443 3481 2446 3494
rect 2456 3466 2459 3519
rect 2523 3509 2526 3519
rect 2463 3494 2467 3498
rect 2464 3479 2467 3488
rect 2419 3452 2422 3464
rect 2460 3462 2461 3466
rect 2470 3452 2473 3505
rect 2476 3485 2479 3490
rect 2485 3479 2488 3488
rect 2501 3481 2504 3494
rect 2522 3479 2525 3488
rect 2521 3452 2524 3462
rect 2396 3418 2400 3422
rect 2396 3399 2400 3414
rect 2412 3411 2416 3427
rect 2428 3426 2432 3431
rect 2428 3418 2432 3422
rect 2428 3399 2432 3414
rect 2412 3395 2416 3396
rect 2428 3391 2432 3395
rect 2288 3367 2291 3377
rect 2295 3337 2298 3346
rect 2311 3339 2314 3352
rect 2324 3324 2327 3377
rect 2391 3367 2394 3377
rect 2331 3352 2335 3356
rect 2332 3337 2335 3346
rect 2287 3310 2290 3322
rect 2328 3320 2329 3324
rect 2338 3310 2341 3363
rect 2406 3352 2409 3384
rect 2344 3343 2347 3348
rect 2353 3337 2356 3346
rect 2369 3339 2372 3352
rect 2390 3337 2393 3346
rect 2406 3337 2409 3346
rect 2389 3310 2392 3320
rect 2281 3261 2284 3299
rect 2288 3281 2291 3291
rect 2295 3251 2298 3260
rect 2311 3253 2314 3266
rect 2324 3238 2327 3291
rect 2391 3281 2394 3291
rect 2331 3266 2335 3270
rect 2332 3251 2335 3260
rect 2287 3224 2290 3236
rect 2328 3234 2329 3238
rect 2338 3224 2341 3277
rect 2344 3257 2347 3262
rect 2353 3251 2356 3260
rect 2369 3253 2372 3266
rect 2390 3251 2393 3260
rect 2406 3251 2409 3260
rect 2389 3224 2392 3234
rect 2281 3121 2284 3213
rect 2406 3210 2409 3247
rect 2288 3141 2291 3151
rect 2295 3111 2298 3120
rect 2311 3113 2314 3126
rect 2324 3098 2327 3151
rect 2391 3141 2394 3151
rect 2331 3126 2335 3130
rect 2332 3111 2335 3120
rect 2287 3084 2290 3096
rect 2328 3094 2329 3098
rect 2338 3084 2341 3137
rect 2406 3126 2409 3158
rect 2344 3117 2347 3122
rect 2353 3111 2356 3120
rect 2369 3113 2372 3126
rect 2390 3111 2393 3120
rect 2406 3111 2409 3120
rect 2389 3084 2392 3094
rect 2404 2956 2407 3005
rect 2404 2912 2407 2952
rect 2412 2949 2416 3391
rect 2420 3367 2423 3377
rect 2427 3337 2430 3346
rect 2443 3339 2446 3352
rect 2456 3324 2459 3377
rect 2523 3367 2526 3377
rect 2463 3352 2467 3356
rect 2464 3337 2467 3346
rect 2419 3310 2422 3322
rect 2460 3320 2461 3324
rect 2470 3310 2473 3363
rect 2476 3343 2479 3348
rect 2485 3337 2488 3346
rect 2501 3339 2504 3352
rect 2522 3337 2525 3346
rect 2521 3310 2524 3320
rect 2420 3281 2423 3291
rect 2427 3251 2430 3260
rect 2443 3253 2446 3266
rect 2456 3238 2459 3291
rect 2523 3281 2526 3291
rect 2463 3266 2467 3270
rect 2464 3251 2467 3260
rect 2419 3224 2422 3236
rect 2460 3234 2461 3238
rect 2470 3224 2473 3277
rect 2476 3257 2479 3262
rect 2485 3251 2488 3260
rect 2501 3253 2504 3266
rect 2522 3251 2525 3260
rect 2521 3224 2524 3234
rect 2529 3203 2533 3936
rect 2553 3931 2557 3936
rect 2678 3916 2684 3970
rect 2678 3842 2684 3912
rect 2678 3710 2684 3838
rect 2678 3578 2684 3706
rect 2552 3509 2555 3519
rect 2538 3479 2541 3488
rect 2559 3479 2562 3488
rect 2575 3481 2578 3494
rect 2538 3438 2541 3475
rect 2588 3466 2591 3519
rect 2655 3509 2658 3519
rect 2678 3516 2684 3574
rect 2595 3494 2599 3498
rect 2596 3479 2599 3488
rect 2551 3452 2554 3464
rect 2592 3462 2593 3466
rect 2602 3452 2605 3505
rect 2608 3485 2611 3490
rect 2617 3479 2620 3488
rect 2633 3481 2636 3494
rect 2654 3479 2657 3488
rect 2670 3479 2673 3490
rect 2653 3452 2656 3462
rect 2670 3445 2673 3475
rect 2670 3411 2673 3441
rect 2678 3446 2684 3512
rect 2678 3404 2684 3442
rect 2538 3352 2541 3384
rect 2552 3367 2555 3377
rect 2538 3337 2541 3346
rect 2559 3337 2562 3346
rect 2575 3339 2578 3352
rect 2588 3324 2591 3377
rect 2655 3367 2658 3377
rect 2595 3352 2599 3356
rect 2596 3337 2599 3346
rect 2551 3310 2554 3322
rect 2592 3320 2593 3324
rect 2602 3310 2605 3363
rect 2670 3352 2673 3399
rect 2608 3343 2611 3348
rect 2617 3337 2620 3346
rect 2633 3339 2636 3352
rect 2654 3337 2657 3346
rect 2670 3337 2673 3348
rect 2653 3310 2656 3320
rect 2670 3303 2673 3333
rect 2678 3374 2684 3400
rect 2552 3281 2555 3291
rect 2538 3251 2541 3260
rect 2559 3251 2562 3260
rect 2575 3253 2578 3266
rect 2538 3210 2541 3247
rect 2588 3238 2591 3291
rect 2655 3281 2658 3291
rect 2678 3288 2684 3370
rect 2595 3266 2599 3270
rect 2596 3251 2599 3260
rect 2551 3224 2554 3236
rect 2592 3234 2593 3238
rect 2602 3224 2605 3277
rect 2608 3257 2611 3262
rect 2617 3251 2620 3260
rect 2633 3253 2636 3266
rect 2654 3251 2657 3260
rect 2670 3251 2673 3262
rect 2653 3224 2656 3234
rect 2670 3217 2673 3247
rect 2513 3192 2517 3195
rect 2513 3173 2517 3188
rect 2529 3185 2533 3199
rect 2545 3199 2549 3203
rect 2545 3192 2549 3195
rect 2545 3173 2549 3188
rect 2670 3185 2673 3213
rect 2529 3169 2533 3170
rect 2545 3165 2549 3169
rect 2420 3141 2423 3151
rect 2427 3111 2430 3120
rect 2443 3113 2446 3126
rect 2456 3098 2459 3151
rect 2523 3141 2526 3151
rect 2463 3126 2467 3130
rect 2464 3111 2467 3120
rect 2419 3084 2422 3096
rect 2460 3094 2461 3098
rect 2470 3084 2473 3137
rect 2476 3117 2479 3122
rect 2485 3111 2488 3120
rect 2501 3113 2504 3126
rect 2522 3111 2525 3120
rect 2521 3084 2524 3094
rect 2420 3029 2423 3039
rect 2427 2999 2430 3008
rect 2443 3001 2446 3014
rect 2456 2986 2459 3039
rect 2523 3029 2526 3039
rect 2463 3014 2467 3018
rect 2464 2999 2467 3008
rect 2419 2972 2422 2984
rect 2460 2982 2461 2986
rect 2470 2972 2473 3025
rect 2476 3005 2479 3010
rect 2485 2999 2488 3008
rect 2501 3001 2504 3014
rect 2522 2999 2525 3008
rect 2521 2972 2524 2982
rect 2404 2897 2407 2906
rect 2288 2527 2291 2537
rect 2295 2497 2298 2506
rect 2311 2499 2314 2512
rect 2324 2484 2327 2537
rect 2391 2527 2394 2537
rect 2331 2512 2335 2516
rect 2332 2497 2335 2506
rect 2287 2470 2290 2482
rect 2328 2480 2329 2484
rect 2338 2470 2341 2523
rect 2344 2503 2347 2508
rect 2353 2497 2356 2506
rect 2369 2499 2372 2512
rect 2390 2497 2393 2506
rect 2406 2497 2409 2506
rect 2389 2470 2392 2480
rect 2281 2365 2284 2459
rect 2406 2456 2409 2493
rect 2412 2449 2416 2945
rect 2529 2958 2533 3165
rect 2538 3126 2541 3158
rect 2552 3141 2555 3151
rect 2538 3111 2541 3120
rect 2559 3111 2562 3120
rect 2575 3113 2578 3126
rect 2588 3098 2591 3151
rect 2655 3141 2658 3151
rect 2595 3126 2599 3130
rect 2596 3111 2599 3120
rect 2551 3084 2554 3096
rect 2592 3094 2593 3098
rect 2602 3084 2605 3137
rect 2670 3126 2673 3173
rect 2608 3117 2611 3122
rect 2617 3111 2620 3120
rect 2633 3113 2636 3126
rect 2654 3111 2657 3120
rect 2670 3118 2673 3122
rect 2678 3148 2684 3284
rect 2670 3111 2673 3114
rect 2653 3084 2656 3094
rect 2678 3069 2684 3144
rect 2678 3036 2684 3065
rect 2538 3006 2541 3008
rect 2538 2999 2541 3002
rect 2538 2965 2541 2995
rect 2678 2992 2684 3032
rect 2419 2927 2422 2937
rect 2420 2897 2423 2906
rect 2441 2899 2444 2912
rect 2457 2897 2460 2906
rect 2466 2903 2469 2908
rect 2421 2870 2424 2880
rect 2472 2870 2475 2923
rect 2478 2912 2482 2916
rect 2478 2897 2481 2906
rect 2486 2884 2489 2937
rect 2522 2927 2525 2937
rect 2499 2899 2502 2912
rect 2515 2897 2518 2906
rect 2484 2880 2485 2884
rect 2523 2870 2526 2882
rect 2420 2527 2423 2537
rect 2427 2497 2430 2506
rect 2443 2499 2446 2512
rect 2456 2484 2459 2537
rect 2523 2527 2526 2537
rect 2463 2512 2467 2516
rect 2464 2497 2467 2506
rect 2419 2470 2422 2482
rect 2460 2480 2461 2484
rect 2470 2470 2473 2523
rect 2476 2503 2479 2508
rect 2485 2497 2488 2506
rect 2501 2499 2504 2512
rect 2522 2497 2525 2506
rect 2521 2470 2524 2480
rect 2396 2436 2400 2441
rect 2396 2417 2400 2432
rect 2412 2429 2416 2445
rect 2428 2445 2432 2449
rect 2428 2436 2432 2441
rect 2428 2417 2432 2432
rect 2412 2413 2416 2414
rect 2428 2409 2432 2413
rect 2288 2385 2291 2395
rect 2295 2355 2298 2364
rect 2311 2357 2314 2370
rect 2324 2342 2327 2395
rect 2391 2385 2394 2395
rect 2331 2370 2335 2374
rect 2332 2355 2335 2364
rect 2287 2328 2290 2340
rect 2328 2338 2329 2342
rect 2338 2328 2341 2381
rect 2406 2370 2409 2402
rect 2344 2361 2347 2366
rect 2353 2355 2356 2364
rect 2369 2357 2372 2370
rect 2390 2355 2393 2364
rect 2406 2355 2409 2364
rect 2389 2328 2392 2338
rect 2281 2279 2284 2317
rect 2288 2299 2291 2309
rect 2295 2269 2298 2278
rect 2311 2271 2314 2284
rect 2324 2256 2327 2309
rect 2391 2299 2394 2309
rect 2331 2284 2335 2288
rect 2332 2269 2335 2278
rect 2287 2242 2290 2254
rect 2328 2252 2329 2256
rect 2338 2242 2341 2295
rect 2344 2275 2347 2280
rect 2353 2269 2356 2278
rect 2369 2271 2372 2284
rect 2390 2269 2393 2278
rect 2406 2269 2409 2278
rect 2389 2242 2392 2252
rect 2281 2139 2284 2231
rect 2406 2228 2409 2265
rect 2288 2159 2291 2169
rect 2295 2129 2298 2138
rect 2311 2131 2314 2144
rect 2324 2116 2327 2169
rect 2391 2159 2394 2169
rect 2331 2144 2335 2148
rect 2332 2129 2335 2138
rect 2287 2102 2290 2114
rect 2328 2112 2329 2116
rect 2338 2102 2341 2155
rect 2406 2144 2409 2176
rect 2344 2135 2347 2140
rect 2353 2129 2356 2138
rect 2369 2131 2372 2144
rect 2390 2129 2393 2138
rect 2406 2129 2409 2138
rect 2389 2102 2392 2112
rect 2412 2088 2416 2409
rect 2420 2385 2423 2395
rect 2427 2355 2430 2364
rect 2443 2357 2446 2370
rect 2456 2342 2459 2395
rect 2523 2385 2526 2395
rect 2463 2370 2467 2374
rect 2464 2355 2467 2364
rect 2419 2328 2422 2340
rect 2460 2338 2461 2342
rect 2470 2328 2473 2381
rect 2476 2361 2479 2366
rect 2485 2355 2488 2364
rect 2501 2357 2504 2370
rect 2522 2355 2525 2364
rect 2521 2328 2524 2338
rect 2420 2299 2423 2309
rect 2427 2269 2430 2278
rect 2443 2271 2446 2284
rect 2456 2256 2459 2309
rect 2523 2299 2526 2309
rect 2463 2284 2467 2288
rect 2464 2269 2467 2278
rect 2419 2242 2422 2254
rect 2460 2252 2461 2256
rect 2470 2242 2473 2295
rect 2476 2275 2479 2280
rect 2485 2269 2488 2278
rect 2501 2271 2504 2284
rect 2522 2269 2525 2278
rect 2521 2242 2524 2252
rect 2529 2221 2533 2954
rect 2553 2949 2557 2954
rect 2678 2934 2684 2988
rect 2678 2860 2684 2930
rect 2678 2728 2684 2856
rect 2678 2596 2684 2724
rect 2552 2527 2555 2537
rect 2538 2497 2541 2506
rect 2559 2497 2562 2506
rect 2575 2499 2578 2512
rect 2538 2456 2541 2493
rect 2588 2484 2591 2537
rect 2655 2527 2658 2537
rect 2678 2534 2684 2592
rect 2595 2512 2599 2516
rect 2596 2497 2599 2506
rect 2551 2470 2554 2482
rect 2592 2480 2593 2484
rect 2602 2470 2605 2523
rect 2608 2503 2611 2508
rect 2617 2497 2620 2506
rect 2633 2499 2636 2512
rect 2654 2497 2657 2506
rect 2670 2497 2673 2508
rect 2653 2470 2656 2480
rect 2670 2463 2673 2493
rect 2670 2429 2673 2459
rect 2678 2464 2684 2530
rect 2678 2422 2684 2460
rect 2538 2370 2541 2402
rect 2552 2385 2555 2395
rect 2538 2355 2541 2364
rect 2559 2355 2562 2364
rect 2575 2357 2578 2370
rect 2588 2342 2591 2395
rect 2655 2385 2658 2395
rect 2595 2370 2599 2374
rect 2596 2355 2599 2364
rect 2551 2328 2554 2340
rect 2592 2338 2593 2342
rect 2602 2328 2605 2381
rect 2670 2370 2673 2417
rect 2608 2361 2611 2366
rect 2617 2355 2620 2364
rect 2633 2357 2636 2370
rect 2654 2355 2657 2364
rect 2670 2355 2673 2366
rect 2653 2328 2656 2338
rect 2670 2321 2673 2351
rect 2678 2392 2684 2418
rect 2552 2299 2555 2309
rect 2538 2269 2541 2278
rect 2559 2269 2562 2278
rect 2575 2271 2578 2284
rect 2538 2228 2541 2265
rect 2588 2256 2591 2309
rect 2655 2299 2658 2309
rect 2678 2306 2684 2388
rect 2595 2284 2599 2288
rect 2596 2269 2599 2278
rect 2551 2242 2554 2254
rect 2592 2252 2593 2256
rect 2602 2242 2605 2295
rect 2608 2275 2611 2280
rect 2617 2269 2620 2278
rect 2633 2271 2636 2284
rect 2654 2269 2657 2278
rect 2670 2269 2673 2280
rect 2653 2242 2656 2252
rect 2670 2235 2673 2265
rect 2513 2210 2517 2213
rect 2513 2191 2517 2206
rect 2529 2203 2533 2217
rect 2545 2217 2549 2221
rect 2545 2210 2549 2213
rect 2545 2191 2549 2206
rect 2670 2203 2673 2231
rect 2529 2187 2533 2188
rect 2545 2183 2549 2187
rect 2420 2159 2423 2169
rect 2427 2129 2430 2138
rect 2443 2131 2446 2144
rect 2456 2116 2459 2169
rect 2523 2159 2526 2169
rect 2463 2144 2467 2148
rect 2464 2129 2467 2138
rect 2419 2102 2422 2114
rect 2460 2112 2461 2116
rect 2470 2102 2473 2155
rect 2476 2135 2479 2140
rect 2485 2129 2488 2138
rect 2501 2131 2504 2144
rect 2522 2129 2525 2138
rect 2521 2102 2524 2112
rect 2529 2088 2533 2183
rect 2538 2144 2541 2176
rect 2552 2159 2555 2169
rect 2538 2129 2541 2138
rect 2559 2129 2562 2138
rect 2575 2131 2578 2144
rect 2588 2116 2591 2169
rect 2655 2159 2658 2169
rect 2595 2144 2599 2148
rect 2596 2129 2599 2138
rect 2551 2102 2554 2114
rect 2592 2112 2593 2116
rect 2602 2102 2605 2155
rect 2670 2144 2673 2191
rect 2608 2135 2611 2140
rect 2617 2129 2620 2138
rect 2633 2131 2636 2144
rect 2654 2129 2657 2138
rect 2670 2136 2673 2140
rect 2678 2166 2684 2302
rect 2670 2129 2673 2132
rect 2653 2102 2656 2112
rect 2678 2088 2684 2162
rect 2690 3994 2696 4098
rect 2690 3961 2696 3990
rect 2690 3908 2696 3957
rect 2690 3859 2696 3904
rect 2690 3776 2696 3855
rect 2690 3644 2696 3772
rect 2690 3512 2696 3640
rect 2690 3459 2696 3508
rect 2690 3347 2696 3455
rect 2690 3317 2696 3343
rect 2690 3261 2696 3313
rect 2690 3231 2696 3257
rect 2690 3091 2696 3227
rect 2690 3012 2696 3087
rect 2690 2979 2696 3008
rect 2690 2926 2696 2975
rect 2690 2877 2696 2922
rect 2690 2794 2696 2873
rect 2690 2662 2696 2790
rect 2690 2530 2696 2658
rect 2690 2477 2696 2526
rect 2690 2365 2696 2473
rect 2690 2335 2696 2361
rect 2690 2279 2696 2331
rect 2690 2249 2696 2275
rect 2690 2109 2696 2245
rect 2690 2088 2696 2105
rect 2702 3915 2708 4098
rect 2702 3901 2708 3911
rect 2702 3783 2708 3897
rect 2702 3769 2708 3779
rect 2702 3651 2708 3765
rect 2702 3637 2708 3647
rect 2702 3505 2708 3633
rect 2702 3431 2708 3501
rect 2702 2933 2708 3427
rect 2702 2919 2708 2929
rect 2702 2801 2708 2915
rect 2702 2787 2708 2797
rect 2702 2669 2708 2783
rect 2702 2655 2708 2665
rect 2702 2523 2708 2651
rect 2702 2449 2708 2519
rect 2702 2088 2708 2445
rect 2714 3967 2720 4098
rect 2714 3835 2720 3963
rect 2714 3717 2720 3831
rect 2714 3703 2720 3713
rect 2714 3585 2720 3699
rect 2714 3571 2720 3581
rect 2714 3439 2720 3567
rect 2714 2985 2720 3435
rect 2714 2853 2720 2981
rect 2714 2735 2720 2849
rect 2714 2721 2720 2731
rect 2714 2603 2720 2717
rect 2714 2589 2720 2599
rect 2714 2457 2720 2585
rect 2714 2088 2720 2453
rect 2726 3987 2732 4098
rect 2726 3954 2732 3983
rect 2726 3852 2732 3950
rect 2726 3453 2732 3848
rect 2726 3340 2732 3449
rect 2726 3310 2732 3336
rect 2726 3254 2732 3306
rect 2726 3224 2732 3250
rect 2726 3084 2732 3220
rect 2726 3005 2732 3080
rect 2726 2972 2732 3001
rect 2726 2870 2732 2968
rect 2726 2471 2732 2866
rect 2726 2358 2732 2467
rect 2726 2328 2732 2354
rect 2726 2272 2732 2324
rect 2726 2242 2732 2268
rect 2726 2102 2732 2238
rect 2726 2088 2732 2098
rect 2738 4058 2744 4098
rect 2738 4025 2744 4054
rect 2738 3923 2744 4021
rect 2738 3523 2744 3919
rect 2738 3411 2744 3519
rect 2738 3381 2744 3407
rect 2738 3325 2744 3377
rect 2738 3295 2744 3321
rect 2738 3155 2744 3291
rect 2738 3076 2744 3151
rect 2738 3043 2744 3072
rect 2738 2941 2744 3039
rect 2738 2541 2744 2937
rect 2738 2429 2744 2537
rect 2738 2399 2744 2425
rect 2738 2343 2744 2395
rect 2738 2313 2744 2339
rect 2738 2173 2744 2309
rect 2738 2088 2744 2169
rect 2750 3425 2756 4098
rect 2772 4044 2775 4054
rect 2761 4024 2765 4025
rect 2779 4014 2782 4023
rect 2795 4016 2798 4029
rect 2808 4001 2811 4054
rect 2875 4044 2878 4054
rect 2904 4044 2907 4054
rect 2815 4029 2819 4033
rect 2816 4014 2819 4023
rect 2771 3987 2774 3999
rect 2812 3997 2813 4001
rect 2822 3987 2825 4040
rect 2828 4020 2831 4025
rect 2837 4014 2840 4023
rect 2853 4016 2856 4029
rect 2874 4014 2877 4023
rect 2890 4023 2893 4025
rect 2890 4020 2897 4023
rect 2890 4014 2893 4020
rect 2911 4014 2914 4023
rect 2927 4016 2930 4029
rect 2873 3987 2876 3997
rect 2890 3980 2893 4010
rect 2940 4001 2943 4054
rect 3007 4044 3010 4054
rect 3036 4044 3039 4054
rect 2947 4029 2951 4033
rect 2948 4014 2951 4023
rect 2903 3987 2906 3999
rect 2944 3997 2945 4001
rect 2954 3987 2957 4040
rect 2960 4020 2963 4025
rect 2969 4014 2972 4023
rect 2985 4016 2988 4029
rect 3006 4014 3009 4023
rect 3022 4023 3025 4025
rect 3022 4020 3029 4023
rect 3022 4014 3025 4020
rect 3043 4014 3046 4023
rect 3059 4016 3062 4029
rect 3005 3987 3008 3997
rect 2890 3977 2942 3980
rect 2770 3957 2773 3970
rect 2796 3960 2799 3963
rect 2803 3957 2806 3970
rect 2820 3957 2823 3970
rect 2770 3908 2773 3923
rect 2784 3915 2787 3919
rect 2802 3908 2805 3923
rect 2821 3908 2824 3923
rect 2827 3922 2830 3963
rect 2843 3915 2846 3956
rect 2849 3923 2852 3963
rect 2868 3915 2871 3956
rect 2877 3957 2880 3970
rect 2893 3957 2896 3970
rect 2914 3960 2917 3963
rect 2921 3957 2924 3970
rect 2939 3966 2942 3977
rect 3022 3974 3025 4010
rect 3072 4001 3075 4054
rect 3139 4044 3142 4054
rect 3168 4044 3171 4054
rect 3079 4029 3083 4033
rect 3080 4014 3083 4023
rect 3035 3987 3038 3999
rect 3076 3997 3077 4001
rect 3086 3987 3089 4040
rect 3092 4020 3095 4025
rect 3101 4014 3104 4023
rect 3117 4016 3120 4029
rect 3138 4014 3141 4023
rect 3154 4023 3157 4025
rect 3154 4020 3161 4023
rect 3154 4014 3157 4020
rect 3175 4014 3178 4023
rect 3191 4016 3194 4029
rect 3137 3987 3140 3997
rect 3154 3980 3157 4002
rect 3204 4001 3207 4054
rect 3271 4044 3274 4054
rect 3211 4029 3215 4033
rect 3212 4014 3215 4023
rect 3167 3987 3170 3999
rect 3208 3997 3209 4001
rect 3218 3987 3221 4040
rect 3224 4020 3227 4025
rect 3233 4014 3236 4023
rect 3249 4016 3252 4029
rect 3270 4014 3273 4023
rect 3286 4023 3289 4025
rect 3286 4020 3290 4023
rect 3286 4014 3289 4020
rect 3286 4006 3289 4010
rect 3269 3987 3272 3997
rect 3020 3969 3025 3974
rect 3082 3976 3157 3980
rect 2939 3963 2984 3966
rect 2939 3953 2942 3963
rect 2957 3950 2977 3953
rect 2974 3931 2977 3950
rect 2877 3908 2880 3923
rect 2892 3908 2895 3923
rect 2899 3915 2903 3918
rect 2920 3908 2923 3923
rect 2770 3889 2773 3904
rect 2784 3893 2787 3897
rect 2802 3889 2805 3904
rect 2821 3889 2824 3904
rect 2770 3842 2773 3855
rect 2796 3849 2799 3852
rect 2770 3825 2773 3838
rect 2780 3835 2784 3845
rect 2803 3842 2806 3855
rect 2820 3842 2823 3855
rect 2827 3849 2830 3890
rect 2843 3856 2846 3897
rect 2849 3849 2852 3889
rect 2868 3856 2871 3897
rect 2877 3889 2880 3904
rect 2892 3889 2895 3904
rect 2899 3894 2903 3897
rect 2920 3889 2923 3904
rect 2877 3842 2880 3855
rect 2796 3828 2799 3831
rect 2803 3825 2806 3838
rect 2820 3825 2823 3838
rect 2770 3776 2773 3791
rect 2784 3783 2787 3787
rect 2802 3776 2805 3791
rect 2821 3776 2824 3791
rect 2827 3790 2830 3831
rect 2843 3783 2846 3824
rect 2849 3791 2852 3831
rect 2868 3783 2871 3824
rect 2877 3825 2880 3838
rect 2893 3842 2896 3855
rect 2914 3849 2917 3852
rect 2921 3842 2924 3855
rect 2974 3855 2977 3927
rect 2985 3891 2988 3963
rect 3020 3966 3023 3969
rect 3020 3963 3065 3966
rect 3020 3953 3023 3963
rect 2893 3825 2896 3838
rect 2914 3828 2917 3831
rect 2921 3825 2924 3838
rect 2974 3821 2977 3851
rect 2985 3835 2988 3887
rect 2992 3875 2996 3941
rect 2980 3831 2984 3834
rect 2973 3818 2977 3821
rect 2974 3799 2977 3818
rect 2877 3776 2880 3791
rect 2892 3776 2895 3791
rect 2899 3783 2903 3786
rect 2920 3776 2923 3791
rect 2770 3757 2773 3772
rect 2784 3761 2787 3765
rect 2802 3757 2805 3772
rect 2821 3757 2824 3772
rect 2770 3710 2773 3723
rect 2796 3717 2799 3720
rect 2770 3693 2773 3706
rect 2803 3710 2806 3723
rect 2820 3710 2823 3723
rect 2827 3717 2830 3758
rect 2843 3724 2846 3765
rect 2849 3717 2852 3757
rect 2868 3724 2871 3765
rect 2877 3757 2880 3772
rect 2892 3757 2895 3772
rect 2899 3762 2903 3765
rect 2920 3757 2923 3772
rect 2877 3710 2880 3723
rect 2796 3696 2799 3699
rect 2803 3693 2806 3706
rect 2820 3693 2823 3706
rect 2770 3644 2773 3659
rect 2784 3651 2787 3655
rect 2802 3644 2805 3659
rect 2821 3644 2824 3659
rect 2827 3658 2830 3699
rect 2843 3651 2846 3692
rect 2849 3659 2852 3699
rect 2868 3651 2871 3692
rect 2877 3693 2880 3706
rect 2893 3710 2896 3723
rect 2914 3717 2917 3720
rect 2921 3710 2924 3723
rect 2974 3724 2977 3795
rect 2985 3760 2988 3831
rect 2893 3693 2896 3706
rect 2914 3696 2917 3699
rect 2921 3693 2924 3706
rect 2974 3667 2977 3720
rect 2985 3703 2988 3756
rect 2992 3744 2996 3809
rect 2980 3699 2984 3702
rect 3023 3702 3026 3953
rect 3038 3950 3058 3953
rect 3055 3931 3058 3950
rect 3055 3855 3058 3927
rect 3066 3891 3069 3963
rect 3073 3875 3077 3941
rect 3082 3842 3085 3976
rect 3286 3973 3289 4002
rect 3110 3970 3217 3973
rect 3044 3838 3085 3842
rect 3044 3834 3047 3838
rect 3044 3831 3089 3834
rect 3044 3821 3047 3831
rect 3062 3818 3082 3821
rect 3044 3816 3047 3817
rect 3079 3799 3082 3818
rect 3079 3724 3082 3795
rect 3090 3760 3093 3831
rect 3097 3744 3101 3809
rect 2877 3644 2880 3659
rect 2892 3644 2895 3659
rect 2899 3651 2903 3654
rect 2920 3644 2923 3659
rect 2770 3625 2773 3640
rect 2784 3629 2787 3633
rect 2802 3625 2805 3640
rect 2821 3625 2824 3640
rect 2770 3578 2773 3591
rect 2796 3585 2799 3588
rect 2770 3561 2773 3574
rect 2803 3578 2806 3591
rect 2820 3578 2823 3591
rect 2827 3585 2830 3626
rect 2843 3592 2846 3633
rect 2849 3585 2852 3625
rect 2868 3592 2871 3633
rect 2877 3625 2880 3640
rect 2892 3625 2895 3640
rect 2899 3630 2903 3633
rect 2920 3625 2923 3640
rect 2877 3578 2880 3591
rect 2796 3564 2799 3567
rect 2803 3561 2806 3574
rect 2820 3561 2823 3574
rect 2770 3512 2773 3527
rect 2784 3519 2787 3523
rect 2770 3493 2773 3508
rect 2793 3505 2797 3515
rect 2802 3512 2805 3527
rect 2821 3512 2824 3527
rect 2827 3526 2830 3567
rect 2843 3519 2846 3560
rect 2849 3527 2852 3567
rect 2868 3519 2871 3560
rect 2877 3561 2880 3574
rect 2893 3578 2896 3591
rect 2914 3585 2917 3588
rect 2921 3578 2924 3591
rect 2974 3589 2977 3663
rect 2985 3625 2988 3699
rect 3020 3699 3065 3702
rect 3020 3689 3023 3699
rect 3038 3686 3058 3689
rect 2893 3561 2896 3574
rect 2914 3564 2917 3567
rect 2921 3561 2924 3574
rect 2974 3535 2977 3585
rect 2985 3571 2988 3621
rect 2992 3609 2996 3677
rect 3055 3667 3058 3686
rect 3055 3589 3058 3663
rect 3066 3625 3069 3699
rect 3110 3702 3113 3970
rect 3221 3970 3289 3973
rect 3325 3965 3330 4141
rect 3229 3725 3242 3957
rect 3337 3952 3341 4151
rect 3623 4091 3629 4167
rect 3623 4051 3629 4087
rect 3275 3831 3279 3948
rect 3349 3938 3352 3987
rect 3349 3894 3352 3934
rect 3357 3931 3361 4040
rect 3365 4011 3368 4021
rect 3372 3981 3375 3990
rect 3388 3983 3391 3996
rect 3401 3968 3404 4021
rect 3468 4011 3471 4021
rect 3408 3996 3412 4000
rect 3409 3981 3412 3990
rect 3364 3954 3367 3966
rect 3405 3964 3406 3968
rect 3415 3954 3418 4007
rect 3421 3987 3424 3992
rect 3430 3981 3433 3990
rect 3446 3983 3449 3996
rect 3467 3981 3470 3990
rect 3466 3954 3469 3964
rect 3349 3879 3352 3888
rect 3357 3847 3361 3927
rect 3474 3940 3478 4040
rect 3623 4018 3629 4047
rect 3483 3988 3486 3990
rect 3483 3981 3486 3984
rect 3483 3947 3486 3977
rect 3623 3974 3629 4014
rect 3364 3909 3367 3919
rect 3365 3879 3368 3888
rect 3386 3881 3389 3894
rect 3402 3879 3405 3888
rect 3411 3885 3414 3890
rect 3366 3852 3369 3862
rect 3417 3852 3420 3905
rect 3423 3894 3427 3898
rect 3423 3879 3426 3888
rect 3431 3866 3434 3919
rect 3467 3909 3470 3919
rect 3444 3881 3447 3894
rect 3460 3879 3463 3888
rect 3429 3862 3430 3866
rect 3468 3852 3471 3864
rect 3474 3848 3478 3936
rect 3498 3931 3502 3936
rect 3623 3916 3629 3970
rect 3623 3842 3629 3912
rect 3275 3805 3278 3827
rect 3275 3802 3320 3805
rect 3275 3792 3278 3802
rect 3253 3788 3274 3792
rect 3293 3789 3313 3792
rect 3229 3711 3244 3725
rect 3229 3707 3240 3711
rect 3110 3699 3155 3702
rect 3110 3689 3113 3699
rect 3128 3686 3148 3689
rect 3073 3609 3077 3677
rect 3145 3667 3148 3686
rect 3145 3589 3148 3663
rect 3156 3625 3159 3699
rect 3163 3609 3167 3677
rect 2980 3567 2984 3570
rect 2877 3512 2880 3527
rect 2892 3512 2895 3527
rect 2899 3519 2903 3522
rect 2920 3512 2923 3527
rect 2784 3497 2787 3501
rect 2802 3493 2805 3508
rect 2821 3493 2824 3508
rect 2770 3446 2773 3459
rect 2796 3453 2799 3456
rect 2778 3439 2782 3449
rect 2803 3446 2806 3459
rect 2820 3446 2823 3459
rect 2827 3453 2830 3494
rect 2843 3460 2846 3501
rect 2849 3453 2852 3493
rect 2868 3460 2871 3501
rect 2877 3493 2880 3508
rect 2892 3493 2895 3508
rect 2899 3498 2903 3501
rect 2920 3493 2923 3508
rect 2877 3446 2880 3459
rect 2893 3446 2896 3459
rect 2914 3453 2917 3456
rect 2921 3446 2924 3459
rect 2974 3453 2977 3531
rect 2985 3489 2988 3567
rect 2992 3473 2996 3545
rect 3004 3446 3008 3459
rect 3013 3439 3016 3449
rect 3023 3432 3026 3501
rect 3045 3497 3048 3501
rect 3063 3493 3066 3508
rect 3082 3493 3085 3508
rect 3030 3446 3034 3459
rect 3057 3453 3060 3456
rect 3064 3446 3067 3459
rect 3081 3446 3084 3459
rect 3088 3453 3091 3494
rect 3104 3460 3107 3501
rect 3110 3453 3113 3493
rect 3129 3460 3132 3501
rect 3138 3493 3141 3508
rect 3153 3493 3156 3508
rect 3160 3498 3164 3501
rect 3181 3493 3184 3508
rect 3138 3446 3141 3459
rect 3154 3446 3157 3459
rect 3175 3453 3178 3456
rect 3182 3446 3185 3459
rect 3198 3440 3202 3676
rect 3240 3581 3244 3707
rect 3253 3662 3256 3788
rect 3275 3783 3278 3788
rect 3275 3780 3297 3783
rect 3310 3770 3313 3789
rect 3310 3690 3313 3766
rect 3321 3726 3324 3802
rect 3328 3710 3332 3780
rect 3507 3719 3511 3760
rect 3574 3733 3579 3772
rect 3275 3672 3320 3675
rect 3275 3662 3278 3672
rect 3293 3659 3313 3662
rect 3253 3653 3256 3658
rect 3253 3650 3297 3653
rect 3310 3640 3313 3659
rect 3240 3577 3242 3581
rect 3310 3560 3313 3636
rect 3321 3596 3324 3672
rect 3328 3580 3332 3650
rect 3402 3593 3406 3630
rect 3574 3603 3579 3729
rect 3574 3540 3579 3599
rect 3582 3744 3586 3809
rect 3582 3683 3586 3740
rect 3582 3553 3586 3679
rect 3582 3540 3586 3549
rect 3590 3728 3594 3772
rect 3590 3540 3594 3724
rect 3623 3744 3629 3838
rect 3623 3710 3629 3740
rect 3623 3578 3629 3706
rect 3357 3531 3361 3532
rect 3474 3530 3478 3531
rect 3233 3509 3236 3519
rect 3240 3479 3243 3488
rect 3256 3481 3259 3494
rect 3269 3466 3272 3519
rect 3336 3509 3339 3519
rect 3276 3494 3280 3498
rect 3277 3479 3280 3488
rect 3232 3452 3235 3464
rect 3273 3462 3274 3466
rect 3283 3452 3286 3505
rect 3289 3485 3292 3490
rect 3298 3479 3301 3488
rect 3314 3481 3317 3494
rect 3335 3479 3338 3488
rect 3351 3479 3354 3488
rect 3334 3452 3337 3462
rect 3191 3428 3192 3431
rect 2750 2443 2756 3421
rect 3056 3318 3060 3400
rect 3071 3397 3074 3407
rect 3078 3367 3081 3376
rect 3094 3369 3097 3382
rect 3107 3354 3110 3407
rect 3174 3397 3177 3407
rect 3114 3382 3118 3386
rect 3115 3367 3118 3376
rect 3070 3340 3073 3352
rect 3111 3350 3112 3354
rect 3121 3340 3124 3393
rect 3189 3382 3192 3428
rect 3127 3373 3130 3378
rect 3136 3367 3139 3376
rect 3152 3369 3155 3382
rect 3173 3367 3176 3376
rect 3189 3367 3192 3376
rect 3172 3340 3175 3350
rect 3189 3333 3192 3363
rect 3064 3291 3067 3328
rect 3071 3311 3074 3321
rect 3078 3281 3081 3290
rect 3094 3283 3097 3296
rect 3107 3268 3110 3321
rect 3174 3311 3177 3321
rect 3114 3296 3118 3300
rect 3115 3281 3118 3290
rect 3070 3254 3073 3266
rect 3111 3264 3112 3268
rect 3121 3254 3124 3307
rect 3127 3287 3130 3292
rect 3136 3281 3139 3290
rect 3152 3283 3155 3296
rect 3173 3281 3176 3290
rect 3189 3291 3192 3292
rect 3210 3294 3214 3436
rect 3226 3347 3229 3441
rect 3351 3438 3354 3475
rect 3357 3431 3361 3526
rect 3365 3509 3368 3519
rect 3372 3479 3375 3488
rect 3388 3481 3391 3494
rect 3401 3466 3404 3519
rect 3468 3509 3471 3519
rect 3408 3494 3412 3498
rect 3409 3479 3412 3488
rect 3364 3452 3367 3464
rect 3405 3462 3406 3466
rect 3415 3452 3418 3505
rect 3421 3485 3424 3490
rect 3430 3479 3433 3488
rect 3446 3481 3449 3494
rect 3467 3479 3470 3488
rect 3466 3452 3469 3462
rect 3341 3418 3345 3422
rect 3341 3399 3345 3414
rect 3357 3411 3361 3427
rect 3373 3426 3377 3431
rect 3373 3418 3377 3422
rect 3373 3399 3377 3414
rect 3357 3395 3361 3396
rect 3373 3391 3377 3395
rect 3233 3367 3236 3377
rect 3240 3337 3243 3346
rect 3256 3339 3259 3352
rect 3269 3324 3272 3377
rect 3336 3367 3339 3377
rect 3276 3352 3280 3356
rect 3277 3337 3280 3346
rect 3232 3310 3235 3322
rect 3273 3320 3274 3324
rect 3283 3310 3286 3363
rect 3351 3352 3354 3384
rect 3289 3343 3292 3348
rect 3298 3337 3301 3346
rect 3314 3339 3317 3352
rect 3335 3337 3338 3346
rect 3351 3337 3354 3346
rect 3334 3310 3337 3320
rect 3189 3286 3192 3287
rect 3172 3254 3175 3264
rect 3210 3192 3214 3274
rect 3226 3261 3229 3299
rect 3233 3281 3236 3291
rect 3240 3251 3243 3260
rect 3256 3253 3259 3266
rect 3269 3238 3272 3291
rect 3336 3281 3339 3291
rect 3276 3266 3280 3270
rect 3277 3251 3280 3260
rect 3232 3224 3235 3236
rect 3273 3234 3274 3238
rect 3283 3224 3286 3277
rect 3289 3257 3292 3262
rect 3298 3251 3301 3260
rect 3314 3253 3317 3266
rect 3335 3251 3338 3260
rect 3351 3251 3354 3260
rect 3334 3224 3337 3234
rect 3226 3121 3229 3213
rect 3351 3210 3354 3247
rect 3233 3141 3236 3151
rect 3240 3111 3243 3120
rect 3256 3113 3259 3126
rect 3269 3098 3272 3151
rect 3336 3141 3339 3151
rect 3276 3126 3280 3130
rect 3277 3111 3280 3120
rect 3232 3084 3235 3096
rect 3273 3094 3274 3098
rect 3283 3084 3286 3137
rect 3351 3126 3354 3158
rect 3289 3117 3292 3122
rect 3298 3111 3301 3120
rect 3314 3113 3317 3126
rect 3335 3111 3338 3120
rect 3351 3111 3354 3120
rect 3334 3084 3337 3094
rect 2772 3062 2775 3072
rect 2779 3032 2782 3041
rect 2795 3034 2798 3047
rect 2808 3019 2811 3072
rect 2875 3062 2878 3072
rect 2904 3062 2907 3072
rect 2815 3047 2819 3051
rect 2816 3032 2819 3041
rect 2771 3005 2774 3017
rect 2812 3015 2813 3019
rect 2822 3005 2825 3058
rect 2828 3038 2831 3043
rect 2837 3032 2840 3041
rect 2853 3034 2856 3047
rect 2874 3032 2877 3041
rect 2890 3041 2893 3043
rect 2890 3038 2897 3041
rect 2890 3032 2893 3038
rect 2911 3032 2914 3041
rect 2927 3034 2930 3047
rect 2873 3005 2876 3015
rect 2890 2998 2893 3028
rect 2940 3019 2943 3072
rect 3007 3062 3010 3072
rect 3036 3062 3039 3072
rect 2947 3047 2951 3051
rect 2948 3032 2951 3041
rect 2903 3005 2906 3017
rect 2944 3015 2945 3019
rect 2954 3005 2957 3058
rect 2960 3038 2963 3043
rect 2969 3032 2972 3041
rect 2985 3034 2988 3047
rect 3006 3032 3009 3041
rect 3022 3041 3025 3043
rect 3022 3038 3029 3041
rect 3022 3032 3025 3038
rect 3043 3032 3046 3041
rect 3059 3034 3062 3047
rect 3005 3005 3008 3015
rect 2890 2995 2942 2998
rect 2770 2975 2773 2988
rect 2796 2978 2799 2981
rect 2803 2975 2806 2988
rect 2820 2975 2823 2988
rect 2770 2926 2773 2941
rect 2784 2933 2787 2937
rect 2802 2926 2805 2941
rect 2821 2926 2824 2941
rect 2827 2940 2830 2981
rect 2843 2933 2846 2974
rect 2849 2941 2852 2981
rect 2868 2933 2871 2974
rect 2877 2975 2880 2988
rect 2893 2975 2896 2988
rect 2914 2978 2917 2981
rect 2921 2975 2924 2988
rect 2939 2984 2942 2995
rect 3022 2992 3025 3028
rect 3072 3019 3075 3072
rect 3139 3062 3142 3072
rect 3168 3062 3171 3072
rect 3079 3047 3083 3051
rect 3080 3032 3083 3041
rect 3035 3005 3038 3017
rect 3076 3015 3077 3019
rect 3086 3005 3089 3058
rect 3092 3038 3095 3043
rect 3101 3032 3104 3041
rect 3117 3034 3120 3047
rect 3138 3032 3141 3041
rect 3154 3041 3157 3043
rect 3154 3038 3161 3041
rect 3154 3032 3157 3038
rect 3175 3032 3178 3041
rect 3191 3034 3194 3047
rect 3137 3005 3140 3015
rect 3154 2998 3157 3020
rect 3204 3019 3207 3072
rect 3271 3062 3274 3072
rect 3211 3047 3215 3051
rect 3212 3032 3215 3041
rect 3167 3005 3170 3017
rect 3208 3015 3209 3019
rect 3218 3005 3221 3058
rect 3224 3038 3227 3043
rect 3233 3032 3236 3041
rect 3249 3034 3252 3047
rect 3270 3032 3273 3041
rect 3286 3041 3289 3043
rect 3286 3038 3290 3041
rect 3286 3032 3289 3038
rect 3286 3024 3289 3028
rect 3269 3005 3272 3015
rect 3020 2987 3025 2992
rect 3082 2994 3157 2998
rect 2939 2981 2984 2984
rect 2939 2971 2942 2981
rect 2957 2968 2977 2971
rect 2974 2949 2977 2968
rect 2877 2926 2880 2941
rect 2892 2926 2895 2941
rect 2899 2933 2903 2936
rect 2920 2926 2923 2941
rect 2770 2907 2773 2922
rect 2784 2911 2787 2915
rect 2802 2907 2805 2922
rect 2821 2907 2824 2922
rect 2770 2860 2773 2873
rect 2796 2867 2799 2870
rect 2770 2843 2773 2856
rect 2780 2853 2784 2863
rect 2803 2860 2806 2873
rect 2820 2860 2823 2873
rect 2827 2867 2830 2908
rect 2843 2874 2846 2915
rect 2849 2867 2852 2907
rect 2868 2874 2871 2915
rect 2877 2907 2880 2922
rect 2892 2907 2895 2922
rect 2899 2912 2903 2915
rect 2920 2907 2923 2922
rect 2877 2860 2880 2873
rect 2796 2846 2799 2849
rect 2803 2843 2806 2856
rect 2820 2843 2823 2856
rect 2770 2794 2773 2809
rect 2784 2801 2787 2805
rect 2802 2794 2805 2809
rect 2821 2794 2824 2809
rect 2827 2808 2830 2849
rect 2843 2801 2846 2842
rect 2849 2809 2852 2849
rect 2868 2801 2871 2842
rect 2877 2843 2880 2856
rect 2893 2860 2896 2873
rect 2914 2867 2917 2870
rect 2921 2860 2924 2873
rect 2974 2873 2977 2945
rect 2985 2909 2988 2981
rect 3020 2984 3023 2987
rect 3020 2981 3065 2984
rect 3020 2971 3023 2981
rect 2893 2843 2896 2856
rect 2914 2846 2917 2849
rect 2921 2843 2924 2856
rect 2974 2839 2977 2869
rect 2985 2853 2988 2905
rect 2992 2893 2996 2959
rect 2980 2849 2984 2852
rect 2973 2836 2977 2839
rect 2974 2817 2977 2836
rect 2877 2794 2880 2809
rect 2892 2794 2895 2809
rect 2899 2801 2903 2804
rect 2920 2794 2923 2809
rect 2770 2775 2773 2790
rect 2784 2779 2787 2783
rect 2802 2775 2805 2790
rect 2821 2775 2824 2790
rect 2770 2728 2773 2741
rect 2796 2735 2799 2738
rect 2770 2711 2773 2724
rect 2803 2728 2806 2741
rect 2820 2728 2823 2741
rect 2827 2735 2830 2776
rect 2843 2742 2846 2783
rect 2849 2735 2852 2775
rect 2868 2742 2871 2783
rect 2877 2775 2880 2790
rect 2892 2775 2895 2790
rect 2899 2780 2903 2783
rect 2920 2775 2923 2790
rect 2877 2728 2880 2741
rect 2796 2714 2799 2717
rect 2803 2711 2806 2724
rect 2820 2711 2823 2724
rect 2770 2662 2773 2677
rect 2784 2669 2787 2673
rect 2802 2662 2805 2677
rect 2821 2662 2824 2677
rect 2827 2676 2830 2717
rect 2843 2669 2846 2710
rect 2849 2677 2852 2717
rect 2868 2669 2871 2710
rect 2877 2711 2880 2724
rect 2893 2728 2896 2741
rect 2914 2735 2917 2738
rect 2921 2728 2924 2741
rect 2974 2742 2977 2813
rect 2985 2778 2988 2849
rect 2893 2711 2896 2724
rect 2914 2714 2917 2717
rect 2921 2711 2924 2724
rect 2974 2685 2977 2738
rect 2985 2721 2988 2774
rect 2992 2762 2996 2827
rect 2980 2717 2984 2720
rect 3023 2720 3026 2971
rect 3038 2968 3058 2971
rect 3055 2949 3058 2968
rect 3055 2873 3058 2945
rect 3066 2909 3069 2981
rect 3073 2893 3077 2959
rect 3082 2860 3085 2994
rect 3286 2991 3289 3020
rect 3110 2988 3217 2991
rect 3044 2856 3085 2860
rect 3044 2852 3047 2856
rect 3044 2849 3089 2852
rect 3044 2839 3047 2849
rect 3062 2836 3082 2839
rect 3044 2834 3047 2835
rect 3079 2817 3082 2836
rect 3079 2742 3082 2813
rect 3090 2778 3093 2849
rect 3097 2762 3101 2827
rect 2877 2662 2880 2677
rect 2892 2662 2895 2677
rect 2899 2669 2903 2672
rect 2920 2662 2923 2677
rect 2770 2643 2773 2658
rect 2784 2647 2787 2651
rect 2802 2643 2805 2658
rect 2821 2643 2824 2658
rect 2770 2596 2773 2609
rect 2796 2603 2799 2606
rect 2770 2579 2773 2592
rect 2803 2596 2806 2609
rect 2820 2596 2823 2609
rect 2827 2603 2830 2644
rect 2843 2610 2846 2651
rect 2849 2603 2852 2643
rect 2868 2610 2871 2651
rect 2877 2643 2880 2658
rect 2892 2643 2895 2658
rect 2899 2648 2903 2651
rect 2920 2643 2923 2658
rect 2877 2596 2880 2609
rect 2796 2582 2799 2585
rect 2803 2579 2806 2592
rect 2820 2579 2823 2592
rect 2770 2530 2773 2545
rect 2784 2537 2787 2541
rect 2770 2511 2773 2526
rect 2793 2523 2797 2533
rect 2802 2530 2805 2545
rect 2821 2530 2824 2545
rect 2827 2544 2830 2585
rect 2843 2537 2846 2578
rect 2849 2545 2852 2585
rect 2868 2537 2871 2578
rect 2877 2579 2880 2592
rect 2893 2596 2896 2609
rect 2914 2603 2917 2606
rect 2921 2596 2924 2609
rect 2974 2607 2977 2681
rect 2985 2643 2988 2717
rect 3020 2717 3065 2720
rect 3020 2707 3023 2717
rect 3038 2704 3058 2707
rect 2893 2579 2896 2592
rect 2914 2582 2917 2585
rect 2921 2579 2924 2592
rect 2974 2553 2977 2603
rect 2985 2589 2988 2639
rect 2992 2627 2996 2695
rect 3055 2685 3058 2704
rect 3055 2607 3058 2681
rect 3066 2643 3069 2717
rect 3110 2720 3113 2988
rect 3221 2988 3289 2991
rect 3349 2956 3352 3005
rect 3349 2912 3352 2952
rect 3357 2949 3361 3391
rect 3365 3367 3368 3377
rect 3372 3337 3375 3346
rect 3388 3339 3391 3352
rect 3401 3324 3404 3377
rect 3468 3367 3471 3377
rect 3408 3352 3412 3356
rect 3409 3337 3412 3346
rect 3364 3310 3367 3322
rect 3405 3320 3406 3324
rect 3415 3310 3418 3363
rect 3421 3343 3424 3348
rect 3430 3337 3433 3346
rect 3446 3339 3449 3352
rect 3467 3337 3470 3346
rect 3466 3310 3469 3320
rect 3365 3281 3368 3291
rect 3372 3251 3375 3260
rect 3388 3253 3391 3266
rect 3401 3238 3404 3291
rect 3468 3281 3471 3291
rect 3408 3266 3412 3270
rect 3409 3251 3412 3260
rect 3364 3224 3367 3236
rect 3405 3234 3406 3238
rect 3415 3224 3418 3277
rect 3421 3257 3424 3262
rect 3430 3251 3433 3260
rect 3446 3253 3449 3266
rect 3467 3251 3470 3260
rect 3466 3224 3469 3234
rect 3474 3203 3478 3525
rect 3497 3509 3500 3519
rect 3483 3479 3486 3488
rect 3504 3479 3507 3488
rect 3520 3481 3523 3494
rect 3483 3438 3486 3475
rect 3533 3466 3536 3519
rect 3600 3509 3603 3519
rect 3623 3516 3629 3574
rect 3540 3494 3544 3498
rect 3541 3479 3544 3488
rect 3496 3452 3499 3464
rect 3537 3462 3538 3466
rect 3547 3452 3550 3505
rect 3553 3485 3556 3490
rect 3562 3479 3565 3488
rect 3578 3481 3581 3494
rect 3599 3479 3602 3488
rect 3615 3479 3618 3490
rect 3598 3452 3601 3462
rect 3615 3445 3618 3475
rect 3615 3411 3618 3441
rect 3623 3446 3629 3512
rect 3623 3404 3629 3442
rect 3483 3352 3486 3384
rect 3497 3367 3500 3377
rect 3483 3337 3486 3346
rect 3504 3337 3507 3346
rect 3520 3339 3523 3352
rect 3533 3324 3536 3377
rect 3600 3367 3603 3377
rect 3540 3352 3544 3356
rect 3541 3337 3544 3346
rect 3496 3310 3499 3322
rect 3537 3320 3538 3324
rect 3547 3310 3550 3363
rect 3615 3352 3618 3399
rect 3553 3343 3556 3348
rect 3562 3337 3565 3346
rect 3578 3339 3581 3352
rect 3599 3337 3602 3346
rect 3615 3337 3618 3348
rect 3598 3310 3601 3320
rect 3615 3303 3618 3333
rect 3623 3374 3629 3400
rect 3497 3281 3500 3291
rect 3483 3251 3486 3260
rect 3504 3251 3507 3260
rect 3520 3253 3523 3266
rect 3483 3210 3486 3247
rect 3533 3238 3536 3291
rect 3600 3281 3603 3291
rect 3623 3288 3629 3370
rect 3540 3266 3544 3270
rect 3541 3251 3544 3260
rect 3496 3224 3499 3236
rect 3537 3234 3538 3238
rect 3547 3224 3550 3277
rect 3553 3257 3556 3262
rect 3562 3251 3565 3260
rect 3578 3253 3581 3266
rect 3599 3251 3602 3260
rect 3615 3251 3618 3262
rect 3598 3224 3601 3234
rect 3615 3217 3618 3247
rect 3458 3192 3462 3195
rect 3458 3173 3462 3188
rect 3474 3185 3478 3199
rect 3490 3199 3494 3203
rect 3490 3192 3494 3195
rect 3490 3173 3494 3188
rect 3615 3185 3618 3213
rect 3474 3169 3478 3170
rect 3490 3165 3494 3169
rect 3365 3141 3368 3151
rect 3372 3111 3375 3120
rect 3388 3113 3391 3126
rect 3401 3098 3404 3151
rect 3468 3141 3471 3151
rect 3408 3126 3412 3130
rect 3409 3111 3412 3120
rect 3364 3084 3367 3096
rect 3405 3094 3406 3098
rect 3415 3084 3418 3137
rect 3421 3117 3424 3122
rect 3430 3111 3433 3120
rect 3446 3113 3449 3126
rect 3467 3111 3470 3120
rect 3466 3084 3469 3094
rect 3365 3029 3368 3039
rect 3372 2999 3375 3008
rect 3388 3001 3391 3014
rect 3401 2986 3404 3039
rect 3468 3029 3471 3039
rect 3408 3014 3412 3018
rect 3409 2999 3412 3008
rect 3364 2972 3367 2984
rect 3405 2982 3406 2986
rect 3415 2972 3418 3025
rect 3421 3005 3424 3010
rect 3430 2999 3433 3008
rect 3446 3001 3449 3014
rect 3467 2999 3470 3008
rect 3466 2972 3469 2982
rect 3349 2897 3352 2906
rect 3110 2717 3155 2720
rect 3110 2707 3113 2717
rect 3128 2704 3148 2707
rect 3073 2627 3077 2695
rect 3145 2685 3148 2704
rect 3145 2607 3148 2681
rect 3156 2643 3159 2717
rect 3163 2627 3167 2695
rect 2980 2585 2984 2588
rect 2877 2530 2880 2545
rect 2892 2530 2895 2545
rect 2899 2537 2903 2540
rect 2920 2530 2923 2545
rect 2784 2515 2787 2519
rect 2802 2511 2805 2526
rect 2821 2511 2824 2526
rect 2770 2464 2773 2477
rect 2796 2471 2799 2474
rect 2778 2457 2782 2467
rect 2803 2464 2806 2477
rect 2820 2464 2823 2477
rect 2827 2471 2830 2512
rect 2843 2478 2846 2519
rect 2849 2471 2852 2511
rect 2868 2478 2871 2519
rect 2877 2511 2880 2526
rect 2892 2511 2895 2526
rect 2899 2516 2903 2519
rect 2920 2511 2923 2526
rect 2877 2464 2880 2477
rect 2893 2464 2896 2477
rect 2914 2471 2917 2474
rect 2921 2464 2924 2477
rect 2974 2471 2977 2549
rect 2985 2507 2988 2585
rect 2992 2491 2996 2563
rect 3004 2464 3008 2477
rect 3013 2457 3016 2467
rect 3023 2450 3026 2519
rect 3045 2515 3048 2519
rect 3063 2511 3066 2526
rect 3082 2511 3085 2526
rect 3030 2464 3034 2477
rect 3057 2471 3060 2474
rect 3064 2464 3067 2477
rect 3081 2464 3084 2477
rect 3088 2471 3091 2512
rect 3104 2478 3107 2519
rect 3110 2471 3113 2511
rect 3129 2478 3132 2519
rect 3138 2511 3141 2526
rect 3153 2511 3156 2526
rect 3160 2516 3164 2519
rect 3181 2511 3184 2526
rect 3138 2464 3141 2477
rect 3154 2464 3157 2477
rect 3175 2471 3178 2474
rect 3182 2464 3185 2477
rect 3198 2458 3202 2694
rect 3233 2527 3236 2537
rect 3240 2497 3243 2506
rect 3256 2499 3259 2512
rect 3269 2484 3272 2537
rect 3336 2527 3339 2537
rect 3276 2512 3280 2516
rect 3277 2497 3280 2506
rect 3232 2470 3235 2482
rect 3273 2480 3274 2484
rect 3283 2470 3286 2523
rect 3289 2503 3292 2508
rect 3298 2497 3301 2506
rect 3314 2499 3317 2512
rect 3335 2497 3338 2506
rect 3351 2497 3354 2506
rect 3334 2470 3337 2480
rect 3191 2446 3192 2449
rect 2750 2088 2756 2439
rect 3056 2336 3060 2418
rect 3071 2415 3074 2425
rect 3078 2385 3081 2394
rect 3094 2387 3097 2400
rect 3107 2372 3110 2425
rect 3174 2415 3177 2425
rect 3114 2400 3118 2404
rect 3115 2385 3118 2394
rect 3070 2358 3073 2370
rect 3111 2368 3112 2372
rect 3121 2358 3124 2411
rect 3189 2400 3192 2446
rect 3127 2391 3130 2396
rect 3136 2385 3139 2394
rect 3152 2387 3155 2400
rect 3173 2385 3176 2394
rect 3189 2385 3192 2394
rect 3172 2358 3175 2368
rect 3189 2351 3192 2381
rect 3064 2309 3067 2346
rect 3071 2329 3074 2339
rect 3078 2299 3081 2308
rect 3094 2301 3097 2314
rect 3107 2286 3110 2339
rect 3174 2329 3177 2339
rect 3114 2314 3118 2318
rect 3115 2299 3118 2308
rect 3070 2272 3073 2284
rect 3111 2282 3112 2286
rect 3121 2272 3124 2325
rect 3127 2305 3130 2310
rect 3136 2299 3139 2308
rect 3152 2301 3155 2314
rect 3173 2299 3176 2308
rect 3189 2309 3192 2310
rect 3210 2312 3214 2454
rect 3226 2365 3229 2459
rect 3351 2456 3354 2493
rect 3357 2449 3361 2945
rect 3474 2958 3478 3165
rect 3483 3126 3486 3158
rect 3497 3141 3500 3151
rect 3483 3111 3486 3120
rect 3504 3111 3507 3120
rect 3520 3113 3523 3126
rect 3533 3098 3536 3151
rect 3600 3141 3603 3151
rect 3540 3126 3544 3130
rect 3541 3111 3544 3120
rect 3496 3084 3499 3096
rect 3537 3094 3538 3098
rect 3547 3084 3550 3137
rect 3615 3126 3618 3173
rect 3553 3117 3556 3122
rect 3562 3111 3565 3120
rect 3578 3113 3581 3126
rect 3599 3111 3602 3120
rect 3615 3118 3618 3122
rect 3623 3148 3629 3284
rect 3615 3111 3618 3114
rect 3598 3084 3601 3094
rect 3623 3069 3629 3144
rect 3623 3036 3629 3065
rect 3483 3007 3486 3008
rect 3483 3002 3487 3003
rect 3483 2999 3486 3002
rect 3483 2965 3486 2995
rect 3623 2992 3629 3032
rect 3364 2927 3367 2937
rect 3365 2897 3368 2906
rect 3386 2899 3389 2912
rect 3402 2897 3405 2906
rect 3411 2903 3414 2908
rect 3366 2870 3369 2880
rect 3417 2870 3420 2923
rect 3423 2912 3427 2916
rect 3423 2897 3426 2906
rect 3431 2884 3434 2937
rect 3467 2927 3470 2937
rect 3444 2899 3447 2912
rect 3460 2897 3463 2906
rect 3429 2880 3430 2884
rect 3468 2870 3471 2882
rect 3365 2527 3368 2537
rect 3372 2497 3375 2506
rect 3388 2499 3391 2512
rect 3401 2484 3404 2537
rect 3468 2527 3471 2537
rect 3408 2512 3412 2516
rect 3409 2497 3412 2506
rect 3364 2470 3367 2482
rect 3405 2480 3406 2484
rect 3415 2470 3418 2523
rect 3421 2503 3424 2508
rect 3430 2497 3433 2506
rect 3446 2499 3449 2512
rect 3467 2497 3470 2506
rect 3466 2470 3469 2480
rect 3341 2436 3345 2441
rect 3341 2417 3345 2432
rect 3357 2429 3361 2445
rect 3373 2445 3377 2449
rect 3373 2436 3377 2441
rect 3373 2417 3377 2432
rect 3357 2413 3361 2414
rect 3373 2409 3377 2413
rect 3233 2385 3236 2395
rect 3240 2355 3243 2364
rect 3256 2357 3259 2370
rect 3269 2342 3272 2395
rect 3336 2385 3339 2395
rect 3276 2370 3280 2374
rect 3277 2355 3280 2364
rect 3232 2328 3235 2340
rect 3273 2338 3274 2342
rect 3283 2328 3286 2381
rect 3351 2370 3354 2402
rect 3289 2361 3292 2366
rect 3298 2355 3301 2364
rect 3314 2357 3317 2370
rect 3335 2355 3338 2364
rect 3351 2355 3354 2364
rect 3334 2328 3337 2338
rect 3189 2304 3192 2305
rect 3172 2272 3175 2282
rect 3210 2210 3214 2292
rect 3226 2279 3229 2317
rect 3233 2299 3236 2309
rect 3240 2269 3243 2278
rect 3256 2271 3259 2284
rect 3269 2256 3272 2309
rect 3336 2299 3339 2309
rect 3276 2284 3280 2288
rect 3277 2269 3280 2278
rect 3232 2242 3235 2254
rect 3273 2252 3274 2256
rect 3283 2242 3286 2295
rect 3289 2275 3292 2280
rect 3298 2269 3301 2278
rect 3314 2271 3317 2284
rect 3335 2269 3338 2278
rect 3351 2269 3354 2278
rect 3334 2242 3337 2252
rect 3226 2139 3229 2231
rect 3351 2228 3354 2265
rect 3233 2159 3236 2169
rect 3240 2129 3243 2138
rect 3256 2131 3259 2144
rect 3269 2116 3272 2169
rect 3336 2159 3339 2169
rect 3276 2144 3280 2148
rect 3277 2129 3280 2138
rect 3232 2102 3235 2114
rect 3273 2112 3274 2116
rect 3283 2102 3286 2155
rect 3351 2144 3354 2176
rect 3289 2135 3292 2140
rect 3298 2129 3301 2138
rect 3314 2131 3317 2144
rect 3335 2129 3338 2138
rect 3351 2129 3354 2138
rect 3334 2102 3337 2112
rect 3357 2088 3361 2409
rect 3365 2385 3368 2395
rect 3372 2355 3375 2364
rect 3388 2357 3391 2370
rect 3401 2342 3404 2395
rect 3468 2385 3471 2395
rect 3408 2370 3412 2374
rect 3409 2355 3412 2364
rect 3364 2328 3367 2340
rect 3405 2338 3406 2342
rect 3415 2328 3418 2381
rect 3421 2361 3424 2366
rect 3430 2355 3433 2364
rect 3446 2357 3449 2370
rect 3467 2355 3470 2364
rect 3466 2328 3469 2338
rect 3365 2299 3368 2309
rect 3372 2269 3375 2278
rect 3388 2271 3391 2284
rect 3401 2256 3404 2309
rect 3468 2299 3471 2309
rect 3408 2284 3412 2288
rect 3409 2269 3412 2278
rect 3364 2242 3367 2254
rect 3405 2252 3406 2256
rect 3415 2242 3418 2295
rect 3421 2275 3424 2280
rect 3430 2269 3433 2278
rect 3446 2271 3449 2284
rect 3467 2269 3470 2278
rect 3466 2242 3469 2252
rect 3474 2221 3478 2954
rect 3498 2949 3502 2954
rect 3623 2934 3629 2988
rect 3623 2860 3629 2930
rect 3623 2728 3629 2856
rect 3623 2596 3629 2724
rect 3497 2527 3500 2537
rect 3483 2497 3486 2506
rect 3504 2497 3507 2506
rect 3520 2499 3523 2512
rect 3483 2456 3486 2493
rect 3533 2484 3536 2537
rect 3600 2527 3603 2537
rect 3623 2534 3629 2592
rect 3540 2512 3544 2516
rect 3541 2497 3544 2506
rect 3496 2470 3499 2482
rect 3537 2480 3538 2484
rect 3547 2470 3550 2523
rect 3553 2503 3556 2508
rect 3562 2497 3565 2506
rect 3578 2499 3581 2512
rect 3599 2497 3602 2506
rect 3615 2497 3618 2508
rect 3598 2470 3601 2480
rect 3615 2463 3618 2493
rect 3615 2429 3618 2459
rect 3623 2464 3629 2530
rect 3623 2422 3629 2460
rect 3483 2370 3486 2402
rect 3497 2385 3500 2395
rect 3483 2355 3486 2364
rect 3504 2355 3507 2364
rect 3520 2357 3523 2370
rect 3533 2342 3536 2395
rect 3600 2385 3603 2395
rect 3540 2370 3544 2374
rect 3541 2355 3544 2364
rect 3496 2328 3499 2340
rect 3537 2338 3538 2342
rect 3547 2328 3550 2381
rect 3615 2370 3618 2417
rect 3553 2361 3556 2366
rect 3562 2355 3565 2364
rect 3578 2357 3581 2370
rect 3599 2355 3602 2364
rect 3615 2355 3618 2366
rect 3598 2328 3601 2338
rect 3615 2321 3618 2351
rect 3623 2392 3629 2418
rect 3497 2299 3500 2309
rect 3483 2269 3486 2278
rect 3504 2269 3507 2278
rect 3520 2271 3523 2284
rect 3483 2228 3486 2265
rect 3533 2256 3536 2309
rect 3600 2299 3603 2309
rect 3623 2306 3629 2388
rect 3540 2284 3544 2288
rect 3541 2269 3544 2278
rect 3496 2242 3499 2254
rect 3537 2252 3538 2256
rect 3547 2242 3550 2295
rect 3553 2275 3556 2280
rect 3562 2269 3565 2278
rect 3578 2271 3581 2284
rect 3599 2269 3602 2278
rect 3615 2269 3618 2280
rect 3598 2242 3601 2252
rect 3615 2235 3618 2265
rect 3458 2210 3462 2213
rect 3458 2191 3462 2206
rect 3474 2203 3478 2217
rect 3490 2217 3494 2221
rect 3490 2210 3494 2213
rect 3490 2191 3494 2206
rect 3615 2203 3618 2231
rect 3474 2187 3478 2188
rect 3490 2183 3494 2187
rect 3365 2159 3368 2169
rect 3372 2129 3375 2138
rect 3388 2131 3391 2144
rect 3401 2116 3404 2169
rect 3468 2159 3471 2169
rect 3408 2144 3412 2148
rect 3409 2129 3412 2138
rect 3364 2102 3367 2114
rect 3405 2112 3406 2116
rect 3415 2102 3418 2155
rect 3421 2135 3424 2140
rect 3430 2129 3433 2138
rect 3446 2131 3449 2144
rect 3467 2129 3470 2138
rect 3466 2102 3469 2112
rect 3474 2088 3478 2183
rect 3483 2144 3486 2176
rect 3497 2159 3500 2169
rect 3483 2129 3486 2138
rect 3504 2129 3507 2138
rect 3520 2131 3523 2144
rect 3533 2116 3536 2169
rect 3600 2159 3603 2169
rect 3540 2144 3544 2148
rect 3541 2129 3544 2138
rect 3496 2102 3499 2114
rect 3537 2112 3538 2116
rect 3547 2102 3550 2155
rect 3615 2144 3618 2191
rect 3553 2135 3556 2140
rect 3562 2129 3565 2138
rect 3578 2131 3581 2144
rect 3599 2129 3602 2138
rect 3615 2136 3618 2140
rect 3623 2166 3629 2302
rect 3615 2129 3618 2132
rect 3598 2102 3601 2112
rect 3623 2088 3629 2162
rect 3635 4099 3641 4174
rect 3635 3994 3641 4095
rect 3635 3961 3641 3990
rect 3635 3908 3641 3957
rect 3635 3859 3641 3904
rect 3635 3776 3641 3855
rect 3635 3737 3641 3772
rect 3635 3644 3641 3733
rect 3635 3512 3641 3640
rect 3635 3459 3641 3508
rect 3635 3347 3641 3455
rect 3635 3317 3641 3343
rect 3635 3261 3641 3313
rect 3635 3231 3641 3257
rect 3635 3091 3641 3227
rect 3635 3012 3641 3087
rect 3635 2979 3641 3008
rect 3635 2926 3641 2975
rect 3635 2877 3641 2922
rect 3635 2794 3641 2873
rect 3635 2662 3641 2790
rect 3635 2530 3641 2658
rect 3635 2477 3641 2526
rect 3635 2365 3641 2473
rect 3635 2335 3641 2361
rect 3635 2279 3641 2331
rect 3635 2249 3641 2275
rect 3635 2109 3641 2245
rect 3635 2088 3641 2105
rect 3647 4107 3653 4182
rect 3647 3915 3653 4103
rect 3647 3901 3653 3911
rect 3647 3783 3653 3897
rect 3647 3769 3653 3779
rect 3647 3719 3653 3765
rect 3647 3651 3653 3715
rect 3647 3637 3653 3647
rect 3647 3505 3653 3633
rect 3647 3431 3653 3501
rect 3647 2933 3653 3427
rect 3647 2919 3653 2929
rect 3647 2801 3653 2915
rect 3647 2787 3653 2797
rect 3647 2669 3653 2783
rect 3647 2655 3653 2665
rect 3647 2523 3653 2651
rect 3647 2449 3653 2519
rect 3647 2088 3653 2445
rect 3659 4115 3665 4189
rect 3659 3967 3665 4111
rect 3659 3835 3665 3963
rect 3659 3756 3665 3831
rect 3659 3717 3665 3752
rect 3659 3703 3665 3713
rect 3659 3585 3665 3699
rect 3659 3571 3665 3581
rect 3659 3439 3665 3567
rect 3659 2985 3665 3435
rect 3659 2853 3665 2981
rect 3659 2735 3665 2849
rect 3659 2721 3665 2731
rect 3659 2603 3665 2717
rect 3659 2589 3665 2599
rect 3659 2457 3665 2585
rect 3659 2088 3665 2453
rect 3671 4123 3677 4196
rect 3671 3987 3677 4119
rect 3671 3954 3677 3983
rect 3671 3852 3677 3950
rect 3671 3593 3677 3848
rect 3671 3453 3677 3589
rect 3671 3340 3677 3449
rect 3671 3310 3677 3336
rect 3671 3254 3677 3306
rect 3671 3224 3677 3250
rect 3671 3084 3677 3220
rect 3671 3005 3677 3080
rect 3671 2972 3677 3001
rect 3671 2870 3677 2968
rect 3671 2471 3677 2866
rect 3671 2358 3677 2467
rect 3671 2328 3677 2354
rect 3671 2272 3677 2324
rect 3671 2242 3677 2268
rect 3671 2102 3677 2238
rect 3671 2088 3677 2098
rect 3683 4058 3689 4204
rect 3683 4025 3689 4054
rect 3683 3923 3689 4021
rect 3683 3623 3689 3919
rect 3683 3523 3689 3619
rect 3683 3411 3689 3519
rect 3683 3381 3689 3407
rect 3683 3325 3689 3377
rect 3683 3295 3689 3321
rect 3683 3155 3689 3291
rect 3683 3076 3689 3151
rect 3683 3043 3689 3072
rect 3683 2941 3689 3039
rect 3683 2541 3689 2937
rect 3683 2429 3689 2537
rect 3683 2399 3689 2425
rect 3683 2343 3689 2395
rect 3683 2313 3689 2339
rect 3683 2173 3689 2309
rect 3683 2088 3689 2169
rect 3695 3728 3701 4159
rect 3717 4044 3720 4054
rect 3724 4014 3727 4023
rect 3740 4016 3743 4029
rect 3753 4001 3756 4054
rect 3820 4044 3823 4054
rect 3849 4044 3852 4054
rect 3760 4029 3764 4033
rect 3761 4014 3764 4023
rect 3716 3987 3719 3999
rect 3757 3997 3758 4001
rect 3767 3987 3770 4040
rect 3773 4020 3776 4025
rect 3782 4014 3785 4023
rect 3798 4016 3801 4029
rect 3819 4014 3822 4023
rect 3835 4023 3838 4025
rect 3835 4020 3842 4023
rect 3835 4014 3838 4020
rect 3856 4014 3859 4023
rect 3872 4016 3875 4029
rect 3818 3987 3821 3997
rect 3835 3980 3838 4010
rect 3885 4001 3888 4054
rect 3952 4044 3955 4054
rect 3981 4044 3984 4054
rect 3892 4029 3896 4033
rect 3893 4014 3896 4023
rect 3848 3987 3851 3999
rect 3889 3997 3890 4001
rect 3899 3987 3902 4040
rect 3905 4020 3908 4025
rect 3914 4014 3917 4023
rect 3930 4016 3933 4029
rect 3951 4014 3954 4023
rect 3967 4023 3970 4025
rect 3967 4020 3974 4023
rect 3967 4014 3970 4020
rect 3988 4014 3991 4023
rect 4004 4016 4007 4029
rect 3950 3987 3953 3997
rect 3835 3977 3887 3980
rect 3715 3957 3718 3970
rect 3741 3960 3744 3963
rect 3748 3957 3751 3970
rect 3765 3957 3768 3970
rect 3715 3908 3718 3923
rect 3729 3915 3732 3919
rect 3747 3908 3750 3923
rect 3766 3908 3769 3923
rect 3772 3922 3775 3963
rect 3788 3915 3791 3956
rect 3794 3923 3797 3963
rect 3813 3915 3816 3956
rect 3822 3957 3825 3970
rect 3838 3957 3841 3970
rect 3859 3960 3862 3963
rect 3866 3957 3869 3970
rect 3884 3966 3887 3977
rect 3967 3974 3970 4010
rect 4017 4001 4020 4054
rect 4084 4044 4087 4054
rect 4113 4044 4116 4054
rect 4024 4029 4028 4033
rect 4025 4014 4028 4023
rect 3980 3987 3983 3999
rect 4021 3997 4022 4001
rect 4031 3987 4034 4040
rect 4037 4020 4040 4025
rect 4046 4014 4049 4023
rect 4062 4016 4065 4029
rect 4083 4014 4086 4023
rect 4099 4023 4102 4025
rect 4099 4020 4106 4023
rect 4099 4014 4102 4020
rect 4120 4014 4123 4023
rect 4136 4016 4139 4029
rect 4082 3987 4085 3997
rect 4099 3980 4102 4002
rect 4149 4001 4152 4054
rect 4216 4044 4219 4054
rect 4156 4029 4160 4033
rect 4157 4014 4160 4023
rect 4112 3987 4115 3999
rect 4153 3997 4154 4001
rect 4163 3987 4166 4040
rect 4169 4020 4172 4025
rect 4178 4014 4181 4023
rect 4194 4016 4197 4029
rect 4215 4014 4218 4023
rect 4231 4023 4234 4025
rect 4231 4020 4235 4023
rect 4231 4014 4234 4020
rect 4231 4006 4234 4010
rect 4214 3987 4217 3997
rect 3965 3969 3970 3974
rect 4027 3976 4102 3980
rect 3884 3963 3929 3966
rect 3884 3953 3887 3963
rect 3902 3950 3922 3953
rect 3919 3931 3922 3950
rect 3822 3908 3825 3923
rect 3837 3908 3840 3923
rect 3844 3915 3848 3918
rect 3865 3908 3868 3923
rect 3715 3889 3718 3904
rect 3729 3893 3732 3897
rect 3747 3889 3750 3904
rect 3766 3889 3769 3904
rect 3715 3842 3718 3855
rect 3741 3849 3744 3852
rect 3715 3825 3718 3838
rect 3725 3835 3729 3845
rect 3748 3842 3751 3855
rect 3765 3842 3768 3855
rect 3772 3849 3775 3890
rect 3788 3856 3791 3897
rect 3794 3849 3797 3889
rect 3813 3856 3816 3897
rect 3822 3889 3825 3904
rect 3837 3889 3840 3904
rect 3844 3894 3848 3897
rect 3865 3889 3868 3904
rect 3822 3842 3825 3855
rect 3741 3828 3744 3831
rect 3748 3825 3751 3838
rect 3765 3825 3768 3838
rect 3715 3776 3718 3791
rect 3729 3783 3732 3787
rect 3747 3776 3750 3791
rect 3766 3776 3769 3791
rect 3772 3790 3775 3831
rect 3788 3783 3791 3824
rect 3794 3791 3797 3831
rect 3813 3783 3816 3824
rect 3822 3825 3825 3838
rect 3838 3842 3841 3855
rect 3859 3849 3862 3852
rect 3866 3842 3869 3855
rect 3919 3855 3922 3927
rect 3930 3891 3933 3963
rect 3965 3966 3968 3969
rect 3965 3963 4010 3966
rect 3965 3953 3968 3963
rect 3838 3825 3841 3838
rect 3859 3828 3862 3831
rect 3866 3825 3869 3838
rect 3919 3821 3922 3851
rect 3930 3835 3933 3887
rect 3937 3875 3941 3941
rect 3925 3831 3929 3834
rect 3918 3818 3922 3821
rect 3919 3799 3922 3818
rect 3822 3776 3825 3791
rect 3837 3776 3840 3791
rect 3844 3783 3848 3786
rect 3865 3776 3868 3791
rect 3715 3757 3718 3772
rect 3729 3761 3732 3765
rect 3747 3757 3750 3772
rect 3766 3757 3769 3772
rect 3695 3425 3701 3724
rect 3715 3710 3718 3723
rect 3741 3717 3744 3720
rect 3715 3693 3718 3706
rect 3748 3710 3751 3723
rect 3765 3710 3768 3723
rect 3772 3717 3775 3758
rect 3788 3724 3791 3765
rect 3794 3717 3797 3757
rect 3813 3724 3816 3765
rect 3822 3757 3825 3772
rect 3837 3757 3840 3772
rect 3844 3762 3848 3765
rect 3865 3757 3868 3772
rect 3822 3710 3825 3723
rect 3741 3696 3744 3699
rect 3748 3693 3751 3706
rect 3765 3693 3768 3706
rect 3715 3644 3718 3659
rect 3729 3651 3732 3655
rect 3747 3644 3750 3659
rect 3766 3644 3769 3659
rect 3772 3658 3775 3699
rect 3788 3651 3791 3692
rect 3794 3659 3797 3699
rect 3813 3651 3816 3692
rect 3822 3693 3825 3706
rect 3838 3710 3841 3723
rect 3859 3717 3862 3720
rect 3866 3710 3869 3723
rect 3919 3724 3922 3795
rect 3930 3760 3933 3831
rect 3838 3693 3841 3706
rect 3859 3696 3862 3699
rect 3866 3693 3869 3706
rect 3919 3667 3922 3720
rect 3930 3703 3933 3756
rect 3937 3744 3941 3809
rect 3925 3699 3929 3702
rect 3968 3702 3971 3953
rect 3983 3950 4003 3953
rect 4000 3931 4003 3950
rect 4000 3855 4003 3927
rect 4011 3891 4014 3963
rect 4018 3875 4022 3941
rect 4027 3842 4030 3976
rect 4231 3973 4234 4002
rect 4055 3970 4162 3973
rect 3989 3838 4030 3842
rect 3989 3834 3992 3838
rect 3989 3831 4034 3834
rect 3989 3821 3992 3831
rect 4007 3818 4027 3821
rect 3989 3816 3992 3817
rect 4024 3799 4027 3818
rect 4024 3724 4027 3795
rect 4035 3760 4038 3831
rect 4042 3744 4046 3809
rect 3822 3644 3825 3659
rect 3837 3644 3840 3659
rect 3844 3651 3848 3654
rect 3865 3644 3868 3659
rect 3715 3625 3718 3640
rect 3729 3629 3732 3633
rect 3747 3625 3750 3640
rect 3766 3625 3769 3640
rect 3715 3578 3718 3591
rect 3741 3585 3744 3588
rect 3715 3561 3718 3574
rect 3748 3578 3751 3591
rect 3765 3578 3768 3591
rect 3772 3585 3775 3626
rect 3788 3592 3791 3633
rect 3794 3585 3797 3625
rect 3813 3592 3816 3633
rect 3822 3625 3825 3640
rect 3837 3625 3840 3640
rect 3844 3630 3848 3633
rect 3865 3625 3868 3640
rect 3822 3578 3825 3591
rect 3741 3564 3744 3567
rect 3748 3561 3751 3574
rect 3765 3561 3768 3574
rect 3715 3512 3718 3527
rect 3729 3519 3732 3523
rect 3715 3493 3718 3508
rect 3738 3505 3742 3515
rect 3747 3512 3750 3527
rect 3766 3512 3769 3527
rect 3772 3526 3775 3567
rect 3788 3519 3791 3560
rect 3794 3527 3797 3567
rect 3813 3519 3816 3560
rect 3822 3561 3825 3574
rect 3838 3578 3841 3591
rect 3859 3585 3862 3588
rect 3866 3578 3869 3591
rect 3919 3589 3922 3663
rect 3930 3625 3933 3699
rect 3965 3699 4010 3702
rect 3965 3689 3968 3699
rect 3983 3686 4003 3689
rect 3838 3561 3841 3574
rect 3859 3564 3862 3567
rect 3866 3561 3869 3574
rect 3919 3535 3922 3585
rect 3930 3571 3933 3621
rect 3937 3609 3941 3677
rect 4000 3667 4003 3686
rect 4000 3589 4003 3663
rect 4011 3625 4014 3699
rect 4055 3702 4058 3970
rect 4166 3970 4234 3973
rect 4055 3699 4100 3702
rect 4055 3689 4058 3699
rect 4073 3686 4093 3689
rect 4018 3609 4022 3677
rect 4090 3667 4093 3686
rect 4090 3589 4093 3663
rect 4101 3625 4104 3699
rect 4108 3609 4112 3677
rect 3925 3567 3929 3570
rect 3822 3512 3825 3527
rect 3837 3512 3840 3527
rect 3844 3519 3848 3522
rect 3865 3512 3868 3527
rect 3729 3497 3732 3501
rect 3747 3493 3750 3508
rect 3766 3493 3769 3508
rect 3715 3446 3718 3459
rect 3741 3453 3744 3456
rect 3723 3439 3727 3449
rect 3748 3446 3751 3459
rect 3765 3446 3768 3459
rect 3772 3453 3775 3494
rect 3788 3460 3791 3501
rect 3794 3453 3797 3493
rect 3813 3460 3816 3501
rect 3822 3493 3825 3508
rect 3837 3493 3840 3508
rect 3844 3498 3848 3501
rect 3865 3493 3868 3508
rect 3822 3446 3825 3459
rect 3838 3446 3841 3459
rect 3859 3453 3862 3456
rect 3866 3446 3869 3459
rect 3919 3453 3922 3531
rect 3930 3489 3933 3567
rect 3937 3473 3941 3545
rect 3949 3446 3953 3459
rect 3958 3439 3961 3449
rect 3968 3432 3971 3501
rect 3990 3497 3993 3501
rect 4008 3493 4011 3508
rect 4027 3493 4030 3508
rect 3975 3446 3979 3459
rect 4002 3453 4005 3456
rect 4009 3446 4012 3459
rect 4026 3446 4029 3459
rect 4033 3453 4036 3494
rect 4049 3460 4052 3501
rect 4055 3453 4058 3493
rect 4074 3460 4077 3501
rect 4083 3493 4086 3508
rect 4098 3493 4101 3508
rect 4105 3498 4109 3501
rect 4126 3493 4129 3508
rect 4083 3446 4086 3459
rect 4099 3446 4102 3459
rect 4120 3453 4123 3456
rect 4127 3446 4130 3459
rect 4143 3440 4147 3676
rect 4136 3428 4137 3431
rect 3695 2443 3701 3421
rect 4001 3318 4005 3400
rect 4016 3397 4019 3407
rect 4023 3367 4026 3376
rect 4039 3369 4042 3382
rect 4052 3354 4055 3407
rect 4119 3397 4122 3407
rect 4059 3382 4063 3386
rect 4060 3367 4063 3376
rect 4015 3340 4018 3352
rect 4056 3350 4057 3354
rect 4066 3340 4069 3393
rect 4134 3382 4137 3428
rect 4072 3373 4075 3378
rect 4081 3367 4084 3376
rect 4097 3369 4100 3382
rect 4118 3367 4121 3376
rect 4134 3367 4137 3376
rect 4117 3340 4120 3350
rect 4134 3333 4137 3363
rect 4009 3291 4012 3328
rect 4016 3311 4019 3321
rect 4023 3281 4026 3290
rect 4039 3283 4042 3296
rect 4052 3268 4055 3321
rect 4119 3311 4122 3321
rect 4059 3296 4063 3300
rect 4060 3281 4063 3290
rect 4015 3254 4018 3266
rect 4056 3264 4057 3268
rect 4066 3254 4069 3307
rect 4072 3287 4075 3292
rect 4081 3281 4084 3290
rect 4097 3283 4100 3296
rect 4118 3281 4121 3290
rect 4134 3291 4137 3292
rect 4155 3294 4159 3436
rect 4134 3286 4137 3287
rect 4117 3254 4120 3264
rect 4155 3192 4159 3274
rect 3717 3062 3720 3072
rect 3724 3032 3727 3041
rect 3740 3034 3743 3047
rect 3753 3019 3756 3072
rect 3820 3062 3823 3072
rect 3849 3062 3852 3072
rect 3760 3047 3764 3051
rect 3761 3032 3764 3041
rect 3716 3005 3719 3017
rect 3757 3015 3758 3019
rect 3767 3005 3770 3058
rect 3773 3038 3776 3043
rect 3782 3032 3785 3041
rect 3798 3034 3801 3047
rect 3819 3032 3822 3041
rect 3835 3041 3838 3043
rect 3835 3038 3842 3041
rect 3835 3032 3838 3038
rect 3856 3032 3859 3041
rect 3872 3034 3875 3047
rect 3818 3005 3821 3015
rect 3835 2998 3838 3028
rect 3885 3019 3888 3072
rect 3952 3062 3955 3072
rect 3981 3062 3984 3072
rect 3892 3047 3896 3051
rect 3893 3032 3896 3041
rect 3848 3005 3851 3017
rect 3889 3015 3890 3019
rect 3899 3005 3902 3058
rect 3905 3038 3908 3043
rect 3914 3032 3917 3041
rect 3930 3034 3933 3047
rect 3951 3032 3954 3041
rect 3967 3041 3970 3043
rect 3967 3038 3974 3041
rect 3967 3032 3970 3038
rect 3988 3032 3991 3041
rect 4004 3034 4007 3047
rect 3950 3005 3953 3015
rect 3835 2995 3887 2998
rect 3715 2975 3718 2988
rect 3741 2978 3744 2981
rect 3748 2975 3751 2988
rect 3765 2975 3768 2988
rect 3715 2926 3718 2941
rect 3729 2933 3732 2937
rect 3747 2926 3750 2941
rect 3766 2926 3769 2941
rect 3772 2940 3775 2981
rect 3788 2933 3791 2974
rect 3794 2941 3797 2981
rect 3813 2933 3816 2974
rect 3822 2975 3825 2988
rect 3838 2975 3841 2988
rect 3859 2978 3862 2981
rect 3866 2975 3869 2988
rect 3884 2984 3887 2995
rect 3967 2992 3970 3028
rect 4017 3019 4020 3072
rect 4084 3062 4087 3072
rect 4113 3062 4116 3072
rect 4024 3047 4028 3051
rect 4025 3032 4028 3041
rect 3980 3005 3983 3017
rect 4021 3015 4022 3019
rect 4031 3005 4034 3058
rect 4037 3038 4040 3043
rect 4046 3032 4049 3041
rect 4062 3034 4065 3047
rect 4083 3032 4086 3041
rect 4099 3041 4102 3043
rect 4099 3038 4106 3041
rect 4099 3032 4102 3038
rect 4120 3032 4123 3041
rect 4136 3034 4139 3047
rect 4082 3005 4085 3015
rect 4099 2998 4102 3020
rect 4149 3019 4152 3072
rect 4216 3062 4219 3072
rect 4156 3047 4160 3051
rect 4157 3032 4160 3041
rect 4112 3005 4115 3017
rect 4153 3015 4154 3019
rect 4163 3005 4166 3058
rect 4169 3038 4172 3043
rect 4178 3032 4181 3041
rect 4194 3034 4197 3047
rect 4215 3032 4218 3041
rect 4231 3041 4234 3043
rect 4231 3038 4235 3041
rect 4231 3032 4234 3038
rect 4231 3024 4234 3028
rect 4214 3005 4217 3015
rect 3965 2987 3970 2992
rect 4027 2994 4102 2998
rect 3884 2981 3929 2984
rect 3884 2971 3887 2981
rect 3902 2968 3922 2971
rect 3919 2949 3922 2968
rect 3822 2926 3825 2941
rect 3837 2926 3840 2941
rect 3844 2933 3848 2936
rect 3865 2926 3868 2941
rect 3715 2907 3718 2922
rect 3729 2911 3732 2915
rect 3747 2907 3750 2922
rect 3766 2907 3769 2922
rect 3715 2860 3718 2873
rect 3741 2867 3744 2870
rect 3715 2843 3718 2856
rect 3725 2853 3729 2863
rect 3748 2860 3751 2873
rect 3765 2860 3768 2873
rect 3772 2867 3775 2908
rect 3788 2874 3791 2915
rect 3794 2867 3797 2907
rect 3813 2874 3816 2915
rect 3822 2907 3825 2922
rect 3837 2907 3840 2922
rect 3844 2912 3848 2915
rect 3865 2907 3868 2922
rect 3822 2860 3825 2873
rect 3741 2846 3744 2849
rect 3748 2843 3751 2856
rect 3765 2843 3768 2856
rect 3715 2794 3718 2809
rect 3729 2801 3732 2805
rect 3747 2794 3750 2809
rect 3766 2794 3769 2809
rect 3772 2808 3775 2849
rect 3788 2801 3791 2842
rect 3794 2809 3797 2849
rect 3813 2801 3816 2842
rect 3822 2843 3825 2856
rect 3838 2860 3841 2873
rect 3859 2867 3862 2870
rect 3866 2860 3869 2873
rect 3919 2873 3922 2945
rect 3930 2909 3933 2981
rect 3965 2984 3968 2987
rect 3965 2981 4010 2984
rect 3965 2971 3968 2981
rect 3838 2843 3841 2856
rect 3859 2846 3862 2849
rect 3866 2843 3869 2856
rect 3919 2839 3922 2869
rect 3930 2853 3933 2905
rect 3937 2893 3941 2959
rect 3925 2849 3929 2852
rect 3918 2836 3922 2839
rect 3919 2817 3922 2836
rect 3822 2794 3825 2809
rect 3837 2794 3840 2809
rect 3844 2801 3848 2804
rect 3865 2794 3868 2809
rect 3715 2775 3718 2790
rect 3729 2779 3732 2783
rect 3747 2775 3750 2790
rect 3766 2775 3769 2790
rect 3715 2728 3718 2741
rect 3741 2735 3744 2738
rect 3715 2711 3718 2724
rect 3748 2728 3751 2741
rect 3765 2728 3768 2741
rect 3772 2735 3775 2776
rect 3788 2742 3791 2783
rect 3794 2735 3797 2775
rect 3813 2742 3816 2783
rect 3822 2775 3825 2790
rect 3837 2775 3840 2790
rect 3844 2780 3848 2783
rect 3865 2775 3868 2790
rect 3822 2728 3825 2741
rect 3741 2714 3744 2717
rect 3748 2711 3751 2724
rect 3765 2711 3768 2724
rect 3715 2662 3718 2677
rect 3729 2669 3732 2673
rect 3747 2662 3750 2677
rect 3766 2662 3769 2677
rect 3772 2676 3775 2717
rect 3788 2669 3791 2710
rect 3794 2677 3797 2717
rect 3813 2669 3816 2710
rect 3822 2711 3825 2724
rect 3838 2728 3841 2741
rect 3859 2735 3862 2738
rect 3866 2728 3869 2741
rect 3919 2742 3922 2813
rect 3930 2778 3933 2849
rect 3838 2711 3841 2724
rect 3859 2714 3862 2717
rect 3866 2711 3869 2724
rect 3919 2685 3922 2738
rect 3930 2721 3933 2774
rect 3937 2762 3941 2827
rect 3925 2717 3929 2720
rect 3968 2720 3971 2971
rect 3983 2968 4003 2971
rect 4000 2949 4003 2968
rect 4000 2873 4003 2945
rect 4011 2909 4014 2981
rect 4018 2893 4022 2959
rect 4027 2860 4030 2994
rect 4231 2991 4234 3020
rect 4055 2988 4162 2991
rect 3989 2856 4030 2860
rect 3989 2852 3992 2856
rect 3989 2849 4034 2852
rect 3989 2839 3992 2849
rect 4007 2836 4027 2839
rect 3989 2834 3992 2835
rect 4024 2817 4027 2836
rect 4024 2742 4027 2813
rect 4035 2778 4038 2849
rect 4042 2762 4046 2827
rect 3822 2662 3825 2677
rect 3837 2662 3840 2677
rect 3844 2669 3848 2672
rect 3865 2662 3868 2677
rect 3715 2643 3718 2658
rect 3729 2647 3732 2651
rect 3747 2643 3750 2658
rect 3766 2643 3769 2658
rect 3715 2596 3718 2609
rect 3741 2603 3744 2606
rect 3715 2579 3718 2592
rect 3748 2596 3751 2609
rect 3765 2596 3768 2609
rect 3772 2603 3775 2644
rect 3788 2610 3791 2651
rect 3794 2603 3797 2643
rect 3813 2610 3816 2651
rect 3822 2643 3825 2658
rect 3837 2643 3840 2658
rect 3844 2648 3848 2651
rect 3865 2643 3868 2658
rect 3822 2596 3825 2609
rect 3741 2582 3744 2585
rect 3748 2579 3751 2592
rect 3765 2579 3768 2592
rect 3715 2530 3718 2545
rect 3729 2537 3732 2541
rect 3715 2511 3718 2526
rect 3738 2523 3742 2533
rect 3747 2530 3750 2545
rect 3766 2530 3769 2545
rect 3772 2544 3775 2585
rect 3788 2537 3791 2578
rect 3794 2545 3797 2585
rect 3813 2537 3816 2578
rect 3822 2579 3825 2592
rect 3838 2596 3841 2609
rect 3859 2603 3862 2606
rect 3866 2596 3869 2609
rect 3919 2607 3922 2681
rect 3930 2643 3933 2717
rect 3965 2717 4010 2720
rect 3965 2707 3968 2717
rect 3983 2704 4003 2707
rect 3838 2579 3841 2592
rect 3859 2582 3862 2585
rect 3866 2579 3869 2592
rect 3919 2553 3922 2603
rect 3930 2589 3933 2639
rect 3937 2627 3941 2695
rect 4000 2685 4003 2704
rect 4000 2607 4003 2681
rect 4011 2643 4014 2717
rect 4055 2720 4058 2988
rect 4166 2988 4234 2991
rect 4055 2717 4100 2720
rect 4055 2707 4058 2717
rect 4073 2704 4093 2707
rect 4018 2627 4022 2695
rect 4090 2685 4093 2704
rect 4090 2607 4093 2681
rect 4101 2643 4104 2717
rect 4108 2627 4112 2695
rect 3925 2585 3929 2588
rect 3822 2530 3825 2545
rect 3837 2530 3840 2545
rect 3844 2537 3848 2540
rect 3865 2530 3868 2545
rect 3729 2515 3732 2519
rect 3747 2511 3750 2526
rect 3766 2511 3769 2526
rect 3715 2464 3718 2477
rect 3741 2471 3744 2474
rect 3723 2457 3727 2467
rect 3748 2464 3751 2477
rect 3765 2464 3768 2477
rect 3772 2471 3775 2512
rect 3788 2478 3791 2519
rect 3794 2471 3797 2511
rect 3813 2478 3816 2519
rect 3822 2511 3825 2526
rect 3837 2511 3840 2526
rect 3844 2516 3848 2519
rect 3865 2511 3868 2526
rect 3822 2464 3825 2477
rect 3838 2464 3841 2477
rect 3859 2471 3862 2474
rect 3866 2464 3869 2477
rect 3919 2471 3922 2549
rect 3930 2507 3933 2585
rect 3937 2491 3941 2563
rect 3949 2464 3953 2477
rect 3958 2457 3961 2467
rect 3968 2450 3971 2519
rect 3990 2515 3993 2519
rect 4008 2511 4011 2526
rect 4027 2511 4030 2526
rect 3975 2464 3979 2477
rect 4002 2471 4005 2474
rect 4009 2464 4012 2477
rect 4026 2464 4029 2477
rect 4033 2471 4036 2512
rect 4049 2478 4052 2519
rect 4055 2471 4058 2511
rect 4074 2478 4077 2519
rect 4083 2511 4086 2526
rect 4098 2511 4101 2526
rect 4105 2516 4109 2519
rect 4126 2511 4129 2526
rect 4083 2464 4086 2477
rect 4099 2464 4102 2477
rect 4120 2471 4123 2474
rect 4127 2464 4130 2477
rect 4143 2458 4147 2694
rect 4291 2670 4300 2694
rect 4136 2446 4137 2449
rect 3695 2088 3701 2439
rect 4001 2336 4005 2418
rect 4016 2415 4019 2425
rect 4023 2385 4026 2394
rect 4039 2387 4042 2400
rect 4052 2372 4055 2425
rect 4119 2415 4122 2425
rect 4059 2400 4063 2404
rect 4060 2385 4063 2394
rect 4015 2358 4018 2370
rect 4056 2368 4057 2372
rect 4066 2358 4069 2411
rect 4134 2400 4137 2446
rect 4072 2391 4075 2396
rect 4081 2385 4084 2394
rect 4097 2387 4100 2400
rect 4118 2385 4121 2394
rect 4134 2385 4137 2394
rect 4117 2358 4120 2368
rect 4134 2351 4137 2381
rect 4009 2309 4012 2346
rect 4016 2329 4019 2339
rect 4023 2299 4026 2308
rect 4039 2301 4042 2314
rect 4052 2286 4055 2339
rect 4119 2329 4122 2339
rect 4059 2314 4063 2318
rect 4060 2299 4063 2308
rect 4015 2272 4018 2284
rect 4056 2282 4057 2286
rect 4066 2272 4069 2325
rect 4072 2305 4075 2310
rect 4081 2299 4084 2308
rect 4097 2301 4100 2314
rect 4118 2299 4121 2308
rect 4134 2309 4137 2310
rect 4155 2312 4159 2454
rect 4134 2304 4137 2305
rect 4117 2272 4120 2282
rect 4155 2210 4159 2292
<< m3contact >>
rect 2081 4443 2086 4448
rect 2172 4326 2176 4330
rect 2281 3481 2285 3485
rect 2538 3984 2542 3988
rect 2537 3881 2541 3885
rect 2281 2499 2285 2503
rect 2670 3114 2674 3118
rect 2538 3002 2542 3006
rect 2537 2899 2541 2903
rect 2670 2132 2674 2136
rect 2761 4020 2765 4024
rect 2801 3937 2806 3942
rect 2812 3933 2817 3938
rect 2835 3942 2840 3947
rect 2859 3937 2864 3942
rect 2874 3941 2879 3947
rect 2904 3937 2909 3942
rect 2933 3936 2938 3941
rect 2888 3931 2893 3936
rect 2917 3931 2921 3936
rect 2959 3930 2964 3935
rect 2765 3877 2770 3882
rect 2801 3870 2806 3875
rect 2812 3874 2817 3879
rect 2835 3865 2840 3870
rect 2859 3870 2864 3875
rect 2888 3876 2893 3881
rect 2917 3876 2921 3881
rect 2874 3865 2879 3871
rect 2904 3870 2909 3875
rect 2933 3871 2938 3876
rect 2959 3871 2964 3876
rect 2764 3808 2769 3813
rect 2801 3805 2806 3810
rect 2812 3801 2817 3806
rect 2835 3810 2840 3815
rect 2859 3805 2864 3810
rect 3015 3936 3020 3941
rect 2874 3809 2879 3815
rect 2904 3805 2909 3810
rect 2933 3804 2938 3809
rect 2888 3799 2893 3804
rect 2917 3799 2921 3804
rect 2959 3798 2964 3803
rect 2765 3745 2770 3750
rect 2801 3738 2806 3743
rect 2812 3742 2817 3747
rect 2835 3733 2840 3738
rect 2859 3738 2864 3743
rect 2888 3744 2893 3749
rect 2917 3744 2921 3749
rect 2874 3733 2879 3739
rect 2904 3738 2909 3743
rect 2933 3739 2938 3744
rect 2958 3740 2963 3745
rect 2764 3676 2769 3681
rect 2801 3673 2806 3678
rect 2812 3669 2817 3674
rect 2835 3678 2840 3683
rect 2859 3673 2864 3678
rect 2874 3677 2879 3683
rect 2904 3673 2909 3678
rect 2933 3672 2938 3677
rect 2888 3667 2893 3672
rect 2917 3667 2921 3672
rect 2959 3666 2964 3671
rect 3015 3812 3020 3817
rect 3040 3930 3045 3935
rect 3039 3871 3044 3876
rect 3100 3936 3105 3941
rect 3064 3798 3069 3803
rect 3064 3740 3069 3745
rect 2765 3613 2770 3618
rect 2801 3606 2806 3611
rect 2812 3610 2817 3615
rect 2835 3601 2840 3606
rect 2859 3606 2864 3611
rect 2888 3612 2893 3617
rect 2917 3612 2921 3617
rect 2874 3601 2879 3607
rect 2904 3606 2909 3611
rect 2933 3607 2938 3612
rect 2959 3605 2964 3610
rect 2764 3544 2769 3549
rect 2801 3541 2806 3546
rect 2812 3537 2817 3542
rect 2835 3546 2840 3551
rect 2859 3541 2864 3546
rect 2874 3545 2879 3551
rect 2904 3541 2909 3546
rect 2933 3540 2938 3545
rect 2888 3535 2893 3540
rect 2917 3535 2921 3540
rect 2959 3534 2964 3539
rect 3015 3672 3020 3677
rect 3040 3666 3045 3671
rect 3039 3605 3044 3610
rect 3217 3969 3221 3973
rect 3122 3809 3127 3814
rect 3483 3984 3487 3988
rect 3482 3881 3486 3885
rect 3357 3842 3362 3847
rect 3474 3843 3479 3848
rect 3097 3681 3102 3686
rect 3131 3674 3136 3679
rect 3128 3601 3133 3606
rect 2765 3481 2770 3486
rect 2801 3474 2806 3479
rect 2812 3478 2817 3483
rect 2835 3469 2840 3474
rect 2859 3474 2864 3479
rect 2888 3480 2893 3485
rect 2917 3480 2921 3485
rect 2874 3469 2879 3475
rect 2904 3474 2909 3479
rect 2933 3475 2938 3480
rect 2958 3469 2963 3474
rect 3015 3548 3020 3553
rect 3003 3480 3008 3485
rect 3062 3474 3067 3479
rect 3073 3478 3078 3483
rect 3096 3469 3101 3474
rect 3120 3474 3125 3479
rect 3149 3480 3154 3485
rect 3178 3480 3182 3485
rect 3135 3469 3140 3475
rect 3165 3474 3170 3479
rect 3190 3480 3195 3485
rect 3357 3526 3362 3531
rect 3226 3481 3230 3485
rect 3064 3369 3068 3373
rect 3474 3525 3479 3530
rect 3189 3287 3193 3291
rect 2761 3038 2765 3042
rect 2763 2958 2768 2963
rect 2801 2955 2806 2960
rect 2812 2951 2817 2956
rect 2835 2960 2840 2965
rect 2859 2955 2864 2960
rect 2874 2959 2879 2965
rect 2904 2955 2909 2960
rect 2933 2954 2938 2959
rect 2888 2949 2893 2954
rect 2917 2949 2921 2954
rect 2959 2948 2964 2953
rect 2765 2895 2770 2900
rect 2801 2888 2806 2893
rect 2812 2892 2817 2897
rect 2835 2883 2840 2888
rect 2859 2888 2864 2893
rect 2888 2894 2893 2899
rect 2917 2894 2921 2899
rect 2874 2883 2879 2889
rect 2904 2888 2909 2893
rect 2933 2889 2938 2894
rect 2959 2889 2964 2894
rect 2764 2826 2769 2831
rect 2801 2823 2806 2828
rect 2812 2819 2817 2824
rect 2835 2828 2840 2833
rect 2859 2823 2864 2828
rect 3015 2954 3020 2959
rect 2874 2827 2879 2833
rect 2904 2823 2909 2828
rect 2933 2822 2938 2827
rect 2888 2817 2893 2822
rect 2917 2817 2921 2822
rect 2959 2816 2964 2821
rect 2765 2763 2770 2768
rect 2801 2756 2806 2761
rect 2812 2760 2817 2765
rect 2835 2751 2840 2756
rect 2859 2756 2864 2761
rect 2888 2762 2893 2767
rect 2917 2762 2921 2767
rect 2874 2751 2879 2757
rect 2904 2756 2909 2761
rect 2933 2757 2938 2762
rect 2958 2758 2963 2763
rect 2764 2694 2769 2699
rect 2801 2691 2806 2696
rect 2812 2687 2817 2692
rect 2835 2696 2840 2701
rect 2859 2691 2864 2696
rect 2874 2695 2879 2701
rect 2904 2691 2909 2696
rect 2933 2690 2938 2695
rect 2888 2685 2893 2690
rect 2917 2685 2921 2690
rect 2959 2684 2964 2689
rect 3015 2830 3020 2835
rect 3040 2948 3045 2953
rect 3039 2889 3044 2894
rect 3100 2954 3105 2959
rect 3064 2816 3069 2821
rect 3064 2758 3069 2763
rect 2765 2631 2770 2636
rect 2801 2624 2806 2629
rect 2812 2628 2817 2633
rect 2835 2619 2840 2624
rect 2859 2624 2864 2629
rect 2888 2630 2893 2635
rect 2917 2630 2921 2635
rect 2874 2619 2879 2625
rect 2904 2624 2909 2629
rect 2933 2625 2938 2630
rect 2959 2623 2964 2628
rect 2764 2562 2769 2567
rect 2801 2559 2806 2564
rect 2812 2555 2817 2560
rect 2835 2564 2840 2569
rect 2859 2559 2864 2564
rect 2874 2563 2879 2569
rect 2904 2559 2909 2564
rect 2933 2558 2938 2563
rect 2888 2553 2893 2558
rect 2917 2553 2921 2558
rect 2959 2552 2964 2557
rect 3015 2690 3020 2695
rect 3040 2684 3045 2689
rect 3039 2623 3044 2628
rect 3217 2987 3221 2991
rect 3122 2827 3127 2832
rect 3097 2699 3102 2704
rect 3131 2692 3136 2697
rect 3128 2619 3133 2624
rect 2765 2499 2770 2504
rect 2801 2492 2806 2497
rect 2812 2496 2817 2501
rect 2835 2487 2840 2492
rect 2859 2492 2864 2497
rect 2888 2498 2893 2503
rect 2917 2498 2921 2503
rect 2874 2487 2879 2493
rect 2904 2492 2909 2497
rect 2933 2493 2938 2498
rect 2958 2487 2963 2492
rect 3015 2566 3020 2571
rect 3003 2498 3008 2503
rect 3062 2492 3067 2497
rect 3073 2496 3078 2501
rect 3096 2487 3101 2492
rect 3120 2492 3125 2497
rect 3149 2498 3154 2503
rect 3178 2498 3182 2503
rect 3135 2487 3140 2493
rect 3165 2492 3170 2497
rect 3190 2498 3195 2503
rect 3226 2499 3230 2503
rect 3064 2387 3068 2391
rect 3615 3114 3619 3118
rect 3483 3003 3487 3007
rect 3189 2305 3193 2309
rect 3482 2899 3486 2903
rect 3615 2132 3619 2136
rect 3706 4020 3710 4024
rect 3707 3940 3712 3945
rect 3746 3937 3751 3942
rect 3757 3933 3762 3938
rect 3780 3942 3785 3947
rect 3804 3937 3809 3942
rect 3819 3941 3824 3947
rect 3849 3937 3854 3942
rect 3878 3936 3883 3941
rect 3833 3931 3838 3936
rect 3862 3931 3866 3936
rect 3904 3930 3909 3935
rect 3710 3877 3715 3882
rect 3746 3870 3751 3875
rect 3757 3874 3762 3879
rect 3780 3865 3785 3870
rect 3804 3870 3809 3875
rect 3833 3876 3838 3881
rect 3862 3876 3866 3881
rect 3819 3865 3824 3871
rect 3849 3870 3854 3875
rect 3878 3871 3883 3876
rect 3904 3871 3909 3876
rect 3709 3808 3714 3813
rect 3746 3805 3751 3810
rect 3757 3801 3762 3806
rect 3780 3810 3785 3815
rect 3804 3805 3809 3810
rect 3960 3936 3965 3941
rect 3819 3809 3824 3815
rect 3849 3805 3854 3810
rect 3878 3804 3883 3809
rect 3833 3799 3838 3804
rect 3862 3799 3866 3804
rect 3904 3798 3909 3803
rect 3710 3745 3715 3750
rect 3746 3738 3751 3743
rect 3757 3742 3762 3747
rect 3780 3733 3785 3738
rect 3804 3738 3809 3743
rect 3833 3744 3838 3749
rect 3862 3744 3866 3749
rect 3819 3733 3824 3739
rect 3849 3738 3854 3743
rect 3878 3739 3883 3744
rect 3903 3740 3908 3745
rect 3709 3676 3714 3681
rect 3746 3673 3751 3678
rect 3757 3669 3762 3674
rect 3780 3678 3785 3683
rect 3804 3673 3809 3678
rect 3819 3677 3824 3683
rect 3849 3673 3854 3678
rect 3878 3672 3883 3677
rect 3833 3667 3838 3672
rect 3862 3667 3866 3672
rect 3904 3666 3909 3671
rect 3960 3812 3965 3817
rect 3985 3930 3990 3935
rect 3984 3871 3989 3876
rect 4045 3936 4050 3941
rect 4009 3798 4014 3803
rect 4009 3740 4014 3745
rect 3710 3613 3715 3618
rect 3746 3606 3751 3611
rect 3757 3610 3762 3615
rect 3780 3601 3785 3606
rect 3804 3606 3809 3611
rect 3833 3612 3838 3617
rect 3862 3612 3866 3617
rect 3819 3601 3824 3607
rect 3849 3606 3854 3611
rect 3878 3607 3883 3612
rect 3904 3605 3909 3610
rect 3709 3544 3714 3549
rect 3746 3541 3751 3546
rect 3757 3537 3762 3542
rect 3780 3546 3785 3551
rect 3804 3541 3809 3546
rect 3819 3545 3824 3551
rect 3849 3541 3854 3546
rect 3878 3540 3883 3545
rect 3833 3535 3838 3540
rect 3862 3535 3866 3540
rect 3904 3534 3909 3539
rect 3960 3672 3965 3677
rect 3985 3666 3990 3671
rect 3984 3605 3989 3610
rect 4162 3969 4166 3973
rect 4067 3809 4072 3814
rect 4042 3681 4047 3686
rect 4076 3674 4081 3679
rect 4073 3601 4078 3606
rect 3710 3481 3715 3486
rect 3746 3474 3751 3479
rect 3757 3478 3762 3483
rect 3780 3469 3785 3474
rect 3804 3474 3809 3479
rect 3833 3480 3838 3485
rect 3862 3480 3866 3485
rect 3819 3469 3824 3475
rect 3849 3474 3854 3479
rect 3878 3475 3883 3480
rect 3903 3469 3908 3474
rect 3960 3548 3965 3553
rect 3948 3480 3953 3485
rect 4007 3474 4012 3479
rect 4018 3478 4023 3483
rect 4041 3469 4046 3474
rect 4065 3474 4070 3479
rect 4094 3480 4099 3485
rect 4123 3480 4127 3485
rect 4080 3469 4085 3475
rect 4110 3474 4115 3479
rect 4135 3480 4140 3485
rect 4009 3369 4013 3373
rect 4134 3287 4138 3291
rect 3706 3038 3710 3042
rect 3708 2958 3713 2963
rect 3746 2955 3751 2960
rect 3757 2951 3762 2956
rect 3780 2960 3785 2965
rect 3804 2955 3809 2960
rect 3819 2959 3824 2965
rect 3849 2955 3854 2960
rect 3878 2954 3883 2959
rect 3833 2949 3838 2954
rect 3862 2949 3866 2954
rect 3904 2948 3909 2953
rect 3710 2895 3715 2900
rect 3746 2888 3751 2893
rect 3757 2892 3762 2897
rect 3780 2883 3785 2888
rect 3804 2888 3809 2893
rect 3833 2894 3838 2899
rect 3862 2894 3866 2899
rect 3819 2883 3824 2889
rect 3849 2888 3854 2893
rect 3878 2889 3883 2894
rect 3904 2889 3909 2894
rect 3709 2826 3714 2831
rect 3746 2823 3751 2828
rect 3757 2819 3762 2824
rect 3780 2828 3785 2833
rect 3804 2823 3809 2828
rect 3960 2954 3965 2959
rect 3819 2827 3824 2833
rect 3849 2823 3854 2828
rect 3878 2822 3883 2827
rect 3833 2817 3838 2822
rect 3862 2817 3866 2822
rect 3904 2816 3909 2821
rect 3710 2763 3715 2768
rect 3746 2756 3751 2761
rect 3757 2760 3762 2765
rect 3780 2751 3785 2756
rect 3804 2756 3809 2761
rect 3833 2762 3838 2767
rect 3862 2762 3866 2767
rect 3819 2751 3824 2757
rect 3849 2756 3854 2761
rect 3878 2757 3883 2762
rect 3903 2758 3908 2763
rect 3709 2694 3714 2699
rect 3746 2691 3751 2696
rect 3757 2687 3762 2692
rect 3780 2696 3785 2701
rect 3804 2691 3809 2696
rect 3819 2695 3824 2701
rect 3849 2691 3854 2696
rect 3878 2690 3883 2695
rect 3833 2685 3838 2690
rect 3862 2685 3866 2690
rect 3904 2684 3909 2689
rect 3960 2830 3965 2835
rect 3985 2948 3990 2953
rect 3984 2889 3989 2894
rect 4045 2954 4050 2959
rect 4009 2816 4014 2821
rect 4009 2758 4014 2763
rect 3710 2631 3715 2636
rect 3746 2624 3751 2629
rect 3757 2628 3762 2633
rect 3780 2619 3785 2624
rect 3804 2624 3809 2629
rect 3833 2630 3838 2635
rect 3862 2630 3866 2635
rect 3819 2619 3824 2625
rect 3849 2624 3854 2629
rect 3878 2625 3883 2630
rect 3904 2623 3909 2628
rect 3709 2562 3714 2567
rect 3746 2559 3751 2564
rect 3757 2555 3762 2560
rect 3780 2564 3785 2569
rect 3804 2559 3809 2564
rect 3819 2563 3824 2569
rect 3849 2559 3854 2564
rect 3878 2558 3883 2563
rect 3833 2553 3838 2558
rect 3862 2553 3866 2558
rect 3904 2552 3909 2557
rect 3960 2690 3965 2695
rect 3985 2684 3990 2689
rect 3984 2623 3989 2628
rect 4162 2987 4166 2991
rect 4067 2827 4072 2832
rect 4042 2699 4047 2704
rect 4076 2692 4081 2697
rect 4073 2619 4078 2624
rect 3710 2499 3715 2504
rect 3746 2492 3751 2497
rect 3757 2496 3762 2501
rect 3780 2487 3785 2492
rect 3804 2492 3809 2497
rect 3833 2498 3838 2503
rect 3862 2498 3866 2503
rect 3819 2487 3824 2493
rect 3849 2492 3854 2497
rect 3878 2493 3883 2498
rect 3903 2487 3908 2492
rect 3960 2566 3965 2571
rect 3948 2498 3953 2503
rect 4007 2492 4012 2497
rect 4018 2496 4023 2501
rect 4041 2487 4046 2492
rect 4065 2492 4070 2497
rect 4094 2498 4099 2503
rect 4123 2498 4127 2503
rect 4080 2487 4085 2493
rect 4110 2492 4115 2497
rect 4135 2498 4140 2503
rect 4009 2387 4013 2391
rect 4134 2305 4138 2309
<< metal3 >>
rect 2080 4448 2088 4450
rect 2080 4443 2081 4448
rect 2086 4443 2088 4448
rect 2080 4442 2088 4443
rect 2171 4330 2177 4331
rect 2171 4326 2172 4330
rect 2176 4326 2177 4330
rect 2171 4325 2177 4326
rect 2760 4024 2766 4025
rect 2760 4020 2761 4024
rect 2765 4020 2766 4024
rect 2760 4019 2766 4020
rect 3705 4024 3711 4025
rect 3705 4020 3706 4024
rect 3710 4020 3711 4024
rect 3705 4019 3711 4020
rect 2760 3989 2765 4019
rect 3705 3989 3710 4019
rect 2537 3988 2765 3989
rect 2537 3984 2538 3988
rect 2542 3984 2765 3988
rect 3482 3988 3710 3989
rect 3482 3984 3483 3988
rect 3487 3984 3710 3988
rect 2537 3983 2543 3984
rect 3482 3983 3488 3984
rect 3216 3973 3222 3974
rect 3216 3969 3217 3973
rect 3221 3969 3222 3973
rect 3216 3968 3222 3969
rect 4161 3973 4167 3974
rect 4161 3969 4162 3973
rect 4166 3969 4167 3973
rect 4161 3968 4167 3969
rect 2801 3947 2841 3948
rect 2801 3943 2835 3947
rect 2800 3942 2807 3943
rect 2800 3937 2801 3942
rect 2806 3937 2807 3942
rect 2834 3942 2835 3943
rect 2840 3942 2841 3947
rect 2873 3947 2909 3952
rect 2834 3941 2841 3942
rect 2858 3942 2865 3943
rect 2800 3936 2807 3937
rect 2811 3938 2818 3939
rect 2811 3933 2812 3938
rect 2817 3933 2818 3938
rect 2858 3937 2859 3942
rect 2864 3937 2865 3942
rect 2873 3941 2874 3947
rect 2879 3946 2909 3947
rect 2879 3941 2880 3946
rect 2904 3943 2909 3946
rect 2873 3940 2880 3941
rect 2903 3942 2910 3943
rect 2903 3937 2904 3942
rect 2909 3937 2910 3942
rect 2932 3941 2939 3942
rect 2858 3936 2865 3937
rect 2887 3936 2894 3937
rect 2903 3936 2910 3937
rect 2916 3936 2922 3937
rect 2859 3933 2864 3936
rect 2811 3928 2864 3933
rect 2887 3931 2888 3936
rect 2893 3931 2894 3936
rect 2916 3931 2917 3936
rect 2921 3931 2922 3936
rect 2887 3930 2922 3931
rect 2888 3926 2922 3930
rect 2932 3936 2933 3941
rect 2938 3936 2939 3941
rect 3014 3941 3021 3942
rect 3014 3936 3015 3941
rect 3020 3936 3021 3941
rect 3099 3941 3106 3942
rect 3099 3936 3100 3941
rect 3105 3936 3106 3941
rect 2932 3935 2939 3936
rect 2958 3935 2965 3936
rect 3014 3935 3021 3936
rect 3039 3935 3046 3936
rect 3099 3935 3106 3936
rect 2932 3930 2959 3935
rect 2964 3930 2965 3935
rect 3015 3930 3040 3935
rect 3045 3930 3046 3935
rect 2932 3909 2937 3930
rect 2958 3929 2965 3930
rect 3039 3929 3046 3930
rect 3096 3930 3105 3935
rect 2765 3903 2937 3909
rect 2536 3885 2542 3886
rect 2536 3881 2537 3885
rect 2541 3881 2674 3885
rect 2765 3883 2770 3903
rect 2536 3880 2674 3881
rect 2280 3485 2286 3486
rect 2280 3481 2281 3485
rect 2285 3481 2286 3485
rect 2280 3480 2286 3481
rect 2669 3119 2674 3880
rect 2764 3882 2771 3883
rect 2764 3877 2765 3882
rect 2770 3877 2771 3882
rect 2764 3876 2771 3877
rect 2811 3879 2864 3884
rect 2888 3882 2922 3886
rect 2800 3875 2807 3876
rect 2800 3870 2801 3875
rect 2806 3870 2807 3875
rect 2811 3874 2812 3879
rect 2817 3874 2818 3879
rect 2859 3876 2864 3879
rect 2887 3881 2922 3882
rect 2887 3876 2888 3881
rect 2893 3876 2894 3881
rect 2916 3876 2917 3881
rect 2921 3876 2922 3881
rect 2811 3873 2818 3874
rect 2858 3875 2865 3876
rect 2887 3875 2894 3876
rect 2903 3875 2910 3876
rect 2916 3875 2922 3876
rect 2932 3876 2939 3877
rect 2958 3876 2965 3877
rect 3038 3876 3045 3877
rect 2800 3869 2807 3870
rect 2834 3870 2841 3871
rect 2834 3869 2835 3870
rect 2801 3865 2835 3869
rect 2840 3865 2841 3870
rect 2858 3870 2859 3875
rect 2864 3870 2865 3875
rect 2858 3869 2865 3870
rect 2873 3871 2880 3872
rect 2801 3864 2841 3865
rect 2873 3865 2874 3871
rect 2879 3866 2880 3871
rect 2903 3870 2904 3875
rect 2909 3870 2910 3875
rect 2932 3871 2933 3876
rect 2938 3871 2959 3876
rect 2964 3871 2965 3876
rect 2932 3870 2939 3871
rect 2958 3870 2965 3871
rect 3015 3871 3039 3876
rect 3044 3871 3045 3876
rect 2903 3869 2910 3870
rect 2904 3866 2909 3869
rect 2879 3865 2909 3866
rect 2873 3860 2909 3865
rect 2933 3843 2938 3870
rect 2764 3837 2938 3843
rect 2764 3814 2769 3837
rect 2801 3815 2841 3816
rect 2763 3813 2770 3814
rect 2763 3808 2764 3813
rect 2769 3808 2770 3813
rect 2801 3811 2835 3815
rect 2763 3807 2770 3808
rect 2800 3810 2807 3811
rect 2800 3805 2801 3810
rect 2806 3805 2807 3810
rect 2834 3810 2835 3811
rect 2840 3810 2841 3815
rect 2873 3815 2909 3820
rect 3015 3818 3020 3871
rect 3038 3870 3045 3871
rect 3096 3842 3101 3930
rect 3058 3837 3101 3842
rect 2834 3809 2841 3810
rect 2858 3810 2865 3811
rect 2800 3804 2807 3805
rect 2811 3806 2818 3807
rect 2811 3801 2812 3806
rect 2817 3801 2818 3806
rect 2858 3805 2859 3810
rect 2864 3805 2865 3810
rect 2873 3809 2874 3815
rect 2879 3814 2909 3815
rect 2879 3809 2880 3814
rect 2904 3811 2909 3814
rect 3014 3817 3021 3818
rect 3014 3812 3015 3817
rect 3020 3812 3021 3817
rect 3014 3811 3021 3812
rect 2873 3808 2880 3809
rect 2903 3810 2910 3811
rect 2903 3805 2904 3810
rect 2909 3805 2910 3810
rect 2932 3809 2939 3810
rect 2858 3804 2865 3805
rect 2887 3804 2894 3805
rect 2903 3804 2910 3805
rect 2916 3804 2922 3805
rect 2859 3801 2864 3804
rect 2811 3796 2864 3801
rect 2887 3799 2888 3804
rect 2893 3799 2894 3804
rect 2916 3799 2917 3804
rect 2921 3799 2922 3804
rect 2887 3798 2922 3799
rect 2888 3794 2922 3798
rect 2932 3804 2933 3809
rect 2938 3804 2939 3809
rect 3058 3804 3063 3837
rect 3121 3814 3128 3815
rect 3121 3809 3122 3814
rect 3127 3809 3128 3814
rect 3121 3808 3128 3809
rect 2932 3803 2939 3804
rect 2958 3803 2965 3804
rect 2932 3798 2959 3803
rect 2964 3798 2965 3803
rect 3058 3803 3070 3804
rect 3058 3798 3064 3803
rect 3069 3798 3070 3803
rect 2932 3777 2937 3798
rect 2958 3797 2965 3798
rect 3063 3797 3070 3798
rect 2765 3771 2937 3777
rect 2765 3751 2770 3771
rect 2764 3750 2771 3751
rect 2764 3745 2765 3750
rect 2770 3745 2771 3750
rect 2764 3744 2771 3745
rect 2811 3747 2864 3752
rect 2888 3750 2922 3754
rect 2800 3743 2807 3744
rect 2800 3738 2801 3743
rect 2806 3738 2807 3743
rect 2811 3742 2812 3747
rect 2817 3742 2818 3747
rect 2859 3744 2864 3747
rect 2887 3749 2922 3750
rect 2887 3744 2888 3749
rect 2893 3744 2894 3749
rect 2916 3744 2917 3749
rect 2921 3744 2922 3749
rect 2957 3745 2964 3746
rect 3063 3745 3070 3746
rect 2811 3741 2818 3742
rect 2858 3743 2865 3744
rect 2887 3743 2894 3744
rect 2903 3743 2910 3744
rect 2916 3743 2922 3744
rect 2932 3744 2958 3745
rect 2800 3737 2807 3738
rect 2834 3738 2841 3739
rect 2834 3737 2835 3738
rect 2801 3733 2835 3737
rect 2840 3733 2841 3738
rect 2858 3738 2859 3743
rect 2864 3738 2865 3743
rect 2858 3737 2865 3738
rect 2873 3739 2880 3740
rect 2801 3732 2841 3733
rect 2873 3733 2874 3739
rect 2879 3734 2880 3739
rect 2903 3738 2904 3743
rect 2909 3738 2910 3743
rect 2903 3737 2910 3738
rect 2932 3739 2933 3744
rect 2938 3740 2958 3744
rect 2963 3740 2964 3745
rect 2938 3739 2939 3740
rect 2957 3739 2964 3740
rect 3059 3740 3064 3745
rect 3069 3740 3070 3745
rect 3059 3739 3070 3740
rect 2932 3738 2939 3739
rect 2904 3734 2909 3737
rect 2879 3733 2909 3734
rect 2873 3728 2909 3733
rect 2932 3711 2937 3738
rect 2764 3705 2937 3711
rect 3059 3711 3064 3739
rect 3059 3706 3102 3711
rect 2764 3682 2769 3705
rect 2801 3683 2841 3684
rect 2763 3681 2770 3682
rect 2763 3676 2764 3681
rect 2769 3676 2770 3681
rect 2801 3679 2835 3683
rect 2763 3675 2770 3676
rect 2800 3678 2807 3679
rect 2800 3673 2801 3678
rect 2806 3673 2807 3678
rect 2834 3678 2835 3679
rect 2840 3678 2841 3683
rect 2873 3683 2909 3688
rect 3097 3687 3102 3706
rect 2834 3677 2841 3678
rect 2858 3678 2865 3679
rect 2800 3672 2807 3673
rect 2811 3674 2818 3675
rect 2811 3669 2812 3674
rect 2817 3669 2818 3674
rect 2858 3673 2859 3678
rect 2864 3673 2865 3678
rect 2873 3677 2874 3683
rect 2879 3682 2909 3683
rect 2879 3677 2880 3682
rect 2904 3679 2909 3682
rect 3096 3686 3103 3687
rect 3096 3681 3097 3686
rect 3102 3681 3103 3686
rect 3096 3680 3103 3681
rect 3122 3679 3127 3808
rect 3130 3679 3137 3680
rect 2873 3676 2880 3677
rect 2903 3678 2910 3679
rect 2903 3673 2904 3678
rect 2909 3673 2910 3678
rect 2932 3677 2939 3678
rect 2858 3672 2865 3673
rect 2887 3672 2894 3673
rect 2903 3672 2910 3673
rect 2916 3672 2922 3673
rect 2859 3669 2864 3672
rect 2811 3664 2864 3669
rect 2887 3667 2888 3672
rect 2893 3667 2894 3672
rect 2916 3667 2917 3672
rect 2921 3667 2922 3672
rect 2887 3666 2922 3667
rect 2888 3662 2922 3666
rect 2932 3672 2933 3677
rect 2938 3672 2939 3677
rect 3014 3677 3021 3678
rect 3014 3672 3015 3677
rect 3020 3672 3021 3677
rect 3110 3674 3131 3679
rect 3136 3674 3137 3679
rect 3110 3673 3122 3674
rect 3130 3673 3137 3674
rect 2932 3671 2939 3672
rect 2958 3671 2965 3672
rect 3014 3671 3021 3672
rect 3039 3671 3046 3672
rect 2932 3666 2959 3671
rect 2964 3666 2965 3671
rect 3015 3666 3040 3671
rect 3045 3666 3046 3671
rect 2932 3645 2937 3666
rect 2958 3665 2965 3666
rect 3039 3665 3046 3666
rect 3110 3665 3115 3673
rect 2765 3639 2937 3645
rect 3077 3644 3115 3665
rect 2765 3619 2770 3639
rect 2764 3618 2771 3619
rect 2764 3613 2765 3618
rect 2770 3613 2771 3618
rect 2764 3612 2771 3613
rect 2811 3615 2864 3620
rect 2888 3618 2922 3622
rect 2800 3611 2807 3612
rect 2800 3606 2801 3611
rect 2806 3606 2807 3611
rect 2811 3610 2812 3615
rect 2817 3610 2818 3615
rect 2859 3612 2864 3615
rect 2887 3617 2922 3618
rect 2887 3612 2888 3617
rect 2893 3612 2894 3617
rect 2916 3612 2917 3617
rect 2921 3612 2922 3617
rect 2811 3609 2818 3610
rect 2858 3611 2865 3612
rect 2887 3611 2894 3612
rect 2903 3611 2910 3612
rect 2916 3611 2922 3612
rect 2932 3612 2939 3613
rect 2800 3605 2807 3606
rect 2834 3606 2841 3607
rect 2834 3605 2835 3606
rect 2801 3601 2835 3605
rect 2840 3601 2841 3606
rect 2858 3606 2859 3611
rect 2864 3606 2865 3611
rect 2858 3605 2865 3606
rect 2873 3607 2880 3608
rect 2801 3600 2841 3601
rect 2873 3601 2874 3607
rect 2879 3602 2880 3607
rect 2903 3606 2904 3611
rect 2909 3606 2910 3611
rect 2932 3607 2933 3612
rect 2938 3610 2939 3612
rect 2958 3610 2965 3611
rect 3038 3610 3045 3611
rect 2938 3607 2959 3610
rect 2932 3606 2959 3607
rect 2903 3605 2910 3606
rect 2933 3605 2959 3606
rect 2964 3605 2965 3610
rect 2904 3602 2909 3605
rect 2879 3601 2909 3602
rect 2873 3596 2909 3601
rect 2933 3579 2938 3605
rect 2958 3604 2965 3605
rect 3015 3605 3039 3610
rect 3044 3605 3045 3610
rect 2764 3573 2938 3579
rect 2764 3550 2769 3573
rect 2801 3551 2841 3552
rect 2763 3549 2770 3550
rect 2763 3544 2764 3549
rect 2769 3544 2770 3549
rect 2801 3547 2835 3551
rect 2763 3543 2770 3544
rect 2800 3546 2807 3547
rect 2800 3541 2801 3546
rect 2806 3541 2807 3546
rect 2834 3546 2835 3547
rect 2840 3546 2841 3551
rect 2873 3551 2909 3556
rect 3015 3554 3020 3605
rect 3038 3604 3045 3605
rect 2834 3545 2841 3546
rect 2858 3546 2865 3547
rect 2800 3540 2807 3541
rect 2811 3542 2818 3543
rect 2811 3537 2812 3542
rect 2817 3537 2818 3542
rect 2858 3541 2859 3546
rect 2864 3541 2865 3546
rect 2873 3545 2874 3551
rect 2879 3550 2909 3551
rect 2879 3545 2880 3550
rect 2904 3547 2909 3550
rect 3014 3553 3021 3554
rect 3014 3548 3015 3553
rect 3020 3548 3021 3553
rect 3014 3547 3021 3548
rect 2873 3544 2880 3545
rect 2903 3546 2910 3547
rect 2903 3541 2904 3546
rect 2909 3541 2910 3546
rect 2932 3545 2939 3546
rect 2858 3540 2865 3541
rect 2887 3540 2894 3541
rect 2903 3540 2910 3541
rect 2916 3540 2922 3541
rect 2859 3537 2864 3540
rect 2811 3532 2864 3537
rect 2887 3535 2888 3540
rect 2893 3535 2894 3540
rect 2916 3535 2917 3540
rect 2921 3535 2922 3540
rect 2887 3534 2922 3535
rect 2888 3530 2922 3534
rect 2932 3540 2933 3545
rect 2938 3540 2939 3545
rect 2932 3539 2939 3540
rect 2958 3539 2965 3540
rect 2932 3534 2959 3539
rect 2964 3534 2965 3539
rect 3077 3535 3082 3644
rect 3127 3606 3134 3607
rect 3127 3601 3128 3606
rect 3133 3601 3134 3606
rect 3127 3600 3134 3601
rect 3034 3534 3082 3535
rect 2932 3513 2937 3534
rect 2958 3533 2965 3534
rect 2765 3507 2937 3513
rect 3003 3529 3082 3534
rect 3128 3538 3133 3600
rect 3128 3532 3195 3538
rect 2765 3487 2770 3507
rect 2764 3486 2771 3487
rect 2764 3481 2765 3486
rect 2770 3481 2771 3486
rect 2764 3480 2771 3481
rect 2811 3483 2864 3488
rect 2888 3486 2922 3490
rect 3003 3486 3008 3529
rect 2800 3479 2807 3480
rect 2800 3474 2801 3479
rect 2806 3474 2807 3479
rect 2811 3478 2812 3483
rect 2817 3478 2818 3483
rect 2859 3480 2864 3483
rect 2887 3485 2922 3486
rect 2887 3480 2888 3485
rect 2893 3480 2894 3485
rect 2916 3480 2917 3485
rect 2921 3480 2922 3485
rect 3002 3485 3009 3486
rect 2811 3477 2818 3478
rect 2858 3479 2865 3480
rect 2887 3479 2894 3480
rect 2903 3479 2910 3480
rect 2916 3479 2922 3480
rect 2932 3480 2939 3481
rect 2800 3473 2807 3474
rect 2834 3474 2841 3475
rect 2834 3473 2835 3474
rect 2801 3469 2835 3473
rect 2840 3469 2841 3474
rect 2858 3474 2859 3479
rect 2864 3474 2865 3479
rect 2858 3473 2865 3474
rect 2873 3475 2880 3476
rect 2801 3468 2841 3469
rect 2873 3469 2874 3475
rect 2879 3470 2880 3475
rect 2903 3474 2904 3479
rect 2909 3474 2910 3479
rect 2932 3475 2933 3480
rect 2938 3475 2939 3480
rect 3002 3480 3003 3485
rect 3008 3480 3009 3485
rect 3072 3483 3125 3488
rect 3149 3486 3183 3490
rect 3190 3486 3195 3532
rect 3002 3479 3009 3480
rect 3061 3479 3068 3480
rect 2932 3474 2939 3475
rect 2957 3474 2964 3475
rect 2903 3473 2910 3474
rect 2904 3470 2909 3473
rect 2879 3469 2909 3470
rect 2873 3464 2909 3469
rect 2934 3469 2958 3474
rect 2963 3469 2964 3474
rect 3061 3474 3062 3479
rect 3067 3474 3068 3479
rect 3072 3478 3073 3483
rect 3078 3478 3079 3483
rect 3120 3480 3125 3483
rect 3148 3485 3183 3486
rect 3148 3480 3149 3485
rect 3154 3480 3155 3485
rect 3177 3480 3178 3485
rect 3182 3480 3183 3485
rect 3072 3477 3079 3478
rect 3119 3479 3126 3480
rect 3148 3479 3155 3480
rect 3164 3479 3171 3480
rect 3177 3479 3183 3480
rect 3189 3485 3196 3486
rect 3189 3480 3190 3485
rect 3195 3480 3196 3485
rect 3189 3479 3196 3480
rect 3061 3473 3068 3474
rect 3095 3474 3102 3475
rect 3095 3473 3096 3474
rect 2669 3118 2675 3119
rect 2669 3114 2670 3118
rect 2674 3114 2675 3118
rect 2669 3113 2675 3114
rect 2934 3101 2939 3469
rect 2957 3468 2964 3469
rect 3062 3469 3096 3473
rect 3101 3469 3102 3474
rect 3119 3474 3120 3479
rect 3125 3474 3126 3479
rect 3119 3473 3126 3474
rect 3134 3475 3141 3476
rect 3062 3468 3102 3469
rect 3134 3469 3135 3475
rect 3140 3470 3141 3475
rect 3164 3474 3165 3479
rect 3170 3474 3171 3479
rect 3164 3473 3171 3474
rect 3165 3470 3170 3473
rect 3140 3469 3170 3470
rect 3134 3464 3170 3469
rect 3217 3441 3222 3968
rect 3746 3947 3786 3948
rect 3706 3945 3713 3946
rect 3684 3940 3707 3945
rect 3712 3940 3713 3945
rect 3746 3943 3780 3947
rect 3481 3885 3487 3886
rect 3481 3881 3482 3885
rect 3486 3881 3619 3885
rect 3481 3880 3619 3881
rect 3473 3848 3480 3849
rect 3356 3847 3363 3848
rect 3356 3842 3357 3847
rect 3362 3842 3363 3847
rect 3473 3843 3474 3848
rect 3479 3843 3480 3848
rect 3473 3842 3480 3843
rect 3356 3841 3363 3842
rect 3357 3532 3362 3841
rect 3356 3531 3363 3532
rect 3474 3531 3479 3842
rect 3356 3526 3357 3531
rect 3362 3526 3363 3531
rect 3356 3525 3363 3526
rect 3473 3530 3480 3531
rect 3473 3525 3474 3530
rect 3479 3525 3480 3530
rect 3473 3524 3480 3525
rect 3225 3485 3231 3486
rect 3225 3481 3226 3485
rect 3230 3481 3231 3485
rect 3225 3480 3231 3481
rect 3064 3436 3222 3441
rect 3064 3374 3069 3436
rect 3063 3373 3069 3374
rect 3063 3369 3064 3373
rect 3068 3369 3069 3373
rect 3063 3368 3069 3369
rect 3226 3311 3231 3480
rect 3189 3306 3231 3311
rect 3189 3292 3194 3306
rect 3188 3291 3194 3292
rect 3188 3287 3189 3291
rect 3193 3287 3194 3291
rect 3188 3286 3194 3287
rect 3614 3119 3619 3880
rect 3614 3118 3620 3119
rect 3614 3114 3615 3118
rect 3619 3114 3620 3118
rect 3614 3113 3620 3114
rect 3684 3101 3689 3940
rect 3706 3939 3713 3940
rect 3745 3942 3752 3943
rect 3745 3937 3746 3942
rect 3751 3937 3752 3942
rect 3779 3942 3780 3943
rect 3785 3942 3786 3947
rect 3818 3947 3854 3952
rect 3779 3941 3786 3942
rect 3803 3942 3810 3943
rect 3745 3936 3752 3937
rect 3756 3938 3763 3939
rect 3756 3933 3757 3938
rect 3762 3933 3763 3938
rect 3803 3937 3804 3942
rect 3809 3937 3810 3942
rect 3818 3941 3819 3947
rect 3824 3946 3854 3947
rect 3824 3941 3825 3946
rect 3849 3943 3854 3946
rect 3818 3940 3825 3941
rect 3848 3942 3855 3943
rect 3848 3937 3849 3942
rect 3854 3937 3855 3942
rect 3877 3941 3884 3942
rect 3803 3936 3810 3937
rect 3832 3936 3839 3937
rect 3848 3936 3855 3937
rect 3861 3936 3867 3937
rect 3804 3933 3809 3936
rect 3756 3928 3809 3933
rect 3832 3931 3833 3936
rect 3838 3931 3839 3936
rect 3861 3931 3862 3936
rect 3866 3931 3867 3936
rect 3832 3930 3867 3931
rect 3833 3926 3867 3930
rect 3877 3936 3878 3941
rect 3883 3936 3884 3941
rect 3959 3941 3966 3942
rect 3959 3936 3960 3941
rect 3965 3936 3966 3941
rect 4044 3941 4051 3942
rect 4044 3936 4045 3941
rect 4050 3936 4051 3941
rect 3877 3935 3884 3936
rect 3903 3935 3910 3936
rect 3959 3935 3966 3936
rect 3984 3935 3991 3936
rect 4044 3935 4051 3936
rect 3877 3930 3904 3935
rect 3909 3930 3910 3935
rect 3960 3930 3985 3935
rect 3990 3930 3991 3935
rect 3877 3909 3882 3930
rect 3903 3929 3910 3930
rect 3984 3929 3991 3930
rect 4041 3930 4050 3935
rect 3710 3903 3882 3909
rect 3710 3883 3715 3903
rect 3709 3882 3716 3883
rect 3709 3877 3710 3882
rect 3715 3877 3716 3882
rect 3709 3876 3716 3877
rect 3756 3879 3809 3884
rect 3833 3882 3867 3886
rect 3745 3875 3752 3876
rect 3745 3870 3746 3875
rect 3751 3870 3752 3875
rect 3756 3874 3757 3879
rect 3762 3874 3763 3879
rect 3804 3876 3809 3879
rect 3832 3881 3867 3882
rect 3832 3876 3833 3881
rect 3838 3876 3839 3881
rect 3861 3876 3862 3881
rect 3866 3876 3867 3881
rect 3756 3873 3763 3874
rect 3803 3875 3810 3876
rect 3832 3875 3839 3876
rect 3848 3875 3855 3876
rect 3861 3875 3867 3876
rect 3877 3876 3884 3877
rect 3903 3876 3910 3877
rect 3983 3876 3990 3877
rect 3745 3869 3752 3870
rect 3779 3870 3786 3871
rect 3779 3869 3780 3870
rect 3746 3865 3780 3869
rect 3785 3865 3786 3870
rect 3803 3870 3804 3875
rect 3809 3870 3810 3875
rect 3803 3869 3810 3870
rect 3818 3871 3825 3872
rect 3746 3864 3786 3865
rect 3818 3865 3819 3871
rect 3824 3866 3825 3871
rect 3848 3870 3849 3875
rect 3854 3870 3855 3875
rect 3877 3871 3878 3876
rect 3883 3871 3904 3876
rect 3909 3871 3910 3876
rect 3877 3870 3884 3871
rect 3903 3870 3910 3871
rect 3960 3871 3984 3876
rect 3989 3871 3990 3876
rect 3848 3869 3855 3870
rect 3849 3866 3854 3869
rect 3824 3865 3854 3866
rect 3818 3860 3854 3865
rect 3878 3843 3883 3870
rect 3709 3837 3883 3843
rect 3709 3814 3714 3837
rect 3746 3815 3786 3816
rect 3708 3813 3715 3814
rect 3708 3808 3709 3813
rect 3714 3808 3715 3813
rect 3746 3811 3780 3815
rect 3708 3807 3715 3808
rect 3745 3810 3752 3811
rect 3745 3805 3746 3810
rect 3751 3805 3752 3810
rect 3779 3810 3780 3811
rect 3785 3810 3786 3815
rect 3818 3815 3854 3820
rect 3960 3818 3965 3871
rect 3983 3870 3990 3871
rect 4041 3842 4046 3930
rect 4003 3837 4046 3842
rect 3779 3809 3786 3810
rect 3803 3810 3810 3811
rect 3745 3804 3752 3805
rect 3756 3806 3763 3807
rect 3756 3801 3757 3806
rect 3762 3801 3763 3806
rect 3803 3805 3804 3810
rect 3809 3805 3810 3810
rect 3818 3809 3819 3815
rect 3824 3814 3854 3815
rect 3824 3809 3825 3814
rect 3849 3811 3854 3814
rect 3959 3817 3966 3818
rect 3959 3812 3960 3817
rect 3965 3812 3966 3817
rect 3959 3811 3966 3812
rect 3818 3808 3825 3809
rect 3848 3810 3855 3811
rect 3848 3805 3849 3810
rect 3854 3805 3855 3810
rect 3877 3809 3884 3810
rect 3803 3804 3810 3805
rect 3832 3804 3839 3805
rect 3848 3804 3855 3805
rect 3861 3804 3867 3805
rect 3804 3801 3809 3804
rect 3756 3796 3809 3801
rect 3832 3799 3833 3804
rect 3838 3799 3839 3804
rect 3861 3799 3862 3804
rect 3866 3799 3867 3804
rect 3832 3798 3867 3799
rect 3833 3794 3867 3798
rect 3877 3804 3878 3809
rect 3883 3804 3884 3809
rect 4003 3804 4008 3837
rect 4066 3814 4073 3815
rect 4066 3809 4067 3814
rect 4072 3809 4073 3814
rect 4066 3808 4073 3809
rect 3877 3803 3884 3804
rect 3903 3803 3910 3804
rect 3877 3798 3904 3803
rect 3909 3798 3910 3803
rect 4003 3803 4015 3804
rect 4003 3798 4009 3803
rect 4014 3798 4015 3803
rect 3877 3777 3882 3798
rect 3903 3797 3910 3798
rect 4008 3797 4015 3798
rect 3710 3771 3882 3777
rect 3710 3751 3715 3771
rect 3709 3750 3716 3751
rect 3709 3745 3710 3750
rect 3715 3745 3716 3750
rect 3709 3744 3716 3745
rect 3756 3747 3809 3752
rect 3833 3750 3867 3754
rect 3745 3743 3752 3744
rect 3745 3738 3746 3743
rect 3751 3738 3752 3743
rect 3756 3742 3757 3747
rect 3762 3742 3763 3747
rect 3804 3744 3809 3747
rect 3832 3749 3867 3750
rect 3832 3744 3833 3749
rect 3838 3744 3839 3749
rect 3861 3744 3862 3749
rect 3866 3744 3867 3749
rect 3902 3745 3909 3746
rect 4008 3745 4015 3746
rect 3756 3741 3763 3742
rect 3803 3743 3810 3744
rect 3832 3743 3839 3744
rect 3848 3743 3855 3744
rect 3861 3743 3867 3744
rect 3877 3744 3903 3745
rect 3745 3737 3752 3738
rect 3779 3738 3786 3739
rect 3779 3737 3780 3738
rect 3746 3733 3780 3737
rect 3785 3733 3786 3738
rect 3803 3738 3804 3743
rect 3809 3738 3810 3743
rect 3803 3737 3810 3738
rect 3818 3739 3825 3740
rect 3746 3732 3786 3733
rect 3818 3733 3819 3739
rect 3824 3734 3825 3739
rect 3848 3738 3849 3743
rect 3854 3738 3855 3743
rect 3848 3737 3855 3738
rect 3877 3739 3878 3744
rect 3883 3740 3903 3744
rect 3908 3740 3909 3745
rect 3883 3739 3884 3740
rect 3902 3739 3909 3740
rect 4004 3740 4009 3745
rect 4014 3740 4015 3745
rect 4004 3739 4015 3740
rect 3877 3738 3884 3739
rect 3849 3734 3854 3737
rect 3824 3733 3854 3734
rect 3818 3728 3854 3733
rect 3877 3711 3882 3738
rect 3709 3705 3882 3711
rect 4004 3711 4009 3739
rect 4004 3706 4047 3711
rect 3709 3682 3714 3705
rect 3746 3683 3786 3684
rect 3708 3681 3715 3682
rect 3708 3676 3709 3681
rect 3714 3676 3715 3681
rect 3746 3679 3780 3683
rect 3708 3675 3715 3676
rect 3745 3678 3752 3679
rect 3745 3673 3746 3678
rect 3751 3673 3752 3678
rect 3779 3678 3780 3679
rect 3785 3678 3786 3683
rect 3818 3683 3854 3688
rect 4042 3687 4047 3706
rect 3779 3677 3786 3678
rect 3803 3678 3810 3679
rect 3745 3672 3752 3673
rect 3756 3674 3763 3675
rect 3756 3669 3757 3674
rect 3762 3669 3763 3674
rect 3803 3673 3804 3678
rect 3809 3673 3810 3678
rect 3818 3677 3819 3683
rect 3824 3682 3854 3683
rect 3824 3677 3825 3682
rect 3849 3679 3854 3682
rect 4041 3686 4048 3687
rect 4041 3681 4042 3686
rect 4047 3681 4048 3686
rect 4041 3680 4048 3681
rect 4067 3679 4072 3808
rect 4075 3679 4082 3680
rect 3818 3676 3825 3677
rect 3848 3678 3855 3679
rect 3848 3673 3849 3678
rect 3854 3673 3855 3678
rect 3877 3677 3884 3678
rect 3803 3672 3810 3673
rect 3832 3672 3839 3673
rect 3848 3672 3855 3673
rect 3861 3672 3867 3673
rect 3804 3669 3809 3672
rect 3756 3664 3809 3669
rect 3832 3667 3833 3672
rect 3838 3667 3839 3672
rect 3861 3667 3862 3672
rect 3866 3667 3867 3672
rect 3832 3666 3867 3667
rect 3833 3662 3867 3666
rect 3877 3672 3878 3677
rect 3883 3672 3884 3677
rect 3959 3677 3966 3678
rect 3959 3672 3960 3677
rect 3965 3672 3966 3677
rect 4055 3674 4076 3679
rect 4081 3674 4082 3679
rect 4055 3673 4067 3674
rect 4075 3673 4082 3674
rect 3877 3671 3884 3672
rect 3903 3671 3910 3672
rect 3959 3671 3966 3672
rect 3984 3671 3991 3672
rect 3877 3666 3904 3671
rect 3909 3666 3910 3671
rect 3960 3666 3985 3671
rect 3990 3666 3991 3671
rect 3877 3645 3882 3666
rect 3903 3665 3910 3666
rect 3984 3665 3991 3666
rect 4055 3665 4060 3673
rect 3710 3639 3882 3645
rect 4022 3644 4060 3665
rect 3710 3619 3715 3639
rect 3709 3618 3716 3619
rect 3709 3613 3710 3618
rect 3715 3613 3716 3618
rect 3709 3612 3716 3613
rect 3756 3615 3809 3620
rect 3833 3618 3867 3622
rect 3745 3611 3752 3612
rect 3745 3606 3746 3611
rect 3751 3606 3752 3611
rect 3756 3610 3757 3615
rect 3762 3610 3763 3615
rect 3804 3612 3809 3615
rect 3832 3617 3867 3618
rect 3832 3612 3833 3617
rect 3838 3612 3839 3617
rect 3861 3612 3862 3617
rect 3866 3612 3867 3617
rect 3756 3609 3763 3610
rect 3803 3611 3810 3612
rect 3832 3611 3839 3612
rect 3848 3611 3855 3612
rect 3861 3611 3867 3612
rect 3877 3612 3884 3613
rect 3745 3605 3752 3606
rect 3779 3606 3786 3607
rect 3779 3605 3780 3606
rect 3746 3601 3780 3605
rect 3785 3601 3786 3606
rect 3803 3606 3804 3611
rect 3809 3606 3810 3611
rect 3803 3605 3810 3606
rect 3818 3607 3825 3608
rect 3746 3600 3786 3601
rect 3818 3601 3819 3607
rect 3824 3602 3825 3607
rect 3848 3606 3849 3611
rect 3854 3606 3855 3611
rect 3877 3607 3878 3612
rect 3883 3610 3884 3612
rect 3903 3610 3910 3611
rect 3983 3610 3990 3611
rect 3883 3607 3904 3610
rect 3877 3606 3904 3607
rect 3848 3605 3855 3606
rect 3878 3605 3904 3606
rect 3909 3605 3910 3610
rect 3849 3602 3854 3605
rect 3824 3601 3854 3602
rect 3818 3596 3854 3601
rect 3878 3579 3883 3605
rect 3903 3604 3910 3605
rect 3960 3605 3984 3610
rect 3989 3605 3990 3610
rect 3709 3573 3883 3579
rect 3709 3550 3714 3573
rect 3746 3551 3786 3552
rect 3708 3549 3715 3550
rect 3708 3544 3709 3549
rect 3714 3544 3715 3549
rect 3746 3547 3780 3551
rect 3708 3543 3715 3544
rect 3745 3546 3752 3547
rect 3745 3541 3746 3546
rect 3751 3541 3752 3546
rect 3779 3546 3780 3547
rect 3785 3546 3786 3551
rect 3818 3551 3854 3556
rect 3960 3554 3965 3605
rect 3983 3604 3990 3605
rect 3779 3545 3786 3546
rect 3803 3546 3810 3547
rect 3745 3540 3752 3541
rect 3756 3542 3763 3543
rect 3756 3537 3757 3542
rect 3762 3537 3763 3542
rect 3803 3541 3804 3546
rect 3809 3541 3810 3546
rect 3818 3545 3819 3551
rect 3824 3550 3854 3551
rect 3824 3545 3825 3550
rect 3849 3547 3854 3550
rect 3959 3553 3966 3554
rect 3959 3548 3960 3553
rect 3965 3548 3966 3553
rect 3959 3547 3966 3548
rect 3818 3544 3825 3545
rect 3848 3546 3855 3547
rect 3848 3541 3849 3546
rect 3854 3541 3855 3546
rect 3877 3545 3884 3546
rect 3803 3540 3810 3541
rect 3832 3540 3839 3541
rect 3848 3540 3855 3541
rect 3861 3540 3867 3541
rect 3804 3537 3809 3540
rect 3756 3532 3809 3537
rect 3832 3535 3833 3540
rect 3838 3535 3839 3540
rect 3861 3535 3862 3540
rect 3866 3535 3867 3540
rect 3832 3534 3867 3535
rect 3833 3530 3867 3534
rect 3877 3540 3878 3545
rect 3883 3540 3884 3545
rect 3877 3539 3884 3540
rect 3903 3539 3910 3540
rect 3877 3534 3904 3539
rect 3909 3534 3910 3539
rect 4022 3535 4027 3644
rect 4072 3606 4079 3607
rect 4072 3601 4073 3606
rect 4078 3601 4079 3606
rect 4072 3600 4079 3601
rect 3979 3534 4027 3535
rect 3877 3513 3882 3534
rect 3903 3533 3910 3534
rect 3710 3507 3882 3513
rect 3948 3529 4027 3534
rect 4073 3538 4078 3600
rect 4073 3532 4140 3538
rect 3710 3487 3715 3507
rect 3709 3486 3716 3487
rect 3709 3481 3710 3486
rect 3715 3481 3716 3486
rect 3709 3480 3716 3481
rect 3756 3483 3809 3488
rect 3833 3486 3867 3490
rect 3948 3486 3953 3529
rect 3745 3479 3752 3480
rect 3745 3474 3746 3479
rect 3751 3474 3752 3479
rect 3756 3478 3757 3483
rect 3762 3478 3763 3483
rect 3804 3480 3809 3483
rect 3832 3485 3867 3486
rect 3832 3480 3833 3485
rect 3838 3480 3839 3485
rect 3861 3480 3862 3485
rect 3866 3480 3867 3485
rect 3947 3485 3954 3486
rect 3756 3477 3763 3478
rect 3803 3479 3810 3480
rect 3832 3479 3839 3480
rect 3848 3479 3855 3480
rect 3861 3479 3867 3480
rect 3877 3480 3884 3481
rect 3745 3473 3752 3474
rect 3779 3474 3786 3475
rect 3779 3473 3780 3474
rect 3746 3469 3780 3473
rect 3785 3469 3786 3474
rect 3803 3474 3804 3479
rect 3809 3474 3810 3479
rect 3803 3473 3810 3474
rect 3818 3475 3825 3476
rect 3746 3468 3786 3469
rect 3818 3469 3819 3475
rect 3824 3470 3825 3475
rect 3848 3474 3849 3479
rect 3854 3474 3855 3479
rect 3877 3475 3878 3480
rect 3883 3475 3884 3480
rect 3947 3480 3948 3485
rect 3953 3480 3954 3485
rect 4017 3483 4070 3488
rect 4094 3486 4128 3490
rect 4135 3486 4140 3532
rect 3947 3479 3954 3480
rect 4006 3479 4013 3480
rect 3877 3474 3884 3475
rect 3902 3474 3909 3475
rect 3848 3473 3855 3474
rect 3849 3470 3854 3473
rect 3824 3469 3854 3470
rect 3818 3464 3854 3469
rect 3879 3469 3903 3474
rect 3908 3469 3909 3474
rect 4006 3474 4007 3479
rect 4012 3474 4013 3479
rect 4017 3478 4018 3483
rect 4023 3478 4024 3483
rect 4065 3480 4070 3483
rect 4093 3485 4128 3486
rect 4093 3480 4094 3485
rect 4099 3480 4100 3485
rect 4122 3480 4123 3485
rect 4127 3480 4128 3485
rect 4017 3477 4024 3478
rect 4064 3479 4071 3480
rect 4093 3479 4100 3480
rect 4109 3479 4116 3480
rect 4122 3479 4128 3480
rect 4134 3485 4141 3486
rect 4134 3480 4135 3485
rect 4140 3480 4141 3485
rect 4134 3479 4141 3480
rect 4006 3473 4013 3474
rect 4040 3474 4047 3475
rect 4040 3473 4041 3474
rect 3879 3338 3884 3469
rect 3902 3468 3909 3469
rect 4007 3469 4041 3473
rect 4046 3469 4047 3474
rect 4064 3474 4065 3479
rect 4070 3474 4071 3479
rect 4064 3473 4071 3474
rect 4079 3475 4086 3476
rect 4007 3468 4047 3469
rect 4079 3469 4080 3475
rect 4085 3470 4086 3475
rect 4109 3474 4110 3479
rect 4115 3474 4116 3479
rect 4109 3473 4116 3474
rect 4110 3470 4115 3473
rect 4085 3469 4115 3470
rect 4079 3464 4115 3469
rect 4162 3441 4167 3968
rect 4009 3436 4167 3441
rect 4009 3374 4014 3436
rect 4008 3373 4014 3374
rect 4008 3369 4009 3373
rect 4013 3369 4014 3373
rect 4008 3368 4014 3369
rect 3879 3332 4190 3338
rect 4133 3291 4139 3292
rect 4133 3287 4134 3291
rect 4138 3287 4139 3291
rect 4133 3286 4139 3287
rect 2934 3095 3689 3101
rect 4134 3082 4139 3286
rect 2281 3077 4139 3082
rect 2281 2504 2286 3077
rect 2675 3042 2766 3043
rect 2675 3038 2761 3042
rect 2765 3038 2766 3042
rect 2676 3007 2681 3038
rect 2760 3037 2766 3038
rect 3705 3042 3711 3043
rect 3705 3038 3706 3042
rect 3710 3038 3711 3042
rect 3705 3037 3711 3038
rect 2537 3006 2681 3007
rect 2537 3002 2538 3006
rect 2542 3002 2681 3006
rect 3482 3007 3488 3008
rect 3705 3007 3710 3037
rect 2537 3001 2543 3002
rect 2763 2999 3243 3004
rect 3482 3003 3483 3007
rect 3487 3003 3710 3007
rect 4185 3004 4190 3332
rect 3482 3002 3710 3003
rect 3848 2999 4190 3004
rect 2763 2964 2768 2999
rect 3238 2994 3876 2999
rect 3216 2991 3222 2992
rect 3216 2987 3217 2991
rect 3221 2987 3222 2991
rect 3216 2986 3222 2987
rect 4161 2991 4167 2992
rect 4161 2987 4162 2991
rect 4166 2987 4167 2991
rect 4161 2986 4167 2987
rect 2801 2965 2841 2966
rect 2762 2963 2769 2964
rect 2762 2958 2763 2963
rect 2768 2958 2769 2963
rect 2801 2961 2835 2965
rect 2762 2957 2769 2958
rect 2800 2960 2807 2961
rect 2800 2955 2801 2960
rect 2806 2955 2807 2960
rect 2834 2960 2835 2961
rect 2840 2960 2841 2965
rect 2873 2965 2909 2970
rect 2834 2959 2841 2960
rect 2858 2960 2865 2961
rect 2800 2954 2807 2955
rect 2811 2956 2818 2957
rect 2811 2951 2812 2956
rect 2817 2951 2818 2956
rect 2858 2955 2859 2960
rect 2864 2955 2865 2960
rect 2873 2959 2874 2965
rect 2879 2964 2909 2965
rect 2879 2959 2880 2964
rect 2904 2961 2909 2964
rect 2873 2958 2880 2959
rect 2903 2960 2910 2961
rect 2903 2955 2904 2960
rect 2909 2955 2910 2960
rect 2932 2959 2939 2960
rect 2858 2954 2865 2955
rect 2887 2954 2894 2955
rect 2903 2954 2910 2955
rect 2916 2954 2922 2955
rect 2859 2951 2864 2954
rect 2811 2946 2864 2951
rect 2887 2949 2888 2954
rect 2893 2949 2894 2954
rect 2916 2949 2917 2954
rect 2921 2949 2922 2954
rect 2887 2948 2922 2949
rect 2888 2944 2922 2948
rect 2932 2954 2933 2959
rect 2938 2954 2939 2959
rect 3014 2959 3021 2960
rect 3014 2954 3015 2959
rect 3020 2954 3021 2959
rect 3099 2959 3106 2960
rect 3099 2954 3100 2959
rect 3105 2954 3106 2959
rect 2932 2953 2939 2954
rect 2958 2953 2965 2954
rect 3014 2953 3021 2954
rect 3039 2953 3046 2954
rect 3099 2953 3106 2954
rect 2932 2948 2959 2953
rect 2964 2948 2965 2953
rect 3015 2948 3040 2953
rect 3045 2948 3046 2953
rect 2932 2927 2937 2948
rect 2958 2947 2965 2948
rect 3039 2947 3046 2948
rect 3096 2948 3105 2953
rect 2765 2921 2937 2927
rect 2536 2903 2542 2904
rect 2536 2899 2537 2903
rect 2541 2899 2674 2903
rect 2765 2901 2770 2921
rect 2536 2898 2674 2899
rect 2280 2503 2286 2504
rect 2280 2499 2281 2503
rect 2285 2499 2286 2503
rect 2280 2498 2286 2499
rect 2669 2137 2674 2898
rect 2764 2900 2771 2901
rect 2764 2895 2765 2900
rect 2770 2895 2771 2900
rect 2764 2894 2771 2895
rect 2811 2897 2864 2902
rect 2888 2900 2922 2904
rect 2800 2893 2807 2894
rect 2800 2888 2801 2893
rect 2806 2888 2807 2893
rect 2811 2892 2812 2897
rect 2817 2892 2818 2897
rect 2859 2894 2864 2897
rect 2887 2899 2922 2900
rect 2887 2894 2888 2899
rect 2893 2894 2894 2899
rect 2916 2894 2917 2899
rect 2921 2894 2922 2899
rect 2811 2891 2818 2892
rect 2858 2893 2865 2894
rect 2887 2893 2894 2894
rect 2903 2893 2910 2894
rect 2916 2893 2922 2894
rect 2932 2894 2939 2895
rect 2958 2894 2965 2895
rect 3038 2894 3045 2895
rect 2800 2887 2807 2888
rect 2834 2888 2841 2889
rect 2834 2887 2835 2888
rect 2801 2883 2835 2887
rect 2840 2883 2841 2888
rect 2858 2888 2859 2893
rect 2864 2888 2865 2893
rect 2858 2887 2865 2888
rect 2873 2889 2880 2890
rect 2801 2882 2841 2883
rect 2873 2883 2874 2889
rect 2879 2884 2880 2889
rect 2903 2888 2904 2893
rect 2909 2888 2910 2893
rect 2932 2889 2933 2894
rect 2938 2889 2959 2894
rect 2964 2889 2965 2894
rect 2932 2888 2939 2889
rect 2958 2888 2965 2889
rect 3015 2889 3039 2894
rect 3044 2889 3045 2894
rect 2903 2887 2910 2888
rect 2904 2884 2909 2887
rect 2879 2883 2909 2884
rect 2873 2878 2909 2883
rect 2933 2861 2938 2888
rect 2764 2855 2938 2861
rect 2764 2832 2769 2855
rect 2801 2833 2841 2834
rect 2763 2831 2770 2832
rect 2763 2826 2764 2831
rect 2769 2826 2770 2831
rect 2801 2829 2835 2833
rect 2763 2825 2770 2826
rect 2800 2828 2807 2829
rect 2800 2823 2801 2828
rect 2806 2823 2807 2828
rect 2834 2828 2835 2829
rect 2840 2828 2841 2833
rect 2873 2833 2909 2838
rect 3015 2836 3020 2889
rect 3038 2888 3045 2889
rect 3096 2860 3101 2948
rect 3058 2855 3101 2860
rect 2834 2827 2841 2828
rect 2858 2828 2865 2829
rect 2800 2822 2807 2823
rect 2811 2824 2818 2825
rect 2811 2819 2812 2824
rect 2817 2819 2818 2824
rect 2858 2823 2859 2828
rect 2864 2823 2865 2828
rect 2873 2827 2874 2833
rect 2879 2832 2909 2833
rect 2879 2827 2880 2832
rect 2904 2829 2909 2832
rect 3014 2835 3021 2836
rect 3014 2830 3015 2835
rect 3020 2830 3021 2835
rect 3014 2829 3021 2830
rect 2873 2826 2880 2827
rect 2903 2828 2910 2829
rect 2903 2823 2904 2828
rect 2909 2823 2910 2828
rect 2932 2827 2939 2828
rect 2858 2822 2865 2823
rect 2887 2822 2894 2823
rect 2903 2822 2910 2823
rect 2916 2822 2922 2823
rect 2859 2819 2864 2822
rect 2811 2814 2864 2819
rect 2887 2817 2888 2822
rect 2893 2817 2894 2822
rect 2916 2817 2917 2822
rect 2921 2817 2922 2822
rect 2887 2816 2922 2817
rect 2888 2812 2922 2816
rect 2932 2822 2933 2827
rect 2938 2822 2939 2827
rect 3058 2822 3063 2855
rect 3121 2832 3128 2833
rect 3121 2827 3122 2832
rect 3127 2827 3128 2832
rect 3121 2826 3128 2827
rect 2932 2821 2939 2822
rect 2958 2821 2965 2822
rect 2932 2816 2959 2821
rect 2964 2816 2965 2821
rect 3058 2821 3070 2822
rect 3058 2816 3064 2821
rect 3069 2816 3070 2821
rect 2932 2795 2937 2816
rect 2958 2815 2965 2816
rect 3063 2815 3070 2816
rect 2765 2789 2937 2795
rect 2765 2769 2770 2789
rect 2764 2768 2771 2769
rect 2764 2763 2765 2768
rect 2770 2763 2771 2768
rect 2764 2762 2771 2763
rect 2811 2765 2864 2770
rect 2888 2768 2922 2772
rect 2800 2761 2807 2762
rect 2800 2756 2801 2761
rect 2806 2756 2807 2761
rect 2811 2760 2812 2765
rect 2817 2760 2818 2765
rect 2859 2762 2864 2765
rect 2887 2767 2922 2768
rect 2887 2762 2888 2767
rect 2893 2762 2894 2767
rect 2916 2762 2917 2767
rect 2921 2762 2922 2767
rect 2957 2763 2964 2764
rect 3063 2763 3070 2764
rect 2811 2759 2818 2760
rect 2858 2761 2865 2762
rect 2887 2761 2894 2762
rect 2903 2761 2910 2762
rect 2916 2761 2922 2762
rect 2932 2762 2958 2763
rect 2800 2755 2807 2756
rect 2834 2756 2841 2757
rect 2834 2755 2835 2756
rect 2801 2751 2835 2755
rect 2840 2751 2841 2756
rect 2858 2756 2859 2761
rect 2864 2756 2865 2761
rect 2858 2755 2865 2756
rect 2873 2757 2880 2758
rect 2801 2750 2841 2751
rect 2873 2751 2874 2757
rect 2879 2752 2880 2757
rect 2903 2756 2904 2761
rect 2909 2756 2910 2761
rect 2903 2755 2910 2756
rect 2932 2757 2933 2762
rect 2938 2758 2958 2762
rect 2963 2758 2964 2763
rect 2938 2757 2939 2758
rect 2957 2757 2964 2758
rect 3059 2758 3064 2763
rect 3069 2758 3070 2763
rect 3059 2757 3070 2758
rect 2932 2756 2939 2757
rect 2904 2752 2909 2755
rect 2879 2751 2909 2752
rect 2873 2746 2909 2751
rect 2932 2729 2937 2756
rect 2764 2723 2937 2729
rect 3059 2729 3064 2757
rect 3059 2724 3102 2729
rect 2764 2700 2769 2723
rect 2801 2701 2841 2702
rect 2763 2699 2770 2700
rect 2763 2694 2764 2699
rect 2769 2694 2770 2699
rect 2801 2697 2835 2701
rect 2763 2693 2770 2694
rect 2800 2696 2807 2697
rect 2800 2691 2801 2696
rect 2806 2691 2807 2696
rect 2834 2696 2835 2697
rect 2840 2696 2841 2701
rect 2873 2701 2909 2706
rect 3097 2705 3102 2724
rect 2834 2695 2841 2696
rect 2858 2696 2865 2697
rect 2800 2690 2807 2691
rect 2811 2692 2818 2693
rect 2811 2687 2812 2692
rect 2817 2687 2818 2692
rect 2858 2691 2859 2696
rect 2864 2691 2865 2696
rect 2873 2695 2874 2701
rect 2879 2700 2909 2701
rect 2879 2695 2880 2700
rect 2904 2697 2909 2700
rect 3096 2704 3103 2705
rect 3096 2699 3097 2704
rect 3102 2699 3103 2704
rect 3096 2698 3103 2699
rect 3122 2697 3127 2826
rect 3130 2697 3137 2698
rect 2873 2694 2880 2695
rect 2903 2696 2910 2697
rect 2903 2691 2904 2696
rect 2909 2691 2910 2696
rect 2932 2695 2939 2696
rect 2858 2690 2865 2691
rect 2887 2690 2894 2691
rect 2903 2690 2910 2691
rect 2916 2690 2922 2691
rect 2859 2687 2864 2690
rect 2811 2682 2864 2687
rect 2887 2685 2888 2690
rect 2893 2685 2894 2690
rect 2916 2685 2917 2690
rect 2921 2685 2922 2690
rect 2887 2684 2922 2685
rect 2888 2680 2922 2684
rect 2932 2690 2933 2695
rect 2938 2690 2939 2695
rect 3014 2695 3021 2696
rect 3014 2690 3015 2695
rect 3020 2690 3021 2695
rect 3110 2692 3131 2697
rect 3136 2692 3137 2697
rect 3110 2691 3122 2692
rect 3130 2691 3137 2692
rect 2932 2689 2939 2690
rect 2958 2689 2965 2690
rect 3014 2689 3021 2690
rect 3039 2689 3046 2690
rect 2932 2684 2959 2689
rect 2964 2684 2965 2689
rect 3015 2684 3040 2689
rect 3045 2684 3046 2689
rect 2932 2663 2937 2684
rect 2958 2683 2965 2684
rect 3039 2683 3046 2684
rect 3110 2683 3115 2691
rect 2765 2657 2937 2663
rect 3077 2662 3115 2683
rect 2765 2637 2770 2657
rect 2764 2636 2771 2637
rect 2764 2631 2765 2636
rect 2770 2631 2771 2636
rect 2764 2630 2771 2631
rect 2811 2633 2864 2638
rect 2888 2636 2922 2640
rect 2800 2629 2807 2630
rect 2800 2624 2801 2629
rect 2806 2624 2807 2629
rect 2811 2628 2812 2633
rect 2817 2628 2818 2633
rect 2859 2630 2864 2633
rect 2887 2635 2922 2636
rect 2887 2630 2888 2635
rect 2893 2630 2894 2635
rect 2916 2630 2917 2635
rect 2921 2630 2922 2635
rect 2811 2627 2818 2628
rect 2858 2629 2865 2630
rect 2887 2629 2894 2630
rect 2903 2629 2910 2630
rect 2916 2629 2922 2630
rect 2932 2630 2939 2631
rect 2800 2623 2807 2624
rect 2834 2624 2841 2625
rect 2834 2623 2835 2624
rect 2801 2619 2835 2623
rect 2840 2619 2841 2624
rect 2858 2624 2859 2629
rect 2864 2624 2865 2629
rect 2858 2623 2865 2624
rect 2873 2625 2880 2626
rect 2801 2618 2841 2619
rect 2873 2619 2874 2625
rect 2879 2620 2880 2625
rect 2903 2624 2904 2629
rect 2909 2624 2910 2629
rect 2932 2625 2933 2630
rect 2938 2628 2939 2630
rect 2958 2628 2965 2629
rect 3038 2628 3045 2629
rect 2938 2625 2959 2628
rect 2932 2624 2959 2625
rect 2903 2623 2910 2624
rect 2933 2623 2959 2624
rect 2964 2623 2965 2628
rect 2904 2620 2909 2623
rect 2879 2619 2909 2620
rect 2873 2614 2909 2619
rect 2933 2597 2938 2623
rect 2958 2622 2965 2623
rect 3015 2623 3039 2628
rect 3044 2623 3045 2628
rect 2764 2591 2938 2597
rect 2764 2568 2769 2591
rect 2801 2569 2841 2570
rect 2763 2567 2770 2568
rect 2763 2562 2764 2567
rect 2769 2562 2770 2567
rect 2801 2565 2835 2569
rect 2763 2561 2770 2562
rect 2800 2564 2807 2565
rect 2800 2559 2801 2564
rect 2806 2559 2807 2564
rect 2834 2564 2835 2565
rect 2840 2564 2841 2569
rect 2873 2569 2909 2574
rect 3015 2572 3020 2623
rect 3038 2622 3045 2623
rect 2834 2563 2841 2564
rect 2858 2564 2865 2565
rect 2800 2558 2807 2559
rect 2811 2560 2818 2561
rect 2811 2555 2812 2560
rect 2817 2555 2818 2560
rect 2858 2559 2859 2564
rect 2864 2559 2865 2564
rect 2873 2563 2874 2569
rect 2879 2568 2909 2569
rect 2879 2563 2880 2568
rect 2904 2565 2909 2568
rect 3014 2571 3021 2572
rect 3014 2566 3015 2571
rect 3020 2566 3021 2571
rect 3014 2565 3021 2566
rect 2873 2562 2880 2563
rect 2903 2564 2910 2565
rect 2903 2559 2904 2564
rect 2909 2559 2910 2564
rect 2932 2563 2939 2564
rect 2858 2558 2865 2559
rect 2887 2558 2894 2559
rect 2903 2558 2910 2559
rect 2916 2558 2922 2559
rect 2859 2555 2864 2558
rect 2811 2550 2864 2555
rect 2887 2553 2888 2558
rect 2893 2553 2894 2558
rect 2916 2553 2917 2558
rect 2921 2553 2922 2558
rect 2887 2552 2922 2553
rect 2888 2548 2922 2552
rect 2932 2558 2933 2563
rect 2938 2558 2939 2563
rect 2932 2557 2939 2558
rect 2958 2557 2965 2558
rect 2932 2552 2959 2557
rect 2964 2552 2965 2557
rect 3077 2553 3082 2662
rect 3127 2624 3134 2625
rect 3127 2619 3128 2624
rect 3133 2619 3134 2624
rect 3127 2618 3134 2619
rect 3034 2552 3082 2553
rect 2932 2531 2937 2552
rect 2958 2551 2965 2552
rect 2765 2525 2937 2531
rect 3003 2547 3082 2552
rect 3128 2556 3133 2618
rect 3128 2550 3195 2556
rect 2765 2505 2770 2525
rect 2764 2504 2771 2505
rect 2764 2499 2765 2504
rect 2770 2499 2771 2504
rect 2764 2498 2771 2499
rect 2811 2501 2864 2506
rect 2888 2504 2922 2508
rect 3003 2504 3008 2547
rect 2800 2497 2807 2498
rect 2800 2492 2801 2497
rect 2806 2492 2807 2497
rect 2811 2496 2812 2501
rect 2817 2496 2818 2501
rect 2859 2498 2864 2501
rect 2887 2503 2922 2504
rect 2887 2498 2888 2503
rect 2893 2498 2894 2503
rect 2916 2498 2917 2503
rect 2921 2498 2922 2503
rect 3002 2503 3009 2504
rect 2811 2495 2818 2496
rect 2858 2497 2865 2498
rect 2887 2497 2894 2498
rect 2903 2497 2910 2498
rect 2916 2497 2922 2498
rect 2932 2498 2939 2499
rect 2800 2491 2807 2492
rect 2834 2492 2841 2493
rect 2834 2491 2835 2492
rect 2801 2487 2835 2491
rect 2840 2487 2841 2492
rect 2858 2492 2859 2497
rect 2864 2492 2865 2497
rect 2858 2491 2865 2492
rect 2873 2493 2880 2494
rect 2801 2486 2841 2487
rect 2873 2487 2874 2493
rect 2879 2488 2880 2493
rect 2903 2492 2904 2497
rect 2909 2492 2910 2497
rect 2932 2493 2933 2498
rect 2938 2493 2939 2498
rect 3002 2498 3003 2503
rect 3008 2498 3009 2503
rect 3072 2501 3125 2506
rect 3149 2504 3183 2508
rect 3190 2504 3195 2550
rect 3002 2497 3009 2498
rect 3061 2497 3068 2498
rect 2932 2492 2939 2493
rect 2957 2492 2964 2493
rect 2903 2491 2910 2492
rect 2904 2488 2909 2491
rect 2879 2487 2909 2488
rect 2873 2482 2909 2487
rect 2934 2487 2958 2492
rect 2963 2487 2964 2492
rect 3061 2492 3062 2497
rect 3067 2492 3068 2497
rect 3072 2496 3073 2501
rect 3078 2496 3079 2501
rect 3120 2498 3125 2501
rect 3148 2503 3183 2504
rect 3148 2498 3149 2503
rect 3154 2498 3155 2503
rect 3177 2498 3178 2503
rect 3182 2498 3183 2503
rect 3072 2495 3079 2496
rect 3119 2497 3126 2498
rect 3148 2497 3155 2498
rect 3164 2497 3171 2498
rect 3177 2497 3183 2498
rect 3189 2503 3196 2504
rect 3189 2498 3190 2503
rect 3195 2498 3196 2503
rect 3189 2497 3196 2498
rect 3061 2491 3068 2492
rect 3095 2492 3102 2493
rect 3095 2491 3096 2492
rect 2669 2136 2675 2137
rect 2669 2132 2670 2136
rect 2674 2132 2675 2136
rect 2669 2131 2675 2132
rect 2934 2134 2939 2487
rect 2957 2486 2964 2487
rect 3062 2487 3096 2491
rect 3101 2487 3102 2492
rect 3119 2492 3120 2497
rect 3125 2492 3126 2497
rect 3119 2491 3126 2492
rect 3134 2493 3141 2494
rect 3062 2486 3102 2487
rect 3134 2487 3135 2493
rect 3140 2488 3141 2493
rect 3164 2492 3165 2497
rect 3170 2492 3171 2497
rect 3164 2491 3171 2492
rect 3165 2488 3170 2491
rect 3140 2487 3170 2488
rect 3134 2482 3170 2487
rect 3217 2459 3222 2986
rect 3746 2965 3786 2966
rect 3707 2963 3714 2964
rect 3684 2958 3708 2963
rect 3713 2958 3714 2963
rect 3746 2961 3780 2965
rect 3481 2903 3487 2904
rect 3481 2899 3482 2903
rect 3486 2899 3619 2903
rect 3481 2898 3619 2899
rect 3225 2503 3231 2504
rect 3225 2499 3226 2503
rect 3230 2499 3231 2503
rect 3225 2498 3231 2499
rect 3064 2454 3222 2459
rect 3064 2392 3069 2454
rect 3063 2391 3069 2392
rect 3063 2387 3064 2391
rect 3068 2387 3069 2391
rect 3063 2386 3069 2387
rect 3226 2329 3231 2498
rect 3189 2324 3231 2329
rect 3189 2310 3194 2324
rect 3188 2309 3194 2310
rect 3188 2305 3189 2309
rect 3193 2305 3194 2309
rect 3188 2304 3194 2305
rect 3614 2137 3619 2898
rect 3614 2136 3620 2137
rect 2934 2129 2979 2134
rect 3614 2132 3615 2136
rect 3619 2132 3620 2136
rect 3614 2131 3620 2132
rect 3684 2125 3689 2958
rect 3707 2957 3714 2958
rect 3745 2960 3752 2961
rect 3745 2955 3746 2960
rect 3751 2955 3752 2960
rect 3779 2960 3780 2961
rect 3785 2960 3786 2965
rect 3818 2965 3854 2970
rect 3779 2959 3786 2960
rect 3803 2960 3810 2961
rect 3745 2954 3752 2955
rect 3756 2956 3763 2957
rect 3756 2951 3757 2956
rect 3762 2951 3763 2956
rect 3803 2955 3804 2960
rect 3809 2955 3810 2960
rect 3818 2959 3819 2965
rect 3824 2964 3854 2965
rect 3824 2959 3825 2964
rect 3849 2961 3854 2964
rect 3818 2958 3825 2959
rect 3848 2960 3855 2961
rect 3848 2955 3849 2960
rect 3854 2955 3855 2960
rect 3877 2959 3884 2960
rect 3803 2954 3810 2955
rect 3832 2954 3839 2955
rect 3848 2954 3855 2955
rect 3861 2954 3867 2955
rect 3804 2951 3809 2954
rect 3756 2946 3809 2951
rect 3832 2949 3833 2954
rect 3838 2949 3839 2954
rect 3861 2949 3862 2954
rect 3866 2949 3867 2954
rect 3832 2948 3867 2949
rect 3833 2944 3867 2948
rect 3877 2954 3878 2959
rect 3883 2954 3884 2959
rect 3959 2959 3966 2960
rect 3959 2954 3960 2959
rect 3965 2954 3966 2959
rect 4044 2959 4051 2960
rect 4044 2954 4045 2959
rect 4050 2954 4051 2959
rect 3877 2953 3884 2954
rect 3903 2953 3910 2954
rect 3959 2953 3966 2954
rect 3984 2953 3991 2954
rect 4044 2953 4051 2954
rect 3877 2948 3904 2953
rect 3909 2948 3910 2953
rect 3960 2948 3985 2953
rect 3990 2948 3991 2953
rect 3877 2927 3882 2948
rect 3903 2947 3910 2948
rect 3984 2947 3991 2948
rect 4041 2948 4050 2953
rect 3710 2921 3882 2927
rect 3710 2901 3715 2921
rect 3709 2900 3716 2901
rect 3709 2895 3710 2900
rect 3715 2895 3716 2900
rect 3709 2894 3716 2895
rect 3756 2897 3809 2902
rect 3833 2900 3867 2904
rect 3745 2893 3752 2894
rect 3745 2888 3746 2893
rect 3751 2888 3752 2893
rect 3756 2892 3757 2897
rect 3762 2892 3763 2897
rect 3804 2894 3809 2897
rect 3832 2899 3867 2900
rect 3832 2894 3833 2899
rect 3838 2894 3839 2899
rect 3861 2894 3862 2899
rect 3866 2894 3867 2899
rect 3756 2891 3763 2892
rect 3803 2893 3810 2894
rect 3832 2893 3839 2894
rect 3848 2893 3855 2894
rect 3861 2893 3867 2894
rect 3877 2894 3884 2895
rect 3903 2894 3910 2895
rect 3983 2894 3990 2895
rect 3745 2887 3752 2888
rect 3779 2888 3786 2889
rect 3779 2887 3780 2888
rect 3746 2883 3780 2887
rect 3785 2883 3786 2888
rect 3803 2888 3804 2893
rect 3809 2888 3810 2893
rect 3803 2887 3810 2888
rect 3818 2889 3825 2890
rect 3746 2882 3786 2883
rect 3818 2883 3819 2889
rect 3824 2884 3825 2889
rect 3848 2888 3849 2893
rect 3854 2888 3855 2893
rect 3877 2889 3878 2894
rect 3883 2889 3904 2894
rect 3909 2889 3910 2894
rect 3877 2888 3884 2889
rect 3903 2888 3910 2889
rect 3960 2889 3984 2894
rect 3989 2889 3990 2894
rect 3848 2887 3855 2888
rect 3849 2884 3854 2887
rect 3824 2883 3854 2884
rect 3818 2878 3854 2883
rect 3878 2861 3883 2888
rect 3709 2855 3883 2861
rect 3709 2832 3714 2855
rect 3746 2833 3786 2834
rect 3708 2831 3715 2832
rect 3708 2826 3709 2831
rect 3714 2826 3715 2831
rect 3746 2829 3780 2833
rect 3708 2825 3715 2826
rect 3745 2828 3752 2829
rect 3745 2823 3746 2828
rect 3751 2823 3752 2828
rect 3779 2828 3780 2829
rect 3785 2828 3786 2833
rect 3818 2833 3854 2838
rect 3960 2836 3965 2889
rect 3983 2888 3990 2889
rect 4041 2860 4046 2948
rect 4003 2855 4046 2860
rect 3779 2827 3786 2828
rect 3803 2828 3810 2829
rect 3745 2822 3752 2823
rect 3756 2824 3763 2825
rect 3756 2819 3757 2824
rect 3762 2819 3763 2824
rect 3803 2823 3804 2828
rect 3809 2823 3810 2828
rect 3818 2827 3819 2833
rect 3824 2832 3854 2833
rect 3824 2827 3825 2832
rect 3849 2829 3854 2832
rect 3959 2835 3966 2836
rect 3959 2830 3960 2835
rect 3965 2830 3966 2835
rect 3959 2829 3966 2830
rect 3818 2826 3825 2827
rect 3848 2828 3855 2829
rect 3848 2823 3849 2828
rect 3854 2823 3855 2828
rect 3877 2827 3884 2828
rect 3803 2822 3810 2823
rect 3832 2822 3839 2823
rect 3848 2822 3855 2823
rect 3861 2822 3867 2823
rect 3804 2819 3809 2822
rect 3756 2814 3809 2819
rect 3832 2817 3833 2822
rect 3838 2817 3839 2822
rect 3861 2817 3862 2822
rect 3866 2817 3867 2822
rect 3832 2816 3867 2817
rect 3833 2812 3867 2816
rect 3877 2822 3878 2827
rect 3883 2822 3884 2827
rect 4003 2822 4008 2855
rect 4066 2832 4073 2833
rect 4066 2827 4067 2832
rect 4072 2827 4073 2832
rect 4066 2826 4073 2827
rect 3877 2821 3884 2822
rect 3903 2821 3910 2822
rect 3877 2816 3904 2821
rect 3909 2816 3910 2821
rect 4003 2821 4015 2822
rect 4003 2816 4009 2821
rect 4014 2816 4015 2821
rect 3877 2795 3882 2816
rect 3903 2815 3910 2816
rect 4008 2815 4015 2816
rect 3710 2789 3882 2795
rect 3710 2769 3715 2789
rect 3709 2768 3716 2769
rect 3709 2763 3710 2768
rect 3715 2763 3716 2768
rect 3709 2762 3716 2763
rect 3756 2765 3809 2770
rect 3833 2768 3867 2772
rect 3745 2761 3752 2762
rect 3745 2756 3746 2761
rect 3751 2756 3752 2761
rect 3756 2760 3757 2765
rect 3762 2760 3763 2765
rect 3804 2762 3809 2765
rect 3832 2767 3867 2768
rect 3832 2762 3833 2767
rect 3838 2762 3839 2767
rect 3861 2762 3862 2767
rect 3866 2762 3867 2767
rect 3902 2763 3909 2764
rect 4008 2763 4015 2764
rect 3756 2759 3763 2760
rect 3803 2761 3810 2762
rect 3832 2761 3839 2762
rect 3848 2761 3855 2762
rect 3861 2761 3867 2762
rect 3877 2762 3903 2763
rect 3745 2755 3752 2756
rect 3779 2756 3786 2757
rect 3779 2755 3780 2756
rect 3746 2751 3780 2755
rect 3785 2751 3786 2756
rect 3803 2756 3804 2761
rect 3809 2756 3810 2761
rect 3803 2755 3810 2756
rect 3818 2757 3825 2758
rect 3746 2750 3786 2751
rect 3818 2751 3819 2757
rect 3824 2752 3825 2757
rect 3848 2756 3849 2761
rect 3854 2756 3855 2761
rect 3848 2755 3855 2756
rect 3877 2757 3878 2762
rect 3883 2758 3903 2762
rect 3908 2758 3909 2763
rect 3883 2757 3884 2758
rect 3902 2757 3909 2758
rect 4004 2758 4009 2763
rect 4014 2758 4015 2763
rect 4004 2757 4015 2758
rect 3877 2756 3884 2757
rect 3849 2752 3854 2755
rect 3824 2751 3854 2752
rect 3818 2746 3854 2751
rect 3877 2729 3882 2756
rect 3709 2723 3882 2729
rect 4004 2729 4009 2757
rect 4004 2724 4047 2729
rect 3709 2700 3714 2723
rect 3746 2701 3786 2702
rect 3708 2699 3715 2700
rect 3708 2694 3709 2699
rect 3714 2694 3715 2699
rect 3746 2697 3780 2701
rect 3708 2693 3715 2694
rect 3745 2696 3752 2697
rect 3745 2691 3746 2696
rect 3751 2691 3752 2696
rect 3779 2696 3780 2697
rect 3785 2696 3786 2701
rect 3818 2701 3854 2706
rect 4042 2705 4047 2724
rect 3779 2695 3786 2696
rect 3803 2696 3810 2697
rect 3745 2690 3752 2691
rect 3756 2692 3763 2693
rect 3756 2687 3757 2692
rect 3762 2687 3763 2692
rect 3803 2691 3804 2696
rect 3809 2691 3810 2696
rect 3818 2695 3819 2701
rect 3824 2700 3854 2701
rect 3824 2695 3825 2700
rect 3849 2697 3854 2700
rect 4041 2704 4048 2705
rect 4041 2699 4042 2704
rect 4047 2699 4048 2704
rect 4041 2698 4048 2699
rect 4067 2697 4072 2826
rect 4075 2697 4082 2698
rect 3818 2694 3825 2695
rect 3848 2696 3855 2697
rect 3848 2691 3849 2696
rect 3854 2691 3855 2696
rect 3877 2695 3884 2696
rect 3803 2690 3810 2691
rect 3832 2690 3839 2691
rect 3848 2690 3855 2691
rect 3861 2690 3867 2691
rect 3804 2687 3809 2690
rect 3756 2682 3809 2687
rect 3832 2685 3833 2690
rect 3838 2685 3839 2690
rect 3861 2685 3862 2690
rect 3866 2685 3867 2690
rect 3832 2684 3867 2685
rect 3833 2680 3867 2684
rect 3877 2690 3878 2695
rect 3883 2690 3884 2695
rect 3959 2695 3966 2696
rect 3959 2690 3960 2695
rect 3965 2690 3966 2695
rect 4055 2692 4076 2697
rect 4081 2692 4082 2697
rect 4055 2691 4067 2692
rect 4075 2691 4082 2692
rect 3877 2689 3884 2690
rect 3903 2689 3910 2690
rect 3959 2689 3966 2690
rect 3984 2689 3991 2690
rect 3877 2684 3904 2689
rect 3909 2684 3910 2689
rect 3960 2684 3985 2689
rect 3990 2684 3991 2689
rect 3877 2663 3882 2684
rect 3903 2683 3910 2684
rect 3984 2683 3991 2684
rect 4055 2683 4060 2691
rect 3710 2657 3882 2663
rect 4022 2662 4060 2683
rect 3710 2637 3715 2657
rect 3709 2636 3716 2637
rect 3709 2631 3710 2636
rect 3715 2631 3716 2636
rect 3709 2630 3716 2631
rect 3756 2633 3809 2638
rect 3833 2636 3867 2640
rect 3745 2629 3752 2630
rect 3745 2624 3746 2629
rect 3751 2624 3752 2629
rect 3756 2628 3757 2633
rect 3762 2628 3763 2633
rect 3804 2630 3809 2633
rect 3832 2635 3867 2636
rect 3832 2630 3833 2635
rect 3838 2630 3839 2635
rect 3861 2630 3862 2635
rect 3866 2630 3867 2635
rect 3756 2627 3763 2628
rect 3803 2629 3810 2630
rect 3832 2629 3839 2630
rect 3848 2629 3855 2630
rect 3861 2629 3867 2630
rect 3877 2630 3884 2631
rect 3745 2623 3752 2624
rect 3779 2624 3786 2625
rect 3779 2623 3780 2624
rect 3746 2619 3780 2623
rect 3785 2619 3786 2624
rect 3803 2624 3804 2629
rect 3809 2624 3810 2629
rect 3803 2623 3810 2624
rect 3818 2625 3825 2626
rect 3746 2618 3786 2619
rect 3818 2619 3819 2625
rect 3824 2620 3825 2625
rect 3848 2624 3849 2629
rect 3854 2624 3855 2629
rect 3877 2625 3878 2630
rect 3883 2628 3884 2630
rect 3903 2628 3910 2629
rect 3983 2628 3990 2629
rect 3883 2625 3904 2628
rect 3877 2624 3904 2625
rect 3848 2623 3855 2624
rect 3878 2623 3904 2624
rect 3909 2623 3910 2628
rect 3849 2620 3854 2623
rect 3824 2619 3854 2620
rect 3818 2614 3854 2619
rect 3878 2597 3883 2623
rect 3903 2622 3910 2623
rect 3960 2623 3984 2628
rect 3989 2623 3990 2628
rect 3709 2591 3883 2597
rect 3709 2568 3714 2591
rect 3746 2569 3786 2570
rect 3708 2567 3715 2568
rect 3708 2562 3709 2567
rect 3714 2562 3715 2567
rect 3746 2565 3780 2569
rect 3708 2561 3715 2562
rect 3745 2564 3752 2565
rect 3745 2559 3746 2564
rect 3751 2559 3752 2564
rect 3779 2564 3780 2565
rect 3785 2564 3786 2569
rect 3818 2569 3854 2574
rect 3960 2572 3965 2623
rect 3983 2622 3990 2623
rect 3779 2563 3786 2564
rect 3803 2564 3810 2565
rect 3745 2558 3752 2559
rect 3756 2560 3763 2561
rect 3756 2555 3757 2560
rect 3762 2555 3763 2560
rect 3803 2559 3804 2564
rect 3809 2559 3810 2564
rect 3818 2563 3819 2569
rect 3824 2568 3854 2569
rect 3824 2563 3825 2568
rect 3849 2565 3854 2568
rect 3959 2571 3966 2572
rect 3959 2566 3960 2571
rect 3965 2566 3966 2571
rect 3959 2565 3966 2566
rect 3818 2562 3825 2563
rect 3848 2564 3855 2565
rect 3848 2559 3849 2564
rect 3854 2559 3855 2564
rect 3877 2563 3884 2564
rect 3803 2558 3810 2559
rect 3832 2558 3839 2559
rect 3848 2558 3855 2559
rect 3861 2558 3867 2559
rect 3804 2555 3809 2558
rect 3756 2550 3809 2555
rect 3832 2553 3833 2558
rect 3838 2553 3839 2558
rect 3861 2553 3862 2558
rect 3866 2553 3867 2558
rect 3832 2552 3867 2553
rect 3833 2548 3867 2552
rect 3877 2558 3878 2563
rect 3883 2558 3884 2563
rect 3877 2557 3884 2558
rect 3903 2557 3910 2558
rect 3877 2552 3904 2557
rect 3909 2552 3910 2557
rect 4022 2553 4027 2662
rect 4072 2624 4079 2625
rect 4072 2619 4073 2624
rect 4078 2619 4079 2624
rect 4072 2618 4079 2619
rect 3979 2552 4027 2553
rect 3877 2531 3882 2552
rect 3903 2551 3910 2552
rect 3710 2525 3882 2531
rect 3948 2547 4027 2552
rect 4073 2556 4078 2618
rect 4073 2550 4140 2556
rect 3710 2505 3715 2525
rect 3709 2504 3716 2505
rect 3709 2499 3710 2504
rect 3715 2499 3716 2504
rect 3709 2498 3716 2499
rect 3756 2501 3809 2506
rect 3833 2504 3867 2508
rect 3948 2504 3953 2547
rect 3745 2497 3752 2498
rect 3745 2492 3746 2497
rect 3751 2492 3752 2497
rect 3756 2496 3757 2501
rect 3762 2496 3763 2501
rect 3804 2498 3809 2501
rect 3832 2503 3867 2504
rect 3832 2498 3833 2503
rect 3838 2498 3839 2503
rect 3861 2498 3862 2503
rect 3866 2498 3867 2503
rect 3947 2503 3954 2504
rect 3756 2495 3763 2496
rect 3803 2497 3810 2498
rect 3832 2497 3839 2498
rect 3848 2497 3855 2498
rect 3861 2497 3867 2498
rect 3877 2498 3884 2499
rect 3745 2491 3752 2492
rect 3779 2492 3786 2493
rect 3779 2491 3780 2492
rect 3746 2487 3780 2491
rect 3785 2487 3786 2492
rect 3803 2492 3804 2497
rect 3809 2492 3810 2497
rect 3803 2491 3810 2492
rect 3818 2493 3825 2494
rect 3746 2486 3786 2487
rect 3818 2487 3819 2493
rect 3824 2488 3825 2493
rect 3848 2492 3849 2497
rect 3854 2492 3855 2497
rect 3877 2493 3878 2498
rect 3883 2493 3884 2498
rect 3947 2498 3948 2503
rect 3953 2498 3954 2503
rect 4017 2501 4070 2506
rect 4094 2504 4128 2508
rect 4135 2504 4140 2550
rect 3947 2497 3954 2498
rect 4006 2497 4013 2498
rect 3877 2492 3884 2493
rect 3902 2492 3909 2493
rect 3848 2491 3855 2492
rect 3849 2488 3854 2491
rect 3824 2487 3854 2488
rect 3879 2487 3903 2492
rect 3908 2487 3909 2492
rect 4006 2492 4007 2497
rect 4012 2492 4013 2497
rect 4017 2496 4018 2501
rect 4023 2496 4024 2501
rect 4065 2498 4070 2501
rect 4093 2503 4128 2504
rect 4093 2498 4094 2503
rect 4099 2498 4100 2503
rect 4122 2498 4123 2503
rect 4127 2498 4128 2503
rect 4017 2495 4024 2496
rect 4064 2497 4071 2498
rect 4093 2497 4100 2498
rect 4109 2497 4116 2498
rect 4122 2497 4128 2498
rect 4134 2503 4141 2504
rect 4134 2498 4135 2503
rect 4140 2498 4141 2503
rect 4134 2497 4141 2498
rect 4006 2491 4013 2492
rect 4040 2492 4047 2493
rect 4040 2491 4041 2492
rect 3818 2482 3854 2487
rect 3902 2486 3909 2487
rect 4007 2487 4041 2491
rect 4046 2487 4047 2492
rect 4064 2492 4065 2497
rect 4070 2492 4071 2497
rect 4064 2491 4071 2492
rect 4079 2493 4086 2494
rect 4007 2486 4047 2487
rect 4079 2487 4080 2493
rect 4085 2488 4086 2493
rect 4109 2492 4110 2497
rect 4115 2492 4116 2497
rect 4109 2491 4116 2492
rect 4110 2488 4115 2491
rect 4085 2487 4115 2488
rect 4079 2482 4115 2487
rect 4162 2459 4167 2986
rect 4009 2454 4167 2459
rect 4180 2503 4236 2508
rect 4009 2392 4014 2454
rect 4008 2391 4014 2392
rect 4008 2387 4009 2391
rect 4013 2387 4014 2391
rect 4008 2386 4014 2387
rect 4180 2329 4185 2503
rect 4134 2324 4185 2329
rect 4134 2310 4139 2324
rect 4133 2309 4139 2310
rect 4133 2305 4134 2309
rect 4138 2305 4139 2309
rect 4133 2304 4139 2305
rect 2934 2120 3689 2125
use BlankPad  t0
timestamp 1006127261
transform 1 0 960 0 1 4368
box -11 -51 298 632
use GNDPad  t1
timestamp 1509371954
transform 1 0 1258 0 1 4352
box 0 -35 309 648
use InPad  t2
timestamp 1509371954
transform 1 0 1599 0 1 4683
box -32 -366 277 317
use InPad  t3
timestamp 1509371954
transform 1 0 1908 0 1 4683
box -32 -366 277 317
use InPad  t4
timestamp 1509371954
transform 1 0 2217 0 1 4683
box -32 -366 277 317
use InPad  InPad_0
timestamp 1509371954
transform 1 0 2526 0 1 4683
box -32 -366 277 317
use InPad  InPad_1
timestamp 1509371954
transform 1 0 2835 0 1 4683
box -32 -366 277 317
use GNDPad  GNDPad_0
timestamp 1509371954
transform 1 0 3112 0 1 4352
box 0 -35 309 648
use VddPad  t8
timestamp 1509371954
transform 1 0 3421 0 1 4352
box 0 -35 309 648
use InPad  InPad_2
timestamp 1509371954
transform 1 0 3762 0 1 4683
box -32 -366 277 317
use Corner  crt
timestamp 1012241868
transform 0 1 4369 -1 0 4825
box -143 -333 774 618
use Corner  clt
timestamp 1012241868
transform 1 0 175 0 1 4369
box -143 -333 774 618
use BlankPad  l9
timestamp 1006127261
transform 0 -1 632 1 0 3740
box -11 -51 298 632
use BlankPad  l8
timestamp 1006127261
transform 0 -1 632 1 0 3431
box -11 -51 298 632
use BlankPad  l7
timestamp 1006127261
transform 0 -1 632 1 0 3122
box -11 -51 298 632
use BlankPad  l6
timestamp 1006127261
transform 0 -1 632 1 0 2813
box -11 -51 298 632
use BlankPad  l5
timestamp 1006127261
transform 0 -1 632 1 0 2504
box -11 -51 298 632
use BlankPad  l4
timestamp 1006127261
transform 0 -1 632 1 0 2195
box -11 -51 298 632
use BlankPad  l3
timestamp 1006127261
transform 0 -1 632 1 0 1886
box -11 -51 298 632
use BlankPad  l2
timestamp 1006127261
transform 0 -1 632 1 0 1577
box -11 -51 298 632
use BlankPad  l1
timestamp 1006127261
transform 0 -1 632 1 0 1268
box -11 -51 298 632
use BlankPad  r9
timestamp 1006127261
transform 0 1 4368 -1 0 4040
box -11 -51 298 632
use BlankPad  r8
timestamp 1006127261
transform 0 1 4368 -1 0 3731
box -11 -51 298 632
use BlankPad  r7
timestamp 1006127261
transform 0 1 4368 -1 0 3422
box -11 -51 298 632
use BlankPad  r6
timestamp 1006127261
transform 0 1 4368 -1 0 3113
box -11 -51 298 632
use OutPad  OutPad_0
timestamp 1012172318
transform 0 1 4343 1 0 2489
box 17 -26 326 657
use BlankPad  r5
timestamp 1006127261
transform 0 1 4368 1 0 2208
box -11 -51 298 632
use BlankPad  r3
timestamp 1006127261
transform 0 1 4368 -1 0 2186
box -11 -51 298 632
use BlankPad  r2
timestamp 1006127261
transform 0 1 4368 -1 0 1877
box -11 -51 298 632
use BlankPad  r1
timestamp 1006127261
transform 0 1 4368 -1 0 1568
box -11 -51 298 632
use BlankPad  r0
timestamp 1006127261
transform 0 1 4368 -1 0 1259
box -11 -51 298 632
use BlankPad  l0
timestamp 1006127261
transform 0 -1 632 1 0 959
box -11 -51 298 632
use Corner  clb
timestamp 1012241868
transform 0 -1 631 1 0 175
box -143 -333 774 618
use BlankPad  b0
timestamp 1006127261
transform -1 0 1260 0 -1 632
box -11 -51 298 632
use BlankPad  b1
timestamp 1006127261
transform -1 0 1569 0 -1 632
box -11 -51 298 632
use BlankPad  b2
timestamp 1006127261
transform -1 0 1878 0 -1 632
box -11 -51 298 632
use BlankPad  b3
timestamp 1006127261
transform -1 0 2187 0 -1 632
box -11 -51 298 632
use BlankPad  b4
timestamp 1006127261
transform -1 0 2496 0 -1 632
box -11 -51 298 632
use BlankPad  b5
timestamp 1006127261
transform -1 0 2805 0 -1 632
box -11 -51 298 632
use BlankPad  b6
timestamp 1006127261
transform -1 0 3114 0 -1 632
box -11 -51 298 632
use BlankPad  b7
timestamp 1006127261
transform -1 0 3423 0 -1 632
box -11 -51 298 632
use BlankPad  b8
timestamp 1006127261
transform -1 0 3732 0 -1 632
box -11 -51 298 632
use Corner  crb
timestamp 1012241868
transform -1 0 4825 0 -1 631
box -143 -333 774 618
use BlankPad  b9
timestamp 1006127261
transform -1 0 4041 0 -1 632
box -11 -51 298 632
<< labels >>
rlabel metal1 1716 4857 1720 4857 1 p0
rlabel metal1 2031 4873 2031 4873 1 p1
rlabel metal1 2340 4865 2340 4865 1 p2
rlabel metal1 3267 4862 3267 4862 1 p5
rlabel metal1 1417 4883 1419 4884 1 p6
rlabel metal1 3571 4861 3572 4861 1 p7
rlabel metal1 2637 4868 2637 4868 1 p3
rlabel metal1 2951 4862 2951 4862 1 p4
rlabel metal2 2954 4304 2967 4317 1 mode
rlabel metal2 3229 3828 3242 3841 1 clk
rlabel metal2 3574 3708 3578 3725 1 GND!
rlabel metal2 3582 3718 3586 3735 1 Vdd!
rlabel metal2 3590 3718 3594 3735 1 reset_b
rlabel metal1 3302 3599 3305 3603 1 GND!
rlabel metal1 3301 3549 3305 3553 1 Vdd!
rlabel metal1 3300 3577 3304 3580 1 clk
rlabel metal1 3302 3729 3305 3733 1 GND!
rlabel metal1 3300 3707 3304 3710 1 clk
rlabel metal1 3301 3679 3305 3683 1 Vdd!
rlabel metal1 3251 3658 3252 3661 3 enable
rlabel metal1 3301 3809 3305 3813 1 Vdd!
rlabel metal2 2692 4063 2692 4063 1 GND!
rlabel metal2 2680 4063 2680 4063 1 Vdd!
rlabel metal1 2529 3919 2532 3923 6 clk
rlabel metal1 2527 3848 2530 3852 8 ~clk
rlabel metal1 2528 3855 2531 3859 1 GND!
rlabel metal1 2529 3912 2532 3916 1 Vdd!
rlabel metal1 2413 4021 2416 4025 4 clk
rlabel metal1 2415 3950 2418 3954 2 ~clk
rlabel metal1 2414 3957 2417 3961 1 GND!
rlabel metal1 2413 4014 2416 4018 1 Vdd!
rlabel metal2 2705 4062 2705 4062 4 f_clk_b
rlabel metal2 2717 4061 2717 4061 5 f_clk
rlabel metal2 2741 4062 2741 4062 5 p_clk
rlabel metal2 2729 4062 2729 4062 5 p_clk_b
rlabel metal1 2545 3519 2548 3523 4 clk
rlabel metal1 2547 3448 2550 3452 2 ~clk
rlabel metal1 2546 3455 2549 3459 1 GND!
rlabel metal1 2545 3512 2548 3516 1 Vdd!
rlabel metal1 2413 3519 2416 3523 4 clk
rlabel metal1 2415 3448 2418 3452 2 ~clk
rlabel metal1 2414 3455 2417 3459 1 GND!
rlabel metal1 2413 3512 2416 3516 1 Vdd!
rlabel metal1 2281 3519 2284 3523 4 clk
rlabel metal1 2283 3448 2286 3452 2 ~clk
rlabel metal1 2282 3455 2285 3459 1 GND!
rlabel metal1 2281 3512 2284 3516 1 Vdd!
rlabel metal2 3637 4063 3637 4063 1 GND!
rlabel metal2 3625 4063 3625 4063 1 Vdd!
rlabel polysilicon 3371 3933 3371 3933 1 CB1
rlabel metal1 3479 3887 3479 3887 1 D
rlabel metal1 3474 3919 3477 3923 6 clk
rlabel metal1 3472 3848 3475 3852 8 ~clk
rlabel metal1 3473 3855 3476 3859 1 GND!
rlabel metal1 3474 3912 3477 3916 1 Vdd!
rlabel polysilicon 3488 3941 3488 3941 1 CB2
rlabel metal1 3358 4021 3361 4025 4 clk
rlabel metal1 3360 3950 3363 3954 2 ~clk
rlabel metal1 3359 3957 3362 3961 1 GND!
rlabel metal1 3358 4014 3361 4018 1 Vdd!
rlabel metal2 3650 4062 3650 4062 4 f_clk_b
rlabel metal2 3662 4061 3662 4061 5 f_clk
rlabel metal2 3674 4062 3674 4062 5 p_clk_b
rlabel metal1 3490 3519 3493 3523 4 clk
rlabel metal1 3492 3448 3495 3452 2 ~clk
rlabel metal1 3491 3455 3494 3459 1 GND!
rlabel metal1 3490 3512 3493 3516 1 Vdd!
rlabel metal1 3358 3519 3361 3523 4 clk
rlabel metal1 3360 3448 3363 3452 2 ~clk
rlabel metal1 3359 3455 3362 3459 1 GND!
rlabel metal1 3358 3512 3361 3516 1 Vdd!
rlabel metal1 3226 3519 3229 3523 4 clk
rlabel metal1 3228 3448 3231 3452 2 ~clk
rlabel metal1 3227 3455 3230 3459 1 GND!
rlabel metal1 3226 3512 3229 3516 1 Vdd!
rlabel polysilicon 3204 3430 3204 3430 1 CB3
rlabel metal1 2897 4047 2900 4051 1 Vdd!
rlabel metal1 3019 3449 3022 3453 1 clk
rlabel metal1 3016 3501 3020 3505 1 ~clk
rlabel metal1 3015 3508 3019 3512 1 GND!
rlabel metal1 3026 3442 3030 3446 1 Vdd!
rlabel metal2 3082 3974 3085 3980 1 select2
rlabel metal2 3022 3974 3025 3981 1 select1
rlabel metal2 2939 3975 2942 3980 1 select0
rlabel m3contact 2762 4020 2765 4023 3 ctrl_reg
rlabel metal1 3161 4047 3164 4051 1 Vdd!
rlabel metal1 3162 3990 3165 3994 1 GND!
rlabel metal1 3163 3983 3166 3987 2 ~clk
rlabel metal1 3161 4054 3164 4058 4 clk
rlabel metal1 3029 4054 3032 4058 4 clk
rlabel metal1 3031 3983 3034 3987 2 ~clk
rlabel metal1 3030 3990 3033 3994 1 GND!
rlabel metal1 3029 4047 3032 4051 1 Vdd!
rlabel metal1 2897 4054 2900 4058 4 clk
rlabel metal1 2899 3983 2902 3987 2 ~clk
rlabel metal1 2898 3990 2901 3994 1 GND!
rlabel metal1 2765 4054 2768 4058 4 clk
rlabel metal1 2767 3983 2770 3987 2 ~clk
rlabel metal1 2766 3990 2769 3994 1 GND!
rlabel metal1 2765 4047 2768 4051 1 Vdd!
rlabel metal2 3110 3965 3113 3970 1 select_out
rlabel metal1 3047 3904 3050 3908 1 GND!
rlabel metal1 2966 3904 2969 3908 1 GND!
rlabel metal1 3046 3970 3050 3974 1 Vdd!
rlabel metal1 2965 3970 2969 3974 1 Vdd!
rlabel metal1 3115 3809 3118 3812 7 Y
rlabel metal1 3046 3838 3050 3842 1 Vdd!
rlabel metal1 2965 3838 2969 3842 1 Vdd!
rlabel metal1 3071 3772 3074 3776 1 GND!
rlabel metal1 2966 3772 2969 3776 1 GND!
rlabel metal1 3046 3706 3050 3710 1 Vdd!
rlabel metal1 2965 3706 2969 3710 1 Vdd!
rlabel metal1 3136 3706 3140 3710 1 Vdd!
rlabel metal1 2966 3640 2969 3644 1 GND!
rlabel metal1 3047 3640 3050 3644 1 GND!
rlabel metal1 3137 3640 3140 3644 1 GND!
rlabel metal1 2965 3574 2969 3578 1 Vdd!
rlabel metal1 3046 3574 3050 3578 1 Vdd!
rlabel metal1 3136 3574 3140 3578 1 Vdd!
rlabel metal1 2966 3508 2969 3512 1 GND!
rlabel metal1 2965 3442 2969 3446 1 Vdd!
rlabel polysilicon 3009 3472 3011 3475 5 D
rlabel polysilicon 3027 3481 3029 3484 5 reset
rlabel metal1 2763 3699 2767 3703 3 clk
rlabel metal1 2763 3706 2767 3710 3 Vdd!
rlabel metal1 2763 3647 2767 3651 3 ~clk
rlabel metal1 2763 3581 2767 3585 3 clk
rlabel metal1 2763 3633 2767 3637 3 ~clk
rlabel metal1 2763 3640 2767 3644 3 GND!
rlabel metal1 2763 3567 2767 3571 3 clk
rlabel metal1 2763 3574 2767 3578 3 Vdd!
rlabel metal1 2763 3515 2767 3519 3 ~clk
rlabel metal1 2763 3442 2767 3446 3 Vdd!
rlabel metal1 2763 3501 2767 3505 3 ~clk
rlabel metal1 2763 3508 2767 3512 3 GND!
rlabel metal1 2763 3772 2767 3776 3 GND!
rlabel metal1 2763 3765 2767 3769 3 ~clk
rlabel metal1 2763 3713 2767 3717 3 clk
rlabel metal1 2763 3779 2767 3783 3 ~clk
rlabel metal1 2763 3838 2767 3842 3 Vdd!
rlabel metal1 2763 3831 2767 3835 3 clk
rlabel metal1 2763 3904 2767 3908 3 GND!
rlabel metal1 2763 3897 2767 3901 3 ~clk
rlabel metal1 2763 3911 2767 3915 3 ~clk
rlabel metal1 2763 3970 2767 3974 3 Vdd!
rlabel metal1 2763 3963 2767 3967 3 clk
rlabel metal1 2282 2473 2285 2477 1 GND!
rlabel metal1 2283 2466 2286 2470 2 ~clk
rlabel metal1 2413 2530 2416 2534 1 Vdd!
rlabel metal1 2414 2473 2417 2477 1 GND!
rlabel metal1 2415 2466 2418 2470 2 ~clk
rlabel metal1 2413 2537 2416 2541 4 clk
rlabel metal1 2545 2530 2548 2534 1 Vdd!
rlabel metal1 2546 2473 2549 2477 1 GND!
rlabel metal1 2547 2466 2550 2470 2 ~clk
rlabel metal1 2545 2537 2548 2541 4 clk
rlabel metal2 2729 3080 2729 3080 5 p_clk_b
rlabel metal2 2741 3080 2741 3080 5 p_clk
rlabel metal2 2717 3079 2717 3079 5 f_clk
rlabel metal2 2705 3080 2705 3080 4 f_clk_b
rlabel metal1 2413 3032 2416 3036 1 Vdd!
rlabel metal1 2414 2975 2417 2979 1 GND!
rlabel metal1 2415 2968 2418 2972 2 ~clk
rlabel metal1 2413 3039 2416 3043 4 clk
rlabel polysilicon 2543 2959 2543 2959 1 CB2
rlabel metal1 2529 2930 2532 2934 1 Vdd!
rlabel metal1 2528 2873 2531 2877 1 GND!
rlabel metal1 2527 2866 2530 2870 8 ~clk
rlabel metal1 2529 2937 2532 2941 6 clk
rlabel metal2 2680 3081 2680 3081 1 Vdd!
rlabel metal2 2692 3081 2692 3081 1 GND!
rlabel metal1 2281 3144 2284 3148 1 Vdd!
rlabel metal1 2282 3087 2285 3091 1 GND!
rlabel metal1 2283 3080 2286 3084 2 ~clk
rlabel metal1 2281 3151 2284 3155 4 clk
rlabel metal1 2413 3144 2416 3148 1 Vdd!
rlabel metal1 2414 3087 2417 3091 1 GND!
rlabel metal1 2415 3080 2418 3084 2 ~clk
rlabel metal1 2413 3151 2416 3155 4 clk
rlabel metal1 2545 3144 2548 3148 1 Vdd!
rlabel metal1 2546 3087 2549 3091 1 GND!
rlabel metal1 2547 3080 2550 3084 2 ~clk
rlabel metal1 2545 3151 2548 3155 4 clk
rlabel metal1 2281 3284 2284 3288 1 Vdd!
rlabel metal1 2282 3227 2285 3231 1 GND!
rlabel metal1 2283 3220 2286 3224 2 ~clk
rlabel metal1 2281 3291 2284 3295 4 clk
rlabel metal1 2413 3284 2416 3288 1 Vdd!
rlabel metal1 2414 3227 2417 3231 1 GND!
rlabel metal1 2415 3220 2418 3224 2 ~clk
rlabel metal1 2413 3291 2416 3295 4 clk
rlabel metal1 2545 3284 2548 3288 1 Vdd!
rlabel metal1 2546 3227 2549 3231 1 GND!
rlabel metal1 2547 3220 2550 3224 2 ~clk
rlabel metal1 2545 3291 2548 3295 4 clk
rlabel metal1 2545 3377 2548 3381 4 clk
rlabel metal1 2547 3306 2550 3310 2 ~clk
rlabel metal1 2546 3313 2549 3317 1 GND!
rlabel metal1 2545 3370 2548 3374 1 Vdd!
rlabel metal1 2413 3377 2416 3381 4 clk
rlabel metal1 2415 3306 2418 3310 2 ~clk
rlabel metal1 2414 3313 2417 3317 1 GND!
rlabel metal1 2413 3370 2416 3374 1 Vdd!
rlabel metal1 2281 3377 2284 3381 4 clk
rlabel metal1 2283 3306 2286 3310 2 ~clk
rlabel metal1 2282 3313 2285 3317 1 GND!
rlabel metal1 2281 3370 2284 3374 1 Vdd!
rlabel metal2 3098 2819 3098 2819 2 Core
rlabel metal1 2763 2981 2767 2985 3 clk
rlabel metal1 2763 2988 2767 2992 3 Vdd!
rlabel metal1 2763 2929 2767 2933 3 ~clk
rlabel metal1 2763 2915 2767 2919 3 ~clk
rlabel metal1 2763 2922 2767 2926 3 GND!
rlabel metal1 2763 2849 2767 2853 3 clk
rlabel metal1 2763 2856 2767 2860 3 Vdd!
rlabel metal1 2763 2797 2767 2801 3 ~clk
rlabel metal1 2763 2731 2767 2735 3 clk
rlabel metal1 2763 2783 2767 2787 3 ~clk
rlabel metal1 2763 2790 2767 2794 3 GND!
rlabel metal1 2763 2526 2767 2530 3 GND!
rlabel metal1 2763 2519 2767 2523 3 ~clk
rlabel metal1 2763 2460 2767 2464 3 Vdd!
rlabel metal1 2763 2533 2767 2537 3 ~clk
rlabel metal1 2763 2592 2767 2596 3 Vdd!
rlabel metal1 2763 2585 2767 2589 3 clk
rlabel metal1 2763 2658 2767 2662 3 GND!
rlabel metal1 2763 2651 2767 2655 3 ~clk
rlabel metal1 2763 2599 2767 2603 3 clk
rlabel metal1 2763 2665 2767 2669 3 ~clk
rlabel metal1 2763 2724 2767 2728 3 Vdd!
rlabel metal1 2763 2717 2767 2721 3 clk
rlabel polysilicon 3027 2499 3029 2502 5 reset
rlabel polysilicon 3009 2490 3011 2493 5 D
rlabel metal1 2965 2460 2969 2464 1 Vdd!
rlabel metal1 2966 2526 2969 2530 1 GND!
rlabel metal1 3136 2592 3140 2596 1 Vdd!
rlabel metal1 3046 2592 3050 2596 1 Vdd!
rlabel metal1 2965 2592 2969 2596 1 Vdd!
rlabel metal1 3137 2658 3140 2662 1 GND!
rlabel metal1 3047 2658 3050 2662 1 GND!
rlabel metal1 2966 2658 2969 2662 1 GND!
rlabel metal1 3136 2724 3140 2728 1 Vdd!
rlabel metal1 2965 2724 2969 2728 1 Vdd!
rlabel metal1 3046 2724 3050 2728 1 Vdd!
rlabel metal1 2966 2790 2969 2794 1 GND!
rlabel metal1 3071 2790 3074 2794 1 GND!
rlabel metal1 2965 2856 2969 2860 1 Vdd!
rlabel metal1 3046 2856 3050 2860 1 Vdd!
rlabel metal1 3115 2827 3118 2830 7 Y
rlabel metal1 2965 2988 2969 2992 1 Vdd!
rlabel metal1 3046 2988 3050 2992 1 Vdd!
rlabel metal1 2966 2922 2969 2926 1 GND!
rlabel metal1 3047 2922 3050 2926 1 GND!
rlabel metal2 3110 2983 3113 2988 1 select_out
rlabel metal1 2765 3065 2768 3069 1 Vdd!
rlabel metal1 2766 3008 2769 3012 1 GND!
rlabel metal1 2767 3001 2770 3005 2 ~clk
rlabel metal1 2765 3072 2768 3076 4 clk
rlabel metal1 2898 3008 2901 3012 1 GND!
rlabel metal1 2899 3001 2902 3005 2 ~clk
rlabel metal1 2897 3072 2900 3076 4 clk
rlabel metal1 3029 3065 3032 3069 1 Vdd!
rlabel metal1 3030 3008 3033 3012 1 GND!
rlabel metal1 3031 3001 3034 3005 2 ~clk
rlabel metal1 3029 3072 3032 3076 4 clk
rlabel metal1 3161 3072 3164 3076 4 clk
rlabel metal1 3163 3001 3166 3005 2 ~clk
rlabel metal1 3162 3008 3165 3012 1 GND!
rlabel metal1 3161 3065 3164 3069 1 Vdd!
rlabel metal2 2939 2993 2942 2998 1 select0
rlabel metal2 3022 2992 3025 2999 1 select1
rlabel metal2 3082 2992 3085 2998 1 select2
rlabel metal1 3026 2460 3030 2464 1 Vdd!
rlabel metal1 3015 2526 3019 2530 1 GND!
rlabel metal1 3016 2519 3020 2523 1 ~clk
rlabel metal1 3019 2467 3022 2471 1 clk
rlabel metal1 2897 3065 2900 3069 1 Vdd!
rlabel metal1 3226 2530 3229 2534 1 Vdd!
rlabel metal1 3227 2473 3230 2477 1 GND!
rlabel metal1 3228 2466 3231 2470 2 ~clk
rlabel metal1 3226 2537 3229 2541 4 clk
rlabel metal1 3358 2530 3361 2534 1 Vdd!
rlabel metal1 3359 2473 3362 2477 1 GND!
rlabel metal1 3360 2466 3363 2470 2 ~clk
rlabel metal1 3358 2537 3361 2541 4 clk
rlabel metal1 3490 2530 3493 2534 1 Vdd!
rlabel metal1 3491 2473 3494 2477 1 GND!
rlabel metal1 3492 2466 3495 2470 2 ~clk
rlabel metal1 3490 2537 3493 2541 4 clk
rlabel metal2 3674 3080 3674 3080 5 p_clk_b
rlabel metal2 3662 3079 3662 3079 5 f_clk
rlabel metal2 3650 3080 3650 3080 4 f_clk_b
rlabel metal1 3358 3032 3361 3036 1 Vdd!
rlabel metal1 3359 2975 3362 2979 1 GND!
rlabel metal1 3360 2968 3363 2972 2 ~clk
rlabel metal1 3358 3039 3361 3043 4 clk
rlabel polysilicon 3488 2959 3488 2959 1 CB2
rlabel metal1 3474 2930 3477 2934 1 Vdd!
rlabel metal1 3473 2873 3476 2877 1 GND!
rlabel metal1 3472 2866 3475 2870 8 ~clk
rlabel metal1 3474 2937 3477 2941 6 clk
rlabel polysilicon 3371 2951 3371 2951 1 CB1
rlabel metal2 3625 3081 3625 3081 1 Vdd!
rlabel metal2 3637 3081 3637 3081 1 GND!
rlabel metal1 3226 3144 3229 3148 1 Vdd!
rlabel metal1 3227 3087 3230 3091 1 GND!
rlabel metal1 3228 3080 3231 3084 2 ~clk
rlabel metal1 3226 3151 3229 3155 4 clk
rlabel metal1 3358 3144 3361 3148 1 Vdd!
rlabel metal1 3359 3087 3362 3091 1 GND!
rlabel metal1 3360 3080 3363 3084 2 ~clk
rlabel metal1 3358 3151 3361 3155 4 clk
rlabel metal1 3490 3144 3493 3148 1 Vdd!
rlabel metal1 3491 3087 3494 3091 1 GND!
rlabel metal1 3492 3080 3495 3084 2 ~clk
rlabel metal1 3490 3151 3493 3155 4 clk
rlabel metal1 3226 3284 3229 3288 1 Vdd!
rlabel metal1 3227 3227 3230 3231 1 GND!
rlabel metal1 3228 3220 3231 3224 2 ~clk
rlabel metal1 3226 3291 3229 3295 4 clk
rlabel metal1 3358 3284 3361 3288 1 Vdd!
rlabel metal1 3359 3227 3362 3231 1 GND!
rlabel metal1 3360 3220 3363 3224 2 ~clk
rlabel metal1 3358 3291 3361 3295 4 clk
rlabel metal1 3490 3284 3493 3288 1 Vdd!
rlabel metal1 3491 3227 3494 3231 1 GND!
rlabel metal1 3492 3220 3495 3224 2 ~clk
rlabel metal1 3490 3291 3493 3295 4 clk
rlabel metal1 3490 3377 3493 3381 4 clk
rlabel metal1 3492 3306 3495 3310 2 ~clk
rlabel metal1 3491 3313 3494 3317 1 GND!
rlabel metal1 3490 3370 3493 3374 1 Vdd!
rlabel metal1 3358 3377 3361 3381 4 clk
rlabel metal1 3360 3306 3363 3310 2 ~clk
rlabel metal1 3359 3313 3362 3317 1 GND!
rlabel metal1 3358 3370 3361 3374 1 Vdd!
rlabel metal1 3226 3377 3229 3381 4 clk
rlabel metal1 3228 3306 3231 3310 2 ~clk
rlabel metal1 3227 3313 3230 3317 1 GND!
rlabel metal1 3226 3370 3229 3374 1 Vdd!
rlabel polysilicon 3216 3284 3216 3284 1 CB4
rlabel metal1 3064 3321 3067 3325 4 clk
rlabel metal1 3066 3250 3069 3254 2 ~clk
rlabel metal1 3065 3257 3068 3261 1 GND!
rlabel metal1 3064 3314 3067 3318 1 Vdd!
rlabel metal1 3064 3400 3067 3404 1 Vdd!
rlabel metal1 3065 3343 3068 3347 1 GND!
rlabel metal1 3066 3336 3069 3340 2 ~clk
rlabel metal1 3064 3407 3067 3411 4 clk
rlabel metal1 2281 2388 2284 2392 1 Vdd!
rlabel metal1 2282 2331 2285 2335 1 GND!
rlabel metal1 2283 2324 2286 2328 2 ~clk
rlabel metal1 2281 2395 2284 2399 4 clk
rlabel metal1 2413 2388 2416 2392 1 Vdd!
rlabel metal1 2414 2331 2417 2335 1 GND!
rlabel metal1 2415 2324 2418 2328 2 ~clk
rlabel metal1 2413 2395 2416 2399 4 clk
rlabel metal1 2545 2388 2548 2392 1 Vdd!
rlabel metal1 2546 2331 2549 2335 1 GND!
rlabel metal1 2547 2324 2550 2328 2 ~clk
rlabel metal1 2545 2395 2548 2399 4 clk
rlabel metal1 2545 2309 2548 2313 4 clk
rlabel metal1 2547 2238 2550 2242 2 ~clk
rlabel metal1 2546 2245 2549 2249 1 GND!
rlabel metal1 2545 2302 2548 2306 1 Vdd!
rlabel metal1 2413 2309 2416 2313 4 clk
rlabel metal1 2415 2238 2418 2242 2 ~clk
rlabel metal1 2414 2245 2417 2249 1 GND!
rlabel metal1 2413 2302 2416 2306 1 Vdd!
rlabel metal1 2281 2309 2284 2313 4 clk
rlabel metal1 2283 2238 2286 2242 2 ~clk
rlabel metal1 2282 2245 2285 2249 1 GND!
rlabel metal1 2281 2302 2284 2306 1 Vdd!
rlabel metal1 2545 2169 2548 2173 4 clk
rlabel metal1 2547 2098 2550 2102 2 ~clk
rlabel metal1 2546 2105 2549 2109 1 GND!
rlabel metal1 2545 2162 2548 2166 1 Vdd!
rlabel metal1 2413 2169 2416 2173 4 clk
rlabel metal1 2415 2098 2418 2102 2 ~clk
rlabel metal1 2414 2105 2417 2109 1 GND!
rlabel metal1 2413 2162 2416 2166 1 Vdd!
rlabel metal1 2281 2169 2284 2173 4 clk
rlabel metal1 2283 2098 2286 2102 2 ~clk
rlabel metal1 2282 2105 2285 2109 1 GND!
rlabel metal1 2281 2162 2284 2166 1 Vdd!
rlabel metal1 3064 2425 3067 2429 4 clk
rlabel metal1 3066 2354 3069 2358 2 ~clk
rlabel metal1 3065 2361 3068 2365 1 GND!
rlabel metal1 3064 2332 3067 2336 1 Vdd!
rlabel metal1 3065 2275 3068 2279 1 GND!
rlabel metal1 3066 2268 3069 2272 2 ~clk
rlabel metal1 3064 2339 3067 2343 4 clk
rlabel metal1 3226 2388 3229 2392 1 Vdd!
rlabel metal1 3227 2331 3230 2335 1 GND!
rlabel metal1 3228 2324 3231 2328 2 ~clk
rlabel metal1 3226 2395 3229 2399 4 clk
rlabel metal1 3358 2388 3361 2392 1 Vdd!
rlabel metal1 3359 2331 3362 2335 1 GND!
rlabel metal1 3360 2324 3363 2328 2 ~clk
rlabel metal1 3358 2395 3361 2399 4 clk
rlabel metal1 3490 2388 3493 2392 1 Vdd!
rlabel metal1 3491 2331 3494 2335 1 GND!
rlabel metal1 3492 2324 3495 2328 2 ~clk
rlabel metal1 3490 2395 3493 2399 4 clk
rlabel metal1 3490 2309 3493 2313 4 clk
rlabel metal1 3492 2238 3495 2242 2 ~clk
rlabel metal1 3491 2245 3494 2249 1 GND!
rlabel metal1 3490 2302 3493 2306 1 Vdd!
rlabel metal1 3358 2309 3361 2313 4 clk
rlabel metal1 3360 2238 3363 2242 2 ~clk
rlabel metal1 3359 2245 3362 2249 1 GND!
rlabel metal1 3358 2302 3361 2306 1 Vdd!
rlabel metal1 3226 2309 3229 2313 4 clk
rlabel metal1 3228 2238 3231 2242 2 ~clk
rlabel metal1 3227 2245 3230 2249 1 GND!
rlabel metal1 3226 2302 3229 2306 1 Vdd!
rlabel metal1 3490 2169 3493 2173 4 clk
rlabel metal1 3492 2098 3495 2102 2 ~clk
rlabel metal1 3491 2105 3494 2109 1 GND!
rlabel metal1 3490 2162 3493 2166 1 Vdd!
rlabel metal1 3358 2169 3361 2173 4 clk
rlabel metal1 3360 2098 3363 2102 2 ~clk
rlabel metal1 3359 2105 3362 2109 1 GND!
rlabel metal1 3358 2162 3361 2166 1 Vdd!
rlabel metal1 3226 2169 3229 2173 4 clk
rlabel metal1 3228 2098 3231 2102 2 ~clk
rlabel metal1 3227 2105 3230 2109 1 GND!
rlabel metal1 3226 2162 3229 2166 1 Vdd!
rlabel metal1 3077 2418 3080 2422 1 Vdd!
rlabel metal2 3686 4062 3686 4062 5 p_clk
rlabel metal2 3686 3080 3686 3080 5 p_clk
rlabel metal1 4140 3679 4140 3679 1 out
rlabel metal1 3842 4047 3845 4051 1 Vdd!
rlabel metal1 3964 3449 3967 3453 1 clk
rlabel metal1 3961 3501 3965 3505 1 ~clk
rlabel metal1 3960 3508 3964 3512 1 GND!
rlabel metal1 3971 3442 3975 3446 1 Vdd!
rlabel metal2 4027 3974 4030 3980 1 select2
rlabel metal2 3967 3974 3970 3981 1 select1
rlabel metal2 3884 3975 3887 3980 1 select0
rlabel m3contact 3707 4020 3710 4023 3 ctrl_reg
rlabel metal1 4106 4047 4109 4051 1 Vdd!
rlabel metal1 4107 3990 4110 3994 1 GND!
rlabel metal1 4108 3983 4111 3987 2 ~clk
rlabel metal1 4106 4054 4109 4058 4 clk
rlabel metal1 3974 4054 3977 4058 4 clk
rlabel metal1 3976 3983 3979 3987 2 ~clk
rlabel metal1 3975 3990 3978 3994 1 GND!
rlabel metal1 3974 4047 3977 4051 1 Vdd!
rlabel metal1 3842 4054 3845 4058 4 clk
rlabel metal1 3844 3983 3847 3987 2 ~clk
rlabel metal1 3843 3990 3846 3994 1 GND!
rlabel metal1 3710 4054 3713 4058 4 clk
rlabel metal1 3712 3983 3715 3987 2 ~clk
rlabel metal1 3711 3990 3714 3994 1 GND!
rlabel metal1 3710 4047 3713 4051 1 Vdd!
rlabel metal2 4055 3965 4058 3970 1 select_out
rlabel metal1 3992 3904 3995 3908 1 GND!
rlabel metal1 3911 3904 3914 3908 1 GND!
rlabel metal1 3991 3970 3995 3974 1 Vdd!
rlabel metal1 3910 3970 3914 3974 1 Vdd!
rlabel metal1 4060 3809 4063 3812 7 Y
rlabel metal1 3991 3838 3995 3842 1 Vdd!
rlabel metal1 3910 3838 3914 3842 1 Vdd!
rlabel metal1 4016 3772 4019 3776 1 GND!
rlabel metal1 3911 3772 3914 3776 1 GND!
rlabel metal1 3991 3706 3995 3710 1 Vdd!
rlabel metal1 3910 3706 3914 3710 1 Vdd!
rlabel metal1 4081 3706 4085 3710 1 Vdd!
rlabel metal1 3911 3640 3914 3644 1 GND!
rlabel metal1 3992 3640 3995 3644 1 GND!
rlabel metal1 4082 3640 4085 3644 1 GND!
rlabel metal1 3910 3574 3914 3578 1 Vdd!
rlabel metal1 3991 3574 3995 3578 1 Vdd!
rlabel metal1 4081 3574 4085 3578 1 Vdd!
rlabel metal1 3911 3508 3914 3512 1 GND!
rlabel metal1 3910 3442 3914 3446 1 Vdd!
rlabel polysilicon 3972 3481 3974 3484 5 reset
rlabel metal1 3708 3699 3712 3703 3 clk
rlabel metal1 3708 3706 3712 3710 3 Vdd!
rlabel metal1 3708 3647 3712 3651 3 ~clk
rlabel metal1 3708 3581 3712 3585 3 clk
rlabel metal1 3708 3633 3712 3637 3 ~clk
rlabel metal1 3708 3640 3712 3644 3 GND!
rlabel metal1 3708 3567 3712 3571 3 clk
rlabel metal1 3708 3574 3712 3578 3 Vdd!
rlabel metal1 3708 3515 3712 3519 3 ~clk
rlabel metal1 3708 3442 3712 3446 3 Vdd!
rlabel metal1 3708 3501 3712 3505 3 ~clk
rlabel metal1 3708 3508 3712 3512 3 GND!
rlabel metal1 3708 3772 3712 3776 3 GND!
rlabel metal1 3708 3765 3712 3769 3 ~clk
rlabel metal1 3708 3713 3712 3717 3 clk
rlabel metal1 3708 3779 3712 3783 3 ~clk
rlabel metal1 3708 3838 3712 3842 3 Vdd!
rlabel metal1 3708 3831 3712 3835 3 clk
rlabel metal1 3708 3904 3712 3908 3 GND!
rlabel metal1 3708 3897 3712 3901 3 ~clk
rlabel metal1 3708 3911 3712 3915 3 ~clk
rlabel metal1 3708 3970 3712 3974 3 Vdd!
rlabel metal1 3708 3963 3712 3967 3 clk
rlabel metal1 3708 2981 3712 2985 3 clk
rlabel metal1 3708 2988 3712 2992 3 Vdd!
rlabel metal1 3708 2929 3712 2933 3 ~clk
rlabel metal1 3708 2915 3712 2919 3 ~clk
rlabel metal1 3708 2922 3712 2926 3 GND!
rlabel metal1 3708 2849 3712 2853 3 clk
rlabel metal1 3708 2856 3712 2860 3 Vdd!
rlabel metal1 3708 2797 3712 2801 3 ~clk
rlabel metal1 3708 2731 3712 2735 3 clk
rlabel metal1 3708 2783 3712 2787 3 ~clk
rlabel metal1 3708 2790 3712 2794 3 GND!
rlabel metal1 3708 2526 3712 2530 3 GND!
rlabel metal1 3708 2519 3712 2523 3 ~clk
rlabel metal1 3708 2460 3712 2464 3 Vdd!
rlabel metal1 3708 2533 3712 2537 3 ~clk
rlabel metal1 3708 2592 3712 2596 3 Vdd!
rlabel metal1 3708 2585 3712 2589 3 clk
rlabel metal1 3708 2658 3712 2662 3 GND!
rlabel metal1 3708 2651 3712 2655 3 ~clk
rlabel metal1 3708 2599 3712 2603 3 clk
rlabel metal1 3708 2665 3712 2669 3 ~clk
rlabel metal1 3708 2724 3712 2728 3 Vdd!
rlabel metal1 3708 2717 3712 2721 3 clk
rlabel polysilicon 3972 2499 3974 2502 5 reset
rlabel polysilicon 3954 2490 3956 2493 5 D
rlabel metal1 3910 2460 3914 2464 1 Vdd!
rlabel metal1 3911 2526 3914 2530 1 GND!
rlabel metal1 4081 2592 4085 2596 1 Vdd!
rlabel metal1 3991 2592 3995 2596 1 Vdd!
rlabel metal1 3910 2592 3914 2596 1 Vdd!
rlabel metal1 4082 2658 4085 2662 1 GND!
rlabel metal1 3992 2658 3995 2662 1 GND!
rlabel metal1 3911 2658 3914 2662 1 GND!
rlabel metal1 4081 2724 4085 2728 1 Vdd!
rlabel metal1 3910 2724 3914 2728 1 Vdd!
rlabel metal1 3991 2724 3995 2728 1 Vdd!
rlabel metal1 3911 2790 3914 2794 1 GND!
rlabel metal1 4016 2790 4019 2794 1 GND!
rlabel metal1 3910 2856 3914 2860 1 Vdd!
rlabel metal1 3991 2856 3995 2860 1 Vdd!
rlabel metal1 4060 2827 4063 2830 7 Y
rlabel metal1 3910 2988 3914 2992 1 Vdd!
rlabel metal1 3991 2988 3995 2992 1 Vdd!
rlabel metal1 3911 2922 3914 2926 1 GND!
rlabel metal1 3992 2922 3995 2926 1 GND!
rlabel metal2 4055 2983 4058 2988 1 select_out
rlabel metal1 3710 3065 3713 3069 1 Vdd!
rlabel metal1 3711 3008 3714 3012 1 GND!
rlabel metal1 3712 3001 3715 3005 2 ~clk
rlabel metal1 3710 3072 3713 3076 4 clk
rlabel metal1 3843 3008 3846 3012 1 GND!
rlabel metal1 3844 3001 3847 3005 2 ~clk
rlabel metal1 3842 3072 3845 3076 4 clk
rlabel metal1 3974 3065 3977 3069 1 Vdd!
rlabel metal1 3975 3008 3978 3012 1 GND!
rlabel metal1 3976 3001 3979 3005 2 ~clk
rlabel metal1 3974 3072 3977 3076 4 clk
rlabel metal1 4106 3072 4109 3076 4 clk
rlabel metal1 4108 3001 4111 3005 2 ~clk
rlabel metal1 4107 3008 4110 3012 1 GND!
rlabel metal1 4106 3065 4109 3069 1 Vdd!
rlabel m3contact 3707 3038 3710 3041 3 ctrl_reg
rlabel metal2 3884 2993 3887 2998 1 select0
rlabel metal2 3967 2992 3970 2999 1 select1
rlabel metal2 4027 2992 4030 2998 1 select2
rlabel metal1 3971 2460 3975 2464 1 Vdd!
rlabel metal1 3960 2526 3964 2530 1 GND!
rlabel metal1 3961 2519 3965 2523 1 ~clk
rlabel metal1 3964 2467 3967 2471 1 clk
rlabel metal1 3842 3065 3845 3069 1 Vdd!
rlabel polysilicon 4149 2448 4149 2448 1 CB3
rlabel metal1 4009 3321 4012 3325 4 clk
rlabel metal1 4011 3250 4014 3254 2 ~clk
rlabel metal1 4010 3257 4013 3261 1 GND!
rlabel metal1 4009 3314 4012 3318 1 Vdd!
rlabel metal1 4009 3400 4012 3404 1 Vdd!
rlabel metal1 4010 3343 4013 3347 1 GND!
rlabel metal1 4011 3336 4014 3340 2 ~clk
rlabel metal1 4009 3407 4012 3411 4 clk
rlabel metal1 4009 2425 4012 2429 4 clk
rlabel metal1 4011 2354 4014 2358 2 ~clk
rlabel metal1 4010 2361 4013 2365 1 GND!
rlabel metal1 4009 2418 4012 2422 1 Vdd!
rlabel metal1 4009 2332 4012 2336 1 Vdd!
rlabel metal1 4010 2275 4013 2279 1 GND!
rlabel metal1 4011 2268 4014 2272 2 ~clk
rlabel metal1 4009 2339 4012 2343 4 clk
rlabel polysilicon 4161 2302 4161 2302 1 CB4
rlabel metal2 3695 4058 3701 4062 1 reset_b
rlabel space 4740 2533 5000 2793 1 OUT
rlabel space 3445 4741 3705 5001 1 Vdd!
rlabel space 3138 4741 3398 5001 1 GND!
rlabel space 2827 4744 3087 5004 1 MODE
rlabel space 3762 4749 3996 4987 1 RESET_b
rlabel space 2534 4752 2768 4990 1 clk
rlabel space 2223 4758 2457 4996 1 DATA
rlabel space 1912 4765 2146 5003 1 PROGRAM
<< end >>
