magic
tech scmos
timestamp 1607749400
<< ntransistor >>
rect 12 24 14 28
rect 28 24 30 28
rect 47 24 49 28
rect 70 24 72 28
rect 75 24 77 28
rect 101 24 103 28
rect 129 24 131 28
rect 149 24 151 28
rect 154 24 156 28
rect 181 24 183 28
<< ptransistor >>
rect 12 43 14 51
rect 28 43 30 51
rect 47 44 49 52
rect 70 43 72 51
rect 75 43 77 51
rect 101 43 103 51
rect 129 44 131 52
rect 149 43 151 51
rect 154 43 156 51
rect 181 43 183 51
<< ndiffusion >>
rect 11 24 12 28
rect 14 24 15 28
rect 27 24 28 28
rect 30 24 31 28
rect 46 24 47 28
rect 49 24 50 28
rect 65 24 70 28
rect 72 24 75 28
rect 77 24 78 28
rect 99 24 101 28
rect 103 24 104 28
rect 128 24 129 28
rect 131 24 132 28
rect 144 24 149 28
rect 151 24 154 28
rect 156 24 157 28
rect 180 24 181 28
rect 183 24 184 28
<< pdiffusion >>
rect 11 43 12 51
rect 14 43 15 51
rect 27 43 28 51
rect 30 43 31 51
rect 46 44 47 52
rect 49 44 50 52
rect 65 43 70 51
rect 72 43 75 51
rect 77 43 78 51
rect 99 43 101 51
rect 103 43 104 51
rect 128 44 129 52
rect 131 44 132 52
rect 144 43 149 51
rect 151 43 154 51
rect 156 43 157 51
rect 180 43 181 51
rect 183 43 184 51
<< ndcontact >>
rect 7 24 11 28
rect 15 24 19 28
rect 23 24 27 28
rect 31 24 35 28
rect 42 24 46 28
rect 50 24 54 28
rect 61 24 65 28
rect 78 24 82 28
rect 95 24 99 28
rect 104 24 108 28
rect 124 24 128 28
rect 132 24 136 28
rect 140 24 144 28
rect 157 24 161 28
rect 176 24 180 28
rect 184 24 188 28
<< pdcontact >>
rect 7 43 11 51
rect 15 43 19 51
rect 23 43 27 51
rect 31 43 35 51
rect 42 44 46 52
rect 50 44 54 52
rect 61 43 65 51
rect 78 43 82 51
rect 95 43 99 51
rect 104 43 108 51
rect 124 44 128 52
rect 132 44 136 52
rect 140 43 144 51
rect 157 43 161 51
rect 176 43 180 51
rect 184 43 188 51
<< psubstratepcontact >>
rect 0 8 4 12
rect 18 8 22 12
rect 38 8 42 12
rect 51 8 55 12
rect 87 8 91 12
rect 113 8 117 12
rect 133 8 137 12
<< nsubstratencontact >>
rect 0 61 4 65
rect 18 61 22 65
rect 38 61 42 65
rect 51 61 55 65
rect 87 61 91 65
rect 113 61 117 65
rect 133 61 137 65
<< polysilicon >>
rect 28 58 30 61
rect 75 58 77 61
rect 101 58 103 61
rect 154 58 156 61
rect 28 54 29 58
rect 101 54 102 58
rect 12 51 14 53
rect 28 51 30 54
rect 47 52 49 54
rect 70 51 72 53
rect 75 51 77 54
rect 101 51 103 54
rect 129 52 131 54
rect 12 28 14 43
rect 28 41 30 43
rect 28 28 30 30
rect 47 28 49 44
rect 149 51 151 53
rect 154 51 156 54
rect 181 51 183 53
rect 70 37 72 43
rect 75 41 77 43
rect 101 41 103 43
rect 66 33 72 37
rect 70 28 72 33
rect 75 28 77 30
rect 101 28 103 30
rect 129 28 131 44
rect 149 37 151 43
rect 154 41 156 43
rect 145 33 151 37
rect 149 28 151 33
rect 154 28 156 30
rect 181 28 183 43
rect 12 22 14 24
rect 28 20 30 24
rect 47 22 49 24
rect 70 22 72 24
rect 29 16 30 20
rect 75 19 77 24
rect 101 20 103 24
rect 129 22 131 24
rect 149 22 151 24
rect 28 13 30 16
rect 76 15 77 19
rect 102 16 103 20
rect 154 19 156 24
rect 181 22 183 24
rect 75 13 77 15
rect 101 12 103 16
rect 155 15 156 19
rect 154 13 156 15
<< polycontact >>
rect 29 54 33 58
rect 75 54 79 58
rect 102 54 106 58
rect 154 54 158 58
rect 8 33 12 37
rect 43 34 47 38
rect 62 33 66 37
rect 125 34 129 38
rect 141 33 145 37
rect 177 33 181 37
rect 25 16 29 20
rect 72 15 76 19
rect 97 16 102 20
rect 151 15 155 19
<< metal1 >>
rect 0 70 34 74
rect 38 70 64 74
rect 68 70 89 74
rect 93 70 164 74
rect 168 70 188 74
rect 4 61 18 65
rect 22 61 38 65
rect 42 61 51 65
rect 55 61 87 65
rect 91 61 113 65
rect 117 61 133 65
rect 137 61 188 65
rect 7 51 10 61
rect 33 54 34 58
rect 42 52 45 61
rect 3 33 8 36
rect 16 36 19 43
rect 23 36 26 43
rect 16 33 26 36
rect 16 28 19 33
rect 23 28 26 33
rect 32 38 35 43
rect 32 36 38 38
rect 42 36 43 38
rect 32 34 43 36
rect 51 37 54 44
rect 61 51 64 61
rect 79 54 82 58
rect 106 54 107 58
rect 124 52 127 61
rect 79 39 82 43
rect 51 35 62 37
rect 32 28 35 34
rect 51 33 57 35
rect 51 28 54 33
rect 61 33 62 35
rect 80 35 82 39
rect 79 28 82 35
rect 95 38 98 43
rect 105 38 108 43
rect 105 34 117 38
rect 121 34 125 38
rect 133 37 136 44
rect 140 51 143 61
rect 158 54 164 58
rect 176 51 179 61
rect 158 38 161 43
rect 95 28 98 34
rect 105 28 108 34
rect 133 33 134 37
rect 138 33 141 36
rect 160 34 161 38
rect 133 28 136 33
rect 158 28 161 34
rect 173 33 177 37
rect 185 28 188 43
rect 7 12 10 24
rect 24 16 25 20
rect 42 12 45 24
rect 61 12 64 24
rect 71 15 72 19
rect 96 16 97 20
rect 124 12 127 24
rect 140 12 143 24
rect 150 15 151 19
rect 176 12 179 24
rect 4 8 18 12
rect 22 8 38 12
rect 42 8 51 12
rect 55 8 87 12
rect 91 8 113 12
rect 117 8 133 12
rect 137 8 188 12
rect 0 0 20 4
rect 24 0 83 4
rect 87 0 108 4
rect 112 0 146 4
rect 150 0 188 4
<< m2contact >>
rect 34 70 38 74
rect 64 70 68 74
rect 89 70 93 74
rect 164 70 168 74
rect 34 54 38 58
rect 38 36 42 40
rect 82 54 86 58
rect 107 54 111 58
rect 57 31 61 35
rect 76 35 80 39
rect 95 34 99 38
rect 117 34 121 38
rect 164 54 168 58
rect 134 33 138 37
rect 156 34 160 38
rect 169 33 173 37
rect 20 16 24 20
rect 67 15 71 19
rect 89 16 96 20
rect 146 15 150 19
rect 20 0 24 4
rect 83 0 87 4
rect 108 0 112 4
rect 146 0 150 4
<< metal2 >>
rect 34 58 38 70
rect 20 4 24 16
rect 64 15 67 70
rect 83 4 86 54
rect 89 20 92 70
rect 164 58 168 70
rect 108 4 111 54
rect 146 4 150 15
<< m3contact >>
rect 42 35 47 40
rect 56 26 61 31
rect 71 34 76 39
rect 99 34 104 39
rect 117 38 122 43
rect 151 34 156 39
rect 135 28 140 33
rect 168 28 173 33
<< metal3 >>
rect 117 45 156 50
rect 42 41 76 45
rect 117 44 126 45
rect 134 44 156 45
rect 41 40 76 41
rect 116 43 123 44
rect 41 35 42 40
rect 47 35 48 40
rect 41 34 48 35
rect 70 39 77 40
rect 70 34 71 39
rect 76 34 77 39
rect 70 33 77 34
rect 98 39 105 40
rect 98 34 99 39
rect 104 34 105 39
rect 116 38 117 43
rect 122 38 123 43
rect 151 40 156 44
rect 116 37 123 38
rect 150 39 157 40
rect 150 34 151 39
rect 156 34 157 39
rect 98 33 105 34
rect 134 33 141 34
rect 150 33 157 34
rect 167 33 174 34
rect 55 31 62 32
rect 55 26 56 31
rect 61 30 62 31
rect 99 30 104 33
rect 61 26 104 30
rect 134 28 135 33
rect 140 28 141 33
rect 167 28 168 33
rect 173 28 174 33
rect 134 27 174 28
rect 55 25 104 26
rect 135 23 174 27
<< labels >>
rlabel metal1 3 33 7 36 1 D
rlabel metal1 0 70 3 74 4 clk
rlabel metal1 0 0 3 4 2 ~clk
rlabel metal1 7 61 10 65 1 Vdd!
rlabel metal1 8 8 11 12 1 GND!
rlabel metal1 95 36 98 39 1 test2
rlabel metal1 105 34 108 37 1 test1
rlabel metal1 185 31 188 38 7 Q
<< end >>
