magic
tech scmos
timestamp 1608257877
<< ntransistor >>
rect 14 12 16 19
<< ptransistor >>
rect 14 39 16 53
<< ndiffusion >>
rect 13 12 14 19
rect 16 12 17 19
<< pdiffusion >>
rect 13 39 14 53
rect 16 39 17 53
<< ndcontact >>
rect -3 12 13 19
rect 17 12 33 19
<< pdcontact >>
rect -3 39 13 53
rect 17 39 33 53
<< polysilicon >>
rect 14 53 16 56
rect 14 31 16 39
rect 14 19 16 27
rect 14 10 16 12
<< polycontact >>
rect 12 27 16 31
<< metal1 >>
rect -10 60 39 64
rect -3 53 0 60
rect 2 27 12 31
rect 30 19 33 39
rect -3 5 0 12
rect -13 1 36 5
<< end >>
