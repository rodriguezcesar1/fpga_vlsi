magic
tech scmos
timestamp 1605552145
<< ntransistor >>
rect 13 530 21 532
rect 62 530 66 532
rect 13 522 21 524
rect 62 522 66 524
rect 13 514 21 516
rect 62 514 66 516
rect 13 506 21 508
rect 62 506 66 508
rect 13 490 21 492
rect 62 490 66 492
rect 13 482 21 484
rect 62 482 66 484
rect 13 474 21 476
rect 62 474 66 476
rect 13 466 21 468
rect 62 466 66 468
rect 13 450 21 452
rect 62 450 66 452
rect 13 442 21 444
rect 62 442 66 444
rect 13 434 21 436
rect 62 434 66 436
rect 13 426 21 428
rect 62 426 66 428
rect 13 410 21 412
rect 62 410 66 412
rect 13 402 21 404
rect 62 402 66 404
rect 13 394 21 396
rect 62 394 66 396
rect 13 386 21 388
rect 62 386 66 388
rect 13 370 21 372
rect 62 370 66 372
rect 13 362 21 364
rect 62 362 66 364
rect 13 354 21 356
rect 62 354 66 356
rect 13 346 21 348
rect 62 346 66 348
rect 13 330 21 332
rect 62 330 66 332
rect 13 322 21 324
rect 62 322 66 324
rect 13 314 21 316
rect 62 314 66 316
rect 13 306 21 308
rect 62 306 66 308
rect 13 290 21 292
rect 62 290 66 292
rect 13 282 21 284
rect 62 282 66 284
rect 13 274 21 276
rect 62 274 66 276
rect 13 266 21 268
rect 62 266 66 268
rect 13 250 21 252
rect 62 250 66 252
rect 13 242 21 244
rect 62 242 66 244
rect 13 234 21 236
rect 62 234 66 236
rect 13 226 21 228
rect 62 226 66 228
rect 13 210 21 212
rect 62 210 66 212
rect 13 202 21 204
rect 62 202 66 204
rect 13 194 21 196
rect 62 194 66 196
rect 13 186 21 188
rect 62 186 66 188
rect 13 170 21 172
rect 62 170 66 172
rect 13 162 21 164
rect 62 162 66 164
rect 13 154 21 156
rect 62 154 66 156
rect 13 146 21 148
rect 62 146 66 148
rect 13 130 21 132
rect 62 130 66 132
rect 13 122 21 124
rect 62 122 66 124
rect 13 114 21 116
rect 62 114 66 116
rect 13 106 21 108
rect 62 106 66 108
rect 13 90 21 92
rect 62 90 66 92
rect 13 82 21 84
rect 62 82 66 84
rect 13 74 21 76
rect 62 74 66 76
rect 13 66 21 68
rect 62 66 66 68
rect 13 50 21 52
rect 62 50 66 52
rect 13 42 21 44
rect 62 42 66 44
rect 13 34 21 36
rect 62 34 66 36
rect 13 26 21 28
rect 62 26 66 28
rect 13 10 21 12
rect 62 10 66 12
rect 13 2 21 4
rect 62 2 66 4
rect 13 -6 21 -4
rect 62 -6 66 -4
rect 13 -14 21 -12
rect 62 -14 66 -12
rect 13 -30 21 -28
rect 62 -30 66 -28
rect 13 -38 21 -36
rect 62 -38 66 -36
rect 13 -46 21 -44
rect 62 -46 66 -44
rect 13 -54 21 -52
rect 62 -54 66 -52
rect 13 -70 21 -68
rect 62 -70 66 -68
rect 13 -78 21 -76
rect 62 -78 66 -76
rect 13 -86 21 -84
rect 62 -86 66 -84
rect 13 -94 21 -92
rect 62 -94 66 -92
<< ptransistor >>
rect 33 530 37 532
rect 46 530 50 532
rect 33 522 37 524
rect 46 522 50 524
rect 33 514 37 516
rect 46 514 50 516
rect 33 506 37 508
rect 46 506 50 508
rect 33 490 37 492
rect 46 490 50 492
rect 33 482 37 484
rect 46 482 50 484
rect 33 474 37 476
rect 46 474 50 476
rect 33 466 37 468
rect 46 466 50 468
rect 33 450 37 452
rect 46 450 50 452
rect 33 442 37 444
rect 46 442 50 444
rect 33 434 37 436
rect 46 434 50 436
rect 33 426 37 428
rect 46 426 50 428
rect 33 410 37 412
rect 46 410 50 412
rect 33 402 37 404
rect 46 402 50 404
rect 33 394 37 396
rect 46 394 50 396
rect 33 386 37 388
rect 46 386 50 388
rect 33 370 37 372
rect 46 370 50 372
rect 33 362 37 364
rect 46 362 50 364
rect 33 354 37 356
rect 46 354 50 356
rect 33 346 37 348
rect 46 346 50 348
rect 33 330 37 332
rect 46 330 50 332
rect 33 322 37 324
rect 46 322 50 324
rect 33 314 37 316
rect 46 314 50 316
rect 33 306 37 308
rect 46 306 50 308
rect 33 290 37 292
rect 46 290 50 292
rect 33 282 37 284
rect 46 282 50 284
rect 33 274 37 276
rect 46 274 50 276
rect 33 266 37 268
rect 46 266 50 268
rect 33 250 37 252
rect 46 250 50 252
rect 33 242 37 244
rect 46 242 50 244
rect 33 234 37 236
rect 46 234 50 236
rect 33 226 37 228
rect 46 226 50 228
rect 33 210 37 212
rect 46 210 50 212
rect 33 202 37 204
rect 46 202 50 204
rect 33 194 37 196
rect 46 194 50 196
rect 33 186 37 188
rect 46 186 50 188
rect 33 170 37 172
rect 46 170 50 172
rect 33 162 37 164
rect 46 162 50 164
rect 33 154 37 156
rect 46 154 50 156
rect 33 146 37 148
rect 46 146 50 148
rect 33 130 37 132
rect 46 130 50 132
rect 33 122 37 124
rect 46 122 50 124
rect 33 114 37 116
rect 46 114 50 116
rect 33 106 37 108
rect 46 106 50 108
rect 33 90 37 92
rect 46 90 50 92
rect 33 82 37 84
rect 46 82 50 84
rect 33 74 37 76
rect 46 74 50 76
rect 33 66 37 68
rect 46 66 50 68
rect 33 50 37 52
rect 46 50 50 52
rect 33 42 37 44
rect 46 42 50 44
rect 33 34 37 36
rect 46 34 50 36
rect 33 26 37 28
rect 46 26 50 28
rect 33 10 37 12
rect 46 10 50 12
rect 33 2 37 4
rect 46 2 50 4
rect 33 -6 37 -4
rect 46 -6 50 -4
rect 33 -14 37 -12
rect 46 -14 50 -12
rect 33 -30 37 -28
rect 46 -30 50 -28
rect 33 -38 37 -36
rect 46 -38 50 -36
rect 33 -46 37 -44
rect 46 -46 50 -44
rect 33 -54 37 -52
rect 46 -54 50 -52
rect 33 -70 37 -68
rect 46 -70 50 -68
rect 33 -78 37 -76
rect 46 -78 50 -76
rect 33 -86 37 -84
rect 46 -86 50 -84
rect 33 -94 37 -92
rect 46 -94 50 -92
<< ndiffusion >>
rect 13 532 21 533
rect 62 532 66 533
rect 13 524 21 530
rect 62 529 66 530
rect 62 524 66 525
rect 13 516 21 522
rect 62 521 66 522
rect 62 516 66 517
rect 13 508 21 514
rect 62 513 66 514
rect 62 508 66 509
rect 13 505 21 506
rect 62 505 66 506
rect 13 492 21 493
rect 62 492 66 493
rect 13 484 21 490
rect 62 489 66 490
rect 62 484 66 485
rect 13 476 21 482
rect 62 481 66 482
rect 62 476 66 477
rect 13 468 21 474
rect 62 473 66 474
rect 62 468 66 469
rect 13 465 21 466
rect 62 465 66 466
rect 13 452 21 453
rect 62 452 66 453
rect 13 444 21 450
rect 62 449 66 450
rect 62 444 66 445
rect 13 436 21 442
rect 62 441 66 442
rect 62 436 66 437
rect 13 428 21 434
rect 62 433 66 434
rect 62 428 66 429
rect 13 425 21 426
rect 62 425 66 426
rect 13 412 21 413
rect 62 412 66 413
rect 13 404 21 410
rect 62 409 66 410
rect 62 404 66 405
rect 13 396 21 402
rect 62 401 66 402
rect 62 396 66 397
rect 13 388 21 394
rect 62 393 66 394
rect 62 388 66 389
rect 13 385 21 386
rect 62 385 66 386
rect 13 372 21 373
rect 62 372 66 373
rect 13 364 21 370
rect 62 369 66 370
rect 62 364 66 365
rect 13 356 21 362
rect 62 361 66 362
rect 62 356 66 357
rect 13 348 21 354
rect 62 353 66 354
rect 62 348 66 349
rect 13 345 21 346
rect 62 345 66 346
rect 13 332 21 333
rect 62 332 66 333
rect 13 324 21 330
rect 62 329 66 330
rect 62 324 66 325
rect 13 316 21 322
rect 62 321 66 322
rect 62 316 66 317
rect 13 308 21 314
rect 62 313 66 314
rect 62 308 66 309
rect 13 305 21 306
rect 62 305 66 306
rect 13 292 21 293
rect 62 292 66 293
rect 13 284 21 290
rect 62 289 66 290
rect 62 284 66 285
rect 13 276 21 282
rect 62 281 66 282
rect 62 276 66 277
rect 13 268 21 274
rect 62 273 66 274
rect 62 268 66 269
rect 13 265 21 266
rect 62 265 66 266
rect 13 252 21 253
rect 62 252 66 253
rect 13 244 21 250
rect 62 249 66 250
rect 62 244 66 245
rect 13 236 21 242
rect 62 241 66 242
rect 62 236 66 237
rect 13 228 21 234
rect 62 233 66 234
rect 62 228 66 229
rect 13 225 21 226
rect 62 225 66 226
rect 13 212 21 213
rect 62 212 66 213
rect 13 204 21 210
rect 62 209 66 210
rect 62 204 66 205
rect 13 196 21 202
rect 62 201 66 202
rect 62 196 66 197
rect 13 188 21 194
rect 62 193 66 194
rect 62 188 66 189
rect 13 185 21 186
rect 62 185 66 186
rect 13 172 21 173
rect 62 172 66 173
rect 13 164 21 170
rect 62 169 66 170
rect 62 164 66 165
rect 13 156 21 162
rect 62 161 66 162
rect 62 156 66 157
rect 13 148 21 154
rect 62 153 66 154
rect 62 148 66 149
rect 13 145 21 146
rect 62 145 66 146
rect 13 132 21 133
rect 62 132 66 133
rect 13 124 21 130
rect 62 129 66 130
rect 62 124 66 125
rect 13 116 21 122
rect 62 121 66 122
rect 62 116 66 117
rect 13 108 21 114
rect 62 113 66 114
rect 62 108 66 109
rect 13 105 21 106
rect 62 105 66 106
rect 13 92 21 93
rect 62 92 66 93
rect 13 84 21 90
rect 62 89 66 90
rect 62 84 66 85
rect 13 76 21 82
rect 62 81 66 82
rect 62 76 66 77
rect 13 68 21 74
rect 62 73 66 74
rect 62 68 66 69
rect 13 65 21 66
rect 62 65 66 66
rect 13 52 21 53
rect 62 52 66 53
rect 13 44 21 50
rect 62 49 66 50
rect 62 44 66 45
rect 13 36 21 42
rect 62 41 66 42
rect 62 36 66 37
rect 13 28 21 34
rect 62 33 66 34
rect 62 28 66 29
rect 13 25 21 26
rect 62 25 66 26
rect 13 12 21 13
rect 62 12 66 13
rect 13 4 21 10
rect 62 9 66 10
rect 62 4 66 5
rect 13 -4 21 2
rect 62 1 66 2
rect 62 -4 66 -3
rect 13 -12 21 -6
rect 62 -7 66 -6
rect 62 -12 66 -11
rect 13 -15 21 -14
rect 62 -15 66 -14
rect 13 -28 21 -27
rect 62 -28 66 -27
rect 13 -36 21 -30
rect 62 -31 66 -30
rect 62 -36 66 -35
rect 13 -44 21 -38
rect 62 -39 66 -38
rect 62 -44 66 -43
rect 13 -52 21 -46
rect 62 -47 66 -46
rect 62 -52 66 -51
rect 13 -55 21 -54
rect 62 -55 66 -54
rect 13 -68 21 -67
rect 62 -68 66 -67
rect 13 -76 21 -70
rect 62 -71 66 -70
rect 62 -76 66 -75
rect 13 -84 21 -78
rect 62 -79 66 -78
rect 62 -84 66 -83
rect 13 -92 21 -86
rect 62 -87 66 -86
rect 62 -92 66 -91
rect 13 -95 21 -94
rect 62 -95 66 -94
<< pdiffusion >>
rect 33 532 37 533
rect 46 532 50 533
rect 33 529 37 530
rect 33 524 37 525
rect 46 529 50 530
rect 46 524 50 525
rect 33 521 37 522
rect 33 516 37 517
rect 46 521 50 522
rect 46 516 50 517
rect 33 513 37 514
rect 33 508 37 509
rect 46 513 50 514
rect 46 508 50 509
rect 33 505 37 506
rect 46 505 50 506
rect 33 492 37 493
rect 46 492 50 493
rect 33 489 37 490
rect 33 484 37 485
rect 46 489 50 490
rect 46 484 50 485
rect 33 481 37 482
rect 33 476 37 477
rect 46 481 50 482
rect 46 476 50 477
rect 33 473 37 474
rect 33 468 37 469
rect 46 473 50 474
rect 46 468 50 469
rect 33 465 37 466
rect 46 465 50 466
rect 33 452 37 453
rect 46 452 50 453
rect 33 449 37 450
rect 33 444 37 445
rect 46 449 50 450
rect 46 444 50 445
rect 33 441 37 442
rect 33 436 37 437
rect 46 441 50 442
rect 46 436 50 437
rect 33 433 37 434
rect 33 428 37 429
rect 46 433 50 434
rect 46 428 50 429
rect 33 425 37 426
rect 46 425 50 426
rect 33 412 37 413
rect 46 412 50 413
rect 33 409 37 410
rect 33 404 37 405
rect 46 409 50 410
rect 46 404 50 405
rect 33 401 37 402
rect 33 396 37 397
rect 46 401 50 402
rect 46 396 50 397
rect 33 393 37 394
rect 33 388 37 389
rect 46 393 50 394
rect 46 388 50 389
rect 33 385 37 386
rect 46 385 50 386
rect 33 372 37 373
rect 46 372 50 373
rect 33 369 37 370
rect 33 364 37 365
rect 46 369 50 370
rect 46 364 50 365
rect 33 361 37 362
rect 33 356 37 357
rect 46 361 50 362
rect 46 356 50 357
rect 33 353 37 354
rect 33 348 37 349
rect 46 353 50 354
rect 46 348 50 349
rect 33 345 37 346
rect 46 345 50 346
rect 33 332 37 333
rect 46 332 50 333
rect 33 329 37 330
rect 33 324 37 325
rect 46 329 50 330
rect 46 324 50 325
rect 33 321 37 322
rect 33 316 37 317
rect 46 321 50 322
rect 46 316 50 317
rect 33 313 37 314
rect 33 308 37 309
rect 46 313 50 314
rect 46 308 50 309
rect 33 305 37 306
rect 46 305 50 306
rect 33 292 37 293
rect 46 292 50 293
rect 33 289 37 290
rect 33 284 37 285
rect 46 289 50 290
rect 46 284 50 285
rect 33 281 37 282
rect 33 276 37 277
rect 46 281 50 282
rect 46 276 50 277
rect 33 273 37 274
rect 33 268 37 269
rect 46 273 50 274
rect 46 268 50 269
rect 33 265 37 266
rect 46 265 50 266
rect 33 252 37 253
rect 46 252 50 253
rect 33 249 37 250
rect 33 244 37 245
rect 46 249 50 250
rect 46 244 50 245
rect 33 241 37 242
rect 33 236 37 237
rect 46 241 50 242
rect 46 236 50 237
rect 33 233 37 234
rect 33 228 37 229
rect 46 233 50 234
rect 46 228 50 229
rect 33 225 37 226
rect 46 225 50 226
rect 33 212 37 213
rect 46 212 50 213
rect 33 209 37 210
rect 33 204 37 205
rect 46 209 50 210
rect 46 204 50 205
rect 33 201 37 202
rect 33 196 37 197
rect 46 201 50 202
rect 46 196 50 197
rect 33 193 37 194
rect 33 188 37 189
rect 46 193 50 194
rect 46 188 50 189
rect 33 185 37 186
rect 46 185 50 186
rect 33 172 37 173
rect 46 172 50 173
rect 33 169 37 170
rect 33 164 37 165
rect 46 169 50 170
rect 46 164 50 165
rect 33 161 37 162
rect 33 156 37 157
rect 46 161 50 162
rect 46 156 50 157
rect 33 153 37 154
rect 33 148 37 149
rect 46 153 50 154
rect 46 148 50 149
rect 33 145 37 146
rect 46 145 50 146
rect 33 132 37 133
rect 46 132 50 133
rect 33 129 37 130
rect 33 124 37 125
rect 46 129 50 130
rect 46 124 50 125
rect 33 121 37 122
rect 33 116 37 117
rect 46 121 50 122
rect 46 116 50 117
rect 33 113 37 114
rect 33 108 37 109
rect 46 113 50 114
rect 46 108 50 109
rect 33 105 37 106
rect 46 105 50 106
rect 33 92 37 93
rect 46 92 50 93
rect 33 89 37 90
rect 33 84 37 85
rect 46 89 50 90
rect 46 84 50 85
rect 33 81 37 82
rect 33 76 37 77
rect 46 81 50 82
rect 46 76 50 77
rect 33 73 37 74
rect 33 68 37 69
rect 46 73 50 74
rect 46 68 50 69
rect 33 65 37 66
rect 46 65 50 66
rect 33 52 37 53
rect 46 52 50 53
rect 33 49 37 50
rect 33 44 37 45
rect 46 49 50 50
rect 46 44 50 45
rect 33 41 37 42
rect 33 36 37 37
rect 46 41 50 42
rect 46 36 50 37
rect 33 33 37 34
rect 33 28 37 29
rect 46 33 50 34
rect 46 28 50 29
rect 33 25 37 26
rect 46 25 50 26
rect 33 12 37 13
rect 46 12 50 13
rect 33 9 37 10
rect 33 4 37 5
rect 46 9 50 10
rect 46 4 50 5
rect 33 1 37 2
rect 33 -4 37 -3
rect 46 1 50 2
rect 46 -4 50 -3
rect 33 -7 37 -6
rect 33 -12 37 -11
rect 46 -7 50 -6
rect 46 -12 50 -11
rect 33 -15 37 -14
rect 46 -15 50 -14
rect 33 -28 37 -27
rect 46 -28 50 -27
rect 33 -31 37 -30
rect 33 -36 37 -35
rect 46 -31 50 -30
rect 46 -36 50 -35
rect 33 -39 37 -38
rect 33 -44 37 -43
rect 46 -39 50 -38
rect 46 -44 50 -43
rect 33 -47 37 -46
rect 33 -52 37 -51
rect 46 -47 50 -46
rect 46 -52 50 -51
rect 33 -55 37 -54
rect 46 -55 50 -54
rect 33 -68 37 -67
rect 46 -68 50 -67
rect 33 -71 37 -70
rect 33 -76 37 -75
rect 46 -71 50 -70
rect 46 -76 50 -75
rect 33 -79 37 -78
rect 33 -84 37 -83
rect 46 -79 50 -78
rect 46 -84 50 -83
rect 33 -87 37 -86
rect 33 -92 37 -91
rect 46 -87 50 -86
rect 46 -92 50 -91
rect 33 -95 37 -94
rect 46 -95 50 -94
<< ndcontact >>
rect 13 533 21 537
rect 62 533 66 537
rect 62 525 66 529
rect 62 517 66 521
rect 62 509 66 513
rect 13 501 21 505
rect 62 501 66 505
rect 13 493 21 497
rect 62 493 66 497
rect 62 485 66 489
rect 62 477 66 481
rect 62 469 66 473
rect 13 461 21 465
rect 62 461 66 465
rect 13 453 21 457
rect 62 453 66 457
rect 62 445 66 449
rect 62 437 66 441
rect 62 429 66 433
rect 13 421 21 425
rect 62 421 66 425
rect 13 413 21 417
rect 62 413 66 417
rect 62 405 66 409
rect 62 397 66 401
rect 62 389 66 393
rect 13 381 21 385
rect 62 381 66 385
rect 13 373 21 377
rect 62 373 66 377
rect 62 365 66 369
rect 62 357 66 361
rect 62 349 66 353
rect 13 341 21 345
rect 62 341 66 345
rect 13 333 21 337
rect 62 333 66 337
rect 62 325 66 329
rect 62 317 66 321
rect 62 309 66 313
rect 13 301 21 305
rect 62 301 66 305
rect 13 293 21 297
rect 62 293 66 297
rect 62 285 66 289
rect 62 277 66 281
rect 62 269 66 273
rect 13 261 21 265
rect 62 261 66 265
rect 13 253 21 257
rect 62 253 66 257
rect 62 245 66 249
rect 62 237 66 241
rect 62 229 66 233
rect 13 221 21 225
rect 62 221 66 225
rect 13 213 21 217
rect 62 213 66 217
rect 62 205 66 209
rect 62 197 66 201
rect 62 189 66 193
rect 13 181 21 185
rect 62 181 66 185
rect 13 173 21 177
rect 62 173 66 177
rect 62 165 66 169
rect 62 157 66 161
rect 62 149 66 153
rect 13 141 21 145
rect 62 141 66 145
rect 13 133 21 137
rect 62 133 66 137
rect 62 125 66 129
rect 62 117 66 121
rect 62 109 66 113
rect 13 101 21 105
rect 62 101 66 105
rect 13 93 21 97
rect 62 93 66 97
rect 62 85 66 89
rect 62 77 66 81
rect 62 69 66 73
rect 13 61 21 65
rect 62 61 66 65
rect 13 53 21 57
rect 62 53 66 57
rect 62 45 66 49
rect 62 37 66 41
rect 62 29 66 33
rect 13 21 21 25
rect 62 21 66 25
rect 13 13 21 17
rect 62 13 66 17
rect 62 5 66 9
rect 62 -3 66 1
rect 62 -11 66 -7
rect 13 -19 21 -15
rect 62 -19 66 -15
rect 13 -27 21 -23
rect 62 -27 66 -23
rect 62 -35 66 -31
rect 62 -43 66 -39
rect 62 -51 66 -47
rect 13 -59 21 -55
rect 62 -59 66 -55
rect 13 -67 21 -63
rect 62 -67 66 -63
rect 62 -75 66 -71
rect 62 -83 66 -79
rect 62 -91 66 -87
rect 13 -99 21 -95
rect 62 -99 66 -95
<< pdcontact >>
rect 33 533 37 537
rect 46 533 50 537
rect 33 525 37 529
rect 46 525 50 529
rect 33 517 37 521
rect 46 517 50 521
rect 33 509 37 513
rect 46 509 50 513
rect 33 501 37 505
rect 46 501 50 505
rect 33 493 37 497
rect 46 493 50 497
rect 33 485 37 489
rect 46 485 50 489
rect 33 477 37 481
rect 46 477 50 481
rect 33 469 37 473
rect 46 469 50 473
rect 33 461 37 465
rect 46 461 50 465
rect 33 453 37 457
rect 46 453 50 457
rect 33 445 37 449
rect 46 445 50 449
rect 33 437 37 441
rect 46 437 50 441
rect 33 429 37 433
rect 46 429 50 433
rect 33 421 37 425
rect 46 421 50 425
rect 33 413 37 417
rect 46 413 50 417
rect 33 405 37 409
rect 46 405 50 409
rect 33 397 37 401
rect 46 397 50 401
rect 33 389 37 393
rect 46 389 50 393
rect 33 381 37 385
rect 46 381 50 385
rect 33 373 37 377
rect 46 373 50 377
rect 33 365 37 369
rect 46 365 50 369
rect 33 357 37 361
rect 46 357 50 361
rect 33 349 37 353
rect 46 349 50 353
rect 33 341 37 345
rect 46 341 50 345
rect 33 333 37 337
rect 46 333 50 337
rect 33 325 37 329
rect 46 325 50 329
rect 33 317 37 321
rect 46 317 50 321
rect 33 309 37 313
rect 46 309 50 313
rect 33 301 37 305
rect 46 301 50 305
rect 33 293 37 297
rect 46 293 50 297
rect 33 285 37 289
rect 46 285 50 289
rect 33 277 37 281
rect 46 277 50 281
rect 33 269 37 273
rect 46 269 50 273
rect 33 261 37 265
rect 46 261 50 265
rect 33 253 37 257
rect 46 253 50 257
rect 33 245 37 249
rect 46 245 50 249
rect 33 237 37 241
rect 46 237 50 241
rect 33 229 37 233
rect 46 229 50 233
rect 33 221 37 225
rect 46 221 50 225
rect 33 213 37 217
rect 46 213 50 217
rect 33 205 37 209
rect 46 205 50 209
rect 33 197 37 201
rect 46 197 50 201
rect 33 189 37 193
rect 46 189 50 193
rect 33 181 37 185
rect 46 181 50 185
rect 33 173 37 177
rect 46 173 50 177
rect 33 165 37 169
rect 46 165 50 169
rect 33 157 37 161
rect 46 157 50 161
rect 33 149 37 153
rect 46 149 50 153
rect 33 141 37 145
rect 46 141 50 145
rect 33 133 37 137
rect 46 133 50 137
rect 33 125 37 129
rect 46 125 50 129
rect 33 117 37 121
rect 46 117 50 121
rect 33 109 37 113
rect 46 109 50 113
rect 33 101 37 105
rect 46 101 50 105
rect 33 93 37 97
rect 46 93 50 97
rect 33 85 37 89
rect 46 85 50 89
rect 33 77 37 81
rect 46 77 50 81
rect 33 69 37 73
rect 46 69 50 73
rect 33 61 37 65
rect 46 61 50 65
rect 33 53 37 57
rect 46 53 50 57
rect 33 45 37 49
rect 46 45 50 49
rect 33 37 37 41
rect 46 37 50 41
rect 33 29 37 33
rect 46 29 50 33
rect 33 21 37 25
rect 46 21 50 25
rect 33 13 37 17
rect 46 13 50 17
rect 33 5 37 9
rect 46 5 50 9
rect 33 -3 37 1
rect 46 -3 50 1
rect 33 -11 37 -7
rect 46 -11 50 -7
rect 33 -19 37 -15
rect 46 -19 50 -15
rect 33 -27 37 -23
rect 46 -27 50 -23
rect 33 -35 37 -31
rect 46 -35 50 -31
rect 33 -43 37 -39
rect 46 -43 50 -39
rect 33 -51 37 -47
rect 46 -51 50 -47
rect 33 -59 37 -55
rect 46 -59 50 -55
rect 33 -67 37 -63
rect 46 -67 50 -63
rect 33 -75 37 -71
rect 46 -75 50 -71
rect 33 -83 37 -79
rect 46 -83 50 -79
rect 33 -91 37 -87
rect 46 -91 50 -87
rect 33 -99 37 -95
rect 46 -99 50 -95
<< polysilicon >>
rect -45 530 13 532
rect 21 530 33 532
rect 37 530 39 532
rect 44 530 46 532
rect 50 530 62 532
rect 66 530 68 532
rect 51 524 53 530
rect -31 522 13 524
rect 21 522 33 524
rect 37 522 39 524
rect 44 522 46 524
rect 50 522 62 524
rect 66 522 68 524
rect 51 516 53 522
rect -17 514 13 516
rect 21 514 33 516
rect 37 514 39 516
rect 44 514 46 516
rect 50 514 62 516
rect 66 514 68 516
rect 51 508 53 514
rect -3 506 13 508
rect 21 506 33 508
rect 37 506 39 508
rect 44 506 46 508
rect 50 506 62 508
rect 66 506 68 508
rect 51 500 53 506
rect 29 498 53 500
rect -45 490 13 492
rect 21 490 33 492
rect 37 490 39 492
rect 44 490 46 492
rect 50 490 62 492
rect 66 490 68 492
rect 51 484 53 490
rect -31 482 13 484
rect 21 482 33 484
rect 37 482 39 484
rect 44 482 46 484
rect 50 482 62 484
rect 66 482 68 484
rect 51 476 53 482
rect -17 474 13 476
rect 21 474 33 476
rect 37 474 39 476
rect 44 474 46 476
rect 50 474 62 476
rect 66 474 68 476
rect 51 468 53 474
rect 4 466 13 468
rect 21 466 33 468
rect 37 466 39 468
rect 44 466 46 468
rect 50 466 62 468
rect 66 466 68 468
rect 51 460 53 466
rect 29 458 53 460
rect -45 450 13 452
rect 21 450 33 452
rect 37 450 39 452
rect 44 450 46 452
rect 50 450 62 452
rect 66 450 68 452
rect 51 444 53 450
rect -31 442 13 444
rect 21 442 33 444
rect 37 442 39 444
rect 44 442 46 444
rect 50 442 62 444
rect 66 442 68 444
rect 51 436 53 442
rect -10 434 13 436
rect 21 434 33 436
rect 37 434 39 436
rect 44 434 46 436
rect 50 434 62 436
rect 66 434 68 436
rect 51 428 53 434
rect -3 426 13 428
rect 21 426 33 428
rect 37 426 39 428
rect 44 426 46 428
rect 50 426 62 428
rect 66 426 68 428
rect 51 420 53 426
rect 29 418 53 420
rect -45 410 13 412
rect 21 410 33 412
rect 37 410 39 412
rect 44 410 46 412
rect 50 410 62 412
rect 66 410 68 412
rect 51 404 53 410
rect -31 402 13 404
rect 21 402 33 404
rect 37 402 39 404
rect 44 402 46 404
rect 50 402 62 404
rect 66 402 68 404
rect 51 396 53 402
rect -10 394 13 396
rect 21 394 33 396
rect 37 394 39 396
rect 44 394 46 396
rect 50 394 62 396
rect 66 394 68 396
rect 51 388 53 394
rect 4 386 13 388
rect 21 386 33 388
rect 37 386 39 388
rect 44 386 46 388
rect 50 386 62 388
rect 66 386 68 388
rect 51 380 53 386
rect 29 378 53 380
rect -45 370 13 372
rect 21 370 33 372
rect 37 370 39 372
rect 44 370 46 372
rect 50 370 62 372
rect 66 370 68 372
rect 51 364 53 370
rect -24 362 13 364
rect 21 362 33 364
rect 37 362 39 364
rect 44 362 46 364
rect 50 362 62 364
rect 66 362 68 364
rect 51 356 53 362
rect -17 354 13 356
rect 21 354 33 356
rect 37 354 39 356
rect 44 354 46 356
rect 50 354 62 356
rect 66 354 68 356
rect 51 348 53 354
rect -3 346 13 348
rect 21 346 33 348
rect 37 346 39 348
rect 44 346 46 348
rect 50 346 62 348
rect 66 346 68 348
rect 51 340 53 346
rect 29 338 53 340
rect -45 330 13 332
rect 21 330 33 332
rect 37 330 39 332
rect 44 330 46 332
rect 50 330 62 332
rect 66 330 68 332
rect 51 324 53 330
rect -24 322 13 324
rect 21 322 33 324
rect 37 322 39 324
rect 44 322 46 324
rect 50 322 62 324
rect 66 322 68 324
rect 51 316 53 322
rect -17 314 13 316
rect 21 314 33 316
rect 37 314 39 316
rect 44 314 46 316
rect 50 314 62 316
rect 66 314 68 316
rect 51 308 53 314
rect 4 306 13 308
rect 21 306 33 308
rect 37 306 39 308
rect 44 306 46 308
rect 50 306 62 308
rect 66 306 68 308
rect 51 300 53 306
rect 29 298 53 300
rect -45 290 13 292
rect 21 290 33 292
rect 37 290 39 292
rect 44 290 46 292
rect 50 290 62 292
rect 66 290 68 292
rect 51 284 53 290
rect -24 282 13 284
rect 21 282 33 284
rect 37 282 39 284
rect 44 282 46 284
rect 50 282 62 284
rect 66 282 68 284
rect 51 276 53 282
rect -10 274 13 276
rect 21 274 33 276
rect 37 274 39 276
rect 44 274 46 276
rect 50 274 62 276
rect 66 274 68 276
rect 51 268 53 274
rect -3 266 13 268
rect 21 266 33 268
rect 37 266 39 268
rect 44 266 46 268
rect 50 266 62 268
rect 66 266 68 268
rect 51 260 53 266
rect 29 258 53 260
rect -45 250 13 252
rect 21 250 33 252
rect 37 250 39 252
rect 44 250 46 252
rect 50 250 62 252
rect 66 250 68 252
rect 51 244 53 250
rect -24 242 13 244
rect 21 242 33 244
rect 37 242 39 244
rect 44 242 46 244
rect 50 242 62 244
rect 66 242 68 244
rect 51 236 53 242
rect -10 234 13 236
rect 21 234 33 236
rect 37 234 39 236
rect 44 234 46 236
rect 50 234 62 236
rect 66 234 68 236
rect 51 228 53 234
rect 4 226 13 228
rect 21 226 33 228
rect 37 226 39 228
rect 44 226 46 228
rect 50 226 62 228
rect 66 226 68 228
rect 51 220 53 226
rect 29 218 53 220
rect -38 210 13 212
rect 21 210 33 212
rect 37 210 39 212
rect 44 210 46 212
rect 50 210 62 212
rect 66 210 68 212
rect 51 204 53 210
rect -31 202 13 204
rect 21 202 33 204
rect 37 202 39 204
rect 44 202 46 204
rect 50 202 62 204
rect 66 202 68 204
rect 51 196 53 202
rect -17 194 13 196
rect 21 194 33 196
rect 37 194 39 196
rect 44 194 46 196
rect 50 194 62 196
rect 66 194 68 196
rect 51 188 53 194
rect -3 186 13 188
rect 21 186 33 188
rect 37 186 39 188
rect 44 186 46 188
rect 50 186 62 188
rect 66 186 68 188
rect 51 180 53 186
rect 29 178 53 180
rect -38 170 13 172
rect 21 170 33 172
rect 37 170 39 172
rect 44 170 46 172
rect 50 170 62 172
rect 66 170 68 172
rect 51 164 53 170
rect -31 162 13 164
rect 21 162 33 164
rect 37 162 39 164
rect 44 162 46 164
rect 50 162 62 164
rect 66 162 68 164
rect 51 156 53 162
rect -17 154 13 156
rect 21 154 33 156
rect 37 154 39 156
rect 44 154 46 156
rect 50 154 62 156
rect 66 154 68 156
rect 51 148 53 154
rect 4 146 13 148
rect 21 146 33 148
rect 37 146 39 148
rect 44 146 46 148
rect 50 146 62 148
rect 66 146 68 148
rect 51 140 53 146
rect 29 138 53 140
rect -38 130 13 132
rect 21 130 33 132
rect 37 130 39 132
rect 44 130 46 132
rect 50 130 62 132
rect 66 130 68 132
rect 51 124 53 130
rect -31 122 13 124
rect 21 122 33 124
rect 37 122 39 124
rect 44 122 46 124
rect 50 122 62 124
rect 66 122 68 124
rect 51 116 53 122
rect -10 114 13 116
rect 21 114 33 116
rect 37 114 39 116
rect 44 114 46 116
rect 50 114 62 116
rect 66 114 68 116
rect 51 108 53 114
rect -3 106 13 108
rect 21 106 33 108
rect 37 106 39 108
rect 44 106 46 108
rect 50 106 62 108
rect 66 106 68 108
rect 51 100 53 106
rect 29 98 53 100
rect -38 90 13 92
rect 21 90 33 92
rect 37 90 39 92
rect 44 90 46 92
rect 50 90 62 92
rect 66 90 68 92
rect 51 84 53 90
rect -31 82 13 84
rect 21 82 33 84
rect 37 82 39 84
rect 44 82 46 84
rect 50 82 62 84
rect 66 82 68 84
rect 51 76 53 82
rect -10 74 13 76
rect 21 74 33 76
rect 37 74 39 76
rect 44 74 46 76
rect 50 74 62 76
rect 66 74 68 76
rect 51 68 53 74
rect 4 66 13 68
rect 21 66 33 68
rect 37 66 39 68
rect 44 66 46 68
rect 50 66 62 68
rect 66 66 68 68
rect 51 60 53 66
rect 29 58 53 60
rect -38 50 13 52
rect 21 50 33 52
rect 37 50 39 52
rect 44 50 46 52
rect 50 50 62 52
rect 66 50 68 52
rect 51 44 53 50
rect -24 42 13 44
rect 21 42 33 44
rect 37 42 39 44
rect 44 42 46 44
rect 50 42 62 44
rect 66 42 68 44
rect 51 36 53 42
rect -17 34 13 36
rect 21 34 33 36
rect 37 34 39 36
rect 44 34 46 36
rect 50 34 62 36
rect 66 34 68 36
rect 51 28 53 34
rect -3 26 13 28
rect 21 26 33 28
rect 37 26 39 28
rect 44 26 46 28
rect 50 26 62 28
rect 66 26 68 28
rect 51 20 53 26
rect 29 18 53 20
rect -38 10 13 12
rect 21 10 33 12
rect 37 10 39 12
rect 44 10 46 12
rect 50 10 62 12
rect 66 10 68 12
rect 51 4 53 10
rect -24 2 13 4
rect 21 2 33 4
rect 37 2 39 4
rect 44 2 46 4
rect 50 2 62 4
rect 66 2 68 4
rect 51 -4 53 2
rect -17 -6 13 -4
rect 21 -6 33 -4
rect 37 -6 39 -4
rect 44 -6 46 -4
rect 50 -6 62 -4
rect 66 -6 68 -4
rect 51 -12 53 -6
rect 4 -14 13 -12
rect 21 -14 33 -12
rect 37 -14 39 -12
rect 44 -14 46 -12
rect 50 -14 62 -12
rect 66 -14 68 -12
rect 51 -20 53 -14
rect 29 -22 53 -20
rect -38 -30 13 -28
rect 21 -30 33 -28
rect 37 -30 39 -28
rect 44 -30 46 -28
rect 50 -30 62 -28
rect 66 -30 68 -28
rect 51 -36 53 -30
rect -24 -38 13 -36
rect 21 -38 33 -36
rect 37 -38 39 -36
rect 44 -38 46 -36
rect 50 -38 62 -36
rect 66 -38 68 -36
rect 51 -44 53 -38
rect -10 -46 13 -44
rect 21 -46 33 -44
rect 37 -46 39 -44
rect 44 -46 46 -44
rect 50 -46 62 -44
rect 66 -46 68 -44
rect 51 -52 53 -46
rect -3 -54 13 -52
rect 21 -54 33 -52
rect 37 -54 39 -52
rect 44 -54 46 -52
rect 50 -54 62 -52
rect 66 -54 68 -52
rect 51 -60 53 -54
rect 29 -62 53 -60
rect -38 -70 13 -68
rect 21 -70 33 -68
rect 37 -70 39 -68
rect 44 -70 46 -68
rect 50 -70 62 -68
rect 66 -70 68 -68
rect 51 -76 53 -70
rect -24 -78 13 -76
rect 21 -78 33 -76
rect 37 -78 39 -76
rect 44 -78 46 -76
rect 50 -78 62 -76
rect 66 -78 68 -76
rect 51 -84 53 -78
rect -10 -86 13 -84
rect 21 -86 33 -84
rect 37 -86 39 -84
rect 44 -86 46 -84
rect 50 -86 62 -84
rect 66 -86 68 -84
rect 51 -92 53 -86
rect 4 -94 13 -92
rect 21 -94 33 -92
rect 37 -94 39 -92
rect 44 -94 46 -92
rect 50 -94 62 -92
rect 66 -94 68 -92
rect 51 -100 53 -94
rect 29 -102 53 -100
<< polycontact >>
rect -49 529 -45 533
rect -35 521 -31 525
rect -21 513 -17 517
rect -7 505 -3 509
rect 25 497 29 501
rect -49 489 -45 493
rect -35 481 -31 485
rect -21 473 -17 477
rect 0 465 4 469
rect 25 457 29 461
rect -49 449 -45 453
rect -35 441 -31 445
rect -14 433 -10 437
rect -7 425 -3 429
rect 25 417 29 421
rect -49 409 -45 413
rect -35 401 -31 405
rect -14 393 -10 397
rect 0 385 4 389
rect 25 377 29 381
rect -49 369 -45 373
rect -28 361 -24 365
rect -21 353 -17 357
rect -7 345 -3 349
rect 25 337 29 341
rect -49 329 -45 333
rect -28 321 -24 325
rect -21 313 -17 317
rect 0 305 4 309
rect 25 297 29 301
rect -49 289 -45 293
rect -28 281 -24 285
rect -14 273 -10 277
rect -7 265 -3 269
rect 25 257 29 261
rect -49 249 -45 253
rect -28 241 -24 245
rect -14 233 -10 237
rect 0 225 4 229
rect 25 217 29 221
rect -42 209 -38 213
rect -35 201 -31 205
rect -21 193 -17 197
rect -7 185 -3 189
rect 25 177 29 181
rect -42 169 -38 173
rect -35 161 -31 165
rect -21 153 -17 157
rect 0 145 4 149
rect 25 137 29 141
rect -42 129 -38 133
rect -35 121 -31 125
rect -14 113 -10 117
rect -7 105 -3 109
rect 25 97 29 101
rect -42 89 -38 93
rect -35 81 -31 85
rect -14 73 -10 77
rect 0 65 4 69
rect 25 57 29 61
rect -42 49 -38 53
rect -28 41 -24 45
rect -21 33 -17 37
rect -7 25 -3 29
rect 25 17 29 21
rect -42 9 -38 13
rect -28 1 -24 5
rect -21 -7 -17 -3
rect 0 -15 4 -11
rect 25 -23 29 -19
rect -42 -31 -38 -27
rect -28 -39 -24 -35
rect -14 -47 -10 -43
rect -7 -55 -3 -51
rect 25 -63 29 -59
rect -42 -71 -38 -67
rect -28 -79 -24 -75
rect -14 -87 -10 -83
rect 0 -95 4 -91
rect 25 -103 29 -99
<< metal1 >>
rect -49 533 -45 541
rect -49 493 -45 529
rect -49 453 -45 489
rect -49 413 -45 449
rect -49 373 -45 409
rect -49 333 -45 369
rect -49 293 -45 329
rect -49 253 -45 289
rect -49 -103 -45 249
rect -42 213 -38 541
rect -42 173 -38 209
rect -42 133 -38 169
rect -42 93 -38 129
rect -42 53 -38 89
rect -42 13 -38 49
rect -42 -27 -38 9
rect -42 -67 -38 -31
rect -42 -103 -38 -71
rect -35 525 -31 541
rect -35 485 -31 521
rect -35 445 -31 481
rect -35 405 -31 441
rect -35 205 -31 401
rect -35 165 -31 201
rect -35 125 -31 161
rect -35 85 -31 121
rect -35 -103 -31 81
rect -28 365 -24 541
rect -28 325 -24 361
rect -28 285 -24 321
rect -28 245 -24 281
rect -28 45 -24 241
rect -28 5 -24 41
rect -28 -35 -24 1
rect -28 -75 -24 -39
rect -28 -103 -24 -79
rect -21 517 -17 541
rect -21 477 -17 513
rect -21 357 -17 473
rect -21 317 -17 353
rect -21 197 -17 313
rect -21 157 -17 193
rect -21 37 -17 153
rect -21 -3 -17 33
rect -21 -103 -17 -7
rect -14 437 -10 541
rect -14 397 -10 433
rect -14 277 -10 393
rect -14 237 -10 273
rect -14 117 -10 233
rect -14 77 -10 113
rect -14 -43 -10 73
rect -14 -83 -10 -47
rect -14 -103 -10 -87
rect -7 509 -3 541
rect -7 429 -3 505
rect -7 349 -3 425
rect -7 269 -3 345
rect -7 189 -3 265
rect -7 109 -3 185
rect -7 29 -3 105
rect -7 -51 -3 25
rect -7 -103 -3 -55
rect 0 469 4 541
rect 0 389 4 465
rect 0 309 4 385
rect 0 229 4 305
rect 0 149 4 225
rect 0 69 4 145
rect 0 -11 4 65
rect 0 -91 4 -15
rect 0 -103 4 -95
rect 7 537 10 541
rect 40 537 43 541
rect 69 537 72 541
rect 7 533 13 537
rect 37 533 46 537
rect 7 497 10 533
rect 25 525 33 529
rect 25 513 29 525
rect 40 521 43 533
rect 54 529 58 537
rect 66 533 72 537
rect 50 525 62 529
rect 37 517 46 521
rect 25 509 33 513
rect 25 505 29 509
rect 40 505 43 517
rect 54 513 58 525
rect 69 521 72 533
rect 66 517 72 521
rect 50 509 62 513
rect 69 505 72 517
rect 21 501 29 505
rect 37 501 46 505
rect 66 501 72 505
rect 40 497 43 501
rect 69 497 72 501
rect 7 493 13 497
rect 37 493 46 497
rect 7 457 10 493
rect 25 485 33 489
rect 25 473 29 485
rect 40 481 43 493
rect 54 489 58 497
rect 66 493 72 497
rect 50 485 62 489
rect 37 477 46 481
rect 25 469 33 473
rect 25 465 29 469
rect 40 465 43 477
rect 54 473 58 485
rect 69 481 72 493
rect 66 477 72 481
rect 50 469 62 473
rect 69 465 72 477
rect 21 461 29 465
rect 37 461 46 465
rect 66 461 72 465
rect 40 457 43 461
rect 69 457 72 461
rect 7 453 13 457
rect 37 453 46 457
rect 7 417 10 453
rect 25 445 33 449
rect 25 433 29 445
rect 40 441 43 453
rect 54 449 58 457
rect 66 453 72 457
rect 50 445 62 449
rect 37 437 46 441
rect 25 429 33 433
rect 25 425 29 429
rect 40 425 43 437
rect 54 433 58 445
rect 69 441 72 453
rect 66 437 72 441
rect 50 429 62 433
rect 69 425 72 437
rect 21 421 29 425
rect 37 421 46 425
rect 66 421 72 425
rect 40 417 43 421
rect 69 417 72 421
rect 7 413 13 417
rect 37 413 46 417
rect 7 377 10 413
rect 25 405 33 409
rect 25 393 29 405
rect 40 401 43 413
rect 54 409 58 417
rect 66 413 72 417
rect 50 405 62 409
rect 37 397 46 401
rect 25 389 33 393
rect 25 385 29 389
rect 40 385 43 397
rect 54 393 58 405
rect 69 401 72 413
rect 66 397 72 401
rect 50 389 62 393
rect 69 385 72 397
rect 21 381 29 385
rect 37 381 46 385
rect 66 381 72 385
rect 40 377 43 381
rect 69 377 72 381
rect 7 373 13 377
rect 37 373 46 377
rect 7 337 10 373
rect 25 365 33 369
rect 25 353 29 365
rect 40 361 43 373
rect 54 369 58 377
rect 66 373 72 377
rect 50 365 62 369
rect 37 357 46 361
rect 25 349 33 353
rect 25 345 29 349
rect 40 345 43 357
rect 54 353 58 365
rect 69 361 72 373
rect 66 357 72 361
rect 50 349 62 353
rect 69 345 72 357
rect 21 341 29 345
rect 37 341 46 345
rect 66 341 72 345
rect 40 337 43 341
rect 69 337 72 341
rect 7 333 13 337
rect 37 333 46 337
rect 7 297 10 333
rect 25 325 33 329
rect 25 313 29 325
rect 40 321 43 333
rect 54 329 58 337
rect 66 333 72 337
rect 50 325 62 329
rect 37 317 46 321
rect 25 309 33 313
rect 25 305 29 309
rect 40 305 43 317
rect 54 313 58 325
rect 69 321 72 333
rect 66 317 72 321
rect 50 309 62 313
rect 69 305 72 317
rect 21 301 29 305
rect 37 301 46 305
rect 66 301 72 305
rect 40 297 43 301
rect 69 297 72 301
rect 7 293 13 297
rect 37 293 46 297
rect 7 257 10 293
rect 25 285 33 289
rect 25 273 29 285
rect 40 281 43 293
rect 54 289 58 297
rect 66 293 72 297
rect 50 285 62 289
rect 37 277 46 281
rect 25 269 33 273
rect 25 265 29 269
rect 40 265 43 277
rect 54 273 58 285
rect 69 281 72 293
rect 66 277 72 281
rect 50 269 62 273
rect 69 265 72 277
rect 21 261 29 265
rect 37 261 46 265
rect 66 261 72 265
rect 40 257 43 261
rect 69 257 72 261
rect 7 253 13 257
rect 37 253 46 257
rect 7 217 10 253
rect 25 245 33 249
rect 25 233 29 245
rect 40 241 43 253
rect 54 249 58 257
rect 66 253 72 257
rect 50 245 62 249
rect 37 237 46 241
rect 25 229 33 233
rect 25 225 29 229
rect 40 225 43 237
rect 54 233 58 245
rect 69 241 72 253
rect 66 237 72 241
rect 50 229 62 233
rect 69 225 72 237
rect 21 221 29 225
rect 37 221 46 225
rect 66 221 72 225
rect 40 217 43 221
rect 69 217 72 221
rect 7 213 13 217
rect 37 213 46 217
rect 7 177 10 213
rect 25 205 33 209
rect 25 193 29 205
rect 40 201 43 213
rect 54 209 58 217
rect 66 213 72 217
rect 50 205 62 209
rect 37 197 46 201
rect 25 189 33 193
rect 25 185 29 189
rect 40 185 43 197
rect 54 193 58 205
rect 69 201 72 213
rect 66 197 72 201
rect 50 189 62 193
rect 69 185 72 197
rect 21 181 29 185
rect 37 181 46 185
rect 66 181 72 185
rect 40 177 43 181
rect 69 177 72 181
rect 7 173 13 177
rect 37 173 46 177
rect 7 137 10 173
rect 25 165 33 169
rect 25 153 29 165
rect 40 161 43 173
rect 54 169 58 177
rect 66 173 72 177
rect 50 165 62 169
rect 37 157 46 161
rect 25 149 33 153
rect 25 145 29 149
rect 40 145 43 157
rect 54 153 58 165
rect 69 161 72 173
rect 66 157 72 161
rect 50 149 62 153
rect 69 145 72 157
rect 21 141 29 145
rect 37 141 46 145
rect 66 141 72 145
rect 40 137 43 141
rect 69 137 72 141
rect 7 133 13 137
rect 37 133 46 137
rect 7 97 10 133
rect 25 125 33 129
rect 25 113 29 125
rect 40 121 43 133
rect 54 129 58 137
rect 66 133 72 137
rect 50 125 62 129
rect 37 117 46 121
rect 25 109 33 113
rect 25 105 29 109
rect 40 105 43 117
rect 54 113 58 125
rect 69 121 72 133
rect 66 117 72 121
rect 50 109 62 113
rect 69 105 72 117
rect 21 101 29 105
rect 37 101 46 105
rect 66 101 72 105
rect 40 97 43 101
rect 69 97 72 101
rect 7 93 13 97
rect 37 93 46 97
rect 7 57 10 93
rect 25 85 33 89
rect 25 73 29 85
rect 40 81 43 93
rect 54 89 58 97
rect 66 93 72 97
rect 50 85 62 89
rect 37 77 46 81
rect 25 69 33 73
rect 25 65 29 69
rect 40 65 43 77
rect 54 73 58 85
rect 69 81 72 93
rect 66 77 72 81
rect 50 69 62 73
rect 69 65 72 77
rect 21 61 29 65
rect 37 61 46 65
rect 66 61 72 65
rect 40 57 43 61
rect 69 57 72 61
rect 7 53 13 57
rect 37 53 46 57
rect 7 17 10 53
rect 25 45 33 49
rect 25 33 29 45
rect 40 41 43 53
rect 54 49 58 57
rect 66 53 72 57
rect 50 45 62 49
rect 37 37 46 41
rect 25 29 33 33
rect 25 25 29 29
rect 40 25 43 37
rect 54 33 58 45
rect 69 41 72 53
rect 66 37 72 41
rect 50 29 62 33
rect 69 25 72 37
rect 21 21 29 25
rect 37 21 46 25
rect 66 21 72 25
rect 40 17 43 21
rect 69 17 72 21
rect 7 13 13 17
rect 37 13 46 17
rect 7 -23 10 13
rect 25 5 33 9
rect 25 -7 29 5
rect 40 1 43 13
rect 54 9 58 17
rect 66 13 72 17
rect 50 5 62 9
rect 37 -3 46 1
rect 25 -11 33 -7
rect 25 -15 29 -11
rect 40 -15 43 -3
rect 54 -7 58 5
rect 69 1 72 13
rect 66 -3 72 1
rect 50 -11 62 -7
rect 69 -15 72 -3
rect 21 -19 29 -15
rect 37 -19 46 -15
rect 66 -19 72 -15
rect 40 -23 43 -19
rect 69 -23 72 -19
rect 7 -27 13 -23
rect 37 -27 46 -23
rect 7 -63 10 -27
rect 25 -35 33 -31
rect 25 -47 29 -35
rect 40 -39 43 -27
rect 54 -31 58 -23
rect 66 -27 72 -23
rect 50 -35 62 -31
rect 37 -43 46 -39
rect 25 -51 33 -47
rect 25 -55 29 -51
rect 40 -55 43 -43
rect 54 -47 58 -35
rect 69 -39 72 -27
rect 66 -43 72 -39
rect 50 -51 62 -47
rect 69 -55 72 -43
rect 21 -59 29 -55
rect 37 -59 46 -55
rect 66 -59 72 -55
rect 40 -63 43 -59
rect 69 -63 72 -59
rect 7 -67 13 -63
rect 37 -67 46 -63
rect 7 -103 10 -67
rect 25 -75 33 -71
rect 25 -87 29 -75
rect 40 -79 43 -67
rect 54 -71 58 -63
rect 66 -67 72 -63
rect 50 -75 62 -71
rect 37 -83 46 -79
rect 25 -91 33 -87
rect 25 -95 29 -91
rect 40 -95 43 -83
rect 54 -87 58 -75
rect 69 -79 72 -67
rect 66 -83 72 -79
rect 50 -91 62 -87
rect 69 -95 72 -83
rect 21 -99 29 -95
rect 37 -99 46 -95
rect 66 -99 72 -95
rect 40 -103 43 -99
rect 69 -103 72 -99
<< m2contact >>
rect 54 537 58 541
rect 54 497 58 501
rect 54 457 58 461
rect 54 417 58 421
rect 54 377 58 381
rect 54 337 58 341
rect 54 297 58 301
rect 54 257 58 261
rect 54 217 58 221
rect 54 177 58 181
rect 54 137 58 141
rect 54 97 58 101
rect 54 57 58 61
rect 54 17 58 21
rect 54 -23 58 -19
rect 54 -63 58 -59
<< metal2 >>
rect 58 537 73 541
rect 58 497 73 501
rect 58 457 73 461
rect 58 417 73 421
rect 58 377 73 381
rect 58 337 73 341
rect 58 297 73 301
rect 58 257 73 261
rect 58 217 73 221
rect 58 177 73 181
rect 58 137 73 141
rect 58 97 73 101
rect 58 57 73 61
rect 58 17 73 21
rect 58 -23 73 -19
rect 58 -63 73 -59
<< labels >>
rlabel metal1 2 -101 2 -101 1 A
rlabel metal1 8 -101 8 -101 1 GND
rlabel metal1 41 -99 41 -99 1 Vdd
rlabel metal1 70 -102 70 -102 8 GND
rlabel metal1 -5 -101 -5 -101 1 A_b
rlabel metal1 -12 -101 -12 -101 1 B
rlabel metal1 -19 -101 -19 -101 1 B_b
rlabel metal1 -26 -101 -26 -101 1 C
rlabel metal1 -32 -101 -32 -101 1 C_b
rlabel metal1 -40 -101 -40 -101 1 D
rlabel metal1 -47 -101 -47 -101 2 D_b
rlabel metal2 67 539 67 539 5 w0
rlabel metal2 67 499 67 499 1 w1
rlabel metal2 67 459 67 459 1 w2
rlabel metal2 67 419 67 419 1 w3
rlabel metal2 67 379 67 379 1 w4
rlabel metal2 67 339 67 339 1 w5
rlabel metal2 67 299 67 299 1 w6
rlabel metal2 68 259 68 259 7 w7
rlabel metal2 68 219 68 219 7 w8
rlabel metal2 68 179 68 179 7 w9
rlabel metal2 68 139 68 139 7 w10
rlabel metal2 68 99 68 99 7 w11
rlabel metal2 68 59 68 59 7 w12
rlabel metal2 68 19 68 19 7 w13
rlabel metal2 68 -21 68 -21 7 w14
rlabel metal2 68 -61 68 -61 7 w15
<< end >>
