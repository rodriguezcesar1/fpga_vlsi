magic
tech scmos
timestamp 1608146812
<< ntransistor >>
rect 7 387 9 391
rect 33 383 35 387
rect 38 383 40 387
rect 88 387 90 391
rect 114 383 116 387
rect 119 383 121 387
rect 61 379 63 383
rect -167 374 -165 378
rect -151 374 -149 378
rect -135 374 -133 378
rect -112 374 -110 378
rect -107 374 -105 378
rect -81 374 -79 378
rect -60 374 -58 378
rect -40 374 -38 378
rect -35 374 -33 378
rect -17 374 -15 378
rect 142 379 144 383
rect -167 328 -165 332
rect -151 328 -149 332
rect -135 328 -133 332
rect -112 328 -110 332
rect -107 328 -105 332
rect -81 328 -79 332
rect -60 328 -58 332
rect -40 328 -38 332
rect -35 328 -33 332
rect -17 328 -15 332
rect 33 327 35 331
rect 38 327 40 331
rect 114 327 116 331
rect 119 327 121 331
rect 33 251 35 255
rect 38 251 40 255
rect 112 255 114 259
rect 138 251 140 255
rect 143 251 145 255
rect 61 247 63 251
rect -167 242 -165 246
rect -151 242 -149 246
rect -135 242 -133 246
rect -112 242 -110 246
rect -107 242 -105 246
rect -81 242 -79 246
rect -60 242 -58 246
rect -40 242 -38 246
rect -35 242 -33 246
rect -17 242 -15 246
rect 166 247 168 251
rect -167 196 -165 200
rect -151 196 -149 200
rect -135 196 -133 200
rect -112 196 -110 200
rect -107 196 -105 200
rect -81 196 -79 200
rect -60 196 -58 200
rect -40 196 -38 200
rect -35 196 -33 200
rect -17 196 -15 200
rect 33 196 35 200
rect 38 196 40 200
rect 138 196 140 200
rect 143 196 145 200
rect 33 119 35 123
rect 38 119 40 123
rect 88 123 90 127
rect 114 119 116 123
rect 119 119 121 123
rect 178 123 180 127
rect 204 119 206 123
rect 209 119 211 123
rect 61 115 63 119
rect -167 110 -165 114
rect -151 110 -149 114
rect -135 110 -133 114
rect -112 110 -110 114
rect -107 110 -105 114
rect -81 110 -79 114
rect -60 110 -58 114
rect -40 110 -38 114
rect -35 110 -33 114
rect -17 110 -15 114
rect 142 115 144 119
rect 232 115 234 119
rect -167 64 -165 68
rect -151 64 -149 68
rect -135 64 -133 68
rect -112 64 -110 68
rect -107 64 -105 68
rect -81 64 -79 68
rect -60 64 -58 68
rect -40 64 -38 68
rect -35 64 -33 68
rect -17 64 -15 68
rect 33 61 35 65
rect 38 61 40 65
rect 114 61 116 65
rect 119 61 121 65
rect 204 61 206 65
rect 209 61 211 65
rect 33 -13 35 -9
rect 38 -13 40 -9
rect 61 -17 63 -13
rect -167 -22 -165 -18
rect -151 -22 -149 -18
rect -135 -22 -133 -18
rect -112 -22 -110 -18
rect -107 -22 -105 -18
rect -81 -22 -79 -18
rect -60 -22 -58 -18
rect -40 -22 -38 -18
rect -35 -22 -33 -18
rect -17 -22 -15 -18
rect -167 -68 -165 -64
rect -151 -68 -149 -64
rect -135 -68 -133 -64
rect -112 -68 -110 -64
rect -107 -68 -105 -64
rect -81 -68 -79 -64
rect -60 -68 -58 -64
rect -40 -68 -38 -64
rect -35 -68 -33 -64
rect -17 -68 -15 -64
rect 67 -68 69 -64
rect 85 -68 87 -64
rect 101 -68 103 -64
rect 117 -68 119 -64
rect 140 -68 142 -64
rect 145 -68 147 -64
rect 171 -68 173 -64
rect 192 -68 194 -64
rect 212 -68 214 -64
rect 217 -68 219 -64
rect 235 -68 237 -64
rect 33 -75 35 -71
rect 38 -75 40 -71
<< ptransistor >>
rect 7 405 9 413
rect -167 392 -165 400
rect -151 392 -149 400
rect -135 392 -133 400
rect -112 392 -110 400
rect -107 392 -105 400
rect -81 392 -79 400
rect -60 392 -58 400
rect -40 392 -38 400
rect -35 392 -33 400
rect -17 392 -15 400
rect 33 399 35 407
rect 38 399 40 407
rect 61 405 63 413
rect 88 405 90 413
rect 114 399 116 407
rect 119 399 121 407
rect 142 405 144 413
rect -167 306 -165 314
rect -151 306 -149 314
rect -135 306 -133 314
rect -112 306 -110 314
rect -107 306 -105 314
rect -81 306 -79 314
rect -60 306 -58 314
rect -40 306 -38 314
rect -35 306 -33 314
rect -17 306 -15 314
rect 33 307 35 315
rect 38 307 40 315
rect 114 307 116 315
rect 119 307 121 315
rect -167 260 -165 268
rect -151 260 -149 268
rect -135 260 -133 268
rect -112 260 -110 268
rect -107 260 -105 268
rect -81 260 -79 268
rect -60 260 -58 268
rect -40 260 -38 268
rect -35 260 -33 268
rect -17 260 -15 268
rect 33 267 35 275
rect 38 267 40 275
rect 61 273 63 281
rect 112 273 114 281
rect 138 267 140 275
rect 143 267 145 275
rect 166 273 168 281
rect -167 174 -165 182
rect -151 174 -149 182
rect -135 174 -133 182
rect -112 174 -110 182
rect -107 174 -105 182
rect -81 174 -79 182
rect -60 174 -58 182
rect -40 174 -38 182
rect -35 174 -33 182
rect -17 174 -15 182
rect 33 176 35 184
rect 38 176 40 184
rect 138 176 140 184
rect 143 176 145 184
rect -167 128 -165 136
rect -151 128 -149 136
rect -135 128 -133 136
rect -112 128 -110 136
rect -107 128 -105 136
rect -81 128 -79 136
rect -60 128 -58 136
rect -40 128 -38 136
rect -35 128 -33 136
rect -17 128 -15 136
rect 33 135 35 143
rect 38 135 40 143
rect 61 141 63 149
rect 88 141 90 149
rect 114 135 116 143
rect 119 135 121 143
rect 142 141 144 149
rect 178 141 180 149
rect 204 135 206 143
rect 209 135 211 143
rect 232 141 234 149
rect -167 42 -165 50
rect -151 42 -149 50
rect -135 42 -133 50
rect -112 42 -110 50
rect -107 42 -105 50
rect -81 42 -79 50
rect -60 42 -58 50
rect -40 42 -38 50
rect -35 42 -33 50
rect -17 42 -15 50
rect 33 41 35 49
rect 38 41 40 49
rect 114 41 116 49
rect 119 41 121 49
rect 204 41 206 49
rect 209 41 211 49
rect -167 -4 -165 4
rect -151 -4 -149 4
rect -135 -4 -133 4
rect -112 -4 -110 4
rect -107 -4 -105 4
rect -81 -4 -79 4
rect -60 -4 -58 4
rect -40 -4 -38 4
rect -35 -4 -33 4
rect -17 -4 -15 4
rect 33 3 35 11
rect 38 3 40 11
rect 61 9 63 17
rect -167 -90 -165 -82
rect -151 -90 -149 -82
rect -135 -90 -133 -82
rect -112 -90 -110 -82
rect -107 -90 -105 -82
rect -81 -90 -79 -82
rect -60 -90 -58 -82
rect -40 -90 -38 -82
rect -35 -90 -33 -82
rect -17 -90 -15 -82
rect 33 -95 35 -87
rect 38 -95 40 -87
rect 67 -90 69 -82
rect 85 -90 87 -82
rect 101 -90 103 -82
rect 117 -90 119 -82
rect 140 -90 142 -82
rect 145 -90 147 -82
rect 171 -90 173 -82
rect 192 -90 194 -82
rect 212 -90 214 -82
rect 217 -90 219 -82
rect 235 -90 237 -82
<< ndiffusion >>
rect 6 387 7 391
rect 9 387 10 391
rect 30 383 33 387
rect 35 383 38 387
rect 40 383 41 387
rect 87 387 88 391
rect 90 387 91 391
rect 111 383 114 387
rect 116 383 119 387
rect 121 383 122 387
rect 60 379 61 383
rect 63 379 64 383
rect -168 374 -167 378
rect -165 374 -164 378
rect -152 374 -151 378
rect -149 374 -148 378
rect -136 374 -135 378
rect -133 374 -132 378
rect -117 374 -112 378
rect -110 374 -107 378
rect -105 374 -104 378
rect -83 374 -81 378
rect -79 374 -78 378
rect -61 374 -60 378
rect -58 374 -57 378
rect -45 374 -40 378
rect -38 374 -35 378
rect -33 374 -32 378
rect -18 374 -17 378
rect -15 374 -14 378
rect 141 379 142 383
rect 144 379 145 383
rect -168 328 -167 332
rect -165 328 -164 332
rect -152 328 -151 332
rect -149 328 -148 332
rect -136 328 -135 332
rect -133 328 -132 332
rect -117 328 -112 332
rect -110 328 -107 332
rect -105 328 -104 332
rect -83 328 -81 332
rect -79 328 -78 332
rect -61 328 -60 332
rect -58 328 -57 332
rect -45 328 -40 332
rect -38 328 -35 332
rect -33 328 -32 332
rect -18 328 -17 332
rect -15 328 -14 332
rect 30 327 33 331
rect 35 327 38 331
rect 40 327 41 331
rect 111 327 114 331
rect 116 327 119 331
rect 121 327 122 331
rect 30 251 33 255
rect 35 251 38 255
rect 40 251 41 255
rect 111 255 112 259
rect 114 255 115 259
rect 135 251 138 255
rect 140 251 143 255
rect 145 251 146 255
rect 60 247 61 251
rect 63 247 64 251
rect -168 242 -167 246
rect -165 242 -164 246
rect -152 242 -151 246
rect -149 242 -148 246
rect -136 242 -135 246
rect -133 242 -132 246
rect -117 242 -112 246
rect -110 242 -107 246
rect -105 242 -104 246
rect -83 242 -81 246
rect -79 242 -78 246
rect -61 242 -60 246
rect -58 242 -57 246
rect -45 242 -40 246
rect -38 242 -35 246
rect -33 242 -32 246
rect -18 242 -17 246
rect -15 242 -14 246
rect 165 247 166 251
rect 168 247 169 251
rect -168 196 -167 200
rect -165 196 -164 200
rect -152 196 -151 200
rect -149 196 -148 200
rect -136 196 -135 200
rect -133 196 -132 200
rect -117 196 -112 200
rect -110 196 -107 200
rect -105 196 -104 200
rect -83 196 -81 200
rect -79 196 -78 200
rect -61 196 -60 200
rect -58 196 -57 200
rect -45 196 -40 200
rect -38 196 -35 200
rect -33 196 -32 200
rect -18 196 -17 200
rect -15 196 -14 200
rect 30 196 33 200
rect 35 196 38 200
rect 40 196 41 200
rect 135 196 138 200
rect 140 196 143 200
rect 145 196 146 200
rect 30 119 33 123
rect 35 119 38 123
rect 40 119 41 123
rect 87 123 88 127
rect 90 123 91 127
rect 111 119 114 123
rect 116 119 119 123
rect 121 119 122 123
rect 177 123 178 127
rect 180 123 181 127
rect 201 119 204 123
rect 206 119 209 123
rect 211 119 212 123
rect 60 115 61 119
rect 63 115 64 119
rect -168 110 -167 114
rect -165 110 -164 114
rect -152 110 -151 114
rect -149 110 -148 114
rect -136 110 -135 114
rect -133 110 -132 114
rect -117 110 -112 114
rect -110 110 -107 114
rect -105 110 -104 114
rect -83 110 -81 114
rect -79 110 -78 114
rect -61 110 -60 114
rect -58 110 -57 114
rect -45 110 -40 114
rect -38 110 -35 114
rect -33 110 -32 114
rect -18 110 -17 114
rect -15 110 -14 114
rect 141 115 142 119
rect 144 115 145 119
rect 231 115 232 119
rect 234 115 235 119
rect -168 64 -167 68
rect -165 64 -164 68
rect -152 64 -151 68
rect -149 64 -148 68
rect -136 64 -135 68
rect -133 64 -132 68
rect -117 64 -112 68
rect -110 64 -107 68
rect -105 64 -104 68
rect -83 64 -81 68
rect -79 64 -78 68
rect -61 64 -60 68
rect -58 64 -57 68
rect -45 64 -40 68
rect -38 64 -35 68
rect -33 64 -32 68
rect -18 64 -17 68
rect -15 64 -14 68
rect 30 61 33 65
rect 35 61 38 65
rect 40 61 41 65
rect 111 61 114 65
rect 116 61 119 65
rect 121 61 122 65
rect 201 61 204 65
rect 206 61 209 65
rect 211 61 212 65
rect 30 -13 33 -9
rect 35 -13 38 -9
rect 40 -13 41 -9
rect 60 -17 61 -13
rect 63 -17 64 -13
rect -168 -22 -167 -18
rect -165 -22 -164 -18
rect -152 -22 -151 -18
rect -149 -22 -148 -18
rect -136 -22 -135 -18
rect -133 -22 -132 -18
rect -117 -22 -112 -18
rect -110 -22 -107 -18
rect -105 -22 -104 -18
rect -83 -22 -81 -18
rect -79 -22 -78 -18
rect -61 -22 -60 -18
rect -58 -22 -57 -18
rect -45 -22 -40 -18
rect -38 -22 -35 -18
rect -33 -22 -32 -18
rect -18 -22 -17 -18
rect -15 -22 -14 -18
rect -168 -68 -167 -64
rect -165 -68 -164 -64
rect -152 -68 -151 -64
rect -149 -68 -148 -64
rect -136 -68 -135 -64
rect -133 -68 -132 -64
rect -117 -68 -112 -64
rect -110 -68 -107 -64
rect -105 -68 -104 -64
rect -83 -68 -81 -64
rect -79 -68 -78 -64
rect -61 -68 -60 -64
rect -58 -68 -57 -64
rect -45 -68 -40 -64
rect -38 -68 -35 -64
rect -33 -68 -32 -64
rect -18 -68 -17 -64
rect -15 -68 -14 -64
rect 66 -68 67 -64
rect 69 -68 70 -64
rect 74 -68 80 -64
rect 84 -68 85 -64
rect 87 -68 88 -64
rect 100 -68 101 -64
rect 103 -68 104 -64
rect 116 -68 117 -64
rect 119 -68 120 -64
rect 135 -68 140 -64
rect 142 -68 145 -64
rect 147 -68 148 -64
rect 169 -68 171 -64
rect 173 -68 174 -64
rect 191 -68 192 -64
rect 194 -68 195 -64
rect 207 -68 212 -64
rect 214 -68 217 -64
rect 219 -68 220 -64
rect 234 -68 235 -64
rect 237 -68 238 -64
rect 30 -75 33 -71
rect 35 -75 38 -71
rect 40 -75 41 -71
<< pdiffusion >>
rect 6 405 7 413
rect 9 405 10 413
rect -168 392 -167 400
rect -165 392 -164 400
rect -152 392 -151 400
rect -149 392 -148 400
rect -136 392 -135 400
rect -133 392 -132 400
rect -117 392 -112 400
rect -110 392 -107 400
rect -105 392 -104 400
rect -83 392 -81 400
rect -79 392 -78 400
rect -61 392 -60 400
rect -58 392 -57 400
rect -45 392 -40 400
rect -38 392 -35 400
rect -33 392 -32 400
rect -18 392 -17 400
rect -15 392 -14 400
rect 30 399 33 407
rect 35 399 38 407
rect 40 399 41 407
rect 60 405 61 413
rect 63 405 64 413
rect 87 405 88 413
rect 90 405 91 413
rect 111 399 114 407
rect 116 399 119 407
rect 121 399 122 407
rect 141 405 142 413
rect 144 405 145 413
rect -168 306 -167 314
rect -165 306 -164 314
rect -152 306 -151 314
rect -149 306 -148 314
rect -136 306 -135 314
rect -133 306 -132 314
rect -117 306 -112 314
rect -110 306 -107 314
rect -105 306 -104 314
rect -83 306 -81 314
rect -79 306 -78 314
rect -61 306 -60 314
rect -58 306 -57 314
rect -45 306 -40 314
rect -38 306 -35 314
rect -33 306 -32 314
rect -18 306 -17 314
rect -15 306 -14 314
rect 30 307 33 315
rect 35 307 38 315
rect 40 307 41 315
rect 111 307 114 315
rect 116 307 119 315
rect 121 307 122 315
rect -168 260 -167 268
rect -165 260 -164 268
rect -152 260 -151 268
rect -149 260 -148 268
rect -136 260 -135 268
rect -133 260 -132 268
rect -117 260 -112 268
rect -110 260 -107 268
rect -105 260 -104 268
rect -83 260 -81 268
rect -79 260 -78 268
rect -61 260 -60 268
rect -58 260 -57 268
rect -45 260 -40 268
rect -38 260 -35 268
rect -33 260 -32 268
rect -18 260 -17 268
rect -15 260 -14 268
rect 30 267 33 275
rect 35 267 38 275
rect 40 267 41 275
rect 60 273 61 281
rect 63 273 64 281
rect 111 273 112 281
rect 114 273 115 281
rect 135 267 138 275
rect 140 267 143 275
rect 145 267 146 275
rect 165 273 166 281
rect 168 273 169 281
rect -168 174 -167 182
rect -165 174 -164 182
rect -152 174 -151 182
rect -149 174 -148 182
rect -136 174 -135 182
rect -133 174 -132 182
rect -117 174 -112 182
rect -110 174 -107 182
rect -105 174 -104 182
rect -83 174 -81 182
rect -79 174 -78 182
rect -61 174 -60 182
rect -58 174 -57 182
rect -45 174 -40 182
rect -38 174 -35 182
rect -33 174 -32 182
rect -18 174 -17 182
rect -15 174 -14 182
rect 30 176 33 184
rect 35 176 38 184
rect 40 176 41 184
rect 135 176 138 184
rect 140 176 143 184
rect 145 176 146 184
rect -168 128 -167 136
rect -165 128 -164 136
rect -152 128 -151 136
rect -149 128 -148 136
rect -136 128 -135 136
rect -133 128 -132 136
rect -117 128 -112 136
rect -110 128 -107 136
rect -105 128 -104 136
rect -83 128 -81 136
rect -79 128 -78 136
rect -61 128 -60 136
rect -58 128 -57 136
rect -45 128 -40 136
rect -38 128 -35 136
rect -33 128 -32 136
rect -18 128 -17 136
rect -15 128 -14 136
rect 30 135 33 143
rect 35 135 38 143
rect 40 135 41 143
rect 60 141 61 149
rect 63 141 64 149
rect 87 141 88 149
rect 90 141 91 149
rect 111 135 114 143
rect 116 135 119 143
rect 121 135 122 143
rect 141 141 142 149
rect 144 141 145 149
rect 177 141 178 149
rect 180 141 181 149
rect 201 135 204 143
rect 206 135 209 143
rect 211 135 212 143
rect 231 141 232 149
rect 234 141 235 149
rect -168 42 -167 50
rect -165 42 -164 50
rect -152 42 -151 50
rect -149 42 -148 50
rect -136 42 -135 50
rect -133 42 -132 50
rect -117 42 -112 50
rect -110 42 -107 50
rect -105 42 -104 50
rect -83 42 -81 50
rect -79 42 -78 50
rect -61 42 -60 50
rect -58 42 -57 50
rect -45 42 -40 50
rect -38 42 -35 50
rect -33 42 -32 50
rect -18 42 -17 50
rect -15 42 -14 50
rect 30 41 33 49
rect 35 41 38 49
rect 40 41 41 49
rect 111 41 114 49
rect 116 41 119 49
rect 121 41 122 49
rect 201 41 204 49
rect 206 41 209 49
rect 211 41 212 49
rect -168 -4 -167 4
rect -165 -4 -164 4
rect -152 -4 -151 4
rect -149 -4 -148 4
rect -136 -4 -135 4
rect -133 -4 -132 4
rect -117 -4 -112 4
rect -110 -4 -107 4
rect -105 -4 -104 4
rect -83 -4 -81 4
rect -79 -4 -78 4
rect -61 -4 -60 4
rect -58 -4 -57 4
rect -45 -4 -40 4
rect -38 -4 -35 4
rect -33 -4 -32 4
rect -18 -4 -17 4
rect -15 -4 -14 4
rect 30 3 33 11
rect 35 3 38 11
rect 40 3 41 11
rect 60 9 61 17
rect 63 9 64 17
rect -168 -90 -167 -82
rect -165 -90 -164 -82
rect -152 -90 -151 -82
rect -149 -90 -148 -82
rect -136 -90 -135 -82
rect -133 -90 -132 -82
rect -117 -90 -112 -82
rect -110 -90 -107 -82
rect -105 -90 -104 -82
rect -83 -90 -81 -82
rect -79 -90 -78 -82
rect -61 -90 -60 -82
rect -58 -90 -57 -82
rect -45 -90 -40 -82
rect -38 -90 -35 -82
rect -33 -90 -32 -82
rect -18 -90 -17 -82
rect -15 -90 -14 -82
rect 30 -95 33 -87
rect 35 -95 38 -87
rect 40 -95 41 -87
rect 66 -90 67 -82
rect 69 -90 70 -82
rect 74 -90 80 -82
rect 84 -90 85 -82
rect 87 -90 88 -82
rect 100 -90 101 -82
rect 103 -90 104 -82
rect 116 -90 117 -82
rect 119 -90 120 -82
rect 135 -90 140 -82
rect 142 -90 145 -82
rect 147 -90 148 -82
rect 169 -90 171 -82
rect 173 -90 174 -82
rect 191 -90 192 -82
rect 194 -90 195 -82
rect 207 -90 212 -82
rect 214 -90 217 -82
rect 219 -90 220 -82
rect 234 -90 235 -82
rect 237 -90 238 -82
<< ndcontact >>
rect 2 387 6 391
rect 10 387 14 391
rect 26 383 30 387
rect 41 383 45 387
rect 83 387 87 391
rect 91 387 95 391
rect 107 383 111 387
rect 122 383 126 387
rect 56 379 60 383
rect 64 379 68 383
rect -172 374 -168 378
rect -164 374 -160 378
rect -156 374 -152 378
rect -148 374 -144 378
rect -140 374 -136 378
rect -132 374 -128 378
rect -121 374 -117 378
rect -104 374 -100 378
rect -87 374 -83 378
rect -78 374 -74 378
rect -65 374 -61 378
rect -57 374 -53 378
rect -49 374 -45 378
rect -32 374 -28 378
rect -22 374 -18 378
rect -14 374 -10 378
rect 137 379 141 383
rect 145 379 149 383
rect -172 328 -168 332
rect -164 328 -160 332
rect -156 328 -152 332
rect -148 328 -144 332
rect -140 328 -136 332
rect -132 328 -128 332
rect -121 328 -117 332
rect -104 328 -100 332
rect -87 328 -83 332
rect -78 328 -74 332
rect -65 328 -61 332
rect -57 328 -53 332
rect -49 328 -45 332
rect -32 328 -28 332
rect -22 328 -18 332
rect -14 328 -10 332
rect 26 327 30 331
rect 41 327 45 331
rect 107 327 111 331
rect 122 327 126 331
rect 26 251 30 255
rect 41 251 45 255
rect 107 255 111 259
rect 115 255 119 259
rect 131 251 135 255
rect 146 251 150 255
rect 56 247 60 251
rect 64 247 68 251
rect -172 242 -168 246
rect -164 242 -160 246
rect -156 242 -152 246
rect -148 242 -144 246
rect -140 242 -136 246
rect -132 242 -128 246
rect -121 242 -117 246
rect -104 242 -100 246
rect -87 242 -83 246
rect -78 242 -74 246
rect -65 242 -61 246
rect -57 242 -53 246
rect -49 242 -45 246
rect -32 242 -28 246
rect -22 242 -18 246
rect -14 242 -10 246
rect 161 247 165 251
rect 169 247 173 251
rect -172 196 -168 200
rect -164 196 -160 200
rect -156 196 -152 200
rect -148 196 -144 200
rect -140 196 -136 200
rect -132 196 -128 200
rect -121 196 -117 200
rect -104 196 -100 200
rect -87 196 -83 200
rect -78 196 -74 200
rect -65 196 -61 200
rect -57 196 -53 200
rect -49 196 -45 200
rect -32 196 -28 200
rect -22 196 -18 200
rect -14 196 -10 200
rect 26 196 30 200
rect 41 196 45 200
rect 131 196 135 200
rect 146 196 150 200
rect 26 119 30 123
rect 41 119 45 123
rect 83 123 87 127
rect 91 123 95 127
rect 107 119 111 123
rect 122 119 126 123
rect 173 123 177 127
rect 181 123 185 127
rect 197 119 201 123
rect 212 119 216 123
rect 56 115 60 119
rect 64 115 68 119
rect -172 110 -168 114
rect -164 110 -160 114
rect -156 110 -152 114
rect -148 110 -144 114
rect -140 110 -136 114
rect -132 110 -128 114
rect -121 110 -117 114
rect -104 110 -100 114
rect -87 110 -83 114
rect -78 110 -74 114
rect -65 110 -61 114
rect -57 110 -53 114
rect -49 110 -45 114
rect -32 110 -28 114
rect -22 110 -18 114
rect -14 110 -10 114
rect 137 115 141 119
rect 145 115 149 119
rect 227 115 231 119
rect 235 115 239 119
rect -172 64 -168 68
rect -164 64 -160 68
rect -156 64 -152 68
rect -148 64 -144 68
rect -140 64 -136 68
rect -132 64 -128 68
rect -121 64 -117 68
rect -104 64 -100 68
rect -87 64 -83 68
rect -78 64 -74 68
rect -65 64 -61 68
rect -57 64 -53 68
rect -49 64 -45 68
rect -32 64 -28 68
rect -22 64 -18 68
rect -14 64 -10 68
rect 26 61 30 65
rect 41 61 45 65
rect 107 61 111 65
rect 122 61 126 65
rect 197 61 201 65
rect 212 61 216 65
rect 26 -13 30 -9
rect 41 -13 45 -9
rect 56 -17 60 -13
rect 64 -17 68 -13
rect -172 -22 -168 -18
rect -164 -22 -160 -18
rect -156 -22 -152 -18
rect -148 -22 -144 -18
rect -140 -22 -136 -18
rect -132 -22 -128 -18
rect -121 -22 -117 -18
rect -104 -22 -100 -18
rect -87 -22 -83 -18
rect -78 -22 -74 -18
rect -65 -22 -61 -18
rect -57 -22 -53 -18
rect -49 -22 -45 -18
rect -32 -22 -28 -18
rect -22 -22 -18 -18
rect -14 -22 -10 -18
rect -172 -68 -168 -64
rect -164 -68 -160 -64
rect -156 -68 -152 -64
rect -148 -68 -144 -64
rect -140 -68 -136 -64
rect -132 -68 -128 -64
rect -121 -68 -117 -64
rect -104 -68 -100 -64
rect -87 -68 -83 -64
rect -78 -68 -74 -64
rect -65 -68 -61 -64
rect -57 -68 -53 -64
rect -49 -68 -45 -64
rect -32 -68 -28 -64
rect -22 -68 -18 -64
rect -14 -68 -10 -64
rect 62 -68 66 -64
rect 70 -68 74 -64
rect 80 -68 84 -64
rect 88 -68 92 -64
rect 96 -68 100 -64
rect 104 -68 108 -64
rect 112 -68 116 -64
rect 120 -68 124 -64
rect 131 -68 135 -64
rect 148 -68 152 -64
rect 165 -68 169 -64
rect 174 -68 178 -64
rect 187 -68 191 -64
rect 195 -68 199 -64
rect 203 -68 207 -64
rect 220 -68 224 -64
rect 230 -68 234 -64
rect 238 -68 242 -64
rect 26 -75 30 -71
rect 41 -75 45 -71
<< pdcontact >>
rect 2 405 6 413
rect 10 405 14 413
rect -172 392 -168 400
rect -164 392 -160 400
rect -156 392 -152 400
rect -148 392 -144 400
rect -140 392 -136 400
rect -132 392 -128 400
rect -121 392 -117 400
rect -104 392 -100 400
rect -87 392 -83 400
rect -78 392 -74 400
rect -65 392 -61 400
rect -57 392 -53 400
rect -49 392 -45 400
rect -32 392 -28 400
rect -22 392 -18 400
rect -14 392 -10 400
rect 26 399 30 407
rect 41 399 45 407
rect 56 405 60 413
rect 64 405 68 413
rect 83 405 87 413
rect 91 405 95 413
rect 107 399 111 407
rect 122 399 126 407
rect 137 405 141 413
rect 145 405 149 413
rect -172 306 -168 314
rect -164 306 -160 314
rect -156 306 -152 314
rect -148 306 -144 314
rect -140 306 -136 314
rect -132 306 -128 314
rect -121 306 -117 314
rect -104 306 -100 314
rect -87 306 -83 314
rect -78 306 -74 314
rect -65 306 -61 314
rect -57 306 -53 314
rect -49 306 -45 314
rect -32 306 -28 314
rect -22 306 -18 314
rect -14 306 -10 314
rect 26 307 30 315
rect 41 307 45 315
rect 107 307 111 315
rect 122 307 126 315
rect -172 260 -168 268
rect -164 260 -160 268
rect -156 260 -152 268
rect -148 260 -144 268
rect -140 260 -136 268
rect -132 260 -128 268
rect -121 260 -117 268
rect -104 260 -100 268
rect -87 260 -83 268
rect -78 260 -74 268
rect -65 260 -61 268
rect -57 260 -53 268
rect -49 260 -45 268
rect -32 260 -28 268
rect -22 260 -18 268
rect -14 260 -10 268
rect 26 267 30 275
rect 41 267 45 275
rect 56 273 60 281
rect 64 273 68 281
rect 107 273 111 281
rect 115 273 119 281
rect 131 267 135 275
rect 146 267 150 275
rect 161 273 165 281
rect 169 273 173 281
rect -172 174 -168 182
rect -164 174 -160 182
rect -156 174 -152 182
rect -148 174 -144 182
rect -140 174 -136 182
rect -132 174 -128 182
rect -121 174 -117 182
rect -104 174 -100 182
rect -87 174 -83 182
rect -78 174 -74 182
rect -65 174 -61 182
rect -57 174 -53 182
rect -49 174 -45 182
rect -32 174 -28 182
rect -22 174 -18 182
rect -14 174 -10 182
rect 26 176 30 184
rect 41 176 45 184
rect 131 176 135 184
rect 146 176 150 184
rect -172 128 -168 136
rect -164 128 -160 136
rect -156 128 -152 136
rect -148 128 -144 136
rect -140 128 -136 136
rect -132 128 -128 136
rect -121 128 -117 136
rect -104 128 -100 136
rect -87 128 -83 136
rect -78 128 -74 136
rect -65 128 -61 136
rect -57 128 -53 136
rect -49 128 -45 136
rect -32 128 -28 136
rect -22 128 -18 136
rect -14 128 -10 136
rect 26 135 30 143
rect 41 135 45 143
rect 56 141 60 149
rect 64 141 68 149
rect 83 141 87 149
rect 91 141 95 149
rect 107 135 111 143
rect 122 135 126 143
rect 137 141 141 149
rect 145 141 149 149
rect 173 141 177 149
rect 181 141 185 149
rect 197 135 201 143
rect 212 135 216 143
rect 227 141 231 149
rect 235 141 239 149
rect -172 42 -168 50
rect -164 42 -160 50
rect -156 42 -152 50
rect -148 42 -144 50
rect -140 42 -136 50
rect -132 42 -128 50
rect -121 42 -117 50
rect -104 42 -100 50
rect -87 42 -83 50
rect -78 42 -74 50
rect -65 42 -61 50
rect -57 42 -53 50
rect -49 42 -45 50
rect -32 42 -28 50
rect -22 42 -18 50
rect -14 42 -10 50
rect 26 41 30 49
rect 41 41 45 49
rect 107 41 111 49
rect 122 41 126 49
rect 197 41 201 49
rect 212 41 216 49
rect -172 -4 -168 4
rect -164 -4 -160 4
rect -156 -4 -152 4
rect -148 -4 -144 4
rect -140 -4 -136 4
rect -132 -4 -128 4
rect -121 -4 -117 4
rect -104 -4 -100 4
rect -87 -4 -83 4
rect -78 -4 -74 4
rect -65 -4 -61 4
rect -57 -4 -53 4
rect -49 -4 -45 4
rect -32 -4 -28 4
rect -22 -4 -18 4
rect -14 -4 -10 4
rect 26 3 30 11
rect 41 3 45 11
rect 56 9 60 17
rect 64 9 68 17
rect -172 -90 -168 -82
rect -164 -90 -160 -82
rect -156 -90 -152 -82
rect -148 -90 -144 -82
rect -140 -90 -136 -82
rect -132 -90 -128 -82
rect -121 -90 -117 -82
rect -104 -90 -100 -82
rect -87 -90 -83 -82
rect -78 -90 -74 -82
rect -65 -90 -61 -82
rect -57 -90 -53 -82
rect -49 -90 -45 -82
rect -32 -90 -28 -82
rect -22 -90 -18 -82
rect -14 -90 -10 -82
rect 26 -95 30 -87
rect 41 -95 45 -87
rect 62 -90 66 -82
rect 70 -90 74 -82
rect 80 -90 84 -82
rect 88 -90 92 -82
rect 96 -90 100 -82
rect 104 -90 108 -82
rect 112 -90 116 -82
rect 120 -90 124 -82
rect 131 -90 135 -82
rect 148 -90 152 -82
rect 165 -90 169 -82
rect 174 -90 178 -82
rect 187 -90 191 -82
rect 195 -90 199 -82
rect 203 -90 207 -82
rect 220 -90 224 -82
rect 230 -90 234 -82
rect 238 -90 242 -82
<< psubstratepcontact >>
rect -166 351 -162 355
rect -131 351 -127 355
rect -5 351 -1 355
rect 19 351 23 355
rect 73 351 80 355
rect 100 351 104 355
rect 154 351 158 355
rect -166 219 -162 223
rect -131 219 -127 223
rect -5 219 -1 223
rect 19 219 23 223
rect 73 219 77 223
rect 100 219 104 223
rect 124 219 128 223
rect -166 87 -162 91
rect -131 87 -127 91
rect -5 87 -1 91
rect 19 87 23 91
rect 73 87 80 91
rect 100 87 104 91
rect 154 87 158 91
rect 190 87 194 91
rect 244 87 248 91
rect -166 -45 -162 -41
rect -131 -45 -127 -41
rect -5 -45 -1 -41
rect 19 -45 23 -41
rect 92 -52 96 -48
rect 121 -52 125 -48
rect 157 -52 161 -48
rect 196 -52 200 -48
rect 73 -111 77 -107
<< nsubstratencontact >>
rect -157 417 -153 421
rect -128 417 -124 421
rect -103 417 -99 421
rect -61 417 -57 421
rect -5 417 -1 421
rect 19 417 23 421
rect 73 417 77 421
rect 100 417 104 421
rect 154 417 158 421
rect -157 285 -153 289
rect -128 285 -124 289
rect -103 285 -99 289
rect -61 285 -57 289
rect -5 285 -1 289
rect 19 285 23 289
rect 73 285 77 289
rect 100 285 104 289
rect 162 285 166 289
rect -157 153 -153 157
rect -128 153 -124 157
rect -103 153 -99 157
rect -61 153 -57 157
rect -5 153 -1 157
rect 19 153 23 157
rect 73 153 77 157
rect 100 153 104 157
rect 154 153 158 157
rect 162 153 166 157
rect 190 153 194 157
rect 244 153 248 157
rect -157 21 -153 25
rect -128 21 -124 25
rect -103 21 -99 25
rect -61 21 -57 25
rect -5 21 -1 25
rect 19 21 23 25
rect 73 21 77 25
rect 100 21 104 25
rect 190 21 194 25
rect 89 -104 93 -100
rect 121 -104 125 -100
rect 157 -104 161 -100
rect 196 -104 200 -100
rect -157 -111 -153 -107
rect -128 -111 -124 -107
rect -103 -111 -99 -107
rect -61 -111 -57 -107
rect 19 -111 23 -107
<< polysilicon >>
rect 7 413 9 415
rect -151 407 -149 410
rect -107 407 -105 410
rect -81 407 -79 410
rect -35 407 -33 410
rect -81 403 -80 407
rect 33 407 35 411
rect 61 413 63 415
rect 88 413 90 415
rect 38 407 40 410
rect -167 400 -165 402
rect -151 400 -149 403
rect -135 400 -133 402
rect -112 400 -110 402
rect -107 400 -105 403
rect -81 400 -79 403
rect -60 400 -58 403
rect -40 400 -38 402
rect -35 400 -33 403
rect -17 400 -15 402
rect -167 378 -165 392
rect -151 390 -149 392
rect -151 378 -149 380
rect -135 378 -133 392
rect -112 387 -110 392
rect -107 390 -105 392
rect -81 390 -79 392
rect -116 383 -110 387
rect -112 378 -110 383
rect -107 378 -105 380
rect -81 378 -79 380
rect -60 378 -58 392
rect -40 387 -38 392
rect -35 390 -33 392
rect -44 383 -38 387
rect -40 378 -38 383
rect -35 378 -33 380
rect -17 378 -15 392
rect 7 391 9 405
rect 114 407 116 411
rect 142 413 144 415
rect 119 407 121 410
rect 33 396 35 399
rect 38 397 40 399
rect 34 392 35 396
rect 33 387 35 392
rect 38 387 40 389
rect 7 385 9 387
rect 61 383 63 405
rect 88 391 90 405
rect 114 396 116 399
rect 119 397 121 399
rect 115 392 116 396
rect 114 387 116 392
rect 119 387 121 389
rect 88 385 90 387
rect 142 383 144 405
rect 33 381 35 383
rect 38 378 40 383
rect 114 381 116 383
rect 61 377 63 379
rect 119 378 121 383
rect 142 377 144 379
rect -167 372 -165 374
rect -151 370 -149 374
rect -135 372 -133 374
rect -112 372 -110 374
rect -150 366 -149 370
rect -107 369 -105 374
rect -81 370 -79 374
rect -60 372 -58 374
rect -40 372 -38 374
rect -151 363 -149 366
rect -106 365 -105 369
rect -80 366 -79 370
rect -35 369 -33 374
rect -17 372 -15 374
rect -107 363 -105 365
rect -81 362 -79 366
rect -34 365 -33 369
rect -35 363 -33 365
rect -151 340 -149 343
rect -107 341 -105 343
rect -150 336 -149 340
rect -106 337 -105 341
rect -81 340 -79 344
rect -35 341 -33 343
rect -167 332 -165 334
rect -151 332 -149 336
rect -135 332 -133 334
rect -112 332 -110 334
rect -107 332 -105 337
rect -80 336 -79 340
rect -34 337 -33 341
rect -81 332 -79 336
rect -60 332 -58 334
rect -40 332 -38 334
rect -35 332 -33 337
rect -17 332 -15 334
rect 33 331 35 334
rect 38 331 40 334
rect 114 331 116 334
rect 119 331 121 334
rect -167 314 -165 328
rect -151 326 -149 328
rect -151 314 -149 316
rect -135 314 -133 328
rect -112 323 -110 328
rect -107 326 -105 328
rect -81 326 -79 328
rect -116 319 -110 323
rect -112 314 -110 319
rect -107 314 -105 316
rect -81 314 -79 316
rect -60 314 -58 328
rect -40 323 -38 328
rect -35 326 -33 328
rect -44 319 -38 323
rect -40 314 -38 319
rect -35 314 -33 316
rect -17 314 -15 328
rect 33 315 35 327
rect 38 325 40 327
rect 38 315 40 317
rect 114 315 116 327
rect 119 325 121 327
rect 119 315 121 317
rect -167 304 -165 306
rect -151 303 -149 306
rect -135 304 -133 306
rect -112 304 -110 306
rect -107 303 -105 306
rect -81 303 -79 306
rect -60 303 -58 306
rect -40 304 -38 306
rect -35 303 -33 306
rect -17 304 -15 306
rect 33 305 35 307
rect -81 299 -80 303
rect 38 302 40 307
rect 114 305 116 307
rect 119 302 121 307
rect -151 296 -149 299
rect -107 296 -105 299
rect -81 296 -79 299
rect -35 296 -33 299
rect -151 275 -149 278
rect -107 275 -105 278
rect -81 275 -79 278
rect -35 275 -33 278
rect 33 275 35 279
rect 61 281 63 283
rect 112 281 114 283
rect 38 275 40 278
rect -81 271 -80 275
rect -167 268 -165 270
rect -151 268 -149 271
rect -135 268 -133 270
rect -112 268 -110 270
rect -107 268 -105 271
rect -81 268 -79 271
rect -60 268 -58 271
rect -40 268 -38 270
rect -35 268 -33 271
rect -17 268 -15 270
rect 138 275 140 279
rect 166 281 168 283
rect 143 275 145 278
rect 33 264 35 267
rect 38 265 40 267
rect 34 260 35 264
rect -167 246 -165 260
rect -151 258 -149 260
rect -151 246 -149 248
rect -135 246 -133 260
rect -112 255 -110 260
rect -107 258 -105 260
rect -81 258 -79 260
rect -116 251 -110 255
rect -112 246 -110 251
rect -107 246 -105 248
rect -81 246 -79 248
rect -60 246 -58 260
rect -40 255 -38 260
rect -35 258 -33 260
rect -44 251 -38 255
rect -40 246 -38 251
rect -35 246 -33 248
rect -17 246 -15 260
rect 33 255 35 260
rect 38 255 40 257
rect 61 251 63 273
rect 112 259 114 273
rect 138 264 140 267
rect 143 265 145 267
rect 139 260 140 264
rect 138 255 140 260
rect 143 255 145 257
rect 112 253 114 255
rect 166 251 168 273
rect 33 249 35 251
rect 38 246 40 251
rect 138 249 140 251
rect 61 245 63 247
rect 143 246 145 251
rect 166 245 168 247
rect -167 240 -165 242
rect -151 238 -149 242
rect -135 240 -133 242
rect -112 240 -110 242
rect -150 234 -149 238
rect -107 237 -105 242
rect -81 238 -79 242
rect -60 240 -58 242
rect -40 240 -38 242
rect -151 231 -149 234
rect -106 233 -105 237
rect -80 234 -79 238
rect -35 237 -33 242
rect -17 240 -15 242
rect -107 231 -105 233
rect -81 230 -79 234
rect -34 233 -33 237
rect -35 231 -33 233
rect -151 208 -149 211
rect -107 209 -105 211
rect -150 204 -149 208
rect -106 205 -105 209
rect -81 208 -79 212
rect -35 209 -33 211
rect -167 200 -165 202
rect -151 200 -149 204
rect -135 200 -133 202
rect -112 200 -110 202
rect -107 200 -105 205
rect -80 204 -79 208
rect -34 205 -33 209
rect -81 200 -79 204
rect -60 200 -58 202
rect -40 200 -38 202
rect -35 200 -33 205
rect -17 200 -15 202
rect 33 200 35 203
rect 38 200 40 203
rect 138 200 140 203
rect 143 200 145 203
rect -167 182 -165 196
rect -151 194 -149 196
rect -151 182 -149 184
rect -135 182 -133 196
rect -112 191 -110 196
rect -107 194 -105 196
rect -81 194 -79 196
rect -116 187 -110 191
rect -112 182 -110 187
rect -107 182 -105 184
rect -81 182 -79 184
rect -60 182 -58 196
rect -40 191 -38 196
rect -35 194 -33 196
rect -44 187 -38 191
rect -40 182 -38 187
rect -35 182 -33 184
rect -17 182 -15 196
rect 33 184 35 196
rect 38 194 40 196
rect 38 184 40 186
rect 138 184 140 196
rect 143 194 145 196
rect 143 184 145 186
rect 33 174 35 176
rect -167 172 -165 174
rect -151 171 -149 174
rect -135 172 -133 174
rect -112 172 -110 174
rect -107 171 -105 174
rect -81 171 -79 174
rect -60 171 -58 174
rect -40 172 -38 174
rect -35 171 -33 174
rect -17 172 -15 174
rect 38 171 40 176
rect 138 174 140 176
rect 143 171 145 176
rect -81 167 -80 171
rect -151 164 -149 167
rect -107 164 -105 167
rect -81 164 -79 167
rect -35 164 -33 167
rect -151 143 -149 146
rect -107 143 -105 146
rect -81 143 -79 146
rect -35 143 -33 146
rect 33 143 35 147
rect 61 149 63 151
rect 88 149 90 151
rect 38 143 40 146
rect -81 139 -80 143
rect -167 136 -165 138
rect -151 136 -149 139
rect -135 136 -133 138
rect -112 136 -110 138
rect -107 136 -105 139
rect -81 136 -79 139
rect -60 136 -58 139
rect -40 136 -38 138
rect -35 136 -33 139
rect -17 136 -15 138
rect 114 143 116 147
rect 142 149 144 151
rect 178 149 180 151
rect 119 143 121 146
rect 33 132 35 135
rect 38 133 40 135
rect 34 128 35 132
rect -167 114 -165 128
rect -151 126 -149 128
rect -151 114 -149 116
rect -135 114 -133 128
rect -112 123 -110 128
rect -107 126 -105 128
rect -81 126 -79 128
rect -116 119 -110 123
rect -112 114 -110 119
rect -107 114 -105 116
rect -81 114 -79 116
rect -60 114 -58 128
rect -40 123 -38 128
rect -35 126 -33 128
rect -44 119 -38 123
rect -40 114 -38 119
rect -35 114 -33 116
rect -17 114 -15 128
rect 33 123 35 128
rect 38 123 40 125
rect 61 119 63 141
rect 88 127 90 141
rect 204 143 206 147
rect 232 149 234 151
rect 209 143 211 146
rect 114 132 116 135
rect 119 133 121 135
rect 115 128 116 132
rect 114 123 116 128
rect 119 123 121 125
rect 88 121 90 123
rect 142 119 144 141
rect 178 127 180 141
rect 204 132 206 135
rect 209 133 211 135
rect 205 128 206 132
rect 204 123 206 128
rect 209 123 211 125
rect 178 121 180 123
rect 232 119 234 141
rect 33 117 35 119
rect 38 114 40 119
rect 114 117 116 119
rect 61 113 63 115
rect 119 114 121 119
rect 204 117 206 119
rect 142 113 144 115
rect 209 114 211 119
rect 232 113 234 115
rect -167 108 -165 110
rect -151 106 -149 110
rect -135 108 -133 110
rect -112 108 -110 110
rect -150 102 -149 106
rect -107 105 -105 110
rect -81 106 -79 110
rect -60 108 -58 110
rect -40 108 -38 110
rect -151 99 -149 102
rect -106 101 -105 105
rect -80 102 -79 106
rect -35 105 -33 110
rect -17 108 -15 110
rect -107 99 -105 101
rect -81 98 -79 102
rect -34 101 -33 105
rect -35 99 -33 101
rect -151 76 -149 79
rect -107 77 -105 79
rect -150 72 -149 76
rect -106 73 -105 77
rect -81 76 -79 80
rect -35 77 -33 79
rect -167 68 -165 70
rect -151 68 -149 72
rect -135 68 -133 70
rect -112 68 -110 70
rect -107 68 -105 73
rect -80 72 -79 76
rect -34 73 -33 77
rect -81 68 -79 72
rect -60 68 -58 70
rect -40 68 -38 70
rect -35 68 -33 73
rect -17 68 -15 70
rect 33 65 35 68
rect 38 65 40 68
rect 114 65 116 68
rect 119 65 121 68
rect 204 65 206 68
rect 209 65 211 68
rect -167 50 -165 64
rect -151 62 -149 64
rect -151 50 -149 52
rect -135 50 -133 64
rect -112 59 -110 64
rect -107 62 -105 64
rect -81 62 -79 64
rect -116 55 -110 59
rect -112 50 -110 55
rect -107 50 -105 52
rect -81 50 -79 52
rect -60 50 -58 64
rect -40 59 -38 64
rect -35 62 -33 64
rect -44 55 -38 59
rect -40 50 -38 55
rect -35 50 -33 52
rect -17 50 -15 64
rect 33 49 35 61
rect 38 59 40 61
rect 38 49 40 51
rect 114 49 116 61
rect 119 59 121 61
rect 119 49 121 51
rect 204 49 206 61
rect 209 59 211 61
rect 209 49 211 51
rect -167 40 -165 42
rect -151 39 -149 42
rect -135 40 -133 42
rect -112 40 -110 42
rect -107 39 -105 42
rect -81 39 -79 42
rect -60 39 -58 42
rect -40 40 -38 42
rect -35 39 -33 42
rect -17 40 -15 42
rect 33 39 35 41
rect -81 35 -80 39
rect 38 36 40 41
rect 114 39 116 41
rect 119 36 121 41
rect 204 39 206 41
rect 209 36 211 41
rect -151 32 -149 35
rect -107 32 -105 35
rect -81 32 -79 35
rect -35 32 -33 35
rect -151 11 -149 14
rect -107 11 -105 14
rect -81 11 -79 14
rect -35 11 -33 14
rect 33 11 35 15
rect 61 17 63 19
rect 38 11 40 14
rect -81 7 -80 11
rect -167 4 -165 6
rect -151 4 -149 7
rect -135 4 -133 6
rect -112 4 -110 6
rect -107 4 -105 7
rect -81 4 -79 7
rect -60 4 -58 7
rect -40 4 -38 6
rect -35 4 -33 7
rect -17 4 -15 6
rect 33 0 35 3
rect 38 1 40 3
rect 34 -4 35 0
rect -167 -18 -165 -4
rect -151 -6 -149 -4
rect -151 -18 -149 -16
rect -135 -18 -133 -4
rect -112 -9 -110 -4
rect -107 -6 -105 -4
rect -81 -6 -79 -4
rect -116 -13 -110 -9
rect -112 -18 -110 -13
rect -107 -18 -105 -16
rect -81 -18 -79 -16
rect -60 -18 -58 -4
rect -40 -9 -38 -4
rect -35 -6 -33 -4
rect -44 -13 -38 -9
rect -40 -18 -38 -13
rect -35 -18 -33 -16
rect -17 -18 -15 -4
rect 33 -9 35 -4
rect 38 -9 40 -7
rect 61 -13 63 9
rect 33 -15 35 -13
rect 38 -18 40 -13
rect 61 -19 63 -17
rect -167 -24 -165 -22
rect -151 -26 -149 -22
rect -135 -24 -133 -22
rect -112 -24 -110 -22
rect -150 -30 -149 -26
rect -107 -27 -105 -22
rect -81 -26 -79 -22
rect -60 -24 -58 -22
rect -40 -24 -38 -22
rect -151 -33 -149 -30
rect -106 -31 -105 -27
rect -80 -30 -79 -26
rect -35 -27 -33 -22
rect -17 -24 -15 -22
rect -107 -33 -105 -31
rect -81 -34 -79 -30
rect -34 -31 -33 -27
rect -35 -33 -33 -31
rect -151 -56 -149 -53
rect -107 -55 -105 -53
rect -150 -60 -149 -56
rect -106 -59 -105 -55
rect -81 -56 -79 -52
rect -35 -55 -33 -53
rect -167 -64 -165 -62
rect -151 -64 -149 -60
rect -135 -64 -133 -62
rect -112 -64 -110 -62
rect -107 -64 -105 -59
rect -80 -60 -79 -56
rect -34 -59 -33 -55
rect 101 -56 103 -53
rect 145 -55 147 -53
rect -81 -64 -79 -60
rect -60 -64 -58 -62
rect -40 -64 -38 -62
rect -35 -64 -33 -59
rect 102 -60 103 -56
rect 146 -59 147 -55
rect 171 -56 173 -52
rect 217 -55 219 -53
rect -17 -64 -15 -62
rect 67 -64 69 -61
rect 85 -64 87 -61
rect 101 -64 103 -60
rect 117 -64 119 -62
rect 140 -64 142 -62
rect 145 -64 147 -59
rect 172 -60 173 -56
rect 218 -59 219 -55
rect 171 -64 173 -60
rect 192 -64 194 -62
rect 212 -64 214 -62
rect 217 -64 219 -59
rect 235 -64 237 -62
rect -167 -82 -165 -68
rect -151 -70 -149 -68
rect -151 -82 -149 -80
rect -135 -82 -133 -68
rect -112 -73 -110 -68
rect -107 -70 -105 -68
rect -81 -70 -79 -68
rect -116 -77 -110 -73
rect -112 -82 -110 -77
rect -107 -82 -105 -80
rect -81 -82 -79 -80
rect -60 -82 -58 -68
rect -40 -73 -38 -68
rect -35 -70 -33 -68
rect -44 -77 -38 -73
rect -40 -82 -38 -77
rect -35 -82 -33 -80
rect -17 -82 -15 -68
rect 33 -71 35 -68
rect 38 -71 40 -68
rect 67 -73 69 -68
rect 33 -87 35 -75
rect 38 -77 40 -75
rect 67 -82 69 -77
rect 85 -82 87 -68
rect 101 -70 103 -68
rect 101 -82 103 -80
rect 117 -82 119 -68
rect 140 -73 142 -68
rect 145 -70 147 -68
rect 171 -70 173 -68
rect 136 -77 142 -73
rect 140 -82 142 -77
rect 145 -82 147 -80
rect 171 -82 173 -80
rect 192 -82 194 -68
rect 212 -73 214 -68
rect 217 -70 219 -68
rect 208 -77 214 -73
rect 212 -82 214 -77
rect 217 -82 219 -80
rect 235 -82 237 -68
rect 38 -87 40 -85
rect -167 -92 -165 -90
rect -151 -93 -149 -90
rect -135 -92 -133 -90
rect -112 -92 -110 -90
rect -107 -93 -105 -90
rect -81 -93 -79 -90
rect -60 -93 -58 -90
rect -40 -92 -38 -90
rect -35 -93 -33 -90
rect -17 -92 -15 -90
rect -81 -97 -80 -93
rect 67 -93 69 -90
rect 85 -93 87 -90
rect 101 -93 103 -90
rect 117 -92 119 -90
rect 140 -92 142 -90
rect 145 -93 147 -90
rect 171 -93 173 -90
rect 192 -93 194 -90
rect 212 -92 214 -90
rect 217 -93 219 -90
rect 235 -92 237 -90
rect 33 -97 35 -95
rect -151 -100 -149 -97
rect -107 -100 -105 -97
rect -81 -100 -79 -97
rect -35 -100 -33 -97
rect 38 -100 40 -95
rect 171 -97 172 -93
rect 101 -100 103 -97
rect 145 -100 147 -97
rect 171 -100 173 -97
rect 217 -100 219 -97
<< polycontact >>
rect -151 403 -147 407
rect -107 403 -103 407
rect -80 403 -76 407
rect -35 403 -31 407
rect 38 410 42 414
rect 3 396 7 400
rect -171 383 -167 387
rect -139 384 -135 388
rect -120 383 -116 387
rect -64 384 -60 388
rect -48 383 -44 387
rect -21 383 -17 387
rect 119 410 123 414
rect 30 392 34 396
rect 57 388 61 392
rect 84 396 88 400
rect 111 392 115 396
rect 138 388 142 392
rect 36 374 40 378
rect 117 374 121 378
rect -154 366 -150 370
rect -110 365 -106 369
rect -85 366 -80 370
rect -38 365 -34 369
rect -154 336 -150 340
rect -110 337 -106 341
rect -85 336 -80 340
rect -38 337 -34 341
rect 38 334 42 338
rect 119 334 123 338
rect -171 319 -167 323
rect -139 318 -135 322
rect -120 319 -116 323
rect -64 318 -60 322
rect -48 319 -44 323
rect -21 319 -17 323
rect 27 318 33 322
rect 108 318 114 322
rect -151 299 -147 303
rect -107 299 -103 303
rect -80 299 -76 303
rect -35 299 -31 303
rect 36 298 40 302
rect 117 298 121 302
rect 38 278 42 282
rect -151 271 -147 275
rect -107 271 -103 275
rect -80 271 -76 275
rect -35 271 -31 275
rect 143 278 147 282
rect 30 260 34 264
rect -171 251 -167 255
rect -139 252 -135 256
rect -120 251 -116 255
rect -64 252 -60 256
rect -48 251 -44 255
rect -21 251 -17 255
rect 57 256 61 260
rect 108 264 112 268
rect 135 260 139 264
rect 162 256 166 260
rect 36 242 40 246
rect 141 242 145 246
rect -154 234 -150 238
rect -110 233 -106 237
rect -85 234 -80 238
rect -38 233 -34 237
rect -154 204 -150 208
rect -110 205 -106 209
rect -85 204 -80 208
rect -38 205 -34 209
rect 38 203 42 207
rect 143 203 147 207
rect -171 187 -167 191
rect -139 186 -135 190
rect -120 187 -116 191
rect -64 186 -60 190
rect -48 187 -44 191
rect -21 187 -17 191
rect 27 187 33 191
rect 132 187 138 191
rect -151 167 -147 171
rect -107 167 -103 171
rect -80 167 -76 171
rect -35 167 -31 171
rect 36 167 40 171
rect 141 167 145 171
rect 38 146 42 150
rect -151 139 -147 143
rect -107 139 -103 143
rect -80 139 -76 143
rect -35 139 -31 143
rect 119 146 123 150
rect 30 128 34 132
rect -171 119 -167 123
rect -139 120 -135 124
rect -120 119 -116 123
rect -64 120 -60 124
rect -48 119 -44 123
rect -21 119 -17 123
rect 57 124 61 128
rect 84 132 88 136
rect 209 146 213 150
rect 111 128 115 132
rect 138 124 142 128
rect 174 132 178 136
rect 201 128 205 132
rect 228 124 232 128
rect 36 110 40 114
rect 117 110 121 114
rect 207 110 211 114
rect -154 102 -150 106
rect -110 101 -106 105
rect -85 102 -80 106
rect -38 101 -34 105
rect -154 72 -150 76
rect -110 73 -106 77
rect -85 72 -80 76
rect -38 73 -34 77
rect 38 68 42 72
rect 119 68 123 72
rect 209 68 213 72
rect -171 55 -167 59
rect -139 54 -135 58
rect -120 55 -116 59
rect -64 54 -60 58
rect -48 55 -44 59
rect -21 55 -17 59
rect 27 52 33 56
rect 108 52 114 56
rect 198 52 204 56
rect -151 35 -147 39
rect -107 35 -103 39
rect -80 35 -76 39
rect -35 35 -31 39
rect 36 32 40 36
rect 117 32 121 36
rect 207 32 211 36
rect 38 14 42 18
rect -151 7 -147 11
rect -107 7 -103 11
rect -80 7 -76 11
rect -35 7 -31 11
rect 30 -4 34 0
rect -171 -13 -167 -9
rect -139 -12 -135 -8
rect -120 -13 -116 -9
rect -64 -12 -60 -8
rect -48 -13 -44 -9
rect -21 -13 -17 -9
rect 57 -8 61 -4
rect 36 -22 40 -18
rect -154 -30 -150 -26
rect -110 -31 -106 -27
rect -85 -30 -80 -26
rect -38 -31 -34 -27
rect -154 -60 -150 -56
rect -110 -59 -106 -55
rect -85 -60 -80 -56
rect -38 -59 -34 -55
rect 98 -60 102 -56
rect 142 -59 146 -55
rect 167 -60 172 -56
rect 214 -59 218 -55
rect 38 -68 42 -64
rect -171 -77 -167 -73
rect -139 -78 -135 -74
rect -120 -77 -116 -73
rect -64 -78 -60 -74
rect -48 -77 -44 -73
rect -21 -77 -17 -73
rect 27 -84 33 -80
rect 65 -77 69 -73
rect 113 -78 117 -74
rect 132 -77 136 -73
rect 188 -78 192 -74
rect 204 -77 208 -73
rect 231 -77 235 -73
rect -151 -97 -147 -93
rect -107 -97 -103 -93
rect -80 -97 -76 -93
rect -35 -97 -31 -93
rect 101 -97 105 -93
rect 145 -97 149 -93
rect 172 -97 176 -93
rect 217 -97 221 -93
rect 36 -104 40 -100
<< metal1 >>
rect -179 417 -173 421
rect -169 417 -157 421
rect -153 417 -139 421
rect -135 417 -128 421
rect -124 417 -122 421
rect -118 417 -103 421
rect -99 417 -66 421
rect -62 417 -61 421
rect -57 417 -49 421
rect -45 417 -21 421
rect -17 417 -5 421
rect -1 417 19 421
rect 23 417 73 421
rect 77 417 100 421
rect 104 417 154 421
rect 158 417 177 421
rect -179 410 -146 414
rect -142 410 -115 414
rect -111 410 -93 414
rect -89 410 -28 414
rect -24 410 -10 414
rect 2 413 5 417
rect -103 403 -100 407
rect -76 403 -75 407
rect -31 403 -29 407
rect 11 400 14 405
rect 26 407 29 417
rect 56 413 59 417
rect 83 413 86 417
rect -176 383 -171 386
rect -163 386 -160 392
rect -156 386 -153 392
rect -163 383 -153 386
rect -163 378 -160 383
rect -156 378 -153 383
rect -147 388 -144 392
rect -147 384 -145 388
rect -141 384 -139 388
rect -131 387 -128 392
rect -103 389 -100 392
rect -131 385 -120 387
rect -147 378 -144 384
rect -131 383 -125 385
rect -131 378 -128 383
rect -121 383 -120 385
rect -102 385 -100 389
rect -103 378 -100 385
rect 0 396 3 399
rect 42 396 45 399
rect -87 388 -84 392
rect -77 388 -74 392
rect -77 384 -68 388
rect -56 387 -53 392
rect -31 388 -28 392
rect -87 378 -84 384
rect -77 378 -74 384
rect -56 383 -55 387
rect -51 383 -48 386
rect -29 384 -28 388
rect -13 387 -10 392
rect 11 391 14 396
rect 19 392 30 395
rect 42 393 50 396
rect -56 378 -53 383
rect -31 378 -28 384
rect -13 378 -10 383
rect -111 365 -110 369
rect -86 366 -85 370
rect -39 365 -38 369
rect -179 358 -158 362
rect -154 358 -99 362
rect -95 358 -74 362
rect -70 358 -43 362
rect -39 358 -10 362
rect 2 355 5 387
rect 19 386 22 392
rect 42 387 45 393
rect 54 388 57 391
rect 65 391 68 405
rect 92 400 95 405
rect 107 407 110 417
rect 137 413 140 417
rect 76 396 77 399
rect 81 396 84 399
rect 123 396 126 399
rect 65 388 73 391
rect 92 391 95 396
rect 65 383 68 388
rect 73 384 77 388
rect 100 392 111 395
rect 123 393 131 396
rect 17 377 22 382
rect 26 355 29 383
rect 56 355 59 379
rect 83 355 86 387
rect 100 386 103 392
rect 123 387 126 393
rect 135 388 138 391
rect 146 391 149 405
rect 146 388 158 391
rect 146 383 149 388
rect 98 377 103 382
rect 107 355 110 383
rect 137 355 140 379
rect -179 351 -172 355
rect -168 351 -166 355
rect -162 351 -158 355
rect -154 351 -140 355
rect -136 351 -131 355
rect -127 351 -122 355
rect -118 351 -99 355
rect -95 351 -65 355
rect -61 351 -50 355
rect -46 351 -22 355
rect -18 351 -5 355
rect -1 351 19 355
rect 23 351 73 355
rect 80 351 100 355
rect 104 351 154 355
rect -179 344 -158 348
rect -154 344 -99 348
rect -95 344 -74 348
rect -70 344 -43 348
rect -39 344 -10 348
rect -111 337 -110 341
rect -86 336 -85 340
rect -39 337 -38 341
rect -163 323 -160 328
rect -156 323 -153 328
rect -173 320 -171 323
rect -163 320 -153 323
rect -163 314 -160 320
rect -156 314 -153 320
rect -147 322 -144 328
rect -131 323 -128 328
rect -147 318 -145 322
rect -141 318 -139 322
rect -131 321 -125 323
rect -121 321 -120 323
rect -131 319 -120 321
rect -103 321 -100 328
rect -147 314 -144 318
rect -131 314 -128 319
rect -102 317 -100 321
rect -103 314 -100 317
rect -87 322 -84 328
rect -77 322 -74 328
rect -56 323 -53 328
rect -77 318 -68 322
rect -56 319 -55 323
rect -51 320 -48 323
rect -31 322 -28 328
rect -13 323 -10 328
rect 26 331 29 351
rect 107 331 110 351
rect -87 314 -84 318
rect -77 314 -74 318
rect -56 314 -53 319
rect -29 318 -28 322
rect -31 314 -28 318
rect -13 314 -10 319
rect 17 318 22 323
rect 26 319 27 322
rect 42 321 45 327
rect 42 318 50 321
rect 97 318 102 323
rect 106 319 108 322
rect 123 321 126 327
rect 123 318 131 321
rect 42 315 45 318
rect 123 315 126 318
rect -103 299 -100 303
rect -76 299 -75 303
rect -31 299 -29 303
rect -179 292 -146 296
rect -142 292 -115 296
rect -111 292 -93 296
rect -89 292 -28 296
rect -24 292 -10 296
rect 26 289 29 307
rect 107 289 110 307
rect -179 285 -173 289
rect -169 285 -157 289
rect -153 285 -139 289
rect -135 285 -128 289
rect -124 285 -122 289
rect -118 285 -103 289
rect -99 285 -66 289
rect -62 285 -61 289
rect -57 285 -49 289
rect -45 285 -21 289
rect -17 285 -5 289
rect -1 285 19 289
rect 23 285 73 289
rect 77 285 100 289
rect 104 285 162 289
rect 166 285 177 289
rect -179 278 -146 282
rect -142 278 -115 282
rect -111 278 -93 282
rect -89 278 -28 282
rect -24 278 -10 282
rect 26 275 29 285
rect 56 281 59 285
rect 107 281 110 285
rect -103 271 -100 275
rect -76 271 -75 275
rect -31 271 -29 275
rect -174 251 -171 254
rect -163 254 -160 260
rect -156 254 -153 260
rect -163 251 -153 254
rect -163 246 -160 251
rect -156 246 -153 251
rect -147 256 -144 260
rect -147 252 -145 256
rect -141 252 -139 256
rect -131 255 -128 260
rect -103 257 -100 260
rect -131 253 -120 255
rect -147 246 -144 252
rect -131 251 -125 253
rect -131 246 -128 251
rect -121 251 -120 253
rect -102 253 -100 257
rect -103 246 -100 253
rect 42 264 45 267
rect -87 256 -84 260
rect -77 256 -74 260
rect -77 252 -68 256
rect -56 255 -53 260
rect -31 256 -28 260
rect -87 246 -84 252
rect -77 246 -74 252
rect -56 251 -55 255
rect -51 251 -48 254
rect -29 252 -28 256
rect -13 255 -10 260
rect 19 260 30 263
rect 42 261 50 264
rect -56 246 -53 251
rect -31 246 -28 252
rect 19 254 22 260
rect 42 255 45 261
rect 54 256 57 259
rect 65 259 68 273
rect 116 268 119 273
rect 131 275 134 285
rect 161 281 164 285
rect 100 264 101 267
rect 105 264 108 267
rect 147 264 150 267
rect 73 259 78 264
rect 116 259 119 264
rect 65 256 73 259
rect -13 246 -10 251
rect 65 251 68 256
rect 124 260 135 263
rect 147 261 155 264
rect 17 245 22 250
rect -111 233 -110 237
rect -86 234 -85 238
rect -39 233 -38 237
rect -179 226 -158 230
rect -154 226 -99 230
rect -95 226 -74 230
rect -70 226 -43 230
rect -39 226 -10 230
rect 26 223 29 251
rect 56 223 59 247
rect 107 223 110 255
rect 124 254 127 260
rect 147 255 150 261
rect 159 256 162 259
rect 170 259 173 273
rect 170 256 176 259
rect 170 251 173 256
rect 122 245 127 250
rect 131 223 134 251
rect 161 223 164 247
rect -179 219 -172 223
rect -168 219 -166 223
rect -162 219 -158 223
rect -154 219 -140 223
rect -136 219 -131 223
rect -127 219 -122 223
rect -118 219 -99 223
rect -95 219 -65 223
rect -61 219 -50 223
rect -46 219 -22 223
rect -18 219 -5 223
rect -1 219 19 223
rect 23 219 73 223
rect 77 219 100 223
rect 104 219 124 223
rect 128 219 176 223
rect -179 212 -158 216
rect -154 212 -99 216
rect -95 212 -74 216
rect -70 212 -43 216
rect -39 212 -10 216
rect -111 205 -110 209
rect -86 204 -85 208
rect -39 205 -38 209
rect 26 200 29 219
rect 131 200 134 219
rect -163 191 -160 196
rect -156 191 -153 196
rect -173 188 -171 191
rect -163 188 -153 191
rect -163 182 -160 188
rect -156 182 -153 188
rect -147 190 -144 196
rect -131 191 -128 196
rect -147 186 -145 190
rect -141 186 -139 190
rect -131 189 -125 191
rect -121 189 -120 191
rect -131 187 -120 189
rect -103 189 -100 196
rect -147 182 -144 186
rect -131 182 -128 187
rect -102 185 -100 189
rect -103 182 -100 185
rect -87 190 -84 196
rect -77 190 -74 196
rect -56 191 -53 196
rect -77 186 -68 190
rect -56 187 -55 191
rect -51 188 -48 191
rect -31 190 -28 196
rect -13 191 -10 196
rect -87 182 -84 186
rect -77 182 -74 186
rect -56 182 -53 187
rect -29 186 -28 190
rect 16 187 21 192
rect 25 188 27 191
rect 42 190 45 196
rect 42 187 50 190
rect 122 187 127 192
rect 131 188 132 191
rect 147 190 150 196
rect 147 187 155 190
rect -31 182 -28 186
rect -13 182 -10 187
rect 42 184 45 187
rect 147 184 150 187
rect -103 167 -100 171
rect -76 167 -75 171
rect -31 167 -29 171
rect -179 160 -146 164
rect -142 160 -115 164
rect -111 160 -93 164
rect -89 160 -28 164
rect -24 160 -10 164
rect 26 157 29 176
rect 131 157 134 176
rect -179 153 -173 157
rect -169 153 -157 157
rect -153 153 -139 157
rect -135 153 -128 157
rect -124 153 -122 157
rect -118 153 -103 157
rect -99 153 -66 157
rect -62 153 -61 157
rect -57 153 -49 157
rect -45 153 -21 157
rect -17 153 -5 157
rect -1 153 19 157
rect 23 153 73 157
rect 77 153 100 157
rect 104 153 154 157
rect 158 153 162 157
rect 166 153 190 157
rect 194 153 244 157
rect -179 146 -146 150
rect -142 146 -115 150
rect -111 146 -93 150
rect -89 146 -28 150
rect -24 146 -10 150
rect 26 143 29 153
rect 56 149 59 153
rect 83 149 86 153
rect -103 139 -100 143
rect -76 139 -75 143
rect -31 139 -29 143
rect -174 119 -171 122
rect -163 122 -160 128
rect -156 122 -153 128
rect -163 119 -153 122
rect -163 114 -160 119
rect -156 114 -153 119
rect -147 124 -144 128
rect -147 120 -145 124
rect -141 120 -139 124
rect -131 123 -128 128
rect -103 125 -100 128
rect -131 121 -120 123
rect -147 114 -144 120
rect -131 119 -125 121
rect -131 114 -128 119
rect -121 119 -120 121
rect -102 121 -100 125
rect -103 114 -100 121
rect 42 132 45 135
rect -87 124 -84 128
rect -77 124 -74 128
rect -77 120 -68 124
rect -56 123 -53 128
rect -31 124 -28 128
rect -87 114 -84 120
rect -77 114 -74 120
rect -56 119 -55 123
rect -51 119 -48 122
rect -29 120 -28 124
rect -13 123 -10 128
rect 19 128 30 131
rect 42 129 50 132
rect -56 114 -53 119
rect -31 114 -28 120
rect 19 122 22 128
rect 42 123 45 129
rect 54 124 57 127
rect 65 127 68 141
rect 92 136 95 141
rect 107 143 110 153
rect 137 149 140 153
rect 173 149 176 153
rect 76 132 77 135
rect 81 132 84 135
rect 123 132 126 135
rect 65 124 73 127
rect 92 127 95 132
rect -13 114 -10 119
rect 65 119 68 124
rect 73 120 77 124
rect 100 128 111 131
rect 123 129 131 132
rect 17 113 22 118
rect -111 101 -110 105
rect -86 102 -85 106
rect -39 101 -38 105
rect -179 94 -158 98
rect -154 94 -99 98
rect -95 94 -74 98
rect -70 94 -43 98
rect -39 94 -10 98
rect 26 91 29 119
rect 56 91 59 115
rect 83 91 86 123
rect 100 122 103 128
rect 123 123 126 129
rect 135 124 138 127
rect 146 127 149 141
rect 182 136 185 141
rect 197 143 200 153
rect 227 149 230 153
rect 171 132 174 135
rect 213 132 216 135
rect 146 124 155 127
rect 182 127 185 132
rect 146 119 149 124
rect 98 113 103 118
rect 107 91 110 119
rect 189 130 201 131
rect 193 128 201 130
rect 213 129 221 132
rect 213 123 216 129
rect 225 124 228 127
rect 236 127 239 141
rect 236 124 248 127
rect 137 91 140 115
rect 173 91 176 123
rect 236 119 239 124
rect 197 91 200 119
rect 227 91 230 115
rect -179 87 -172 91
rect -168 87 -166 91
rect -162 87 -158 91
rect -154 87 -140 91
rect -136 87 -131 91
rect -127 87 -122 91
rect -118 87 -99 91
rect -95 87 -65 91
rect -61 87 -50 91
rect -46 87 -22 91
rect -18 87 -5 91
rect -1 87 19 91
rect 23 87 73 91
rect 80 87 100 91
rect 104 87 154 91
rect 158 87 190 91
rect 194 87 244 91
rect -179 80 -158 84
rect -154 80 -99 84
rect -95 80 -74 84
rect -70 80 -43 84
rect -39 80 -10 84
rect -111 73 -110 77
rect -86 72 -85 76
rect -39 73 -38 77
rect -163 59 -160 64
rect -156 59 -153 64
rect -173 56 -171 59
rect -163 56 -153 59
rect -163 50 -160 56
rect -156 50 -153 56
rect -147 58 -144 64
rect -131 59 -128 64
rect -147 54 -145 58
rect -141 54 -139 58
rect -131 57 -125 59
rect -121 57 -120 59
rect -131 55 -120 57
rect -103 57 -100 64
rect -147 50 -144 54
rect -131 50 -128 55
rect -102 53 -100 57
rect -103 50 -100 53
rect -87 58 -84 64
rect -77 58 -74 64
rect -56 59 -53 64
rect -77 54 -68 58
rect -56 55 -55 59
rect -51 56 -48 59
rect -31 58 -28 64
rect -13 59 -10 64
rect 26 65 29 87
rect 107 65 110 87
rect 197 65 200 87
rect -87 50 -84 54
rect -77 50 -74 54
rect -56 50 -53 55
rect -29 54 -28 58
rect -31 50 -28 54
rect -13 50 -10 55
rect 17 52 22 57
rect 26 53 27 56
rect 42 55 45 61
rect 42 52 50 55
rect 97 52 102 57
rect 106 53 108 56
rect 123 55 126 61
rect 123 52 131 55
rect 190 53 198 56
rect 213 55 216 61
rect 213 52 221 55
rect 42 49 45 52
rect 123 49 126 52
rect 213 49 216 52
rect -103 35 -100 39
rect -76 35 -75 39
rect -31 35 -29 39
rect -179 28 -146 32
rect -142 28 -115 32
rect -111 28 -93 32
rect -89 28 -28 32
rect -24 28 -10 32
rect 26 25 29 41
rect 107 25 110 41
rect 197 25 200 41
rect -179 21 -173 25
rect -169 21 -157 25
rect -153 21 -139 25
rect -135 21 -128 25
rect -124 21 -122 25
rect -118 21 -103 25
rect -99 21 -66 25
rect -62 21 -61 25
rect -57 21 -49 25
rect -45 21 -21 25
rect -17 21 -5 25
rect -1 21 19 25
rect 23 21 73 25
rect 77 21 100 25
rect 104 21 190 25
rect 194 21 248 25
rect -179 14 -146 18
rect -142 14 -115 18
rect -111 14 -93 18
rect -89 14 -28 18
rect -24 14 -10 18
rect 26 11 29 21
rect 56 17 59 21
rect -103 7 -100 11
rect -76 7 -75 11
rect -31 7 -29 11
rect -174 -13 -171 -10
rect -163 -10 -160 -4
rect -156 -10 -153 -4
rect -163 -13 -153 -10
rect -163 -18 -160 -13
rect -156 -18 -153 -13
rect -147 -8 -144 -4
rect -147 -12 -145 -8
rect -141 -12 -139 -8
rect -131 -9 -128 -4
rect -103 -7 -100 -4
rect -131 -11 -120 -9
rect -147 -18 -144 -12
rect -131 -13 -125 -11
rect -131 -18 -128 -13
rect -121 -13 -120 -11
rect -102 -11 -100 -7
rect -103 -18 -100 -11
rect 42 0 45 3
rect -87 -8 -84 -4
rect -77 -8 -74 -4
rect -77 -12 -68 -8
rect -56 -9 -53 -4
rect -31 -8 -28 -4
rect -87 -18 -84 -12
rect -77 -18 -74 -12
rect -56 -13 -55 -9
rect -51 -13 -48 -10
rect -29 -12 -28 -8
rect -13 -9 -10 -4
rect 19 -4 30 -1
rect 42 -3 50 0
rect -56 -18 -53 -13
rect -31 -18 -28 -12
rect 19 -10 22 -4
rect 42 -9 45 -3
rect 54 -8 57 -5
rect 65 -5 68 9
rect 73 -5 78 0
rect 65 -8 73 -5
rect -13 -18 -10 -13
rect 65 -13 68 -8
rect 17 -19 22 -14
rect -111 -31 -110 -27
rect -86 -30 -85 -26
rect -39 -31 -38 -27
rect -179 -38 -158 -34
rect -154 -38 -99 -34
rect -95 -38 -74 -34
rect -70 -38 -43 -34
rect -39 -38 -10 -34
rect 26 -41 29 -13
rect 56 -41 59 -17
rect -179 -45 -172 -41
rect -168 -45 -166 -41
rect -162 -45 -158 -41
rect -154 -45 -140 -41
rect -136 -45 -131 -41
rect -127 -45 -122 -41
rect -118 -45 -99 -41
rect -95 -45 -65 -41
rect -61 -45 -50 -41
rect -46 -45 -22 -41
rect -18 -45 -5 -41
rect -1 -45 19 -41
rect 23 -45 94 -41
rect 98 -45 153 -41
rect 157 -45 178 -41
rect 182 -45 209 -41
rect 213 -45 242 -41
rect -179 -52 -158 -48
rect -154 -52 -99 -48
rect -95 -52 -74 -48
rect -70 -52 -43 -48
rect -39 -52 -10 -48
rect -111 -59 -110 -55
rect -86 -60 -85 -56
rect -39 -59 -38 -55
rect -163 -73 -160 -68
rect -156 -73 -153 -68
rect -173 -76 -171 -73
rect -163 -76 -153 -73
rect -163 -82 -160 -76
rect -156 -82 -153 -76
rect -147 -74 -144 -68
rect -131 -73 -128 -68
rect -147 -78 -145 -74
rect -141 -78 -139 -74
rect -131 -75 -125 -73
rect -121 -75 -120 -73
rect -131 -77 -120 -75
rect -103 -75 -100 -68
rect -147 -82 -144 -78
rect -131 -82 -128 -77
rect -102 -79 -100 -75
rect -103 -82 -100 -79
rect -87 -74 -84 -68
rect -77 -74 -74 -68
rect -56 -73 -53 -68
rect -77 -78 -68 -74
rect -56 -77 -55 -73
rect -51 -76 -48 -73
rect -31 -74 -28 -68
rect -13 -73 -10 -68
rect 26 -71 29 -45
rect 62 -52 92 -48
rect 96 -52 121 -48
rect 125 -52 157 -48
rect 161 -52 196 -48
rect 200 -52 242 -48
rect 62 -64 65 -52
rect 112 -64 115 -52
rect 131 -64 134 -52
rect 141 -59 142 -55
rect 166 -60 167 -56
rect 187 -64 190 -52
rect 203 -64 206 -52
rect 213 -59 214 -55
rect 230 -64 233 -52
rect -87 -82 -84 -78
rect -77 -82 -74 -78
rect -56 -82 -53 -77
rect -29 -78 -28 -74
rect 89 -73 92 -68
rect 96 -73 99 -68
rect -31 -82 -28 -78
rect -13 -82 -10 -77
rect 16 -84 21 -79
rect 25 -83 27 -80
rect 42 -81 45 -75
rect 74 -76 99 -73
rect 42 -84 50 -81
rect 42 -87 45 -84
rect -103 -97 -100 -93
rect -76 -97 -75 -93
rect -31 -97 -29 -93
rect 74 -90 77 -76
rect 96 -82 99 -76
rect 105 -74 108 -68
rect 121 -73 124 -68
rect 105 -78 107 -74
rect 111 -78 113 -74
rect 121 -75 127 -73
rect 131 -75 132 -73
rect 121 -77 132 -75
rect 149 -75 152 -68
rect 105 -82 108 -78
rect 121 -82 124 -77
rect 150 -79 152 -75
rect 149 -82 152 -79
rect 165 -74 168 -68
rect 175 -74 178 -68
rect 196 -73 199 -68
rect 175 -78 184 -74
rect 196 -77 197 -73
rect 201 -76 204 -73
rect 221 -74 224 -68
rect 165 -82 168 -78
rect 175 -82 178 -78
rect 196 -82 199 -77
rect 223 -78 224 -74
rect 239 -74 242 -68
rect 221 -82 224 -78
rect 239 -82 242 -78
rect -179 -104 -146 -100
rect -142 -104 -115 -100
rect -111 -104 -93 -100
rect -89 -104 -28 -100
rect -24 -104 -10 -100
rect 26 -107 29 -95
rect 62 -100 66 -90
rect 89 -100 92 -90
rect 112 -100 115 -90
rect 131 -100 134 -90
rect 149 -97 152 -93
rect 176 -97 177 -93
rect 187 -100 190 -90
rect 203 -100 206 -90
rect 221 -97 223 -93
rect 230 -100 233 -90
rect 62 -104 89 -100
rect 93 -104 121 -100
rect 125 -104 157 -100
rect 161 -104 196 -100
rect 200 -104 242 -100
rect -179 -111 -173 -107
rect -169 -111 -157 -107
rect -153 -111 -139 -107
rect -135 -111 -128 -107
rect -124 -111 -122 -107
rect -118 -111 -103 -107
rect -99 -111 -66 -107
rect -62 -111 -61 -107
rect -57 -111 -49 -107
rect -45 -111 -21 -107
rect -17 -111 19 -107
rect 23 -111 73 -107
rect 77 -111 105 -107
rect 109 -111 134 -107
rect 138 -111 159 -107
rect 163 -111 223 -107
rect 227 -111 242 -107
<< m2contact >>
rect -173 417 -169 421
rect -139 417 -135 421
rect -122 417 -118 421
rect -66 417 -62 421
rect -49 417 -45 421
rect -21 417 -17 421
rect -146 410 -142 414
rect -115 410 -111 414
rect -93 410 -89 414
rect -28 410 -24 414
rect -172 400 -168 404
rect -147 403 -143 407
rect -140 400 -136 404
rect -122 400 -118 404
rect -100 403 -96 407
rect -75 403 -71 407
rect -65 400 -61 404
rect -49 400 -45 404
rect -29 403 -25 407
rect -22 400 -18 404
rect 42 410 46 414
rect -145 384 -141 388
rect -125 381 -121 385
rect -106 385 -102 389
rect -4 396 0 400
rect 11 396 15 400
rect -87 384 -83 388
rect -68 384 -64 388
rect -55 383 -51 387
rect -33 384 -29 388
rect -25 383 -21 387
rect -13 383 -9 387
rect -172 370 -168 374
rect -140 370 -136 374
rect -122 370 -118 374
rect -65 370 -61 374
rect -50 370 -46 374
rect -22 370 -18 374
rect -158 366 -154 370
rect -115 365 -111 369
rect -93 366 -86 370
rect -43 365 -39 369
rect -158 358 -154 362
rect -99 358 -95 362
rect -74 358 -70 362
rect -43 358 -39 362
rect 50 388 54 396
rect 123 410 127 414
rect 77 396 81 400
rect 92 396 96 400
rect 73 388 77 392
rect 19 382 23 386
rect 32 374 36 378
rect 131 388 135 396
rect 158 388 162 392
rect 100 382 104 386
rect 113 374 117 378
rect -172 351 -168 355
rect -158 351 -154 355
rect -140 351 -136 355
rect -122 351 -118 355
rect -99 351 -95 355
rect -65 351 -61 355
rect -50 351 -46 355
rect -22 351 -18 355
rect -158 344 -154 348
rect -99 344 -95 348
rect -74 344 -70 348
rect -43 344 -39 348
rect -158 336 -154 340
rect -115 337 -111 341
rect -93 336 -86 340
rect -43 337 -39 341
rect -172 332 -168 336
rect -140 332 -136 336
rect -122 332 -118 336
rect -65 332 -61 336
rect -50 332 -46 336
rect -22 332 -18 336
rect -177 320 -173 324
rect -145 318 -141 322
rect -125 321 -121 325
rect -106 317 -102 321
rect -87 318 -83 322
rect -68 318 -64 322
rect -55 319 -51 323
rect 42 334 46 338
rect 123 334 127 338
rect -33 318 -29 322
rect -25 319 -21 323
rect -13 319 -9 323
rect 22 319 26 323
rect 50 318 54 322
rect 102 319 106 323
rect 131 318 135 322
rect -172 302 -168 306
rect -147 299 -143 303
rect -140 302 -136 306
rect -122 302 -118 306
rect -100 299 -96 303
rect -75 299 -71 303
rect -65 302 -61 306
rect -49 302 -45 306
rect -29 299 -25 303
rect -22 302 -18 306
rect -146 292 -142 296
rect -115 292 -111 296
rect -93 292 -89 296
rect -28 292 -24 296
rect 32 298 36 302
rect 113 298 117 302
rect -173 285 -169 289
rect -139 285 -135 289
rect -122 285 -118 289
rect -66 285 -62 289
rect -49 285 -45 289
rect -21 285 -17 289
rect -146 278 -142 282
rect -115 278 -111 282
rect -93 278 -89 282
rect -28 278 -24 282
rect 42 278 46 282
rect -172 268 -168 272
rect -147 271 -143 275
rect -140 268 -136 272
rect -122 268 -118 272
rect -100 271 -96 275
rect -75 271 -71 275
rect -65 268 -61 272
rect -49 268 -45 272
rect -29 271 -25 275
rect -22 268 -18 272
rect -178 251 -174 255
rect -145 252 -141 256
rect -125 249 -121 253
rect -106 253 -102 257
rect -87 252 -83 256
rect -68 252 -64 256
rect -55 251 -51 255
rect -33 252 -29 256
rect -25 251 -21 255
rect -13 251 -9 255
rect 50 256 54 264
rect 147 278 151 282
rect 101 264 105 268
rect 116 264 120 268
rect 19 250 23 254
rect 73 255 77 259
rect -172 238 -168 242
rect -140 238 -136 242
rect -122 238 -118 242
rect -65 238 -61 242
rect -50 238 -46 242
rect -22 238 -18 242
rect -158 234 -154 238
rect -115 233 -111 237
rect -93 234 -86 238
rect -43 233 -39 237
rect -158 226 -154 230
rect -99 226 -95 230
rect -74 226 -70 230
rect -43 226 -39 230
rect 32 242 36 246
rect 155 256 159 264
rect 176 256 180 260
rect 124 250 128 254
rect 137 242 141 246
rect -172 219 -168 223
rect -158 219 -154 223
rect -140 219 -136 223
rect -122 219 -118 223
rect -99 219 -95 223
rect -65 219 -61 223
rect -50 219 -46 223
rect -22 219 -18 223
rect -158 212 -154 216
rect -99 212 -95 216
rect -74 212 -70 216
rect -43 212 -39 216
rect -158 204 -154 208
rect -115 205 -111 209
rect -93 204 -86 208
rect -43 205 -39 209
rect -172 200 -168 204
rect -140 200 -136 204
rect -122 200 -118 204
rect -65 200 -61 204
rect -50 200 -46 204
rect -22 200 -18 204
rect 42 203 46 207
rect 147 203 151 207
rect -177 188 -173 192
rect -145 186 -141 190
rect -125 189 -121 193
rect -106 185 -102 189
rect -87 186 -83 190
rect -68 186 -64 190
rect -55 187 -51 191
rect -33 186 -29 190
rect -25 187 -21 191
rect -13 187 -9 191
rect 21 188 25 192
rect 50 187 54 191
rect 127 188 131 192
rect 155 187 159 191
rect -172 170 -168 174
rect -147 167 -143 171
rect -140 170 -136 174
rect -122 170 -118 174
rect -100 167 -96 171
rect -75 167 -71 171
rect -65 170 -61 174
rect -49 170 -45 174
rect -29 167 -25 171
rect -22 170 -18 174
rect -146 160 -142 164
rect -115 160 -111 164
rect -93 160 -89 164
rect -28 160 -24 164
rect 32 167 36 171
rect 137 167 141 171
rect -173 153 -169 157
rect -139 153 -135 157
rect -122 153 -118 157
rect -66 153 -62 157
rect -49 153 -45 157
rect -21 153 -17 157
rect -146 146 -142 150
rect -115 146 -111 150
rect -93 146 -89 150
rect -28 146 -24 150
rect 42 146 46 150
rect -172 136 -168 140
rect -147 139 -143 143
rect -140 136 -136 140
rect -122 136 -118 140
rect -100 139 -96 143
rect -75 139 -71 143
rect -65 136 -61 140
rect -49 136 -45 140
rect -29 139 -25 143
rect -22 136 -18 140
rect -178 119 -174 123
rect -145 120 -141 124
rect -125 117 -121 121
rect -106 121 -102 125
rect -87 120 -83 124
rect -68 120 -64 124
rect -55 119 -51 123
rect -33 120 -29 124
rect -25 119 -21 123
rect -13 119 -9 123
rect 50 124 54 132
rect 123 146 127 150
rect 77 132 81 136
rect 92 132 96 136
rect 73 124 77 128
rect 19 118 23 122
rect -172 106 -168 110
rect -140 106 -136 110
rect -122 106 -118 110
rect -65 106 -61 110
rect -50 106 -46 110
rect -22 106 -18 110
rect -158 102 -154 106
rect -115 101 -111 105
rect -93 102 -86 106
rect -43 101 -39 105
rect -158 94 -154 98
rect -99 94 -95 98
rect -74 94 -70 98
rect -43 94 -39 98
rect 32 110 36 114
rect 131 124 135 132
rect 213 146 217 150
rect 167 132 171 136
rect 182 132 186 136
rect 155 124 159 128
rect 100 118 104 122
rect 189 126 193 130
rect 221 124 225 132
rect 113 110 117 114
rect 203 110 207 114
rect -172 87 -168 91
rect -158 87 -154 91
rect -140 87 -136 91
rect -122 87 -118 91
rect -99 87 -95 91
rect -65 87 -61 91
rect -50 87 -46 91
rect -22 87 -18 91
rect -158 80 -154 84
rect -99 80 -95 84
rect -74 80 -70 84
rect -43 80 -39 84
rect -158 72 -154 76
rect -115 73 -111 77
rect -93 72 -86 76
rect -43 73 -39 77
rect -172 68 -168 72
rect -140 68 -136 72
rect -122 68 -118 72
rect -65 68 -61 72
rect -50 68 -46 72
rect -22 68 -18 72
rect -177 56 -173 60
rect -145 54 -141 58
rect -125 57 -121 61
rect -106 53 -102 57
rect -87 54 -83 58
rect -68 54 -64 58
rect -55 55 -51 59
rect 42 68 46 72
rect 123 68 127 72
rect 213 68 217 72
rect -33 54 -29 58
rect -25 55 -21 59
rect -13 55 -9 59
rect 22 53 26 57
rect 50 52 54 56
rect 102 53 106 57
rect 131 52 135 56
rect 186 53 190 57
rect 221 52 225 56
rect -172 38 -168 42
rect -147 35 -143 39
rect -140 38 -136 42
rect -122 38 -118 42
rect -100 35 -96 39
rect -75 35 -71 39
rect -65 38 -61 42
rect -49 38 -45 42
rect -29 35 -25 39
rect -22 38 -18 42
rect -146 28 -142 32
rect -115 28 -111 32
rect -93 28 -89 32
rect -28 28 -24 32
rect 32 32 36 36
rect 113 32 117 36
rect 203 32 207 36
rect -173 21 -169 25
rect -139 21 -135 25
rect -122 21 -118 25
rect -66 21 -62 25
rect -49 21 -45 25
rect -21 21 -17 25
rect -146 14 -142 18
rect -115 14 -111 18
rect -93 14 -89 18
rect -28 14 -24 18
rect 42 14 46 18
rect -172 4 -168 8
rect -147 7 -143 11
rect -140 4 -136 8
rect -122 4 -118 8
rect -100 7 -96 11
rect -75 7 -71 11
rect -65 4 -61 8
rect -49 4 -45 8
rect -29 7 -25 11
rect -22 4 -18 8
rect -178 -13 -174 -9
rect -145 -12 -141 -8
rect -125 -15 -121 -11
rect -106 -11 -102 -7
rect -87 -12 -83 -8
rect -68 -12 -64 -8
rect -55 -13 -51 -9
rect -33 -12 -29 -8
rect -25 -13 -21 -9
rect -13 -13 -9 -9
rect 50 -8 54 0
rect 19 -14 23 -10
rect 73 -9 77 -5
rect -172 -26 -168 -22
rect -140 -26 -136 -22
rect -122 -26 -118 -22
rect -65 -26 -61 -22
rect -50 -26 -46 -22
rect -22 -26 -18 -22
rect -158 -30 -154 -26
rect -115 -31 -111 -27
rect -93 -30 -86 -26
rect -43 -31 -39 -27
rect -158 -38 -154 -34
rect -99 -38 -95 -34
rect -74 -38 -70 -34
rect -43 -38 -39 -34
rect 32 -22 36 -18
rect -172 -45 -168 -41
rect -158 -45 -154 -41
rect -140 -45 -136 -41
rect -122 -45 -118 -41
rect -99 -45 -95 -41
rect -65 -45 -61 -41
rect -50 -45 -46 -41
rect -22 -45 -18 -41
rect 94 -45 98 -41
rect 153 -45 157 -41
rect 178 -45 182 -41
rect 209 -45 213 -41
rect -158 -52 -154 -48
rect -99 -52 -95 -48
rect -74 -52 -70 -48
rect -43 -52 -39 -48
rect -158 -60 -154 -56
rect -115 -59 -111 -55
rect -93 -60 -86 -56
rect -43 -59 -39 -55
rect -172 -64 -168 -60
rect -140 -64 -136 -60
rect -122 -64 -118 -60
rect -65 -64 -61 -60
rect -50 -64 -46 -60
rect -22 -64 -18 -60
rect -177 -76 -173 -72
rect -145 -78 -141 -74
rect -125 -75 -121 -71
rect -106 -79 -102 -75
rect -87 -78 -83 -74
rect -68 -78 -64 -74
rect -55 -77 -51 -73
rect 94 -60 98 -56
rect 137 -59 141 -55
rect 159 -60 166 -56
rect 209 -59 213 -55
rect 42 -68 46 -64
rect -33 -78 -29 -74
rect -25 -77 -21 -73
rect -13 -77 -9 -73
rect 21 -83 25 -79
rect 61 -77 65 -73
rect 50 -84 54 -80
rect -172 -94 -168 -90
rect -147 -97 -143 -93
rect -140 -94 -136 -90
rect -122 -94 -118 -90
rect -100 -97 -96 -93
rect -75 -97 -71 -93
rect -65 -94 -61 -90
rect -49 -94 -45 -90
rect -29 -97 -25 -93
rect -22 -94 -18 -90
rect 107 -78 111 -74
rect 127 -75 131 -71
rect 146 -79 150 -75
rect 165 -78 169 -74
rect 184 -78 188 -74
rect 197 -77 201 -73
rect 219 -78 223 -74
rect 227 -77 231 -73
rect 239 -78 243 -74
rect -146 -104 -142 -100
rect -115 -104 -111 -100
rect -93 -104 -89 -100
rect -28 -104 -24 -100
rect 105 -97 109 -93
rect 152 -97 156 -93
rect 177 -97 181 -93
rect 223 -97 227 -93
rect 32 -104 36 -100
rect -173 -111 -169 -107
rect -139 -111 -135 -107
rect -122 -111 -118 -107
rect -66 -111 -62 -107
rect -49 -111 -45 -107
rect -21 -111 -17 -107
rect 105 -111 109 -107
rect 134 -111 138 -107
rect 159 -111 163 -107
rect 223 -111 227 -107
<< metal2 >>
rect -172 404 -169 417
rect -146 407 -143 410
rect -139 404 -136 417
rect -122 404 -119 417
rect -172 355 -169 370
rect -158 362 -155 366
rect -140 355 -137 370
rect -121 355 -118 370
rect -115 369 -112 410
rect -99 362 -96 403
rect -93 370 -90 410
rect -74 362 -71 403
rect -65 404 -62 417
rect -49 404 -46 417
rect -28 407 -25 410
rect -21 404 -18 417
rect -3 413 0 426
rect -3 410 42 413
rect -3 400 0 410
rect 15 397 35 400
rect 32 378 35 397
rect -65 355 -62 370
rect -50 355 -47 370
rect -43 362 -39 365
rect -22 355 -19 370
rect -172 336 -169 351
rect -158 340 -155 344
rect -140 336 -137 351
rect -121 336 -118 351
rect -172 289 -169 302
rect -146 296 -143 299
rect -172 272 -169 285
rect -139 289 -136 302
rect -122 289 -119 302
rect -115 296 -112 337
rect -99 303 -96 344
rect -93 296 -90 336
rect -74 303 -71 344
rect -65 336 -62 351
rect -50 336 -47 351
rect -43 341 -39 344
rect -22 336 -19 351
rect -65 289 -62 302
rect -146 275 -143 278
rect -139 272 -136 285
rect -122 272 -119 285
rect -172 223 -169 238
rect -158 230 -155 234
rect -140 223 -137 238
rect -121 223 -118 238
rect -115 237 -112 278
rect -99 230 -96 271
rect -93 238 -90 278
rect -74 230 -71 271
rect -65 272 -62 285
rect -49 289 -46 302
rect -28 296 -25 299
rect -21 289 -18 302
rect 32 302 35 374
rect 43 338 46 410
rect 78 413 81 426
rect 78 410 123 413
rect 78 400 81 410
rect -49 272 -46 285
rect -28 275 -25 278
rect -21 272 -18 285
rect 32 268 35 298
rect 43 282 46 334
rect 50 322 54 388
rect 38 278 42 281
rect 31 265 35 268
rect 32 246 35 265
rect -65 223 -62 238
rect -50 223 -47 238
rect -43 230 -39 233
rect -22 223 -19 238
rect -172 204 -169 219
rect -158 208 -155 212
rect -140 204 -137 219
rect -121 204 -118 219
rect -172 157 -169 170
rect -146 164 -143 167
rect -172 140 -169 153
rect -139 157 -136 170
rect -122 157 -119 170
rect -115 164 -112 205
rect -99 171 -96 212
rect -93 164 -90 204
rect -74 171 -71 212
rect -65 204 -62 219
rect -50 204 -47 219
rect -43 209 -39 212
rect -22 204 -19 219
rect -65 157 -62 170
rect -146 143 -143 146
rect -139 140 -136 153
rect -122 140 -119 153
rect -172 91 -169 106
rect -158 98 -155 102
rect -140 91 -137 106
rect -121 91 -118 106
rect -115 105 -112 146
rect -99 98 -96 139
rect -93 106 -90 146
rect -74 98 -71 139
rect -65 140 -62 153
rect -49 157 -46 170
rect -28 164 -25 167
rect -21 157 -18 170
rect 32 171 35 242
rect 43 207 46 278
rect -49 140 -46 153
rect -28 143 -25 146
rect -21 140 -18 153
rect 32 114 35 167
rect 43 150 46 203
rect 50 191 54 256
rect 38 146 42 149
rect 81 149 84 400
rect 96 397 116 400
rect 113 378 116 397
rect 113 302 116 374
rect 124 338 127 410
rect 131 322 135 388
rect 140 289 143 426
rect 102 285 143 289
rect 102 281 105 285
rect 102 278 147 281
rect 102 268 105 278
rect 120 265 140 268
rect 102 263 105 264
rect 137 246 140 265
rect 137 171 140 242
rect 148 207 151 278
rect 155 191 159 256
rect -65 91 -62 106
rect -50 91 -47 106
rect -43 98 -39 101
rect -22 91 -19 106
rect -172 72 -169 87
rect -158 76 -155 80
rect -140 72 -137 87
rect -121 72 -118 87
rect -172 25 -169 38
rect -146 32 -143 35
rect -172 8 -169 21
rect -139 25 -136 38
rect -122 25 -119 38
rect -115 32 -112 73
rect -99 39 -96 80
rect -93 32 -90 72
rect -74 39 -71 80
rect -65 72 -62 87
rect -50 72 -47 87
rect -43 77 -39 80
rect -22 72 -19 87
rect -65 25 -62 38
rect -146 11 -143 14
rect -139 8 -136 21
rect -122 8 -119 21
rect -172 -41 -169 -26
rect -158 -34 -155 -30
rect -140 -41 -137 -26
rect -121 -41 -118 -26
rect -115 -27 -112 14
rect -99 -34 -96 7
rect -93 -26 -90 14
rect -74 -34 -71 7
rect -65 8 -62 21
rect -49 25 -46 38
rect -28 32 -25 35
rect -21 25 -18 38
rect 32 36 35 110
rect 43 72 46 146
rect 78 146 123 149
rect 78 136 81 146
rect 96 133 116 136
rect -49 8 -46 21
rect -28 11 -25 14
rect -21 8 -18 21
rect 32 -18 35 32
rect 43 18 46 68
rect 50 56 54 124
rect 113 114 116 133
rect 113 36 116 110
rect 124 72 127 146
rect 168 149 171 426
rect 168 146 213 149
rect 168 136 171 146
rect 186 133 206 136
rect 131 56 135 124
rect 203 114 206 133
rect 203 36 206 110
rect 214 72 217 146
rect 221 56 225 124
rect 38 14 42 17
rect -65 -41 -62 -26
rect -50 -41 -47 -26
rect -43 -34 -39 -31
rect -22 -41 -19 -26
rect -172 -60 -169 -45
rect -158 -56 -155 -52
rect -140 -60 -137 -45
rect -121 -60 -118 -45
rect -172 -107 -169 -94
rect -146 -100 -143 -97
rect -139 -107 -136 -94
rect -122 -107 -119 -94
rect -115 -100 -112 -59
rect -99 -93 -96 -52
rect -93 -100 -90 -60
rect -74 -93 -71 -52
rect -65 -60 -62 -45
rect -50 -60 -47 -45
rect -43 -55 -39 -52
rect -22 -60 -19 -45
rect -65 -107 -62 -94
rect -49 -107 -46 -94
rect -28 -100 -25 -97
rect -21 -107 -18 -94
rect 32 -100 35 -22
rect 43 -64 46 14
rect 50 -80 54 -8
rect 94 -56 97 -45
rect 106 -107 109 -97
rect 134 -107 137 -55
rect 153 -93 156 -45
rect 159 -107 162 -60
rect 178 -93 181 -45
rect 209 -55 213 -45
rect 224 -107 227 -97
<< m3contact >>
rect -141 384 -136 389
rect -130 380 -125 385
rect -107 389 -102 394
rect -83 384 -78 389
rect -68 388 -63 394
rect -38 384 -33 389
rect -9 383 -4 388
rect -54 378 -49 383
rect -25 378 -21 383
rect 17 377 22 382
rect -177 324 -172 329
rect -141 317 -136 322
rect -130 321 -125 326
rect -107 312 -102 317
rect -83 317 -78 322
rect -54 323 -49 328
rect -25 323 -21 328
rect -68 312 -63 318
rect -38 317 -33 322
rect -9 318 -4 323
rect 17 318 22 323
rect -178 255 -173 260
rect -141 252 -136 257
rect -130 248 -125 253
rect -107 257 -102 262
rect -83 252 -78 257
rect 73 383 78 388
rect -68 256 -63 262
rect -38 252 -33 257
rect -9 251 -4 256
rect -54 246 -49 251
rect -25 246 -21 251
rect 17 245 22 250
rect -177 192 -172 197
rect -141 185 -136 190
rect -130 189 -125 194
rect -107 180 -102 185
rect -83 185 -78 190
rect -54 191 -49 196
rect -25 191 -21 196
rect -68 180 -63 186
rect -38 185 -33 190
rect -9 186 -4 191
rect 16 187 21 192
rect -178 123 -173 128
rect -141 120 -136 125
rect -130 116 -125 121
rect -107 125 -102 130
rect -83 120 -78 125
rect -68 124 -63 130
rect -38 120 -33 125
rect -9 119 -4 124
rect -54 114 -49 119
rect -25 114 -21 119
rect 17 113 22 118
rect 73 259 78 264
rect 98 377 103 382
rect 97 318 102 323
rect 158 383 163 388
rect 122 245 127 250
rect 122 187 127 192
rect -177 60 -172 65
rect -141 53 -136 58
rect -130 57 -125 62
rect -107 48 -102 53
rect -83 53 -78 58
rect -54 59 -49 64
rect -25 59 -21 64
rect -68 48 -63 54
rect -38 53 -33 58
rect -9 54 -4 59
rect 17 52 22 57
rect -178 -9 -173 -4
rect -141 -12 -136 -7
rect -130 -16 -125 -11
rect -107 -7 -102 -2
rect -83 -12 -78 -7
rect -68 -8 -63 -2
rect -38 -12 -33 -7
rect -9 -13 -4 -8
rect -54 -18 -49 -13
rect -25 -18 -21 -13
rect 17 -19 22 -14
rect 73 119 78 124
rect 98 113 103 118
rect 97 52 102 57
rect 180 256 185 261
rect 155 128 160 133
rect 189 121 194 126
rect 186 48 191 53
rect -177 -72 -172 -67
rect -141 -79 -136 -74
rect -130 -75 -125 -70
rect -107 -84 -102 -79
rect -83 -79 -78 -74
rect -54 -73 -49 -68
rect -25 -73 -21 -68
rect -68 -84 -63 -78
rect -38 -79 -33 -74
rect -9 -78 -4 -73
rect 16 -84 21 -79
rect 73 -5 78 0
rect 61 -73 66 -68
rect 126 -71 131 -66
rect 111 -79 116 -74
rect 141 -79 146 -74
rect 169 -79 174 -74
rect 198 -73 203 -68
rect 227 -73 231 -68
rect 184 -84 189 -78
rect 214 -79 219 -74
rect 243 -78 248 -73
<< metal3 >>
rect -141 394 -101 395
rect -141 390 -107 394
rect -142 389 -135 390
rect -142 384 -141 389
rect -136 384 -135 389
rect -108 389 -107 390
rect -102 389 -101 394
rect -69 394 -33 399
rect -108 388 -101 389
rect -84 389 -77 390
rect -142 383 -135 384
rect -131 385 -124 386
rect -131 380 -130 385
rect -125 380 -124 385
rect -84 384 -83 389
rect -78 384 -77 389
rect -69 388 -68 394
rect -63 393 -33 394
rect -63 388 -62 393
rect -38 390 -33 393
rect -69 387 -62 388
rect -39 389 -32 390
rect -39 384 -38 389
rect -33 384 -32 389
rect -10 388 -3 389
rect -84 383 -77 384
rect -55 383 -48 384
rect -39 383 -32 384
rect -26 383 -20 384
rect -83 380 -78 383
rect -131 375 -78 380
rect -55 378 -54 383
rect -49 378 -48 383
rect -26 378 -25 383
rect -21 378 -20 383
rect -55 377 -20 378
rect -54 373 -20 377
rect -10 383 -9 388
rect -4 383 -3 388
rect 72 388 79 389
rect 72 383 73 388
rect 78 383 79 388
rect 157 388 164 389
rect 157 383 158 388
rect 163 383 164 388
rect -10 382 -3 383
rect 16 382 23 383
rect 72 382 79 383
rect 97 382 104 383
rect 157 382 164 383
rect -10 377 17 382
rect 22 377 23 382
rect 73 377 98 382
rect 103 377 104 382
rect -10 356 -5 377
rect 16 376 23 377
rect 97 376 104 377
rect 154 377 163 382
rect -177 350 -5 356
rect -177 330 -172 350
rect -178 329 -171 330
rect -178 324 -177 329
rect -172 324 -171 329
rect -178 323 -171 324
rect -131 326 -78 331
rect -54 329 -20 333
rect -142 322 -135 323
rect -142 317 -141 322
rect -136 317 -135 322
rect -131 321 -130 326
rect -125 321 -124 326
rect -83 323 -78 326
rect -55 328 -20 329
rect -55 323 -54 328
rect -49 323 -48 328
rect -26 323 -25 328
rect -21 323 -20 328
rect -131 320 -124 321
rect -84 322 -77 323
rect -55 322 -48 323
rect -39 322 -32 323
rect -26 322 -20 323
rect -10 323 -3 324
rect 16 323 23 324
rect 96 323 103 324
rect -142 316 -135 317
rect -108 317 -101 318
rect -108 316 -107 317
rect -141 312 -107 316
rect -102 312 -101 317
rect -84 317 -83 322
rect -78 317 -77 322
rect -84 316 -77 317
rect -69 318 -62 319
rect -141 311 -101 312
rect -69 312 -68 318
rect -63 313 -62 318
rect -39 317 -38 322
rect -33 317 -32 322
rect -10 318 -9 323
rect -4 318 17 323
rect 22 318 23 323
rect -10 317 -3 318
rect 16 317 23 318
rect 73 318 97 323
rect 102 318 103 323
rect -39 316 -32 317
rect -38 313 -33 316
rect -63 312 -33 313
rect -69 307 -33 312
rect -9 290 -4 317
rect -178 284 -4 290
rect -178 261 -173 284
rect -141 262 -101 263
rect -179 260 -172 261
rect -179 255 -178 260
rect -173 255 -172 260
rect -141 258 -107 262
rect -179 254 -172 255
rect -142 257 -135 258
rect -142 252 -141 257
rect -136 252 -135 257
rect -108 257 -107 258
rect -102 257 -101 262
rect -69 262 -33 267
rect 73 265 78 318
rect 96 317 103 318
rect 154 289 159 377
rect 116 284 159 289
rect -108 256 -101 257
rect -84 257 -77 258
rect -142 251 -135 252
rect -131 253 -124 254
rect -131 248 -130 253
rect -125 248 -124 253
rect -84 252 -83 257
rect -78 252 -77 257
rect -69 256 -68 262
rect -63 261 -33 262
rect -63 256 -62 261
rect -38 258 -33 261
rect 72 264 79 265
rect 72 259 73 264
rect 78 259 79 264
rect 72 258 79 259
rect -69 255 -62 256
rect -39 257 -32 258
rect -39 252 -38 257
rect -33 252 -32 257
rect -10 256 -3 257
rect -84 251 -77 252
rect -55 251 -48 252
rect -39 251 -32 252
rect -26 251 -20 252
rect -83 248 -78 251
rect -131 243 -78 248
rect -55 246 -54 251
rect -49 246 -48 251
rect -26 246 -25 251
rect -21 246 -20 251
rect -55 245 -20 246
rect -54 241 -20 245
rect -10 251 -9 256
rect -4 251 -3 256
rect 116 251 121 284
rect 179 261 186 262
rect 179 256 180 261
rect 185 256 186 261
rect 179 255 186 256
rect -10 250 -3 251
rect 16 250 23 251
rect -10 245 17 250
rect 22 245 23 250
rect 116 250 128 251
rect 116 245 122 250
rect 127 245 128 250
rect -10 224 -5 245
rect 16 244 23 245
rect 121 244 128 245
rect -177 218 -5 224
rect -177 198 -172 218
rect -178 197 -171 198
rect -178 192 -177 197
rect -172 192 -171 197
rect -178 191 -171 192
rect -131 194 -78 199
rect -54 197 -20 201
rect -142 190 -135 191
rect -142 185 -141 190
rect -136 185 -135 190
rect -131 189 -130 194
rect -125 189 -124 194
rect -83 191 -78 194
rect -55 196 -20 197
rect -55 191 -54 196
rect -49 191 -48 196
rect -26 191 -25 196
rect -21 191 -20 196
rect 15 192 22 193
rect 121 192 128 193
rect -131 188 -124 189
rect -84 190 -77 191
rect -55 190 -48 191
rect -39 190 -32 191
rect -26 190 -20 191
rect -10 191 16 192
rect -142 184 -135 185
rect -108 185 -101 186
rect -108 184 -107 185
rect -141 180 -107 184
rect -102 180 -101 185
rect -84 185 -83 190
rect -78 185 -77 190
rect -84 184 -77 185
rect -69 186 -62 187
rect -141 179 -101 180
rect -69 180 -68 186
rect -63 181 -62 186
rect -39 185 -38 190
rect -33 185 -32 190
rect -39 184 -32 185
rect -10 186 -9 191
rect -4 187 16 191
rect 21 187 22 192
rect -4 186 -3 187
rect 15 186 22 187
rect 117 187 122 192
rect 127 187 128 192
rect 117 186 128 187
rect -10 185 -3 186
rect -38 181 -33 184
rect -63 180 -33 181
rect -69 175 -33 180
rect -10 158 -5 185
rect -178 152 -5 158
rect 117 158 122 186
rect 117 153 160 158
rect -178 129 -173 152
rect -141 130 -101 131
rect -179 128 -172 129
rect -179 123 -178 128
rect -173 123 -172 128
rect -141 126 -107 130
rect -179 122 -172 123
rect -142 125 -135 126
rect -142 120 -141 125
rect -136 120 -135 125
rect -108 125 -107 126
rect -102 125 -101 130
rect -69 130 -33 135
rect 155 134 160 153
rect -108 124 -101 125
rect -84 125 -77 126
rect -142 119 -135 120
rect -131 121 -124 122
rect -131 116 -130 121
rect -125 116 -124 121
rect -84 120 -83 125
rect -78 120 -77 125
rect -69 124 -68 130
rect -63 129 -33 130
rect -63 124 -62 129
rect -38 126 -33 129
rect 154 133 161 134
rect 154 128 155 133
rect 160 128 161 133
rect 154 127 161 128
rect 180 126 185 255
rect 188 126 195 127
rect -69 123 -62 124
rect -39 125 -32 126
rect -39 120 -38 125
rect -33 120 -32 125
rect -10 124 -3 125
rect -84 119 -77 120
rect -55 119 -48 120
rect -39 119 -32 120
rect -26 119 -20 120
rect -83 116 -78 119
rect -131 111 -78 116
rect -55 114 -54 119
rect -49 114 -48 119
rect -26 114 -25 119
rect -21 114 -20 119
rect -55 113 -20 114
rect -54 109 -20 113
rect -10 119 -9 124
rect -4 119 -3 124
rect 72 124 79 125
rect 72 119 73 124
rect 78 119 79 124
rect 168 121 189 126
rect 194 121 195 126
rect 168 120 180 121
rect 188 120 195 121
rect -10 118 -3 119
rect 16 118 23 119
rect 72 118 79 119
rect 97 118 104 119
rect -10 113 17 118
rect 22 113 23 118
rect 73 113 98 118
rect 103 113 104 118
rect -10 92 -5 113
rect 16 112 23 113
rect 97 112 104 113
rect 168 112 173 120
rect -177 86 -5 92
rect 135 91 173 112
rect -177 66 -172 86
rect -178 65 -171 66
rect -178 60 -177 65
rect -172 60 -171 65
rect -178 59 -171 60
rect -131 62 -78 67
rect -54 65 -20 69
rect -142 58 -135 59
rect -142 53 -141 58
rect -136 53 -135 58
rect -131 57 -130 62
rect -125 57 -124 62
rect -83 59 -78 62
rect -55 64 -20 65
rect -55 59 -54 64
rect -49 59 -48 64
rect -26 59 -25 64
rect -21 59 -20 64
rect -131 56 -124 57
rect -84 58 -77 59
rect -55 58 -48 59
rect -39 58 -32 59
rect -26 58 -20 59
rect -10 59 -3 60
rect -142 52 -135 53
rect -108 53 -101 54
rect -108 52 -107 53
rect -141 48 -107 52
rect -102 48 -101 53
rect -84 53 -83 58
rect -78 53 -77 58
rect -84 52 -77 53
rect -69 54 -62 55
rect -141 47 -101 48
rect -69 48 -68 54
rect -63 49 -62 54
rect -39 53 -38 58
rect -33 53 -32 58
rect -10 54 -9 59
rect -4 57 -3 59
rect 16 57 23 58
rect 96 57 103 58
rect -4 54 17 57
rect -10 53 17 54
rect -39 52 -32 53
rect -9 52 17 53
rect 22 52 23 57
rect -38 49 -33 52
rect -63 48 -33 49
rect -69 43 -33 48
rect -9 26 -4 52
rect 16 51 23 52
rect 73 52 97 57
rect 102 52 103 57
rect -178 20 -4 26
rect -178 -3 -173 20
rect -141 -2 -101 -1
rect -179 -4 -172 -3
rect -179 -9 -178 -4
rect -173 -9 -172 -4
rect -141 -6 -107 -2
rect -179 -10 -172 -9
rect -142 -7 -135 -6
rect -142 -12 -141 -7
rect -136 -12 -135 -7
rect -108 -7 -107 -6
rect -102 -7 -101 -2
rect -69 -2 -33 3
rect 73 1 78 52
rect 96 51 103 52
rect -108 -8 -101 -7
rect -84 -7 -77 -6
rect -142 -13 -135 -12
rect -131 -11 -124 -10
rect -131 -16 -130 -11
rect -125 -16 -124 -11
rect -84 -12 -83 -7
rect -78 -12 -77 -7
rect -69 -8 -68 -2
rect -63 -3 -33 -2
rect -63 -8 -62 -3
rect -38 -6 -33 -3
rect 72 0 79 1
rect 72 -5 73 0
rect 78 -5 79 0
rect 72 -6 79 -5
rect -69 -9 -62 -8
rect -39 -7 -32 -6
rect -39 -12 -38 -7
rect -33 -12 -32 -7
rect -10 -8 -3 -7
rect -84 -13 -77 -12
rect -55 -13 -48 -12
rect -39 -13 -32 -12
rect -26 -13 -20 -12
rect -83 -16 -78 -13
rect -131 -21 -78 -16
rect -55 -18 -54 -13
rect -49 -18 -48 -13
rect -26 -18 -25 -13
rect -21 -18 -20 -13
rect -55 -19 -20 -18
rect -54 -23 -20 -19
rect -10 -13 -9 -8
rect -4 -13 -3 -8
rect -10 -14 -3 -13
rect 16 -14 23 -13
rect -10 -19 17 -14
rect 22 -19 23 -14
rect 135 -18 140 91
rect 185 53 192 54
rect 185 48 186 53
rect 191 48 192 53
rect 185 47 192 48
rect 92 -19 140 -18
rect -10 -40 -5 -19
rect 16 -20 23 -19
rect -177 -46 -5 -40
rect 61 -24 140 -19
rect 186 -15 191 47
rect 186 -21 248 -15
rect -177 -66 -172 -46
rect -178 -67 -171 -66
rect -178 -72 -177 -67
rect -172 -72 -171 -67
rect -178 -73 -171 -72
rect -131 -70 -78 -65
rect -54 -67 -20 -63
rect 61 -67 66 -24
rect 125 -66 174 -65
rect -142 -74 -135 -73
rect -142 -79 -141 -74
rect -136 -79 -135 -74
rect -131 -75 -130 -70
rect -125 -75 -124 -70
rect -83 -73 -78 -70
rect -55 -68 -20 -67
rect -55 -73 -54 -68
rect -49 -73 -48 -68
rect -26 -73 -25 -68
rect -21 -73 -20 -68
rect 60 -68 67 -67
rect -131 -76 -124 -75
rect -84 -74 -77 -73
rect -55 -74 -48 -73
rect -39 -74 -32 -73
rect -26 -74 -20 -73
rect -10 -73 -3 -72
rect -142 -80 -135 -79
rect -108 -79 -101 -78
rect -108 -80 -107 -79
rect -141 -84 -107 -80
rect -102 -84 -101 -79
rect -84 -79 -83 -74
rect -78 -79 -77 -74
rect -84 -80 -77 -79
rect -69 -78 -62 -77
rect -141 -85 -101 -84
rect -69 -84 -68 -78
rect -63 -83 -62 -78
rect -39 -79 -38 -74
rect -33 -79 -32 -74
rect -10 -78 -9 -73
rect -4 -78 -3 -73
rect 60 -73 61 -68
rect 66 -73 67 -68
rect 125 -71 126 -66
rect 131 -70 174 -66
rect 198 -67 232 -63
rect 131 -71 132 -70
rect 125 -72 132 -71
rect 169 -73 174 -70
rect 197 -68 232 -67
rect 197 -73 198 -68
rect 203 -73 204 -68
rect 226 -73 227 -68
rect 231 -73 232 -68
rect 243 -72 248 -21
rect 60 -74 67 -73
rect 110 -74 117 -73
rect -10 -79 -3 -78
rect 15 -79 22 -78
rect -39 -80 -32 -79
rect -38 -83 -33 -80
rect -63 -84 -33 -83
rect -8 -84 16 -79
rect 21 -84 22 -79
rect 110 -79 111 -74
rect 116 -79 117 -74
rect 110 -80 117 -79
rect 140 -74 147 -73
rect 140 -79 141 -74
rect 146 -79 147 -74
rect 140 -80 147 -79
rect 168 -74 175 -73
rect 197 -74 204 -73
rect 213 -74 220 -73
rect 226 -74 232 -73
rect 242 -73 249 -72
rect 168 -79 169 -74
rect 174 -79 175 -74
rect 168 -80 175 -79
rect 183 -78 190 -77
rect -69 -89 -33 -84
rect 15 -85 22 -84
rect 111 -85 146 -80
rect 183 -84 184 -78
rect 189 -83 190 -78
rect 213 -79 214 -74
rect 219 -79 220 -74
rect 242 -78 243 -73
rect 248 -78 249 -73
rect 242 -79 249 -78
rect 213 -80 220 -79
rect 214 -83 219 -80
rect 189 -84 219 -83
rect 183 -89 219 -84
<< labels >>
rlabel metal1 -13 381 -10 388 7 Q
rlabel metal1 -176 383 -172 386 1 D
rlabel metal1 -179 410 -175 414 3 clk
rlabel metal1 -179 417 -175 421 3 Vdd!
rlabel metal1 -179 358 -175 362 3 ~clk
rlabel metal1 -13 318 -10 325 7 Q
rlabel metal1 -179 292 -175 296 3 clk
rlabel metal1 -179 344 -175 348 3 ~clk
rlabel metal1 -179 351 -175 355 3 GND!
rlabel metal1 -176 320 -172 323 5 D
rlabel metal1 -13 249 -10 256 7 Q
rlabel metal1 -176 251 -172 254 1 D
rlabel metal1 -179 278 -175 282 3 clk
rlabel metal1 -179 285 -175 289 3 Vdd!
rlabel metal1 -179 226 -175 230 3 ~clk
rlabel metal1 -13 186 -10 193 7 Q
rlabel metal1 -179 160 -175 164 3 clk
rlabel metal1 -179 212 -175 216 3 ~clk
rlabel metal1 -179 219 -175 223 3 GND!
rlabel metal1 -176 188 -172 191 5 D
rlabel metal1 -176 -76 -172 -73 5 D
rlabel metal1 -179 -45 -175 -41 3 GND!
rlabel metal1 -179 -52 -175 -48 3 ~clk
rlabel metal1 -179 -111 -175 -107 3 Vdd!
rlabel metal1 -179 -104 -175 -100 3 clk
rlabel metal1 -13 -78 -10 -71 7 Q
rlabel metal1 -179 -38 -175 -34 3 ~clk
rlabel metal1 -179 21 -175 25 3 Vdd!
rlabel metal1 -179 14 -175 18 3 clk
rlabel metal1 -176 -13 -172 -10 1 D
rlabel metal1 -13 -15 -10 -8 7 Q
rlabel metal1 -176 56 -172 59 5 D
rlabel metal1 -179 87 -175 91 3 GND!
rlabel metal1 -179 80 -175 84 3 ~clk
rlabel metal1 -179 28 -175 32 3 clk
rlabel metal1 -13 54 -10 61 7 Q
rlabel metal1 -179 94 -175 98 3 ~clk
rlabel metal1 -179 153 -175 157 3 Vdd!
rlabel metal1 -179 146 -175 150 3 clk
rlabel metal1 -176 119 -172 122 1 D
rlabel metal1 -13 117 -10 124 7 Q
rlabel metal1 86 -104 89 -100 5 Vdd!
rlabel polysilicon 85 -72 87 -69 5 reset
rlabel polysilicon 67 -81 69 -78 5 D
rlabel metal1 89 -45 92 -41 4 ~clk
rlabel metal1 89 -111 92 -107 2 clk
rlabel metal1 81 -52 88 -48 5 GND!
rlabel metal3 8 -84 10 -79 1 a7
rlabel metal1 23 -111 27 -107 1 Vdd!
rlabel metal1 24 -45 27 -41 1 GND!
rlabel metal1 194 21 198 25 1 Vdd!
rlabel metal3 11 -19 13 -14 1 a6
rlabel metal1 104 21 108 25 1 Vdd!
rlabel metal1 23 21 27 25 1 Vdd!
rlabel metal3 9 52 11 57 1 a5
rlabel metal1 195 87 198 91 1 GND!
rlabel metal1 105 87 108 91 1 GND!
rlabel metal1 24 87 27 91 1 GND!
rlabel metal1 245 124 248 127 7 out
rlabel metal1 194 153 198 157 1 Vdd!
rlabel metal3 11 113 13 118 1 a4
rlabel metal1 23 153 27 157 1 Vdd!
rlabel metal1 104 153 108 157 1 Vdd!
rlabel metal3 8 187 10 192 1 a3
rlabel metal1 24 219 27 223 1 GND!
rlabel metal1 129 219 132 223 1 GND!
rlabel metal1 23 285 27 289 1 Vdd!
rlabel metal3 11 245 13 250 1 a2
rlabel metal1 104 285 108 289 1 Vdd!
rlabel metal1 173 256 176 259 7 Y
rlabel metal3 9 318 11 323 1 a1
rlabel metal1 23 417 27 421 1 Vdd!
rlabel metal3 11 377 13 382 1 a0
rlabel metal1 104 417 108 421 1 Vdd!
rlabel metal2 -3 422 0 426 4 select0
rlabel metal2 78 422 81 426 5 select1
rlabel metal2 140 422 143 426 5 select2
rlabel metal2 168 421 171 426 5 select_out
rlabel metal1 24 351 27 355 1 GND!
rlabel metal1 105 351 108 355 1 GND!
<< end >>
