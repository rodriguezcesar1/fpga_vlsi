magic
tech scmos
timestamp 1607764455
<< ntransistor >>
rect -6 23 -4 27
rect 12 23 14 27
rect 28 23 30 27
rect 44 23 46 27
rect 67 23 69 27
rect 72 23 74 27
rect 98 23 100 27
rect 119 23 121 27
rect 139 23 141 27
rect 144 23 146 27
rect 162 23 164 27
<< ptransistor >>
rect -6 41 -4 49
rect 12 41 14 49
rect 28 41 30 49
rect 44 41 46 49
rect 67 41 69 49
rect 72 41 74 49
rect 98 41 100 49
rect 119 41 121 49
rect 139 41 141 49
rect 144 41 146 49
rect 162 41 164 49
<< ndiffusion >>
rect -7 23 -6 27
rect -4 23 -3 27
rect 1 23 7 27
rect 11 23 12 27
rect 14 23 15 27
rect 27 23 28 27
rect 30 23 31 27
rect 43 23 44 27
rect 46 23 47 27
rect 62 23 67 27
rect 69 23 72 27
rect 74 23 75 27
rect 96 23 98 27
rect 100 23 101 27
rect 118 23 119 27
rect 121 23 122 27
rect 134 23 139 27
rect 141 23 144 27
rect 146 23 147 27
rect 161 23 162 27
rect 164 23 165 27
<< pdiffusion >>
rect -7 41 -6 49
rect -4 41 -3 49
rect 1 41 7 49
rect 11 41 12 49
rect 14 41 15 49
rect 27 41 28 49
rect 30 41 31 49
rect 43 41 44 49
rect 46 41 47 49
rect 62 41 67 49
rect 69 41 72 49
rect 74 41 75 49
rect 96 41 98 49
rect 100 41 101 49
rect 118 41 119 49
rect 121 41 122 49
rect 134 41 139 49
rect 141 41 144 49
rect 146 41 147 49
rect 161 41 162 49
rect 164 41 165 49
<< ndcontact >>
rect -11 23 -7 27
rect -3 23 1 27
rect 7 23 11 27
rect 15 23 19 27
rect 23 23 27 27
rect 31 23 35 27
rect 39 23 43 27
rect 47 23 51 27
rect 58 23 62 27
rect 75 23 79 27
rect 92 23 96 27
rect 101 23 105 27
rect 114 23 118 27
rect 122 23 126 27
rect 130 23 134 27
rect 147 23 151 27
rect 157 23 161 27
rect 165 23 169 27
<< pdcontact >>
rect -11 41 -7 49
rect -3 41 1 49
rect 7 41 11 49
rect 15 41 19 49
rect 23 41 27 49
rect 31 41 35 49
rect 39 41 43 49
rect 47 41 51 49
rect 58 41 62 49
rect 75 41 79 49
rect 92 41 96 49
rect 101 41 105 49
rect 114 41 118 49
rect 122 41 126 49
rect 130 41 134 49
rect 147 41 151 49
rect 157 41 161 49
rect 165 41 169 49
<< psubstratepcontact >>
rect 19 7 23 11
rect 48 7 52 11
rect 84 7 88 11
rect 123 7 127 11
<< nsubstratencontact >>
rect 16 59 20 63
rect 48 59 52 63
rect 84 59 88 63
rect 123 59 127 63
<< polysilicon >>
rect 28 56 30 59
rect 72 56 74 59
rect 98 56 100 59
rect 144 56 146 59
rect 98 52 99 56
rect -6 49 -4 52
rect 12 49 14 52
rect 28 49 30 52
rect 44 49 46 51
rect 67 49 69 51
rect 72 49 74 52
rect 98 49 100 52
rect 119 49 121 52
rect 139 49 141 51
rect 144 49 146 52
rect 162 49 164 51
rect -6 27 -4 41
rect 12 27 14 41
rect 28 39 30 41
rect 28 27 30 29
rect 44 27 46 41
rect 67 36 69 41
rect 72 39 74 41
rect 98 39 100 41
rect 63 32 69 36
rect 67 27 69 32
rect 72 27 74 29
rect 98 27 100 29
rect 119 27 121 41
rect 139 36 141 41
rect 144 39 146 41
rect 135 32 141 36
rect 139 27 141 32
rect 144 27 146 29
rect 162 27 164 41
rect -6 20 -4 23
rect 12 20 14 23
rect 28 19 30 23
rect 44 21 46 23
rect 67 21 69 23
rect 29 15 30 19
rect 72 18 74 23
rect 98 19 100 23
rect 119 21 121 23
rect 139 21 141 23
rect 28 12 30 15
rect 73 14 74 18
rect 99 15 100 19
rect 144 18 146 23
rect 162 21 164 23
rect 72 12 74 14
rect 98 11 100 15
rect 145 14 146 18
rect 144 12 146 14
<< polycontact >>
rect 28 52 32 56
rect 72 52 76 56
rect 99 52 103 56
rect 144 52 148 56
rect 40 33 44 37
rect 59 32 63 36
rect 115 33 119 37
rect 131 32 135 36
rect 158 32 162 36
rect 25 15 29 19
rect 69 14 73 18
rect 94 15 99 19
rect 141 14 145 18
<< metal1 >>
rect -11 66 32 70
rect 36 66 61 70
rect 65 66 86 70
rect 90 66 150 70
rect 154 66 169 70
rect -11 59 16 63
rect 20 59 48 63
rect 52 59 84 63
rect 88 59 123 63
rect 127 59 169 63
rect -11 49 -7 59
rect 16 49 19 59
rect 39 49 42 59
rect 58 49 61 59
rect 76 52 79 56
rect 103 52 104 56
rect 114 49 117 59
rect 130 49 133 59
rect 148 52 150 56
rect 157 49 160 59
rect 1 35 4 49
rect 23 35 26 41
rect 1 32 26 35
rect 16 27 19 32
rect 23 27 26 32
rect 32 37 35 41
rect 32 33 34 37
rect 38 33 40 37
rect 48 36 51 41
rect 76 38 79 41
rect 48 34 59 36
rect 32 27 35 33
rect 48 32 54 34
rect 48 27 51 32
rect 58 32 59 34
rect 77 34 79 38
rect 76 27 79 34
rect 92 37 95 41
rect 102 37 105 41
rect 102 33 111 37
rect 123 36 126 41
rect 148 37 151 41
rect 92 27 95 33
rect 102 27 105 33
rect 123 32 124 36
rect 128 32 131 35
rect 150 33 151 37
rect 123 27 126 32
rect 148 27 151 33
rect 166 27 169 41
rect -11 11 -8 23
rect 39 11 42 23
rect 58 11 61 23
rect 68 14 69 18
rect 93 15 94 19
rect 114 11 117 23
rect 130 11 133 23
rect 140 14 141 18
rect 157 11 160 23
rect -11 7 19 11
rect 23 7 48 11
rect 52 7 84 11
rect 88 7 123 11
rect 127 7 169 11
rect -11 0 21 4
rect 25 0 80 4
rect 84 0 105 4
rect 109 0 136 4
rect 140 0 169 4
<< m2contact >>
rect 32 66 36 70
rect 61 66 65 70
rect 86 66 90 70
rect 150 66 154 70
rect 32 52 36 56
rect 79 52 83 56
rect 104 52 108 56
rect 150 52 154 56
rect 34 33 38 37
rect 54 30 58 34
rect 73 34 77 38
rect 92 33 96 37
rect 111 33 115 37
rect 124 32 128 36
rect 146 33 150 37
rect 154 32 158 36
rect 21 15 25 19
rect 64 14 68 18
rect 86 15 93 19
rect 136 14 140 18
rect 21 0 25 4
rect 80 0 84 4
rect 105 0 109 4
rect 136 0 140 4
<< metal2 >>
rect 33 56 36 66
rect 21 4 24 15
rect 61 14 64 66
rect 80 4 83 52
rect 86 19 89 66
rect 151 56 154 66
rect 105 4 108 52
rect 136 4 140 14
<< m3contact >>
rect 38 33 43 38
rect 53 25 58 30
rect 68 33 73 38
rect 96 33 101 38
rect 111 37 116 43
rect 141 33 146 38
rect 125 27 130 32
rect 154 27 158 32
<< metal3 >>
rect 38 39 73 44
rect 110 43 146 48
rect 37 38 44 39
rect 37 33 38 38
rect 43 33 44 38
rect 37 32 44 33
rect 67 38 74 39
rect 67 33 68 38
rect 73 33 74 38
rect 67 32 74 33
rect 95 38 102 39
rect 95 33 96 38
rect 101 33 102 38
rect 110 37 111 43
rect 116 42 146 43
rect 116 37 117 42
rect 141 39 146 42
rect 110 36 117 37
rect 140 38 147 39
rect 140 33 141 38
rect 146 33 147 38
rect 95 32 102 33
rect 124 32 131 33
rect 140 32 147 33
rect 153 32 159 33
rect 52 30 59 31
rect 52 25 53 30
rect 58 29 59 30
rect 96 29 101 32
rect 58 25 101 29
rect 124 27 125 32
rect 130 27 131 32
rect 153 27 154 32
rect 158 27 159 32
rect 124 26 159 27
rect 52 24 101 25
rect 125 22 159 26
<< labels >>
rlabel metal1 166 30 169 37 7 Q
rlabel metal1 8 7 15 11 1 GND!
rlabel metal1 16 66 19 70 4 clk
rlabel metal1 16 0 19 4 2 ~clk
rlabel polysilicon -6 37 -4 40 1 D
rlabel polysilicon 12 28 14 31 1 reset
rlabel metal1 13 59 16 63 1 Vdd!
<< end >>
