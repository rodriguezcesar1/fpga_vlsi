magic
tech scmos
timestamp 1607750431
<< ntransistor >>
rect 134 487 136 491
rect 160 483 162 487
rect 165 483 167 487
rect 215 487 217 491
rect 241 483 243 487
rect 246 483 248 487
rect 188 479 190 483
rect 269 479 271 483
rect 160 453 162 457
rect 165 453 167 457
rect 241 453 243 457
rect 246 453 248 457
rect 160 383 162 387
rect 165 383 167 387
rect 239 387 241 391
rect 265 383 267 387
rect 270 383 272 387
rect 188 379 190 383
rect 293 379 295 383
rect 160 353 162 357
rect 165 353 167 357
rect 265 353 267 357
rect 270 353 272 357
rect 160 283 162 287
rect 165 283 167 287
rect 215 287 217 291
rect 241 283 243 287
rect 246 283 248 287
rect 188 279 190 283
rect 269 279 271 283
rect 160 253 162 257
rect 165 253 167 257
rect 241 253 243 257
rect 246 253 248 257
rect 160 183 162 187
rect 165 183 167 187
rect 188 179 190 183
rect 160 153 162 157
rect 165 153 167 157
<< ptransistor >>
rect 134 505 136 513
rect 160 499 162 507
rect 165 499 167 507
rect 188 505 190 513
rect 215 505 217 513
rect 241 499 243 507
rect 246 499 248 507
rect 269 505 271 513
rect 160 433 162 441
rect 165 433 167 441
rect 241 433 243 441
rect 246 433 248 441
rect 160 399 162 407
rect 165 399 167 407
rect 188 405 190 413
rect 239 405 241 413
rect 265 399 267 407
rect 270 399 272 407
rect 293 405 295 413
rect 160 333 162 341
rect 165 333 167 341
rect 265 333 267 341
rect 270 333 272 341
rect 160 299 162 307
rect 165 299 167 307
rect 188 305 190 313
rect 215 305 217 313
rect 241 299 243 307
rect 246 299 248 307
rect 269 305 271 313
rect 160 233 162 241
rect 165 233 167 241
rect 241 233 243 241
rect 246 233 248 241
rect 160 199 162 207
rect 165 199 167 207
rect 188 205 190 213
rect 160 133 162 141
rect 165 133 167 141
<< ndiffusion >>
rect 133 487 134 491
rect 136 487 137 491
rect 157 483 160 487
rect 162 483 165 487
rect 167 483 168 487
rect 214 487 215 491
rect 217 487 218 491
rect 238 483 241 487
rect 243 483 246 487
rect 248 483 249 487
rect 187 479 188 483
rect 190 479 191 483
rect 268 479 269 483
rect 271 479 272 483
rect 157 453 160 457
rect 162 453 165 457
rect 167 453 168 457
rect 238 453 241 457
rect 243 453 246 457
rect 248 453 249 457
rect 157 383 160 387
rect 162 383 165 387
rect 167 383 168 387
rect 238 387 239 391
rect 241 387 242 391
rect 262 383 265 387
rect 267 383 270 387
rect 272 383 273 387
rect 187 379 188 383
rect 190 379 191 383
rect 292 379 293 383
rect 295 379 296 383
rect 157 353 160 357
rect 162 353 165 357
rect 167 353 168 357
rect 262 353 265 357
rect 267 353 270 357
rect 272 353 273 357
rect 157 283 160 287
rect 162 283 165 287
rect 167 283 168 287
rect 214 287 215 291
rect 217 287 218 291
rect 238 283 241 287
rect 243 283 246 287
rect 248 283 249 287
rect 187 279 188 283
rect 190 279 191 283
rect 268 279 269 283
rect 271 279 272 283
rect 157 253 160 257
rect 162 253 165 257
rect 167 253 168 257
rect 238 253 241 257
rect 243 253 246 257
rect 248 253 249 257
rect 157 183 160 187
rect 162 183 165 187
rect 167 183 168 187
rect 187 179 188 183
rect 190 179 191 183
rect 157 153 160 157
rect 162 153 165 157
rect 167 153 168 157
<< pdiffusion >>
rect 133 505 134 513
rect 136 505 137 513
rect 157 499 160 507
rect 162 499 165 507
rect 167 499 168 507
rect 187 505 188 513
rect 190 505 191 513
rect 214 505 215 513
rect 217 505 218 513
rect 238 499 241 507
rect 243 499 246 507
rect 248 499 249 507
rect 268 505 269 513
rect 271 505 272 513
rect 157 433 160 441
rect 162 433 165 441
rect 167 433 168 441
rect 238 433 241 441
rect 243 433 246 441
rect 248 433 249 441
rect 157 399 160 407
rect 162 399 165 407
rect 167 399 168 407
rect 187 405 188 413
rect 190 405 191 413
rect 238 405 239 413
rect 241 405 242 413
rect 262 399 265 407
rect 267 399 270 407
rect 272 399 273 407
rect 292 405 293 413
rect 295 405 296 413
rect 157 333 160 341
rect 162 333 165 341
rect 167 333 168 341
rect 262 333 265 341
rect 267 333 270 341
rect 272 333 273 341
rect 157 299 160 307
rect 162 299 165 307
rect 167 299 168 307
rect 187 305 188 313
rect 190 305 191 313
rect 214 305 215 313
rect 217 305 218 313
rect 238 299 241 307
rect 243 299 246 307
rect 248 299 249 307
rect 268 305 269 313
rect 271 305 272 313
rect 157 233 160 241
rect 162 233 165 241
rect 167 233 168 241
rect 238 233 241 241
rect 243 233 246 241
rect 248 233 249 241
rect 157 199 160 207
rect 162 199 165 207
rect 167 199 168 207
rect 187 205 188 213
rect 190 205 191 213
rect 157 133 160 141
rect 162 133 165 141
rect 167 133 168 141
<< ndcontact >>
rect 129 487 133 491
rect 137 487 141 491
rect 153 483 157 487
rect 168 483 172 487
rect 210 487 214 491
rect 218 487 222 491
rect 234 483 238 487
rect 249 483 253 487
rect 183 479 187 483
rect 191 479 195 483
rect 264 479 268 483
rect 272 479 276 483
rect 153 453 157 457
rect 168 453 172 457
rect 234 453 238 457
rect 249 453 253 457
rect 153 383 157 387
rect 168 383 172 387
rect 234 387 238 391
rect 242 387 246 391
rect 258 383 262 387
rect 273 383 277 387
rect 183 379 187 383
rect 191 379 195 383
rect 288 379 292 383
rect 296 379 300 383
rect 153 353 157 357
rect 168 353 172 357
rect 258 353 262 357
rect 273 353 277 357
rect 153 283 157 287
rect 168 283 172 287
rect 210 287 214 291
rect 218 287 222 291
rect 234 283 238 287
rect 249 283 253 287
rect 183 279 187 283
rect 191 279 195 283
rect 264 279 268 283
rect 272 279 276 283
rect 153 253 157 257
rect 168 253 172 257
rect 234 253 238 257
rect 249 253 253 257
rect 153 183 157 187
rect 168 183 172 187
rect 183 179 187 183
rect 191 179 195 183
rect 153 153 157 157
rect 168 153 172 157
<< pdcontact >>
rect 129 505 133 513
rect 137 505 141 513
rect 153 499 157 507
rect 168 499 172 507
rect 183 505 187 513
rect 191 505 195 513
rect 210 505 214 513
rect 218 505 222 513
rect 234 499 238 507
rect 249 499 253 507
rect 264 505 268 513
rect 272 505 276 513
rect 153 433 157 441
rect 168 433 172 441
rect 234 433 238 441
rect 249 433 253 441
rect 153 399 157 407
rect 168 399 172 407
rect 183 405 187 413
rect 191 405 195 413
rect 234 405 238 413
rect 242 405 246 413
rect 258 399 262 407
rect 273 399 277 407
rect 288 405 292 413
rect 296 405 300 413
rect 153 333 157 341
rect 168 333 172 341
rect 258 333 262 341
rect 273 333 277 341
rect 153 299 157 307
rect 168 299 172 307
rect 183 305 187 313
rect 191 305 195 313
rect 210 305 214 313
rect 218 305 222 313
rect 234 299 238 307
rect 249 299 253 307
rect 264 305 268 313
rect 272 305 276 313
rect 153 233 157 241
rect 168 233 172 241
rect 234 233 238 241
rect 249 233 253 241
rect 153 199 157 207
rect 168 199 172 207
rect 183 205 187 213
rect 191 205 195 213
rect 153 133 157 141
rect 168 133 172 141
<< psubstratepcontact >>
rect 122 467 126 471
rect 146 467 150 471
rect 200 467 207 471
rect 227 467 231 471
rect 281 467 285 471
rect 122 367 126 371
rect 146 367 150 371
rect 200 367 204 371
rect 227 367 231 371
rect 251 367 255 371
rect 122 267 126 271
rect 146 267 150 271
rect 200 267 207 271
rect 227 267 231 271
rect 281 267 285 271
rect 122 167 126 171
rect 146 167 150 171
rect 200 167 204 171
<< nsubstratencontact >>
rect 122 517 126 521
rect 146 517 150 521
rect 200 517 204 521
rect 227 517 231 521
rect 281 517 285 521
rect 122 417 126 421
rect 146 417 150 421
rect 200 417 204 421
rect 227 417 231 421
rect 289 417 293 421
rect 122 317 126 321
rect 146 317 150 321
rect 200 317 204 321
rect 227 317 231 321
rect 281 317 285 321
rect 289 317 293 321
rect 122 217 126 221
rect 146 217 150 221
rect 200 217 204 221
rect 227 217 231 221
rect 146 117 150 121
<< polysilicon >>
rect 134 513 136 515
rect 160 507 162 511
rect 188 513 190 515
rect 215 513 217 515
rect 165 507 167 510
rect 134 491 136 505
rect 241 507 243 511
rect 269 513 271 515
rect 246 507 248 510
rect 160 496 162 499
rect 165 497 167 499
rect 161 492 162 496
rect 160 487 162 492
rect 165 487 167 489
rect 134 485 136 487
rect 188 483 190 505
rect 215 491 217 505
rect 241 496 243 499
rect 246 497 248 499
rect 242 492 243 496
rect 241 487 243 492
rect 246 487 248 489
rect 215 485 217 487
rect 269 483 271 505
rect 160 481 162 483
rect 165 478 167 483
rect 241 481 243 483
rect 188 477 190 479
rect 246 478 248 483
rect 269 477 271 479
rect 160 457 162 460
rect 165 457 167 460
rect 241 457 243 460
rect 246 457 248 460
rect 160 441 162 453
rect 165 451 167 453
rect 165 441 167 443
rect 241 441 243 453
rect 246 451 248 453
rect 246 441 248 443
rect 160 431 162 433
rect 165 428 167 433
rect 241 431 243 433
rect 246 428 248 433
rect 160 407 162 411
rect 188 413 190 415
rect 239 413 241 415
rect 165 407 167 410
rect 265 407 267 411
rect 293 413 295 415
rect 270 407 272 410
rect 160 396 162 399
rect 165 397 167 399
rect 161 392 162 396
rect 160 387 162 392
rect 165 387 167 389
rect 188 383 190 405
rect 239 391 241 405
rect 265 396 267 399
rect 270 397 272 399
rect 266 392 267 396
rect 265 387 267 392
rect 270 387 272 389
rect 239 385 241 387
rect 293 383 295 405
rect 160 381 162 383
rect 165 378 167 383
rect 265 381 267 383
rect 188 377 190 379
rect 270 378 272 383
rect 293 377 295 379
rect 160 357 162 360
rect 165 357 167 360
rect 265 357 267 360
rect 270 357 272 360
rect 160 341 162 353
rect 165 351 167 353
rect 165 341 167 343
rect 265 341 267 353
rect 270 351 272 353
rect 270 341 272 343
rect 160 331 162 333
rect 165 328 167 333
rect 265 331 267 333
rect 270 328 272 333
rect 160 307 162 311
rect 188 313 190 315
rect 215 313 217 315
rect 165 307 167 310
rect 241 307 243 311
rect 269 313 271 315
rect 246 307 248 310
rect 160 296 162 299
rect 165 297 167 299
rect 161 292 162 296
rect 160 287 162 292
rect 165 287 167 289
rect 188 283 190 305
rect 215 291 217 305
rect 241 296 243 299
rect 246 297 248 299
rect 242 292 243 296
rect 241 287 243 292
rect 246 287 248 289
rect 215 285 217 287
rect 269 283 271 305
rect 160 281 162 283
rect 165 278 167 283
rect 241 281 243 283
rect 188 277 190 279
rect 246 278 248 283
rect 269 277 271 279
rect 160 257 162 260
rect 165 257 167 260
rect 241 257 243 260
rect 246 257 248 260
rect 160 241 162 253
rect 165 251 167 253
rect 165 241 167 243
rect 241 241 243 253
rect 246 251 248 253
rect 246 241 248 243
rect 160 231 162 233
rect 165 228 167 233
rect 241 231 243 233
rect 246 228 248 233
rect 160 207 162 211
rect 188 213 190 215
rect 165 207 167 210
rect 160 196 162 199
rect 165 197 167 199
rect 161 192 162 196
rect 160 187 162 192
rect 165 187 167 189
rect 188 183 190 205
rect 160 181 162 183
rect 165 178 167 183
rect 188 177 190 179
rect 160 157 162 160
rect 165 157 167 160
rect 160 141 162 153
rect 165 151 167 153
rect 165 141 167 143
rect 160 131 162 133
rect 165 128 167 133
<< polycontact >>
rect 165 510 169 514
rect 130 496 134 500
rect 246 510 250 514
rect 157 492 161 496
rect 184 488 188 492
rect 211 496 215 500
rect 238 492 242 496
rect 265 488 269 492
rect 163 474 167 478
rect 244 474 248 478
rect 165 460 169 464
rect 246 460 250 464
rect 154 444 160 448
rect 235 444 241 448
rect 163 424 167 428
rect 244 424 248 428
rect 165 410 169 414
rect 270 410 274 414
rect 157 392 161 396
rect 184 388 188 392
rect 235 396 239 400
rect 262 392 266 396
rect 289 388 293 392
rect 163 374 167 378
rect 268 374 272 378
rect 165 360 169 364
rect 270 360 274 364
rect 154 344 160 348
rect 259 344 265 348
rect 163 324 167 328
rect 268 324 272 328
rect 165 310 169 314
rect 246 310 250 314
rect 157 292 161 296
rect 184 288 188 292
rect 211 296 215 300
rect 238 292 242 296
rect 265 288 269 292
rect 163 274 167 278
rect 244 274 248 278
rect 165 260 169 264
rect 246 260 250 264
rect 154 244 160 248
rect 235 244 241 248
rect 163 224 167 228
rect 244 224 248 228
rect 165 210 169 214
rect 157 192 161 196
rect 184 188 188 192
rect 163 174 167 178
rect 165 160 169 164
rect 154 144 160 148
rect 163 124 167 128
<< metal1 >>
rect 126 517 146 521
rect 150 517 200 521
rect 204 517 227 521
rect 231 517 281 521
rect 285 517 304 521
rect 129 513 132 517
rect 138 500 141 505
rect 153 507 156 517
rect 183 513 186 517
rect 210 513 213 517
rect 127 496 130 499
rect 169 496 172 499
rect 138 491 141 496
rect 146 492 157 495
rect 169 493 177 496
rect 129 471 132 487
rect 146 486 149 492
rect 169 487 172 493
rect 181 488 184 491
rect 192 491 195 505
rect 219 500 222 505
rect 234 507 237 517
rect 264 513 267 517
rect 203 496 204 499
rect 208 496 211 499
rect 250 496 253 499
rect 192 488 200 491
rect 219 491 222 496
rect 192 483 195 488
rect 200 484 204 488
rect 227 492 238 495
rect 250 493 258 496
rect 144 477 149 482
rect 153 471 156 483
rect 183 471 186 479
rect 210 471 213 487
rect 227 486 230 492
rect 250 487 253 493
rect 262 488 265 491
rect 273 491 276 505
rect 273 488 285 491
rect 273 483 276 488
rect 225 477 230 482
rect 234 471 237 483
rect 264 471 267 479
rect 126 467 146 471
rect 150 467 200 471
rect 207 467 227 471
rect 231 467 281 471
rect 153 457 156 467
rect 234 457 237 467
rect 144 444 149 449
rect 153 445 154 448
rect 169 447 172 453
rect 169 444 177 447
rect 224 444 229 449
rect 233 445 235 448
rect 250 447 253 453
rect 250 444 258 447
rect 169 441 172 444
rect 250 441 253 444
rect 153 421 156 433
rect 234 421 237 433
rect 126 417 146 421
rect 150 417 200 421
rect 204 417 227 421
rect 231 417 289 421
rect 293 417 304 421
rect 153 407 156 417
rect 183 413 186 417
rect 234 413 237 417
rect 169 396 172 399
rect 146 392 157 395
rect 169 393 177 396
rect 146 386 149 392
rect 169 387 172 393
rect 181 388 184 391
rect 192 391 195 405
rect 243 400 246 405
rect 258 407 261 417
rect 288 413 291 417
rect 227 396 228 399
rect 232 396 235 399
rect 274 396 277 399
rect 200 391 205 396
rect 243 391 246 396
rect 192 388 200 391
rect 192 383 195 388
rect 251 392 262 395
rect 274 393 282 396
rect 144 377 149 382
rect 153 371 156 383
rect 183 371 186 379
rect 234 371 237 387
rect 251 386 254 392
rect 274 387 277 393
rect 286 388 289 391
rect 297 391 300 405
rect 297 388 303 391
rect 297 383 300 388
rect 249 377 254 382
rect 258 371 261 383
rect 288 371 291 379
rect 126 367 146 371
rect 150 367 200 371
rect 204 367 227 371
rect 231 367 251 371
rect 255 367 303 371
rect 153 357 156 367
rect 258 357 261 367
rect 143 344 148 349
rect 152 345 154 348
rect 169 347 172 353
rect 169 344 177 347
rect 249 344 254 349
rect 258 345 259 348
rect 274 347 277 353
rect 274 344 282 347
rect 169 341 172 344
rect 274 341 277 344
rect 153 321 156 333
rect 258 321 261 333
rect 126 317 146 321
rect 150 317 200 321
rect 204 317 227 321
rect 231 317 281 321
rect 285 317 289 321
rect 293 317 304 321
rect 153 307 156 317
rect 183 313 186 317
rect 210 313 213 317
rect 169 296 172 299
rect 146 292 157 295
rect 169 293 177 296
rect 146 286 149 292
rect 169 287 172 293
rect 181 288 184 291
rect 192 291 195 305
rect 219 300 222 305
rect 234 307 237 317
rect 264 313 267 317
rect 203 296 204 299
rect 208 296 211 299
rect 250 296 253 299
rect 192 288 200 291
rect 219 291 222 296
rect 192 283 195 288
rect 200 284 204 288
rect 227 292 238 295
rect 250 293 258 296
rect 144 277 149 282
rect 153 271 156 283
rect 183 271 186 279
rect 210 271 213 287
rect 227 286 230 292
rect 250 287 253 293
rect 262 288 265 291
rect 273 291 276 305
rect 273 288 282 291
rect 273 283 276 288
rect 225 277 230 282
rect 234 271 237 283
rect 264 271 267 279
rect 126 267 146 271
rect 150 267 200 271
rect 207 267 227 271
rect 231 267 281 271
rect 153 257 156 267
rect 234 257 237 267
rect 144 244 149 249
rect 153 245 154 248
rect 169 247 172 253
rect 169 244 177 247
rect 224 244 229 249
rect 233 245 235 248
rect 250 247 253 253
rect 250 244 258 247
rect 169 241 172 244
rect 250 241 253 244
rect 153 221 156 233
rect 234 221 237 233
rect 126 217 146 221
rect 150 217 200 221
rect 204 217 227 221
rect 231 217 285 221
rect 153 207 156 217
rect 183 213 186 217
rect 169 196 172 199
rect 146 192 157 195
rect 169 193 177 196
rect 146 186 149 192
rect 169 187 172 193
rect 181 188 184 191
rect 192 191 195 205
rect 200 191 205 196
rect 192 188 200 191
rect 192 183 195 188
rect 144 177 149 182
rect 153 171 156 183
rect 183 171 186 179
rect 126 167 146 171
rect 150 167 200 171
rect 204 167 290 171
rect 153 157 156 167
rect 143 144 148 149
rect 152 145 154 148
rect 169 147 172 153
rect 169 144 177 147
rect 169 141 172 144
rect 153 121 156 133
rect 122 117 146 121
rect 150 117 289 121
<< m2contact >>
rect 169 510 173 514
rect 123 496 127 500
rect 138 496 142 500
rect 177 488 181 496
rect 250 510 254 514
rect 204 496 208 500
rect 219 496 223 500
rect 200 488 204 492
rect 146 482 150 486
rect 159 474 163 478
rect 258 488 262 496
rect 285 488 289 492
rect 227 482 231 486
rect 240 474 244 478
rect 169 460 173 464
rect 250 460 254 464
rect 149 445 153 449
rect 177 444 181 448
rect 229 445 233 449
rect 258 444 262 448
rect 159 424 163 428
rect 240 424 244 428
rect 169 410 173 414
rect 177 388 181 396
rect 274 410 278 414
rect 228 396 232 400
rect 243 396 247 400
rect 146 382 150 386
rect 200 387 204 391
rect 159 374 163 378
rect 282 388 286 396
rect 251 382 255 386
rect 264 374 268 378
rect 169 360 173 364
rect 274 360 278 364
rect 148 345 152 349
rect 177 344 181 348
rect 254 345 258 349
rect 282 344 286 348
rect 159 324 163 328
rect 264 324 268 328
rect 169 310 173 314
rect 177 288 181 296
rect 250 310 254 314
rect 204 296 208 300
rect 219 296 223 300
rect 200 288 204 292
rect 146 282 150 286
rect 159 274 163 278
rect 258 288 262 296
rect 282 288 286 292
rect 227 282 231 286
rect 240 274 244 278
rect 169 260 173 264
rect 250 260 254 264
rect 149 245 153 249
rect 177 244 181 248
rect 229 245 233 249
rect 258 244 262 248
rect 159 224 163 228
rect 240 224 244 228
rect 169 210 173 214
rect 177 188 181 196
rect 146 182 150 186
rect 200 187 204 191
rect 159 174 163 178
rect 169 160 173 164
rect 148 145 152 149
rect 177 144 181 148
rect 159 124 163 128
<< metal2 >>
rect 124 513 127 526
rect 124 510 169 513
rect 124 500 127 510
rect 142 497 162 500
rect 159 478 162 497
rect 159 428 162 474
rect 170 464 173 510
rect 205 513 208 526
rect 205 510 250 513
rect 205 500 208 510
rect 159 400 162 424
rect 170 414 173 460
rect 177 448 181 488
rect 165 410 169 413
rect 158 397 162 400
rect 159 378 162 397
rect 159 328 162 374
rect 170 364 173 410
rect 159 278 162 324
rect 170 314 173 360
rect 177 348 181 388
rect 165 310 169 313
rect 208 313 211 500
rect 223 497 243 500
rect 240 478 243 497
rect 240 428 243 474
rect 251 464 254 510
rect 258 448 262 488
rect 267 421 270 526
rect 229 417 270 421
rect 229 413 232 417
rect 229 410 274 413
rect 229 400 232 410
rect 247 397 267 400
rect 229 395 232 396
rect 264 378 267 397
rect 264 328 267 374
rect 275 364 278 410
rect 282 348 286 388
rect 159 228 162 274
rect 170 264 173 310
rect 205 310 250 313
rect 205 300 208 310
rect 223 297 243 300
rect 159 178 162 224
rect 170 214 173 260
rect 177 248 181 288
rect 240 278 243 297
rect 240 228 243 274
rect 251 264 254 310
rect 258 248 262 288
rect 165 210 169 213
rect 159 128 162 174
rect 170 164 173 210
rect 177 148 181 188
<< m3contact >>
rect 144 477 149 482
rect 144 444 149 449
rect 200 483 205 488
rect 144 377 149 382
rect 143 344 148 349
rect 144 277 149 282
rect 200 391 205 396
rect 225 477 230 482
rect 224 444 229 449
rect 285 483 290 488
rect 249 377 254 382
rect 249 344 254 349
rect 144 244 149 249
rect 144 177 149 182
rect 200 283 205 288
rect 225 277 230 282
rect 224 244 229 249
rect 282 292 287 297
rect 143 144 148 149
rect 200 191 205 196
<< metal3 >>
rect 199 488 206 489
rect 199 483 200 488
rect 205 483 206 488
rect 284 488 291 489
rect 284 483 285 488
rect 290 483 291 488
rect 143 482 150 483
rect 199 482 206 483
rect 224 482 231 483
rect 284 482 291 483
rect 138 477 144 482
rect 149 477 150 482
rect 200 477 225 482
rect 230 477 231 482
rect 143 476 150 477
rect 224 476 231 477
rect 281 477 290 482
rect 143 449 150 450
rect 223 449 230 450
rect 136 444 144 449
rect 149 444 150 449
rect 143 443 150 444
rect 200 444 224 449
rect 229 444 230 449
rect 200 397 205 444
rect 223 443 230 444
rect 281 421 286 477
rect 243 416 286 421
rect 199 396 206 397
rect 199 391 200 396
rect 205 391 206 396
rect 199 390 206 391
rect 243 383 248 416
rect 143 382 150 383
rect 138 377 144 382
rect 149 377 150 382
rect 243 382 255 383
rect 243 377 249 382
rect 254 377 255 382
rect 143 376 150 377
rect 248 376 255 377
rect 142 349 149 350
rect 248 349 255 350
rect 135 344 143 349
rect 148 344 149 349
rect 142 343 149 344
rect 244 344 249 349
rect 254 344 255 349
rect 244 343 255 344
rect 244 322 249 343
rect 244 317 287 322
rect 282 298 287 317
rect 281 297 288 298
rect 281 292 282 297
rect 287 292 288 297
rect 281 291 288 292
rect 199 288 206 289
rect 199 283 200 288
rect 205 283 206 288
rect 143 282 150 283
rect 199 282 206 283
rect 224 282 231 283
rect 138 277 144 282
rect 149 277 150 282
rect 200 277 225 282
rect 230 277 231 282
rect 143 276 150 277
rect 224 276 231 277
rect 143 249 150 250
rect 223 249 230 250
rect 136 244 144 249
rect 149 244 150 249
rect 143 243 150 244
rect 200 244 224 249
rect 229 244 230 249
rect 200 197 205 244
rect 223 243 230 244
rect 199 196 206 197
rect 199 191 200 196
rect 205 191 206 196
rect 199 190 206 191
rect 143 182 150 183
rect 138 177 144 182
rect 149 177 150 182
rect 143 176 150 177
rect 142 149 149 150
rect 135 144 143 149
rect 148 144 149 149
rect 142 143 149 144
<< labels >>
rlabel metal1 150 117 154 121 1 Vdd!
rlabel metal1 150 217 154 221 1 Vdd!
rlabel metal1 151 267 154 271 1 GND!
rlabel metal1 151 167 154 171 1 GND!
rlabel metal1 232 267 235 271 1 GND!
rlabel metal1 231 317 235 321 1 Vdd!
rlabel metal1 231 217 235 221 1 Vdd!
rlabel metal1 150 317 154 321 1 Vdd!
rlabel metal1 150 517 154 521 1 Vdd!
rlabel metal1 150 417 154 421 1 Vdd!
rlabel metal1 151 467 154 471 1 GND!
rlabel metal1 151 367 154 371 1 GND!
rlabel metal3 138 477 140 482 1 a0
rlabel metal3 136 444 138 449 1 a1
rlabel metal3 138 377 140 382 1 a2
rlabel metal3 135 344 137 349 1 a3
rlabel metal1 232 467 235 471 1 GND!
rlabel metal1 231 517 235 521 1 Vdd!
rlabel metal1 231 417 235 421 1 Vdd!
rlabel metal1 256 367 259 371 1 GND!
rlabel metal1 300 388 303 391 7 Y
rlabel metal3 138 277 140 282 1 a4
rlabel metal3 136 244 138 249 1 a5
rlabel metal3 138 177 140 182 1 a6
rlabel metal3 135 144 137 149 1 a7
rlabel metal2 124 522 127 526 4 select0
rlabel metal2 205 522 208 526 5 select1
rlabel metal2 267 522 270 526 5 select2
<< end >>
