magic
tech scmos
timestamp 1608340715
<< ntransistor >>
rect 497 1914 499 1918
rect 502 1914 504 1918
rect 518 1914 520 1918
rect 534 1914 536 1918
rect 539 1914 541 1918
rect 560 1914 562 1918
rect 576 1914 578 1918
rect 592 1914 594 1918
rect 597 1914 599 1918
rect 613 1914 615 1918
rect 629 1914 631 1918
rect 634 1914 636 1918
rect 650 1914 652 1918
rect 666 1914 668 1918
rect 671 1914 673 1918
rect 692 1914 694 1918
rect 708 1914 710 1918
rect 724 1914 726 1918
rect 729 1914 731 1918
rect 745 1914 747 1918
rect 761 1914 763 1918
rect 766 1914 768 1918
rect 782 1914 784 1918
rect 798 1914 800 1918
rect 803 1914 805 1918
rect 824 1914 826 1918
rect 840 1914 842 1918
rect 856 1914 858 1918
rect 861 1914 863 1918
rect 877 1914 879 1918
rect 893 1914 895 1918
rect 898 1914 900 1918
rect 914 1914 916 1918
rect 930 1914 932 1918
rect 935 1914 937 1918
rect 956 1914 958 1918
rect 972 1914 974 1918
rect 988 1914 990 1918
rect 993 1914 995 1918
rect 1009 1914 1011 1918
rect 1430 1914 1432 1918
rect 1435 1914 1437 1918
rect 1451 1914 1453 1918
rect 1467 1914 1469 1918
rect 1472 1914 1474 1918
rect 1493 1914 1495 1918
rect 1509 1914 1511 1918
rect 1525 1914 1527 1918
rect 1530 1914 1532 1918
rect 1546 1914 1548 1918
rect 1562 1914 1564 1918
rect 1567 1914 1569 1918
rect 1583 1914 1585 1918
rect 1599 1914 1601 1918
rect 1604 1914 1606 1918
rect 1625 1914 1627 1918
rect 1641 1914 1643 1918
rect 1657 1914 1659 1918
rect 1662 1914 1664 1918
rect 1678 1914 1680 1918
rect 1694 1914 1696 1918
rect 1699 1914 1701 1918
rect 1715 1914 1717 1918
rect 1731 1914 1733 1918
rect 1736 1914 1738 1918
rect 1757 1914 1759 1918
rect 1773 1914 1775 1918
rect 1789 1914 1791 1918
rect 1794 1914 1796 1918
rect 1810 1914 1812 1918
rect 1826 1914 1828 1918
rect 1831 1914 1833 1918
rect 1847 1914 1849 1918
rect 1863 1914 1865 1918
rect 1868 1914 1870 1918
rect 1889 1914 1891 1918
rect 1905 1914 1907 1918
rect 1921 1914 1923 1918
rect 1926 1914 1928 1918
rect 1942 1914 1944 1918
rect 157 1881 159 1885
rect 162 1881 164 1885
rect 178 1881 180 1885
rect 194 1881 196 1885
rect 199 1881 201 1885
rect 220 1881 222 1885
rect 236 1881 238 1885
rect 252 1881 254 1885
rect 257 1881 259 1885
rect 273 1881 275 1885
rect 1090 1881 1092 1885
rect 1095 1881 1097 1885
rect 1111 1881 1113 1885
rect 1127 1881 1129 1885
rect 1132 1881 1134 1885
rect 1153 1881 1155 1885
rect 1169 1881 1171 1885
rect 1185 1881 1187 1885
rect 1190 1881 1192 1885
rect 1206 1881 1208 1885
rect 281 1844 283 1848
rect 676 1848 678 1852
rect 702 1844 704 1848
rect 707 1844 709 1848
rect 757 1848 759 1852
rect 783 1844 785 1848
rect 788 1844 790 1848
rect 730 1840 732 1844
rect 164 1835 166 1839
rect 502 1835 504 1839
rect 518 1835 520 1839
rect 534 1835 536 1839
rect 557 1835 559 1839
rect 562 1835 564 1839
rect 588 1835 590 1839
rect 609 1835 611 1839
rect 629 1835 631 1839
rect 634 1835 636 1839
rect 652 1835 654 1839
rect 811 1840 813 1844
rect 1214 1844 1216 1848
rect 1609 1848 1611 1852
rect 1635 1844 1637 1848
rect 1640 1844 1642 1848
rect 1690 1848 1692 1852
rect 1716 1844 1718 1848
rect 1721 1844 1723 1848
rect 1663 1840 1665 1844
rect 1097 1835 1099 1839
rect 1435 1835 1437 1839
rect 1451 1835 1453 1839
rect 1467 1835 1469 1839
rect 1490 1835 1492 1839
rect 1495 1835 1497 1839
rect 1521 1835 1523 1839
rect 1542 1835 1544 1839
rect 1562 1835 1564 1839
rect 1567 1835 1569 1839
rect 1585 1835 1587 1839
rect 1744 1840 1746 1844
rect 502 1789 504 1793
rect 518 1789 520 1793
rect 534 1789 536 1793
rect 557 1789 559 1793
rect 562 1789 564 1793
rect 588 1789 590 1793
rect 609 1789 611 1793
rect 629 1789 631 1793
rect 634 1789 636 1793
rect 652 1789 654 1793
rect 148 1779 150 1783
rect 164 1779 166 1783
rect 169 1779 171 1783
rect 185 1779 187 1783
rect 201 1779 203 1783
rect 222 1779 224 1783
rect 227 1779 229 1783
rect 243 1779 245 1783
rect 259 1779 261 1783
rect 264 1779 266 1783
rect 702 1788 704 1792
rect 707 1788 709 1792
rect 783 1788 785 1792
rect 788 1788 790 1792
rect 1435 1789 1437 1793
rect 1451 1789 1453 1793
rect 1467 1789 1469 1793
rect 1490 1789 1492 1793
rect 1495 1789 1497 1793
rect 1521 1789 1523 1793
rect 1542 1789 1544 1793
rect 1562 1789 1564 1793
rect 1567 1789 1569 1793
rect 1585 1789 1587 1793
rect 1081 1779 1083 1783
rect 1097 1779 1099 1783
rect 1102 1779 1104 1783
rect 1118 1779 1120 1783
rect 1134 1779 1136 1783
rect 1155 1779 1157 1783
rect 1160 1779 1162 1783
rect 1176 1779 1178 1783
rect 1192 1779 1194 1783
rect 1197 1779 1199 1783
rect 1635 1788 1637 1792
rect 1640 1788 1642 1792
rect 1716 1788 1718 1792
rect 1721 1788 1723 1792
rect 702 1712 704 1716
rect 707 1712 709 1716
rect 781 1716 783 1720
rect 807 1712 809 1716
rect 812 1712 814 1716
rect 730 1708 732 1712
rect 502 1703 504 1707
rect 518 1703 520 1707
rect 534 1703 536 1707
rect 557 1703 559 1707
rect 562 1703 564 1707
rect 588 1703 590 1707
rect 609 1703 611 1707
rect 629 1703 631 1707
rect 634 1703 636 1707
rect 652 1703 654 1707
rect 835 1708 837 1712
rect 1635 1712 1637 1716
rect 1640 1712 1642 1716
rect 1714 1716 1716 1720
rect 1740 1712 1742 1716
rect 1745 1712 1747 1716
rect 1663 1708 1665 1712
rect 1435 1703 1437 1707
rect 1451 1703 1453 1707
rect 1467 1703 1469 1707
rect 1490 1703 1492 1707
rect 1495 1703 1497 1707
rect 1521 1703 1523 1707
rect 1542 1703 1544 1707
rect 1562 1703 1564 1707
rect 1567 1703 1569 1707
rect 1585 1703 1587 1707
rect 1768 1708 1770 1712
rect 502 1657 504 1661
rect 518 1657 520 1661
rect 534 1657 536 1661
rect 557 1657 559 1661
rect 562 1657 564 1661
rect 588 1657 590 1661
rect 609 1657 611 1661
rect 629 1657 631 1661
rect 634 1657 636 1661
rect 652 1657 654 1661
rect 702 1657 704 1661
rect 707 1657 709 1661
rect 807 1657 809 1661
rect 812 1657 814 1661
rect 1435 1657 1437 1661
rect 1451 1657 1453 1661
rect 1467 1657 1469 1661
rect 1490 1657 1492 1661
rect 1495 1657 1497 1661
rect 1521 1657 1523 1661
rect 1542 1657 1544 1661
rect 1562 1657 1564 1661
rect 1567 1657 1569 1661
rect 1585 1657 1587 1661
rect 1635 1657 1637 1661
rect 1640 1657 1642 1661
rect 1740 1657 1742 1661
rect 1745 1657 1747 1661
rect 702 1580 704 1584
rect 707 1580 709 1584
rect 757 1584 759 1588
rect 783 1580 785 1584
rect 788 1580 790 1584
rect 847 1584 849 1588
rect 873 1580 875 1584
rect 878 1580 880 1584
rect 730 1576 732 1580
rect 502 1571 504 1575
rect 518 1571 520 1575
rect 534 1571 536 1575
rect 557 1571 559 1575
rect 562 1571 564 1575
rect 588 1571 590 1575
rect 609 1571 611 1575
rect 629 1571 631 1575
rect 634 1571 636 1575
rect 652 1571 654 1575
rect 811 1576 813 1580
rect 901 1576 903 1580
rect 1635 1580 1637 1584
rect 1640 1580 1642 1584
rect 1690 1584 1692 1588
rect 1716 1580 1718 1584
rect 1721 1580 1723 1584
rect 1780 1584 1782 1588
rect 1806 1580 1808 1584
rect 1811 1580 1813 1584
rect 1663 1576 1665 1580
rect 1435 1571 1437 1575
rect 1451 1571 1453 1575
rect 1467 1571 1469 1575
rect 1490 1571 1492 1575
rect 1495 1571 1497 1575
rect 1521 1571 1523 1575
rect 1542 1571 1544 1575
rect 1562 1571 1564 1575
rect 1567 1571 1569 1575
rect 1585 1571 1587 1575
rect 1744 1576 1746 1580
rect 1834 1576 1836 1580
rect 502 1525 504 1529
rect 518 1525 520 1529
rect 534 1525 536 1529
rect 557 1525 559 1529
rect 562 1525 564 1529
rect 588 1525 590 1529
rect 609 1525 611 1529
rect 629 1525 631 1529
rect 634 1525 636 1529
rect 652 1525 654 1529
rect 702 1522 704 1526
rect 707 1522 709 1526
rect 783 1522 785 1526
rect 788 1522 790 1526
rect 873 1522 875 1526
rect 878 1522 880 1526
rect 1435 1525 1437 1529
rect 1451 1525 1453 1529
rect 1467 1525 1469 1529
rect 1490 1525 1492 1529
rect 1495 1525 1497 1529
rect 1521 1525 1523 1529
rect 1542 1525 1544 1529
rect 1562 1525 1564 1529
rect 1567 1525 1569 1529
rect 1585 1525 1587 1529
rect 1635 1522 1637 1526
rect 1640 1522 1642 1526
rect 1716 1522 1718 1526
rect 1721 1522 1723 1526
rect 1806 1522 1808 1526
rect 1811 1522 1813 1526
rect 702 1448 704 1452
rect 707 1448 709 1452
rect 730 1444 732 1448
rect 502 1439 504 1443
rect 518 1439 520 1443
rect 534 1439 536 1443
rect 557 1439 559 1443
rect 562 1439 564 1443
rect 588 1439 590 1443
rect 609 1439 611 1443
rect 629 1439 631 1443
rect 634 1439 636 1443
rect 652 1439 654 1443
rect 1635 1448 1637 1452
rect 1640 1448 1642 1452
rect 1663 1444 1665 1448
rect 1435 1439 1437 1443
rect 1451 1439 1453 1443
rect 1467 1439 1469 1443
rect 1490 1439 1492 1443
rect 1495 1439 1497 1443
rect 1521 1439 1523 1443
rect 1542 1439 1544 1443
rect 1562 1439 1564 1443
rect 1567 1439 1569 1443
rect 1585 1439 1587 1443
rect 502 1393 504 1397
rect 518 1393 520 1397
rect 534 1393 536 1397
rect 557 1393 559 1397
rect 562 1393 564 1397
rect 588 1393 590 1397
rect 609 1393 611 1397
rect 629 1393 631 1397
rect 634 1393 636 1397
rect 652 1393 654 1397
rect 736 1393 738 1397
rect 754 1393 756 1397
rect 779 1393 781 1397
rect 795 1393 797 1397
rect 818 1393 820 1397
rect 823 1393 825 1397
rect 849 1393 851 1397
rect 870 1393 872 1397
rect 890 1393 892 1397
rect 895 1393 897 1397
rect 913 1393 915 1397
rect 25 1379 27 1383
rect 30 1379 32 1383
rect 46 1379 48 1383
rect 62 1379 64 1383
rect 67 1379 69 1383
rect 88 1379 90 1383
rect 104 1379 106 1383
rect 120 1379 122 1383
rect 125 1379 127 1383
rect 141 1379 143 1383
rect 157 1379 159 1383
rect 162 1379 164 1383
rect 178 1379 180 1383
rect 194 1379 196 1383
rect 199 1379 201 1383
rect 220 1379 222 1383
rect 236 1379 238 1383
rect 252 1379 254 1383
rect 257 1379 259 1383
rect 273 1379 275 1383
rect 289 1379 291 1383
rect 294 1379 296 1383
rect 310 1379 312 1383
rect 326 1379 328 1383
rect 331 1379 333 1383
rect 352 1379 354 1383
rect 368 1379 370 1383
rect 384 1379 386 1383
rect 389 1379 391 1383
rect 405 1379 407 1383
rect 702 1386 704 1390
rect 707 1386 709 1390
rect 1435 1393 1437 1397
rect 1451 1393 1453 1397
rect 1467 1393 1469 1397
rect 1490 1393 1492 1397
rect 1495 1393 1497 1397
rect 1521 1393 1523 1397
rect 1542 1393 1544 1397
rect 1562 1393 1564 1397
rect 1567 1393 1569 1397
rect 1585 1393 1587 1397
rect 1669 1393 1671 1397
rect 1687 1393 1689 1397
rect 1712 1393 1714 1397
rect 1728 1393 1730 1397
rect 1751 1393 1753 1397
rect 1756 1393 1758 1397
rect 1782 1393 1784 1397
rect 1803 1393 1805 1397
rect 1823 1393 1825 1397
rect 1828 1393 1830 1397
rect 1846 1393 1848 1397
rect 958 1379 960 1383
rect 963 1379 965 1383
rect 979 1379 981 1383
rect 995 1379 997 1383
rect 1000 1379 1002 1383
rect 1021 1379 1023 1383
rect 1037 1379 1039 1383
rect 1053 1379 1055 1383
rect 1058 1379 1060 1383
rect 1074 1379 1076 1383
rect 1090 1379 1092 1383
rect 1095 1379 1097 1383
rect 1111 1379 1113 1383
rect 1127 1379 1129 1383
rect 1132 1379 1134 1383
rect 1153 1379 1155 1383
rect 1169 1379 1171 1383
rect 1185 1379 1187 1383
rect 1190 1379 1192 1383
rect 1206 1379 1208 1383
rect 1222 1379 1224 1383
rect 1227 1379 1229 1383
rect 1243 1379 1245 1383
rect 1259 1379 1261 1383
rect 1264 1379 1266 1383
rect 1285 1379 1287 1383
rect 1301 1379 1303 1383
rect 1317 1379 1319 1383
rect 1322 1379 1324 1383
rect 1338 1379 1340 1383
rect 1635 1386 1637 1390
rect 1640 1386 1642 1390
rect 140 1335 142 1339
rect 164 1335 166 1339
rect 925 1337 929 1339
rect 1073 1335 1075 1339
rect 1097 1335 1099 1339
rect 1858 1337 1862 1339
rect 160 1324 162 1328
rect 1093 1324 1095 1328
rect 151 1310 155 1312
rect 1084 1310 1088 1312
rect 140 1301 142 1305
rect 164 1301 166 1305
rect 1073 1301 1075 1305
rect 1097 1301 1099 1305
rect 796 1269 798 1273
rect 801 1269 803 1273
rect 817 1269 819 1273
rect 833 1269 835 1273
rect 838 1269 840 1273
rect 859 1269 861 1273
rect 875 1269 877 1273
rect 891 1269 893 1273
rect 896 1269 898 1273
rect 912 1269 914 1273
rect 1729 1269 1731 1273
rect 1734 1269 1736 1273
rect 1750 1269 1752 1273
rect 1766 1269 1768 1273
rect 1771 1269 1773 1273
rect 1792 1269 1794 1273
rect 1808 1269 1810 1273
rect 1824 1269 1826 1273
rect 1829 1269 1831 1273
rect 1845 1269 1847 1273
rect 25 1239 27 1243
rect 30 1239 32 1243
rect 46 1239 48 1243
rect 62 1239 64 1243
rect 67 1239 69 1243
rect 88 1239 90 1243
rect 104 1239 106 1243
rect 120 1239 122 1243
rect 125 1239 127 1243
rect 141 1239 143 1243
rect 157 1239 159 1243
rect 162 1239 164 1243
rect 178 1239 180 1243
rect 194 1239 196 1243
rect 199 1239 201 1243
rect 220 1239 222 1243
rect 236 1239 238 1243
rect 252 1239 254 1243
rect 257 1239 259 1243
rect 273 1239 275 1243
rect 289 1239 291 1243
rect 294 1239 296 1243
rect 310 1239 312 1243
rect 326 1239 328 1243
rect 331 1239 333 1243
rect 352 1239 354 1243
rect 368 1239 370 1243
rect 384 1239 386 1243
rect 389 1239 391 1243
rect 405 1239 407 1243
rect 958 1239 960 1243
rect 963 1239 965 1243
rect 979 1239 981 1243
rect 995 1239 997 1243
rect 1000 1239 1002 1243
rect 1021 1239 1023 1243
rect 1037 1239 1039 1243
rect 1053 1239 1055 1243
rect 1058 1239 1060 1243
rect 1074 1239 1076 1243
rect 1090 1239 1092 1243
rect 1095 1239 1097 1243
rect 1111 1239 1113 1243
rect 1127 1239 1129 1243
rect 1132 1239 1134 1243
rect 1153 1239 1155 1243
rect 1169 1239 1171 1243
rect 1185 1239 1187 1243
rect 1190 1239 1192 1243
rect 1206 1239 1208 1243
rect 1222 1239 1224 1243
rect 1227 1239 1229 1243
rect 1243 1239 1245 1243
rect 1259 1239 1261 1243
rect 1264 1239 1266 1243
rect 1285 1239 1287 1243
rect 1301 1239 1303 1243
rect 1317 1239 1319 1243
rect 1322 1239 1324 1243
rect 1338 1239 1340 1243
rect 937 1193 941 1195
rect 1870 1193 1874 1195
rect 796 1183 798 1187
rect 801 1183 803 1187
rect 817 1183 819 1187
rect 833 1183 835 1187
rect 838 1183 840 1187
rect 859 1183 861 1187
rect 875 1183 877 1187
rect 891 1183 893 1187
rect 896 1183 898 1187
rect 912 1183 914 1187
rect 1729 1183 1731 1187
rect 1734 1183 1736 1187
rect 1750 1183 1752 1187
rect 1766 1183 1768 1187
rect 1771 1183 1773 1187
rect 1792 1183 1794 1187
rect 1808 1183 1810 1187
rect 1824 1183 1826 1187
rect 1829 1183 1831 1187
rect 1845 1183 1847 1187
rect 25 1153 27 1157
rect 30 1153 32 1157
rect 46 1153 48 1157
rect 62 1153 64 1157
rect 67 1153 69 1157
rect 88 1153 90 1157
rect 104 1153 106 1157
rect 120 1153 122 1157
rect 125 1153 127 1157
rect 141 1153 143 1157
rect 157 1153 159 1157
rect 162 1153 164 1157
rect 178 1153 180 1157
rect 194 1153 196 1157
rect 199 1153 201 1157
rect 220 1153 222 1157
rect 236 1153 238 1157
rect 252 1153 254 1157
rect 257 1153 259 1157
rect 273 1153 275 1157
rect 289 1153 291 1157
rect 294 1153 296 1157
rect 310 1153 312 1157
rect 326 1153 328 1157
rect 331 1153 333 1157
rect 352 1153 354 1157
rect 368 1153 370 1157
rect 384 1153 386 1157
rect 389 1153 391 1157
rect 405 1153 407 1157
rect 958 1153 960 1157
rect 963 1153 965 1157
rect 979 1153 981 1157
rect 995 1153 997 1157
rect 1000 1153 1002 1157
rect 1021 1153 1023 1157
rect 1037 1153 1039 1157
rect 1053 1153 1055 1157
rect 1058 1153 1060 1157
rect 1074 1153 1076 1157
rect 1090 1153 1092 1157
rect 1095 1153 1097 1157
rect 1111 1153 1113 1157
rect 1127 1153 1129 1157
rect 1132 1153 1134 1157
rect 1153 1153 1155 1157
rect 1169 1153 1171 1157
rect 1185 1153 1187 1157
rect 1190 1153 1192 1157
rect 1206 1153 1208 1157
rect 1222 1153 1224 1157
rect 1227 1153 1229 1157
rect 1243 1153 1245 1157
rect 1259 1153 1261 1157
rect 1264 1153 1266 1157
rect 1285 1153 1287 1157
rect 1301 1153 1303 1157
rect 1317 1153 1319 1157
rect 1322 1153 1324 1157
rect 1338 1153 1340 1157
rect 257 1109 259 1113
rect 281 1109 283 1113
rect 1190 1109 1192 1113
rect 1214 1109 1216 1113
rect 277 1098 279 1102
rect 1210 1098 1212 1102
rect 268 1084 272 1086
rect 1201 1084 1205 1086
rect 257 1075 259 1079
rect 281 1075 283 1079
rect 1190 1075 1192 1079
rect 1214 1075 1216 1079
rect 25 1013 27 1017
rect 30 1013 32 1017
rect 46 1013 48 1017
rect 62 1013 64 1017
rect 67 1013 69 1017
rect 88 1013 90 1017
rect 104 1013 106 1017
rect 120 1013 122 1017
rect 125 1013 127 1017
rect 141 1013 143 1017
rect 157 1013 159 1017
rect 162 1013 164 1017
rect 178 1013 180 1017
rect 194 1013 196 1017
rect 199 1013 201 1017
rect 220 1013 222 1017
rect 236 1013 238 1017
rect 252 1013 254 1017
rect 257 1013 259 1017
rect 273 1013 275 1017
rect 289 1013 291 1017
rect 294 1013 296 1017
rect 310 1013 312 1017
rect 326 1013 328 1017
rect 331 1013 333 1017
rect 352 1013 354 1017
rect 368 1013 370 1017
rect 384 1013 386 1017
rect 389 1013 391 1017
rect 405 1013 407 1017
rect 958 1013 960 1017
rect 963 1013 965 1017
rect 979 1013 981 1017
rect 995 1013 997 1017
rect 1000 1013 1002 1017
rect 1021 1013 1023 1017
rect 1037 1013 1039 1017
rect 1053 1013 1055 1017
rect 1058 1013 1060 1017
rect 1074 1013 1076 1017
rect 1090 1013 1092 1017
rect 1095 1013 1097 1017
rect 1111 1013 1113 1017
rect 1127 1013 1129 1017
rect 1132 1013 1134 1017
rect 1153 1013 1155 1017
rect 1169 1013 1171 1017
rect 1185 1013 1187 1017
rect 1190 1013 1192 1017
rect 1206 1013 1208 1017
rect 1222 1013 1224 1017
rect 1227 1013 1229 1017
rect 1243 1013 1245 1017
rect 1259 1013 1261 1017
rect 1264 1013 1266 1017
rect 1285 1013 1287 1017
rect 1301 1013 1303 1017
rect 1317 1013 1319 1017
rect 1322 1013 1324 1017
rect 1338 1013 1340 1017
rect 497 934 499 938
rect 502 934 504 938
rect 518 934 520 938
rect 534 934 536 938
rect 539 934 541 938
rect 560 934 562 938
rect 576 934 578 938
rect 592 934 594 938
rect 597 934 599 938
rect 613 934 615 938
rect 629 934 631 938
rect 634 934 636 938
rect 650 934 652 938
rect 666 934 668 938
rect 671 934 673 938
rect 692 934 694 938
rect 708 934 710 938
rect 724 934 726 938
rect 729 934 731 938
rect 745 934 747 938
rect 761 934 763 938
rect 766 934 768 938
rect 782 934 784 938
rect 798 934 800 938
rect 803 934 805 938
rect 824 934 826 938
rect 840 934 842 938
rect 856 934 858 938
rect 861 934 863 938
rect 877 934 879 938
rect 893 934 895 938
rect 898 934 900 938
rect 914 934 916 938
rect 930 934 932 938
rect 935 934 937 938
rect 956 934 958 938
rect 972 934 974 938
rect 988 934 990 938
rect 993 934 995 938
rect 1009 934 1011 938
rect 1430 934 1432 938
rect 1435 934 1437 938
rect 1451 934 1453 938
rect 1467 934 1469 938
rect 1472 934 1474 938
rect 1493 934 1495 938
rect 1509 934 1511 938
rect 1525 934 1527 938
rect 1530 934 1532 938
rect 1546 934 1548 938
rect 1562 934 1564 938
rect 1567 934 1569 938
rect 1583 934 1585 938
rect 1599 934 1601 938
rect 1604 934 1606 938
rect 1625 934 1627 938
rect 1641 934 1643 938
rect 1657 934 1659 938
rect 1662 934 1664 938
rect 1678 934 1680 938
rect 1694 934 1696 938
rect 1699 934 1701 938
rect 1715 934 1717 938
rect 1731 934 1733 938
rect 1736 934 1738 938
rect 1757 934 1759 938
rect 1773 934 1775 938
rect 1789 934 1791 938
rect 1794 934 1796 938
rect 1810 934 1812 938
rect 1826 934 1828 938
rect 1831 934 1833 938
rect 1847 934 1849 938
rect 1863 934 1865 938
rect 1868 934 1870 938
rect 1889 934 1891 938
rect 1905 934 1907 938
rect 1921 934 1923 938
rect 1926 934 1928 938
rect 1942 934 1944 938
rect 157 901 159 905
rect 162 901 164 905
rect 178 901 180 905
rect 194 901 196 905
rect 199 901 201 905
rect 220 901 222 905
rect 236 901 238 905
rect 252 901 254 905
rect 257 901 259 905
rect 273 901 275 905
rect 1090 901 1092 905
rect 1095 901 1097 905
rect 1111 901 1113 905
rect 1127 901 1129 905
rect 1132 901 1134 905
rect 1153 901 1155 905
rect 1169 901 1171 905
rect 1185 901 1187 905
rect 1190 901 1192 905
rect 1206 901 1208 905
rect 281 864 283 868
rect 676 868 678 872
rect 702 864 704 868
rect 707 864 709 868
rect 757 868 759 872
rect 783 864 785 868
rect 788 864 790 868
rect 730 860 732 864
rect 164 855 166 859
rect 502 855 504 859
rect 518 855 520 859
rect 534 855 536 859
rect 557 855 559 859
rect 562 855 564 859
rect 588 855 590 859
rect 609 855 611 859
rect 629 855 631 859
rect 634 855 636 859
rect 652 855 654 859
rect 811 860 813 864
rect 1214 864 1216 868
rect 1609 868 1611 872
rect 1635 864 1637 868
rect 1640 864 1642 868
rect 1690 868 1692 872
rect 1716 864 1718 868
rect 1721 864 1723 868
rect 1663 860 1665 864
rect 1097 855 1099 859
rect 1435 855 1437 859
rect 1451 855 1453 859
rect 1467 855 1469 859
rect 1490 855 1492 859
rect 1495 855 1497 859
rect 1521 855 1523 859
rect 1542 855 1544 859
rect 1562 855 1564 859
rect 1567 855 1569 859
rect 1585 855 1587 859
rect 1744 860 1746 864
rect 502 809 504 813
rect 518 809 520 813
rect 534 809 536 813
rect 557 809 559 813
rect 562 809 564 813
rect 588 809 590 813
rect 609 809 611 813
rect 629 809 631 813
rect 634 809 636 813
rect 652 809 654 813
rect 148 799 150 803
rect 164 799 166 803
rect 169 799 171 803
rect 185 799 187 803
rect 201 799 203 803
rect 222 799 224 803
rect 227 799 229 803
rect 243 799 245 803
rect 259 799 261 803
rect 264 799 266 803
rect 702 808 704 812
rect 707 808 709 812
rect 783 808 785 812
rect 788 808 790 812
rect 1435 809 1437 813
rect 1451 809 1453 813
rect 1467 809 1469 813
rect 1490 809 1492 813
rect 1495 809 1497 813
rect 1521 809 1523 813
rect 1542 809 1544 813
rect 1562 809 1564 813
rect 1567 809 1569 813
rect 1585 809 1587 813
rect 1081 799 1083 803
rect 1097 799 1099 803
rect 1102 799 1104 803
rect 1118 799 1120 803
rect 1134 799 1136 803
rect 1155 799 1157 803
rect 1160 799 1162 803
rect 1176 799 1178 803
rect 1192 799 1194 803
rect 1197 799 1199 803
rect 1635 808 1637 812
rect 1640 808 1642 812
rect 1716 808 1718 812
rect 1721 808 1723 812
rect 702 732 704 736
rect 707 732 709 736
rect 781 736 783 740
rect 807 732 809 736
rect 812 732 814 736
rect 730 728 732 732
rect 502 723 504 727
rect 518 723 520 727
rect 534 723 536 727
rect 557 723 559 727
rect 562 723 564 727
rect 588 723 590 727
rect 609 723 611 727
rect 629 723 631 727
rect 634 723 636 727
rect 652 723 654 727
rect 835 728 837 732
rect 1635 732 1637 736
rect 1640 732 1642 736
rect 1714 736 1716 740
rect 1740 732 1742 736
rect 1745 732 1747 736
rect 1663 728 1665 732
rect 1435 723 1437 727
rect 1451 723 1453 727
rect 1467 723 1469 727
rect 1490 723 1492 727
rect 1495 723 1497 727
rect 1521 723 1523 727
rect 1542 723 1544 727
rect 1562 723 1564 727
rect 1567 723 1569 727
rect 1585 723 1587 727
rect 1768 728 1770 732
rect 502 677 504 681
rect 518 677 520 681
rect 534 677 536 681
rect 557 677 559 681
rect 562 677 564 681
rect 588 677 590 681
rect 609 677 611 681
rect 629 677 631 681
rect 634 677 636 681
rect 652 677 654 681
rect 702 677 704 681
rect 707 677 709 681
rect 807 677 809 681
rect 812 677 814 681
rect 1435 677 1437 681
rect 1451 677 1453 681
rect 1467 677 1469 681
rect 1490 677 1492 681
rect 1495 677 1497 681
rect 1521 677 1523 681
rect 1542 677 1544 681
rect 1562 677 1564 681
rect 1567 677 1569 681
rect 1585 677 1587 681
rect 1635 677 1637 681
rect 1640 677 1642 681
rect 1740 677 1742 681
rect 1745 677 1747 681
rect 702 600 704 604
rect 707 600 709 604
rect 757 604 759 608
rect 783 600 785 604
rect 788 600 790 604
rect 847 604 849 608
rect 873 600 875 604
rect 878 600 880 604
rect 730 596 732 600
rect 502 591 504 595
rect 518 591 520 595
rect 534 591 536 595
rect 557 591 559 595
rect 562 591 564 595
rect 588 591 590 595
rect 609 591 611 595
rect 629 591 631 595
rect 634 591 636 595
rect 652 591 654 595
rect 811 596 813 600
rect 901 596 903 600
rect 1635 600 1637 604
rect 1640 600 1642 604
rect 1690 604 1692 608
rect 1716 600 1718 604
rect 1721 600 1723 604
rect 1780 604 1782 608
rect 1806 600 1808 604
rect 1811 600 1813 604
rect 1663 596 1665 600
rect 1435 591 1437 595
rect 1451 591 1453 595
rect 1467 591 1469 595
rect 1490 591 1492 595
rect 1495 591 1497 595
rect 1521 591 1523 595
rect 1542 591 1544 595
rect 1562 591 1564 595
rect 1567 591 1569 595
rect 1585 591 1587 595
rect 1744 596 1746 600
rect 1834 596 1836 600
rect 502 545 504 549
rect 518 545 520 549
rect 534 545 536 549
rect 557 545 559 549
rect 562 545 564 549
rect 588 545 590 549
rect 609 545 611 549
rect 629 545 631 549
rect 634 545 636 549
rect 652 545 654 549
rect 702 542 704 546
rect 707 542 709 546
rect 783 542 785 546
rect 788 542 790 546
rect 873 542 875 546
rect 878 542 880 546
rect 1435 545 1437 549
rect 1451 545 1453 549
rect 1467 545 1469 549
rect 1490 545 1492 549
rect 1495 545 1497 549
rect 1521 545 1523 549
rect 1542 545 1544 549
rect 1562 545 1564 549
rect 1567 545 1569 549
rect 1585 545 1587 549
rect 1635 542 1637 546
rect 1640 542 1642 546
rect 1716 542 1718 546
rect 1721 542 1723 546
rect 1806 542 1808 546
rect 1811 542 1813 546
rect 702 468 704 472
rect 707 468 709 472
rect 730 464 732 468
rect 502 459 504 463
rect 518 459 520 463
rect 534 459 536 463
rect 557 459 559 463
rect 562 459 564 463
rect 588 459 590 463
rect 609 459 611 463
rect 629 459 631 463
rect 634 459 636 463
rect 652 459 654 463
rect 1635 468 1637 472
rect 1640 468 1642 472
rect 1663 464 1665 468
rect 1435 459 1437 463
rect 1451 459 1453 463
rect 1467 459 1469 463
rect 1490 459 1492 463
rect 1495 459 1497 463
rect 1521 459 1523 463
rect 1542 459 1544 463
rect 1562 459 1564 463
rect 1567 459 1569 463
rect 1585 459 1587 463
rect 502 413 504 417
rect 518 413 520 417
rect 534 413 536 417
rect 557 413 559 417
rect 562 413 564 417
rect 588 413 590 417
rect 609 413 611 417
rect 629 413 631 417
rect 634 413 636 417
rect 652 413 654 417
rect 736 413 738 417
rect 754 413 756 417
rect 779 413 781 417
rect 795 413 797 417
rect 818 413 820 417
rect 823 413 825 417
rect 849 413 851 417
rect 870 413 872 417
rect 890 413 892 417
rect 895 413 897 417
rect 913 413 915 417
rect 25 399 27 403
rect 30 399 32 403
rect 46 399 48 403
rect 62 399 64 403
rect 67 399 69 403
rect 88 399 90 403
rect 104 399 106 403
rect 120 399 122 403
rect 125 399 127 403
rect 141 399 143 403
rect 157 399 159 403
rect 162 399 164 403
rect 178 399 180 403
rect 194 399 196 403
rect 199 399 201 403
rect 220 399 222 403
rect 236 399 238 403
rect 252 399 254 403
rect 257 399 259 403
rect 273 399 275 403
rect 289 399 291 403
rect 294 399 296 403
rect 310 399 312 403
rect 326 399 328 403
rect 331 399 333 403
rect 352 399 354 403
rect 368 399 370 403
rect 384 399 386 403
rect 389 399 391 403
rect 405 399 407 403
rect 702 406 704 410
rect 707 406 709 410
rect 1435 413 1437 417
rect 1451 413 1453 417
rect 1467 413 1469 417
rect 1490 413 1492 417
rect 1495 413 1497 417
rect 1521 413 1523 417
rect 1542 413 1544 417
rect 1562 413 1564 417
rect 1567 413 1569 417
rect 1585 413 1587 417
rect 1669 413 1671 417
rect 1687 413 1689 417
rect 1712 413 1714 417
rect 1728 413 1730 417
rect 1751 413 1753 417
rect 1756 413 1758 417
rect 1782 413 1784 417
rect 1803 413 1805 417
rect 1823 413 1825 417
rect 1828 413 1830 417
rect 1846 413 1848 417
rect 958 399 960 403
rect 963 399 965 403
rect 979 399 981 403
rect 995 399 997 403
rect 1000 399 1002 403
rect 1021 399 1023 403
rect 1037 399 1039 403
rect 1053 399 1055 403
rect 1058 399 1060 403
rect 1074 399 1076 403
rect 1090 399 1092 403
rect 1095 399 1097 403
rect 1111 399 1113 403
rect 1127 399 1129 403
rect 1132 399 1134 403
rect 1153 399 1155 403
rect 1169 399 1171 403
rect 1185 399 1187 403
rect 1190 399 1192 403
rect 1206 399 1208 403
rect 1222 399 1224 403
rect 1227 399 1229 403
rect 1243 399 1245 403
rect 1259 399 1261 403
rect 1264 399 1266 403
rect 1285 399 1287 403
rect 1301 399 1303 403
rect 1317 399 1319 403
rect 1322 399 1324 403
rect 1338 399 1340 403
rect 1635 406 1637 410
rect 1640 406 1642 410
rect 140 355 142 359
rect 164 355 166 359
rect 925 357 929 359
rect 1073 355 1075 359
rect 1097 355 1099 359
rect 1858 357 1862 359
rect 160 344 162 348
rect 1093 344 1095 348
rect 151 330 155 332
rect 1084 330 1088 332
rect 140 321 142 325
rect 164 321 166 325
rect 1073 321 1075 325
rect 1097 321 1099 325
rect 796 289 798 293
rect 801 289 803 293
rect 817 289 819 293
rect 833 289 835 293
rect 838 289 840 293
rect 859 289 861 293
rect 875 289 877 293
rect 891 289 893 293
rect 896 289 898 293
rect 912 289 914 293
rect 1729 289 1731 293
rect 1734 289 1736 293
rect 1750 289 1752 293
rect 1766 289 1768 293
rect 1771 289 1773 293
rect 1792 289 1794 293
rect 1808 289 1810 293
rect 1824 289 1826 293
rect 1829 289 1831 293
rect 1845 289 1847 293
rect 25 259 27 263
rect 30 259 32 263
rect 46 259 48 263
rect 62 259 64 263
rect 67 259 69 263
rect 88 259 90 263
rect 104 259 106 263
rect 120 259 122 263
rect 125 259 127 263
rect 141 259 143 263
rect 157 259 159 263
rect 162 259 164 263
rect 178 259 180 263
rect 194 259 196 263
rect 199 259 201 263
rect 220 259 222 263
rect 236 259 238 263
rect 252 259 254 263
rect 257 259 259 263
rect 273 259 275 263
rect 289 259 291 263
rect 294 259 296 263
rect 310 259 312 263
rect 326 259 328 263
rect 331 259 333 263
rect 352 259 354 263
rect 368 259 370 263
rect 384 259 386 263
rect 389 259 391 263
rect 405 259 407 263
rect 958 259 960 263
rect 963 259 965 263
rect 979 259 981 263
rect 995 259 997 263
rect 1000 259 1002 263
rect 1021 259 1023 263
rect 1037 259 1039 263
rect 1053 259 1055 263
rect 1058 259 1060 263
rect 1074 259 1076 263
rect 1090 259 1092 263
rect 1095 259 1097 263
rect 1111 259 1113 263
rect 1127 259 1129 263
rect 1132 259 1134 263
rect 1153 259 1155 263
rect 1169 259 1171 263
rect 1185 259 1187 263
rect 1190 259 1192 263
rect 1206 259 1208 263
rect 1222 259 1224 263
rect 1227 259 1229 263
rect 1243 259 1245 263
rect 1259 259 1261 263
rect 1264 259 1266 263
rect 1285 259 1287 263
rect 1301 259 1303 263
rect 1317 259 1319 263
rect 1322 259 1324 263
rect 1338 259 1340 263
rect 937 213 941 215
rect 1870 213 1874 215
rect 796 203 798 207
rect 801 203 803 207
rect 817 203 819 207
rect 833 203 835 207
rect 838 203 840 207
rect 859 203 861 207
rect 875 203 877 207
rect 891 203 893 207
rect 896 203 898 207
rect 912 203 914 207
rect 1729 203 1731 207
rect 1734 203 1736 207
rect 1750 203 1752 207
rect 1766 203 1768 207
rect 1771 203 1773 207
rect 1792 203 1794 207
rect 1808 203 1810 207
rect 1824 203 1826 207
rect 1829 203 1831 207
rect 1845 203 1847 207
rect 25 173 27 177
rect 30 173 32 177
rect 46 173 48 177
rect 62 173 64 177
rect 67 173 69 177
rect 88 173 90 177
rect 104 173 106 177
rect 120 173 122 177
rect 125 173 127 177
rect 141 173 143 177
rect 157 173 159 177
rect 162 173 164 177
rect 178 173 180 177
rect 194 173 196 177
rect 199 173 201 177
rect 220 173 222 177
rect 236 173 238 177
rect 252 173 254 177
rect 257 173 259 177
rect 273 173 275 177
rect 289 173 291 177
rect 294 173 296 177
rect 310 173 312 177
rect 326 173 328 177
rect 331 173 333 177
rect 352 173 354 177
rect 368 173 370 177
rect 384 173 386 177
rect 389 173 391 177
rect 405 173 407 177
rect 958 173 960 177
rect 963 173 965 177
rect 979 173 981 177
rect 995 173 997 177
rect 1000 173 1002 177
rect 1021 173 1023 177
rect 1037 173 1039 177
rect 1053 173 1055 177
rect 1058 173 1060 177
rect 1074 173 1076 177
rect 1090 173 1092 177
rect 1095 173 1097 177
rect 1111 173 1113 177
rect 1127 173 1129 177
rect 1132 173 1134 177
rect 1153 173 1155 177
rect 1169 173 1171 177
rect 1185 173 1187 177
rect 1190 173 1192 177
rect 1206 173 1208 177
rect 1222 173 1224 177
rect 1227 173 1229 177
rect 1243 173 1245 177
rect 1259 173 1261 177
rect 1264 173 1266 177
rect 1285 173 1287 177
rect 1301 173 1303 177
rect 1317 173 1319 177
rect 1322 173 1324 177
rect 1338 173 1340 177
rect 257 129 259 133
rect 281 129 283 133
rect 1190 129 1192 133
rect 1214 129 1216 133
rect 277 118 279 122
rect 1210 118 1212 122
rect 268 104 272 106
rect 1201 104 1205 106
rect 257 95 259 99
rect 281 95 283 99
rect 1190 95 1192 99
rect 1214 95 1216 99
rect 25 33 27 37
rect 30 33 32 37
rect 46 33 48 37
rect 62 33 64 37
rect 67 33 69 37
rect 88 33 90 37
rect 104 33 106 37
rect 120 33 122 37
rect 125 33 127 37
rect 141 33 143 37
rect 157 33 159 37
rect 162 33 164 37
rect 178 33 180 37
rect 194 33 196 37
rect 199 33 201 37
rect 220 33 222 37
rect 236 33 238 37
rect 252 33 254 37
rect 257 33 259 37
rect 273 33 275 37
rect 289 33 291 37
rect 294 33 296 37
rect 310 33 312 37
rect 326 33 328 37
rect 331 33 333 37
rect 352 33 354 37
rect 368 33 370 37
rect 384 33 386 37
rect 389 33 391 37
rect 405 33 407 37
rect 958 33 960 37
rect 963 33 965 37
rect 979 33 981 37
rect 995 33 997 37
rect 1000 33 1002 37
rect 1021 33 1023 37
rect 1037 33 1039 37
rect 1053 33 1055 37
rect 1058 33 1060 37
rect 1074 33 1076 37
rect 1090 33 1092 37
rect 1095 33 1097 37
rect 1111 33 1113 37
rect 1127 33 1129 37
rect 1132 33 1134 37
rect 1153 33 1155 37
rect 1169 33 1171 37
rect 1185 33 1187 37
rect 1190 33 1192 37
rect 1206 33 1208 37
rect 1222 33 1224 37
rect 1227 33 1229 37
rect 1243 33 1245 37
rect 1259 33 1261 37
rect 1264 33 1266 37
rect 1285 33 1287 37
rect 1301 33 1303 37
rect 1317 33 1319 37
rect 1322 33 1324 37
rect 1338 33 1340 37
<< ptransistor >>
rect 497 1937 499 1945
rect 502 1937 504 1945
rect 518 1937 520 1945
rect 534 1937 536 1945
rect 539 1937 541 1945
rect 560 1937 562 1945
rect 576 1937 578 1945
rect 592 1937 594 1945
rect 597 1937 599 1945
rect 613 1937 615 1945
rect 629 1937 631 1945
rect 634 1937 636 1945
rect 650 1937 652 1945
rect 666 1937 668 1945
rect 671 1937 673 1945
rect 692 1937 694 1945
rect 708 1937 710 1945
rect 724 1937 726 1945
rect 729 1937 731 1945
rect 745 1937 747 1945
rect 761 1937 763 1945
rect 766 1937 768 1945
rect 782 1937 784 1945
rect 798 1937 800 1945
rect 803 1937 805 1945
rect 824 1937 826 1945
rect 840 1937 842 1945
rect 856 1937 858 1945
rect 861 1937 863 1945
rect 877 1937 879 1945
rect 893 1937 895 1945
rect 898 1937 900 1945
rect 914 1937 916 1945
rect 930 1937 932 1945
rect 935 1937 937 1945
rect 956 1937 958 1945
rect 972 1937 974 1945
rect 988 1937 990 1945
rect 993 1937 995 1945
rect 1009 1937 1011 1945
rect 1430 1937 1432 1945
rect 1435 1937 1437 1945
rect 1451 1937 1453 1945
rect 1467 1937 1469 1945
rect 1472 1937 1474 1945
rect 1493 1937 1495 1945
rect 1509 1937 1511 1945
rect 1525 1937 1527 1945
rect 1530 1937 1532 1945
rect 1546 1937 1548 1945
rect 1562 1937 1564 1945
rect 1567 1937 1569 1945
rect 1583 1937 1585 1945
rect 1599 1937 1601 1945
rect 1604 1937 1606 1945
rect 1625 1937 1627 1945
rect 1641 1937 1643 1945
rect 1657 1937 1659 1945
rect 1662 1937 1664 1945
rect 1678 1937 1680 1945
rect 1694 1937 1696 1945
rect 1699 1937 1701 1945
rect 1715 1937 1717 1945
rect 1731 1937 1733 1945
rect 1736 1937 1738 1945
rect 1757 1937 1759 1945
rect 1773 1937 1775 1945
rect 1789 1937 1791 1945
rect 1794 1937 1796 1945
rect 1810 1937 1812 1945
rect 1826 1937 1828 1945
rect 1831 1937 1833 1945
rect 1847 1937 1849 1945
rect 1863 1937 1865 1945
rect 1868 1937 1870 1945
rect 1889 1937 1891 1945
rect 1905 1937 1907 1945
rect 1921 1937 1923 1945
rect 1926 1937 1928 1945
rect 1942 1937 1944 1945
rect 157 1904 159 1912
rect 162 1904 164 1912
rect 178 1904 180 1912
rect 194 1904 196 1912
rect 199 1904 201 1912
rect 220 1904 222 1912
rect 236 1904 238 1912
rect 252 1904 254 1912
rect 257 1904 259 1912
rect 273 1904 275 1912
rect 1090 1904 1092 1912
rect 1095 1904 1097 1912
rect 1111 1904 1113 1912
rect 1127 1904 1129 1912
rect 1132 1904 1134 1912
rect 1153 1904 1155 1912
rect 1169 1904 1171 1912
rect 1185 1904 1187 1912
rect 1190 1904 1192 1912
rect 1206 1904 1208 1912
rect 676 1866 678 1874
rect 502 1853 504 1861
rect 518 1853 520 1861
rect 534 1853 536 1861
rect 557 1853 559 1861
rect 562 1853 564 1861
rect 588 1853 590 1861
rect 609 1853 611 1861
rect 629 1853 631 1861
rect 634 1853 636 1861
rect 652 1853 654 1861
rect 702 1860 704 1868
rect 707 1860 709 1868
rect 730 1866 732 1874
rect 757 1866 759 1874
rect 783 1860 785 1868
rect 788 1860 790 1868
rect 811 1866 813 1874
rect 1609 1866 1611 1874
rect 1435 1853 1437 1861
rect 1451 1853 1453 1861
rect 1467 1853 1469 1861
rect 1490 1853 1492 1861
rect 1495 1853 1497 1861
rect 1521 1853 1523 1861
rect 1542 1853 1544 1861
rect 1562 1853 1564 1861
rect 1567 1853 1569 1861
rect 1585 1853 1587 1861
rect 1635 1860 1637 1868
rect 1640 1860 1642 1868
rect 1663 1866 1665 1874
rect 1690 1866 1692 1874
rect 1716 1860 1718 1868
rect 1721 1860 1723 1868
rect 1744 1866 1746 1874
rect 148 1802 150 1810
rect 164 1802 166 1810
rect 169 1802 171 1810
rect 185 1802 187 1810
rect 201 1802 203 1810
rect 222 1802 224 1810
rect 227 1802 229 1810
rect 243 1802 245 1810
rect 259 1802 261 1810
rect 264 1802 266 1810
rect 1081 1802 1083 1810
rect 1097 1802 1099 1810
rect 1102 1802 1104 1810
rect 1118 1802 1120 1810
rect 1134 1802 1136 1810
rect 1155 1802 1157 1810
rect 1160 1802 1162 1810
rect 1176 1802 1178 1810
rect 1192 1802 1194 1810
rect 1197 1802 1199 1810
rect 502 1767 504 1775
rect 518 1767 520 1775
rect 534 1767 536 1775
rect 557 1767 559 1775
rect 562 1767 564 1775
rect 588 1767 590 1775
rect 609 1767 611 1775
rect 629 1767 631 1775
rect 634 1767 636 1775
rect 652 1767 654 1775
rect 702 1768 704 1776
rect 707 1768 709 1776
rect 783 1768 785 1776
rect 788 1768 790 1776
rect 1435 1767 1437 1775
rect 1451 1767 1453 1775
rect 1467 1767 1469 1775
rect 1490 1767 1492 1775
rect 1495 1767 1497 1775
rect 1521 1767 1523 1775
rect 1542 1767 1544 1775
rect 1562 1767 1564 1775
rect 1567 1767 1569 1775
rect 1585 1767 1587 1775
rect 1635 1768 1637 1776
rect 1640 1768 1642 1776
rect 1716 1768 1718 1776
rect 1721 1768 1723 1776
rect 502 1721 504 1729
rect 518 1721 520 1729
rect 534 1721 536 1729
rect 557 1721 559 1729
rect 562 1721 564 1729
rect 588 1721 590 1729
rect 609 1721 611 1729
rect 629 1721 631 1729
rect 634 1721 636 1729
rect 652 1721 654 1729
rect 702 1728 704 1736
rect 707 1728 709 1736
rect 730 1734 732 1742
rect 781 1734 783 1742
rect 807 1728 809 1736
rect 812 1728 814 1736
rect 835 1734 837 1742
rect 1435 1721 1437 1729
rect 1451 1721 1453 1729
rect 1467 1721 1469 1729
rect 1490 1721 1492 1729
rect 1495 1721 1497 1729
rect 1521 1721 1523 1729
rect 1542 1721 1544 1729
rect 1562 1721 1564 1729
rect 1567 1721 1569 1729
rect 1585 1721 1587 1729
rect 1635 1728 1637 1736
rect 1640 1728 1642 1736
rect 1663 1734 1665 1742
rect 1714 1734 1716 1742
rect 1740 1728 1742 1736
rect 1745 1728 1747 1736
rect 1768 1734 1770 1742
rect 502 1635 504 1643
rect 518 1635 520 1643
rect 534 1635 536 1643
rect 557 1635 559 1643
rect 562 1635 564 1643
rect 588 1635 590 1643
rect 609 1635 611 1643
rect 629 1635 631 1643
rect 634 1635 636 1643
rect 652 1635 654 1643
rect 702 1637 704 1645
rect 707 1637 709 1645
rect 807 1637 809 1645
rect 812 1637 814 1645
rect 1435 1635 1437 1643
rect 1451 1635 1453 1643
rect 1467 1635 1469 1643
rect 1490 1635 1492 1643
rect 1495 1635 1497 1643
rect 1521 1635 1523 1643
rect 1542 1635 1544 1643
rect 1562 1635 1564 1643
rect 1567 1635 1569 1643
rect 1585 1635 1587 1643
rect 1635 1637 1637 1645
rect 1640 1637 1642 1645
rect 1740 1637 1742 1645
rect 1745 1637 1747 1645
rect 502 1589 504 1597
rect 518 1589 520 1597
rect 534 1589 536 1597
rect 557 1589 559 1597
rect 562 1589 564 1597
rect 588 1589 590 1597
rect 609 1589 611 1597
rect 629 1589 631 1597
rect 634 1589 636 1597
rect 652 1589 654 1597
rect 702 1596 704 1604
rect 707 1596 709 1604
rect 730 1602 732 1610
rect 757 1602 759 1610
rect 783 1596 785 1604
rect 788 1596 790 1604
rect 811 1602 813 1610
rect 847 1602 849 1610
rect 873 1596 875 1604
rect 878 1596 880 1604
rect 901 1602 903 1610
rect 1435 1589 1437 1597
rect 1451 1589 1453 1597
rect 1467 1589 1469 1597
rect 1490 1589 1492 1597
rect 1495 1589 1497 1597
rect 1521 1589 1523 1597
rect 1542 1589 1544 1597
rect 1562 1589 1564 1597
rect 1567 1589 1569 1597
rect 1585 1589 1587 1597
rect 1635 1596 1637 1604
rect 1640 1596 1642 1604
rect 1663 1602 1665 1610
rect 1690 1602 1692 1610
rect 1716 1596 1718 1604
rect 1721 1596 1723 1604
rect 1744 1602 1746 1610
rect 1780 1602 1782 1610
rect 1806 1596 1808 1604
rect 1811 1596 1813 1604
rect 1834 1602 1836 1610
rect 502 1503 504 1511
rect 518 1503 520 1511
rect 534 1503 536 1511
rect 557 1503 559 1511
rect 562 1503 564 1511
rect 588 1503 590 1511
rect 609 1503 611 1511
rect 629 1503 631 1511
rect 634 1503 636 1511
rect 652 1503 654 1511
rect 702 1502 704 1510
rect 707 1502 709 1510
rect 783 1502 785 1510
rect 788 1502 790 1510
rect 873 1502 875 1510
rect 878 1502 880 1510
rect 1435 1503 1437 1511
rect 1451 1503 1453 1511
rect 1467 1503 1469 1511
rect 1490 1503 1492 1511
rect 1495 1503 1497 1511
rect 1521 1503 1523 1511
rect 1542 1503 1544 1511
rect 1562 1503 1564 1511
rect 1567 1503 1569 1511
rect 1585 1503 1587 1511
rect 1635 1502 1637 1510
rect 1640 1502 1642 1510
rect 1716 1502 1718 1510
rect 1721 1502 1723 1510
rect 1806 1502 1808 1510
rect 1811 1502 1813 1510
rect 502 1457 504 1465
rect 518 1457 520 1465
rect 534 1457 536 1465
rect 557 1457 559 1465
rect 562 1457 564 1465
rect 588 1457 590 1465
rect 609 1457 611 1465
rect 629 1457 631 1465
rect 634 1457 636 1465
rect 652 1457 654 1465
rect 702 1464 704 1472
rect 707 1464 709 1472
rect 730 1470 732 1478
rect 1435 1457 1437 1465
rect 1451 1457 1453 1465
rect 1467 1457 1469 1465
rect 1490 1457 1492 1465
rect 1495 1457 1497 1465
rect 1521 1457 1523 1465
rect 1542 1457 1544 1465
rect 1562 1457 1564 1465
rect 1567 1457 1569 1465
rect 1585 1457 1587 1465
rect 1635 1464 1637 1472
rect 1640 1464 1642 1472
rect 1663 1470 1665 1478
rect 25 1402 27 1410
rect 30 1402 32 1410
rect 46 1402 48 1410
rect 62 1402 64 1410
rect 67 1402 69 1410
rect 88 1402 90 1410
rect 104 1402 106 1410
rect 120 1402 122 1410
rect 125 1402 127 1410
rect 141 1402 143 1410
rect 157 1402 159 1410
rect 162 1402 164 1410
rect 178 1402 180 1410
rect 194 1402 196 1410
rect 199 1402 201 1410
rect 220 1402 222 1410
rect 236 1402 238 1410
rect 252 1402 254 1410
rect 257 1402 259 1410
rect 273 1402 275 1410
rect 289 1402 291 1410
rect 294 1402 296 1410
rect 310 1402 312 1410
rect 326 1402 328 1410
rect 331 1402 333 1410
rect 352 1402 354 1410
rect 368 1402 370 1410
rect 384 1402 386 1410
rect 389 1402 391 1410
rect 405 1402 407 1410
rect 958 1402 960 1410
rect 963 1402 965 1410
rect 979 1402 981 1410
rect 995 1402 997 1410
rect 1000 1402 1002 1410
rect 1021 1402 1023 1410
rect 1037 1402 1039 1410
rect 1053 1402 1055 1410
rect 1058 1402 1060 1410
rect 1074 1402 1076 1410
rect 1090 1402 1092 1410
rect 1095 1402 1097 1410
rect 1111 1402 1113 1410
rect 1127 1402 1129 1410
rect 1132 1402 1134 1410
rect 1153 1402 1155 1410
rect 1169 1402 1171 1410
rect 1185 1402 1187 1410
rect 1190 1402 1192 1410
rect 1206 1402 1208 1410
rect 1222 1402 1224 1410
rect 1227 1402 1229 1410
rect 1243 1402 1245 1410
rect 1259 1402 1261 1410
rect 1264 1402 1266 1410
rect 1285 1402 1287 1410
rect 1301 1402 1303 1410
rect 1317 1402 1319 1410
rect 1322 1402 1324 1410
rect 1338 1402 1340 1410
rect 502 1371 504 1379
rect 518 1371 520 1379
rect 534 1371 536 1379
rect 557 1371 559 1379
rect 562 1371 564 1379
rect 588 1371 590 1379
rect 609 1371 611 1379
rect 629 1371 631 1379
rect 634 1371 636 1379
rect 652 1371 654 1379
rect 702 1366 704 1374
rect 707 1366 709 1374
rect 736 1371 738 1379
rect 754 1371 756 1379
rect 779 1371 781 1379
rect 795 1371 797 1379
rect 818 1371 820 1379
rect 823 1371 825 1379
rect 849 1371 851 1379
rect 870 1371 872 1379
rect 890 1371 892 1379
rect 895 1371 897 1379
rect 913 1371 915 1379
rect 1435 1371 1437 1379
rect 1451 1371 1453 1379
rect 1467 1371 1469 1379
rect 1490 1371 1492 1379
rect 1495 1371 1497 1379
rect 1521 1371 1523 1379
rect 1542 1371 1544 1379
rect 1562 1371 1564 1379
rect 1567 1371 1569 1379
rect 1585 1371 1587 1379
rect 1635 1366 1637 1374
rect 1640 1366 1642 1374
rect 1669 1371 1671 1379
rect 1687 1371 1689 1379
rect 1712 1371 1714 1379
rect 1728 1371 1730 1379
rect 1751 1371 1753 1379
rect 1756 1371 1758 1379
rect 1782 1371 1784 1379
rect 1803 1371 1805 1379
rect 1823 1371 1825 1379
rect 1828 1371 1830 1379
rect 1846 1371 1848 1379
rect 796 1292 798 1300
rect 801 1292 803 1300
rect 817 1292 819 1300
rect 833 1292 835 1300
rect 838 1292 840 1300
rect 859 1292 861 1300
rect 875 1292 877 1300
rect 891 1292 893 1300
rect 896 1292 898 1300
rect 912 1292 914 1300
rect 1729 1292 1731 1300
rect 1734 1292 1736 1300
rect 1750 1292 1752 1300
rect 1766 1292 1768 1300
rect 1771 1292 1773 1300
rect 1792 1292 1794 1300
rect 1808 1292 1810 1300
rect 1824 1292 1826 1300
rect 1829 1292 1831 1300
rect 1845 1292 1847 1300
rect 25 1262 27 1270
rect 30 1262 32 1270
rect 46 1262 48 1270
rect 62 1262 64 1270
rect 67 1262 69 1270
rect 88 1262 90 1270
rect 104 1262 106 1270
rect 120 1262 122 1270
rect 125 1262 127 1270
rect 141 1262 143 1270
rect 157 1262 159 1270
rect 162 1262 164 1270
rect 178 1262 180 1270
rect 194 1262 196 1270
rect 199 1262 201 1270
rect 220 1262 222 1270
rect 236 1262 238 1270
rect 252 1262 254 1270
rect 257 1262 259 1270
rect 273 1262 275 1270
rect 289 1262 291 1270
rect 294 1262 296 1270
rect 310 1262 312 1270
rect 326 1262 328 1270
rect 331 1262 333 1270
rect 352 1262 354 1270
rect 368 1262 370 1270
rect 384 1262 386 1270
rect 389 1262 391 1270
rect 405 1262 407 1270
rect 958 1262 960 1270
rect 963 1262 965 1270
rect 979 1262 981 1270
rect 995 1262 997 1270
rect 1000 1262 1002 1270
rect 1021 1262 1023 1270
rect 1037 1262 1039 1270
rect 1053 1262 1055 1270
rect 1058 1262 1060 1270
rect 1074 1262 1076 1270
rect 1090 1262 1092 1270
rect 1095 1262 1097 1270
rect 1111 1262 1113 1270
rect 1127 1262 1129 1270
rect 1132 1262 1134 1270
rect 1153 1262 1155 1270
rect 1169 1262 1171 1270
rect 1185 1262 1187 1270
rect 1190 1262 1192 1270
rect 1206 1262 1208 1270
rect 1222 1262 1224 1270
rect 1227 1262 1229 1270
rect 1243 1262 1245 1270
rect 1259 1262 1261 1270
rect 1264 1262 1266 1270
rect 1285 1262 1287 1270
rect 1301 1262 1303 1270
rect 1317 1262 1319 1270
rect 1322 1262 1324 1270
rect 1338 1262 1340 1270
rect 796 1206 798 1214
rect 801 1206 803 1214
rect 817 1206 819 1214
rect 833 1206 835 1214
rect 838 1206 840 1214
rect 859 1206 861 1214
rect 875 1206 877 1214
rect 891 1206 893 1214
rect 896 1206 898 1214
rect 912 1206 914 1214
rect 1729 1206 1731 1214
rect 1734 1206 1736 1214
rect 1750 1206 1752 1214
rect 1766 1206 1768 1214
rect 1771 1206 1773 1214
rect 1792 1206 1794 1214
rect 1808 1206 1810 1214
rect 1824 1206 1826 1214
rect 1829 1206 1831 1214
rect 1845 1206 1847 1214
rect 25 1176 27 1184
rect 30 1176 32 1184
rect 46 1176 48 1184
rect 62 1176 64 1184
rect 67 1176 69 1184
rect 88 1176 90 1184
rect 104 1176 106 1184
rect 120 1176 122 1184
rect 125 1176 127 1184
rect 141 1176 143 1184
rect 157 1176 159 1184
rect 162 1176 164 1184
rect 178 1176 180 1184
rect 194 1176 196 1184
rect 199 1176 201 1184
rect 220 1176 222 1184
rect 236 1176 238 1184
rect 252 1176 254 1184
rect 257 1176 259 1184
rect 273 1176 275 1184
rect 289 1176 291 1184
rect 294 1176 296 1184
rect 310 1176 312 1184
rect 326 1176 328 1184
rect 331 1176 333 1184
rect 352 1176 354 1184
rect 368 1176 370 1184
rect 384 1176 386 1184
rect 389 1176 391 1184
rect 405 1176 407 1184
rect 958 1176 960 1184
rect 963 1176 965 1184
rect 979 1176 981 1184
rect 995 1176 997 1184
rect 1000 1176 1002 1184
rect 1021 1176 1023 1184
rect 1037 1176 1039 1184
rect 1053 1176 1055 1184
rect 1058 1176 1060 1184
rect 1074 1176 1076 1184
rect 1090 1176 1092 1184
rect 1095 1176 1097 1184
rect 1111 1176 1113 1184
rect 1127 1176 1129 1184
rect 1132 1176 1134 1184
rect 1153 1176 1155 1184
rect 1169 1176 1171 1184
rect 1185 1176 1187 1184
rect 1190 1176 1192 1184
rect 1206 1176 1208 1184
rect 1222 1176 1224 1184
rect 1227 1176 1229 1184
rect 1243 1176 1245 1184
rect 1259 1176 1261 1184
rect 1264 1176 1266 1184
rect 1285 1176 1287 1184
rect 1301 1176 1303 1184
rect 1317 1176 1319 1184
rect 1322 1176 1324 1184
rect 1338 1176 1340 1184
rect 25 1036 27 1044
rect 30 1036 32 1044
rect 46 1036 48 1044
rect 62 1036 64 1044
rect 67 1036 69 1044
rect 88 1036 90 1044
rect 104 1036 106 1044
rect 120 1036 122 1044
rect 125 1036 127 1044
rect 141 1036 143 1044
rect 157 1036 159 1044
rect 162 1036 164 1044
rect 178 1036 180 1044
rect 194 1036 196 1044
rect 199 1036 201 1044
rect 220 1036 222 1044
rect 236 1036 238 1044
rect 252 1036 254 1044
rect 257 1036 259 1044
rect 273 1036 275 1044
rect 289 1036 291 1044
rect 294 1036 296 1044
rect 310 1036 312 1044
rect 326 1036 328 1044
rect 331 1036 333 1044
rect 352 1036 354 1044
rect 368 1036 370 1044
rect 384 1036 386 1044
rect 389 1036 391 1044
rect 405 1036 407 1044
rect 958 1036 960 1044
rect 963 1036 965 1044
rect 979 1036 981 1044
rect 995 1036 997 1044
rect 1000 1036 1002 1044
rect 1021 1036 1023 1044
rect 1037 1036 1039 1044
rect 1053 1036 1055 1044
rect 1058 1036 1060 1044
rect 1074 1036 1076 1044
rect 1090 1036 1092 1044
rect 1095 1036 1097 1044
rect 1111 1036 1113 1044
rect 1127 1036 1129 1044
rect 1132 1036 1134 1044
rect 1153 1036 1155 1044
rect 1169 1036 1171 1044
rect 1185 1036 1187 1044
rect 1190 1036 1192 1044
rect 1206 1036 1208 1044
rect 1222 1036 1224 1044
rect 1227 1036 1229 1044
rect 1243 1036 1245 1044
rect 1259 1036 1261 1044
rect 1264 1036 1266 1044
rect 1285 1036 1287 1044
rect 1301 1036 1303 1044
rect 1317 1036 1319 1044
rect 1322 1036 1324 1044
rect 1338 1036 1340 1044
rect 497 957 499 965
rect 502 957 504 965
rect 518 957 520 965
rect 534 957 536 965
rect 539 957 541 965
rect 560 957 562 965
rect 576 957 578 965
rect 592 957 594 965
rect 597 957 599 965
rect 613 957 615 965
rect 629 957 631 965
rect 634 957 636 965
rect 650 957 652 965
rect 666 957 668 965
rect 671 957 673 965
rect 692 957 694 965
rect 708 957 710 965
rect 724 957 726 965
rect 729 957 731 965
rect 745 957 747 965
rect 761 957 763 965
rect 766 957 768 965
rect 782 957 784 965
rect 798 957 800 965
rect 803 957 805 965
rect 824 957 826 965
rect 840 957 842 965
rect 856 957 858 965
rect 861 957 863 965
rect 877 957 879 965
rect 893 957 895 965
rect 898 957 900 965
rect 914 957 916 965
rect 930 957 932 965
rect 935 957 937 965
rect 956 957 958 965
rect 972 957 974 965
rect 988 957 990 965
rect 993 957 995 965
rect 1009 957 1011 965
rect 1430 957 1432 965
rect 1435 957 1437 965
rect 1451 957 1453 965
rect 1467 957 1469 965
rect 1472 957 1474 965
rect 1493 957 1495 965
rect 1509 957 1511 965
rect 1525 957 1527 965
rect 1530 957 1532 965
rect 1546 957 1548 965
rect 1562 957 1564 965
rect 1567 957 1569 965
rect 1583 957 1585 965
rect 1599 957 1601 965
rect 1604 957 1606 965
rect 1625 957 1627 965
rect 1641 957 1643 965
rect 1657 957 1659 965
rect 1662 957 1664 965
rect 1678 957 1680 965
rect 1694 957 1696 965
rect 1699 957 1701 965
rect 1715 957 1717 965
rect 1731 957 1733 965
rect 1736 957 1738 965
rect 1757 957 1759 965
rect 1773 957 1775 965
rect 1789 957 1791 965
rect 1794 957 1796 965
rect 1810 957 1812 965
rect 1826 957 1828 965
rect 1831 957 1833 965
rect 1847 957 1849 965
rect 1863 957 1865 965
rect 1868 957 1870 965
rect 1889 957 1891 965
rect 1905 957 1907 965
rect 1921 957 1923 965
rect 1926 957 1928 965
rect 1942 957 1944 965
rect 157 924 159 932
rect 162 924 164 932
rect 178 924 180 932
rect 194 924 196 932
rect 199 924 201 932
rect 220 924 222 932
rect 236 924 238 932
rect 252 924 254 932
rect 257 924 259 932
rect 273 924 275 932
rect 1090 924 1092 932
rect 1095 924 1097 932
rect 1111 924 1113 932
rect 1127 924 1129 932
rect 1132 924 1134 932
rect 1153 924 1155 932
rect 1169 924 1171 932
rect 1185 924 1187 932
rect 1190 924 1192 932
rect 1206 924 1208 932
rect 676 886 678 894
rect 502 873 504 881
rect 518 873 520 881
rect 534 873 536 881
rect 557 873 559 881
rect 562 873 564 881
rect 588 873 590 881
rect 609 873 611 881
rect 629 873 631 881
rect 634 873 636 881
rect 652 873 654 881
rect 702 880 704 888
rect 707 880 709 888
rect 730 886 732 894
rect 757 886 759 894
rect 783 880 785 888
rect 788 880 790 888
rect 811 886 813 894
rect 1609 886 1611 894
rect 1435 873 1437 881
rect 1451 873 1453 881
rect 1467 873 1469 881
rect 1490 873 1492 881
rect 1495 873 1497 881
rect 1521 873 1523 881
rect 1542 873 1544 881
rect 1562 873 1564 881
rect 1567 873 1569 881
rect 1585 873 1587 881
rect 1635 880 1637 888
rect 1640 880 1642 888
rect 1663 886 1665 894
rect 1690 886 1692 894
rect 1716 880 1718 888
rect 1721 880 1723 888
rect 1744 886 1746 894
rect 148 822 150 830
rect 164 822 166 830
rect 169 822 171 830
rect 185 822 187 830
rect 201 822 203 830
rect 222 822 224 830
rect 227 822 229 830
rect 243 822 245 830
rect 259 822 261 830
rect 264 822 266 830
rect 1081 822 1083 830
rect 1097 822 1099 830
rect 1102 822 1104 830
rect 1118 822 1120 830
rect 1134 822 1136 830
rect 1155 822 1157 830
rect 1160 822 1162 830
rect 1176 822 1178 830
rect 1192 822 1194 830
rect 1197 822 1199 830
rect 502 787 504 795
rect 518 787 520 795
rect 534 787 536 795
rect 557 787 559 795
rect 562 787 564 795
rect 588 787 590 795
rect 609 787 611 795
rect 629 787 631 795
rect 634 787 636 795
rect 652 787 654 795
rect 702 788 704 796
rect 707 788 709 796
rect 783 788 785 796
rect 788 788 790 796
rect 1435 787 1437 795
rect 1451 787 1453 795
rect 1467 787 1469 795
rect 1490 787 1492 795
rect 1495 787 1497 795
rect 1521 787 1523 795
rect 1542 787 1544 795
rect 1562 787 1564 795
rect 1567 787 1569 795
rect 1585 787 1587 795
rect 1635 788 1637 796
rect 1640 788 1642 796
rect 1716 788 1718 796
rect 1721 788 1723 796
rect 502 741 504 749
rect 518 741 520 749
rect 534 741 536 749
rect 557 741 559 749
rect 562 741 564 749
rect 588 741 590 749
rect 609 741 611 749
rect 629 741 631 749
rect 634 741 636 749
rect 652 741 654 749
rect 702 748 704 756
rect 707 748 709 756
rect 730 754 732 762
rect 781 754 783 762
rect 807 748 809 756
rect 812 748 814 756
rect 835 754 837 762
rect 1435 741 1437 749
rect 1451 741 1453 749
rect 1467 741 1469 749
rect 1490 741 1492 749
rect 1495 741 1497 749
rect 1521 741 1523 749
rect 1542 741 1544 749
rect 1562 741 1564 749
rect 1567 741 1569 749
rect 1585 741 1587 749
rect 1635 748 1637 756
rect 1640 748 1642 756
rect 1663 754 1665 762
rect 1714 754 1716 762
rect 1740 748 1742 756
rect 1745 748 1747 756
rect 1768 754 1770 762
rect 502 655 504 663
rect 518 655 520 663
rect 534 655 536 663
rect 557 655 559 663
rect 562 655 564 663
rect 588 655 590 663
rect 609 655 611 663
rect 629 655 631 663
rect 634 655 636 663
rect 652 655 654 663
rect 702 657 704 665
rect 707 657 709 665
rect 807 657 809 665
rect 812 657 814 665
rect 1435 655 1437 663
rect 1451 655 1453 663
rect 1467 655 1469 663
rect 1490 655 1492 663
rect 1495 655 1497 663
rect 1521 655 1523 663
rect 1542 655 1544 663
rect 1562 655 1564 663
rect 1567 655 1569 663
rect 1585 655 1587 663
rect 1635 657 1637 665
rect 1640 657 1642 665
rect 1740 657 1742 665
rect 1745 657 1747 665
rect 502 609 504 617
rect 518 609 520 617
rect 534 609 536 617
rect 557 609 559 617
rect 562 609 564 617
rect 588 609 590 617
rect 609 609 611 617
rect 629 609 631 617
rect 634 609 636 617
rect 652 609 654 617
rect 702 616 704 624
rect 707 616 709 624
rect 730 622 732 630
rect 757 622 759 630
rect 783 616 785 624
rect 788 616 790 624
rect 811 622 813 630
rect 847 622 849 630
rect 873 616 875 624
rect 878 616 880 624
rect 901 622 903 630
rect 1435 609 1437 617
rect 1451 609 1453 617
rect 1467 609 1469 617
rect 1490 609 1492 617
rect 1495 609 1497 617
rect 1521 609 1523 617
rect 1542 609 1544 617
rect 1562 609 1564 617
rect 1567 609 1569 617
rect 1585 609 1587 617
rect 1635 616 1637 624
rect 1640 616 1642 624
rect 1663 622 1665 630
rect 1690 622 1692 630
rect 1716 616 1718 624
rect 1721 616 1723 624
rect 1744 622 1746 630
rect 1780 622 1782 630
rect 1806 616 1808 624
rect 1811 616 1813 624
rect 1834 622 1836 630
rect 502 523 504 531
rect 518 523 520 531
rect 534 523 536 531
rect 557 523 559 531
rect 562 523 564 531
rect 588 523 590 531
rect 609 523 611 531
rect 629 523 631 531
rect 634 523 636 531
rect 652 523 654 531
rect 702 522 704 530
rect 707 522 709 530
rect 783 522 785 530
rect 788 522 790 530
rect 873 522 875 530
rect 878 522 880 530
rect 1435 523 1437 531
rect 1451 523 1453 531
rect 1467 523 1469 531
rect 1490 523 1492 531
rect 1495 523 1497 531
rect 1521 523 1523 531
rect 1542 523 1544 531
rect 1562 523 1564 531
rect 1567 523 1569 531
rect 1585 523 1587 531
rect 1635 522 1637 530
rect 1640 522 1642 530
rect 1716 522 1718 530
rect 1721 522 1723 530
rect 1806 522 1808 530
rect 1811 522 1813 530
rect 502 477 504 485
rect 518 477 520 485
rect 534 477 536 485
rect 557 477 559 485
rect 562 477 564 485
rect 588 477 590 485
rect 609 477 611 485
rect 629 477 631 485
rect 634 477 636 485
rect 652 477 654 485
rect 702 484 704 492
rect 707 484 709 492
rect 730 490 732 498
rect 1435 477 1437 485
rect 1451 477 1453 485
rect 1467 477 1469 485
rect 1490 477 1492 485
rect 1495 477 1497 485
rect 1521 477 1523 485
rect 1542 477 1544 485
rect 1562 477 1564 485
rect 1567 477 1569 485
rect 1585 477 1587 485
rect 1635 484 1637 492
rect 1640 484 1642 492
rect 1663 490 1665 498
rect 25 422 27 430
rect 30 422 32 430
rect 46 422 48 430
rect 62 422 64 430
rect 67 422 69 430
rect 88 422 90 430
rect 104 422 106 430
rect 120 422 122 430
rect 125 422 127 430
rect 141 422 143 430
rect 157 422 159 430
rect 162 422 164 430
rect 178 422 180 430
rect 194 422 196 430
rect 199 422 201 430
rect 220 422 222 430
rect 236 422 238 430
rect 252 422 254 430
rect 257 422 259 430
rect 273 422 275 430
rect 289 422 291 430
rect 294 422 296 430
rect 310 422 312 430
rect 326 422 328 430
rect 331 422 333 430
rect 352 422 354 430
rect 368 422 370 430
rect 384 422 386 430
rect 389 422 391 430
rect 405 422 407 430
rect 958 422 960 430
rect 963 422 965 430
rect 979 422 981 430
rect 995 422 997 430
rect 1000 422 1002 430
rect 1021 422 1023 430
rect 1037 422 1039 430
rect 1053 422 1055 430
rect 1058 422 1060 430
rect 1074 422 1076 430
rect 1090 422 1092 430
rect 1095 422 1097 430
rect 1111 422 1113 430
rect 1127 422 1129 430
rect 1132 422 1134 430
rect 1153 422 1155 430
rect 1169 422 1171 430
rect 1185 422 1187 430
rect 1190 422 1192 430
rect 1206 422 1208 430
rect 1222 422 1224 430
rect 1227 422 1229 430
rect 1243 422 1245 430
rect 1259 422 1261 430
rect 1264 422 1266 430
rect 1285 422 1287 430
rect 1301 422 1303 430
rect 1317 422 1319 430
rect 1322 422 1324 430
rect 1338 422 1340 430
rect 502 391 504 399
rect 518 391 520 399
rect 534 391 536 399
rect 557 391 559 399
rect 562 391 564 399
rect 588 391 590 399
rect 609 391 611 399
rect 629 391 631 399
rect 634 391 636 399
rect 652 391 654 399
rect 702 386 704 394
rect 707 386 709 394
rect 736 391 738 399
rect 754 391 756 399
rect 779 391 781 399
rect 795 391 797 399
rect 818 391 820 399
rect 823 391 825 399
rect 849 391 851 399
rect 870 391 872 399
rect 890 391 892 399
rect 895 391 897 399
rect 913 391 915 399
rect 1435 391 1437 399
rect 1451 391 1453 399
rect 1467 391 1469 399
rect 1490 391 1492 399
rect 1495 391 1497 399
rect 1521 391 1523 399
rect 1542 391 1544 399
rect 1562 391 1564 399
rect 1567 391 1569 399
rect 1585 391 1587 399
rect 1635 386 1637 394
rect 1640 386 1642 394
rect 1669 391 1671 399
rect 1687 391 1689 399
rect 1712 391 1714 399
rect 1728 391 1730 399
rect 1751 391 1753 399
rect 1756 391 1758 399
rect 1782 391 1784 399
rect 1803 391 1805 399
rect 1823 391 1825 399
rect 1828 391 1830 399
rect 1846 391 1848 399
rect 796 312 798 320
rect 801 312 803 320
rect 817 312 819 320
rect 833 312 835 320
rect 838 312 840 320
rect 859 312 861 320
rect 875 312 877 320
rect 891 312 893 320
rect 896 312 898 320
rect 912 312 914 320
rect 1729 312 1731 320
rect 1734 312 1736 320
rect 1750 312 1752 320
rect 1766 312 1768 320
rect 1771 312 1773 320
rect 1792 312 1794 320
rect 1808 312 1810 320
rect 1824 312 1826 320
rect 1829 312 1831 320
rect 1845 312 1847 320
rect 25 282 27 290
rect 30 282 32 290
rect 46 282 48 290
rect 62 282 64 290
rect 67 282 69 290
rect 88 282 90 290
rect 104 282 106 290
rect 120 282 122 290
rect 125 282 127 290
rect 141 282 143 290
rect 157 282 159 290
rect 162 282 164 290
rect 178 282 180 290
rect 194 282 196 290
rect 199 282 201 290
rect 220 282 222 290
rect 236 282 238 290
rect 252 282 254 290
rect 257 282 259 290
rect 273 282 275 290
rect 289 282 291 290
rect 294 282 296 290
rect 310 282 312 290
rect 326 282 328 290
rect 331 282 333 290
rect 352 282 354 290
rect 368 282 370 290
rect 384 282 386 290
rect 389 282 391 290
rect 405 282 407 290
rect 958 282 960 290
rect 963 282 965 290
rect 979 282 981 290
rect 995 282 997 290
rect 1000 282 1002 290
rect 1021 282 1023 290
rect 1037 282 1039 290
rect 1053 282 1055 290
rect 1058 282 1060 290
rect 1074 282 1076 290
rect 1090 282 1092 290
rect 1095 282 1097 290
rect 1111 282 1113 290
rect 1127 282 1129 290
rect 1132 282 1134 290
rect 1153 282 1155 290
rect 1169 282 1171 290
rect 1185 282 1187 290
rect 1190 282 1192 290
rect 1206 282 1208 290
rect 1222 282 1224 290
rect 1227 282 1229 290
rect 1243 282 1245 290
rect 1259 282 1261 290
rect 1264 282 1266 290
rect 1285 282 1287 290
rect 1301 282 1303 290
rect 1317 282 1319 290
rect 1322 282 1324 290
rect 1338 282 1340 290
rect 796 226 798 234
rect 801 226 803 234
rect 817 226 819 234
rect 833 226 835 234
rect 838 226 840 234
rect 859 226 861 234
rect 875 226 877 234
rect 891 226 893 234
rect 896 226 898 234
rect 912 226 914 234
rect 1729 226 1731 234
rect 1734 226 1736 234
rect 1750 226 1752 234
rect 1766 226 1768 234
rect 1771 226 1773 234
rect 1792 226 1794 234
rect 1808 226 1810 234
rect 1824 226 1826 234
rect 1829 226 1831 234
rect 1845 226 1847 234
rect 25 196 27 204
rect 30 196 32 204
rect 46 196 48 204
rect 62 196 64 204
rect 67 196 69 204
rect 88 196 90 204
rect 104 196 106 204
rect 120 196 122 204
rect 125 196 127 204
rect 141 196 143 204
rect 157 196 159 204
rect 162 196 164 204
rect 178 196 180 204
rect 194 196 196 204
rect 199 196 201 204
rect 220 196 222 204
rect 236 196 238 204
rect 252 196 254 204
rect 257 196 259 204
rect 273 196 275 204
rect 289 196 291 204
rect 294 196 296 204
rect 310 196 312 204
rect 326 196 328 204
rect 331 196 333 204
rect 352 196 354 204
rect 368 196 370 204
rect 384 196 386 204
rect 389 196 391 204
rect 405 196 407 204
rect 958 196 960 204
rect 963 196 965 204
rect 979 196 981 204
rect 995 196 997 204
rect 1000 196 1002 204
rect 1021 196 1023 204
rect 1037 196 1039 204
rect 1053 196 1055 204
rect 1058 196 1060 204
rect 1074 196 1076 204
rect 1090 196 1092 204
rect 1095 196 1097 204
rect 1111 196 1113 204
rect 1127 196 1129 204
rect 1132 196 1134 204
rect 1153 196 1155 204
rect 1169 196 1171 204
rect 1185 196 1187 204
rect 1190 196 1192 204
rect 1206 196 1208 204
rect 1222 196 1224 204
rect 1227 196 1229 204
rect 1243 196 1245 204
rect 1259 196 1261 204
rect 1264 196 1266 204
rect 1285 196 1287 204
rect 1301 196 1303 204
rect 1317 196 1319 204
rect 1322 196 1324 204
rect 1338 196 1340 204
rect 25 56 27 64
rect 30 56 32 64
rect 46 56 48 64
rect 62 56 64 64
rect 67 56 69 64
rect 88 56 90 64
rect 104 56 106 64
rect 120 56 122 64
rect 125 56 127 64
rect 141 56 143 64
rect 157 56 159 64
rect 162 56 164 64
rect 178 56 180 64
rect 194 56 196 64
rect 199 56 201 64
rect 220 56 222 64
rect 236 56 238 64
rect 252 56 254 64
rect 257 56 259 64
rect 273 56 275 64
rect 289 56 291 64
rect 294 56 296 64
rect 310 56 312 64
rect 326 56 328 64
rect 331 56 333 64
rect 352 56 354 64
rect 368 56 370 64
rect 384 56 386 64
rect 389 56 391 64
rect 405 56 407 64
rect 958 56 960 64
rect 963 56 965 64
rect 979 56 981 64
rect 995 56 997 64
rect 1000 56 1002 64
rect 1021 56 1023 64
rect 1037 56 1039 64
rect 1053 56 1055 64
rect 1058 56 1060 64
rect 1074 56 1076 64
rect 1090 56 1092 64
rect 1095 56 1097 64
rect 1111 56 1113 64
rect 1127 56 1129 64
rect 1132 56 1134 64
rect 1153 56 1155 64
rect 1169 56 1171 64
rect 1185 56 1187 64
rect 1190 56 1192 64
rect 1206 56 1208 64
rect 1222 56 1224 64
rect 1227 56 1229 64
rect 1243 56 1245 64
rect 1259 56 1261 64
rect 1264 56 1266 64
rect 1285 56 1287 64
rect 1301 56 1303 64
rect 1317 56 1319 64
rect 1322 56 1324 64
rect 1338 56 1340 64
<< ndiffusion >>
rect 496 1914 497 1918
rect 499 1914 502 1918
rect 504 1914 505 1918
rect 517 1914 518 1918
rect 520 1914 521 1918
rect 533 1914 534 1918
rect 536 1914 539 1918
rect 541 1914 542 1918
rect 559 1914 560 1918
rect 562 1914 563 1918
rect 575 1914 576 1918
rect 578 1914 579 1918
rect 591 1914 592 1918
rect 594 1914 597 1918
rect 599 1914 600 1918
rect 612 1914 613 1918
rect 615 1914 616 1918
rect 628 1914 629 1918
rect 631 1914 634 1918
rect 636 1914 637 1918
rect 649 1914 650 1918
rect 652 1914 653 1918
rect 665 1914 666 1918
rect 668 1914 671 1918
rect 673 1914 674 1918
rect 691 1914 692 1918
rect 694 1914 695 1918
rect 707 1914 708 1918
rect 710 1914 711 1918
rect 723 1914 724 1918
rect 726 1914 729 1918
rect 731 1914 732 1918
rect 744 1914 745 1918
rect 747 1914 748 1918
rect 760 1914 761 1918
rect 763 1914 766 1918
rect 768 1914 769 1918
rect 781 1914 782 1918
rect 784 1914 785 1918
rect 797 1914 798 1918
rect 800 1914 803 1918
rect 805 1914 806 1918
rect 823 1914 824 1918
rect 826 1914 827 1918
rect 839 1914 840 1918
rect 842 1914 843 1918
rect 855 1914 856 1918
rect 858 1914 861 1918
rect 863 1914 864 1918
rect 876 1914 877 1918
rect 879 1914 880 1918
rect 892 1914 893 1918
rect 895 1914 898 1918
rect 900 1914 901 1918
rect 913 1914 914 1918
rect 916 1914 917 1918
rect 929 1914 930 1918
rect 932 1914 935 1918
rect 937 1914 938 1918
rect 955 1914 956 1918
rect 958 1914 959 1918
rect 971 1914 972 1918
rect 974 1914 975 1918
rect 987 1914 988 1918
rect 990 1914 993 1918
rect 995 1914 996 1918
rect 1008 1914 1009 1918
rect 1011 1914 1012 1918
rect 1429 1914 1430 1918
rect 1432 1914 1435 1918
rect 1437 1914 1438 1918
rect 1450 1914 1451 1918
rect 1453 1914 1454 1918
rect 1466 1914 1467 1918
rect 1469 1914 1472 1918
rect 1474 1914 1475 1918
rect 1492 1914 1493 1918
rect 1495 1914 1496 1918
rect 1508 1914 1509 1918
rect 1511 1914 1512 1918
rect 1524 1914 1525 1918
rect 1527 1914 1530 1918
rect 1532 1914 1533 1918
rect 1545 1914 1546 1918
rect 1548 1914 1549 1918
rect 1561 1914 1562 1918
rect 1564 1914 1567 1918
rect 1569 1914 1570 1918
rect 1582 1914 1583 1918
rect 1585 1914 1586 1918
rect 1598 1914 1599 1918
rect 1601 1914 1604 1918
rect 1606 1914 1607 1918
rect 1624 1914 1625 1918
rect 1627 1914 1628 1918
rect 1640 1914 1641 1918
rect 1643 1914 1644 1918
rect 1656 1914 1657 1918
rect 1659 1914 1662 1918
rect 1664 1914 1665 1918
rect 1677 1914 1678 1918
rect 1680 1914 1681 1918
rect 1693 1914 1694 1918
rect 1696 1914 1699 1918
rect 1701 1914 1702 1918
rect 1714 1914 1715 1918
rect 1717 1914 1718 1918
rect 1730 1914 1731 1918
rect 1733 1914 1736 1918
rect 1738 1914 1739 1918
rect 1756 1914 1757 1918
rect 1759 1914 1760 1918
rect 1772 1914 1773 1918
rect 1775 1914 1776 1918
rect 1788 1914 1789 1918
rect 1791 1914 1794 1918
rect 1796 1914 1797 1918
rect 1809 1914 1810 1918
rect 1812 1914 1813 1918
rect 1825 1914 1826 1918
rect 1828 1914 1831 1918
rect 1833 1914 1834 1918
rect 1846 1914 1847 1918
rect 1849 1914 1850 1918
rect 1862 1914 1863 1918
rect 1865 1914 1868 1918
rect 1870 1914 1871 1918
rect 1888 1914 1889 1918
rect 1891 1914 1892 1918
rect 1904 1914 1905 1918
rect 1907 1914 1908 1918
rect 1920 1914 1921 1918
rect 1923 1914 1926 1918
rect 1928 1914 1929 1918
rect 1941 1914 1942 1918
rect 1944 1914 1945 1918
rect 156 1881 157 1885
rect 159 1881 162 1885
rect 164 1881 165 1885
rect 177 1881 178 1885
rect 180 1881 181 1885
rect 193 1881 194 1885
rect 196 1881 199 1885
rect 201 1881 202 1885
rect 219 1881 220 1885
rect 222 1881 223 1885
rect 235 1881 236 1885
rect 238 1881 239 1885
rect 251 1881 252 1885
rect 254 1881 257 1885
rect 259 1881 260 1885
rect 272 1881 273 1885
rect 275 1881 276 1885
rect 1089 1881 1090 1885
rect 1092 1881 1095 1885
rect 1097 1881 1098 1885
rect 1110 1881 1111 1885
rect 1113 1881 1114 1885
rect 1126 1881 1127 1885
rect 1129 1881 1132 1885
rect 1134 1881 1135 1885
rect 1152 1881 1153 1885
rect 1155 1881 1156 1885
rect 1168 1881 1169 1885
rect 1171 1881 1172 1885
rect 1184 1881 1185 1885
rect 1187 1881 1190 1885
rect 1192 1881 1193 1885
rect 1205 1881 1206 1885
rect 1208 1881 1209 1885
rect 280 1844 281 1848
rect 283 1844 284 1848
rect 675 1848 676 1852
rect 678 1848 679 1852
rect 699 1844 702 1848
rect 704 1844 707 1848
rect 709 1844 710 1848
rect 756 1848 757 1852
rect 759 1848 760 1852
rect 780 1844 783 1848
rect 785 1844 788 1848
rect 790 1844 791 1848
rect 729 1840 730 1844
rect 732 1840 733 1844
rect 163 1835 164 1839
rect 166 1835 167 1839
rect 501 1835 502 1839
rect 504 1835 505 1839
rect 517 1835 518 1839
rect 520 1835 521 1839
rect 533 1835 534 1839
rect 536 1835 537 1839
rect 552 1835 557 1839
rect 559 1835 562 1839
rect 564 1835 565 1839
rect 586 1835 588 1839
rect 590 1835 591 1839
rect 608 1835 609 1839
rect 611 1835 612 1839
rect 624 1835 629 1839
rect 631 1835 634 1839
rect 636 1835 637 1839
rect 651 1835 652 1839
rect 654 1835 655 1839
rect 810 1840 811 1844
rect 813 1840 814 1844
rect 1213 1844 1214 1848
rect 1216 1844 1217 1848
rect 1608 1848 1609 1852
rect 1611 1848 1612 1852
rect 1632 1844 1635 1848
rect 1637 1844 1640 1848
rect 1642 1844 1643 1848
rect 1689 1848 1690 1852
rect 1692 1848 1693 1852
rect 1713 1844 1716 1848
rect 1718 1844 1721 1848
rect 1723 1844 1724 1848
rect 1662 1840 1663 1844
rect 1665 1840 1666 1844
rect 1096 1835 1097 1839
rect 1099 1835 1100 1839
rect 1434 1835 1435 1839
rect 1437 1835 1438 1839
rect 1450 1835 1451 1839
rect 1453 1835 1454 1839
rect 1466 1835 1467 1839
rect 1469 1835 1470 1839
rect 1485 1835 1490 1839
rect 1492 1835 1495 1839
rect 1497 1835 1498 1839
rect 1519 1835 1521 1839
rect 1523 1835 1524 1839
rect 1541 1835 1542 1839
rect 1544 1835 1545 1839
rect 1557 1835 1562 1839
rect 1564 1835 1567 1839
rect 1569 1835 1570 1839
rect 1584 1835 1585 1839
rect 1587 1835 1588 1839
rect 1743 1840 1744 1844
rect 1746 1840 1747 1844
rect 501 1789 502 1793
rect 504 1789 505 1793
rect 517 1789 518 1793
rect 520 1789 521 1793
rect 533 1789 534 1793
rect 536 1789 537 1793
rect 552 1789 557 1793
rect 559 1789 562 1793
rect 564 1789 565 1793
rect 586 1789 588 1793
rect 590 1789 591 1793
rect 608 1789 609 1793
rect 611 1789 612 1793
rect 624 1789 629 1793
rect 631 1789 634 1793
rect 636 1789 637 1793
rect 651 1789 652 1793
rect 654 1789 655 1793
rect 147 1779 148 1783
rect 150 1779 151 1783
rect 163 1779 164 1783
rect 166 1779 169 1783
rect 171 1779 172 1783
rect 184 1779 185 1783
rect 187 1779 188 1783
rect 200 1779 201 1783
rect 203 1779 204 1783
rect 221 1779 222 1783
rect 224 1779 227 1783
rect 229 1779 230 1783
rect 242 1779 243 1783
rect 245 1779 246 1783
rect 258 1779 259 1783
rect 261 1779 264 1783
rect 266 1779 267 1783
rect 699 1788 702 1792
rect 704 1788 707 1792
rect 709 1788 710 1792
rect 780 1788 783 1792
rect 785 1788 788 1792
rect 790 1788 791 1792
rect 1434 1789 1435 1793
rect 1437 1789 1438 1793
rect 1450 1789 1451 1793
rect 1453 1789 1454 1793
rect 1466 1789 1467 1793
rect 1469 1789 1470 1793
rect 1485 1789 1490 1793
rect 1492 1789 1495 1793
rect 1497 1789 1498 1793
rect 1519 1789 1521 1793
rect 1523 1789 1524 1793
rect 1541 1789 1542 1793
rect 1544 1789 1545 1793
rect 1557 1789 1562 1793
rect 1564 1789 1567 1793
rect 1569 1789 1570 1793
rect 1584 1789 1585 1793
rect 1587 1789 1588 1793
rect 1080 1779 1081 1783
rect 1083 1779 1084 1783
rect 1096 1779 1097 1783
rect 1099 1779 1102 1783
rect 1104 1779 1105 1783
rect 1117 1779 1118 1783
rect 1120 1779 1121 1783
rect 1133 1779 1134 1783
rect 1136 1779 1137 1783
rect 1154 1779 1155 1783
rect 1157 1779 1160 1783
rect 1162 1779 1163 1783
rect 1175 1779 1176 1783
rect 1178 1779 1179 1783
rect 1191 1779 1192 1783
rect 1194 1779 1197 1783
rect 1199 1779 1200 1783
rect 1632 1788 1635 1792
rect 1637 1788 1640 1792
rect 1642 1788 1643 1792
rect 1713 1788 1716 1792
rect 1718 1788 1721 1792
rect 1723 1788 1724 1792
rect 699 1712 702 1716
rect 704 1712 707 1716
rect 709 1712 710 1716
rect 780 1716 781 1720
rect 783 1716 784 1720
rect 804 1712 807 1716
rect 809 1712 812 1716
rect 814 1712 815 1716
rect 729 1708 730 1712
rect 732 1708 733 1712
rect 501 1703 502 1707
rect 504 1703 505 1707
rect 517 1703 518 1707
rect 520 1703 521 1707
rect 533 1703 534 1707
rect 536 1703 537 1707
rect 552 1703 557 1707
rect 559 1703 562 1707
rect 564 1703 565 1707
rect 586 1703 588 1707
rect 590 1703 591 1707
rect 608 1703 609 1707
rect 611 1703 612 1707
rect 624 1703 629 1707
rect 631 1703 634 1707
rect 636 1703 637 1707
rect 651 1703 652 1707
rect 654 1703 655 1707
rect 834 1708 835 1712
rect 837 1708 838 1712
rect 1632 1712 1635 1716
rect 1637 1712 1640 1716
rect 1642 1712 1643 1716
rect 1713 1716 1714 1720
rect 1716 1716 1717 1720
rect 1737 1712 1740 1716
rect 1742 1712 1745 1716
rect 1747 1712 1748 1716
rect 1662 1708 1663 1712
rect 1665 1708 1666 1712
rect 1434 1703 1435 1707
rect 1437 1703 1438 1707
rect 1450 1703 1451 1707
rect 1453 1703 1454 1707
rect 1466 1703 1467 1707
rect 1469 1703 1470 1707
rect 1485 1703 1490 1707
rect 1492 1703 1495 1707
rect 1497 1703 1498 1707
rect 1519 1703 1521 1707
rect 1523 1703 1524 1707
rect 1541 1703 1542 1707
rect 1544 1703 1545 1707
rect 1557 1703 1562 1707
rect 1564 1703 1567 1707
rect 1569 1703 1570 1707
rect 1584 1703 1585 1707
rect 1587 1703 1588 1707
rect 1767 1708 1768 1712
rect 1770 1708 1771 1712
rect 501 1657 502 1661
rect 504 1657 505 1661
rect 517 1657 518 1661
rect 520 1657 521 1661
rect 533 1657 534 1661
rect 536 1657 537 1661
rect 552 1657 557 1661
rect 559 1657 562 1661
rect 564 1657 565 1661
rect 586 1657 588 1661
rect 590 1657 591 1661
rect 608 1657 609 1661
rect 611 1657 612 1661
rect 624 1657 629 1661
rect 631 1657 634 1661
rect 636 1657 637 1661
rect 651 1657 652 1661
rect 654 1657 655 1661
rect 699 1657 702 1661
rect 704 1657 707 1661
rect 709 1657 710 1661
rect 804 1657 807 1661
rect 809 1657 812 1661
rect 814 1657 815 1661
rect 1434 1657 1435 1661
rect 1437 1657 1438 1661
rect 1450 1657 1451 1661
rect 1453 1657 1454 1661
rect 1466 1657 1467 1661
rect 1469 1657 1470 1661
rect 1485 1657 1490 1661
rect 1492 1657 1495 1661
rect 1497 1657 1498 1661
rect 1519 1657 1521 1661
rect 1523 1657 1524 1661
rect 1541 1657 1542 1661
rect 1544 1657 1545 1661
rect 1557 1657 1562 1661
rect 1564 1657 1567 1661
rect 1569 1657 1570 1661
rect 1584 1657 1585 1661
rect 1587 1657 1588 1661
rect 1632 1657 1635 1661
rect 1637 1657 1640 1661
rect 1642 1657 1643 1661
rect 1737 1657 1740 1661
rect 1742 1657 1745 1661
rect 1747 1657 1748 1661
rect 699 1580 702 1584
rect 704 1580 707 1584
rect 709 1580 710 1584
rect 756 1584 757 1588
rect 759 1584 760 1588
rect 780 1580 783 1584
rect 785 1580 788 1584
rect 790 1580 791 1584
rect 846 1584 847 1588
rect 849 1584 850 1588
rect 870 1580 873 1584
rect 875 1580 878 1584
rect 880 1580 881 1584
rect 729 1576 730 1580
rect 732 1576 733 1580
rect 501 1571 502 1575
rect 504 1571 505 1575
rect 517 1571 518 1575
rect 520 1571 521 1575
rect 533 1571 534 1575
rect 536 1571 537 1575
rect 552 1571 557 1575
rect 559 1571 562 1575
rect 564 1571 565 1575
rect 586 1571 588 1575
rect 590 1571 591 1575
rect 608 1571 609 1575
rect 611 1571 612 1575
rect 624 1571 629 1575
rect 631 1571 634 1575
rect 636 1571 637 1575
rect 651 1571 652 1575
rect 654 1571 655 1575
rect 810 1576 811 1580
rect 813 1576 814 1580
rect 900 1576 901 1580
rect 903 1576 904 1580
rect 1632 1580 1635 1584
rect 1637 1580 1640 1584
rect 1642 1580 1643 1584
rect 1689 1584 1690 1588
rect 1692 1584 1693 1588
rect 1713 1580 1716 1584
rect 1718 1580 1721 1584
rect 1723 1580 1724 1584
rect 1779 1584 1780 1588
rect 1782 1584 1783 1588
rect 1803 1580 1806 1584
rect 1808 1580 1811 1584
rect 1813 1580 1814 1584
rect 1662 1576 1663 1580
rect 1665 1576 1666 1580
rect 1434 1571 1435 1575
rect 1437 1571 1438 1575
rect 1450 1571 1451 1575
rect 1453 1571 1454 1575
rect 1466 1571 1467 1575
rect 1469 1571 1470 1575
rect 1485 1571 1490 1575
rect 1492 1571 1495 1575
rect 1497 1571 1498 1575
rect 1519 1571 1521 1575
rect 1523 1571 1524 1575
rect 1541 1571 1542 1575
rect 1544 1571 1545 1575
rect 1557 1571 1562 1575
rect 1564 1571 1567 1575
rect 1569 1571 1570 1575
rect 1584 1571 1585 1575
rect 1587 1571 1588 1575
rect 1743 1576 1744 1580
rect 1746 1576 1747 1580
rect 1833 1576 1834 1580
rect 1836 1576 1837 1580
rect 501 1525 502 1529
rect 504 1525 505 1529
rect 517 1525 518 1529
rect 520 1525 521 1529
rect 533 1525 534 1529
rect 536 1525 537 1529
rect 552 1525 557 1529
rect 559 1525 562 1529
rect 564 1525 565 1529
rect 586 1525 588 1529
rect 590 1525 591 1529
rect 608 1525 609 1529
rect 611 1525 612 1529
rect 624 1525 629 1529
rect 631 1525 634 1529
rect 636 1525 637 1529
rect 651 1525 652 1529
rect 654 1525 655 1529
rect 699 1522 702 1526
rect 704 1522 707 1526
rect 709 1522 710 1526
rect 780 1522 783 1526
rect 785 1522 788 1526
rect 790 1522 791 1526
rect 870 1522 873 1526
rect 875 1522 878 1526
rect 880 1522 881 1526
rect 1434 1525 1435 1529
rect 1437 1525 1438 1529
rect 1450 1525 1451 1529
rect 1453 1525 1454 1529
rect 1466 1525 1467 1529
rect 1469 1525 1470 1529
rect 1485 1525 1490 1529
rect 1492 1525 1495 1529
rect 1497 1525 1498 1529
rect 1519 1525 1521 1529
rect 1523 1525 1524 1529
rect 1541 1525 1542 1529
rect 1544 1525 1545 1529
rect 1557 1525 1562 1529
rect 1564 1525 1567 1529
rect 1569 1525 1570 1529
rect 1584 1525 1585 1529
rect 1587 1525 1588 1529
rect 1632 1522 1635 1526
rect 1637 1522 1640 1526
rect 1642 1522 1643 1526
rect 1713 1522 1716 1526
rect 1718 1522 1721 1526
rect 1723 1522 1724 1526
rect 1803 1522 1806 1526
rect 1808 1522 1811 1526
rect 1813 1522 1814 1526
rect 699 1448 702 1452
rect 704 1448 707 1452
rect 709 1448 710 1452
rect 729 1444 730 1448
rect 732 1444 733 1448
rect 501 1439 502 1443
rect 504 1439 505 1443
rect 517 1439 518 1443
rect 520 1439 521 1443
rect 533 1439 534 1443
rect 536 1439 537 1443
rect 552 1439 557 1443
rect 559 1439 562 1443
rect 564 1439 565 1443
rect 586 1439 588 1443
rect 590 1439 591 1443
rect 608 1439 609 1443
rect 611 1439 612 1443
rect 624 1439 629 1443
rect 631 1439 634 1443
rect 636 1439 637 1443
rect 651 1439 652 1443
rect 654 1439 655 1443
rect 1632 1448 1635 1452
rect 1637 1448 1640 1452
rect 1642 1448 1643 1452
rect 1662 1444 1663 1448
rect 1665 1444 1666 1448
rect 1434 1439 1435 1443
rect 1437 1439 1438 1443
rect 1450 1439 1451 1443
rect 1453 1439 1454 1443
rect 1466 1439 1467 1443
rect 1469 1439 1470 1443
rect 1485 1439 1490 1443
rect 1492 1439 1495 1443
rect 1497 1439 1498 1443
rect 1519 1439 1521 1443
rect 1523 1439 1524 1443
rect 1541 1439 1542 1443
rect 1544 1439 1545 1443
rect 1557 1439 1562 1443
rect 1564 1439 1567 1443
rect 1569 1439 1570 1443
rect 1584 1439 1585 1443
rect 1587 1439 1588 1443
rect 501 1393 502 1397
rect 504 1393 505 1397
rect 517 1393 518 1397
rect 520 1393 521 1397
rect 533 1393 534 1397
rect 536 1393 537 1397
rect 552 1393 557 1397
rect 559 1393 562 1397
rect 564 1393 565 1397
rect 586 1393 588 1397
rect 590 1393 591 1397
rect 608 1393 609 1397
rect 611 1393 612 1397
rect 624 1393 629 1397
rect 631 1393 634 1397
rect 636 1393 637 1397
rect 651 1393 652 1397
rect 654 1393 655 1397
rect 735 1393 736 1397
rect 738 1393 739 1397
rect 743 1393 749 1397
rect 753 1393 754 1397
rect 756 1393 757 1397
rect 778 1393 779 1397
rect 781 1393 782 1397
rect 794 1393 795 1397
rect 797 1393 798 1397
rect 813 1393 818 1397
rect 820 1393 823 1397
rect 825 1393 826 1397
rect 847 1393 849 1397
rect 851 1393 852 1397
rect 869 1393 870 1397
rect 872 1393 873 1397
rect 885 1393 890 1397
rect 892 1393 895 1397
rect 897 1393 898 1397
rect 912 1393 913 1397
rect 915 1393 916 1397
rect 24 1379 25 1383
rect 27 1379 30 1383
rect 32 1379 33 1383
rect 45 1379 46 1383
rect 48 1379 49 1383
rect 61 1379 62 1383
rect 64 1379 67 1383
rect 69 1379 70 1383
rect 87 1379 88 1383
rect 90 1379 91 1383
rect 103 1379 104 1383
rect 106 1379 107 1383
rect 119 1379 120 1383
rect 122 1379 125 1383
rect 127 1379 128 1383
rect 140 1379 141 1383
rect 143 1379 144 1383
rect 156 1379 157 1383
rect 159 1379 162 1383
rect 164 1379 165 1383
rect 177 1379 178 1383
rect 180 1379 181 1383
rect 193 1379 194 1383
rect 196 1379 199 1383
rect 201 1379 202 1383
rect 219 1379 220 1383
rect 222 1379 223 1383
rect 235 1379 236 1383
rect 238 1379 239 1383
rect 251 1379 252 1383
rect 254 1379 257 1383
rect 259 1379 260 1383
rect 272 1379 273 1383
rect 275 1379 276 1383
rect 288 1379 289 1383
rect 291 1379 294 1383
rect 296 1379 297 1383
rect 309 1379 310 1383
rect 312 1379 313 1383
rect 325 1379 326 1383
rect 328 1379 331 1383
rect 333 1379 334 1383
rect 351 1379 352 1383
rect 354 1379 355 1383
rect 367 1379 368 1383
rect 370 1379 371 1383
rect 383 1379 384 1383
rect 386 1379 389 1383
rect 391 1379 392 1383
rect 404 1379 405 1383
rect 407 1379 408 1383
rect 699 1386 702 1390
rect 704 1386 707 1390
rect 709 1386 710 1390
rect 1434 1393 1435 1397
rect 1437 1393 1438 1397
rect 1450 1393 1451 1397
rect 1453 1393 1454 1397
rect 1466 1393 1467 1397
rect 1469 1393 1470 1397
rect 1485 1393 1490 1397
rect 1492 1393 1495 1397
rect 1497 1393 1498 1397
rect 1519 1393 1521 1397
rect 1523 1393 1524 1397
rect 1541 1393 1542 1397
rect 1544 1393 1545 1397
rect 1557 1393 1562 1397
rect 1564 1393 1567 1397
rect 1569 1393 1570 1397
rect 1584 1393 1585 1397
rect 1587 1393 1588 1397
rect 1668 1393 1669 1397
rect 1671 1393 1672 1397
rect 1676 1393 1682 1397
rect 1686 1393 1687 1397
rect 1689 1393 1690 1397
rect 1711 1393 1712 1397
rect 1714 1393 1715 1397
rect 1727 1393 1728 1397
rect 1730 1393 1731 1397
rect 1746 1393 1751 1397
rect 1753 1393 1756 1397
rect 1758 1393 1759 1397
rect 1780 1393 1782 1397
rect 1784 1393 1785 1397
rect 1802 1393 1803 1397
rect 1805 1393 1806 1397
rect 1818 1393 1823 1397
rect 1825 1393 1828 1397
rect 1830 1393 1831 1397
rect 1845 1393 1846 1397
rect 1848 1393 1849 1397
rect 957 1379 958 1383
rect 960 1379 963 1383
rect 965 1379 966 1383
rect 978 1379 979 1383
rect 981 1379 982 1383
rect 994 1379 995 1383
rect 997 1379 1000 1383
rect 1002 1379 1003 1383
rect 1020 1379 1021 1383
rect 1023 1379 1024 1383
rect 1036 1379 1037 1383
rect 1039 1379 1040 1383
rect 1052 1379 1053 1383
rect 1055 1379 1058 1383
rect 1060 1379 1061 1383
rect 1073 1379 1074 1383
rect 1076 1379 1077 1383
rect 1089 1379 1090 1383
rect 1092 1379 1095 1383
rect 1097 1379 1098 1383
rect 1110 1379 1111 1383
rect 1113 1379 1114 1383
rect 1126 1379 1127 1383
rect 1129 1379 1132 1383
rect 1134 1379 1135 1383
rect 1152 1379 1153 1383
rect 1155 1379 1156 1383
rect 1168 1379 1169 1383
rect 1171 1379 1172 1383
rect 1184 1379 1185 1383
rect 1187 1379 1190 1383
rect 1192 1379 1193 1383
rect 1205 1379 1206 1383
rect 1208 1379 1209 1383
rect 1221 1379 1222 1383
rect 1224 1379 1227 1383
rect 1229 1379 1230 1383
rect 1242 1379 1243 1383
rect 1245 1379 1246 1383
rect 1258 1379 1259 1383
rect 1261 1379 1264 1383
rect 1266 1379 1267 1383
rect 1284 1379 1285 1383
rect 1287 1379 1288 1383
rect 1300 1379 1301 1383
rect 1303 1379 1304 1383
rect 1316 1379 1317 1383
rect 1319 1379 1322 1383
rect 1324 1379 1325 1383
rect 1337 1379 1338 1383
rect 1340 1379 1341 1383
rect 1632 1386 1635 1390
rect 1637 1386 1640 1390
rect 1642 1386 1643 1390
rect 139 1335 140 1339
rect 142 1335 143 1339
rect 163 1335 164 1339
rect 166 1335 167 1339
rect 925 1339 929 1340
rect 925 1336 929 1337
rect 1072 1335 1073 1339
rect 1075 1335 1076 1339
rect 1096 1335 1097 1339
rect 1099 1335 1100 1339
rect 1858 1339 1862 1340
rect 1858 1336 1862 1337
rect 159 1324 160 1328
rect 162 1324 163 1328
rect 1092 1324 1093 1328
rect 1095 1324 1096 1328
rect 151 1312 155 1313
rect 151 1309 155 1310
rect 1084 1312 1088 1313
rect 1084 1309 1088 1310
rect 139 1301 140 1305
rect 142 1301 143 1305
rect 163 1301 164 1305
rect 166 1301 167 1305
rect 1072 1301 1073 1305
rect 1075 1301 1076 1305
rect 1096 1301 1097 1305
rect 1099 1301 1100 1305
rect 795 1269 796 1273
rect 798 1269 801 1273
rect 803 1269 804 1273
rect 816 1269 817 1273
rect 819 1269 820 1273
rect 832 1269 833 1273
rect 835 1269 838 1273
rect 840 1269 841 1273
rect 858 1269 859 1273
rect 861 1269 862 1273
rect 874 1269 875 1273
rect 877 1269 878 1273
rect 890 1269 891 1273
rect 893 1269 896 1273
rect 898 1269 899 1273
rect 911 1269 912 1273
rect 914 1269 915 1273
rect 1728 1269 1729 1273
rect 1731 1269 1734 1273
rect 1736 1269 1737 1273
rect 1749 1269 1750 1273
rect 1752 1269 1753 1273
rect 1765 1269 1766 1273
rect 1768 1269 1771 1273
rect 1773 1269 1774 1273
rect 1791 1269 1792 1273
rect 1794 1269 1795 1273
rect 1807 1269 1808 1273
rect 1810 1269 1811 1273
rect 1823 1269 1824 1273
rect 1826 1269 1829 1273
rect 1831 1269 1832 1273
rect 1844 1269 1845 1273
rect 1847 1269 1848 1273
rect 24 1239 25 1243
rect 27 1239 30 1243
rect 32 1239 33 1243
rect 45 1239 46 1243
rect 48 1239 49 1243
rect 61 1239 62 1243
rect 64 1239 67 1243
rect 69 1239 70 1243
rect 87 1239 88 1243
rect 90 1239 91 1243
rect 103 1239 104 1243
rect 106 1239 107 1243
rect 119 1239 120 1243
rect 122 1239 125 1243
rect 127 1239 128 1243
rect 140 1239 141 1243
rect 143 1239 144 1243
rect 156 1239 157 1243
rect 159 1239 162 1243
rect 164 1239 165 1243
rect 177 1239 178 1243
rect 180 1239 181 1243
rect 193 1239 194 1243
rect 196 1239 199 1243
rect 201 1239 202 1243
rect 219 1239 220 1243
rect 222 1239 223 1243
rect 235 1239 236 1243
rect 238 1239 239 1243
rect 251 1239 252 1243
rect 254 1239 257 1243
rect 259 1239 260 1243
rect 272 1239 273 1243
rect 275 1239 276 1243
rect 288 1239 289 1243
rect 291 1239 294 1243
rect 296 1239 297 1243
rect 309 1239 310 1243
rect 312 1239 313 1243
rect 325 1239 326 1243
rect 328 1239 331 1243
rect 333 1239 334 1243
rect 351 1239 352 1243
rect 354 1239 355 1243
rect 367 1239 368 1243
rect 370 1239 371 1243
rect 383 1239 384 1243
rect 386 1239 389 1243
rect 391 1239 392 1243
rect 404 1239 405 1243
rect 407 1239 408 1243
rect 957 1239 958 1243
rect 960 1239 963 1243
rect 965 1239 966 1243
rect 978 1239 979 1243
rect 981 1239 982 1243
rect 994 1239 995 1243
rect 997 1239 1000 1243
rect 1002 1239 1003 1243
rect 1020 1239 1021 1243
rect 1023 1239 1024 1243
rect 1036 1239 1037 1243
rect 1039 1239 1040 1243
rect 1052 1239 1053 1243
rect 1055 1239 1058 1243
rect 1060 1239 1061 1243
rect 1073 1239 1074 1243
rect 1076 1239 1077 1243
rect 1089 1239 1090 1243
rect 1092 1239 1095 1243
rect 1097 1239 1098 1243
rect 1110 1239 1111 1243
rect 1113 1239 1114 1243
rect 1126 1239 1127 1243
rect 1129 1239 1132 1243
rect 1134 1239 1135 1243
rect 1152 1239 1153 1243
rect 1155 1239 1156 1243
rect 1168 1239 1169 1243
rect 1171 1239 1172 1243
rect 1184 1239 1185 1243
rect 1187 1239 1190 1243
rect 1192 1239 1193 1243
rect 1205 1239 1206 1243
rect 1208 1239 1209 1243
rect 1221 1239 1222 1243
rect 1224 1239 1227 1243
rect 1229 1239 1230 1243
rect 1242 1239 1243 1243
rect 1245 1239 1246 1243
rect 1258 1239 1259 1243
rect 1261 1239 1264 1243
rect 1266 1239 1267 1243
rect 1284 1239 1285 1243
rect 1287 1239 1288 1243
rect 1300 1239 1301 1243
rect 1303 1239 1304 1243
rect 1316 1239 1317 1243
rect 1319 1239 1322 1243
rect 1324 1239 1325 1243
rect 1337 1239 1338 1243
rect 1340 1239 1341 1243
rect 937 1195 941 1196
rect 937 1192 941 1193
rect 1870 1195 1874 1196
rect 1870 1192 1874 1193
rect 795 1183 796 1187
rect 798 1183 801 1187
rect 803 1183 804 1187
rect 816 1183 817 1187
rect 819 1183 820 1187
rect 832 1183 833 1187
rect 835 1183 838 1187
rect 840 1183 841 1187
rect 858 1183 859 1187
rect 861 1183 862 1187
rect 874 1183 875 1187
rect 877 1183 878 1187
rect 890 1183 891 1187
rect 893 1183 896 1187
rect 898 1183 899 1187
rect 911 1183 912 1187
rect 914 1183 915 1187
rect 1728 1183 1729 1187
rect 1731 1183 1734 1187
rect 1736 1183 1737 1187
rect 1749 1183 1750 1187
rect 1752 1183 1753 1187
rect 1765 1183 1766 1187
rect 1768 1183 1771 1187
rect 1773 1183 1774 1187
rect 1791 1183 1792 1187
rect 1794 1183 1795 1187
rect 1807 1183 1808 1187
rect 1810 1183 1811 1187
rect 1823 1183 1824 1187
rect 1826 1183 1829 1187
rect 1831 1183 1832 1187
rect 1844 1183 1845 1187
rect 1847 1183 1848 1187
rect 24 1153 25 1157
rect 27 1153 30 1157
rect 32 1153 33 1157
rect 45 1153 46 1157
rect 48 1153 49 1157
rect 61 1153 62 1157
rect 64 1153 67 1157
rect 69 1153 70 1157
rect 87 1153 88 1157
rect 90 1153 91 1157
rect 103 1153 104 1157
rect 106 1153 107 1157
rect 119 1153 120 1157
rect 122 1153 125 1157
rect 127 1153 128 1157
rect 140 1153 141 1157
rect 143 1153 144 1157
rect 156 1153 157 1157
rect 159 1153 162 1157
rect 164 1153 165 1157
rect 177 1153 178 1157
rect 180 1153 181 1157
rect 193 1153 194 1157
rect 196 1153 199 1157
rect 201 1153 202 1157
rect 219 1153 220 1157
rect 222 1153 223 1157
rect 235 1153 236 1157
rect 238 1153 239 1157
rect 251 1153 252 1157
rect 254 1153 257 1157
rect 259 1153 260 1157
rect 272 1153 273 1157
rect 275 1153 276 1157
rect 288 1153 289 1157
rect 291 1153 294 1157
rect 296 1153 297 1157
rect 309 1153 310 1157
rect 312 1153 313 1157
rect 325 1153 326 1157
rect 328 1153 331 1157
rect 333 1153 334 1157
rect 351 1153 352 1157
rect 354 1153 355 1157
rect 367 1153 368 1157
rect 370 1153 371 1157
rect 383 1153 384 1157
rect 386 1153 389 1157
rect 391 1153 392 1157
rect 404 1153 405 1157
rect 407 1153 408 1157
rect 957 1153 958 1157
rect 960 1153 963 1157
rect 965 1153 966 1157
rect 978 1153 979 1157
rect 981 1153 982 1157
rect 994 1153 995 1157
rect 997 1153 1000 1157
rect 1002 1153 1003 1157
rect 1020 1153 1021 1157
rect 1023 1153 1024 1157
rect 1036 1153 1037 1157
rect 1039 1153 1040 1157
rect 1052 1153 1053 1157
rect 1055 1153 1058 1157
rect 1060 1153 1061 1157
rect 1073 1153 1074 1157
rect 1076 1153 1077 1157
rect 1089 1153 1090 1157
rect 1092 1153 1095 1157
rect 1097 1153 1098 1157
rect 1110 1153 1111 1157
rect 1113 1153 1114 1157
rect 1126 1153 1127 1157
rect 1129 1153 1132 1157
rect 1134 1153 1135 1157
rect 1152 1153 1153 1157
rect 1155 1153 1156 1157
rect 1168 1153 1169 1157
rect 1171 1153 1172 1157
rect 1184 1153 1185 1157
rect 1187 1153 1190 1157
rect 1192 1153 1193 1157
rect 1205 1153 1206 1157
rect 1208 1153 1209 1157
rect 1221 1153 1222 1157
rect 1224 1153 1227 1157
rect 1229 1153 1230 1157
rect 1242 1153 1243 1157
rect 1245 1153 1246 1157
rect 1258 1153 1259 1157
rect 1261 1153 1264 1157
rect 1266 1153 1267 1157
rect 1284 1153 1285 1157
rect 1287 1153 1288 1157
rect 1300 1153 1301 1157
rect 1303 1153 1304 1157
rect 1316 1153 1317 1157
rect 1319 1153 1322 1157
rect 1324 1153 1325 1157
rect 1337 1153 1338 1157
rect 1340 1153 1341 1157
rect 256 1109 257 1113
rect 259 1109 260 1113
rect 280 1109 281 1113
rect 283 1109 284 1113
rect 1189 1109 1190 1113
rect 1192 1109 1193 1113
rect 1213 1109 1214 1113
rect 1216 1109 1217 1113
rect 276 1098 277 1102
rect 279 1098 280 1102
rect 1209 1098 1210 1102
rect 1212 1098 1213 1102
rect 268 1086 272 1087
rect 268 1083 272 1084
rect 1201 1086 1205 1087
rect 1201 1083 1205 1084
rect 256 1075 257 1079
rect 259 1075 260 1079
rect 280 1075 281 1079
rect 283 1075 284 1079
rect 1189 1075 1190 1079
rect 1192 1075 1193 1079
rect 1213 1075 1214 1079
rect 1216 1075 1217 1079
rect 24 1013 25 1017
rect 27 1013 30 1017
rect 32 1013 33 1017
rect 45 1013 46 1017
rect 48 1013 49 1017
rect 61 1013 62 1017
rect 64 1013 67 1017
rect 69 1013 70 1017
rect 87 1013 88 1017
rect 90 1013 91 1017
rect 103 1013 104 1017
rect 106 1013 107 1017
rect 119 1013 120 1017
rect 122 1013 125 1017
rect 127 1013 128 1017
rect 140 1013 141 1017
rect 143 1013 144 1017
rect 156 1013 157 1017
rect 159 1013 162 1017
rect 164 1013 165 1017
rect 177 1013 178 1017
rect 180 1013 181 1017
rect 193 1013 194 1017
rect 196 1013 199 1017
rect 201 1013 202 1017
rect 219 1013 220 1017
rect 222 1013 223 1017
rect 235 1013 236 1017
rect 238 1013 239 1017
rect 251 1013 252 1017
rect 254 1013 257 1017
rect 259 1013 260 1017
rect 272 1013 273 1017
rect 275 1013 276 1017
rect 288 1013 289 1017
rect 291 1013 294 1017
rect 296 1013 297 1017
rect 309 1013 310 1017
rect 312 1013 313 1017
rect 325 1013 326 1017
rect 328 1013 331 1017
rect 333 1013 334 1017
rect 351 1013 352 1017
rect 354 1013 355 1017
rect 367 1013 368 1017
rect 370 1013 371 1017
rect 383 1013 384 1017
rect 386 1013 389 1017
rect 391 1013 392 1017
rect 404 1013 405 1017
rect 407 1013 408 1017
rect 957 1013 958 1017
rect 960 1013 963 1017
rect 965 1013 966 1017
rect 978 1013 979 1017
rect 981 1013 982 1017
rect 994 1013 995 1017
rect 997 1013 1000 1017
rect 1002 1013 1003 1017
rect 1020 1013 1021 1017
rect 1023 1013 1024 1017
rect 1036 1013 1037 1017
rect 1039 1013 1040 1017
rect 1052 1013 1053 1017
rect 1055 1013 1058 1017
rect 1060 1013 1061 1017
rect 1073 1013 1074 1017
rect 1076 1013 1077 1017
rect 1089 1013 1090 1017
rect 1092 1013 1095 1017
rect 1097 1013 1098 1017
rect 1110 1013 1111 1017
rect 1113 1013 1114 1017
rect 1126 1013 1127 1017
rect 1129 1013 1132 1017
rect 1134 1013 1135 1017
rect 1152 1013 1153 1017
rect 1155 1013 1156 1017
rect 1168 1013 1169 1017
rect 1171 1013 1172 1017
rect 1184 1013 1185 1017
rect 1187 1013 1190 1017
rect 1192 1013 1193 1017
rect 1205 1013 1206 1017
rect 1208 1013 1209 1017
rect 1221 1013 1222 1017
rect 1224 1013 1227 1017
rect 1229 1013 1230 1017
rect 1242 1013 1243 1017
rect 1245 1013 1246 1017
rect 1258 1013 1259 1017
rect 1261 1013 1264 1017
rect 1266 1013 1267 1017
rect 1284 1013 1285 1017
rect 1287 1013 1288 1017
rect 1300 1013 1301 1017
rect 1303 1013 1304 1017
rect 1316 1013 1317 1017
rect 1319 1013 1322 1017
rect 1324 1013 1325 1017
rect 1337 1013 1338 1017
rect 1340 1013 1341 1017
rect 496 934 497 938
rect 499 934 502 938
rect 504 934 505 938
rect 517 934 518 938
rect 520 934 521 938
rect 533 934 534 938
rect 536 934 539 938
rect 541 934 542 938
rect 559 934 560 938
rect 562 934 563 938
rect 575 934 576 938
rect 578 934 579 938
rect 591 934 592 938
rect 594 934 597 938
rect 599 934 600 938
rect 612 934 613 938
rect 615 934 616 938
rect 628 934 629 938
rect 631 934 634 938
rect 636 934 637 938
rect 649 934 650 938
rect 652 934 653 938
rect 665 934 666 938
rect 668 934 671 938
rect 673 934 674 938
rect 691 934 692 938
rect 694 934 695 938
rect 707 934 708 938
rect 710 934 711 938
rect 723 934 724 938
rect 726 934 729 938
rect 731 934 732 938
rect 744 934 745 938
rect 747 934 748 938
rect 760 934 761 938
rect 763 934 766 938
rect 768 934 769 938
rect 781 934 782 938
rect 784 934 785 938
rect 797 934 798 938
rect 800 934 803 938
rect 805 934 806 938
rect 823 934 824 938
rect 826 934 827 938
rect 839 934 840 938
rect 842 934 843 938
rect 855 934 856 938
rect 858 934 861 938
rect 863 934 864 938
rect 876 934 877 938
rect 879 934 880 938
rect 892 934 893 938
rect 895 934 898 938
rect 900 934 901 938
rect 913 934 914 938
rect 916 934 917 938
rect 929 934 930 938
rect 932 934 935 938
rect 937 934 938 938
rect 955 934 956 938
rect 958 934 959 938
rect 971 934 972 938
rect 974 934 975 938
rect 987 934 988 938
rect 990 934 993 938
rect 995 934 996 938
rect 1008 934 1009 938
rect 1011 934 1012 938
rect 1429 934 1430 938
rect 1432 934 1435 938
rect 1437 934 1438 938
rect 1450 934 1451 938
rect 1453 934 1454 938
rect 1466 934 1467 938
rect 1469 934 1472 938
rect 1474 934 1475 938
rect 1492 934 1493 938
rect 1495 934 1496 938
rect 1508 934 1509 938
rect 1511 934 1512 938
rect 1524 934 1525 938
rect 1527 934 1530 938
rect 1532 934 1533 938
rect 1545 934 1546 938
rect 1548 934 1549 938
rect 1561 934 1562 938
rect 1564 934 1567 938
rect 1569 934 1570 938
rect 1582 934 1583 938
rect 1585 934 1586 938
rect 1598 934 1599 938
rect 1601 934 1604 938
rect 1606 934 1607 938
rect 1624 934 1625 938
rect 1627 934 1628 938
rect 1640 934 1641 938
rect 1643 934 1644 938
rect 1656 934 1657 938
rect 1659 934 1662 938
rect 1664 934 1665 938
rect 1677 934 1678 938
rect 1680 934 1681 938
rect 1693 934 1694 938
rect 1696 934 1699 938
rect 1701 934 1702 938
rect 1714 934 1715 938
rect 1717 934 1718 938
rect 1730 934 1731 938
rect 1733 934 1736 938
rect 1738 934 1739 938
rect 1756 934 1757 938
rect 1759 934 1760 938
rect 1772 934 1773 938
rect 1775 934 1776 938
rect 1788 934 1789 938
rect 1791 934 1794 938
rect 1796 934 1797 938
rect 1809 934 1810 938
rect 1812 934 1813 938
rect 1825 934 1826 938
rect 1828 934 1831 938
rect 1833 934 1834 938
rect 1846 934 1847 938
rect 1849 934 1850 938
rect 1862 934 1863 938
rect 1865 934 1868 938
rect 1870 934 1871 938
rect 1888 934 1889 938
rect 1891 934 1892 938
rect 1904 934 1905 938
rect 1907 934 1908 938
rect 1920 934 1921 938
rect 1923 934 1926 938
rect 1928 934 1929 938
rect 1941 934 1942 938
rect 1944 934 1945 938
rect 156 901 157 905
rect 159 901 162 905
rect 164 901 165 905
rect 177 901 178 905
rect 180 901 181 905
rect 193 901 194 905
rect 196 901 199 905
rect 201 901 202 905
rect 219 901 220 905
rect 222 901 223 905
rect 235 901 236 905
rect 238 901 239 905
rect 251 901 252 905
rect 254 901 257 905
rect 259 901 260 905
rect 272 901 273 905
rect 275 901 276 905
rect 1089 901 1090 905
rect 1092 901 1095 905
rect 1097 901 1098 905
rect 1110 901 1111 905
rect 1113 901 1114 905
rect 1126 901 1127 905
rect 1129 901 1132 905
rect 1134 901 1135 905
rect 1152 901 1153 905
rect 1155 901 1156 905
rect 1168 901 1169 905
rect 1171 901 1172 905
rect 1184 901 1185 905
rect 1187 901 1190 905
rect 1192 901 1193 905
rect 1205 901 1206 905
rect 1208 901 1209 905
rect 280 864 281 868
rect 283 864 284 868
rect 675 868 676 872
rect 678 868 679 872
rect 699 864 702 868
rect 704 864 707 868
rect 709 864 710 868
rect 756 868 757 872
rect 759 868 760 872
rect 780 864 783 868
rect 785 864 788 868
rect 790 864 791 868
rect 729 860 730 864
rect 732 860 733 864
rect 163 855 164 859
rect 166 855 167 859
rect 501 855 502 859
rect 504 855 505 859
rect 517 855 518 859
rect 520 855 521 859
rect 533 855 534 859
rect 536 855 537 859
rect 552 855 557 859
rect 559 855 562 859
rect 564 855 565 859
rect 586 855 588 859
rect 590 855 591 859
rect 608 855 609 859
rect 611 855 612 859
rect 624 855 629 859
rect 631 855 634 859
rect 636 855 637 859
rect 651 855 652 859
rect 654 855 655 859
rect 810 860 811 864
rect 813 860 814 864
rect 1213 864 1214 868
rect 1216 864 1217 868
rect 1608 868 1609 872
rect 1611 868 1612 872
rect 1632 864 1635 868
rect 1637 864 1640 868
rect 1642 864 1643 868
rect 1689 868 1690 872
rect 1692 868 1693 872
rect 1713 864 1716 868
rect 1718 864 1721 868
rect 1723 864 1724 868
rect 1662 860 1663 864
rect 1665 860 1666 864
rect 1096 855 1097 859
rect 1099 855 1100 859
rect 1434 855 1435 859
rect 1437 855 1438 859
rect 1450 855 1451 859
rect 1453 855 1454 859
rect 1466 855 1467 859
rect 1469 855 1470 859
rect 1485 855 1490 859
rect 1492 855 1495 859
rect 1497 855 1498 859
rect 1519 855 1521 859
rect 1523 855 1524 859
rect 1541 855 1542 859
rect 1544 855 1545 859
rect 1557 855 1562 859
rect 1564 855 1567 859
rect 1569 855 1570 859
rect 1584 855 1585 859
rect 1587 855 1588 859
rect 1743 860 1744 864
rect 1746 860 1747 864
rect 501 809 502 813
rect 504 809 505 813
rect 517 809 518 813
rect 520 809 521 813
rect 533 809 534 813
rect 536 809 537 813
rect 552 809 557 813
rect 559 809 562 813
rect 564 809 565 813
rect 586 809 588 813
rect 590 809 591 813
rect 608 809 609 813
rect 611 809 612 813
rect 624 809 629 813
rect 631 809 634 813
rect 636 809 637 813
rect 651 809 652 813
rect 654 809 655 813
rect 147 799 148 803
rect 150 799 151 803
rect 163 799 164 803
rect 166 799 169 803
rect 171 799 172 803
rect 184 799 185 803
rect 187 799 188 803
rect 200 799 201 803
rect 203 799 204 803
rect 221 799 222 803
rect 224 799 227 803
rect 229 799 230 803
rect 242 799 243 803
rect 245 799 246 803
rect 258 799 259 803
rect 261 799 264 803
rect 266 799 267 803
rect 699 808 702 812
rect 704 808 707 812
rect 709 808 710 812
rect 780 808 783 812
rect 785 808 788 812
rect 790 808 791 812
rect 1434 809 1435 813
rect 1437 809 1438 813
rect 1450 809 1451 813
rect 1453 809 1454 813
rect 1466 809 1467 813
rect 1469 809 1470 813
rect 1485 809 1490 813
rect 1492 809 1495 813
rect 1497 809 1498 813
rect 1519 809 1521 813
rect 1523 809 1524 813
rect 1541 809 1542 813
rect 1544 809 1545 813
rect 1557 809 1562 813
rect 1564 809 1567 813
rect 1569 809 1570 813
rect 1584 809 1585 813
rect 1587 809 1588 813
rect 1080 799 1081 803
rect 1083 799 1084 803
rect 1096 799 1097 803
rect 1099 799 1102 803
rect 1104 799 1105 803
rect 1117 799 1118 803
rect 1120 799 1121 803
rect 1133 799 1134 803
rect 1136 799 1137 803
rect 1154 799 1155 803
rect 1157 799 1160 803
rect 1162 799 1163 803
rect 1175 799 1176 803
rect 1178 799 1179 803
rect 1191 799 1192 803
rect 1194 799 1197 803
rect 1199 799 1200 803
rect 1632 808 1635 812
rect 1637 808 1640 812
rect 1642 808 1643 812
rect 1713 808 1716 812
rect 1718 808 1721 812
rect 1723 808 1724 812
rect 699 732 702 736
rect 704 732 707 736
rect 709 732 710 736
rect 780 736 781 740
rect 783 736 784 740
rect 804 732 807 736
rect 809 732 812 736
rect 814 732 815 736
rect 729 728 730 732
rect 732 728 733 732
rect 501 723 502 727
rect 504 723 505 727
rect 517 723 518 727
rect 520 723 521 727
rect 533 723 534 727
rect 536 723 537 727
rect 552 723 557 727
rect 559 723 562 727
rect 564 723 565 727
rect 586 723 588 727
rect 590 723 591 727
rect 608 723 609 727
rect 611 723 612 727
rect 624 723 629 727
rect 631 723 634 727
rect 636 723 637 727
rect 651 723 652 727
rect 654 723 655 727
rect 834 728 835 732
rect 837 728 838 732
rect 1632 732 1635 736
rect 1637 732 1640 736
rect 1642 732 1643 736
rect 1713 736 1714 740
rect 1716 736 1717 740
rect 1737 732 1740 736
rect 1742 732 1745 736
rect 1747 732 1748 736
rect 1662 728 1663 732
rect 1665 728 1666 732
rect 1434 723 1435 727
rect 1437 723 1438 727
rect 1450 723 1451 727
rect 1453 723 1454 727
rect 1466 723 1467 727
rect 1469 723 1470 727
rect 1485 723 1490 727
rect 1492 723 1495 727
rect 1497 723 1498 727
rect 1519 723 1521 727
rect 1523 723 1524 727
rect 1541 723 1542 727
rect 1544 723 1545 727
rect 1557 723 1562 727
rect 1564 723 1567 727
rect 1569 723 1570 727
rect 1584 723 1585 727
rect 1587 723 1588 727
rect 1767 728 1768 732
rect 1770 728 1771 732
rect 501 677 502 681
rect 504 677 505 681
rect 517 677 518 681
rect 520 677 521 681
rect 533 677 534 681
rect 536 677 537 681
rect 552 677 557 681
rect 559 677 562 681
rect 564 677 565 681
rect 586 677 588 681
rect 590 677 591 681
rect 608 677 609 681
rect 611 677 612 681
rect 624 677 629 681
rect 631 677 634 681
rect 636 677 637 681
rect 651 677 652 681
rect 654 677 655 681
rect 699 677 702 681
rect 704 677 707 681
rect 709 677 710 681
rect 804 677 807 681
rect 809 677 812 681
rect 814 677 815 681
rect 1434 677 1435 681
rect 1437 677 1438 681
rect 1450 677 1451 681
rect 1453 677 1454 681
rect 1466 677 1467 681
rect 1469 677 1470 681
rect 1485 677 1490 681
rect 1492 677 1495 681
rect 1497 677 1498 681
rect 1519 677 1521 681
rect 1523 677 1524 681
rect 1541 677 1542 681
rect 1544 677 1545 681
rect 1557 677 1562 681
rect 1564 677 1567 681
rect 1569 677 1570 681
rect 1584 677 1585 681
rect 1587 677 1588 681
rect 1632 677 1635 681
rect 1637 677 1640 681
rect 1642 677 1643 681
rect 1737 677 1740 681
rect 1742 677 1745 681
rect 1747 677 1748 681
rect 699 600 702 604
rect 704 600 707 604
rect 709 600 710 604
rect 756 604 757 608
rect 759 604 760 608
rect 780 600 783 604
rect 785 600 788 604
rect 790 600 791 604
rect 846 604 847 608
rect 849 604 850 608
rect 870 600 873 604
rect 875 600 878 604
rect 880 600 881 604
rect 729 596 730 600
rect 732 596 733 600
rect 501 591 502 595
rect 504 591 505 595
rect 517 591 518 595
rect 520 591 521 595
rect 533 591 534 595
rect 536 591 537 595
rect 552 591 557 595
rect 559 591 562 595
rect 564 591 565 595
rect 586 591 588 595
rect 590 591 591 595
rect 608 591 609 595
rect 611 591 612 595
rect 624 591 629 595
rect 631 591 634 595
rect 636 591 637 595
rect 651 591 652 595
rect 654 591 655 595
rect 810 596 811 600
rect 813 596 814 600
rect 900 596 901 600
rect 903 596 904 600
rect 1632 600 1635 604
rect 1637 600 1640 604
rect 1642 600 1643 604
rect 1689 604 1690 608
rect 1692 604 1693 608
rect 1713 600 1716 604
rect 1718 600 1721 604
rect 1723 600 1724 604
rect 1779 604 1780 608
rect 1782 604 1783 608
rect 1803 600 1806 604
rect 1808 600 1811 604
rect 1813 600 1814 604
rect 1662 596 1663 600
rect 1665 596 1666 600
rect 1434 591 1435 595
rect 1437 591 1438 595
rect 1450 591 1451 595
rect 1453 591 1454 595
rect 1466 591 1467 595
rect 1469 591 1470 595
rect 1485 591 1490 595
rect 1492 591 1495 595
rect 1497 591 1498 595
rect 1519 591 1521 595
rect 1523 591 1524 595
rect 1541 591 1542 595
rect 1544 591 1545 595
rect 1557 591 1562 595
rect 1564 591 1567 595
rect 1569 591 1570 595
rect 1584 591 1585 595
rect 1587 591 1588 595
rect 1743 596 1744 600
rect 1746 596 1747 600
rect 1833 596 1834 600
rect 1836 596 1837 600
rect 501 545 502 549
rect 504 545 505 549
rect 517 545 518 549
rect 520 545 521 549
rect 533 545 534 549
rect 536 545 537 549
rect 552 545 557 549
rect 559 545 562 549
rect 564 545 565 549
rect 586 545 588 549
rect 590 545 591 549
rect 608 545 609 549
rect 611 545 612 549
rect 624 545 629 549
rect 631 545 634 549
rect 636 545 637 549
rect 651 545 652 549
rect 654 545 655 549
rect 699 542 702 546
rect 704 542 707 546
rect 709 542 710 546
rect 780 542 783 546
rect 785 542 788 546
rect 790 542 791 546
rect 870 542 873 546
rect 875 542 878 546
rect 880 542 881 546
rect 1434 545 1435 549
rect 1437 545 1438 549
rect 1450 545 1451 549
rect 1453 545 1454 549
rect 1466 545 1467 549
rect 1469 545 1470 549
rect 1485 545 1490 549
rect 1492 545 1495 549
rect 1497 545 1498 549
rect 1519 545 1521 549
rect 1523 545 1524 549
rect 1541 545 1542 549
rect 1544 545 1545 549
rect 1557 545 1562 549
rect 1564 545 1567 549
rect 1569 545 1570 549
rect 1584 545 1585 549
rect 1587 545 1588 549
rect 1632 542 1635 546
rect 1637 542 1640 546
rect 1642 542 1643 546
rect 1713 542 1716 546
rect 1718 542 1721 546
rect 1723 542 1724 546
rect 1803 542 1806 546
rect 1808 542 1811 546
rect 1813 542 1814 546
rect 699 468 702 472
rect 704 468 707 472
rect 709 468 710 472
rect 729 464 730 468
rect 732 464 733 468
rect 501 459 502 463
rect 504 459 505 463
rect 517 459 518 463
rect 520 459 521 463
rect 533 459 534 463
rect 536 459 537 463
rect 552 459 557 463
rect 559 459 562 463
rect 564 459 565 463
rect 586 459 588 463
rect 590 459 591 463
rect 608 459 609 463
rect 611 459 612 463
rect 624 459 629 463
rect 631 459 634 463
rect 636 459 637 463
rect 651 459 652 463
rect 654 459 655 463
rect 1632 468 1635 472
rect 1637 468 1640 472
rect 1642 468 1643 472
rect 1662 464 1663 468
rect 1665 464 1666 468
rect 1434 459 1435 463
rect 1437 459 1438 463
rect 1450 459 1451 463
rect 1453 459 1454 463
rect 1466 459 1467 463
rect 1469 459 1470 463
rect 1485 459 1490 463
rect 1492 459 1495 463
rect 1497 459 1498 463
rect 1519 459 1521 463
rect 1523 459 1524 463
rect 1541 459 1542 463
rect 1544 459 1545 463
rect 1557 459 1562 463
rect 1564 459 1567 463
rect 1569 459 1570 463
rect 1584 459 1585 463
rect 1587 459 1588 463
rect 501 413 502 417
rect 504 413 505 417
rect 517 413 518 417
rect 520 413 521 417
rect 533 413 534 417
rect 536 413 537 417
rect 552 413 557 417
rect 559 413 562 417
rect 564 413 565 417
rect 586 413 588 417
rect 590 413 591 417
rect 608 413 609 417
rect 611 413 612 417
rect 624 413 629 417
rect 631 413 634 417
rect 636 413 637 417
rect 651 413 652 417
rect 654 413 655 417
rect 735 413 736 417
rect 738 413 739 417
rect 743 413 749 417
rect 753 413 754 417
rect 756 413 757 417
rect 778 413 779 417
rect 781 413 782 417
rect 794 413 795 417
rect 797 413 798 417
rect 813 413 818 417
rect 820 413 823 417
rect 825 413 826 417
rect 847 413 849 417
rect 851 413 852 417
rect 869 413 870 417
rect 872 413 873 417
rect 885 413 890 417
rect 892 413 895 417
rect 897 413 898 417
rect 912 413 913 417
rect 915 413 916 417
rect 24 399 25 403
rect 27 399 30 403
rect 32 399 33 403
rect 45 399 46 403
rect 48 399 49 403
rect 61 399 62 403
rect 64 399 67 403
rect 69 399 70 403
rect 87 399 88 403
rect 90 399 91 403
rect 103 399 104 403
rect 106 399 107 403
rect 119 399 120 403
rect 122 399 125 403
rect 127 399 128 403
rect 140 399 141 403
rect 143 399 144 403
rect 156 399 157 403
rect 159 399 162 403
rect 164 399 165 403
rect 177 399 178 403
rect 180 399 181 403
rect 193 399 194 403
rect 196 399 199 403
rect 201 399 202 403
rect 219 399 220 403
rect 222 399 223 403
rect 235 399 236 403
rect 238 399 239 403
rect 251 399 252 403
rect 254 399 257 403
rect 259 399 260 403
rect 272 399 273 403
rect 275 399 276 403
rect 288 399 289 403
rect 291 399 294 403
rect 296 399 297 403
rect 309 399 310 403
rect 312 399 313 403
rect 325 399 326 403
rect 328 399 331 403
rect 333 399 334 403
rect 351 399 352 403
rect 354 399 355 403
rect 367 399 368 403
rect 370 399 371 403
rect 383 399 384 403
rect 386 399 389 403
rect 391 399 392 403
rect 404 399 405 403
rect 407 399 408 403
rect 699 406 702 410
rect 704 406 707 410
rect 709 406 710 410
rect 1434 413 1435 417
rect 1437 413 1438 417
rect 1450 413 1451 417
rect 1453 413 1454 417
rect 1466 413 1467 417
rect 1469 413 1470 417
rect 1485 413 1490 417
rect 1492 413 1495 417
rect 1497 413 1498 417
rect 1519 413 1521 417
rect 1523 413 1524 417
rect 1541 413 1542 417
rect 1544 413 1545 417
rect 1557 413 1562 417
rect 1564 413 1567 417
rect 1569 413 1570 417
rect 1584 413 1585 417
rect 1587 413 1588 417
rect 1668 413 1669 417
rect 1671 413 1672 417
rect 1676 413 1682 417
rect 1686 413 1687 417
rect 1689 413 1690 417
rect 1711 413 1712 417
rect 1714 413 1715 417
rect 1727 413 1728 417
rect 1730 413 1731 417
rect 1746 413 1751 417
rect 1753 413 1756 417
rect 1758 413 1759 417
rect 1780 413 1782 417
rect 1784 413 1785 417
rect 1802 413 1803 417
rect 1805 413 1806 417
rect 1818 413 1823 417
rect 1825 413 1828 417
rect 1830 413 1831 417
rect 1845 413 1846 417
rect 1848 413 1849 417
rect 957 399 958 403
rect 960 399 963 403
rect 965 399 966 403
rect 978 399 979 403
rect 981 399 982 403
rect 994 399 995 403
rect 997 399 1000 403
rect 1002 399 1003 403
rect 1020 399 1021 403
rect 1023 399 1024 403
rect 1036 399 1037 403
rect 1039 399 1040 403
rect 1052 399 1053 403
rect 1055 399 1058 403
rect 1060 399 1061 403
rect 1073 399 1074 403
rect 1076 399 1077 403
rect 1089 399 1090 403
rect 1092 399 1095 403
rect 1097 399 1098 403
rect 1110 399 1111 403
rect 1113 399 1114 403
rect 1126 399 1127 403
rect 1129 399 1132 403
rect 1134 399 1135 403
rect 1152 399 1153 403
rect 1155 399 1156 403
rect 1168 399 1169 403
rect 1171 399 1172 403
rect 1184 399 1185 403
rect 1187 399 1190 403
rect 1192 399 1193 403
rect 1205 399 1206 403
rect 1208 399 1209 403
rect 1221 399 1222 403
rect 1224 399 1227 403
rect 1229 399 1230 403
rect 1242 399 1243 403
rect 1245 399 1246 403
rect 1258 399 1259 403
rect 1261 399 1264 403
rect 1266 399 1267 403
rect 1284 399 1285 403
rect 1287 399 1288 403
rect 1300 399 1301 403
rect 1303 399 1304 403
rect 1316 399 1317 403
rect 1319 399 1322 403
rect 1324 399 1325 403
rect 1337 399 1338 403
rect 1340 399 1341 403
rect 1632 406 1635 410
rect 1637 406 1640 410
rect 1642 406 1643 410
rect 139 355 140 359
rect 142 355 143 359
rect 163 355 164 359
rect 166 355 167 359
rect 925 359 929 360
rect 925 356 929 357
rect 1072 355 1073 359
rect 1075 355 1076 359
rect 1096 355 1097 359
rect 1099 355 1100 359
rect 1858 359 1862 360
rect 1858 356 1862 357
rect 159 344 160 348
rect 162 344 163 348
rect 1092 344 1093 348
rect 1095 344 1096 348
rect 151 332 155 333
rect 151 329 155 330
rect 1084 332 1088 333
rect 1084 329 1088 330
rect 139 321 140 325
rect 142 321 143 325
rect 163 321 164 325
rect 166 321 167 325
rect 1072 321 1073 325
rect 1075 321 1076 325
rect 1096 321 1097 325
rect 1099 321 1100 325
rect 795 289 796 293
rect 798 289 801 293
rect 803 289 804 293
rect 816 289 817 293
rect 819 289 820 293
rect 832 289 833 293
rect 835 289 838 293
rect 840 289 841 293
rect 858 289 859 293
rect 861 289 862 293
rect 874 289 875 293
rect 877 289 878 293
rect 890 289 891 293
rect 893 289 896 293
rect 898 289 899 293
rect 911 289 912 293
rect 914 289 915 293
rect 1728 289 1729 293
rect 1731 289 1734 293
rect 1736 289 1737 293
rect 1749 289 1750 293
rect 1752 289 1753 293
rect 1765 289 1766 293
rect 1768 289 1771 293
rect 1773 289 1774 293
rect 1791 289 1792 293
rect 1794 289 1795 293
rect 1807 289 1808 293
rect 1810 289 1811 293
rect 1823 289 1824 293
rect 1826 289 1829 293
rect 1831 289 1832 293
rect 1844 289 1845 293
rect 1847 289 1848 293
rect 24 259 25 263
rect 27 259 30 263
rect 32 259 33 263
rect 45 259 46 263
rect 48 259 49 263
rect 61 259 62 263
rect 64 259 67 263
rect 69 259 70 263
rect 87 259 88 263
rect 90 259 91 263
rect 103 259 104 263
rect 106 259 107 263
rect 119 259 120 263
rect 122 259 125 263
rect 127 259 128 263
rect 140 259 141 263
rect 143 259 144 263
rect 156 259 157 263
rect 159 259 162 263
rect 164 259 165 263
rect 177 259 178 263
rect 180 259 181 263
rect 193 259 194 263
rect 196 259 199 263
rect 201 259 202 263
rect 219 259 220 263
rect 222 259 223 263
rect 235 259 236 263
rect 238 259 239 263
rect 251 259 252 263
rect 254 259 257 263
rect 259 259 260 263
rect 272 259 273 263
rect 275 259 276 263
rect 288 259 289 263
rect 291 259 294 263
rect 296 259 297 263
rect 309 259 310 263
rect 312 259 313 263
rect 325 259 326 263
rect 328 259 331 263
rect 333 259 334 263
rect 351 259 352 263
rect 354 259 355 263
rect 367 259 368 263
rect 370 259 371 263
rect 383 259 384 263
rect 386 259 389 263
rect 391 259 392 263
rect 404 259 405 263
rect 407 259 408 263
rect 957 259 958 263
rect 960 259 963 263
rect 965 259 966 263
rect 978 259 979 263
rect 981 259 982 263
rect 994 259 995 263
rect 997 259 1000 263
rect 1002 259 1003 263
rect 1020 259 1021 263
rect 1023 259 1024 263
rect 1036 259 1037 263
rect 1039 259 1040 263
rect 1052 259 1053 263
rect 1055 259 1058 263
rect 1060 259 1061 263
rect 1073 259 1074 263
rect 1076 259 1077 263
rect 1089 259 1090 263
rect 1092 259 1095 263
rect 1097 259 1098 263
rect 1110 259 1111 263
rect 1113 259 1114 263
rect 1126 259 1127 263
rect 1129 259 1132 263
rect 1134 259 1135 263
rect 1152 259 1153 263
rect 1155 259 1156 263
rect 1168 259 1169 263
rect 1171 259 1172 263
rect 1184 259 1185 263
rect 1187 259 1190 263
rect 1192 259 1193 263
rect 1205 259 1206 263
rect 1208 259 1209 263
rect 1221 259 1222 263
rect 1224 259 1227 263
rect 1229 259 1230 263
rect 1242 259 1243 263
rect 1245 259 1246 263
rect 1258 259 1259 263
rect 1261 259 1264 263
rect 1266 259 1267 263
rect 1284 259 1285 263
rect 1287 259 1288 263
rect 1300 259 1301 263
rect 1303 259 1304 263
rect 1316 259 1317 263
rect 1319 259 1322 263
rect 1324 259 1325 263
rect 1337 259 1338 263
rect 1340 259 1341 263
rect 937 215 941 216
rect 937 212 941 213
rect 1870 215 1874 216
rect 1870 212 1874 213
rect 795 203 796 207
rect 798 203 801 207
rect 803 203 804 207
rect 816 203 817 207
rect 819 203 820 207
rect 832 203 833 207
rect 835 203 838 207
rect 840 203 841 207
rect 858 203 859 207
rect 861 203 862 207
rect 874 203 875 207
rect 877 203 878 207
rect 890 203 891 207
rect 893 203 896 207
rect 898 203 899 207
rect 911 203 912 207
rect 914 203 915 207
rect 1728 203 1729 207
rect 1731 203 1734 207
rect 1736 203 1737 207
rect 1749 203 1750 207
rect 1752 203 1753 207
rect 1765 203 1766 207
rect 1768 203 1771 207
rect 1773 203 1774 207
rect 1791 203 1792 207
rect 1794 203 1795 207
rect 1807 203 1808 207
rect 1810 203 1811 207
rect 1823 203 1824 207
rect 1826 203 1829 207
rect 1831 203 1832 207
rect 1844 203 1845 207
rect 1847 203 1848 207
rect 24 173 25 177
rect 27 173 30 177
rect 32 173 33 177
rect 45 173 46 177
rect 48 173 49 177
rect 61 173 62 177
rect 64 173 67 177
rect 69 173 70 177
rect 87 173 88 177
rect 90 173 91 177
rect 103 173 104 177
rect 106 173 107 177
rect 119 173 120 177
rect 122 173 125 177
rect 127 173 128 177
rect 140 173 141 177
rect 143 173 144 177
rect 156 173 157 177
rect 159 173 162 177
rect 164 173 165 177
rect 177 173 178 177
rect 180 173 181 177
rect 193 173 194 177
rect 196 173 199 177
rect 201 173 202 177
rect 219 173 220 177
rect 222 173 223 177
rect 235 173 236 177
rect 238 173 239 177
rect 251 173 252 177
rect 254 173 257 177
rect 259 173 260 177
rect 272 173 273 177
rect 275 173 276 177
rect 288 173 289 177
rect 291 173 294 177
rect 296 173 297 177
rect 309 173 310 177
rect 312 173 313 177
rect 325 173 326 177
rect 328 173 331 177
rect 333 173 334 177
rect 351 173 352 177
rect 354 173 355 177
rect 367 173 368 177
rect 370 173 371 177
rect 383 173 384 177
rect 386 173 389 177
rect 391 173 392 177
rect 404 173 405 177
rect 407 173 408 177
rect 957 173 958 177
rect 960 173 963 177
rect 965 173 966 177
rect 978 173 979 177
rect 981 173 982 177
rect 994 173 995 177
rect 997 173 1000 177
rect 1002 173 1003 177
rect 1020 173 1021 177
rect 1023 173 1024 177
rect 1036 173 1037 177
rect 1039 173 1040 177
rect 1052 173 1053 177
rect 1055 173 1058 177
rect 1060 173 1061 177
rect 1073 173 1074 177
rect 1076 173 1077 177
rect 1089 173 1090 177
rect 1092 173 1095 177
rect 1097 173 1098 177
rect 1110 173 1111 177
rect 1113 173 1114 177
rect 1126 173 1127 177
rect 1129 173 1132 177
rect 1134 173 1135 177
rect 1152 173 1153 177
rect 1155 173 1156 177
rect 1168 173 1169 177
rect 1171 173 1172 177
rect 1184 173 1185 177
rect 1187 173 1190 177
rect 1192 173 1193 177
rect 1205 173 1206 177
rect 1208 173 1209 177
rect 1221 173 1222 177
rect 1224 173 1227 177
rect 1229 173 1230 177
rect 1242 173 1243 177
rect 1245 173 1246 177
rect 1258 173 1259 177
rect 1261 173 1264 177
rect 1266 173 1267 177
rect 1284 173 1285 177
rect 1287 173 1288 177
rect 1300 173 1301 177
rect 1303 173 1304 177
rect 1316 173 1317 177
rect 1319 173 1322 177
rect 1324 173 1325 177
rect 1337 173 1338 177
rect 1340 173 1341 177
rect 256 129 257 133
rect 259 129 260 133
rect 280 129 281 133
rect 283 129 284 133
rect 1189 129 1190 133
rect 1192 129 1193 133
rect 1213 129 1214 133
rect 1216 129 1217 133
rect 276 118 277 122
rect 279 118 280 122
rect 1209 118 1210 122
rect 1212 118 1213 122
rect 268 106 272 107
rect 268 103 272 104
rect 1201 106 1205 107
rect 1201 103 1205 104
rect 256 95 257 99
rect 259 95 260 99
rect 280 95 281 99
rect 283 95 284 99
rect 1189 95 1190 99
rect 1192 95 1193 99
rect 1213 95 1214 99
rect 1216 95 1217 99
rect 24 33 25 37
rect 27 33 30 37
rect 32 33 33 37
rect 45 33 46 37
rect 48 33 49 37
rect 61 33 62 37
rect 64 33 67 37
rect 69 33 70 37
rect 87 33 88 37
rect 90 33 91 37
rect 103 33 104 37
rect 106 33 107 37
rect 119 33 120 37
rect 122 33 125 37
rect 127 33 128 37
rect 140 33 141 37
rect 143 33 144 37
rect 156 33 157 37
rect 159 33 162 37
rect 164 33 165 37
rect 177 33 178 37
rect 180 33 181 37
rect 193 33 194 37
rect 196 33 199 37
rect 201 33 202 37
rect 219 33 220 37
rect 222 33 223 37
rect 235 33 236 37
rect 238 33 239 37
rect 251 33 252 37
rect 254 33 257 37
rect 259 33 260 37
rect 272 33 273 37
rect 275 33 276 37
rect 288 33 289 37
rect 291 33 294 37
rect 296 33 297 37
rect 309 33 310 37
rect 312 33 313 37
rect 325 33 326 37
rect 328 33 331 37
rect 333 33 334 37
rect 351 33 352 37
rect 354 33 355 37
rect 367 33 368 37
rect 370 33 371 37
rect 383 33 384 37
rect 386 33 389 37
rect 391 33 392 37
rect 404 33 405 37
rect 407 33 408 37
rect 957 33 958 37
rect 960 33 963 37
rect 965 33 966 37
rect 978 33 979 37
rect 981 33 982 37
rect 994 33 995 37
rect 997 33 1000 37
rect 1002 33 1003 37
rect 1020 33 1021 37
rect 1023 33 1024 37
rect 1036 33 1037 37
rect 1039 33 1040 37
rect 1052 33 1053 37
rect 1055 33 1058 37
rect 1060 33 1061 37
rect 1073 33 1074 37
rect 1076 33 1077 37
rect 1089 33 1090 37
rect 1092 33 1095 37
rect 1097 33 1098 37
rect 1110 33 1111 37
rect 1113 33 1114 37
rect 1126 33 1127 37
rect 1129 33 1132 37
rect 1134 33 1135 37
rect 1152 33 1153 37
rect 1155 33 1156 37
rect 1168 33 1169 37
rect 1171 33 1172 37
rect 1184 33 1185 37
rect 1187 33 1190 37
rect 1192 33 1193 37
rect 1205 33 1206 37
rect 1208 33 1209 37
rect 1221 33 1222 37
rect 1224 33 1227 37
rect 1229 33 1230 37
rect 1242 33 1243 37
rect 1245 33 1246 37
rect 1258 33 1259 37
rect 1261 33 1264 37
rect 1266 33 1267 37
rect 1284 33 1285 37
rect 1287 33 1288 37
rect 1300 33 1301 37
rect 1303 33 1304 37
rect 1316 33 1317 37
rect 1319 33 1322 37
rect 1324 33 1325 37
rect 1337 33 1338 37
rect 1340 33 1341 37
<< pdiffusion >>
rect 496 1937 497 1945
rect 499 1937 502 1945
rect 504 1937 505 1945
rect 517 1937 518 1945
rect 520 1941 521 1945
rect 520 1937 525 1941
rect 533 1937 534 1945
rect 536 1937 539 1945
rect 541 1937 542 1945
rect 559 1937 560 1945
rect 562 1937 563 1945
rect 575 1937 576 1945
rect 578 1941 579 1945
rect 578 1937 583 1941
rect 591 1937 592 1945
rect 594 1937 597 1945
rect 599 1937 600 1945
rect 612 1937 613 1945
rect 615 1937 616 1945
rect 628 1937 629 1945
rect 631 1937 634 1945
rect 636 1937 637 1945
rect 649 1937 650 1945
rect 652 1941 653 1945
rect 652 1937 657 1941
rect 665 1937 666 1945
rect 668 1937 671 1945
rect 673 1937 674 1945
rect 691 1937 692 1945
rect 694 1937 695 1945
rect 707 1937 708 1945
rect 710 1941 711 1945
rect 710 1937 715 1941
rect 723 1937 724 1945
rect 726 1937 729 1945
rect 731 1937 732 1945
rect 744 1937 745 1945
rect 747 1937 748 1945
rect 760 1937 761 1945
rect 763 1937 766 1945
rect 768 1937 769 1945
rect 781 1937 782 1945
rect 784 1941 785 1945
rect 784 1937 789 1941
rect 797 1937 798 1945
rect 800 1937 803 1945
rect 805 1937 806 1945
rect 823 1937 824 1945
rect 826 1937 827 1945
rect 839 1937 840 1945
rect 842 1941 843 1945
rect 842 1937 847 1941
rect 855 1937 856 1945
rect 858 1937 861 1945
rect 863 1937 864 1945
rect 876 1937 877 1945
rect 879 1937 880 1945
rect 892 1937 893 1945
rect 895 1937 898 1945
rect 900 1937 901 1945
rect 913 1937 914 1945
rect 916 1941 917 1945
rect 916 1937 921 1941
rect 929 1937 930 1945
rect 932 1937 935 1945
rect 937 1937 938 1945
rect 955 1937 956 1945
rect 958 1937 959 1945
rect 971 1937 972 1945
rect 974 1941 975 1945
rect 974 1937 979 1941
rect 987 1937 988 1945
rect 990 1937 993 1945
rect 995 1937 996 1945
rect 1008 1937 1009 1945
rect 1011 1937 1012 1945
rect 1429 1937 1430 1945
rect 1432 1937 1435 1945
rect 1437 1937 1438 1945
rect 1450 1937 1451 1945
rect 1453 1941 1454 1945
rect 1453 1937 1458 1941
rect 1466 1937 1467 1945
rect 1469 1937 1472 1945
rect 1474 1937 1475 1945
rect 1492 1937 1493 1945
rect 1495 1937 1496 1945
rect 1508 1937 1509 1945
rect 1511 1941 1512 1945
rect 1511 1937 1516 1941
rect 1524 1937 1525 1945
rect 1527 1937 1530 1945
rect 1532 1937 1533 1945
rect 1545 1937 1546 1945
rect 1548 1937 1549 1945
rect 1561 1937 1562 1945
rect 1564 1937 1567 1945
rect 1569 1937 1570 1945
rect 1582 1937 1583 1945
rect 1585 1941 1586 1945
rect 1585 1937 1590 1941
rect 1598 1937 1599 1945
rect 1601 1937 1604 1945
rect 1606 1937 1607 1945
rect 1624 1937 1625 1945
rect 1627 1937 1628 1945
rect 1640 1937 1641 1945
rect 1643 1941 1644 1945
rect 1643 1937 1648 1941
rect 1656 1937 1657 1945
rect 1659 1937 1662 1945
rect 1664 1937 1665 1945
rect 1677 1937 1678 1945
rect 1680 1937 1681 1945
rect 1693 1937 1694 1945
rect 1696 1937 1699 1945
rect 1701 1937 1702 1945
rect 1714 1937 1715 1945
rect 1717 1941 1718 1945
rect 1717 1937 1722 1941
rect 1730 1937 1731 1945
rect 1733 1937 1736 1945
rect 1738 1937 1739 1945
rect 1756 1937 1757 1945
rect 1759 1937 1760 1945
rect 1772 1937 1773 1945
rect 1775 1941 1776 1945
rect 1775 1937 1780 1941
rect 1788 1937 1789 1945
rect 1791 1937 1794 1945
rect 1796 1937 1797 1945
rect 1809 1937 1810 1945
rect 1812 1937 1813 1945
rect 1825 1937 1826 1945
rect 1828 1937 1831 1945
rect 1833 1937 1834 1945
rect 1846 1937 1847 1945
rect 1849 1941 1850 1945
rect 1849 1937 1854 1941
rect 1862 1937 1863 1945
rect 1865 1937 1868 1945
rect 1870 1937 1871 1945
rect 1888 1937 1889 1945
rect 1891 1937 1892 1945
rect 1904 1937 1905 1945
rect 1907 1941 1908 1945
rect 1907 1937 1912 1941
rect 1920 1937 1921 1945
rect 1923 1937 1926 1945
rect 1928 1937 1929 1945
rect 1941 1937 1942 1945
rect 1944 1937 1945 1945
rect 156 1904 157 1912
rect 159 1904 162 1912
rect 164 1904 165 1912
rect 177 1904 178 1912
rect 180 1908 181 1912
rect 180 1904 185 1908
rect 193 1904 194 1912
rect 196 1904 199 1912
rect 201 1904 202 1912
rect 219 1904 220 1912
rect 222 1904 223 1912
rect 235 1904 236 1912
rect 238 1908 239 1912
rect 238 1904 243 1908
rect 251 1904 252 1912
rect 254 1904 257 1912
rect 259 1904 260 1912
rect 272 1904 273 1912
rect 275 1904 276 1912
rect 1089 1904 1090 1912
rect 1092 1904 1095 1912
rect 1097 1904 1098 1912
rect 1110 1904 1111 1912
rect 1113 1908 1114 1912
rect 1113 1904 1118 1908
rect 1126 1904 1127 1912
rect 1129 1904 1132 1912
rect 1134 1904 1135 1912
rect 1152 1904 1153 1912
rect 1155 1904 1156 1912
rect 1168 1904 1169 1912
rect 1171 1908 1172 1912
rect 1171 1904 1176 1908
rect 1184 1904 1185 1912
rect 1187 1904 1190 1912
rect 1192 1904 1193 1912
rect 1205 1904 1206 1912
rect 1208 1904 1209 1912
rect 675 1866 676 1874
rect 678 1866 679 1874
rect 501 1853 502 1861
rect 504 1853 505 1861
rect 517 1853 518 1861
rect 520 1853 521 1861
rect 533 1853 534 1861
rect 536 1853 537 1861
rect 552 1853 557 1861
rect 559 1853 562 1861
rect 564 1853 565 1861
rect 586 1853 588 1861
rect 590 1853 591 1861
rect 608 1853 609 1861
rect 611 1853 612 1861
rect 624 1853 629 1861
rect 631 1853 634 1861
rect 636 1853 637 1861
rect 651 1853 652 1861
rect 654 1853 655 1861
rect 699 1860 702 1868
rect 704 1860 707 1868
rect 709 1860 710 1868
rect 729 1866 730 1874
rect 732 1866 733 1874
rect 756 1866 757 1874
rect 759 1866 760 1874
rect 780 1860 783 1868
rect 785 1860 788 1868
rect 790 1860 791 1868
rect 810 1866 811 1874
rect 813 1866 814 1874
rect 1608 1866 1609 1874
rect 1611 1866 1612 1874
rect 1434 1853 1435 1861
rect 1437 1853 1438 1861
rect 1450 1853 1451 1861
rect 1453 1853 1454 1861
rect 1466 1853 1467 1861
rect 1469 1853 1470 1861
rect 1485 1853 1490 1861
rect 1492 1853 1495 1861
rect 1497 1853 1498 1861
rect 1519 1853 1521 1861
rect 1523 1853 1524 1861
rect 1541 1853 1542 1861
rect 1544 1853 1545 1861
rect 1557 1853 1562 1861
rect 1564 1853 1567 1861
rect 1569 1853 1570 1861
rect 1584 1853 1585 1861
rect 1587 1853 1588 1861
rect 1632 1860 1635 1868
rect 1637 1860 1640 1868
rect 1642 1860 1643 1868
rect 1662 1866 1663 1874
rect 1665 1866 1666 1874
rect 1689 1866 1690 1874
rect 1692 1866 1693 1874
rect 1713 1860 1716 1868
rect 1718 1860 1721 1868
rect 1723 1860 1724 1868
rect 1743 1866 1744 1874
rect 1746 1866 1747 1874
rect 147 1802 148 1810
rect 150 1802 151 1810
rect 163 1802 164 1810
rect 166 1802 169 1810
rect 171 1802 172 1810
rect 184 1806 185 1810
rect 180 1802 185 1806
rect 187 1802 188 1810
rect 200 1802 201 1810
rect 203 1802 204 1810
rect 221 1802 222 1810
rect 224 1802 227 1810
rect 229 1802 230 1810
rect 242 1806 243 1810
rect 238 1802 243 1806
rect 245 1802 246 1810
rect 258 1802 259 1810
rect 261 1802 264 1810
rect 266 1802 267 1810
rect 1080 1802 1081 1810
rect 1083 1802 1084 1810
rect 1096 1802 1097 1810
rect 1099 1802 1102 1810
rect 1104 1802 1105 1810
rect 1117 1806 1118 1810
rect 1113 1802 1118 1806
rect 1120 1802 1121 1810
rect 1133 1802 1134 1810
rect 1136 1802 1137 1810
rect 1154 1802 1155 1810
rect 1157 1802 1160 1810
rect 1162 1802 1163 1810
rect 1175 1806 1176 1810
rect 1171 1802 1176 1806
rect 1178 1802 1179 1810
rect 1191 1802 1192 1810
rect 1194 1802 1197 1810
rect 1199 1802 1200 1810
rect 501 1767 502 1775
rect 504 1767 505 1775
rect 517 1767 518 1775
rect 520 1767 521 1775
rect 533 1767 534 1775
rect 536 1767 537 1775
rect 552 1767 557 1775
rect 559 1767 562 1775
rect 564 1767 565 1775
rect 586 1767 588 1775
rect 590 1767 591 1775
rect 608 1767 609 1775
rect 611 1767 612 1775
rect 624 1767 629 1775
rect 631 1767 634 1775
rect 636 1767 637 1775
rect 651 1767 652 1775
rect 654 1767 655 1775
rect 699 1768 702 1776
rect 704 1768 707 1776
rect 709 1768 710 1776
rect 780 1768 783 1776
rect 785 1768 788 1776
rect 790 1768 791 1776
rect 1434 1767 1435 1775
rect 1437 1767 1438 1775
rect 1450 1767 1451 1775
rect 1453 1767 1454 1775
rect 1466 1767 1467 1775
rect 1469 1767 1470 1775
rect 1485 1767 1490 1775
rect 1492 1767 1495 1775
rect 1497 1767 1498 1775
rect 1519 1767 1521 1775
rect 1523 1767 1524 1775
rect 1541 1767 1542 1775
rect 1544 1767 1545 1775
rect 1557 1767 1562 1775
rect 1564 1767 1567 1775
rect 1569 1767 1570 1775
rect 1584 1767 1585 1775
rect 1587 1767 1588 1775
rect 1632 1768 1635 1776
rect 1637 1768 1640 1776
rect 1642 1768 1643 1776
rect 1713 1768 1716 1776
rect 1718 1768 1721 1776
rect 1723 1768 1724 1776
rect 501 1721 502 1729
rect 504 1721 505 1729
rect 517 1721 518 1729
rect 520 1721 521 1729
rect 533 1721 534 1729
rect 536 1721 537 1729
rect 552 1721 557 1729
rect 559 1721 562 1729
rect 564 1721 565 1729
rect 586 1721 588 1729
rect 590 1721 591 1729
rect 608 1721 609 1729
rect 611 1721 612 1729
rect 624 1721 629 1729
rect 631 1721 634 1729
rect 636 1721 637 1729
rect 651 1721 652 1729
rect 654 1721 655 1729
rect 699 1728 702 1736
rect 704 1728 707 1736
rect 709 1728 710 1736
rect 729 1734 730 1742
rect 732 1734 733 1742
rect 780 1734 781 1742
rect 783 1734 784 1742
rect 804 1728 807 1736
rect 809 1728 812 1736
rect 814 1728 815 1736
rect 834 1734 835 1742
rect 837 1734 838 1742
rect 1434 1721 1435 1729
rect 1437 1721 1438 1729
rect 1450 1721 1451 1729
rect 1453 1721 1454 1729
rect 1466 1721 1467 1729
rect 1469 1721 1470 1729
rect 1485 1721 1490 1729
rect 1492 1721 1495 1729
rect 1497 1721 1498 1729
rect 1519 1721 1521 1729
rect 1523 1721 1524 1729
rect 1541 1721 1542 1729
rect 1544 1721 1545 1729
rect 1557 1721 1562 1729
rect 1564 1721 1567 1729
rect 1569 1721 1570 1729
rect 1584 1721 1585 1729
rect 1587 1721 1588 1729
rect 1632 1728 1635 1736
rect 1637 1728 1640 1736
rect 1642 1728 1643 1736
rect 1662 1734 1663 1742
rect 1665 1734 1666 1742
rect 1713 1734 1714 1742
rect 1716 1734 1717 1742
rect 1737 1728 1740 1736
rect 1742 1728 1745 1736
rect 1747 1728 1748 1736
rect 1767 1734 1768 1742
rect 1770 1734 1771 1742
rect 501 1635 502 1643
rect 504 1635 505 1643
rect 517 1635 518 1643
rect 520 1635 521 1643
rect 533 1635 534 1643
rect 536 1635 537 1643
rect 552 1635 557 1643
rect 559 1635 562 1643
rect 564 1635 565 1643
rect 586 1635 588 1643
rect 590 1635 591 1643
rect 608 1635 609 1643
rect 611 1635 612 1643
rect 624 1635 629 1643
rect 631 1635 634 1643
rect 636 1635 637 1643
rect 651 1635 652 1643
rect 654 1635 655 1643
rect 699 1637 702 1645
rect 704 1637 707 1645
rect 709 1637 710 1645
rect 804 1637 807 1645
rect 809 1637 812 1645
rect 814 1637 815 1645
rect 1434 1635 1435 1643
rect 1437 1635 1438 1643
rect 1450 1635 1451 1643
rect 1453 1635 1454 1643
rect 1466 1635 1467 1643
rect 1469 1635 1470 1643
rect 1485 1635 1490 1643
rect 1492 1635 1495 1643
rect 1497 1635 1498 1643
rect 1519 1635 1521 1643
rect 1523 1635 1524 1643
rect 1541 1635 1542 1643
rect 1544 1635 1545 1643
rect 1557 1635 1562 1643
rect 1564 1635 1567 1643
rect 1569 1635 1570 1643
rect 1584 1635 1585 1643
rect 1587 1635 1588 1643
rect 1632 1637 1635 1645
rect 1637 1637 1640 1645
rect 1642 1637 1643 1645
rect 1737 1637 1740 1645
rect 1742 1637 1745 1645
rect 1747 1637 1748 1645
rect 501 1589 502 1597
rect 504 1589 505 1597
rect 517 1589 518 1597
rect 520 1589 521 1597
rect 533 1589 534 1597
rect 536 1589 537 1597
rect 552 1589 557 1597
rect 559 1589 562 1597
rect 564 1589 565 1597
rect 586 1589 588 1597
rect 590 1589 591 1597
rect 608 1589 609 1597
rect 611 1589 612 1597
rect 624 1589 629 1597
rect 631 1589 634 1597
rect 636 1589 637 1597
rect 651 1589 652 1597
rect 654 1589 655 1597
rect 699 1596 702 1604
rect 704 1596 707 1604
rect 709 1596 710 1604
rect 729 1602 730 1610
rect 732 1602 733 1610
rect 756 1602 757 1610
rect 759 1602 760 1610
rect 780 1596 783 1604
rect 785 1596 788 1604
rect 790 1596 791 1604
rect 810 1602 811 1610
rect 813 1602 814 1610
rect 846 1602 847 1610
rect 849 1602 850 1610
rect 870 1596 873 1604
rect 875 1596 878 1604
rect 880 1596 881 1604
rect 900 1602 901 1610
rect 903 1602 904 1610
rect 1434 1589 1435 1597
rect 1437 1589 1438 1597
rect 1450 1589 1451 1597
rect 1453 1589 1454 1597
rect 1466 1589 1467 1597
rect 1469 1589 1470 1597
rect 1485 1589 1490 1597
rect 1492 1589 1495 1597
rect 1497 1589 1498 1597
rect 1519 1589 1521 1597
rect 1523 1589 1524 1597
rect 1541 1589 1542 1597
rect 1544 1589 1545 1597
rect 1557 1589 1562 1597
rect 1564 1589 1567 1597
rect 1569 1589 1570 1597
rect 1584 1589 1585 1597
rect 1587 1589 1588 1597
rect 1632 1596 1635 1604
rect 1637 1596 1640 1604
rect 1642 1596 1643 1604
rect 1662 1602 1663 1610
rect 1665 1602 1666 1610
rect 1689 1602 1690 1610
rect 1692 1602 1693 1610
rect 1713 1596 1716 1604
rect 1718 1596 1721 1604
rect 1723 1596 1724 1604
rect 1743 1602 1744 1610
rect 1746 1602 1747 1610
rect 1779 1602 1780 1610
rect 1782 1602 1783 1610
rect 1803 1596 1806 1604
rect 1808 1596 1811 1604
rect 1813 1596 1814 1604
rect 1833 1602 1834 1610
rect 1836 1602 1837 1610
rect 501 1503 502 1511
rect 504 1503 505 1511
rect 517 1503 518 1511
rect 520 1503 521 1511
rect 533 1503 534 1511
rect 536 1503 537 1511
rect 552 1503 557 1511
rect 559 1503 562 1511
rect 564 1503 565 1511
rect 586 1503 588 1511
rect 590 1503 591 1511
rect 608 1503 609 1511
rect 611 1503 612 1511
rect 624 1503 629 1511
rect 631 1503 634 1511
rect 636 1503 637 1511
rect 651 1503 652 1511
rect 654 1503 655 1511
rect 699 1502 702 1510
rect 704 1502 707 1510
rect 709 1502 710 1510
rect 780 1502 783 1510
rect 785 1502 788 1510
rect 790 1502 791 1510
rect 870 1502 873 1510
rect 875 1502 878 1510
rect 880 1502 881 1510
rect 1434 1503 1435 1511
rect 1437 1503 1438 1511
rect 1450 1503 1451 1511
rect 1453 1503 1454 1511
rect 1466 1503 1467 1511
rect 1469 1503 1470 1511
rect 1485 1503 1490 1511
rect 1492 1503 1495 1511
rect 1497 1503 1498 1511
rect 1519 1503 1521 1511
rect 1523 1503 1524 1511
rect 1541 1503 1542 1511
rect 1544 1503 1545 1511
rect 1557 1503 1562 1511
rect 1564 1503 1567 1511
rect 1569 1503 1570 1511
rect 1584 1503 1585 1511
rect 1587 1503 1588 1511
rect 1632 1502 1635 1510
rect 1637 1502 1640 1510
rect 1642 1502 1643 1510
rect 1713 1502 1716 1510
rect 1718 1502 1721 1510
rect 1723 1502 1724 1510
rect 1803 1502 1806 1510
rect 1808 1502 1811 1510
rect 1813 1502 1814 1510
rect 501 1457 502 1465
rect 504 1457 505 1465
rect 517 1457 518 1465
rect 520 1457 521 1465
rect 533 1457 534 1465
rect 536 1457 537 1465
rect 552 1457 557 1465
rect 559 1457 562 1465
rect 564 1457 565 1465
rect 586 1457 588 1465
rect 590 1457 591 1465
rect 608 1457 609 1465
rect 611 1457 612 1465
rect 624 1457 629 1465
rect 631 1457 634 1465
rect 636 1457 637 1465
rect 651 1457 652 1465
rect 654 1457 655 1465
rect 699 1464 702 1472
rect 704 1464 707 1472
rect 709 1464 710 1472
rect 729 1470 730 1478
rect 732 1470 733 1478
rect 1434 1457 1435 1465
rect 1437 1457 1438 1465
rect 1450 1457 1451 1465
rect 1453 1457 1454 1465
rect 1466 1457 1467 1465
rect 1469 1457 1470 1465
rect 1485 1457 1490 1465
rect 1492 1457 1495 1465
rect 1497 1457 1498 1465
rect 1519 1457 1521 1465
rect 1523 1457 1524 1465
rect 1541 1457 1542 1465
rect 1544 1457 1545 1465
rect 1557 1457 1562 1465
rect 1564 1457 1567 1465
rect 1569 1457 1570 1465
rect 1584 1457 1585 1465
rect 1587 1457 1588 1465
rect 1632 1464 1635 1472
rect 1637 1464 1640 1472
rect 1642 1464 1643 1472
rect 1662 1470 1663 1478
rect 1665 1470 1666 1478
rect 24 1402 25 1410
rect 27 1402 30 1410
rect 32 1402 33 1410
rect 45 1402 46 1410
rect 48 1406 49 1410
rect 48 1402 53 1406
rect 61 1402 62 1410
rect 64 1402 67 1410
rect 69 1402 70 1410
rect 87 1402 88 1410
rect 90 1402 91 1410
rect 103 1402 104 1410
rect 106 1406 107 1410
rect 106 1402 111 1406
rect 119 1402 120 1410
rect 122 1402 125 1410
rect 127 1402 128 1410
rect 140 1402 141 1410
rect 143 1402 144 1410
rect 156 1402 157 1410
rect 159 1402 162 1410
rect 164 1402 165 1410
rect 177 1402 178 1410
rect 180 1406 181 1410
rect 180 1402 185 1406
rect 193 1402 194 1410
rect 196 1402 199 1410
rect 201 1402 202 1410
rect 219 1402 220 1410
rect 222 1402 223 1410
rect 235 1402 236 1410
rect 238 1406 239 1410
rect 238 1402 243 1406
rect 251 1402 252 1410
rect 254 1402 257 1410
rect 259 1402 260 1410
rect 272 1402 273 1410
rect 275 1402 276 1410
rect 288 1402 289 1410
rect 291 1402 294 1410
rect 296 1402 297 1410
rect 309 1402 310 1410
rect 312 1406 313 1410
rect 312 1402 317 1406
rect 325 1402 326 1410
rect 328 1402 331 1410
rect 333 1402 334 1410
rect 351 1402 352 1410
rect 354 1402 355 1410
rect 367 1402 368 1410
rect 370 1406 371 1410
rect 370 1402 375 1406
rect 383 1402 384 1410
rect 386 1402 389 1410
rect 391 1402 392 1410
rect 404 1402 405 1410
rect 407 1402 408 1410
rect 957 1402 958 1410
rect 960 1402 963 1410
rect 965 1402 966 1410
rect 978 1402 979 1410
rect 981 1406 982 1410
rect 981 1402 986 1406
rect 994 1402 995 1410
rect 997 1402 1000 1410
rect 1002 1402 1003 1410
rect 1020 1402 1021 1410
rect 1023 1402 1024 1410
rect 1036 1402 1037 1410
rect 1039 1406 1040 1410
rect 1039 1402 1044 1406
rect 1052 1402 1053 1410
rect 1055 1402 1058 1410
rect 1060 1402 1061 1410
rect 1073 1402 1074 1410
rect 1076 1402 1077 1410
rect 1089 1402 1090 1410
rect 1092 1402 1095 1410
rect 1097 1402 1098 1410
rect 1110 1402 1111 1410
rect 1113 1406 1114 1410
rect 1113 1402 1118 1406
rect 1126 1402 1127 1410
rect 1129 1402 1132 1410
rect 1134 1402 1135 1410
rect 1152 1402 1153 1410
rect 1155 1402 1156 1410
rect 1168 1402 1169 1410
rect 1171 1406 1172 1410
rect 1171 1402 1176 1406
rect 1184 1402 1185 1410
rect 1187 1402 1190 1410
rect 1192 1402 1193 1410
rect 1205 1402 1206 1410
rect 1208 1402 1209 1410
rect 1221 1402 1222 1410
rect 1224 1402 1227 1410
rect 1229 1402 1230 1410
rect 1242 1402 1243 1410
rect 1245 1406 1246 1410
rect 1245 1402 1250 1406
rect 1258 1402 1259 1410
rect 1261 1402 1264 1410
rect 1266 1402 1267 1410
rect 1284 1402 1285 1410
rect 1287 1402 1288 1410
rect 1300 1402 1301 1410
rect 1303 1406 1304 1410
rect 1303 1402 1308 1406
rect 1316 1402 1317 1410
rect 1319 1402 1322 1410
rect 1324 1402 1325 1410
rect 1337 1402 1338 1410
rect 1340 1402 1341 1410
rect 501 1371 502 1379
rect 504 1371 505 1379
rect 517 1371 518 1379
rect 520 1371 521 1379
rect 533 1371 534 1379
rect 536 1371 537 1379
rect 552 1371 557 1379
rect 559 1371 562 1379
rect 564 1371 565 1379
rect 586 1371 588 1379
rect 590 1371 591 1379
rect 608 1371 609 1379
rect 611 1371 612 1379
rect 624 1371 629 1379
rect 631 1371 634 1379
rect 636 1371 637 1379
rect 651 1371 652 1379
rect 654 1371 655 1379
rect 699 1366 702 1374
rect 704 1366 707 1374
rect 709 1366 710 1374
rect 735 1371 736 1379
rect 738 1371 739 1379
rect 743 1371 749 1379
rect 753 1371 754 1379
rect 756 1371 757 1379
rect 778 1371 779 1379
rect 781 1371 782 1379
rect 794 1371 795 1379
rect 797 1371 798 1379
rect 813 1371 818 1379
rect 820 1371 823 1379
rect 825 1371 826 1379
rect 847 1371 849 1379
rect 851 1371 852 1379
rect 869 1371 870 1379
rect 872 1371 873 1379
rect 885 1371 890 1379
rect 892 1371 895 1379
rect 897 1371 898 1379
rect 912 1371 913 1379
rect 915 1371 916 1379
rect 1434 1371 1435 1379
rect 1437 1371 1438 1379
rect 1450 1371 1451 1379
rect 1453 1371 1454 1379
rect 1466 1371 1467 1379
rect 1469 1371 1470 1379
rect 1485 1371 1490 1379
rect 1492 1371 1495 1379
rect 1497 1371 1498 1379
rect 1519 1371 1521 1379
rect 1523 1371 1524 1379
rect 1541 1371 1542 1379
rect 1544 1371 1545 1379
rect 1557 1371 1562 1379
rect 1564 1371 1567 1379
rect 1569 1371 1570 1379
rect 1584 1371 1585 1379
rect 1587 1371 1588 1379
rect 1632 1366 1635 1374
rect 1637 1366 1640 1374
rect 1642 1366 1643 1374
rect 1668 1371 1669 1379
rect 1671 1371 1672 1379
rect 1676 1371 1682 1379
rect 1686 1371 1687 1379
rect 1689 1371 1690 1379
rect 1711 1371 1712 1379
rect 1714 1371 1715 1379
rect 1727 1371 1728 1379
rect 1730 1371 1731 1379
rect 1746 1371 1751 1379
rect 1753 1371 1756 1379
rect 1758 1371 1759 1379
rect 1780 1371 1782 1379
rect 1784 1371 1785 1379
rect 1802 1371 1803 1379
rect 1805 1371 1806 1379
rect 1818 1371 1823 1379
rect 1825 1371 1828 1379
rect 1830 1371 1831 1379
rect 1845 1371 1846 1379
rect 1848 1371 1849 1379
rect 795 1292 796 1300
rect 798 1292 801 1300
rect 803 1292 804 1300
rect 816 1292 817 1300
rect 819 1296 820 1300
rect 819 1292 824 1296
rect 832 1292 833 1300
rect 835 1292 838 1300
rect 840 1292 841 1300
rect 858 1292 859 1300
rect 861 1292 862 1300
rect 874 1292 875 1300
rect 877 1296 878 1300
rect 877 1292 882 1296
rect 890 1292 891 1300
rect 893 1292 896 1300
rect 898 1292 899 1300
rect 911 1292 912 1300
rect 914 1292 915 1300
rect 1728 1292 1729 1300
rect 1731 1292 1734 1300
rect 1736 1292 1737 1300
rect 1749 1292 1750 1300
rect 1752 1296 1753 1300
rect 1752 1292 1757 1296
rect 1765 1292 1766 1300
rect 1768 1292 1771 1300
rect 1773 1292 1774 1300
rect 1791 1292 1792 1300
rect 1794 1292 1795 1300
rect 1807 1292 1808 1300
rect 1810 1296 1811 1300
rect 1810 1292 1815 1296
rect 1823 1292 1824 1300
rect 1826 1292 1829 1300
rect 1831 1292 1832 1300
rect 1844 1292 1845 1300
rect 1847 1292 1848 1300
rect 24 1262 25 1270
rect 27 1262 30 1270
rect 32 1262 33 1270
rect 45 1262 46 1270
rect 48 1266 49 1270
rect 48 1262 53 1266
rect 61 1262 62 1270
rect 64 1262 67 1270
rect 69 1262 70 1270
rect 87 1262 88 1270
rect 90 1262 91 1270
rect 103 1262 104 1270
rect 106 1266 107 1270
rect 106 1262 111 1266
rect 119 1262 120 1270
rect 122 1262 125 1270
rect 127 1262 128 1270
rect 140 1262 141 1270
rect 143 1262 144 1270
rect 156 1262 157 1270
rect 159 1262 162 1270
rect 164 1262 165 1270
rect 177 1262 178 1270
rect 180 1266 181 1270
rect 180 1262 185 1266
rect 193 1262 194 1270
rect 196 1262 199 1270
rect 201 1262 202 1270
rect 219 1262 220 1270
rect 222 1262 223 1270
rect 235 1262 236 1270
rect 238 1266 239 1270
rect 238 1262 243 1266
rect 251 1262 252 1270
rect 254 1262 257 1270
rect 259 1262 260 1270
rect 272 1262 273 1270
rect 275 1262 276 1270
rect 288 1262 289 1270
rect 291 1262 294 1270
rect 296 1262 297 1270
rect 309 1262 310 1270
rect 312 1266 313 1270
rect 312 1262 317 1266
rect 325 1262 326 1270
rect 328 1262 331 1270
rect 333 1262 334 1270
rect 351 1262 352 1270
rect 354 1262 355 1270
rect 367 1262 368 1270
rect 370 1266 371 1270
rect 370 1262 375 1266
rect 383 1262 384 1270
rect 386 1262 389 1270
rect 391 1262 392 1270
rect 404 1262 405 1270
rect 407 1262 408 1270
rect 957 1262 958 1270
rect 960 1262 963 1270
rect 965 1262 966 1270
rect 978 1262 979 1270
rect 981 1266 982 1270
rect 981 1262 986 1266
rect 994 1262 995 1270
rect 997 1262 1000 1270
rect 1002 1262 1003 1270
rect 1020 1262 1021 1270
rect 1023 1262 1024 1270
rect 1036 1262 1037 1270
rect 1039 1266 1040 1270
rect 1039 1262 1044 1266
rect 1052 1262 1053 1270
rect 1055 1262 1058 1270
rect 1060 1262 1061 1270
rect 1073 1262 1074 1270
rect 1076 1262 1077 1270
rect 1089 1262 1090 1270
rect 1092 1262 1095 1270
rect 1097 1262 1098 1270
rect 1110 1262 1111 1270
rect 1113 1266 1114 1270
rect 1113 1262 1118 1266
rect 1126 1262 1127 1270
rect 1129 1262 1132 1270
rect 1134 1262 1135 1270
rect 1152 1262 1153 1270
rect 1155 1262 1156 1270
rect 1168 1262 1169 1270
rect 1171 1266 1172 1270
rect 1171 1262 1176 1266
rect 1184 1262 1185 1270
rect 1187 1262 1190 1270
rect 1192 1262 1193 1270
rect 1205 1262 1206 1270
rect 1208 1262 1209 1270
rect 1221 1262 1222 1270
rect 1224 1262 1227 1270
rect 1229 1262 1230 1270
rect 1242 1262 1243 1270
rect 1245 1266 1246 1270
rect 1245 1262 1250 1266
rect 1258 1262 1259 1270
rect 1261 1262 1264 1270
rect 1266 1262 1267 1270
rect 1284 1262 1285 1270
rect 1287 1262 1288 1270
rect 1300 1262 1301 1270
rect 1303 1266 1304 1270
rect 1303 1262 1308 1266
rect 1316 1262 1317 1270
rect 1319 1262 1322 1270
rect 1324 1262 1325 1270
rect 1337 1262 1338 1270
rect 1340 1262 1341 1270
rect 795 1206 796 1214
rect 798 1206 801 1214
rect 803 1206 804 1214
rect 816 1206 817 1214
rect 819 1210 820 1214
rect 819 1206 824 1210
rect 832 1206 833 1214
rect 835 1206 838 1214
rect 840 1206 841 1214
rect 858 1206 859 1214
rect 861 1206 862 1214
rect 874 1206 875 1214
rect 877 1210 878 1214
rect 877 1206 882 1210
rect 890 1206 891 1214
rect 893 1206 896 1214
rect 898 1206 899 1214
rect 911 1206 912 1214
rect 914 1206 915 1214
rect 1728 1206 1729 1214
rect 1731 1206 1734 1214
rect 1736 1206 1737 1214
rect 1749 1206 1750 1214
rect 1752 1210 1753 1214
rect 1752 1206 1757 1210
rect 1765 1206 1766 1214
rect 1768 1206 1771 1214
rect 1773 1206 1774 1214
rect 1791 1206 1792 1214
rect 1794 1206 1795 1214
rect 1807 1206 1808 1214
rect 1810 1210 1811 1214
rect 1810 1206 1815 1210
rect 1823 1206 1824 1214
rect 1826 1206 1829 1214
rect 1831 1206 1832 1214
rect 1844 1206 1845 1214
rect 1847 1206 1848 1214
rect 24 1176 25 1184
rect 27 1176 30 1184
rect 32 1176 33 1184
rect 45 1176 46 1184
rect 48 1180 49 1184
rect 48 1176 53 1180
rect 61 1176 62 1184
rect 64 1176 67 1184
rect 69 1176 70 1184
rect 87 1176 88 1184
rect 90 1176 91 1184
rect 103 1176 104 1184
rect 106 1180 107 1184
rect 106 1176 111 1180
rect 119 1176 120 1184
rect 122 1176 125 1184
rect 127 1176 128 1184
rect 140 1176 141 1184
rect 143 1176 144 1184
rect 156 1176 157 1184
rect 159 1176 162 1184
rect 164 1176 165 1184
rect 177 1176 178 1184
rect 180 1180 181 1184
rect 180 1176 185 1180
rect 193 1176 194 1184
rect 196 1176 199 1184
rect 201 1176 202 1184
rect 219 1176 220 1184
rect 222 1176 223 1184
rect 235 1176 236 1184
rect 238 1180 239 1184
rect 238 1176 243 1180
rect 251 1176 252 1184
rect 254 1176 257 1184
rect 259 1176 260 1184
rect 272 1176 273 1184
rect 275 1176 276 1184
rect 288 1176 289 1184
rect 291 1176 294 1184
rect 296 1176 297 1184
rect 309 1176 310 1184
rect 312 1180 313 1184
rect 312 1176 317 1180
rect 325 1176 326 1184
rect 328 1176 331 1184
rect 333 1176 334 1184
rect 351 1176 352 1184
rect 354 1176 355 1184
rect 367 1176 368 1184
rect 370 1180 371 1184
rect 370 1176 375 1180
rect 383 1176 384 1184
rect 386 1176 389 1184
rect 391 1176 392 1184
rect 404 1176 405 1184
rect 407 1176 408 1184
rect 957 1176 958 1184
rect 960 1176 963 1184
rect 965 1176 966 1184
rect 978 1176 979 1184
rect 981 1180 982 1184
rect 981 1176 986 1180
rect 994 1176 995 1184
rect 997 1176 1000 1184
rect 1002 1176 1003 1184
rect 1020 1176 1021 1184
rect 1023 1176 1024 1184
rect 1036 1176 1037 1184
rect 1039 1180 1040 1184
rect 1039 1176 1044 1180
rect 1052 1176 1053 1184
rect 1055 1176 1058 1184
rect 1060 1176 1061 1184
rect 1073 1176 1074 1184
rect 1076 1176 1077 1184
rect 1089 1176 1090 1184
rect 1092 1176 1095 1184
rect 1097 1176 1098 1184
rect 1110 1176 1111 1184
rect 1113 1180 1114 1184
rect 1113 1176 1118 1180
rect 1126 1176 1127 1184
rect 1129 1176 1132 1184
rect 1134 1176 1135 1184
rect 1152 1176 1153 1184
rect 1155 1176 1156 1184
rect 1168 1176 1169 1184
rect 1171 1180 1172 1184
rect 1171 1176 1176 1180
rect 1184 1176 1185 1184
rect 1187 1176 1190 1184
rect 1192 1176 1193 1184
rect 1205 1176 1206 1184
rect 1208 1176 1209 1184
rect 1221 1176 1222 1184
rect 1224 1176 1227 1184
rect 1229 1176 1230 1184
rect 1242 1176 1243 1184
rect 1245 1180 1246 1184
rect 1245 1176 1250 1180
rect 1258 1176 1259 1184
rect 1261 1176 1264 1184
rect 1266 1176 1267 1184
rect 1284 1176 1285 1184
rect 1287 1176 1288 1184
rect 1300 1176 1301 1184
rect 1303 1180 1304 1184
rect 1303 1176 1308 1180
rect 1316 1176 1317 1184
rect 1319 1176 1322 1184
rect 1324 1176 1325 1184
rect 1337 1176 1338 1184
rect 1340 1176 1341 1184
rect 24 1036 25 1044
rect 27 1036 30 1044
rect 32 1036 33 1044
rect 45 1036 46 1044
rect 48 1040 49 1044
rect 48 1036 53 1040
rect 61 1036 62 1044
rect 64 1036 67 1044
rect 69 1036 70 1044
rect 87 1036 88 1044
rect 90 1036 91 1044
rect 103 1036 104 1044
rect 106 1040 107 1044
rect 106 1036 111 1040
rect 119 1036 120 1044
rect 122 1036 125 1044
rect 127 1036 128 1044
rect 140 1036 141 1044
rect 143 1036 144 1044
rect 156 1036 157 1044
rect 159 1036 162 1044
rect 164 1036 165 1044
rect 177 1036 178 1044
rect 180 1040 181 1044
rect 180 1036 185 1040
rect 193 1036 194 1044
rect 196 1036 199 1044
rect 201 1036 202 1044
rect 219 1036 220 1044
rect 222 1036 223 1044
rect 235 1036 236 1044
rect 238 1040 239 1044
rect 238 1036 243 1040
rect 251 1036 252 1044
rect 254 1036 257 1044
rect 259 1036 260 1044
rect 272 1036 273 1044
rect 275 1036 276 1044
rect 288 1036 289 1044
rect 291 1036 294 1044
rect 296 1036 297 1044
rect 309 1036 310 1044
rect 312 1040 313 1044
rect 312 1036 317 1040
rect 325 1036 326 1044
rect 328 1036 331 1044
rect 333 1036 334 1044
rect 351 1036 352 1044
rect 354 1036 355 1044
rect 367 1036 368 1044
rect 370 1040 371 1044
rect 370 1036 375 1040
rect 383 1036 384 1044
rect 386 1036 389 1044
rect 391 1036 392 1044
rect 404 1036 405 1044
rect 407 1036 408 1044
rect 957 1036 958 1044
rect 960 1036 963 1044
rect 965 1036 966 1044
rect 978 1036 979 1044
rect 981 1040 982 1044
rect 981 1036 986 1040
rect 994 1036 995 1044
rect 997 1036 1000 1044
rect 1002 1036 1003 1044
rect 1020 1036 1021 1044
rect 1023 1036 1024 1044
rect 1036 1036 1037 1044
rect 1039 1040 1040 1044
rect 1039 1036 1044 1040
rect 1052 1036 1053 1044
rect 1055 1036 1058 1044
rect 1060 1036 1061 1044
rect 1073 1036 1074 1044
rect 1076 1036 1077 1044
rect 1089 1036 1090 1044
rect 1092 1036 1095 1044
rect 1097 1036 1098 1044
rect 1110 1036 1111 1044
rect 1113 1040 1114 1044
rect 1113 1036 1118 1040
rect 1126 1036 1127 1044
rect 1129 1036 1132 1044
rect 1134 1036 1135 1044
rect 1152 1036 1153 1044
rect 1155 1036 1156 1044
rect 1168 1036 1169 1044
rect 1171 1040 1172 1044
rect 1171 1036 1176 1040
rect 1184 1036 1185 1044
rect 1187 1036 1190 1044
rect 1192 1036 1193 1044
rect 1205 1036 1206 1044
rect 1208 1036 1209 1044
rect 1221 1036 1222 1044
rect 1224 1036 1227 1044
rect 1229 1036 1230 1044
rect 1242 1036 1243 1044
rect 1245 1040 1246 1044
rect 1245 1036 1250 1040
rect 1258 1036 1259 1044
rect 1261 1036 1264 1044
rect 1266 1036 1267 1044
rect 1284 1036 1285 1044
rect 1287 1036 1288 1044
rect 1300 1036 1301 1044
rect 1303 1040 1304 1044
rect 1303 1036 1308 1040
rect 1316 1036 1317 1044
rect 1319 1036 1322 1044
rect 1324 1036 1325 1044
rect 1337 1036 1338 1044
rect 1340 1036 1341 1044
rect 496 957 497 965
rect 499 957 502 965
rect 504 957 505 965
rect 517 957 518 965
rect 520 961 521 965
rect 520 957 525 961
rect 533 957 534 965
rect 536 957 539 965
rect 541 957 542 965
rect 559 957 560 965
rect 562 957 563 965
rect 575 957 576 965
rect 578 961 579 965
rect 578 957 583 961
rect 591 957 592 965
rect 594 957 597 965
rect 599 957 600 965
rect 612 957 613 965
rect 615 957 616 965
rect 628 957 629 965
rect 631 957 634 965
rect 636 957 637 965
rect 649 957 650 965
rect 652 961 653 965
rect 652 957 657 961
rect 665 957 666 965
rect 668 957 671 965
rect 673 957 674 965
rect 691 957 692 965
rect 694 957 695 965
rect 707 957 708 965
rect 710 961 711 965
rect 710 957 715 961
rect 723 957 724 965
rect 726 957 729 965
rect 731 957 732 965
rect 744 957 745 965
rect 747 957 748 965
rect 760 957 761 965
rect 763 957 766 965
rect 768 957 769 965
rect 781 957 782 965
rect 784 961 785 965
rect 784 957 789 961
rect 797 957 798 965
rect 800 957 803 965
rect 805 957 806 965
rect 823 957 824 965
rect 826 957 827 965
rect 839 957 840 965
rect 842 961 843 965
rect 842 957 847 961
rect 855 957 856 965
rect 858 957 861 965
rect 863 957 864 965
rect 876 957 877 965
rect 879 957 880 965
rect 892 957 893 965
rect 895 957 898 965
rect 900 957 901 965
rect 913 957 914 965
rect 916 961 917 965
rect 916 957 921 961
rect 929 957 930 965
rect 932 957 935 965
rect 937 957 938 965
rect 955 957 956 965
rect 958 957 959 965
rect 971 957 972 965
rect 974 961 975 965
rect 974 957 979 961
rect 987 957 988 965
rect 990 957 993 965
rect 995 957 996 965
rect 1008 957 1009 965
rect 1011 957 1012 965
rect 1429 957 1430 965
rect 1432 957 1435 965
rect 1437 957 1438 965
rect 1450 957 1451 965
rect 1453 961 1454 965
rect 1453 957 1458 961
rect 1466 957 1467 965
rect 1469 957 1472 965
rect 1474 957 1475 965
rect 1492 957 1493 965
rect 1495 957 1496 965
rect 1508 957 1509 965
rect 1511 961 1512 965
rect 1511 957 1516 961
rect 1524 957 1525 965
rect 1527 957 1530 965
rect 1532 957 1533 965
rect 1545 957 1546 965
rect 1548 957 1549 965
rect 1561 957 1562 965
rect 1564 957 1567 965
rect 1569 957 1570 965
rect 1582 957 1583 965
rect 1585 961 1586 965
rect 1585 957 1590 961
rect 1598 957 1599 965
rect 1601 957 1604 965
rect 1606 957 1607 965
rect 1624 957 1625 965
rect 1627 957 1628 965
rect 1640 957 1641 965
rect 1643 961 1644 965
rect 1643 957 1648 961
rect 1656 957 1657 965
rect 1659 957 1662 965
rect 1664 957 1665 965
rect 1677 957 1678 965
rect 1680 957 1681 965
rect 1693 957 1694 965
rect 1696 957 1699 965
rect 1701 957 1702 965
rect 1714 957 1715 965
rect 1717 961 1718 965
rect 1717 957 1722 961
rect 1730 957 1731 965
rect 1733 957 1736 965
rect 1738 957 1739 965
rect 1756 957 1757 965
rect 1759 957 1760 965
rect 1772 957 1773 965
rect 1775 961 1776 965
rect 1775 957 1780 961
rect 1788 957 1789 965
rect 1791 957 1794 965
rect 1796 957 1797 965
rect 1809 957 1810 965
rect 1812 957 1813 965
rect 1825 957 1826 965
rect 1828 957 1831 965
rect 1833 957 1834 965
rect 1846 957 1847 965
rect 1849 961 1850 965
rect 1849 957 1854 961
rect 1862 957 1863 965
rect 1865 957 1868 965
rect 1870 957 1871 965
rect 1888 957 1889 965
rect 1891 957 1892 965
rect 1904 957 1905 965
rect 1907 961 1908 965
rect 1907 957 1912 961
rect 1920 957 1921 965
rect 1923 957 1926 965
rect 1928 957 1929 965
rect 1941 957 1942 965
rect 1944 957 1945 965
rect 156 924 157 932
rect 159 924 162 932
rect 164 924 165 932
rect 177 924 178 932
rect 180 928 181 932
rect 180 924 185 928
rect 193 924 194 932
rect 196 924 199 932
rect 201 924 202 932
rect 219 924 220 932
rect 222 924 223 932
rect 235 924 236 932
rect 238 928 239 932
rect 238 924 243 928
rect 251 924 252 932
rect 254 924 257 932
rect 259 924 260 932
rect 272 924 273 932
rect 275 924 276 932
rect 1089 924 1090 932
rect 1092 924 1095 932
rect 1097 924 1098 932
rect 1110 924 1111 932
rect 1113 928 1114 932
rect 1113 924 1118 928
rect 1126 924 1127 932
rect 1129 924 1132 932
rect 1134 924 1135 932
rect 1152 924 1153 932
rect 1155 924 1156 932
rect 1168 924 1169 932
rect 1171 928 1172 932
rect 1171 924 1176 928
rect 1184 924 1185 932
rect 1187 924 1190 932
rect 1192 924 1193 932
rect 1205 924 1206 932
rect 1208 924 1209 932
rect 675 886 676 894
rect 678 886 679 894
rect 501 873 502 881
rect 504 873 505 881
rect 517 873 518 881
rect 520 873 521 881
rect 533 873 534 881
rect 536 873 537 881
rect 552 873 557 881
rect 559 873 562 881
rect 564 873 565 881
rect 586 873 588 881
rect 590 873 591 881
rect 608 873 609 881
rect 611 873 612 881
rect 624 873 629 881
rect 631 873 634 881
rect 636 873 637 881
rect 651 873 652 881
rect 654 873 655 881
rect 699 880 702 888
rect 704 880 707 888
rect 709 880 710 888
rect 729 886 730 894
rect 732 886 733 894
rect 756 886 757 894
rect 759 886 760 894
rect 780 880 783 888
rect 785 880 788 888
rect 790 880 791 888
rect 810 886 811 894
rect 813 886 814 894
rect 1608 886 1609 894
rect 1611 886 1612 894
rect 1434 873 1435 881
rect 1437 873 1438 881
rect 1450 873 1451 881
rect 1453 873 1454 881
rect 1466 873 1467 881
rect 1469 873 1470 881
rect 1485 873 1490 881
rect 1492 873 1495 881
rect 1497 873 1498 881
rect 1519 873 1521 881
rect 1523 873 1524 881
rect 1541 873 1542 881
rect 1544 873 1545 881
rect 1557 873 1562 881
rect 1564 873 1567 881
rect 1569 873 1570 881
rect 1584 873 1585 881
rect 1587 873 1588 881
rect 1632 880 1635 888
rect 1637 880 1640 888
rect 1642 880 1643 888
rect 1662 886 1663 894
rect 1665 886 1666 894
rect 1689 886 1690 894
rect 1692 886 1693 894
rect 1713 880 1716 888
rect 1718 880 1721 888
rect 1723 880 1724 888
rect 1743 886 1744 894
rect 1746 886 1747 894
rect 147 822 148 830
rect 150 822 151 830
rect 163 822 164 830
rect 166 822 169 830
rect 171 822 172 830
rect 184 826 185 830
rect 180 822 185 826
rect 187 822 188 830
rect 200 822 201 830
rect 203 822 204 830
rect 221 822 222 830
rect 224 822 227 830
rect 229 822 230 830
rect 242 826 243 830
rect 238 822 243 826
rect 245 822 246 830
rect 258 822 259 830
rect 261 822 264 830
rect 266 822 267 830
rect 1080 822 1081 830
rect 1083 822 1084 830
rect 1096 822 1097 830
rect 1099 822 1102 830
rect 1104 822 1105 830
rect 1117 826 1118 830
rect 1113 822 1118 826
rect 1120 822 1121 830
rect 1133 822 1134 830
rect 1136 822 1137 830
rect 1154 822 1155 830
rect 1157 822 1160 830
rect 1162 822 1163 830
rect 1175 826 1176 830
rect 1171 822 1176 826
rect 1178 822 1179 830
rect 1191 822 1192 830
rect 1194 822 1197 830
rect 1199 822 1200 830
rect 501 787 502 795
rect 504 787 505 795
rect 517 787 518 795
rect 520 787 521 795
rect 533 787 534 795
rect 536 787 537 795
rect 552 787 557 795
rect 559 787 562 795
rect 564 787 565 795
rect 586 787 588 795
rect 590 787 591 795
rect 608 787 609 795
rect 611 787 612 795
rect 624 787 629 795
rect 631 787 634 795
rect 636 787 637 795
rect 651 787 652 795
rect 654 787 655 795
rect 699 788 702 796
rect 704 788 707 796
rect 709 788 710 796
rect 780 788 783 796
rect 785 788 788 796
rect 790 788 791 796
rect 1434 787 1435 795
rect 1437 787 1438 795
rect 1450 787 1451 795
rect 1453 787 1454 795
rect 1466 787 1467 795
rect 1469 787 1470 795
rect 1485 787 1490 795
rect 1492 787 1495 795
rect 1497 787 1498 795
rect 1519 787 1521 795
rect 1523 787 1524 795
rect 1541 787 1542 795
rect 1544 787 1545 795
rect 1557 787 1562 795
rect 1564 787 1567 795
rect 1569 787 1570 795
rect 1584 787 1585 795
rect 1587 787 1588 795
rect 1632 788 1635 796
rect 1637 788 1640 796
rect 1642 788 1643 796
rect 1713 788 1716 796
rect 1718 788 1721 796
rect 1723 788 1724 796
rect 501 741 502 749
rect 504 741 505 749
rect 517 741 518 749
rect 520 741 521 749
rect 533 741 534 749
rect 536 741 537 749
rect 552 741 557 749
rect 559 741 562 749
rect 564 741 565 749
rect 586 741 588 749
rect 590 741 591 749
rect 608 741 609 749
rect 611 741 612 749
rect 624 741 629 749
rect 631 741 634 749
rect 636 741 637 749
rect 651 741 652 749
rect 654 741 655 749
rect 699 748 702 756
rect 704 748 707 756
rect 709 748 710 756
rect 729 754 730 762
rect 732 754 733 762
rect 780 754 781 762
rect 783 754 784 762
rect 804 748 807 756
rect 809 748 812 756
rect 814 748 815 756
rect 834 754 835 762
rect 837 754 838 762
rect 1434 741 1435 749
rect 1437 741 1438 749
rect 1450 741 1451 749
rect 1453 741 1454 749
rect 1466 741 1467 749
rect 1469 741 1470 749
rect 1485 741 1490 749
rect 1492 741 1495 749
rect 1497 741 1498 749
rect 1519 741 1521 749
rect 1523 741 1524 749
rect 1541 741 1542 749
rect 1544 741 1545 749
rect 1557 741 1562 749
rect 1564 741 1567 749
rect 1569 741 1570 749
rect 1584 741 1585 749
rect 1587 741 1588 749
rect 1632 748 1635 756
rect 1637 748 1640 756
rect 1642 748 1643 756
rect 1662 754 1663 762
rect 1665 754 1666 762
rect 1713 754 1714 762
rect 1716 754 1717 762
rect 1737 748 1740 756
rect 1742 748 1745 756
rect 1747 748 1748 756
rect 1767 754 1768 762
rect 1770 754 1771 762
rect 501 655 502 663
rect 504 655 505 663
rect 517 655 518 663
rect 520 655 521 663
rect 533 655 534 663
rect 536 655 537 663
rect 552 655 557 663
rect 559 655 562 663
rect 564 655 565 663
rect 586 655 588 663
rect 590 655 591 663
rect 608 655 609 663
rect 611 655 612 663
rect 624 655 629 663
rect 631 655 634 663
rect 636 655 637 663
rect 651 655 652 663
rect 654 655 655 663
rect 699 657 702 665
rect 704 657 707 665
rect 709 657 710 665
rect 804 657 807 665
rect 809 657 812 665
rect 814 657 815 665
rect 1434 655 1435 663
rect 1437 655 1438 663
rect 1450 655 1451 663
rect 1453 655 1454 663
rect 1466 655 1467 663
rect 1469 655 1470 663
rect 1485 655 1490 663
rect 1492 655 1495 663
rect 1497 655 1498 663
rect 1519 655 1521 663
rect 1523 655 1524 663
rect 1541 655 1542 663
rect 1544 655 1545 663
rect 1557 655 1562 663
rect 1564 655 1567 663
rect 1569 655 1570 663
rect 1584 655 1585 663
rect 1587 655 1588 663
rect 1632 657 1635 665
rect 1637 657 1640 665
rect 1642 657 1643 665
rect 1737 657 1740 665
rect 1742 657 1745 665
rect 1747 657 1748 665
rect 501 609 502 617
rect 504 609 505 617
rect 517 609 518 617
rect 520 609 521 617
rect 533 609 534 617
rect 536 609 537 617
rect 552 609 557 617
rect 559 609 562 617
rect 564 609 565 617
rect 586 609 588 617
rect 590 609 591 617
rect 608 609 609 617
rect 611 609 612 617
rect 624 609 629 617
rect 631 609 634 617
rect 636 609 637 617
rect 651 609 652 617
rect 654 609 655 617
rect 699 616 702 624
rect 704 616 707 624
rect 709 616 710 624
rect 729 622 730 630
rect 732 622 733 630
rect 756 622 757 630
rect 759 622 760 630
rect 780 616 783 624
rect 785 616 788 624
rect 790 616 791 624
rect 810 622 811 630
rect 813 622 814 630
rect 846 622 847 630
rect 849 622 850 630
rect 870 616 873 624
rect 875 616 878 624
rect 880 616 881 624
rect 900 622 901 630
rect 903 622 904 630
rect 1434 609 1435 617
rect 1437 609 1438 617
rect 1450 609 1451 617
rect 1453 609 1454 617
rect 1466 609 1467 617
rect 1469 609 1470 617
rect 1485 609 1490 617
rect 1492 609 1495 617
rect 1497 609 1498 617
rect 1519 609 1521 617
rect 1523 609 1524 617
rect 1541 609 1542 617
rect 1544 609 1545 617
rect 1557 609 1562 617
rect 1564 609 1567 617
rect 1569 609 1570 617
rect 1584 609 1585 617
rect 1587 609 1588 617
rect 1632 616 1635 624
rect 1637 616 1640 624
rect 1642 616 1643 624
rect 1662 622 1663 630
rect 1665 622 1666 630
rect 1689 622 1690 630
rect 1692 622 1693 630
rect 1713 616 1716 624
rect 1718 616 1721 624
rect 1723 616 1724 624
rect 1743 622 1744 630
rect 1746 622 1747 630
rect 1779 622 1780 630
rect 1782 622 1783 630
rect 1803 616 1806 624
rect 1808 616 1811 624
rect 1813 616 1814 624
rect 1833 622 1834 630
rect 1836 622 1837 630
rect 501 523 502 531
rect 504 523 505 531
rect 517 523 518 531
rect 520 523 521 531
rect 533 523 534 531
rect 536 523 537 531
rect 552 523 557 531
rect 559 523 562 531
rect 564 523 565 531
rect 586 523 588 531
rect 590 523 591 531
rect 608 523 609 531
rect 611 523 612 531
rect 624 523 629 531
rect 631 523 634 531
rect 636 523 637 531
rect 651 523 652 531
rect 654 523 655 531
rect 699 522 702 530
rect 704 522 707 530
rect 709 522 710 530
rect 780 522 783 530
rect 785 522 788 530
rect 790 522 791 530
rect 870 522 873 530
rect 875 522 878 530
rect 880 522 881 530
rect 1434 523 1435 531
rect 1437 523 1438 531
rect 1450 523 1451 531
rect 1453 523 1454 531
rect 1466 523 1467 531
rect 1469 523 1470 531
rect 1485 523 1490 531
rect 1492 523 1495 531
rect 1497 523 1498 531
rect 1519 523 1521 531
rect 1523 523 1524 531
rect 1541 523 1542 531
rect 1544 523 1545 531
rect 1557 523 1562 531
rect 1564 523 1567 531
rect 1569 523 1570 531
rect 1584 523 1585 531
rect 1587 523 1588 531
rect 1632 522 1635 530
rect 1637 522 1640 530
rect 1642 522 1643 530
rect 1713 522 1716 530
rect 1718 522 1721 530
rect 1723 522 1724 530
rect 1803 522 1806 530
rect 1808 522 1811 530
rect 1813 522 1814 530
rect 501 477 502 485
rect 504 477 505 485
rect 517 477 518 485
rect 520 477 521 485
rect 533 477 534 485
rect 536 477 537 485
rect 552 477 557 485
rect 559 477 562 485
rect 564 477 565 485
rect 586 477 588 485
rect 590 477 591 485
rect 608 477 609 485
rect 611 477 612 485
rect 624 477 629 485
rect 631 477 634 485
rect 636 477 637 485
rect 651 477 652 485
rect 654 477 655 485
rect 699 484 702 492
rect 704 484 707 492
rect 709 484 710 492
rect 729 490 730 498
rect 732 490 733 498
rect 1434 477 1435 485
rect 1437 477 1438 485
rect 1450 477 1451 485
rect 1453 477 1454 485
rect 1466 477 1467 485
rect 1469 477 1470 485
rect 1485 477 1490 485
rect 1492 477 1495 485
rect 1497 477 1498 485
rect 1519 477 1521 485
rect 1523 477 1524 485
rect 1541 477 1542 485
rect 1544 477 1545 485
rect 1557 477 1562 485
rect 1564 477 1567 485
rect 1569 477 1570 485
rect 1584 477 1585 485
rect 1587 477 1588 485
rect 1632 484 1635 492
rect 1637 484 1640 492
rect 1642 484 1643 492
rect 1662 490 1663 498
rect 1665 490 1666 498
rect 24 422 25 430
rect 27 422 30 430
rect 32 422 33 430
rect 45 422 46 430
rect 48 426 49 430
rect 48 422 53 426
rect 61 422 62 430
rect 64 422 67 430
rect 69 422 70 430
rect 87 422 88 430
rect 90 422 91 430
rect 103 422 104 430
rect 106 426 107 430
rect 106 422 111 426
rect 119 422 120 430
rect 122 422 125 430
rect 127 422 128 430
rect 140 422 141 430
rect 143 422 144 430
rect 156 422 157 430
rect 159 422 162 430
rect 164 422 165 430
rect 177 422 178 430
rect 180 426 181 430
rect 180 422 185 426
rect 193 422 194 430
rect 196 422 199 430
rect 201 422 202 430
rect 219 422 220 430
rect 222 422 223 430
rect 235 422 236 430
rect 238 426 239 430
rect 238 422 243 426
rect 251 422 252 430
rect 254 422 257 430
rect 259 422 260 430
rect 272 422 273 430
rect 275 422 276 430
rect 288 422 289 430
rect 291 422 294 430
rect 296 422 297 430
rect 309 422 310 430
rect 312 426 313 430
rect 312 422 317 426
rect 325 422 326 430
rect 328 422 331 430
rect 333 422 334 430
rect 351 422 352 430
rect 354 422 355 430
rect 367 422 368 430
rect 370 426 371 430
rect 370 422 375 426
rect 383 422 384 430
rect 386 422 389 430
rect 391 422 392 430
rect 404 422 405 430
rect 407 422 408 430
rect 957 422 958 430
rect 960 422 963 430
rect 965 422 966 430
rect 978 422 979 430
rect 981 426 982 430
rect 981 422 986 426
rect 994 422 995 430
rect 997 422 1000 430
rect 1002 422 1003 430
rect 1020 422 1021 430
rect 1023 422 1024 430
rect 1036 422 1037 430
rect 1039 426 1040 430
rect 1039 422 1044 426
rect 1052 422 1053 430
rect 1055 422 1058 430
rect 1060 422 1061 430
rect 1073 422 1074 430
rect 1076 422 1077 430
rect 1089 422 1090 430
rect 1092 422 1095 430
rect 1097 422 1098 430
rect 1110 422 1111 430
rect 1113 426 1114 430
rect 1113 422 1118 426
rect 1126 422 1127 430
rect 1129 422 1132 430
rect 1134 422 1135 430
rect 1152 422 1153 430
rect 1155 422 1156 430
rect 1168 422 1169 430
rect 1171 426 1172 430
rect 1171 422 1176 426
rect 1184 422 1185 430
rect 1187 422 1190 430
rect 1192 422 1193 430
rect 1205 422 1206 430
rect 1208 422 1209 430
rect 1221 422 1222 430
rect 1224 422 1227 430
rect 1229 422 1230 430
rect 1242 422 1243 430
rect 1245 426 1246 430
rect 1245 422 1250 426
rect 1258 422 1259 430
rect 1261 422 1264 430
rect 1266 422 1267 430
rect 1284 422 1285 430
rect 1287 422 1288 430
rect 1300 422 1301 430
rect 1303 426 1304 430
rect 1303 422 1308 426
rect 1316 422 1317 430
rect 1319 422 1322 430
rect 1324 422 1325 430
rect 1337 422 1338 430
rect 1340 422 1341 430
rect 501 391 502 399
rect 504 391 505 399
rect 517 391 518 399
rect 520 391 521 399
rect 533 391 534 399
rect 536 391 537 399
rect 552 391 557 399
rect 559 391 562 399
rect 564 391 565 399
rect 586 391 588 399
rect 590 391 591 399
rect 608 391 609 399
rect 611 391 612 399
rect 624 391 629 399
rect 631 391 634 399
rect 636 391 637 399
rect 651 391 652 399
rect 654 391 655 399
rect 699 386 702 394
rect 704 386 707 394
rect 709 386 710 394
rect 735 391 736 399
rect 738 391 739 399
rect 743 391 749 399
rect 753 391 754 399
rect 756 391 757 399
rect 778 391 779 399
rect 781 391 782 399
rect 794 391 795 399
rect 797 391 798 399
rect 813 391 818 399
rect 820 391 823 399
rect 825 391 826 399
rect 847 391 849 399
rect 851 391 852 399
rect 869 391 870 399
rect 872 391 873 399
rect 885 391 890 399
rect 892 391 895 399
rect 897 391 898 399
rect 912 391 913 399
rect 915 391 916 399
rect 1434 391 1435 399
rect 1437 391 1438 399
rect 1450 391 1451 399
rect 1453 391 1454 399
rect 1466 391 1467 399
rect 1469 391 1470 399
rect 1485 391 1490 399
rect 1492 391 1495 399
rect 1497 391 1498 399
rect 1519 391 1521 399
rect 1523 391 1524 399
rect 1541 391 1542 399
rect 1544 391 1545 399
rect 1557 391 1562 399
rect 1564 391 1567 399
rect 1569 391 1570 399
rect 1584 391 1585 399
rect 1587 391 1588 399
rect 1632 386 1635 394
rect 1637 386 1640 394
rect 1642 386 1643 394
rect 1668 391 1669 399
rect 1671 391 1672 399
rect 1676 391 1682 399
rect 1686 391 1687 399
rect 1689 391 1690 399
rect 1711 391 1712 399
rect 1714 391 1715 399
rect 1727 391 1728 399
rect 1730 391 1731 399
rect 1746 391 1751 399
rect 1753 391 1756 399
rect 1758 391 1759 399
rect 1780 391 1782 399
rect 1784 391 1785 399
rect 1802 391 1803 399
rect 1805 391 1806 399
rect 1818 391 1823 399
rect 1825 391 1828 399
rect 1830 391 1831 399
rect 1845 391 1846 399
rect 1848 391 1849 399
rect 795 312 796 320
rect 798 312 801 320
rect 803 312 804 320
rect 816 312 817 320
rect 819 316 820 320
rect 819 312 824 316
rect 832 312 833 320
rect 835 312 838 320
rect 840 312 841 320
rect 858 312 859 320
rect 861 312 862 320
rect 874 312 875 320
rect 877 316 878 320
rect 877 312 882 316
rect 890 312 891 320
rect 893 312 896 320
rect 898 312 899 320
rect 911 312 912 320
rect 914 312 915 320
rect 1728 312 1729 320
rect 1731 312 1734 320
rect 1736 312 1737 320
rect 1749 312 1750 320
rect 1752 316 1753 320
rect 1752 312 1757 316
rect 1765 312 1766 320
rect 1768 312 1771 320
rect 1773 312 1774 320
rect 1791 312 1792 320
rect 1794 312 1795 320
rect 1807 312 1808 320
rect 1810 316 1811 320
rect 1810 312 1815 316
rect 1823 312 1824 320
rect 1826 312 1829 320
rect 1831 312 1832 320
rect 1844 312 1845 320
rect 1847 312 1848 320
rect 24 282 25 290
rect 27 282 30 290
rect 32 282 33 290
rect 45 282 46 290
rect 48 286 49 290
rect 48 282 53 286
rect 61 282 62 290
rect 64 282 67 290
rect 69 282 70 290
rect 87 282 88 290
rect 90 282 91 290
rect 103 282 104 290
rect 106 286 107 290
rect 106 282 111 286
rect 119 282 120 290
rect 122 282 125 290
rect 127 282 128 290
rect 140 282 141 290
rect 143 282 144 290
rect 156 282 157 290
rect 159 282 162 290
rect 164 282 165 290
rect 177 282 178 290
rect 180 286 181 290
rect 180 282 185 286
rect 193 282 194 290
rect 196 282 199 290
rect 201 282 202 290
rect 219 282 220 290
rect 222 282 223 290
rect 235 282 236 290
rect 238 286 239 290
rect 238 282 243 286
rect 251 282 252 290
rect 254 282 257 290
rect 259 282 260 290
rect 272 282 273 290
rect 275 282 276 290
rect 288 282 289 290
rect 291 282 294 290
rect 296 282 297 290
rect 309 282 310 290
rect 312 286 313 290
rect 312 282 317 286
rect 325 282 326 290
rect 328 282 331 290
rect 333 282 334 290
rect 351 282 352 290
rect 354 282 355 290
rect 367 282 368 290
rect 370 286 371 290
rect 370 282 375 286
rect 383 282 384 290
rect 386 282 389 290
rect 391 282 392 290
rect 404 282 405 290
rect 407 282 408 290
rect 957 282 958 290
rect 960 282 963 290
rect 965 282 966 290
rect 978 282 979 290
rect 981 286 982 290
rect 981 282 986 286
rect 994 282 995 290
rect 997 282 1000 290
rect 1002 282 1003 290
rect 1020 282 1021 290
rect 1023 282 1024 290
rect 1036 282 1037 290
rect 1039 286 1040 290
rect 1039 282 1044 286
rect 1052 282 1053 290
rect 1055 282 1058 290
rect 1060 282 1061 290
rect 1073 282 1074 290
rect 1076 282 1077 290
rect 1089 282 1090 290
rect 1092 282 1095 290
rect 1097 282 1098 290
rect 1110 282 1111 290
rect 1113 286 1114 290
rect 1113 282 1118 286
rect 1126 282 1127 290
rect 1129 282 1132 290
rect 1134 282 1135 290
rect 1152 282 1153 290
rect 1155 282 1156 290
rect 1168 282 1169 290
rect 1171 286 1172 290
rect 1171 282 1176 286
rect 1184 282 1185 290
rect 1187 282 1190 290
rect 1192 282 1193 290
rect 1205 282 1206 290
rect 1208 282 1209 290
rect 1221 282 1222 290
rect 1224 282 1227 290
rect 1229 282 1230 290
rect 1242 282 1243 290
rect 1245 286 1246 290
rect 1245 282 1250 286
rect 1258 282 1259 290
rect 1261 282 1264 290
rect 1266 282 1267 290
rect 1284 282 1285 290
rect 1287 282 1288 290
rect 1300 282 1301 290
rect 1303 286 1304 290
rect 1303 282 1308 286
rect 1316 282 1317 290
rect 1319 282 1322 290
rect 1324 282 1325 290
rect 1337 282 1338 290
rect 1340 282 1341 290
rect 795 226 796 234
rect 798 226 801 234
rect 803 226 804 234
rect 816 226 817 234
rect 819 230 820 234
rect 819 226 824 230
rect 832 226 833 234
rect 835 226 838 234
rect 840 226 841 234
rect 858 226 859 234
rect 861 226 862 234
rect 874 226 875 234
rect 877 230 878 234
rect 877 226 882 230
rect 890 226 891 234
rect 893 226 896 234
rect 898 226 899 234
rect 911 226 912 234
rect 914 226 915 234
rect 1728 226 1729 234
rect 1731 226 1734 234
rect 1736 226 1737 234
rect 1749 226 1750 234
rect 1752 230 1753 234
rect 1752 226 1757 230
rect 1765 226 1766 234
rect 1768 226 1771 234
rect 1773 226 1774 234
rect 1791 226 1792 234
rect 1794 226 1795 234
rect 1807 226 1808 234
rect 1810 230 1811 234
rect 1810 226 1815 230
rect 1823 226 1824 234
rect 1826 226 1829 234
rect 1831 226 1832 234
rect 1844 226 1845 234
rect 1847 226 1848 234
rect 24 196 25 204
rect 27 196 30 204
rect 32 196 33 204
rect 45 196 46 204
rect 48 200 49 204
rect 48 196 53 200
rect 61 196 62 204
rect 64 196 67 204
rect 69 196 70 204
rect 87 196 88 204
rect 90 196 91 204
rect 103 196 104 204
rect 106 200 107 204
rect 106 196 111 200
rect 119 196 120 204
rect 122 196 125 204
rect 127 196 128 204
rect 140 196 141 204
rect 143 196 144 204
rect 156 196 157 204
rect 159 196 162 204
rect 164 196 165 204
rect 177 196 178 204
rect 180 200 181 204
rect 180 196 185 200
rect 193 196 194 204
rect 196 196 199 204
rect 201 196 202 204
rect 219 196 220 204
rect 222 196 223 204
rect 235 196 236 204
rect 238 200 239 204
rect 238 196 243 200
rect 251 196 252 204
rect 254 196 257 204
rect 259 196 260 204
rect 272 196 273 204
rect 275 196 276 204
rect 288 196 289 204
rect 291 196 294 204
rect 296 196 297 204
rect 309 196 310 204
rect 312 200 313 204
rect 312 196 317 200
rect 325 196 326 204
rect 328 196 331 204
rect 333 196 334 204
rect 351 196 352 204
rect 354 196 355 204
rect 367 196 368 204
rect 370 200 371 204
rect 370 196 375 200
rect 383 196 384 204
rect 386 196 389 204
rect 391 196 392 204
rect 404 196 405 204
rect 407 196 408 204
rect 957 196 958 204
rect 960 196 963 204
rect 965 196 966 204
rect 978 196 979 204
rect 981 200 982 204
rect 981 196 986 200
rect 994 196 995 204
rect 997 196 1000 204
rect 1002 196 1003 204
rect 1020 196 1021 204
rect 1023 196 1024 204
rect 1036 196 1037 204
rect 1039 200 1040 204
rect 1039 196 1044 200
rect 1052 196 1053 204
rect 1055 196 1058 204
rect 1060 196 1061 204
rect 1073 196 1074 204
rect 1076 196 1077 204
rect 1089 196 1090 204
rect 1092 196 1095 204
rect 1097 196 1098 204
rect 1110 196 1111 204
rect 1113 200 1114 204
rect 1113 196 1118 200
rect 1126 196 1127 204
rect 1129 196 1132 204
rect 1134 196 1135 204
rect 1152 196 1153 204
rect 1155 196 1156 204
rect 1168 196 1169 204
rect 1171 200 1172 204
rect 1171 196 1176 200
rect 1184 196 1185 204
rect 1187 196 1190 204
rect 1192 196 1193 204
rect 1205 196 1206 204
rect 1208 196 1209 204
rect 1221 196 1222 204
rect 1224 196 1227 204
rect 1229 196 1230 204
rect 1242 196 1243 204
rect 1245 200 1246 204
rect 1245 196 1250 200
rect 1258 196 1259 204
rect 1261 196 1264 204
rect 1266 196 1267 204
rect 1284 196 1285 204
rect 1287 196 1288 204
rect 1300 196 1301 204
rect 1303 200 1304 204
rect 1303 196 1308 200
rect 1316 196 1317 204
rect 1319 196 1322 204
rect 1324 196 1325 204
rect 1337 196 1338 204
rect 1340 196 1341 204
rect 24 56 25 64
rect 27 56 30 64
rect 32 56 33 64
rect 45 56 46 64
rect 48 60 49 64
rect 48 56 53 60
rect 61 56 62 64
rect 64 56 67 64
rect 69 56 70 64
rect 87 56 88 64
rect 90 56 91 64
rect 103 56 104 64
rect 106 60 107 64
rect 106 56 111 60
rect 119 56 120 64
rect 122 56 125 64
rect 127 56 128 64
rect 140 56 141 64
rect 143 56 144 64
rect 156 56 157 64
rect 159 56 162 64
rect 164 56 165 64
rect 177 56 178 64
rect 180 60 181 64
rect 180 56 185 60
rect 193 56 194 64
rect 196 56 199 64
rect 201 56 202 64
rect 219 56 220 64
rect 222 56 223 64
rect 235 56 236 64
rect 238 60 239 64
rect 238 56 243 60
rect 251 56 252 64
rect 254 56 257 64
rect 259 56 260 64
rect 272 56 273 64
rect 275 56 276 64
rect 288 56 289 64
rect 291 56 294 64
rect 296 56 297 64
rect 309 56 310 64
rect 312 60 313 64
rect 312 56 317 60
rect 325 56 326 64
rect 328 56 331 64
rect 333 56 334 64
rect 351 56 352 64
rect 354 56 355 64
rect 367 56 368 64
rect 370 60 371 64
rect 370 56 375 60
rect 383 56 384 64
rect 386 56 389 64
rect 391 56 392 64
rect 404 56 405 64
rect 407 56 408 64
rect 957 56 958 64
rect 960 56 963 64
rect 965 56 966 64
rect 978 56 979 64
rect 981 60 982 64
rect 981 56 986 60
rect 994 56 995 64
rect 997 56 1000 64
rect 1002 56 1003 64
rect 1020 56 1021 64
rect 1023 56 1024 64
rect 1036 56 1037 64
rect 1039 60 1040 64
rect 1039 56 1044 60
rect 1052 56 1053 64
rect 1055 56 1058 64
rect 1060 56 1061 64
rect 1073 56 1074 64
rect 1076 56 1077 64
rect 1089 56 1090 64
rect 1092 56 1095 64
rect 1097 56 1098 64
rect 1110 56 1111 64
rect 1113 60 1114 64
rect 1113 56 1118 60
rect 1126 56 1127 64
rect 1129 56 1132 64
rect 1134 56 1135 64
rect 1152 56 1153 64
rect 1155 56 1156 64
rect 1168 56 1169 64
rect 1171 60 1172 64
rect 1171 56 1176 60
rect 1184 56 1185 64
rect 1187 56 1190 64
rect 1192 56 1193 64
rect 1205 56 1206 64
rect 1208 56 1209 64
rect 1221 56 1222 64
rect 1224 56 1227 64
rect 1229 56 1230 64
rect 1242 56 1243 64
rect 1245 60 1246 64
rect 1245 56 1250 60
rect 1258 56 1259 64
rect 1261 56 1264 64
rect 1266 56 1267 64
rect 1284 56 1285 64
rect 1287 56 1288 64
rect 1300 56 1301 64
rect 1303 60 1304 64
rect 1303 56 1308 60
rect 1316 56 1317 64
rect 1319 56 1322 64
rect 1324 56 1325 64
rect 1337 56 1338 64
rect 1340 56 1341 64
<< ndcontact >>
rect 492 1914 496 1918
rect 505 1914 509 1918
rect 513 1914 517 1918
rect 521 1914 525 1918
rect 529 1914 533 1918
rect 542 1914 546 1918
rect 555 1914 559 1918
rect 563 1914 567 1918
rect 571 1914 575 1918
rect 579 1914 583 1918
rect 587 1914 591 1918
rect 600 1914 604 1918
rect 608 1914 612 1918
rect 616 1914 620 1918
rect 624 1914 628 1918
rect 637 1914 641 1918
rect 645 1914 649 1918
rect 653 1914 657 1918
rect 661 1914 665 1918
rect 674 1914 678 1918
rect 687 1914 691 1918
rect 695 1914 699 1918
rect 703 1914 707 1918
rect 711 1914 715 1918
rect 719 1914 723 1918
rect 732 1914 736 1918
rect 740 1914 744 1918
rect 748 1914 752 1918
rect 756 1914 760 1918
rect 769 1914 773 1918
rect 777 1914 781 1918
rect 785 1914 789 1918
rect 793 1914 797 1918
rect 806 1914 810 1918
rect 819 1914 823 1918
rect 827 1914 831 1918
rect 835 1914 839 1918
rect 843 1914 847 1918
rect 851 1914 855 1918
rect 864 1914 868 1918
rect 872 1914 876 1918
rect 880 1914 884 1918
rect 888 1914 892 1918
rect 901 1914 905 1918
rect 909 1914 913 1918
rect 917 1914 921 1918
rect 925 1914 929 1918
rect 938 1914 942 1918
rect 951 1914 955 1918
rect 959 1914 963 1918
rect 967 1914 971 1918
rect 975 1914 979 1918
rect 983 1914 987 1918
rect 996 1914 1000 1918
rect 1004 1914 1008 1918
rect 1012 1914 1016 1918
rect 1425 1914 1429 1918
rect 1438 1914 1442 1918
rect 1446 1914 1450 1918
rect 1454 1914 1458 1918
rect 1462 1914 1466 1918
rect 1475 1914 1479 1918
rect 1488 1914 1492 1918
rect 1496 1914 1500 1918
rect 1504 1914 1508 1918
rect 1512 1914 1516 1918
rect 1520 1914 1524 1918
rect 1533 1914 1537 1918
rect 1541 1914 1545 1918
rect 1549 1914 1553 1918
rect 1557 1914 1561 1918
rect 1570 1914 1574 1918
rect 1578 1914 1582 1918
rect 1586 1914 1590 1918
rect 1594 1914 1598 1918
rect 1607 1914 1611 1918
rect 1620 1914 1624 1918
rect 1628 1914 1632 1918
rect 1636 1914 1640 1918
rect 1644 1914 1648 1918
rect 1652 1914 1656 1918
rect 1665 1914 1669 1918
rect 1673 1914 1677 1918
rect 1681 1914 1685 1918
rect 1689 1914 1693 1918
rect 1702 1914 1706 1918
rect 1710 1914 1714 1918
rect 1718 1914 1722 1918
rect 1726 1914 1730 1918
rect 1739 1914 1743 1918
rect 1752 1914 1756 1918
rect 1760 1914 1764 1918
rect 1768 1914 1772 1918
rect 1776 1914 1780 1918
rect 1784 1914 1788 1918
rect 1797 1914 1801 1918
rect 1805 1914 1809 1918
rect 1813 1914 1817 1918
rect 1821 1914 1825 1918
rect 1834 1914 1838 1918
rect 1842 1914 1846 1918
rect 1850 1914 1854 1918
rect 1858 1914 1862 1918
rect 1871 1914 1875 1918
rect 1884 1914 1888 1918
rect 1892 1914 1896 1918
rect 1900 1914 1904 1918
rect 1908 1914 1912 1918
rect 1916 1914 1920 1918
rect 1929 1914 1933 1918
rect 1937 1914 1941 1918
rect 1945 1914 1949 1918
rect 152 1881 156 1885
rect 165 1881 169 1885
rect 173 1881 177 1885
rect 181 1881 185 1885
rect 189 1881 193 1885
rect 202 1881 206 1885
rect 215 1881 219 1885
rect 223 1881 227 1885
rect 231 1881 235 1885
rect 239 1881 243 1885
rect 247 1881 251 1885
rect 260 1881 264 1885
rect 268 1881 272 1885
rect 276 1881 280 1885
rect 1085 1881 1089 1885
rect 1098 1881 1102 1885
rect 1106 1881 1110 1885
rect 1114 1881 1118 1885
rect 1122 1881 1126 1885
rect 1135 1881 1139 1885
rect 1148 1881 1152 1885
rect 1156 1881 1160 1885
rect 1164 1881 1168 1885
rect 1172 1881 1176 1885
rect 1180 1881 1184 1885
rect 1193 1881 1197 1885
rect 1201 1881 1205 1885
rect 1209 1881 1213 1885
rect 276 1844 280 1848
rect 284 1844 288 1848
rect 671 1848 675 1852
rect 679 1848 683 1852
rect 695 1844 699 1848
rect 710 1844 714 1848
rect 752 1848 756 1852
rect 760 1848 764 1852
rect 776 1844 780 1848
rect 791 1844 795 1848
rect 725 1840 729 1844
rect 733 1840 737 1844
rect 159 1835 163 1839
rect 167 1835 171 1839
rect 497 1835 501 1839
rect 505 1835 509 1839
rect 513 1835 517 1839
rect 521 1835 525 1839
rect 529 1835 533 1839
rect 537 1835 541 1839
rect 548 1835 552 1839
rect 565 1835 569 1839
rect 582 1835 586 1839
rect 591 1835 595 1839
rect 604 1835 608 1839
rect 612 1835 616 1839
rect 620 1835 624 1839
rect 637 1835 641 1839
rect 647 1835 651 1839
rect 655 1835 659 1839
rect 806 1840 810 1844
rect 814 1840 818 1844
rect 1209 1844 1213 1848
rect 1217 1844 1221 1848
rect 1604 1848 1608 1852
rect 1612 1848 1616 1852
rect 1628 1844 1632 1848
rect 1643 1844 1647 1848
rect 1685 1848 1689 1852
rect 1693 1848 1697 1852
rect 1709 1844 1713 1848
rect 1724 1844 1728 1848
rect 1658 1840 1662 1844
rect 1666 1840 1670 1844
rect 1092 1835 1096 1839
rect 1100 1835 1104 1839
rect 1430 1835 1434 1839
rect 1438 1835 1442 1839
rect 1446 1835 1450 1839
rect 1454 1835 1458 1839
rect 1462 1835 1466 1839
rect 1470 1835 1474 1839
rect 1481 1835 1485 1839
rect 1498 1835 1502 1839
rect 1515 1835 1519 1839
rect 1524 1835 1528 1839
rect 1537 1835 1541 1839
rect 1545 1835 1549 1839
rect 1553 1835 1557 1839
rect 1570 1835 1574 1839
rect 1580 1835 1584 1839
rect 1588 1835 1592 1839
rect 1739 1840 1743 1844
rect 1747 1840 1751 1844
rect 497 1789 501 1793
rect 505 1789 509 1793
rect 513 1789 517 1793
rect 521 1789 525 1793
rect 529 1789 533 1793
rect 537 1789 541 1793
rect 548 1789 552 1793
rect 565 1789 569 1793
rect 582 1789 586 1793
rect 591 1789 595 1793
rect 604 1789 608 1793
rect 612 1789 616 1793
rect 620 1789 624 1793
rect 637 1789 641 1793
rect 647 1789 651 1793
rect 655 1789 659 1793
rect 143 1779 147 1783
rect 151 1779 155 1783
rect 159 1779 163 1783
rect 172 1779 176 1783
rect 180 1779 184 1783
rect 188 1779 192 1783
rect 196 1779 200 1783
rect 204 1779 208 1783
rect 217 1779 221 1783
rect 230 1779 234 1783
rect 238 1779 242 1783
rect 246 1779 250 1783
rect 254 1779 258 1783
rect 267 1779 271 1783
rect 695 1788 699 1792
rect 710 1788 714 1792
rect 776 1788 780 1792
rect 791 1788 795 1792
rect 1430 1789 1434 1793
rect 1438 1789 1442 1793
rect 1446 1789 1450 1793
rect 1454 1789 1458 1793
rect 1462 1789 1466 1793
rect 1470 1789 1474 1793
rect 1481 1789 1485 1793
rect 1498 1789 1502 1793
rect 1515 1789 1519 1793
rect 1524 1789 1528 1793
rect 1537 1789 1541 1793
rect 1545 1789 1549 1793
rect 1553 1789 1557 1793
rect 1570 1789 1574 1793
rect 1580 1789 1584 1793
rect 1588 1789 1592 1793
rect 1076 1779 1080 1783
rect 1084 1779 1088 1783
rect 1092 1779 1096 1783
rect 1105 1779 1109 1783
rect 1113 1779 1117 1783
rect 1121 1779 1125 1783
rect 1129 1779 1133 1783
rect 1137 1779 1141 1783
rect 1150 1779 1154 1783
rect 1163 1779 1167 1783
rect 1171 1779 1175 1783
rect 1179 1779 1183 1783
rect 1187 1779 1191 1783
rect 1200 1779 1204 1783
rect 1628 1788 1632 1792
rect 1643 1788 1647 1792
rect 1709 1788 1713 1792
rect 1724 1788 1728 1792
rect 695 1712 699 1716
rect 710 1712 714 1716
rect 776 1716 780 1720
rect 784 1716 788 1720
rect 800 1712 804 1716
rect 815 1712 819 1716
rect 725 1708 729 1712
rect 733 1708 737 1712
rect 497 1703 501 1707
rect 505 1703 509 1707
rect 513 1703 517 1707
rect 521 1703 525 1707
rect 529 1703 533 1707
rect 537 1703 541 1707
rect 548 1703 552 1707
rect 565 1703 569 1707
rect 582 1703 586 1707
rect 591 1703 595 1707
rect 604 1703 608 1707
rect 612 1703 616 1707
rect 620 1703 624 1707
rect 637 1703 641 1707
rect 647 1703 651 1707
rect 655 1703 659 1707
rect 830 1708 834 1712
rect 838 1708 842 1712
rect 1628 1712 1632 1716
rect 1643 1712 1647 1716
rect 1709 1716 1713 1720
rect 1717 1716 1721 1720
rect 1733 1712 1737 1716
rect 1748 1712 1752 1716
rect 1658 1708 1662 1712
rect 1666 1708 1670 1712
rect 1430 1703 1434 1707
rect 1438 1703 1442 1707
rect 1446 1703 1450 1707
rect 1454 1703 1458 1707
rect 1462 1703 1466 1707
rect 1470 1703 1474 1707
rect 1481 1703 1485 1707
rect 1498 1703 1502 1707
rect 1515 1703 1519 1707
rect 1524 1703 1528 1707
rect 1537 1703 1541 1707
rect 1545 1703 1549 1707
rect 1553 1703 1557 1707
rect 1570 1703 1574 1707
rect 1580 1703 1584 1707
rect 1588 1703 1592 1707
rect 1763 1708 1767 1712
rect 1771 1708 1775 1712
rect 497 1657 501 1661
rect 505 1657 509 1661
rect 513 1657 517 1661
rect 521 1657 525 1661
rect 529 1657 533 1661
rect 537 1657 541 1661
rect 548 1657 552 1661
rect 565 1657 569 1661
rect 582 1657 586 1661
rect 591 1657 595 1661
rect 604 1657 608 1661
rect 612 1657 616 1661
rect 620 1657 624 1661
rect 637 1657 641 1661
rect 647 1657 651 1661
rect 655 1657 659 1661
rect 695 1657 699 1661
rect 710 1657 714 1661
rect 800 1657 804 1661
rect 815 1657 819 1661
rect 1430 1657 1434 1661
rect 1438 1657 1442 1661
rect 1446 1657 1450 1661
rect 1454 1657 1458 1661
rect 1462 1657 1466 1661
rect 1470 1657 1474 1661
rect 1481 1657 1485 1661
rect 1498 1657 1502 1661
rect 1515 1657 1519 1661
rect 1524 1657 1528 1661
rect 1537 1657 1541 1661
rect 1545 1657 1549 1661
rect 1553 1657 1557 1661
rect 1570 1657 1574 1661
rect 1580 1657 1584 1661
rect 1588 1657 1592 1661
rect 1628 1657 1632 1661
rect 1643 1657 1647 1661
rect 1733 1657 1737 1661
rect 1748 1657 1752 1661
rect 695 1580 699 1584
rect 710 1580 714 1584
rect 752 1584 756 1588
rect 760 1584 764 1588
rect 776 1580 780 1584
rect 791 1580 795 1584
rect 842 1584 846 1588
rect 850 1584 854 1588
rect 866 1580 870 1584
rect 881 1580 885 1584
rect 725 1576 729 1580
rect 733 1576 737 1580
rect 497 1571 501 1575
rect 505 1571 509 1575
rect 513 1571 517 1575
rect 521 1571 525 1575
rect 529 1571 533 1575
rect 537 1571 541 1575
rect 548 1571 552 1575
rect 565 1571 569 1575
rect 582 1571 586 1575
rect 591 1571 595 1575
rect 604 1571 608 1575
rect 612 1571 616 1575
rect 620 1571 624 1575
rect 637 1571 641 1575
rect 647 1571 651 1575
rect 655 1571 659 1575
rect 806 1576 810 1580
rect 814 1576 818 1580
rect 896 1576 900 1580
rect 904 1576 908 1580
rect 1628 1580 1632 1584
rect 1643 1580 1647 1584
rect 1685 1584 1689 1588
rect 1693 1584 1697 1588
rect 1709 1580 1713 1584
rect 1724 1580 1728 1584
rect 1775 1584 1779 1588
rect 1783 1584 1787 1588
rect 1799 1580 1803 1584
rect 1814 1580 1818 1584
rect 1658 1576 1662 1580
rect 1666 1576 1670 1580
rect 1430 1571 1434 1575
rect 1438 1571 1442 1575
rect 1446 1571 1450 1575
rect 1454 1571 1458 1575
rect 1462 1571 1466 1575
rect 1470 1571 1474 1575
rect 1481 1571 1485 1575
rect 1498 1571 1502 1575
rect 1515 1571 1519 1575
rect 1524 1571 1528 1575
rect 1537 1571 1541 1575
rect 1545 1571 1549 1575
rect 1553 1571 1557 1575
rect 1570 1571 1574 1575
rect 1580 1571 1584 1575
rect 1588 1571 1592 1575
rect 1739 1576 1743 1580
rect 1747 1576 1751 1580
rect 1829 1576 1833 1580
rect 1837 1576 1841 1580
rect 497 1525 501 1529
rect 505 1525 509 1529
rect 513 1525 517 1529
rect 521 1525 525 1529
rect 529 1525 533 1529
rect 537 1525 541 1529
rect 548 1525 552 1529
rect 565 1525 569 1529
rect 582 1525 586 1529
rect 591 1525 595 1529
rect 604 1525 608 1529
rect 612 1525 616 1529
rect 620 1525 624 1529
rect 637 1525 641 1529
rect 647 1525 651 1529
rect 655 1525 659 1529
rect 695 1522 699 1526
rect 710 1522 714 1526
rect 776 1522 780 1526
rect 791 1522 795 1526
rect 866 1522 870 1526
rect 881 1522 885 1526
rect 1430 1525 1434 1529
rect 1438 1525 1442 1529
rect 1446 1525 1450 1529
rect 1454 1525 1458 1529
rect 1462 1525 1466 1529
rect 1470 1525 1474 1529
rect 1481 1525 1485 1529
rect 1498 1525 1502 1529
rect 1515 1525 1519 1529
rect 1524 1525 1528 1529
rect 1537 1525 1541 1529
rect 1545 1525 1549 1529
rect 1553 1525 1557 1529
rect 1570 1525 1574 1529
rect 1580 1525 1584 1529
rect 1588 1525 1592 1529
rect 1628 1522 1632 1526
rect 1643 1522 1647 1526
rect 1709 1522 1713 1526
rect 1724 1522 1728 1526
rect 1799 1522 1803 1526
rect 1814 1522 1818 1526
rect 695 1448 699 1452
rect 710 1448 714 1452
rect 725 1444 729 1448
rect 733 1444 737 1448
rect 497 1439 501 1443
rect 505 1439 509 1443
rect 513 1439 517 1443
rect 521 1439 525 1443
rect 529 1439 533 1443
rect 537 1439 541 1443
rect 548 1439 552 1443
rect 565 1439 569 1443
rect 582 1439 586 1443
rect 591 1439 595 1443
rect 604 1439 608 1443
rect 612 1439 616 1443
rect 620 1439 624 1443
rect 637 1439 641 1443
rect 647 1439 651 1443
rect 655 1439 659 1443
rect 1628 1448 1632 1452
rect 1643 1448 1647 1452
rect 1658 1444 1662 1448
rect 1666 1444 1670 1448
rect 1430 1439 1434 1443
rect 1438 1439 1442 1443
rect 1446 1439 1450 1443
rect 1454 1439 1458 1443
rect 1462 1439 1466 1443
rect 1470 1439 1474 1443
rect 1481 1439 1485 1443
rect 1498 1439 1502 1443
rect 1515 1439 1519 1443
rect 1524 1439 1528 1443
rect 1537 1439 1541 1443
rect 1545 1439 1549 1443
rect 1553 1439 1557 1443
rect 1570 1439 1574 1443
rect 1580 1439 1584 1443
rect 1588 1439 1592 1443
rect 497 1393 501 1397
rect 505 1393 509 1397
rect 513 1393 517 1397
rect 521 1393 525 1397
rect 529 1393 533 1397
rect 537 1393 541 1397
rect 548 1393 552 1397
rect 565 1393 569 1397
rect 582 1393 586 1397
rect 591 1393 595 1397
rect 604 1393 608 1397
rect 612 1393 616 1397
rect 620 1393 624 1397
rect 637 1393 641 1397
rect 647 1393 651 1397
rect 655 1393 659 1397
rect 731 1393 735 1397
rect 739 1393 743 1397
rect 749 1393 753 1397
rect 757 1393 761 1397
rect 766 1393 770 1397
rect 774 1393 778 1397
rect 782 1393 786 1397
rect 790 1393 794 1397
rect 798 1393 802 1397
rect 809 1393 813 1397
rect 826 1393 830 1397
rect 843 1393 847 1397
rect 852 1393 856 1397
rect 865 1393 869 1397
rect 873 1393 877 1397
rect 881 1393 885 1397
rect 898 1393 902 1397
rect 908 1393 912 1397
rect 916 1393 920 1397
rect 20 1379 24 1383
rect 33 1379 37 1383
rect 41 1379 45 1383
rect 49 1379 53 1383
rect 57 1379 61 1383
rect 70 1379 74 1383
rect 83 1379 87 1383
rect 91 1379 95 1383
rect 99 1379 103 1383
rect 107 1379 111 1383
rect 115 1379 119 1383
rect 128 1379 132 1383
rect 136 1379 140 1383
rect 144 1379 148 1383
rect 152 1379 156 1383
rect 165 1379 169 1383
rect 173 1379 177 1383
rect 181 1379 185 1383
rect 189 1379 193 1383
rect 202 1379 206 1383
rect 215 1379 219 1383
rect 223 1379 227 1383
rect 231 1379 235 1383
rect 239 1379 243 1383
rect 247 1379 251 1383
rect 260 1379 264 1383
rect 268 1379 272 1383
rect 276 1379 280 1383
rect 284 1379 288 1383
rect 297 1379 301 1383
rect 305 1379 309 1383
rect 313 1379 317 1383
rect 321 1379 325 1383
rect 334 1379 338 1383
rect 347 1379 351 1383
rect 355 1379 359 1383
rect 363 1379 367 1383
rect 371 1379 375 1383
rect 379 1379 383 1383
rect 392 1379 396 1383
rect 400 1379 404 1383
rect 408 1379 412 1383
rect 695 1386 699 1390
rect 710 1386 714 1390
rect 1430 1393 1434 1397
rect 1438 1393 1442 1397
rect 1446 1393 1450 1397
rect 1454 1393 1458 1397
rect 1462 1393 1466 1397
rect 1470 1393 1474 1397
rect 1481 1393 1485 1397
rect 1498 1393 1502 1397
rect 1515 1393 1519 1397
rect 1524 1393 1528 1397
rect 1537 1393 1541 1397
rect 1545 1393 1549 1397
rect 1553 1393 1557 1397
rect 1570 1393 1574 1397
rect 1580 1393 1584 1397
rect 1588 1393 1592 1397
rect 1664 1393 1668 1397
rect 1672 1393 1676 1397
rect 1682 1393 1686 1397
rect 1690 1393 1694 1397
rect 1699 1393 1703 1397
rect 1707 1393 1711 1397
rect 1715 1393 1719 1397
rect 1723 1393 1727 1397
rect 1731 1393 1735 1397
rect 1742 1393 1746 1397
rect 1759 1393 1763 1397
rect 1776 1393 1780 1397
rect 1785 1393 1789 1397
rect 1798 1393 1802 1397
rect 1806 1393 1810 1397
rect 1814 1393 1818 1397
rect 1831 1393 1835 1397
rect 1841 1393 1845 1397
rect 1849 1393 1853 1397
rect 953 1379 957 1383
rect 966 1379 970 1383
rect 974 1379 978 1383
rect 982 1379 986 1383
rect 990 1379 994 1383
rect 1003 1379 1007 1383
rect 1016 1379 1020 1383
rect 1024 1379 1028 1383
rect 1032 1379 1036 1383
rect 1040 1379 1044 1383
rect 1048 1379 1052 1383
rect 1061 1379 1065 1383
rect 1069 1379 1073 1383
rect 1077 1379 1081 1383
rect 1085 1379 1089 1383
rect 1098 1379 1102 1383
rect 1106 1379 1110 1383
rect 1114 1379 1118 1383
rect 1122 1379 1126 1383
rect 1135 1379 1139 1383
rect 1148 1379 1152 1383
rect 1156 1379 1160 1383
rect 1164 1379 1168 1383
rect 1172 1379 1176 1383
rect 1180 1379 1184 1383
rect 1193 1379 1197 1383
rect 1201 1379 1205 1383
rect 1209 1379 1213 1383
rect 1217 1379 1221 1383
rect 1230 1379 1234 1383
rect 1238 1379 1242 1383
rect 1246 1379 1250 1383
rect 1254 1379 1258 1383
rect 1267 1379 1271 1383
rect 1280 1379 1284 1383
rect 1288 1379 1292 1383
rect 1296 1379 1300 1383
rect 1304 1379 1308 1383
rect 1312 1379 1316 1383
rect 1325 1379 1329 1383
rect 1333 1379 1337 1383
rect 1341 1379 1345 1383
rect 1628 1386 1632 1390
rect 1643 1386 1647 1390
rect 925 1340 929 1344
rect 135 1335 139 1339
rect 143 1335 147 1339
rect 159 1335 163 1339
rect 167 1335 171 1339
rect 1858 1340 1862 1344
rect 925 1332 929 1336
rect 1068 1335 1072 1339
rect 1076 1335 1080 1339
rect 1092 1335 1096 1339
rect 1100 1335 1104 1339
rect 1858 1332 1862 1336
rect 155 1324 159 1328
rect 163 1324 167 1328
rect 1088 1324 1092 1328
rect 1096 1324 1100 1328
rect 151 1313 155 1317
rect 1084 1313 1088 1317
rect 151 1305 155 1309
rect 135 1301 139 1305
rect 143 1301 147 1305
rect 159 1301 163 1305
rect 167 1301 171 1305
rect 1084 1305 1088 1309
rect 1068 1301 1072 1305
rect 1076 1301 1080 1305
rect 1092 1301 1096 1305
rect 1100 1301 1104 1305
rect 791 1269 795 1273
rect 804 1269 808 1273
rect 812 1269 816 1273
rect 820 1269 824 1273
rect 828 1269 832 1273
rect 841 1269 845 1273
rect 854 1269 858 1273
rect 862 1269 866 1273
rect 870 1269 874 1273
rect 878 1269 882 1273
rect 886 1269 890 1273
rect 899 1269 903 1273
rect 907 1269 911 1273
rect 915 1269 919 1273
rect 1724 1269 1728 1273
rect 1737 1269 1741 1273
rect 1745 1269 1749 1273
rect 1753 1269 1757 1273
rect 1761 1269 1765 1273
rect 1774 1269 1778 1273
rect 1787 1269 1791 1273
rect 1795 1269 1799 1273
rect 1803 1269 1807 1273
rect 1811 1269 1815 1273
rect 1819 1269 1823 1273
rect 1832 1269 1836 1273
rect 1840 1269 1844 1273
rect 1848 1269 1852 1273
rect 20 1239 24 1243
rect 33 1239 37 1243
rect 41 1239 45 1243
rect 49 1239 53 1243
rect 57 1239 61 1243
rect 70 1239 74 1243
rect 83 1239 87 1243
rect 91 1239 95 1243
rect 99 1239 103 1243
rect 107 1239 111 1243
rect 115 1239 119 1243
rect 128 1239 132 1243
rect 136 1239 140 1243
rect 144 1239 148 1243
rect 152 1239 156 1243
rect 165 1239 169 1243
rect 173 1239 177 1243
rect 181 1239 185 1243
rect 189 1239 193 1243
rect 202 1239 206 1243
rect 215 1239 219 1243
rect 223 1239 227 1243
rect 231 1239 235 1243
rect 239 1239 243 1243
rect 247 1239 251 1243
rect 260 1239 264 1243
rect 268 1239 272 1243
rect 276 1239 280 1243
rect 284 1239 288 1243
rect 297 1239 301 1243
rect 305 1239 309 1243
rect 313 1239 317 1243
rect 321 1239 325 1243
rect 334 1239 338 1243
rect 347 1239 351 1243
rect 355 1239 359 1243
rect 363 1239 367 1243
rect 371 1239 375 1243
rect 379 1239 383 1243
rect 392 1239 396 1243
rect 400 1239 404 1243
rect 408 1239 412 1243
rect 953 1239 957 1243
rect 966 1239 970 1243
rect 974 1239 978 1243
rect 982 1239 986 1243
rect 990 1239 994 1243
rect 1003 1239 1007 1243
rect 1016 1239 1020 1243
rect 1024 1239 1028 1243
rect 1032 1239 1036 1243
rect 1040 1239 1044 1243
rect 1048 1239 1052 1243
rect 1061 1239 1065 1243
rect 1069 1239 1073 1243
rect 1077 1239 1081 1243
rect 1085 1239 1089 1243
rect 1098 1239 1102 1243
rect 1106 1239 1110 1243
rect 1114 1239 1118 1243
rect 1122 1239 1126 1243
rect 1135 1239 1139 1243
rect 1148 1239 1152 1243
rect 1156 1239 1160 1243
rect 1164 1239 1168 1243
rect 1172 1239 1176 1243
rect 1180 1239 1184 1243
rect 1193 1239 1197 1243
rect 1201 1239 1205 1243
rect 1209 1239 1213 1243
rect 1217 1239 1221 1243
rect 1230 1239 1234 1243
rect 1238 1239 1242 1243
rect 1246 1239 1250 1243
rect 1254 1239 1258 1243
rect 1267 1239 1271 1243
rect 1280 1239 1284 1243
rect 1288 1239 1292 1243
rect 1296 1239 1300 1243
rect 1304 1239 1308 1243
rect 1312 1239 1316 1243
rect 1325 1239 1329 1243
rect 1333 1239 1337 1243
rect 1341 1239 1345 1243
rect 937 1196 941 1200
rect 937 1188 941 1192
rect 1870 1196 1874 1200
rect 1870 1188 1874 1192
rect 791 1183 795 1187
rect 804 1183 808 1187
rect 812 1183 816 1187
rect 820 1183 824 1187
rect 828 1183 832 1187
rect 841 1183 845 1187
rect 854 1183 858 1187
rect 862 1183 866 1187
rect 870 1183 874 1187
rect 878 1183 882 1187
rect 886 1183 890 1187
rect 899 1183 903 1187
rect 907 1183 911 1187
rect 915 1183 919 1187
rect 1724 1183 1728 1187
rect 1737 1183 1741 1187
rect 1745 1183 1749 1187
rect 1753 1183 1757 1187
rect 1761 1183 1765 1187
rect 1774 1183 1778 1187
rect 1787 1183 1791 1187
rect 1795 1183 1799 1187
rect 1803 1183 1807 1187
rect 1811 1183 1815 1187
rect 1819 1183 1823 1187
rect 1832 1183 1836 1187
rect 1840 1183 1844 1187
rect 1848 1183 1852 1187
rect 20 1153 24 1157
rect 33 1153 37 1157
rect 41 1153 45 1157
rect 49 1153 53 1157
rect 57 1153 61 1157
rect 70 1153 74 1157
rect 83 1153 87 1157
rect 91 1153 95 1157
rect 99 1153 103 1157
rect 107 1153 111 1157
rect 115 1153 119 1157
rect 128 1153 132 1157
rect 136 1153 140 1157
rect 144 1153 148 1157
rect 152 1153 156 1157
rect 165 1153 169 1157
rect 173 1153 177 1157
rect 181 1153 185 1157
rect 189 1153 193 1157
rect 202 1153 206 1157
rect 215 1153 219 1157
rect 223 1153 227 1157
rect 231 1153 235 1157
rect 239 1153 243 1157
rect 247 1153 251 1157
rect 260 1153 264 1157
rect 268 1153 272 1157
rect 276 1153 280 1157
rect 284 1153 288 1157
rect 297 1153 301 1157
rect 305 1153 309 1157
rect 313 1153 317 1157
rect 321 1153 325 1157
rect 334 1153 338 1157
rect 347 1153 351 1157
rect 355 1153 359 1157
rect 363 1153 367 1157
rect 371 1153 375 1157
rect 379 1153 383 1157
rect 392 1153 396 1157
rect 400 1153 404 1157
rect 408 1153 412 1157
rect 953 1153 957 1157
rect 966 1153 970 1157
rect 974 1153 978 1157
rect 982 1153 986 1157
rect 990 1153 994 1157
rect 1003 1153 1007 1157
rect 1016 1153 1020 1157
rect 1024 1153 1028 1157
rect 1032 1153 1036 1157
rect 1040 1153 1044 1157
rect 1048 1153 1052 1157
rect 1061 1153 1065 1157
rect 1069 1153 1073 1157
rect 1077 1153 1081 1157
rect 1085 1153 1089 1157
rect 1098 1153 1102 1157
rect 1106 1153 1110 1157
rect 1114 1153 1118 1157
rect 1122 1153 1126 1157
rect 1135 1153 1139 1157
rect 1148 1153 1152 1157
rect 1156 1153 1160 1157
rect 1164 1153 1168 1157
rect 1172 1153 1176 1157
rect 1180 1153 1184 1157
rect 1193 1153 1197 1157
rect 1201 1153 1205 1157
rect 1209 1153 1213 1157
rect 1217 1153 1221 1157
rect 1230 1153 1234 1157
rect 1238 1153 1242 1157
rect 1246 1153 1250 1157
rect 1254 1153 1258 1157
rect 1267 1153 1271 1157
rect 1280 1153 1284 1157
rect 1288 1153 1292 1157
rect 1296 1153 1300 1157
rect 1304 1153 1308 1157
rect 1312 1153 1316 1157
rect 1325 1153 1329 1157
rect 1333 1153 1337 1157
rect 1341 1153 1345 1157
rect 252 1109 256 1113
rect 260 1109 264 1113
rect 276 1109 280 1113
rect 284 1109 288 1113
rect 1185 1109 1189 1113
rect 1193 1109 1197 1113
rect 1209 1109 1213 1113
rect 1217 1109 1221 1113
rect 272 1098 276 1102
rect 280 1098 284 1102
rect 1205 1098 1209 1102
rect 1213 1098 1217 1102
rect 268 1087 272 1091
rect 1201 1087 1205 1091
rect 268 1079 272 1083
rect 1201 1079 1205 1083
rect 252 1075 256 1079
rect 260 1075 264 1079
rect 276 1075 280 1079
rect 284 1075 288 1079
rect 1185 1075 1189 1079
rect 1193 1075 1197 1079
rect 1209 1075 1213 1079
rect 1217 1075 1221 1079
rect 20 1013 24 1017
rect 33 1013 37 1017
rect 41 1013 45 1017
rect 49 1013 53 1017
rect 57 1013 61 1017
rect 70 1013 74 1017
rect 83 1013 87 1017
rect 91 1013 95 1017
rect 99 1013 103 1017
rect 107 1013 111 1017
rect 115 1013 119 1017
rect 128 1013 132 1017
rect 136 1013 140 1017
rect 144 1013 148 1017
rect 152 1013 156 1017
rect 165 1013 169 1017
rect 173 1013 177 1017
rect 181 1013 185 1017
rect 189 1013 193 1017
rect 202 1013 206 1017
rect 215 1013 219 1017
rect 223 1013 227 1017
rect 231 1013 235 1017
rect 239 1013 243 1017
rect 247 1013 251 1017
rect 260 1013 264 1017
rect 268 1013 272 1017
rect 276 1013 280 1017
rect 284 1013 288 1017
rect 297 1013 301 1017
rect 305 1013 309 1017
rect 313 1013 317 1017
rect 321 1013 325 1017
rect 334 1013 338 1017
rect 347 1013 351 1017
rect 355 1013 359 1017
rect 363 1013 367 1017
rect 371 1013 375 1017
rect 379 1013 383 1017
rect 392 1013 396 1017
rect 400 1013 404 1017
rect 408 1013 412 1017
rect 953 1013 957 1017
rect 966 1013 970 1017
rect 974 1013 978 1017
rect 982 1013 986 1017
rect 990 1013 994 1017
rect 1003 1013 1007 1017
rect 1016 1013 1020 1017
rect 1024 1013 1028 1017
rect 1032 1013 1036 1017
rect 1040 1013 1044 1017
rect 1048 1013 1052 1017
rect 1061 1013 1065 1017
rect 1069 1013 1073 1017
rect 1077 1013 1081 1017
rect 1085 1013 1089 1017
rect 1098 1013 1102 1017
rect 1106 1013 1110 1017
rect 1114 1013 1118 1017
rect 1122 1013 1126 1017
rect 1135 1013 1139 1017
rect 1148 1013 1152 1017
rect 1156 1013 1160 1017
rect 1164 1013 1168 1017
rect 1172 1013 1176 1017
rect 1180 1013 1184 1017
rect 1193 1013 1197 1017
rect 1201 1013 1205 1017
rect 1209 1013 1213 1017
rect 1217 1013 1221 1017
rect 1230 1013 1234 1017
rect 1238 1013 1242 1017
rect 1246 1013 1250 1017
rect 1254 1013 1258 1017
rect 1267 1013 1271 1017
rect 1280 1013 1284 1017
rect 1288 1013 1292 1017
rect 1296 1013 1300 1017
rect 1304 1013 1308 1017
rect 1312 1013 1316 1017
rect 1325 1013 1329 1017
rect 1333 1013 1337 1017
rect 1341 1013 1345 1017
rect 492 934 496 938
rect 505 934 509 938
rect 513 934 517 938
rect 521 934 525 938
rect 529 934 533 938
rect 542 934 546 938
rect 555 934 559 938
rect 563 934 567 938
rect 571 934 575 938
rect 579 934 583 938
rect 587 934 591 938
rect 600 934 604 938
rect 608 934 612 938
rect 616 934 620 938
rect 624 934 628 938
rect 637 934 641 938
rect 645 934 649 938
rect 653 934 657 938
rect 661 934 665 938
rect 674 934 678 938
rect 687 934 691 938
rect 695 934 699 938
rect 703 934 707 938
rect 711 934 715 938
rect 719 934 723 938
rect 732 934 736 938
rect 740 934 744 938
rect 748 934 752 938
rect 756 934 760 938
rect 769 934 773 938
rect 777 934 781 938
rect 785 934 789 938
rect 793 934 797 938
rect 806 934 810 938
rect 819 934 823 938
rect 827 934 831 938
rect 835 934 839 938
rect 843 934 847 938
rect 851 934 855 938
rect 864 934 868 938
rect 872 934 876 938
rect 880 934 884 938
rect 888 934 892 938
rect 901 934 905 938
rect 909 934 913 938
rect 917 934 921 938
rect 925 934 929 938
rect 938 934 942 938
rect 951 934 955 938
rect 959 934 963 938
rect 967 934 971 938
rect 975 934 979 938
rect 983 934 987 938
rect 996 934 1000 938
rect 1004 934 1008 938
rect 1012 934 1016 938
rect 1425 934 1429 938
rect 1438 934 1442 938
rect 1446 934 1450 938
rect 1454 934 1458 938
rect 1462 934 1466 938
rect 1475 934 1479 938
rect 1488 934 1492 938
rect 1496 934 1500 938
rect 1504 934 1508 938
rect 1512 934 1516 938
rect 1520 934 1524 938
rect 1533 934 1537 938
rect 1541 934 1545 938
rect 1549 934 1553 938
rect 1557 934 1561 938
rect 1570 934 1574 938
rect 1578 934 1582 938
rect 1586 934 1590 938
rect 1594 934 1598 938
rect 1607 934 1611 938
rect 1620 934 1624 938
rect 1628 934 1632 938
rect 1636 934 1640 938
rect 1644 934 1648 938
rect 1652 934 1656 938
rect 1665 934 1669 938
rect 1673 934 1677 938
rect 1681 934 1685 938
rect 1689 934 1693 938
rect 1702 934 1706 938
rect 1710 934 1714 938
rect 1718 934 1722 938
rect 1726 934 1730 938
rect 1739 934 1743 938
rect 1752 934 1756 938
rect 1760 934 1764 938
rect 1768 934 1772 938
rect 1776 934 1780 938
rect 1784 934 1788 938
rect 1797 934 1801 938
rect 1805 934 1809 938
rect 1813 934 1817 938
rect 1821 934 1825 938
rect 1834 934 1838 938
rect 1842 934 1846 938
rect 1850 934 1854 938
rect 1858 934 1862 938
rect 1871 934 1875 938
rect 1884 934 1888 938
rect 1892 934 1896 938
rect 1900 934 1904 938
rect 1908 934 1912 938
rect 1916 934 1920 938
rect 1929 934 1933 938
rect 1937 934 1941 938
rect 1945 934 1949 938
rect 152 901 156 905
rect 165 901 169 905
rect 173 901 177 905
rect 181 901 185 905
rect 189 901 193 905
rect 202 901 206 905
rect 215 901 219 905
rect 223 901 227 905
rect 231 901 235 905
rect 239 901 243 905
rect 247 901 251 905
rect 260 901 264 905
rect 268 901 272 905
rect 276 901 280 905
rect 1085 901 1089 905
rect 1098 901 1102 905
rect 1106 901 1110 905
rect 1114 901 1118 905
rect 1122 901 1126 905
rect 1135 901 1139 905
rect 1148 901 1152 905
rect 1156 901 1160 905
rect 1164 901 1168 905
rect 1172 901 1176 905
rect 1180 901 1184 905
rect 1193 901 1197 905
rect 1201 901 1205 905
rect 1209 901 1213 905
rect 276 864 280 868
rect 284 864 288 868
rect 671 868 675 872
rect 679 868 683 872
rect 695 864 699 868
rect 710 864 714 868
rect 752 868 756 872
rect 760 868 764 872
rect 776 864 780 868
rect 791 864 795 868
rect 725 860 729 864
rect 733 860 737 864
rect 159 855 163 859
rect 167 855 171 859
rect 497 855 501 859
rect 505 855 509 859
rect 513 855 517 859
rect 521 855 525 859
rect 529 855 533 859
rect 537 855 541 859
rect 548 855 552 859
rect 565 855 569 859
rect 582 855 586 859
rect 591 855 595 859
rect 604 855 608 859
rect 612 855 616 859
rect 620 855 624 859
rect 637 855 641 859
rect 647 855 651 859
rect 655 855 659 859
rect 806 860 810 864
rect 814 860 818 864
rect 1209 864 1213 868
rect 1217 864 1221 868
rect 1604 868 1608 872
rect 1612 868 1616 872
rect 1628 864 1632 868
rect 1643 864 1647 868
rect 1685 868 1689 872
rect 1693 868 1697 872
rect 1709 864 1713 868
rect 1724 864 1728 868
rect 1658 860 1662 864
rect 1666 860 1670 864
rect 1092 855 1096 859
rect 1100 855 1104 859
rect 1430 855 1434 859
rect 1438 855 1442 859
rect 1446 855 1450 859
rect 1454 855 1458 859
rect 1462 855 1466 859
rect 1470 855 1474 859
rect 1481 855 1485 859
rect 1498 855 1502 859
rect 1515 855 1519 859
rect 1524 855 1528 859
rect 1537 855 1541 859
rect 1545 855 1549 859
rect 1553 855 1557 859
rect 1570 855 1574 859
rect 1580 855 1584 859
rect 1588 855 1592 859
rect 1739 860 1743 864
rect 1747 860 1751 864
rect 497 809 501 813
rect 505 809 509 813
rect 513 809 517 813
rect 521 809 525 813
rect 529 809 533 813
rect 537 809 541 813
rect 548 809 552 813
rect 565 809 569 813
rect 582 809 586 813
rect 591 809 595 813
rect 604 809 608 813
rect 612 809 616 813
rect 620 809 624 813
rect 637 809 641 813
rect 647 809 651 813
rect 655 809 659 813
rect 143 799 147 803
rect 151 799 155 803
rect 159 799 163 803
rect 172 799 176 803
rect 180 799 184 803
rect 188 799 192 803
rect 196 799 200 803
rect 204 799 208 803
rect 217 799 221 803
rect 230 799 234 803
rect 238 799 242 803
rect 246 799 250 803
rect 254 799 258 803
rect 267 799 271 803
rect 695 808 699 812
rect 710 808 714 812
rect 776 808 780 812
rect 791 808 795 812
rect 1430 809 1434 813
rect 1438 809 1442 813
rect 1446 809 1450 813
rect 1454 809 1458 813
rect 1462 809 1466 813
rect 1470 809 1474 813
rect 1481 809 1485 813
rect 1498 809 1502 813
rect 1515 809 1519 813
rect 1524 809 1528 813
rect 1537 809 1541 813
rect 1545 809 1549 813
rect 1553 809 1557 813
rect 1570 809 1574 813
rect 1580 809 1584 813
rect 1588 809 1592 813
rect 1076 799 1080 803
rect 1084 799 1088 803
rect 1092 799 1096 803
rect 1105 799 1109 803
rect 1113 799 1117 803
rect 1121 799 1125 803
rect 1129 799 1133 803
rect 1137 799 1141 803
rect 1150 799 1154 803
rect 1163 799 1167 803
rect 1171 799 1175 803
rect 1179 799 1183 803
rect 1187 799 1191 803
rect 1200 799 1204 803
rect 1628 808 1632 812
rect 1643 808 1647 812
rect 1709 808 1713 812
rect 1724 808 1728 812
rect 695 732 699 736
rect 710 732 714 736
rect 776 736 780 740
rect 784 736 788 740
rect 800 732 804 736
rect 815 732 819 736
rect 725 728 729 732
rect 733 728 737 732
rect 497 723 501 727
rect 505 723 509 727
rect 513 723 517 727
rect 521 723 525 727
rect 529 723 533 727
rect 537 723 541 727
rect 548 723 552 727
rect 565 723 569 727
rect 582 723 586 727
rect 591 723 595 727
rect 604 723 608 727
rect 612 723 616 727
rect 620 723 624 727
rect 637 723 641 727
rect 647 723 651 727
rect 655 723 659 727
rect 830 728 834 732
rect 838 728 842 732
rect 1628 732 1632 736
rect 1643 732 1647 736
rect 1709 736 1713 740
rect 1717 736 1721 740
rect 1733 732 1737 736
rect 1748 732 1752 736
rect 1658 728 1662 732
rect 1666 728 1670 732
rect 1430 723 1434 727
rect 1438 723 1442 727
rect 1446 723 1450 727
rect 1454 723 1458 727
rect 1462 723 1466 727
rect 1470 723 1474 727
rect 1481 723 1485 727
rect 1498 723 1502 727
rect 1515 723 1519 727
rect 1524 723 1528 727
rect 1537 723 1541 727
rect 1545 723 1549 727
rect 1553 723 1557 727
rect 1570 723 1574 727
rect 1580 723 1584 727
rect 1588 723 1592 727
rect 1763 728 1767 732
rect 1771 728 1775 732
rect 497 677 501 681
rect 505 677 509 681
rect 513 677 517 681
rect 521 677 525 681
rect 529 677 533 681
rect 537 677 541 681
rect 548 677 552 681
rect 565 677 569 681
rect 582 677 586 681
rect 591 677 595 681
rect 604 677 608 681
rect 612 677 616 681
rect 620 677 624 681
rect 637 677 641 681
rect 647 677 651 681
rect 655 677 659 681
rect 695 677 699 681
rect 710 677 714 681
rect 800 677 804 681
rect 815 677 819 681
rect 1430 677 1434 681
rect 1438 677 1442 681
rect 1446 677 1450 681
rect 1454 677 1458 681
rect 1462 677 1466 681
rect 1470 677 1474 681
rect 1481 677 1485 681
rect 1498 677 1502 681
rect 1515 677 1519 681
rect 1524 677 1528 681
rect 1537 677 1541 681
rect 1545 677 1549 681
rect 1553 677 1557 681
rect 1570 677 1574 681
rect 1580 677 1584 681
rect 1588 677 1592 681
rect 1628 677 1632 681
rect 1643 677 1647 681
rect 1733 677 1737 681
rect 1748 677 1752 681
rect 695 600 699 604
rect 710 600 714 604
rect 752 604 756 608
rect 760 604 764 608
rect 776 600 780 604
rect 791 600 795 604
rect 842 604 846 608
rect 850 604 854 608
rect 866 600 870 604
rect 881 600 885 604
rect 725 596 729 600
rect 733 596 737 600
rect 497 591 501 595
rect 505 591 509 595
rect 513 591 517 595
rect 521 591 525 595
rect 529 591 533 595
rect 537 591 541 595
rect 548 591 552 595
rect 565 591 569 595
rect 582 591 586 595
rect 591 591 595 595
rect 604 591 608 595
rect 612 591 616 595
rect 620 591 624 595
rect 637 591 641 595
rect 647 591 651 595
rect 655 591 659 595
rect 806 596 810 600
rect 814 596 818 600
rect 896 596 900 600
rect 904 596 908 600
rect 1628 600 1632 604
rect 1643 600 1647 604
rect 1685 604 1689 608
rect 1693 604 1697 608
rect 1709 600 1713 604
rect 1724 600 1728 604
rect 1775 604 1779 608
rect 1783 604 1787 608
rect 1799 600 1803 604
rect 1814 600 1818 604
rect 1658 596 1662 600
rect 1666 596 1670 600
rect 1430 591 1434 595
rect 1438 591 1442 595
rect 1446 591 1450 595
rect 1454 591 1458 595
rect 1462 591 1466 595
rect 1470 591 1474 595
rect 1481 591 1485 595
rect 1498 591 1502 595
rect 1515 591 1519 595
rect 1524 591 1528 595
rect 1537 591 1541 595
rect 1545 591 1549 595
rect 1553 591 1557 595
rect 1570 591 1574 595
rect 1580 591 1584 595
rect 1588 591 1592 595
rect 1739 596 1743 600
rect 1747 596 1751 600
rect 1829 596 1833 600
rect 1837 596 1841 600
rect 497 545 501 549
rect 505 545 509 549
rect 513 545 517 549
rect 521 545 525 549
rect 529 545 533 549
rect 537 545 541 549
rect 548 545 552 549
rect 565 545 569 549
rect 582 545 586 549
rect 591 545 595 549
rect 604 545 608 549
rect 612 545 616 549
rect 620 545 624 549
rect 637 545 641 549
rect 647 545 651 549
rect 655 545 659 549
rect 695 542 699 546
rect 710 542 714 546
rect 776 542 780 546
rect 791 542 795 546
rect 866 542 870 546
rect 881 542 885 546
rect 1430 545 1434 549
rect 1438 545 1442 549
rect 1446 545 1450 549
rect 1454 545 1458 549
rect 1462 545 1466 549
rect 1470 545 1474 549
rect 1481 545 1485 549
rect 1498 545 1502 549
rect 1515 545 1519 549
rect 1524 545 1528 549
rect 1537 545 1541 549
rect 1545 545 1549 549
rect 1553 545 1557 549
rect 1570 545 1574 549
rect 1580 545 1584 549
rect 1588 545 1592 549
rect 1628 542 1632 546
rect 1643 542 1647 546
rect 1709 542 1713 546
rect 1724 542 1728 546
rect 1799 542 1803 546
rect 1814 542 1818 546
rect 695 468 699 472
rect 710 468 714 472
rect 725 464 729 468
rect 733 464 737 468
rect 497 459 501 463
rect 505 459 509 463
rect 513 459 517 463
rect 521 459 525 463
rect 529 459 533 463
rect 537 459 541 463
rect 548 459 552 463
rect 565 459 569 463
rect 582 459 586 463
rect 591 459 595 463
rect 604 459 608 463
rect 612 459 616 463
rect 620 459 624 463
rect 637 459 641 463
rect 647 459 651 463
rect 655 459 659 463
rect 1628 468 1632 472
rect 1643 468 1647 472
rect 1658 464 1662 468
rect 1666 464 1670 468
rect 1430 459 1434 463
rect 1438 459 1442 463
rect 1446 459 1450 463
rect 1454 459 1458 463
rect 1462 459 1466 463
rect 1470 459 1474 463
rect 1481 459 1485 463
rect 1498 459 1502 463
rect 1515 459 1519 463
rect 1524 459 1528 463
rect 1537 459 1541 463
rect 1545 459 1549 463
rect 1553 459 1557 463
rect 1570 459 1574 463
rect 1580 459 1584 463
rect 1588 459 1592 463
rect 497 413 501 417
rect 505 413 509 417
rect 513 413 517 417
rect 521 413 525 417
rect 529 413 533 417
rect 537 413 541 417
rect 548 413 552 417
rect 565 413 569 417
rect 582 413 586 417
rect 591 413 595 417
rect 604 413 608 417
rect 612 413 616 417
rect 620 413 624 417
rect 637 413 641 417
rect 647 413 651 417
rect 655 413 659 417
rect 731 413 735 417
rect 739 413 743 417
rect 749 413 753 417
rect 757 413 761 417
rect 766 413 770 417
rect 774 413 778 417
rect 782 413 786 417
rect 790 413 794 417
rect 798 413 802 417
rect 809 413 813 417
rect 826 413 830 417
rect 843 413 847 417
rect 852 413 856 417
rect 865 413 869 417
rect 873 413 877 417
rect 881 413 885 417
rect 898 413 902 417
rect 908 413 912 417
rect 916 413 920 417
rect 20 399 24 403
rect 33 399 37 403
rect 41 399 45 403
rect 49 399 53 403
rect 57 399 61 403
rect 70 399 74 403
rect 83 399 87 403
rect 91 399 95 403
rect 99 399 103 403
rect 107 399 111 403
rect 115 399 119 403
rect 128 399 132 403
rect 136 399 140 403
rect 144 399 148 403
rect 152 399 156 403
rect 165 399 169 403
rect 173 399 177 403
rect 181 399 185 403
rect 189 399 193 403
rect 202 399 206 403
rect 215 399 219 403
rect 223 399 227 403
rect 231 399 235 403
rect 239 399 243 403
rect 247 399 251 403
rect 260 399 264 403
rect 268 399 272 403
rect 276 399 280 403
rect 284 399 288 403
rect 297 399 301 403
rect 305 399 309 403
rect 313 399 317 403
rect 321 399 325 403
rect 334 399 338 403
rect 347 399 351 403
rect 355 399 359 403
rect 363 399 367 403
rect 371 399 375 403
rect 379 399 383 403
rect 392 399 396 403
rect 400 399 404 403
rect 408 399 412 403
rect 695 406 699 410
rect 710 406 714 410
rect 1430 413 1434 417
rect 1438 413 1442 417
rect 1446 413 1450 417
rect 1454 413 1458 417
rect 1462 413 1466 417
rect 1470 413 1474 417
rect 1481 413 1485 417
rect 1498 413 1502 417
rect 1515 413 1519 417
rect 1524 413 1528 417
rect 1537 413 1541 417
rect 1545 413 1549 417
rect 1553 413 1557 417
rect 1570 413 1574 417
rect 1580 413 1584 417
rect 1588 413 1592 417
rect 1664 413 1668 417
rect 1672 413 1676 417
rect 1682 413 1686 417
rect 1690 413 1694 417
rect 1699 413 1703 417
rect 1707 413 1711 417
rect 1715 413 1719 417
rect 1723 413 1727 417
rect 1731 413 1735 417
rect 1742 413 1746 417
rect 1759 413 1763 417
rect 1776 413 1780 417
rect 1785 413 1789 417
rect 1798 413 1802 417
rect 1806 413 1810 417
rect 1814 413 1818 417
rect 1831 413 1835 417
rect 1841 413 1845 417
rect 1849 413 1853 417
rect 953 399 957 403
rect 966 399 970 403
rect 974 399 978 403
rect 982 399 986 403
rect 990 399 994 403
rect 1003 399 1007 403
rect 1016 399 1020 403
rect 1024 399 1028 403
rect 1032 399 1036 403
rect 1040 399 1044 403
rect 1048 399 1052 403
rect 1061 399 1065 403
rect 1069 399 1073 403
rect 1077 399 1081 403
rect 1085 399 1089 403
rect 1098 399 1102 403
rect 1106 399 1110 403
rect 1114 399 1118 403
rect 1122 399 1126 403
rect 1135 399 1139 403
rect 1148 399 1152 403
rect 1156 399 1160 403
rect 1164 399 1168 403
rect 1172 399 1176 403
rect 1180 399 1184 403
rect 1193 399 1197 403
rect 1201 399 1205 403
rect 1209 399 1213 403
rect 1217 399 1221 403
rect 1230 399 1234 403
rect 1238 399 1242 403
rect 1246 399 1250 403
rect 1254 399 1258 403
rect 1267 399 1271 403
rect 1280 399 1284 403
rect 1288 399 1292 403
rect 1296 399 1300 403
rect 1304 399 1308 403
rect 1312 399 1316 403
rect 1325 399 1329 403
rect 1333 399 1337 403
rect 1341 399 1345 403
rect 1628 406 1632 410
rect 1643 406 1647 410
rect 925 360 929 364
rect 135 355 139 359
rect 143 355 147 359
rect 159 355 163 359
rect 167 355 171 359
rect 1858 360 1862 364
rect 925 352 929 356
rect 1068 355 1072 359
rect 1076 355 1080 359
rect 1092 355 1096 359
rect 1100 355 1104 359
rect 1858 352 1862 356
rect 155 344 159 348
rect 163 344 167 348
rect 1088 344 1092 348
rect 1096 344 1100 348
rect 151 333 155 337
rect 1084 333 1088 337
rect 151 325 155 329
rect 135 321 139 325
rect 143 321 147 325
rect 159 321 163 325
rect 167 321 171 325
rect 1084 325 1088 329
rect 1068 321 1072 325
rect 1076 321 1080 325
rect 1092 321 1096 325
rect 1100 321 1104 325
rect 791 289 795 293
rect 804 289 808 293
rect 812 289 816 293
rect 820 289 824 293
rect 828 289 832 293
rect 841 289 845 293
rect 854 289 858 293
rect 862 289 866 293
rect 870 289 874 293
rect 878 289 882 293
rect 886 289 890 293
rect 899 289 903 293
rect 907 289 911 293
rect 915 289 919 293
rect 1724 289 1728 293
rect 1737 289 1741 293
rect 1745 289 1749 293
rect 1753 289 1757 293
rect 1761 289 1765 293
rect 1774 289 1778 293
rect 1787 289 1791 293
rect 1795 289 1799 293
rect 1803 289 1807 293
rect 1811 289 1815 293
rect 1819 289 1823 293
rect 1832 289 1836 293
rect 1840 289 1844 293
rect 1848 289 1852 293
rect 20 259 24 263
rect 33 259 37 263
rect 41 259 45 263
rect 49 259 53 263
rect 57 259 61 263
rect 70 259 74 263
rect 83 259 87 263
rect 91 259 95 263
rect 99 259 103 263
rect 107 259 111 263
rect 115 259 119 263
rect 128 259 132 263
rect 136 259 140 263
rect 144 259 148 263
rect 152 259 156 263
rect 165 259 169 263
rect 173 259 177 263
rect 181 259 185 263
rect 189 259 193 263
rect 202 259 206 263
rect 215 259 219 263
rect 223 259 227 263
rect 231 259 235 263
rect 239 259 243 263
rect 247 259 251 263
rect 260 259 264 263
rect 268 259 272 263
rect 276 259 280 263
rect 284 259 288 263
rect 297 259 301 263
rect 305 259 309 263
rect 313 259 317 263
rect 321 259 325 263
rect 334 259 338 263
rect 347 259 351 263
rect 355 259 359 263
rect 363 259 367 263
rect 371 259 375 263
rect 379 259 383 263
rect 392 259 396 263
rect 400 259 404 263
rect 408 259 412 263
rect 953 259 957 263
rect 966 259 970 263
rect 974 259 978 263
rect 982 259 986 263
rect 990 259 994 263
rect 1003 259 1007 263
rect 1016 259 1020 263
rect 1024 259 1028 263
rect 1032 259 1036 263
rect 1040 259 1044 263
rect 1048 259 1052 263
rect 1061 259 1065 263
rect 1069 259 1073 263
rect 1077 259 1081 263
rect 1085 259 1089 263
rect 1098 259 1102 263
rect 1106 259 1110 263
rect 1114 259 1118 263
rect 1122 259 1126 263
rect 1135 259 1139 263
rect 1148 259 1152 263
rect 1156 259 1160 263
rect 1164 259 1168 263
rect 1172 259 1176 263
rect 1180 259 1184 263
rect 1193 259 1197 263
rect 1201 259 1205 263
rect 1209 259 1213 263
rect 1217 259 1221 263
rect 1230 259 1234 263
rect 1238 259 1242 263
rect 1246 259 1250 263
rect 1254 259 1258 263
rect 1267 259 1271 263
rect 1280 259 1284 263
rect 1288 259 1292 263
rect 1296 259 1300 263
rect 1304 259 1308 263
rect 1312 259 1316 263
rect 1325 259 1329 263
rect 1333 259 1337 263
rect 1341 259 1345 263
rect 937 216 941 220
rect 937 208 941 212
rect 1870 216 1874 220
rect 1870 208 1874 212
rect 791 203 795 207
rect 804 203 808 207
rect 812 203 816 207
rect 820 203 824 207
rect 828 203 832 207
rect 841 203 845 207
rect 854 203 858 207
rect 862 203 866 207
rect 870 203 874 207
rect 878 203 882 207
rect 886 203 890 207
rect 899 203 903 207
rect 907 203 911 207
rect 915 203 919 207
rect 1724 203 1728 207
rect 1737 203 1741 207
rect 1745 203 1749 207
rect 1753 203 1757 207
rect 1761 203 1765 207
rect 1774 203 1778 207
rect 1787 203 1791 207
rect 1795 203 1799 207
rect 1803 203 1807 207
rect 1811 203 1815 207
rect 1819 203 1823 207
rect 1832 203 1836 207
rect 1840 203 1844 207
rect 1848 203 1852 207
rect 20 173 24 177
rect 33 173 37 177
rect 41 173 45 177
rect 49 173 53 177
rect 57 173 61 177
rect 70 173 74 177
rect 83 173 87 177
rect 91 173 95 177
rect 99 173 103 177
rect 107 173 111 177
rect 115 173 119 177
rect 128 173 132 177
rect 136 173 140 177
rect 144 173 148 177
rect 152 173 156 177
rect 165 173 169 177
rect 173 173 177 177
rect 181 173 185 177
rect 189 173 193 177
rect 202 173 206 177
rect 215 173 219 177
rect 223 173 227 177
rect 231 173 235 177
rect 239 173 243 177
rect 247 173 251 177
rect 260 173 264 177
rect 268 173 272 177
rect 276 173 280 177
rect 284 173 288 177
rect 297 173 301 177
rect 305 173 309 177
rect 313 173 317 177
rect 321 173 325 177
rect 334 173 338 177
rect 347 173 351 177
rect 355 173 359 177
rect 363 173 367 177
rect 371 173 375 177
rect 379 173 383 177
rect 392 173 396 177
rect 400 173 404 177
rect 408 173 412 177
rect 953 173 957 177
rect 966 173 970 177
rect 974 173 978 177
rect 982 173 986 177
rect 990 173 994 177
rect 1003 173 1007 177
rect 1016 173 1020 177
rect 1024 173 1028 177
rect 1032 173 1036 177
rect 1040 173 1044 177
rect 1048 173 1052 177
rect 1061 173 1065 177
rect 1069 173 1073 177
rect 1077 173 1081 177
rect 1085 173 1089 177
rect 1098 173 1102 177
rect 1106 173 1110 177
rect 1114 173 1118 177
rect 1122 173 1126 177
rect 1135 173 1139 177
rect 1148 173 1152 177
rect 1156 173 1160 177
rect 1164 173 1168 177
rect 1172 173 1176 177
rect 1180 173 1184 177
rect 1193 173 1197 177
rect 1201 173 1205 177
rect 1209 173 1213 177
rect 1217 173 1221 177
rect 1230 173 1234 177
rect 1238 173 1242 177
rect 1246 173 1250 177
rect 1254 173 1258 177
rect 1267 173 1271 177
rect 1280 173 1284 177
rect 1288 173 1292 177
rect 1296 173 1300 177
rect 1304 173 1308 177
rect 1312 173 1316 177
rect 1325 173 1329 177
rect 1333 173 1337 177
rect 1341 173 1345 177
rect 252 129 256 133
rect 260 129 264 133
rect 276 129 280 133
rect 284 129 288 133
rect 1185 129 1189 133
rect 1193 129 1197 133
rect 1209 129 1213 133
rect 1217 129 1221 133
rect 272 118 276 122
rect 280 118 284 122
rect 1205 118 1209 122
rect 1213 118 1217 122
rect 268 107 272 111
rect 1201 107 1205 111
rect 268 99 272 103
rect 1201 99 1205 103
rect 252 95 256 99
rect 260 95 264 99
rect 276 95 280 99
rect 284 95 288 99
rect 1185 95 1189 99
rect 1193 95 1197 99
rect 1209 95 1213 99
rect 1217 95 1221 99
rect 20 33 24 37
rect 33 33 37 37
rect 41 33 45 37
rect 49 33 53 37
rect 57 33 61 37
rect 70 33 74 37
rect 83 33 87 37
rect 91 33 95 37
rect 99 33 103 37
rect 107 33 111 37
rect 115 33 119 37
rect 128 33 132 37
rect 136 33 140 37
rect 144 33 148 37
rect 152 33 156 37
rect 165 33 169 37
rect 173 33 177 37
rect 181 33 185 37
rect 189 33 193 37
rect 202 33 206 37
rect 215 33 219 37
rect 223 33 227 37
rect 231 33 235 37
rect 239 33 243 37
rect 247 33 251 37
rect 260 33 264 37
rect 268 33 272 37
rect 276 33 280 37
rect 284 33 288 37
rect 297 33 301 37
rect 305 33 309 37
rect 313 33 317 37
rect 321 33 325 37
rect 334 33 338 37
rect 347 33 351 37
rect 355 33 359 37
rect 363 33 367 37
rect 371 33 375 37
rect 379 33 383 37
rect 392 33 396 37
rect 400 33 404 37
rect 408 33 412 37
rect 953 33 957 37
rect 966 33 970 37
rect 974 33 978 37
rect 982 33 986 37
rect 990 33 994 37
rect 1003 33 1007 37
rect 1016 33 1020 37
rect 1024 33 1028 37
rect 1032 33 1036 37
rect 1040 33 1044 37
rect 1048 33 1052 37
rect 1061 33 1065 37
rect 1069 33 1073 37
rect 1077 33 1081 37
rect 1085 33 1089 37
rect 1098 33 1102 37
rect 1106 33 1110 37
rect 1114 33 1118 37
rect 1122 33 1126 37
rect 1135 33 1139 37
rect 1148 33 1152 37
rect 1156 33 1160 37
rect 1164 33 1168 37
rect 1172 33 1176 37
rect 1180 33 1184 37
rect 1193 33 1197 37
rect 1201 33 1205 37
rect 1209 33 1213 37
rect 1217 33 1221 37
rect 1230 33 1234 37
rect 1238 33 1242 37
rect 1246 33 1250 37
rect 1254 33 1258 37
rect 1267 33 1271 37
rect 1280 33 1284 37
rect 1288 33 1292 37
rect 1296 33 1300 37
rect 1304 33 1308 37
rect 1312 33 1316 37
rect 1325 33 1329 37
rect 1333 33 1337 37
rect 1341 33 1345 37
<< pdcontact >>
rect 492 1937 496 1945
rect 505 1937 509 1945
rect 513 1937 517 1945
rect 521 1941 525 1945
rect 529 1937 533 1945
rect 542 1937 546 1945
rect 555 1937 559 1945
rect 563 1937 567 1945
rect 571 1937 575 1945
rect 579 1941 583 1945
rect 587 1937 591 1945
rect 600 1937 604 1945
rect 608 1937 612 1945
rect 616 1937 620 1945
rect 624 1937 628 1945
rect 637 1937 641 1945
rect 645 1937 649 1945
rect 653 1941 657 1945
rect 661 1937 665 1945
rect 674 1937 678 1945
rect 687 1937 691 1945
rect 695 1937 699 1945
rect 703 1937 707 1945
rect 711 1941 715 1945
rect 719 1937 723 1945
rect 732 1937 736 1945
rect 740 1937 744 1945
rect 748 1937 752 1945
rect 756 1937 760 1945
rect 769 1937 773 1945
rect 777 1937 781 1945
rect 785 1941 789 1945
rect 793 1937 797 1945
rect 806 1937 810 1945
rect 819 1937 823 1945
rect 827 1937 831 1945
rect 835 1937 839 1945
rect 843 1941 847 1945
rect 851 1937 855 1945
rect 864 1937 868 1945
rect 872 1937 876 1945
rect 880 1937 884 1945
rect 888 1937 892 1945
rect 901 1937 905 1945
rect 909 1937 913 1945
rect 917 1941 921 1945
rect 925 1937 929 1945
rect 938 1937 942 1945
rect 951 1937 955 1945
rect 959 1937 963 1945
rect 967 1937 971 1945
rect 975 1941 979 1945
rect 983 1937 987 1945
rect 996 1937 1000 1945
rect 1004 1937 1008 1945
rect 1012 1937 1016 1945
rect 1425 1937 1429 1945
rect 1438 1937 1442 1945
rect 1446 1937 1450 1945
rect 1454 1941 1458 1945
rect 1462 1937 1466 1945
rect 1475 1937 1479 1945
rect 1488 1937 1492 1945
rect 1496 1937 1500 1945
rect 1504 1937 1508 1945
rect 1512 1941 1516 1945
rect 1520 1937 1524 1945
rect 1533 1937 1537 1945
rect 1541 1937 1545 1945
rect 1549 1937 1553 1945
rect 1557 1937 1561 1945
rect 1570 1937 1574 1945
rect 1578 1937 1582 1945
rect 1586 1941 1590 1945
rect 1594 1937 1598 1945
rect 1607 1937 1611 1945
rect 1620 1937 1624 1945
rect 1628 1937 1632 1945
rect 1636 1937 1640 1945
rect 1644 1941 1648 1945
rect 1652 1937 1656 1945
rect 1665 1937 1669 1945
rect 1673 1937 1677 1945
rect 1681 1937 1685 1945
rect 1689 1937 1693 1945
rect 1702 1937 1706 1945
rect 1710 1937 1714 1945
rect 1718 1941 1722 1945
rect 1726 1937 1730 1945
rect 1739 1937 1743 1945
rect 1752 1937 1756 1945
rect 1760 1937 1764 1945
rect 1768 1937 1772 1945
rect 1776 1941 1780 1945
rect 1784 1937 1788 1945
rect 1797 1937 1801 1945
rect 1805 1937 1809 1945
rect 1813 1937 1817 1945
rect 1821 1937 1825 1945
rect 1834 1937 1838 1945
rect 1842 1937 1846 1945
rect 1850 1941 1854 1945
rect 1858 1937 1862 1945
rect 1871 1937 1875 1945
rect 1884 1937 1888 1945
rect 1892 1937 1896 1945
rect 1900 1937 1904 1945
rect 1908 1941 1912 1945
rect 1916 1937 1920 1945
rect 1929 1937 1933 1945
rect 1937 1937 1941 1945
rect 1945 1937 1949 1945
rect 152 1904 156 1912
rect 165 1904 169 1912
rect 173 1904 177 1912
rect 181 1908 185 1912
rect 189 1904 193 1912
rect 202 1904 206 1912
rect 215 1904 219 1912
rect 223 1904 227 1912
rect 231 1904 235 1912
rect 239 1908 243 1912
rect 247 1904 251 1912
rect 260 1904 264 1912
rect 268 1904 272 1912
rect 276 1904 280 1912
rect 1085 1904 1089 1912
rect 1098 1904 1102 1912
rect 1106 1904 1110 1912
rect 1114 1908 1118 1912
rect 1122 1904 1126 1912
rect 1135 1904 1139 1912
rect 1148 1904 1152 1912
rect 1156 1904 1160 1912
rect 1164 1904 1168 1912
rect 1172 1908 1176 1912
rect 1180 1904 1184 1912
rect 1193 1904 1197 1912
rect 1201 1904 1205 1912
rect 1209 1904 1213 1912
rect 671 1866 675 1874
rect 679 1866 683 1874
rect 497 1853 501 1861
rect 505 1853 509 1861
rect 513 1853 517 1861
rect 521 1853 525 1861
rect 529 1853 533 1861
rect 537 1853 541 1861
rect 548 1853 552 1861
rect 565 1853 569 1861
rect 582 1853 586 1861
rect 591 1853 595 1861
rect 604 1853 608 1861
rect 612 1853 616 1861
rect 620 1853 624 1861
rect 637 1853 641 1861
rect 647 1853 651 1861
rect 655 1853 659 1861
rect 695 1860 699 1868
rect 710 1860 714 1868
rect 725 1866 729 1874
rect 733 1866 737 1874
rect 752 1866 756 1874
rect 760 1866 764 1874
rect 776 1860 780 1868
rect 791 1860 795 1868
rect 806 1866 810 1874
rect 814 1866 818 1874
rect 1604 1866 1608 1874
rect 1612 1866 1616 1874
rect 1430 1853 1434 1861
rect 1438 1853 1442 1861
rect 1446 1853 1450 1861
rect 1454 1853 1458 1861
rect 1462 1853 1466 1861
rect 1470 1853 1474 1861
rect 1481 1853 1485 1861
rect 1498 1853 1502 1861
rect 1515 1853 1519 1861
rect 1524 1853 1528 1861
rect 1537 1853 1541 1861
rect 1545 1853 1549 1861
rect 1553 1853 1557 1861
rect 1570 1853 1574 1861
rect 1580 1853 1584 1861
rect 1588 1853 1592 1861
rect 1628 1860 1632 1868
rect 1643 1860 1647 1868
rect 1658 1866 1662 1874
rect 1666 1866 1670 1874
rect 1685 1866 1689 1874
rect 1693 1866 1697 1874
rect 1709 1860 1713 1868
rect 1724 1860 1728 1868
rect 1739 1866 1743 1874
rect 1747 1866 1751 1874
rect 143 1802 147 1810
rect 151 1802 155 1810
rect 159 1802 163 1810
rect 172 1802 176 1810
rect 180 1806 184 1810
rect 188 1802 192 1810
rect 196 1802 200 1810
rect 204 1802 208 1810
rect 217 1802 221 1810
rect 230 1802 234 1810
rect 238 1806 242 1810
rect 246 1802 250 1810
rect 254 1802 258 1810
rect 267 1802 271 1810
rect 1076 1802 1080 1810
rect 1084 1802 1088 1810
rect 1092 1802 1096 1810
rect 1105 1802 1109 1810
rect 1113 1806 1117 1810
rect 1121 1802 1125 1810
rect 1129 1802 1133 1810
rect 1137 1802 1141 1810
rect 1150 1802 1154 1810
rect 1163 1802 1167 1810
rect 1171 1806 1175 1810
rect 1179 1802 1183 1810
rect 1187 1802 1191 1810
rect 1200 1802 1204 1810
rect 497 1767 501 1775
rect 505 1767 509 1775
rect 513 1767 517 1775
rect 521 1767 525 1775
rect 529 1767 533 1775
rect 537 1767 541 1775
rect 548 1767 552 1775
rect 565 1767 569 1775
rect 582 1767 586 1775
rect 591 1767 595 1775
rect 604 1767 608 1775
rect 612 1767 616 1775
rect 620 1767 624 1775
rect 637 1767 641 1775
rect 647 1767 651 1775
rect 655 1767 659 1775
rect 695 1768 699 1776
rect 710 1768 714 1776
rect 776 1768 780 1776
rect 791 1768 795 1776
rect 1430 1767 1434 1775
rect 1438 1767 1442 1775
rect 1446 1767 1450 1775
rect 1454 1767 1458 1775
rect 1462 1767 1466 1775
rect 1470 1767 1474 1775
rect 1481 1767 1485 1775
rect 1498 1767 1502 1775
rect 1515 1767 1519 1775
rect 1524 1767 1528 1775
rect 1537 1767 1541 1775
rect 1545 1767 1549 1775
rect 1553 1767 1557 1775
rect 1570 1767 1574 1775
rect 1580 1767 1584 1775
rect 1588 1767 1592 1775
rect 1628 1768 1632 1776
rect 1643 1768 1647 1776
rect 1709 1768 1713 1776
rect 1724 1768 1728 1776
rect 497 1721 501 1729
rect 505 1721 509 1729
rect 513 1721 517 1729
rect 521 1721 525 1729
rect 529 1721 533 1729
rect 537 1721 541 1729
rect 548 1721 552 1729
rect 565 1721 569 1729
rect 582 1721 586 1729
rect 591 1721 595 1729
rect 604 1721 608 1729
rect 612 1721 616 1729
rect 620 1721 624 1729
rect 637 1721 641 1729
rect 647 1721 651 1729
rect 655 1721 659 1729
rect 695 1728 699 1736
rect 710 1728 714 1736
rect 725 1734 729 1742
rect 733 1734 737 1742
rect 776 1734 780 1742
rect 784 1734 788 1742
rect 800 1728 804 1736
rect 815 1728 819 1736
rect 830 1734 834 1742
rect 838 1734 842 1742
rect 1430 1721 1434 1729
rect 1438 1721 1442 1729
rect 1446 1721 1450 1729
rect 1454 1721 1458 1729
rect 1462 1721 1466 1729
rect 1470 1721 1474 1729
rect 1481 1721 1485 1729
rect 1498 1721 1502 1729
rect 1515 1721 1519 1729
rect 1524 1721 1528 1729
rect 1537 1721 1541 1729
rect 1545 1721 1549 1729
rect 1553 1721 1557 1729
rect 1570 1721 1574 1729
rect 1580 1721 1584 1729
rect 1588 1721 1592 1729
rect 1628 1728 1632 1736
rect 1643 1728 1647 1736
rect 1658 1734 1662 1742
rect 1666 1734 1670 1742
rect 1709 1734 1713 1742
rect 1717 1734 1721 1742
rect 1733 1728 1737 1736
rect 1748 1728 1752 1736
rect 1763 1734 1767 1742
rect 1771 1734 1775 1742
rect 497 1635 501 1643
rect 505 1635 509 1643
rect 513 1635 517 1643
rect 521 1635 525 1643
rect 529 1635 533 1643
rect 537 1635 541 1643
rect 548 1635 552 1643
rect 565 1635 569 1643
rect 582 1635 586 1643
rect 591 1635 595 1643
rect 604 1635 608 1643
rect 612 1635 616 1643
rect 620 1635 624 1643
rect 637 1635 641 1643
rect 647 1635 651 1643
rect 655 1635 659 1643
rect 695 1637 699 1645
rect 710 1637 714 1645
rect 800 1637 804 1645
rect 815 1637 819 1645
rect 1430 1635 1434 1643
rect 1438 1635 1442 1643
rect 1446 1635 1450 1643
rect 1454 1635 1458 1643
rect 1462 1635 1466 1643
rect 1470 1635 1474 1643
rect 1481 1635 1485 1643
rect 1498 1635 1502 1643
rect 1515 1635 1519 1643
rect 1524 1635 1528 1643
rect 1537 1635 1541 1643
rect 1545 1635 1549 1643
rect 1553 1635 1557 1643
rect 1570 1635 1574 1643
rect 1580 1635 1584 1643
rect 1588 1635 1592 1643
rect 1628 1637 1632 1645
rect 1643 1637 1647 1645
rect 1733 1637 1737 1645
rect 1748 1637 1752 1645
rect 497 1589 501 1597
rect 505 1589 509 1597
rect 513 1589 517 1597
rect 521 1589 525 1597
rect 529 1589 533 1597
rect 537 1589 541 1597
rect 548 1589 552 1597
rect 565 1589 569 1597
rect 582 1589 586 1597
rect 591 1589 595 1597
rect 604 1589 608 1597
rect 612 1589 616 1597
rect 620 1589 624 1597
rect 637 1589 641 1597
rect 647 1589 651 1597
rect 655 1589 659 1597
rect 695 1596 699 1604
rect 710 1596 714 1604
rect 725 1602 729 1610
rect 733 1602 737 1610
rect 752 1602 756 1610
rect 760 1602 764 1610
rect 776 1596 780 1604
rect 791 1596 795 1604
rect 806 1602 810 1610
rect 814 1602 818 1610
rect 842 1602 846 1610
rect 850 1602 854 1610
rect 866 1596 870 1604
rect 881 1596 885 1604
rect 896 1602 900 1610
rect 904 1602 908 1610
rect 1430 1589 1434 1597
rect 1438 1589 1442 1597
rect 1446 1589 1450 1597
rect 1454 1589 1458 1597
rect 1462 1589 1466 1597
rect 1470 1589 1474 1597
rect 1481 1589 1485 1597
rect 1498 1589 1502 1597
rect 1515 1589 1519 1597
rect 1524 1589 1528 1597
rect 1537 1589 1541 1597
rect 1545 1589 1549 1597
rect 1553 1589 1557 1597
rect 1570 1589 1574 1597
rect 1580 1589 1584 1597
rect 1588 1589 1592 1597
rect 1628 1596 1632 1604
rect 1643 1596 1647 1604
rect 1658 1602 1662 1610
rect 1666 1602 1670 1610
rect 1685 1602 1689 1610
rect 1693 1602 1697 1610
rect 1709 1596 1713 1604
rect 1724 1596 1728 1604
rect 1739 1602 1743 1610
rect 1747 1602 1751 1610
rect 1775 1602 1779 1610
rect 1783 1602 1787 1610
rect 1799 1596 1803 1604
rect 1814 1596 1818 1604
rect 1829 1602 1833 1610
rect 1837 1602 1841 1610
rect 497 1503 501 1511
rect 505 1503 509 1511
rect 513 1503 517 1511
rect 521 1503 525 1511
rect 529 1503 533 1511
rect 537 1503 541 1511
rect 548 1503 552 1511
rect 565 1503 569 1511
rect 582 1503 586 1511
rect 591 1503 595 1511
rect 604 1503 608 1511
rect 612 1503 616 1511
rect 620 1503 624 1511
rect 637 1503 641 1511
rect 647 1503 651 1511
rect 655 1503 659 1511
rect 695 1502 699 1510
rect 710 1502 714 1510
rect 776 1502 780 1510
rect 791 1502 795 1510
rect 866 1502 870 1510
rect 881 1502 885 1510
rect 1430 1503 1434 1511
rect 1438 1503 1442 1511
rect 1446 1503 1450 1511
rect 1454 1503 1458 1511
rect 1462 1503 1466 1511
rect 1470 1503 1474 1511
rect 1481 1503 1485 1511
rect 1498 1503 1502 1511
rect 1515 1503 1519 1511
rect 1524 1503 1528 1511
rect 1537 1503 1541 1511
rect 1545 1503 1549 1511
rect 1553 1503 1557 1511
rect 1570 1503 1574 1511
rect 1580 1503 1584 1511
rect 1588 1503 1592 1511
rect 1628 1502 1632 1510
rect 1643 1502 1647 1510
rect 1709 1502 1713 1510
rect 1724 1502 1728 1510
rect 1799 1502 1803 1510
rect 1814 1502 1818 1510
rect 497 1457 501 1465
rect 505 1457 509 1465
rect 513 1457 517 1465
rect 521 1457 525 1465
rect 529 1457 533 1465
rect 537 1457 541 1465
rect 548 1457 552 1465
rect 565 1457 569 1465
rect 582 1457 586 1465
rect 591 1457 595 1465
rect 604 1457 608 1465
rect 612 1457 616 1465
rect 620 1457 624 1465
rect 637 1457 641 1465
rect 647 1457 651 1465
rect 655 1457 659 1465
rect 695 1464 699 1472
rect 710 1464 714 1472
rect 725 1470 729 1478
rect 733 1470 737 1478
rect 1430 1457 1434 1465
rect 1438 1457 1442 1465
rect 1446 1457 1450 1465
rect 1454 1457 1458 1465
rect 1462 1457 1466 1465
rect 1470 1457 1474 1465
rect 1481 1457 1485 1465
rect 1498 1457 1502 1465
rect 1515 1457 1519 1465
rect 1524 1457 1528 1465
rect 1537 1457 1541 1465
rect 1545 1457 1549 1465
rect 1553 1457 1557 1465
rect 1570 1457 1574 1465
rect 1580 1457 1584 1465
rect 1588 1457 1592 1465
rect 1628 1464 1632 1472
rect 1643 1464 1647 1472
rect 1658 1470 1662 1478
rect 1666 1470 1670 1478
rect 20 1402 24 1410
rect 33 1402 37 1410
rect 41 1402 45 1410
rect 49 1406 53 1410
rect 57 1402 61 1410
rect 70 1402 74 1410
rect 83 1402 87 1410
rect 91 1402 95 1410
rect 99 1402 103 1410
rect 107 1406 111 1410
rect 115 1402 119 1410
rect 128 1402 132 1410
rect 136 1402 140 1410
rect 144 1402 148 1410
rect 152 1402 156 1410
rect 165 1402 169 1410
rect 173 1402 177 1410
rect 181 1406 185 1410
rect 189 1402 193 1410
rect 202 1402 206 1410
rect 215 1402 219 1410
rect 223 1402 227 1410
rect 231 1402 235 1410
rect 239 1406 243 1410
rect 247 1402 251 1410
rect 260 1402 264 1410
rect 268 1402 272 1410
rect 276 1402 280 1410
rect 284 1402 288 1410
rect 297 1402 301 1410
rect 305 1402 309 1410
rect 313 1406 317 1410
rect 321 1402 325 1410
rect 334 1402 338 1410
rect 347 1402 351 1410
rect 355 1402 359 1410
rect 363 1402 367 1410
rect 371 1406 375 1410
rect 379 1402 383 1410
rect 392 1402 396 1410
rect 400 1402 404 1410
rect 408 1402 412 1410
rect 953 1402 957 1410
rect 966 1402 970 1410
rect 974 1402 978 1410
rect 982 1406 986 1410
rect 990 1402 994 1410
rect 1003 1402 1007 1410
rect 1016 1402 1020 1410
rect 1024 1402 1028 1410
rect 1032 1402 1036 1410
rect 1040 1406 1044 1410
rect 1048 1402 1052 1410
rect 1061 1402 1065 1410
rect 1069 1402 1073 1410
rect 1077 1402 1081 1410
rect 1085 1402 1089 1410
rect 1098 1402 1102 1410
rect 1106 1402 1110 1410
rect 1114 1406 1118 1410
rect 1122 1402 1126 1410
rect 1135 1402 1139 1410
rect 1148 1402 1152 1410
rect 1156 1402 1160 1410
rect 1164 1402 1168 1410
rect 1172 1406 1176 1410
rect 1180 1402 1184 1410
rect 1193 1402 1197 1410
rect 1201 1402 1205 1410
rect 1209 1402 1213 1410
rect 1217 1402 1221 1410
rect 1230 1402 1234 1410
rect 1238 1402 1242 1410
rect 1246 1406 1250 1410
rect 1254 1402 1258 1410
rect 1267 1402 1271 1410
rect 1280 1402 1284 1410
rect 1288 1402 1292 1410
rect 1296 1402 1300 1410
rect 1304 1406 1308 1410
rect 1312 1402 1316 1410
rect 1325 1402 1329 1410
rect 1333 1402 1337 1410
rect 1341 1402 1345 1410
rect 497 1371 501 1379
rect 505 1371 509 1379
rect 513 1371 517 1379
rect 521 1371 525 1379
rect 529 1371 533 1379
rect 537 1371 541 1379
rect 548 1371 552 1379
rect 565 1371 569 1379
rect 582 1371 586 1379
rect 591 1371 595 1379
rect 604 1371 608 1379
rect 612 1371 616 1379
rect 620 1371 624 1379
rect 637 1371 641 1379
rect 647 1371 651 1379
rect 655 1371 659 1379
rect 695 1366 699 1374
rect 710 1366 714 1374
rect 731 1371 735 1379
rect 739 1371 743 1379
rect 749 1371 753 1379
rect 757 1371 761 1379
rect 766 1371 770 1379
rect 774 1371 778 1379
rect 782 1371 786 1379
rect 790 1371 794 1379
rect 798 1371 802 1379
rect 809 1371 813 1379
rect 826 1371 830 1379
rect 843 1371 847 1379
rect 852 1371 856 1379
rect 865 1371 869 1379
rect 873 1371 877 1379
rect 881 1371 885 1379
rect 898 1371 902 1379
rect 908 1371 912 1379
rect 916 1371 920 1379
rect 1430 1371 1434 1379
rect 1438 1371 1442 1379
rect 1446 1371 1450 1379
rect 1454 1371 1458 1379
rect 1462 1371 1466 1379
rect 1470 1371 1474 1379
rect 1481 1371 1485 1379
rect 1498 1371 1502 1379
rect 1515 1371 1519 1379
rect 1524 1371 1528 1379
rect 1537 1371 1541 1379
rect 1545 1371 1549 1379
rect 1553 1371 1557 1379
rect 1570 1371 1574 1379
rect 1580 1371 1584 1379
rect 1588 1371 1592 1379
rect 1628 1366 1632 1374
rect 1643 1366 1647 1374
rect 1664 1371 1668 1379
rect 1672 1371 1676 1379
rect 1682 1371 1686 1379
rect 1690 1371 1694 1379
rect 1699 1371 1703 1379
rect 1707 1371 1711 1379
rect 1715 1371 1719 1379
rect 1723 1371 1727 1379
rect 1731 1371 1735 1379
rect 1742 1371 1746 1379
rect 1759 1371 1763 1379
rect 1776 1371 1780 1379
rect 1785 1371 1789 1379
rect 1798 1371 1802 1379
rect 1806 1371 1810 1379
rect 1814 1371 1818 1379
rect 1831 1371 1835 1379
rect 1841 1371 1845 1379
rect 1849 1371 1853 1379
rect 791 1292 795 1300
rect 804 1292 808 1300
rect 812 1292 816 1300
rect 820 1296 824 1300
rect 828 1292 832 1300
rect 841 1292 845 1300
rect 854 1292 858 1300
rect 862 1292 866 1300
rect 870 1292 874 1300
rect 878 1296 882 1300
rect 886 1292 890 1300
rect 899 1292 903 1300
rect 907 1292 911 1300
rect 915 1292 919 1300
rect 1724 1292 1728 1300
rect 1737 1292 1741 1300
rect 1745 1292 1749 1300
rect 1753 1296 1757 1300
rect 1761 1292 1765 1300
rect 1774 1292 1778 1300
rect 1787 1292 1791 1300
rect 1795 1292 1799 1300
rect 1803 1292 1807 1300
rect 1811 1296 1815 1300
rect 1819 1292 1823 1300
rect 1832 1292 1836 1300
rect 1840 1292 1844 1300
rect 1848 1292 1852 1300
rect 20 1262 24 1270
rect 33 1262 37 1270
rect 41 1262 45 1270
rect 49 1266 53 1270
rect 57 1262 61 1270
rect 70 1262 74 1270
rect 83 1262 87 1270
rect 91 1262 95 1270
rect 99 1262 103 1270
rect 107 1266 111 1270
rect 115 1262 119 1270
rect 128 1262 132 1270
rect 136 1262 140 1270
rect 144 1262 148 1270
rect 152 1262 156 1270
rect 165 1262 169 1270
rect 173 1262 177 1270
rect 181 1266 185 1270
rect 189 1262 193 1270
rect 202 1262 206 1270
rect 215 1262 219 1270
rect 223 1262 227 1270
rect 231 1262 235 1270
rect 239 1266 243 1270
rect 247 1262 251 1270
rect 260 1262 264 1270
rect 268 1262 272 1270
rect 276 1262 280 1270
rect 284 1262 288 1270
rect 297 1262 301 1270
rect 305 1262 309 1270
rect 313 1266 317 1270
rect 321 1262 325 1270
rect 334 1262 338 1270
rect 347 1262 351 1270
rect 355 1262 359 1270
rect 363 1262 367 1270
rect 371 1266 375 1270
rect 379 1262 383 1270
rect 392 1262 396 1270
rect 400 1262 404 1270
rect 408 1262 412 1270
rect 953 1262 957 1270
rect 966 1262 970 1270
rect 974 1262 978 1270
rect 982 1266 986 1270
rect 990 1262 994 1270
rect 1003 1262 1007 1270
rect 1016 1262 1020 1270
rect 1024 1262 1028 1270
rect 1032 1262 1036 1270
rect 1040 1266 1044 1270
rect 1048 1262 1052 1270
rect 1061 1262 1065 1270
rect 1069 1262 1073 1270
rect 1077 1262 1081 1270
rect 1085 1262 1089 1270
rect 1098 1262 1102 1270
rect 1106 1262 1110 1270
rect 1114 1266 1118 1270
rect 1122 1262 1126 1270
rect 1135 1262 1139 1270
rect 1148 1262 1152 1270
rect 1156 1262 1160 1270
rect 1164 1262 1168 1270
rect 1172 1266 1176 1270
rect 1180 1262 1184 1270
rect 1193 1262 1197 1270
rect 1201 1262 1205 1270
rect 1209 1262 1213 1270
rect 1217 1262 1221 1270
rect 1230 1262 1234 1270
rect 1238 1262 1242 1270
rect 1246 1266 1250 1270
rect 1254 1262 1258 1270
rect 1267 1262 1271 1270
rect 1280 1262 1284 1270
rect 1288 1262 1292 1270
rect 1296 1262 1300 1270
rect 1304 1266 1308 1270
rect 1312 1262 1316 1270
rect 1325 1262 1329 1270
rect 1333 1262 1337 1270
rect 1341 1262 1345 1270
rect 791 1206 795 1214
rect 804 1206 808 1214
rect 812 1206 816 1214
rect 820 1210 824 1214
rect 828 1206 832 1214
rect 841 1206 845 1214
rect 854 1206 858 1214
rect 862 1206 866 1214
rect 870 1206 874 1214
rect 878 1210 882 1214
rect 886 1206 890 1214
rect 899 1206 903 1214
rect 907 1206 911 1214
rect 915 1206 919 1214
rect 1724 1206 1728 1214
rect 1737 1206 1741 1214
rect 1745 1206 1749 1214
rect 1753 1210 1757 1214
rect 1761 1206 1765 1214
rect 1774 1206 1778 1214
rect 1787 1206 1791 1214
rect 1795 1206 1799 1214
rect 1803 1206 1807 1214
rect 1811 1210 1815 1214
rect 1819 1206 1823 1214
rect 1832 1206 1836 1214
rect 1840 1206 1844 1214
rect 1848 1206 1852 1214
rect 20 1176 24 1184
rect 33 1176 37 1184
rect 41 1176 45 1184
rect 49 1180 53 1184
rect 57 1176 61 1184
rect 70 1176 74 1184
rect 83 1176 87 1184
rect 91 1176 95 1184
rect 99 1176 103 1184
rect 107 1180 111 1184
rect 115 1176 119 1184
rect 128 1176 132 1184
rect 136 1176 140 1184
rect 144 1176 148 1184
rect 152 1176 156 1184
rect 165 1176 169 1184
rect 173 1176 177 1184
rect 181 1180 185 1184
rect 189 1176 193 1184
rect 202 1176 206 1184
rect 215 1176 219 1184
rect 223 1176 227 1184
rect 231 1176 235 1184
rect 239 1180 243 1184
rect 247 1176 251 1184
rect 260 1176 264 1184
rect 268 1176 272 1184
rect 276 1176 280 1184
rect 284 1176 288 1184
rect 297 1176 301 1184
rect 305 1176 309 1184
rect 313 1180 317 1184
rect 321 1176 325 1184
rect 334 1176 338 1184
rect 347 1176 351 1184
rect 355 1176 359 1184
rect 363 1176 367 1184
rect 371 1180 375 1184
rect 379 1176 383 1184
rect 392 1176 396 1184
rect 400 1176 404 1184
rect 408 1176 412 1184
rect 953 1176 957 1184
rect 966 1176 970 1184
rect 974 1176 978 1184
rect 982 1180 986 1184
rect 990 1176 994 1184
rect 1003 1176 1007 1184
rect 1016 1176 1020 1184
rect 1024 1176 1028 1184
rect 1032 1176 1036 1184
rect 1040 1180 1044 1184
rect 1048 1176 1052 1184
rect 1061 1176 1065 1184
rect 1069 1176 1073 1184
rect 1077 1176 1081 1184
rect 1085 1176 1089 1184
rect 1098 1176 1102 1184
rect 1106 1176 1110 1184
rect 1114 1180 1118 1184
rect 1122 1176 1126 1184
rect 1135 1176 1139 1184
rect 1148 1176 1152 1184
rect 1156 1176 1160 1184
rect 1164 1176 1168 1184
rect 1172 1180 1176 1184
rect 1180 1176 1184 1184
rect 1193 1176 1197 1184
rect 1201 1176 1205 1184
rect 1209 1176 1213 1184
rect 1217 1176 1221 1184
rect 1230 1176 1234 1184
rect 1238 1176 1242 1184
rect 1246 1180 1250 1184
rect 1254 1176 1258 1184
rect 1267 1176 1271 1184
rect 1280 1176 1284 1184
rect 1288 1176 1292 1184
rect 1296 1176 1300 1184
rect 1304 1180 1308 1184
rect 1312 1176 1316 1184
rect 1325 1176 1329 1184
rect 1333 1176 1337 1184
rect 1341 1176 1345 1184
rect 20 1036 24 1044
rect 33 1036 37 1044
rect 41 1036 45 1044
rect 49 1040 53 1044
rect 57 1036 61 1044
rect 70 1036 74 1044
rect 83 1036 87 1044
rect 91 1036 95 1044
rect 99 1036 103 1044
rect 107 1040 111 1044
rect 115 1036 119 1044
rect 128 1036 132 1044
rect 136 1036 140 1044
rect 144 1036 148 1044
rect 152 1036 156 1044
rect 165 1036 169 1044
rect 173 1036 177 1044
rect 181 1040 185 1044
rect 189 1036 193 1044
rect 202 1036 206 1044
rect 215 1036 219 1044
rect 223 1036 227 1044
rect 231 1036 235 1044
rect 239 1040 243 1044
rect 247 1036 251 1044
rect 260 1036 264 1044
rect 268 1036 272 1044
rect 276 1036 280 1044
rect 284 1036 288 1044
rect 297 1036 301 1044
rect 305 1036 309 1044
rect 313 1040 317 1044
rect 321 1036 325 1044
rect 334 1036 338 1044
rect 347 1036 351 1044
rect 355 1036 359 1044
rect 363 1036 367 1044
rect 371 1040 375 1044
rect 379 1036 383 1044
rect 392 1036 396 1044
rect 400 1036 404 1044
rect 408 1036 412 1044
rect 953 1036 957 1044
rect 966 1036 970 1044
rect 974 1036 978 1044
rect 982 1040 986 1044
rect 990 1036 994 1044
rect 1003 1036 1007 1044
rect 1016 1036 1020 1044
rect 1024 1036 1028 1044
rect 1032 1036 1036 1044
rect 1040 1040 1044 1044
rect 1048 1036 1052 1044
rect 1061 1036 1065 1044
rect 1069 1036 1073 1044
rect 1077 1036 1081 1044
rect 1085 1036 1089 1044
rect 1098 1036 1102 1044
rect 1106 1036 1110 1044
rect 1114 1040 1118 1044
rect 1122 1036 1126 1044
rect 1135 1036 1139 1044
rect 1148 1036 1152 1044
rect 1156 1036 1160 1044
rect 1164 1036 1168 1044
rect 1172 1040 1176 1044
rect 1180 1036 1184 1044
rect 1193 1036 1197 1044
rect 1201 1036 1205 1044
rect 1209 1036 1213 1044
rect 1217 1036 1221 1044
rect 1230 1036 1234 1044
rect 1238 1036 1242 1044
rect 1246 1040 1250 1044
rect 1254 1036 1258 1044
rect 1267 1036 1271 1044
rect 1280 1036 1284 1044
rect 1288 1036 1292 1044
rect 1296 1036 1300 1044
rect 1304 1040 1308 1044
rect 1312 1036 1316 1044
rect 1325 1036 1329 1044
rect 1333 1036 1337 1044
rect 1341 1036 1345 1044
rect 492 957 496 965
rect 505 957 509 965
rect 513 957 517 965
rect 521 961 525 965
rect 529 957 533 965
rect 542 957 546 965
rect 555 957 559 965
rect 563 957 567 965
rect 571 957 575 965
rect 579 961 583 965
rect 587 957 591 965
rect 600 957 604 965
rect 608 957 612 965
rect 616 957 620 965
rect 624 957 628 965
rect 637 957 641 965
rect 645 957 649 965
rect 653 961 657 965
rect 661 957 665 965
rect 674 957 678 965
rect 687 957 691 965
rect 695 957 699 965
rect 703 957 707 965
rect 711 961 715 965
rect 719 957 723 965
rect 732 957 736 965
rect 740 957 744 965
rect 748 957 752 965
rect 756 957 760 965
rect 769 957 773 965
rect 777 957 781 965
rect 785 961 789 965
rect 793 957 797 965
rect 806 957 810 965
rect 819 957 823 965
rect 827 957 831 965
rect 835 957 839 965
rect 843 961 847 965
rect 851 957 855 965
rect 864 957 868 965
rect 872 957 876 965
rect 880 957 884 965
rect 888 957 892 965
rect 901 957 905 965
rect 909 957 913 965
rect 917 961 921 965
rect 925 957 929 965
rect 938 957 942 965
rect 951 957 955 965
rect 959 957 963 965
rect 967 957 971 965
rect 975 961 979 965
rect 983 957 987 965
rect 996 957 1000 965
rect 1004 957 1008 965
rect 1012 957 1016 965
rect 1425 957 1429 965
rect 1438 957 1442 965
rect 1446 957 1450 965
rect 1454 961 1458 965
rect 1462 957 1466 965
rect 1475 957 1479 965
rect 1488 957 1492 965
rect 1496 957 1500 965
rect 1504 957 1508 965
rect 1512 961 1516 965
rect 1520 957 1524 965
rect 1533 957 1537 965
rect 1541 957 1545 965
rect 1549 957 1553 965
rect 1557 957 1561 965
rect 1570 957 1574 965
rect 1578 957 1582 965
rect 1586 961 1590 965
rect 1594 957 1598 965
rect 1607 957 1611 965
rect 1620 957 1624 965
rect 1628 957 1632 965
rect 1636 957 1640 965
rect 1644 961 1648 965
rect 1652 957 1656 965
rect 1665 957 1669 965
rect 1673 957 1677 965
rect 1681 957 1685 965
rect 1689 957 1693 965
rect 1702 957 1706 965
rect 1710 957 1714 965
rect 1718 961 1722 965
rect 1726 957 1730 965
rect 1739 957 1743 965
rect 1752 957 1756 965
rect 1760 957 1764 965
rect 1768 957 1772 965
rect 1776 961 1780 965
rect 1784 957 1788 965
rect 1797 957 1801 965
rect 1805 957 1809 965
rect 1813 957 1817 965
rect 1821 957 1825 965
rect 1834 957 1838 965
rect 1842 957 1846 965
rect 1850 961 1854 965
rect 1858 957 1862 965
rect 1871 957 1875 965
rect 1884 957 1888 965
rect 1892 957 1896 965
rect 1900 957 1904 965
rect 1908 961 1912 965
rect 1916 957 1920 965
rect 1929 957 1933 965
rect 1937 957 1941 965
rect 1945 957 1949 965
rect 152 924 156 932
rect 165 924 169 932
rect 173 924 177 932
rect 181 928 185 932
rect 189 924 193 932
rect 202 924 206 932
rect 215 924 219 932
rect 223 924 227 932
rect 231 924 235 932
rect 239 928 243 932
rect 247 924 251 932
rect 260 924 264 932
rect 268 924 272 932
rect 276 924 280 932
rect 1085 924 1089 932
rect 1098 924 1102 932
rect 1106 924 1110 932
rect 1114 928 1118 932
rect 1122 924 1126 932
rect 1135 924 1139 932
rect 1148 924 1152 932
rect 1156 924 1160 932
rect 1164 924 1168 932
rect 1172 928 1176 932
rect 1180 924 1184 932
rect 1193 924 1197 932
rect 1201 924 1205 932
rect 1209 924 1213 932
rect 671 886 675 894
rect 679 886 683 894
rect 497 873 501 881
rect 505 873 509 881
rect 513 873 517 881
rect 521 873 525 881
rect 529 873 533 881
rect 537 873 541 881
rect 548 873 552 881
rect 565 873 569 881
rect 582 873 586 881
rect 591 873 595 881
rect 604 873 608 881
rect 612 873 616 881
rect 620 873 624 881
rect 637 873 641 881
rect 647 873 651 881
rect 655 873 659 881
rect 695 880 699 888
rect 710 880 714 888
rect 725 886 729 894
rect 733 886 737 894
rect 752 886 756 894
rect 760 886 764 894
rect 776 880 780 888
rect 791 880 795 888
rect 806 886 810 894
rect 814 886 818 894
rect 1604 886 1608 894
rect 1612 886 1616 894
rect 1430 873 1434 881
rect 1438 873 1442 881
rect 1446 873 1450 881
rect 1454 873 1458 881
rect 1462 873 1466 881
rect 1470 873 1474 881
rect 1481 873 1485 881
rect 1498 873 1502 881
rect 1515 873 1519 881
rect 1524 873 1528 881
rect 1537 873 1541 881
rect 1545 873 1549 881
rect 1553 873 1557 881
rect 1570 873 1574 881
rect 1580 873 1584 881
rect 1588 873 1592 881
rect 1628 880 1632 888
rect 1643 880 1647 888
rect 1658 886 1662 894
rect 1666 886 1670 894
rect 1685 886 1689 894
rect 1693 886 1697 894
rect 1709 880 1713 888
rect 1724 880 1728 888
rect 1739 886 1743 894
rect 1747 886 1751 894
rect 143 822 147 830
rect 151 822 155 830
rect 159 822 163 830
rect 172 822 176 830
rect 180 826 184 830
rect 188 822 192 830
rect 196 822 200 830
rect 204 822 208 830
rect 217 822 221 830
rect 230 822 234 830
rect 238 826 242 830
rect 246 822 250 830
rect 254 822 258 830
rect 267 822 271 830
rect 1076 822 1080 830
rect 1084 822 1088 830
rect 1092 822 1096 830
rect 1105 822 1109 830
rect 1113 826 1117 830
rect 1121 822 1125 830
rect 1129 822 1133 830
rect 1137 822 1141 830
rect 1150 822 1154 830
rect 1163 822 1167 830
rect 1171 826 1175 830
rect 1179 822 1183 830
rect 1187 822 1191 830
rect 1200 822 1204 830
rect 497 787 501 795
rect 505 787 509 795
rect 513 787 517 795
rect 521 787 525 795
rect 529 787 533 795
rect 537 787 541 795
rect 548 787 552 795
rect 565 787 569 795
rect 582 787 586 795
rect 591 787 595 795
rect 604 787 608 795
rect 612 787 616 795
rect 620 787 624 795
rect 637 787 641 795
rect 647 787 651 795
rect 655 787 659 795
rect 695 788 699 796
rect 710 788 714 796
rect 776 788 780 796
rect 791 788 795 796
rect 1430 787 1434 795
rect 1438 787 1442 795
rect 1446 787 1450 795
rect 1454 787 1458 795
rect 1462 787 1466 795
rect 1470 787 1474 795
rect 1481 787 1485 795
rect 1498 787 1502 795
rect 1515 787 1519 795
rect 1524 787 1528 795
rect 1537 787 1541 795
rect 1545 787 1549 795
rect 1553 787 1557 795
rect 1570 787 1574 795
rect 1580 787 1584 795
rect 1588 787 1592 795
rect 1628 788 1632 796
rect 1643 788 1647 796
rect 1709 788 1713 796
rect 1724 788 1728 796
rect 497 741 501 749
rect 505 741 509 749
rect 513 741 517 749
rect 521 741 525 749
rect 529 741 533 749
rect 537 741 541 749
rect 548 741 552 749
rect 565 741 569 749
rect 582 741 586 749
rect 591 741 595 749
rect 604 741 608 749
rect 612 741 616 749
rect 620 741 624 749
rect 637 741 641 749
rect 647 741 651 749
rect 655 741 659 749
rect 695 748 699 756
rect 710 748 714 756
rect 725 754 729 762
rect 733 754 737 762
rect 776 754 780 762
rect 784 754 788 762
rect 800 748 804 756
rect 815 748 819 756
rect 830 754 834 762
rect 838 754 842 762
rect 1430 741 1434 749
rect 1438 741 1442 749
rect 1446 741 1450 749
rect 1454 741 1458 749
rect 1462 741 1466 749
rect 1470 741 1474 749
rect 1481 741 1485 749
rect 1498 741 1502 749
rect 1515 741 1519 749
rect 1524 741 1528 749
rect 1537 741 1541 749
rect 1545 741 1549 749
rect 1553 741 1557 749
rect 1570 741 1574 749
rect 1580 741 1584 749
rect 1588 741 1592 749
rect 1628 748 1632 756
rect 1643 748 1647 756
rect 1658 754 1662 762
rect 1666 754 1670 762
rect 1709 754 1713 762
rect 1717 754 1721 762
rect 1733 748 1737 756
rect 1748 748 1752 756
rect 1763 754 1767 762
rect 1771 754 1775 762
rect 497 655 501 663
rect 505 655 509 663
rect 513 655 517 663
rect 521 655 525 663
rect 529 655 533 663
rect 537 655 541 663
rect 548 655 552 663
rect 565 655 569 663
rect 582 655 586 663
rect 591 655 595 663
rect 604 655 608 663
rect 612 655 616 663
rect 620 655 624 663
rect 637 655 641 663
rect 647 655 651 663
rect 655 655 659 663
rect 695 657 699 665
rect 710 657 714 665
rect 800 657 804 665
rect 815 657 819 665
rect 1430 655 1434 663
rect 1438 655 1442 663
rect 1446 655 1450 663
rect 1454 655 1458 663
rect 1462 655 1466 663
rect 1470 655 1474 663
rect 1481 655 1485 663
rect 1498 655 1502 663
rect 1515 655 1519 663
rect 1524 655 1528 663
rect 1537 655 1541 663
rect 1545 655 1549 663
rect 1553 655 1557 663
rect 1570 655 1574 663
rect 1580 655 1584 663
rect 1588 655 1592 663
rect 1628 657 1632 665
rect 1643 657 1647 665
rect 1733 657 1737 665
rect 1748 657 1752 665
rect 497 609 501 617
rect 505 609 509 617
rect 513 609 517 617
rect 521 609 525 617
rect 529 609 533 617
rect 537 609 541 617
rect 548 609 552 617
rect 565 609 569 617
rect 582 609 586 617
rect 591 609 595 617
rect 604 609 608 617
rect 612 609 616 617
rect 620 609 624 617
rect 637 609 641 617
rect 647 609 651 617
rect 655 609 659 617
rect 695 616 699 624
rect 710 616 714 624
rect 725 622 729 630
rect 733 622 737 630
rect 752 622 756 630
rect 760 622 764 630
rect 776 616 780 624
rect 791 616 795 624
rect 806 622 810 630
rect 814 622 818 630
rect 842 622 846 630
rect 850 622 854 630
rect 866 616 870 624
rect 881 616 885 624
rect 896 622 900 630
rect 904 622 908 630
rect 1430 609 1434 617
rect 1438 609 1442 617
rect 1446 609 1450 617
rect 1454 609 1458 617
rect 1462 609 1466 617
rect 1470 609 1474 617
rect 1481 609 1485 617
rect 1498 609 1502 617
rect 1515 609 1519 617
rect 1524 609 1528 617
rect 1537 609 1541 617
rect 1545 609 1549 617
rect 1553 609 1557 617
rect 1570 609 1574 617
rect 1580 609 1584 617
rect 1588 609 1592 617
rect 1628 616 1632 624
rect 1643 616 1647 624
rect 1658 622 1662 630
rect 1666 622 1670 630
rect 1685 622 1689 630
rect 1693 622 1697 630
rect 1709 616 1713 624
rect 1724 616 1728 624
rect 1739 622 1743 630
rect 1747 622 1751 630
rect 1775 622 1779 630
rect 1783 622 1787 630
rect 1799 616 1803 624
rect 1814 616 1818 624
rect 1829 622 1833 630
rect 1837 622 1841 630
rect 497 523 501 531
rect 505 523 509 531
rect 513 523 517 531
rect 521 523 525 531
rect 529 523 533 531
rect 537 523 541 531
rect 548 523 552 531
rect 565 523 569 531
rect 582 523 586 531
rect 591 523 595 531
rect 604 523 608 531
rect 612 523 616 531
rect 620 523 624 531
rect 637 523 641 531
rect 647 523 651 531
rect 655 523 659 531
rect 695 522 699 530
rect 710 522 714 530
rect 776 522 780 530
rect 791 522 795 530
rect 866 522 870 530
rect 881 522 885 530
rect 1430 523 1434 531
rect 1438 523 1442 531
rect 1446 523 1450 531
rect 1454 523 1458 531
rect 1462 523 1466 531
rect 1470 523 1474 531
rect 1481 523 1485 531
rect 1498 523 1502 531
rect 1515 523 1519 531
rect 1524 523 1528 531
rect 1537 523 1541 531
rect 1545 523 1549 531
rect 1553 523 1557 531
rect 1570 523 1574 531
rect 1580 523 1584 531
rect 1588 523 1592 531
rect 1628 522 1632 530
rect 1643 522 1647 530
rect 1709 522 1713 530
rect 1724 522 1728 530
rect 1799 522 1803 530
rect 1814 522 1818 530
rect 497 477 501 485
rect 505 477 509 485
rect 513 477 517 485
rect 521 477 525 485
rect 529 477 533 485
rect 537 477 541 485
rect 548 477 552 485
rect 565 477 569 485
rect 582 477 586 485
rect 591 477 595 485
rect 604 477 608 485
rect 612 477 616 485
rect 620 477 624 485
rect 637 477 641 485
rect 647 477 651 485
rect 655 477 659 485
rect 695 484 699 492
rect 710 484 714 492
rect 725 490 729 498
rect 733 490 737 498
rect 1430 477 1434 485
rect 1438 477 1442 485
rect 1446 477 1450 485
rect 1454 477 1458 485
rect 1462 477 1466 485
rect 1470 477 1474 485
rect 1481 477 1485 485
rect 1498 477 1502 485
rect 1515 477 1519 485
rect 1524 477 1528 485
rect 1537 477 1541 485
rect 1545 477 1549 485
rect 1553 477 1557 485
rect 1570 477 1574 485
rect 1580 477 1584 485
rect 1588 477 1592 485
rect 1628 484 1632 492
rect 1643 484 1647 492
rect 1658 490 1662 498
rect 1666 490 1670 498
rect 20 422 24 430
rect 33 422 37 430
rect 41 422 45 430
rect 49 426 53 430
rect 57 422 61 430
rect 70 422 74 430
rect 83 422 87 430
rect 91 422 95 430
rect 99 422 103 430
rect 107 426 111 430
rect 115 422 119 430
rect 128 422 132 430
rect 136 422 140 430
rect 144 422 148 430
rect 152 422 156 430
rect 165 422 169 430
rect 173 422 177 430
rect 181 426 185 430
rect 189 422 193 430
rect 202 422 206 430
rect 215 422 219 430
rect 223 422 227 430
rect 231 422 235 430
rect 239 426 243 430
rect 247 422 251 430
rect 260 422 264 430
rect 268 422 272 430
rect 276 422 280 430
rect 284 422 288 430
rect 297 422 301 430
rect 305 422 309 430
rect 313 426 317 430
rect 321 422 325 430
rect 334 422 338 430
rect 347 422 351 430
rect 355 422 359 430
rect 363 422 367 430
rect 371 426 375 430
rect 379 422 383 430
rect 392 422 396 430
rect 400 422 404 430
rect 408 422 412 430
rect 953 422 957 430
rect 966 422 970 430
rect 974 422 978 430
rect 982 426 986 430
rect 990 422 994 430
rect 1003 422 1007 430
rect 1016 422 1020 430
rect 1024 422 1028 430
rect 1032 422 1036 430
rect 1040 426 1044 430
rect 1048 422 1052 430
rect 1061 422 1065 430
rect 1069 422 1073 430
rect 1077 422 1081 430
rect 1085 422 1089 430
rect 1098 422 1102 430
rect 1106 422 1110 430
rect 1114 426 1118 430
rect 1122 422 1126 430
rect 1135 422 1139 430
rect 1148 422 1152 430
rect 1156 422 1160 430
rect 1164 422 1168 430
rect 1172 426 1176 430
rect 1180 422 1184 430
rect 1193 422 1197 430
rect 1201 422 1205 430
rect 1209 422 1213 430
rect 1217 422 1221 430
rect 1230 422 1234 430
rect 1238 422 1242 430
rect 1246 426 1250 430
rect 1254 422 1258 430
rect 1267 422 1271 430
rect 1280 422 1284 430
rect 1288 422 1292 430
rect 1296 422 1300 430
rect 1304 426 1308 430
rect 1312 422 1316 430
rect 1325 422 1329 430
rect 1333 422 1337 430
rect 1341 422 1345 430
rect 497 391 501 399
rect 505 391 509 399
rect 513 391 517 399
rect 521 391 525 399
rect 529 391 533 399
rect 537 391 541 399
rect 548 391 552 399
rect 565 391 569 399
rect 582 391 586 399
rect 591 391 595 399
rect 604 391 608 399
rect 612 391 616 399
rect 620 391 624 399
rect 637 391 641 399
rect 647 391 651 399
rect 655 391 659 399
rect 695 386 699 394
rect 710 386 714 394
rect 731 391 735 399
rect 739 391 743 399
rect 749 391 753 399
rect 757 391 761 399
rect 766 391 770 399
rect 774 391 778 399
rect 782 391 786 399
rect 790 391 794 399
rect 798 391 802 399
rect 809 391 813 399
rect 826 391 830 399
rect 843 391 847 399
rect 852 391 856 399
rect 865 391 869 399
rect 873 391 877 399
rect 881 391 885 399
rect 898 391 902 399
rect 908 391 912 399
rect 916 391 920 399
rect 1430 391 1434 399
rect 1438 391 1442 399
rect 1446 391 1450 399
rect 1454 391 1458 399
rect 1462 391 1466 399
rect 1470 391 1474 399
rect 1481 391 1485 399
rect 1498 391 1502 399
rect 1515 391 1519 399
rect 1524 391 1528 399
rect 1537 391 1541 399
rect 1545 391 1549 399
rect 1553 391 1557 399
rect 1570 391 1574 399
rect 1580 391 1584 399
rect 1588 391 1592 399
rect 1628 386 1632 394
rect 1643 386 1647 394
rect 1664 391 1668 399
rect 1672 391 1676 399
rect 1682 391 1686 399
rect 1690 391 1694 399
rect 1699 391 1703 399
rect 1707 391 1711 399
rect 1715 391 1719 399
rect 1723 391 1727 399
rect 1731 391 1735 399
rect 1742 391 1746 399
rect 1759 391 1763 399
rect 1776 391 1780 399
rect 1785 391 1789 399
rect 1798 391 1802 399
rect 1806 391 1810 399
rect 1814 391 1818 399
rect 1831 391 1835 399
rect 1841 391 1845 399
rect 1849 391 1853 399
rect 791 312 795 320
rect 804 312 808 320
rect 812 312 816 320
rect 820 316 824 320
rect 828 312 832 320
rect 841 312 845 320
rect 854 312 858 320
rect 862 312 866 320
rect 870 312 874 320
rect 878 316 882 320
rect 886 312 890 320
rect 899 312 903 320
rect 907 312 911 320
rect 915 312 919 320
rect 1724 312 1728 320
rect 1737 312 1741 320
rect 1745 312 1749 320
rect 1753 316 1757 320
rect 1761 312 1765 320
rect 1774 312 1778 320
rect 1787 312 1791 320
rect 1795 312 1799 320
rect 1803 312 1807 320
rect 1811 316 1815 320
rect 1819 312 1823 320
rect 1832 312 1836 320
rect 1840 312 1844 320
rect 1848 312 1852 320
rect 20 282 24 290
rect 33 282 37 290
rect 41 282 45 290
rect 49 286 53 290
rect 57 282 61 290
rect 70 282 74 290
rect 83 282 87 290
rect 91 282 95 290
rect 99 282 103 290
rect 107 286 111 290
rect 115 282 119 290
rect 128 282 132 290
rect 136 282 140 290
rect 144 282 148 290
rect 152 282 156 290
rect 165 282 169 290
rect 173 282 177 290
rect 181 286 185 290
rect 189 282 193 290
rect 202 282 206 290
rect 215 282 219 290
rect 223 282 227 290
rect 231 282 235 290
rect 239 286 243 290
rect 247 282 251 290
rect 260 282 264 290
rect 268 282 272 290
rect 276 282 280 290
rect 284 282 288 290
rect 297 282 301 290
rect 305 282 309 290
rect 313 286 317 290
rect 321 282 325 290
rect 334 282 338 290
rect 347 282 351 290
rect 355 282 359 290
rect 363 282 367 290
rect 371 286 375 290
rect 379 282 383 290
rect 392 282 396 290
rect 400 282 404 290
rect 408 282 412 290
rect 953 282 957 290
rect 966 282 970 290
rect 974 282 978 290
rect 982 286 986 290
rect 990 282 994 290
rect 1003 282 1007 290
rect 1016 282 1020 290
rect 1024 282 1028 290
rect 1032 282 1036 290
rect 1040 286 1044 290
rect 1048 282 1052 290
rect 1061 282 1065 290
rect 1069 282 1073 290
rect 1077 282 1081 290
rect 1085 282 1089 290
rect 1098 282 1102 290
rect 1106 282 1110 290
rect 1114 286 1118 290
rect 1122 282 1126 290
rect 1135 282 1139 290
rect 1148 282 1152 290
rect 1156 282 1160 290
rect 1164 282 1168 290
rect 1172 286 1176 290
rect 1180 282 1184 290
rect 1193 282 1197 290
rect 1201 282 1205 290
rect 1209 282 1213 290
rect 1217 282 1221 290
rect 1230 282 1234 290
rect 1238 282 1242 290
rect 1246 286 1250 290
rect 1254 282 1258 290
rect 1267 282 1271 290
rect 1280 282 1284 290
rect 1288 282 1292 290
rect 1296 282 1300 290
rect 1304 286 1308 290
rect 1312 282 1316 290
rect 1325 282 1329 290
rect 1333 282 1337 290
rect 1341 282 1345 290
rect 791 226 795 234
rect 804 226 808 234
rect 812 226 816 234
rect 820 230 824 234
rect 828 226 832 234
rect 841 226 845 234
rect 854 226 858 234
rect 862 226 866 234
rect 870 226 874 234
rect 878 230 882 234
rect 886 226 890 234
rect 899 226 903 234
rect 907 226 911 234
rect 915 226 919 234
rect 1724 226 1728 234
rect 1737 226 1741 234
rect 1745 226 1749 234
rect 1753 230 1757 234
rect 1761 226 1765 234
rect 1774 226 1778 234
rect 1787 226 1791 234
rect 1795 226 1799 234
rect 1803 226 1807 234
rect 1811 230 1815 234
rect 1819 226 1823 234
rect 1832 226 1836 234
rect 1840 226 1844 234
rect 1848 226 1852 234
rect 20 196 24 204
rect 33 196 37 204
rect 41 196 45 204
rect 49 200 53 204
rect 57 196 61 204
rect 70 196 74 204
rect 83 196 87 204
rect 91 196 95 204
rect 99 196 103 204
rect 107 200 111 204
rect 115 196 119 204
rect 128 196 132 204
rect 136 196 140 204
rect 144 196 148 204
rect 152 196 156 204
rect 165 196 169 204
rect 173 196 177 204
rect 181 200 185 204
rect 189 196 193 204
rect 202 196 206 204
rect 215 196 219 204
rect 223 196 227 204
rect 231 196 235 204
rect 239 200 243 204
rect 247 196 251 204
rect 260 196 264 204
rect 268 196 272 204
rect 276 196 280 204
rect 284 196 288 204
rect 297 196 301 204
rect 305 196 309 204
rect 313 200 317 204
rect 321 196 325 204
rect 334 196 338 204
rect 347 196 351 204
rect 355 196 359 204
rect 363 196 367 204
rect 371 200 375 204
rect 379 196 383 204
rect 392 196 396 204
rect 400 196 404 204
rect 408 196 412 204
rect 953 196 957 204
rect 966 196 970 204
rect 974 196 978 204
rect 982 200 986 204
rect 990 196 994 204
rect 1003 196 1007 204
rect 1016 196 1020 204
rect 1024 196 1028 204
rect 1032 196 1036 204
rect 1040 200 1044 204
rect 1048 196 1052 204
rect 1061 196 1065 204
rect 1069 196 1073 204
rect 1077 196 1081 204
rect 1085 196 1089 204
rect 1098 196 1102 204
rect 1106 196 1110 204
rect 1114 200 1118 204
rect 1122 196 1126 204
rect 1135 196 1139 204
rect 1148 196 1152 204
rect 1156 196 1160 204
rect 1164 196 1168 204
rect 1172 200 1176 204
rect 1180 196 1184 204
rect 1193 196 1197 204
rect 1201 196 1205 204
rect 1209 196 1213 204
rect 1217 196 1221 204
rect 1230 196 1234 204
rect 1238 196 1242 204
rect 1246 200 1250 204
rect 1254 196 1258 204
rect 1267 196 1271 204
rect 1280 196 1284 204
rect 1288 196 1292 204
rect 1296 196 1300 204
rect 1304 200 1308 204
rect 1312 196 1316 204
rect 1325 196 1329 204
rect 1333 196 1337 204
rect 1341 196 1345 204
rect 20 56 24 64
rect 33 56 37 64
rect 41 56 45 64
rect 49 60 53 64
rect 57 56 61 64
rect 70 56 74 64
rect 83 56 87 64
rect 91 56 95 64
rect 99 56 103 64
rect 107 60 111 64
rect 115 56 119 64
rect 128 56 132 64
rect 136 56 140 64
rect 144 56 148 64
rect 152 56 156 64
rect 165 56 169 64
rect 173 56 177 64
rect 181 60 185 64
rect 189 56 193 64
rect 202 56 206 64
rect 215 56 219 64
rect 223 56 227 64
rect 231 56 235 64
rect 239 60 243 64
rect 247 56 251 64
rect 260 56 264 64
rect 268 56 272 64
rect 276 56 280 64
rect 284 56 288 64
rect 297 56 301 64
rect 305 56 309 64
rect 313 60 317 64
rect 321 56 325 64
rect 334 56 338 64
rect 347 56 351 64
rect 355 56 359 64
rect 363 56 367 64
rect 371 60 375 64
rect 379 56 383 64
rect 392 56 396 64
rect 400 56 404 64
rect 408 56 412 64
rect 953 56 957 64
rect 966 56 970 64
rect 974 56 978 64
rect 982 60 986 64
rect 990 56 994 64
rect 1003 56 1007 64
rect 1016 56 1020 64
rect 1024 56 1028 64
rect 1032 56 1036 64
rect 1040 60 1044 64
rect 1048 56 1052 64
rect 1061 56 1065 64
rect 1069 56 1073 64
rect 1077 56 1081 64
rect 1085 56 1089 64
rect 1098 56 1102 64
rect 1106 56 1110 64
rect 1114 60 1118 64
rect 1122 56 1126 64
rect 1135 56 1139 64
rect 1148 56 1152 64
rect 1156 56 1160 64
rect 1164 56 1168 64
rect 1172 60 1176 64
rect 1180 56 1184 64
rect 1193 56 1197 64
rect 1201 56 1205 64
rect 1209 56 1213 64
rect 1217 56 1221 64
rect 1230 56 1234 64
rect 1238 56 1242 64
rect 1246 60 1250 64
rect 1254 56 1258 64
rect 1267 56 1271 64
rect 1280 56 1284 64
rect 1288 56 1292 64
rect 1296 56 1300 64
rect 1304 60 1308 64
rect 1312 56 1316 64
rect 1325 56 1329 64
rect 1333 56 1337 64
rect 1341 56 1345 64
<< psubstratepcontact >>
rect 522 1898 526 1902
rect 550 1898 554 1902
rect 580 1898 584 1902
rect 654 1898 658 1902
rect 682 1898 686 1902
rect 712 1898 716 1902
rect 786 1898 790 1902
rect 814 1898 818 1902
rect 844 1898 848 1902
rect 918 1898 922 1902
rect 946 1898 950 1902
rect 976 1898 980 1902
rect 1455 1898 1459 1902
rect 1483 1898 1487 1902
rect 1513 1898 1517 1902
rect 1587 1898 1591 1902
rect 1615 1898 1619 1902
rect 1645 1898 1649 1902
rect 1719 1898 1723 1902
rect 1747 1898 1751 1902
rect 1777 1898 1781 1902
rect 1851 1898 1855 1902
rect 1879 1898 1883 1902
rect 1909 1898 1913 1902
rect 182 1865 186 1869
rect 210 1865 214 1869
rect 240 1865 244 1869
rect 1115 1865 1119 1869
rect 1143 1865 1147 1869
rect 1173 1865 1177 1869
rect 503 1812 507 1816
rect 538 1812 542 1816
rect 664 1812 668 1816
rect 688 1812 692 1816
rect 742 1812 749 1816
rect 769 1812 773 1816
rect 823 1812 827 1816
rect 1436 1812 1440 1816
rect 1471 1812 1475 1816
rect 1597 1812 1601 1816
rect 1621 1812 1625 1816
rect 1675 1812 1682 1816
rect 1702 1812 1706 1816
rect 1756 1812 1760 1816
rect 179 1763 183 1767
rect 209 1763 213 1767
rect 237 1763 241 1767
rect 1112 1763 1116 1767
rect 1142 1763 1146 1767
rect 1170 1763 1174 1767
rect 503 1680 507 1684
rect 538 1680 542 1684
rect 664 1680 668 1684
rect 688 1680 692 1684
rect 742 1680 746 1684
rect 769 1680 773 1684
rect 793 1680 797 1684
rect 1436 1680 1440 1684
rect 1471 1680 1475 1684
rect 1597 1680 1601 1684
rect 1621 1680 1625 1684
rect 1675 1680 1679 1684
rect 1702 1680 1706 1684
rect 1726 1680 1730 1684
rect 503 1548 507 1552
rect 538 1548 542 1552
rect 664 1548 668 1552
rect 688 1548 692 1552
rect 742 1548 749 1552
rect 769 1548 773 1552
rect 823 1548 827 1552
rect 859 1548 863 1552
rect 913 1548 917 1552
rect 1436 1548 1440 1552
rect 1471 1548 1475 1552
rect 1597 1548 1601 1552
rect 1621 1548 1625 1552
rect 1675 1548 1682 1552
rect 1702 1548 1706 1552
rect 1756 1548 1760 1552
rect 1792 1548 1796 1552
rect 1846 1548 1850 1552
rect 503 1416 507 1420
rect 538 1416 542 1420
rect 664 1416 668 1420
rect 688 1416 692 1420
rect 799 1416 803 1420
rect 1436 1416 1440 1420
rect 1471 1416 1475 1420
rect 1597 1416 1601 1420
rect 1621 1416 1625 1420
rect 1732 1416 1736 1420
rect 50 1363 54 1367
rect 78 1363 82 1367
rect 108 1363 112 1367
rect 182 1363 186 1367
rect 210 1363 214 1367
rect 240 1363 244 1367
rect 314 1363 318 1367
rect 342 1363 346 1367
rect 372 1363 376 1367
rect 983 1363 987 1367
rect 1011 1363 1015 1367
rect 1041 1363 1045 1367
rect 1115 1363 1119 1367
rect 1143 1363 1147 1367
rect 1173 1363 1177 1367
rect 1247 1363 1251 1367
rect 1275 1363 1279 1367
rect 1305 1363 1309 1367
rect 821 1253 825 1257
rect 849 1253 853 1257
rect 879 1253 883 1257
rect 1754 1253 1758 1257
rect 1782 1253 1786 1257
rect 1812 1253 1816 1257
rect 50 1223 54 1227
rect 78 1223 82 1227
rect 108 1223 112 1227
rect 182 1223 186 1227
rect 210 1223 214 1227
rect 240 1223 244 1227
rect 314 1223 318 1227
rect 342 1223 346 1227
rect 372 1223 376 1227
rect 983 1223 987 1227
rect 1011 1223 1015 1227
rect 1041 1223 1045 1227
rect 1115 1223 1119 1227
rect 1143 1223 1147 1227
rect 1173 1223 1177 1227
rect 1247 1223 1251 1227
rect 1275 1223 1279 1227
rect 1305 1223 1309 1227
rect 821 1167 825 1171
rect 849 1167 853 1171
rect 879 1167 883 1171
rect 1754 1167 1758 1171
rect 1782 1167 1786 1171
rect 1812 1167 1816 1171
rect 50 1137 54 1141
rect 78 1137 82 1141
rect 108 1137 112 1141
rect 182 1137 186 1141
rect 210 1137 214 1141
rect 240 1137 244 1141
rect 314 1137 318 1141
rect 342 1137 346 1141
rect 372 1137 376 1141
rect 983 1137 987 1141
rect 1011 1137 1015 1141
rect 1041 1137 1045 1141
rect 1115 1137 1119 1141
rect 1143 1137 1147 1141
rect 1173 1137 1177 1141
rect 1247 1137 1251 1141
rect 1275 1137 1279 1141
rect 1305 1137 1309 1141
rect 50 997 54 1001
rect 78 997 82 1001
rect 108 997 112 1001
rect 182 997 186 1001
rect 210 997 214 1001
rect 240 997 244 1001
rect 314 997 318 1001
rect 342 997 346 1001
rect 372 997 376 1001
rect 983 997 987 1001
rect 1011 997 1015 1001
rect 1041 997 1045 1001
rect 1115 997 1119 1001
rect 1143 997 1147 1001
rect 1173 997 1177 1001
rect 1247 997 1251 1001
rect 1275 997 1279 1001
rect 1305 997 1309 1001
rect 522 918 526 922
rect 550 918 554 922
rect 580 918 584 922
rect 654 918 658 922
rect 682 918 686 922
rect 712 918 716 922
rect 786 918 790 922
rect 814 918 818 922
rect 844 918 848 922
rect 918 918 922 922
rect 946 918 950 922
rect 976 918 980 922
rect 1455 918 1459 922
rect 1483 918 1487 922
rect 1513 918 1517 922
rect 1587 918 1591 922
rect 1615 918 1619 922
rect 1645 918 1649 922
rect 1719 918 1723 922
rect 1747 918 1751 922
rect 1777 918 1781 922
rect 1851 918 1855 922
rect 1879 918 1883 922
rect 1909 918 1913 922
rect 182 885 186 889
rect 210 885 214 889
rect 240 885 244 889
rect 1115 885 1119 889
rect 1143 885 1147 889
rect 1173 885 1177 889
rect 503 832 507 836
rect 538 832 542 836
rect 664 832 668 836
rect 688 832 692 836
rect 742 832 749 836
rect 769 832 773 836
rect 823 832 827 836
rect 1436 832 1440 836
rect 1471 832 1475 836
rect 1597 832 1601 836
rect 1621 832 1625 836
rect 1675 832 1682 836
rect 1702 832 1706 836
rect 1756 832 1760 836
rect 179 783 183 787
rect 209 783 213 787
rect 237 783 241 787
rect 1112 783 1116 787
rect 1142 783 1146 787
rect 1170 783 1174 787
rect 503 700 507 704
rect 538 700 542 704
rect 664 700 668 704
rect 688 700 692 704
rect 742 700 746 704
rect 769 700 773 704
rect 793 700 797 704
rect 1436 700 1440 704
rect 1471 700 1475 704
rect 1597 700 1601 704
rect 1621 700 1625 704
rect 1675 700 1679 704
rect 1702 700 1706 704
rect 1726 700 1730 704
rect 503 568 507 572
rect 538 568 542 572
rect 664 568 668 572
rect 688 568 692 572
rect 742 568 749 572
rect 769 568 773 572
rect 823 568 827 572
rect 859 568 863 572
rect 913 568 917 572
rect 1436 568 1440 572
rect 1471 568 1475 572
rect 1597 568 1601 572
rect 1621 568 1625 572
rect 1675 568 1682 572
rect 1702 568 1706 572
rect 1756 568 1760 572
rect 1792 568 1796 572
rect 1846 568 1850 572
rect 503 436 507 440
rect 538 436 542 440
rect 664 436 668 440
rect 688 436 692 440
rect 799 436 803 440
rect 1436 436 1440 440
rect 1471 436 1475 440
rect 1597 436 1601 440
rect 1621 436 1625 440
rect 1732 436 1736 440
rect 50 383 54 387
rect 78 383 82 387
rect 108 383 112 387
rect 182 383 186 387
rect 210 383 214 387
rect 240 383 244 387
rect 314 383 318 387
rect 342 383 346 387
rect 372 383 376 387
rect 983 383 987 387
rect 1011 383 1015 387
rect 1041 383 1045 387
rect 1115 383 1119 387
rect 1143 383 1147 387
rect 1173 383 1177 387
rect 1247 383 1251 387
rect 1275 383 1279 387
rect 1305 383 1309 387
rect 821 273 825 277
rect 849 273 853 277
rect 879 273 883 277
rect 1754 273 1758 277
rect 1782 273 1786 277
rect 1812 273 1816 277
rect 50 243 54 247
rect 78 243 82 247
rect 108 243 112 247
rect 182 243 186 247
rect 210 243 214 247
rect 240 243 244 247
rect 314 243 318 247
rect 342 243 346 247
rect 372 243 376 247
rect 983 243 987 247
rect 1011 243 1015 247
rect 1041 243 1045 247
rect 1115 243 1119 247
rect 1143 243 1147 247
rect 1173 243 1177 247
rect 1247 243 1251 247
rect 1275 243 1279 247
rect 1305 243 1309 247
rect 821 187 825 191
rect 849 187 853 191
rect 879 187 883 191
rect 1754 187 1758 191
rect 1782 187 1786 191
rect 1812 187 1816 191
rect 50 157 54 161
rect 78 157 82 161
rect 108 157 112 161
rect 182 157 186 161
rect 210 157 214 161
rect 240 157 244 161
rect 314 157 318 161
rect 342 157 346 161
rect 372 157 376 161
rect 983 157 987 161
rect 1011 157 1015 161
rect 1041 157 1045 161
rect 1115 157 1119 161
rect 1143 157 1147 161
rect 1173 157 1177 161
rect 1247 157 1251 161
rect 1275 157 1279 161
rect 1305 157 1309 161
rect 50 17 54 21
rect 78 17 82 21
rect 108 17 112 21
rect 182 17 186 21
rect 210 17 214 21
rect 240 17 244 21
rect 314 17 318 21
rect 342 17 346 21
rect 372 17 376 21
rect 983 17 987 21
rect 1011 17 1015 21
rect 1041 17 1045 21
rect 1115 17 1119 21
rect 1143 17 1147 21
rect 1173 17 1177 21
rect 1247 17 1251 21
rect 1275 17 1279 21
rect 1305 17 1309 21
<< nsubstratencontact >>
rect 522 1955 526 1959
rect 550 1955 554 1959
rect 580 1955 584 1959
rect 617 1955 621 1959
rect 654 1955 658 1959
rect 682 1955 686 1959
rect 712 1955 716 1959
rect 749 1955 753 1959
rect 786 1955 790 1959
rect 814 1955 818 1959
rect 844 1955 848 1959
rect 881 1955 885 1959
rect 918 1955 922 1959
rect 946 1955 950 1959
rect 976 1955 980 1959
rect 1013 1955 1017 1959
rect 1455 1955 1459 1959
rect 1483 1955 1487 1959
rect 1513 1955 1517 1959
rect 1550 1955 1554 1959
rect 1587 1955 1591 1959
rect 1615 1955 1619 1959
rect 1645 1955 1649 1959
rect 1682 1955 1686 1959
rect 1719 1955 1723 1959
rect 1747 1955 1751 1959
rect 1777 1955 1781 1959
rect 1814 1955 1818 1959
rect 1851 1955 1855 1959
rect 1879 1955 1883 1959
rect 1909 1955 1913 1959
rect 1946 1955 1950 1959
rect 182 1922 186 1926
rect 210 1922 214 1926
rect 240 1922 244 1926
rect 277 1922 281 1926
rect 1115 1922 1119 1926
rect 1143 1922 1147 1926
rect 1173 1922 1177 1926
rect 1210 1922 1214 1926
rect 512 1878 516 1882
rect 541 1878 545 1882
rect 566 1878 570 1882
rect 608 1878 612 1882
rect 664 1878 668 1882
rect 688 1878 692 1882
rect 742 1878 746 1882
rect 769 1878 773 1882
rect 823 1878 827 1882
rect 1445 1878 1449 1882
rect 1474 1878 1478 1882
rect 1499 1878 1503 1882
rect 1541 1878 1545 1882
rect 1597 1878 1601 1882
rect 1621 1878 1625 1882
rect 1675 1878 1679 1882
rect 1702 1878 1706 1882
rect 1756 1878 1760 1882
rect 142 1820 146 1824
rect 179 1820 183 1824
rect 209 1820 213 1824
rect 237 1820 241 1824
rect 1075 1820 1079 1824
rect 1112 1820 1116 1824
rect 1142 1820 1146 1824
rect 1170 1820 1174 1824
rect 512 1746 516 1750
rect 541 1746 545 1750
rect 566 1746 570 1750
rect 608 1746 612 1750
rect 664 1746 668 1750
rect 688 1746 692 1750
rect 742 1746 746 1750
rect 769 1746 773 1750
rect 831 1746 835 1750
rect 1445 1746 1449 1750
rect 1474 1746 1478 1750
rect 1499 1746 1503 1750
rect 1541 1746 1545 1750
rect 1597 1746 1601 1750
rect 1621 1746 1625 1750
rect 1675 1746 1679 1750
rect 1702 1746 1706 1750
rect 1764 1746 1768 1750
rect 512 1614 516 1618
rect 541 1614 545 1618
rect 566 1614 570 1618
rect 608 1614 612 1618
rect 664 1614 668 1618
rect 688 1614 692 1618
rect 742 1614 746 1618
rect 769 1614 773 1618
rect 823 1614 827 1618
rect 831 1614 835 1618
rect 859 1614 863 1618
rect 913 1614 917 1618
rect 1445 1614 1449 1618
rect 1474 1614 1478 1618
rect 1499 1614 1503 1618
rect 1541 1614 1545 1618
rect 1597 1614 1601 1618
rect 1621 1614 1625 1618
rect 1675 1614 1679 1618
rect 1702 1614 1706 1618
rect 1756 1614 1760 1618
rect 1764 1614 1768 1618
rect 1792 1614 1796 1618
rect 1846 1614 1850 1618
rect 512 1482 516 1486
rect 541 1482 545 1486
rect 566 1482 570 1486
rect 608 1482 612 1486
rect 664 1482 668 1486
rect 688 1482 692 1486
rect 742 1482 746 1486
rect 769 1482 773 1486
rect 859 1482 863 1486
rect 1445 1482 1449 1486
rect 1474 1482 1478 1486
rect 1499 1482 1503 1486
rect 1541 1482 1545 1486
rect 1597 1482 1601 1486
rect 1621 1482 1625 1486
rect 1675 1482 1679 1486
rect 1702 1482 1706 1486
rect 1792 1482 1796 1486
rect 50 1420 54 1424
rect 78 1420 82 1424
rect 108 1420 112 1424
rect 145 1420 149 1424
rect 182 1420 186 1424
rect 210 1420 214 1424
rect 240 1420 244 1424
rect 277 1420 281 1424
rect 314 1420 318 1424
rect 342 1420 346 1424
rect 372 1420 376 1424
rect 409 1420 413 1424
rect 983 1420 987 1424
rect 1011 1420 1015 1424
rect 1041 1420 1045 1424
rect 1078 1420 1082 1424
rect 1115 1420 1119 1424
rect 1143 1420 1147 1424
rect 1173 1420 1177 1424
rect 1210 1420 1214 1424
rect 1247 1420 1251 1424
rect 1275 1420 1279 1424
rect 1305 1420 1309 1424
rect 1342 1420 1346 1424
rect 512 1350 516 1354
rect 541 1350 545 1354
rect 566 1350 570 1354
rect 608 1350 612 1354
rect 688 1350 692 1354
rect 742 1350 746 1354
rect 773 1350 777 1354
rect 802 1350 806 1354
rect 827 1350 831 1354
rect 869 1350 873 1354
rect 1445 1350 1449 1354
rect 1474 1350 1478 1354
rect 1499 1350 1503 1354
rect 1541 1350 1545 1354
rect 1621 1350 1625 1354
rect 1675 1350 1679 1354
rect 1706 1350 1710 1354
rect 1735 1350 1739 1354
rect 1760 1350 1764 1354
rect 1802 1350 1806 1354
rect 821 1310 825 1314
rect 849 1310 853 1314
rect 879 1310 883 1314
rect 916 1310 920 1314
rect 1754 1310 1758 1314
rect 1782 1310 1786 1314
rect 1812 1310 1816 1314
rect 1849 1310 1853 1314
rect 50 1280 54 1284
rect 78 1280 82 1284
rect 108 1280 112 1284
rect 145 1280 149 1284
rect 182 1280 186 1284
rect 210 1280 214 1284
rect 240 1280 244 1284
rect 277 1280 281 1284
rect 314 1280 318 1284
rect 342 1280 346 1284
rect 372 1280 376 1284
rect 409 1280 413 1284
rect 983 1280 987 1284
rect 1011 1280 1015 1284
rect 1041 1280 1045 1284
rect 1078 1280 1082 1284
rect 1115 1280 1119 1284
rect 1143 1280 1147 1284
rect 1173 1280 1177 1284
rect 1210 1280 1214 1284
rect 1247 1280 1251 1284
rect 1275 1280 1279 1284
rect 1305 1280 1309 1284
rect 1342 1280 1346 1284
rect 821 1224 825 1228
rect 849 1224 853 1228
rect 879 1224 883 1228
rect 916 1224 920 1228
rect 1754 1224 1758 1228
rect 1782 1224 1786 1228
rect 1812 1224 1816 1228
rect 1849 1224 1853 1228
rect 50 1194 54 1198
rect 78 1194 82 1198
rect 108 1194 112 1198
rect 145 1194 149 1198
rect 182 1194 186 1198
rect 210 1194 214 1198
rect 240 1194 244 1198
rect 277 1194 281 1198
rect 314 1194 318 1198
rect 342 1194 346 1198
rect 372 1194 376 1198
rect 409 1194 413 1198
rect 983 1194 987 1198
rect 1011 1194 1015 1198
rect 1041 1194 1045 1198
rect 1078 1194 1082 1198
rect 1115 1194 1119 1198
rect 1143 1194 1147 1198
rect 1173 1194 1177 1198
rect 1210 1194 1214 1198
rect 1247 1194 1251 1198
rect 1275 1194 1279 1198
rect 1305 1194 1309 1198
rect 1342 1194 1346 1198
rect 50 1054 54 1058
rect 78 1054 82 1058
rect 108 1054 112 1058
rect 145 1054 149 1058
rect 182 1054 186 1058
rect 210 1054 214 1058
rect 240 1054 244 1058
rect 277 1054 281 1058
rect 314 1054 318 1058
rect 342 1054 346 1058
rect 372 1054 376 1058
rect 409 1054 413 1058
rect 983 1054 987 1058
rect 1011 1054 1015 1058
rect 1041 1054 1045 1058
rect 1078 1054 1082 1058
rect 1115 1054 1119 1058
rect 1143 1054 1147 1058
rect 1173 1054 1177 1058
rect 1210 1054 1214 1058
rect 1247 1054 1251 1058
rect 1275 1054 1279 1058
rect 1305 1054 1309 1058
rect 1342 1054 1346 1058
rect 522 975 526 979
rect 550 975 554 979
rect 580 975 584 979
rect 617 975 621 979
rect 654 975 658 979
rect 682 975 686 979
rect 712 975 716 979
rect 749 975 753 979
rect 786 975 790 979
rect 814 975 818 979
rect 844 975 848 979
rect 881 975 885 979
rect 918 975 922 979
rect 946 975 950 979
rect 976 975 980 979
rect 1013 975 1017 979
rect 1455 975 1459 979
rect 1483 975 1487 979
rect 1513 975 1517 979
rect 1550 975 1554 979
rect 1587 975 1591 979
rect 1615 975 1619 979
rect 1645 975 1649 979
rect 1682 975 1686 979
rect 1719 975 1723 979
rect 1747 975 1751 979
rect 1777 975 1781 979
rect 1814 975 1818 979
rect 1851 975 1855 979
rect 1879 975 1883 979
rect 1909 975 1913 979
rect 1946 975 1950 979
rect 182 942 186 946
rect 210 942 214 946
rect 240 942 244 946
rect 277 942 281 946
rect 1115 942 1119 946
rect 1143 942 1147 946
rect 1173 942 1177 946
rect 1210 942 1214 946
rect 512 898 516 902
rect 541 898 545 902
rect 566 898 570 902
rect 608 898 612 902
rect 664 898 668 902
rect 688 898 692 902
rect 742 898 746 902
rect 769 898 773 902
rect 823 898 827 902
rect 1445 898 1449 902
rect 1474 898 1478 902
rect 1499 898 1503 902
rect 1541 898 1545 902
rect 1597 898 1601 902
rect 1621 898 1625 902
rect 1675 898 1679 902
rect 1702 898 1706 902
rect 1756 898 1760 902
rect 142 840 146 844
rect 179 840 183 844
rect 209 840 213 844
rect 237 840 241 844
rect 1075 840 1079 844
rect 1112 840 1116 844
rect 1142 840 1146 844
rect 1170 840 1174 844
rect 512 766 516 770
rect 541 766 545 770
rect 566 766 570 770
rect 608 766 612 770
rect 664 766 668 770
rect 688 766 692 770
rect 742 766 746 770
rect 769 766 773 770
rect 831 766 835 770
rect 1445 766 1449 770
rect 1474 766 1478 770
rect 1499 766 1503 770
rect 1541 766 1545 770
rect 1597 766 1601 770
rect 1621 766 1625 770
rect 1675 766 1679 770
rect 1702 766 1706 770
rect 1764 766 1768 770
rect 512 634 516 638
rect 541 634 545 638
rect 566 634 570 638
rect 608 634 612 638
rect 664 634 668 638
rect 688 634 692 638
rect 742 634 746 638
rect 769 634 773 638
rect 823 634 827 638
rect 831 634 835 638
rect 859 634 863 638
rect 913 634 917 638
rect 1445 634 1449 638
rect 1474 634 1478 638
rect 1499 634 1503 638
rect 1541 634 1545 638
rect 1597 634 1601 638
rect 1621 634 1625 638
rect 1675 634 1679 638
rect 1702 634 1706 638
rect 1756 634 1760 638
rect 1764 634 1768 638
rect 1792 634 1796 638
rect 1846 634 1850 638
rect 512 502 516 506
rect 541 502 545 506
rect 566 502 570 506
rect 608 502 612 506
rect 664 502 668 506
rect 688 502 692 506
rect 742 502 746 506
rect 769 502 773 506
rect 859 502 863 506
rect 1445 502 1449 506
rect 1474 502 1478 506
rect 1499 502 1503 506
rect 1541 502 1545 506
rect 1597 502 1601 506
rect 1621 502 1625 506
rect 1675 502 1679 506
rect 1702 502 1706 506
rect 1792 502 1796 506
rect 50 440 54 444
rect 78 440 82 444
rect 108 440 112 444
rect 145 440 149 444
rect 182 440 186 444
rect 210 440 214 444
rect 240 440 244 444
rect 277 440 281 444
rect 314 440 318 444
rect 342 440 346 444
rect 372 440 376 444
rect 409 440 413 444
rect 983 440 987 444
rect 1011 440 1015 444
rect 1041 440 1045 444
rect 1078 440 1082 444
rect 1115 440 1119 444
rect 1143 440 1147 444
rect 1173 440 1177 444
rect 1210 440 1214 444
rect 1247 440 1251 444
rect 1275 440 1279 444
rect 1305 440 1309 444
rect 1342 440 1346 444
rect 512 370 516 374
rect 541 370 545 374
rect 566 370 570 374
rect 608 370 612 374
rect 688 370 692 374
rect 742 370 746 374
rect 773 370 777 374
rect 802 370 806 374
rect 827 370 831 374
rect 869 370 873 374
rect 1445 370 1449 374
rect 1474 370 1478 374
rect 1499 370 1503 374
rect 1541 370 1545 374
rect 1621 370 1625 374
rect 1675 370 1679 374
rect 1706 370 1710 374
rect 1735 370 1739 374
rect 1760 370 1764 374
rect 1802 370 1806 374
rect 821 330 825 334
rect 849 330 853 334
rect 879 330 883 334
rect 916 330 920 334
rect 1754 330 1758 334
rect 1782 330 1786 334
rect 1812 330 1816 334
rect 1849 330 1853 334
rect 50 300 54 304
rect 78 300 82 304
rect 108 300 112 304
rect 145 300 149 304
rect 182 300 186 304
rect 210 300 214 304
rect 240 300 244 304
rect 277 300 281 304
rect 314 300 318 304
rect 342 300 346 304
rect 372 300 376 304
rect 409 300 413 304
rect 983 300 987 304
rect 1011 300 1015 304
rect 1041 300 1045 304
rect 1078 300 1082 304
rect 1115 300 1119 304
rect 1143 300 1147 304
rect 1173 300 1177 304
rect 1210 300 1214 304
rect 1247 300 1251 304
rect 1275 300 1279 304
rect 1305 300 1309 304
rect 1342 300 1346 304
rect 821 244 825 248
rect 849 244 853 248
rect 879 244 883 248
rect 916 244 920 248
rect 1754 244 1758 248
rect 1782 244 1786 248
rect 1812 244 1816 248
rect 1849 244 1853 248
rect 50 214 54 218
rect 78 214 82 218
rect 108 214 112 218
rect 145 214 149 218
rect 182 214 186 218
rect 210 214 214 218
rect 240 214 244 218
rect 277 214 281 218
rect 314 214 318 218
rect 342 214 346 218
rect 372 214 376 218
rect 409 214 413 218
rect 983 214 987 218
rect 1011 214 1015 218
rect 1041 214 1045 218
rect 1078 214 1082 218
rect 1115 214 1119 218
rect 1143 214 1147 218
rect 1173 214 1177 218
rect 1210 214 1214 218
rect 1247 214 1251 218
rect 1275 214 1279 218
rect 1305 214 1309 218
rect 1342 214 1346 218
rect 50 74 54 78
rect 78 74 82 78
rect 108 74 112 78
rect 145 74 149 78
rect 182 74 186 78
rect 210 74 214 78
rect 240 74 244 78
rect 277 74 281 78
rect 314 74 318 78
rect 342 74 346 78
rect 372 74 376 78
rect 409 74 413 78
rect 983 74 987 78
rect 1011 74 1015 78
rect 1041 74 1045 78
rect 1078 74 1082 78
rect 1115 74 1119 78
rect 1143 74 1147 78
rect 1173 74 1177 78
rect 1210 74 1214 78
rect 1247 74 1251 78
rect 1275 74 1279 78
rect 1305 74 1309 78
rect 1342 74 1346 78
<< polysilicon >>
rect 497 1945 499 1947
rect 502 1945 504 1948
rect 518 1945 520 1947
rect 534 1945 536 1947
rect 539 1945 541 1948
rect 560 1945 562 1948
rect 576 1945 578 1948
rect 592 1945 594 1947
rect 597 1945 599 1948
rect 613 1945 615 1947
rect 629 1945 631 1947
rect 634 1945 636 1948
rect 650 1945 652 1947
rect 666 1945 668 1947
rect 671 1945 673 1948
rect 692 1945 694 1948
rect 708 1945 710 1948
rect 724 1945 726 1947
rect 729 1945 731 1948
rect 745 1945 747 1947
rect 761 1945 763 1947
rect 766 1945 768 1948
rect 782 1945 784 1947
rect 798 1945 800 1947
rect 803 1945 805 1948
rect 824 1945 826 1948
rect 840 1945 842 1948
rect 856 1945 858 1947
rect 861 1945 863 1948
rect 877 1945 879 1947
rect 893 1945 895 1947
rect 898 1945 900 1948
rect 914 1945 916 1947
rect 930 1945 932 1947
rect 935 1945 937 1948
rect 956 1945 958 1948
rect 972 1945 974 1948
rect 988 1945 990 1947
rect 993 1945 995 1948
rect 1009 1945 1011 1947
rect 1430 1945 1432 1947
rect 1435 1945 1437 1948
rect 1451 1945 1453 1947
rect 1467 1945 1469 1947
rect 1472 1945 1474 1948
rect 1493 1945 1495 1948
rect 1509 1945 1511 1948
rect 1525 1945 1527 1947
rect 1530 1945 1532 1948
rect 1546 1945 1548 1947
rect 1562 1945 1564 1947
rect 1567 1945 1569 1948
rect 1583 1945 1585 1947
rect 1599 1945 1601 1947
rect 1604 1945 1606 1948
rect 1625 1945 1627 1948
rect 1641 1945 1643 1948
rect 1657 1945 1659 1947
rect 1662 1945 1664 1948
rect 1678 1945 1680 1947
rect 1694 1945 1696 1947
rect 1699 1945 1701 1948
rect 1715 1945 1717 1947
rect 1731 1945 1733 1947
rect 1736 1945 1738 1948
rect 1757 1945 1759 1948
rect 1773 1945 1775 1948
rect 1789 1945 1791 1947
rect 1794 1945 1796 1948
rect 1810 1945 1812 1947
rect 1826 1945 1828 1947
rect 1831 1945 1833 1948
rect 1847 1945 1849 1947
rect 1863 1945 1865 1947
rect 1868 1945 1870 1948
rect 1889 1945 1891 1948
rect 1905 1945 1907 1948
rect 1921 1945 1923 1947
rect 1926 1945 1928 1948
rect 1942 1945 1944 1947
rect 497 1932 499 1937
rect 502 1935 504 1937
rect 497 1918 499 1928
rect 502 1918 504 1925
rect 518 1918 520 1937
rect 534 1928 536 1937
rect 539 1935 541 1937
rect 560 1935 562 1937
rect 576 1934 578 1937
rect 534 1918 536 1921
rect 539 1918 541 1920
rect 560 1918 562 1920
rect 576 1918 578 1930
rect 592 1928 594 1937
rect 597 1935 599 1937
rect 613 1929 615 1937
rect 629 1932 631 1937
rect 634 1935 636 1937
rect 592 1918 594 1921
rect 597 1918 599 1920
rect 613 1918 615 1925
rect 629 1918 631 1928
rect 634 1918 636 1925
rect 650 1918 652 1937
rect 666 1928 668 1937
rect 671 1935 673 1937
rect 692 1935 694 1937
rect 708 1934 710 1937
rect 666 1918 668 1921
rect 671 1918 673 1920
rect 692 1918 694 1920
rect 708 1918 710 1930
rect 724 1928 726 1937
rect 729 1935 731 1937
rect 745 1929 747 1937
rect 761 1932 763 1937
rect 766 1935 768 1937
rect 724 1918 726 1921
rect 729 1918 731 1920
rect 745 1918 747 1925
rect 761 1918 763 1928
rect 766 1918 768 1925
rect 782 1918 784 1937
rect 798 1928 800 1937
rect 803 1935 805 1937
rect 824 1935 826 1937
rect 840 1934 842 1937
rect 798 1918 800 1921
rect 803 1918 805 1920
rect 824 1918 826 1920
rect 840 1918 842 1930
rect 856 1928 858 1937
rect 861 1935 863 1937
rect 877 1929 879 1937
rect 893 1932 895 1937
rect 898 1935 900 1937
rect 856 1918 858 1921
rect 861 1918 863 1920
rect 877 1918 879 1925
rect 893 1918 895 1928
rect 898 1918 900 1925
rect 914 1918 916 1937
rect 930 1928 932 1937
rect 935 1935 937 1937
rect 956 1935 958 1937
rect 972 1934 974 1937
rect 930 1918 932 1921
rect 935 1918 937 1920
rect 956 1918 958 1920
rect 972 1918 974 1930
rect 988 1928 990 1937
rect 993 1935 995 1937
rect 1009 1929 1011 1937
rect 1430 1932 1432 1937
rect 1435 1935 1437 1937
rect 988 1918 990 1921
rect 993 1918 995 1920
rect 1009 1918 1011 1925
rect 157 1912 159 1914
rect 162 1912 164 1915
rect 178 1912 180 1914
rect 194 1912 196 1914
rect 199 1912 201 1915
rect 220 1912 222 1915
rect 236 1912 238 1915
rect 252 1912 254 1914
rect 257 1912 259 1915
rect 1430 1918 1432 1928
rect 1435 1918 1437 1925
rect 1451 1918 1453 1937
rect 1467 1928 1469 1937
rect 1472 1935 1474 1937
rect 1493 1935 1495 1937
rect 1509 1934 1511 1937
rect 1467 1918 1469 1921
rect 1472 1918 1474 1920
rect 1493 1918 1495 1920
rect 1509 1918 1511 1930
rect 1525 1928 1527 1937
rect 1530 1935 1532 1937
rect 1546 1929 1548 1937
rect 1562 1932 1564 1937
rect 1567 1935 1569 1937
rect 1525 1918 1527 1921
rect 1530 1918 1532 1920
rect 1546 1918 1548 1925
rect 1562 1918 1564 1928
rect 1567 1918 1569 1925
rect 1583 1918 1585 1937
rect 1599 1928 1601 1937
rect 1604 1935 1606 1937
rect 1625 1935 1627 1937
rect 1641 1934 1643 1937
rect 1599 1918 1601 1921
rect 1604 1918 1606 1920
rect 1625 1918 1627 1920
rect 1641 1918 1643 1930
rect 1657 1928 1659 1937
rect 1662 1935 1664 1937
rect 1678 1929 1680 1937
rect 1694 1932 1696 1937
rect 1699 1935 1701 1937
rect 1657 1918 1659 1921
rect 1662 1918 1664 1920
rect 1678 1918 1680 1925
rect 1694 1918 1696 1928
rect 1699 1918 1701 1925
rect 1715 1918 1717 1937
rect 1731 1928 1733 1937
rect 1736 1935 1738 1937
rect 1757 1935 1759 1937
rect 1773 1934 1775 1937
rect 1731 1918 1733 1921
rect 1736 1918 1738 1920
rect 1757 1918 1759 1920
rect 1773 1918 1775 1930
rect 1789 1928 1791 1937
rect 1794 1935 1796 1937
rect 1810 1929 1812 1937
rect 1826 1932 1828 1937
rect 1831 1935 1833 1937
rect 1789 1918 1791 1921
rect 1794 1918 1796 1920
rect 1810 1918 1812 1925
rect 1826 1918 1828 1928
rect 1831 1918 1833 1925
rect 1847 1918 1849 1937
rect 1863 1928 1865 1937
rect 1868 1935 1870 1937
rect 1889 1935 1891 1937
rect 1905 1934 1907 1937
rect 1863 1918 1865 1921
rect 1868 1918 1870 1920
rect 1889 1918 1891 1920
rect 1905 1918 1907 1930
rect 1921 1928 1923 1937
rect 1926 1935 1928 1937
rect 1942 1929 1944 1937
rect 1921 1918 1923 1921
rect 1926 1918 1928 1920
rect 1942 1918 1944 1925
rect 273 1912 275 1914
rect 497 1912 499 1914
rect 502 1911 504 1914
rect 518 1912 520 1914
rect 534 1912 536 1914
rect 539 1909 541 1914
rect 560 1909 562 1914
rect 576 1912 578 1914
rect 592 1912 594 1914
rect 597 1909 599 1914
rect 613 1912 615 1914
rect 629 1912 631 1914
rect 634 1911 636 1914
rect 650 1912 652 1914
rect 666 1912 668 1914
rect 671 1909 673 1914
rect 692 1909 694 1914
rect 708 1912 710 1914
rect 724 1912 726 1914
rect 729 1909 731 1914
rect 745 1912 747 1914
rect 761 1912 763 1914
rect 766 1911 768 1914
rect 782 1912 784 1914
rect 798 1912 800 1914
rect 803 1909 805 1914
rect 824 1909 826 1914
rect 840 1912 842 1914
rect 856 1912 858 1914
rect 861 1909 863 1914
rect 877 1912 879 1914
rect 893 1912 895 1914
rect 898 1911 900 1914
rect 914 1912 916 1914
rect 930 1912 932 1914
rect 935 1909 937 1914
rect 956 1909 958 1914
rect 972 1912 974 1914
rect 988 1912 990 1914
rect 993 1909 995 1914
rect 1009 1912 1011 1914
rect 1090 1912 1092 1914
rect 1095 1912 1097 1915
rect 1111 1912 1113 1914
rect 1127 1912 1129 1914
rect 1132 1912 1134 1915
rect 1153 1912 1155 1915
rect 1169 1912 1171 1915
rect 1185 1912 1187 1914
rect 1190 1912 1192 1915
rect 1206 1912 1208 1914
rect 1430 1912 1432 1914
rect 1435 1911 1437 1914
rect 1451 1912 1453 1914
rect 1467 1912 1469 1914
rect 1472 1909 1474 1914
rect 1493 1909 1495 1914
rect 1509 1912 1511 1914
rect 1525 1912 1527 1914
rect 1530 1909 1532 1914
rect 1546 1912 1548 1914
rect 1562 1912 1564 1914
rect 1567 1911 1569 1914
rect 1583 1912 1585 1914
rect 1599 1912 1601 1914
rect 1604 1909 1606 1914
rect 1625 1909 1627 1914
rect 1641 1912 1643 1914
rect 1657 1912 1659 1914
rect 1662 1909 1664 1914
rect 1678 1912 1680 1914
rect 1694 1912 1696 1914
rect 1699 1911 1701 1914
rect 1715 1912 1717 1914
rect 1731 1912 1733 1914
rect 1736 1909 1738 1914
rect 1757 1909 1759 1914
rect 1773 1912 1775 1914
rect 1789 1912 1791 1914
rect 1794 1909 1796 1914
rect 1810 1912 1812 1914
rect 1826 1912 1828 1914
rect 1831 1911 1833 1914
rect 1847 1912 1849 1914
rect 1863 1912 1865 1914
rect 1868 1909 1870 1914
rect 1889 1909 1891 1914
rect 1905 1912 1907 1914
rect 1921 1912 1923 1914
rect 1926 1909 1928 1914
rect 1942 1912 1944 1914
rect 157 1899 159 1904
rect 162 1902 164 1904
rect 157 1885 159 1895
rect 162 1885 164 1892
rect 178 1885 180 1904
rect 194 1895 196 1904
rect 199 1902 201 1904
rect 220 1902 222 1904
rect 236 1901 238 1904
rect 194 1885 196 1888
rect 199 1885 201 1887
rect 220 1885 222 1887
rect 236 1885 238 1897
rect 252 1895 254 1904
rect 257 1902 259 1904
rect 252 1885 254 1888
rect 257 1885 259 1887
rect 273 1885 275 1904
rect 1090 1899 1092 1904
rect 1095 1902 1097 1904
rect 1090 1885 1092 1895
rect 1095 1885 1097 1892
rect 1111 1885 1113 1904
rect 1127 1895 1129 1904
rect 1132 1902 1134 1904
rect 1153 1902 1155 1904
rect 1169 1901 1171 1904
rect 1127 1885 1129 1888
rect 1132 1885 1134 1887
rect 1153 1885 1155 1887
rect 1169 1885 1171 1897
rect 1185 1895 1187 1904
rect 1190 1902 1192 1904
rect 1185 1885 1187 1888
rect 1190 1885 1192 1887
rect 1206 1885 1208 1904
rect 157 1879 159 1881
rect 162 1878 164 1881
rect 178 1879 180 1881
rect 194 1879 196 1881
rect 199 1876 201 1881
rect 220 1876 222 1881
rect 236 1879 238 1881
rect 252 1879 254 1881
rect 257 1876 259 1881
rect 273 1879 275 1881
rect 1090 1879 1092 1881
rect 1095 1878 1097 1881
rect 1111 1879 1113 1881
rect 1127 1879 1129 1881
rect 676 1874 678 1876
rect 518 1868 520 1871
rect 562 1868 564 1871
rect 588 1868 590 1871
rect 634 1868 636 1871
rect 588 1864 589 1868
rect 702 1868 704 1872
rect 730 1874 732 1876
rect 757 1874 759 1876
rect 707 1868 709 1871
rect 502 1861 504 1863
rect 518 1861 520 1864
rect 534 1861 536 1863
rect 557 1861 559 1863
rect 562 1861 564 1864
rect 588 1861 590 1864
rect 609 1861 611 1864
rect 629 1861 631 1863
rect 634 1861 636 1864
rect 652 1861 654 1863
rect 281 1848 283 1851
rect 281 1842 283 1844
rect 164 1839 166 1842
rect 502 1839 504 1853
rect 518 1851 520 1853
rect 518 1839 520 1841
rect 534 1839 536 1853
rect 557 1848 559 1853
rect 562 1851 564 1853
rect 588 1851 590 1853
rect 553 1844 559 1848
rect 557 1839 559 1844
rect 562 1839 564 1841
rect 588 1839 590 1841
rect 609 1839 611 1853
rect 629 1848 631 1853
rect 634 1851 636 1853
rect 625 1844 631 1848
rect 629 1839 631 1844
rect 634 1839 636 1841
rect 652 1839 654 1853
rect 676 1852 678 1866
rect 783 1868 785 1872
rect 811 1874 813 1876
rect 1132 1876 1134 1881
rect 1153 1876 1155 1881
rect 1169 1879 1171 1881
rect 1185 1879 1187 1881
rect 1190 1876 1192 1881
rect 1206 1879 1208 1881
rect 788 1868 790 1871
rect 702 1857 704 1860
rect 707 1858 709 1860
rect 703 1853 704 1857
rect 702 1848 704 1853
rect 707 1848 709 1850
rect 676 1846 678 1848
rect 730 1844 732 1866
rect 757 1852 759 1866
rect 1609 1874 1611 1876
rect 783 1857 785 1860
rect 788 1858 790 1860
rect 784 1853 785 1857
rect 783 1848 785 1853
rect 788 1848 790 1850
rect 757 1846 759 1848
rect 811 1844 813 1866
rect 1451 1868 1453 1871
rect 1495 1868 1497 1871
rect 1521 1868 1523 1871
rect 1567 1868 1569 1871
rect 1521 1864 1522 1868
rect 1635 1868 1637 1872
rect 1663 1874 1665 1876
rect 1690 1874 1692 1876
rect 1640 1868 1642 1871
rect 1435 1861 1437 1863
rect 1451 1861 1453 1864
rect 1467 1861 1469 1863
rect 1490 1861 1492 1863
rect 1495 1861 1497 1864
rect 1521 1861 1523 1864
rect 1542 1861 1544 1864
rect 1562 1861 1564 1863
rect 1567 1861 1569 1864
rect 1585 1861 1587 1863
rect 1214 1848 1216 1851
rect 702 1842 704 1844
rect 707 1839 709 1844
rect 783 1842 785 1844
rect 730 1838 732 1840
rect 788 1839 790 1844
rect 1214 1842 1216 1844
rect 811 1838 813 1840
rect 1097 1839 1099 1842
rect 1435 1839 1437 1853
rect 1451 1851 1453 1853
rect 1451 1839 1453 1841
rect 1467 1839 1469 1853
rect 1490 1848 1492 1853
rect 1495 1851 1497 1853
rect 1521 1851 1523 1853
rect 1486 1844 1492 1848
rect 1490 1839 1492 1844
rect 1495 1839 1497 1841
rect 1521 1839 1523 1841
rect 1542 1839 1544 1853
rect 1562 1848 1564 1853
rect 1567 1851 1569 1853
rect 1558 1844 1564 1848
rect 1562 1839 1564 1844
rect 1567 1839 1569 1841
rect 1585 1839 1587 1853
rect 1609 1852 1611 1866
rect 1716 1868 1718 1872
rect 1744 1874 1746 1876
rect 1721 1868 1723 1871
rect 1635 1857 1637 1860
rect 1640 1858 1642 1860
rect 1636 1853 1637 1857
rect 1635 1848 1637 1853
rect 1640 1848 1642 1850
rect 1609 1846 1611 1848
rect 1663 1844 1665 1866
rect 1690 1852 1692 1866
rect 1716 1857 1718 1860
rect 1721 1858 1723 1860
rect 1717 1853 1718 1857
rect 1716 1848 1718 1853
rect 1721 1848 1723 1850
rect 1690 1846 1692 1848
rect 1744 1844 1746 1866
rect 1635 1842 1637 1844
rect 1640 1839 1642 1844
rect 1716 1842 1718 1844
rect 1663 1838 1665 1840
rect 1721 1839 1723 1844
rect 1744 1838 1746 1840
rect 164 1833 166 1835
rect 502 1833 504 1835
rect 518 1831 520 1835
rect 534 1833 536 1835
rect 557 1833 559 1835
rect 519 1827 520 1831
rect 562 1830 564 1835
rect 588 1831 590 1835
rect 609 1833 611 1835
rect 629 1833 631 1835
rect 518 1824 520 1827
rect 563 1826 564 1830
rect 589 1827 590 1831
rect 634 1830 636 1835
rect 652 1833 654 1835
rect 1097 1833 1099 1835
rect 1435 1833 1437 1835
rect 1451 1831 1453 1835
rect 1467 1833 1469 1835
rect 1490 1833 1492 1835
rect 562 1824 564 1826
rect 588 1823 590 1827
rect 635 1826 636 1830
rect 1452 1827 1453 1831
rect 1495 1830 1497 1835
rect 1521 1831 1523 1835
rect 1542 1833 1544 1835
rect 1562 1833 1564 1835
rect 634 1824 636 1826
rect 1451 1824 1453 1827
rect 1496 1826 1497 1830
rect 1522 1827 1523 1831
rect 1567 1830 1569 1835
rect 1585 1833 1587 1835
rect 1495 1824 1497 1826
rect 1521 1823 1523 1827
rect 1568 1826 1569 1830
rect 1567 1824 1569 1826
rect 148 1810 150 1812
rect 164 1810 166 1813
rect 169 1810 171 1812
rect 185 1810 187 1813
rect 201 1810 203 1813
rect 222 1810 224 1813
rect 227 1810 229 1812
rect 243 1810 245 1812
rect 259 1810 261 1813
rect 264 1810 266 1812
rect 1081 1810 1083 1812
rect 1097 1810 1099 1813
rect 1102 1810 1104 1812
rect 1118 1810 1120 1813
rect 1134 1810 1136 1813
rect 1155 1810 1157 1813
rect 1160 1810 1162 1812
rect 1176 1810 1178 1812
rect 1192 1810 1194 1813
rect 1197 1810 1199 1812
rect 148 1783 150 1802
rect 164 1800 166 1802
rect 169 1793 171 1802
rect 185 1799 187 1802
rect 201 1800 203 1802
rect 222 1800 224 1802
rect 164 1783 166 1785
rect 169 1783 171 1786
rect 185 1783 187 1795
rect 227 1793 229 1802
rect 201 1783 203 1785
rect 222 1783 224 1785
rect 227 1783 229 1786
rect 243 1783 245 1802
rect 259 1800 261 1802
rect 264 1797 266 1802
rect 518 1801 520 1804
rect 562 1802 564 1804
rect 519 1797 520 1801
rect 563 1798 564 1802
rect 588 1801 590 1805
rect 634 1802 636 1804
rect 502 1793 504 1795
rect 518 1793 520 1797
rect 534 1793 536 1795
rect 557 1793 559 1795
rect 562 1793 564 1798
rect 589 1797 590 1801
rect 635 1798 636 1802
rect 588 1793 590 1797
rect 609 1793 611 1795
rect 629 1793 631 1795
rect 634 1793 636 1798
rect 652 1793 654 1795
rect 259 1783 261 1790
rect 264 1783 266 1793
rect 702 1792 704 1795
rect 707 1792 709 1795
rect 783 1792 785 1795
rect 788 1792 790 1795
rect 148 1777 150 1779
rect 164 1774 166 1779
rect 169 1777 171 1779
rect 185 1777 187 1779
rect 201 1774 203 1779
rect 222 1774 224 1779
rect 227 1777 229 1779
rect 243 1777 245 1779
rect 259 1776 261 1779
rect 264 1777 266 1779
rect 502 1775 504 1789
rect 518 1787 520 1789
rect 518 1775 520 1777
rect 534 1775 536 1789
rect 557 1784 559 1789
rect 562 1787 564 1789
rect 588 1787 590 1789
rect 553 1780 559 1784
rect 557 1775 559 1780
rect 562 1775 564 1777
rect 588 1775 590 1777
rect 609 1775 611 1789
rect 629 1784 631 1789
rect 634 1787 636 1789
rect 625 1780 631 1784
rect 629 1775 631 1780
rect 634 1775 636 1777
rect 652 1775 654 1789
rect 702 1776 704 1788
rect 707 1786 709 1788
rect 707 1776 709 1778
rect 783 1776 785 1788
rect 788 1786 790 1788
rect 1081 1783 1083 1802
rect 1097 1800 1099 1802
rect 1102 1793 1104 1802
rect 1118 1799 1120 1802
rect 1134 1800 1136 1802
rect 1155 1800 1157 1802
rect 1097 1783 1099 1785
rect 1102 1783 1104 1786
rect 1118 1783 1120 1795
rect 1160 1793 1162 1802
rect 1134 1783 1136 1785
rect 1155 1783 1157 1785
rect 1160 1783 1162 1786
rect 1176 1783 1178 1802
rect 1192 1800 1194 1802
rect 1197 1797 1199 1802
rect 1451 1801 1453 1804
rect 1495 1802 1497 1804
rect 1452 1797 1453 1801
rect 1496 1798 1497 1802
rect 1521 1801 1523 1805
rect 1567 1802 1569 1804
rect 1435 1793 1437 1795
rect 1451 1793 1453 1797
rect 1467 1793 1469 1795
rect 1490 1793 1492 1795
rect 1495 1793 1497 1798
rect 1522 1797 1523 1801
rect 1568 1798 1569 1802
rect 1521 1793 1523 1797
rect 1542 1793 1544 1795
rect 1562 1793 1564 1795
rect 1567 1793 1569 1798
rect 1585 1793 1587 1795
rect 1192 1783 1194 1790
rect 1197 1783 1199 1793
rect 1635 1792 1637 1795
rect 1640 1792 1642 1795
rect 1716 1792 1718 1795
rect 1721 1792 1723 1795
rect 788 1776 790 1778
rect 1081 1777 1083 1779
rect 1097 1774 1099 1779
rect 1102 1777 1104 1779
rect 1118 1777 1120 1779
rect 1134 1774 1136 1779
rect 1155 1774 1157 1779
rect 1160 1777 1162 1779
rect 1176 1777 1178 1779
rect 1192 1776 1194 1779
rect 1197 1777 1199 1779
rect 1435 1775 1437 1789
rect 1451 1787 1453 1789
rect 1451 1775 1453 1777
rect 1467 1775 1469 1789
rect 1490 1784 1492 1789
rect 1495 1787 1497 1789
rect 1521 1787 1523 1789
rect 1486 1780 1492 1784
rect 1490 1775 1492 1780
rect 1495 1775 1497 1777
rect 1521 1775 1523 1777
rect 1542 1775 1544 1789
rect 1562 1784 1564 1789
rect 1567 1787 1569 1789
rect 1558 1780 1564 1784
rect 1562 1775 1564 1780
rect 1567 1775 1569 1777
rect 1585 1775 1587 1789
rect 1635 1776 1637 1788
rect 1640 1786 1642 1788
rect 1640 1776 1642 1778
rect 1716 1776 1718 1788
rect 1721 1786 1723 1788
rect 1721 1776 1723 1778
rect 502 1765 504 1767
rect 518 1764 520 1767
rect 534 1765 536 1767
rect 557 1765 559 1767
rect 562 1764 564 1767
rect 588 1764 590 1767
rect 609 1764 611 1767
rect 629 1765 631 1767
rect 634 1764 636 1767
rect 652 1765 654 1767
rect 702 1766 704 1768
rect 588 1760 589 1764
rect 707 1763 709 1768
rect 783 1766 785 1768
rect 788 1763 790 1768
rect 1435 1765 1437 1767
rect 1451 1764 1453 1767
rect 1467 1765 1469 1767
rect 1490 1765 1492 1767
rect 1495 1764 1497 1767
rect 1521 1764 1523 1767
rect 1542 1764 1544 1767
rect 1562 1765 1564 1767
rect 1567 1764 1569 1767
rect 1585 1765 1587 1767
rect 1635 1766 1637 1768
rect 518 1757 520 1760
rect 562 1757 564 1760
rect 588 1757 590 1760
rect 634 1757 636 1760
rect 1521 1760 1522 1764
rect 1640 1763 1642 1768
rect 1716 1766 1718 1768
rect 1721 1763 1723 1768
rect 1451 1757 1453 1760
rect 1495 1757 1497 1760
rect 1521 1757 1523 1760
rect 1567 1757 1569 1760
rect 518 1736 520 1739
rect 562 1736 564 1739
rect 588 1736 590 1739
rect 634 1736 636 1739
rect 702 1736 704 1740
rect 730 1742 732 1744
rect 781 1742 783 1744
rect 707 1736 709 1739
rect 588 1732 589 1736
rect 502 1729 504 1731
rect 518 1729 520 1732
rect 534 1729 536 1731
rect 557 1729 559 1731
rect 562 1729 564 1732
rect 588 1729 590 1732
rect 609 1729 611 1732
rect 629 1729 631 1731
rect 634 1729 636 1732
rect 652 1729 654 1731
rect 807 1736 809 1740
rect 835 1742 837 1744
rect 812 1736 814 1739
rect 702 1725 704 1728
rect 707 1726 709 1728
rect 703 1721 704 1725
rect 502 1707 504 1721
rect 518 1719 520 1721
rect 518 1707 520 1709
rect 534 1707 536 1721
rect 557 1716 559 1721
rect 562 1719 564 1721
rect 588 1719 590 1721
rect 553 1712 559 1716
rect 557 1707 559 1712
rect 562 1707 564 1709
rect 588 1707 590 1709
rect 609 1707 611 1721
rect 629 1716 631 1721
rect 634 1719 636 1721
rect 625 1712 631 1716
rect 629 1707 631 1712
rect 634 1707 636 1709
rect 652 1707 654 1721
rect 702 1716 704 1721
rect 707 1716 709 1718
rect 730 1712 732 1734
rect 781 1720 783 1734
rect 1451 1736 1453 1739
rect 1495 1736 1497 1739
rect 1521 1736 1523 1739
rect 1567 1736 1569 1739
rect 1635 1736 1637 1740
rect 1663 1742 1665 1744
rect 1714 1742 1716 1744
rect 1640 1736 1642 1739
rect 807 1725 809 1728
rect 812 1726 814 1728
rect 808 1721 809 1725
rect 807 1716 809 1721
rect 812 1716 814 1718
rect 781 1714 783 1716
rect 835 1712 837 1734
rect 1521 1732 1522 1736
rect 1435 1729 1437 1731
rect 1451 1729 1453 1732
rect 1467 1729 1469 1731
rect 1490 1729 1492 1731
rect 1495 1729 1497 1732
rect 1521 1729 1523 1732
rect 1542 1729 1544 1732
rect 1562 1729 1564 1731
rect 1567 1729 1569 1732
rect 1585 1729 1587 1731
rect 1740 1736 1742 1740
rect 1768 1742 1770 1744
rect 1745 1736 1747 1739
rect 1635 1725 1637 1728
rect 1640 1726 1642 1728
rect 1636 1721 1637 1725
rect 702 1710 704 1712
rect 707 1707 709 1712
rect 807 1710 809 1712
rect 730 1706 732 1708
rect 812 1707 814 1712
rect 835 1706 837 1708
rect 1435 1707 1437 1721
rect 1451 1719 1453 1721
rect 1451 1707 1453 1709
rect 1467 1707 1469 1721
rect 1490 1716 1492 1721
rect 1495 1719 1497 1721
rect 1521 1719 1523 1721
rect 1486 1712 1492 1716
rect 1490 1707 1492 1712
rect 1495 1707 1497 1709
rect 1521 1707 1523 1709
rect 1542 1707 1544 1721
rect 1562 1716 1564 1721
rect 1567 1719 1569 1721
rect 1558 1712 1564 1716
rect 1562 1707 1564 1712
rect 1567 1707 1569 1709
rect 1585 1707 1587 1721
rect 1635 1716 1637 1721
rect 1640 1716 1642 1718
rect 1663 1712 1665 1734
rect 1714 1720 1716 1734
rect 1740 1725 1742 1728
rect 1745 1726 1747 1728
rect 1741 1721 1742 1725
rect 1740 1716 1742 1721
rect 1745 1716 1747 1718
rect 1714 1714 1716 1716
rect 1768 1712 1770 1734
rect 1635 1710 1637 1712
rect 1640 1707 1642 1712
rect 1740 1710 1742 1712
rect 1663 1706 1665 1708
rect 1745 1707 1747 1712
rect 1768 1706 1770 1708
rect 502 1701 504 1703
rect 518 1699 520 1703
rect 534 1701 536 1703
rect 557 1701 559 1703
rect 519 1695 520 1699
rect 562 1698 564 1703
rect 588 1699 590 1703
rect 609 1701 611 1703
rect 629 1701 631 1703
rect 518 1692 520 1695
rect 563 1694 564 1698
rect 589 1695 590 1699
rect 634 1698 636 1703
rect 652 1701 654 1703
rect 1435 1701 1437 1703
rect 1451 1699 1453 1703
rect 1467 1701 1469 1703
rect 1490 1701 1492 1703
rect 562 1692 564 1694
rect 588 1691 590 1695
rect 635 1694 636 1698
rect 1452 1695 1453 1699
rect 1495 1698 1497 1703
rect 1521 1699 1523 1703
rect 1542 1701 1544 1703
rect 1562 1701 1564 1703
rect 634 1692 636 1694
rect 1451 1692 1453 1695
rect 1496 1694 1497 1698
rect 1522 1695 1523 1699
rect 1567 1698 1569 1703
rect 1585 1701 1587 1703
rect 1495 1692 1497 1694
rect 1521 1691 1523 1695
rect 1568 1694 1569 1698
rect 1567 1692 1569 1694
rect 518 1669 520 1672
rect 562 1670 564 1672
rect 519 1665 520 1669
rect 563 1666 564 1670
rect 588 1669 590 1673
rect 634 1670 636 1672
rect 502 1661 504 1663
rect 518 1661 520 1665
rect 534 1661 536 1663
rect 557 1661 559 1663
rect 562 1661 564 1666
rect 589 1665 590 1669
rect 635 1666 636 1670
rect 1451 1669 1453 1672
rect 1495 1670 1497 1672
rect 588 1661 590 1665
rect 609 1661 611 1663
rect 629 1661 631 1663
rect 634 1661 636 1666
rect 1452 1665 1453 1669
rect 1496 1666 1497 1670
rect 1521 1669 1523 1673
rect 1567 1670 1569 1672
rect 652 1661 654 1663
rect 702 1661 704 1664
rect 707 1661 709 1664
rect 807 1661 809 1664
rect 812 1661 814 1664
rect 1435 1661 1437 1663
rect 1451 1661 1453 1665
rect 1467 1661 1469 1663
rect 1490 1661 1492 1663
rect 1495 1661 1497 1666
rect 1522 1665 1523 1669
rect 1568 1666 1569 1670
rect 1521 1661 1523 1665
rect 1542 1661 1544 1663
rect 1562 1661 1564 1663
rect 1567 1661 1569 1666
rect 1585 1661 1587 1663
rect 1635 1661 1637 1664
rect 1640 1661 1642 1664
rect 1740 1661 1742 1664
rect 1745 1661 1747 1664
rect 502 1643 504 1657
rect 518 1655 520 1657
rect 518 1643 520 1645
rect 534 1643 536 1657
rect 557 1652 559 1657
rect 562 1655 564 1657
rect 588 1655 590 1657
rect 553 1648 559 1652
rect 557 1643 559 1648
rect 562 1643 564 1645
rect 588 1643 590 1645
rect 609 1643 611 1657
rect 629 1652 631 1657
rect 634 1655 636 1657
rect 625 1648 631 1652
rect 629 1643 631 1648
rect 634 1643 636 1645
rect 652 1643 654 1657
rect 702 1645 704 1657
rect 707 1655 709 1657
rect 707 1645 709 1647
rect 807 1645 809 1657
rect 812 1655 814 1657
rect 812 1645 814 1647
rect 1435 1643 1437 1657
rect 1451 1655 1453 1657
rect 1451 1643 1453 1645
rect 1467 1643 1469 1657
rect 1490 1652 1492 1657
rect 1495 1655 1497 1657
rect 1521 1655 1523 1657
rect 1486 1648 1492 1652
rect 1490 1643 1492 1648
rect 1495 1643 1497 1645
rect 1521 1643 1523 1645
rect 1542 1643 1544 1657
rect 1562 1652 1564 1657
rect 1567 1655 1569 1657
rect 1558 1648 1564 1652
rect 1562 1643 1564 1648
rect 1567 1643 1569 1645
rect 1585 1643 1587 1657
rect 1635 1645 1637 1657
rect 1640 1655 1642 1657
rect 1640 1645 1642 1647
rect 1740 1645 1742 1657
rect 1745 1655 1747 1657
rect 1745 1645 1747 1647
rect 702 1635 704 1637
rect 502 1633 504 1635
rect 518 1632 520 1635
rect 534 1633 536 1635
rect 557 1633 559 1635
rect 562 1632 564 1635
rect 588 1632 590 1635
rect 609 1632 611 1635
rect 629 1633 631 1635
rect 634 1632 636 1635
rect 652 1633 654 1635
rect 707 1632 709 1637
rect 807 1635 809 1637
rect 812 1632 814 1637
rect 1635 1635 1637 1637
rect 1435 1633 1437 1635
rect 588 1628 589 1632
rect 1451 1632 1453 1635
rect 1467 1633 1469 1635
rect 1490 1633 1492 1635
rect 1495 1632 1497 1635
rect 1521 1632 1523 1635
rect 1542 1632 1544 1635
rect 1562 1633 1564 1635
rect 1567 1632 1569 1635
rect 1585 1633 1587 1635
rect 1640 1632 1642 1637
rect 1740 1635 1742 1637
rect 1745 1632 1747 1637
rect 1521 1628 1522 1632
rect 518 1625 520 1628
rect 562 1625 564 1628
rect 588 1625 590 1628
rect 634 1625 636 1628
rect 1451 1625 1453 1628
rect 1495 1625 1497 1628
rect 1521 1625 1523 1628
rect 1567 1625 1569 1628
rect 518 1604 520 1607
rect 562 1604 564 1607
rect 588 1604 590 1607
rect 634 1604 636 1607
rect 702 1604 704 1608
rect 730 1610 732 1612
rect 757 1610 759 1612
rect 707 1604 709 1607
rect 588 1600 589 1604
rect 502 1597 504 1599
rect 518 1597 520 1600
rect 534 1597 536 1599
rect 557 1597 559 1599
rect 562 1597 564 1600
rect 588 1597 590 1600
rect 609 1597 611 1600
rect 629 1597 631 1599
rect 634 1597 636 1600
rect 652 1597 654 1599
rect 783 1604 785 1608
rect 811 1610 813 1612
rect 847 1610 849 1612
rect 788 1604 790 1607
rect 702 1593 704 1596
rect 707 1594 709 1596
rect 703 1589 704 1593
rect 502 1575 504 1589
rect 518 1587 520 1589
rect 518 1575 520 1577
rect 534 1575 536 1589
rect 557 1584 559 1589
rect 562 1587 564 1589
rect 588 1587 590 1589
rect 553 1580 559 1584
rect 557 1575 559 1580
rect 562 1575 564 1577
rect 588 1575 590 1577
rect 609 1575 611 1589
rect 629 1584 631 1589
rect 634 1587 636 1589
rect 625 1580 631 1584
rect 629 1575 631 1580
rect 634 1575 636 1577
rect 652 1575 654 1589
rect 702 1584 704 1589
rect 707 1584 709 1586
rect 730 1580 732 1602
rect 757 1588 759 1602
rect 873 1604 875 1608
rect 901 1610 903 1612
rect 878 1604 880 1607
rect 783 1593 785 1596
rect 788 1594 790 1596
rect 784 1589 785 1593
rect 783 1584 785 1589
rect 788 1584 790 1586
rect 757 1582 759 1584
rect 811 1580 813 1602
rect 847 1588 849 1602
rect 1451 1604 1453 1607
rect 1495 1604 1497 1607
rect 1521 1604 1523 1607
rect 1567 1604 1569 1607
rect 1635 1604 1637 1608
rect 1663 1610 1665 1612
rect 1690 1610 1692 1612
rect 1640 1604 1642 1607
rect 873 1593 875 1596
rect 878 1594 880 1596
rect 874 1589 875 1593
rect 873 1584 875 1589
rect 878 1584 880 1586
rect 847 1582 849 1584
rect 901 1580 903 1602
rect 1521 1600 1522 1604
rect 1435 1597 1437 1599
rect 1451 1597 1453 1600
rect 1467 1597 1469 1599
rect 1490 1597 1492 1599
rect 1495 1597 1497 1600
rect 1521 1597 1523 1600
rect 1542 1597 1544 1600
rect 1562 1597 1564 1599
rect 1567 1597 1569 1600
rect 1585 1597 1587 1599
rect 1716 1604 1718 1608
rect 1744 1610 1746 1612
rect 1780 1610 1782 1612
rect 1721 1604 1723 1607
rect 1635 1593 1637 1596
rect 1640 1594 1642 1596
rect 1636 1589 1637 1593
rect 702 1578 704 1580
rect 707 1575 709 1580
rect 783 1578 785 1580
rect 730 1574 732 1576
rect 788 1575 790 1580
rect 873 1578 875 1580
rect 811 1574 813 1576
rect 878 1575 880 1580
rect 901 1574 903 1576
rect 1435 1575 1437 1589
rect 1451 1587 1453 1589
rect 1451 1575 1453 1577
rect 1467 1575 1469 1589
rect 1490 1584 1492 1589
rect 1495 1587 1497 1589
rect 1521 1587 1523 1589
rect 1486 1580 1492 1584
rect 1490 1575 1492 1580
rect 1495 1575 1497 1577
rect 1521 1575 1523 1577
rect 1542 1575 1544 1589
rect 1562 1584 1564 1589
rect 1567 1587 1569 1589
rect 1558 1580 1564 1584
rect 1562 1575 1564 1580
rect 1567 1575 1569 1577
rect 1585 1575 1587 1589
rect 1635 1584 1637 1589
rect 1640 1584 1642 1586
rect 1663 1580 1665 1602
rect 1690 1588 1692 1602
rect 1806 1604 1808 1608
rect 1834 1610 1836 1612
rect 1811 1604 1813 1607
rect 1716 1593 1718 1596
rect 1721 1594 1723 1596
rect 1717 1589 1718 1593
rect 1716 1584 1718 1589
rect 1721 1584 1723 1586
rect 1690 1582 1692 1584
rect 1744 1580 1746 1602
rect 1780 1588 1782 1602
rect 1806 1593 1808 1596
rect 1811 1594 1813 1596
rect 1807 1589 1808 1593
rect 1806 1584 1808 1589
rect 1811 1584 1813 1586
rect 1780 1582 1782 1584
rect 1834 1580 1836 1602
rect 1635 1578 1637 1580
rect 1640 1575 1642 1580
rect 1716 1578 1718 1580
rect 1663 1574 1665 1576
rect 1721 1575 1723 1580
rect 1806 1578 1808 1580
rect 1744 1574 1746 1576
rect 1811 1575 1813 1580
rect 1834 1574 1836 1576
rect 502 1569 504 1571
rect 518 1567 520 1571
rect 534 1569 536 1571
rect 557 1569 559 1571
rect 519 1563 520 1567
rect 562 1566 564 1571
rect 588 1567 590 1571
rect 609 1569 611 1571
rect 629 1569 631 1571
rect 518 1560 520 1563
rect 563 1562 564 1566
rect 589 1563 590 1567
rect 634 1566 636 1571
rect 652 1569 654 1571
rect 1435 1569 1437 1571
rect 1451 1567 1453 1571
rect 1467 1569 1469 1571
rect 1490 1569 1492 1571
rect 562 1560 564 1562
rect 588 1559 590 1563
rect 635 1562 636 1566
rect 1452 1563 1453 1567
rect 1495 1566 1497 1571
rect 1521 1567 1523 1571
rect 1542 1569 1544 1571
rect 1562 1569 1564 1571
rect 634 1560 636 1562
rect 1451 1560 1453 1563
rect 1496 1562 1497 1566
rect 1522 1563 1523 1567
rect 1567 1566 1569 1571
rect 1585 1569 1587 1571
rect 1495 1560 1497 1562
rect 1521 1559 1523 1563
rect 1568 1562 1569 1566
rect 1567 1560 1569 1562
rect 518 1537 520 1540
rect 562 1538 564 1540
rect 519 1533 520 1537
rect 563 1534 564 1538
rect 588 1537 590 1541
rect 634 1538 636 1540
rect 502 1529 504 1531
rect 518 1529 520 1533
rect 534 1529 536 1531
rect 557 1529 559 1531
rect 562 1529 564 1534
rect 589 1533 590 1537
rect 635 1534 636 1538
rect 1451 1537 1453 1540
rect 1495 1538 1497 1540
rect 588 1529 590 1533
rect 609 1529 611 1531
rect 629 1529 631 1531
rect 634 1529 636 1534
rect 1452 1533 1453 1537
rect 1496 1534 1497 1538
rect 1521 1537 1523 1541
rect 1567 1538 1569 1540
rect 652 1529 654 1531
rect 1435 1529 1437 1531
rect 1451 1529 1453 1533
rect 1467 1529 1469 1531
rect 1490 1529 1492 1531
rect 1495 1529 1497 1534
rect 1522 1533 1523 1537
rect 1568 1534 1569 1538
rect 1521 1529 1523 1533
rect 1542 1529 1544 1531
rect 1562 1529 1564 1531
rect 1567 1529 1569 1534
rect 1585 1529 1587 1531
rect 702 1526 704 1529
rect 707 1526 709 1529
rect 783 1526 785 1529
rect 788 1526 790 1529
rect 873 1526 875 1529
rect 878 1526 880 1529
rect 502 1511 504 1525
rect 518 1523 520 1525
rect 518 1511 520 1513
rect 534 1511 536 1525
rect 557 1520 559 1525
rect 562 1523 564 1525
rect 588 1523 590 1525
rect 553 1516 559 1520
rect 557 1511 559 1516
rect 562 1511 564 1513
rect 588 1511 590 1513
rect 609 1511 611 1525
rect 629 1520 631 1525
rect 634 1523 636 1525
rect 625 1516 631 1520
rect 629 1511 631 1516
rect 634 1511 636 1513
rect 652 1511 654 1525
rect 1635 1526 1637 1529
rect 1640 1526 1642 1529
rect 1716 1526 1718 1529
rect 1721 1526 1723 1529
rect 1806 1526 1808 1529
rect 1811 1526 1813 1529
rect 702 1510 704 1522
rect 707 1520 709 1522
rect 707 1510 709 1512
rect 783 1510 785 1522
rect 788 1520 790 1522
rect 788 1510 790 1512
rect 873 1510 875 1522
rect 878 1520 880 1522
rect 878 1510 880 1512
rect 1435 1511 1437 1525
rect 1451 1523 1453 1525
rect 1451 1511 1453 1513
rect 1467 1511 1469 1525
rect 1490 1520 1492 1525
rect 1495 1523 1497 1525
rect 1521 1523 1523 1525
rect 1486 1516 1492 1520
rect 1490 1511 1492 1516
rect 1495 1511 1497 1513
rect 1521 1511 1523 1513
rect 1542 1511 1544 1525
rect 1562 1520 1564 1525
rect 1567 1523 1569 1525
rect 1558 1516 1564 1520
rect 1562 1511 1564 1516
rect 1567 1511 1569 1513
rect 1585 1511 1587 1525
rect 502 1501 504 1503
rect 518 1500 520 1503
rect 534 1501 536 1503
rect 557 1501 559 1503
rect 562 1500 564 1503
rect 588 1500 590 1503
rect 609 1500 611 1503
rect 629 1501 631 1503
rect 634 1500 636 1503
rect 652 1501 654 1503
rect 1635 1510 1637 1522
rect 1640 1520 1642 1522
rect 1640 1510 1642 1512
rect 1716 1510 1718 1522
rect 1721 1520 1723 1522
rect 1721 1510 1723 1512
rect 1806 1510 1808 1522
rect 1811 1520 1813 1522
rect 1811 1510 1813 1512
rect 702 1500 704 1502
rect 588 1496 589 1500
rect 707 1497 709 1502
rect 783 1500 785 1502
rect 788 1497 790 1502
rect 873 1500 875 1502
rect 878 1497 880 1502
rect 1435 1501 1437 1503
rect 518 1493 520 1496
rect 562 1493 564 1496
rect 588 1493 590 1496
rect 634 1493 636 1496
rect 1451 1500 1453 1503
rect 1467 1501 1469 1503
rect 1490 1501 1492 1503
rect 1495 1500 1497 1503
rect 1521 1500 1523 1503
rect 1542 1500 1544 1503
rect 1562 1501 1564 1503
rect 1567 1500 1569 1503
rect 1585 1501 1587 1503
rect 1635 1500 1637 1502
rect 1521 1496 1522 1500
rect 1640 1497 1642 1502
rect 1716 1500 1718 1502
rect 1721 1497 1723 1502
rect 1806 1500 1808 1502
rect 1811 1497 1813 1502
rect 1451 1493 1453 1496
rect 1495 1493 1497 1496
rect 1521 1493 1523 1496
rect 1567 1493 1569 1496
rect 518 1472 520 1475
rect 562 1472 564 1475
rect 588 1472 590 1475
rect 634 1472 636 1475
rect 702 1472 704 1476
rect 730 1478 732 1480
rect 707 1472 709 1475
rect 588 1468 589 1472
rect 502 1465 504 1467
rect 518 1465 520 1468
rect 534 1465 536 1467
rect 557 1465 559 1467
rect 562 1465 564 1468
rect 588 1465 590 1468
rect 609 1465 611 1468
rect 629 1465 631 1467
rect 634 1465 636 1468
rect 652 1465 654 1467
rect 1451 1472 1453 1475
rect 1495 1472 1497 1475
rect 1521 1472 1523 1475
rect 1567 1472 1569 1475
rect 1635 1472 1637 1476
rect 1663 1478 1665 1480
rect 1640 1472 1642 1475
rect 702 1461 704 1464
rect 707 1462 709 1464
rect 703 1457 704 1461
rect 502 1443 504 1457
rect 518 1455 520 1457
rect 518 1443 520 1445
rect 534 1443 536 1457
rect 557 1452 559 1457
rect 562 1455 564 1457
rect 588 1455 590 1457
rect 553 1448 559 1452
rect 557 1443 559 1448
rect 562 1443 564 1445
rect 588 1443 590 1445
rect 609 1443 611 1457
rect 629 1452 631 1457
rect 634 1455 636 1457
rect 625 1448 631 1452
rect 629 1443 631 1448
rect 634 1443 636 1445
rect 652 1443 654 1457
rect 702 1452 704 1457
rect 707 1452 709 1454
rect 730 1448 732 1470
rect 1521 1468 1522 1472
rect 1435 1465 1437 1467
rect 1451 1465 1453 1468
rect 1467 1465 1469 1467
rect 1490 1465 1492 1467
rect 1495 1465 1497 1468
rect 1521 1465 1523 1468
rect 1542 1465 1544 1468
rect 1562 1465 1564 1467
rect 1567 1465 1569 1468
rect 1585 1465 1587 1467
rect 1635 1461 1637 1464
rect 1640 1462 1642 1464
rect 1636 1457 1637 1461
rect 702 1446 704 1448
rect 707 1443 709 1448
rect 730 1442 732 1444
rect 1435 1443 1437 1457
rect 1451 1455 1453 1457
rect 1451 1443 1453 1445
rect 1467 1443 1469 1457
rect 1490 1452 1492 1457
rect 1495 1455 1497 1457
rect 1521 1455 1523 1457
rect 1486 1448 1492 1452
rect 1490 1443 1492 1448
rect 1495 1443 1497 1445
rect 1521 1443 1523 1445
rect 1542 1443 1544 1457
rect 1562 1452 1564 1457
rect 1567 1455 1569 1457
rect 1558 1448 1564 1452
rect 1562 1443 1564 1448
rect 1567 1443 1569 1445
rect 1585 1443 1587 1457
rect 1635 1452 1637 1457
rect 1640 1452 1642 1454
rect 1663 1448 1665 1470
rect 1635 1446 1637 1448
rect 1640 1443 1642 1448
rect 1663 1442 1665 1444
rect 502 1437 504 1439
rect 518 1435 520 1439
rect 534 1437 536 1439
rect 557 1437 559 1439
rect 519 1431 520 1435
rect 562 1434 564 1439
rect 588 1435 590 1439
rect 609 1437 611 1439
rect 629 1437 631 1439
rect 518 1428 520 1431
rect 563 1430 564 1434
rect 589 1431 590 1435
rect 634 1434 636 1439
rect 652 1437 654 1439
rect 1435 1437 1437 1439
rect 1451 1435 1453 1439
rect 1467 1437 1469 1439
rect 1490 1437 1492 1439
rect 562 1428 564 1430
rect 588 1427 590 1431
rect 635 1430 636 1434
rect 1452 1431 1453 1435
rect 1495 1434 1497 1439
rect 1521 1435 1523 1439
rect 1542 1437 1544 1439
rect 1562 1437 1564 1439
rect 634 1428 636 1430
rect 1451 1428 1453 1431
rect 1496 1430 1497 1434
rect 1522 1431 1523 1435
rect 1567 1434 1569 1439
rect 1585 1437 1587 1439
rect 1495 1428 1497 1430
rect 1521 1427 1523 1431
rect 1568 1430 1569 1434
rect 1567 1428 1569 1430
rect 25 1410 27 1412
rect 30 1410 32 1413
rect 46 1410 48 1412
rect 62 1410 64 1412
rect 67 1410 69 1413
rect 88 1410 90 1413
rect 104 1410 106 1413
rect 120 1410 122 1412
rect 125 1410 127 1413
rect 141 1410 143 1412
rect 157 1410 159 1412
rect 162 1410 164 1413
rect 178 1410 180 1412
rect 194 1410 196 1412
rect 199 1410 201 1413
rect 220 1410 222 1413
rect 236 1410 238 1413
rect 252 1410 254 1412
rect 257 1410 259 1413
rect 273 1410 275 1412
rect 289 1410 291 1412
rect 294 1410 296 1413
rect 310 1410 312 1412
rect 326 1410 328 1412
rect 331 1410 333 1413
rect 352 1410 354 1413
rect 368 1410 370 1413
rect 384 1410 386 1412
rect 389 1410 391 1413
rect 405 1410 407 1412
rect 958 1410 960 1412
rect 963 1410 965 1413
rect 979 1410 981 1412
rect 995 1410 997 1412
rect 1000 1410 1002 1413
rect 1021 1410 1023 1413
rect 1037 1410 1039 1413
rect 1053 1410 1055 1412
rect 1058 1410 1060 1413
rect 1074 1410 1076 1412
rect 1090 1410 1092 1412
rect 1095 1410 1097 1413
rect 1111 1410 1113 1412
rect 1127 1410 1129 1412
rect 1132 1410 1134 1413
rect 1153 1410 1155 1413
rect 1169 1410 1171 1413
rect 1185 1410 1187 1412
rect 1190 1410 1192 1413
rect 1206 1410 1208 1412
rect 1222 1410 1224 1412
rect 1227 1410 1229 1413
rect 1243 1410 1245 1412
rect 1259 1410 1261 1412
rect 1264 1410 1266 1413
rect 1285 1410 1287 1413
rect 1301 1410 1303 1413
rect 1317 1410 1319 1412
rect 1322 1410 1324 1413
rect 1338 1410 1340 1412
rect 518 1405 520 1408
rect 562 1406 564 1408
rect 25 1397 27 1402
rect 30 1400 32 1402
rect 25 1383 27 1393
rect 30 1383 32 1390
rect 46 1383 48 1402
rect 62 1393 64 1402
rect 67 1400 69 1402
rect 88 1400 90 1402
rect 104 1399 106 1402
rect 62 1383 64 1386
rect 67 1383 69 1385
rect 88 1383 90 1385
rect 104 1383 106 1395
rect 120 1393 122 1402
rect 125 1400 127 1402
rect 120 1383 122 1386
rect 125 1383 127 1385
rect 141 1383 143 1402
rect 157 1399 159 1402
rect 162 1400 164 1402
rect 157 1383 159 1395
rect 162 1383 164 1390
rect 178 1383 180 1402
rect 194 1393 196 1402
rect 199 1400 201 1402
rect 220 1400 222 1402
rect 236 1399 238 1402
rect 194 1383 196 1386
rect 199 1383 201 1385
rect 220 1383 222 1385
rect 236 1383 238 1395
rect 252 1393 254 1402
rect 257 1400 259 1402
rect 252 1383 254 1386
rect 257 1383 259 1385
rect 273 1383 275 1402
rect 289 1399 291 1402
rect 294 1400 296 1402
rect 289 1383 291 1395
rect 294 1383 296 1390
rect 310 1383 312 1402
rect 326 1393 328 1402
rect 331 1400 333 1402
rect 352 1400 354 1402
rect 368 1399 370 1402
rect 326 1383 328 1386
rect 331 1383 333 1385
rect 352 1383 354 1385
rect 368 1383 370 1395
rect 384 1393 386 1402
rect 389 1400 391 1402
rect 405 1394 407 1402
rect 519 1401 520 1405
rect 563 1402 564 1406
rect 588 1405 590 1409
rect 634 1406 636 1408
rect 502 1397 504 1399
rect 518 1397 520 1401
rect 534 1397 536 1399
rect 557 1397 559 1399
rect 562 1397 564 1402
rect 589 1401 590 1405
rect 635 1402 636 1406
rect 779 1405 781 1408
rect 823 1406 825 1408
rect 588 1397 590 1401
rect 609 1397 611 1399
rect 629 1397 631 1399
rect 634 1397 636 1402
rect 780 1401 781 1405
rect 824 1402 825 1406
rect 849 1405 851 1409
rect 895 1406 897 1408
rect 652 1397 654 1399
rect 736 1397 738 1400
rect 754 1397 756 1400
rect 779 1397 781 1401
rect 795 1397 797 1399
rect 818 1397 820 1399
rect 823 1397 825 1402
rect 850 1401 851 1405
rect 896 1402 897 1406
rect 1451 1405 1453 1408
rect 1495 1406 1497 1408
rect 849 1397 851 1401
rect 870 1397 872 1399
rect 890 1397 892 1399
rect 895 1397 897 1402
rect 913 1397 915 1399
rect 958 1397 960 1402
rect 963 1400 965 1402
rect 384 1383 386 1386
rect 389 1383 391 1385
rect 405 1383 407 1390
rect 502 1379 504 1393
rect 518 1391 520 1393
rect 518 1379 520 1381
rect 534 1379 536 1393
rect 557 1388 559 1393
rect 562 1391 564 1393
rect 588 1391 590 1393
rect 553 1384 559 1388
rect 557 1379 559 1384
rect 562 1379 564 1381
rect 588 1379 590 1381
rect 609 1379 611 1393
rect 629 1388 631 1393
rect 634 1391 636 1393
rect 625 1384 631 1388
rect 629 1379 631 1384
rect 634 1379 636 1381
rect 652 1379 654 1393
rect 702 1390 704 1393
rect 707 1390 709 1393
rect 736 1388 738 1393
rect 25 1377 27 1379
rect 30 1376 32 1379
rect 46 1377 48 1379
rect 62 1377 64 1379
rect 67 1374 69 1379
rect 88 1374 90 1379
rect 104 1377 106 1379
rect 120 1377 122 1379
rect 125 1374 127 1379
rect 141 1377 143 1379
rect 157 1377 159 1379
rect 162 1376 164 1379
rect 178 1377 180 1379
rect 194 1377 196 1379
rect 199 1374 201 1379
rect 220 1374 222 1379
rect 236 1377 238 1379
rect 252 1377 254 1379
rect 257 1374 259 1379
rect 273 1377 275 1379
rect 289 1377 291 1379
rect 294 1376 296 1379
rect 310 1377 312 1379
rect 326 1377 328 1379
rect 331 1374 333 1379
rect 352 1374 354 1379
rect 368 1377 370 1379
rect 384 1377 386 1379
rect 389 1374 391 1379
rect 405 1377 407 1379
rect 702 1374 704 1386
rect 707 1384 709 1386
rect 736 1379 738 1384
rect 754 1379 756 1393
rect 779 1391 781 1393
rect 779 1379 781 1381
rect 795 1379 797 1393
rect 818 1388 820 1393
rect 823 1391 825 1393
rect 849 1391 851 1393
rect 814 1384 820 1388
rect 818 1379 820 1384
rect 823 1379 825 1381
rect 849 1379 851 1381
rect 870 1379 872 1393
rect 890 1388 892 1393
rect 895 1391 897 1393
rect 886 1384 892 1388
rect 890 1379 892 1384
rect 895 1379 897 1381
rect 913 1379 915 1393
rect 958 1383 960 1393
rect 963 1383 965 1390
rect 979 1383 981 1402
rect 995 1393 997 1402
rect 1000 1400 1002 1402
rect 1021 1400 1023 1402
rect 1037 1399 1039 1402
rect 995 1383 997 1386
rect 1000 1383 1002 1385
rect 1021 1383 1023 1385
rect 1037 1383 1039 1395
rect 1053 1393 1055 1402
rect 1058 1400 1060 1402
rect 1053 1383 1055 1386
rect 1058 1383 1060 1385
rect 1074 1383 1076 1402
rect 1090 1399 1092 1402
rect 1095 1400 1097 1402
rect 1090 1383 1092 1395
rect 1095 1383 1097 1390
rect 1111 1383 1113 1402
rect 1127 1393 1129 1402
rect 1132 1400 1134 1402
rect 1153 1400 1155 1402
rect 1169 1399 1171 1402
rect 1127 1383 1129 1386
rect 1132 1383 1134 1385
rect 1153 1383 1155 1385
rect 1169 1383 1171 1395
rect 1185 1393 1187 1402
rect 1190 1400 1192 1402
rect 1185 1383 1187 1386
rect 1190 1383 1192 1385
rect 1206 1383 1208 1402
rect 1222 1399 1224 1402
rect 1227 1400 1229 1402
rect 1222 1383 1224 1395
rect 1227 1383 1229 1390
rect 1243 1383 1245 1402
rect 1259 1393 1261 1402
rect 1264 1400 1266 1402
rect 1285 1400 1287 1402
rect 1301 1399 1303 1402
rect 1259 1383 1261 1386
rect 1264 1383 1266 1385
rect 1285 1383 1287 1385
rect 1301 1383 1303 1395
rect 1317 1393 1319 1402
rect 1322 1400 1324 1402
rect 1338 1394 1340 1402
rect 1452 1401 1453 1405
rect 1496 1402 1497 1406
rect 1521 1405 1523 1409
rect 1567 1406 1569 1408
rect 1435 1397 1437 1399
rect 1451 1397 1453 1401
rect 1467 1397 1469 1399
rect 1490 1397 1492 1399
rect 1495 1397 1497 1402
rect 1522 1401 1523 1405
rect 1568 1402 1569 1406
rect 1712 1405 1714 1408
rect 1756 1406 1758 1408
rect 1521 1397 1523 1401
rect 1542 1397 1544 1399
rect 1562 1397 1564 1399
rect 1567 1397 1569 1402
rect 1713 1401 1714 1405
rect 1757 1402 1758 1406
rect 1782 1405 1784 1409
rect 1828 1406 1830 1408
rect 1585 1397 1587 1399
rect 1669 1397 1671 1400
rect 1687 1397 1689 1400
rect 1712 1397 1714 1401
rect 1728 1397 1730 1399
rect 1751 1397 1753 1399
rect 1756 1397 1758 1402
rect 1783 1401 1784 1405
rect 1829 1402 1830 1406
rect 1782 1397 1784 1401
rect 1803 1397 1805 1399
rect 1823 1397 1825 1399
rect 1828 1397 1830 1402
rect 1846 1397 1848 1399
rect 1317 1383 1319 1386
rect 1322 1383 1324 1385
rect 1338 1383 1340 1390
rect 1435 1379 1437 1393
rect 1451 1391 1453 1393
rect 1451 1379 1453 1381
rect 1467 1379 1469 1393
rect 1490 1388 1492 1393
rect 1495 1391 1497 1393
rect 1521 1391 1523 1393
rect 1486 1384 1492 1388
rect 1490 1379 1492 1384
rect 1495 1379 1497 1381
rect 1521 1379 1523 1381
rect 1542 1379 1544 1393
rect 1562 1388 1564 1393
rect 1567 1391 1569 1393
rect 1558 1384 1564 1388
rect 1562 1379 1564 1384
rect 1567 1379 1569 1381
rect 1585 1379 1587 1393
rect 1635 1390 1637 1393
rect 1640 1390 1642 1393
rect 1669 1388 1671 1393
rect 707 1374 709 1376
rect 502 1369 504 1371
rect 518 1368 520 1371
rect 534 1369 536 1371
rect 557 1369 559 1371
rect 562 1368 564 1371
rect 588 1368 590 1371
rect 609 1368 611 1371
rect 629 1369 631 1371
rect 634 1368 636 1371
rect 652 1369 654 1371
rect 588 1364 589 1368
rect 958 1377 960 1379
rect 963 1376 965 1379
rect 979 1377 981 1379
rect 995 1377 997 1379
rect 1000 1374 1002 1379
rect 1021 1374 1023 1379
rect 1037 1377 1039 1379
rect 1053 1377 1055 1379
rect 1058 1374 1060 1379
rect 1074 1377 1076 1379
rect 1090 1377 1092 1379
rect 736 1368 738 1371
rect 754 1368 756 1371
rect 779 1368 781 1371
rect 795 1369 797 1371
rect 818 1369 820 1371
rect 823 1368 825 1371
rect 849 1368 851 1371
rect 870 1368 872 1371
rect 890 1369 892 1371
rect 895 1368 897 1371
rect 913 1369 915 1371
rect 1095 1376 1097 1379
rect 1111 1377 1113 1379
rect 1127 1377 1129 1379
rect 1132 1374 1134 1379
rect 1153 1374 1155 1379
rect 1169 1377 1171 1379
rect 1185 1377 1187 1379
rect 1190 1374 1192 1379
rect 1206 1377 1208 1379
rect 1222 1377 1224 1379
rect 1227 1376 1229 1379
rect 1243 1377 1245 1379
rect 1259 1377 1261 1379
rect 1264 1374 1266 1379
rect 1285 1374 1287 1379
rect 1301 1377 1303 1379
rect 1317 1377 1319 1379
rect 1322 1374 1324 1379
rect 1338 1377 1340 1379
rect 1635 1374 1637 1386
rect 1640 1384 1642 1386
rect 1669 1379 1671 1384
rect 1687 1379 1689 1393
rect 1712 1391 1714 1393
rect 1712 1379 1714 1381
rect 1728 1379 1730 1393
rect 1751 1388 1753 1393
rect 1756 1391 1758 1393
rect 1782 1391 1784 1393
rect 1747 1384 1753 1388
rect 1751 1379 1753 1384
rect 1756 1379 1758 1381
rect 1782 1379 1784 1381
rect 1803 1379 1805 1393
rect 1823 1388 1825 1393
rect 1828 1391 1830 1393
rect 1819 1384 1825 1388
rect 1823 1379 1825 1384
rect 1828 1379 1830 1381
rect 1846 1379 1848 1393
rect 1640 1374 1642 1376
rect 1435 1369 1437 1371
rect 1451 1368 1453 1371
rect 1467 1369 1469 1371
rect 1490 1369 1492 1371
rect 1495 1368 1497 1371
rect 1521 1368 1523 1371
rect 1542 1368 1544 1371
rect 1562 1369 1564 1371
rect 1567 1368 1569 1371
rect 1585 1369 1587 1371
rect 702 1364 704 1366
rect 518 1361 520 1364
rect 562 1361 564 1364
rect 588 1361 590 1364
rect 634 1361 636 1364
rect 707 1361 709 1366
rect 849 1364 850 1368
rect 779 1361 781 1364
rect 823 1361 825 1364
rect 849 1361 851 1364
rect 895 1361 897 1364
rect 1521 1364 1522 1368
rect 1669 1368 1671 1371
rect 1687 1368 1689 1371
rect 1712 1368 1714 1371
rect 1728 1369 1730 1371
rect 1751 1369 1753 1371
rect 1756 1368 1758 1371
rect 1782 1368 1784 1371
rect 1803 1368 1805 1371
rect 1823 1369 1825 1371
rect 1828 1368 1830 1371
rect 1846 1369 1848 1371
rect 1635 1364 1637 1366
rect 1451 1361 1453 1364
rect 1495 1361 1497 1364
rect 1521 1361 1523 1364
rect 1567 1361 1569 1364
rect 1640 1361 1642 1366
rect 1782 1364 1783 1368
rect 1712 1361 1714 1364
rect 1756 1361 1758 1364
rect 1782 1361 1784 1364
rect 1828 1361 1830 1364
rect 140 1339 142 1342
rect 164 1339 166 1342
rect 1073 1339 1075 1342
rect 1097 1339 1099 1342
rect 922 1337 925 1339
rect 929 1337 932 1339
rect 140 1333 142 1335
rect 164 1333 166 1335
rect 1855 1337 1858 1339
rect 1862 1337 1865 1339
rect 1073 1333 1075 1335
rect 1097 1333 1099 1335
rect 160 1328 162 1330
rect 1093 1328 1095 1330
rect 160 1321 162 1324
rect 1093 1321 1095 1324
rect 149 1310 151 1312
rect 155 1310 174 1312
rect 1082 1310 1084 1312
rect 1088 1310 1107 1312
rect 140 1305 142 1307
rect 164 1305 166 1307
rect 1073 1305 1075 1307
rect 1097 1305 1099 1307
rect 140 1298 142 1301
rect 164 1298 166 1301
rect 796 1300 798 1302
rect 801 1300 803 1303
rect 817 1300 819 1302
rect 833 1300 835 1302
rect 838 1300 840 1303
rect 859 1300 861 1303
rect 875 1300 877 1303
rect 891 1300 893 1302
rect 896 1300 898 1303
rect 912 1300 914 1302
rect 1073 1298 1075 1301
rect 1097 1298 1099 1301
rect 1729 1300 1731 1302
rect 1734 1300 1736 1303
rect 1750 1300 1752 1302
rect 1766 1300 1768 1302
rect 1771 1300 1773 1303
rect 1792 1300 1794 1303
rect 1808 1300 1810 1303
rect 1824 1300 1826 1302
rect 1829 1300 1831 1303
rect 1845 1300 1847 1302
rect 796 1287 798 1292
rect 801 1290 803 1292
rect 796 1273 798 1283
rect 801 1273 803 1280
rect 817 1273 819 1292
rect 833 1283 835 1292
rect 838 1290 840 1292
rect 859 1290 861 1292
rect 875 1289 877 1292
rect 833 1273 835 1276
rect 838 1273 840 1275
rect 859 1273 861 1275
rect 875 1273 877 1285
rect 891 1283 893 1292
rect 896 1290 898 1292
rect 891 1273 893 1276
rect 896 1273 898 1275
rect 912 1273 914 1292
rect 1729 1287 1731 1292
rect 1734 1290 1736 1292
rect 1729 1273 1731 1283
rect 1734 1273 1736 1280
rect 1750 1273 1752 1292
rect 1766 1283 1768 1292
rect 1771 1290 1773 1292
rect 1792 1290 1794 1292
rect 1808 1289 1810 1292
rect 1766 1273 1768 1276
rect 1771 1273 1773 1275
rect 1792 1273 1794 1275
rect 1808 1273 1810 1285
rect 1824 1283 1826 1292
rect 1829 1290 1831 1292
rect 1824 1273 1826 1276
rect 1829 1273 1831 1275
rect 1845 1273 1847 1292
rect 25 1270 27 1272
rect 30 1270 32 1273
rect 46 1270 48 1272
rect 62 1270 64 1272
rect 67 1270 69 1273
rect 88 1270 90 1273
rect 104 1270 106 1273
rect 120 1270 122 1272
rect 125 1270 127 1273
rect 141 1270 143 1272
rect 157 1270 159 1272
rect 162 1270 164 1273
rect 178 1270 180 1272
rect 194 1270 196 1272
rect 199 1270 201 1273
rect 220 1270 222 1273
rect 236 1270 238 1273
rect 252 1270 254 1272
rect 257 1270 259 1273
rect 273 1270 275 1272
rect 289 1270 291 1272
rect 294 1270 296 1273
rect 310 1270 312 1272
rect 326 1270 328 1272
rect 331 1270 333 1273
rect 352 1270 354 1273
rect 368 1270 370 1273
rect 384 1270 386 1272
rect 389 1270 391 1273
rect 405 1270 407 1272
rect 958 1270 960 1272
rect 963 1270 965 1273
rect 979 1270 981 1272
rect 995 1270 997 1272
rect 1000 1270 1002 1273
rect 1021 1270 1023 1273
rect 1037 1270 1039 1273
rect 1053 1270 1055 1272
rect 1058 1270 1060 1273
rect 1074 1270 1076 1272
rect 1090 1270 1092 1272
rect 1095 1270 1097 1273
rect 1111 1270 1113 1272
rect 1127 1270 1129 1272
rect 1132 1270 1134 1273
rect 1153 1270 1155 1273
rect 1169 1270 1171 1273
rect 1185 1270 1187 1272
rect 1190 1270 1192 1273
rect 1206 1270 1208 1272
rect 1222 1270 1224 1272
rect 1227 1270 1229 1273
rect 1243 1270 1245 1272
rect 1259 1270 1261 1272
rect 1264 1270 1266 1273
rect 1285 1270 1287 1273
rect 1301 1270 1303 1273
rect 1317 1270 1319 1272
rect 1322 1270 1324 1273
rect 1338 1270 1340 1272
rect 796 1267 798 1269
rect 801 1266 803 1269
rect 817 1267 819 1269
rect 833 1267 835 1269
rect 838 1264 840 1269
rect 859 1264 861 1269
rect 875 1267 877 1269
rect 891 1267 893 1269
rect 896 1264 898 1269
rect 912 1267 914 1269
rect 25 1257 27 1262
rect 30 1260 32 1262
rect 25 1243 27 1253
rect 30 1243 32 1250
rect 46 1243 48 1262
rect 62 1253 64 1262
rect 67 1260 69 1262
rect 88 1260 90 1262
rect 104 1259 106 1262
rect 62 1243 64 1246
rect 67 1243 69 1245
rect 88 1243 90 1245
rect 104 1243 106 1255
rect 120 1253 122 1262
rect 125 1260 127 1262
rect 120 1243 122 1246
rect 125 1243 127 1245
rect 141 1243 143 1262
rect 157 1259 159 1262
rect 162 1260 164 1262
rect 157 1243 159 1255
rect 162 1243 164 1250
rect 178 1243 180 1262
rect 194 1253 196 1262
rect 199 1260 201 1262
rect 220 1260 222 1262
rect 236 1259 238 1262
rect 194 1243 196 1246
rect 199 1243 201 1245
rect 220 1243 222 1245
rect 236 1243 238 1255
rect 252 1253 254 1262
rect 257 1260 259 1262
rect 252 1243 254 1246
rect 257 1243 259 1245
rect 273 1243 275 1262
rect 289 1259 291 1262
rect 294 1260 296 1262
rect 289 1243 291 1255
rect 294 1243 296 1250
rect 310 1243 312 1262
rect 326 1253 328 1262
rect 331 1260 333 1262
rect 352 1260 354 1262
rect 368 1259 370 1262
rect 326 1243 328 1246
rect 331 1243 333 1245
rect 352 1243 354 1245
rect 368 1243 370 1255
rect 384 1253 386 1262
rect 389 1260 391 1262
rect 405 1254 407 1262
rect 1729 1267 1731 1269
rect 1734 1266 1736 1269
rect 1750 1267 1752 1269
rect 1766 1267 1768 1269
rect 1771 1264 1773 1269
rect 1792 1264 1794 1269
rect 1808 1267 1810 1269
rect 1824 1267 1826 1269
rect 1829 1264 1831 1269
rect 1845 1267 1847 1269
rect 958 1257 960 1262
rect 963 1260 965 1262
rect 384 1243 386 1246
rect 389 1243 391 1245
rect 405 1243 407 1250
rect 958 1243 960 1253
rect 963 1243 965 1250
rect 979 1243 981 1262
rect 995 1253 997 1262
rect 1000 1260 1002 1262
rect 1021 1260 1023 1262
rect 1037 1259 1039 1262
rect 995 1243 997 1246
rect 1000 1243 1002 1245
rect 1021 1243 1023 1245
rect 1037 1243 1039 1255
rect 1053 1253 1055 1262
rect 1058 1260 1060 1262
rect 1053 1243 1055 1246
rect 1058 1243 1060 1245
rect 1074 1243 1076 1262
rect 1090 1259 1092 1262
rect 1095 1260 1097 1262
rect 1090 1243 1092 1255
rect 1095 1243 1097 1250
rect 1111 1243 1113 1262
rect 1127 1253 1129 1262
rect 1132 1260 1134 1262
rect 1153 1260 1155 1262
rect 1169 1259 1171 1262
rect 1127 1243 1129 1246
rect 1132 1243 1134 1245
rect 1153 1243 1155 1245
rect 1169 1243 1171 1255
rect 1185 1253 1187 1262
rect 1190 1260 1192 1262
rect 1185 1243 1187 1246
rect 1190 1243 1192 1245
rect 1206 1243 1208 1262
rect 1222 1259 1224 1262
rect 1227 1260 1229 1262
rect 1222 1243 1224 1255
rect 1227 1243 1229 1250
rect 1243 1243 1245 1262
rect 1259 1253 1261 1262
rect 1264 1260 1266 1262
rect 1285 1260 1287 1262
rect 1301 1259 1303 1262
rect 1259 1243 1261 1246
rect 1264 1243 1266 1245
rect 1285 1243 1287 1245
rect 1301 1243 1303 1255
rect 1317 1253 1319 1262
rect 1322 1260 1324 1262
rect 1338 1254 1340 1262
rect 1317 1243 1319 1246
rect 1322 1243 1324 1245
rect 1338 1243 1340 1250
rect 25 1237 27 1239
rect 30 1236 32 1239
rect 46 1237 48 1239
rect 62 1237 64 1239
rect 67 1234 69 1239
rect 88 1234 90 1239
rect 104 1237 106 1239
rect 120 1237 122 1239
rect 125 1234 127 1239
rect 141 1237 143 1239
rect 157 1237 159 1239
rect 162 1236 164 1239
rect 178 1237 180 1239
rect 194 1237 196 1239
rect 199 1234 201 1239
rect 220 1234 222 1239
rect 236 1237 238 1239
rect 252 1237 254 1239
rect 257 1234 259 1239
rect 273 1237 275 1239
rect 289 1237 291 1239
rect 294 1236 296 1239
rect 310 1237 312 1239
rect 326 1237 328 1239
rect 331 1234 333 1239
rect 352 1234 354 1239
rect 368 1237 370 1239
rect 384 1237 386 1239
rect 389 1234 391 1239
rect 405 1237 407 1239
rect 958 1237 960 1239
rect 963 1236 965 1239
rect 979 1237 981 1239
rect 995 1237 997 1239
rect 1000 1234 1002 1239
rect 1021 1234 1023 1239
rect 1037 1237 1039 1239
rect 1053 1237 1055 1239
rect 1058 1234 1060 1239
rect 1074 1237 1076 1239
rect 1090 1237 1092 1239
rect 1095 1236 1097 1239
rect 1111 1237 1113 1239
rect 1127 1237 1129 1239
rect 1132 1234 1134 1239
rect 1153 1234 1155 1239
rect 1169 1237 1171 1239
rect 1185 1237 1187 1239
rect 1190 1234 1192 1239
rect 1206 1237 1208 1239
rect 1222 1237 1224 1239
rect 1227 1236 1229 1239
rect 1243 1237 1245 1239
rect 1259 1237 1261 1239
rect 1264 1234 1266 1239
rect 1285 1234 1287 1239
rect 1301 1237 1303 1239
rect 1317 1237 1319 1239
rect 1322 1234 1324 1239
rect 1338 1237 1340 1239
rect 796 1214 798 1216
rect 801 1214 803 1217
rect 817 1214 819 1216
rect 833 1214 835 1216
rect 838 1214 840 1217
rect 859 1214 861 1217
rect 875 1214 877 1217
rect 891 1214 893 1216
rect 896 1214 898 1217
rect 912 1214 914 1216
rect 1729 1214 1731 1216
rect 1734 1214 1736 1217
rect 1750 1214 1752 1216
rect 1766 1214 1768 1216
rect 1771 1214 1773 1217
rect 1792 1214 1794 1217
rect 1808 1214 1810 1217
rect 1824 1214 1826 1216
rect 1829 1214 1831 1217
rect 1845 1214 1847 1216
rect 796 1201 798 1206
rect 801 1204 803 1206
rect 796 1187 798 1197
rect 801 1187 803 1194
rect 817 1187 819 1206
rect 833 1197 835 1206
rect 838 1204 840 1206
rect 859 1204 861 1206
rect 875 1203 877 1206
rect 833 1187 835 1190
rect 838 1187 840 1189
rect 859 1187 861 1189
rect 875 1187 877 1199
rect 891 1197 893 1206
rect 896 1204 898 1206
rect 891 1187 893 1190
rect 896 1187 898 1189
rect 912 1187 914 1206
rect 1729 1201 1731 1206
rect 1734 1204 1736 1206
rect 934 1193 937 1195
rect 941 1193 944 1195
rect 1729 1187 1731 1197
rect 1734 1187 1736 1194
rect 1750 1187 1752 1206
rect 1766 1197 1768 1206
rect 1771 1204 1773 1206
rect 1792 1204 1794 1206
rect 1808 1203 1810 1206
rect 1766 1187 1768 1190
rect 1771 1187 1773 1189
rect 1792 1187 1794 1189
rect 1808 1187 1810 1199
rect 1824 1197 1826 1206
rect 1829 1204 1831 1206
rect 1824 1187 1826 1190
rect 1829 1187 1831 1189
rect 1845 1187 1847 1206
rect 1867 1193 1870 1195
rect 1874 1193 1877 1195
rect 25 1184 27 1186
rect 30 1184 32 1187
rect 46 1184 48 1186
rect 62 1184 64 1186
rect 67 1184 69 1187
rect 88 1184 90 1187
rect 104 1184 106 1187
rect 120 1184 122 1186
rect 125 1184 127 1187
rect 141 1184 143 1186
rect 157 1184 159 1186
rect 162 1184 164 1187
rect 178 1184 180 1186
rect 194 1184 196 1186
rect 199 1184 201 1187
rect 220 1184 222 1187
rect 236 1184 238 1187
rect 252 1184 254 1186
rect 257 1184 259 1187
rect 273 1184 275 1186
rect 289 1184 291 1186
rect 294 1184 296 1187
rect 310 1184 312 1186
rect 326 1184 328 1186
rect 331 1184 333 1187
rect 352 1184 354 1187
rect 368 1184 370 1187
rect 384 1184 386 1186
rect 389 1184 391 1187
rect 405 1184 407 1186
rect 958 1184 960 1186
rect 963 1184 965 1187
rect 979 1184 981 1186
rect 995 1184 997 1186
rect 1000 1184 1002 1187
rect 1021 1184 1023 1187
rect 1037 1184 1039 1187
rect 1053 1184 1055 1186
rect 1058 1184 1060 1187
rect 1074 1184 1076 1186
rect 1090 1184 1092 1186
rect 1095 1184 1097 1187
rect 1111 1184 1113 1186
rect 1127 1184 1129 1186
rect 1132 1184 1134 1187
rect 1153 1184 1155 1187
rect 1169 1184 1171 1187
rect 1185 1184 1187 1186
rect 1190 1184 1192 1187
rect 1206 1184 1208 1186
rect 1222 1184 1224 1186
rect 1227 1184 1229 1187
rect 1243 1184 1245 1186
rect 1259 1184 1261 1186
rect 1264 1184 1266 1187
rect 1285 1184 1287 1187
rect 1301 1184 1303 1187
rect 1317 1184 1319 1186
rect 1322 1184 1324 1187
rect 1338 1184 1340 1186
rect 796 1181 798 1183
rect 801 1180 803 1183
rect 817 1181 819 1183
rect 833 1181 835 1183
rect 838 1178 840 1183
rect 859 1178 861 1183
rect 875 1181 877 1183
rect 891 1181 893 1183
rect 896 1178 898 1183
rect 912 1181 914 1183
rect 25 1171 27 1176
rect 30 1174 32 1176
rect 25 1157 27 1167
rect 30 1157 32 1164
rect 46 1157 48 1176
rect 62 1167 64 1176
rect 67 1174 69 1176
rect 88 1174 90 1176
rect 104 1173 106 1176
rect 62 1157 64 1160
rect 67 1157 69 1159
rect 88 1157 90 1159
rect 104 1157 106 1169
rect 120 1167 122 1176
rect 125 1174 127 1176
rect 120 1157 122 1160
rect 125 1157 127 1159
rect 141 1157 143 1176
rect 157 1173 159 1176
rect 162 1174 164 1176
rect 157 1157 159 1169
rect 162 1157 164 1164
rect 178 1157 180 1176
rect 194 1167 196 1176
rect 199 1174 201 1176
rect 220 1174 222 1176
rect 236 1173 238 1176
rect 194 1157 196 1160
rect 199 1157 201 1159
rect 220 1157 222 1159
rect 236 1157 238 1169
rect 252 1167 254 1176
rect 257 1174 259 1176
rect 252 1157 254 1160
rect 257 1157 259 1159
rect 273 1157 275 1176
rect 289 1173 291 1176
rect 294 1174 296 1176
rect 289 1157 291 1169
rect 294 1157 296 1164
rect 310 1157 312 1176
rect 326 1167 328 1176
rect 331 1174 333 1176
rect 352 1174 354 1176
rect 368 1173 370 1176
rect 326 1157 328 1160
rect 331 1157 333 1159
rect 352 1157 354 1159
rect 368 1157 370 1169
rect 384 1167 386 1176
rect 389 1174 391 1176
rect 405 1168 407 1176
rect 1729 1181 1731 1183
rect 1734 1180 1736 1183
rect 1750 1181 1752 1183
rect 1766 1181 1768 1183
rect 1771 1178 1773 1183
rect 1792 1178 1794 1183
rect 1808 1181 1810 1183
rect 1824 1181 1826 1183
rect 1829 1178 1831 1183
rect 1845 1181 1847 1183
rect 958 1171 960 1176
rect 963 1174 965 1176
rect 384 1157 386 1160
rect 389 1157 391 1159
rect 405 1157 407 1164
rect 958 1157 960 1167
rect 963 1157 965 1164
rect 979 1157 981 1176
rect 995 1167 997 1176
rect 1000 1174 1002 1176
rect 1021 1174 1023 1176
rect 1037 1173 1039 1176
rect 995 1157 997 1160
rect 1000 1157 1002 1159
rect 1021 1157 1023 1159
rect 1037 1157 1039 1169
rect 1053 1167 1055 1176
rect 1058 1174 1060 1176
rect 1053 1157 1055 1160
rect 1058 1157 1060 1159
rect 1074 1157 1076 1176
rect 1090 1173 1092 1176
rect 1095 1174 1097 1176
rect 1090 1157 1092 1169
rect 1095 1157 1097 1164
rect 1111 1157 1113 1176
rect 1127 1167 1129 1176
rect 1132 1174 1134 1176
rect 1153 1174 1155 1176
rect 1169 1173 1171 1176
rect 1127 1157 1129 1160
rect 1132 1157 1134 1159
rect 1153 1157 1155 1159
rect 1169 1157 1171 1169
rect 1185 1167 1187 1176
rect 1190 1174 1192 1176
rect 1185 1157 1187 1160
rect 1190 1157 1192 1159
rect 1206 1157 1208 1176
rect 1222 1173 1224 1176
rect 1227 1174 1229 1176
rect 1222 1157 1224 1169
rect 1227 1157 1229 1164
rect 1243 1157 1245 1176
rect 1259 1167 1261 1176
rect 1264 1174 1266 1176
rect 1285 1174 1287 1176
rect 1301 1173 1303 1176
rect 1259 1157 1261 1160
rect 1264 1157 1266 1159
rect 1285 1157 1287 1159
rect 1301 1157 1303 1169
rect 1317 1167 1319 1176
rect 1322 1174 1324 1176
rect 1338 1168 1340 1176
rect 1317 1157 1319 1160
rect 1322 1157 1324 1159
rect 1338 1157 1340 1164
rect 25 1151 27 1153
rect 30 1150 32 1153
rect 46 1151 48 1153
rect 62 1151 64 1153
rect 67 1148 69 1153
rect 88 1148 90 1153
rect 104 1151 106 1153
rect 120 1151 122 1153
rect 125 1148 127 1153
rect 141 1151 143 1153
rect 157 1151 159 1153
rect 162 1150 164 1153
rect 178 1151 180 1153
rect 194 1151 196 1153
rect 199 1148 201 1153
rect 220 1148 222 1153
rect 236 1151 238 1153
rect 252 1151 254 1153
rect 257 1148 259 1153
rect 273 1151 275 1153
rect 289 1151 291 1153
rect 294 1150 296 1153
rect 310 1151 312 1153
rect 326 1151 328 1153
rect 331 1148 333 1153
rect 352 1148 354 1153
rect 368 1151 370 1153
rect 384 1151 386 1153
rect 389 1148 391 1153
rect 405 1151 407 1153
rect 958 1151 960 1153
rect 963 1150 965 1153
rect 979 1151 981 1153
rect 995 1151 997 1153
rect 1000 1148 1002 1153
rect 1021 1148 1023 1153
rect 1037 1151 1039 1153
rect 1053 1151 1055 1153
rect 1058 1148 1060 1153
rect 1074 1151 1076 1153
rect 1090 1151 1092 1153
rect 1095 1150 1097 1153
rect 1111 1151 1113 1153
rect 1127 1151 1129 1153
rect 1132 1148 1134 1153
rect 1153 1148 1155 1153
rect 1169 1151 1171 1153
rect 1185 1151 1187 1153
rect 1190 1148 1192 1153
rect 1206 1151 1208 1153
rect 1222 1151 1224 1153
rect 1227 1150 1229 1153
rect 1243 1151 1245 1153
rect 1259 1151 1261 1153
rect 1264 1148 1266 1153
rect 1285 1148 1287 1153
rect 1301 1151 1303 1153
rect 1317 1151 1319 1153
rect 1322 1148 1324 1153
rect 1338 1151 1340 1153
rect 257 1113 259 1116
rect 281 1113 283 1116
rect 1190 1113 1192 1116
rect 1214 1113 1216 1116
rect 257 1107 259 1109
rect 281 1107 283 1109
rect 1190 1107 1192 1109
rect 1214 1107 1216 1109
rect 277 1102 279 1104
rect 1210 1102 1212 1104
rect 277 1095 279 1098
rect 1210 1095 1212 1098
rect 266 1084 268 1086
rect 272 1084 291 1086
rect 1199 1084 1201 1086
rect 1205 1084 1224 1086
rect 257 1079 259 1081
rect 281 1079 283 1081
rect 1190 1079 1192 1081
rect 1214 1079 1216 1081
rect 257 1072 259 1075
rect 281 1072 283 1075
rect 1190 1072 1192 1075
rect 1214 1072 1216 1075
rect 25 1044 27 1046
rect 30 1044 32 1047
rect 46 1044 48 1046
rect 62 1044 64 1046
rect 67 1044 69 1047
rect 88 1044 90 1047
rect 104 1044 106 1047
rect 120 1044 122 1046
rect 125 1044 127 1047
rect 141 1044 143 1046
rect 157 1044 159 1046
rect 162 1044 164 1047
rect 178 1044 180 1046
rect 194 1044 196 1046
rect 199 1044 201 1047
rect 220 1044 222 1047
rect 236 1044 238 1047
rect 252 1044 254 1046
rect 257 1044 259 1047
rect 273 1044 275 1046
rect 289 1044 291 1046
rect 294 1044 296 1047
rect 310 1044 312 1046
rect 326 1044 328 1046
rect 331 1044 333 1047
rect 352 1044 354 1047
rect 368 1044 370 1047
rect 384 1044 386 1046
rect 389 1044 391 1047
rect 405 1044 407 1046
rect 958 1044 960 1046
rect 963 1044 965 1047
rect 979 1044 981 1046
rect 995 1044 997 1046
rect 1000 1044 1002 1047
rect 1021 1044 1023 1047
rect 1037 1044 1039 1047
rect 1053 1044 1055 1046
rect 1058 1044 1060 1047
rect 1074 1044 1076 1046
rect 1090 1044 1092 1046
rect 1095 1044 1097 1047
rect 1111 1044 1113 1046
rect 1127 1044 1129 1046
rect 1132 1044 1134 1047
rect 1153 1044 1155 1047
rect 1169 1044 1171 1047
rect 1185 1044 1187 1046
rect 1190 1044 1192 1047
rect 1206 1044 1208 1046
rect 1222 1044 1224 1046
rect 1227 1044 1229 1047
rect 1243 1044 1245 1046
rect 1259 1044 1261 1046
rect 1264 1044 1266 1047
rect 1285 1044 1287 1047
rect 1301 1044 1303 1047
rect 1317 1044 1319 1046
rect 1322 1044 1324 1047
rect 1338 1044 1340 1046
rect 25 1031 27 1036
rect 30 1034 32 1036
rect 25 1017 27 1027
rect 30 1017 32 1024
rect 46 1017 48 1036
rect 62 1027 64 1036
rect 67 1034 69 1036
rect 88 1034 90 1036
rect 104 1033 106 1036
rect 62 1017 64 1020
rect 67 1017 69 1019
rect 88 1017 90 1019
rect 104 1017 106 1029
rect 120 1027 122 1036
rect 125 1034 127 1036
rect 120 1017 122 1020
rect 125 1017 127 1019
rect 141 1017 143 1036
rect 157 1033 159 1036
rect 162 1034 164 1036
rect 157 1017 159 1029
rect 162 1017 164 1024
rect 178 1017 180 1036
rect 194 1027 196 1036
rect 199 1034 201 1036
rect 220 1034 222 1036
rect 236 1033 238 1036
rect 194 1017 196 1020
rect 199 1017 201 1019
rect 220 1017 222 1019
rect 236 1017 238 1029
rect 252 1027 254 1036
rect 257 1034 259 1036
rect 252 1017 254 1020
rect 257 1017 259 1019
rect 273 1017 275 1036
rect 289 1033 291 1036
rect 294 1034 296 1036
rect 289 1017 291 1029
rect 294 1017 296 1024
rect 310 1017 312 1036
rect 326 1027 328 1036
rect 331 1034 333 1036
rect 352 1034 354 1036
rect 368 1033 370 1036
rect 326 1017 328 1020
rect 331 1017 333 1019
rect 352 1017 354 1019
rect 368 1017 370 1029
rect 384 1027 386 1036
rect 389 1034 391 1036
rect 405 1028 407 1036
rect 958 1031 960 1036
rect 963 1034 965 1036
rect 384 1017 386 1020
rect 389 1017 391 1019
rect 405 1017 407 1024
rect 958 1017 960 1027
rect 963 1017 965 1024
rect 979 1017 981 1036
rect 995 1027 997 1036
rect 1000 1034 1002 1036
rect 1021 1034 1023 1036
rect 1037 1033 1039 1036
rect 995 1017 997 1020
rect 1000 1017 1002 1019
rect 1021 1017 1023 1019
rect 1037 1017 1039 1029
rect 1053 1027 1055 1036
rect 1058 1034 1060 1036
rect 1053 1017 1055 1020
rect 1058 1017 1060 1019
rect 1074 1017 1076 1036
rect 1090 1033 1092 1036
rect 1095 1034 1097 1036
rect 1090 1017 1092 1029
rect 1095 1017 1097 1024
rect 1111 1017 1113 1036
rect 1127 1027 1129 1036
rect 1132 1034 1134 1036
rect 1153 1034 1155 1036
rect 1169 1033 1171 1036
rect 1127 1017 1129 1020
rect 1132 1017 1134 1019
rect 1153 1017 1155 1019
rect 1169 1017 1171 1029
rect 1185 1027 1187 1036
rect 1190 1034 1192 1036
rect 1185 1017 1187 1020
rect 1190 1017 1192 1019
rect 1206 1017 1208 1036
rect 1222 1033 1224 1036
rect 1227 1034 1229 1036
rect 1222 1017 1224 1029
rect 1227 1017 1229 1024
rect 1243 1017 1245 1036
rect 1259 1027 1261 1036
rect 1264 1034 1266 1036
rect 1285 1034 1287 1036
rect 1301 1033 1303 1036
rect 1259 1017 1261 1020
rect 1264 1017 1266 1019
rect 1285 1017 1287 1019
rect 1301 1017 1303 1029
rect 1317 1027 1319 1036
rect 1322 1034 1324 1036
rect 1338 1028 1340 1036
rect 1317 1017 1319 1020
rect 1322 1017 1324 1019
rect 1338 1017 1340 1024
rect 25 1011 27 1013
rect 30 1010 32 1013
rect 46 1011 48 1013
rect 62 1011 64 1013
rect 67 1008 69 1013
rect 88 1008 90 1013
rect 104 1011 106 1013
rect 120 1011 122 1013
rect 125 1008 127 1013
rect 141 1011 143 1013
rect 157 1011 159 1013
rect 162 1010 164 1013
rect 178 1011 180 1013
rect 194 1011 196 1013
rect 199 1008 201 1013
rect 220 1008 222 1013
rect 236 1011 238 1013
rect 252 1011 254 1013
rect 257 1008 259 1013
rect 273 1011 275 1013
rect 289 1011 291 1013
rect 294 1010 296 1013
rect 310 1011 312 1013
rect 326 1011 328 1013
rect 331 1008 333 1013
rect 352 1008 354 1013
rect 368 1011 370 1013
rect 384 1011 386 1013
rect 389 1008 391 1013
rect 405 1011 407 1013
rect 958 1011 960 1013
rect 963 1010 965 1013
rect 979 1011 981 1013
rect 995 1011 997 1013
rect 1000 1008 1002 1013
rect 1021 1008 1023 1013
rect 1037 1011 1039 1013
rect 1053 1011 1055 1013
rect 1058 1008 1060 1013
rect 1074 1011 1076 1013
rect 1090 1011 1092 1013
rect 1095 1010 1097 1013
rect 1111 1011 1113 1013
rect 1127 1011 1129 1013
rect 1132 1008 1134 1013
rect 1153 1008 1155 1013
rect 1169 1011 1171 1013
rect 1185 1011 1187 1013
rect 1190 1008 1192 1013
rect 1206 1011 1208 1013
rect 1222 1011 1224 1013
rect 1227 1010 1229 1013
rect 1243 1011 1245 1013
rect 1259 1011 1261 1013
rect 1264 1008 1266 1013
rect 1285 1008 1287 1013
rect 1301 1011 1303 1013
rect 1317 1011 1319 1013
rect 1322 1008 1324 1013
rect 1338 1011 1340 1013
rect 497 965 499 967
rect 502 965 504 968
rect 518 965 520 967
rect 534 965 536 967
rect 539 965 541 968
rect 560 965 562 968
rect 576 965 578 968
rect 592 965 594 967
rect 597 965 599 968
rect 613 965 615 967
rect 629 965 631 967
rect 634 965 636 968
rect 650 965 652 967
rect 666 965 668 967
rect 671 965 673 968
rect 692 965 694 968
rect 708 965 710 968
rect 724 965 726 967
rect 729 965 731 968
rect 745 965 747 967
rect 761 965 763 967
rect 766 965 768 968
rect 782 965 784 967
rect 798 965 800 967
rect 803 965 805 968
rect 824 965 826 968
rect 840 965 842 968
rect 856 965 858 967
rect 861 965 863 968
rect 877 965 879 967
rect 893 965 895 967
rect 898 965 900 968
rect 914 965 916 967
rect 930 965 932 967
rect 935 965 937 968
rect 956 965 958 968
rect 972 965 974 968
rect 988 965 990 967
rect 993 965 995 968
rect 1009 965 1011 967
rect 1430 965 1432 967
rect 1435 965 1437 968
rect 1451 965 1453 967
rect 1467 965 1469 967
rect 1472 965 1474 968
rect 1493 965 1495 968
rect 1509 965 1511 968
rect 1525 965 1527 967
rect 1530 965 1532 968
rect 1546 965 1548 967
rect 1562 965 1564 967
rect 1567 965 1569 968
rect 1583 965 1585 967
rect 1599 965 1601 967
rect 1604 965 1606 968
rect 1625 965 1627 968
rect 1641 965 1643 968
rect 1657 965 1659 967
rect 1662 965 1664 968
rect 1678 965 1680 967
rect 1694 965 1696 967
rect 1699 965 1701 968
rect 1715 965 1717 967
rect 1731 965 1733 967
rect 1736 965 1738 968
rect 1757 965 1759 968
rect 1773 965 1775 968
rect 1789 965 1791 967
rect 1794 965 1796 968
rect 1810 965 1812 967
rect 1826 965 1828 967
rect 1831 965 1833 968
rect 1847 965 1849 967
rect 1863 965 1865 967
rect 1868 965 1870 968
rect 1889 965 1891 968
rect 1905 965 1907 968
rect 1921 965 1923 967
rect 1926 965 1928 968
rect 1942 965 1944 967
rect 497 952 499 957
rect 502 955 504 957
rect 497 938 499 948
rect 502 938 504 945
rect 518 938 520 957
rect 534 948 536 957
rect 539 955 541 957
rect 560 955 562 957
rect 576 954 578 957
rect 534 938 536 941
rect 539 938 541 940
rect 560 938 562 940
rect 576 938 578 950
rect 592 948 594 957
rect 597 955 599 957
rect 613 949 615 957
rect 629 952 631 957
rect 634 955 636 957
rect 592 938 594 941
rect 597 938 599 940
rect 613 938 615 945
rect 629 938 631 948
rect 634 938 636 945
rect 650 938 652 957
rect 666 948 668 957
rect 671 955 673 957
rect 692 955 694 957
rect 708 954 710 957
rect 666 938 668 941
rect 671 938 673 940
rect 692 938 694 940
rect 708 938 710 950
rect 724 948 726 957
rect 729 955 731 957
rect 745 949 747 957
rect 761 952 763 957
rect 766 955 768 957
rect 724 938 726 941
rect 729 938 731 940
rect 745 938 747 945
rect 761 938 763 948
rect 766 938 768 945
rect 782 938 784 957
rect 798 948 800 957
rect 803 955 805 957
rect 824 955 826 957
rect 840 954 842 957
rect 798 938 800 941
rect 803 938 805 940
rect 824 938 826 940
rect 840 938 842 950
rect 856 948 858 957
rect 861 955 863 957
rect 877 949 879 957
rect 893 952 895 957
rect 898 955 900 957
rect 856 938 858 941
rect 861 938 863 940
rect 877 938 879 945
rect 893 938 895 948
rect 898 938 900 945
rect 914 938 916 957
rect 930 948 932 957
rect 935 955 937 957
rect 956 955 958 957
rect 972 954 974 957
rect 930 938 932 941
rect 935 938 937 940
rect 956 938 958 940
rect 972 938 974 950
rect 988 948 990 957
rect 993 955 995 957
rect 1009 949 1011 957
rect 1430 952 1432 957
rect 1435 955 1437 957
rect 988 938 990 941
rect 993 938 995 940
rect 1009 938 1011 945
rect 157 932 159 934
rect 162 932 164 935
rect 178 932 180 934
rect 194 932 196 934
rect 199 932 201 935
rect 220 932 222 935
rect 236 932 238 935
rect 252 932 254 934
rect 257 932 259 935
rect 1430 938 1432 948
rect 1435 938 1437 945
rect 1451 938 1453 957
rect 1467 948 1469 957
rect 1472 955 1474 957
rect 1493 955 1495 957
rect 1509 954 1511 957
rect 1467 938 1469 941
rect 1472 938 1474 940
rect 1493 938 1495 940
rect 1509 938 1511 950
rect 1525 948 1527 957
rect 1530 955 1532 957
rect 1546 949 1548 957
rect 1562 952 1564 957
rect 1567 955 1569 957
rect 1525 938 1527 941
rect 1530 938 1532 940
rect 1546 938 1548 945
rect 1562 938 1564 948
rect 1567 938 1569 945
rect 1583 938 1585 957
rect 1599 948 1601 957
rect 1604 955 1606 957
rect 1625 955 1627 957
rect 1641 954 1643 957
rect 1599 938 1601 941
rect 1604 938 1606 940
rect 1625 938 1627 940
rect 1641 938 1643 950
rect 1657 948 1659 957
rect 1662 955 1664 957
rect 1678 949 1680 957
rect 1694 952 1696 957
rect 1699 955 1701 957
rect 1657 938 1659 941
rect 1662 938 1664 940
rect 1678 938 1680 945
rect 1694 938 1696 948
rect 1699 938 1701 945
rect 1715 938 1717 957
rect 1731 948 1733 957
rect 1736 955 1738 957
rect 1757 955 1759 957
rect 1773 954 1775 957
rect 1731 938 1733 941
rect 1736 938 1738 940
rect 1757 938 1759 940
rect 1773 938 1775 950
rect 1789 948 1791 957
rect 1794 955 1796 957
rect 1810 949 1812 957
rect 1826 952 1828 957
rect 1831 955 1833 957
rect 1789 938 1791 941
rect 1794 938 1796 940
rect 1810 938 1812 945
rect 1826 938 1828 948
rect 1831 938 1833 945
rect 1847 938 1849 957
rect 1863 948 1865 957
rect 1868 955 1870 957
rect 1889 955 1891 957
rect 1905 954 1907 957
rect 1863 938 1865 941
rect 1868 938 1870 940
rect 1889 938 1891 940
rect 1905 938 1907 950
rect 1921 948 1923 957
rect 1926 955 1928 957
rect 1942 949 1944 957
rect 1921 938 1923 941
rect 1926 938 1928 940
rect 1942 938 1944 945
rect 273 932 275 934
rect 497 932 499 934
rect 502 931 504 934
rect 518 932 520 934
rect 534 932 536 934
rect 539 929 541 934
rect 560 929 562 934
rect 576 932 578 934
rect 592 932 594 934
rect 597 929 599 934
rect 613 932 615 934
rect 629 932 631 934
rect 634 931 636 934
rect 650 932 652 934
rect 666 932 668 934
rect 671 929 673 934
rect 692 929 694 934
rect 708 932 710 934
rect 724 932 726 934
rect 729 929 731 934
rect 745 932 747 934
rect 761 932 763 934
rect 766 931 768 934
rect 782 932 784 934
rect 798 932 800 934
rect 803 929 805 934
rect 824 929 826 934
rect 840 932 842 934
rect 856 932 858 934
rect 861 929 863 934
rect 877 932 879 934
rect 893 932 895 934
rect 898 931 900 934
rect 914 932 916 934
rect 930 932 932 934
rect 935 929 937 934
rect 956 929 958 934
rect 972 932 974 934
rect 988 932 990 934
rect 993 929 995 934
rect 1009 932 1011 934
rect 1090 932 1092 934
rect 1095 932 1097 935
rect 1111 932 1113 934
rect 1127 932 1129 934
rect 1132 932 1134 935
rect 1153 932 1155 935
rect 1169 932 1171 935
rect 1185 932 1187 934
rect 1190 932 1192 935
rect 1206 932 1208 934
rect 1430 932 1432 934
rect 1435 931 1437 934
rect 1451 932 1453 934
rect 1467 932 1469 934
rect 1472 929 1474 934
rect 1493 929 1495 934
rect 1509 932 1511 934
rect 1525 932 1527 934
rect 1530 929 1532 934
rect 1546 932 1548 934
rect 1562 932 1564 934
rect 1567 931 1569 934
rect 1583 932 1585 934
rect 1599 932 1601 934
rect 1604 929 1606 934
rect 1625 929 1627 934
rect 1641 932 1643 934
rect 1657 932 1659 934
rect 1662 929 1664 934
rect 1678 932 1680 934
rect 1694 932 1696 934
rect 1699 931 1701 934
rect 1715 932 1717 934
rect 1731 932 1733 934
rect 1736 929 1738 934
rect 1757 929 1759 934
rect 1773 932 1775 934
rect 1789 932 1791 934
rect 1794 929 1796 934
rect 1810 932 1812 934
rect 1826 932 1828 934
rect 1831 931 1833 934
rect 1847 932 1849 934
rect 1863 932 1865 934
rect 1868 929 1870 934
rect 1889 929 1891 934
rect 1905 932 1907 934
rect 1921 932 1923 934
rect 1926 929 1928 934
rect 1942 932 1944 934
rect 157 919 159 924
rect 162 922 164 924
rect 157 905 159 915
rect 162 905 164 912
rect 178 905 180 924
rect 194 915 196 924
rect 199 922 201 924
rect 220 922 222 924
rect 236 921 238 924
rect 194 905 196 908
rect 199 905 201 907
rect 220 905 222 907
rect 236 905 238 917
rect 252 915 254 924
rect 257 922 259 924
rect 252 905 254 908
rect 257 905 259 907
rect 273 905 275 924
rect 1090 919 1092 924
rect 1095 922 1097 924
rect 1090 905 1092 915
rect 1095 905 1097 912
rect 1111 905 1113 924
rect 1127 915 1129 924
rect 1132 922 1134 924
rect 1153 922 1155 924
rect 1169 921 1171 924
rect 1127 905 1129 908
rect 1132 905 1134 907
rect 1153 905 1155 907
rect 1169 905 1171 917
rect 1185 915 1187 924
rect 1190 922 1192 924
rect 1185 905 1187 908
rect 1190 905 1192 907
rect 1206 905 1208 924
rect 157 899 159 901
rect 162 898 164 901
rect 178 899 180 901
rect 194 899 196 901
rect 199 896 201 901
rect 220 896 222 901
rect 236 899 238 901
rect 252 899 254 901
rect 257 896 259 901
rect 273 899 275 901
rect 1090 899 1092 901
rect 1095 898 1097 901
rect 1111 899 1113 901
rect 1127 899 1129 901
rect 676 894 678 896
rect 518 888 520 891
rect 562 888 564 891
rect 588 888 590 891
rect 634 888 636 891
rect 588 884 589 888
rect 702 888 704 892
rect 730 894 732 896
rect 757 894 759 896
rect 707 888 709 891
rect 502 881 504 883
rect 518 881 520 884
rect 534 881 536 883
rect 557 881 559 883
rect 562 881 564 884
rect 588 881 590 884
rect 609 881 611 884
rect 629 881 631 883
rect 634 881 636 884
rect 652 881 654 883
rect 281 868 283 871
rect 281 862 283 864
rect 164 859 166 862
rect 502 859 504 873
rect 518 871 520 873
rect 518 859 520 861
rect 534 859 536 873
rect 557 868 559 873
rect 562 871 564 873
rect 588 871 590 873
rect 553 864 559 868
rect 557 859 559 864
rect 562 859 564 861
rect 588 859 590 861
rect 609 859 611 873
rect 629 868 631 873
rect 634 871 636 873
rect 625 864 631 868
rect 629 859 631 864
rect 634 859 636 861
rect 652 859 654 873
rect 676 872 678 886
rect 783 888 785 892
rect 811 894 813 896
rect 1132 896 1134 901
rect 1153 896 1155 901
rect 1169 899 1171 901
rect 1185 899 1187 901
rect 1190 896 1192 901
rect 1206 899 1208 901
rect 788 888 790 891
rect 702 877 704 880
rect 707 878 709 880
rect 703 873 704 877
rect 702 868 704 873
rect 707 868 709 870
rect 676 866 678 868
rect 730 864 732 886
rect 757 872 759 886
rect 1609 894 1611 896
rect 783 877 785 880
rect 788 878 790 880
rect 784 873 785 877
rect 783 868 785 873
rect 788 868 790 870
rect 757 866 759 868
rect 811 864 813 886
rect 1451 888 1453 891
rect 1495 888 1497 891
rect 1521 888 1523 891
rect 1567 888 1569 891
rect 1521 884 1522 888
rect 1635 888 1637 892
rect 1663 894 1665 896
rect 1690 894 1692 896
rect 1640 888 1642 891
rect 1435 881 1437 883
rect 1451 881 1453 884
rect 1467 881 1469 883
rect 1490 881 1492 883
rect 1495 881 1497 884
rect 1521 881 1523 884
rect 1542 881 1544 884
rect 1562 881 1564 883
rect 1567 881 1569 884
rect 1585 881 1587 883
rect 1214 868 1216 871
rect 702 862 704 864
rect 707 859 709 864
rect 783 862 785 864
rect 730 858 732 860
rect 788 859 790 864
rect 1214 862 1216 864
rect 811 858 813 860
rect 1097 859 1099 862
rect 1435 859 1437 873
rect 1451 871 1453 873
rect 1451 859 1453 861
rect 1467 859 1469 873
rect 1490 868 1492 873
rect 1495 871 1497 873
rect 1521 871 1523 873
rect 1486 864 1492 868
rect 1490 859 1492 864
rect 1495 859 1497 861
rect 1521 859 1523 861
rect 1542 859 1544 873
rect 1562 868 1564 873
rect 1567 871 1569 873
rect 1558 864 1564 868
rect 1562 859 1564 864
rect 1567 859 1569 861
rect 1585 859 1587 873
rect 1609 872 1611 886
rect 1716 888 1718 892
rect 1744 894 1746 896
rect 1721 888 1723 891
rect 1635 877 1637 880
rect 1640 878 1642 880
rect 1636 873 1637 877
rect 1635 868 1637 873
rect 1640 868 1642 870
rect 1609 866 1611 868
rect 1663 864 1665 886
rect 1690 872 1692 886
rect 1716 877 1718 880
rect 1721 878 1723 880
rect 1717 873 1718 877
rect 1716 868 1718 873
rect 1721 868 1723 870
rect 1690 866 1692 868
rect 1744 864 1746 886
rect 1635 862 1637 864
rect 1640 859 1642 864
rect 1716 862 1718 864
rect 1663 858 1665 860
rect 1721 859 1723 864
rect 1744 858 1746 860
rect 164 853 166 855
rect 502 853 504 855
rect 518 851 520 855
rect 534 853 536 855
rect 557 853 559 855
rect 519 847 520 851
rect 562 850 564 855
rect 588 851 590 855
rect 609 853 611 855
rect 629 853 631 855
rect 518 844 520 847
rect 563 846 564 850
rect 589 847 590 851
rect 634 850 636 855
rect 652 853 654 855
rect 1097 853 1099 855
rect 1435 853 1437 855
rect 1451 851 1453 855
rect 1467 853 1469 855
rect 1490 853 1492 855
rect 562 844 564 846
rect 588 843 590 847
rect 635 846 636 850
rect 1452 847 1453 851
rect 1495 850 1497 855
rect 1521 851 1523 855
rect 1542 853 1544 855
rect 1562 853 1564 855
rect 634 844 636 846
rect 1451 844 1453 847
rect 1496 846 1497 850
rect 1522 847 1523 851
rect 1567 850 1569 855
rect 1585 853 1587 855
rect 1495 844 1497 846
rect 1521 843 1523 847
rect 1568 846 1569 850
rect 1567 844 1569 846
rect 148 830 150 832
rect 164 830 166 833
rect 169 830 171 832
rect 185 830 187 833
rect 201 830 203 833
rect 222 830 224 833
rect 227 830 229 832
rect 243 830 245 832
rect 259 830 261 833
rect 264 830 266 832
rect 1081 830 1083 832
rect 1097 830 1099 833
rect 1102 830 1104 832
rect 1118 830 1120 833
rect 1134 830 1136 833
rect 1155 830 1157 833
rect 1160 830 1162 832
rect 1176 830 1178 832
rect 1192 830 1194 833
rect 1197 830 1199 832
rect 148 803 150 822
rect 164 820 166 822
rect 169 813 171 822
rect 185 819 187 822
rect 201 820 203 822
rect 222 820 224 822
rect 164 803 166 805
rect 169 803 171 806
rect 185 803 187 815
rect 227 813 229 822
rect 201 803 203 805
rect 222 803 224 805
rect 227 803 229 806
rect 243 803 245 822
rect 259 820 261 822
rect 264 817 266 822
rect 518 821 520 824
rect 562 822 564 824
rect 519 817 520 821
rect 563 818 564 822
rect 588 821 590 825
rect 634 822 636 824
rect 502 813 504 815
rect 518 813 520 817
rect 534 813 536 815
rect 557 813 559 815
rect 562 813 564 818
rect 589 817 590 821
rect 635 818 636 822
rect 588 813 590 817
rect 609 813 611 815
rect 629 813 631 815
rect 634 813 636 818
rect 652 813 654 815
rect 259 803 261 810
rect 264 803 266 813
rect 702 812 704 815
rect 707 812 709 815
rect 783 812 785 815
rect 788 812 790 815
rect 148 797 150 799
rect 164 794 166 799
rect 169 797 171 799
rect 185 797 187 799
rect 201 794 203 799
rect 222 794 224 799
rect 227 797 229 799
rect 243 797 245 799
rect 259 796 261 799
rect 264 797 266 799
rect 502 795 504 809
rect 518 807 520 809
rect 518 795 520 797
rect 534 795 536 809
rect 557 804 559 809
rect 562 807 564 809
rect 588 807 590 809
rect 553 800 559 804
rect 557 795 559 800
rect 562 795 564 797
rect 588 795 590 797
rect 609 795 611 809
rect 629 804 631 809
rect 634 807 636 809
rect 625 800 631 804
rect 629 795 631 800
rect 634 795 636 797
rect 652 795 654 809
rect 702 796 704 808
rect 707 806 709 808
rect 707 796 709 798
rect 783 796 785 808
rect 788 806 790 808
rect 1081 803 1083 822
rect 1097 820 1099 822
rect 1102 813 1104 822
rect 1118 819 1120 822
rect 1134 820 1136 822
rect 1155 820 1157 822
rect 1097 803 1099 805
rect 1102 803 1104 806
rect 1118 803 1120 815
rect 1160 813 1162 822
rect 1134 803 1136 805
rect 1155 803 1157 805
rect 1160 803 1162 806
rect 1176 803 1178 822
rect 1192 820 1194 822
rect 1197 817 1199 822
rect 1451 821 1453 824
rect 1495 822 1497 824
rect 1452 817 1453 821
rect 1496 818 1497 822
rect 1521 821 1523 825
rect 1567 822 1569 824
rect 1435 813 1437 815
rect 1451 813 1453 817
rect 1467 813 1469 815
rect 1490 813 1492 815
rect 1495 813 1497 818
rect 1522 817 1523 821
rect 1568 818 1569 822
rect 1521 813 1523 817
rect 1542 813 1544 815
rect 1562 813 1564 815
rect 1567 813 1569 818
rect 1585 813 1587 815
rect 1192 803 1194 810
rect 1197 803 1199 813
rect 1635 812 1637 815
rect 1640 812 1642 815
rect 1716 812 1718 815
rect 1721 812 1723 815
rect 788 796 790 798
rect 1081 797 1083 799
rect 1097 794 1099 799
rect 1102 797 1104 799
rect 1118 797 1120 799
rect 1134 794 1136 799
rect 1155 794 1157 799
rect 1160 797 1162 799
rect 1176 797 1178 799
rect 1192 796 1194 799
rect 1197 797 1199 799
rect 1435 795 1437 809
rect 1451 807 1453 809
rect 1451 795 1453 797
rect 1467 795 1469 809
rect 1490 804 1492 809
rect 1495 807 1497 809
rect 1521 807 1523 809
rect 1486 800 1492 804
rect 1490 795 1492 800
rect 1495 795 1497 797
rect 1521 795 1523 797
rect 1542 795 1544 809
rect 1562 804 1564 809
rect 1567 807 1569 809
rect 1558 800 1564 804
rect 1562 795 1564 800
rect 1567 795 1569 797
rect 1585 795 1587 809
rect 1635 796 1637 808
rect 1640 806 1642 808
rect 1640 796 1642 798
rect 1716 796 1718 808
rect 1721 806 1723 808
rect 1721 796 1723 798
rect 502 785 504 787
rect 518 784 520 787
rect 534 785 536 787
rect 557 785 559 787
rect 562 784 564 787
rect 588 784 590 787
rect 609 784 611 787
rect 629 785 631 787
rect 634 784 636 787
rect 652 785 654 787
rect 702 786 704 788
rect 588 780 589 784
rect 707 783 709 788
rect 783 786 785 788
rect 788 783 790 788
rect 1435 785 1437 787
rect 1451 784 1453 787
rect 1467 785 1469 787
rect 1490 785 1492 787
rect 1495 784 1497 787
rect 1521 784 1523 787
rect 1542 784 1544 787
rect 1562 785 1564 787
rect 1567 784 1569 787
rect 1585 785 1587 787
rect 1635 786 1637 788
rect 518 777 520 780
rect 562 777 564 780
rect 588 777 590 780
rect 634 777 636 780
rect 1521 780 1522 784
rect 1640 783 1642 788
rect 1716 786 1718 788
rect 1721 783 1723 788
rect 1451 777 1453 780
rect 1495 777 1497 780
rect 1521 777 1523 780
rect 1567 777 1569 780
rect 518 756 520 759
rect 562 756 564 759
rect 588 756 590 759
rect 634 756 636 759
rect 702 756 704 760
rect 730 762 732 764
rect 781 762 783 764
rect 707 756 709 759
rect 588 752 589 756
rect 502 749 504 751
rect 518 749 520 752
rect 534 749 536 751
rect 557 749 559 751
rect 562 749 564 752
rect 588 749 590 752
rect 609 749 611 752
rect 629 749 631 751
rect 634 749 636 752
rect 652 749 654 751
rect 807 756 809 760
rect 835 762 837 764
rect 812 756 814 759
rect 702 745 704 748
rect 707 746 709 748
rect 703 741 704 745
rect 502 727 504 741
rect 518 739 520 741
rect 518 727 520 729
rect 534 727 536 741
rect 557 736 559 741
rect 562 739 564 741
rect 588 739 590 741
rect 553 732 559 736
rect 557 727 559 732
rect 562 727 564 729
rect 588 727 590 729
rect 609 727 611 741
rect 629 736 631 741
rect 634 739 636 741
rect 625 732 631 736
rect 629 727 631 732
rect 634 727 636 729
rect 652 727 654 741
rect 702 736 704 741
rect 707 736 709 738
rect 730 732 732 754
rect 781 740 783 754
rect 1451 756 1453 759
rect 1495 756 1497 759
rect 1521 756 1523 759
rect 1567 756 1569 759
rect 1635 756 1637 760
rect 1663 762 1665 764
rect 1714 762 1716 764
rect 1640 756 1642 759
rect 807 745 809 748
rect 812 746 814 748
rect 808 741 809 745
rect 807 736 809 741
rect 812 736 814 738
rect 781 734 783 736
rect 835 732 837 754
rect 1521 752 1522 756
rect 1435 749 1437 751
rect 1451 749 1453 752
rect 1467 749 1469 751
rect 1490 749 1492 751
rect 1495 749 1497 752
rect 1521 749 1523 752
rect 1542 749 1544 752
rect 1562 749 1564 751
rect 1567 749 1569 752
rect 1585 749 1587 751
rect 1740 756 1742 760
rect 1768 762 1770 764
rect 1745 756 1747 759
rect 1635 745 1637 748
rect 1640 746 1642 748
rect 1636 741 1637 745
rect 702 730 704 732
rect 707 727 709 732
rect 807 730 809 732
rect 730 726 732 728
rect 812 727 814 732
rect 835 726 837 728
rect 1435 727 1437 741
rect 1451 739 1453 741
rect 1451 727 1453 729
rect 1467 727 1469 741
rect 1490 736 1492 741
rect 1495 739 1497 741
rect 1521 739 1523 741
rect 1486 732 1492 736
rect 1490 727 1492 732
rect 1495 727 1497 729
rect 1521 727 1523 729
rect 1542 727 1544 741
rect 1562 736 1564 741
rect 1567 739 1569 741
rect 1558 732 1564 736
rect 1562 727 1564 732
rect 1567 727 1569 729
rect 1585 727 1587 741
rect 1635 736 1637 741
rect 1640 736 1642 738
rect 1663 732 1665 754
rect 1714 740 1716 754
rect 1740 745 1742 748
rect 1745 746 1747 748
rect 1741 741 1742 745
rect 1740 736 1742 741
rect 1745 736 1747 738
rect 1714 734 1716 736
rect 1768 732 1770 754
rect 1635 730 1637 732
rect 1640 727 1642 732
rect 1740 730 1742 732
rect 1663 726 1665 728
rect 1745 727 1747 732
rect 1768 726 1770 728
rect 502 721 504 723
rect 518 719 520 723
rect 534 721 536 723
rect 557 721 559 723
rect 519 715 520 719
rect 562 718 564 723
rect 588 719 590 723
rect 609 721 611 723
rect 629 721 631 723
rect 518 712 520 715
rect 563 714 564 718
rect 589 715 590 719
rect 634 718 636 723
rect 652 721 654 723
rect 1435 721 1437 723
rect 1451 719 1453 723
rect 1467 721 1469 723
rect 1490 721 1492 723
rect 562 712 564 714
rect 588 711 590 715
rect 635 714 636 718
rect 1452 715 1453 719
rect 1495 718 1497 723
rect 1521 719 1523 723
rect 1542 721 1544 723
rect 1562 721 1564 723
rect 634 712 636 714
rect 1451 712 1453 715
rect 1496 714 1497 718
rect 1522 715 1523 719
rect 1567 718 1569 723
rect 1585 721 1587 723
rect 1495 712 1497 714
rect 1521 711 1523 715
rect 1568 714 1569 718
rect 1567 712 1569 714
rect 518 689 520 692
rect 562 690 564 692
rect 519 685 520 689
rect 563 686 564 690
rect 588 689 590 693
rect 634 690 636 692
rect 502 681 504 683
rect 518 681 520 685
rect 534 681 536 683
rect 557 681 559 683
rect 562 681 564 686
rect 589 685 590 689
rect 635 686 636 690
rect 1451 689 1453 692
rect 1495 690 1497 692
rect 588 681 590 685
rect 609 681 611 683
rect 629 681 631 683
rect 634 681 636 686
rect 1452 685 1453 689
rect 1496 686 1497 690
rect 1521 689 1523 693
rect 1567 690 1569 692
rect 652 681 654 683
rect 702 681 704 684
rect 707 681 709 684
rect 807 681 809 684
rect 812 681 814 684
rect 1435 681 1437 683
rect 1451 681 1453 685
rect 1467 681 1469 683
rect 1490 681 1492 683
rect 1495 681 1497 686
rect 1522 685 1523 689
rect 1568 686 1569 690
rect 1521 681 1523 685
rect 1542 681 1544 683
rect 1562 681 1564 683
rect 1567 681 1569 686
rect 1585 681 1587 683
rect 1635 681 1637 684
rect 1640 681 1642 684
rect 1740 681 1742 684
rect 1745 681 1747 684
rect 502 663 504 677
rect 518 675 520 677
rect 518 663 520 665
rect 534 663 536 677
rect 557 672 559 677
rect 562 675 564 677
rect 588 675 590 677
rect 553 668 559 672
rect 557 663 559 668
rect 562 663 564 665
rect 588 663 590 665
rect 609 663 611 677
rect 629 672 631 677
rect 634 675 636 677
rect 625 668 631 672
rect 629 663 631 668
rect 634 663 636 665
rect 652 663 654 677
rect 702 665 704 677
rect 707 675 709 677
rect 707 665 709 667
rect 807 665 809 677
rect 812 675 814 677
rect 812 665 814 667
rect 1435 663 1437 677
rect 1451 675 1453 677
rect 1451 663 1453 665
rect 1467 663 1469 677
rect 1490 672 1492 677
rect 1495 675 1497 677
rect 1521 675 1523 677
rect 1486 668 1492 672
rect 1490 663 1492 668
rect 1495 663 1497 665
rect 1521 663 1523 665
rect 1542 663 1544 677
rect 1562 672 1564 677
rect 1567 675 1569 677
rect 1558 668 1564 672
rect 1562 663 1564 668
rect 1567 663 1569 665
rect 1585 663 1587 677
rect 1635 665 1637 677
rect 1640 675 1642 677
rect 1640 665 1642 667
rect 1740 665 1742 677
rect 1745 675 1747 677
rect 1745 665 1747 667
rect 702 655 704 657
rect 502 653 504 655
rect 518 652 520 655
rect 534 653 536 655
rect 557 653 559 655
rect 562 652 564 655
rect 588 652 590 655
rect 609 652 611 655
rect 629 653 631 655
rect 634 652 636 655
rect 652 653 654 655
rect 707 652 709 657
rect 807 655 809 657
rect 812 652 814 657
rect 1635 655 1637 657
rect 1435 653 1437 655
rect 588 648 589 652
rect 1451 652 1453 655
rect 1467 653 1469 655
rect 1490 653 1492 655
rect 1495 652 1497 655
rect 1521 652 1523 655
rect 1542 652 1544 655
rect 1562 653 1564 655
rect 1567 652 1569 655
rect 1585 653 1587 655
rect 1640 652 1642 657
rect 1740 655 1742 657
rect 1745 652 1747 657
rect 1521 648 1522 652
rect 518 645 520 648
rect 562 645 564 648
rect 588 645 590 648
rect 634 645 636 648
rect 1451 645 1453 648
rect 1495 645 1497 648
rect 1521 645 1523 648
rect 1567 645 1569 648
rect 518 624 520 627
rect 562 624 564 627
rect 588 624 590 627
rect 634 624 636 627
rect 702 624 704 628
rect 730 630 732 632
rect 757 630 759 632
rect 707 624 709 627
rect 588 620 589 624
rect 502 617 504 619
rect 518 617 520 620
rect 534 617 536 619
rect 557 617 559 619
rect 562 617 564 620
rect 588 617 590 620
rect 609 617 611 620
rect 629 617 631 619
rect 634 617 636 620
rect 652 617 654 619
rect 783 624 785 628
rect 811 630 813 632
rect 847 630 849 632
rect 788 624 790 627
rect 702 613 704 616
rect 707 614 709 616
rect 703 609 704 613
rect 502 595 504 609
rect 518 607 520 609
rect 518 595 520 597
rect 534 595 536 609
rect 557 604 559 609
rect 562 607 564 609
rect 588 607 590 609
rect 553 600 559 604
rect 557 595 559 600
rect 562 595 564 597
rect 588 595 590 597
rect 609 595 611 609
rect 629 604 631 609
rect 634 607 636 609
rect 625 600 631 604
rect 629 595 631 600
rect 634 595 636 597
rect 652 595 654 609
rect 702 604 704 609
rect 707 604 709 606
rect 730 600 732 622
rect 757 608 759 622
rect 873 624 875 628
rect 901 630 903 632
rect 878 624 880 627
rect 783 613 785 616
rect 788 614 790 616
rect 784 609 785 613
rect 783 604 785 609
rect 788 604 790 606
rect 757 602 759 604
rect 811 600 813 622
rect 847 608 849 622
rect 1451 624 1453 627
rect 1495 624 1497 627
rect 1521 624 1523 627
rect 1567 624 1569 627
rect 1635 624 1637 628
rect 1663 630 1665 632
rect 1690 630 1692 632
rect 1640 624 1642 627
rect 873 613 875 616
rect 878 614 880 616
rect 874 609 875 613
rect 873 604 875 609
rect 878 604 880 606
rect 847 602 849 604
rect 901 600 903 622
rect 1521 620 1522 624
rect 1435 617 1437 619
rect 1451 617 1453 620
rect 1467 617 1469 619
rect 1490 617 1492 619
rect 1495 617 1497 620
rect 1521 617 1523 620
rect 1542 617 1544 620
rect 1562 617 1564 619
rect 1567 617 1569 620
rect 1585 617 1587 619
rect 1716 624 1718 628
rect 1744 630 1746 632
rect 1780 630 1782 632
rect 1721 624 1723 627
rect 1635 613 1637 616
rect 1640 614 1642 616
rect 1636 609 1637 613
rect 702 598 704 600
rect 707 595 709 600
rect 783 598 785 600
rect 730 594 732 596
rect 788 595 790 600
rect 873 598 875 600
rect 811 594 813 596
rect 878 595 880 600
rect 901 594 903 596
rect 1435 595 1437 609
rect 1451 607 1453 609
rect 1451 595 1453 597
rect 1467 595 1469 609
rect 1490 604 1492 609
rect 1495 607 1497 609
rect 1521 607 1523 609
rect 1486 600 1492 604
rect 1490 595 1492 600
rect 1495 595 1497 597
rect 1521 595 1523 597
rect 1542 595 1544 609
rect 1562 604 1564 609
rect 1567 607 1569 609
rect 1558 600 1564 604
rect 1562 595 1564 600
rect 1567 595 1569 597
rect 1585 595 1587 609
rect 1635 604 1637 609
rect 1640 604 1642 606
rect 1663 600 1665 622
rect 1690 608 1692 622
rect 1806 624 1808 628
rect 1834 630 1836 632
rect 1811 624 1813 627
rect 1716 613 1718 616
rect 1721 614 1723 616
rect 1717 609 1718 613
rect 1716 604 1718 609
rect 1721 604 1723 606
rect 1690 602 1692 604
rect 1744 600 1746 622
rect 1780 608 1782 622
rect 1806 613 1808 616
rect 1811 614 1813 616
rect 1807 609 1808 613
rect 1806 604 1808 609
rect 1811 604 1813 606
rect 1780 602 1782 604
rect 1834 600 1836 622
rect 1635 598 1637 600
rect 1640 595 1642 600
rect 1716 598 1718 600
rect 1663 594 1665 596
rect 1721 595 1723 600
rect 1806 598 1808 600
rect 1744 594 1746 596
rect 1811 595 1813 600
rect 1834 594 1836 596
rect 502 589 504 591
rect 518 587 520 591
rect 534 589 536 591
rect 557 589 559 591
rect 519 583 520 587
rect 562 586 564 591
rect 588 587 590 591
rect 609 589 611 591
rect 629 589 631 591
rect 518 580 520 583
rect 563 582 564 586
rect 589 583 590 587
rect 634 586 636 591
rect 652 589 654 591
rect 1435 589 1437 591
rect 1451 587 1453 591
rect 1467 589 1469 591
rect 1490 589 1492 591
rect 562 580 564 582
rect 588 579 590 583
rect 635 582 636 586
rect 1452 583 1453 587
rect 1495 586 1497 591
rect 1521 587 1523 591
rect 1542 589 1544 591
rect 1562 589 1564 591
rect 634 580 636 582
rect 1451 580 1453 583
rect 1496 582 1497 586
rect 1522 583 1523 587
rect 1567 586 1569 591
rect 1585 589 1587 591
rect 1495 580 1497 582
rect 1521 579 1523 583
rect 1568 582 1569 586
rect 1567 580 1569 582
rect 518 557 520 560
rect 562 558 564 560
rect 519 553 520 557
rect 563 554 564 558
rect 588 557 590 561
rect 634 558 636 560
rect 502 549 504 551
rect 518 549 520 553
rect 534 549 536 551
rect 557 549 559 551
rect 562 549 564 554
rect 589 553 590 557
rect 635 554 636 558
rect 1451 557 1453 560
rect 1495 558 1497 560
rect 588 549 590 553
rect 609 549 611 551
rect 629 549 631 551
rect 634 549 636 554
rect 1452 553 1453 557
rect 1496 554 1497 558
rect 1521 557 1523 561
rect 1567 558 1569 560
rect 652 549 654 551
rect 1435 549 1437 551
rect 1451 549 1453 553
rect 1467 549 1469 551
rect 1490 549 1492 551
rect 1495 549 1497 554
rect 1522 553 1523 557
rect 1568 554 1569 558
rect 1521 549 1523 553
rect 1542 549 1544 551
rect 1562 549 1564 551
rect 1567 549 1569 554
rect 1585 549 1587 551
rect 702 546 704 549
rect 707 546 709 549
rect 783 546 785 549
rect 788 546 790 549
rect 873 546 875 549
rect 878 546 880 549
rect 502 531 504 545
rect 518 543 520 545
rect 518 531 520 533
rect 534 531 536 545
rect 557 540 559 545
rect 562 543 564 545
rect 588 543 590 545
rect 553 536 559 540
rect 557 531 559 536
rect 562 531 564 533
rect 588 531 590 533
rect 609 531 611 545
rect 629 540 631 545
rect 634 543 636 545
rect 625 536 631 540
rect 629 531 631 536
rect 634 531 636 533
rect 652 531 654 545
rect 1635 546 1637 549
rect 1640 546 1642 549
rect 1716 546 1718 549
rect 1721 546 1723 549
rect 1806 546 1808 549
rect 1811 546 1813 549
rect 702 530 704 542
rect 707 540 709 542
rect 707 530 709 532
rect 783 530 785 542
rect 788 540 790 542
rect 788 530 790 532
rect 873 530 875 542
rect 878 540 880 542
rect 878 530 880 532
rect 1435 531 1437 545
rect 1451 543 1453 545
rect 1451 531 1453 533
rect 1467 531 1469 545
rect 1490 540 1492 545
rect 1495 543 1497 545
rect 1521 543 1523 545
rect 1486 536 1492 540
rect 1490 531 1492 536
rect 1495 531 1497 533
rect 1521 531 1523 533
rect 1542 531 1544 545
rect 1562 540 1564 545
rect 1567 543 1569 545
rect 1558 536 1564 540
rect 1562 531 1564 536
rect 1567 531 1569 533
rect 1585 531 1587 545
rect 502 521 504 523
rect 518 520 520 523
rect 534 521 536 523
rect 557 521 559 523
rect 562 520 564 523
rect 588 520 590 523
rect 609 520 611 523
rect 629 521 631 523
rect 634 520 636 523
rect 652 521 654 523
rect 1635 530 1637 542
rect 1640 540 1642 542
rect 1640 530 1642 532
rect 1716 530 1718 542
rect 1721 540 1723 542
rect 1721 530 1723 532
rect 1806 530 1808 542
rect 1811 540 1813 542
rect 1811 530 1813 532
rect 702 520 704 522
rect 588 516 589 520
rect 707 517 709 522
rect 783 520 785 522
rect 788 517 790 522
rect 873 520 875 522
rect 878 517 880 522
rect 1435 521 1437 523
rect 518 513 520 516
rect 562 513 564 516
rect 588 513 590 516
rect 634 513 636 516
rect 1451 520 1453 523
rect 1467 521 1469 523
rect 1490 521 1492 523
rect 1495 520 1497 523
rect 1521 520 1523 523
rect 1542 520 1544 523
rect 1562 521 1564 523
rect 1567 520 1569 523
rect 1585 521 1587 523
rect 1635 520 1637 522
rect 1521 516 1522 520
rect 1640 517 1642 522
rect 1716 520 1718 522
rect 1721 517 1723 522
rect 1806 520 1808 522
rect 1811 517 1813 522
rect 1451 513 1453 516
rect 1495 513 1497 516
rect 1521 513 1523 516
rect 1567 513 1569 516
rect 518 492 520 495
rect 562 492 564 495
rect 588 492 590 495
rect 634 492 636 495
rect 702 492 704 496
rect 730 498 732 500
rect 707 492 709 495
rect 588 488 589 492
rect 502 485 504 487
rect 518 485 520 488
rect 534 485 536 487
rect 557 485 559 487
rect 562 485 564 488
rect 588 485 590 488
rect 609 485 611 488
rect 629 485 631 487
rect 634 485 636 488
rect 652 485 654 487
rect 1451 492 1453 495
rect 1495 492 1497 495
rect 1521 492 1523 495
rect 1567 492 1569 495
rect 1635 492 1637 496
rect 1663 498 1665 500
rect 1640 492 1642 495
rect 702 481 704 484
rect 707 482 709 484
rect 703 477 704 481
rect 502 463 504 477
rect 518 475 520 477
rect 518 463 520 465
rect 534 463 536 477
rect 557 472 559 477
rect 562 475 564 477
rect 588 475 590 477
rect 553 468 559 472
rect 557 463 559 468
rect 562 463 564 465
rect 588 463 590 465
rect 609 463 611 477
rect 629 472 631 477
rect 634 475 636 477
rect 625 468 631 472
rect 629 463 631 468
rect 634 463 636 465
rect 652 463 654 477
rect 702 472 704 477
rect 707 472 709 474
rect 730 468 732 490
rect 1521 488 1522 492
rect 1435 485 1437 487
rect 1451 485 1453 488
rect 1467 485 1469 487
rect 1490 485 1492 487
rect 1495 485 1497 488
rect 1521 485 1523 488
rect 1542 485 1544 488
rect 1562 485 1564 487
rect 1567 485 1569 488
rect 1585 485 1587 487
rect 1635 481 1637 484
rect 1640 482 1642 484
rect 1636 477 1637 481
rect 702 466 704 468
rect 707 463 709 468
rect 730 462 732 464
rect 1435 463 1437 477
rect 1451 475 1453 477
rect 1451 463 1453 465
rect 1467 463 1469 477
rect 1490 472 1492 477
rect 1495 475 1497 477
rect 1521 475 1523 477
rect 1486 468 1492 472
rect 1490 463 1492 468
rect 1495 463 1497 465
rect 1521 463 1523 465
rect 1542 463 1544 477
rect 1562 472 1564 477
rect 1567 475 1569 477
rect 1558 468 1564 472
rect 1562 463 1564 468
rect 1567 463 1569 465
rect 1585 463 1587 477
rect 1635 472 1637 477
rect 1640 472 1642 474
rect 1663 468 1665 490
rect 1635 466 1637 468
rect 1640 463 1642 468
rect 1663 462 1665 464
rect 502 457 504 459
rect 518 455 520 459
rect 534 457 536 459
rect 557 457 559 459
rect 519 451 520 455
rect 562 454 564 459
rect 588 455 590 459
rect 609 457 611 459
rect 629 457 631 459
rect 518 448 520 451
rect 563 450 564 454
rect 589 451 590 455
rect 634 454 636 459
rect 652 457 654 459
rect 1435 457 1437 459
rect 1451 455 1453 459
rect 1467 457 1469 459
rect 1490 457 1492 459
rect 562 448 564 450
rect 588 447 590 451
rect 635 450 636 454
rect 1452 451 1453 455
rect 1495 454 1497 459
rect 1521 455 1523 459
rect 1542 457 1544 459
rect 1562 457 1564 459
rect 634 448 636 450
rect 1451 448 1453 451
rect 1496 450 1497 454
rect 1522 451 1523 455
rect 1567 454 1569 459
rect 1585 457 1587 459
rect 1495 448 1497 450
rect 1521 447 1523 451
rect 1568 450 1569 454
rect 1567 448 1569 450
rect 25 430 27 432
rect 30 430 32 433
rect 46 430 48 432
rect 62 430 64 432
rect 67 430 69 433
rect 88 430 90 433
rect 104 430 106 433
rect 120 430 122 432
rect 125 430 127 433
rect 141 430 143 432
rect 157 430 159 432
rect 162 430 164 433
rect 178 430 180 432
rect 194 430 196 432
rect 199 430 201 433
rect 220 430 222 433
rect 236 430 238 433
rect 252 430 254 432
rect 257 430 259 433
rect 273 430 275 432
rect 289 430 291 432
rect 294 430 296 433
rect 310 430 312 432
rect 326 430 328 432
rect 331 430 333 433
rect 352 430 354 433
rect 368 430 370 433
rect 384 430 386 432
rect 389 430 391 433
rect 405 430 407 432
rect 958 430 960 432
rect 963 430 965 433
rect 979 430 981 432
rect 995 430 997 432
rect 1000 430 1002 433
rect 1021 430 1023 433
rect 1037 430 1039 433
rect 1053 430 1055 432
rect 1058 430 1060 433
rect 1074 430 1076 432
rect 1090 430 1092 432
rect 1095 430 1097 433
rect 1111 430 1113 432
rect 1127 430 1129 432
rect 1132 430 1134 433
rect 1153 430 1155 433
rect 1169 430 1171 433
rect 1185 430 1187 432
rect 1190 430 1192 433
rect 1206 430 1208 432
rect 1222 430 1224 432
rect 1227 430 1229 433
rect 1243 430 1245 432
rect 1259 430 1261 432
rect 1264 430 1266 433
rect 1285 430 1287 433
rect 1301 430 1303 433
rect 1317 430 1319 432
rect 1322 430 1324 433
rect 1338 430 1340 432
rect 518 425 520 428
rect 562 426 564 428
rect 25 417 27 422
rect 30 420 32 422
rect 25 403 27 413
rect 30 403 32 410
rect 46 403 48 422
rect 62 413 64 422
rect 67 420 69 422
rect 88 420 90 422
rect 104 419 106 422
rect 62 403 64 406
rect 67 403 69 405
rect 88 403 90 405
rect 104 403 106 415
rect 120 413 122 422
rect 125 420 127 422
rect 120 403 122 406
rect 125 403 127 405
rect 141 403 143 422
rect 157 419 159 422
rect 162 420 164 422
rect 157 403 159 415
rect 162 403 164 410
rect 178 403 180 422
rect 194 413 196 422
rect 199 420 201 422
rect 220 420 222 422
rect 236 419 238 422
rect 194 403 196 406
rect 199 403 201 405
rect 220 403 222 405
rect 236 403 238 415
rect 252 413 254 422
rect 257 420 259 422
rect 252 403 254 406
rect 257 403 259 405
rect 273 403 275 422
rect 289 419 291 422
rect 294 420 296 422
rect 289 403 291 415
rect 294 403 296 410
rect 310 403 312 422
rect 326 413 328 422
rect 331 420 333 422
rect 352 420 354 422
rect 368 419 370 422
rect 326 403 328 406
rect 331 403 333 405
rect 352 403 354 405
rect 368 403 370 415
rect 384 413 386 422
rect 389 420 391 422
rect 405 414 407 422
rect 519 421 520 425
rect 563 422 564 426
rect 588 425 590 429
rect 634 426 636 428
rect 502 417 504 419
rect 518 417 520 421
rect 534 417 536 419
rect 557 417 559 419
rect 562 417 564 422
rect 589 421 590 425
rect 635 422 636 426
rect 779 425 781 428
rect 823 426 825 428
rect 588 417 590 421
rect 609 417 611 419
rect 629 417 631 419
rect 634 417 636 422
rect 780 421 781 425
rect 824 422 825 426
rect 849 425 851 429
rect 895 426 897 428
rect 652 417 654 419
rect 736 417 738 420
rect 754 417 756 420
rect 779 417 781 421
rect 795 417 797 419
rect 818 417 820 419
rect 823 417 825 422
rect 850 421 851 425
rect 896 422 897 426
rect 1451 425 1453 428
rect 1495 426 1497 428
rect 849 417 851 421
rect 870 417 872 419
rect 890 417 892 419
rect 895 417 897 422
rect 913 417 915 419
rect 958 417 960 422
rect 963 420 965 422
rect 384 403 386 406
rect 389 403 391 405
rect 405 403 407 410
rect 502 399 504 413
rect 518 411 520 413
rect 518 399 520 401
rect 534 399 536 413
rect 557 408 559 413
rect 562 411 564 413
rect 588 411 590 413
rect 553 404 559 408
rect 557 399 559 404
rect 562 399 564 401
rect 588 399 590 401
rect 609 399 611 413
rect 629 408 631 413
rect 634 411 636 413
rect 625 404 631 408
rect 629 399 631 404
rect 634 399 636 401
rect 652 399 654 413
rect 702 410 704 413
rect 707 410 709 413
rect 736 408 738 413
rect 25 397 27 399
rect 30 396 32 399
rect 46 397 48 399
rect 62 397 64 399
rect 67 394 69 399
rect 88 394 90 399
rect 104 397 106 399
rect 120 397 122 399
rect 125 394 127 399
rect 141 397 143 399
rect 157 397 159 399
rect 162 396 164 399
rect 178 397 180 399
rect 194 397 196 399
rect 199 394 201 399
rect 220 394 222 399
rect 236 397 238 399
rect 252 397 254 399
rect 257 394 259 399
rect 273 397 275 399
rect 289 397 291 399
rect 294 396 296 399
rect 310 397 312 399
rect 326 397 328 399
rect 331 394 333 399
rect 352 394 354 399
rect 368 397 370 399
rect 384 397 386 399
rect 389 394 391 399
rect 405 397 407 399
rect 702 394 704 406
rect 707 404 709 406
rect 736 399 738 404
rect 754 399 756 413
rect 779 411 781 413
rect 779 399 781 401
rect 795 399 797 413
rect 818 408 820 413
rect 823 411 825 413
rect 849 411 851 413
rect 814 404 820 408
rect 818 399 820 404
rect 823 399 825 401
rect 849 399 851 401
rect 870 399 872 413
rect 890 408 892 413
rect 895 411 897 413
rect 886 404 892 408
rect 890 399 892 404
rect 895 399 897 401
rect 913 399 915 413
rect 958 403 960 413
rect 963 403 965 410
rect 979 403 981 422
rect 995 413 997 422
rect 1000 420 1002 422
rect 1021 420 1023 422
rect 1037 419 1039 422
rect 995 403 997 406
rect 1000 403 1002 405
rect 1021 403 1023 405
rect 1037 403 1039 415
rect 1053 413 1055 422
rect 1058 420 1060 422
rect 1053 403 1055 406
rect 1058 403 1060 405
rect 1074 403 1076 422
rect 1090 419 1092 422
rect 1095 420 1097 422
rect 1090 403 1092 415
rect 1095 403 1097 410
rect 1111 403 1113 422
rect 1127 413 1129 422
rect 1132 420 1134 422
rect 1153 420 1155 422
rect 1169 419 1171 422
rect 1127 403 1129 406
rect 1132 403 1134 405
rect 1153 403 1155 405
rect 1169 403 1171 415
rect 1185 413 1187 422
rect 1190 420 1192 422
rect 1185 403 1187 406
rect 1190 403 1192 405
rect 1206 403 1208 422
rect 1222 419 1224 422
rect 1227 420 1229 422
rect 1222 403 1224 415
rect 1227 403 1229 410
rect 1243 403 1245 422
rect 1259 413 1261 422
rect 1264 420 1266 422
rect 1285 420 1287 422
rect 1301 419 1303 422
rect 1259 403 1261 406
rect 1264 403 1266 405
rect 1285 403 1287 405
rect 1301 403 1303 415
rect 1317 413 1319 422
rect 1322 420 1324 422
rect 1338 414 1340 422
rect 1452 421 1453 425
rect 1496 422 1497 426
rect 1521 425 1523 429
rect 1567 426 1569 428
rect 1435 417 1437 419
rect 1451 417 1453 421
rect 1467 417 1469 419
rect 1490 417 1492 419
rect 1495 417 1497 422
rect 1522 421 1523 425
rect 1568 422 1569 426
rect 1712 425 1714 428
rect 1756 426 1758 428
rect 1521 417 1523 421
rect 1542 417 1544 419
rect 1562 417 1564 419
rect 1567 417 1569 422
rect 1713 421 1714 425
rect 1757 422 1758 426
rect 1782 425 1784 429
rect 1828 426 1830 428
rect 1585 417 1587 419
rect 1669 417 1671 420
rect 1687 417 1689 420
rect 1712 417 1714 421
rect 1728 417 1730 419
rect 1751 417 1753 419
rect 1756 417 1758 422
rect 1783 421 1784 425
rect 1829 422 1830 426
rect 1782 417 1784 421
rect 1803 417 1805 419
rect 1823 417 1825 419
rect 1828 417 1830 422
rect 1846 417 1848 419
rect 1317 403 1319 406
rect 1322 403 1324 405
rect 1338 403 1340 410
rect 1435 399 1437 413
rect 1451 411 1453 413
rect 1451 399 1453 401
rect 1467 399 1469 413
rect 1490 408 1492 413
rect 1495 411 1497 413
rect 1521 411 1523 413
rect 1486 404 1492 408
rect 1490 399 1492 404
rect 1495 399 1497 401
rect 1521 399 1523 401
rect 1542 399 1544 413
rect 1562 408 1564 413
rect 1567 411 1569 413
rect 1558 404 1564 408
rect 1562 399 1564 404
rect 1567 399 1569 401
rect 1585 399 1587 413
rect 1635 410 1637 413
rect 1640 410 1642 413
rect 1669 408 1671 413
rect 707 394 709 396
rect 502 389 504 391
rect 518 388 520 391
rect 534 389 536 391
rect 557 389 559 391
rect 562 388 564 391
rect 588 388 590 391
rect 609 388 611 391
rect 629 389 631 391
rect 634 388 636 391
rect 652 389 654 391
rect 588 384 589 388
rect 958 397 960 399
rect 963 396 965 399
rect 979 397 981 399
rect 995 397 997 399
rect 1000 394 1002 399
rect 1021 394 1023 399
rect 1037 397 1039 399
rect 1053 397 1055 399
rect 1058 394 1060 399
rect 1074 397 1076 399
rect 1090 397 1092 399
rect 736 388 738 391
rect 754 388 756 391
rect 779 388 781 391
rect 795 389 797 391
rect 818 389 820 391
rect 823 388 825 391
rect 849 388 851 391
rect 870 388 872 391
rect 890 389 892 391
rect 895 388 897 391
rect 913 389 915 391
rect 1095 396 1097 399
rect 1111 397 1113 399
rect 1127 397 1129 399
rect 1132 394 1134 399
rect 1153 394 1155 399
rect 1169 397 1171 399
rect 1185 397 1187 399
rect 1190 394 1192 399
rect 1206 397 1208 399
rect 1222 397 1224 399
rect 1227 396 1229 399
rect 1243 397 1245 399
rect 1259 397 1261 399
rect 1264 394 1266 399
rect 1285 394 1287 399
rect 1301 397 1303 399
rect 1317 397 1319 399
rect 1322 394 1324 399
rect 1338 397 1340 399
rect 1635 394 1637 406
rect 1640 404 1642 406
rect 1669 399 1671 404
rect 1687 399 1689 413
rect 1712 411 1714 413
rect 1712 399 1714 401
rect 1728 399 1730 413
rect 1751 408 1753 413
rect 1756 411 1758 413
rect 1782 411 1784 413
rect 1747 404 1753 408
rect 1751 399 1753 404
rect 1756 399 1758 401
rect 1782 399 1784 401
rect 1803 399 1805 413
rect 1823 408 1825 413
rect 1828 411 1830 413
rect 1819 404 1825 408
rect 1823 399 1825 404
rect 1828 399 1830 401
rect 1846 399 1848 413
rect 1640 394 1642 396
rect 1435 389 1437 391
rect 1451 388 1453 391
rect 1467 389 1469 391
rect 1490 389 1492 391
rect 1495 388 1497 391
rect 1521 388 1523 391
rect 1542 388 1544 391
rect 1562 389 1564 391
rect 1567 388 1569 391
rect 1585 389 1587 391
rect 702 384 704 386
rect 518 381 520 384
rect 562 381 564 384
rect 588 381 590 384
rect 634 381 636 384
rect 707 381 709 386
rect 849 384 850 388
rect 779 381 781 384
rect 823 381 825 384
rect 849 381 851 384
rect 895 381 897 384
rect 1521 384 1522 388
rect 1669 388 1671 391
rect 1687 388 1689 391
rect 1712 388 1714 391
rect 1728 389 1730 391
rect 1751 389 1753 391
rect 1756 388 1758 391
rect 1782 388 1784 391
rect 1803 388 1805 391
rect 1823 389 1825 391
rect 1828 388 1830 391
rect 1846 389 1848 391
rect 1635 384 1637 386
rect 1451 381 1453 384
rect 1495 381 1497 384
rect 1521 381 1523 384
rect 1567 381 1569 384
rect 1640 381 1642 386
rect 1782 384 1783 388
rect 1712 381 1714 384
rect 1756 381 1758 384
rect 1782 381 1784 384
rect 1828 381 1830 384
rect 140 359 142 362
rect 164 359 166 362
rect 1073 359 1075 362
rect 1097 359 1099 362
rect 922 357 925 359
rect 929 357 932 359
rect 140 353 142 355
rect 164 353 166 355
rect 1855 357 1858 359
rect 1862 357 1865 359
rect 1073 353 1075 355
rect 1097 353 1099 355
rect 160 348 162 350
rect 1093 348 1095 350
rect 160 341 162 344
rect 1093 341 1095 344
rect 149 330 151 332
rect 155 330 174 332
rect 1082 330 1084 332
rect 1088 330 1107 332
rect 140 325 142 327
rect 164 325 166 327
rect 1073 325 1075 327
rect 1097 325 1099 327
rect 140 318 142 321
rect 164 318 166 321
rect 796 320 798 322
rect 801 320 803 323
rect 817 320 819 322
rect 833 320 835 322
rect 838 320 840 323
rect 859 320 861 323
rect 875 320 877 323
rect 891 320 893 322
rect 896 320 898 323
rect 912 320 914 322
rect 1073 318 1075 321
rect 1097 318 1099 321
rect 1729 320 1731 322
rect 1734 320 1736 323
rect 1750 320 1752 322
rect 1766 320 1768 322
rect 1771 320 1773 323
rect 1792 320 1794 323
rect 1808 320 1810 323
rect 1824 320 1826 322
rect 1829 320 1831 323
rect 1845 320 1847 322
rect 796 307 798 312
rect 801 310 803 312
rect 796 293 798 303
rect 801 293 803 300
rect 817 293 819 312
rect 833 303 835 312
rect 838 310 840 312
rect 859 310 861 312
rect 875 309 877 312
rect 833 293 835 296
rect 838 293 840 295
rect 859 293 861 295
rect 875 293 877 305
rect 891 303 893 312
rect 896 310 898 312
rect 891 293 893 296
rect 896 293 898 295
rect 912 293 914 312
rect 1729 307 1731 312
rect 1734 310 1736 312
rect 1729 293 1731 303
rect 1734 293 1736 300
rect 1750 293 1752 312
rect 1766 303 1768 312
rect 1771 310 1773 312
rect 1792 310 1794 312
rect 1808 309 1810 312
rect 1766 293 1768 296
rect 1771 293 1773 295
rect 1792 293 1794 295
rect 1808 293 1810 305
rect 1824 303 1826 312
rect 1829 310 1831 312
rect 1824 293 1826 296
rect 1829 293 1831 295
rect 1845 293 1847 312
rect 25 290 27 292
rect 30 290 32 293
rect 46 290 48 292
rect 62 290 64 292
rect 67 290 69 293
rect 88 290 90 293
rect 104 290 106 293
rect 120 290 122 292
rect 125 290 127 293
rect 141 290 143 292
rect 157 290 159 292
rect 162 290 164 293
rect 178 290 180 292
rect 194 290 196 292
rect 199 290 201 293
rect 220 290 222 293
rect 236 290 238 293
rect 252 290 254 292
rect 257 290 259 293
rect 273 290 275 292
rect 289 290 291 292
rect 294 290 296 293
rect 310 290 312 292
rect 326 290 328 292
rect 331 290 333 293
rect 352 290 354 293
rect 368 290 370 293
rect 384 290 386 292
rect 389 290 391 293
rect 405 290 407 292
rect 958 290 960 292
rect 963 290 965 293
rect 979 290 981 292
rect 995 290 997 292
rect 1000 290 1002 293
rect 1021 290 1023 293
rect 1037 290 1039 293
rect 1053 290 1055 292
rect 1058 290 1060 293
rect 1074 290 1076 292
rect 1090 290 1092 292
rect 1095 290 1097 293
rect 1111 290 1113 292
rect 1127 290 1129 292
rect 1132 290 1134 293
rect 1153 290 1155 293
rect 1169 290 1171 293
rect 1185 290 1187 292
rect 1190 290 1192 293
rect 1206 290 1208 292
rect 1222 290 1224 292
rect 1227 290 1229 293
rect 1243 290 1245 292
rect 1259 290 1261 292
rect 1264 290 1266 293
rect 1285 290 1287 293
rect 1301 290 1303 293
rect 1317 290 1319 292
rect 1322 290 1324 293
rect 1338 290 1340 292
rect 796 287 798 289
rect 801 286 803 289
rect 817 287 819 289
rect 833 287 835 289
rect 838 284 840 289
rect 859 284 861 289
rect 875 287 877 289
rect 891 287 893 289
rect 896 284 898 289
rect 912 287 914 289
rect 25 277 27 282
rect 30 280 32 282
rect 25 263 27 273
rect 30 263 32 270
rect 46 263 48 282
rect 62 273 64 282
rect 67 280 69 282
rect 88 280 90 282
rect 104 279 106 282
rect 62 263 64 266
rect 67 263 69 265
rect 88 263 90 265
rect 104 263 106 275
rect 120 273 122 282
rect 125 280 127 282
rect 120 263 122 266
rect 125 263 127 265
rect 141 263 143 282
rect 157 279 159 282
rect 162 280 164 282
rect 157 263 159 275
rect 162 263 164 270
rect 178 263 180 282
rect 194 273 196 282
rect 199 280 201 282
rect 220 280 222 282
rect 236 279 238 282
rect 194 263 196 266
rect 199 263 201 265
rect 220 263 222 265
rect 236 263 238 275
rect 252 273 254 282
rect 257 280 259 282
rect 252 263 254 266
rect 257 263 259 265
rect 273 263 275 282
rect 289 279 291 282
rect 294 280 296 282
rect 289 263 291 275
rect 294 263 296 270
rect 310 263 312 282
rect 326 273 328 282
rect 331 280 333 282
rect 352 280 354 282
rect 368 279 370 282
rect 326 263 328 266
rect 331 263 333 265
rect 352 263 354 265
rect 368 263 370 275
rect 384 273 386 282
rect 389 280 391 282
rect 405 274 407 282
rect 1729 287 1731 289
rect 1734 286 1736 289
rect 1750 287 1752 289
rect 1766 287 1768 289
rect 1771 284 1773 289
rect 1792 284 1794 289
rect 1808 287 1810 289
rect 1824 287 1826 289
rect 1829 284 1831 289
rect 1845 287 1847 289
rect 958 277 960 282
rect 963 280 965 282
rect 384 263 386 266
rect 389 263 391 265
rect 405 263 407 270
rect 958 263 960 273
rect 963 263 965 270
rect 979 263 981 282
rect 995 273 997 282
rect 1000 280 1002 282
rect 1021 280 1023 282
rect 1037 279 1039 282
rect 995 263 997 266
rect 1000 263 1002 265
rect 1021 263 1023 265
rect 1037 263 1039 275
rect 1053 273 1055 282
rect 1058 280 1060 282
rect 1053 263 1055 266
rect 1058 263 1060 265
rect 1074 263 1076 282
rect 1090 279 1092 282
rect 1095 280 1097 282
rect 1090 263 1092 275
rect 1095 263 1097 270
rect 1111 263 1113 282
rect 1127 273 1129 282
rect 1132 280 1134 282
rect 1153 280 1155 282
rect 1169 279 1171 282
rect 1127 263 1129 266
rect 1132 263 1134 265
rect 1153 263 1155 265
rect 1169 263 1171 275
rect 1185 273 1187 282
rect 1190 280 1192 282
rect 1185 263 1187 266
rect 1190 263 1192 265
rect 1206 263 1208 282
rect 1222 279 1224 282
rect 1227 280 1229 282
rect 1222 263 1224 275
rect 1227 263 1229 270
rect 1243 263 1245 282
rect 1259 273 1261 282
rect 1264 280 1266 282
rect 1285 280 1287 282
rect 1301 279 1303 282
rect 1259 263 1261 266
rect 1264 263 1266 265
rect 1285 263 1287 265
rect 1301 263 1303 275
rect 1317 273 1319 282
rect 1322 280 1324 282
rect 1338 274 1340 282
rect 1317 263 1319 266
rect 1322 263 1324 265
rect 1338 263 1340 270
rect 25 257 27 259
rect 30 256 32 259
rect 46 257 48 259
rect 62 257 64 259
rect 67 254 69 259
rect 88 254 90 259
rect 104 257 106 259
rect 120 257 122 259
rect 125 254 127 259
rect 141 257 143 259
rect 157 257 159 259
rect 162 256 164 259
rect 178 257 180 259
rect 194 257 196 259
rect 199 254 201 259
rect 220 254 222 259
rect 236 257 238 259
rect 252 257 254 259
rect 257 254 259 259
rect 273 257 275 259
rect 289 257 291 259
rect 294 256 296 259
rect 310 257 312 259
rect 326 257 328 259
rect 331 254 333 259
rect 352 254 354 259
rect 368 257 370 259
rect 384 257 386 259
rect 389 254 391 259
rect 405 257 407 259
rect 958 257 960 259
rect 963 256 965 259
rect 979 257 981 259
rect 995 257 997 259
rect 1000 254 1002 259
rect 1021 254 1023 259
rect 1037 257 1039 259
rect 1053 257 1055 259
rect 1058 254 1060 259
rect 1074 257 1076 259
rect 1090 257 1092 259
rect 1095 256 1097 259
rect 1111 257 1113 259
rect 1127 257 1129 259
rect 1132 254 1134 259
rect 1153 254 1155 259
rect 1169 257 1171 259
rect 1185 257 1187 259
rect 1190 254 1192 259
rect 1206 257 1208 259
rect 1222 257 1224 259
rect 1227 256 1229 259
rect 1243 257 1245 259
rect 1259 257 1261 259
rect 1264 254 1266 259
rect 1285 254 1287 259
rect 1301 257 1303 259
rect 1317 257 1319 259
rect 1322 254 1324 259
rect 1338 257 1340 259
rect 796 234 798 236
rect 801 234 803 237
rect 817 234 819 236
rect 833 234 835 236
rect 838 234 840 237
rect 859 234 861 237
rect 875 234 877 237
rect 891 234 893 236
rect 896 234 898 237
rect 912 234 914 236
rect 1729 234 1731 236
rect 1734 234 1736 237
rect 1750 234 1752 236
rect 1766 234 1768 236
rect 1771 234 1773 237
rect 1792 234 1794 237
rect 1808 234 1810 237
rect 1824 234 1826 236
rect 1829 234 1831 237
rect 1845 234 1847 236
rect 796 221 798 226
rect 801 224 803 226
rect 796 207 798 217
rect 801 207 803 214
rect 817 207 819 226
rect 833 217 835 226
rect 838 224 840 226
rect 859 224 861 226
rect 875 223 877 226
rect 833 207 835 210
rect 838 207 840 209
rect 859 207 861 209
rect 875 207 877 219
rect 891 217 893 226
rect 896 224 898 226
rect 891 207 893 210
rect 896 207 898 209
rect 912 207 914 226
rect 1729 221 1731 226
rect 1734 224 1736 226
rect 934 213 937 215
rect 941 213 944 215
rect 1729 207 1731 217
rect 1734 207 1736 214
rect 1750 207 1752 226
rect 1766 217 1768 226
rect 1771 224 1773 226
rect 1792 224 1794 226
rect 1808 223 1810 226
rect 1766 207 1768 210
rect 1771 207 1773 209
rect 1792 207 1794 209
rect 1808 207 1810 219
rect 1824 217 1826 226
rect 1829 224 1831 226
rect 1824 207 1826 210
rect 1829 207 1831 209
rect 1845 207 1847 226
rect 1867 213 1870 215
rect 1874 213 1877 215
rect 25 204 27 206
rect 30 204 32 207
rect 46 204 48 206
rect 62 204 64 206
rect 67 204 69 207
rect 88 204 90 207
rect 104 204 106 207
rect 120 204 122 206
rect 125 204 127 207
rect 141 204 143 206
rect 157 204 159 206
rect 162 204 164 207
rect 178 204 180 206
rect 194 204 196 206
rect 199 204 201 207
rect 220 204 222 207
rect 236 204 238 207
rect 252 204 254 206
rect 257 204 259 207
rect 273 204 275 206
rect 289 204 291 206
rect 294 204 296 207
rect 310 204 312 206
rect 326 204 328 206
rect 331 204 333 207
rect 352 204 354 207
rect 368 204 370 207
rect 384 204 386 206
rect 389 204 391 207
rect 405 204 407 206
rect 958 204 960 206
rect 963 204 965 207
rect 979 204 981 206
rect 995 204 997 206
rect 1000 204 1002 207
rect 1021 204 1023 207
rect 1037 204 1039 207
rect 1053 204 1055 206
rect 1058 204 1060 207
rect 1074 204 1076 206
rect 1090 204 1092 206
rect 1095 204 1097 207
rect 1111 204 1113 206
rect 1127 204 1129 206
rect 1132 204 1134 207
rect 1153 204 1155 207
rect 1169 204 1171 207
rect 1185 204 1187 206
rect 1190 204 1192 207
rect 1206 204 1208 206
rect 1222 204 1224 206
rect 1227 204 1229 207
rect 1243 204 1245 206
rect 1259 204 1261 206
rect 1264 204 1266 207
rect 1285 204 1287 207
rect 1301 204 1303 207
rect 1317 204 1319 206
rect 1322 204 1324 207
rect 1338 204 1340 206
rect 796 201 798 203
rect 801 200 803 203
rect 817 201 819 203
rect 833 201 835 203
rect 838 198 840 203
rect 859 198 861 203
rect 875 201 877 203
rect 891 201 893 203
rect 896 198 898 203
rect 912 201 914 203
rect 25 191 27 196
rect 30 194 32 196
rect 25 177 27 187
rect 30 177 32 184
rect 46 177 48 196
rect 62 187 64 196
rect 67 194 69 196
rect 88 194 90 196
rect 104 193 106 196
rect 62 177 64 180
rect 67 177 69 179
rect 88 177 90 179
rect 104 177 106 189
rect 120 187 122 196
rect 125 194 127 196
rect 120 177 122 180
rect 125 177 127 179
rect 141 177 143 196
rect 157 193 159 196
rect 162 194 164 196
rect 157 177 159 189
rect 162 177 164 184
rect 178 177 180 196
rect 194 187 196 196
rect 199 194 201 196
rect 220 194 222 196
rect 236 193 238 196
rect 194 177 196 180
rect 199 177 201 179
rect 220 177 222 179
rect 236 177 238 189
rect 252 187 254 196
rect 257 194 259 196
rect 252 177 254 180
rect 257 177 259 179
rect 273 177 275 196
rect 289 193 291 196
rect 294 194 296 196
rect 289 177 291 189
rect 294 177 296 184
rect 310 177 312 196
rect 326 187 328 196
rect 331 194 333 196
rect 352 194 354 196
rect 368 193 370 196
rect 326 177 328 180
rect 331 177 333 179
rect 352 177 354 179
rect 368 177 370 189
rect 384 187 386 196
rect 389 194 391 196
rect 405 188 407 196
rect 1729 201 1731 203
rect 1734 200 1736 203
rect 1750 201 1752 203
rect 1766 201 1768 203
rect 1771 198 1773 203
rect 1792 198 1794 203
rect 1808 201 1810 203
rect 1824 201 1826 203
rect 1829 198 1831 203
rect 1845 201 1847 203
rect 958 191 960 196
rect 963 194 965 196
rect 384 177 386 180
rect 389 177 391 179
rect 405 177 407 184
rect 958 177 960 187
rect 963 177 965 184
rect 979 177 981 196
rect 995 187 997 196
rect 1000 194 1002 196
rect 1021 194 1023 196
rect 1037 193 1039 196
rect 995 177 997 180
rect 1000 177 1002 179
rect 1021 177 1023 179
rect 1037 177 1039 189
rect 1053 187 1055 196
rect 1058 194 1060 196
rect 1053 177 1055 180
rect 1058 177 1060 179
rect 1074 177 1076 196
rect 1090 193 1092 196
rect 1095 194 1097 196
rect 1090 177 1092 189
rect 1095 177 1097 184
rect 1111 177 1113 196
rect 1127 187 1129 196
rect 1132 194 1134 196
rect 1153 194 1155 196
rect 1169 193 1171 196
rect 1127 177 1129 180
rect 1132 177 1134 179
rect 1153 177 1155 179
rect 1169 177 1171 189
rect 1185 187 1187 196
rect 1190 194 1192 196
rect 1185 177 1187 180
rect 1190 177 1192 179
rect 1206 177 1208 196
rect 1222 193 1224 196
rect 1227 194 1229 196
rect 1222 177 1224 189
rect 1227 177 1229 184
rect 1243 177 1245 196
rect 1259 187 1261 196
rect 1264 194 1266 196
rect 1285 194 1287 196
rect 1301 193 1303 196
rect 1259 177 1261 180
rect 1264 177 1266 179
rect 1285 177 1287 179
rect 1301 177 1303 189
rect 1317 187 1319 196
rect 1322 194 1324 196
rect 1338 188 1340 196
rect 1317 177 1319 180
rect 1322 177 1324 179
rect 1338 177 1340 184
rect 25 171 27 173
rect 30 170 32 173
rect 46 171 48 173
rect 62 171 64 173
rect 67 168 69 173
rect 88 168 90 173
rect 104 171 106 173
rect 120 171 122 173
rect 125 168 127 173
rect 141 171 143 173
rect 157 171 159 173
rect 162 170 164 173
rect 178 171 180 173
rect 194 171 196 173
rect 199 168 201 173
rect 220 168 222 173
rect 236 171 238 173
rect 252 171 254 173
rect 257 168 259 173
rect 273 171 275 173
rect 289 171 291 173
rect 294 170 296 173
rect 310 171 312 173
rect 326 171 328 173
rect 331 168 333 173
rect 352 168 354 173
rect 368 171 370 173
rect 384 171 386 173
rect 389 168 391 173
rect 405 171 407 173
rect 958 171 960 173
rect 963 170 965 173
rect 979 171 981 173
rect 995 171 997 173
rect 1000 168 1002 173
rect 1021 168 1023 173
rect 1037 171 1039 173
rect 1053 171 1055 173
rect 1058 168 1060 173
rect 1074 171 1076 173
rect 1090 171 1092 173
rect 1095 170 1097 173
rect 1111 171 1113 173
rect 1127 171 1129 173
rect 1132 168 1134 173
rect 1153 168 1155 173
rect 1169 171 1171 173
rect 1185 171 1187 173
rect 1190 168 1192 173
rect 1206 171 1208 173
rect 1222 171 1224 173
rect 1227 170 1229 173
rect 1243 171 1245 173
rect 1259 171 1261 173
rect 1264 168 1266 173
rect 1285 168 1287 173
rect 1301 171 1303 173
rect 1317 171 1319 173
rect 1322 168 1324 173
rect 1338 171 1340 173
rect 257 133 259 136
rect 281 133 283 136
rect 1190 133 1192 136
rect 1214 133 1216 136
rect 257 127 259 129
rect 281 127 283 129
rect 1190 127 1192 129
rect 1214 127 1216 129
rect 277 122 279 124
rect 1210 122 1212 124
rect 277 115 279 118
rect 1210 115 1212 118
rect 266 104 268 106
rect 272 104 291 106
rect 1199 104 1201 106
rect 1205 104 1224 106
rect 257 99 259 101
rect 281 99 283 101
rect 1190 99 1192 101
rect 1214 99 1216 101
rect 257 92 259 95
rect 281 92 283 95
rect 1190 92 1192 95
rect 1214 92 1216 95
rect 25 64 27 66
rect 30 64 32 67
rect 46 64 48 66
rect 62 64 64 66
rect 67 64 69 67
rect 88 64 90 67
rect 104 64 106 67
rect 120 64 122 66
rect 125 64 127 67
rect 141 64 143 66
rect 157 64 159 66
rect 162 64 164 67
rect 178 64 180 66
rect 194 64 196 66
rect 199 64 201 67
rect 220 64 222 67
rect 236 64 238 67
rect 252 64 254 66
rect 257 64 259 67
rect 273 64 275 66
rect 289 64 291 66
rect 294 64 296 67
rect 310 64 312 66
rect 326 64 328 66
rect 331 64 333 67
rect 352 64 354 67
rect 368 64 370 67
rect 384 64 386 66
rect 389 64 391 67
rect 405 64 407 66
rect 958 64 960 66
rect 963 64 965 67
rect 979 64 981 66
rect 995 64 997 66
rect 1000 64 1002 67
rect 1021 64 1023 67
rect 1037 64 1039 67
rect 1053 64 1055 66
rect 1058 64 1060 67
rect 1074 64 1076 66
rect 1090 64 1092 66
rect 1095 64 1097 67
rect 1111 64 1113 66
rect 1127 64 1129 66
rect 1132 64 1134 67
rect 1153 64 1155 67
rect 1169 64 1171 67
rect 1185 64 1187 66
rect 1190 64 1192 67
rect 1206 64 1208 66
rect 1222 64 1224 66
rect 1227 64 1229 67
rect 1243 64 1245 66
rect 1259 64 1261 66
rect 1264 64 1266 67
rect 1285 64 1287 67
rect 1301 64 1303 67
rect 1317 64 1319 66
rect 1322 64 1324 67
rect 1338 64 1340 66
rect 25 51 27 56
rect 30 54 32 56
rect 25 37 27 47
rect 30 37 32 44
rect 46 37 48 56
rect 62 47 64 56
rect 67 54 69 56
rect 88 54 90 56
rect 104 53 106 56
rect 62 37 64 40
rect 67 37 69 39
rect 88 37 90 39
rect 104 37 106 49
rect 120 47 122 56
rect 125 54 127 56
rect 120 37 122 40
rect 125 37 127 39
rect 141 37 143 56
rect 157 53 159 56
rect 162 54 164 56
rect 157 37 159 49
rect 162 37 164 44
rect 178 37 180 56
rect 194 47 196 56
rect 199 54 201 56
rect 220 54 222 56
rect 236 53 238 56
rect 194 37 196 40
rect 199 37 201 39
rect 220 37 222 39
rect 236 37 238 49
rect 252 47 254 56
rect 257 54 259 56
rect 252 37 254 40
rect 257 37 259 39
rect 273 37 275 56
rect 289 53 291 56
rect 294 54 296 56
rect 289 37 291 49
rect 294 37 296 44
rect 310 37 312 56
rect 326 47 328 56
rect 331 54 333 56
rect 352 54 354 56
rect 368 53 370 56
rect 326 37 328 40
rect 331 37 333 39
rect 352 37 354 39
rect 368 37 370 49
rect 384 47 386 56
rect 389 54 391 56
rect 405 48 407 56
rect 958 51 960 56
rect 963 54 965 56
rect 384 37 386 40
rect 389 37 391 39
rect 405 37 407 44
rect 958 37 960 47
rect 963 37 965 44
rect 979 37 981 56
rect 995 47 997 56
rect 1000 54 1002 56
rect 1021 54 1023 56
rect 1037 53 1039 56
rect 995 37 997 40
rect 1000 37 1002 39
rect 1021 37 1023 39
rect 1037 37 1039 49
rect 1053 47 1055 56
rect 1058 54 1060 56
rect 1053 37 1055 40
rect 1058 37 1060 39
rect 1074 37 1076 56
rect 1090 53 1092 56
rect 1095 54 1097 56
rect 1090 37 1092 49
rect 1095 37 1097 44
rect 1111 37 1113 56
rect 1127 47 1129 56
rect 1132 54 1134 56
rect 1153 54 1155 56
rect 1169 53 1171 56
rect 1127 37 1129 40
rect 1132 37 1134 39
rect 1153 37 1155 39
rect 1169 37 1171 49
rect 1185 47 1187 56
rect 1190 54 1192 56
rect 1185 37 1187 40
rect 1190 37 1192 39
rect 1206 37 1208 56
rect 1222 53 1224 56
rect 1227 54 1229 56
rect 1222 37 1224 49
rect 1227 37 1229 44
rect 1243 37 1245 56
rect 1259 47 1261 56
rect 1264 54 1266 56
rect 1285 54 1287 56
rect 1301 53 1303 56
rect 1259 37 1261 40
rect 1264 37 1266 39
rect 1285 37 1287 39
rect 1301 37 1303 49
rect 1317 47 1319 56
rect 1322 54 1324 56
rect 1338 48 1340 56
rect 1317 37 1319 40
rect 1322 37 1324 39
rect 1338 37 1340 44
rect 25 31 27 33
rect 30 30 32 33
rect 46 31 48 33
rect 62 31 64 33
rect 67 28 69 33
rect 88 28 90 33
rect 104 31 106 33
rect 120 31 122 33
rect 125 28 127 33
rect 141 31 143 33
rect 157 31 159 33
rect 162 30 164 33
rect 178 31 180 33
rect 194 31 196 33
rect 199 28 201 33
rect 220 28 222 33
rect 236 31 238 33
rect 252 31 254 33
rect 257 28 259 33
rect 273 31 275 33
rect 289 31 291 33
rect 294 30 296 33
rect 310 31 312 33
rect 326 31 328 33
rect 331 28 333 33
rect 352 28 354 33
rect 368 31 370 33
rect 384 31 386 33
rect 389 28 391 33
rect 405 31 407 33
rect 958 31 960 33
rect 963 30 965 33
rect 979 31 981 33
rect 995 31 997 33
rect 1000 28 1002 33
rect 1021 28 1023 33
rect 1037 31 1039 33
rect 1053 31 1055 33
rect 1058 28 1060 33
rect 1074 31 1076 33
rect 1090 31 1092 33
rect 1095 30 1097 33
rect 1111 31 1113 33
rect 1127 31 1129 33
rect 1132 28 1134 33
rect 1153 28 1155 33
rect 1169 31 1171 33
rect 1185 31 1187 33
rect 1190 28 1192 33
rect 1206 31 1208 33
rect 1222 31 1224 33
rect 1227 30 1229 33
rect 1243 31 1245 33
rect 1259 31 1261 33
rect 1264 28 1266 33
rect 1285 28 1287 33
rect 1301 31 1303 33
rect 1317 31 1319 33
rect 1322 28 1324 33
rect 1338 31 1340 33
<< polycontact >>
rect 502 1948 506 1952
rect 539 1948 543 1952
rect 559 1948 563 1952
rect 597 1948 601 1952
rect 634 1948 638 1952
rect 671 1948 675 1952
rect 691 1948 695 1952
rect 729 1948 733 1952
rect 766 1948 770 1952
rect 803 1948 807 1952
rect 823 1948 827 1952
rect 861 1948 865 1952
rect 898 1948 902 1952
rect 935 1948 939 1952
rect 955 1948 959 1952
rect 993 1948 997 1952
rect 1435 1948 1439 1952
rect 1472 1948 1476 1952
rect 1492 1948 1496 1952
rect 1530 1948 1534 1952
rect 1567 1948 1571 1952
rect 1604 1948 1608 1952
rect 1624 1948 1628 1952
rect 1662 1948 1666 1952
rect 1699 1948 1703 1952
rect 1736 1948 1740 1952
rect 1756 1948 1760 1952
rect 1794 1948 1798 1952
rect 1831 1948 1835 1952
rect 1868 1948 1872 1952
rect 1888 1948 1892 1952
rect 1926 1948 1930 1952
rect 496 1928 500 1932
rect 514 1930 518 1934
rect 162 1915 166 1919
rect 199 1915 203 1919
rect 219 1915 223 1919
rect 257 1915 261 1919
rect 574 1930 578 1934
rect 532 1921 536 1928
rect 590 1921 594 1928
rect 611 1925 615 1929
rect 628 1928 632 1932
rect 646 1930 650 1934
rect 706 1930 710 1934
rect 664 1921 668 1928
rect 722 1921 726 1928
rect 743 1925 747 1929
rect 760 1928 764 1932
rect 778 1930 782 1934
rect 838 1930 842 1934
rect 796 1921 800 1928
rect 854 1921 858 1928
rect 875 1925 879 1929
rect 892 1928 896 1932
rect 910 1930 914 1934
rect 970 1930 974 1934
rect 928 1921 932 1928
rect 986 1921 990 1928
rect 1007 1925 1011 1929
rect 1429 1928 1433 1932
rect 1447 1930 1451 1934
rect 1095 1915 1099 1919
rect 1132 1915 1136 1919
rect 1152 1915 1156 1919
rect 1190 1915 1194 1919
rect 1507 1930 1511 1934
rect 1465 1921 1469 1928
rect 1523 1921 1527 1928
rect 1544 1925 1548 1929
rect 1561 1928 1565 1932
rect 1579 1930 1583 1934
rect 1639 1930 1643 1934
rect 1597 1921 1601 1928
rect 1655 1921 1659 1928
rect 1676 1925 1680 1929
rect 1693 1928 1697 1932
rect 1711 1930 1715 1934
rect 1771 1930 1775 1934
rect 1729 1921 1733 1928
rect 1787 1921 1791 1928
rect 1808 1925 1812 1929
rect 1825 1928 1829 1932
rect 1843 1930 1847 1934
rect 1903 1930 1907 1934
rect 1861 1921 1865 1928
rect 1919 1921 1923 1928
rect 1940 1925 1944 1929
rect 502 1907 506 1911
rect 539 1905 543 1909
rect 559 1905 563 1909
rect 595 1905 599 1909
rect 634 1907 638 1911
rect 671 1905 675 1909
rect 691 1905 695 1909
rect 727 1905 731 1909
rect 766 1907 770 1911
rect 803 1905 807 1909
rect 823 1905 827 1909
rect 859 1905 863 1909
rect 898 1907 902 1911
rect 935 1905 939 1909
rect 955 1905 959 1909
rect 991 1905 995 1909
rect 1435 1907 1439 1911
rect 1472 1905 1476 1909
rect 1492 1905 1496 1909
rect 1528 1905 1532 1909
rect 1567 1907 1571 1911
rect 1604 1905 1608 1909
rect 1624 1905 1628 1909
rect 1660 1905 1664 1909
rect 1699 1907 1703 1911
rect 1736 1905 1740 1909
rect 1756 1905 1760 1909
rect 1792 1905 1796 1909
rect 1831 1907 1835 1911
rect 1868 1905 1872 1909
rect 1888 1905 1892 1909
rect 1924 1905 1928 1909
rect 156 1895 160 1899
rect 174 1897 178 1901
rect 234 1897 238 1901
rect 192 1888 196 1895
rect 250 1888 254 1895
rect 269 1892 273 1896
rect 1089 1895 1093 1899
rect 1107 1897 1111 1901
rect 1167 1897 1171 1901
rect 1125 1888 1129 1895
rect 1183 1888 1187 1895
rect 1202 1892 1206 1896
rect 162 1874 166 1878
rect 199 1872 203 1876
rect 219 1872 223 1876
rect 255 1872 259 1876
rect 518 1864 522 1868
rect 562 1864 566 1868
rect 589 1864 593 1868
rect 634 1864 638 1868
rect 707 1871 711 1875
rect 280 1851 284 1855
rect 672 1857 676 1861
rect 163 1842 167 1846
rect 498 1844 502 1848
rect 530 1845 534 1849
rect 549 1844 553 1848
rect 605 1845 609 1849
rect 621 1844 625 1848
rect 648 1844 652 1848
rect 788 1871 792 1875
rect 1095 1874 1099 1878
rect 699 1853 703 1857
rect 726 1849 730 1853
rect 753 1857 757 1861
rect 1132 1872 1136 1876
rect 1152 1872 1156 1876
rect 1188 1872 1192 1876
rect 780 1853 784 1857
rect 807 1849 811 1853
rect 1451 1864 1455 1868
rect 1495 1864 1499 1868
rect 1522 1864 1526 1868
rect 1567 1864 1571 1868
rect 1640 1871 1644 1875
rect 1213 1851 1217 1855
rect 1605 1857 1609 1861
rect 705 1835 709 1839
rect 1096 1842 1100 1846
rect 1431 1844 1435 1848
rect 786 1835 790 1839
rect 1463 1845 1467 1849
rect 1482 1844 1486 1848
rect 1538 1845 1542 1849
rect 1554 1844 1558 1848
rect 1581 1844 1585 1848
rect 1721 1871 1725 1875
rect 1632 1853 1636 1857
rect 1659 1849 1663 1853
rect 1686 1857 1690 1861
rect 1713 1853 1717 1857
rect 1740 1849 1744 1853
rect 1638 1835 1642 1839
rect 1719 1835 1723 1839
rect 515 1827 519 1831
rect 559 1826 563 1830
rect 584 1827 589 1831
rect 631 1826 635 1830
rect 1448 1827 1452 1831
rect 1492 1826 1496 1830
rect 1517 1827 1522 1831
rect 1564 1826 1568 1830
rect 162 1813 166 1817
rect 200 1813 204 1817
rect 220 1813 224 1817
rect 257 1813 261 1817
rect 1095 1813 1099 1817
rect 1133 1813 1137 1817
rect 1153 1813 1157 1817
rect 1190 1813 1194 1817
rect 150 1790 154 1794
rect 185 1795 189 1799
rect 169 1786 173 1793
rect 227 1786 231 1793
rect 245 1795 249 1799
rect 515 1797 519 1801
rect 559 1798 563 1802
rect 263 1793 267 1797
rect 584 1797 589 1801
rect 631 1798 635 1802
rect 707 1795 711 1799
rect 788 1795 792 1799
rect 498 1780 502 1784
rect 164 1770 168 1774
rect 200 1770 204 1774
rect 220 1770 224 1774
rect 257 1772 261 1776
rect 530 1779 534 1783
rect 549 1780 553 1784
rect 605 1779 609 1783
rect 621 1780 625 1784
rect 648 1780 652 1784
rect 696 1779 702 1783
rect 777 1779 783 1783
rect 1083 1790 1087 1794
rect 1118 1795 1122 1799
rect 1102 1786 1106 1793
rect 1160 1786 1164 1793
rect 1178 1795 1182 1799
rect 1448 1797 1452 1801
rect 1492 1798 1496 1802
rect 1196 1793 1200 1797
rect 1517 1797 1522 1801
rect 1564 1798 1568 1802
rect 1640 1795 1644 1799
rect 1721 1795 1725 1799
rect 1431 1780 1435 1784
rect 1097 1770 1101 1774
rect 1133 1770 1137 1774
rect 1153 1770 1157 1774
rect 1190 1772 1194 1776
rect 1463 1779 1467 1783
rect 1482 1780 1486 1784
rect 1538 1779 1542 1783
rect 1554 1780 1558 1784
rect 1581 1780 1585 1784
rect 1629 1779 1635 1783
rect 1710 1779 1716 1783
rect 518 1760 522 1764
rect 562 1760 566 1764
rect 589 1760 593 1764
rect 634 1760 638 1764
rect 705 1759 709 1763
rect 786 1759 790 1763
rect 1451 1760 1455 1764
rect 1495 1760 1499 1764
rect 1522 1760 1526 1764
rect 1567 1760 1571 1764
rect 1638 1759 1642 1763
rect 1719 1759 1723 1763
rect 707 1739 711 1743
rect 518 1732 522 1736
rect 562 1732 566 1736
rect 589 1732 593 1736
rect 634 1732 638 1736
rect 812 1739 816 1743
rect 699 1721 703 1725
rect 498 1712 502 1716
rect 530 1713 534 1717
rect 549 1712 553 1716
rect 605 1713 609 1717
rect 621 1712 625 1716
rect 648 1712 652 1716
rect 726 1717 730 1721
rect 777 1725 781 1729
rect 1640 1739 1644 1743
rect 804 1721 808 1725
rect 831 1717 835 1721
rect 1451 1732 1455 1736
rect 1495 1732 1499 1736
rect 1522 1732 1526 1736
rect 1567 1732 1571 1736
rect 1745 1739 1749 1743
rect 1632 1721 1636 1725
rect 1431 1712 1435 1716
rect 705 1703 709 1707
rect 810 1703 814 1707
rect 1463 1713 1467 1717
rect 1482 1712 1486 1716
rect 1538 1713 1542 1717
rect 1554 1712 1558 1716
rect 1581 1712 1585 1716
rect 1659 1717 1663 1721
rect 1710 1725 1714 1729
rect 1737 1721 1741 1725
rect 1764 1717 1768 1721
rect 1638 1703 1642 1707
rect 1743 1703 1747 1707
rect 515 1695 519 1699
rect 559 1694 563 1698
rect 584 1695 589 1699
rect 631 1694 635 1698
rect 1448 1695 1452 1699
rect 1492 1694 1496 1698
rect 1517 1695 1522 1699
rect 1564 1694 1568 1698
rect 515 1665 519 1669
rect 559 1666 563 1670
rect 584 1665 589 1669
rect 631 1666 635 1670
rect 707 1664 711 1668
rect 812 1664 816 1668
rect 1448 1665 1452 1669
rect 1492 1666 1496 1670
rect 1517 1665 1522 1669
rect 1564 1666 1568 1670
rect 1640 1664 1644 1668
rect 1745 1664 1749 1668
rect 498 1648 502 1652
rect 530 1647 534 1651
rect 549 1648 553 1652
rect 605 1647 609 1651
rect 621 1648 625 1652
rect 648 1648 652 1652
rect 696 1648 702 1652
rect 801 1648 807 1652
rect 1431 1648 1435 1652
rect 1463 1647 1467 1651
rect 1482 1648 1486 1652
rect 1538 1647 1542 1651
rect 1554 1648 1558 1652
rect 1581 1648 1585 1652
rect 1629 1648 1635 1652
rect 1734 1648 1740 1652
rect 518 1628 522 1632
rect 562 1628 566 1632
rect 589 1628 593 1632
rect 634 1628 638 1632
rect 705 1628 709 1632
rect 810 1628 814 1632
rect 1451 1628 1455 1632
rect 1495 1628 1499 1632
rect 1522 1628 1526 1632
rect 1567 1628 1571 1632
rect 1638 1628 1642 1632
rect 1743 1628 1747 1632
rect 707 1607 711 1611
rect 518 1600 522 1604
rect 562 1600 566 1604
rect 589 1600 593 1604
rect 634 1600 638 1604
rect 788 1607 792 1611
rect 699 1589 703 1593
rect 498 1580 502 1584
rect 530 1581 534 1585
rect 549 1580 553 1584
rect 605 1581 609 1585
rect 621 1580 625 1584
rect 648 1580 652 1584
rect 726 1585 730 1589
rect 753 1593 757 1597
rect 878 1607 882 1611
rect 780 1589 784 1593
rect 807 1585 811 1589
rect 843 1593 847 1597
rect 1640 1607 1644 1611
rect 870 1589 874 1593
rect 897 1585 901 1589
rect 1451 1600 1455 1604
rect 1495 1600 1499 1604
rect 1522 1600 1526 1604
rect 1567 1600 1571 1604
rect 1721 1607 1725 1611
rect 1632 1589 1636 1593
rect 1431 1580 1435 1584
rect 705 1571 709 1575
rect 786 1571 790 1575
rect 876 1571 880 1575
rect 1463 1581 1467 1585
rect 1482 1580 1486 1584
rect 1538 1581 1542 1585
rect 1554 1580 1558 1584
rect 1581 1580 1585 1584
rect 1659 1585 1663 1589
rect 1686 1593 1690 1597
rect 1811 1607 1815 1611
rect 1713 1589 1717 1593
rect 1740 1585 1744 1589
rect 1776 1593 1780 1597
rect 1803 1589 1807 1593
rect 1830 1585 1834 1589
rect 1638 1571 1642 1575
rect 1719 1571 1723 1575
rect 1809 1571 1813 1575
rect 515 1563 519 1567
rect 559 1562 563 1566
rect 584 1563 589 1567
rect 631 1562 635 1566
rect 1448 1563 1452 1567
rect 1492 1562 1496 1566
rect 1517 1563 1522 1567
rect 1564 1562 1568 1566
rect 515 1533 519 1537
rect 559 1534 563 1538
rect 584 1533 589 1537
rect 631 1534 635 1538
rect 1448 1533 1452 1537
rect 1492 1534 1496 1538
rect 707 1529 711 1533
rect 788 1529 792 1533
rect 878 1529 882 1533
rect 1517 1533 1522 1537
rect 1564 1534 1568 1538
rect 1640 1529 1644 1533
rect 1721 1529 1725 1533
rect 1811 1529 1815 1533
rect 498 1516 502 1520
rect 530 1515 534 1519
rect 549 1516 553 1520
rect 605 1515 609 1519
rect 621 1516 625 1520
rect 648 1516 652 1520
rect 696 1513 702 1517
rect 777 1513 783 1517
rect 867 1513 873 1517
rect 1431 1516 1435 1520
rect 1463 1515 1467 1519
rect 1482 1516 1486 1520
rect 1538 1515 1542 1519
rect 1554 1516 1558 1520
rect 1581 1516 1585 1520
rect 1629 1513 1635 1517
rect 1710 1513 1716 1517
rect 1800 1513 1806 1517
rect 518 1496 522 1500
rect 562 1496 566 1500
rect 589 1496 593 1500
rect 634 1496 638 1500
rect 705 1493 709 1497
rect 786 1493 790 1497
rect 876 1493 880 1497
rect 1451 1496 1455 1500
rect 1495 1496 1499 1500
rect 1522 1496 1526 1500
rect 1567 1496 1571 1500
rect 1638 1493 1642 1497
rect 1719 1493 1723 1497
rect 1809 1493 1813 1497
rect 707 1475 711 1479
rect 518 1468 522 1472
rect 562 1468 566 1472
rect 589 1468 593 1472
rect 634 1468 638 1472
rect 1640 1475 1644 1479
rect 699 1457 703 1461
rect 498 1448 502 1452
rect 530 1449 534 1453
rect 549 1448 553 1452
rect 605 1449 609 1453
rect 621 1448 625 1452
rect 648 1448 652 1452
rect 726 1453 730 1457
rect 1451 1468 1455 1472
rect 1495 1468 1499 1472
rect 1522 1468 1526 1472
rect 1567 1468 1571 1472
rect 1632 1457 1636 1461
rect 1431 1448 1435 1452
rect 705 1439 709 1443
rect 1463 1449 1467 1453
rect 1482 1448 1486 1452
rect 1538 1449 1542 1453
rect 1554 1448 1558 1452
rect 1581 1448 1585 1452
rect 1659 1453 1663 1457
rect 1638 1439 1642 1443
rect 515 1431 519 1435
rect 559 1430 563 1434
rect 584 1431 589 1435
rect 631 1430 635 1434
rect 1448 1431 1452 1435
rect 1492 1430 1496 1434
rect 1517 1431 1522 1435
rect 1564 1430 1568 1434
rect 30 1413 34 1417
rect 67 1413 71 1417
rect 87 1413 91 1417
rect 125 1413 129 1417
rect 162 1413 166 1417
rect 199 1413 203 1417
rect 219 1413 223 1417
rect 257 1413 261 1417
rect 294 1413 298 1417
rect 331 1413 335 1417
rect 351 1413 355 1417
rect 389 1413 393 1417
rect 963 1413 967 1417
rect 1000 1413 1004 1417
rect 1020 1413 1024 1417
rect 1058 1413 1062 1417
rect 1095 1413 1099 1417
rect 1132 1413 1136 1417
rect 1152 1413 1156 1417
rect 1190 1413 1194 1417
rect 1227 1413 1231 1417
rect 1264 1413 1268 1417
rect 1284 1413 1288 1417
rect 1322 1413 1326 1417
rect 24 1393 28 1397
rect 42 1395 46 1399
rect 102 1395 106 1399
rect 60 1386 64 1393
rect 118 1386 122 1393
rect 137 1390 141 1394
rect 155 1395 159 1399
rect 174 1395 178 1399
rect 234 1395 238 1399
rect 192 1386 196 1393
rect 250 1386 254 1393
rect 269 1390 273 1394
rect 287 1395 291 1399
rect 306 1395 310 1399
rect 366 1395 370 1399
rect 324 1386 328 1393
rect 515 1401 519 1405
rect 559 1402 563 1406
rect 584 1401 589 1405
rect 631 1402 635 1406
rect 776 1401 780 1405
rect 820 1402 824 1406
rect 845 1401 850 1405
rect 892 1402 896 1406
rect 382 1386 386 1393
rect 403 1390 407 1394
rect 707 1393 711 1397
rect 957 1393 961 1397
rect 975 1395 979 1399
rect 498 1384 502 1388
rect 530 1383 534 1387
rect 549 1384 553 1388
rect 605 1383 609 1387
rect 621 1384 625 1388
rect 648 1384 652 1388
rect 30 1372 34 1376
rect 67 1370 71 1374
rect 87 1370 91 1374
rect 123 1370 127 1374
rect 162 1372 166 1376
rect 199 1370 203 1374
rect 219 1370 223 1374
rect 255 1370 259 1374
rect 294 1372 298 1376
rect 331 1370 335 1374
rect 351 1370 355 1374
rect 387 1370 391 1374
rect 696 1377 702 1381
rect 734 1384 738 1388
rect 791 1383 795 1387
rect 810 1384 814 1388
rect 866 1383 870 1387
rect 882 1384 886 1388
rect 909 1384 913 1388
rect 1035 1395 1039 1399
rect 993 1386 997 1393
rect 1051 1386 1055 1393
rect 1070 1390 1074 1394
rect 1088 1395 1092 1399
rect 1107 1395 1111 1399
rect 1167 1395 1171 1399
rect 1125 1386 1129 1393
rect 1183 1386 1187 1393
rect 1202 1390 1206 1394
rect 1220 1395 1224 1399
rect 1239 1395 1243 1399
rect 1299 1395 1303 1399
rect 1257 1386 1261 1393
rect 1448 1401 1452 1405
rect 1492 1402 1496 1406
rect 1517 1401 1522 1405
rect 1564 1402 1568 1406
rect 1709 1401 1713 1405
rect 1753 1402 1757 1406
rect 1778 1401 1783 1405
rect 1825 1402 1829 1406
rect 1315 1386 1319 1393
rect 1336 1390 1340 1394
rect 1640 1393 1644 1397
rect 1431 1384 1435 1388
rect 1463 1383 1467 1387
rect 1482 1384 1486 1388
rect 1538 1383 1542 1387
rect 1554 1384 1558 1388
rect 1581 1384 1585 1388
rect 518 1364 522 1368
rect 562 1364 566 1368
rect 589 1364 593 1368
rect 634 1364 638 1368
rect 963 1372 967 1376
rect 1000 1370 1004 1374
rect 1020 1370 1024 1374
rect 1056 1370 1060 1374
rect 1095 1372 1099 1376
rect 1132 1370 1136 1374
rect 1152 1370 1156 1374
rect 1188 1370 1192 1374
rect 1227 1372 1231 1376
rect 1264 1370 1268 1374
rect 1284 1370 1288 1374
rect 1320 1370 1324 1374
rect 1629 1377 1635 1381
rect 1667 1384 1671 1388
rect 1724 1383 1728 1387
rect 1743 1384 1747 1388
rect 1799 1383 1803 1387
rect 1815 1384 1819 1388
rect 1842 1384 1846 1388
rect 779 1364 783 1368
rect 823 1364 827 1368
rect 850 1364 854 1368
rect 895 1364 899 1368
rect 1451 1364 1455 1368
rect 1495 1364 1499 1368
rect 1522 1364 1526 1368
rect 1567 1364 1571 1368
rect 1712 1364 1716 1368
rect 1756 1364 1760 1368
rect 1783 1364 1787 1368
rect 1828 1364 1832 1368
rect 705 1357 709 1361
rect 1638 1357 1642 1361
rect 139 1342 143 1346
rect 163 1342 167 1346
rect 1072 1342 1076 1346
rect 1096 1342 1100 1346
rect 918 1336 922 1340
rect 1851 1336 1855 1340
rect 159 1317 163 1321
rect 1092 1317 1096 1321
rect 174 1309 178 1313
rect 1107 1309 1111 1313
rect 801 1303 805 1307
rect 838 1303 842 1307
rect 858 1303 862 1307
rect 896 1303 900 1307
rect 1734 1303 1738 1307
rect 1771 1303 1775 1307
rect 1791 1303 1795 1307
rect 1829 1303 1833 1307
rect 139 1294 143 1298
rect 163 1294 167 1298
rect 1072 1294 1076 1298
rect 1096 1294 1100 1298
rect 795 1283 799 1287
rect 813 1285 817 1289
rect 30 1273 34 1277
rect 67 1273 71 1277
rect 87 1273 91 1277
rect 125 1273 129 1277
rect 162 1273 166 1277
rect 199 1273 203 1277
rect 219 1273 223 1277
rect 257 1273 261 1277
rect 294 1273 298 1277
rect 331 1273 335 1277
rect 351 1273 355 1277
rect 389 1273 393 1277
rect 873 1285 877 1289
rect 831 1276 835 1283
rect 889 1276 893 1283
rect 908 1280 912 1284
rect 1728 1283 1732 1287
rect 1746 1285 1750 1289
rect 963 1273 967 1277
rect 1000 1273 1004 1277
rect 1020 1273 1024 1277
rect 1058 1273 1062 1277
rect 1095 1273 1099 1277
rect 1132 1273 1136 1277
rect 1152 1273 1156 1277
rect 1190 1273 1194 1277
rect 1227 1273 1231 1277
rect 1264 1273 1268 1277
rect 1284 1273 1288 1277
rect 1322 1273 1326 1277
rect 1806 1285 1810 1289
rect 1764 1276 1768 1283
rect 1822 1276 1826 1283
rect 1841 1280 1845 1284
rect 801 1262 805 1266
rect 24 1253 28 1257
rect 42 1255 46 1259
rect 102 1255 106 1259
rect 60 1246 64 1253
rect 118 1246 122 1253
rect 137 1250 141 1254
rect 155 1255 159 1259
rect 174 1255 178 1259
rect 234 1255 238 1259
rect 192 1246 196 1253
rect 250 1246 254 1253
rect 269 1250 273 1254
rect 287 1255 291 1259
rect 306 1255 310 1259
rect 366 1255 370 1259
rect 324 1246 328 1253
rect 838 1260 842 1264
rect 858 1260 862 1264
rect 894 1260 898 1264
rect 1734 1262 1738 1266
rect 382 1246 386 1253
rect 403 1250 407 1254
rect 957 1253 961 1257
rect 975 1255 979 1259
rect 1035 1255 1039 1259
rect 993 1246 997 1253
rect 1051 1246 1055 1253
rect 1070 1250 1074 1254
rect 1088 1255 1092 1259
rect 1107 1255 1111 1259
rect 1167 1255 1171 1259
rect 1125 1246 1129 1253
rect 1183 1246 1187 1253
rect 1202 1250 1206 1254
rect 1220 1255 1224 1259
rect 1239 1255 1243 1259
rect 1299 1255 1303 1259
rect 1257 1246 1261 1253
rect 1771 1260 1775 1264
rect 1791 1260 1795 1264
rect 1827 1260 1831 1264
rect 1315 1246 1319 1253
rect 1336 1250 1340 1254
rect 30 1232 34 1236
rect 67 1230 71 1234
rect 87 1230 91 1234
rect 123 1230 127 1234
rect 162 1232 166 1236
rect 199 1230 203 1234
rect 219 1230 223 1234
rect 255 1230 259 1234
rect 294 1232 298 1236
rect 331 1230 335 1234
rect 351 1230 355 1234
rect 387 1230 391 1234
rect 963 1232 967 1236
rect 1000 1230 1004 1234
rect 1020 1230 1024 1234
rect 1056 1230 1060 1234
rect 1095 1232 1099 1236
rect 1132 1230 1136 1234
rect 1152 1230 1156 1234
rect 1188 1230 1192 1234
rect 1227 1232 1231 1236
rect 1264 1230 1268 1234
rect 1284 1230 1288 1234
rect 1320 1230 1324 1234
rect 801 1217 805 1221
rect 838 1217 842 1221
rect 858 1217 862 1221
rect 896 1217 900 1221
rect 1734 1217 1738 1221
rect 1771 1217 1775 1221
rect 1791 1217 1795 1221
rect 1829 1217 1833 1221
rect 795 1197 799 1201
rect 813 1199 817 1203
rect 30 1187 34 1191
rect 67 1187 71 1191
rect 87 1187 91 1191
rect 125 1187 129 1191
rect 162 1187 166 1191
rect 199 1187 203 1191
rect 219 1187 223 1191
rect 257 1187 261 1191
rect 294 1187 298 1191
rect 331 1187 335 1191
rect 351 1187 355 1191
rect 389 1187 393 1191
rect 873 1199 877 1203
rect 831 1190 835 1197
rect 889 1190 893 1197
rect 908 1194 912 1198
rect 930 1192 934 1196
rect 1728 1197 1732 1201
rect 1746 1199 1750 1203
rect 963 1187 967 1191
rect 1000 1187 1004 1191
rect 1020 1187 1024 1191
rect 1058 1187 1062 1191
rect 1095 1187 1099 1191
rect 1132 1187 1136 1191
rect 1152 1187 1156 1191
rect 1190 1187 1194 1191
rect 1227 1187 1231 1191
rect 1264 1187 1268 1191
rect 1284 1187 1288 1191
rect 1322 1187 1326 1191
rect 1806 1199 1810 1203
rect 1764 1190 1768 1197
rect 1822 1190 1826 1197
rect 1841 1194 1845 1198
rect 1863 1192 1867 1196
rect 801 1176 805 1180
rect 24 1167 28 1171
rect 42 1169 46 1173
rect 102 1169 106 1173
rect 60 1160 64 1167
rect 118 1160 122 1167
rect 137 1164 141 1168
rect 155 1169 159 1173
rect 174 1169 178 1173
rect 234 1169 238 1173
rect 192 1160 196 1167
rect 250 1160 254 1167
rect 269 1164 273 1168
rect 287 1169 291 1173
rect 306 1169 310 1173
rect 366 1169 370 1173
rect 324 1160 328 1167
rect 838 1174 842 1178
rect 858 1174 862 1178
rect 894 1174 898 1178
rect 1734 1176 1738 1180
rect 382 1160 386 1167
rect 403 1164 407 1168
rect 957 1167 961 1171
rect 975 1169 979 1173
rect 1035 1169 1039 1173
rect 993 1160 997 1167
rect 1051 1160 1055 1167
rect 1070 1164 1074 1168
rect 1088 1169 1092 1173
rect 1107 1169 1111 1173
rect 1167 1169 1171 1173
rect 1125 1160 1129 1167
rect 1183 1160 1187 1167
rect 1202 1164 1206 1168
rect 1220 1169 1224 1173
rect 1239 1169 1243 1173
rect 1299 1169 1303 1173
rect 1257 1160 1261 1167
rect 1771 1174 1775 1178
rect 1791 1174 1795 1178
rect 1827 1174 1831 1178
rect 1315 1160 1319 1167
rect 1336 1164 1340 1168
rect 30 1146 34 1150
rect 67 1144 71 1148
rect 87 1144 91 1148
rect 123 1144 127 1148
rect 162 1146 166 1150
rect 199 1144 203 1148
rect 219 1144 223 1148
rect 255 1144 259 1148
rect 294 1146 298 1150
rect 331 1144 335 1148
rect 351 1144 355 1148
rect 387 1144 391 1148
rect 963 1146 967 1150
rect 1000 1144 1004 1148
rect 1020 1144 1024 1148
rect 1056 1144 1060 1148
rect 1095 1146 1099 1150
rect 1132 1144 1136 1148
rect 1152 1144 1156 1148
rect 1188 1144 1192 1148
rect 1227 1146 1231 1150
rect 1264 1144 1268 1148
rect 1284 1144 1288 1148
rect 1320 1144 1324 1148
rect 256 1116 260 1120
rect 280 1116 284 1120
rect 1189 1116 1193 1120
rect 1213 1116 1217 1120
rect 276 1091 280 1095
rect 1209 1091 1213 1095
rect 291 1083 295 1087
rect 1224 1083 1228 1087
rect 256 1068 260 1072
rect 280 1068 284 1072
rect 1189 1068 1193 1072
rect 1213 1068 1217 1072
rect 30 1047 34 1051
rect 67 1047 71 1051
rect 87 1047 91 1051
rect 125 1047 129 1051
rect 162 1047 166 1051
rect 199 1047 203 1051
rect 219 1047 223 1051
rect 257 1047 261 1051
rect 294 1047 298 1051
rect 331 1047 335 1051
rect 351 1047 355 1051
rect 389 1047 393 1051
rect 963 1047 967 1051
rect 1000 1047 1004 1051
rect 1020 1047 1024 1051
rect 1058 1047 1062 1051
rect 1095 1047 1099 1051
rect 1132 1047 1136 1051
rect 1152 1047 1156 1051
rect 1190 1047 1194 1051
rect 1227 1047 1231 1051
rect 1264 1047 1268 1051
rect 1284 1047 1288 1051
rect 1322 1047 1326 1051
rect 24 1027 28 1031
rect 42 1029 46 1033
rect 102 1029 106 1033
rect 60 1020 64 1027
rect 118 1020 122 1027
rect 137 1024 141 1028
rect 155 1029 159 1033
rect 174 1029 178 1033
rect 234 1029 238 1033
rect 192 1020 196 1027
rect 250 1020 254 1027
rect 269 1024 273 1028
rect 287 1029 291 1033
rect 306 1029 310 1033
rect 366 1029 370 1033
rect 324 1020 328 1027
rect 382 1020 386 1027
rect 403 1024 407 1028
rect 957 1027 961 1031
rect 975 1029 979 1033
rect 1035 1029 1039 1033
rect 993 1020 997 1027
rect 1051 1020 1055 1027
rect 1070 1024 1074 1028
rect 1088 1029 1092 1033
rect 1107 1029 1111 1033
rect 1167 1029 1171 1033
rect 1125 1020 1129 1027
rect 1183 1020 1187 1027
rect 1202 1024 1206 1028
rect 1220 1029 1224 1033
rect 1239 1029 1243 1033
rect 1299 1029 1303 1033
rect 1257 1020 1261 1027
rect 1315 1020 1319 1027
rect 1336 1024 1340 1028
rect 30 1006 34 1010
rect 67 1004 71 1008
rect 87 1004 91 1008
rect 123 1004 127 1008
rect 162 1006 166 1010
rect 199 1004 203 1008
rect 219 1004 223 1008
rect 255 1004 259 1008
rect 294 1006 298 1010
rect 331 1004 335 1008
rect 351 1004 355 1008
rect 387 1004 391 1008
rect 963 1006 967 1010
rect 1000 1004 1004 1008
rect 1020 1004 1024 1008
rect 1056 1004 1060 1008
rect 1095 1006 1099 1010
rect 1132 1004 1136 1008
rect 1152 1004 1156 1008
rect 1188 1004 1192 1008
rect 1227 1006 1231 1010
rect 1264 1004 1268 1008
rect 1284 1004 1288 1008
rect 1320 1004 1324 1008
rect 502 968 506 972
rect 539 968 543 972
rect 559 968 563 972
rect 597 968 601 972
rect 634 968 638 972
rect 671 968 675 972
rect 691 968 695 972
rect 729 968 733 972
rect 766 968 770 972
rect 803 968 807 972
rect 823 968 827 972
rect 861 968 865 972
rect 898 968 902 972
rect 935 968 939 972
rect 955 968 959 972
rect 993 968 997 972
rect 1435 968 1439 972
rect 1472 968 1476 972
rect 1492 968 1496 972
rect 1530 968 1534 972
rect 1567 968 1571 972
rect 1604 968 1608 972
rect 1624 968 1628 972
rect 1662 968 1666 972
rect 1699 968 1703 972
rect 1736 968 1740 972
rect 1756 968 1760 972
rect 1794 968 1798 972
rect 1831 968 1835 972
rect 1868 968 1872 972
rect 1888 968 1892 972
rect 1926 968 1930 972
rect 496 948 500 952
rect 514 950 518 954
rect 162 935 166 939
rect 199 935 203 939
rect 219 935 223 939
rect 257 935 261 939
rect 574 950 578 954
rect 532 941 536 948
rect 590 941 594 948
rect 611 945 615 949
rect 628 948 632 952
rect 646 950 650 954
rect 706 950 710 954
rect 664 941 668 948
rect 722 941 726 948
rect 743 945 747 949
rect 760 948 764 952
rect 778 950 782 954
rect 838 950 842 954
rect 796 941 800 948
rect 854 941 858 948
rect 875 945 879 949
rect 892 948 896 952
rect 910 950 914 954
rect 970 950 974 954
rect 928 941 932 948
rect 986 941 990 948
rect 1007 945 1011 949
rect 1429 948 1433 952
rect 1447 950 1451 954
rect 1095 935 1099 939
rect 1132 935 1136 939
rect 1152 935 1156 939
rect 1190 935 1194 939
rect 1507 950 1511 954
rect 1465 941 1469 948
rect 1523 941 1527 948
rect 1544 945 1548 949
rect 1561 948 1565 952
rect 1579 950 1583 954
rect 1639 950 1643 954
rect 1597 941 1601 948
rect 1655 941 1659 948
rect 1676 945 1680 949
rect 1693 948 1697 952
rect 1711 950 1715 954
rect 1771 950 1775 954
rect 1729 941 1733 948
rect 1787 941 1791 948
rect 1808 945 1812 949
rect 1825 948 1829 952
rect 1843 950 1847 954
rect 1903 950 1907 954
rect 1861 941 1865 948
rect 1919 941 1923 948
rect 1940 945 1944 949
rect 502 927 506 931
rect 539 925 543 929
rect 559 925 563 929
rect 595 925 599 929
rect 634 927 638 931
rect 671 925 675 929
rect 691 925 695 929
rect 727 925 731 929
rect 766 927 770 931
rect 803 925 807 929
rect 823 925 827 929
rect 859 925 863 929
rect 898 927 902 931
rect 935 925 939 929
rect 955 925 959 929
rect 991 925 995 929
rect 1435 927 1439 931
rect 1472 925 1476 929
rect 1492 925 1496 929
rect 1528 925 1532 929
rect 1567 927 1571 931
rect 1604 925 1608 929
rect 1624 925 1628 929
rect 1660 925 1664 929
rect 1699 927 1703 931
rect 1736 925 1740 929
rect 1756 925 1760 929
rect 1792 925 1796 929
rect 1831 927 1835 931
rect 1868 925 1872 929
rect 1888 925 1892 929
rect 1924 925 1928 929
rect 156 915 160 919
rect 174 917 178 921
rect 234 917 238 921
rect 192 908 196 915
rect 250 908 254 915
rect 269 912 273 916
rect 1089 915 1093 919
rect 1107 917 1111 921
rect 1167 917 1171 921
rect 1125 908 1129 915
rect 1183 908 1187 915
rect 1202 912 1206 916
rect 162 894 166 898
rect 199 892 203 896
rect 219 892 223 896
rect 255 892 259 896
rect 518 884 522 888
rect 562 884 566 888
rect 589 884 593 888
rect 634 884 638 888
rect 707 891 711 895
rect 280 871 284 875
rect 672 877 676 881
rect 163 862 167 866
rect 498 864 502 868
rect 530 865 534 869
rect 549 864 553 868
rect 605 865 609 869
rect 621 864 625 868
rect 648 864 652 868
rect 788 891 792 895
rect 1095 894 1099 898
rect 699 873 703 877
rect 726 869 730 873
rect 753 877 757 881
rect 1132 892 1136 896
rect 1152 892 1156 896
rect 1188 892 1192 896
rect 780 873 784 877
rect 807 869 811 873
rect 1451 884 1455 888
rect 1495 884 1499 888
rect 1522 884 1526 888
rect 1567 884 1571 888
rect 1640 891 1644 895
rect 1213 871 1217 875
rect 1605 877 1609 881
rect 705 855 709 859
rect 1096 862 1100 866
rect 1431 864 1435 868
rect 786 855 790 859
rect 1463 865 1467 869
rect 1482 864 1486 868
rect 1538 865 1542 869
rect 1554 864 1558 868
rect 1581 864 1585 868
rect 1721 891 1725 895
rect 1632 873 1636 877
rect 1659 869 1663 873
rect 1686 877 1690 881
rect 1713 873 1717 877
rect 1740 869 1744 873
rect 1638 855 1642 859
rect 1719 855 1723 859
rect 515 847 519 851
rect 559 846 563 850
rect 584 847 589 851
rect 631 846 635 850
rect 1448 847 1452 851
rect 1492 846 1496 850
rect 1517 847 1522 851
rect 1564 846 1568 850
rect 162 833 166 837
rect 200 833 204 837
rect 220 833 224 837
rect 257 833 261 837
rect 1095 833 1099 837
rect 1133 833 1137 837
rect 1153 833 1157 837
rect 1190 833 1194 837
rect 150 810 154 814
rect 185 815 189 819
rect 169 806 173 813
rect 227 806 231 813
rect 245 815 249 819
rect 515 817 519 821
rect 559 818 563 822
rect 263 813 267 817
rect 584 817 589 821
rect 631 818 635 822
rect 707 815 711 819
rect 788 815 792 819
rect 498 800 502 804
rect 164 790 168 794
rect 200 790 204 794
rect 220 790 224 794
rect 257 792 261 796
rect 530 799 534 803
rect 549 800 553 804
rect 605 799 609 803
rect 621 800 625 804
rect 648 800 652 804
rect 696 799 702 803
rect 777 799 783 803
rect 1083 810 1087 814
rect 1118 815 1122 819
rect 1102 806 1106 813
rect 1160 806 1164 813
rect 1178 815 1182 819
rect 1448 817 1452 821
rect 1492 818 1496 822
rect 1196 813 1200 817
rect 1517 817 1522 821
rect 1564 818 1568 822
rect 1640 815 1644 819
rect 1721 815 1725 819
rect 1431 800 1435 804
rect 1097 790 1101 794
rect 1133 790 1137 794
rect 1153 790 1157 794
rect 1190 792 1194 796
rect 1463 799 1467 803
rect 1482 800 1486 804
rect 1538 799 1542 803
rect 1554 800 1558 804
rect 1581 800 1585 804
rect 1629 799 1635 803
rect 1710 799 1716 803
rect 518 780 522 784
rect 562 780 566 784
rect 589 780 593 784
rect 634 780 638 784
rect 705 779 709 783
rect 786 779 790 783
rect 1451 780 1455 784
rect 1495 780 1499 784
rect 1522 780 1526 784
rect 1567 780 1571 784
rect 1638 779 1642 783
rect 1719 779 1723 783
rect 707 759 711 763
rect 518 752 522 756
rect 562 752 566 756
rect 589 752 593 756
rect 634 752 638 756
rect 812 759 816 763
rect 699 741 703 745
rect 498 732 502 736
rect 530 733 534 737
rect 549 732 553 736
rect 605 733 609 737
rect 621 732 625 736
rect 648 732 652 736
rect 726 737 730 741
rect 777 745 781 749
rect 1640 759 1644 763
rect 804 741 808 745
rect 831 737 835 741
rect 1451 752 1455 756
rect 1495 752 1499 756
rect 1522 752 1526 756
rect 1567 752 1571 756
rect 1745 759 1749 763
rect 1632 741 1636 745
rect 1431 732 1435 736
rect 705 723 709 727
rect 810 723 814 727
rect 1463 733 1467 737
rect 1482 732 1486 736
rect 1538 733 1542 737
rect 1554 732 1558 736
rect 1581 732 1585 736
rect 1659 737 1663 741
rect 1710 745 1714 749
rect 1737 741 1741 745
rect 1764 737 1768 741
rect 1638 723 1642 727
rect 1743 723 1747 727
rect 515 715 519 719
rect 559 714 563 718
rect 584 715 589 719
rect 631 714 635 718
rect 1448 715 1452 719
rect 1492 714 1496 718
rect 1517 715 1522 719
rect 1564 714 1568 718
rect 515 685 519 689
rect 559 686 563 690
rect 584 685 589 689
rect 631 686 635 690
rect 707 684 711 688
rect 812 684 816 688
rect 1448 685 1452 689
rect 1492 686 1496 690
rect 1517 685 1522 689
rect 1564 686 1568 690
rect 1640 684 1644 688
rect 1745 684 1749 688
rect 498 668 502 672
rect 530 667 534 671
rect 549 668 553 672
rect 605 667 609 671
rect 621 668 625 672
rect 648 668 652 672
rect 696 668 702 672
rect 801 668 807 672
rect 1431 668 1435 672
rect 1463 667 1467 671
rect 1482 668 1486 672
rect 1538 667 1542 671
rect 1554 668 1558 672
rect 1581 668 1585 672
rect 1629 668 1635 672
rect 1734 668 1740 672
rect 518 648 522 652
rect 562 648 566 652
rect 589 648 593 652
rect 634 648 638 652
rect 705 648 709 652
rect 810 648 814 652
rect 1451 648 1455 652
rect 1495 648 1499 652
rect 1522 648 1526 652
rect 1567 648 1571 652
rect 1638 648 1642 652
rect 1743 648 1747 652
rect 707 627 711 631
rect 518 620 522 624
rect 562 620 566 624
rect 589 620 593 624
rect 634 620 638 624
rect 788 627 792 631
rect 699 609 703 613
rect 498 600 502 604
rect 530 601 534 605
rect 549 600 553 604
rect 605 601 609 605
rect 621 600 625 604
rect 648 600 652 604
rect 726 605 730 609
rect 753 613 757 617
rect 878 627 882 631
rect 780 609 784 613
rect 807 605 811 609
rect 843 613 847 617
rect 1640 627 1644 631
rect 870 609 874 613
rect 897 605 901 609
rect 1451 620 1455 624
rect 1495 620 1499 624
rect 1522 620 1526 624
rect 1567 620 1571 624
rect 1721 627 1725 631
rect 1632 609 1636 613
rect 1431 600 1435 604
rect 705 591 709 595
rect 786 591 790 595
rect 876 591 880 595
rect 1463 601 1467 605
rect 1482 600 1486 604
rect 1538 601 1542 605
rect 1554 600 1558 604
rect 1581 600 1585 604
rect 1659 605 1663 609
rect 1686 613 1690 617
rect 1811 627 1815 631
rect 1713 609 1717 613
rect 1740 605 1744 609
rect 1776 613 1780 617
rect 1803 609 1807 613
rect 1830 605 1834 609
rect 1638 591 1642 595
rect 1719 591 1723 595
rect 1809 591 1813 595
rect 515 583 519 587
rect 559 582 563 586
rect 584 583 589 587
rect 631 582 635 586
rect 1448 583 1452 587
rect 1492 582 1496 586
rect 1517 583 1522 587
rect 1564 582 1568 586
rect 515 553 519 557
rect 559 554 563 558
rect 584 553 589 557
rect 631 554 635 558
rect 1448 553 1452 557
rect 1492 554 1496 558
rect 707 549 711 553
rect 788 549 792 553
rect 878 549 882 553
rect 1517 553 1522 557
rect 1564 554 1568 558
rect 1640 549 1644 553
rect 1721 549 1725 553
rect 1811 549 1815 553
rect 498 536 502 540
rect 530 535 534 539
rect 549 536 553 540
rect 605 535 609 539
rect 621 536 625 540
rect 648 536 652 540
rect 696 533 702 537
rect 777 533 783 537
rect 867 533 873 537
rect 1431 536 1435 540
rect 1463 535 1467 539
rect 1482 536 1486 540
rect 1538 535 1542 539
rect 1554 536 1558 540
rect 1581 536 1585 540
rect 1629 533 1635 537
rect 1710 533 1716 537
rect 1800 533 1806 537
rect 518 516 522 520
rect 562 516 566 520
rect 589 516 593 520
rect 634 516 638 520
rect 705 513 709 517
rect 786 513 790 517
rect 876 513 880 517
rect 1451 516 1455 520
rect 1495 516 1499 520
rect 1522 516 1526 520
rect 1567 516 1571 520
rect 1638 513 1642 517
rect 1719 513 1723 517
rect 1809 513 1813 517
rect 707 495 711 499
rect 518 488 522 492
rect 562 488 566 492
rect 589 488 593 492
rect 634 488 638 492
rect 1640 495 1644 499
rect 699 477 703 481
rect 498 468 502 472
rect 530 469 534 473
rect 549 468 553 472
rect 605 469 609 473
rect 621 468 625 472
rect 648 468 652 472
rect 726 473 730 477
rect 1451 488 1455 492
rect 1495 488 1499 492
rect 1522 488 1526 492
rect 1567 488 1571 492
rect 1632 477 1636 481
rect 1431 468 1435 472
rect 705 459 709 463
rect 1463 469 1467 473
rect 1482 468 1486 472
rect 1538 469 1542 473
rect 1554 468 1558 472
rect 1581 468 1585 472
rect 1659 473 1663 477
rect 1638 459 1642 463
rect 515 451 519 455
rect 559 450 563 454
rect 584 451 589 455
rect 631 450 635 454
rect 1448 451 1452 455
rect 1492 450 1496 454
rect 1517 451 1522 455
rect 1564 450 1568 454
rect 30 433 34 437
rect 67 433 71 437
rect 87 433 91 437
rect 125 433 129 437
rect 162 433 166 437
rect 199 433 203 437
rect 219 433 223 437
rect 257 433 261 437
rect 294 433 298 437
rect 331 433 335 437
rect 351 433 355 437
rect 389 433 393 437
rect 963 433 967 437
rect 1000 433 1004 437
rect 1020 433 1024 437
rect 1058 433 1062 437
rect 1095 433 1099 437
rect 1132 433 1136 437
rect 1152 433 1156 437
rect 1190 433 1194 437
rect 1227 433 1231 437
rect 1264 433 1268 437
rect 1284 433 1288 437
rect 1322 433 1326 437
rect 24 413 28 417
rect 42 415 46 419
rect 102 415 106 419
rect 60 406 64 413
rect 118 406 122 413
rect 137 410 141 414
rect 155 415 159 419
rect 174 415 178 419
rect 234 415 238 419
rect 192 406 196 413
rect 250 406 254 413
rect 269 410 273 414
rect 287 415 291 419
rect 306 415 310 419
rect 366 415 370 419
rect 324 406 328 413
rect 515 421 519 425
rect 559 422 563 426
rect 584 421 589 425
rect 631 422 635 426
rect 776 421 780 425
rect 820 422 824 426
rect 845 421 850 425
rect 892 422 896 426
rect 382 406 386 413
rect 403 410 407 414
rect 707 413 711 417
rect 957 413 961 417
rect 975 415 979 419
rect 498 404 502 408
rect 530 403 534 407
rect 549 404 553 408
rect 605 403 609 407
rect 621 404 625 408
rect 648 404 652 408
rect 30 392 34 396
rect 67 390 71 394
rect 87 390 91 394
rect 123 390 127 394
rect 162 392 166 396
rect 199 390 203 394
rect 219 390 223 394
rect 255 390 259 394
rect 294 392 298 396
rect 331 390 335 394
rect 351 390 355 394
rect 387 390 391 394
rect 696 397 702 401
rect 734 404 738 408
rect 791 403 795 407
rect 810 404 814 408
rect 866 403 870 407
rect 882 404 886 408
rect 909 404 913 408
rect 1035 415 1039 419
rect 993 406 997 413
rect 1051 406 1055 413
rect 1070 410 1074 414
rect 1088 415 1092 419
rect 1107 415 1111 419
rect 1167 415 1171 419
rect 1125 406 1129 413
rect 1183 406 1187 413
rect 1202 410 1206 414
rect 1220 415 1224 419
rect 1239 415 1243 419
rect 1299 415 1303 419
rect 1257 406 1261 413
rect 1448 421 1452 425
rect 1492 422 1496 426
rect 1517 421 1522 425
rect 1564 422 1568 426
rect 1709 421 1713 425
rect 1753 422 1757 426
rect 1778 421 1783 425
rect 1825 422 1829 426
rect 1315 406 1319 413
rect 1336 410 1340 414
rect 1640 413 1644 417
rect 1431 404 1435 408
rect 1463 403 1467 407
rect 1482 404 1486 408
rect 1538 403 1542 407
rect 1554 404 1558 408
rect 1581 404 1585 408
rect 518 384 522 388
rect 562 384 566 388
rect 589 384 593 388
rect 634 384 638 388
rect 963 392 967 396
rect 1000 390 1004 394
rect 1020 390 1024 394
rect 1056 390 1060 394
rect 1095 392 1099 396
rect 1132 390 1136 394
rect 1152 390 1156 394
rect 1188 390 1192 394
rect 1227 392 1231 396
rect 1264 390 1268 394
rect 1284 390 1288 394
rect 1320 390 1324 394
rect 1629 397 1635 401
rect 1667 404 1671 408
rect 1724 403 1728 407
rect 1743 404 1747 408
rect 1799 403 1803 407
rect 1815 404 1819 408
rect 1842 404 1846 408
rect 779 384 783 388
rect 823 384 827 388
rect 850 384 854 388
rect 895 384 899 388
rect 1451 384 1455 388
rect 1495 384 1499 388
rect 1522 384 1526 388
rect 1567 384 1571 388
rect 1712 384 1716 388
rect 1756 384 1760 388
rect 1783 384 1787 388
rect 1828 384 1832 388
rect 705 377 709 381
rect 1638 377 1642 381
rect 139 362 143 366
rect 163 362 167 366
rect 1072 362 1076 366
rect 1096 362 1100 366
rect 918 356 922 360
rect 1851 356 1855 360
rect 159 337 163 341
rect 1092 337 1096 341
rect 174 329 178 333
rect 1107 329 1111 333
rect 801 323 805 327
rect 838 323 842 327
rect 858 323 862 327
rect 896 323 900 327
rect 1734 323 1738 327
rect 1771 323 1775 327
rect 1791 323 1795 327
rect 1829 323 1833 327
rect 139 314 143 318
rect 163 314 167 318
rect 1072 314 1076 318
rect 1096 314 1100 318
rect 795 303 799 307
rect 813 305 817 309
rect 30 293 34 297
rect 67 293 71 297
rect 87 293 91 297
rect 125 293 129 297
rect 162 293 166 297
rect 199 293 203 297
rect 219 293 223 297
rect 257 293 261 297
rect 294 293 298 297
rect 331 293 335 297
rect 351 293 355 297
rect 389 293 393 297
rect 873 305 877 309
rect 831 296 835 303
rect 889 296 893 303
rect 908 300 912 304
rect 1728 303 1732 307
rect 1746 305 1750 309
rect 963 293 967 297
rect 1000 293 1004 297
rect 1020 293 1024 297
rect 1058 293 1062 297
rect 1095 293 1099 297
rect 1132 293 1136 297
rect 1152 293 1156 297
rect 1190 293 1194 297
rect 1227 293 1231 297
rect 1264 293 1268 297
rect 1284 293 1288 297
rect 1322 293 1326 297
rect 1806 305 1810 309
rect 1764 296 1768 303
rect 1822 296 1826 303
rect 1841 300 1845 304
rect 801 282 805 286
rect 24 273 28 277
rect 42 275 46 279
rect 102 275 106 279
rect 60 266 64 273
rect 118 266 122 273
rect 137 270 141 274
rect 155 275 159 279
rect 174 275 178 279
rect 234 275 238 279
rect 192 266 196 273
rect 250 266 254 273
rect 269 270 273 274
rect 287 275 291 279
rect 306 275 310 279
rect 366 275 370 279
rect 324 266 328 273
rect 838 280 842 284
rect 858 280 862 284
rect 894 280 898 284
rect 1734 282 1738 286
rect 382 266 386 273
rect 403 270 407 274
rect 957 273 961 277
rect 975 275 979 279
rect 1035 275 1039 279
rect 993 266 997 273
rect 1051 266 1055 273
rect 1070 270 1074 274
rect 1088 275 1092 279
rect 1107 275 1111 279
rect 1167 275 1171 279
rect 1125 266 1129 273
rect 1183 266 1187 273
rect 1202 270 1206 274
rect 1220 275 1224 279
rect 1239 275 1243 279
rect 1299 275 1303 279
rect 1257 266 1261 273
rect 1771 280 1775 284
rect 1791 280 1795 284
rect 1827 280 1831 284
rect 1315 266 1319 273
rect 1336 270 1340 274
rect 30 252 34 256
rect 67 250 71 254
rect 87 250 91 254
rect 123 250 127 254
rect 162 252 166 256
rect 199 250 203 254
rect 219 250 223 254
rect 255 250 259 254
rect 294 252 298 256
rect 331 250 335 254
rect 351 250 355 254
rect 387 250 391 254
rect 963 252 967 256
rect 1000 250 1004 254
rect 1020 250 1024 254
rect 1056 250 1060 254
rect 1095 252 1099 256
rect 1132 250 1136 254
rect 1152 250 1156 254
rect 1188 250 1192 254
rect 1227 252 1231 256
rect 1264 250 1268 254
rect 1284 250 1288 254
rect 1320 250 1324 254
rect 801 237 805 241
rect 838 237 842 241
rect 858 237 862 241
rect 896 237 900 241
rect 1734 237 1738 241
rect 1771 237 1775 241
rect 1791 237 1795 241
rect 1829 237 1833 241
rect 795 217 799 221
rect 813 219 817 223
rect 30 207 34 211
rect 67 207 71 211
rect 87 207 91 211
rect 125 207 129 211
rect 162 207 166 211
rect 199 207 203 211
rect 219 207 223 211
rect 257 207 261 211
rect 294 207 298 211
rect 331 207 335 211
rect 351 207 355 211
rect 389 207 393 211
rect 873 219 877 223
rect 831 210 835 217
rect 889 210 893 217
rect 908 214 912 218
rect 930 212 934 216
rect 1728 217 1732 221
rect 1746 219 1750 223
rect 963 207 967 211
rect 1000 207 1004 211
rect 1020 207 1024 211
rect 1058 207 1062 211
rect 1095 207 1099 211
rect 1132 207 1136 211
rect 1152 207 1156 211
rect 1190 207 1194 211
rect 1227 207 1231 211
rect 1264 207 1268 211
rect 1284 207 1288 211
rect 1322 207 1326 211
rect 1806 219 1810 223
rect 1764 210 1768 217
rect 1822 210 1826 217
rect 1841 214 1845 218
rect 1863 212 1867 216
rect 801 196 805 200
rect 24 187 28 191
rect 42 189 46 193
rect 102 189 106 193
rect 60 180 64 187
rect 118 180 122 187
rect 137 184 141 188
rect 155 189 159 193
rect 174 189 178 193
rect 234 189 238 193
rect 192 180 196 187
rect 250 180 254 187
rect 269 184 273 188
rect 287 189 291 193
rect 306 189 310 193
rect 366 189 370 193
rect 324 180 328 187
rect 838 194 842 198
rect 858 194 862 198
rect 894 194 898 198
rect 1734 196 1738 200
rect 382 180 386 187
rect 403 184 407 188
rect 957 187 961 191
rect 975 189 979 193
rect 1035 189 1039 193
rect 993 180 997 187
rect 1051 180 1055 187
rect 1070 184 1074 188
rect 1088 189 1092 193
rect 1107 189 1111 193
rect 1167 189 1171 193
rect 1125 180 1129 187
rect 1183 180 1187 187
rect 1202 184 1206 188
rect 1220 189 1224 193
rect 1239 189 1243 193
rect 1299 189 1303 193
rect 1257 180 1261 187
rect 1771 194 1775 198
rect 1791 194 1795 198
rect 1827 194 1831 198
rect 1315 180 1319 187
rect 1336 184 1340 188
rect 30 166 34 170
rect 67 164 71 168
rect 87 164 91 168
rect 123 164 127 168
rect 162 166 166 170
rect 199 164 203 168
rect 219 164 223 168
rect 255 164 259 168
rect 294 166 298 170
rect 331 164 335 168
rect 351 164 355 168
rect 387 164 391 168
rect 963 166 967 170
rect 1000 164 1004 168
rect 1020 164 1024 168
rect 1056 164 1060 168
rect 1095 166 1099 170
rect 1132 164 1136 168
rect 1152 164 1156 168
rect 1188 164 1192 168
rect 1227 166 1231 170
rect 1264 164 1268 168
rect 1284 164 1288 168
rect 1320 164 1324 168
rect 256 136 260 140
rect 280 136 284 140
rect 1189 136 1193 140
rect 1213 136 1217 140
rect 276 111 280 115
rect 1209 111 1213 115
rect 291 103 295 107
rect 1224 103 1228 107
rect 256 88 260 92
rect 280 88 284 92
rect 1189 88 1193 92
rect 1213 88 1217 92
rect 30 67 34 71
rect 67 67 71 71
rect 87 67 91 71
rect 125 67 129 71
rect 162 67 166 71
rect 199 67 203 71
rect 219 67 223 71
rect 257 67 261 71
rect 294 67 298 71
rect 331 67 335 71
rect 351 67 355 71
rect 389 67 393 71
rect 963 67 967 71
rect 1000 67 1004 71
rect 1020 67 1024 71
rect 1058 67 1062 71
rect 1095 67 1099 71
rect 1132 67 1136 71
rect 1152 67 1156 71
rect 1190 67 1194 71
rect 1227 67 1231 71
rect 1264 67 1268 71
rect 1284 67 1288 71
rect 1322 67 1326 71
rect 24 47 28 51
rect 42 49 46 53
rect 102 49 106 53
rect 60 40 64 47
rect 118 40 122 47
rect 137 44 141 48
rect 155 49 159 53
rect 174 49 178 53
rect 234 49 238 53
rect 192 40 196 47
rect 250 40 254 47
rect 269 44 273 48
rect 287 49 291 53
rect 306 49 310 53
rect 366 49 370 53
rect 324 40 328 47
rect 382 40 386 47
rect 403 44 407 48
rect 957 47 961 51
rect 975 49 979 53
rect 1035 49 1039 53
rect 993 40 997 47
rect 1051 40 1055 47
rect 1070 44 1074 48
rect 1088 49 1092 53
rect 1107 49 1111 53
rect 1167 49 1171 53
rect 1125 40 1129 47
rect 1183 40 1187 47
rect 1202 44 1206 48
rect 1220 49 1224 53
rect 1239 49 1243 53
rect 1299 49 1303 53
rect 1257 40 1261 47
rect 1315 40 1319 47
rect 1336 44 1340 48
rect 30 26 34 30
rect 67 24 71 28
rect 87 24 91 28
rect 123 24 127 28
rect 162 26 166 30
rect 199 24 203 28
rect 219 24 223 28
rect 255 24 259 28
rect 294 26 298 30
rect 331 24 335 28
rect 351 24 355 28
rect 387 24 391 28
rect 963 26 967 30
rect 1000 24 1004 28
rect 1020 24 1024 28
rect 1056 24 1060 28
rect 1095 26 1099 30
rect 1132 24 1136 28
rect 1152 24 1156 28
rect 1188 24 1192 28
rect 1227 26 1231 30
rect 1264 24 1268 28
rect 1284 24 1288 28
rect 1320 24 1324 28
<< metal1 >>
rect 483 1962 498 1966
rect 502 1962 534 1966
rect 538 1962 601 1966
rect 605 1962 630 1966
rect 634 1962 666 1966
rect 670 1962 733 1966
rect 737 1962 762 1966
rect 766 1962 798 1966
rect 802 1962 865 1966
rect 869 1962 894 1966
rect 898 1962 930 1966
rect 934 1962 997 1966
rect 1001 1962 1017 1966
rect 1416 1962 1431 1966
rect 1435 1962 1467 1966
rect 1471 1962 1534 1966
rect 1538 1962 1563 1966
rect 1567 1962 1599 1966
rect 1603 1962 1666 1966
rect 1670 1962 1695 1966
rect 1699 1962 1731 1966
rect 1735 1962 1798 1966
rect 1802 1962 1827 1966
rect 1831 1962 1863 1966
rect 1867 1962 1930 1966
rect 1934 1962 1950 1966
rect 423 1955 522 1959
rect 526 1955 550 1959
rect 554 1955 580 1959
rect 584 1955 617 1959
rect 621 1955 654 1959
rect 658 1955 682 1959
rect 686 1955 712 1959
rect 716 1955 749 1959
rect 753 1955 786 1959
rect 790 1955 814 1959
rect 818 1955 844 1959
rect 848 1955 881 1959
rect 885 1955 918 1959
rect 922 1955 946 1959
rect 950 1955 976 1959
rect 980 1955 1013 1959
rect 1356 1955 1455 1959
rect 1459 1955 1483 1959
rect 1487 1955 1513 1959
rect 1517 1955 1550 1959
rect 1554 1955 1587 1959
rect 1591 1955 1615 1959
rect 1619 1955 1645 1959
rect 1649 1955 1682 1959
rect 1686 1955 1719 1959
rect 1723 1955 1747 1959
rect 1751 1955 1777 1959
rect 1781 1955 1814 1959
rect 1818 1955 1851 1959
rect 1855 1955 1879 1959
rect 1883 1955 1909 1959
rect 1913 1955 1946 1959
rect 492 1945 495 1955
rect 513 1945 516 1955
rect 529 1945 532 1955
rect 543 1948 548 1952
rect 552 1948 559 1952
rect 571 1945 574 1955
rect 587 1945 590 1955
rect 608 1945 611 1955
rect 624 1945 627 1955
rect 645 1945 648 1955
rect 661 1945 664 1955
rect 675 1948 680 1952
rect 684 1948 691 1952
rect 703 1945 706 1955
rect 719 1945 722 1955
rect 740 1945 743 1955
rect 756 1945 759 1955
rect 777 1945 780 1955
rect 793 1945 796 1955
rect 807 1948 812 1952
rect 816 1948 823 1952
rect 835 1945 838 1955
rect 851 1945 854 1955
rect 872 1945 875 1955
rect 888 1945 891 1955
rect 909 1945 912 1955
rect 925 1945 928 1955
rect 939 1948 944 1952
rect 948 1948 955 1952
rect 967 1945 970 1955
rect 983 1945 986 1955
rect 1004 1945 1007 1955
rect 1425 1945 1428 1955
rect 1446 1945 1449 1955
rect 1462 1945 1465 1955
rect 1476 1948 1481 1952
rect 1485 1948 1492 1952
rect 1504 1945 1507 1955
rect 1520 1945 1523 1955
rect 1541 1945 1544 1955
rect 1557 1945 1560 1955
rect 1578 1945 1581 1955
rect 1594 1945 1597 1955
rect 1608 1948 1613 1952
rect 1617 1948 1624 1952
rect 1636 1945 1639 1955
rect 1652 1945 1655 1955
rect 1673 1945 1676 1955
rect 1689 1945 1692 1955
rect 1710 1945 1713 1955
rect 1726 1945 1729 1955
rect 1740 1948 1745 1952
rect 1749 1948 1756 1952
rect 1768 1945 1771 1955
rect 1784 1945 1787 1955
rect 1805 1945 1808 1955
rect 1821 1945 1824 1955
rect 1842 1945 1845 1955
rect 1858 1945 1861 1955
rect 1872 1948 1877 1952
rect 1881 1948 1888 1952
rect 1900 1945 1903 1955
rect 1916 1945 1919 1955
rect 1937 1945 1940 1955
rect 149 1929 158 1933
rect 162 1929 194 1933
rect 198 1929 261 1933
rect 265 1929 477 1933
rect 509 1931 514 1934
rect 518 1931 542 1934
rect 567 1931 574 1934
rect 578 1931 600 1934
rect 149 1922 182 1926
rect 186 1922 210 1926
rect 214 1922 240 1926
rect 244 1922 277 1926
rect 281 1922 417 1926
rect 152 1912 155 1922
rect 173 1912 176 1922
rect 189 1912 192 1922
rect 203 1915 208 1919
rect 212 1915 219 1919
rect 231 1912 234 1922
rect 247 1912 250 1922
rect 268 1912 271 1922
rect 525 1921 532 1924
rect 536 1925 555 1928
rect 555 1918 558 1924
rect 583 1921 590 1924
rect 594 1925 611 1928
rect 641 1931 646 1934
rect 650 1931 674 1934
rect 699 1931 706 1934
rect 710 1931 732 1934
rect 657 1921 664 1924
rect 668 1925 687 1928
rect 687 1918 690 1924
rect 715 1921 722 1924
rect 726 1925 743 1928
rect 773 1931 778 1934
rect 782 1931 806 1934
rect 831 1931 838 1934
rect 842 1931 864 1934
rect 789 1921 796 1924
rect 800 1925 819 1928
rect 819 1918 822 1924
rect 847 1921 854 1924
rect 858 1925 875 1928
rect 905 1931 910 1934
rect 914 1931 938 1934
rect 963 1931 970 1934
rect 974 1931 996 1934
rect 1082 1929 1091 1933
rect 1095 1929 1127 1933
rect 1131 1929 1194 1933
rect 1198 1929 1410 1933
rect 921 1921 928 1924
rect 932 1925 951 1928
rect 147 1895 156 1899
rect 169 1898 174 1901
rect 178 1898 202 1901
rect 227 1898 234 1901
rect 238 1898 260 1901
rect 492 1902 495 1914
rect 513 1902 516 1914
rect 529 1902 532 1914
rect 543 1905 555 1908
rect 571 1902 574 1914
rect 587 1902 590 1914
rect 608 1902 611 1914
rect 624 1902 627 1914
rect 645 1902 648 1914
rect 661 1902 664 1914
rect 675 1905 687 1908
rect 703 1902 706 1914
rect 719 1902 722 1914
rect 740 1902 743 1914
rect 756 1902 759 1914
rect 777 1902 780 1914
rect 793 1902 796 1914
rect 807 1905 819 1908
rect 835 1902 838 1914
rect 851 1902 854 1914
rect 872 1902 875 1914
rect 951 1918 954 1924
rect 979 1921 986 1924
rect 990 1925 1007 1928
rect 1442 1931 1447 1934
rect 1451 1931 1475 1934
rect 1500 1931 1507 1934
rect 1511 1931 1533 1934
rect 1082 1922 1115 1926
rect 1119 1922 1143 1926
rect 1147 1922 1173 1926
rect 1177 1922 1210 1926
rect 1214 1922 1350 1926
rect 888 1902 891 1914
rect 909 1902 912 1914
rect 925 1902 928 1914
rect 939 1905 951 1908
rect 967 1902 970 1914
rect 983 1902 986 1914
rect 1004 1902 1007 1914
rect 1085 1912 1088 1922
rect 1106 1912 1109 1922
rect 1122 1912 1125 1922
rect 1136 1915 1141 1919
rect 1145 1915 1152 1919
rect 1164 1912 1167 1922
rect 1180 1912 1183 1922
rect 1201 1912 1204 1922
rect 1458 1921 1465 1924
rect 1469 1925 1488 1928
rect 1488 1918 1491 1924
rect 1516 1921 1523 1924
rect 1527 1925 1544 1928
rect 1574 1931 1579 1934
rect 1583 1931 1607 1934
rect 1632 1931 1639 1934
rect 1643 1931 1665 1934
rect 1590 1921 1597 1924
rect 1601 1925 1620 1928
rect 1620 1918 1623 1924
rect 1648 1921 1655 1924
rect 1659 1925 1676 1928
rect 1706 1931 1711 1934
rect 1715 1931 1739 1934
rect 1764 1931 1771 1934
rect 1775 1931 1797 1934
rect 1722 1921 1729 1924
rect 1733 1925 1752 1928
rect 1752 1918 1755 1924
rect 1780 1921 1787 1924
rect 1791 1925 1808 1928
rect 1838 1931 1843 1934
rect 1847 1931 1871 1934
rect 1896 1931 1903 1934
rect 1907 1931 1929 1934
rect 1854 1921 1861 1924
rect 1865 1925 1884 1928
rect 435 1898 522 1902
rect 526 1898 550 1902
rect 554 1898 580 1902
rect 584 1898 654 1902
rect 658 1898 682 1902
rect 686 1898 712 1902
rect 716 1898 786 1902
rect 790 1898 814 1902
rect 818 1898 844 1902
rect 848 1898 918 1902
rect 922 1898 946 1902
rect 950 1898 976 1902
rect 980 1898 1017 1902
rect 185 1888 192 1891
rect 196 1892 215 1895
rect 215 1885 218 1891
rect 243 1888 250 1891
rect 254 1892 269 1895
rect 1080 1895 1089 1899
rect 1102 1898 1107 1901
rect 1111 1898 1135 1901
rect 1160 1898 1167 1901
rect 1171 1898 1193 1901
rect 1425 1902 1428 1914
rect 1446 1902 1449 1914
rect 1462 1902 1465 1914
rect 1476 1905 1488 1908
rect 1504 1902 1507 1914
rect 1520 1902 1523 1914
rect 1541 1902 1544 1914
rect 1557 1902 1560 1914
rect 1578 1902 1581 1914
rect 1594 1902 1597 1914
rect 1608 1905 1620 1908
rect 1636 1902 1639 1914
rect 1652 1902 1655 1914
rect 1673 1902 1676 1914
rect 1689 1902 1692 1914
rect 1710 1902 1713 1914
rect 1726 1902 1729 1914
rect 1740 1905 1752 1908
rect 1768 1902 1771 1914
rect 1784 1902 1787 1914
rect 1805 1902 1808 1914
rect 1884 1918 1887 1924
rect 1912 1921 1919 1924
rect 1923 1925 1940 1928
rect 1821 1902 1824 1914
rect 1842 1902 1845 1914
rect 1858 1902 1861 1914
rect 1872 1905 1884 1908
rect 1900 1902 1903 1914
rect 1916 1902 1919 1914
rect 1937 1902 1940 1914
rect 1368 1898 1455 1902
rect 1459 1898 1483 1902
rect 1487 1898 1513 1902
rect 1517 1898 1587 1902
rect 1591 1898 1615 1902
rect 1619 1898 1645 1902
rect 1649 1898 1719 1902
rect 1723 1898 1747 1902
rect 1751 1898 1777 1902
rect 1781 1898 1851 1902
rect 1855 1898 1879 1902
rect 1883 1898 1909 1902
rect 1913 1898 1950 1902
rect 471 1891 498 1895
rect 502 1891 549 1895
rect 553 1891 599 1895
rect 603 1891 630 1895
rect 634 1891 681 1895
rect 685 1891 731 1895
rect 735 1891 762 1895
rect 766 1891 813 1895
rect 817 1891 863 1895
rect 867 1891 894 1895
rect 898 1891 945 1895
rect 949 1891 995 1895
rect 999 1891 1017 1895
rect 1118 1888 1125 1891
rect 1129 1892 1148 1895
rect 152 1869 155 1881
rect 173 1869 176 1881
rect 189 1869 192 1881
rect 203 1872 215 1875
rect 231 1869 234 1881
rect 247 1869 250 1881
rect 268 1869 271 1881
rect 423 1878 496 1882
rect 500 1878 512 1882
rect 516 1878 530 1882
rect 534 1878 541 1882
rect 545 1878 547 1882
rect 551 1878 566 1882
rect 570 1878 603 1882
rect 607 1878 608 1882
rect 612 1878 620 1882
rect 624 1878 648 1882
rect 652 1878 664 1882
rect 668 1878 688 1882
rect 692 1878 742 1882
rect 746 1878 769 1882
rect 773 1878 823 1882
rect 827 1878 846 1882
rect 1148 1885 1151 1891
rect 1176 1888 1183 1891
rect 1187 1892 1202 1895
rect 1404 1891 1431 1895
rect 1435 1891 1482 1895
rect 1486 1891 1532 1895
rect 1536 1891 1563 1895
rect 1567 1891 1614 1895
rect 1618 1891 1664 1895
rect 1668 1891 1695 1895
rect 1699 1891 1746 1895
rect 1750 1891 1796 1895
rect 1800 1891 1827 1895
rect 1831 1891 1878 1895
rect 1882 1891 1928 1895
rect 1932 1891 1950 1895
rect 459 1871 523 1875
rect 527 1871 554 1875
rect 558 1871 576 1875
rect 580 1871 641 1875
rect 645 1871 659 1875
rect 671 1874 674 1878
rect 149 1865 182 1869
rect 186 1865 210 1869
rect 214 1865 240 1869
rect 244 1865 429 1869
rect 149 1858 158 1862
rect 162 1858 209 1862
rect 213 1858 259 1862
rect 263 1858 465 1862
rect 566 1864 569 1868
rect 593 1864 594 1868
rect 638 1864 640 1868
rect 680 1861 683 1866
rect 695 1868 698 1878
rect 725 1874 728 1878
rect 752 1874 755 1878
rect 147 1842 163 1846
rect 272 1844 276 1848
rect 288 1844 292 1848
rect 296 1844 498 1848
rect 506 1847 509 1853
rect 513 1847 516 1853
rect 506 1844 516 1847
rect 506 1839 509 1844
rect 155 1835 159 1839
rect 171 1835 292 1839
rect 513 1839 516 1844
rect 522 1849 525 1853
rect 522 1845 524 1849
rect 528 1845 530 1849
rect 538 1848 541 1853
rect 566 1850 569 1853
rect 538 1846 549 1848
rect 522 1839 525 1845
rect 538 1844 544 1846
rect 538 1839 541 1844
rect 548 1844 549 1846
rect 567 1846 569 1850
rect 566 1839 569 1846
rect 669 1857 672 1860
rect 711 1857 714 1860
rect 582 1849 585 1853
rect 592 1849 595 1853
rect 592 1845 601 1849
rect 613 1848 616 1853
rect 638 1849 641 1853
rect 582 1839 585 1845
rect 592 1839 595 1845
rect 613 1844 614 1848
rect 618 1844 621 1847
rect 640 1845 641 1849
rect 656 1848 659 1853
rect 680 1852 683 1857
rect 688 1853 699 1856
rect 711 1854 719 1857
rect 613 1839 616 1844
rect 638 1839 641 1845
rect 656 1839 659 1844
rect 142 1827 158 1831
rect 162 1827 225 1831
rect 229 1827 261 1831
rect 265 1827 477 1831
rect 558 1826 559 1830
rect 583 1827 584 1831
rect 630 1826 631 1830
rect 146 1820 179 1824
rect 183 1820 209 1824
rect 213 1820 237 1824
rect 241 1820 417 1824
rect 152 1810 155 1820
rect 173 1810 176 1820
rect 189 1810 192 1820
rect 204 1813 211 1817
rect 215 1813 220 1817
rect 231 1810 234 1820
rect 247 1810 250 1820
rect 268 1810 271 1820
rect 447 1819 511 1823
rect 515 1819 570 1823
rect 574 1819 595 1823
rect 599 1819 626 1823
rect 630 1819 659 1823
rect 671 1816 674 1848
rect 688 1847 691 1853
rect 711 1848 714 1854
rect 723 1849 726 1852
rect 734 1852 737 1866
rect 761 1861 764 1866
rect 776 1868 779 1878
rect 806 1874 809 1878
rect 745 1857 746 1860
rect 750 1857 753 1860
rect 1085 1869 1088 1881
rect 1106 1869 1109 1881
rect 1122 1869 1125 1881
rect 1136 1872 1148 1875
rect 1164 1869 1167 1881
rect 1180 1869 1183 1881
rect 1201 1869 1204 1881
rect 1356 1878 1429 1882
rect 1433 1878 1445 1882
rect 1449 1878 1463 1882
rect 1467 1878 1474 1882
rect 1478 1878 1480 1882
rect 1484 1878 1499 1882
rect 1503 1878 1536 1882
rect 1540 1878 1541 1882
rect 1545 1878 1553 1882
rect 1557 1878 1581 1882
rect 1585 1878 1597 1882
rect 1601 1878 1621 1882
rect 1625 1878 1675 1882
rect 1679 1878 1702 1882
rect 1706 1878 1756 1882
rect 1760 1878 1779 1882
rect 1392 1871 1456 1875
rect 1460 1871 1487 1875
rect 1491 1871 1509 1875
rect 1513 1871 1574 1875
rect 1578 1871 1592 1875
rect 1604 1874 1607 1878
rect 792 1857 795 1860
rect 734 1849 742 1852
rect 761 1852 764 1857
rect 734 1844 737 1849
rect 742 1845 746 1849
rect 769 1853 780 1856
rect 792 1854 800 1857
rect 686 1838 691 1843
rect 695 1816 698 1844
rect 725 1816 728 1840
rect 752 1816 755 1848
rect 769 1847 772 1853
rect 792 1848 795 1854
rect 804 1849 807 1852
rect 815 1852 818 1866
rect 1082 1865 1115 1869
rect 1119 1865 1143 1869
rect 1147 1865 1173 1869
rect 1177 1865 1362 1869
rect 1082 1858 1091 1862
rect 1095 1858 1142 1862
rect 1146 1858 1192 1862
rect 1196 1858 1398 1862
rect 1499 1864 1502 1868
rect 1526 1864 1527 1868
rect 1571 1864 1573 1868
rect 1613 1861 1616 1866
rect 1628 1868 1631 1878
rect 1658 1874 1661 1878
rect 1685 1874 1688 1878
rect 815 1849 827 1852
rect 815 1844 818 1849
rect 767 1838 772 1843
rect 776 1816 779 1844
rect 1080 1842 1096 1846
rect 1205 1844 1209 1848
rect 1221 1844 1225 1848
rect 1229 1844 1431 1848
rect 1439 1847 1442 1853
rect 1446 1847 1449 1853
rect 1439 1844 1449 1847
rect 806 1816 809 1840
rect 1439 1839 1442 1844
rect 1088 1835 1092 1839
rect 1104 1835 1225 1839
rect 1446 1839 1449 1844
rect 1455 1849 1458 1853
rect 1455 1845 1457 1849
rect 1461 1845 1463 1849
rect 1471 1848 1474 1853
rect 1499 1850 1502 1853
rect 1471 1846 1482 1848
rect 1455 1839 1458 1845
rect 1471 1844 1477 1846
rect 1471 1839 1474 1844
rect 1481 1844 1482 1846
rect 1500 1846 1502 1850
rect 1499 1839 1502 1846
rect 1602 1857 1605 1860
rect 1644 1857 1647 1860
rect 1515 1849 1518 1853
rect 1525 1849 1528 1853
rect 1525 1845 1534 1849
rect 1546 1848 1549 1853
rect 1571 1849 1574 1853
rect 1515 1839 1518 1845
rect 1525 1839 1528 1845
rect 1546 1844 1547 1848
rect 1551 1844 1554 1847
rect 1573 1845 1574 1849
rect 1589 1848 1592 1853
rect 1613 1852 1616 1857
rect 1621 1853 1632 1856
rect 1644 1854 1652 1857
rect 1546 1839 1549 1844
rect 1571 1839 1574 1845
rect 1589 1839 1592 1844
rect 1075 1827 1091 1831
rect 1095 1827 1158 1831
rect 1162 1827 1194 1831
rect 1198 1827 1410 1831
rect 1491 1826 1492 1830
rect 1516 1827 1517 1831
rect 1563 1826 1564 1830
rect 1079 1820 1112 1824
rect 1116 1820 1142 1824
rect 1146 1820 1170 1824
rect 1174 1820 1350 1824
rect 435 1812 497 1816
rect 501 1812 503 1816
rect 507 1812 511 1816
rect 515 1812 529 1816
rect 533 1812 538 1816
rect 542 1812 547 1816
rect 551 1812 570 1816
rect 574 1812 604 1816
rect 608 1812 619 1816
rect 623 1812 647 1816
rect 651 1812 664 1816
rect 668 1812 688 1816
rect 692 1812 742 1816
rect 749 1812 769 1816
rect 773 1812 823 1816
rect 163 1796 185 1799
rect 189 1796 196 1799
rect 447 1805 511 1809
rect 515 1805 570 1809
rect 574 1805 595 1809
rect 599 1805 626 1809
rect 630 1805 659 1809
rect 221 1796 245 1799
rect 249 1796 254 1799
rect 558 1798 559 1802
rect 583 1797 584 1801
rect 630 1798 631 1802
rect 267 1793 276 1797
rect 154 1790 169 1793
rect 208 1790 227 1793
rect 173 1786 180 1789
rect 205 1783 208 1789
rect 231 1786 238 1789
rect 506 1784 509 1789
rect 513 1784 516 1789
rect 496 1781 498 1784
rect 506 1781 516 1784
rect 152 1767 155 1779
rect 173 1767 176 1779
rect 189 1767 192 1779
rect 208 1770 220 1773
rect 231 1767 234 1779
rect 247 1767 250 1779
rect 268 1767 271 1779
rect 506 1775 509 1781
rect 513 1775 516 1781
rect 522 1783 525 1789
rect 538 1784 541 1789
rect 522 1779 524 1783
rect 528 1779 530 1783
rect 538 1782 544 1784
rect 548 1782 549 1784
rect 538 1780 549 1782
rect 566 1782 569 1789
rect 522 1775 525 1779
rect 538 1775 541 1780
rect 567 1778 569 1782
rect 566 1775 569 1778
rect 582 1783 585 1789
rect 592 1783 595 1789
rect 613 1784 616 1789
rect 592 1779 601 1783
rect 613 1780 614 1784
rect 618 1781 621 1784
rect 638 1783 641 1789
rect 656 1784 659 1789
rect 695 1792 698 1812
rect 776 1792 779 1812
rect 1085 1810 1088 1820
rect 1106 1810 1109 1820
rect 1122 1810 1125 1820
rect 1137 1813 1144 1817
rect 1148 1813 1153 1817
rect 1164 1810 1167 1820
rect 1180 1810 1183 1820
rect 1201 1810 1204 1820
rect 1380 1819 1444 1823
rect 1448 1819 1503 1823
rect 1507 1819 1528 1823
rect 1532 1819 1559 1823
rect 1563 1819 1592 1823
rect 1604 1816 1607 1848
rect 1621 1847 1624 1853
rect 1644 1848 1647 1854
rect 1656 1849 1659 1852
rect 1667 1852 1670 1866
rect 1694 1861 1697 1866
rect 1709 1868 1712 1878
rect 1739 1874 1742 1878
rect 1678 1857 1679 1860
rect 1683 1857 1686 1860
rect 1725 1857 1728 1860
rect 1667 1849 1675 1852
rect 1694 1852 1697 1857
rect 1667 1844 1670 1849
rect 1675 1845 1679 1849
rect 1702 1853 1713 1856
rect 1725 1854 1733 1857
rect 1619 1838 1624 1843
rect 1628 1816 1631 1844
rect 1658 1816 1661 1840
rect 1685 1816 1688 1848
rect 1702 1847 1705 1853
rect 1725 1848 1728 1854
rect 1737 1849 1740 1852
rect 1748 1852 1751 1866
rect 1748 1849 1760 1852
rect 1748 1844 1751 1849
rect 1700 1838 1705 1843
rect 1709 1816 1712 1844
rect 1739 1816 1742 1840
rect 1368 1812 1430 1816
rect 1434 1812 1436 1816
rect 1440 1812 1444 1816
rect 1448 1812 1462 1816
rect 1466 1812 1471 1816
rect 1475 1812 1480 1816
rect 1484 1812 1503 1816
rect 1507 1812 1537 1816
rect 1541 1812 1552 1816
rect 1556 1812 1580 1816
rect 1584 1812 1597 1816
rect 1601 1812 1621 1816
rect 1625 1812 1675 1816
rect 1682 1812 1702 1816
rect 1706 1812 1756 1816
rect 1096 1796 1118 1799
rect 1122 1796 1129 1799
rect 1380 1805 1444 1809
rect 1448 1805 1503 1809
rect 1507 1805 1528 1809
rect 1532 1805 1559 1809
rect 1563 1805 1592 1809
rect 1154 1796 1178 1799
rect 1182 1796 1187 1799
rect 1491 1798 1492 1802
rect 1516 1797 1517 1801
rect 1563 1798 1564 1802
rect 1200 1793 1209 1797
rect 1087 1790 1102 1793
rect 582 1775 585 1779
rect 592 1775 595 1779
rect 613 1775 616 1780
rect 640 1779 641 1783
rect 638 1775 641 1779
rect 656 1775 659 1780
rect 686 1779 691 1784
rect 695 1780 696 1783
rect 711 1782 714 1788
rect 711 1779 719 1782
rect 766 1779 771 1784
rect 775 1780 777 1783
rect 792 1782 795 1788
rect 1141 1790 1160 1793
rect 1106 1786 1113 1789
rect 1138 1783 1141 1789
rect 792 1779 800 1782
rect 1164 1786 1171 1789
rect 1439 1784 1442 1789
rect 1446 1784 1449 1789
rect 1429 1781 1431 1784
rect 1439 1781 1449 1784
rect 711 1776 714 1779
rect 792 1776 795 1779
rect 142 1763 179 1767
rect 183 1763 209 1767
rect 213 1763 237 1767
rect 241 1763 429 1767
rect 566 1760 569 1764
rect 593 1760 594 1764
rect 638 1760 640 1764
rect 142 1756 160 1760
rect 164 1756 210 1760
rect 214 1756 261 1760
rect 265 1756 465 1760
rect 511 1753 523 1757
rect 527 1753 554 1757
rect 558 1753 576 1757
rect 580 1753 641 1757
rect 645 1753 659 1757
rect 695 1750 698 1768
rect 776 1750 779 1768
rect 1085 1767 1088 1779
rect 1106 1767 1109 1779
rect 1122 1767 1125 1779
rect 1141 1770 1153 1773
rect 1164 1767 1167 1779
rect 1180 1767 1183 1779
rect 1201 1767 1204 1779
rect 1439 1775 1442 1781
rect 1446 1775 1449 1781
rect 1455 1783 1458 1789
rect 1471 1784 1474 1789
rect 1455 1779 1457 1783
rect 1461 1779 1463 1783
rect 1471 1782 1477 1784
rect 1481 1782 1482 1784
rect 1471 1780 1482 1782
rect 1499 1782 1502 1789
rect 1455 1775 1458 1779
rect 1471 1775 1474 1780
rect 1500 1778 1502 1782
rect 1499 1775 1502 1778
rect 1515 1783 1518 1789
rect 1525 1783 1528 1789
rect 1546 1784 1549 1789
rect 1525 1779 1534 1783
rect 1546 1780 1547 1784
rect 1551 1781 1554 1784
rect 1571 1783 1574 1789
rect 1589 1784 1592 1789
rect 1628 1792 1631 1812
rect 1709 1792 1712 1812
rect 1515 1775 1518 1779
rect 1525 1775 1528 1779
rect 1546 1775 1549 1780
rect 1573 1779 1574 1783
rect 1571 1775 1574 1779
rect 1589 1775 1592 1780
rect 1619 1779 1624 1784
rect 1628 1780 1629 1783
rect 1644 1782 1647 1788
rect 1644 1779 1652 1782
rect 1699 1779 1704 1784
rect 1708 1780 1710 1783
rect 1725 1782 1728 1788
rect 1725 1779 1733 1782
rect 1644 1776 1647 1779
rect 1725 1776 1728 1779
rect 1075 1763 1112 1767
rect 1116 1763 1142 1767
rect 1146 1763 1170 1767
rect 1174 1763 1362 1767
rect 1499 1760 1502 1764
rect 1526 1760 1527 1764
rect 1571 1760 1573 1764
rect 1075 1756 1093 1760
rect 1097 1756 1143 1760
rect 1147 1756 1194 1760
rect 1198 1756 1398 1760
rect 1444 1753 1456 1757
rect 1460 1753 1487 1757
rect 1491 1753 1509 1757
rect 1513 1753 1574 1757
rect 1578 1753 1592 1757
rect 1628 1750 1631 1768
rect 1709 1750 1712 1768
rect 423 1746 496 1750
rect 500 1746 512 1750
rect 516 1746 530 1750
rect 534 1746 541 1750
rect 545 1746 547 1750
rect 551 1746 566 1750
rect 570 1746 603 1750
rect 607 1746 608 1750
rect 612 1746 620 1750
rect 624 1746 648 1750
rect 652 1746 664 1750
rect 668 1746 688 1750
rect 692 1746 742 1750
rect 746 1746 769 1750
rect 773 1746 831 1750
rect 835 1746 846 1750
rect 1356 1746 1429 1750
rect 1433 1746 1445 1750
rect 1449 1746 1463 1750
rect 1467 1746 1474 1750
rect 1478 1746 1480 1750
rect 1484 1746 1499 1750
rect 1503 1746 1536 1750
rect 1540 1746 1541 1750
rect 1545 1746 1553 1750
rect 1557 1746 1581 1750
rect 1585 1746 1597 1750
rect 1601 1746 1621 1750
rect 1625 1746 1675 1750
rect 1679 1746 1702 1750
rect 1706 1746 1764 1750
rect 1768 1746 1779 1750
rect 459 1739 507 1743
rect 511 1739 523 1743
rect 527 1739 554 1743
rect 558 1739 576 1743
rect 580 1739 641 1743
rect 645 1739 659 1743
rect 695 1736 698 1746
rect 725 1742 728 1746
rect 776 1742 779 1746
rect 566 1732 569 1736
rect 593 1732 594 1736
rect 638 1732 640 1736
rect 495 1712 498 1715
rect 506 1715 509 1721
rect 513 1715 516 1721
rect 506 1712 516 1715
rect 506 1707 509 1712
rect 513 1707 516 1712
rect 522 1717 525 1721
rect 522 1713 524 1717
rect 528 1713 530 1717
rect 538 1716 541 1721
rect 566 1718 569 1721
rect 538 1714 549 1716
rect 522 1707 525 1713
rect 538 1712 544 1714
rect 538 1707 541 1712
rect 548 1712 549 1714
rect 567 1714 569 1718
rect 566 1707 569 1714
rect 711 1725 714 1728
rect 582 1717 585 1721
rect 592 1717 595 1721
rect 592 1713 601 1717
rect 613 1716 616 1721
rect 638 1717 641 1721
rect 582 1707 585 1713
rect 592 1707 595 1713
rect 613 1712 614 1716
rect 618 1712 621 1715
rect 640 1713 641 1717
rect 656 1716 659 1721
rect 688 1721 699 1724
rect 711 1722 719 1725
rect 613 1707 616 1712
rect 638 1707 641 1713
rect 688 1715 691 1721
rect 711 1716 714 1722
rect 723 1717 726 1720
rect 734 1720 737 1734
rect 785 1729 788 1734
rect 800 1736 803 1746
rect 830 1742 833 1746
rect 769 1725 770 1728
rect 774 1725 777 1728
rect 1392 1739 1440 1743
rect 1444 1739 1456 1743
rect 1460 1739 1487 1743
rect 1491 1739 1509 1743
rect 1513 1739 1574 1743
rect 1578 1739 1592 1743
rect 1628 1736 1631 1746
rect 1658 1742 1661 1746
rect 1709 1742 1712 1746
rect 816 1725 819 1728
rect 742 1720 747 1725
rect 785 1720 788 1725
rect 734 1717 742 1720
rect 656 1707 659 1712
rect 734 1712 737 1717
rect 793 1721 804 1724
rect 816 1722 824 1725
rect 686 1706 691 1711
rect 558 1694 559 1698
rect 583 1695 584 1699
rect 630 1694 631 1698
rect 447 1687 511 1691
rect 515 1687 570 1691
rect 574 1687 595 1691
rect 599 1687 626 1691
rect 630 1687 659 1691
rect 695 1684 698 1712
rect 725 1684 728 1708
rect 776 1684 779 1716
rect 793 1715 796 1721
rect 816 1716 819 1722
rect 828 1717 831 1720
rect 839 1720 842 1734
rect 1499 1732 1502 1736
rect 1526 1732 1527 1736
rect 1571 1732 1573 1736
rect 839 1717 845 1720
rect 839 1712 842 1717
rect 1428 1712 1431 1715
rect 1439 1715 1442 1721
rect 1446 1715 1449 1721
rect 1439 1712 1449 1715
rect 791 1706 796 1711
rect 800 1684 803 1712
rect 830 1684 833 1708
rect 1439 1707 1442 1712
rect 1446 1707 1449 1712
rect 1455 1717 1458 1721
rect 1455 1713 1457 1717
rect 1461 1713 1463 1717
rect 1471 1716 1474 1721
rect 1499 1718 1502 1721
rect 1471 1714 1482 1716
rect 1455 1707 1458 1713
rect 1471 1712 1477 1714
rect 1471 1707 1474 1712
rect 1481 1712 1482 1714
rect 1500 1714 1502 1718
rect 1499 1707 1502 1714
rect 1644 1725 1647 1728
rect 1515 1717 1518 1721
rect 1525 1717 1528 1721
rect 1525 1713 1534 1717
rect 1546 1716 1549 1721
rect 1571 1717 1574 1721
rect 1515 1707 1518 1713
rect 1525 1707 1528 1713
rect 1546 1712 1547 1716
rect 1551 1712 1554 1715
rect 1573 1713 1574 1717
rect 1589 1716 1592 1721
rect 1621 1721 1632 1724
rect 1644 1722 1652 1725
rect 1546 1707 1549 1712
rect 1571 1707 1574 1713
rect 1621 1715 1624 1721
rect 1644 1716 1647 1722
rect 1656 1717 1659 1720
rect 1667 1720 1670 1734
rect 1718 1729 1721 1734
rect 1733 1736 1736 1746
rect 1763 1742 1766 1746
rect 1702 1725 1703 1728
rect 1707 1725 1710 1728
rect 1749 1725 1752 1728
rect 1675 1720 1680 1725
rect 1718 1720 1721 1725
rect 1667 1717 1675 1720
rect 1589 1707 1592 1712
rect 1667 1712 1670 1717
rect 1726 1721 1737 1724
rect 1749 1722 1757 1725
rect 1619 1706 1624 1711
rect 1491 1694 1492 1698
rect 1516 1695 1517 1699
rect 1563 1694 1564 1698
rect 1380 1687 1444 1691
rect 1448 1687 1503 1691
rect 1507 1687 1528 1691
rect 1532 1687 1559 1691
rect 1563 1687 1592 1691
rect 1628 1684 1631 1712
rect 1658 1684 1661 1708
rect 1709 1684 1712 1716
rect 1726 1715 1729 1721
rect 1749 1716 1752 1722
rect 1761 1717 1764 1720
rect 1772 1720 1775 1734
rect 1772 1717 1778 1720
rect 1772 1712 1775 1717
rect 1724 1706 1729 1711
rect 1733 1684 1736 1712
rect 1763 1684 1766 1708
rect 435 1680 497 1684
rect 501 1680 503 1684
rect 507 1680 511 1684
rect 515 1680 529 1684
rect 533 1680 538 1684
rect 542 1680 547 1684
rect 551 1680 570 1684
rect 574 1680 604 1684
rect 608 1680 619 1684
rect 623 1680 647 1684
rect 651 1680 664 1684
rect 668 1680 688 1684
rect 692 1680 742 1684
rect 746 1680 769 1684
rect 773 1680 793 1684
rect 797 1680 845 1684
rect 1368 1680 1430 1684
rect 1434 1680 1436 1684
rect 1440 1680 1444 1684
rect 1448 1680 1462 1684
rect 1466 1680 1471 1684
rect 1475 1680 1480 1684
rect 1484 1680 1503 1684
rect 1507 1680 1537 1684
rect 1541 1680 1552 1684
rect 1556 1680 1580 1684
rect 1584 1680 1597 1684
rect 1601 1680 1621 1684
rect 1625 1680 1675 1684
rect 1679 1680 1702 1684
rect 1706 1680 1726 1684
rect 1730 1680 1778 1684
rect 447 1673 511 1677
rect 515 1673 570 1677
rect 574 1673 595 1677
rect 599 1673 626 1677
rect 630 1673 659 1677
rect 558 1666 559 1670
rect 583 1665 584 1669
rect 630 1666 631 1670
rect 695 1661 698 1680
rect 800 1661 803 1680
rect 1380 1673 1444 1677
rect 1448 1673 1503 1677
rect 1507 1673 1528 1677
rect 1532 1673 1559 1677
rect 1563 1673 1592 1677
rect 1491 1666 1492 1670
rect 1516 1665 1517 1669
rect 1563 1666 1564 1670
rect 1628 1661 1631 1680
rect 1733 1661 1736 1680
rect 506 1652 509 1657
rect 513 1652 516 1657
rect 496 1649 498 1652
rect 506 1649 516 1652
rect 506 1643 509 1649
rect 513 1643 516 1649
rect 522 1651 525 1657
rect 538 1652 541 1657
rect 522 1647 524 1651
rect 528 1647 530 1651
rect 538 1650 544 1652
rect 548 1650 549 1652
rect 538 1648 549 1650
rect 566 1650 569 1657
rect 522 1643 525 1647
rect 538 1643 541 1648
rect 567 1646 569 1650
rect 566 1643 569 1646
rect 582 1651 585 1657
rect 592 1651 595 1657
rect 613 1652 616 1657
rect 592 1647 601 1651
rect 613 1648 614 1652
rect 618 1649 621 1652
rect 638 1651 641 1657
rect 656 1652 659 1657
rect 582 1643 585 1647
rect 592 1643 595 1647
rect 613 1643 616 1648
rect 640 1647 641 1651
rect 685 1648 690 1653
rect 694 1649 696 1652
rect 711 1651 714 1657
rect 711 1648 719 1651
rect 791 1648 796 1653
rect 800 1649 801 1652
rect 816 1651 819 1657
rect 816 1648 824 1651
rect 1439 1652 1442 1657
rect 1446 1652 1449 1657
rect 1429 1649 1431 1652
rect 1439 1649 1449 1652
rect 638 1643 641 1647
rect 656 1643 659 1648
rect 711 1645 714 1648
rect 816 1645 819 1648
rect 1439 1643 1442 1649
rect 566 1628 569 1632
rect 593 1628 594 1632
rect 638 1628 640 1632
rect 459 1621 523 1625
rect 527 1621 554 1625
rect 558 1621 576 1625
rect 580 1621 641 1625
rect 645 1621 659 1625
rect 695 1618 698 1637
rect 800 1618 803 1637
rect 1446 1643 1449 1649
rect 1455 1651 1458 1657
rect 1471 1652 1474 1657
rect 1455 1647 1457 1651
rect 1461 1647 1463 1651
rect 1471 1650 1477 1652
rect 1481 1650 1482 1652
rect 1471 1648 1482 1650
rect 1499 1650 1502 1657
rect 1455 1643 1458 1647
rect 1471 1643 1474 1648
rect 1500 1646 1502 1650
rect 1499 1643 1502 1646
rect 1515 1651 1518 1657
rect 1525 1651 1528 1657
rect 1546 1652 1549 1657
rect 1525 1647 1534 1651
rect 1546 1648 1547 1652
rect 1551 1649 1554 1652
rect 1571 1651 1574 1657
rect 1589 1652 1592 1657
rect 1515 1643 1518 1647
rect 1525 1643 1528 1647
rect 1546 1643 1549 1648
rect 1573 1647 1574 1651
rect 1618 1648 1623 1653
rect 1627 1649 1629 1652
rect 1644 1651 1647 1657
rect 1644 1648 1652 1651
rect 1724 1648 1729 1653
rect 1733 1649 1734 1652
rect 1749 1651 1752 1657
rect 1749 1648 1757 1651
rect 1571 1643 1574 1647
rect 1589 1643 1592 1648
rect 1644 1645 1647 1648
rect 1749 1645 1752 1648
rect 1499 1628 1502 1632
rect 1526 1628 1527 1632
rect 1571 1628 1573 1632
rect 1392 1621 1456 1625
rect 1460 1621 1487 1625
rect 1491 1621 1509 1625
rect 1513 1621 1574 1625
rect 1578 1621 1592 1625
rect 1628 1618 1631 1637
rect 1733 1618 1736 1637
rect 423 1614 496 1618
rect 500 1614 512 1618
rect 516 1614 530 1618
rect 534 1614 541 1618
rect 545 1614 547 1618
rect 551 1614 566 1618
rect 570 1614 603 1618
rect 607 1614 608 1618
rect 612 1614 620 1618
rect 624 1614 648 1618
rect 652 1614 664 1618
rect 668 1614 688 1618
rect 692 1614 742 1618
rect 746 1614 769 1618
rect 773 1614 823 1618
rect 827 1614 831 1618
rect 835 1614 859 1618
rect 863 1614 913 1618
rect 1356 1614 1429 1618
rect 1433 1614 1445 1618
rect 1449 1614 1463 1618
rect 1467 1614 1474 1618
rect 1478 1614 1480 1618
rect 1484 1614 1499 1618
rect 1503 1614 1536 1618
rect 1540 1614 1541 1618
rect 1545 1614 1553 1618
rect 1557 1614 1581 1618
rect 1585 1614 1597 1618
rect 1601 1614 1621 1618
rect 1625 1614 1675 1618
rect 1679 1614 1702 1618
rect 1706 1614 1756 1618
rect 1760 1614 1764 1618
rect 1768 1614 1792 1618
rect 1796 1614 1846 1618
rect 459 1607 523 1611
rect 527 1607 554 1611
rect 558 1607 576 1611
rect 580 1607 641 1611
rect 645 1607 659 1611
rect 695 1604 698 1614
rect 725 1610 728 1614
rect 752 1610 755 1614
rect 566 1600 569 1604
rect 593 1600 594 1604
rect 638 1600 640 1604
rect 495 1580 498 1583
rect 506 1583 509 1589
rect 513 1583 516 1589
rect 506 1580 516 1583
rect 506 1575 509 1580
rect 513 1575 516 1580
rect 522 1585 525 1589
rect 522 1581 524 1585
rect 528 1581 530 1585
rect 538 1584 541 1589
rect 566 1586 569 1589
rect 538 1582 549 1584
rect 522 1575 525 1581
rect 538 1580 544 1582
rect 538 1575 541 1580
rect 548 1580 549 1582
rect 567 1582 569 1586
rect 566 1575 569 1582
rect 711 1593 714 1596
rect 582 1585 585 1589
rect 592 1585 595 1589
rect 592 1581 601 1585
rect 613 1584 616 1589
rect 638 1585 641 1589
rect 582 1575 585 1581
rect 592 1575 595 1581
rect 613 1580 614 1584
rect 618 1580 621 1583
rect 640 1581 641 1585
rect 656 1584 659 1589
rect 688 1589 699 1592
rect 711 1590 719 1593
rect 613 1575 616 1580
rect 638 1575 641 1581
rect 688 1583 691 1589
rect 711 1584 714 1590
rect 723 1585 726 1588
rect 734 1588 737 1602
rect 761 1597 764 1602
rect 776 1604 779 1614
rect 806 1610 809 1614
rect 842 1610 845 1614
rect 745 1593 746 1596
rect 750 1593 753 1596
rect 792 1593 795 1596
rect 734 1585 742 1588
rect 761 1588 764 1593
rect 656 1575 659 1580
rect 734 1580 737 1585
rect 742 1581 746 1585
rect 769 1589 780 1592
rect 792 1590 800 1593
rect 686 1574 691 1579
rect 558 1562 559 1566
rect 583 1563 584 1567
rect 630 1562 631 1566
rect 447 1555 511 1559
rect 515 1555 570 1559
rect 574 1555 595 1559
rect 599 1555 626 1559
rect 630 1555 659 1559
rect 695 1552 698 1580
rect 725 1552 728 1576
rect 752 1552 755 1584
rect 769 1583 772 1589
rect 792 1584 795 1590
rect 804 1585 807 1588
rect 815 1588 818 1602
rect 851 1597 854 1602
rect 866 1604 869 1614
rect 896 1610 899 1614
rect 840 1593 843 1596
rect 1392 1607 1456 1611
rect 1460 1607 1487 1611
rect 1491 1607 1509 1611
rect 1513 1607 1574 1611
rect 1578 1607 1592 1611
rect 1628 1604 1631 1614
rect 1658 1610 1661 1614
rect 1685 1610 1688 1614
rect 882 1593 885 1596
rect 815 1585 824 1588
rect 851 1588 854 1593
rect 815 1580 818 1585
rect 767 1574 772 1579
rect 776 1552 779 1580
rect 858 1591 870 1592
rect 862 1589 870 1591
rect 882 1590 890 1593
rect 882 1584 885 1590
rect 894 1585 897 1588
rect 905 1588 908 1602
rect 1499 1600 1502 1604
rect 1526 1600 1527 1604
rect 1571 1600 1573 1604
rect 905 1585 925 1588
rect 806 1552 809 1576
rect 842 1552 845 1584
rect 905 1580 908 1585
rect 1428 1580 1431 1583
rect 1439 1583 1442 1589
rect 1446 1583 1449 1589
rect 1439 1580 1449 1583
rect 866 1552 869 1580
rect 896 1552 899 1576
rect 1439 1575 1442 1580
rect 1446 1575 1449 1580
rect 1455 1585 1458 1589
rect 1455 1581 1457 1585
rect 1461 1581 1463 1585
rect 1471 1584 1474 1589
rect 1499 1586 1502 1589
rect 1471 1582 1482 1584
rect 1455 1575 1458 1581
rect 1471 1580 1477 1582
rect 1471 1575 1474 1580
rect 1481 1580 1482 1582
rect 1500 1582 1502 1586
rect 1499 1575 1502 1582
rect 1644 1593 1647 1596
rect 1515 1585 1518 1589
rect 1525 1585 1528 1589
rect 1525 1581 1534 1585
rect 1546 1584 1549 1589
rect 1571 1585 1574 1589
rect 1515 1575 1518 1581
rect 1525 1575 1528 1581
rect 1546 1580 1547 1584
rect 1551 1580 1554 1583
rect 1573 1581 1574 1585
rect 1589 1584 1592 1589
rect 1621 1589 1632 1592
rect 1644 1590 1652 1593
rect 1546 1575 1549 1580
rect 1571 1575 1574 1581
rect 1621 1583 1624 1589
rect 1644 1584 1647 1590
rect 1656 1585 1659 1588
rect 1667 1588 1670 1602
rect 1694 1597 1697 1602
rect 1709 1604 1712 1614
rect 1739 1610 1742 1614
rect 1775 1610 1778 1614
rect 1678 1593 1679 1596
rect 1683 1593 1686 1596
rect 1725 1593 1728 1596
rect 1667 1585 1675 1588
rect 1694 1588 1697 1593
rect 1589 1575 1592 1580
rect 1667 1580 1670 1585
rect 1675 1581 1679 1585
rect 1702 1589 1713 1592
rect 1725 1590 1733 1593
rect 1619 1574 1624 1579
rect 1491 1562 1492 1566
rect 1516 1563 1517 1567
rect 1563 1562 1564 1566
rect 1380 1555 1444 1559
rect 1448 1555 1503 1559
rect 1507 1555 1528 1559
rect 1532 1555 1559 1559
rect 1563 1555 1592 1559
rect 1628 1552 1631 1580
rect 1658 1552 1661 1576
rect 1685 1552 1688 1584
rect 1702 1583 1705 1589
rect 1725 1584 1728 1590
rect 1737 1585 1740 1588
rect 1748 1588 1751 1602
rect 1784 1597 1787 1602
rect 1799 1604 1802 1614
rect 1829 1610 1832 1614
rect 1773 1593 1776 1596
rect 1815 1593 1818 1596
rect 1748 1585 1757 1588
rect 1784 1588 1787 1593
rect 1748 1580 1751 1585
rect 1700 1574 1705 1579
rect 1709 1552 1712 1580
rect 1791 1591 1803 1592
rect 1795 1589 1803 1591
rect 1815 1590 1823 1593
rect 1815 1584 1818 1590
rect 1827 1585 1830 1588
rect 1838 1588 1841 1602
rect 1838 1585 1858 1588
rect 1739 1552 1742 1576
rect 1775 1552 1778 1584
rect 1838 1580 1841 1585
rect 1799 1552 1802 1580
rect 1829 1552 1832 1576
rect 435 1548 497 1552
rect 501 1548 503 1552
rect 507 1548 511 1552
rect 515 1548 529 1552
rect 533 1548 538 1552
rect 542 1548 547 1552
rect 551 1548 570 1552
rect 574 1548 604 1552
rect 608 1548 619 1552
rect 623 1548 647 1552
rect 651 1548 664 1552
rect 668 1548 688 1552
rect 692 1548 742 1552
rect 749 1548 769 1552
rect 773 1548 823 1552
rect 827 1548 859 1552
rect 863 1548 913 1552
rect 1368 1548 1430 1552
rect 1434 1548 1436 1552
rect 1440 1548 1444 1552
rect 1448 1548 1462 1552
rect 1466 1548 1471 1552
rect 1475 1548 1480 1552
rect 1484 1548 1503 1552
rect 1507 1548 1537 1552
rect 1541 1548 1552 1552
rect 1556 1548 1580 1552
rect 1584 1548 1597 1552
rect 1601 1548 1621 1552
rect 1625 1548 1675 1552
rect 1682 1548 1702 1552
rect 1706 1548 1756 1552
rect 1760 1548 1792 1552
rect 1796 1548 1846 1552
rect 447 1541 511 1545
rect 515 1541 570 1545
rect 574 1541 595 1545
rect 599 1541 626 1545
rect 630 1541 659 1545
rect 558 1534 559 1538
rect 583 1533 584 1537
rect 630 1534 631 1538
rect 506 1520 509 1525
rect 513 1520 516 1525
rect 496 1517 498 1520
rect 506 1517 516 1520
rect 506 1511 509 1517
rect 513 1511 516 1517
rect 522 1519 525 1525
rect 538 1520 541 1525
rect 522 1515 524 1519
rect 528 1515 530 1519
rect 538 1518 544 1520
rect 548 1518 549 1520
rect 538 1516 549 1518
rect 566 1518 569 1525
rect 522 1511 525 1515
rect 538 1511 541 1516
rect 567 1514 569 1518
rect 566 1511 569 1514
rect 582 1519 585 1525
rect 592 1519 595 1525
rect 613 1520 616 1525
rect 592 1515 601 1519
rect 613 1516 614 1520
rect 618 1517 621 1520
rect 638 1519 641 1525
rect 656 1520 659 1525
rect 695 1526 698 1548
rect 776 1526 779 1548
rect 866 1526 869 1548
rect 1380 1541 1444 1545
rect 1448 1541 1503 1545
rect 1507 1541 1528 1545
rect 1532 1541 1559 1545
rect 1563 1541 1592 1545
rect 1491 1534 1492 1538
rect 1516 1533 1517 1537
rect 1563 1534 1564 1538
rect 582 1511 585 1515
rect 592 1511 595 1515
rect 613 1511 616 1516
rect 640 1515 641 1519
rect 638 1511 641 1515
rect 656 1511 659 1516
rect 686 1513 691 1518
rect 695 1514 696 1517
rect 711 1516 714 1522
rect 711 1513 719 1516
rect 766 1513 771 1518
rect 775 1514 777 1517
rect 792 1516 795 1522
rect 792 1513 800 1516
rect 859 1514 867 1517
rect 882 1516 885 1522
rect 1439 1520 1442 1525
rect 1446 1520 1449 1525
rect 1429 1517 1431 1520
rect 882 1513 890 1516
rect 1439 1517 1449 1520
rect 711 1510 714 1513
rect 792 1510 795 1513
rect 882 1510 885 1513
rect 1439 1511 1442 1517
rect 566 1496 569 1500
rect 593 1496 594 1500
rect 638 1496 640 1500
rect 1446 1511 1449 1517
rect 1455 1519 1458 1525
rect 1471 1520 1474 1525
rect 1455 1515 1457 1519
rect 1461 1515 1463 1519
rect 1471 1518 1477 1520
rect 1481 1518 1482 1520
rect 1471 1516 1482 1518
rect 1499 1518 1502 1525
rect 1455 1511 1458 1515
rect 1471 1511 1474 1516
rect 1500 1514 1502 1518
rect 1499 1511 1502 1514
rect 1515 1519 1518 1525
rect 1525 1519 1528 1525
rect 1546 1520 1549 1525
rect 1525 1515 1534 1519
rect 1546 1516 1547 1520
rect 1551 1517 1554 1520
rect 1571 1519 1574 1525
rect 1589 1520 1592 1525
rect 1628 1526 1631 1548
rect 1709 1526 1712 1548
rect 1799 1526 1802 1548
rect 1515 1511 1518 1515
rect 1525 1511 1528 1515
rect 1546 1511 1549 1516
rect 1573 1515 1574 1519
rect 1571 1511 1574 1515
rect 1589 1511 1592 1516
rect 1619 1513 1624 1518
rect 1628 1514 1629 1517
rect 1644 1516 1647 1522
rect 1644 1513 1652 1516
rect 1699 1513 1704 1518
rect 1708 1514 1710 1517
rect 1725 1516 1728 1522
rect 1725 1513 1733 1516
rect 1792 1514 1800 1517
rect 1815 1516 1818 1522
rect 1815 1513 1823 1516
rect 1644 1510 1647 1513
rect 1725 1510 1728 1513
rect 1815 1510 1818 1513
rect 459 1489 523 1493
rect 527 1489 554 1493
rect 558 1489 576 1493
rect 580 1489 641 1493
rect 645 1489 659 1493
rect 695 1486 698 1502
rect 776 1486 779 1502
rect 866 1486 869 1502
rect 1499 1496 1502 1500
rect 1526 1496 1527 1500
rect 1571 1496 1573 1500
rect 1392 1489 1456 1493
rect 1460 1489 1487 1493
rect 1491 1489 1509 1493
rect 1513 1489 1574 1493
rect 1578 1489 1592 1493
rect 1628 1486 1631 1502
rect 1709 1486 1712 1502
rect 1799 1486 1802 1502
rect 423 1482 496 1486
rect 500 1482 512 1486
rect 516 1482 530 1486
rect 534 1482 541 1486
rect 545 1482 547 1486
rect 551 1482 566 1486
rect 570 1482 603 1486
rect 607 1482 608 1486
rect 612 1482 620 1486
rect 624 1482 648 1486
rect 652 1482 664 1486
rect 668 1482 688 1486
rect 692 1482 742 1486
rect 746 1482 769 1486
rect 773 1482 859 1486
rect 863 1482 917 1486
rect 1356 1482 1429 1486
rect 1433 1482 1445 1486
rect 1449 1482 1463 1486
rect 1467 1482 1474 1486
rect 1478 1482 1480 1486
rect 1484 1482 1499 1486
rect 1503 1482 1536 1486
rect 1540 1482 1541 1486
rect 1545 1482 1553 1486
rect 1557 1482 1581 1486
rect 1585 1482 1597 1486
rect 1601 1482 1621 1486
rect 1625 1482 1675 1486
rect 1679 1482 1702 1486
rect 1706 1482 1792 1486
rect 1796 1482 1850 1486
rect 459 1475 523 1479
rect 527 1475 554 1479
rect 558 1475 576 1479
rect 580 1475 641 1479
rect 645 1475 659 1479
rect 695 1472 698 1482
rect 725 1478 728 1482
rect 566 1468 569 1472
rect 593 1468 594 1472
rect 638 1468 640 1472
rect 495 1448 498 1451
rect 506 1451 509 1457
rect 513 1451 516 1457
rect 506 1448 516 1451
rect 506 1443 509 1448
rect 513 1443 516 1448
rect 522 1453 525 1457
rect 522 1449 524 1453
rect 528 1449 530 1453
rect 538 1452 541 1457
rect 566 1454 569 1457
rect 538 1450 549 1452
rect 522 1443 525 1449
rect 538 1448 544 1450
rect 538 1443 541 1448
rect 548 1448 549 1450
rect 567 1450 569 1454
rect 566 1443 569 1450
rect 1392 1475 1456 1479
rect 1460 1475 1487 1479
rect 1491 1475 1509 1479
rect 1513 1475 1574 1479
rect 1578 1475 1592 1479
rect 1628 1472 1631 1482
rect 1658 1478 1661 1482
rect 711 1461 714 1464
rect 582 1453 585 1457
rect 592 1453 595 1457
rect 592 1449 601 1453
rect 613 1452 616 1457
rect 638 1453 641 1457
rect 582 1443 585 1449
rect 592 1443 595 1449
rect 613 1448 614 1452
rect 618 1448 621 1451
rect 640 1449 641 1453
rect 656 1452 659 1457
rect 688 1457 699 1460
rect 711 1458 719 1461
rect 613 1443 616 1448
rect 638 1443 641 1449
rect 688 1451 691 1457
rect 711 1452 714 1458
rect 723 1453 726 1456
rect 734 1456 737 1470
rect 1499 1468 1502 1472
rect 1526 1468 1527 1472
rect 1571 1468 1573 1472
rect 742 1456 747 1461
rect 734 1453 742 1456
rect 656 1443 659 1448
rect 734 1448 737 1453
rect 1428 1448 1431 1451
rect 1439 1451 1442 1457
rect 1446 1451 1449 1457
rect 1439 1448 1449 1451
rect 686 1442 691 1447
rect 17 1427 26 1431
rect 30 1427 62 1431
rect 66 1427 129 1431
rect 133 1427 158 1431
rect 162 1427 194 1431
rect 198 1427 261 1431
rect 265 1427 290 1431
rect 294 1427 326 1431
rect 330 1427 393 1431
rect 397 1427 477 1431
rect 558 1430 559 1434
rect 583 1431 584 1435
rect 630 1430 631 1434
rect 17 1420 50 1424
rect 54 1420 78 1424
rect 82 1420 108 1424
rect 112 1420 145 1424
rect 149 1420 182 1424
rect 186 1420 210 1424
rect 214 1420 240 1424
rect 244 1420 277 1424
rect 281 1420 314 1424
rect 318 1420 342 1424
rect 346 1420 372 1424
rect 376 1420 409 1424
rect 413 1420 417 1424
rect 490 1423 511 1427
rect 515 1423 520 1427
rect 524 1423 570 1427
rect 574 1423 595 1427
rect 599 1423 626 1427
rect 630 1423 659 1427
rect 695 1420 698 1448
rect 725 1420 728 1444
rect 1439 1443 1442 1448
rect 1446 1443 1449 1448
rect 1455 1453 1458 1457
rect 1455 1449 1457 1453
rect 1461 1449 1463 1453
rect 1471 1452 1474 1457
rect 1499 1454 1502 1457
rect 1471 1450 1482 1452
rect 1455 1443 1458 1449
rect 1471 1448 1477 1450
rect 1471 1443 1474 1448
rect 1481 1448 1482 1450
rect 1500 1450 1502 1454
rect 1499 1443 1502 1450
rect 1644 1461 1647 1464
rect 1515 1453 1518 1457
rect 1525 1453 1528 1457
rect 1525 1449 1534 1453
rect 1546 1452 1549 1457
rect 1571 1453 1574 1457
rect 1515 1443 1518 1449
rect 1525 1443 1528 1449
rect 1546 1448 1547 1452
rect 1551 1448 1554 1451
rect 1573 1449 1574 1453
rect 1589 1452 1592 1457
rect 1621 1457 1632 1460
rect 1644 1458 1652 1461
rect 1546 1443 1549 1448
rect 1571 1443 1574 1449
rect 1621 1451 1624 1457
rect 1644 1452 1647 1458
rect 1656 1453 1659 1456
rect 1667 1456 1670 1470
rect 1675 1456 1680 1461
rect 1667 1453 1675 1456
rect 1589 1443 1592 1448
rect 1667 1448 1670 1453
rect 1619 1442 1624 1447
rect 950 1427 959 1431
rect 963 1427 995 1431
rect 999 1427 1062 1431
rect 1066 1427 1091 1431
rect 1095 1427 1127 1431
rect 1131 1427 1194 1431
rect 1198 1427 1223 1431
rect 1227 1427 1259 1431
rect 1263 1427 1326 1431
rect 1330 1427 1410 1431
rect 1491 1430 1492 1434
rect 1516 1431 1517 1435
rect 1563 1430 1564 1434
rect 950 1420 983 1424
rect 987 1420 1011 1424
rect 1015 1420 1041 1424
rect 1045 1420 1078 1424
rect 1082 1420 1115 1424
rect 1119 1420 1143 1424
rect 1147 1420 1173 1424
rect 1177 1420 1210 1424
rect 1214 1420 1247 1424
rect 1251 1420 1275 1424
rect 1279 1420 1305 1424
rect 1309 1420 1342 1424
rect 1346 1420 1350 1424
rect 1423 1423 1444 1427
rect 1448 1423 1453 1427
rect 1457 1423 1503 1427
rect 1507 1423 1528 1427
rect 1532 1423 1559 1427
rect 1563 1423 1592 1427
rect 1628 1420 1631 1448
rect 1658 1420 1661 1444
rect 20 1410 23 1420
rect 41 1410 44 1420
rect 57 1410 60 1420
rect 71 1413 76 1417
rect 80 1413 87 1417
rect 99 1410 102 1420
rect 115 1410 118 1420
rect 136 1410 139 1420
rect 152 1410 155 1420
rect 173 1410 176 1420
rect 189 1410 192 1420
rect 203 1413 208 1417
rect 212 1413 219 1417
rect 231 1410 234 1420
rect 247 1410 250 1420
rect 268 1410 271 1420
rect 284 1410 287 1420
rect 305 1410 308 1420
rect 321 1410 324 1420
rect 335 1413 340 1417
rect 344 1413 351 1417
rect 363 1410 366 1420
rect 379 1410 382 1420
rect 400 1410 403 1420
rect 435 1416 497 1420
rect 501 1416 503 1420
rect 507 1416 511 1420
rect 515 1416 529 1420
rect 533 1416 538 1420
rect 542 1416 547 1420
rect 551 1416 570 1420
rect 574 1416 604 1420
rect 608 1416 619 1420
rect 623 1416 647 1420
rect 651 1416 664 1420
rect 668 1416 688 1420
rect 692 1416 772 1420
rect 776 1416 790 1420
rect 794 1416 799 1420
rect 803 1416 808 1420
rect 812 1416 831 1420
rect 835 1416 865 1420
rect 869 1416 880 1420
rect 884 1416 908 1420
rect 912 1416 921 1420
rect 37 1396 42 1399
rect 46 1396 70 1399
rect 95 1396 102 1399
rect 106 1396 128 1399
rect 148 1396 155 1399
rect 169 1396 174 1399
rect 178 1396 202 1399
rect 227 1396 234 1399
rect 238 1396 260 1399
rect 280 1396 287 1399
rect 301 1396 306 1399
rect 310 1396 334 1399
rect 447 1409 511 1413
rect 515 1409 520 1413
rect 524 1409 570 1413
rect 574 1409 595 1413
rect 599 1409 626 1413
rect 630 1409 659 1413
rect 359 1396 366 1399
rect 370 1396 392 1399
rect 558 1402 559 1406
rect 583 1401 584 1405
rect 630 1402 631 1406
rect 53 1386 60 1389
rect 64 1390 83 1393
rect 83 1383 86 1389
rect 111 1386 118 1389
rect 122 1390 137 1393
rect 185 1386 192 1389
rect 196 1390 215 1393
rect 215 1383 218 1389
rect 243 1386 250 1389
rect 254 1390 269 1393
rect 317 1386 324 1389
rect 328 1390 347 1393
rect 347 1383 350 1389
rect 375 1386 382 1389
rect 386 1390 403 1393
rect 506 1388 509 1393
rect 513 1388 516 1393
rect 496 1385 498 1388
rect 506 1385 516 1388
rect 506 1379 509 1385
rect 20 1367 23 1379
rect 41 1367 44 1379
rect 57 1367 60 1379
rect 71 1370 83 1373
rect 99 1367 102 1379
rect 115 1367 118 1379
rect 136 1367 139 1379
rect 152 1367 155 1379
rect 173 1367 176 1379
rect 189 1367 192 1379
rect 203 1370 215 1373
rect 231 1367 234 1379
rect 247 1367 250 1379
rect 268 1367 271 1379
rect 284 1367 287 1379
rect 305 1367 308 1379
rect 321 1367 324 1379
rect 335 1370 347 1373
rect 363 1367 366 1379
rect 379 1367 382 1379
rect 400 1367 403 1379
rect 513 1379 516 1385
rect 522 1387 525 1393
rect 538 1388 541 1393
rect 522 1383 524 1387
rect 528 1383 530 1387
rect 538 1386 544 1388
rect 548 1386 549 1388
rect 538 1384 549 1386
rect 566 1386 569 1393
rect 522 1379 525 1383
rect 538 1379 541 1384
rect 567 1382 569 1386
rect 566 1379 569 1382
rect 582 1387 585 1393
rect 592 1387 595 1393
rect 613 1388 616 1393
rect 592 1383 601 1387
rect 613 1384 614 1388
rect 618 1385 621 1388
rect 638 1387 641 1393
rect 656 1388 659 1393
rect 695 1390 698 1416
rect 731 1409 750 1413
rect 754 1409 772 1413
rect 776 1409 831 1413
rect 835 1409 856 1413
rect 860 1409 887 1413
rect 891 1409 920 1413
rect 953 1410 956 1420
rect 974 1410 977 1420
rect 990 1410 993 1420
rect 1004 1413 1009 1417
rect 1013 1413 1020 1417
rect 1032 1410 1035 1420
rect 1048 1410 1051 1420
rect 1069 1410 1072 1420
rect 1085 1410 1088 1420
rect 1106 1410 1109 1420
rect 1122 1410 1125 1420
rect 1136 1413 1141 1417
rect 1145 1413 1152 1417
rect 1164 1410 1167 1420
rect 1180 1410 1183 1420
rect 1201 1410 1204 1420
rect 1217 1410 1220 1420
rect 1238 1410 1241 1420
rect 1254 1410 1257 1420
rect 1268 1413 1273 1417
rect 1277 1413 1284 1417
rect 1296 1410 1299 1420
rect 1312 1410 1315 1420
rect 1333 1410 1336 1420
rect 1368 1416 1430 1420
rect 1434 1416 1436 1420
rect 1440 1416 1444 1420
rect 1448 1416 1462 1420
rect 1466 1416 1471 1420
rect 1475 1416 1480 1420
rect 1484 1416 1503 1420
rect 1507 1416 1537 1420
rect 1541 1416 1552 1420
rect 1556 1416 1580 1420
rect 1584 1416 1597 1420
rect 1601 1416 1621 1420
rect 1625 1416 1705 1420
rect 1709 1416 1723 1420
rect 1727 1416 1732 1420
rect 1736 1416 1741 1420
rect 1745 1416 1764 1420
rect 1768 1416 1798 1420
rect 1802 1416 1813 1420
rect 1817 1416 1841 1420
rect 1845 1416 1854 1420
rect 731 1397 734 1409
rect 819 1402 820 1406
rect 844 1401 845 1405
rect 891 1402 892 1406
rect 582 1379 585 1383
rect 592 1379 595 1383
rect 613 1379 616 1384
rect 640 1383 641 1387
rect 758 1388 761 1393
rect 767 1388 770 1393
rect 774 1388 777 1393
rect 638 1379 641 1383
rect 656 1379 659 1384
rect 685 1377 690 1382
rect 694 1378 696 1381
rect 711 1380 714 1386
rect 743 1385 777 1388
rect 711 1377 719 1380
rect 711 1374 714 1377
rect 17 1363 50 1367
rect 54 1363 78 1367
rect 82 1363 108 1367
rect 112 1363 182 1367
rect 186 1363 210 1367
rect 214 1363 240 1367
rect 244 1363 314 1367
rect 318 1363 342 1367
rect 346 1363 372 1367
rect 376 1363 429 1367
rect 566 1364 569 1368
rect 593 1364 594 1368
rect 638 1364 640 1368
rect 743 1371 746 1385
rect 767 1379 770 1385
rect 774 1379 777 1385
rect 783 1387 786 1393
rect 799 1388 802 1393
rect 783 1383 785 1387
rect 789 1383 791 1387
rect 799 1386 805 1388
rect 809 1386 810 1388
rect 799 1384 810 1386
rect 827 1386 830 1393
rect 783 1379 786 1383
rect 799 1379 802 1384
rect 828 1382 830 1386
rect 827 1379 830 1382
rect 970 1396 975 1399
rect 979 1396 1003 1399
rect 1028 1396 1035 1399
rect 1039 1396 1061 1399
rect 1081 1396 1088 1399
rect 1102 1396 1107 1399
rect 1111 1396 1135 1399
rect 1160 1396 1167 1399
rect 1171 1396 1193 1399
rect 1213 1396 1220 1399
rect 1234 1396 1239 1399
rect 1243 1396 1267 1399
rect 1380 1409 1444 1413
rect 1448 1409 1453 1413
rect 1457 1409 1503 1413
rect 1507 1409 1528 1413
rect 1532 1409 1559 1413
rect 1563 1409 1592 1413
rect 1292 1396 1299 1399
rect 1303 1396 1325 1399
rect 1491 1402 1492 1406
rect 1516 1401 1517 1405
rect 1563 1402 1564 1406
rect 843 1387 846 1393
rect 853 1387 856 1393
rect 874 1388 877 1393
rect 853 1383 862 1387
rect 874 1384 875 1388
rect 879 1385 882 1388
rect 899 1387 902 1393
rect 917 1388 920 1393
rect 843 1379 846 1383
rect 853 1379 856 1383
rect 874 1379 877 1384
rect 901 1383 902 1387
rect 899 1379 902 1383
rect 917 1379 920 1384
rect 986 1386 993 1389
rect 997 1390 1016 1393
rect 1016 1383 1019 1389
rect 1044 1386 1051 1389
rect 1055 1390 1070 1393
rect 1118 1386 1125 1389
rect 1129 1390 1148 1393
rect 1148 1383 1151 1389
rect 1176 1386 1183 1389
rect 1187 1390 1202 1393
rect 1250 1386 1257 1389
rect 1261 1390 1280 1393
rect 1280 1383 1283 1389
rect 1308 1386 1315 1389
rect 1319 1390 1336 1393
rect 1439 1388 1442 1393
rect 1446 1388 1449 1393
rect 1429 1385 1431 1388
rect 1439 1385 1449 1388
rect 1439 1379 1442 1385
rect 17 1356 26 1360
rect 30 1356 77 1360
rect 81 1356 127 1360
rect 131 1356 158 1360
rect 162 1356 209 1360
rect 213 1356 259 1360
rect 263 1356 290 1360
rect 294 1356 341 1360
rect 345 1356 391 1360
rect 395 1357 465 1360
rect 509 1357 523 1361
rect 527 1357 554 1361
rect 558 1357 576 1361
rect 580 1357 641 1361
rect 645 1357 659 1361
rect 695 1354 698 1366
rect 827 1364 830 1368
rect 854 1364 855 1368
rect 899 1364 901 1368
rect 953 1367 956 1379
rect 974 1367 977 1379
rect 990 1367 993 1379
rect 1004 1370 1016 1373
rect 1032 1367 1035 1379
rect 1048 1367 1051 1379
rect 1069 1367 1072 1379
rect 1085 1367 1088 1379
rect 1106 1367 1109 1379
rect 1122 1367 1125 1379
rect 1136 1370 1148 1373
rect 1164 1367 1167 1379
rect 1180 1367 1183 1379
rect 1201 1367 1204 1379
rect 1217 1367 1220 1379
rect 1238 1367 1241 1379
rect 1254 1367 1257 1379
rect 1268 1370 1280 1373
rect 1296 1367 1299 1379
rect 1312 1367 1315 1379
rect 1333 1367 1336 1379
rect 1446 1379 1449 1385
rect 1455 1387 1458 1393
rect 1471 1388 1474 1393
rect 1455 1383 1457 1387
rect 1461 1383 1463 1387
rect 1471 1386 1477 1388
rect 1481 1386 1482 1388
rect 1471 1384 1482 1386
rect 1499 1386 1502 1393
rect 1455 1379 1458 1383
rect 1471 1379 1474 1384
rect 1500 1382 1502 1386
rect 1499 1379 1502 1382
rect 1515 1387 1518 1393
rect 1525 1387 1528 1393
rect 1546 1388 1549 1393
rect 1525 1383 1534 1387
rect 1546 1384 1547 1388
rect 1551 1385 1554 1388
rect 1571 1387 1574 1393
rect 1589 1388 1592 1393
rect 1628 1390 1631 1416
rect 1664 1409 1683 1413
rect 1687 1409 1705 1413
rect 1709 1409 1764 1413
rect 1768 1409 1789 1413
rect 1793 1409 1820 1413
rect 1824 1409 1853 1413
rect 1664 1397 1667 1409
rect 1752 1402 1753 1406
rect 1777 1401 1778 1405
rect 1824 1402 1825 1406
rect 1515 1379 1518 1383
rect 1525 1379 1528 1383
rect 1546 1379 1549 1384
rect 1573 1383 1574 1387
rect 1691 1388 1694 1393
rect 1700 1388 1703 1393
rect 1707 1388 1710 1393
rect 1571 1379 1574 1383
rect 1589 1379 1592 1384
rect 1618 1377 1623 1382
rect 1627 1378 1629 1381
rect 1644 1380 1647 1386
rect 1676 1385 1710 1388
rect 1644 1377 1652 1380
rect 1644 1374 1647 1377
rect 950 1363 983 1367
rect 987 1363 1011 1367
rect 1015 1363 1041 1367
rect 1045 1363 1115 1367
rect 1119 1363 1143 1367
rect 1147 1363 1173 1367
rect 1177 1363 1247 1367
rect 1251 1363 1275 1367
rect 1279 1363 1305 1367
rect 1309 1363 1362 1367
rect 1499 1364 1502 1368
rect 1526 1364 1527 1368
rect 1571 1364 1573 1368
rect 1676 1371 1679 1385
rect 1700 1379 1703 1385
rect 1707 1379 1710 1385
rect 1716 1387 1719 1393
rect 1732 1388 1735 1393
rect 1716 1383 1718 1387
rect 1722 1383 1724 1387
rect 1732 1386 1738 1388
rect 1742 1386 1743 1388
rect 1732 1384 1743 1386
rect 1760 1386 1763 1393
rect 1716 1379 1719 1383
rect 1732 1379 1735 1384
rect 1761 1382 1763 1386
rect 1760 1379 1763 1382
rect 1776 1387 1779 1393
rect 1786 1387 1789 1393
rect 1807 1388 1810 1393
rect 1786 1383 1795 1387
rect 1807 1384 1808 1388
rect 1812 1385 1815 1388
rect 1832 1387 1835 1393
rect 1850 1388 1853 1393
rect 1776 1379 1779 1383
rect 1786 1379 1789 1383
rect 1807 1379 1810 1384
rect 1834 1383 1835 1387
rect 1832 1379 1835 1383
rect 1850 1379 1853 1384
rect 735 1357 740 1361
rect 744 1357 784 1361
rect 788 1357 815 1361
rect 819 1357 837 1361
rect 841 1357 902 1361
rect 906 1357 920 1361
rect 950 1356 959 1360
rect 963 1356 1010 1360
rect 1014 1356 1060 1360
rect 1064 1356 1091 1360
rect 1095 1356 1142 1360
rect 1146 1356 1192 1360
rect 1196 1356 1223 1360
rect 1227 1356 1274 1360
rect 1278 1356 1324 1360
rect 1328 1357 1398 1360
rect 1442 1357 1456 1361
rect 1460 1357 1487 1361
rect 1491 1357 1509 1361
rect 1513 1357 1574 1361
rect 1578 1357 1592 1361
rect 1628 1354 1631 1366
rect 1760 1364 1763 1368
rect 1787 1364 1788 1368
rect 1832 1364 1834 1368
rect 1668 1357 1673 1361
rect 1677 1357 1717 1361
rect 1721 1357 1748 1361
rect 1752 1357 1770 1361
rect 1774 1357 1835 1361
rect 1839 1357 1853 1361
rect 24 1350 408 1353
rect 423 1350 496 1354
rect 500 1350 512 1354
rect 516 1350 530 1354
rect 534 1350 541 1354
rect 545 1350 547 1354
rect 551 1350 566 1354
rect 570 1350 603 1354
rect 607 1350 608 1354
rect 612 1350 620 1354
rect 624 1350 648 1354
rect 652 1350 688 1354
rect 692 1350 731 1354
rect 735 1350 742 1354
rect 746 1350 757 1354
rect 761 1350 773 1354
rect 777 1350 791 1354
rect 795 1350 802 1354
rect 806 1350 808 1354
rect 812 1350 827 1354
rect 831 1350 864 1354
rect 868 1350 869 1354
rect 873 1350 881 1354
rect 885 1350 909 1354
rect 913 1350 921 1354
rect 957 1350 1341 1353
rect 1356 1350 1429 1354
rect 1433 1350 1445 1354
rect 1449 1350 1463 1354
rect 1467 1350 1474 1354
rect 1478 1350 1480 1354
rect 1484 1350 1499 1354
rect 1503 1350 1536 1354
rect 1540 1350 1541 1354
rect 1545 1350 1553 1354
rect 1557 1350 1581 1354
rect 1585 1350 1621 1354
rect 1625 1350 1664 1354
rect 1668 1350 1675 1354
rect 1679 1350 1690 1354
rect 1694 1350 1706 1354
rect 1710 1350 1724 1354
rect 1728 1350 1735 1354
rect 1739 1350 1741 1354
rect 1745 1350 1760 1354
rect 1764 1350 1797 1354
rect 1801 1350 1802 1354
rect 1806 1350 1814 1354
rect 1818 1350 1842 1354
rect 1846 1350 1854 1354
rect 167 1343 276 1346
rect 459 1343 505 1347
rect 509 1343 739 1346
rect 929 1344 937 1348
rect 1100 1343 1209 1346
rect 1392 1343 1438 1347
rect 1442 1343 1672 1346
rect 1862 1344 1870 1348
rect 147 1335 151 1339
rect 155 1335 159 1339
rect 447 1336 749 1339
rect 925 1328 929 1332
rect 1080 1335 1084 1339
rect 1088 1335 1092 1339
rect 1380 1336 1682 1339
rect 1858 1328 1862 1332
rect 7 1324 135 1328
rect 139 1324 155 1328
rect 171 1324 1068 1328
rect 1072 1324 1088 1328
rect 1104 1324 1950 1328
rect 163 1317 408 1320
rect 483 1317 797 1321
rect 801 1317 833 1321
rect 837 1317 900 1321
rect 904 1317 920 1321
rect 1096 1317 1341 1320
rect 1416 1317 1730 1321
rect 1734 1317 1766 1321
rect 1770 1317 1833 1321
rect 1837 1317 1853 1321
rect 178 1310 408 1313
rect 423 1310 783 1314
rect 787 1310 821 1314
rect 825 1310 849 1314
rect 853 1310 879 1314
rect 883 1310 916 1314
rect 147 1301 151 1305
rect 155 1301 159 1305
rect 791 1300 794 1310
rect 812 1300 815 1310
rect 828 1300 831 1310
rect 842 1303 847 1307
rect 851 1303 858 1307
rect 870 1300 873 1310
rect 886 1300 889 1310
rect 907 1300 910 1310
rect 1111 1310 1341 1313
rect 1356 1310 1716 1314
rect 1720 1310 1754 1314
rect 1758 1310 1782 1314
rect 1786 1310 1812 1314
rect 1816 1310 1849 1314
rect 1080 1301 1084 1305
rect 1088 1301 1092 1305
rect 1724 1300 1727 1310
rect 1745 1300 1748 1310
rect 1761 1300 1764 1310
rect 1775 1303 1780 1307
rect 1784 1303 1791 1307
rect 1803 1300 1806 1310
rect 1819 1300 1822 1310
rect 1840 1300 1843 1310
rect 167 1294 277 1297
rect 17 1287 26 1291
rect 30 1287 62 1291
rect 66 1287 129 1291
rect 133 1287 158 1291
rect 162 1287 194 1291
rect 198 1287 261 1291
rect 265 1287 290 1291
rect 294 1287 326 1291
rect 330 1287 393 1291
rect 397 1287 477 1291
rect 17 1280 50 1284
rect 54 1280 78 1284
rect 82 1280 108 1284
rect 112 1280 145 1284
rect 149 1280 182 1284
rect 186 1280 210 1284
rect 214 1280 240 1284
rect 244 1280 277 1284
rect 281 1280 314 1284
rect 318 1280 342 1284
rect 346 1280 372 1284
rect 376 1280 409 1284
rect 413 1280 417 1284
rect 808 1286 813 1289
rect 817 1286 841 1289
rect 1100 1294 1210 1297
rect 866 1286 873 1289
rect 877 1286 899 1289
rect 950 1287 959 1291
rect 963 1287 995 1291
rect 999 1287 1062 1291
rect 1066 1287 1091 1291
rect 1095 1287 1127 1291
rect 1131 1287 1194 1291
rect 1198 1287 1223 1291
rect 1227 1287 1259 1291
rect 1263 1287 1326 1291
rect 1330 1287 1410 1291
rect 20 1270 23 1280
rect 41 1270 44 1280
rect 57 1270 60 1280
rect 71 1273 76 1277
rect 80 1273 87 1277
rect 99 1270 102 1280
rect 115 1270 118 1280
rect 136 1270 139 1280
rect 152 1270 155 1280
rect 173 1270 176 1280
rect 189 1270 192 1280
rect 203 1273 208 1277
rect 212 1273 219 1277
rect 231 1270 234 1280
rect 247 1270 250 1280
rect 268 1270 271 1280
rect 284 1270 287 1280
rect 305 1270 308 1280
rect 321 1270 324 1280
rect 335 1273 340 1277
rect 344 1273 351 1277
rect 363 1270 366 1280
rect 379 1270 382 1280
rect 400 1270 403 1280
rect 824 1276 831 1279
rect 835 1280 854 1283
rect 37 1256 42 1259
rect 46 1256 70 1259
rect 95 1256 102 1259
rect 106 1256 128 1259
rect 148 1256 155 1259
rect 169 1256 174 1259
rect 178 1256 202 1259
rect 227 1256 234 1259
rect 238 1256 260 1259
rect 280 1256 287 1259
rect 301 1256 306 1259
rect 310 1256 334 1259
rect 359 1256 366 1259
rect 370 1256 392 1259
rect 854 1273 857 1279
rect 882 1276 889 1279
rect 893 1280 908 1283
rect 950 1280 983 1284
rect 987 1280 1011 1284
rect 1015 1280 1041 1284
rect 1045 1280 1078 1284
rect 1082 1280 1115 1284
rect 1119 1280 1143 1284
rect 1147 1280 1173 1284
rect 1177 1280 1210 1284
rect 1214 1280 1247 1284
rect 1251 1280 1275 1284
rect 1279 1280 1305 1284
rect 1309 1280 1342 1284
rect 1346 1280 1350 1284
rect 1741 1286 1746 1289
rect 1750 1286 1774 1289
rect 1799 1286 1806 1289
rect 1810 1286 1832 1289
rect 953 1270 956 1280
rect 974 1270 977 1280
rect 990 1270 993 1280
rect 1004 1273 1009 1277
rect 1013 1273 1020 1277
rect 1032 1270 1035 1280
rect 1048 1270 1051 1280
rect 1069 1270 1072 1280
rect 1085 1270 1088 1280
rect 1106 1270 1109 1280
rect 1122 1270 1125 1280
rect 1136 1273 1141 1277
rect 1145 1273 1152 1277
rect 1164 1270 1167 1280
rect 1180 1270 1183 1280
rect 1201 1270 1204 1280
rect 1217 1270 1220 1280
rect 1238 1270 1241 1280
rect 1254 1270 1257 1280
rect 1268 1273 1273 1277
rect 1277 1273 1284 1277
rect 1296 1270 1299 1280
rect 1312 1270 1315 1280
rect 1333 1270 1336 1280
rect 1757 1276 1764 1279
rect 1768 1280 1787 1283
rect 791 1257 794 1269
rect 812 1257 815 1269
rect 828 1257 831 1269
rect 842 1260 854 1263
rect 870 1257 873 1269
rect 886 1257 889 1269
rect 907 1257 910 1269
rect 53 1246 60 1249
rect 64 1250 83 1253
rect 83 1243 86 1249
rect 111 1246 118 1249
rect 122 1250 137 1253
rect 185 1246 192 1249
rect 196 1250 215 1253
rect 215 1243 218 1249
rect 243 1246 250 1249
rect 254 1250 269 1253
rect 317 1246 324 1249
rect 328 1250 347 1253
rect 347 1243 350 1249
rect 375 1246 382 1249
rect 386 1250 403 1253
rect 435 1253 821 1257
rect 825 1253 849 1257
rect 853 1253 879 1257
rect 883 1253 920 1257
rect 970 1256 975 1259
rect 979 1256 1003 1259
rect 1028 1256 1035 1259
rect 1039 1256 1061 1259
rect 1081 1256 1088 1259
rect 1102 1256 1107 1259
rect 1111 1256 1135 1259
rect 1160 1256 1167 1259
rect 1171 1256 1193 1259
rect 1213 1256 1220 1259
rect 1234 1256 1239 1259
rect 1243 1256 1267 1259
rect 1292 1256 1299 1259
rect 1303 1256 1325 1259
rect 1787 1273 1790 1279
rect 1815 1276 1822 1279
rect 1826 1280 1841 1283
rect 1724 1257 1727 1269
rect 1745 1257 1748 1269
rect 1761 1257 1764 1269
rect 1775 1260 1787 1263
rect 1803 1257 1806 1269
rect 1819 1257 1822 1269
rect 1840 1257 1843 1269
rect 471 1246 797 1250
rect 801 1246 848 1250
rect 852 1246 898 1250
rect 902 1246 920 1250
rect 986 1246 993 1249
rect 997 1250 1016 1253
rect 20 1227 23 1239
rect 41 1227 44 1239
rect 57 1227 60 1239
rect 71 1230 83 1233
rect 99 1227 102 1239
rect 115 1227 118 1239
rect 136 1227 139 1239
rect 152 1227 155 1239
rect 173 1227 176 1239
rect 189 1227 192 1239
rect 203 1230 215 1233
rect 231 1227 234 1239
rect 247 1227 250 1239
rect 268 1227 271 1239
rect 284 1227 287 1239
rect 305 1227 308 1239
rect 321 1227 324 1239
rect 335 1230 347 1233
rect 363 1227 366 1239
rect 379 1227 382 1239
rect 400 1227 403 1239
rect 794 1239 915 1242
rect 1016 1243 1019 1249
rect 1044 1246 1051 1249
rect 1055 1250 1070 1253
rect 1118 1246 1125 1249
rect 1129 1250 1148 1253
rect 1148 1243 1151 1249
rect 1176 1246 1183 1249
rect 1187 1250 1202 1253
rect 1250 1246 1257 1249
rect 1261 1250 1280 1253
rect 1280 1243 1283 1249
rect 1308 1246 1315 1249
rect 1319 1250 1336 1253
rect 1368 1253 1754 1257
rect 1758 1253 1782 1257
rect 1786 1253 1812 1257
rect 1816 1253 1853 1257
rect 1404 1246 1730 1250
rect 1734 1246 1781 1250
rect 1785 1246 1831 1250
rect 1835 1246 1853 1250
rect 483 1231 797 1235
rect 801 1231 833 1235
rect 837 1231 900 1235
rect 904 1231 920 1235
rect 17 1223 50 1227
rect 54 1223 78 1227
rect 82 1223 108 1227
rect 112 1223 182 1227
rect 186 1223 210 1227
rect 214 1223 240 1227
rect 244 1223 314 1227
rect 318 1223 342 1227
rect 346 1223 372 1227
rect 376 1223 429 1227
rect 787 1224 821 1228
rect 825 1224 849 1228
rect 853 1224 879 1228
rect 883 1224 916 1228
rect 953 1227 956 1239
rect 974 1227 977 1239
rect 990 1227 993 1239
rect 1004 1230 1016 1233
rect 1032 1227 1035 1239
rect 1048 1227 1051 1239
rect 1069 1227 1072 1239
rect 1085 1227 1088 1239
rect 1106 1227 1109 1239
rect 1122 1227 1125 1239
rect 1136 1230 1148 1233
rect 1164 1227 1167 1239
rect 1180 1227 1183 1239
rect 1201 1227 1204 1239
rect 1217 1227 1220 1239
rect 1238 1227 1241 1239
rect 1254 1227 1257 1239
rect 1268 1230 1280 1233
rect 1296 1227 1299 1239
rect 1312 1227 1315 1239
rect 1333 1227 1336 1239
rect 1727 1239 1848 1242
rect 1416 1231 1730 1235
rect 1734 1231 1766 1235
rect 1770 1231 1833 1235
rect 1837 1231 1853 1235
rect 17 1216 26 1220
rect 30 1216 77 1220
rect 81 1216 127 1220
rect 131 1216 158 1220
rect 162 1216 209 1220
rect 213 1216 259 1220
rect 263 1216 290 1220
rect 294 1216 341 1220
rect 345 1216 391 1220
rect 395 1216 465 1220
rect 791 1214 794 1224
rect 812 1214 815 1224
rect 828 1214 831 1224
rect 842 1217 847 1221
rect 851 1217 858 1221
rect 870 1214 873 1224
rect 886 1214 889 1224
rect 907 1214 910 1224
rect 950 1223 983 1227
rect 987 1223 1011 1227
rect 1015 1223 1041 1227
rect 1045 1223 1115 1227
rect 1119 1223 1143 1227
rect 1147 1223 1173 1227
rect 1177 1223 1247 1227
rect 1251 1223 1275 1227
rect 1279 1223 1305 1227
rect 1309 1223 1362 1227
rect 1720 1224 1754 1228
rect 1758 1224 1782 1228
rect 1786 1224 1812 1228
rect 1816 1224 1849 1228
rect 950 1216 959 1220
rect 963 1216 1010 1220
rect 1014 1216 1060 1220
rect 1064 1216 1091 1220
rect 1095 1216 1142 1220
rect 1146 1216 1192 1220
rect 1196 1216 1223 1220
rect 1227 1216 1274 1220
rect 1278 1216 1324 1220
rect 1328 1216 1398 1220
rect 1724 1214 1727 1224
rect 1745 1214 1748 1224
rect 1761 1214 1764 1224
rect 1775 1217 1780 1221
rect 1784 1217 1791 1221
rect 1803 1214 1806 1224
rect 1819 1214 1822 1224
rect 1840 1214 1843 1224
rect 23 1209 408 1212
rect 17 1201 26 1205
rect 30 1201 62 1205
rect 66 1201 129 1205
rect 133 1201 158 1205
rect 162 1201 194 1205
rect 198 1201 261 1205
rect 265 1201 290 1205
rect 294 1201 326 1205
rect 330 1201 393 1205
rect 397 1201 477 1205
rect 17 1194 50 1198
rect 54 1194 78 1198
rect 82 1194 108 1198
rect 112 1194 145 1198
rect 149 1194 182 1198
rect 186 1194 210 1198
rect 214 1194 240 1198
rect 244 1194 277 1198
rect 281 1194 314 1198
rect 318 1194 342 1198
rect 346 1194 372 1198
rect 376 1194 409 1198
rect 413 1194 417 1198
rect 808 1200 813 1203
rect 817 1200 841 1203
rect 956 1209 1341 1212
rect 866 1200 873 1203
rect 877 1200 899 1203
rect 950 1201 959 1205
rect 963 1201 995 1205
rect 999 1201 1062 1205
rect 1066 1201 1091 1205
rect 1095 1201 1127 1205
rect 1131 1201 1194 1205
rect 1198 1201 1223 1205
rect 1227 1201 1259 1205
rect 1263 1201 1326 1205
rect 1330 1201 1410 1205
rect 20 1184 23 1194
rect 41 1184 44 1194
rect 57 1184 60 1194
rect 71 1187 76 1191
rect 80 1187 87 1191
rect 99 1184 102 1194
rect 115 1184 118 1194
rect 136 1184 139 1194
rect 152 1184 155 1194
rect 173 1184 176 1194
rect 189 1184 192 1194
rect 203 1187 208 1191
rect 212 1187 219 1191
rect 231 1184 234 1194
rect 247 1184 250 1194
rect 268 1184 271 1194
rect 284 1184 287 1194
rect 305 1184 308 1194
rect 321 1184 324 1194
rect 335 1187 340 1191
rect 344 1187 351 1191
rect 363 1184 366 1194
rect 379 1184 382 1194
rect 400 1184 403 1194
rect 824 1190 831 1193
rect 835 1194 854 1197
rect 37 1170 42 1173
rect 46 1170 70 1173
rect 95 1170 102 1173
rect 106 1170 128 1173
rect 148 1170 155 1173
rect 169 1170 174 1173
rect 178 1170 202 1173
rect 227 1170 234 1173
rect 238 1170 260 1173
rect 280 1170 287 1173
rect 301 1170 306 1173
rect 310 1170 334 1173
rect 359 1170 366 1173
rect 370 1170 392 1173
rect 854 1187 857 1193
rect 882 1190 889 1193
rect 893 1194 908 1197
rect 919 1192 930 1196
rect 950 1194 983 1198
rect 987 1194 1011 1198
rect 1015 1194 1041 1198
rect 1045 1194 1078 1198
rect 1082 1194 1115 1198
rect 1119 1194 1143 1198
rect 1147 1194 1173 1198
rect 1177 1194 1210 1198
rect 1214 1194 1247 1198
rect 1251 1194 1275 1198
rect 1279 1194 1305 1198
rect 1309 1194 1342 1198
rect 1346 1194 1350 1198
rect 1741 1200 1746 1203
rect 1750 1200 1774 1203
rect 1799 1200 1806 1203
rect 1810 1200 1832 1203
rect 953 1184 956 1194
rect 974 1184 977 1194
rect 990 1184 993 1194
rect 1004 1187 1009 1191
rect 1013 1187 1020 1191
rect 1032 1184 1035 1194
rect 1048 1184 1051 1194
rect 1069 1184 1072 1194
rect 1085 1184 1088 1194
rect 1106 1184 1109 1194
rect 1122 1184 1125 1194
rect 1136 1187 1141 1191
rect 1145 1187 1152 1191
rect 1164 1184 1167 1194
rect 1180 1184 1183 1194
rect 1201 1184 1204 1194
rect 1217 1184 1220 1194
rect 1238 1184 1241 1194
rect 1254 1184 1257 1194
rect 1268 1187 1273 1191
rect 1277 1187 1284 1191
rect 1296 1184 1299 1194
rect 1312 1184 1315 1194
rect 1333 1184 1336 1194
rect 1757 1190 1764 1193
rect 1768 1194 1787 1197
rect 791 1171 794 1183
rect 812 1171 815 1183
rect 828 1171 831 1183
rect 842 1174 854 1177
rect 870 1171 873 1183
rect 886 1171 889 1183
rect 907 1171 910 1183
rect 53 1160 60 1163
rect 64 1164 83 1167
rect 83 1157 86 1163
rect 111 1160 118 1163
rect 122 1164 137 1167
rect 185 1160 192 1163
rect 196 1164 215 1167
rect 215 1157 218 1163
rect 243 1160 250 1163
rect 254 1164 269 1167
rect 317 1160 324 1163
rect 328 1164 347 1167
rect 347 1157 350 1163
rect 375 1160 382 1163
rect 386 1164 403 1167
rect 435 1167 821 1171
rect 825 1167 849 1171
rect 853 1167 879 1171
rect 883 1167 920 1171
rect 970 1170 975 1173
rect 979 1170 1003 1173
rect 1028 1170 1035 1173
rect 1039 1170 1061 1173
rect 1081 1170 1088 1173
rect 1102 1170 1107 1173
rect 1111 1170 1135 1173
rect 1160 1170 1167 1173
rect 1171 1170 1193 1173
rect 1213 1170 1220 1173
rect 1234 1170 1239 1173
rect 1243 1170 1267 1173
rect 1292 1170 1299 1173
rect 1303 1170 1325 1173
rect 1787 1187 1790 1193
rect 1815 1190 1822 1193
rect 1826 1194 1841 1197
rect 1852 1192 1863 1196
rect 1724 1171 1727 1183
rect 1745 1171 1748 1183
rect 1761 1171 1764 1183
rect 1775 1174 1787 1177
rect 1803 1171 1806 1183
rect 1819 1171 1822 1183
rect 1840 1171 1843 1183
rect 471 1160 797 1164
rect 801 1160 848 1164
rect 852 1160 898 1164
rect 902 1160 920 1164
rect 986 1160 993 1163
rect 997 1164 1016 1167
rect 1016 1157 1019 1163
rect 1044 1160 1051 1163
rect 1055 1164 1070 1167
rect 1118 1160 1125 1163
rect 1129 1164 1148 1167
rect 1148 1157 1151 1163
rect 1176 1160 1183 1163
rect 1187 1164 1202 1167
rect 1250 1160 1257 1163
rect 1261 1164 1280 1167
rect 1280 1157 1283 1163
rect 1308 1160 1315 1163
rect 1319 1164 1336 1167
rect 1368 1167 1754 1171
rect 1758 1167 1782 1171
rect 1786 1167 1812 1171
rect 1816 1167 1853 1171
rect 1404 1160 1730 1164
rect 1734 1160 1781 1164
rect 1785 1160 1831 1164
rect 1835 1160 1853 1164
rect 20 1141 23 1153
rect 41 1141 44 1153
rect 57 1141 60 1153
rect 71 1144 83 1147
rect 99 1141 102 1153
rect 115 1141 118 1153
rect 136 1141 139 1153
rect 152 1141 155 1153
rect 173 1141 176 1153
rect 189 1141 192 1153
rect 203 1144 215 1147
rect 231 1141 234 1153
rect 247 1141 250 1153
rect 268 1141 271 1153
rect 284 1141 287 1153
rect 305 1141 308 1153
rect 321 1141 324 1153
rect 335 1144 347 1147
rect 363 1141 366 1153
rect 379 1141 382 1153
rect 400 1141 403 1153
rect 953 1141 956 1153
rect 974 1141 977 1153
rect 990 1141 993 1153
rect 1004 1144 1016 1147
rect 1032 1141 1035 1153
rect 1048 1141 1051 1153
rect 1069 1141 1072 1153
rect 1085 1141 1088 1153
rect 1106 1141 1109 1153
rect 1122 1141 1125 1153
rect 1136 1144 1148 1147
rect 1164 1141 1167 1153
rect 1180 1141 1183 1153
rect 1201 1141 1204 1153
rect 1217 1141 1220 1153
rect 1238 1141 1241 1153
rect 1254 1141 1257 1153
rect 1268 1144 1280 1147
rect 1296 1141 1299 1153
rect 1312 1141 1315 1153
rect 1333 1141 1336 1153
rect 17 1137 50 1141
rect 54 1137 78 1141
rect 82 1137 108 1141
rect 112 1137 182 1141
rect 186 1137 210 1141
rect 214 1137 240 1141
rect 244 1137 314 1141
rect 318 1137 342 1141
rect 346 1137 372 1141
rect 376 1137 429 1141
rect 950 1137 983 1141
rect 987 1137 1011 1141
rect 1015 1137 1041 1141
rect 1045 1137 1115 1141
rect 1119 1137 1143 1141
rect 1147 1137 1173 1141
rect 1177 1137 1247 1141
rect 1251 1137 1275 1141
rect 1279 1137 1305 1141
rect 1309 1137 1362 1141
rect 17 1130 26 1134
rect 30 1130 77 1134
rect 81 1130 127 1134
rect 131 1130 158 1134
rect 162 1130 209 1134
rect 213 1130 259 1134
rect 263 1130 290 1134
rect 294 1130 341 1134
rect 345 1130 391 1134
rect 395 1130 465 1134
rect 950 1130 959 1134
rect 963 1130 1010 1134
rect 1014 1130 1060 1134
rect 1064 1130 1091 1134
rect 1095 1130 1142 1134
rect 1146 1130 1192 1134
rect 1196 1130 1223 1134
rect 1227 1130 1274 1134
rect 1278 1130 1324 1134
rect 1328 1130 1398 1134
rect 23 1124 408 1127
rect 956 1124 1341 1127
rect 148 1117 252 1120
rect 1081 1117 1185 1120
rect 264 1109 268 1113
rect 272 1109 276 1113
rect 1197 1109 1201 1113
rect 1205 1109 1209 1113
rect 7 1098 252 1102
rect 256 1098 272 1102
rect 288 1098 937 1102
rect 941 1098 1185 1102
rect 1189 1098 1205 1102
rect 1221 1098 1870 1102
rect 1874 1098 1952 1102
rect 280 1091 408 1094
rect 1213 1091 1341 1094
rect 295 1084 408 1087
rect 1228 1084 1341 1087
rect 264 1075 268 1079
rect 272 1075 276 1079
rect 1197 1075 1201 1079
rect 1205 1075 1209 1079
rect 148 1068 252 1071
rect 1081 1068 1185 1071
rect 17 1061 26 1065
rect 30 1061 62 1065
rect 66 1061 129 1065
rect 133 1061 158 1065
rect 162 1061 194 1065
rect 198 1061 261 1065
rect 265 1061 290 1065
rect 294 1061 326 1065
rect 330 1061 393 1065
rect 397 1061 477 1065
rect 950 1061 959 1065
rect 963 1061 995 1065
rect 999 1061 1062 1065
rect 1066 1061 1091 1065
rect 1095 1061 1127 1065
rect 1131 1061 1194 1065
rect 1198 1061 1223 1065
rect 1227 1061 1259 1065
rect 1263 1061 1326 1065
rect 1330 1061 1410 1065
rect 17 1054 50 1058
rect 54 1054 78 1058
rect 82 1054 108 1058
rect 112 1054 145 1058
rect 149 1054 182 1058
rect 186 1054 210 1058
rect 214 1054 240 1058
rect 244 1054 277 1058
rect 281 1054 314 1058
rect 318 1054 342 1058
rect 346 1054 372 1058
rect 376 1054 409 1058
rect 413 1054 417 1058
rect 950 1054 983 1058
rect 987 1054 1011 1058
rect 1015 1054 1041 1058
rect 1045 1054 1078 1058
rect 1082 1054 1115 1058
rect 1119 1054 1143 1058
rect 1147 1054 1173 1058
rect 1177 1054 1210 1058
rect 1214 1054 1247 1058
rect 1251 1054 1275 1058
rect 1279 1054 1305 1058
rect 1309 1054 1342 1058
rect 1346 1054 1350 1058
rect 20 1044 23 1054
rect 41 1044 44 1054
rect 57 1044 60 1054
rect 71 1047 76 1051
rect 80 1047 87 1051
rect 99 1044 102 1054
rect 115 1044 118 1054
rect 136 1044 139 1054
rect 152 1044 155 1054
rect 173 1044 176 1054
rect 189 1044 192 1054
rect 203 1047 208 1051
rect 212 1047 219 1051
rect 231 1044 234 1054
rect 247 1044 250 1054
rect 268 1044 271 1054
rect 284 1044 287 1054
rect 305 1044 308 1054
rect 321 1044 324 1054
rect 335 1047 340 1051
rect 344 1047 351 1051
rect 363 1044 366 1054
rect 379 1044 382 1054
rect 400 1044 403 1054
rect 953 1044 956 1054
rect 974 1044 977 1054
rect 990 1044 993 1054
rect 1004 1047 1009 1051
rect 1013 1047 1020 1051
rect 1032 1044 1035 1054
rect 1048 1044 1051 1054
rect 1069 1044 1072 1054
rect 1085 1044 1088 1054
rect 1106 1044 1109 1054
rect 1122 1044 1125 1054
rect 1136 1047 1141 1051
rect 1145 1047 1152 1051
rect 1164 1044 1167 1054
rect 1180 1044 1183 1054
rect 1201 1044 1204 1054
rect 1217 1044 1220 1054
rect 1238 1044 1241 1054
rect 1254 1044 1257 1054
rect 1268 1047 1273 1051
rect 1277 1047 1284 1051
rect 1296 1044 1299 1054
rect 1312 1044 1315 1054
rect 1333 1044 1336 1054
rect 37 1030 42 1033
rect 46 1030 70 1033
rect 95 1030 102 1033
rect 106 1030 128 1033
rect 148 1030 155 1033
rect 169 1030 174 1033
rect 178 1030 202 1033
rect 227 1030 234 1033
rect 238 1030 260 1033
rect 280 1030 287 1033
rect 301 1030 306 1033
rect 310 1030 334 1033
rect 359 1030 366 1033
rect 370 1030 392 1033
rect 53 1020 60 1023
rect 64 1024 83 1027
rect 83 1017 86 1023
rect 111 1020 118 1023
rect 122 1024 137 1027
rect 185 1020 192 1023
rect 196 1024 215 1027
rect 215 1017 218 1023
rect 243 1020 250 1023
rect 254 1024 269 1027
rect 317 1020 324 1023
rect 328 1024 347 1027
rect 347 1017 350 1023
rect 375 1020 382 1023
rect 386 1024 403 1027
rect 970 1030 975 1033
rect 979 1030 1003 1033
rect 1028 1030 1035 1033
rect 1039 1030 1061 1033
rect 1081 1030 1088 1033
rect 1102 1030 1107 1033
rect 1111 1030 1135 1033
rect 1160 1030 1167 1033
rect 1171 1030 1193 1033
rect 1213 1030 1220 1033
rect 1234 1030 1239 1033
rect 1243 1030 1267 1033
rect 1292 1030 1299 1033
rect 1303 1030 1325 1033
rect 986 1020 993 1023
rect 997 1024 1016 1027
rect 1016 1017 1019 1023
rect 1044 1020 1051 1023
rect 1055 1024 1070 1027
rect 1118 1020 1125 1023
rect 1129 1024 1148 1027
rect 1148 1017 1151 1023
rect 1176 1020 1183 1023
rect 1187 1024 1202 1027
rect 1250 1020 1257 1023
rect 1261 1024 1280 1027
rect 1280 1017 1283 1023
rect 1308 1020 1315 1023
rect 1319 1024 1336 1027
rect 20 1001 23 1013
rect 41 1001 44 1013
rect 57 1001 60 1013
rect 71 1004 83 1007
rect 99 1001 102 1013
rect 115 1001 118 1013
rect 136 1001 139 1013
rect 152 1001 155 1013
rect 173 1001 176 1013
rect 189 1001 192 1013
rect 203 1004 215 1007
rect 231 1001 234 1013
rect 247 1001 250 1013
rect 268 1001 271 1013
rect 284 1001 287 1013
rect 305 1001 308 1013
rect 321 1001 324 1013
rect 335 1004 347 1007
rect 363 1001 366 1013
rect 379 1001 382 1013
rect 400 1001 403 1013
rect 953 1001 956 1013
rect 974 1001 977 1013
rect 990 1001 993 1013
rect 1004 1004 1016 1007
rect 1032 1001 1035 1013
rect 1048 1001 1051 1013
rect 1069 1001 1072 1013
rect 1085 1001 1088 1013
rect 1106 1001 1109 1013
rect 1122 1001 1125 1013
rect 1136 1004 1148 1007
rect 1164 1001 1167 1013
rect 1180 1001 1183 1013
rect 1201 1001 1204 1013
rect 1217 1001 1220 1013
rect 1238 1001 1241 1013
rect 1254 1001 1257 1013
rect 1268 1004 1280 1007
rect 1296 1001 1299 1013
rect 1312 1001 1315 1013
rect 1333 1001 1336 1013
rect 17 997 50 1001
rect 54 997 78 1001
rect 82 997 108 1001
rect 112 997 182 1001
rect 186 997 210 1001
rect 214 997 240 1001
rect 244 997 314 1001
rect 318 997 342 1001
rect 346 997 372 1001
rect 376 997 429 1001
rect 950 997 983 1001
rect 987 997 1011 1001
rect 1015 997 1041 1001
rect 1045 997 1115 1001
rect 1119 997 1143 1001
rect 1147 997 1173 1001
rect 1177 997 1247 1001
rect 1251 997 1275 1001
rect 1279 997 1305 1001
rect 1309 997 1362 1001
rect 17 990 26 994
rect 30 990 77 994
rect 81 990 127 994
rect 131 990 158 994
rect 162 990 209 994
rect 213 990 259 994
rect 263 990 290 994
rect 294 990 341 994
rect 345 990 391 994
rect 395 990 465 994
rect 950 990 959 994
rect 963 990 1010 994
rect 1014 990 1060 994
rect 1064 990 1091 994
rect 1095 990 1142 994
rect 1146 990 1192 994
rect 1196 990 1223 994
rect 1227 990 1274 994
rect 1278 990 1324 994
rect 1328 990 1398 994
rect 483 982 498 986
rect 502 982 534 986
rect 538 982 601 986
rect 605 982 630 986
rect 634 982 666 986
rect 670 982 733 986
rect 737 982 762 986
rect 766 982 798 986
rect 802 982 865 986
rect 869 982 894 986
rect 898 982 930 986
rect 934 982 997 986
rect 1001 982 1017 986
rect 1416 982 1431 986
rect 1435 982 1467 986
rect 1471 982 1534 986
rect 1538 982 1563 986
rect 1567 982 1599 986
rect 1603 982 1666 986
rect 1670 982 1695 986
rect 1699 982 1731 986
rect 1735 982 1798 986
rect 1802 982 1827 986
rect 1831 982 1863 986
rect 1867 982 1930 986
rect 1934 982 1950 986
rect 423 975 522 979
rect 526 975 550 979
rect 554 975 580 979
rect 584 975 617 979
rect 621 975 654 979
rect 658 975 682 979
rect 686 975 712 979
rect 716 975 749 979
rect 753 975 786 979
rect 790 975 814 979
rect 818 975 844 979
rect 848 975 881 979
rect 885 975 918 979
rect 922 975 946 979
rect 950 975 976 979
rect 980 975 1013 979
rect 1356 975 1455 979
rect 1459 975 1483 979
rect 1487 975 1513 979
rect 1517 975 1550 979
rect 1554 975 1587 979
rect 1591 975 1615 979
rect 1619 975 1645 979
rect 1649 975 1682 979
rect 1686 975 1719 979
rect 1723 975 1747 979
rect 1751 975 1777 979
rect 1781 975 1814 979
rect 1818 975 1851 979
rect 1855 975 1879 979
rect 1883 975 1909 979
rect 1913 975 1946 979
rect 492 965 495 975
rect 513 965 516 975
rect 529 965 532 975
rect 543 968 548 972
rect 552 968 559 972
rect 571 965 574 975
rect 587 965 590 975
rect 608 965 611 975
rect 624 965 627 975
rect 645 965 648 975
rect 661 965 664 975
rect 675 968 680 972
rect 684 968 691 972
rect 703 965 706 975
rect 719 965 722 975
rect 740 965 743 975
rect 756 965 759 975
rect 777 965 780 975
rect 793 965 796 975
rect 807 968 812 972
rect 816 968 823 972
rect 835 965 838 975
rect 851 965 854 975
rect 872 965 875 975
rect 888 965 891 975
rect 909 965 912 975
rect 925 965 928 975
rect 939 968 944 972
rect 948 968 955 972
rect 967 965 970 975
rect 983 965 986 975
rect 1004 965 1007 975
rect 1425 965 1428 975
rect 1446 965 1449 975
rect 1462 965 1465 975
rect 1476 968 1481 972
rect 1485 968 1492 972
rect 1504 965 1507 975
rect 1520 965 1523 975
rect 1541 965 1544 975
rect 1557 965 1560 975
rect 1578 965 1581 975
rect 1594 965 1597 975
rect 1608 968 1613 972
rect 1617 968 1624 972
rect 1636 965 1639 975
rect 1652 965 1655 975
rect 1673 965 1676 975
rect 1689 965 1692 975
rect 1710 965 1713 975
rect 1726 965 1729 975
rect 1740 968 1745 972
rect 1749 968 1756 972
rect 1768 965 1771 975
rect 1784 965 1787 975
rect 1805 965 1808 975
rect 1821 965 1824 975
rect 1842 965 1845 975
rect 1858 965 1861 975
rect 1872 968 1877 972
rect 1881 968 1888 972
rect 1900 965 1903 975
rect 1916 965 1919 975
rect 1937 965 1940 975
rect 149 949 158 953
rect 162 949 194 953
rect 198 949 261 953
rect 265 949 477 953
rect 509 951 514 954
rect 518 951 542 954
rect 567 951 574 954
rect 578 951 600 954
rect 149 942 182 946
rect 186 942 210 946
rect 214 942 240 946
rect 244 942 277 946
rect 281 942 417 946
rect 152 932 155 942
rect 173 932 176 942
rect 189 932 192 942
rect 203 935 208 939
rect 212 935 219 939
rect 231 932 234 942
rect 247 932 250 942
rect 268 932 271 942
rect 525 941 532 944
rect 536 945 555 948
rect 555 938 558 944
rect 583 941 590 944
rect 594 945 611 948
rect 641 951 646 954
rect 650 951 674 954
rect 699 951 706 954
rect 710 951 732 954
rect 657 941 664 944
rect 668 945 687 948
rect 687 938 690 944
rect 715 941 722 944
rect 726 945 743 948
rect 773 951 778 954
rect 782 951 806 954
rect 831 951 838 954
rect 842 951 864 954
rect 789 941 796 944
rect 800 945 819 948
rect 819 938 822 944
rect 847 941 854 944
rect 858 945 875 948
rect 905 951 910 954
rect 914 951 938 954
rect 963 951 970 954
rect 974 951 996 954
rect 1082 949 1091 953
rect 1095 949 1127 953
rect 1131 949 1194 953
rect 1198 949 1410 953
rect 921 941 928 944
rect 932 945 951 948
rect 147 915 156 919
rect 169 918 174 921
rect 178 918 202 921
rect 227 918 234 921
rect 238 918 260 921
rect 492 922 495 934
rect 513 922 516 934
rect 529 922 532 934
rect 543 925 555 928
rect 571 922 574 934
rect 587 922 590 934
rect 608 922 611 934
rect 624 922 627 934
rect 645 922 648 934
rect 661 922 664 934
rect 675 925 687 928
rect 703 922 706 934
rect 719 922 722 934
rect 740 922 743 934
rect 756 922 759 934
rect 777 922 780 934
rect 793 922 796 934
rect 807 925 819 928
rect 835 922 838 934
rect 851 922 854 934
rect 872 922 875 934
rect 951 938 954 944
rect 979 941 986 944
rect 990 945 1007 948
rect 1442 951 1447 954
rect 1451 951 1475 954
rect 1500 951 1507 954
rect 1511 951 1533 954
rect 1082 942 1115 946
rect 1119 942 1143 946
rect 1147 942 1173 946
rect 1177 942 1210 946
rect 1214 942 1350 946
rect 888 922 891 934
rect 909 922 912 934
rect 925 922 928 934
rect 939 925 951 928
rect 967 922 970 934
rect 983 922 986 934
rect 1004 922 1007 934
rect 1085 932 1088 942
rect 1106 932 1109 942
rect 1122 932 1125 942
rect 1136 935 1141 939
rect 1145 935 1152 939
rect 1164 932 1167 942
rect 1180 932 1183 942
rect 1201 932 1204 942
rect 1458 941 1465 944
rect 1469 945 1488 948
rect 1488 938 1491 944
rect 1516 941 1523 944
rect 1527 945 1544 948
rect 1574 951 1579 954
rect 1583 951 1607 954
rect 1632 951 1639 954
rect 1643 951 1665 954
rect 1590 941 1597 944
rect 1601 945 1620 948
rect 1620 938 1623 944
rect 1648 941 1655 944
rect 1659 945 1676 948
rect 1706 951 1711 954
rect 1715 951 1739 954
rect 1764 951 1771 954
rect 1775 951 1797 954
rect 1722 941 1729 944
rect 1733 945 1752 948
rect 1752 938 1755 944
rect 1780 941 1787 944
rect 1791 945 1808 948
rect 1838 951 1843 954
rect 1847 951 1871 954
rect 1896 951 1903 954
rect 1907 951 1929 954
rect 1854 941 1861 944
rect 1865 945 1884 948
rect 435 918 522 922
rect 526 918 550 922
rect 554 918 580 922
rect 584 918 654 922
rect 658 918 682 922
rect 686 918 712 922
rect 716 918 786 922
rect 790 918 814 922
rect 818 918 844 922
rect 848 918 918 922
rect 922 918 946 922
rect 950 918 976 922
rect 980 918 1017 922
rect 185 908 192 911
rect 196 912 215 915
rect 215 905 218 911
rect 243 908 250 911
rect 254 912 269 915
rect 1080 915 1089 919
rect 1102 918 1107 921
rect 1111 918 1135 921
rect 1160 918 1167 921
rect 1171 918 1193 921
rect 1425 922 1428 934
rect 1446 922 1449 934
rect 1462 922 1465 934
rect 1476 925 1488 928
rect 1504 922 1507 934
rect 1520 922 1523 934
rect 1541 922 1544 934
rect 1557 922 1560 934
rect 1578 922 1581 934
rect 1594 922 1597 934
rect 1608 925 1620 928
rect 1636 922 1639 934
rect 1652 922 1655 934
rect 1673 922 1676 934
rect 1689 922 1692 934
rect 1710 922 1713 934
rect 1726 922 1729 934
rect 1740 925 1752 928
rect 1768 922 1771 934
rect 1784 922 1787 934
rect 1805 922 1808 934
rect 1884 938 1887 944
rect 1912 941 1919 944
rect 1923 945 1940 948
rect 1821 922 1824 934
rect 1842 922 1845 934
rect 1858 922 1861 934
rect 1872 925 1884 928
rect 1900 922 1903 934
rect 1916 922 1919 934
rect 1937 922 1940 934
rect 1368 918 1455 922
rect 1459 918 1483 922
rect 1487 918 1513 922
rect 1517 918 1587 922
rect 1591 918 1615 922
rect 1619 918 1645 922
rect 1649 918 1719 922
rect 1723 918 1747 922
rect 1751 918 1777 922
rect 1781 918 1851 922
rect 1855 918 1879 922
rect 1883 918 1909 922
rect 1913 918 1950 922
rect 471 911 498 915
rect 502 911 549 915
rect 553 911 599 915
rect 603 911 630 915
rect 634 911 681 915
rect 685 911 731 915
rect 735 911 762 915
rect 766 911 813 915
rect 817 911 863 915
rect 867 911 894 915
rect 898 911 945 915
rect 949 911 995 915
rect 999 911 1017 915
rect 1118 908 1125 911
rect 1129 912 1148 915
rect 152 889 155 901
rect 173 889 176 901
rect 189 889 192 901
rect 203 892 215 895
rect 231 889 234 901
rect 247 889 250 901
rect 268 889 271 901
rect 423 898 496 902
rect 500 898 512 902
rect 516 898 530 902
rect 534 898 541 902
rect 545 898 547 902
rect 551 898 566 902
rect 570 898 603 902
rect 607 898 608 902
rect 612 898 620 902
rect 624 898 648 902
rect 652 898 664 902
rect 668 898 688 902
rect 692 898 742 902
rect 746 898 769 902
rect 773 898 823 902
rect 827 898 846 902
rect 1148 905 1151 911
rect 1176 908 1183 911
rect 1187 912 1202 915
rect 1404 911 1431 915
rect 1435 911 1482 915
rect 1486 911 1532 915
rect 1536 911 1563 915
rect 1567 911 1614 915
rect 1618 911 1664 915
rect 1668 911 1695 915
rect 1699 911 1746 915
rect 1750 911 1796 915
rect 1800 911 1827 915
rect 1831 911 1878 915
rect 1882 911 1928 915
rect 1932 911 1950 915
rect 459 891 523 895
rect 527 891 554 895
rect 558 891 576 895
rect 580 891 641 895
rect 645 891 659 895
rect 671 894 674 898
rect 149 885 182 889
rect 186 885 210 889
rect 214 885 240 889
rect 244 885 429 889
rect 149 878 158 882
rect 162 878 209 882
rect 213 878 259 882
rect 263 878 465 882
rect 566 884 569 888
rect 593 884 594 888
rect 638 884 640 888
rect 680 881 683 886
rect 695 888 698 898
rect 725 894 728 898
rect 752 894 755 898
rect 147 862 163 866
rect 272 864 276 868
rect 288 864 292 868
rect 296 864 498 868
rect 506 867 509 873
rect 513 867 516 873
rect 506 864 516 867
rect 506 859 509 864
rect 155 855 159 859
rect 171 855 292 859
rect 513 859 516 864
rect 522 869 525 873
rect 522 865 524 869
rect 528 865 530 869
rect 538 868 541 873
rect 566 870 569 873
rect 538 866 549 868
rect 522 859 525 865
rect 538 864 544 866
rect 538 859 541 864
rect 548 864 549 866
rect 567 866 569 870
rect 566 859 569 866
rect 669 877 672 880
rect 711 877 714 880
rect 582 869 585 873
rect 592 869 595 873
rect 592 865 601 869
rect 613 868 616 873
rect 638 869 641 873
rect 582 859 585 865
rect 592 859 595 865
rect 613 864 614 868
rect 618 864 621 867
rect 640 865 641 869
rect 656 868 659 873
rect 680 872 683 877
rect 688 873 699 876
rect 711 874 719 877
rect 613 859 616 864
rect 638 859 641 865
rect 656 859 659 864
rect 142 847 158 851
rect 162 847 225 851
rect 229 847 261 851
rect 265 847 477 851
rect 558 846 559 850
rect 583 847 584 851
rect 630 846 631 850
rect 146 840 179 844
rect 183 840 209 844
rect 213 840 237 844
rect 241 840 417 844
rect 152 830 155 840
rect 173 830 176 840
rect 189 830 192 840
rect 204 833 211 837
rect 215 833 220 837
rect 231 830 234 840
rect 247 830 250 840
rect 268 830 271 840
rect 447 839 511 843
rect 515 839 570 843
rect 574 839 595 843
rect 599 839 626 843
rect 630 839 659 843
rect 671 836 674 868
rect 688 867 691 873
rect 711 868 714 874
rect 723 869 726 872
rect 734 872 737 886
rect 761 881 764 886
rect 776 888 779 898
rect 806 894 809 898
rect 745 877 746 880
rect 750 877 753 880
rect 1085 889 1088 901
rect 1106 889 1109 901
rect 1122 889 1125 901
rect 1136 892 1148 895
rect 1164 889 1167 901
rect 1180 889 1183 901
rect 1201 889 1204 901
rect 1356 898 1429 902
rect 1433 898 1445 902
rect 1449 898 1463 902
rect 1467 898 1474 902
rect 1478 898 1480 902
rect 1484 898 1499 902
rect 1503 898 1536 902
rect 1540 898 1541 902
rect 1545 898 1553 902
rect 1557 898 1581 902
rect 1585 898 1597 902
rect 1601 898 1621 902
rect 1625 898 1675 902
rect 1679 898 1702 902
rect 1706 898 1756 902
rect 1760 898 1779 902
rect 1392 891 1456 895
rect 1460 891 1487 895
rect 1491 891 1509 895
rect 1513 891 1574 895
rect 1578 891 1592 895
rect 1604 894 1607 898
rect 792 877 795 880
rect 734 869 742 872
rect 761 872 764 877
rect 734 864 737 869
rect 742 865 746 869
rect 769 873 780 876
rect 792 874 800 877
rect 686 858 691 863
rect 695 836 698 864
rect 725 836 728 860
rect 752 836 755 868
rect 769 867 772 873
rect 792 868 795 874
rect 804 869 807 872
rect 815 872 818 886
rect 1082 885 1115 889
rect 1119 885 1143 889
rect 1147 885 1173 889
rect 1177 885 1362 889
rect 1082 878 1091 882
rect 1095 878 1142 882
rect 1146 878 1192 882
rect 1196 878 1398 882
rect 1499 884 1502 888
rect 1526 884 1527 888
rect 1571 884 1573 888
rect 1613 881 1616 886
rect 1628 888 1631 898
rect 1658 894 1661 898
rect 1685 894 1688 898
rect 815 869 827 872
rect 815 864 818 869
rect 767 858 772 863
rect 776 836 779 864
rect 1080 862 1096 866
rect 1205 864 1209 868
rect 1221 864 1225 868
rect 1229 864 1431 868
rect 1439 867 1442 873
rect 1446 867 1449 873
rect 1439 864 1449 867
rect 806 836 809 860
rect 1439 859 1442 864
rect 1088 855 1092 859
rect 1104 855 1225 859
rect 1446 859 1449 864
rect 1455 869 1458 873
rect 1455 865 1457 869
rect 1461 865 1463 869
rect 1471 868 1474 873
rect 1499 870 1502 873
rect 1471 866 1482 868
rect 1455 859 1458 865
rect 1471 864 1477 866
rect 1471 859 1474 864
rect 1481 864 1482 866
rect 1500 866 1502 870
rect 1499 859 1502 866
rect 1602 877 1605 880
rect 1644 877 1647 880
rect 1515 869 1518 873
rect 1525 869 1528 873
rect 1525 865 1534 869
rect 1546 868 1549 873
rect 1571 869 1574 873
rect 1515 859 1518 865
rect 1525 859 1528 865
rect 1546 864 1547 868
rect 1551 864 1554 867
rect 1573 865 1574 869
rect 1589 868 1592 873
rect 1613 872 1616 877
rect 1621 873 1632 876
rect 1644 874 1652 877
rect 1546 859 1549 864
rect 1571 859 1574 865
rect 1589 859 1592 864
rect 1075 847 1091 851
rect 1095 847 1158 851
rect 1162 847 1194 851
rect 1198 847 1410 851
rect 1491 846 1492 850
rect 1516 847 1517 851
rect 1563 846 1564 850
rect 1079 840 1112 844
rect 1116 840 1142 844
rect 1146 840 1170 844
rect 1174 840 1350 844
rect 435 832 497 836
rect 501 832 503 836
rect 507 832 511 836
rect 515 832 529 836
rect 533 832 538 836
rect 542 832 547 836
rect 551 832 570 836
rect 574 832 604 836
rect 608 832 619 836
rect 623 832 647 836
rect 651 832 664 836
rect 668 832 688 836
rect 692 832 742 836
rect 749 832 769 836
rect 773 832 823 836
rect 163 816 185 819
rect 189 816 196 819
rect 447 825 511 829
rect 515 825 570 829
rect 574 825 595 829
rect 599 825 626 829
rect 630 825 659 829
rect 221 816 245 819
rect 249 816 254 819
rect 558 818 559 822
rect 583 817 584 821
rect 630 818 631 822
rect 267 813 276 817
rect 154 810 169 813
rect 208 810 227 813
rect 173 806 180 809
rect 205 803 208 809
rect 231 806 238 809
rect 506 804 509 809
rect 513 804 516 809
rect 496 801 498 804
rect 506 801 516 804
rect 152 787 155 799
rect 173 787 176 799
rect 189 787 192 799
rect 208 790 220 793
rect 231 787 234 799
rect 247 787 250 799
rect 268 787 271 799
rect 506 795 509 801
rect 513 795 516 801
rect 522 803 525 809
rect 538 804 541 809
rect 522 799 524 803
rect 528 799 530 803
rect 538 802 544 804
rect 548 802 549 804
rect 538 800 549 802
rect 566 802 569 809
rect 522 795 525 799
rect 538 795 541 800
rect 567 798 569 802
rect 566 795 569 798
rect 582 803 585 809
rect 592 803 595 809
rect 613 804 616 809
rect 592 799 601 803
rect 613 800 614 804
rect 618 801 621 804
rect 638 803 641 809
rect 656 804 659 809
rect 695 812 698 832
rect 776 812 779 832
rect 1085 830 1088 840
rect 1106 830 1109 840
rect 1122 830 1125 840
rect 1137 833 1144 837
rect 1148 833 1153 837
rect 1164 830 1167 840
rect 1180 830 1183 840
rect 1201 830 1204 840
rect 1380 839 1444 843
rect 1448 839 1503 843
rect 1507 839 1528 843
rect 1532 839 1559 843
rect 1563 839 1592 843
rect 1604 836 1607 868
rect 1621 867 1624 873
rect 1644 868 1647 874
rect 1656 869 1659 872
rect 1667 872 1670 886
rect 1694 881 1697 886
rect 1709 888 1712 898
rect 1739 894 1742 898
rect 1678 877 1679 880
rect 1683 877 1686 880
rect 1725 877 1728 880
rect 1667 869 1675 872
rect 1694 872 1697 877
rect 1667 864 1670 869
rect 1675 865 1679 869
rect 1702 873 1713 876
rect 1725 874 1733 877
rect 1619 858 1624 863
rect 1628 836 1631 864
rect 1658 836 1661 860
rect 1685 836 1688 868
rect 1702 867 1705 873
rect 1725 868 1728 874
rect 1737 869 1740 872
rect 1748 872 1751 886
rect 1748 869 1760 872
rect 1748 864 1751 869
rect 1700 858 1705 863
rect 1709 836 1712 864
rect 1739 836 1742 860
rect 1368 832 1430 836
rect 1434 832 1436 836
rect 1440 832 1444 836
rect 1448 832 1462 836
rect 1466 832 1471 836
rect 1475 832 1480 836
rect 1484 832 1503 836
rect 1507 832 1537 836
rect 1541 832 1552 836
rect 1556 832 1580 836
rect 1584 832 1597 836
rect 1601 832 1621 836
rect 1625 832 1675 836
rect 1682 832 1702 836
rect 1706 832 1756 836
rect 1096 816 1118 819
rect 1122 816 1129 819
rect 1380 825 1444 829
rect 1448 825 1503 829
rect 1507 825 1528 829
rect 1532 825 1559 829
rect 1563 825 1592 829
rect 1154 816 1178 819
rect 1182 816 1187 819
rect 1491 818 1492 822
rect 1516 817 1517 821
rect 1563 818 1564 822
rect 1200 813 1209 817
rect 1087 810 1102 813
rect 582 795 585 799
rect 592 795 595 799
rect 613 795 616 800
rect 640 799 641 803
rect 638 795 641 799
rect 656 795 659 800
rect 686 799 691 804
rect 695 800 696 803
rect 711 802 714 808
rect 711 799 719 802
rect 766 799 771 804
rect 775 800 777 803
rect 792 802 795 808
rect 1141 810 1160 813
rect 1106 806 1113 809
rect 1138 803 1141 809
rect 792 799 800 802
rect 1164 806 1171 809
rect 1439 804 1442 809
rect 1446 804 1449 809
rect 1429 801 1431 804
rect 1439 801 1449 804
rect 711 796 714 799
rect 792 796 795 799
rect 142 783 179 787
rect 183 783 209 787
rect 213 783 237 787
rect 241 783 429 787
rect 566 780 569 784
rect 593 780 594 784
rect 638 780 640 784
rect 142 776 160 780
rect 164 776 210 780
rect 214 776 261 780
rect 265 776 465 780
rect 511 773 523 777
rect 527 773 554 777
rect 558 773 576 777
rect 580 773 641 777
rect 645 773 659 777
rect 695 770 698 788
rect 776 770 779 788
rect 1085 787 1088 799
rect 1106 787 1109 799
rect 1122 787 1125 799
rect 1141 790 1153 793
rect 1164 787 1167 799
rect 1180 787 1183 799
rect 1201 787 1204 799
rect 1439 795 1442 801
rect 1446 795 1449 801
rect 1455 803 1458 809
rect 1471 804 1474 809
rect 1455 799 1457 803
rect 1461 799 1463 803
rect 1471 802 1477 804
rect 1481 802 1482 804
rect 1471 800 1482 802
rect 1499 802 1502 809
rect 1455 795 1458 799
rect 1471 795 1474 800
rect 1500 798 1502 802
rect 1499 795 1502 798
rect 1515 803 1518 809
rect 1525 803 1528 809
rect 1546 804 1549 809
rect 1525 799 1534 803
rect 1546 800 1547 804
rect 1551 801 1554 804
rect 1571 803 1574 809
rect 1589 804 1592 809
rect 1628 812 1631 832
rect 1709 812 1712 832
rect 1515 795 1518 799
rect 1525 795 1528 799
rect 1546 795 1549 800
rect 1573 799 1574 803
rect 1571 795 1574 799
rect 1589 795 1592 800
rect 1619 799 1624 804
rect 1628 800 1629 803
rect 1644 802 1647 808
rect 1644 799 1652 802
rect 1699 799 1704 804
rect 1708 800 1710 803
rect 1725 802 1728 808
rect 1725 799 1733 802
rect 1644 796 1647 799
rect 1725 796 1728 799
rect 1075 783 1112 787
rect 1116 783 1142 787
rect 1146 783 1170 787
rect 1174 783 1362 787
rect 1499 780 1502 784
rect 1526 780 1527 784
rect 1571 780 1573 784
rect 1075 776 1093 780
rect 1097 776 1143 780
rect 1147 776 1194 780
rect 1198 776 1398 780
rect 1444 773 1456 777
rect 1460 773 1487 777
rect 1491 773 1509 777
rect 1513 773 1574 777
rect 1578 773 1592 777
rect 1628 770 1631 788
rect 1709 770 1712 788
rect 423 766 496 770
rect 500 766 512 770
rect 516 766 530 770
rect 534 766 541 770
rect 545 766 547 770
rect 551 766 566 770
rect 570 766 603 770
rect 607 766 608 770
rect 612 766 620 770
rect 624 766 648 770
rect 652 766 664 770
rect 668 766 688 770
rect 692 766 742 770
rect 746 766 769 770
rect 773 766 831 770
rect 835 766 846 770
rect 1356 766 1429 770
rect 1433 766 1445 770
rect 1449 766 1463 770
rect 1467 766 1474 770
rect 1478 766 1480 770
rect 1484 766 1499 770
rect 1503 766 1536 770
rect 1540 766 1541 770
rect 1545 766 1553 770
rect 1557 766 1581 770
rect 1585 766 1597 770
rect 1601 766 1621 770
rect 1625 766 1675 770
rect 1679 766 1702 770
rect 1706 766 1764 770
rect 1768 766 1779 770
rect 459 759 507 763
rect 511 759 523 763
rect 527 759 554 763
rect 558 759 576 763
rect 580 759 641 763
rect 645 759 659 763
rect 695 756 698 766
rect 725 762 728 766
rect 776 762 779 766
rect 566 752 569 756
rect 593 752 594 756
rect 638 752 640 756
rect 495 732 498 735
rect 506 735 509 741
rect 513 735 516 741
rect 506 732 516 735
rect 506 727 509 732
rect 513 727 516 732
rect 522 737 525 741
rect 522 733 524 737
rect 528 733 530 737
rect 538 736 541 741
rect 566 738 569 741
rect 538 734 549 736
rect 522 727 525 733
rect 538 732 544 734
rect 538 727 541 732
rect 548 732 549 734
rect 567 734 569 738
rect 566 727 569 734
rect 711 745 714 748
rect 582 737 585 741
rect 592 737 595 741
rect 592 733 601 737
rect 613 736 616 741
rect 638 737 641 741
rect 582 727 585 733
rect 592 727 595 733
rect 613 732 614 736
rect 618 732 621 735
rect 640 733 641 737
rect 656 736 659 741
rect 688 741 699 744
rect 711 742 719 745
rect 613 727 616 732
rect 638 727 641 733
rect 688 735 691 741
rect 711 736 714 742
rect 723 737 726 740
rect 734 740 737 754
rect 785 749 788 754
rect 800 756 803 766
rect 830 762 833 766
rect 769 745 770 748
rect 774 745 777 748
rect 1392 759 1440 763
rect 1444 759 1456 763
rect 1460 759 1487 763
rect 1491 759 1509 763
rect 1513 759 1574 763
rect 1578 759 1592 763
rect 1628 756 1631 766
rect 1658 762 1661 766
rect 1709 762 1712 766
rect 816 745 819 748
rect 742 740 747 745
rect 785 740 788 745
rect 734 737 742 740
rect 656 727 659 732
rect 734 732 737 737
rect 793 741 804 744
rect 816 742 824 745
rect 686 726 691 731
rect 558 714 559 718
rect 583 715 584 719
rect 630 714 631 718
rect 447 707 511 711
rect 515 707 570 711
rect 574 707 595 711
rect 599 707 626 711
rect 630 707 659 711
rect 695 704 698 732
rect 725 704 728 728
rect 776 704 779 736
rect 793 735 796 741
rect 816 736 819 742
rect 828 737 831 740
rect 839 740 842 754
rect 1499 752 1502 756
rect 1526 752 1527 756
rect 1571 752 1573 756
rect 839 737 845 740
rect 839 732 842 737
rect 1428 732 1431 735
rect 1439 735 1442 741
rect 1446 735 1449 741
rect 1439 732 1449 735
rect 791 726 796 731
rect 800 704 803 732
rect 830 704 833 728
rect 1439 727 1442 732
rect 1446 727 1449 732
rect 1455 737 1458 741
rect 1455 733 1457 737
rect 1461 733 1463 737
rect 1471 736 1474 741
rect 1499 738 1502 741
rect 1471 734 1482 736
rect 1455 727 1458 733
rect 1471 732 1477 734
rect 1471 727 1474 732
rect 1481 732 1482 734
rect 1500 734 1502 738
rect 1499 727 1502 734
rect 1644 745 1647 748
rect 1515 737 1518 741
rect 1525 737 1528 741
rect 1525 733 1534 737
rect 1546 736 1549 741
rect 1571 737 1574 741
rect 1515 727 1518 733
rect 1525 727 1528 733
rect 1546 732 1547 736
rect 1551 732 1554 735
rect 1573 733 1574 737
rect 1589 736 1592 741
rect 1621 741 1632 744
rect 1644 742 1652 745
rect 1546 727 1549 732
rect 1571 727 1574 733
rect 1621 735 1624 741
rect 1644 736 1647 742
rect 1656 737 1659 740
rect 1667 740 1670 754
rect 1718 749 1721 754
rect 1733 756 1736 766
rect 1763 762 1766 766
rect 1702 745 1703 748
rect 1707 745 1710 748
rect 1749 745 1752 748
rect 1675 740 1680 745
rect 1718 740 1721 745
rect 1667 737 1675 740
rect 1589 727 1592 732
rect 1667 732 1670 737
rect 1726 741 1737 744
rect 1749 742 1757 745
rect 1619 726 1624 731
rect 1491 714 1492 718
rect 1516 715 1517 719
rect 1563 714 1564 718
rect 1380 707 1444 711
rect 1448 707 1503 711
rect 1507 707 1528 711
rect 1532 707 1559 711
rect 1563 707 1592 711
rect 1628 704 1631 732
rect 1658 704 1661 728
rect 1709 704 1712 736
rect 1726 735 1729 741
rect 1749 736 1752 742
rect 1761 737 1764 740
rect 1772 740 1775 754
rect 1772 737 1778 740
rect 1772 732 1775 737
rect 1724 726 1729 731
rect 1733 704 1736 732
rect 1763 704 1766 728
rect 435 700 497 704
rect 501 700 503 704
rect 507 700 511 704
rect 515 700 529 704
rect 533 700 538 704
rect 542 700 547 704
rect 551 700 570 704
rect 574 700 604 704
rect 608 700 619 704
rect 623 700 647 704
rect 651 700 664 704
rect 668 700 688 704
rect 692 700 742 704
rect 746 700 769 704
rect 773 700 793 704
rect 797 700 845 704
rect 1368 700 1430 704
rect 1434 700 1436 704
rect 1440 700 1444 704
rect 1448 700 1462 704
rect 1466 700 1471 704
rect 1475 700 1480 704
rect 1484 700 1503 704
rect 1507 700 1537 704
rect 1541 700 1552 704
rect 1556 700 1580 704
rect 1584 700 1597 704
rect 1601 700 1621 704
rect 1625 700 1675 704
rect 1679 700 1702 704
rect 1706 700 1726 704
rect 1730 700 1778 704
rect 447 693 511 697
rect 515 693 570 697
rect 574 693 595 697
rect 599 693 626 697
rect 630 693 659 697
rect 558 686 559 690
rect 583 685 584 689
rect 630 686 631 690
rect 695 681 698 700
rect 800 681 803 700
rect 1380 693 1444 697
rect 1448 693 1503 697
rect 1507 693 1528 697
rect 1532 693 1559 697
rect 1563 693 1592 697
rect 1491 686 1492 690
rect 1516 685 1517 689
rect 1563 686 1564 690
rect 1628 681 1631 700
rect 1733 681 1736 700
rect 506 672 509 677
rect 513 672 516 677
rect 496 669 498 672
rect 506 669 516 672
rect 506 663 509 669
rect 513 663 516 669
rect 522 671 525 677
rect 538 672 541 677
rect 522 667 524 671
rect 528 667 530 671
rect 538 670 544 672
rect 548 670 549 672
rect 538 668 549 670
rect 566 670 569 677
rect 522 663 525 667
rect 538 663 541 668
rect 567 666 569 670
rect 566 663 569 666
rect 582 671 585 677
rect 592 671 595 677
rect 613 672 616 677
rect 592 667 601 671
rect 613 668 614 672
rect 618 669 621 672
rect 638 671 641 677
rect 656 672 659 677
rect 582 663 585 667
rect 592 663 595 667
rect 613 663 616 668
rect 640 667 641 671
rect 685 668 690 673
rect 694 669 696 672
rect 711 671 714 677
rect 711 668 719 671
rect 791 668 796 673
rect 800 669 801 672
rect 816 671 819 677
rect 816 668 824 671
rect 1439 672 1442 677
rect 1446 672 1449 677
rect 1429 669 1431 672
rect 1439 669 1449 672
rect 638 663 641 667
rect 656 663 659 668
rect 711 665 714 668
rect 816 665 819 668
rect 1439 663 1442 669
rect 566 648 569 652
rect 593 648 594 652
rect 638 648 640 652
rect 459 641 523 645
rect 527 641 554 645
rect 558 641 576 645
rect 580 641 641 645
rect 645 641 659 645
rect 695 638 698 657
rect 800 638 803 657
rect 1446 663 1449 669
rect 1455 671 1458 677
rect 1471 672 1474 677
rect 1455 667 1457 671
rect 1461 667 1463 671
rect 1471 670 1477 672
rect 1481 670 1482 672
rect 1471 668 1482 670
rect 1499 670 1502 677
rect 1455 663 1458 667
rect 1471 663 1474 668
rect 1500 666 1502 670
rect 1499 663 1502 666
rect 1515 671 1518 677
rect 1525 671 1528 677
rect 1546 672 1549 677
rect 1525 667 1534 671
rect 1546 668 1547 672
rect 1551 669 1554 672
rect 1571 671 1574 677
rect 1589 672 1592 677
rect 1515 663 1518 667
rect 1525 663 1528 667
rect 1546 663 1549 668
rect 1573 667 1574 671
rect 1618 668 1623 673
rect 1627 669 1629 672
rect 1644 671 1647 677
rect 1644 668 1652 671
rect 1724 668 1729 673
rect 1733 669 1734 672
rect 1749 671 1752 677
rect 1749 668 1757 671
rect 1571 663 1574 667
rect 1589 663 1592 668
rect 1644 665 1647 668
rect 1749 665 1752 668
rect 1499 648 1502 652
rect 1526 648 1527 652
rect 1571 648 1573 652
rect 1392 641 1456 645
rect 1460 641 1487 645
rect 1491 641 1509 645
rect 1513 641 1574 645
rect 1578 641 1592 645
rect 1628 638 1631 657
rect 1733 638 1736 657
rect 423 634 496 638
rect 500 634 512 638
rect 516 634 530 638
rect 534 634 541 638
rect 545 634 547 638
rect 551 634 566 638
rect 570 634 603 638
rect 607 634 608 638
rect 612 634 620 638
rect 624 634 648 638
rect 652 634 664 638
rect 668 634 688 638
rect 692 634 742 638
rect 746 634 769 638
rect 773 634 823 638
rect 827 634 831 638
rect 835 634 859 638
rect 863 634 913 638
rect 1356 634 1429 638
rect 1433 634 1445 638
rect 1449 634 1463 638
rect 1467 634 1474 638
rect 1478 634 1480 638
rect 1484 634 1499 638
rect 1503 634 1536 638
rect 1540 634 1541 638
rect 1545 634 1553 638
rect 1557 634 1581 638
rect 1585 634 1597 638
rect 1601 634 1621 638
rect 1625 634 1675 638
rect 1679 634 1702 638
rect 1706 634 1756 638
rect 1760 634 1764 638
rect 1768 634 1792 638
rect 1796 634 1846 638
rect 459 627 523 631
rect 527 627 554 631
rect 558 627 576 631
rect 580 627 641 631
rect 645 627 659 631
rect 695 624 698 634
rect 725 630 728 634
rect 752 630 755 634
rect 566 620 569 624
rect 593 620 594 624
rect 638 620 640 624
rect 495 600 498 603
rect 506 603 509 609
rect 513 603 516 609
rect 506 600 516 603
rect 506 595 509 600
rect 513 595 516 600
rect 522 605 525 609
rect 522 601 524 605
rect 528 601 530 605
rect 538 604 541 609
rect 566 606 569 609
rect 538 602 549 604
rect 522 595 525 601
rect 538 600 544 602
rect 538 595 541 600
rect 548 600 549 602
rect 567 602 569 606
rect 566 595 569 602
rect 711 613 714 616
rect 582 605 585 609
rect 592 605 595 609
rect 592 601 601 605
rect 613 604 616 609
rect 638 605 641 609
rect 582 595 585 601
rect 592 595 595 601
rect 613 600 614 604
rect 618 600 621 603
rect 640 601 641 605
rect 656 604 659 609
rect 688 609 699 612
rect 711 610 719 613
rect 613 595 616 600
rect 638 595 641 601
rect 688 603 691 609
rect 711 604 714 610
rect 723 605 726 608
rect 734 608 737 622
rect 761 617 764 622
rect 776 624 779 634
rect 806 630 809 634
rect 842 630 845 634
rect 745 613 746 616
rect 750 613 753 616
rect 792 613 795 616
rect 734 605 742 608
rect 761 608 764 613
rect 656 595 659 600
rect 734 600 737 605
rect 742 601 746 605
rect 769 609 780 612
rect 792 610 800 613
rect 686 594 691 599
rect 558 582 559 586
rect 583 583 584 587
rect 630 582 631 586
rect 447 575 511 579
rect 515 575 570 579
rect 574 575 595 579
rect 599 575 626 579
rect 630 575 659 579
rect 695 572 698 600
rect 725 572 728 596
rect 752 572 755 604
rect 769 603 772 609
rect 792 604 795 610
rect 804 605 807 608
rect 815 608 818 622
rect 851 617 854 622
rect 866 624 869 634
rect 896 630 899 634
rect 840 613 843 616
rect 1392 627 1456 631
rect 1460 627 1487 631
rect 1491 627 1509 631
rect 1513 627 1574 631
rect 1578 627 1592 631
rect 1628 624 1631 634
rect 1658 630 1661 634
rect 1685 630 1688 634
rect 882 613 885 616
rect 815 605 824 608
rect 851 608 854 613
rect 815 600 818 605
rect 767 594 772 599
rect 776 572 779 600
rect 858 611 870 612
rect 862 609 870 611
rect 882 610 890 613
rect 882 604 885 610
rect 894 605 897 608
rect 905 608 908 622
rect 1499 620 1502 624
rect 1526 620 1527 624
rect 1571 620 1573 624
rect 905 605 925 608
rect 806 572 809 596
rect 842 572 845 604
rect 905 600 908 605
rect 1428 600 1431 603
rect 1439 603 1442 609
rect 1446 603 1449 609
rect 1439 600 1449 603
rect 866 572 869 600
rect 896 572 899 596
rect 1439 595 1442 600
rect 1446 595 1449 600
rect 1455 605 1458 609
rect 1455 601 1457 605
rect 1461 601 1463 605
rect 1471 604 1474 609
rect 1499 606 1502 609
rect 1471 602 1482 604
rect 1455 595 1458 601
rect 1471 600 1477 602
rect 1471 595 1474 600
rect 1481 600 1482 602
rect 1500 602 1502 606
rect 1499 595 1502 602
rect 1644 613 1647 616
rect 1515 605 1518 609
rect 1525 605 1528 609
rect 1525 601 1534 605
rect 1546 604 1549 609
rect 1571 605 1574 609
rect 1515 595 1518 601
rect 1525 595 1528 601
rect 1546 600 1547 604
rect 1551 600 1554 603
rect 1573 601 1574 605
rect 1589 604 1592 609
rect 1621 609 1632 612
rect 1644 610 1652 613
rect 1546 595 1549 600
rect 1571 595 1574 601
rect 1621 603 1624 609
rect 1644 604 1647 610
rect 1656 605 1659 608
rect 1667 608 1670 622
rect 1694 617 1697 622
rect 1709 624 1712 634
rect 1739 630 1742 634
rect 1775 630 1778 634
rect 1678 613 1679 616
rect 1683 613 1686 616
rect 1725 613 1728 616
rect 1667 605 1675 608
rect 1694 608 1697 613
rect 1589 595 1592 600
rect 1667 600 1670 605
rect 1675 601 1679 605
rect 1702 609 1713 612
rect 1725 610 1733 613
rect 1619 594 1624 599
rect 1491 582 1492 586
rect 1516 583 1517 587
rect 1563 582 1564 586
rect 1380 575 1444 579
rect 1448 575 1503 579
rect 1507 575 1528 579
rect 1532 575 1559 579
rect 1563 575 1592 579
rect 1628 572 1631 600
rect 1658 572 1661 596
rect 1685 572 1688 604
rect 1702 603 1705 609
rect 1725 604 1728 610
rect 1737 605 1740 608
rect 1748 608 1751 622
rect 1784 617 1787 622
rect 1799 624 1802 634
rect 1829 630 1832 634
rect 1773 613 1776 616
rect 1815 613 1818 616
rect 1748 605 1757 608
rect 1784 608 1787 613
rect 1748 600 1751 605
rect 1700 594 1705 599
rect 1709 572 1712 600
rect 1791 611 1803 612
rect 1795 609 1803 611
rect 1815 610 1823 613
rect 1815 604 1818 610
rect 1827 605 1830 608
rect 1838 608 1841 622
rect 1838 605 1858 608
rect 1739 572 1742 596
rect 1775 572 1778 604
rect 1838 600 1841 605
rect 1799 572 1802 600
rect 1829 572 1832 596
rect 435 568 497 572
rect 501 568 503 572
rect 507 568 511 572
rect 515 568 529 572
rect 533 568 538 572
rect 542 568 547 572
rect 551 568 570 572
rect 574 568 604 572
rect 608 568 619 572
rect 623 568 647 572
rect 651 568 664 572
rect 668 568 688 572
rect 692 568 742 572
rect 749 568 769 572
rect 773 568 823 572
rect 827 568 859 572
rect 863 568 913 572
rect 1368 568 1430 572
rect 1434 568 1436 572
rect 1440 568 1444 572
rect 1448 568 1462 572
rect 1466 568 1471 572
rect 1475 568 1480 572
rect 1484 568 1503 572
rect 1507 568 1537 572
rect 1541 568 1552 572
rect 1556 568 1580 572
rect 1584 568 1597 572
rect 1601 568 1621 572
rect 1625 568 1675 572
rect 1682 568 1702 572
rect 1706 568 1756 572
rect 1760 568 1792 572
rect 1796 568 1846 572
rect 447 561 511 565
rect 515 561 570 565
rect 574 561 595 565
rect 599 561 626 565
rect 630 561 659 565
rect 558 554 559 558
rect 583 553 584 557
rect 630 554 631 558
rect 506 540 509 545
rect 513 540 516 545
rect 496 537 498 540
rect 506 537 516 540
rect 506 531 509 537
rect 513 531 516 537
rect 522 539 525 545
rect 538 540 541 545
rect 522 535 524 539
rect 528 535 530 539
rect 538 538 544 540
rect 548 538 549 540
rect 538 536 549 538
rect 566 538 569 545
rect 522 531 525 535
rect 538 531 541 536
rect 567 534 569 538
rect 566 531 569 534
rect 582 539 585 545
rect 592 539 595 545
rect 613 540 616 545
rect 592 535 601 539
rect 613 536 614 540
rect 618 537 621 540
rect 638 539 641 545
rect 656 540 659 545
rect 695 546 698 568
rect 776 546 779 568
rect 866 546 869 568
rect 1380 561 1444 565
rect 1448 561 1503 565
rect 1507 561 1528 565
rect 1532 561 1559 565
rect 1563 561 1592 565
rect 1491 554 1492 558
rect 1516 553 1517 557
rect 1563 554 1564 558
rect 582 531 585 535
rect 592 531 595 535
rect 613 531 616 536
rect 640 535 641 539
rect 638 531 641 535
rect 656 531 659 536
rect 686 533 691 538
rect 695 534 696 537
rect 711 536 714 542
rect 711 533 719 536
rect 766 533 771 538
rect 775 534 777 537
rect 792 536 795 542
rect 792 533 800 536
rect 859 534 867 537
rect 882 536 885 542
rect 1439 540 1442 545
rect 1446 540 1449 545
rect 1429 537 1431 540
rect 882 533 890 536
rect 1439 537 1449 540
rect 711 530 714 533
rect 792 530 795 533
rect 882 530 885 533
rect 1439 531 1442 537
rect 566 516 569 520
rect 593 516 594 520
rect 638 516 640 520
rect 1446 531 1449 537
rect 1455 539 1458 545
rect 1471 540 1474 545
rect 1455 535 1457 539
rect 1461 535 1463 539
rect 1471 538 1477 540
rect 1481 538 1482 540
rect 1471 536 1482 538
rect 1499 538 1502 545
rect 1455 531 1458 535
rect 1471 531 1474 536
rect 1500 534 1502 538
rect 1499 531 1502 534
rect 1515 539 1518 545
rect 1525 539 1528 545
rect 1546 540 1549 545
rect 1525 535 1534 539
rect 1546 536 1547 540
rect 1551 537 1554 540
rect 1571 539 1574 545
rect 1589 540 1592 545
rect 1628 546 1631 568
rect 1709 546 1712 568
rect 1799 546 1802 568
rect 1515 531 1518 535
rect 1525 531 1528 535
rect 1546 531 1549 536
rect 1573 535 1574 539
rect 1571 531 1574 535
rect 1589 531 1592 536
rect 1619 533 1624 538
rect 1628 534 1629 537
rect 1644 536 1647 542
rect 1644 533 1652 536
rect 1699 533 1704 538
rect 1708 534 1710 537
rect 1725 536 1728 542
rect 1725 533 1733 536
rect 1792 534 1800 537
rect 1815 536 1818 542
rect 1815 533 1823 536
rect 1644 530 1647 533
rect 1725 530 1728 533
rect 1815 530 1818 533
rect 459 509 523 513
rect 527 509 554 513
rect 558 509 576 513
rect 580 509 641 513
rect 645 509 659 513
rect 695 506 698 522
rect 776 506 779 522
rect 866 506 869 522
rect 1499 516 1502 520
rect 1526 516 1527 520
rect 1571 516 1573 520
rect 1392 509 1456 513
rect 1460 509 1487 513
rect 1491 509 1509 513
rect 1513 509 1574 513
rect 1578 509 1592 513
rect 1628 506 1631 522
rect 1709 506 1712 522
rect 1799 506 1802 522
rect 423 502 496 506
rect 500 502 512 506
rect 516 502 530 506
rect 534 502 541 506
rect 545 502 547 506
rect 551 502 566 506
rect 570 502 603 506
rect 607 502 608 506
rect 612 502 620 506
rect 624 502 648 506
rect 652 502 664 506
rect 668 502 688 506
rect 692 502 742 506
rect 746 502 769 506
rect 773 502 859 506
rect 863 502 917 506
rect 1356 502 1429 506
rect 1433 502 1445 506
rect 1449 502 1463 506
rect 1467 502 1474 506
rect 1478 502 1480 506
rect 1484 502 1499 506
rect 1503 502 1536 506
rect 1540 502 1541 506
rect 1545 502 1553 506
rect 1557 502 1581 506
rect 1585 502 1597 506
rect 1601 502 1621 506
rect 1625 502 1675 506
rect 1679 502 1702 506
rect 1706 502 1792 506
rect 1796 502 1850 506
rect 459 495 523 499
rect 527 495 554 499
rect 558 495 576 499
rect 580 495 641 499
rect 645 495 659 499
rect 695 492 698 502
rect 725 498 728 502
rect 566 488 569 492
rect 593 488 594 492
rect 638 488 640 492
rect 495 468 498 471
rect 506 471 509 477
rect 513 471 516 477
rect 506 468 516 471
rect 506 463 509 468
rect 513 463 516 468
rect 522 473 525 477
rect 522 469 524 473
rect 528 469 530 473
rect 538 472 541 477
rect 566 474 569 477
rect 538 470 549 472
rect 522 463 525 469
rect 538 468 544 470
rect 538 463 541 468
rect 548 468 549 470
rect 567 470 569 474
rect 566 463 569 470
rect 1392 495 1456 499
rect 1460 495 1487 499
rect 1491 495 1509 499
rect 1513 495 1574 499
rect 1578 495 1592 499
rect 1628 492 1631 502
rect 1658 498 1661 502
rect 711 481 714 484
rect 582 473 585 477
rect 592 473 595 477
rect 592 469 601 473
rect 613 472 616 477
rect 638 473 641 477
rect 582 463 585 469
rect 592 463 595 469
rect 613 468 614 472
rect 618 468 621 471
rect 640 469 641 473
rect 656 472 659 477
rect 688 477 699 480
rect 711 478 719 481
rect 613 463 616 468
rect 638 463 641 469
rect 688 471 691 477
rect 711 472 714 478
rect 723 473 726 476
rect 734 476 737 490
rect 1499 488 1502 492
rect 1526 488 1527 492
rect 1571 488 1573 492
rect 742 476 747 481
rect 734 473 742 476
rect 656 463 659 468
rect 734 468 737 473
rect 1428 468 1431 471
rect 1439 471 1442 477
rect 1446 471 1449 477
rect 1439 468 1449 471
rect 686 462 691 467
rect 17 447 26 451
rect 30 447 62 451
rect 66 447 129 451
rect 133 447 158 451
rect 162 447 194 451
rect 198 447 261 451
rect 265 447 290 451
rect 294 447 326 451
rect 330 447 393 451
rect 397 447 477 451
rect 558 450 559 454
rect 583 451 584 455
rect 630 450 631 454
rect 17 440 50 444
rect 54 440 78 444
rect 82 440 108 444
rect 112 440 145 444
rect 149 440 182 444
rect 186 440 210 444
rect 214 440 240 444
rect 244 440 277 444
rect 281 440 314 444
rect 318 440 342 444
rect 346 440 372 444
rect 376 440 409 444
rect 413 440 417 444
rect 490 443 511 447
rect 515 443 520 447
rect 524 443 570 447
rect 574 443 595 447
rect 599 443 626 447
rect 630 443 659 447
rect 695 440 698 468
rect 725 440 728 464
rect 1439 463 1442 468
rect 1446 463 1449 468
rect 1455 473 1458 477
rect 1455 469 1457 473
rect 1461 469 1463 473
rect 1471 472 1474 477
rect 1499 474 1502 477
rect 1471 470 1482 472
rect 1455 463 1458 469
rect 1471 468 1477 470
rect 1471 463 1474 468
rect 1481 468 1482 470
rect 1500 470 1502 474
rect 1499 463 1502 470
rect 1644 481 1647 484
rect 1515 473 1518 477
rect 1525 473 1528 477
rect 1525 469 1534 473
rect 1546 472 1549 477
rect 1571 473 1574 477
rect 1515 463 1518 469
rect 1525 463 1528 469
rect 1546 468 1547 472
rect 1551 468 1554 471
rect 1573 469 1574 473
rect 1589 472 1592 477
rect 1621 477 1632 480
rect 1644 478 1652 481
rect 1546 463 1549 468
rect 1571 463 1574 469
rect 1621 471 1624 477
rect 1644 472 1647 478
rect 1656 473 1659 476
rect 1667 476 1670 490
rect 1675 476 1680 481
rect 1667 473 1675 476
rect 1589 463 1592 468
rect 1667 468 1670 473
rect 1619 462 1624 467
rect 950 447 959 451
rect 963 447 995 451
rect 999 447 1062 451
rect 1066 447 1091 451
rect 1095 447 1127 451
rect 1131 447 1194 451
rect 1198 447 1223 451
rect 1227 447 1259 451
rect 1263 447 1326 451
rect 1330 447 1410 451
rect 1491 450 1492 454
rect 1516 451 1517 455
rect 1563 450 1564 454
rect 950 440 983 444
rect 987 440 1011 444
rect 1015 440 1041 444
rect 1045 440 1078 444
rect 1082 440 1115 444
rect 1119 440 1143 444
rect 1147 440 1173 444
rect 1177 440 1210 444
rect 1214 440 1247 444
rect 1251 440 1275 444
rect 1279 440 1305 444
rect 1309 440 1342 444
rect 1346 440 1350 444
rect 1423 443 1444 447
rect 1448 443 1453 447
rect 1457 443 1503 447
rect 1507 443 1528 447
rect 1532 443 1559 447
rect 1563 443 1592 447
rect 1628 440 1631 468
rect 1658 440 1661 464
rect 20 430 23 440
rect 41 430 44 440
rect 57 430 60 440
rect 71 433 76 437
rect 80 433 87 437
rect 99 430 102 440
rect 115 430 118 440
rect 136 430 139 440
rect 152 430 155 440
rect 173 430 176 440
rect 189 430 192 440
rect 203 433 208 437
rect 212 433 219 437
rect 231 430 234 440
rect 247 430 250 440
rect 268 430 271 440
rect 284 430 287 440
rect 305 430 308 440
rect 321 430 324 440
rect 335 433 340 437
rect 344 433 351 437
rect 363 430 366 440
rect 379 430 382 440
rect 400 430 403 440
rect 435 436 497 440
rect 501 436 503 440
rect 507 436 511 440
rect 515 436 529 440
rect 533 436 538 440
rect 542 436 547 440
rect 551 436 570 440
rect 574 436 604 440
rect 608 436 619 440
rect 623 436 647 440
rect 651 436 664 440
rect 668 436 688 440
rect 692 436 772 440
rect 776 436 790 440
rect 794 436 799 440
rect 803 436 808 440
rect 812 436 831 440
rect 835 436 865 440
rect 869 436 880 440
rect 884 436 908 440
rect 912 436 921 440
rect 37 416 42 419
rect 46 416 70 419
rect 95 416 102 419
rect 106 416 128 419
rect 148 416 155 419
rect 169 416 174 419
rect 178 416 202 419
rect 227 416 234 419
rect 238 416 260 419
rect 280 416 287 419
rect 301 416 306 419
rect 310 416 334 419
rect 447 429 511 433
rect 515 429 520 433
rect 524 429 570 433
rect 574 429 595 433
rect 599 429 626 433
rect 630 429 659 433
rect 359 416 366 419
rect 370 416 392 419
rect 558 422 559 426
rect 583 421 584 425
rect 630 422 631 426
rect 53 406 60 409
rect 64 410 83 413
rect 83 403 86 409
rect 111 406 118 409
rect 122 410 137 413
rect 185 406 192 409
rect 196 410 215 413
rect 215 403 218 409
rect 243 406 250 409
rect 254 410 269 413
rect 317 406 324 409
rect 328 410 347 413
rect 347 403 350 409
rect 375 406 382 409
rect 386 410 403 413
rect 506 408 509 413
rect 513 408 516 413
rect 496 405 498 408
rect 506 405 516 408
rect 506 399 509 405
rect 20 387 23 399
rect 41 387 44 399
rect 57 387 60 399
rect 71 390 83 393
rect 99 387 102 399
rect 115 387 118 399
rect 136 387 139 399
rect 152 387 155 399
rect 173 387 176 399
rect 189 387 192 399
rect 203 390 215 393
rect 231 387 234 399
rect 247 387 250 399
rect 268 387 271 399
rect 284 387 287 399
rect 305 387 308 399
rect 321 387 324 399
rect 335 390 347 393
rect 363 387 366 399
rect 379 387 382 399
rect 400 387 403 399
rect 513 399 516 405
rect 522 407 525 413
rect 538 408 541 413
rect 522 403 524 407
rect 528 403 530 407
rect 538 406 544 408
rect 548 406 549 408
rect 538 404 549 406
rect 566 406 569 413
rect 522 399 525 403
rect 538 399 541 404
rect 567 402 569 406
rect 566 399 569 402
rect 582 407 585 413
rect 592 407 595 413
rect 613 408 616 413
rect 592 403 601 407
rect 613 404 614 408
rect 618 405 621 408
rect 638 407 641 413
rect 656 408 659 413
rect 695 410 698 436
rect 731 429 750 433
rect 754 429 772 433
rect 776 429 831 433
rect 835 429 856 433
rect 860 429 887 433
rect 891 429 920 433
rect 953 430 956 440
rect 974 430 977 440
rect 990 430 993 440
rect 1004 433 1009 437
rect 1013 433 1020 437
rect 1032 430 1035 440
rect 1048 430 1051 440
rect 1069 430 1072 440
rect 1085 430 1088 440
rect 1106 430 1109 440
rect 1122 430 1125 440
rect 1136 433 1141 437
rect 1145 433 1152 437
rect 1164 430 1167 440
rect 1180 430 1183 440
rect 1201 430 1204 440
rect 1217 430 1220 440
rect 1238 430 1241 440
rect 1254 430 1257 440
rect 1268 433 1273 437
rect 1277 433 1284 437
rect 1296 430 1299 440
rect 1312 430 1315 440
rect 1333 430 1336 440
rect 1368 436 1430 440
rect 1434 436 1436 440
rect 1440 436 1444 440
rect 1448 436 1462 440
rect 1466 436 1471 440
rect 1475 436 1480 440
rect 1484 436 1503 440
rect 1507 436 1537 440
rect 1541 436 1552 440
rect 1556 436 1580 440
rect 1584 436 1597 440
rect 1601 436 1621 440
rect 1625 436 1705 440
rect 1709 436 1723 440
rect 1727 436 1732 440
rect 1736 436 1741 440
rect 1745 436 1764 440
rect 1768 436 1798 440
rect 1802 436 1813 440
rect 1817 436 1841 440
rect 1845 436 1854 440
rect 731 417 734 429
rect 819 422 820 426
rect 844 421 845 425
rect 891 422 892 426
rect 582 399 585 403
rect 592 399 595 403
rect 613 399 616 404
rect 640 403 641 407
rect 758 408 761 413
rect 767 408 770 413
rect 774 408 777 413
rect 638 399 641 403
rect 656 399 659 404
rect 685 397 690 402
rect 694 398 696 401
rect 711 400 714 406
rect 743 405 777 408
rect 711 397 719 400
rect 711 394 714 397
rect 17 383 50 387
rect 54 383 78 387
rect 82 383 108 387
rect 112 383 182 387
rect 186 383 210 387
rect 214 383 240 387
rect 244 383 314 387
rect 318 383 342 387
rect 346 383 372 387
rect 376 383 429 387
rect 566 384 569 388
rect 593 384 594 388
rect 638 384 640 388
rect 743 391 746 405
rect 767 399 770 405
rect 774 399 777 405
rect 783 407 786 413
rect 799 408 802 413
rect 783 403 785 407
rect 789 403 791 407
rect 799 406 805 408
rect 809 406 810 408
rect 799 404 810 406
rect 827 406 830 413
rect 783 399 786 403
rect 799 399 802 404
rect 828 402 830 406
rect 827 399 830 402
rect 970 416 975 419
rect 979 416 1003 419
rect 1028 416 1035 419
rect 1039 416 1061 419
rect 1081 416 1088 419
rect 1102 416 1107 419
rect 1111 416 1135 419
rect 1160 416 1167 419
rect 1171 416 1193 419
rect 1213 416 1220 419
rect 1234 416 1239 419
rect 1243 416 1267 419
rect 1380 429 1444 433
rect 1448 429 1453 433
rect 1457 429 1503 433
rect 1507 429 1528 433
rect 1532 429 1559 433
rect 1563 429 1592 433
rect 1292 416 1299 419
rect 1303 416 1325 419
rect 1491 422 1492 426
rect 1516 421 1517 425
rect 1563 422 1564 426
rect 843 407 846 413
rect 853 407 856 413
rect 874 408 877 413
rect 853 403 862 407
rect 874 404 875 408
rect 879 405 882 408
rect 899 407 902 413
rect 917 408 920 413
rect 843 399 846 403
rect 853 399 856 403
rect 874 399 877 404
rect 901 403 902 407
rect 899 399 902 403
rect 917 399 920 404
rect 986 406 993 409
rect 997 410 1016 413
rect 1016 403 1019 409
rect 1044 406 1051 409
rect 1055 410 1070 413
rect 1118 406 1125 409
rect 1129 410 1148 413
rect 1148 403 1151 409
rect 1176 406 1183 409
rect 1187 410 1202 413
rect 1250 406 1257 409
rect 1261 410 1280 413
rect 1280 403 1283 409
rect 1308 406 1315 409
rect 1319 410 1336 413
rect 1439 408 1442 413
rect 1446 408 1449 413
rect 1429 405 1431 408
rect 1439 405 1449 408
rect 1439 399 1442 405
rect 17 376 26 380
rect 30 376 77 380
rect 81 376 127 380
rect 131 376 158 380
rect 162 376 209 380
rect 213 376 259 380
rect 263 376 290 380
rect 294 376 341 380
rect 345 376 391 380
rect 395 377 465 380
rect 509 377 523 381
rect 527 377 554 381
rect 558 377 576 381
rect 580 377 641 381
rect 645 377 659 381
rect 695 374 698 386
rect 827 384 830 388
rect 854 384 855 388
rect 899 384 901 388
rect 953 387 956 399
rect 974 387 977 399
rect 990 387 993 399
rect 1004 390 1016 393
rect 1032 387 1035 399
rect 1048 387 1051 399
rect 1069 387 1072 399
rect 1085 387 1088 399
rect 1106 387 1109 399
rect 1122 387 1125 399
rect 1136 390 1148 393
rect 1164 387 1167 399
rect 1180 387 1183 399
rect 1201 387 1204 399
rect 1217 387 1220 399
rect 1238 387 1241 399
rect 1254 387 1257 399
rect 1268 390 1280 393
rect 1296 387 1299 399
rect 1312 387 1315 399
rect 1333 387 1336 399
rect 1446 399 1449 405
rect 1455 407 1458 413
rect 1471 408 1474 413
rect 1455 403 1457 407
rect 1461 403 1463 407
rect 1471 406 1477 408
rect 1481 406 1482 408
rect 1471 404 1482 406
rect 1499 406 1502 413
rect 1455 399 1458 403
rect 1471 399 1474 404
rect 1500 402 1502 406
rect 1499 399 1502 402
rect 1515 407 1518 413
rect 1525 407 1528 413
rect 1546 408 1549 413
rect 1525 403 1534 407
rect 1546 404 1547 408
rect 1551 405 1554 408
rect 1571 407 1574 413
rect 1589 408 1592 413
rect 1628 410 1631 436
rect 1664 429 1683 433
rect 1687 429 1705 433
rect 1709 429 1764 433
rect 1768 429 1789 433
rect 1793 429 1820 433
rect 1824 429 1853 433
rect 1664 417 1667 429
rect 1752 422 1753 426
rect 1777 421 1778 425
rect 1824 422 1825 426
rect 1515 399 1518 403
rect 1525 399 1528 403
rect 1546 399 1549 404
rect 1573 403 1574 407
rect 1691 408 1694 413
rect 1700 408 1703 413
rect 1707 408 1710 413
rect 1571 399 1574 403
rect 1589 399 1592 404
rect 1618 397 1623 402
rect 1627 398 1629 401
rect 1644 400 1647 406
rect 1676 405 1710 408
rect 1644 397 1652 400
rect 1644 394 1647 397
rect 950 383 983 387
rect 987 383 1011 387
rect 1015 383 1041 387
rect 1045 383 1115 387
rect 1119 383 1143 387
rect 1147 383 1173 387
rect 1177 383 1247 387
rect 1251 383 1275 387
rect 1279 383 1305 387
rect 1309 383 1362 387
rect 1499 384 1502 388
rect 1526 384 1527 388
rect 1571 384 1573 388
rect 1676 391 1679 405
rect 1700 399 1703 405
rect 1707 399 1710 405
rect 1716 407 1719 413
rect 1732 408 1735 413
rect 1716 403 1718 407
rect 1722 403 1724 407
rect 1732 406 1738 408
rect 1742 406 1743 408
rect 1732 404 1743 406
rect 1760 406 1763 413
rect 1716 399 1719 403
rect 1732 399 1735 404
rect 1761 402 1763 406
rect 1760 399 1763 402
rect 1776 407 1779 413
rect 1786 407 1789 413
rect 1807 408 1810 413
rect 1786 403 1795 407
rect 1807 404 1808 408
rect 1812 405 1815 408
rect 1832 407 1835 413
rect 1850 408 1853 413
rect 1776 399 1779 403
rect 1786 399 1789 403
rect 1807 399 1810 404
rect 1834 403 1835 407
rect 1832 399 1835 403
rect 1850 399 1853 404
rect 735 377 740 381
rect 744 377 784 381
rect 788 377 815 381
rect 819 377 837 381
rect 841 377 902 381
rect 906 377 920 381
rect 950 376 959 380
rect 963 376 1010 380
rect 1014 376 1060 380
rect 1064 376 1091 380
rect 1095 376 1142 380
rect 1146 376 1192 380
rect 1196 376 1223 380
rect 1227 376 1274 380
rect 1278 376 1324 380
rect 1328 377 1398 380
rect 1442 377 1456 381
rect 1460 377 1487 381
rect 1491 377 1509 381
rect 1513 377 1574 381
rect 1578 377 1592 381
rect 1628 374 1631 386
rect 1760 384 1763 388
rect 1787 384 1788 388
rect 1832 384 1834 388
rect 1668 377 1673 381
rect 1677 377 1717 381
rect 1721 377 1748 381
rect 1752 377 1770 381
rect 1774 377 1835 381
rect 1839 377 1853 381
rect 24 370 408 373
rect 423 370 496 374
rect 500 370 512 374
rect 516 370 530 374
rect 534 370 541 374
rect 545 370 547 374
rect 551 370 566 374
rect 570 370 603 374
rect 607 370 608 374
rect 612 370 620 374
rect 624 370 648 374
rect 652 370 688 374
rect 692 370 731 374
rect 735 370 742 374
rect 746 370 757 374
rect 761 370 773 374
rect 777 370 791 374
rect 795 370 802 374
rect 806 370 808 374
rect 812 370 827 374
rect 831 370 864 374
rect 868 370 869 374
rect 873 370 881 374
rect 885 370 909 374
rect 913 370 921 374
rect 957 370 1341 373
rect 1356 370 1429 374
rect 1433 370 1445 374
rect 1449 370 1463 374
rect 1467 370 1474 374
rect 1478 370 1480 374
rect 1484 370 1499 374
rect 1503 370 1536 374
rect 1540 370 1541 374
rect 1545 370 1553 374
rect 1557 370 1581 374
rect 1585 370 1621 374
rect 1625 370 1664 374
rect 1668 370 1675 374
rect 1679 370 1690 374
rect 1694 370 1706 374
rect 1710 370 1724 374
rect 1728 370 1735 374
rect 1739 370 1741 374
rect 1745 370 1760 374
rect 1764 370 1797 374
rect 1801 370 1802 374
rect 1806 370 1814 374
rect 1818 370 1842 374
rect 1846 370 1854 374
rect 167 363 276 366
rect 459 363 505 367
rect 509 363 739 366
rect 929 364 937 368
rect 1100 363 1209 366
rect 1392 363 1438 367
rect 1442 363 1672 366
rect 1862 364 1870 368
rect 147 355 151 359
rect 155 355 159 359
rect 447 356 749 359
rect 925 348 929 352
rect 1080 355 1084 359
rect 1088 355 1092 359
rect 1380 356 1682 359
rect 1858 348 1862 352
rect 3 344 135 348
rect 139 344 155 348
rect 171 344 1068 348
rect 1072 344 1088 348
rect 1104 344 1950 348
rect 163 337 408 340
rect 483 337 797 341
rect 801 337 833 341
rect 837 337 900 341
rect 904 337 920 341
rect 1096 337 1341 340
rect 1416 337 1730 341
rect 1734 337 1766 341
rect 1770 337 1833 341
rect 1837 337 1853 341
rect 178 330 408 333
rect 423 330 783 334
rect 787 330 821 334
rect 825 330 849 334
rect 853 330 879 334
rect 883 330 916 334
rect 147 321 151 325
rect 155 321 159 325
rect 791 320 794 330
rect 812 320 815 330
rect 828 320 831 330
rect 842 323 847 327
rect 851 323 858 327
rect 870 320 873 330
rect 886 320 889 330
rect 907 320 910 330
rect 1111 330 1341 333
rect 1356 330 1716 334
rect 1720 330 1754 334
rect 1758 330 1782 334
rect 1786 330 1812 334
rect 1816 330 1849 334
rect 1080 321 1084 325
rect 1088 321 1092 325
rect 1724 320 1727 330
rect 1745 320 1748 330
rect 1761 320 1764 330
rect 1775 323 1780 327
rect 1784 323 1791 327
rect 1803 320 1806 330
rect 1819 320 1822 330
rect 1840 320 1843 330
rect 167 314 277 317
rect 17 307 26 311
rect 30 307 62 311
rect 66 307 129 311
rect 133 307 158 311
rect 162 307 194 311
rect 198 307 261 311
rect 265 307 290 311
rect 294 307 326 311
rect 330 307 393 311
rect 397 307 477 311
rect 17 300 50 304
rect 54 300 78 304
rect 82 300 108 304
rect 112 300 145 304
rect 149 300 182 304
rect 186 300 210 304
rect 214 300 240 304
rect 244 300 277 304
rect 281 300 314 304
rect 318 300 342 304
rect 346 300 372 304
rect 376 300 409 304
rect 413 300 417 304
rect 808 306 813 309
rect 817 306 841 309
rect 1100 314 1210 317
rect 866 306 873 309
rect 877 306 899 309
rect 950 307 959 311
rect 963 307 995 311
rect 999 307 1062 311
rect 1066 307 1091 311
rect 1095 307 1127 311
rect 1131 307 1194 311
rect 1198 307 1223 311
rect 1227 307 1259 311
rect 1263 307 1326 311
rect 1330 307 1410 311
rect 20 290 23 300
rect 41 290 44 300
rect 57 290 60 300
rect 71 293 76 297
rect 80 293 87 297
rect 99 290 102 300
rect 115 290 118 300
rect 136 290 139 300
rect 152 290 155 300
rect 173 290 176 300
rect 189 290 192 300
rect 203 293 208 297
rect 212 293 219 297
rect 231 290 234 300
rect 247 290 250 300
rect 268 290 271 300
rect 284 290 287 300
rect 305 290 308 300
rect 321 290 324 300
rect 335 293 340 297
rect 344 293 351 297
rect 363 290 366 300
rect 379 290 382 300
rect 400 290 403 300
rect 824 296 831 299
rect 835 300 854 303
rect 37 276 42 279
rect 46 276 70 279
rect 95 276 102 279
rect 106 276 128 279
rect 148 276 155 279
rect 169 276 174 279
rect 178 276 202 279
rect 227 276 234 279
rect 238 276 260 279
rect 280 276 287 279
rect 301 276 306 279
rect 310 276 334 279
rect 359 276 366 279
rect 370 276 392 279
rect 854 293 857 299
rect 882 296 889 299
rect 893 300 908 303
rect 950 300 983 304
rect 987 300 1011 304
rect 1015 300 1041 304
rect 1045 300 1078 304
rect 1082 300 1115 304
rect 1119 300 1143 304
rect 1147 300 1173 304
rect 1177 300 1210 304
rect 1214 300 1247 304
rect 1251 300 1275 304
rect 1279 300 1305 304
rect 1309 300 1342 304
rect 1346 300 1350 304
rect 1741 306 1746 309
rect 1750 306 1774 309
rect 1799 306 1806 309
rect 1810 306 1832 309
rect 953 290 956 300
rect 974 290 977 300
rect 990 290 993 300
rect 1004 293 1009 297
rect 1013 293 1020 297
rect 1032 290 1035 300
rect 1048 290 1051 300
rect 1069 290 1072 300
rect 1085 290 1088 300
rect 1106 290 1109 300
rect 1122 290 1125 300
rect 1136 293 1141 297
rect 1145 293 1152 297
rect 1164 290 1167 300
rect 1180 290 1183 300
rect 1201 290 1204 300
rect 1217 290 1220 300
rect 1238 290 1241 300
rect 1254 290 1257 300
rect 1268 293 1273 297
rect 1277 293 1284 297
rect 1296 290 1299 300
rect 1312 290 1315 300
rect 1333 290 1336 300
rect 1757 296 1764 299
rect 1768 300 1787 303
rect 791 277 794 289
rect 812 277 815 289
rect 828 277 831 289
rect 842 280 854 283
rect 870 277 873 289
rect 886 277 889 289
rect 907 277 910 289
rect 53 266 60 269
rect 64 270 83 273
rect 83 263 86 269
rect 111 266 118 269
rect 122 270 137 273
rect 185 266 192 269
rect 196 270 215 273
rect 215 263 218 269
rect 243 266 250 269
rect 254 270 269 273
rect 317 266 324 269
rect 328 270 347 273
rect 347 263 350 269
rect 375 266 382 269
rect 386 270 403 273
rect 435 273 821 277
rect 825 273 849 277
rect 853 273 879 277
rect 883 273 920 277
rect 970 276 975 279
rect 979 276 1003 279
rect 1028 276 1035 279
rect 1039 276 1061 279
rect 1081 276 1088 279
rect 1102 276 1107 279
rect 1111 276 1135 279
rect 1160 276 1167 279
rect 1171 276 1193 279
rect 1213 276 1220 279
rect 1234 276 1239 279
rect 1243 276 1267 279
rect 1292 276 1299 279
rect 1303 276 1325 279
rect 1787 293 1790 299
rect 1815 296 1822 299
rect 1826 300 1841 303
rect 1724 277 1727 289
rect 1745 277 1748 289
rect 1761 277 1764 289
rect 1775 280 1787 283
rect 1803 277 1806 289
rect 1819 277 1822 289
rect 1840 277 1843 289
rect 471 266 797 270
rect 801 266 848 270
rect 852 266 898 270
rect 902 266 920 270
rect 986 266 993 269
rect 997 270 1016 273
rect 20 247 23 259
rect 41 247 44 259
rect 57 247 60 259
rect 71 250 83 253
rect 99 247 102 259
rect 115 247 118 259
rect 136 247 139 259
rect 152 247 155 259
rect 173 247 176 259
rect 189 247 192 259
rect 203 250 215 253
rect 231 247 234 259
rect 247 247 250 259
rect 268 247 271 259
rect 284 247 287 259
rect 305 247 308 259
rect 321 247 324 259
rect 335 250 347 253
rect 363 247 366 259
rect 379 247 382 259
rect 400 247 403 259
rect 794 259 915 262
rect 1016 263 1019 269
rect 1044 266 1051 269
rect 1055 270 1070 273
rect 1118 266 1125 269
rect 1129 270 1148 273
rect 1148 263 1151 269
rect 1176 266 1183 269
rect 1187 270 1202 273
rect 1250 266 1257 269
rect 1261 270 1280 273
rect 1280 263 1283 269
rect 1308 266 1315 269
rect 1319 270 1336 273
rect 1368 273 1754 277
rect 1758 273 1782 277
rect 1786 273 1812 277
rect 1816 273 1853 277
rect 1404 266 1730 270
rect 1734 266 1781 270
rect 1785 266 1831 270
rect 1835 266 1853 270
rect 483 251 797 255
rect 801 251 833 255
rect 837 251 900 255
rect 904 251 920 255
rect 17 243 50 247
rect 54 243 78 247
rect 82 243 108 247
rect 112 243 182 247
rect 186 243 210 247
rect 214 243 240 247
rect 244 243 314 247
rect 318 243 342 247
rect 346 243 372 247
rect 376 243 429 247
rect 787 244 821 248
rect 825 244 849 248
rect 853 244 879 248
rect 883 244 916 248
rect 953 247 956 259
rect 974 247 977 259
rect 990 247 993 259
rect 1004 250 1016 253
rect 1032 247 1035 259
rect 1048 247 1051 259
rect 1069 247 1072 259
rect 1085 247 1088 259
rect 1106 247 1109 259
rect 1122 247 1125 259
rect 1136 250 1148 253
rect 1164 247 1167 259
rect 1180 247 1183 259
rect 1201 247 1204 259
rect 1217 247 1220 259
rect 1238 247 1241 259
rect 1254 247 1257 259
rect 1268 250 1280 253
rect 1296 247 1299 259
rect 1312 247 1315 259
rect 1333 247 1336 259
rect 1727 259 1848 262
rect 1416 251 1730 255
rect 1734 251 1766 255
rect 1770 251 1833 255
rect 1837 251 1853 255
rect 17 236 26 240
rect 30 236 77 240
rect 81 236 127 240
rect 131 236 158 240
rect 162 236 209 240
rect 213 236 259 240
rect 263 236 290 240
rect 294 236 341 240
rect 345 236 391 240
rect 395 236 465 240
rect 791 234 794 244
rect 812 234 815 244
rect 828 234 831 244
rect 842 237 847 241
rect 851 237 858 241
rect 870 234 873 244
rect 886 234 889 244
rect 907 234 910 244
rect 950 243 983 247
rect 987 243 1011 247
rect 1015 243 1041 247
rect 1045 243 1115 247
rect 1119 243 1143 247
rect 1147 243 1173 247
rect 1177 243 1247 247
rect 1251 243 1275 247
rect 1279 243 1305 247
rect 1309 243 1362 247
rect 1720 244 1754 248
rect 1758 244 1782 248
rect 1786 244 1812 248
rect 1816 244 1849 248
rect 950 236 959 240
rect 963 236 1010 240
rect 1014 236 1060 240
rect 1064 236 1091 240
rect 1095 236 1142 240
rect 1146 236 1192 240
rect 1196 236 1223 240
rect 1227 236 1274 240
rect 1278 236 1324 240
rect 1328 236 1398 240
rect 1724 234 1727 244
rect 1745 234 1748 244
rect 1761 234 1764 244
rect 1775 237 1780 241
rect 1784 237 1791 241
rect 1803 234 1806 244
rect 1819 234 1822 244
rect 1840 234 1843 244
rect 23 229 408 232
rect 17 221 26 225
rect 30 221 62 225
rect 66 221 129 225
rect 133 221 158 225
rect 162 221 194 225
rect 198 221 261 225
rect 265 221 290 225
rect 294 221 326 225
rect 330 221 393 225
rect 397 221 477 225
rect 17 214 50 218
rect 54 214 78 218
rect 82 214 108 218
rect 112 214 145 218
rect 149 214 182 218
rect 186 214 210 218
rect 214 214 240 218
rect 244 214 277 218
rect 281 214 314 218
rect 318 214 342 218
rect 346 214 372 218
rect 376 214 409 218
rect 413 214 417 218
rect 808 220 813 223
rect 817 220 841 223
rect 956 229 1341 232
rect 866 220 873 223
rect 877 220 899 223
rect 950 221 959 225
rect 963 221 995 225
rect 999 221 1062 225
rect 1066 221 1091 225
rect 1095 221 1127 225
rect 1131 221 1194 225
rect 1198 221 1223 225
rect 1227 221 1259 225
rect 1263 221 1326 225
rect 1330 221 1410 225
rect 20 204 23 214
rect 41 204 44 214
rect 57 204 60 214
rect 71 207 76 211
rect 80 207 87 211
rect 99 204 102 214
rect 115 204 118 214
rect 136 204 139 214
rect 152 204 155 214
rect 173 204 176 214
rect 189 204 192 214
rect 203 207 208 211
rect 212 207 219 211
rect 231 204 234 214
rect 247 204 250 214
rect 268 204 271 214
rect 284 204 287 214
rect 305 204 308 214
rect 321 204 324 214
rect 335 207 340 211
rect 344 207 351 211
rect 363 204 366 214
rect 379 204 382 214
rect 400 204 403 214
rect 824 210 831 213
rect 835 214 854 217
rect 37 190 42 193
rect 46 190 70 193
rect 95 190 102 193
rect 106 190 128 193
rect 148 190 155 193
rect 169 190 174 193
rect 178 190 202 193
rect 227 190 234 193
rect 238 190 260 193
rect 280 190 287 193
rect 301 190 306 193
rect 310 190 334 193
rect 359 190 366 193
rect 370 190 392 193
rect 854 207 857 213
rect 882 210 889 213
rect 893 214 908 217
rect 919 212 930 216
rect 950 214 983 218
rect 987 214 1011 218
rect 1015 214 1041 218
rect 1045 214 1078 218
rect 1082 214 1115 218
rect 1119 214 1143 218
rect 1147 214 1173 218
rect 1177 214 1210 218
rect 1214 214 1247 218
rect 1251 214 1275 218
rect 1279 214 1305 218
rect 1309 214 1342 218
rect 1346 214 1350 218
rect 1741 220 1746 223
rect 1750 220 1774 223
rect 1799 220 1806 223
rect 1810 220 1832 223
rect 953 204 956 214
rect 974 204 977 214
rect 990 204 993 214
rect 1004 207 1009 211
rect 1013 207 1020 211
rect 1032 204 1035 214
rect 1048 204 1051 214
rect 1069 204 1072 214
rect 1085 204 1088 214
rect 1106 204 1109 214
rect 1122 204 1125 214
rect 1136 207 1141 211
rect 1145 207 1152 211
rect 1164 204 1167 214
rect 1180 204 1183 214
rect 1201 204 1204 214
rect 1217 204 1220 214
rect 1238 204 1241 214
rect 1254 204 1257 214
rect 1268 207 1273 211
rect 1277 207 1284 211
rect 1296 204 1299 214
rect 1312 204 1315 214
rect 1333 204 1336 214
rect 1757 210 1764 213
rect 1768 214 1787 217
rect 791 191 794 203
rect 812 191 815 203
rect 828 191 831 203
rect 842 194 854 197
rect 870 191 873 203
rect 886 191 889 203
rect 907 191 910 203
rect 53 180 60 183
rect 64 184 83 187
rect 83 177 86 183
rect 111 180 118 183
rect 122 184 137 187
rect 185 180 192 183
rect 196 184 215 187
rect 215 177 218 183
rect 243 180 250 183
rect 254 184 269 187
rect 317 180 324 183
rect 328 184 347 187
rect 347 177 350 183
rect 375 180 382 183
rect 386 184 403 187
rect 435 187 821 191
rect 825 187 849 191
rect 853 187 879 191
rect 883 187 920 191
rect 970 190 975 193
rect 979 190 1003 193
rect 1028 190 1035 193
rect 1039 190 1061 193
rect 1081 190 1088 193
rect 1102 190 1107 193
rect 1111 190 1135 193
rect 1160 190 1167 193
rect 1171 190 1193 193
rect 1213 190 1220 193
rect 1234 190 1239 193
rect 1243 190 1267 193
rect 1292 190 1299 193
rect 1303 190 1325 193
rect 1787 207 1790 213
rect 1815 210 1822 213
rect 1826 214 1841 217
rect 1852 212 1863 216
rect 1724 191 1727 203
rect 1745 191 1748 203
rect 1761 191 1764 203
rect 1775 194 1787 197
rect 1803 191 1806 203
rect 1819 191 1822 203
rect 1840 191 1843 203
rect 471 180 797 184
rect 801 180 848 184
rect 852 180 898 184
rect 902 180 920 184
rect 986 180 993 183
rect 997 184 1016 187
rect 1016 177 1019 183
rect 1044 180 1051 183
rect 1055 184 1070 187
rect 1118 180 1125 183
rect 1129 184 1148 187
rect 1148 177 1151 183
rect 1176 180 1183 183
rect 1187 184 1202 187
rect 1250 180 1257 183
rect 1261 184 1280 187
rect 1280 177 1283 183
rect 1308 180 1315 183
rect 1319 184 1336 187
rect 1368 187 1754 191
rect 1758 187 1782 191
rect 1786 187 1812 191
rect 1816 187 1853 191
rect 1404 180 1730 184
rect 1734 180 1781 184
rect 1785 180 1831 184
rect 1835 180 1853 184
rect 20 161 23 173
rect 41 161 44 173
rect 57 161 60 173
rect 71 164 83 167
rect 99 161 102 173
rect 115 161 118 173
rect 136 161 139 173
rect 152 161 155 173
rect 173 161 176 173
rect 189 161 192 173
rect 203 164 215 167
rect 231 161 234 173
rect 247 161 250 173
rect 268 161 271 173
rect 284 161 287 173
rect 305 161 308 173
rect 321 161 324 173
rect 335 164 347 167
rect 363 161 366 173
rect 379 161 382 173
rect 400 161 403 173
rect 953 161 956 173
rect 974 161 977 173
rect 990 161 993 173
rect 1004 164 1016 167
rect 1032 161 1035 173
rect 1048 161 1051 173
rect 1069 161 1072 173
rect 1085 161 1088 173
rect 1106 161 1109 173
rect 1122 161 1125 173
rect 1136 164 1148 167
rect 1164 161 1167 173
rect 1180 161 1183 173
rect 1201 161 1204 173
rect 1217 161 1220 173
rect 1238 161 1241 173
rect 1254 161 1257 173
rect 1268 164 1280 167
rect 1296 161 1299 173
rect 1312 161 1315 173
rect 1333 161 1336 173
rect 17 157 50 161
rect 54 157 78 161
rect 82 157 108 161
rect 112 157 182 161
rect 186 157 210 161
rect 214 157 240 161
rect 244 157 314 161
rect 318 157 342 161
rect 346 157 372 161
rect 376 157 429 161
rect 950 157 983 161
rect 987 157 1011 161
rect 1015 157 1041 161
rect 1045 157 1115 161
rect 1119 157 1143 161
rect 1147 157 1173 161
rect 1177 157 1247 161
rect 1251 157 1275 161
rect 1279 157 1305 161
rect 1309 157 1362 161
rect 17 150 26 154
rect 30 150 77 154
rect 81 150 127 154
rect 131 150 158 154
rect 162 150 209 154
rect 213 150 259 154
rect 263 150 290 154
rect 294 150 341 154
rect 345 150 391 154
rect 395 150 465 154
rect 950 150 959 154
rect 963 150 1010 154
rect 1014 150 1060 154
rect 1064 150 1091 154
rect 1095 150 1142 154
rect 1146 150 1192 154
rect 1196 150 1223 154
rect 1227 150 1274 154
rect 1278 150 1324 154
rect 1328 150 1398 154
rect 23 144 408 147
rect 956 144 1341 147
rect 148 137 252 140
rect 1081 137 1185 140
rect 264 129 268 133
rect 272 129 276 133
rect 1197 129 1201 133
rect 1205 129 1209 133
rect 0 118 252 122
rect 256 118 272 122
rect 288 118 937 122
rect 941 118 1185 122
rect 1189 118 1205 122
rect 1221 118 1870 122
rect 1874 118 1957 122
rect 280 111 408 114
rect 1213 111 1341 114
rect 295 104 408 107
rect 1228 104 1341 107
rect 264 95 268 99
rect 272 95 276 99
rect 1197 95 1201 99
rect 1205 95 1209 99
rect 148 88 252 91
rect 1081 88 1185 91
rect 17 81 26 85
rect 30 81 62 85
rect 66 81 129 85
rect 133 81 158 85
rect 162 81 194 85
rect 198 81 261 85
rect 265 81 290 85
rect 294 81 326 85
rect 330 81 393 85
rect 397 81 477 85
rect 950 81 959 85
rect 963 81 995 85
rect 999 81 1062 85
rect 1066 81 1091 85
rect 1095 81 1127 85
rect 1131 81 1194 85
rect 1198 81 1223 85
rect 1227 81 1259 85
rect 1263 81 1326 85
rect 1330 81 1410 85
rect 17 74 50 78
rect 54 74 78 78
rect 82 74 108 78
rect 112 74 145 78
rect 149 74 182 78
rect 186 74 210 78
rect 214 74 240 78
rect 244 74 277 78
rect 281 74 314 78
rect 318 74 342 78
rect 346 74 372 78
rect 376 74 409 78
rect 413 74 417 78
rect 950 74 983 78
rect 987 74 1011 78
rect 1015 74 1041 78
rect 1045 74 1078 78
rect 1082 74 1115 78
rect 1119 74 1143 78
rect 1147 74 1173 78
rect 1177 74 1210 78
rect 1214 74 1247 78
rect 1251 74 1275 78
rect 1279 74 1305 78
rect 1309 74 1342 78
rect 1346 74 1350 78
rect 20 64 23 74
rect 41 64 44 74
rect 57 64 60 74
rect 71 67 76 71
rect 80 67 87 71
rect 99 64 102 74
rect 115 64 118 74
rect 136 64 139 74
rect 152 64 155 74
rect 173 64 176 74
rect 189 64 192 74
rect 203 67 208 71
rect 212 67 219 71
rect 231 64 234 74
rect 247 64 250 74
rect 268 64 271 74
rect 284 64 287 74
rect 305 64 308 74
rect 321 64 324 74
rect 335 67 340 71
rect 344 67 351 71
rect 363 64 366 74
rect 379 64 382 74
rect 400 64 403 74
rect 953 64 956 74
rect 974 64 977 74
rect 990 64 993 74
rect 1004 67 1009 71
rect 1013 67 1020 71
rect 1032 64 1035 74
rect 1048 64 1051 74
rect 1069 64 1072 74
rect 1085 64 1088 74
rect 1106 64 1109 74
rect 1122 64 1125 74
rect 1136 67 1141 71
rect 1145 67 1152 71
rect 1164 64 1167 74
rect 1180 64 1183 74
rect 1201 64 1204 74
rect 1217 64 1220 74
rect 1238 64 1241 74
rect 1254 64 1257 74
rect 1268 67 1273 71
rect 1277 67 1284 71
rect 1296 64 1299 74
rect 1312 64 1315 74
rect 1333 64 1336 74
rect 37 50 42 53
rect 46 50 70 53
rect 95 50 102 53
rect 106 50 128 53
rect 148 50 155 53
rect 169 50 174 53
rect 178 50 202 53
rect 227 50 234 53
rect 238 50 260 53
rect 280 50 287 53
rect 301 50 306 53
rect 310 50 334 53
rect 359 50 366 53
rect 370 50 392 53
rect 53 40 60 43
rect 64 44 83 47
rect 83 37 86 43
rect 111 40 118 43
rect 122 44 137 47
rect 185 40 192 43
rect 196 44 215 47
rect 215 37 218 43
rect 243 40 250 43
rect 254 44 269 47
rect 317 40 324 43
rect 328 44 347 47
rect 347 37 350 43
rect 375 40 382 43
rect 386 44 403 47
rect 970 50 975 53
rect 979 50 1003 53
rect 1028 50 1035 53
rect 1039 50 1061 53
rect 1081 50 1088 53
rect 1102 50 1107 53
rect 1111 50 1135 53
rect 1160 50 1167 53
rect 1171 50 1193 53
rect 1213 50 1220 53
rect 1234 50 1239 53
rect 1243 50 1267 53
rect 1292 50 1299 53
rect 1303 50 1325 53
rect 986 40 993 43
rect 997 44 1016 47
rect 1016 37 1019 43
rect 1044 40 1051 43
rect 1055 44 1070 47
rect 1118 40 1125 43
rect 1129 44 1148 47
rect 1148 37 1151 43
rect 1176 40 1183 43
rect 1187 44 1202 47
rect 1250 40 1257 43
rect 1261 44 1280 47
rect 1280 37 1283 43
rect 1308 40 1315 43
rect 1319 44 1336 47
rect 20 21 23 33
rect 41 21 44 33
rect 57 21 60 33
rect 71 24 83 27
rect 99 21 102 33
rect 115 21 118 33
rect 136 21 139 33
rect 152 21 155 33
rect 173 21 176 33
rect 189 21 192 33
rect 203 24 215 27
rect 231 21 234 33
rect 247 21 250 33
rect 268 21 271 33
rect 284 21 287 33
rect 305 21 308 33
rect 321 21 324 33
rect 335 24 347 27
rect 363 21 366 33
rect 379 21 382 33
rect 400 21 403 33
rect 953 21 956 33
rect 974 21 977 33
rect 990 21 993 33
rect 1004 24 1016 27
rect 1032 21 1035 33
rect 1048 21 1051 33
rect 1069 21 1072 33
rect 1085 21 1088 33
rect 1106 21 1109 33
rect 1122 21 1125 33
rect 1136 24 1148 27
rect 1164 21 1167 33
rect 1180 21 1183 33
rect 1201 21 1204 33
rect 1217 21 1220 33
rect 1238 21 1241 33
rect 1254 21 1257 33
rect 1268 24 1280 27
rect 1296 21 1299 33
rect 1312 21 1315 33
rect 1333 21 1336 33
rect 17 17 50 21
rect 54 17 78 21
rect 82 17 108 21
rect 112 17 182 21
rect 186 17 210 21
rect 214 17 240 21
rect 244 17 314 21
rect 318 17 342 21
rect 346 17 372 21
rect 376 17 429 21
rect 950 17 983 21
rect 987 17 1011 21
rect 1015 17 1041 21
rect 1045 17 1115 21
rect 1119 17 1143 21
rect 1147 17 1173 21
rect 1177 17 1247 21
rect 1251 17 1275 21
rect 1279 17 1305 21
rect 1309 17 1362 21
rect 17 10 26 14
rect 30 10 77 14
rect 81 10 127 14
rect 131 10 158 14
rect 162 10 209 14
rect 213 10 259 14
rect 263 10 290 14
rect 294 10 341 14
rect 345 10 391 14
rect 395 10 465 14
rect 950 10 959 14
rect 963 10 1010 14
rect 1014 10 1060 14
rect 1064 10 1091 14
rect 1095 10 1142 14
rect 1146 10 1192 14
rect 1196 10 1223 14
rect 1227 10 1274 14
rect 1278 10 1324 14
rect 1328 10 1398 14
<< m2contact >>
rect 477 1962 483 1966
rect 498 1962 502 1966
rect 534 1962 538 1966
rect 601 1962 605 1966
rect 630 1962 634 1966
rect 666 1962 670 1966
rect 733 1962 737 1966
rect 762 1962 766 1966
rect 798 1962 802 1966
rect 865 1962 869 1966
rect 894 1962 898 1966
rect 930 1962 934 1966
rect 997 1962 1001 1966
rect 1410 1962 1416 1966
rect 1431 1962 1435 1966
rect 1467 1962 1471 1966
rect 1534 1962 1538 1966
rect 1563 1962 1567 1966
rect 1599 1962 1603 1966
rect 1666 1962 1670 1966
rect 1695 1962 1699 1966
rect 1731 1962 1735 1966
rect 1798 1962 1802 1966
rect 1827 1962 1831 1966
rect 1863 1962 1867 1966
rect 1930 1962 1934 1966
rect 417 1955 423 1959
rect 1350 1955 1356 1959
rect 498 1948 502 1952
rect 548 1948 552 1952
rect 601 1948 605 1952
rect 630 1948 634 1952
rect 680 1948 684 1952
rect 733 1948 737 1952
rect 762 1948 766 1952
rect 812 1948 816 1952
rect 865 1948 869 1952
rect 894 1948 898 1952
rect 944 1948 948 1952
rect 997 1948 1001 1952
rect 1431 1948 1435 1952
rect 1481 1948 1485 1952
rect 1534 1948 1538 1952
rect 1563 1948 1567 1952
rect 1613 1948 1617 1952
rect 1666 1948 1670 1952
rect 1695 1948 1699 1952
rect 1745 1948 1749 1952
rect 1798 1948 1802 1952
rect 1827 1948 1831 1952
rect 1877 1948 1881 1952
rect 1930 1948 1934 1952
rect 521 1937 525 1941
rect 158 1929 162 1933
rect 194 1929 198 1933
rect 261 1929 265 1933
rect 477 1929 483 1933
rect 492 1928 496 1932
rect 505 1931 509 1937
rect 542 1931 546 1937
rect 555 1933 559 1937
rect 579 1937 583 1941
rect 653 1937 657 1941
rect 563 1931 567 1937
rect 600 1931 604 1937
rect 616 1933 620 1937
rect 417 1922 423 1926
rect 158 1915 162 1919
rect 208 1915 212 1919
rect 261 1915 265 1919
rect 505 1918 509 1922
rect 521 1918 525 1924
rect 555 1924 559 1928
rect 542 1918 546 1922
rect 563 1918 567 1922
rect 579 1918 583 1924
rect 624 1928 628 1932
rect 637 1931 641 1937
rect 674 1931 678 1937
rect 687 1933 691 1937
rect 711 1937 715 1941
rect 785 1937 789 1941
rect 695 1931 699 1937
rect 732 1931 736 1937
rect 748 1933 752 1937
rect 600 1918 604 1922
rect 616 1918 620 1922
rect 637 1918 641 1922
rect 653 1918 657 1924
rect 687 1924 691 1928
rect 674 1918 678 1922
rect 695 1918 699 1922
rect 711 1918 715 1924
rect 756 1928 760 1932
rect 769 1931 773 1937
rect 806 1931 810 1937
rect 819 1933 823 1937
rect 843 1937 847 1941
rect 917 1937 921 1941
rect 827 1931 831 1937
rect 864 1931 868 1937
rect 880 1933 884 1937
rect 732 1918 736 1922
rect 748 1918 752 1922
rect 769 1918 773 1922
rect 785 1918 789 1924
rect 819 1924 823 1928
rect 806 1918 810 1922
rect 827 1918 831 1922
rect 843 1918 847 1924
rect 888 1928 892 1932
rect 901 1931 905 1937
rect 938 1931 942 1937
rect 951 1933 955 1937
rect 975 1937 979 1941
rect 1454 1937 1458 1941
rect 959 1931 963 1937
rect 996 1931 1000 1937
rect 1012 1933 1016 1937
rect 1091 1929 1095 1933
rect 1127 1929 1131 1933
rect 1194 1929 1198 1933
rect 1410 1929 1416 1933
rect 864 1918 868 1922
rect 880 1918 884 1922
rect 901 1918 905 1922
rect 917 1918 921 1924
rect 951 1924 955 1928
rect 938 1918 942 1922
rect 181 1904 185 1908
rect 143 1895 147 1899
rect 165 1898 169 1904
rect 202 1898 206 1904
rect 215 1900 219 1904
rect 239 1904 243 1908
rect 223 1898 227 1904
rect 260 1898 264 1904
rect 276 1898 280 1904
rect 498 1907 502 1911
rect 535 1905 539 1909
rect 555 1905 559 1909
rect 599 1905 603 1909
rect 630 1907 634 1911
rect 667 1905 671 1909
rect 687 1905 691 1909
rect 731 1905 735 1909
rect 762 1907 766 1911
rect 799 1905 803 1909
rect 819 1905 823 1909
rect 863 1905 867 1909
rect 880 1910 884 1914
rect 959 1918 963 1922
rect 975 1918 979 1924
rect 1425 1928 1429 1932
rect 1438 1931 1442 1937
rect 1475 1931 1479 1937
rect 1488 1933 1492 1937
rect 1512 1937 1516 1941
rect 1586 1937 1590 1941
rect 1496 1931 1500 1937
rect 1533 1931 1537 1937
rect 1549 1933 1553 1937
rect 1350 1922 1356 1926
rect 996 1918 1000 1922
rect 1012 1918 1016 1922
rect 894 1907 898 1911
rect 931 1905 935 1909
rect 951 1905 955 1909
rect 995 1905 999 1909
rect 1012 1910 1016 1914
rect 1091 1915 1095 1919
rect 1141 1915 1145 1919
rect 1194 1915 1198 1919
rect 1438 1918 1442 1922
rect 1454 1918 1458 1924
rect 1488 1924 1492 1928
rect 1475 1918 1479 1922
rect 1496 1918 1500 1922
rect 1512 1918 1516 1924
rect 1557 1928 1561 1932
rect 1570 1931 1574 1937
rect 1607 1931 1611 1937
rect 1620 1933 1624 1937
rect 1644 1937 1648 1941
rect 1718 1937 1722 1941
rect 1628 1931 1632 1937
rect 1665 1931 1669 1937
rect 1681 1933 1685 1937
rect 1533 1918 1537 1922
rect 1549 1918 1553 1922
rect 1570 1918 1574 1922
rect 1586 1918 1590 1924
rect 1620 1924 1624 1928
rect 1607 1918 1611 1922
rect 1628 1918 1632 1922
rect 1644 1918 1648 1924
rect 1689 1928 1693 1932
rect 1702 1931 1706 1937
rect 1739 1931 1743 1937
rect 1752 1933 1756 1937
rect 1776 1937 1780 1941
rect 1850 1937 1854 1941
rect 1760 1931 1764 1937
rect 1797 1931 1801 1937
rect 1813 1933 1817 1937
rect 1665 1918 1669 1922
rect 1681 1918 1685 1922
rect 1702 1918 1706 1922
rect 1718 1918 1722 1924
rect 1752 1924 1756 1928
rect 1739 1918 1743 1922
rect 1760 1918 1764 1922
rect 1776 1918 1780 1924
rect 1821 1928 1825 1932
rect 1834 1931 1838 1937
rect 1871 1931 1875 1937
rect 1884 1933 1888 1937
rect 1908 1937 1912 1941
rect 1892 1931 1896 1937
rect 1929 1931 1933 1937
rect 1945 1933 1949 1937
rect 1797 1918 1801 1922
rect 1813 1918 1817 1922
rect 1834 1918 1838 1922
rect 1850 1918 1854 1924
rect 1884 1924 1888 1928
rect 1871 1918 1875 1922
rect 1114 1904 1118 1908
rect 429 1898 435 1902
rect 165 1885 169 1889
rect 181 1885 185 1891
rect 215 1891 219 1895
rect 202 1885 206 1889
rect 223 1885 227 1889
rect 239 1885 243 1891
rect 1076 1895 1080 1899
rect 1098 1898 1102 1904
rect 1135 1898 1139 1904
rect 1148 1900 1152 1904
rect 1172 1904 1176 1908
rect 1156 1898 1160 1904
rect 1193 1898 1197 1904
rect 1209 1898 1213 1904
rect 1431 1907 1435 1911
rect 1468 1905 1472 1909
rect 1488 1905 1492 1909
rect 1532 1905 1536 1909
rect 1563 1907 1567 1911
rect 1600 1905 1604 1909
rect 1620 1905 1624 1909
rect 1664 1905 1668 1909
rect 1695 1907 1699 1911
rect 1732 1905 1736 1909
rect 1752 1905 1756 1909
rect 1796 1905 1800 1909
rect 1813 1910 1817 1914
rect 1892 1918 1896 1922
rect 1908 1918 1912 1924
rect 1929 1918 1933 1922
rect 1945 1918 1949 1922
rect 1827 1907 1831 1911
rect 1864 1905 1868 1909
rect 1884 1905 1888 1909
rect 1928 1905 1932 1909
rect 1945 1910 1949 1914
rect 1362 1898 1368 1902
rect 465 1891 471 1895
rect 498 1891 502 1895
rect 549 1891 553 1895
rect 599 1891 603 1895
rect 630 1891 634 1895
rect 681 1891 685 1895
rect 731 1891 735 1895
rect 762 1891 766 1895
rect 813 1891 817 1895
rect 863 1891 867 1895
rect 894 1891 898 1895
rect 945 1891 949 1895
rect 995 1891 999 1895
rect 260 1885 264 1889
rect 276 1885 280 1889
rect 1098 1885 1102 1889
rect 1114 1885 1118 1891
rect 1148 1891 1152 1895
rect 1135 1885 1139 1889
rect 158 1874 162 1878
rect 195 1872 199 1876
rect 215 1872 219 1876
rect 259 1872 263 1876
rect 417 1878 423 1882
rect 496 1878 500 1882
rect 530 1878 534 1882
rect 547 1878 551 1882
rect 603 1878 607 1882
rect 620 1878 624 1882
rect 648 1878 652 1882
rect 1156 1885 1160 1889
rect 1172 1885 1176 1891
rect 1398 1891 1404 1895
rect 1431 1891 1435 1895
rect 1482 1891 1486 1895
rect 1532 1891 1536 1895
rect 1563 1891 1567 1895
rect 1614 1891 1618 1895
rect 1664 1891 1668 1895
rect 1695 1891 1699 1895
rect 1746 1891 1750 1895
rect 1796 1891 1800 1895
rect 1827 1891 1831 1895
rect 1878 1891 1882 1895
rect 1928 1891 1932 1895
rect 1193 1885 1197 1889
rect 1209 1885 1213 1889
rect 453 1871 459 1875
rect 523 1871 527 1875
rect 554 1871 558 1875
rect 576 1871 580 1875
rect 641 1871 645 1875
rect 429 1865 435 1869
rect 158 1858 162 1862
rect 209 1858 213 1862
rect 259 1858 263 1862
rect 465 1858 471 1862
rect 497 1861 501 1865
rect 522 1864 526 1868
rect 529 1861 533 1865
rect 547 1861 551 1865
rect 569 1864 573 1868
rect 594 1864 598 1868
rect 604 1861 608 1865
rect 620 1861 624 1865
rect 640 1864 644 1868
rect 647 1861 651 1865
rect 711 1871 715 1875
rect 276 1851 280 1855
rect 143 1842 147 1846
rect 268 1844 272 1848
rect 292 1844 296 1848
rect 151 1835 155 1839
rect 292 1835 296 1839
rect 524 1845 528 1849
rect 544 1842 548 1846
rect 563 1846 567 1850
rect 665 1857 669 1861
rect 680 1857 684 1861
rect 582 1845 586 1849
rect 601 1845 605 1849
rect 614 1844 618 1848
rect 636 1845 640 1849
rect 644 1844 648 1848
rect 656 1844 660 1848
rect 497 1831 501 1835
rect 529 1831 533 1835
rect 547 1831 551 1835
rect 604 1831 608 1835
rect 619 1831 623 1835
rect 647 1831 651 1835
rect 158 1827 162 1831
rect 225 1827 229 1831
rect 261 1827 265 1831
rect 477 1827 483 1831
rect 511 1827 515 1831
rect 554 1826 558 1830
rect 576 1827 583 1831
rect 626 1826 630 1830
rect 417 1820 423 1824
rect 158 1813 162 1817
rect 211 1813 215 1817
rect 261 1813 265 1817
rect 441 1819 447 1823
rect 511 1819 515 1823
rect 570 1819 574 1823
rect 595 1819 599 1823
rect 626 1819 630 1823
rect 719 1849 723 1857
rect 792 1871 796 1875
rect 746 1857 750 1861
rect 761 1857 765 1861
rect 1091 1874 1095 1878
rect 1128 1872 1132 1876
rect 1148 1872 1152 1876
rect 1192 1872 1196 1876
rect 1350 1878 1356 1882
rect 1429 1878 1433 1882
rect 1463 1878 1467 1882
rect 1480 1878 1484 1882
rect 1536 1878 1540 1882
rect 1553 1878 1557 1882
rect 1581 1878 1585 1882
rect 1386 1871 1392 1875
rect 1456 1871 1460 1875
rect 1487 1871 1491 1875
rect 1509 1871 1513 1875
rect 1574 1871 1578 1875
rect 742 1849 746 1853
rect 688 1843 692 1847
rect 701 1835 705 1839
rect 800 1849 804 1857
rect 1362 1865 1368 1869
rect 1091 1858 1095 1862
rect 1142 1858 1146 1862
rect 1192 1858 1196 1862
rect 1398 1858 1404 1862
rect 1430 1861 1434 1865
rect 1455 1864 1459 1868
rect 1462 1861 1466 1865
rect 1480 1861 1484 1865
rect 1502 1864 1506 1868
rect 1527 1864 1531 1868
rect 1537 1861 1541 1865
rect 1553 1861 1557 1865
rect 1573 1864 1577 1868
rect 1580 1861 1584 1865
rect 1644 1871 1648 1875
rect 827 1849 831 1853
rect 1209 1851 1213 1855
rect 769 1843 773 1847
rect 1076 1842 1080 1846
rect 1201 1844 1205 1848
rect 1225 1844 1229 1848
rect 782 1835 786 1839
rect 1084 1835 1088 1839
rect 1225 1835 1229 1839
rect 1457 1845 1461 1849
rect 1477 1842 1481 1846
rect 1496 1846 1500 1850
rect 1598 1857 1602 1861
rect 1613 1857 1617 1861
rect 1515 1845 1519 1849
rect 1534 1845 1538 1849
rect 1547 1844 1551 1848
rect 1569 1845 1573 1849
rect 1577 1844 1581 1848
rect 1589 1844 1593 1848
rect 1430 1831 1434 1835
rect 1462 1831 1466 1835
rect 1480 1831 1484 1835
rect 1537 1831 1541 1835
rect 1552 1831 1556 1835
rect 1580 1831 1584 1835
rect 1091 1827 1095 1831
rect 1158 1827 1162 1831
rect 1194 1827 1198 1831
rect 1410 1827 1416 1831
rect 1444 1827 1448 1831
rect 1487 1826 1491 1830
rect 1509 1827 1516 1831
rect 1559 1826 1563 1830
rect 1350 1820 1356 1824
rect 429 1812 435 1816
rect 497 1812 501 1816
rect 511 1812 515 1816
rect 529 1812 533 1816
rect 547 1812 551 1816
rect 570 1812 574 1816
rect 604 1812 608 1816
rect 619 1812 623 1816
rect 647 1812 651 1816
rect 180 1802 184 1806
rect 143 1796 147 1802
rect 159 1796 163 1802
rect 196 1796 200 1802
rect 204 1798 208 1802
rect 238 1802 242 1806
rect 441 1805 447 1809
rect 511 1805 515 1809
rect 570 1805 574 1809
rect 595 1805 599 1809
rect 626 1805 630 1809
rect 217 1796 221 1802
rect 254 1796 258 1802
rect 511 1797 515 1801
rect 554 1798 558 1802
rect 576 1797 583 1801
rect 626 1798 630 1802
rect 276 1793 280 1797
rect 497 1793 501 1797
rect 529 1793 533 1797
rect 547 1793 551 1797
rect 604 1793 608 1797
rect 619 1793 623 1797
rect 647 1793 651 1797
rect 143 1783 147 1787
rect 159 1783 163 1787
rect 204 1789 208 1793
rect 180 1783 184 1789
rect 196 1783 200 1787
rect 217 1783 221 1787
rect 238 1783 242 1789
rect 254 1783 258 1787
rect 492 1781 496 1785
rect 160 1770 164 1774
rect 204 1770 208 1774
rect 224 1770 228 1774
rect 261 1772 265 1776
rect 524 1779 528 1783
rect 544 1782 548 1786
rect 563 1778 567 1782
rect 582 1779 586 1783
rect 601 1779 605 1783
rect 614 1780 618 1784
rect 711 1795 715 1799
rect 1091 1813 1095 1817
rect 1144 1813 1148 1817
rect 1194 1813 1198 1817
rect 1374 1819 1380 1823
rect 1444 1819 1448 1823
rect 1503 1819 1507 1823
rect 1528 1819 1532 1823
rect 1559 1819 1563 1823
rect 1652 1849 1656 1857
rect 1725 1871 1729 1875
rect 1679 1857 1683 1861
rect 1694 1857 1698 1861
rect 1675 1849 1679 1853
rect 1621 1843 1625 1847
rect 1634 1835 1638 1839
rect 1733 1849 1737 1857
rect 1760 1849 1764 1853
rect 1702 1843 1706 1847
rect 1715 1835 1719 1839
rect 1362 1812 1368 1816
rect 1430 1812 1434 1816
rect 1444 1812 1448 1816
rect 1462 1812 1466 1816
rect 1480 1812 1484 1816
rect 1503 1812 1507 1816
rect 1537 1812 1541 1816
rect 1552 1812 1556 1816
rect 1580 1812 1584 1816
rect 1113 1802 1117 1806
rect 792 1795 796 1799
rect 1076 1796 1080 1802
rect 1092 1796 1096 1802
rect 1129 1796 1133 1802
rect 1137 1798 1141 1802
rect 1171 1802 1175 1806
rect 1374 1805 1380 1809
rect 1444 1805 1448 1809
rect 1503 1805 1507 1809
rect 1528 1805 1532 1809
rect 1559 1805 1563 1809
rect 1150 1796 1154 1802
rect 1187 1796 1191 1802
rect 1444 1797 1448 1801
rect 1487 1798 1491 1802
rect 1509 1797 1516 1801
rect 1559 1798 1563 1802
rect 1209 1793 1213 1797
rect 1430 1793 1434 1797
rect 1462 1793 1466 1797
rect 1480 1793 1484 1797
rect 1537 1793 1541 1797
rect 1552 1793 1556 1797
rect 1580 1793 1584 1797
rect 636 1779 640 1783
rect 644 1780 648 1784
rect 656 1780 660 1784
rect 691 1780 695 1784
rect 719 1779 723 1783
rect 771 1780 775 1784
rect 1076 1783 1080 1787
rect 1092 1783 1096 1787
rect 1137 1789 1141 1793
rect 1113 1783 1117 1789
rect 1129 1783 1133 1787
rect 800 1779 804 1783
rect 1150 1783 1154 1787
rect 1171 1783 1175 1789
rect 1187 1783 1191 1787
rect 1425 1781 1429 1785
rect 429 1763 435 1767
rect 497 1763 501 1767
rect 522 1760 526 1764
rect 529 1763 533 1767
rect 547 1763 551 1767
rect 569 1760 573 1764
rect 594 1760 598 1764
rect 604 1763 608 1767
rect 620 1763 624 1767
rect 640 1760 644 1764
rect 647 1763 651 1767
rect 160 1756 164 1760
rect 210 1756 214 1760
rect 261 1756 265 1760
rect 465 1756 471 1760
rect 507 1753 511 1757
rect 523 1753 527 1757
rect 554 1753 558 1757
rect 576 1753 580 1757
rect 641 1753 645 1757
rect 701 1759 705 1763
rect 1093 1770 1097 1774
rect 1137 1770 1141 1774
rect 1157 1770 1161 1774
rect 1194 1772 1198 1776
rect 1457 1779 1461 1783
rect 1477 1782 1481 1786
rect 1496 1778 1500 1782
rect 1515 1779 1519 1783
rect 1534 1779 1538 1783
rect 1547 1780 1551 1784
rect 1644 1795 1648 1799
rect 1725 1795 1729 1799
rect 1569 1779 1573 1783
rect 1577 1780 1581 1784
rect 1589 1780 1593 1784
rect 1624 1780 1628 1784
rect 1652 1779 1656 1783
rect 1704 1780 1708 1784
rect 1733 1779 1737 1783
rect 1362 1763 1368 1767
rect 1430 1763 1434 1767
rect 782 1759 786 1763
rect 1455 1760 1459 1764
rect 1462 1763 1466 1767
rect 1480 1763 1484 1767
rect 1502 1760 1506 1764
rect 1527 1760 1531 1764
rect 1537 1763 1541 1767
rect 1553 1763 1557 1767
rect 1573 1760 1577 1764
rect 1580 1763 1584 1767
rect 1093 1756 1097 1760
rect 1143 1756 1147 1760
rect 1194 1756 1198 1760
rect 1398 1756 1404 1760
rect 1440 1753 1444 1757
rect 1456 1753 1460 1757
rect 1487 1753 1491 1757
rect 1509 1753 1513 1757
rect 1574 1753 1578 1757
rect 1634 1759 1638 1763
rect 1715 1759 1719 1763
rect 417 1746 423 1750
rect 496 1746 500 1750
rect 530 1746 534 1750
rect 547 1746 551 1750
rect 603 1746 607 1750
rect 620 1746 624 1750
rect 648 1746 652 1750
rect 1350 1746 1356 1750
rect 1429 1746 1433 1750
rect 1463 1746 1467 1750
rect 1480 1746 1484 1750
rect 1536 1746 1540 1750
rect 1553 1746 1557 1750
rect 1581 1746 1585 1750
rect 453 1739 459 1743
rect 507 1739 511 1743
rect 523 1739 527 1743
rect 554 1739 558 1743
rect 576 1739 580 1743
rect 641 1739 645 1743
rect 711 1739 715 1743
rect 497 1729 501 1733
rect 522 1732 526 1736
rect 529 1729 533 1733
rect 547 1729 551 1733
rect 569 1732 573 1736
rect 594 1732 598 1736
rect 604 1729 608 1733
rect 620 1729 624 1733
rect 640 1732 644 1736
rect 647 1729 651 1733
rect 491 1712 495 1716
rect 524 1713 528 1717
rect 544 1710 548 1714
rect 563 1714 567 1718
rect 582 1713 586 1717
rect 601 1713 605 1717
rect 614 1712 618 1716
rect 636 1713 640 1717
rect 644 1712 648 1716
rect 656 1712 660 1716
rect 719 1717 723 1725
rect 816 1739 820 1743
rect 770 1725 774 1729
rect 785 1725 789 1729
rect 1386 1739 1392 1743
rect 1440 1739 1444 1743
rect 1456 1739 1460 1743
rect 1487 1739 1491 1743
rect 1509 1739 1513 1743
rect 1574 1739 1578 1743
rect 1644 1739 1648 1743
rect 688 1711 692 1715
rect 742 1716 746 1720
rect 497 1699 501 1703
rect 529 1699 533 1703
rect 547 1699 551 1703
rect 604 1699 608 1703
rect 619 1699 623 1703
rect 647 1699 651 1703
rect 511 1695 515 1699
rect 554 1694 558 1698
rect 576 1695 583 1699
rect 626 1694 630 1698
rect 441 1687 447 1691
rect 511 1687 515 1691
rect 570 1687 574 1691
rect 595 1687 599 1691
rect 626 1687 630 1691
rect 701 1703 705 1707
rect 824 1717 828 1725
rect 1430 1729 1434 1733
rect 1455 1732 1459 1736
rect 1462 1729 1466 1733
rect 1480 1729 1484 1733
rect 1502 1732 1506 1736
rect 1527 1732 1531 1736
rect 1537 1729 1541 1733
rect 1553 1729 1557 1733
rect 1573 1732 1577 1736
rect 1580 1729 1584 1733
rect 845 1717 849 1721
rect 793 1711 797 1715
rect 1424 1712 1428 1716
rect 806 1703 810 1707
rect 1457 1713 1461 1717
rect 1477 1710 1481 1714
rect 1496 1714 1500 1718
rect 1515 1713 1519 1717
rect 1534 1713 1538 1717
rect 1547 1712 1551 1716
rect 1569 1713 1573 1717
rect 1577 1712 1581 1716
rect 1589 1712 1593 1716
rect 1652 1717 1656 1725
rect 1749 1739 1753 1743
rect 1703 1725 1707 1729
rect 1718 1725 1722 1729
rect 1621 1711 1625 1715
rect 1675 1716 1679 1720
rect 1430 1699 1434 1703
rect 1462 1699 1466 1703
rect 1480 1699 1484 1703
rect 1537 1699 1541 1703
rect 1552 1699 1556 1703
rect 1580 1699 1584 1703
rect 1444 1695 1448 1699
rect 1487 1694 1491 1698
rect 1509 1695 1516 1699
rect 1559 1694 1563 1698
rect 1374 1687 1380 1691
rect 1444 1687 1448 1691
rect 1503 1687 1507 1691
rect 1528 1687 1532 1691
rect 1559 1687 1563 1691
rect 1634 1703 1638 1707
rect 1757 1717 1761 1725
rect 1778 1717 1782 1721
rect 1726 1711 1730 1715
rect 1739 1703 1743 1707
rect 429 1680 435 1684
rect 497 1680 501 1684
rect 511 1680 515 1684
rect 529 1680 533 1684
rect 547 1680 551 1684
rect 570 1680 574 1684
rect 604 1680 608 1684
rect 619 1680 623 1684
rect 647 1680 651 1684
rect 1362 1680 1368 1684
rect 1430 1680 1434 1684
rect 1444 1680 1448 1684
rect 1462 1680 1466 1684
rect 1480 1680 1484 1684
rect 1503 1680 1507 1684
rect 1537 1680 1541 1684
rect 1552 1680 1556 1684
rect 1580 1680 1584 1684
rect 441 1673 447 1677
rect 511 1673 515 1677
rect 570 1673 574 1677
rect 595 1673 599 1677
rect 626 1673 630 1677
rect 511 1665 515 1669
rect 554 1666 558 1670
rect 576 1665 583 1669
rect 626 1666 630 1670
rect 497 1661 501 1665
rect 529 1661 533 1665
rect 547 1661 551 1665
rect 604 1661 608 1665
rect 619 1661 623 1665
rect 647 1661 651 1665
rect 711 1664 715 1668
rect 1374 1673 1380 1677
rect 1444 1673 1448 1677
rect 1503 1673 1507 1677
rect 1528 1673 1532 1677
rect 1559 1673 1563 1677
rect 816 1664 820 1668
rect 1444 1665 1448 1669
rect 1487 1666 1491 1670
rect 1509 1665 1516 1669
rect 1559 1666 1563 1670
rect 1430 1661 1434 1665
rect 1462 1661 1466 1665
rect 1480 1661 1484 1665
rect 1537 1661 1541 1665
rect 1552 1661 1556 1665
rect 1580 1661 1584 1665
rect 1644 1664 1648 1668
rect 1749 1664 1753 1668
rect 492 1649 496 1653
rect 524 1647 528 1651
rect 544 1650 548 1654
rect 563 1646 567 1650
rect 582 1647 586 1651
rect 601 1647 605 1651
rect 614 1648 618 1652
rect 636 1647 640 1651
rect 644 1648 648 1652
rect 656 1648 660 1652
rect 690 1649 694 1653
rect 719 1648 723 1652
rect 796 1649 800 1653
rect 824 1648 828 1652
rect 1425 1649 1429 1653
rect 497 1631 501 1635
rect 522 1628 526 1632
rect 529 1631 533 1635
rect 547 1631 551 1635
rect 569 1628 573 1632
rect 594 1628 598 1632
rect 604 1631 608 1635
rect 620 1631 624 1635
rect 640 1628 644 1632
rect 647 1631 651 1635
rect 453 1621 459 1625
rect 523 1621 527 1625
rect 554 1621 558 1625
rect 576 1621 580 1625
rect 641 1621 645 1625
rect 701 1628 705 1632
rect 1457 1647 1461 1651
rect 1477 1650 1481 1654
rect 1496 1646 1500 1650
rect 1515 1647 1519 1651
rect 1534 1647 1538 1651
rect 1547 1648 1551 1652
rect 1569 1647 1573 1651
rect 1577 1648 1581 1652
rect 1589 1648 1593 1652
rect 1623 1649 1627 1653
rect 1652 1648 1656 1652
rect 1729 1649 1733 1653
rect 1757 1648 1761 1652
rect 806 1628 810 1632
rect 1430 1631 1434 1635
rect 1455 1628 1459 1632
rect 1462 1631 1466 1635
rect 1480 1631 1484 1635
rect 1502 1628 1506 1632
rect 1527 1628 1531 1632
rect 1537 1631 1541 1635
rect 1553 1631 1557 1635
rect 1573 1628 1577 1632
rect 1580 1631 1584 1635
rect 1386 1621 1392 1625
rect 1456 1621 1460 1625
rect 1487 1621 1491 1625
rect 1509 1621 1513 1625
rect 1574 1621 1578 1625
rect 1634 1628 1638 1632
rect 1739 1628 1743 1632
rect 417 1614 423 1618
rect 496 1614 500 1618
rect 530 1614 534 1618
rect 547 1614 551 1618
rect 603 1614 607 1618
rect 620 1614 624 1618
rect 648 1614 652 1618
rect 1350 1614 1356 1618
rect 1429 1614 1433 1618
rect 1463 1614 1467 1618
rect 1480 1614 1484 1618
rect 1536 1614 1540 1618
rect 1553 1614 1557 1618
rect 1581 1614 1585 1618
rect 453 1607 459 1611
rect 523 1607 527 1611
rect 554 1607 558 1611
rect 576 1607 580 1611
rect 641 1607 645 1611
rect 711 1607 715 1611
rect 497 1597 501 1601
rect 522 1600 526 1604
rect 529 1597 533 1601
rect 547 1597 551 1601
rect 569 1600 573 1604
rect 594 1600 598 1604
rect 604 1597 608 1601
rect 620 1597 624 1601
rect 640 1600 644 1604
rect 647 1597 651 1601
rect 491 1580 495 1584
rect 524 1581 528 1585
rect 544 1578 548 1582
rect 563 1582 567 1586
rect 582 1581 586 1585
rect 601 1581 605 1585
rect 614 1580 618 1584
rect 636 1581 640 1585
rect 644 1580 648 1584
rect 656 1580 660 1584
rect 719 1585 723 1593
rect 792 1607 796 1611
rect 746 1593 750 1597
rect 761 1593 765 1597
rect 742 1585 746 1589
rect 688 1579 692 1583
rect 497 1567 501 1571
rect 529 1567 533 1571
rect 547 1567 551 1571
rect 604 1567 608 1571
rect 619 1567 623 1571
rect 647 1567 651 1571
rect 511 1563 515 1567
rect 554 1562 558 1566
rect 576 1563 583 1567
rect 626 1562 630 1566
rect 441 1555 447 1559
rect 511 1555 515 1559
rect 570 1555 574 1559
rect 595 1555 599 1559
rect 626 1555 630 1559
rect 701 1571 705 1575
rect 800 1585 804 1593
rect 882 1607 886 1611
rect 836 1593 840 1597
rect 851 1593 855 1597
rect 1386 1607 1392 1611
rect 1456 1607 1460 1611
rect 1487 1607 1491 1611
rect 1509 1607 1513 1611
rect 1574 1607 1578 1611
rect 1644 1607 1648 1611
rect 824 1585 828 1589
rect 769 1579 773 1583
rect 858 1587 862 1591
rect 890 1585 894 1593
rect 1430 1597 1434 1601
rect 1455 1600 1459 1604
rect 1462 1597 1466 1601
rect 1480 1597 1484 1601
rect 1502 1600 1506 1604
rect 1527 1600 1531 1604
rect 1537 1597 1541 1601
rect 1553 1597 1557 1601
rect 1573 1600 1577 1604
rect 1580 1597 1584 1601
rect 782 1571 786 1575
rect 925 1584 929 1588
rect 1424 1580 1428 1584
rect 872 1571 876 1575
rect 1457 1581 1461 1585
rect 1477 1578 1481 1582
rect 1496 1582 1500 1586
rect 1515 1581 1519 1585
rect 1534 1581 1538 1585
rect 1547 1580 1551 1584
rect 1569 1581 1573 1585
rect 1577 1580 1581 1584
rect 1589 1580 1593 1584
rect 1652 1585 1656 1593
rect 1725 1607 1729 1611
rect 1679 1593 1683 1597
rect 1694 1593 1698 1597
rect 1675 1585 1679 1589
rect 1621 1579 1625 1583
rect 1430 1567 1434 1571
rect 1462 1567 1466 1571
rect 1480 1567 1484 1571
rect 1537 1567 1541 1571
rect 1552 1567 1556 1571
rect 1580 1567 1584 1571
rect 1444 1563 1448 1567
rect 1487 1562 1491 1566
rect 1509 1563 1516 1567
rect 1559 1562 1563 1566
rect 1374 1555 1380 1559
rect 1444 1555 1448 1559
rect 1503 1555 1507 1559
rect 1528 1555 1532 1559
rect 1559 1555 1563 1559
rect 1634 1571 1638 1575
rect 1733 1585 1737 1593
rect 1815 1607 1819 1611
rect 1769 1593 1773 1597
rect 1784 1593 1788 1597
rect 1757 1585 1761 1589
rect 1702 1579 1706 1583
rect 1791 1587 1795 1591
rect 1823 1585 1827 1593
rect 1715 1571 1719 1575
rect 1858 1584 1862 1588
rect 1805 1571 1809 1575
rect 429 1548 435 1552
rect 497 1548 501 1552
rect 511 1548 515 1552
rect 529 1548 533 1552
rect 547 1548 551 1552
rect 570 1548 574 1552
rect 604 1548 608 1552
rect 619 1548 623 1552
rect 647 1548 651 1552
rect 1362 1548 1368 1552
rect 1430 1548 1434 1552
rect 1444 1548 1448 1552
rect 1462 1548 1466 1552
rect 1480 1548 1484 1552
rect 1503 1548 1507 1552
rect 1537 1548 1541 1552
rect 1552 1548 1556 1552
rect 1580 1548 1584 1552
rect 441 1541 447 1545
rect 511 1541 515 1545
rect 570 1541 574 1545
rect 595 1541 599 1545
rect 626 1541 630 1545
rect 511 1533 515 1537
rect 554 1534 558 1538
rect 576 1533 583 1537
rect 626 1534 630 1538
rect 497 1529 501 1533
rect 529 1529 533 1533
rect 547 1529 551 1533
rect 604 1529 608 1533
rect 619 1529 623 1533
rect 647 1529 651 1533
rect 492 1517 496 1521
rect 524 1515 528 1519
rect 544 1518 548 1522
rect 563 1514 567 1518
rect 582 1515 586 1519
rect 601 1515 605 1519
rect 614 1516 618 1520
rect 711 1529 715 1533
rect 792 1529 796 1533
rect 1374 1541 1380 1545
rect 1444 1541 1448 1545
rect 1503 1541 1507 1545
rect 1528 1541 1532 1545
rect 1559 1541 1563 1545
rect 1444 1533 1448 1537
rect 1487 1534 1491 1538
rect 1509 1533 1516 1537
rect 1559 1534 1563 1538
rect 882 1529 886 1533
rect 1430 1529 1434 1533
rect 1462 1529 1466 1533
rect 1480 1529 1484 1533
rect 1537 1529 1541 1533
rect 1552 1529 1556 1533
rect 1580 1529 1584 1533
rect 636 1515 640 1519
rect 644 1516 648 1520
rect 656 1516 660 1520
rect 691 1514 695 1518
rect 719 1513 723 1517
rect 771 1514 775 1518
rect 800 1513 804 1517
rect 855 1514 859 1518
rect 1425 1517 1429 1521
rect 890 1513 894 1517
rect 497 1499 501 1503
rect 522 1496 526 1500
rect 529 1499 533 1503
rect 547 1499 551 1503
rect 569 1496 573 1500
rect 594 1496 598 1500
rect 604 1499 608 1503
rect 620 1499 624 1503
rect 640 1496 644 1500
rect 647 1499 651 1503
rect 1457 1515 1461 1519
rect 1477 1518 1481 1522
rect 1496 1514 1500 1518
rect 1515 1515 1519 1519
rect 1534 1515 1538 1519
rect 1547 1516 1551 1520
rect 1644 1529 1648 1533
rect 1725 1529 1729 1533
rect 1815 1529 1819 1533
rect 1569 1515 1573 1519
rect 1577 1516 1581 1520
rect 1589 1516 1593 1520
rect 1624 1514 1628 1518
rect 1652 1513 1656 1517
rect 1704 1514 1708 1518
rect 1733 1513 1737 1517
rect 1788 1514 1792 1518
rect 1823 1513 1827 1517
rect 453 1489 459 1493
rect 523 1489 527 1493
rect 554 1489 558 1493
rect 576 1489 580 1493
rect 641 1489 645 1493
rect 701 1493 705 1497
rect 782 1493 786 1497
rect 1430 1499 1434 1503
rect 872 1493 876 1497
rect 1455 1496 1459 1500
rect 1462 1499 1466 1503
rect 1480 1499 1484 1503
rect 1502 1496 1506 1500
rect 1527 1496 1531 1500
rect 1537 1499 1541 1503
rect 1553 1499 1557 1503
rect 1573 1496 1577 1500
rect 1580 1499 1584 1503
rect 1386 1489 1392 1493
rect 1456 1489 1460 1493
rect 1487 1489 1491 1493
rect 1509 1489 1513 1493
rect 1574 1489 1578 1493
rect 1634 1493 1638 1497
rect 1715 1493 1719 1497
rect 1805 1493 1809 1497
rect 417 1482 423 1486
rect 496 1482 500 1486
rect 530 1482 534 1486
rect 547 1482 551 1486
rect 603 1482 607 1486
rect 620 1482 624 1486
rect 648 1482 652 1486
rect 1350 1482 1356 1486
rect 1429 1482 1433 1486
rect 1463 1482 1467 1486
rect 1480 1482 1484 1486
rect 1536 1482 1540 1486
rect 1553 1482 1557 1486
rect 1581 1482 1585 1486
rect 453 1475 459 1479
rect 523 1475 527 1479
rect 554 1475 558 1479
rect 576 1475 580 1479
rect 641 1475 645 1479
rect 711 1475 715 1479
rect 497 1465 501 1469
rect 522 1468 526 1472
rect 529 1465 533 1469
rect 547 1465 551 1469
rect 569 1468 573 1472
rect 594 1468 598 1472
rect 604 1465 608 1469
rect 620 1465 624 1469
rect 640 1468 644 1472
rect 647 1465 651 1469
rect 491 1448 495 1452
rect 524 1449 528 1453
rect 544 1446 548 1450
rect 563 1450 567 1454
rect 1386 1475 1392 1479
rect 1456 1475 1460 1479
rect 1487 1475 1491 1479
rect 1509 1475 1513 1479
rect 1574 1475 1578 1479
rect 1644 1475 1648 1479
rect 582 1449 586 1453
rect 601 1449 605 1453
rect 614 1448 618 1452
rect 636 1449 640 1453
rect 644 1448 648 1452
rect 656 1448 660 1452
rect 719 1453 723 1461
rect 1430 1465 1434 1469
rect 1455 1468 1459 1472
rect 1462 1465 1466 1469
rect 1480 1465 1484 1469
rect 1502 1468 1506 1472
rect 1527 1468 1531 1472
rect 1537 1465 1541 1469
rect 1553 1465 1557 1469
rect 1573 1468 1577 1472
rect 1580 1465 1584 1469
rect 688 1447 692 1451
rect 742 1452 746 1456
rect 1424 1448 1428 1452
rect 497 1435 501 1439
rect 529 1435 533 1439
rect 547 1435 551 1439
rect 604 1435 608 1439
rect 619 1435 623 1439
rect 647 1435 651 1439
rect 511 1431 515 1435
rect 26 1427 30 1431
rect 62 1427 66 1431
rect 129 1427 133 1431
rect 158 1427 162 1431
rect 194 1427 198 1431
rect 261 1427 265 1431
rect 290 1427 294 1431
rect 326 1427 330 1431
rect 393 1427 397 1431
rect 477 1427 483 1431
rect 554 1430 558 1434
rect 576 1431 583 1435
rect 626 1430 630 1434
rect 417 1420 423 1424
rect 511 1423 515 1427
rect 520 1423 524 1427
rect 570 1423 574 1427
rect 595 1423 599 1427
rect 626 1423 630 1427
rect 701 1439 705 1443
rect 1457 1449 1461 1453
rect 1477 1446 1481 1450
rect 1496 1450 1500 1454
rect 1515 1449 1519 1453
rect 1534 1449 1538 1453
rect 1547 1448 1551 1452
rect 1569 1449 1573 1453
rect 1577 1448 1581 1452
rect 1589 1448 1593 1452
rect 1652 1453 1656 1461
rect 1621 1447 1625 1451
rect 1675 1452 1679 1456
rect 1430 1435 1434 1439
rect 1462 1435 1466 1439
rect 1480 1435 1484 1439
rect 1537 1435 1541 1439
rect 1552 1435 1556 1439
rect 1580 1435 1584 1439
rect 1444 1431 1448 1435
rect 959 1427 963 1431
rect 995 1427 999 1431
rect 1062 1427 1066 1431
rect 1091 1427 1095 1431
rect 1127 1427 1131 1431
rect 1194 1427 1198 1431
rect 1223 1427 1227 1431
rect 1259 1427 1263 1431
rect 1326 1427 1330 1431
rect 1410 1427 1416 1431
rect 1487 1430 1491 1434
rect 1509 1431 1516 1435
rect 1559 1430 1563 1434
rect 1350 1420 1356 1424
rect 1444 1423 1448 1427
rect 1453 1423 1457 1427
rect 1503 1423 1507 1427
rect 1528 1423 1532 1427
rect 1559 1423 1563 1427
rect 1634 1439 1638 1443
rect 26 1413 30 1417
rect 76 1413 80 1417
rect 129 1413 133 1417
rect 158 1413 162 1417
rect 208 1413 212 1417
rect 261 1413 265 1417
rect 290 1413 294 1417
rect 340 1413 344 1417
rect 393 1413 397 1417
rect 429 1416 435 1420
rect 497 1416 501 1420
rect 511 1416 515 1420
rect 529 1416 533 1420
rect 547 1416 551 1420
rect 570 1416 574 1420
rect 604 1416 608 1420
rect 619 1416 623 1420
rect 647 1416 651 1420
rect 772 1416 776 1420
rect 790 1416 794 1420
rect 808 1416 812 1420
rect 831 1416 835 1420
rect 865 1416 869 1420
rect 880 1416 884 1420
rect 908 1416 912 1420
rect 49 1402 53 1406
rect 20 1393 24 1397
rect 33 1396 37 1402
rect 70 1396 74 1402
rect 83 1398 87 1402
rect 107 1402 111 1406
rect 181 1402 185 1406
rect 91 1396 95 1402
rect 128 1396 132 1402
rect 144 1396 148 1402
rect 165 1396 169 1402
rect 202 1396 206 1402
rect 215 1398 219 1402
rect 239 1402 243 1406
rect 313 1402 317 1406
rect 223 1396 227 1402
rect 260 1396 264 1402
rect 276 1396 280 1402
rect 297 1396 301 1402
rect 334 1396 338 1402
rect 347 1398 351 1402
rect 371 1402 375 1406
rect 441 1409 447 1413
rect 511 1409 515 1413
rect 520 1409 524 1413
rect 570 1409 574 1413
rect 595 1409 599 1413
rect 626 1409 630 1413
rect 355 1396 359 1402
rect 392 1396 396 1402
rect 408 1398 412 1402
rect 511 1401 515 1405
rect 554 1402 558 1406
rect 576 1401 583 1405
rect 626 1402 630 1406
rect 497 1397 501 1401
rect 529 1397 533 1401
rect 547 1397 551 1401
rect 604 1397 608 1401
rect 619 1397 623 1401
rect 647 1397 651 1401
rect 33 1383 37 1387
rect 49 1383 53 1389
rect 83 1389 87 1393
rect 70 1383 74 1387
rect 91 1383 95 1387
rect 107 1383 111 1389
rect 128 1383 132 1387
rect 144 1383 148 1387
rect 165 1383 169 1387
rect 181 1383 185 1389
rect 215 1389 219 1393
rect 202 1383 206 1387
rect 223 1383 227 1387
rect 239 1383 243 1389
rect 260 1383 264 1387
rect 276 1383 280 1387
rect 297 1383 301 1387
rect 313 1383 317 1389
rect 347 1389 351 1393
rect 334 1383 338 1387
rect 355 1383 359 1387
rect 371 1383 375 1389
rect 392 1383 396 1387
rect 408 1383 412 1387
rect 492 1385 496 1389
rect 26 1372 30 1376
rect 63 1370 67 1374
rect 83 1370 87 1374
rect 127 1370 131 1374
rect 158 1372 162 1376
rect 195 1370 199 1374
rect 215 1370 219 1374
rect 259 1370 263 1374
rect 290 1372 294 1376
rect 327 1370 331 1374
rect 347 1370 351 1374
rect 391 1370 395 1374
rect 524 1383 528 1387
rect 544 1386 548 1390
rect 563 1382 567 1386
rect 582 1383 586 1387
rect 601 1383 605 1387
rect 614 1384 618 1388
rect 750 1409 754 1413
rect 772 1409 776 1413
rect 831 1409 835 1413
rect 856 1409 860 1413
rect 887 1409 891 1413
rect 959 1413 963 1417
rect 1009 1413 1013 1417
rect 1062 1413 1066 1417
rect 1091 1413 1095 1417
rect 1141 1413 1145 1417
rect 1194 1413 1198 1417
rect 1223 1413 1227 1417
rect 1273 1413 1277 1417
rect 1326 1413 1330 1417
rect 1362 1416 1368 1420
rect 1430 1416 1434 1420
rect 1444 1416 1448 1420
rect 1462 1416 1466 1420
rect 1480 1416 1484 1420
rect 1503 1416 1507 1420
rect 1537 1416 1541 1420
rect 1552 1416 1556 1420
rect 1580 1416 1584 1420
rect 1705 1416 1709 1420
rect 1723 1416 1727 1420
rect 1741 1416 1745 1420
rect 1764 1416 1768 1420
rect 1798 1416 1802 1420
rect 1813 1416 1817 1420
rect 1841 1416 1845 1420
rect 772 1401 776 1405
rect 815 1402 819 1406
rect 837 1401 844 1405
rect 887 1402 891 1406
rect 982 1402 986 1406
rect 790 1397 794 1401
rect 808 1397 812 1401
rect 865 1397 869 1401
rect 880 1397 884 1401
rect 908 1397 912 1401
rect 711 1393 715 1397
rect 636 1383 640 1387
rect 644 1384 648 1388
rect 656 1384 660 1388
rect 690 1378 694 1382
rect 730 1384 734 1388
rect 719 1377 723 1381
rect 497 1367 501 1371
rect 429 1363 435 1367
rect 522 1364 526 1368
rect 529 1367 533 1371
rect 547 1367 551 1371
rect 569 1364 573 1368
rect 594 1364 598 1368
rect 604 1367 608 1371
rect 620 1367 624 1371
rect 640 1364 644 1368
rect 647 1367 651 1371
rect 785 1383 789 1387
rect 805 1386 809 1390
rect 824 1382 828 1386
rect 953 1393 957 1397
rect 966 1396 970 1402
rect 1003 1396 1007 1402
rect 1016 1398 1020 1402
rect 1040 1402 1044 1406
rect 1114 1402 1118 1406
rect 1024 1396 1028 1402
rect 1061 1396 1065 1402
rect 1077 1396 1081 1402
rect 1098 1396 1102 1402
rect 1135 1396 1139 1402
rect 1148 1398 1152 1402
rect 1172 1402 1176 1406
rect 1246 1402 1250 1406
rect 1156 1396 1160 1402
rect 1193 1396 1197 1402
rect 1209 1396 1213 1402
rect 1230 1396 1234 1402
rect 1267 1396 1271 1402
rect 1280 1398 1284 1402
rect 1304 1402 1308 1406
rect 1374 1409 1380 1413
rect 1444 1409 1448 1413
rect 1453 1409 1457 1413
rect 1503 1409 1507 1413
rect 1528 1409 1532 1413
rect 1559 1409 1563 1413
rect 1288 1396 1292 1402
rect 1325 1396 1329 1402
rect 1341 1398 1345 1402
rect 1444 1401 1448 1405
rect 1487 1402 1491 1406
rect 1509 1401 1516 1405
rect 1559 1402 1563 1406
rect 1430 1397 1434 1401
rect 1462 1397 1466 1401
rect 1480 1397 1484 1401
rect 1537 1397 1541 1401
rect 1552 1397 1556 1401
rect 1580 1397 1584 1401
rect 843 1383 847 1387
rect 862 1383 866 1387
rect 875 1384 879 1388
rect 897 1383 901 1387
rect 905 1384 909 1388
rect 917 1384 921 1388
rect 966 1383 970 1387
rect 982 1383 986 1389
rect 1016 1389 1020 1393
rect 1003 1383 1007 1387
rect 1024 1383 1028 1387
rect 1040 1383 1044 1389
rect 1061 1383 1065 1387
rect 1077 1383 1081 1387
rect 1098 1383 1102 1387
rect 1114 1383 1118 1389
rect 1148 1389 1152 1393
rect 1135 1383 1139 1387
rect 1156 1383 1160 1387
rect 1172 1383 1176 1389
rect 1193 1383 1197 1387
rect 1209 1383 1213 1387
rect 1230 1383 1234 1387
rect 1246 1383 1250 1389
rect 1280 1389 1284 1393
rect 1267 1383 1271 1387
rect 1288 1383 1292 1387
rect 1304 1383 1308 1389
rect 1325 1383 1329 1387
rect 1341 1383 1345 1387
rect 1425 1385 1429 1389
rect 731 1367 735 1371
rect 757 1367 761 1371
rect 26 1356 30 1360
rect 77 1356 81 1360
rect 127 1356 131 1360
rect 158 1356 162 1360
rect 209 1356 213 1360
rect 259 1356 263 1360
rect 290 1356 294 1360
rect 341 1356 345 1360
rect 391 1356 395 1360
rect 465 1357 471 1361
rect 505 1357 509 1361
rect 523 1357 527 1361
rect 554 1357 558 1361
rect 576 1357 580 1361
rect 641 1357 645 1361
rect 783 1364 787 1368
rect 790 1367 794 1371
rect 808 1367 812 1371
rect 830 1364 834 1368
rect 855 1364 859 1368
rect 865 1367 869 1371
rect 881 1367 885 1371
rect 901 1364 905 1368
rect 908 1367 912 1371
rect 959 1372 963 1376
rect 996 1370 1000 1374
rect 1016 1370 1020 1374
rect 1060 1370 1064 1374
rect 1091 1372 1095 1376
rect 1128 1370 1132 1374
rect 1148 1370 1152 1374
rect 1192 1370 1196 1374
rect 1223 1372 1227 1376
rect 1260 1370 1264 1374
rect 1280 1370 1284 1374
rect 1324 1370 1328 1374
rect 1457 1383 1461 1387
rect 1477 1386 1481 1390
rect 1496 1382 1500 1386
rect 1515 1383 1519 1387
rect 1534 1383 1538 1387
rect 1547 1384 1551 1388
rect 1683 1409 1687 1413
rect 1705 1409 1709 1413
rect 1764 1409 1768 1413
rect 1789 1409 1793 1413
rect 1820 1409 1824 1413
rect 1705 1401 1709 1405
rect 1748 1402 1752 1406
rect 1770 1401 1777 1405
rect 1820 1402 1824 1406
rect 1723 1397 1727 1401
rect 1741 1397 1745 1401
rect 1798 1397 1802 1401
rect 1813 1397 1817 1401
rect 1841 1397 1845 1401
rect 1644 1393 1648 1397
rect 1569 1383 1573 1387
rect 1577 1384 1581 1388
rect 1589 1384 1593 1388
rect 1623 1378 1627 1382
rect 1663 1384 1667 1388
rect 1652 1377 1656 1381
rect 1430 1367 1434 1371
rect 1362 1363 1368 1367
rect 1455 1364 1459 1368
rect 1462 1367 1466 1371
rect 1480 1367 1484 1371
rect 1502 1364 1506 1368
rect 1527 1364 1531 1368
rect 1537 1367 1541 1371
rect 1553 1367 1557 1371
rect 1573 1364 1577 1368
rect 1580 1367 1584 1371
rect 1718 1383 1722 1387
rect 1738 1386 1742 1390
rect 1757 1382 1761 1386
rect 1776 1383 1780 1387
rect 1795 1383 1799 1387
rect 1808 1384 1812 1388
rect 1830 1383 1834 1387
rect 1838 1384 1842 1388
rect 1850 1384 1854 1388
rect 1664 1367 1668 1371
rect 1690 1367 1694 1371
rect 701 1357 705 1361
rect 740 1357 744 1361
rect 784 1357 788 1361
rect 815 1357 819 1361
rect 837 1357 841 1361
rect 902 1357 906 1361
rect 959 1356 963 1360
rect 1010 1356 1014 1360
rect 1060 1356 1064 1360
rect 1091 1356 1095 1360
rect 1142 1356 1146 1360
rect 1192 1356 1196 1360
rect 1223 1356 1227 1360
rect 1274 1356 1278 1360
rect 1324 1356 1328 1360
rect 1398 1357 1404 1361
rect 1438 1357 1442 1361
rect 1456 1357 1460 1361
rect 1487 1357 1491 1361
rect 1509 1357 1513 1361
rect 1574 1357 1578 1361
rect 1716 1364 1720 1368
rect 1723 1367 1727 1371
rect 1741 1367 1745 1371
rect 1763 1364 1767 1368
rect 1788 1364 1792 1368
rect 1798 1367 1802 1371
rect 1814 1367 1818 1371
rect 1834 1364 1838 1368
rect 1841 1367 1845 1371
rect 1634 1357 1638 1361
rect 1673 1357 1677 1361
rect 1717 1357 1721 1361
rect 1748 1357 1752 1361
rect 1770 1357 1774 1361
rect 1835 1357 1839 1361
rect 20 1349 24 1353
rect 408 1349 412 1353
rect 417 1350 423 1354
rect 496 1350 500 1354
rect 530 1350 534 1354
rect 547 1350 551 1354
rect 603 1350 607 1354
rect 620 1350 624 1354
rect 648 1350 652 1354
rect 731 1350 735 1354
rect 757 1350 761 1354
rect 791 1350 795 1354
rect 808 1350 812 1354
rect 864 1350 868 1354
rect 881 1350 885 1354
rect 909 1350 913 1354
rect 953 1349 957 1353
rect 1341 1349 1345 1353
rect 1350 1350 1356 1354
rect 1429 1350 1433 1354
rect 1463 1350 1467 1354
rect 1480 1350 1484 1354
rect 1536 1350 1540 1354
rect 1553 1350 1557 1354
rect 1581 1350 1585 1354
rect 1664 1350 1668 1354
rect 1690 1350 1694 1354
rect 1724 1350 1728 1354
rect 1741 1350 1745 1354
rect 1797 1350 1801 1354
rect 1814 1350 1818 1354
rect 1842 1350 1846 1354
rect 143 1342 148 1346
rect 276 1342 280 1346
rect 453 1343 459 1347
rect 505 1343 509 1347
rect 739 1343 743 1347
rect 925 1344 929 1348
rect 937 1344 941 1348
rect 1076 1342 1081 1346
rect 1209 1342 1213 1346
rect 1386 1343 1392 1347
rect 1438 1343 1442 1347
rect 1672 1343 1676 1347
rect 1858 1344 1862 1348
rect 1870 1344 1874 1348
rect 151 1335 155 1339
rect 441 1335 447 1339
rect 749 1336 753 1340
rect 914 1336 918 1340
rect 135 1331 139 1335
rect 167 1331 171 1335
rect 1084 1335 1088 1339
rect 1374 1335 1380 1339
rect 1682 1336 1686 1340
rect 1847 1336 1851 1340
rect 1068 1331 1072 1335
rect 1100 1331 1104 1335
rect 135 1324 139 1328
rect 167 1324 171 1328
rect 1068 1324 1072 1328
rect 1100 1324 1104 1328
rect 151 1317 155 1321
rect 408 1317 412 1321
rect 477 1317 483 1321
rect 797 1317 801 1321
rect 833 1317 837 1321
rect 900 1317 904 1321
rect 1084 1317 1088 1321
rect 1341 1317 1345 1321
rect 1410 1317 1416 1321
rect 1730 1317 1734 1321
rect 1766 1317 1770 1321
rect 1833 1317 1837 1321
rect 408 1309 412 1313
rect 417 1310 423 1314
rect 783 1310 787 1314
rect 135 1305 139 1309
rect 167 1305 171 1309
rect 151 1301 155 1305
rect 797 1303 801 1307
rect 847 1303 851 1307
rect 900 1303 904 1307
rect 1341 1309 1345 1313
rect 1350 1310 1356 1314
rect 1716 1310 1720 1314
rect 1068 1305 1072 1309
rect 1100 1305 1104 1309
rect 1084 1301 1088 1305
rect 1730 1303 1734 1307
rect 1780 1303 1784 1307
rect 1833 1303 1837 1307
rect 143 1294 148 1298
rect 277 1294 281 1298
rect 820 1292 824 1296
rect 26 1287 30 1291
rect 62 1287 66 1291
rect 129 1287 133 1291
rect 158 1287 162 1291
rect 194 1287 198 1291
rect 261 1287 265 1291
rect 290 1287 294 1291
rect 326 1287 330 1291
rect 393 1287 397 1291
rect 477 1287 483 1291
rect 417 1280 423 1284
rect 791 1283 795 1287
rect 804 1286 808 1292
rect 841 1286 845 1292
rect 854 1288 858 1292
rect 878 1292 882 1296
rect 1076 1294 1081 1298
rect 1210 1294 1214 1298
rect 1753 1292 1757 1296
rect 862 1286 866 1292
rect 899 1286 903 1292
rect 915 1286 919 1292
rect 959 1287 963 1291
rect 995 1287 999 1291
rect 1062 1287 1066 1291
rect 1091 1287 1095 1291
rect 1127 1287 1131 1291
rect 1194 1287 1198 1291
rect 1223 1287 1227 1291
rect 1259 1287 1263 1291
rect 1326 1287 1330 1291
rect 1410 1287 1416 1291
rect 26 1273 30 1277
rect 76 1273 80 1277
rect 129 1273 133 1277
rect 158 1273 162 1277
rect 208 1273 212 1277
rect 261 1273 265 1277
rect 290 1273 294 1277
rect 340 1273 344 1277
rect 393 1273 397 1277
rect 804 1273 808 1277
rect 820 1273 824 1279
rect 854 1279 858 1283
rect 841 1273 845 1277
rect 49 1262 53 1266
rect 20 1253 24 1257
rect 33 1256 37 1262
rect 70 1256 74 1262
rect 83 1258 87 1262
rect 107 1262 111 1266
rect 181 1262 185 1266
rect 91 1256 95 1262
rect 128 1256 132 1262
rect 144 1256 148 1262
rect 165 1256 169 1262
rect 202 1256 206 1262
rect 215 1258 219 1262
rect 239 1262 243 1266
rect 313 1262 317 1266
rect 223 1256 227 1262
rect 260 1256 264 1262
rect 276 1256 280 1262
rect 297 1256 301 1262
rect 334 1256 338 1262
rect 347 1258 351 1262
rect 371 1262 375 1266
rect 355 1256 359 1262
rect 392 1256 396 1262
rect 408 1258 412 1262
rect 862 1273 866 1277
rect 878 1273 882 1279
rect 1350 1280 1356 1284
rect 1724 1283 1728 1287
rect 1737 1286 1741 1292
rect 1774 1286 1778 1292
rect 1787 1288 1791 1292
rect 1811 1292 1815 1296
rect 1795 1286 1799 1292
rect 1832 1286 1836 1292
rect 1848 1286 1852 1292
rect 899 1273 903 1277
rect 915 1273 919 1277
rect 959 1273 963 1277
rect 1009 1273 1013 1277
rect 1062 1273 1066 1277
rect 1091 1273 1095 1277
rect 1141 1273 1145 1277
rect 1194 1273 1198 1277
rect 1223 1273 1227 1277
rect 1273 1273 1277 1277
rect 1326 1273 1330 1277
rect 1737 1273 1741 1277
rect 1753 1273 1757 1279
rect 1787 1279 1791 1283
rect 1774 1273 1778 1277
rect 797 1262 801 1266
rect 834 1260 838 1264
rect 854 1260 858 1264
rect 898 1260 902 1264
rect 982 1262 986 1266
rect 33 1243 37 1247
rect 49 1243 53 1249
rect 83 1249 87 1253
rect 70 1243 74 1247
rect 91 1243 95 1247
rect 107 1243 111 1249
rect 128 1243 132 1247
rect 144 1243 148 1247
rect 165 1243 169 1247
rect 181 1243 185 1249
rect 215 1249 219 1253
rect 202 1243 206 1247
rect 223 1243 227 1247
rect 239 1243 243 1249
rect 260 1243 264 1247
rect 276 1243 280 1247
rect 297 1243 301 1247
rect 313 1243 317 1249
rect 347 1249 351 1253
rect 334 1243 338 1247
rect 355 1243 359 1247
rect 371 1243 375 1249
rect 429 1253 435 1257
rect 953 1253 957 1257
rect 966 1256 970 1262
rect 1003 1256 1007 1262
rect 1016 1258 1020 1262
rect 1040 1262 1044 1266
rect 1114 1262 1118 1266
rect 1024 1256 1028 1262
rect 1061 1256 1065 1262
rect 1077 1256 1081 1262
rect 1098 1256 1102 1262
rect 1135 1256 1139 1262
rect 1148 1258 1152 1262
rect 1172 1262 1176 1266
rect 1246 1262 1250 1266
rect 1156 1256 1160 1262
rect 1193 1256 1197 1262
rect 1209 1256 1213 1262
rect 1230 1256 1234 1262
rect 1267 1256 1271 1262
rect 1280 1258 1284 1262
rect 1304 1262 1308 1266
rect 1288 1256 1292 1262
rect 1325 1256 1329 1262
rect 1341 1258 1345 1262
rect 1795 1273 1799 1277
rect 1811 1273 1815 1279
rect 1832 1273 1836 1277
rect 1848 1273 1852 1277
rect 1730 1262 1734 1266
rect 1767 1260 1771 1264
rect 1787 1260 1791 1264
rect 1831 1260 1835 1264
rect 392 1243 396 1247
rect 408 1243 412 1247
rect 465 1246 471 1250
rect 797 1246 801 1250
rect 848 1246 852 1250
rect 898 1246 902 1250
rect 966 1243 970 1247
rect 982 1243 986 1249
rect 1016 1249 1020 1253
rect 1003 1243 1007 1247
rect 26 1232 30 1236
rect 63 1230 67 1234
rect 83 1230 87 1234
rect 127 1230 131 1234
rect 158 1232 162 1236
rect 195 1230 199 1234
rect 215 1230 219 1234
rect 259 1230 263 1234
rect 290 1232 294 1236
rect 327 1230 331 1234
rect 347 1230 351 1234
rect 391 1230 395 1234
rect 790 1238 794 1242
rect 915 1239 919 1243
rect 1024 1243 1028 1247
rect 1040 1243 1044 1249
rect 1061 1243 1065 1247
rect 1077 1243 1081 1247
rect 1098 1243 1102 1247
rect 1114 1243 1118 1249
rect 1148 1249 1152 1253
rect 1135 1243 1139 1247
rect 1156 1243 1160 1247
rect 1172 1243 1176 1249
rect 1193 1243 1197 1247
rect 1209 1243 1213 1247
rect 1230 1243 1234 1247
rect 1246 1243 1250 1249
rect 1280 1249 1284 1253
rect 1267 1243 1271 1247
rect 1288 1243 1292 1247
rect 1304 1243 1308 1249
rect 1362 1253 1368 1257
rect 1325 1243 1329 1247
rect 1341 1243 1345 1247
rect 1398 1246 1404 1250
rect 1730 1246 1734 1250
rect 1781 1246 1785 1250
rect 1831 1246 1835 1250
rect 477 1231 483 1235
rect 797 1231 801 1235
rect 833 1231 837 1235
rect 900 1231 904 1235
rect 429 1223 435 1227
rect 783 1224 787 1228
rect 959 1232 963 1236
rect 996 1230 1000 1234
rect 1016 1230 1020 1234
rect 1060 1230 1064 1234
rect 1091 1232 1095 1236
rect 1128 1230 1132 1234
rect 1148 1230 1152 1234
rect 1192 1230 1196 1234
rect 1223 1232 1227 1236
rect 1260 1230 1264 1234
rect 1280 1230 1284 1234
rect 1324 1230 1328 1234
rect 1723 1238 1727 1242
rect 1848 1239 1852 1243
rect 1410 1231 1416 1235
rect 1730 1231 1734 1235
rect 1766 1231 1770 1235
rect 1833 1231 1837 1235
rect 26 1216 30 1220
rect 77 1216 81 1220
rect 127 1216 131 1220
rect 158 1216 162 1220
rect 209 1216 213 1220
rect 259 1216 263 1220
rect 290 1216 294 1220
rect 341 1216 345 1220
rect 391 1216 395 1220
rect 465 1216 471 1220
rect 797 1217 801 1221
rect 847 1217 851 1221
rect 900 1217 904 1221
rect 1362 1223 1368 1227
rect 1716 1224 1720 1228
rect 959 1216 963 1220
rect 1010 1216 1014 1220
rect 1060 1216 1064 1220
rect 1091 1216 1095 1220
rect 1142 1216 1146 1220
rect 1192 1216 1196 1220
rect 1223 1216 1227 1220
rect 1274 1216 1278 1220
rect 1324 1216 1328 1220
rect 1398 1216 1404 1220
rect 1730 1217 1734 1221
rect 1780 1217 1784 1221
rect 1833 1217 1837 1221
rect 19 1209 23 1213
rect 408 1209 412 1213
rect 820 1206 824 1210
rect 26 1201 30 1205
rect 62 1201 66 1205
rect 129 1201 133 1205
rect 158 1201 162 1205
rect 194 1201 198 1205
rect 261 1201 265 1205
rect 290 1201 294 1205
rect 326 1201 330 1205
rect 393 1201 397 1205
rect 477 1201 483 1205
rect 417 1194 423 1198
rect 791 1197 795 1201
rect 804 1200 808 1206
rect 841 1200 845 1206
rect 854 1202 858 1206
rect 878 1206 882 1210
rect 952 1209 956 1213
rect 1341 1209 1345 1213
rect 1753 1206 1757 1210
rect 862 1200 866 1206
rect 899 1200 903 1206
rect 915 1202 919 1206
rect 937 1200 941 1204
rect 959 1201 963 1205
rect 995 1201 999 1205
rect 1062 1201 1066 1205
rect 1091 1201 1095 1205
rect 1127 1201 1131 1205
rect 1194 1201 1198 1205
rect 1223 1201 1227 1205
rect 1259 1201 1263 1205
rect 1326 1201 1330 1205
rect 1410 1201 1416 1205
rect 26 1187 30 1191
rect 76 1187 80 1191
rect 129 1187 133 1191
rect 158 1187 162 1191
rect 208 1187 212 1191
rect 261 1187 265 1191
rect 290 1187 294 1191
rect 340 1187 344 1191
rect 393 1187 397 1191
rect 804 1187 808 1191
rect 820 1187 824 1193
rect 854 1193 858 1197
rect 841 1187 845 1191
rect 49 1176 53 1180
rect 20 1167 24 1171
rect 33 1170 37 1176
rect 70 1170 74 1176
rect 83 1172 87 1176
rect 107 1176 111 1180
rect 181 1176 185 1180
rect 91 1170 95 1176
rect 128 1170 132 1176
rect 144 1170 148 1176
rect 165 1170 169 1176
rect 202 1170 206 1176
rect 215 1172 219 1176
rect 239 1176 243 1180
rect 313 1176 317 1180
rect 223 1170 227 1176
rect 260 1170 264 1176
rect 276 1170 280 1176
rect 297 1170 301 1176
rect 334 1170 338 1176
rect 347 1172 351 1176
rect 371 1176 375 1180
rect 355 1170 359 1176
rect 392 1170 396 1176
rect 408 1172 412 1176
rect 862 1187 866 1191
rect 878 1187 882 1193
rect 899 1187 903 1191
rect 915 1187 919 1196
rect 1350 1194 1356 1198
rect 1724 1197 1728 1201
rect 1737 1200 1741 1206
rect 1774 1200 1778 1206
rect 1787 1202 1791 1206
rect 1811 1206 1815 1210
rect 1795 1200 1799 1206
rect 1832 1200 1836 1206
rect 1848 1202 1852 1206
rect 1870 1200 1874 1204
rect 937 1184 941 1188
rect 959 1187 963 1191
rect 1009 1187 1013 1191
rect 1062 1187 1066 1191
rect 1091 1187 1095 1191
rect 1141 1187 1145 1191
rect 1194 1187 1198 1191
rect 1223 1187 1227 1191
rect 1273 1187 1277 1191
rect 1326 1187 1330 1191
rect 1737 1187 1741 1191
rect 1753 1187 1757 1193
rect 1787 1193 1791 1197
rect 1774 1187 1778 1191
rect 797 1176 801 1180
rect 834 1174 838 1178
rect 854 1174 858 1178
rect 898 1174 902 1178
rect 982 1176 986 1180
rect 33 1157 37 1161
rect 49 1157 53 1163
rect 83 1163 87 1167
rect 70 1157 74 1161
rect 91 1157 95 1161
rect 107 1157 111 1163
rect 128 1157 132 1161
rect 144 1157 148 1161
rect 165 1157 169 1161
rect 181 1157 185 1163
rect 215 1163 219 1167
rect 202 1157 206 1161
rect 223 1157 227 1161
rect 239 1157 243 1163
rect 260 1157 264 1161
rect 276 1157 280 1161
rect 297 1157 301 1161
rect 313 1157 317 1163
rect 347 1163 351 1167
rect 334 1157 338 1161
rect 355 1157 359 1161
rect 371 1157 375 1163
rect 429 1167 435 1171
rect 953 1167 957 1171
rect 966 1170 970 1176
rect 1003 1170 1007 1176
rect 1016 1172 1020 1176
rect 1040 1176 1044 1180
rect 1114 1176 1118 1180
rect 1024 1170 1028 1176
rect 1061 1170 1065 1176
rect 1077 1170 1081 1176
rect 1098 1170 1102 1176
rect 1135 1170 1139 1176
rect 1148 1172 1152 1176
rect 1172 1176 1176 1180
rect 1246 1176 1250 1180
rect 1156 1170 1160 1176
rect 1193 1170 1197 1176
rect 1209 1170 1213 1176
rect 1230 1170 1234 1176
rect 1267 1170 1271 1176
rect 1280 1172 1284 1176
rect 1304 1176 1308 1180
rect 1288 1170 1292 1176
rect 1325 1170 1329 1176
rect 1341 1172 1345 1176
rect 1795 1187 1799 1191
rect 1811 1187 1815 1193
rect 1832 1187 1836 1191
rect 1848 1187 1852 1196
rect 1870 1184 1874 1188
rect 1730 1176 1734 1180
rect 1767 1174 1771 1178
rect 1787 1174 1791 1178
rect 1831 1174 1835 1178
rect 392 1157 396 1161
rect 408 1157 412 1161
rect 465 1160 471 1164
rect 797 1160 801 1164
rect 848 1160 852 1164
rect 898 1160 902 1164
rect 966 1157 970 1161
rect 982 1157 986 1163
rect 1016 1163 1020 1167
rect 1003 1157 1007 1161
rect 1024 1157 1028 1161
rect 1040 1157 1044 1163
rect 1061 1157 1065 1161
rect 1077 1157 1081 1161
rect 1098 1157 1102 1161
rect 1114 1157 1118 1163
rect 1148 1163 1152 1167
rect 1135 1157 1139 1161
rect 1156 1157 1160 1161
rect 1172 1157 1176 1163
rect 1193 1157 1197 1161
rect 1209 1157 1213 1161
rect 1230 1157 1234 1161
rect 1246 1157 1250 1163
rect 1280 1163 1284 1167
rect 1267 1157 1271 1161
rect 1288 1157 1292 1161
rect 1304 1157 1308 1163
rect 1362 1167 1368 1171
rect 1325 1157 1329 1161
rect 1341 1157 1345 1161
rect 1398 1160 1404 1164
rect 1730 1160 1734 1164
rect 1781 1160 1785 1164
rect 1831 1160 1835 1164
rect 26 1146 30 1150
rect 63 1144 67 1148
rect 83 1144 87 1148
rect 127 1144 131 1148
rect 158 1146 162 1150
rect 195 1144 199 1148
rect 215 1144 219 1148
rect 259 1144 263 1148
rect 290 1146 294 1150
rect 327 1144 331 1148
rect 347 1144 351 1148
rect 391 1144 395 1148
rect 959 1146 963 1150
rect 996 1144 1000 1148
rect 1016 1144 1020 1148
rect 1060 1144 1064 1148
rect 1091 1146 1095 1150
rect 1128 1144 1132 1148
rect 1148 1144 1152 1148
rect 1192 1144 1196 1148
rect 1223 1146 1227 1150
rect 1260 1144 1264 1148
rect 1280 1144 1284 1148
rect 1324 1144 1328 1148
rect 429 1137 435 1141
rect 1362 1137 1368 1141
rect 26 1130 30 1134
rect 77 1130 81 1134
rect 127 1130 131 1134
rect 158 1130 162 1134
rect 209 1130 213 1134
rect 259 1130 263 1134
rect 290 1130 294 1134
rect 341 1130 345 1134
rect 391 1130 395 1134
rect 465 1130 471 1134
rect 959 1130 963 1134
rect 1010 1130 1014 1134
rect 1060 1130 1064 1134
rect 1091 1130 1095 1134
rect 1142 1130 1146 1134
rect 1192 1130 1196 1134
rect 1223 1130 1227 1134
rect 1274 1130 1278 1134
rect 1324 1130 1328 1134
rect 1398 1130 1404 1134
rect 19 1123 23 1127
rect 408 1123 412 1127
rect 952 1123 956 1127
rect 1341 1123 1345 1127
rect 144 1116 148 1120
rect 252 1116 256 1120
rect 276 1116 280 1120
rect 1077 1116 1081 1120
rect 1185 1116 1189 1120
rect 1209 1116 1213 1120
rect 268 1109 272 1113
rect 252 1105 256 1109
rect 284 1105 288 1109
rect 1201 1109 1205 1113
rect 1185 1105 1189 1109
rect 1217 1105 1221 1109
rect 252 1098 256 1102
rect 284 1098 288 1102
rect 937 1098 941 1102
rect 1185 1098 1189 1102
rect 1217 1098 1221 1102
rect 1870 1098 1874 1102
rect 268 1091 272 1095
rect 408 1091 412 1095
rect 1201 1091 1205 1095
rect 1341 1091 1345 1095
rect 408 1083 412 1087
rect 1341 1083 1345 1087
rect 252 1079 256 1083
rect 284 1079 288 1083
rect 268 1075 272 1079
rect 1185 1079 1189 1083
rect 1217 1079 1221 1083
rect 1201 1075 1205 1079
rect 144 1068 148 1072
rect 252 1068 256 1072
rect 276 1068 280 1072
rect 1077 1068 1081 1072
rect 1185 1068 1189 1072
rect 1209 1068 1213 1072
rect 26 1061 30 1065
rect 62 1061 66 1065
rect 129 1061 133 1065
rect 158 1061 162 1065
rect 194 1061 198 1065
rect 261 1061 265 1065
rect 290 1061 294 1065
rect 326 1061 330 1065
rect 393 1061 397 1065
rect 477 1061 483 1065
rect 959 1061 963 1065
rect 995 1061 999 1065
rect 1062 1061 1066 1065
rect 1091 1061 1095 1065
rect 1127 1061 1131 1065
rect 1194 1061 1198 1065
rect 1223 1061 1227 1065
rect 1259 1061 1263 1065
rect 1326 1061 1330 1065
rect 1410 1061 1416 1065
rect 417 1054 423 1058
rect 1350 1054 1356 1058
rect 26 1047 30 1051
rect 76 1047 80 1051
rect 129 1047 133 1051
rect 158 1047 162 1051
rect 208 1047 212 1051
rect 261 1047 265 1051
rect 290 1047 294 1051
rect 340 1047 344 1051
rect 393 1047 397 1051
rect 959 1047 963 1051
rect 1009 1047 1013 1051
rect 1062 1047 1066 1051
rect 1091 1047 1095 1051
rect 1141 1047 1145 1051
rect 1194 1047 1198 1051
rect 1223 1047 1227 1051
rect 1273 1047 1277 1051
rect 1326 1047 1330 1051
rect 49 1036 53 1040
rect 20 1027 24 1031
rect 33 1030 37 1036
rect 70 1030 74 1036
rect 83 1032 87 1036
rect 107 1036 111 1040
rect 181 1036 185 1040
rect 91 1030 95 1036
rect 128 1030 132 1036
rect 144 1030 148 1036
rect 165 1030 169 1036
rect 202 1030 206 1036
rect 215 1032 219 1036
rect 239 1036 243 1040
rect 313 1036 317 1040
rect 223 1030 227 1036
rect 260 1030 264 1036
rect 276 1030 280 1036
rect 297 1030 301 1036
rect 334 1030 338 1036
rect 347 1032 351 1036
rect 371 1036 375 1040
rect 982 1036 986 1040
rect 355 1030 359 1036
rect 392 1030 396 1036
rect 408 1032 412 1036
rect 33 1017 37 1021
rect 49 1017 53 1023
rect 83 1023 87 1027
rect 70 1017 74 1021
rect 91 1017 95 1021
rect 107 1017 111 1023
rect 128 1017 132 1021
rect 144 1017 148 1021
rect 165 1017 169 1021
rect 181 1017 185 1023
rect 215 1023 219 1027
rect 202 1017 206 1021
rect 223 1017 227 1021
rect 239 1017 243 1023
rect 260 1017 264 1021
rect 276 1017 280 1021
rect 297 1017 301 1021
rect 313 1017 317 1023
rect 347 1023 351 1027
rect 334 1017 338 1021
rect 355 1017 359 1021
rect 371 1017 375 1023
rect 953 1027 957 1031
rect 966 1030 970 1036
rect 1003 1030 1007 1036
rect 1016 1032 1020 1036
rect 1040 1036 1044 1040
rect 1114 1036 1118 1040
rect 1024 1030 1028 1036
rect 1061 1030 1065 1036
rect 1077 1030 1081 1036
rect 1098 1030 1102 1036
rect 1135 1030 1139 1036
rect 1148 1032 1152 1036
rect 1172 1036 1176 1040
rect 1246 1036 1250 1040
rect 1156 1030 1160 1036
rect 1193 1030 1197 1036
rect 1209 1030 1213 1036
rect 1230 1030 1234 1036
rect 1267 1030 1271 1036
rect 1280 1032 1284 1036
rect 1304 1036 1308 1040
rect 1288 1030 1292 1036
rect 1325 1030 1329 1036
rect 1341 1032 1345 1036
rect 392 1017 396 1021
rect 408 1017 412 1021
rect 966 1017 970 1021
rect 982 1017 986 1023
rect 1016 1023 1020 1027
rect 1003 1017 1007 1021
rect 1024 1017 1028 1021
rect 1040 1017 1044 1023
rect 1061 1017 1065 1021
rect 1077 1017 1081 1021
rect 1098 1017 1102 1021
rect 1114 1017 1118 1023
rect 1148 1023 1152 1027
rect 1135 1017 1139 1021
rect 1156 1017 1160 1021
rect 1172 1017 1176 1023
rect 1193 1017 1197 1021
rect 1209 1017 1213 1021
rect 1230 1017 1234 1021
rect 1246 1017 1250 1023
rect 1280 1023 1284 1027
rect 1267 1017 1271 1021
rect 1288 1017 1292 1021
rect 1304 1017 1308 1023
rect 1325 1017 1329 1021
rect 1341 1017 1345 1021
rect 26 1006 30 1010
rect 63 1004 67 1008
rect 83 1004 87 1008
rect 127 1004 131 1008
rect 158 1006 162 1010
rect 195 1004 199 1008
rect 215 1004 219 1008
rect 259 1004 263 1008
rect 290 1006 294 1010
rect 327 1004 331 1008
rect 347 1004 351 1008
rect 391 1004 395 1008
rect 959 1006 963 1010
rect 996 1004 1000 1008
rect 1016 1004 1020 1008
rect 1060 1004 1064 1008
rect 1091 1006 1095 1010
rect 1128 1004 1132 1008
rect 1148 1004 1152 1008
rect 1192 1004 1196 1008
rect 1223 1006 1227 1010
rect 1260 1004 1264 1008
rect 1280 1004 1284 1008
rect 1324 1004 1328 1008
rect 429 997 435 1001
rect 1362 997 1368 1001
rect 26 990 30 994
rect 77 990 81 994
rect 127 990 131 994
rect 158 990 162 994
rect 209 990 213 994
rect 259 990 263 994
rect 290 990 294 994
rect 341 990 345 994
rect 391 990 395 994
rect 465 990 471 994
rect 959 990 963 994
rect 1010 990 1014 994
rect 1060 990 1064 994
rect 1091 990 1095 994
rect 1142 990 1146 994
rect 1192 990 1196 994
rect 1223 990 1227 994
rect 1274 990 1278 994
rect 1324 990 1328 994
rect 1398 990 1404 994
rect 477 982 483 986
rect 498 982 502 986
rect 534 982 538 986
rect 601 982 605 986
rect 630 982 634 986
rect 666 982 670 986
rect 733 982 737 986
rect 762 982 766 986
rect 798 982 802 986
rect 865 982 869 986
rect 894 982 898 986
rect 930 982 934 986
rect 997 982 1001 986
rect 1410 982 1416 986
rect 1431 982 1435 986
rect 1467 982 1471 986
rect 1534 982 1538 986
rect 1563 982 1567 986
rect 1599 982 1603 986
rect 1666 982 1670 986
rect 1695 982 1699 986
rect 1731 982 1735 986
rect 1798 982 1802 986
rect 1827 982 1831 986
rect 1863 982 1867 986
rect 1930 982 1934 986
rect 417 975 423 979
rect 1350 975 1356 979
rect 498 968 502 972
rect 548 968 552 972
rect 601 968 605 972
rect 630 968 634 972
rect 680 968 684 972
rect 733 968 737 972
rect 762 968 766 972
rect 812 968 816 972
rect 865 968 869 972
rect 894 968 898 972
rect 944 968 948 972
rect 997 968 1001 972
rect 1431 968 1435 972
rect 1481 968 1485 972
rect 1534 968 1538 972
rect 1563 968 1567 972
rect 1613 968 1617 972
rect 1666 968 1670 972
rect 1695 968 1699 972
rect 1745 968 1749 972
rect 1798 968 1802 972
rect 1827 968 1831 972
rect 1877 968 1881 972
rect 1930 968 1934 972
rect 521 957 525 961
rect 158 949 162 953
rect 194 949 198 953
rect 261 949 265 953
rect 477 949 483 953
rect 492 948 496 952
rect 505 951 509 957
rect 542 951 546 957
rect 555 953 559 957
rect 579 957 583 961
rect 653 957 657 961
rect 563 951 567 957
rect 600 951 604 957
rect 616 953 620 957
rect 417 942 423 946
rect 158 935 162 939
rect 208 935 212 939
rect 261 935 265 939
rect 505 938 509 942
rect 521 938 525 944
rect 555 944 559 948
rect 542 938 546 942
rect 563 938 567 942
rect 579 938 583 944
rect 624 948 628 952
rect 637 951 641 957
rect 674 951 678 957
rect 687 953 691 957
rect 711 957 715 961
rect 785 957 789 961
rect 695 951 699 957
rect 732 951 736 957
rect 748 953 752 957
rect 600 938 604 942
rect 616 938 620 942
rect 637 938 641 942
rect 653 938 657 944
rect 687 944 691 948
rect 674 938 678 942
rect 695 938 699 942
rect 711 938 715 944
rect 756 948 760 952
rect 769 951 773 957
rect 806 951 810 957
rect 819 953 823 957
rect 843 957 847 961
rect 917 957 921 961
rect 827 951 831 957
rect 864 951 868 957
rect 880 953 884 957
rect 732 938 736 942
rect 748 938 752 942
rect 769 938 773 942
rect 785 938 789 944
rect 819 944 823 948
rect 806 938 810 942
rect 827 938 831 942
rect 843 938 847 944
rect 888 948 892 952
rect 901 951 905 957
rect 938 951 942 957
rect 951 953 955 957
rect 975 957 979 961
rect 1454 957 1458 961
rect 959 951 963 957
rect 996 951 1000 957
rect 1012 953 1016 957
rect 1091 949 1095 953
rect 1127 949 1131 953
rect 1194 949 1198 953
rect 1410 949 1416 953
rect 864 938 868 942
rect 880 938 884 942
rect 901 938 905 942
rect 917 938 921 944
rect 951 944 955 948
rect 938 938 942 942
rect 181 924 185 928
rect 143 915 147 919
rect 165 918 169 924
rect 202 918 206 924
rect 215 920 219 924
rect 239 924 243 928
rect 223 918 227 924
rect 260 918 264 924
rect 276 918 280 924
rect 498 927 502 931
rect 535 925 539 929
rect 555 925 559 929
rect 599 925 603 929
rect 630 927 634 931
rect 667 925 671 929
rect 687 925 691 929
rect 731 925 735 929
rect 762 927 766 931
rect 799 925 803 929
rect 819 925 823 929
rect 863 925 867 929
rect 880 930 884 934
rect 959 938 963 942
rect 975 938 979 944
rect 1425 948 1429 952
rect 1438 951 1442 957
rect 1475 951 1479 957
rect 1488 953 1492 957
rect 1512 957 1516 961
rect 1586 957 1590 961
rect 1496 951 1500 957
rect 1533 951 1537 957
rect 1549 953 1553 957
rect 1350 942 1356 946
rect 996 938 1000 942
rect 1012 938 1016 942
rect 894 927 898 931
rect 931 925 935 929
rect 951 925 955 929
rect 995 925 999 929
rect 1012 930 1016 934
rect 1091 935 1095 939
rect 1141 935 1145 939
rect 1194 935 1198 939
rect 1438 938 1442 942
rect 1454 938 1458 944
rect 1488 944 1492 948
rect 1475 938 1479 942
rect 1496 938 1500 942
rect 1512 938 1516 944
rect 1557 948 1561 952
rect 1570 951 1574 957
rect 1607 951 1611 957
rect 1620 953 1624 957
rect 1644 957 1648 961
rect 1718 957 1722 961
rect 1628 951 1632 957
rect 1665 951 1669 957
rect 1681 953 1685 957
rect 1533 938 1537 942
rect 1549 938 1553 942
rect 1570 938 1574 942
rect 1586 938 1590 944
rect 1620 944 1624 948
rect 1607 938 1611 942
rect 1628 938 1632 942
rect 1644 938 1648 944
rect 1689 948 1693 952
rect 1702 951 1706 957
rect 1739 951 1743 957
rect 1752 953 1756 957
rect 1776 957 1780 961
rect 1850 957 1854 961
rect 1760 951 1764 957
rect 1797 951 1801 957
rect 1813 953 1817 957
rect 1665 938 1669 942
rect 1681 938 1685 942
rect 1702 938 1706 942
rect 1718 938 1722 944
rect 1752 944 1756 948
rect 1739 938 1743 942
rect 1760 938 1764 942
rect 1776 938 1780 944
rect 1821 948 1825 952
rect 1834 951 1838 957
rect 1871 951 1875 957
rect 1884 953 1888 957
rect 1908 957 1912 961
rect 1892 951 1896 957
rect 1929 951 1933 957
rect 1945 953 1949 957
rect 1797 938 1801 942
rect 1813 938 1817 942
rect 1834 938 1838 942
rect 1850 938 1854 944
rect 1884 944 1888 948
rect 1871 938 1875 942
rect 1114 924 1118 928
rect 429 918 435 922
rect 165 905 169 909
rect 181 905 185 911
rect 215 911 219 915
rect 202 905 206 909
rect 223 905 227 909
rect 239 905 243 911
rect 1076 915 1080 919
rect 1098 918 1102 924
rect 1135 918 1139 924
rect 1148 920 1152 924
rect 1172 924 1176 928
rect 1156 918 1160 924
rect 1193 918 1197 924
rect 1209 918 1213 924
rect 1431 927 1435 931
rect 1468 925 1472 929
rect 1488 925 1492 929
rect 1532 925 1536 929
rect 1563 927 1567 931
rect 1600 925 1604 929
rect 1620 925 1624 929
rect 1664 925 1668 929
rect 1695 927 1699 931
rect 1732 925 1736 929
rect 1752 925 1756 929
rect 1796 925 1800 929
rect 1813 930 1817 934
rect 1892 938 1896 942
rect 1908 938 1912 944
rect 1929 938 1933 942
rect 1945 938 1949 942
rect 1827 927 1831 931
rect 1864 925 1868 929
rect 1884 925 1888 929
rect 1928 925 1932 929
rect 1945 930 1949 934
rect 1362 918 1368 922
rect 465 911 471 915
rect 498 911 502 915
rect 549 911 553 915
rect 599 911 603 915
rect 630 911 634 915
rect 681 911 685 915
rect 731 911 735 915
rect 762 911 766 915
rect 813 911 817 915
rect 863 911 867 915
rect 894 911 898 915
rect 945 911 949 915
rect 995 911 999 915
rect 260 905 264 909
rect 276 905 280 909
rect 1098 905 1102 909
rect 1114 905 1118 911
rect 1148 911 1152 915
rect 1135 905 1139 909
rect 158 894 162 898
rect 195 892 199 896
rect 215 892 219 896
rect 259 892 263 896
rect 417 898 423 902
rect 496 898 500 902
rect 530 898 534 902
rect 547 898 551 902
rect 603 898 607 902
rect 620 898 624 902
rect 648 898 652 902
rect 1156 905 1160 909
rect 1172 905 1176 911
rect 1398 911 1404 915
rect 1431 911 1435 915
rect 1482 911 1486 915
rect 1532 911 1536 915
rect 1563 911 1567 915
rect 1614 911 1618 915
rect 1664 911 1668 915
rect 1695 911 1699 915
rect 1746 911 1750 915
rect 1796 911 1800 915
rect 1827 911 1831 915
rect 1878 911 1882 915
rect 1928 911 1932 915
rect 1193 905 1197 909
rect 1209 905 1213 909
rect 453 891 459 895
rect 523 891 527 895
rect 554 891 558 895
rect 576 891 580 895
rect 641 891 645 895
rect 429 885 435 889
rect 158 878 162 882
rect 209 878 213 882
rect 259 878 263 882
rect 465 878 471 882
rect 497 881 501 885
rect 522 884 526 888
rect 529 881 533 885
rect 547 881 551 885
rect 569 884 573 888
rect 594 884 598 888
rect 604 881 608 885
rect 620 881 624 885
rect 640 884 644 888
rect 647 881 651 885
rect 711 891 715 895
rect 276 871 280 875
rect 143 862 147 866
rect 268 864 272 868
rect 292 864 296 868
rect 151 855 155 859
rect 292 855 296 859
rect 524 865 528 869
rect 544 862 548 866
rect 563 866 567 870
rect 665 877 669 881
rect 680 877 684 881
rect 582 865 586 869
rect 601 865 605 869
rect 614 864 618 868
rect 636 865 640 869
rect 644 864 648 868
rect 656 864 660 868
rect 497 851 501 855
rect 529 851 533 855
rect 547 851 551 855
rect 604 851 608 855
rect 619 851 623 855
rect 647 851 651 855
rect 158 847 162 851
rect 225 847 229 851
rect 261 847 265 851
rect 477 847 483 851
rect 511 847 515 851
rect 554 846 558 850
rect 576 847 583 851
rect 626 846 630 850
rect 417 840 423 844
rect 158 833 162 837
rect 211 833 215 837
rect 261 833 265 837
rect 441 839 447 843
rect 511 839 515 843
rect 570 839 574 843
rect 595 839 599 843
rect 626 839 630 843
rect 719 869 723 877
rect 792 891 796 895
rect 746 877 750 881
rect 761 877 765 881
rect 1091 894 1095 898
rect 1128 892 1132 896
rect 1148 892 1152 896
rect 1192 892 1196 896
rect 1350 898 1356 902
rect 1429 898 1433 902
rect 1463 898 1467 902
rect 1480 898 1484 902
rect 1536 898 1540 902
rect 1553 898 1557 902
rect 1581 898 1585 902
rect 1386 891 1392 895
rect 1456 891 1460 895
rect 1487 891 1491 895
rect 1509 891 1513 895
rect 1574 891 1578 895
rect 742 869 746 873
rect 688 863 692 867
rect 701 855 705 859
rect 800 869 804 877
rect 1362 885 1368 889
rect 1091 878 1095 882
rect 1142 878 1146 882
rect 1192 878 1196 882
rect 1398 878 1404 882
rect 1430 881 1434 885
rect 1455 884 1459 888
rect 1462 881 1466 885
rect 1480 881 1484 885
rect 1502 884 1506 888
rect 1527 884 1531 888
rect 1537 881 1541 885
rect 1553 881 1557 885
rect 1573 884 1577 888
rect 1580 881 1584 885
rect 1644 891 1648 895
rect 827 869 831 873
rect 1209 871 1213 875
rect 769 863 773 867
rect 1076 862 1080 866
rect 1201 864 1205 868
rect 1225 864 1229 868
rect 782 855 786 859
rect 1084 855 1088 859
rect 1225 855 1229 859
rect 1457 865 1461 869
rect 1477 862 1481 866
rect 1496 866 1500 870
rect 1598 877 1602 881
rect 1613 877 1617 881
rect 1515 865 1519 869
rect 1534 865 1538 869
rect 1547 864 1551 868
rect 1569 865 1573 869
rect 1577 864 1581 868
rect 1589 864 1593 868
rect 1430 851 1434 855
rect 1462 851 1466 855
rect 1480 851 1484 855
rect 1537 851 1541 855
rect 1552 851 1556 855
rect 1580 851 1584 855
rect 1091 847 1095 851
rect 1158 847 1162 851
rect 1194 847 1198 851
rect 1410 847 1416 851
rect 1444 847 1448 851
rect 1487 846 1491 850
rect 1509 847 1516 851
rect 1559 846 1563 850
rect 1350 840 1356 844
rect 429 832 435 836
rect 497 832 501 836
rect 511 832 515 836
rect 529 832 533 836
rect 547 832 551 836
rect 570 832 574 836
rect 604 832 608 836
rect 619 832 623 836
rect 647 832 651 836
rect 180 822 184 826
rect 143 816 147 822
rect 159 816 163 822
rect 196 816 200 822
rect 204 818 208 822
rect 238 822 242 826
rect 441 825 447 829
rect 511 825 515 829
rect 570 825 574 829
rect 595 825 599 829
rect 626 825 630 829
rect 217 816 221 822
rect 254 816 258 822
rect 511 817 515 821
rect 554 818 558 822
rect 576 817 583 821
rect 626 818 630 822
rect 276 813 280 817
rect 497 813 501 817
rect 529 813 533 817
rect 547 813 551 817
rect 604 813 608 817
rect 619 813 623 817
rect 647 813 651 817
rect 143 803 147 807
rect 159 803 163 807
rect 204 809 208 813
rect 180 803 184 809
rect 196 803 200 807
rect 217 803 221 807
rect 238 803 242 809
rect 254 803 258 807
rect 492 801 496 805
rect 160 790 164 794
rect 204 790 208 794
rect 224 790 228 794
rect 261 792 265 796
rect 524 799 528 803
rect 544 802 548 806
rect 563 798 567 802
rect 582 799 586 803
rect 601 799 605 803
rect 614 800 618 804
rect 711 815 715 819
rect 1091 833 1095 837
rect 1144 833 1148 837
rect 1194 833 1198 837
rect 1374 839 1380 843
rect 1444 839 1448 843
rect 1503 839 1507 843
rect 1528 839 1532 843
rect 1559 839 1563 843
rect 1652 869 1656 877
rect 1725 891 1729 895
rect 1679 877 1683 881
rect 1694 877 1698 881
rect 1675 869 1679 873
rect 1621 863 1625 867
rect 1634 855 1638 859
rect 1733 869 1737 877
rect 1760 869 1764 873
rect 1702 863 1706 867
rect 1715 855 1719 859
rect 1362 832 1368 836
rect 1430 832 1434 836
rect 1444 832 1448 836
rect 1462 832 1466 836
rect 1480 832 1484 836
rect 1503 832 1507 836
rect 1537 832 1541 836
rect 1552 832 1556 836
rect 1580 832 1584 836
rect 1113 822 1117 826
rect 792 815 796 819
rect 1076 816 1080 822
rect 1092 816 1096 822
rect 1129 816 1133 822
rect 1137 818 1141 822
rect 1171 822 1175 826
rect 1374 825 1380 829
rect 1444 825 1448 829
rect 1503 825 1507 829
rect 1528 825 1532 829
rect 1559 825 1563 829
rect 1150 816 1154 822
rect 1187 816 1191 822
rect 1444 817 1448 821
rect 1487 818 1491 822
rect 1509 817 1516 821
rect 1559 818 1563 822
rect 1209 813 1213 817
rect 1430 813 1434 817
rect 1462 813 1466 817
rect 1480 813 1484 817
rect 1537 813 1541 817
rect 1552 813 1556 817
rect 1580 813 1584 817
rect 636 799 640 803
rect 644 800 648 804
rect 656 800 660 804
rect 691 800 695 804
rect 719 799 723 803
rect 771 800 775 804
rect 1076 803 1080 807
rect 1092 803 1096 807
rect 1137 809 1141 813
rect 1113 803 1117 809
rect 1129 803 1133 807
rect 800 799 804 803
rect 1150 803 1154 807
rect 1171 803 1175 809
rect 1187 803 1191 807
rect 1425 801 1429 805
rect 429 783 435 787
rect 497 783 501 787
rect 522 780 526 784
rect 529 783 533 787
rect 547 783 551 787
rect 569 780 573 784
rect 594 780 598 784
rect 604 783 608 787
rect 620 783 624 787
rect 640 780 644 784
rect 647 783 651 787
rect 160 776 164 780
rect 210 776 214 780
rect 261 776 265 780
rect 465 776 471 780
rect 507 773 511 777
rect 523 773 527 777
rect 554 773 558 777
rect 576 773 580 777
rect 641 773 645 777
rect 701 779 705 783
rect 1093 790 1097 794
rect 1137 790 1141 794
rect 1157 790 1161 794
rect 1194 792 1198 796
rect 1457 799 1461 803
rect 1477 802 1481 806
rect 1496 798 1500 802
rect 1515 799 1519 803
rect 1534 799 1538 803
rect 1547 800 1551 804
rect 1644 815 1648 819
rect 1725 815 1729 819
rect 1569 799 1573 803
rect 1577 800 1581 804
rect 1589 800 1593 804
rect 1624 800 1628 804
rect 1652 799 1656 803
rect 1704 800 1708 804
rect 1733 799 1737 803
rect 1362 783 1368 787
rect 1430 783 1434 787
rect 782 779 786 783
rect 1455 780 1459 784
rect 1462 783 1466 787
rect 1480 783 1484 787
rect 1502 780 1506 784
rect 1527 780 1531 784
rect 1537 783 1541 787
rect 1553 783 1557 787
rect 1573 780 1577 784
rect 1580 783 1584 787
rect 1093 776 1097 780
rect 1143 776 1147 780
rect 1194 776 1198 780
rect 1398 776 1404 780
rect 1440 773 1444 777
rect 1456 773 1460 777
rect 1487 773 1491 777
rect 1509 773 1513 777
rect 1574 773 1578 777
rect 1634 779 1638 783
rect 1715 779 1719 783
rect 417 766 423 770
rect 496 766 500 770
rect 530 766 534 770
rect 547 766 551 770
rect 603 766 607 770
rect 620 766 624 770
rect 648 766 652 770
rect 1350 766 1356 770
rect 1429 766 1433 770
rect 1463 766 1467 770
rect 1480 766 1484 770
rect 1536 766 1540 770
rect 1553 766 1557 770
rect 1581 766 1585 770
rect 453 759 459 763
rect 507 759 511 763
rect 523 759 527 763
rect 554 759 558 763
rect 576 759 580 763
rect 641 759 645 763
rect 711 759 715 763
rect 497 749 501 753
rect 522 752 526 756
rect 529 749 533 753
rect 547 749 551 753
rect 569 752 573 756
rect 594 752 598 756
rect 604 749 608 753
rect 620 749 624 753
rect 640 752 644 756
rect 647 749 651 753
rect 491 732 495 736
rect 524 733 528 737
rect 544 730 548 734
rect 563 734 567 738
rect 582 733 586 737
rect 601 733 605 737
rect 614 732 618 736
rect 636 733 640 737
rect 644 732 648 736
rect 656 732 660 736
rect 719 737 723 745
rect 816 759 820 763
rect 770 745 774 749
rect 785 745 789 749
rect 1386 759 1392 763
rect 1440 759 1444 763
rect 1456 759 1460 763
rect 1487 759 1491 763
rect 1509 759 1513 763
rect 1574 759 1578 763
rect 1644 759 1648 763
rect 688 731 692 735
rect 742 736 746 740
rect 497 719 501 723
rect 529 719 533 723
rect 547 719 551 723
rect 604 719 608 723
rect 619 719 623 723
rect 647 719 651 723
rect 511 715 515 719
rect 554 714 558 718
rect 576 715 583 719
rect 626 714 630 718
rect 441 707 447 711
rect 511 707 515 711
rect 570 707 574 711
rect 595 707 599 711
rect 626 707 630 711
rect 701 723 705 727
rect 824 737 828 745
rect 1430 749 1434 753
rect 1455 752 1459 756
rect 1462 749 1466 753
rect 1480 749 1484 753
rect 1502 752 1506 756
rect 1527 752 1531 756
rect 1537 749 1541 753
rect 1553 749 1557 753
rect 1573 752 1577 756
rect 1580 749 1584 753
rect 845 737 849 741
rect 793 731 797 735
rect 1424 732 1428 736
rect 806 723 810 727
rect 1457 733 1461 737
rect 1477 730 1481 734
rect 1496 734 1500 738
rect 1515 733 1519 737
rect 1534 733 1538 737
rect 1547 732 1551 736
rect 1569 733 1573 737
rect 1577 732 1581 736
rect 1589 732 1593 736
rect 1652 737 1656 745
rect 1749 759 1753 763
rect 1703 745 1707 749
rect 1718 745 1722 749
rect 1621 731 1625 735
rect 1675 736 1679 740
rect 1430 719 1434 723
rect 1462 719 1466 723
rect 1480 719 1484 723
rect 1537 719 1541 723
rect 1552 719 1556 723
rect 1580 719 1584 723
rect 1444 715 1448 719
rect 1487 714 1491 718
rect 1509 715 1516 719
rect 1559 714 1563 718
rect 1374 707 1380 711
rect 1444 707 1448 711
rect 1503 707 1507 711
rect 1528 707 1532 711
rect 1559 707 1563 711
rect 1634 723 1638 727
rect 1757 737 1761 745
rect 1778 737 1782 741
rect 1726 731 1730 735
rect 1739 723 1743 727
rect 429 700 435 704
rect 497 700 501 704
rect 511 700 515 704
rect 529 700 533 704
rect 547 700 551 704
rect 570 700 574 704
rect 604 700 608 704
rect 619 700 623 704
rect 647 700 651 704
rect 1362 700 1368 704
rect 1430 700 1434 704
rect 1444 700 1448 704
rect 1462 700 1466 704
rect 1480 700 1484 704
rect 1503 700 1507 704
rect 1537 700 1541 704
rect 1552 700 1556 704
rect 1580 700 1584 704
rect 441 693 447 697
rect 511 693 515 697
rect 570 693 574 697
rect 595 693 599 697
rect 626 693 630 697
rect 511 685 515 689
rect 554 686 558 690
rect 576 685 583 689
rect 626 686 630 690
rect 497 681 501 685
rect 529 681 533 685
rect 547 681 551 685
rect 604 681 608 685
rect 619 681 623 685
rect 647 681 651 685
rect 711 684 715 688
rect 1374 693 1380 697
rect 1444 693 1448 697
rect 1503 693 1507 697
rect 1528 693 1532 697
rect 1559 693 1563 697
rect 816 684 820 688
rect 1444 685 1448 689
rect 1487 686 1491 690
rect 1509 685 1516 689
rect 1559 686 1563 690
rect 1430 681 1434 685
rect 1462 681 1466 685
rect 1480 681 1484 685
rect 1537 681 1541 685
rect 1552 681 1556 685
rect 1580 681 1584 685
rect 1644 684 1648 688
rect 1749 684 1753 688
rect 492 669 496 673
rect 524 667 528 671
rect 544 670 548 674
rect 563 666 567 670
rect 582 667 586 671
rect 601 667 605 671
rect 614 668 618 672
rect 636 667 640 671
rect 644 668 648 672
rect 656 668 660 672
rect 690 669 694 673
rect 719 668 723 672
rect 796 669 800 673
rect 824 668 828 672
rect 1425 669 1429 673
rect 497 651 501 655
rect 522 648 526 652
rect 529 651 533 655
rect 547 651 551 655
rect 569 648 573 652
rect 594 648 598 652
rect 604 651 608 655
rect 620 651 624 655
rect 640 648 644 652
rect 647 651 651 655
rect 453 641 459 645
rect 523 641 527 645
rect 554 641 558 645
rect 576 641 580 645
rect 641 641 645 645
rect 701 648 705 652
rect 1457 667 1461 671
rect 1477 670 1481 674
rect 1496 666 1500 670
rect 1515 667 1519 671
rect 1534 667 1538 671
rect 1547 668 1551 672
rect 1569 667 1573 671
rect 1577 668 1581 672
rect 1589 668 1593 672
rect 1623 669 1627 673
rect 1652 668 1656 672
rect 1729 669 1733 673
rect 1757 668 1761 672
rect 806 648 810 652
rect 1430 651 1434 655
rect 1455 648 1459 652
rect 1462 651 1466 655
rect 1480 651 1484 655
rect 1502 648 1506 652
rect 1527 648 1531 652
rect 1537 651 1541 655
rect 1553 651 1557 655
rect 1573 648 1577 652
rect 1580 651 1584 655
rect 1386 641 1392 645
rect 1456 641 1460 645
rect 1487 641 1491 645
rect 1509 641 1513 645
rect 1574 641 1578 645
rect 1634 648 1638 652
rect 1739 648 1743 652
rect 417 634 423 638
rect 496 634 500 638
rect 530 634 534 638
rect 547 634 551 638
rect 603 634 607 638
rect 620 634 624 638
rect 648 634 652 638
rect 1350 634 1356 638
rect 1429 634 1433 638
rect 1463 634 1467 638
rect 1480 634 1484 638
rect 1536 634 1540 638
rect 1553 634 1557 638
rect 1581 634 1585 638
rect 453 627 459 631
rect 523 627 527 631
rect 554 627 558 631
rect 576 627 580 631
rect 641 627 645 631
rect 711 627 715 631
rect 497 617 501 621
rect 522 620 526 624
rect 529 617 533 621
rect 547 617 551 621
rect 569 620 573 624
rect 594 620 598 624
rect 604 617 608 621
rect 620 617 624 621
rect 640 620 644 624
rect 647 617 651 621
rect 491 600 495 604
rect 524 601 528 605
rect 544 598 548 602
rect 563 602 567 606
rect 582 601 586 605
rect 601 601 605 605
rect 614 600 618 604
rect 636 601 640 605
rect 644 600 648 604
rect 656 600 660 604
rect 719 605 723 613
rect 792 627 796 631
rect 746 613 750 617
rect 761 613 765 617
rect 742 605 746 609
rect 688 599 692 603
rect 497 587 501 591
rect 529 587 533 591
rect 547 587 551 591
rect 604 587 608 591
rect 619 587 623 591
rect 647 587 651 591
rect 511 583 515 587
rect 554 582 558 586
rect 576 583 583 587
rect 626 582 630 586
rect 441 575 447 579
rect 511 575 515 579
rect 570 575 574 579
rect 595 575 599 579
rect 626 575 630 579
rect 701 591 705 595
rect 800 605 804 613
rect 882 627 886 631
rect 836 613 840 617
rect 851 613 855 617
rect 1386 627 1392 631
rect 1456 627 1460 631
rect 1487 627 1491 631
rect 1509 627 1513 631
rect 1574 627 1578 631
rect 1644 627 1648 631
rect 824 605 828 609
rect 769 599 773 603
rect 858 607 862 611
rect 890 605 894 613
rect 1430 617 1434 621
rect 1455 620 1459 624
rect 1462 617 1466 621
rect 1480 617 1484 621
rect 1502 620 1506 624
rect 1527 620 1531 624
rect 1537 617 1541 621
rect 1553 617 1557 621
rect 1573 620 1577 624
rect 1580 617 1584 621
rect 782 591 786 595
rect 925 604 929 608
rect 1424 600 1428 604
rect 872 591 876 595
rect 1457 601 1461 605
rect 1477 598 1481 602
rect 1496 602 1500 606
rect 1515 601 1519 605
rect 1534 601 1538 605
rect 1547 600 1551 604
rect 1569 601 1573 605
rect 1577 600 1581 604
rect 1589 600 1593 604
rect 1652 605 1656 613
rect 1725 627 1729 631
rect 1679 613 1683 617
rect 1694 613 1698 617
rect 1675 605 1679 609
rect 1621 599 1625 603
rect 1430 587 1434 591
rect 1462 587 1466 591
rect 1480 587 1484 591
rect 1537 587 1541 591
rect 1552 587 1556 591
rect 1580 587 1584 591
rect 1444 583 1448 587
rect 1487 582 1491 586
rect 1509 583 1516 587
rect 1559 582 1563 586
rect 1374 575 1380 579
rect 1444 575 1448 579
rect 1503 575 1507 579
rect 1528 575 1532 579
rect 1559 575 1563 579
rect 1634 591 1638 595
rect 1733 605 1737 613
rect 1815 627 1819 631
rect 1769 613 1773 617
rect 1784 613 1788 617
rect 1757 605 1761 609
rect 1702 599 1706 603
rect 1791 607 1795 611
rect 1823 605 1827 613
rect 1715 591 1719 595
rect 1858 604 1862 608
rect 1805 591 1809 595
rect 429 568 435 572
rect 497 568 501 572
rect 511 568 515 572
rect 529 568 533 572
rect 547 568 551 572
rect 570 568 574 572
rect 604 568 608 572
rect 619 568 623 572
rect 647 568 651 572
rect 1362 568 1368 572
rect 1430 568 1434 572
rect 1444 568 1448 572
rect 1462 568 1466 572
rect 1480 568 1484 572
rect 1503 568 1507 572
rect 1537 568 1541 572
rect 1552 568 1556 572
rect 1580 568 1584 572
rect 441 561 447 565
rect 511 561 515 565
rect 570 561 574 565
rect 595 561 599 565
rect 626 561 630 565
rect 511 553 515 557
rect 554 554 558 558
rect 576 553 583 557
rect 626 554 630 558
rect 497 549 501 553
rect 529 549 533 553
rect 547 549 551 553
rect 604 549 608 553
rect 619 549 623 553
rect 647 549 651 553
rect 492 537 496 541
rect 524 535 528 539
rect 544 538 548 542
rect 563 534 567 538
rect 582 535 586 539
rect 601 535 605 539
rect 614 536 618 540
rect 711 549 715 553
rect 792 549 796 553
rect 1374 561 1380 565
rect 1444 561 1448 565
rect 1503 561 1507 565
rect 1528 561 1532 565
rect 1559 561 1563 565
rect 1444 553 1448 557
rect 1487 554 1491 558
rect 1509 553 1516 557
rect 1559 554 1563 558
rect 882 549 886 553
rect 1430 549 1434 553
rect 1462 549 1466 553
rect 1480 549 1484 553
rect 1537 549 1541 553
rect 1552 549 1556 553
rect 1580 549 1584 553
rect 636 535 640 539
rect 644 536 648 540
rect 656 536 660 540
rect 691 534 695 538
rect 719 533 723 537
rect 771 534 775 538
rect 800 533 804 537
rect 855 534 859 538
rect 1425 537 1429 541
rect 890 533 894 537
rect 497 519 501 523
rect 522 516 526 520
rect 529 519 533 523
rect 547 519 551 523
rect 569 516 573 520
rect 594 516 598 520
rect 604 519 608 523
rect 620 519 624 523
rect 640 516 644 520
rect 647 519 651 523
rect 1457 535 1461 539
rect 1477 538 1481 542
rect 1496 534 1500 538
rect 1515 535 1519 539
rect 1534 535 1538 539
rect 1547 536 1551 540
rect 1644 549 1648 553
rect 1725 549 1729 553
rect 1815 549 1819 553
rect 1569 535 1573 539
rect 1577 536 1581 540
rect 1589 536 1593 540
rect 1624 534 1628 538
rect 1652 533 1656 537
rect 1704 534 1708 538
rect 1733 533 1737 537
rect 1788 534 1792 538
rect 1823 533 1827 537
rect 453 509 459 513
rect 523 509 527 513
rect 554 509 558 513
rect 576 509 580 513
rect 641 509 645 513
rect 701 513 705 517
rect 782 513 786 517
rect 1430 519 1434 523
rect 872 513 876 517
rect 1455 516 1459 520
rect 1462 519 1466 523
rect 1480 519 1484 523
rect 1502 516 1506 520
rect 1527 516 1531 520
rect 1537 519 1541 523
rect 1553 519 1557 523
rect 1573 516 1577 520
rect 1580 519 1584 523
rect 1386 509 1392 513
rect 1456 509 1460 513
rect 1487 509 1491 513
rect 1509 509 1513 513
rect 1574 509 1578 513
rect 1634 513 1638 517
rect 1715 513 1719 517
rect 1805 513 1809 517
rect 417 502 423 506
rect 496 502 500 506
rect 530 502 534 506
rect 547 502 551 506
rect 603 502 607 506
rect 620 502 624 506
rect 648 502 652 506
rect 1350 502 1356 506
rect 1429 502 1433 506
rect 1463 502 1467 506
rect 1480 502 1484 506
rect 1536 502 1540 506
rect 1553 502 1557 506
rect 1581 502 1585 506
rect 453 495 459 499
rect 523 495 527 499
rect 554 495 558 499
rect 576 495 580 499
rect 641 495 645 499
rect 711 495 715 499
rect 497 485 501 489
rect 522 488 526 492
rect 529 485 533 489
rect 547 485 551 489
rect 569 488 573 492
rect 594 488 598 492
rect 604 485 608 489
rect 620 485 624 489
rect 640 488 644 492
rect 647 485 651 489
rect 491 468 495 472
rect 524 469 528 473
rect 544 466 548 470
rect 563 470 567 474
rect 1386 495 1392 499
rect 1456 495 1460 499
rect 1487 495 1491 499
rect 1509 495 1513 499
rect 1574 495 1578 499
rect 1644 495 1648 499
rect 582 469 586 473
rect 601 469 605 473
rect 614 468 618 472
rect 636 469 640 473
rect 644 468 648 472
rect 656 468 660 472
rect 719 473 723 481
rect 1430 485 1434 489
rect 1455 488 1459 492
rect 1462 485 1466 489
rect 1480 485 1484 489
rect 1502 488 1506 492
rect 1527 488 1531 492
rect 1537 485 1541 489
rect 1553 485 1557 489
rect 1573 488 1577 492
rect 1580 485 1584 489
rect 688 467 692 471
rect 742 472 746 476
rect 1424 468 1428 472
rect 497 455 501 459
rect 529 455 533 459
rect 547 455 551 459
rect 604 455 608 459
rect 619 455 623 459
rect 647 455 651 459
rect 511 451 515 455
rect 26 447 30 451
rect 62 447 66 451
rect 129 447 133 451
rect 158 447 162 451
rect 194 447 198 451
rect 261 447 265 451
rect 290 447 294 451
rect 326 447 330 451
rect 393 447 397 451
rect 477 447 483 451
rect 554 450 558 454
rect 576 451 583 455
rect 626 450 630 454
rect 417 440 423 444
rect 511 443 515 447
rect 520 443 524 447
rect 570 443 574 447
rect 595 443 599 447
rect 626 443 630 447
rect 701 459 705 463
rect 1457 469 1461 473
rect 1477 466 1481 470
rect 1496 470 1500 474
rect 1515 469 1519 473
rect 1534 469 1538 473
rect 1547 468 1551 472
rect 1569 469 1573 473
rect 1577 468 1581 472
rect 1589 468 1593 472
rect 1652 473 1656 481
rect 1621 467 1625 471
rect 1675 472 1679 476
rect 1430 455 1434 459
rect 1462 455 1466 459
rect 1480 455 1484 459
rect 1537 455 1541 459
rect 1552 455 1556 459
rect 1580 455 1584 459
rect 1444 451 1448 455
rect 959 447 963 451
rect 995 447 999 451
rect 1062 447 1066 451
rect 1091 447 1095 451
rect 1127 447 1131 451
rect 1194 447 1198 451
rect 1223 447 1227 451
rect 1259 447 1263 451
rect 1326 447 1330 451
rect 1410 447 1416 451
rect 1487 450 1491 454
rect 1509 451 1516 455
rect 1559 450 1563 454
rect 1350 440 1356 444
rect 1444 443 1448 447
rect 1453 443 1457 447
rect 1503 443 1507 447
rect 1528 443 1532 447
rect 1559 443 1563 447
rect 1634 459 1638 463
rect 26 433 30 437
rect 76 433 80 437
rect 129 433 133 437
rect 158 433 162 437
rect 208 433 212 437
rect 261 433 265 437
rect 290 433 294 437
rect 340 433 344 437
rect 393 433 397 437
rect 429 436 435 440
rect 497 436 501 440
rect 511 436 515 440
rect 529 436 533 440
rect 547 436 551 440
rect 570 436 574 440
rect 604 436 608 440
rect 619 436 623 440
rect 647 436 651 440
rect 772 436 776 440
rect 790 436 794 440
rect 808 436 812 440
rect 831 436 835 440
rect 865 436 869 440
rect 880 436 884 440
rect 908 436 912 440
rect 49 422 53 426
rect 20 413 24 417
rect 33 416 37 422
rect 70 416 74 422
rect 83 418 87 422
rect 107 422 111 426
rect 181 422 185 426
rect 91 416 95 422
rect 128 416 132 422
rect 144 416 148 422
rect 165 416 169 422
rect 202 416 206 422
rect 215 418 219 422
rect 239 422 243 426
rect 313 422 317 426
rect 223 416 227 422
rect 260 416 264 422
rect 276 416 280 422
rect 297 416 301 422
rect 334 416 338 422
rect 347 418 351 422
rect 371 422 375 426
rect 441 429 447 433
rect 511 429 515 433
rect 520 429 524 433
rect 570 429 574 433
rect 595 429 599 433
rect 626 429 630 433
rect 355 416 359 422
rect 392 416 396 422
rect 408 418 412 422
rect 511 421 515 425
rect 554 422 558 426
rect 576 421 583 425
rect 626 422 630 426
rect 497 417 501 421
rect 529 417 533 421
rect 547 417 551 421
rect 604 417 608 421
rect 619 417 623 421
rect 647 417 651 421
rect 33 403 37 407
rect 49 403 53 409
rect 83 409 87 413
rect 70 403 74 407
rect 91 403 95 407
rect 107 403 111 409
rect 128 403 132 407
rect 144 403 148 407
rect 165 403 169 407
rect 181 403 185 409
rect 215 409 219 413
rect 202 403 206 407
rect 223 403 227 407
rect 239 403 243 409
rect 260 403 264 407
rect 276 403 280 407
rect 297 403 301 407
rect 313 403 317 409
rect 347 409 351 413
rect 334 403 338 407
rect 355 403 359 407
rect 371 403 375 409
rect 392 403 396 407
rect 408 403 412 407
rect 492 405 496 409
rect 26 392 30 396
rect 63 390 67 394
rect 83 390 87 394
rect 127 390 131 394
rect 158 392 162 396
rect 195 390 199 394
rect 215 390 219 394
rect 259 390 263 394
rect 290 392 294 396
rect 327 390 331 394
rect 347 390 351 394
rect 391 390 395 394
rect 524 403 528 407
rect 544 406 548 410
rect 563 402 567 406
rect 582 403 586 407
rect 601 403 605 407
rect 614 404 618 408
rect 750 429 754 433
rect 772 429 776 433
rect 831 429 835 433
rect 856 429 860 433
rect 887 429 891 433
rect 959 433 963 437
rect 1009 433 1013 437
rect 1062 433 1066 437
rect 1091 433 1095 437
rect 1141 433 1145 437
rect 1194 433 1198 437
rect 1223 433 1227 437
rect 1273 433 1277 437
rect 1326 433 1330 437
rect 1362 436 1368 440
rect 1430 436 1434 440
rect 1444 436 1448 440
rect 1462 436 1466 440
rect 1480 436 1484 440
rect 1503 436 1507 440
rect 1537 436 1541 440
rect 1552 436 1556 440
rect 1580 436 1584 440
rect 1705 436 1709 440
rect 1723 436 1727 440
rect 1741 436 1745 440
rect 1764 436 1768 440
rect 1798 436 1802 440
rect 1813 436 1817 440
rect 1841 436 1845 440
rect 772 421 776 425
rect 815 422 819 426
rect 837 421 844 425
rect 887 422 891 426
rect 982 422 986 426
rect 790 417 794 421
rect 808 417 812 421
rect 865 417 869 421
rect 880 417 884 421
rect 908 417 912 421
rect 711 413 715 417
rect 636 403 640 407
rect 644 404 648 408
rect 656 404 660 408
rect 690 398 694 402
rect 730 404 734 408
rect 719 397 723 401
rect 497 387 501 391
rect 429 383 435 387
rect 522 384 526 388
rect 529 387 533 391
rect 547 387 551 391
rect 569 384 573 388
rect 594 384 598 388
rect 604 387 608 391
rect 620 387 624 391
rect 640 384 644 388
rect 647 387 651 391
rect 785 403 789 407
rect 805 406 809 410
rect 824 402 828 406
rect 953 413 957 417
rect 966 416 970 422
rect 1003 416 1007 422
rect 1016 418 1020 422
rect 1040 422 1044 426
rect 1114 422 1118 426
rect 1024 416 1028 422
rect 1061 416 1065 422
rect 1077 416 1081 422
rect 1098 416 1102 422
rect 1135 416 1139 422
rect 1148 418 1152 422
rect 1172 422 1176 426
rect 1246 422 1250 426
rect 1156 416 1160 422
rect 1193 416 1197 422
rect 1209 416 1213 422
rect 1230 416 1234 422
rect 1267 416 1271 422
rect 1280 418 1284 422
rect 1304 422 1308 426
rect 1374 429 1380 433
rect 1444 429 1448 433
rect 1453 429 1457 433
rect 1503 429 1507 433
rect 1528 429 1532 433
rect 1559 429 1563 433
rect 1288 416 1292 422
rect 1325 416 1329 422
rect 1341 418 1345 422
rect 1444 421 1448 425
rect 1487 422 1491 426
rect 1509 421 1516 425
rect 1559 422 1563 426
rect 1430 417 1434 421
rect 1462 417 1466 421
rect 1480 417 1484 421
rect 1537 417 1541 421
rect 1552 417 1556 421
rect 1580 417 1584 421
rect 843 403 847 407
rect 862 403 866 407
rect 875 404 879 408
rect 897 403 901 407
rect 905 404 909 408
rect 917 404 921 408
rect 966 403 970 407
rect 982 403 986 409
rect 1016 409 1020 413
rect 1003 403 1007 407
rect 1024 403 1028 407
rect 1040 403 1044 409
rect 1061 403 1065 407
rect 1077 403 1081 407
rect 1098 403 1102 407
rect 1114 403 1118 409
rect 1148 409 1152 413
rect 1135 403 1139 407
rect 1156 403 1160 407
rect 1172 403 1176 409
rect 1193 403 1197 407
rect 1209 403 1213 407
rect 1230 403 1234 407
rect 1246 403 1250 409
rect 1280 409 1284 413
rect 1267 403 1271 407
rect 1288 403 1292 407
rect 1304 403 1308 409
rect 1325 403 1329 407
rect 1341 403 1345 407
rect 1425 405 1429 409
rect 731 387 735 391
rect 757 387 761 391
rect 26 376 30 380
rect 77 376 81 380
rect 127 376 131 380
rect 158 376 162 380
rect 209 376 213 380
rect 259 376 263 380
rect 290 376 294 380
rect 341 376 345 380
rect 391 376 395 380
rect 465 377 471 381
rect 505 377 509 381
rect 523 377 527 381
rect 554 377 558 381
rect 576 377 580 381
rect 641 377 645 381
rect 783 384 787 388
rect 790 387 794 391
rect 808 387 812 391
rect 830 384 834 388
rect 855 384 859 388
rect 865 387 869 391
rect 881 387 885 391
rect 901 384 905 388
rect 908 387 912 391
rect 959 392 963 396
rect 996 390 1000 394
rect 1016 390 1020 394
rect 1060 390 1064 394
rect 1091 392 1095 396
rect 1128 390 1132 394
rect 1148 390 1152 394
rect 1192 390 1196 394
rect 1223 392 1227 396
rect 1260 390 1264 394
rect 1280 390 1284 394
rect 1324 390 1328 394
rect 1457 403 1461 407
rect 1477 406 1481 410
rect 1496 402 1500 406
rect 1515 403 1519 407
rect 1534 403 1538 407
rect 1547 404 1551 408
rect 1683 429 1687 433
rect 1705 429 1709 433
rect 1764 429 1768 433
rect 1789 429 1793 433
rect 1820 429 1824 433
rect 1705 421 1709 425
rect 1748 422 1752 426
rect 1770 421 1777 425
rect 1820 422 1824 426
rect 1723 417 1727 421
rect 1741 417 1745 421
rect 1798 417 1802 421
rect 1813 417 1817 421
rect 1841 417 1845 421
rect 1644 413 1648 417
rect 1569 403 1573 407
rect 1577 404 1581 408
rect 1589 404 1593 408
rect 1623 398 1627 402
rect 1663 404 1667 408
rect 1652 397 1656 401
rect 1430 387 1434 391
rect 1362 383 1368 387
rect 1455 384 1459 388
rect 1462 387 1466 391
rect 1480 387 1484 391
rect 1502 384 1506 388
rect 1527 384 1531 388
rect 1537 387 1541 391
rect 1553 387 1557 391
rect 1573 384 1577 388
rect 1580 387 1584 391
rect 1718 403 1722 407
rect 1738 406 1742 410
rect 1757 402 1761 406
rect 1776 403 1780 407
rect 1795 403 1799 407
rect 1808 404 1812 408
rect 1830 403 1834 407
rect 1838 404 1842 408
rect 1850 404 1854 408
rect 1664 387 1668 391
rect 1690 387 1694 391
rect 701 377 705 381
rect 740 377 744 381
rect 784 377 788 381
rect 815 377 819 381
rect 837 377 841 381
rect 902 377 906 381
rect 959 376 963 380
rect 1010 376 1014 380
rect 1060 376 1064 380
rect 1091 376 1095 380
rect 1142 376 1146 380
rect 1192 376 1196 380
rect 1223 376 1227 380
rect 1274 376 1278 380
rect 1324 376 1328 380
rect 1398 377 1404 381
rect 1438 377 1442 381
rect 1456 377 1460 381
rect 1487 377 1491 381
rect 1509 377 1513 381
rect 1574 377 1578 381
rect 1716 384 1720 388
rect 1723 387 1727 391
rect 1741 387 1745 391
rect 1763 384 1767 388
rect 1788 384 1792 388
rect 1798 387 1802 391
rect 1814 387 1818 391
rect 1834 384 1838 388
rect 1841 387 1845 391
rect 1634 377 1638 381
rect 1673 377 1677 381
rect 1717 377 1721 381
rect 1748 377 1752 381
rect 1770 377 1774 381
rect 1835 377 1839 381
rect 20 369 24 373
rect 408 369 412 373
rect 417 370 423 374
rect 496 370 500 374
rect 530 370 534 374
rect 547 370 551 374
rect 603 370 607 374
rect 620 370 624 374
rect 648 370 652 374
rect 731 370 735 374
rect 757 370 761 374
rect 791 370 795 374
rect 808 370 812 374
rect 864 370 868 374
rect 881 370 885 374
rect 909 370 913 374
rect 953 369 957 373
rect 1341 369 1345 373
rect 1350 370 1356 374
rect 1429 370 1433 374
rect 1463 370 1467 374
rect 1480 370 1484 374
rect 1536 370 1540 374
rect 1553 370 1557 374
rect 1581 370 1585 374
rect 1664 370 1668 374
rect 1690 370 1694 374
rect 1724 370 1728 374
rect 1741 370 1745 374
rect 1797 370 1801 374
rect 1814 370 1818 374
rect 1842 370 1846 374
rect 143 362 148 366
rect 276 362 280 366
rect 453 363 459 367
rect 505 363 509 367
rect 739 363 743 367
rect 925 364 929 368
rect 937 364 941 368
rect 1076 362 1081 366
rect 1209 362 1213 366
rect 1386 363 1392 367
rect 1438 363 1442 367
rect 1672 363 1676 367
rect 1858 364 1862 368
rect 1870 364 1874 368
rect 151 355 155 359
rect 441 355 447 359
rect 749 356 753 360
rect 914 356 918 360
rect 135 351 139 355
rect 167 351 171 355
rect 1084 355 1088 359
rect 1374 355 1380 359
rect 1682 356 1686 360
rect 1847 356 1851 360
rect 1068 351 1072 355
rect 1100 351 1104 355
rect 135 344 139 348
rect 167 344 171 348
rect 1068 344 1072 348
rect 1100 344 1104 348
rect 151 337 155 341
rect 408 337 412 341
rect 477 337 483 341
rect 797 337 801 341
rect 833 337 837 341
rect 900 337 904 341
rect 1084 337 1088 341
rect 1341 337 1345 341
rect 1410 337 1416 341
rect 1730 337 1734 341
rect 1766 337 1770 341
rect 1833 337 1837 341
rect 408 329 412 333
rect 417 330 423 334
rect 783 330 787 334
rect 135 325 139 329
rect 167 325 171 329
rect 151 321 155 325
rect 797 323 801 327
rect 847 323 851 327
rect 900 323 904 327
rect 1341 329 1345 333
rect 1350 330 1356 334
rect 1716 330 1720 334
rect 1068 325 1072 329
rect 1100 325 1104 329
rect 1084 321 1088 325
rect 1730 323 1734 327
rect 1780 323 1784 327
rect 1833 323 1837 327
rect 143 314 148 318
rect 277 314 281 318
rect 820 312 824 316
rect 26 307 30 311
rect 62 307 66 311
rect 129 307 133 311
rect 158 307 162 311
rect 194 307 198 311
rect 261 307 265 311
rect 290 307 294 311
rect 326 307 330 311
rect 393 307 397 311
rect 477 307 483 311
rect 417 300 423 304
rect 791 303 795 307
rect 804 306 808 312
rect 841 306 845 312
rect 854 308 858 312
rect 878 312 882 316
rect 1076 314 1081 318
rect 1210 314 1214 318
rect 1753 312 1757 316
rect 862 306 866 312
rect 899 306 903 312
rect 915 306 919 312
rect 959 307 963 311
rect 995 307 999 311
rect 1062 307 1066 311
rect 1091 307 1095 311
rect 1127 307 1131 311
rect 1194 307 1198 311
rect 1223 307 1227 311
rect 1259 307 1263 311
rect 1326 307 1330 311
rect 1410 307 1416 311
rect 26 293 30 297
rect 76 293 80 297
rect 129 293 133 297
rect 158 293 162 297
rect 208 293 212 297
rect 261 293 265 297
rect 290 293 294 297
rect 340 293 344 297
rect 393 293 397 297
rect 804 293 808 297
rect 820 293 824 299
rect 854 299 858 303
rect 841 293 845 297
rect 49 282 53 286
rect 20 273 24 277
rect 33 276 37 282
rect 70 276 74 282
rect 83 278 87 282
rect 107 282 111 286
rect 181 282 185 286
rect 91 276 95 282
rect 128 276 132 282
rect 144 276 148 282
rect 165 276 169 282
rect 202 276 206 282
rect 215 278 219 282
rect 239 282 243 286
rect 313 282 317 286
rect 223 276 227 282
rect 260 276 264 282
rect 276 276 280 282
rect 297 276 301 282
rect 334 276 338 282
rect 347 278 351 282
rect 371 282 375 286
rect 355 276 359 282
rect 392 276 396 282
rect 408 278 412 282
rect 862 293 866 297
rect 878 293 882 299
rect 1350 300 1356 304
rect 1724 303 1728 307
rect 1737 306 1741 312
rect 1774 306 1778 312
rect 1787 308 1791 312
rect 1811 312 1815 316
rect 1795 306 1799 312
rect 1832 306 1836 312
rect 1848 306 1852 312
rect 899 293 903 297
rect 915 293 919 297
rect 959 293 963 297
rect 1009 293 1013 297
rect 1062 293 1066 297
rect 1091 293 1095 297
rect 1141 293 1145 297
rect 1194 293 1198 297
rect 1223 293 1227 297
rect 1273 293 1277 297
rect 1326 293 1330 297
rect 1737 293 1741 297
rect 1753 293 1757 299
rect 1787 299 1791 303
rect 1774 293 1778 297
rect 797 282 801 286
rect 834 280 838 284
rect 854 280 858 284
rect 898 280 902 284
rect 982 282 986 286
rect 33 263 37 267
rect 49 263 53 269
rect 83 269 87 273
rect 70 263 74 267
rect 91 263 95 267
rect 107 263 111 269
rect 128 263 132 267
rect 144 263 148 267
rect 165 263 169 267
rect 181 263 185 269
rect 215 269 219 273
rect 202 263 206 267
rect 223 263 227 267
rect 239 263 243 269
rect 260 263 264 267
rect 276 263 280 267
rect 297 263 301 267
rect 313 263 317 269
rect 347 269 351 273
rect 334 263 338 267
rect 355 263 359 267
rect 371 263 375 269
rect 429 273 435 277
rect 953 273 957 277
rect 966 276 970 282
rect 1003 276 1007 282
rect 1016 278 1020 282
rect 1040 282 1044 286
rect 1114 282 1118 286
rect 1024 276 1028 282
rect 1061 276 1065 282
rect 1077 276 1081 282
rect 1098 276 1102 282
rect 1135 276 1139 282
rect 1148 278 1152 282
rect 1172 282 1176 286
rect 1246 282 1250 286
rect 1156 276 1160 282
rect 1193 276 1197 282
rect 1209 276 1213 282
rect 1230 276 1234 282
rect 1267 276 1271 282
rect 1280 278 1284 282
rect 1304 282 1308 286
rect 1288 276 1292 282
rect 1325 276 1329 282
rect 1341 278 1345 282
rect 1795 293 1799 297
rect 1811 293 1815 299
rect 1832 293 1836 297
rect 1848 293 1852 297
rect 1730 282 1734 286
rect 1767 280 1771 284
rect 1787 280 1791 284
rect 1831 280 1835 284
rect 392 263 396 267
rect 408 263 412 267
rect 465 266 471 270
rect 797 266 801 270
rect 848 266 852 270
rect 898 266 902 270
rect 966 263 970 267
rect 982 263 986 269
rect 1016 269 1020 273
rect 1003 263 1007 267
rect 26 252 30 256
rect 63 250 67 254
rect 83 250 87 254
rect 127 250 131 254
rect 158 252 162 256
rect 195 250 199 254
rect 215 250 219 254
rect 259 250 263 254
rect 290 252 294 256
rect 327 250 331 254
rect 347 250 351 254
rect 391 250 395 254
rect 790 258 794 262
rect 915 259 919 263
rect 1024 263 1028 267
rect 1040 263 1044 269
rect 1061 263 1065 267
rect 1077 263 1081 267
rect 1098 263 1102 267
rect 1114 263 1118 269
rect 1148 269 1152 273
rect 1135 263 1139 267
rect 1156 263 1160 267
rect 1172 263 1176 269
rect 1193 263 1197 267
rect 1209 263 1213 267
rect 1230 263 1234 267
rect 1246 263 1250 269
rect 1280 269 1284 273
rect 1267 263 1271 267
rect 1288 263 1292 267
rect 1304 263 1308 269
rect 1362 273 1368 277
rect 1325 263 1329 267
rect 1341 263 1345 267
rect 1398 266 1404 270
rect 1730 266 1734 270
rect 1781 266 1785 270
rect 1831 266 1835 270
rect 477 251 483 255
rect 797 251 801 255
rect 833 251 837 255
rect 900 251 904 255
rect 429 243 435 247
rect 783 244 787 248
rect 959 252 963 256
rect 996 250 1000 254
rect 1016 250 1020 254
rect 1060 250 1064 254
rect 1091 252 1095 256
rect 1128 250 1132 254
rect 1148 250 1152 254
rect 1192 250 1196 254
rect 1223 252 1227 256
rect 1260 250 1264 254
rect 1280 250 1284 254
rect 1324 250 1328 254
rect 1723 258 1727 262
rect 1848 259 1852 263
rect 1410 251 1416 255
rect 1730 251 1734 255
rect 1766 251 1770 255
rect 1833 251 1837 255
rect 26 236 30 240
rect 77 236 81 240
rect 127 236 131 240
rect 158 236 162 240
rect 209 236 213 240
rect 259 236 263 240
rect 290 236 294 240
rect 341 236 345 240
rect 391 236 395 240
rect 465 236 471 240
rect 797 237 801 241
rect 847 237 851 241
rect 900 237 904 241
rect 1362 243 1368 247
rect 1716 244 1720 248
rect 959 236 963 240
rect 1010 236 1014 240
rect 1060 236 1064 240
rect 1091 236 1095 240
rect 1142 236 1146 240
rect 1192 236 1196 240
rect 1223 236 1227 240
rect 1274 236 1278 240
rect 1324 236 1328 240
rect 1398 236 1404 240
rect 1730 237 1734 241
rect 1780 237 1784 241
rect 1833 237 1837 241
rect 19 229 23 233
rect 408 229 412 233
rect 820 226 824 230
rect 26 221 30 225
rect 62 221 66 225
rect 129 221 133 225
rect 158 221 162 225
rect 194 221 198 225
rect 261 221 265 225
rect 290 221 294 225
rect 326 221 330 225
rect 393 221 397 225
rect 477 221 483 225
rect 417 214 423 218
rect 791 217 795 221
rect 804 220 808 226
rect 841 220 845 226
rect 854 222 858 226
rect 878 226 882 230
rect 952 229 956 233
rect 1341 229 1345 233
rect 1753 226 1757 230
rect 862 220 866 226
rect 899 220 903 226
rect 915 222 919 226
rect 937 220 941 224
rect 959 221 963 225
rect 995 221 999 225
rect 1062 221 1066 225
rect 1091 221 1095 225
rect 1127 221 1131 225
rect 1194 221 1198 225
rect 1223 221 1227 225
rect 1259 221 1263 225
rect 1326 221 1330 225
rect 1410 221 1416 225
rect 26 207 30 211
rect 76 207 80 211
rect 129 207 133 211
rect 158 207 162 211
rect 208 207 212 211
rect 261 207 265 211
rect 290 207 294 211
rect 340 207 344 211
rect 393 207 397 211
rect 804 207 808 211
rect 820 207 824 213
rect 854 213 858 217
rect 841 207 845 211
rect 49 196 53 200
rect 20 187 24 191
rect 33 190 37 196
rect 70 190 74 196
rect 83 192 87 196
rect 107 196 111 200
rect 181 196 185 200
rect 91 190 95 196
rect 128 190 132 196
rect 144 190 148 196
rect 165 190 169 196
rect 202 190 206 196
rect 215 192 219 196
rect 239 196 243 200
rect 313 196 317 200
rect 223 190 227 196
rect 260 190 264 196
rect 276 190 280 196
rect 297 190 301 196
rect 334 190 338 196
rect 347 192 351 196
rect 371 196 375 200
rect 355 190 359 196
rect 392 190 396 196
rect 408 192 412 196
rect 862 207 866 211
rect 878 207 882 213
rect 899 207 903 211
rect 915 207 919 216
rect 1350 214 1356 218
rect 1724 217 1728 221
rect 1737 220 1741 226
rect 1774 220 1778 226
rect 1787 222 1791 226
rect 1811 226 1815 230
rect 1795 220 1799 226
rect 1832 220 1836 226
rect 1848 222 1852 226
rect 1870 220 1874 224
rect 937 204 941 208
rect 959 207 963 211
rect 1009 207 1013 211
rect 1062 207 1066 211
rect 1091 207 1095 211
rect 1141 207 1145 211
rect 1194 207 1198 211
rect 1223 207 1227 211
rect 1273 207 1277 211
rect 1326 207 1330 211
rect 1737 207 1741 211
rect 1753 207 1757 213
rect 1787 213 1791 217
rect 1774 207 1778 211
rect 797 196 801 200
rect 834 194 838 198
rect 854 194 858 198
rect 898 194 902 198
rect 982 196 986 200
rect 33 177 37 181
rect 49 177 53 183
rect 83 183 87 187
rect 70 177 74 181
rect 91 177 95 181
rect 107 177 111 183
rect 128 177 132 181
rect 144 177 148 181
rect 165 177 169 181
rect 181 177 185 183
rect 215 183 219 187
rect 202 177 206 181
rect 223 177 227 181
rect 239 177 243 183
rect 260 177 264 181
rect 276 177 280 181
rect 297 177 301 181
rect 313 177 317 183
rect 347 183 351 187
rect 334 177 338 181
rect 355 177 359 181
rect 371 177 375 183
rect 429 187 435 191
rect 953 187 957 191
rect 966 190 970 196
rect 1003 190 1007 196
rect 1016 192 1020 196
rect 1040 196 1044 200
rect 1114 196 1118 200
rect 1024 190 1028 196
rect 1061 190 1065 196
rect 1077 190 1081 196
rect 1098 190 1102 196
rect 1135 190 1139 196
rect 1148 192 1152 196
rect 1172 196 1176 200
rect 1246 196 1250 200
rect 1156 190 1160 196
rect 1193 190 1197 196
rect 1209 190 1213 196
rect 1230 190 1234 196
rect 1267 190 1271 196
rect 1280 192 1284 196
rect 1304 196 1308 200
rect 1288 190 1292 196
rect 1325 190 1329 196
rect 1341 192 1345 196
rect 1795 207 1799 211
rect 1811 207 1815 213
rect 1832 207 1836 211
rect 1848 207 1852 216
rect 1870 204 1874 208
rect 1730 196 1734 200
rect 1767 194 1771 198
rect 1787 194 1791 198
rect 1831 194 1835 198
rect 392 177 396 181
rect 408 177 412 181
rect 465 180 471 184
rect 797 180 801 184
rect 848 180 852 184
rect 898 180 902 184
rect 966 177 970 181
rect 982 177 986 183
rect 1016 183 1020 187
rect 1003 177 1007 181
rect 1024 177 1028 181
rect 1040 177 1044 183
rect 1061 177 1065 181
rect 1077 177 1081 181
rect 1098 177 1102 181
rect 1114 177 1118 183
rect 1148 183 1152 187
rect 1135 177 1139 181
rect 1156 177 1160 181
rect 1172 177 1176 183
rect 1193 177 1197 181
rect 1209 177 1213 181
rect 1230 177 1234 181
rect 1246 177 1250 183
rect 1280 183 1284 187
rect 1267 177 1271 181
rect 1288 177 1292 181
rect 1304 177 1308 183
rect 1362 187 1368 191
rect 1325 177 1329 181
rect 1341 177 1345 181
rect 1398 180 1404 184
rect 1730 180 1734 184
rect 1781 180 1785 184
rect 1831 180 1835 184
rect 26 166 30 170
rect 63 164 67 168
rect 83 164 87 168
rect 127 164 131 168
rect 158 166 162 170
rect 195 164 199 168
rect 215 164 219 168
rect 259 164 263 168
rect 290 166 294 170
rect 327 164 331 168
rect 347 164 351 168
rect 391 164 395 168
rect 959 166 963 170
rect 996 164 1000 168
rect 1016 164 1020 168
rect 1060 164 1064 168
rect 1091 166 1095 170
rect 1128 164 1132 168
rect 1148 164 1152 168
rect 1192 164 1196 168
rect 1223 166 1227 170
rect 1260 164 1264 168
rect 1280 164 1284 168
rect 1324 164 1328 168
rect 429 157 435 161
rect 1362 157 1368 161
rect 26 150 30 154
rect 77 150 81 154
rect 127 150 131 154
rect 158 150 162 154
rect 209 150 213 154
rect 259 150 263 154
rect 290 150 294 154
rect 341 150 345 154
rect 391 150 395 154
rect 465 150 471 154
rect 959 150 963 154
rect 1010 150 1014 154
rect 1060 150 1064 154
rect 1091 150 1095 154
rect 1142 150 1146 154
rect 1192 150 1196 154
rect 1223 150 1227 154
rect 1274 150 1278 154
rect 1324 150 1328 154
rect 1398 150 1404 154
rect 19 143 23 147
rect 408 143 412 147
rect 952 143 956 147
rect 1341 143 1345 147
rect 144 136 148 140
rect 252 136 256 140
rect 276 136 280 140
rect 1077 136 1081 140
rect 1185 136 1189 140
rect 1209 136 1213 140
rect 268 129 272 133
rect 252 125 256 129
rect 284 125 288 129
rect 1201 129 1205 133
rect 1185 125 1189 129
rect 1217 125 1221 129
rect 252 118 256 122
rect 284 118 288 122
rect 937 118 941 122
rect 1185 118 1189 122
rect 1217 118 1221 122
rect 1870 118 1874 122
rect 268 111 272 115
rect 408 111 412 115
rect 1201 111 1205 115
rect 1341 111 1345 115
rect 408 103 412 107
rect 1341 103 1345 107
rect 252 99 256 103
rect 284 99 288 103
rect 268 95 272 99
rect 1185 99 1189 103
rect 1217 99 1221 103
rect 1201 95 1205 99
rect 144 88 148 92
rect 252 88 256 92
rect 276 88 280 92
rect 1077 88 1081 92
rect 1185 88 1189 92
rect 1209 88 1213 92
rect 26 81 30 85
rect 62 81 66 85
rect 129 81 133 85
rect 158 81 162 85
rect 194 81 198 85
rect 261 81 265 85
rect 290 81 294 85
rect 326 81 330 85
rect 393 81 397 85
rect 477 81 483 85
rect 959 81 963 85
rect 995 81 999 85
rect 1062 81 1066 85
rect 1091 81 1095 85
rect 1127 81 1131 85
rect 1194 81 1198 85
rect 1223 81 1227 85
rect 1259 81 1263 85
rect 1326 81 1330 85
rect 1410 81 1416 85
rect 417 74 423 78
rect 1350 74 1356 78
rect 26 67 30 71
rect 76 67 80 71
rect 129 67 133 71
rect 158 67 162 71
rect 208 67 212 71
rect 261 67 265 71
rect 290 67 294 71
rect 340 67 344 71
rect 393 67 397 71
rect 959 67 963 71
rect 1009 67 1013 71
rect 1062 67 1066 71
rect 1091 67 1095 71
rect 1141 67 1145 71
rect 1194 67 1198 71
rect 1223 67 1227 71
rect 1273 67 1277 71
rect 1326 67 1330 71
rect 49 56 53 60
rect 20 47 24 51
rect 33 50 37 56
rect 70 50 74 56
rect 83 52 87 56
rect 107 56 111 60
rect 181 56 185 60
rect 91 50 95 56
rect 128 50 132 56
rect 144 50 148 56
rect 165 50 169 56
rect 202 50 206 56
rect 215 52 219 56
rect 239 56 243 60
rect 313 56 317 60
rect 223 50 227 56
rect 260 50 264 56
rect 276 50 280 56
rect 297 50 301 56
rect 334 50 338 56
rect 347 52 351 56
rect 371 56 375 60
rect 982 56 986 60
rect 355 50 359 56
rect 392 50 396 56
rect 408 52 412 56
rect 33 37 37 41
rect 49 37 53 43
rect 83 43 87 47
rect 70 37 74 41
rect 91 37 95 41
rect 107 37 111 43
rect 128 37 132 41
rect 144 37 148 41
rect 165 37 169 41
rect 181 37 185 43
rect 215 43 219 47
rect 202 37 206 41
rect 223 37 227 41
rect 239 37 243 43
rect 260 37 264 41
rect 276 37 280 41
rect 297 37 301 41
rect 313 37 317 43
rect 347 43 351 47
rect 334 37 338 41
rect 355 37 359 41
rect 371 37 375 43
rect 953 47 957 51
rect 966 50 970 56
rect 1003 50 1007 56
rect 1016 52 1020 56
rect 1040 56 1044 60
rect 1114 56 1118 60
rect 1024 50 1028 56
rect 1061 50 1065 56
rect 1077 50 1081 56
rect 1098 50 1102 56
rect 1135 50 1139 56
rect 1148 52 1152 56
rect 1172 56 1176 60
rect 1246 56 1250 60
rect 1156 50 1160 56
rect 1193 50 1197 56
rect 1209 50 1213 56
rect 1230 50 1234 56
rect 1267 50 1271 56
rect 1280 52 1284 56
rect 1304 56 1308 60
rect 1288 50 1292 56
rect 1325 50 1329 56
rect 1341 52 1345 56
rect 392 37 396 41
rect 408 37 412 41
rect 966 37 970 41
rect 982 37 986 43
rect 1016 43 1020 47
rect 1003 37 1007 41
rect 1024 37 1028 41
rect 1040 37 1044 43
rect 1061 37 1065 41
rect 1077 37 1081 41
rect 1098 37 1102 41
rect 1114 37 1118 43
rect 1148 43 1152 47
rect 1135 37 1139 41
rect 1156 37 1160 41
rect 1172 37 1176 43
rect 1193 37 1197 41
rect 1209 37 1213 41
rect 1230 37 1234 41
rect 1246 37 1250 43
rect 1280 43 1284 47
rect 1267 37 1271 41
rect 1288 37 1292 41
rect 1304 37 1308 43
rect 1325 37 1329 41
rect 1341 37 1345 41
rect 26 26 30 30
rect 63 24 67 28
rect 83 24 87 28
rect 127 24 131 28
rect 158 26 162 30
rect 195 24 199 28
rect 215 24 219 28
rect 259 24 263 28
rect 290 26 294 30
rect 327 24 331 28
rect 347 24 351 28
rect 391 24 395 28
rect 959 26 963 30
rect 996 24 1000 28
rect 1016 24 1020 28
rect 1060 24 1064 28
rect 1091 26 1095 30
rect 1128 24 1132 28
rect 1148 24 1152 28
rect 1192 24 1196 28
rect 1223 26 1227 30
rect 1260 24 1264 28
rect 1280 24 1284 28
rect 1324 24 1328 28
rect 429 17 435 21
rect 1362 17 1368 21
rect 26 10 30 14
rect 77 10 81 14
rect 127 10 131 14
rect 158 10 162 14
rect 209 10 213 14
rect 259 10 263 14
rect 290 10 294 14
rect 341 10 345 14
rect 391 10 395 14
rect 465 10 471 14
rect 959 10 963 14
rect 1010 10 1014 14
rect 1060 10 1064 14
rect 1091 10 1095 14
rect 1142 10 1146 14
rect 1192 10 1196 14
rect 1223 10 1227 14
rect 1274 10 1278 14
rect 1324 10 1328 14
rect 1398 10 1404 14
<< metal2 >>
rect 143 1846 146 1895
rect 143 1802 146 1842
rect 151 1839 155 1982
rect 159 1919 162 1929
rect 166 1889 169 1898
rect 182 1891 185 1904
rect 195 1876 198 1929
rect 262 1919 265 1929
rect 202 1904 206 1908
rect 203 1889 206 1898
rect 158 1862 161 1874
rect 199 1872 200 1876
rect 209 1862 212 1915
rect 215 1895 218 1900
rect 224 1889 227 1898
rect 240 1891 243 1904
rect 261 1889 264 1898
rect 260 1862 263 1872
rect 143 1787 146 1796
rect 27 1417 30 1427
rect 34 1387 37 1396
rect 50 1389 53 1402
rect 63 1374 66 1427
rect 130 1417 133 1427
rect 70 1402 74 1406
rect 71 1387 74 1396
rect 26 1360 29 1372
rect 67 1370 68 1374
rect 77 1360 80 1413
rect 83 1393 86 1398
rect 92 1387 95 1396
rect 108 1389 111 1402
rect 129 1387 132 1396
rect 145 1387 148 1396
rect 128 1360 131 1370
rect 20 1257 23 1349
rect 145 1346 148 1383
rect 151 1339 155 1835
rect 268 1848 272 1982
rect 417 1959 423 1973
rect 417 1926 423 1955
rect 277 1896 280 1898
rect 277 1889 280 1892
rect 277 1855 280 1885
rect 417 1882 423 1922
rect 158 1817 161 1827
rect 159 1787 162 1796
rect 180 1789 183 1802
rect 196 1787 199 1796
rect 205 1793 208 1798
rect 160 1760 163 1770
rect 211 1760 214 1813
rect 217 1802 221 1806
rect 217 1787 220 1796
rect 225 1774 228 1827
rect 261 1817 264 1827
rect 238 1789 241 1802
rect 254 1787 257 1796
rect 223 1770 224 1774
rect 262 1760 265 1772
rect 159 1417 162 1427
rect 166 1387 169 1396
rect 182 1389 185 1402
rect 195 1374 198 1427
rect 262 1417 265 1427
rect 202 1402 206 1406
rect 203 1387 206 1396
rect 158 1360 161 1372
rect 199 1370 200 1374
rect 209 1360 212 1413
rect 215 1393 218 1398
rect 224 1387 227 1396
rect 240 1389 243 1402
rect 261 1387 264 1396
rect 260 1360 263 1370
rect 135 1328 139 1331
rect 135 1309 139 1324
rect 151 1321 155 1335
rect 167 1335 171 1339
rect 167 1328 171 1331
rect 167 1309 171 1324
rect 151 1305 155 1306
rect 167 1301 171 1305
rect 27 1277 30 1287
rect 34 1247 37 1256
rect 50 1249 53 1262
rect 63 1234 66 1287
rect 130 1277 133 1287
rect 70 1262 74 1266
rect 71 1247 74 1256
rect 26 1220 29 1232
rect 67 1230 68 1234
rect 77 1220 80 1273
rect 145 1262 148 1294
rect 83 1253 86 1258
rect 92 1247 95 1256
rect 108 1249 111 1262
rect 129 1247 132 1256
rect 145 1247 148 1256
rect 128 1220 131 1230
rect 20 1171 23 1209
rect 27 1191 30 1201
rect 34 1161 37 1170
rect 50 1163 53 1176
rect 63 1148 66 1201
rect 130 1191 133 1201
rect 70 1176 74 1180
rect 71 1161 74 1170
rect 26 1134 29 1146
rect 67 1144 68 1148
rect 77 1134 80 1187
rect 83 1167 86 1172
rect 92 1161 95 1170
rect 108 1163 111 1176
rect 129 1161 132 1170
rect 145 1161 148 1170
rect 128 1134 131 1144
rect 20 1031 23 1123
rect 145 1120 148 1157
rect 27 1051 30 1061
rect 34 1021 37 1030
rect 50 1023 53 1036
rect 63 1008 66 1061
rect 130 1051 133 1061
rect 70 1036 74 1040
rect 71 1021 74 1030
rect 26 994 29 1006
rect 67 1004 68 1008
rect 77 994 80 1047
rect 145 1036 148 1068
rect 83 1027 86 1032
rect 92 1021 95 1030
rect 108 1023 111 1036
rect 129 1021 132 1030
rect 145 1021 148 1030
rect 128 994 131 1004
rect 143 866 146 915
rect 143 822 146 862
rect 151 859 155 1301
rect 159 1277 162 1287
rect 166 1247 169 1256
rect 182 1249 185 1262
rect 195 1234 198 1287
rect 262 1277 265 1287
rect 202 1262 206 1266
rect 203 1247 206 1256
rect 158 1220 161 1232
rect 199 1230 200 1234
rect 209 1220 212 1273
rect 215 1253 218 1258
rect 224 1247 227 1256
rect 240 1249 243 1262
rect 261 1247 264 1256
rect 260 1220 263 1230
rect 159 1191 162 1201
rect 166 1161 169 1170
rect 182 1163 185 1176
rect 195 1148 198 1201
rect 262 1191 265 1201
rect 202 1176 206 1180
rect 203 1161 206 1170
rect 158 1134 161 1146
rect 199 1144 200 1148
rect 209 1134 212 1187
rect 215 1167 218 1172
rect 224 1161 227 1170
rect 240 1163 243 1176
rect 261 1161 264 1170
rect 260 1134 263 1144
rect 268 1113 272 1844
rect 292 1839 296 1844
rect 417 1824 423 1878
rect 417 1750 423 1820
rect 417 1618 423 1746
rect 417 1486 423 1614
rect 291 1417 294 1427
rect 277 1387 280 1396
rect 298 1387 301 1396
rect 314 1389 317 1402
rect 277 1346 280 1383
rect 327 1374 330 1427
rect 394 1417 397 1427
rect 417 1424 423 1482
rect 334 1402 338 1406
rect 335 1387 338 1396
rect 290 1360 293 1372
rect 331 1370 332 1374
rect 341 1360 344 1413
rect 347 1393 350 1398
rect 356 1387 359 1396
rect 372 1389 375 1402
rect 393 1387 396 1396
rect 409 1387 412 1398
rect 392 1360 395 1370
rect 409 1353 412 1383
rect 409 1321 412 1349
rect 417 1354 423 1420
rect 417 1314 423 1350
rect 277 1262 280 1294
rect 291 1277 294 1287
rect 277 1247 280 1256
rect 298 1247 301 1256
rect 314 1249 317 1262
rect 327 1234 330 1287
rect 394 1277 397 1287
rect 334 1262 338 1266
rect 335 1247 338 1256
rect 290 1220 293 1232
rect 331 1230 332 1234
rect 341 1220 344 1273
rect 409 1262 412 1309
rect 347 1253 350 1258
rect 356 1247 359 1256
rect 372 1249 375 1262
rect 393 1247 396 1256
rect 409 1247 412 1258
rect 392 1220 395 1230
rect 409 1213 412 1243
rect 417 1284 423 1310
rect 291 1191 294 1201
rect 277 1161 280 1170
rect 298 1161 301 1170
rect 314 1163 317 1176
rect 277 1120 280 1157
rect 327 1148 330 1201
rect 394 1191 397 1201
rect 417 1198 423 1280
rect 334 1176 338 1180
rect 335 1161 338 1170
rect 290 1134 293 1146
rect 331 1144 332 1148
rect 341 1134 344 1187
rect 347 1167 350 1172
rect 356 1161 359 1170
rect 372 1163 375 1176
rect 393 1161 396 1170
rect 409 1161 412 1172
rect 392 1134 395 1144
rect 409 1127 412 1157
rect 252 1102 256 1105
rect 252 1083 256 1098
rect 268 1095 272 1109
rect 284 1109 288 1113
rect 284 1102 288 1105
rect 284 1083 288 1098
rect 409 1095 412 1123
rect 268 1079 272 1080
rect 284 1075 288 1079
rect 159 1051 162 1061
rect 166 1021 169 1030
rect 182 1023 185 1036
rect 195 1008 198 1061
rect 262 1051 265 1061
rect 202 1036 206 1040
rect 203 1021 206 1030
rect 158 994 161 1006
rect 199 1004 200 1008
rect 209 994 212 1047
rect 215 1027 218 1032
rect 224 1021 227 1030
rect 240 1023 243 1036
rect 261 1021 264 1030
rect 260 994 263 1004
rect 159 939 162 949
rect 166 909 169 918
rect 182 911 185 924
rect 195 896 198 949
rect 262 939 265 949
rect 202 924 206 928
rect 203 909 206 918
rect 158 882 161 894
rect 199 892 200 896
rect 209 882 212 935
rect 215 915 218 920
rect 224 909 227 918
rect 240 911 243 924
rect 261 909 264 918
rect 260 882 263 892
rect 143 807 146 816
rect 27 437 30 447
rect 34 407 37 416
rect 50 409 53 422
rect 63 394 66 447
rect 130 437 133 447
rect 70 422 74 426
rect 71 407 74 416
rect 26 380 29 392
rect 67 390 68 394
rect 77 380 80 433
rect 83 413 86 418
rect 92 407 95 416
rect 108 409 111 422
rect 129 407 132 416
rect 145 407 148 416
rect 128 380 131 390
rect 20 277 23 369
rect 145 366 148 403
rect 151 359 155 855
rect 268 868 272 1075
rect 277 1036 280 1068
rect 291 1051 294 1061
rect 277 1021 280 1030
rect 298 1021 301 1030
rect 314 1023 317 1036
rect 327 1008 330 1061
rect 394 1051 397 1061
rect 334 1036 338 1040
rect 335 1021 338 1030
rect 290 994 293 1006
rect 331 1004 332 1008
rect 341 994 344 1047
rect 409 1036 412 1083
rect 347 1027 350 1032
rect 356 1021 359 1030
rect 372 1023 375 1036
rect 393 1021 396 1030
rect 409 1028 412 1032
rect 417 1058 423 1194
rect 409 1021 412 1024
rect 392 994 395 1004
rect 417 979 423 1054
rect 417 946 423 975
rect 277 916 280 918
rect 277 909 280 912
rect 277 875 280 905
rect 417 902 423 942
rect 158 837 161 847
rect 159 807 162 816
rect 180 809 183 822
rect 196 807 199 816
rect 205 813 208 818
rect 160 780 163 790
rect 211 780 214 833
rect 217 822 221 826
rect 217 807 220 816
rect 225 794 228 847
rect 261 837 264 847
rect 238 809 241 822
rect 254 807 257 816
rect 223 790 224 794
rect 262 780 265 792
rect 159 437 162 447
rect 166 407 169 416
rect 182 409 185 422
rect 195 394 198 447
rect 262 437 265 447
rect 202 422 206 426
rect 203 407 206 416
rect 158 380 161 392
rect 199 390 200 394
rect 209 380 212 433
rect 215 413 218 418
rect 224 407 227 416
rect 240 409 243 422
rect 261 407 264 416
rect 260 380 263 390
rect 135 348 139 351
rect 135 329 139 344
rect 151 341 155 355
rect 167 355 171 359
rect 167 348 171 351
rect 167 329 171 344
rect 151 325 155 326
rect 167 321 171 325
rect 27 297 30 307
rect 34 267 37 276
rect 50 269 53 282
rect 63 254 66 307
rect 130 297 133 307
rect 70 282 74 286
rect 71 267 74 276
rect 26 240 29 252
rect 67 250 68 254
rect 77 240 80 293
rect 145 282 148 314
rect 83 273 86 278
rect 92 267 95 276
rect 108 269 111 282
rect 129 267 132 276
rect 145 267 148 276
rect 128 240 131 250
rect 20 191 23 229
rect 27 211 30 221
rect 34 181 37 190
rect 50 183 53 196
rect 63 168 66 221
rect 130 211 133 221
rect 70 196 74 200
rect 71 181 74 190
rect 26 154 29 166
rect 67 164 68 168
rect 77 154 80 207
rect 83 187 86 192
rect 92 181 95 190
rect 108 183 111 196
rect 129 181 132 190
rect 145 181 148 190
rect 128 154 131 164
rect 20 51 23 143
rect 145 140 148 177
rect 27 71 30 81
rect 34 41 37 50
rect 50 43 53 56
rect 63 28 66 81
rect 130 71 133 81
rect 70 56 74 60
rect 71 41 74 50
rect 26 14 29 26
rect 67 24 68 28
rect 77 14 80 67
rect 145 56 148 88
rect 83 47 86 52
rect 92 41 95 50
rect 108 43 111 56
rect 129 41 132 50
rect 145 41 148 50
rect 128 14 131 24
rect 151 0 155 321
rect 159 297 162 307
rect 166 267 169 276
rect 182 269 185 282
rect 195 254 198 307
rect 262 297 265 307
rect 202 282 206 286
rect 203 267 206 276
rect 158 240 161 252
rect 199 250 200 254
rect 209 240 212 293
rect 215 273 218 278
rect 224 267 227 276
rect 240 269 243 282
rect 261 267 264 276
rect 260 240 263 250
rect 159 211 162 221
rect 166 181 169 190
rect 182 183 185 196
rect 195 168 198 221
rect 262 211 265 221
rect 202 196 206 200
rect 203 181 206 190
rect 158 154 161 166
rect 199 164 200 168
rect 209 154 212 207
rect 215 187 218 192
rect 224 181 227 190
rect 240 183 243 196
rect 261 181 264 190
rect 260 154 263 164
rect 268 133 272 864
rect 292 859 296 864
rect 417 844 423 898
rect 417 770 423 840
rect 417 638 423 766
rect 417 506 423 634
rect 291 437 294 447
rect 277 407 280 416
rect 298 407 301 416
rect 314 409 317 422
rect 277 366 280 403
rect 327 394 330 447
rect 394 437 397 447
rect 417 444 423 502
rect 334 422 338 426
rect 335 407 338 416
rect 290 380 293 392
rect 331 390 332 394
rect 341 380 344 433
rect 347 413 350 418
rect 356 407 359 416
rect 372 409 375 422
rect 393 407 396 416
rect 409 407 412 418
rect 392 380 395 390
rect 409 373 412 403
rect 409 341 412 369
rect 417 374 423 440
rect 417 334 423 370
rect 277 282 280 314
rect 291 297 294 307
rect 277 267 280 276
rect 298 267 301 276
rect 314 269 317 282
rect 327 254 330 307
rect 394 297 397 307
rect 334 282 338 286
rect 335 267 338 276
rect 290 240 293 252
rect 331 250 332 254
rect 341 240 344 293
rect 409 282 412 329
rect 347 273 350 278
rect 356 267 359 276
rect 372 269 375 282
rect 393 267 396 276
rect 409 267 412 278
rect 392 240 395 250
rect 409 233 412 263
rect 417 304 423 330
rect 291 211 294 221
rect 277 181 280 190
rect 298 181 301 190
rect 314 183 317 196
rect 277 140 280 177
rect 327 168 330 221
rect 394 211 397 221
rect 417 218 423 300
rect 334 196 338 200
rect 335 181 338 190
rect 290 154 293 166
rect 331 164 332 168
rect 341 154 344 207
rect 347 187 350 192
rect 356 181 359 190
rect 372 183 375 196
rect 393 181 396 190
rect 409 181 412 192
rect 392 154 395 164
rect 409 147 412 177
rect 252 122 256 125
rect 252 103 256 118
rect 268 115 272 129
rect 284 129 288 133
rect 284 122 288 125
rect 284 103 288 118
rect 409 115 412 143
rect 268 99 272 100
rect 284 95 288 99
rect 159 71 162 81
rect 166 41 169 50
rect 182 43 185 56
rect 195 28 198 81
rect 262 71 265 81
rect 202 56 206 60
rect 203 41 206 50
rect 158 14 161 26
rect 199 24 200 28
rect 209 14 212 67
rect 215 47 218 52
rect 224 41 227 50
rect 240 43 243 56
rect 261 41 264 50
rect 260 14 263 24
rect 268 0 272 95
rect 277 56 280 88
rect 291 71 294 81
rect 277 41 280 50
rect 298 41 301 50
rect 314 43 317 56
rect 327 28 330 81
rect 394 71 397 81
rect 334 56 338 60
rect 335 41 338 50
rect 290 14 293 26
rect 331 24 332 28
rect 341 14 344 67
rect 409 56 412 103
rect 347 47 350 52
rect 356 41 359 50
rect 372 43 375 56
rect 393 41 396 50
rect 409 48 412 52
rect 417 78 423 214
rect 409 41 412 44
rect 392 14 395 24
rect 417 0 423 74
rect 429 1902 435 1973
rect 429 1869 435 1898
rect 429 1816 435 1865
rect 429 1767 435 1812
rect 429 1684 435 1763
rect 429 1552 435 1680
rect 429 1420 435 1548
rect 429 1367 435 1416
rect 429 1257 435 1363
rect 429 1227 435 1253
rect 429 1171 435 1223
rect 429 1141 435 1167
rect 429 1001 435 1137
rect 429 922 435 997
rect 429 889 435 918
rect 429 836 435 885
rect 429 787 435 832
rect 429 704 435 783
rect 429 572 435 700
rect 429 440 435 568
rect 429 387 435 436
rect 429 277 435 383
rect 429 247 435 273
rect 429 191 435 243
rect 429 161 435 187
rect 429 21 435 157
rect 429 0 435 17
rect 441 1823 447 1973
rect 441 1809 447 1819
rect 441 1691 447 1805
rect 441 1677 447 1687
rect 441 1559 447 1673
rect 441 1545 447 1555
rect 441 1413 447 1541
rect 441 1339 447 1409
rect 441 843 447 1335
rect 441 829 447 839
rect 441 711 447 825
rect 441 697 447 707
rect 441 579 447 693
rect 441 565 447 575
rect 441 433 447 561
rect 441 359 447 429
rect 441 0 447 355
rect 453 1875 459 1973
rect 453 1743 459 1871
rect 453 1625 459 1739
rect 453 1611 459 1621
rect 453 1493 459 1607
rect 453 1479 459 1489
rect 453 1347 459 1475
rect 453 895 459 1343
rect 453 763 459 891
rect 453 645 459 759
rect 453 631 459 641
rect 453 513 459 627
rect 453 499 459 509
rect 453 367 459 495
rect 453 0 459 363
rect 465 1895 471 1973
rect 465 1862 471 1891
rect 465 1760 471 1858
rect 465 1361 471 1756
rect 465 1250 471 1357
rect 465 1220 471 1246
rect 465 1164 471 1216
rect 465 1134 471 1160
rect 465 994 471 1130
rect 465 915 471 990
rect 465 882 471 911
rect 465 780 471 878
rect 465 381 471 776
rect 465 270 471 377
rect 465 240 471 266
rect 465 184 471 236
rect 465 154 471 180
rect 465 14 471 150
rect 465 0 471 10
rect 477 1966 483 1973
rect 477 1933 483 1962
rect 499 1952 502 1962
rect 477 1831 483 1929
rect 506 1922 509 1931
rect 522 1924 525 1937
rect 535 1909 538 1962
rect 602 1952 605 1962
rect 631 1952 634 1962
rect 542 1937 546 1941
rect 543 1922 546 1931
rect 498 1895 501 1907
rect 539 1905 540 1909
rect 549 1895 552 1948
rect 555 1928 558 1933
rect 564 1922 567 1931
rect 580 1924 583 1937
rect 601 1922 604 1931
rect 617 1931 620 1933
rect 617 1928 624 1931
rect 617 1922 620 1928
rect 638 1922 641 1931
rect 654 1924 657 1937
rect 600 1895 603 1905
rect 617 1888 620 1918
rect 667 1909 670 1962
rect 734 1952 737 1962
rect 763 1952 766 1962
rect 674 1937 678 1941
rect 675 1922 678 1931
rect 630 1895 633 1907
rect 671 1905 672 1909
rect 681 1895 684 1948
rect 687 1928 690 1933
rect 696 1922 699 1931
rect 712 1924 715 1937
rect 733 1922 736 1931
rect 749 1931 752 1933
rect 749 1928 756 1931
rect 749 1922 752 1928
rect 770 1922 773 1931
rect 786 1924 789 1937
rect 732 1895 735 1905
rect 617 1885 669 1888
rect 497 1865 500 1878
rect 523 1868 526 1871
rect 530 1865 533 1878
rect 547 1865 550 1878
rect 477 1431 483 1827
rect 497 1816 500 1831
rect 511 1823 514 1827
rect 529 1816 532 1831
rect 548 1816 551 1831
rect 554 1830 557 1871
rect 570 1823 573 1864
rect 576 1831 579 1871
rect 595 1823 598 1864
rect 604 1865 607 1878
rect 620 1865 623 1878
rect 641 1868 644 1871
rect 648 1865 651 1878
rect 666 1874 669 1885
rect 749 1882 752 1918
rect 799 1909 802 1962
rect 866 1952 869 1962
rect 895 1952 898 1962
rect 806 1937 810 1941
rect 807 1922 810 1931
rect 762 1895 765 1907
rect 803 1905 804 1909
rect 813 1895 816 1948
rect 819 1928 822 1933
rect 828 1922 831 1931
rect 844 1924 847 1937
rect 865 1922 868 1931
rect 881 1931 884 1933
rect 881 1928 888 1931
rect 881 1922 884 1928
rect 902 1922 905 1931
rect 918 1924 921 1937
rect 864 1895 867 1905
rect 881 1888 884 1910
rect 931 1909 934 1962
rect 998 1952 1001 1962
rect 938 1937 942 1941
rect 939 1922 942 1931
rect 894 1895 897 1907
rect 935 1905 936 1909
rect 945 1895 948 1948
rect 951 1928 954 1933
rect 960 1922 963 1931
rect 976 1924 979 1937
rect 997 1922 1000 1931
rect 1013 1931 1016 1933
rect 1013 1928 1017 1931
rect 1013 1922 1016 1928
rect 1013 1914 1016 1918
rect 996 1895 999 1905
rect 747 1877 752 1882
rect 809 1884 884 1888
rect 666 1871 711 1874
rect 666 1861 669 1871
rect 684 1858 704 1861
rect 701 1839 704 1858
rect 604 1816 607 1831
rect 619 1816 622 1831
rect 626 1823 630 1826
rect 647 1816 650 1831
rect 497 1797 500 1812
rect 511 1801 514 1805
rect 529 1797 532 1812
rect 548 1797 551 1812
rect 497 1750 500 1763
rect 523 1757 526 1760
rect 497 1733 500 1746
rect 507 1743 511 1753
rect 530 1750 533 1763
rect 547 1750 550 1763
rect 554 1757 557 1798
rect 570 1764 573 1805
rect 576 1757 579 1797
rect 595 1764 598 1805
rect 604 1797 607 1812
rect 619 1797 622 1812
rect 626 1802 630 1805
rect 647 1797 650 1812
rect 604 1750 607 1763
rect 523 1736 526 1739
rect 530 1733 533 1746
rect 547 1733 550 1746
rect 497 1684 500 1699
rect 511 1691 514 1695
rect 529 1684 532 1699
rect 548 1684 551 1699
rect 554 1698 557 1739
rect 570 1691 573 1732
rect 576 1699 579 1739
rect 595 1691 598 1732
rect 604 1733 607 1746
rect 620 1750 623 1763
rect 641 1757 644 1760
rect 648 1750 651 1763
rect 701 1763 704 1835
rect 712 1799 715 1871
rect 747 1874 750 1877
rect 747 1871 792 1874
rect 747 1861 750 1871
rect 620 1733 623 1746
rect 641 1736 644 1739
rect 648 1733 651 1746
rect 701 1729 704 1759
rect 712 1743 715 1795
rect 719 1783 723 1849
rect 707 1739 711 1742
rect 700 1726 704 1729
rect 701 1707 704 1726
rect 604 1684 607 1699
rect 619 1684 622 1699
rect 626 1691 630 1694
rect 647 1684 650 1699
rect 497 1665 500 1680
rect 511 1669 514 1673
rect 529 1665 532 1680
rect 548 1665 551 1680
rect 497 1618 500 1631
rect 523 1625 526 1628
rect 497 1601 500 1614
rect 530 1618 533 1631
rect 547 1618 550 1631
rect 554 1625 557 1666
rect 570 1632 573 1673
rect 576 1625 579 1665
rect 595 1632 598 1673
rect 604 1665 607 1680
rect 619 1665 622 1680
rect 626 1670 630 1673
rect 647 1665 650 1680
rect 604 1618 607 1631
rect 523 1604 526 1607
rect 530 1601 533 1614
rect 547 1601 550 1614
rect 497 1552 500 1567
rect 511 1559 514 1563
rect 529 1552 532 1567
rect 548 1552 551 1567
rect 554 1566 557 1607
rect 570 1559 573 1600
rect 576 1567 579 1607
rect 595 1559 598 1600
rect 604 1601 607 1614
rect 620 1618 623 1631
rect 641 1625 644 1628
rect 648 1618 651 1631
rect 701 1632 704 1703
rect 712 1668 715 1739
rect 620 1601 623 1614
rect 641 1604 644 1607
rect 648 1601 651 1614
rect 701 1575 704 1628
rect 712 1611 715 1664
rect 719 1652 723 1717
rect 707 1607 711 1610
rect 750 1610 753 1861
rect 765 1858 785 1861
rect 782 1839 785 1858
rect 782 1763 785 1835
rect 793 1799 796 1871
rect 800 1783 804 1849
rect 809 1750 812 1884
rect 1013 1881 1016 1910
rect 837 1878 944 1881
rect 771 1746 812 1750
rect 771 1742 774 1746
rect 771 1739 816 1742
rect 771 1729 774 1739
rect 789 1726 809 1729
rect 771 1724 774 1725
rect 806 1707 809 1726
rect 806 1632 809 1703
rect 817 1668 820 1739
rect 824 1652 828 1717
rect 604 1552 607 1567
rect 619 1552 622 1567
rect 626 1559 630 1562
rect 647 1552 650 1567
rect 497 1533 500 1548
rect 511 1537 514 1541
rect 529 1533 532 1548
rect 548 1533 551 1548
rect 497 1486 500 1499
rect 523 1493 526 1496
rect 497 1469 500 1482
rect 530 1486 533 1499
rect 547 1486 550 1499
rect 554 1493 557 1534
rect 570 1500 573 1541
rect 576 1493 579 1533
rect 595 1500 598 1541
rect 604 1533 607 1548
rect 619 1533 622 1548
rect 626 1538 630 1541
rect 647 1533 650 1548
rect 604 1486 607 1499
rect 523 1472 526 1475
rect 530 1469 533 1482
rect 547 1469 550 1482
rect 477 1321 483 1427
rect 497 1420 500 1435
rect 511 1427 514 1431
rect 497 1401 500 1416
rect 520 1413 524 1423
rect 529 1420 532 1435
rect 548 1420 551 1435
rect 554 1434 557 1475
rect 570 1427 573 1468
rect 576 1435 579 1475
rect 595 1427 598 1468
rect 604 1469 607 1482
rect 620 1486 623 1499
rect 641 1493 644 1496
rect 648 1486 651 1499
rect 701 1497 704 1571
rect 712 1533 715 1607
rect 747 1607 792 1610
rect 747 1597 750 1607
rect 765 1594 785 1597
rect 620 1469 623 1482
rect 641 1472 644 1475
rect 648 1469 651 1482
rect 701 1443 704 1493
rect 712 1479 715 1529
rect 719 1517 723 1585
rect 782 1575 785 1594
rect 782 1497 785 1571
rect 793 1533 796 1607
rect 837 1610 840 1878
rect 948 1878 1016 1881
rect 1076 1846 1079 1895
rect 1076 1802 1079 1842
rect 1084 1839 1088 1982
rect 1092 1919 1095 1929
rect 1099 1889 1102 1898
rect 1115 1891 1118 1904
rect 1128 1876 1131 1929
rect 1195 1919 1198 1929
rect 1135 1904 1139 1908
rect 1136 1889 1139 1898
rect 1091 1862 1094 1874
rect 1132 1872 1133 1876
rect 1142 1862 1145 1915
rect 1148 1895 1151 1900
rect 1157 1889 1160 1898
rect 1173 1891 1176 1904
rect 1194 1889 1197 1898
rect 1193 1862 1196 1872
rect 1076 1787 1079 1796
rect 837 1607 882 1610
rect 837 1597 840 1607
rect 855 1594 875 1597
rect 800 1517 804 1585
rect 872 1575 875 1594
rect 872 1497 875 1571
rect 883 1533 886 1607
rect 890 1517 894 1585
rect 707 1475 711 1478
rect 604 1420 607 1435
rect 619 1420 622 1435
rect 626 1427 630 1430
rect 647 1420 650 1435
rect 511 1405 514 1409
rect 529 1401 532 1416
rect 548 1401 551 1416
rect 497 1354 500 1367
rect 523 1361 526 1364
rect 505 1347 509 1357
rect 530 1354 533 1367
rect 547 1354 550 1367
rect 554 1361 557 1402
rect 570 1368 573 1409
rect 576 1361 579 1401
rect 595 1368 598 1409
rect 604 1401 607 1416
rect 619 1401 622 1416
rect 626 1406 630 1409
rect 647 1401 650 1416
rect 604 1354 607 1367
rect 620 1354 623 1367
rect 641 1361 644 1364
rect 648 1354 651 1367
rect 701 1361 704 1439
rect 712 1397 715 1475
rect 719 1381 723 1453
rect 731 1354 735 1367
rect 740 1347 743 1357
rect 750 1340 753 1409
rect 772 1405 775 1409
rect 790 1401 793 1416
rect 809 1401 812 1416
rect 757 1354 761 1367
rect 784 1361 787 1364
rect 791 1354 794 1367
rect 808 1354 811 1367
rect 815 1361 818 1402
rect 831 1368 834 1409
rect 837 1361 840 1401
rect 856 1368 859 1409
rect 865 1401 868 1416
rect 880 1401 883 1416
rect 887 1406 891 1409
rect 908 1401 911 1416
rect 865 1354 868 1367
rect 881 1354 884 1367
rect 902 1361 905 1364
rect 909 1354 912 1367
rect 925 1348 929 1584
rect 960 1417 963 1427
rect 967 1387 970 1396
rect 983 1389 986 1402
rect 996 1374 999 1427
rect 1063 1417 1066 1427
rect 1003 1402 1007 1406
rect 1004 1387 1007 1396
rect 959 1360 962 1372
rect 1000 1370 1001 1374
rect 1010 1360 1013 1413
rect 1016 1393 1019 1398
rect 1025 1387 1028 1396
rect 1041 1389 1044 1402
rect 1062 1387 1065 1396
rect 1078 1387 1081 1396
rect 1061 1360 1064 1370
rect 918 1336 919 1339
rect 477 1291 483 1317
rect 477 1235 483 1287
rect 477 1205 483 1231
rect 783 1228 787 1310
rect 798 1307 801 1317
rect 805 1277 808 1286
rect 821 1279 824 1292
rect 834 1264 837 1317
rect 901 1307 904 1317
rect 841 1292 845 1296
rect 842 1277 845 1286
rect 797 1250 800 1262
rect 838 1260 839 1264
rect 848 1250 851 1303
rect 916 1292 919 1336
rect 854 1283 857 1288
rect 863 1277 866 1286
rect 879 1279 882 1292
rect 900 1277 903 1286
rect 916 1277 919 1286
rect 899 1250 902 1260
rect 916 1243 919 1273
rect 477 1065 483 1201
rect 791 1201 794 1238
rect 798 1221 801 1231
rect 805 1191 808 1200
rect 821 1193 824 1206
rect 834 1178 837 1231
rect 901 1221 904 1231
rect 841 1206 845 1210
rect 842 1191 845 1200
rect 797 1164 800 1176
rect 838 1174 839 1178
rect 848 1164 851 1217
rect 854 1197 857 1202
rect 863 1191 866 1200
rect 879 1193 882 1206
rect 900 1191 903 1200
rect 916 1201 919 1202
rect 937 1204 941 1344
rect 953 1257 956 1349
rect 1078 1346 1081 1383
rect 1084 1339 1088 1835
rect 1201 1848 1205 1982
rect 1350 1959 1356 1973
rect 1350 1926 1356 1955
rect 1210 1896 1213 1898
rect 1210 1889 1213 1892
rect 1210 1855 1213 1885
rect 1350 1882 1356 1922
rect 1091 1817 1094 1827
rect 1092 1787 1095 1796
rect 1113 1789 1116 1802
rect 1129 1787 1132 1796
rect 1138 1793 1141 1798
rect 1093 1760 1096 1770
rect 1144 1760 1147 1813
rect 1150 1802 1154 1806
rect 1150 1787 1153 1796
rect 1158 1774 1161 1827
rect 1194 1817 1197 1827
rect 1171 1789 1174 1802
rect 1187 1787 1190 1796
rect 1156 1770 1157 1774
rect 1195 1760 1198 1772
rect 1092 1417 1095 1427
rect 1099 1387 1102 1396
rect 1115 1389 1118 1402
rect 1128 1374 1131 1427
rect 1195 1417 1198 1427
rect 1135 1402 1139 1406
rect 1136 1387 1139 1396
rect 1091 1360 1094 1372
rect 1132 1370 1133 1374
rect 1142 1360 1145 1413
rect 1148 1393 1151 1398
rect 1157 1387 1160 1396
rect 1173 1389 1176 1402
rect 1194 1387 1197 1396
rect 1193 1360 1196 1370
rect 1068 1328 1072 1331
rect 1068 1309 1072 1324
rect 1084 1321 1088 1335
rect 1100 1335 1104 1339
rect 1100 1328 1104 1331
rect 1100 1309 1104 1324
rect 1084 1305 1088 1306
rect 1100 1301 1104 1305
rect 960 1277 963 1287
rect 967 1247 970 1256
rect 983 1249 986 1262
rect 996 1234 999 1287
rect 1063 1277 1066 1287
rect 1003 1262 1007 1266
rect 1004 1247 1007 1256
rect 959 1220 962 1232
rect 1000 1230 1001 1234
rect 1010 1220 1013 1273
rect 1078 1262 1081 1294
rect 1016 1253 1019 1258
rect 1025 1247 1028 1256
rect 1041 1249 1044 1262
rect 1062 1247 1065 1256
rect 1078 1247 1081 1256
rect 1061 1220 1064 1230
rect 916 1196 919 1197
rect 899 1164 902 1174
rect 937 1102 941 1184
rect 953 1171 956 1209
rect 960 1191 963 1201
rect 967 1161 970 1170
rect 983 1163 986 1176
rect 996 1148 999 1201
rect 1063 1191 1066 1201
rect 1003 1176 1007 1180
rect 1004 1161 1007 1170
rect 959 1134 962 1146
rect 1000 1144 1001 1148
rect 1010 1134 1013 1187
rect 1016 1167 1019 1172
rect 1025 1161 1028 1170
rect 1041 1163 1044 1176
rect 1062 1161 1065 1170
rect 1078 1161 1081 1170
rect 1061 1134 1064 1144
rect 477 986 483 1061
rect 953 1031 956 1123
rect 1078 1120 1081 1157
rect 960 1051 963 1061
rect 967 1021 970 1030
rect 983 1023 986 1036
rect 996 1008 999 1061
rect 1063 1051 1066 1061
rect 1003 1036 1007 1040
rect 1004 1021 1007 1030
rect 959 994 962 1006
rect 1000 1004 1001 1008
rect 1010 994 1013 1047
rect 1078 1036 1081 1068
rect 1016 1027 1019 1032
rect 1025 1021 1028 1030
rect 1041 1023 1044 1036
rect 1062 1021 1065 1030
rect 1078 1021 1081 1030
rect 1061 994 1064 1004
rect 477 953 483 982
rect 499 972 502 982
rect 477 851 483 949
rect 506 942 509 951
rect 522 944 525 957
rect 535 929 538 982
rect 602 972 605 982
rect 631 972 634 982
rect 542 957 546 961
rect 543 942 546 951
rect 498 915 501 927
rect 539 925 540 929
rect 549 915 552 968
rect 555 948 558 953
rect 564 942 567 951
rect 580 944 583 957
rect 601 942 604 951
rect 617 951 620 953
rect 617 948 624 951
rect 617 942 620 948
rect 638 942 641 951
rect 654 944 657 957
rect 600 915 603 925
rect 617 908 620 938
rect 667 929 670 982
rect 734 972 737 982
rect 763 972 766 982
rect 674 957 678 961
rect 675 942 678 951
rect 630 915 633 927
rect 671 925 672 929
rect 681 915 684 968
rect 687 948 690 953
rect 696 942 699 951
rect 712 944 715 957
rect 733 942 736 951
rect 749 951 752 953
rect 749 948 756 951
rect 749 942 752 948
rect 770 942 773 951
rect 786 944 789 957
rect 732 915 735 925
rect 617 905 669 908
rect 497 885 500 898
rect 523 888 526 891
rect 530 885 533 898
rect 547 885 550 898
rect 477 451 483 847
rect 497 836 500 851
rect 511 843 514 847
rect 529 836 532 851
rect 548 836 551 851
rect 554 850 557 891
rect 570 843 573 884
rect 576 851 579 891
rect 595 843 598 884
rect 604 885 607 898
rect 620 885 623 898
rect 641 888 644 891
rect 648 885 651 898
rect 666 894 669 905
rect 749 902 752 938
rect 799 929 802 982
rect 866 972 869 982
rect 895 972 898 982
rect 806 957 810 961
rect 807 942 810 951
rect 762 915 765 927
rect 803 925 804 929
rect 813 915 816 968
rect 819 948 822 953
rect 828 942 831 951
rect 844 944 847 957
rect 865 942 868 951
rect 881 951 884 953
rect 881 948 888 951
rect 881 942 884 948
rect 902 942 905 951
rect 918 944 921 957
rect 864 915 867 925
rect 881 908 884 930
rect 931 929 934 982
rect 998 972 1001 982
rect 938 957 942 961
rect 939 942 942 951
rect 894 915 897 927
rect 935 925 936 929
rect 945 915 948 968
rect 951 948 954 953
rect 960 942 963 951
rect 976 944 979 957
rect 997 942 1000 951
rect 1013 951 1016 953
rect 1013 948 1017 951
rect 1013 942 1016 948
rect 1013 934 1016 938
rect 996 915 999 925
rect 747 897 752 902
rect 809 904 884 908
rect 666 891 711 894
rect 666 881 669 891
rect 684 878 704 881
rect 701 859 704 878
rect 604 836 607 851
rect 619 836 622 851
rect 626 843 630 846
rect 647 836 650 851
rect 497 817 500 832
rect 511 821 514 825
rect 529 817 532 832
rect 548 817 551 832
rect 497 770 500 783
rect 523 777 526 780
rect 497 753 500 766
rect 507 763 511 773
rect 530 770 533 783
rect 547 770 550 783
rect 554 777 557 818
rect 570 784 573 825
rect 576 777 579 817
rect 595 784 598 825
rect 604 817 607 832
rect 619 817 622 832
rect 626 822 630 825
rect 647 817 650 832
rect 604 770 607 783
rect 523 756 526 759
rect 530 753 533 766
rect 547 753 550 766
rect 497 704 500 719
rect 511 711 514 715
rect 529 704 532 719
rect 548 704 551 719
rect 554 718 557 759
rect 570 711 573 752
rect 576 719 579 759
rect 595 711 598 752
rect 604 753 607 766
rect 620 770 623 783
rect 641 777 644 780
rect 648 770 651 783
rect 701 783 704 855
rect 712 819 715 891
rect 747 894 750 897
rect 747 891 792 894
rect 747 881 750 891
rect 620 753 623 766
rect 641 756 644 759
rect 648 753 651 766
rect 701 749 704 779
rect 712 763 715 815
rect 719 803 723 869
rect 707 759 711 762
rect 700 746 704 749
rect 701 727 704 746
rect 604 704 607 719
rect 619 704 622 719
rect 626 711 630 714
rect 647 704 650 719
rect 497 685 500 700
rect 511 689 514 693
rect 529 685 532 700
rect 548 685 551 700
rect 497 638 500 651
rect 523 645 526 648
rect 497 621 500 634
rect 530 638 533 651
rect 547 638 550 651
rect 554 645 557 686
rect 570 652 573 693
rect 576 645 579 685
rect 595 652 598 693
rect 604 685 607 700
rect 619 685 622 700
rect 626 690 630 693
rect 647 685 650 700
rect 604 638 607 651
rect 523 624 526 627
rect 530 621 533 634
rect 547 621 550 634
rect 497 572 500 587
rect 511 579 514 583
rect 529 572 532 587
rect 548 572 551 587
rect 554 586 557 627
rect 570 579 573 620
rect 576 587 579 627
rect 595 579 598 620
rect 604 621 607 634
rect 620 638 623 651
rect 641 645 644 648
rect 648 638 651 651
rect 701 652 704 723
rect 712 688 715 759
rect 620 621 623 634
rect 641 624 644 627
rect 648 621 651 634
rect 701 595 704 648
rect 712 631 715 684
rect 719 672 723 737
rect 707 627 711 630
rect 750 630 753 881
rect 765 878 785 881
rect 782 859 785 878
rect 782 783 785 855
rect 793 819 796 891
rect 800 803 804 869
rect 809 770 812 904
rect 1013 901 1016 930
rect 837 898 944 901
rect 771 766 812 770
rect 771 762 774 766
rect 771 759 816 762
rect 771 749 774 759
rect 789 746 809 749
rect 771 744 774 745
rect 806 727 809 746
rect 806 652 809 723
rect 817 688 820 759
rect 824 672 828 737
rect 604 572 607 587
rect 619 572 622 587
rect 626 579 630 582
rect 647 572 650 587
rect 497 553 500 568
rect 511 557 514 561
rect 529 553 532 568
rect 548 553 551 568
rect 497 506 500 519
rect 523 513 526 516
rect 497 489 500 502
rect 530 506 533 519
rect 547 506 550 519
rect 554 513 557 554
rect 570 520 573 561
rect 576 513 579 553
rect 595 520 598 561
rect 604 553 607 568
rect 619 553 622 568
rect 626 558 630 561
rect 647 553 650 568
rect 604 506 607 519
rect 523 492 526 495
rect 530 489 533 502
rect 547 489 550 502
rect 477 341 483 447
rect 497 440 500 455
rect 511 447 514 451
rect 497 421 500 436
rect 520 433 524 443
rect 529 440 532 455
rect 548 440 551 455
rect 554 454 557 495
rect 570 447 573 488
rect 576 455 579 495
rect 595 447 598 488
rect 604 489 607 502
rect 620 506 623 519
rect 641 513 644 516
rect 648 506 651 519
rect 701 517 704 591
rect 712 553 715 627
rect 747 627 792 630
rect 747 617 750 627
rect 765 614 785 617
rect 620 489 623 502
rect 641 492 644 495
rect 648 489 651 502
rect 701 463 704 513
rect 712 499 715 549
rect 719 537 723 605
rect 782 595 785 614
rect 782 517 785 591
rect 793 553 796 627
rect 837 630 840 898
rect 948 898 1016 901
rect 1076 866 1079 915
rect 1076 822 1079 862
rect 1084 859 1088 1301
rect 1092 1277 1095 1287
rect 1099 1247 1102 1256
rect 1115 1249 1118 1262
rect 1128 1234 1131 1287
rect 1195 1277 1198 1287
rect 1135 1262 1139 1266
rect 1136 1247 1139 1256
rect 1091 1220 1094 1232
rect 1132 1230 1133 1234
rect 1142 1220 1145 1273
rect 1148 1253 1151 1258
rect 1157 1247 1160 1256
rect 1173 1249 1176 1262
rect 1194 1247 1197 1256
rect 1193 1220 1196 1230
rect 1092 1191 1095 1201
rect 1099 1161 1102 1170
rect 1115 1163 1118 1176
rect 1128 1148 1131 1201
rect 1195 1191 1198 1201
rect 1135 1176 1139 1180
rect 1136 1161 1139 1170
rect 1091 1134 1094 1146
rect 1132 1144 1133 1148
rect 1142 1134 1145 1187
rect 1148 1167 1151 1172
rect 1157 1161 1160 1170
rect 1173 1163 1176 1176
rect 1194 1161 1197 1170
rect 1193 1134 1196 1144
rect 1201 1113 1205 1844
rect 1225 1839 1229 1844
rect 1350 1824 1356 1878
rect 1350 1750 1356 1820
rect 1350 1618 1356 1746
rect 1350 1486 1356 1614
rect 1224 1417 1227 1427
rect 1210 1387 1213 1396
rect 1231 1387 1234 1396
rect 1247 1389 1250 1402
rect 1210 1346 1213 1383
rect 1260 1374 1263 1427
rect 1327 1417 1330 1427
rect 1350 1424 1356 1482
rect 1267 1402 1271 1406
rect 1268 1387 1271 1396
rect 1223 1360 1226 1372
rect 1264 1370 1265 1374
rect 1274 1360 1277 1413
rect 1280 1393 1283 1398
rect 1289 1387 1292 1396
rect 1305 1389 1308 1402
rect 1326 1387 1329 1396
rect 1342 1387 1345 1398
rect 1325 1360 1328 1370
rect 1342 1353 1345 1383
rect 1342 1321 1345 1349
rect 1350 1354 1356 1420
rect 1350 1314 1356 1350
rect 1210 1262 1213 1294
rect 1224 1277 1227 1287
rect 1210 1247 1213 1256
rect 1231 1247 1234 1256
rect 1247 1249 1250 1262
rect 1260 1234 1263 1287
rect 1327 1277 1330 1287
rect 1267 1262 1271 1266
rect 1268 1247 1271 1256
rect 1223 1220 1226 1232
rect 1264 1230 1265 1234
rect 1274 1220 1277 1273
rect 1342 1262 1345 1309
rect 1280 1253 1283 1258
rect 1289 1247 1292 1256
rect 1305 1249 1308 1262
rect 1326 1247 1329 1256
rect 1342 1247 1345 1258
rect 1325 1220 1328 1230
rect 1342 1213 1345 1243
rect 1350 1284 1356 1310
rect 1224 1191 1227 1201
rect 1210 1161 1213 1170
rect 1231 1161 1234 1170
rect 1247 1163 1250 1176
rect 1210 1120 1213 1157
rect 1260 1148 1263 1201
rect 1327 1191 1330 1201
rect 1350 1198 1356 1280
rect 1267 1176 1271 1180
rect 1268 1161 1271 1170
rect 1223 1134 1226 1146
rect 1264 1144 1265 1148
rect 1274 1134 1277 1187
rect 1280 1167 1283 1172
rect 1289 1161 1292 1170
rect 1305 1163 1308 1176
rect 1326 1161 1329 1170
rect 1342 1161 1345 1172
rect 1325 1134 1328 1144
rect 1342 1127 1345 1157
rect 1185 1102 1189 1105
rect 1185 1083 1189 1098
rect 1201 1095 1205 1109
rect 1217 1109 1221 1113
rect 1217 1102 1221 1105
rect 1217 1083 1221 1098
rect 1342 1095 1345 1123
rect 1201 1079 1205 1080
rect 1217 1075 1221 1079
rect 1092 1051 1095 1061
rect 1099 1021 1102 1030
rect 1115 1023 1118 1036
rect 1128 1008 1131 1061
rect 1195 1051 1198 1061
rect 1135 1036 1139 1040
rect 1136 1021 1139 1030
rect 1091 994 1094 1006
rect 1132 1004 1133 1008
rect 1142 994 1145 1047
rect 1148 1027 1151 1032
rect 1157 1021 1160 1030
rect 1173 1023 1176 1036
rect 1194 1021 1197 1030
rect 1193 994 1196 1004
rect 1092 939 1095 949
rect 1099 909 1102 918
rect 1115 911 1118 924
rect 1128 896 1131 949
rect 1195 939 1198 949
rect 1135 924 1139 928
rect 1136 909 1139 918
rect 1091 882 1094 894
rect 1132 892 1133 896
rect 1142 882 1145 935
rect 1148 915 1151 920
rect 1157 909 1160 918
rect 1173 911 1176 924
rect 1194 909 1197 918
rect 1193 882 1196 892
rect 1076 807 1079 816
rect 837 627 882 630
rect 837 617 840 627
rect 855 614 875 617
rect 800 537 804 605
rect 872 595 875 614
rect 872 517 875 591
rect 883 553 886 627
rect 890 537 894 605
rect 707 495 711 498
rect 604 440 607 455
rect 619 440 622 455
rect 626 447 630 450
rect 647 440 650 455
rect 511 425 514 429
rect 529 421 532 436
rect 548 421 551 436
rect 497 374 500 387
rect 523 381 526 384
rect 505 367 509 377
rect 530 374 533 387
rect 547 374 550 387
rect 554 381 557 422
rect 570 388 573 429
rect 576 381 579 421
rect 595 388 598 429
rect 604 421 607 436
rect 619 421 622 436
rect 626 426 630 429
rect 647 421 650 436
rect 604 374 607 387
rect 620 374 623 387
rect 641 381 644 384
rect 648 374 651 387
rect 701 381 704 459
rect 712 417 715 495
rect 719 401 723 473
rect 731 374 735 387
rect 740 367 743 377
rect 750 360 753 429
rect 772 425 775 429
rect 790 421 793 436
rect 809 421 812 436
rect 757 374 761 387
rect 784 381 787 384
rect 791 374 794 387
rect 808 374 811 387
rect 815 381 818 422
rect 831 388 834 429
rect 837 381 840 421
rect 856 388 859 429
rect 865 421 868 436
rect 880 421 883 436
rect 887 426 891 429
rect 908 421 911 436
rect 865 374 868 387
rect 881 374 884 387
rect 902 381 905 384
rect 909 374 912 387
rect 925 368 929 604
rect 960 437 963 447
rect 967 407 970 416
rect 983 409 986 422
rect 996 394 999 447
rect 1063 437 1066 447
rect 1003 422 1007 426
rect 1004 407 1007 416
rect 959 380 962 392
rect 1000 390 1001 394
rect 1010 380 1013 433
rect 1016 413 1019 418
rect 1025 407 1028 416
rect 1041 409 1044 422
rect 1062 407 1065 416
rect 1078 407 1081 416
rect 1061 380 1064 390
rect 918 356 919 359
rect 477 311 483 337
rect 477 255 483 307
rect 477 225 483 251
rect 783 248 787 330
rect 798 327 801 337
rect 805 297 808 306
rect 821 299 824 312
rect 834 284 837 337
rect 901 327 904 337
rect 841 312 845 316
rect 842 297 845 306
rect 797 270 800 282
rect 838 280 839 284
rect 848 270 851 323
rect 916 312 919 356
rect 854 303 857 308
rect 863 297 866 306
rect 879 299 882 312
rect 900 297 903 306
rect 916 297 919 306
rect 899 270 902 280
rect 916 263 919 293
rect 477 85 483 221
rect 791 221 794 258
rect 798 241 801 251
rect 805 211 808 220
rect 821 213 824 226
rect 834 198 837 251
rect 901 241 904 251
rect 841 226 845 230
rect 842 211 845 220
rect 797 184 800 196
rect 838 194 839 198
rect 848 184 851 237
rect 854 217 857 222
rect 863 211 866 220
rect 879 213 882 226
rect 900 211 903 220
rect 916 221 919 222
rect 937 224 941 364
rect 953 277 956 369
rect 1078 366 1081 403
rect 1084 359 1088 855
rect 1201 868 1205 1075
rect 1210 1036 1213 1068
rect 1224 1051 1227 1061
rect 1210 1021 1213 1030
rect 1231 1021 1234 1030
rect 1247 1023 1250 1036
rect 1260 1008 1263 1061
rect 1327 1051 1330 1061
rect 1267 1036 1271 1040
rect 1268 1021 1271 1030
rect 1223 994 1226 1006
rect 1264 1004 1265 1008
rect 1274 994 1277 1047
rect 1342 1036 1345 1083
rect 1280 1027 1283 1032
rect 1289 1021 1292 1030
rect 1305 1023 1308 1036
rect 1326 1021 1329 1030
rect 1342 1028 1345 1032
rect 1350 1058 1356 1194
rect 1342 1021 1345 1024
rect 1325 994 1328 1004
rect 1350 979 1356 1054
rect 1350 946 1356 975
rect 1210 917 1213 918
rect 1210 912 1214 913
rect 1210 909 1213 912
rect 1210 875 1213 905
rect 1350 902 1356 942
rect 1091 837 1094 847
rect 1092 807 1095 816
rect 1113 809 1116 822
rect 1129 807 1132 816
rect 1138 813 1141 818
rect 1093 780 1096 790
rect 1144 780 1147 833
rect 1150 822 1154 826
rect 1150 807 1153 816
rect 1158 794 1161 847
rect 1194 837 1197 847
rect 1171 809 1174 822
rect 1187 807 1190 816
rect 1156 790 1157 794
rect 1195 780 1198 792
rect 1092 437 1095 447
rect 1099 407 1102 416
rect 1115 409 1118 422
rect 1128 394 1131 447
rect 1195 437 1198 447
rect 1135 422 1139 426
rect 1136 407 1139 416
rect 1091 380 1094 392
rect 1132 390 1133 394
rect 1142 380 1145 433
rect 1148 413 1151 418
rect 1157 407 1160 416
rect 1173 409 1176 422
rect 1194 407 1197 416
rect 1193 380 1196 390
rect 1068 348 1072 351
rect 1068 329 1072 344
rect 1084 341 1088 355
rect 1100 355 1104 359
rect 1100 348 1104 351
rect 1100 329 1104 344
rect 1084 325 1088 326
rect 1100 321 1104 325
rect 960 297 963 307
rect 967 267 970 276
rect 983 269 986 282
rect 996 254 999 307
rect 1063 297 1066 307
rect 1003 282 1007 286
rect 1004 267 1007 276
rect 959 240 962 252
rect 1000 250 1001 254
rect 1010 240 1013 293
rect 1078 282 1081 314
rect 1016 273 1019 278
rect 1025 267 1028 276
rect 1041 269 1044 282
rect 1062 267 1065 276
rect 1078 267 1081 276
rect 1061 240 1064 250
rect 916 216 919 217
rect 899 184 902 194
rect 937 122 941 204
rect 953 191 956 229
rect 960 211 963 221
rect 967 181 970 190
rect 983 183 986 196
rect 996 168 999 221
rect 1063 211 1066 221
rect 1003 196 1007 200
rect 1004 181 1007 190
rect 959 154 962 166
rect 1000 164 1001 168
rect 1010 154 1013 207
rect 1016 187 1019 192
rect 1025 181 1028 190
rect 1041 183 1044 196
rect 1062 181 1065 190
rect 1078 181 1081 190
rect 1061 154 1064 164
rect 477 0 483 81
rect 953 51 956 143
rect 1078 140 1081 177
rect 960 71 963 81
rect 967 41 970 50
rect 983 43 986 56
rect 996 28 999 81
rect 1063 71 1066 81
rect 1003 56 1007 60
rect 1004 41 1007 50
rect 959 14 962 26
rect 1000 24 1001 28
rect 1010 14 1013 67
rect 1078 56 1081 88
rect 1016 47 1019 52
rect 1025 41 1028 50
rect 1041 43 1044 56
rect 1062 41 1065 50
rect 1078 41 1081 50
rect 1061 14 1064 24
rect 1084 0 1088 321
rect 1092 297 1095 307
rect 1099 267 1102 276
rect 1115 269 1118 282
rect 1128 254 1131 307
rect 1195 297 1198 307
rect 1135 282 1139 286
rect 1136 267 1139 276
rect 1091 240 1094 252
rect 1132 250 1133 254
rect 1142 240 1145 293
rect 1148 273 1151 278
rect 1157 267 1160 276
rect 1173 269 1176 282
rect 1194 267 1197 276
rect 1193 240 1196 250
rect 1092 211 1095 221
rect 1099 181 1102 190
rect 1115 183 1118 196
rect 1128 168 1131 221
rect 1195 211 1198 221
rect 1135 196 1139 200
rect 1136 181 1139 190
rect 1091 154 1094 166
rect 1132 164 1133 168
rect 1142 154 1145 207
rect 1148 187 1151 192
rect 1157 181 1160 190
rect 1173 183 1176 196
rect 1194 181 1197 190
rect 1193 154 1196 164
rect 1201 133 1205 864
rect 1225 859 1229 864
rect 1350 844 1356 898
rect 1350 770 1356 840
rect 1350 638 1356 766
rect 1350 506 1356 634
rect 1224 437 1227 447
rect 1210 407 1213 416
rect 1231 407 1234 416
rect 1247 409 1250 422
rect 1210 366 1213 403
rect 1260 394 1263 447
rect 1327 437 1330 447
rect 1350 444 1356 502
rect 1267 422 1271 426
rect 1268 407 1271 416
rect 1223 380 1226 392
rect 1264 390 1265 394
rect 1274 380 1277 433
rect 1280 413 1283 418
rect 1289 407 1292 416
rect 1305 409 1308 422
rect 1326 407 1329 416
rect 1342 407 1345 418
rect 1325 380 1328 390
rect 1342 373 1345 403
rect 1342 341 1345 369
rect 1350 374 1356 440
rect 1350 334 1356 370
rect 1210 282 1213 314
rect 1224 297 1227 307
rect 1210 267 1213 276
rect 1231 267 1234 276
rect 1247 269 1250 282
rect 1260 254 1263 307
rect 1327 297 1330 307
rect 1267 282 1271 286
rect 1268 267 1271 276
rect 1223 240 1226 252
rect 1264 250 1265 254
rect 1274 240 1277 293
rect 1342 282 1345 329
rect 1280 273 1283 278
rect 1289 267 1292 276
rect 1305 269 1308 282
rect 1326 267 1329 276
rect 1342 267 1345 278
rect 1325 240 1328 250
rect 1342 233 1345 263
rect 1350 304 1356 330
rect 1224 211 1227 221
rect 1210 181 1213 190
rect 1231 181 1234 190
rect 1247 183 1250 196
rect 1210 140 1213 177
rect 1260 168 1263 221
rect 1327 211 1330 221
rect 1350 218 1356 300
rect 1267 196 1271 200
rect 1268 181 1271 190
rect 1223 154 1226 166
rect 1264 164 1265 168
rect 1274 154 1277 207
rect 1280 187 1283 192
rect 1289 181 1292 190
rect 1305 183 1308 196
rect 1326 181 1329 190
rect 1342 181 1345 192
rect 1325 154 1328 164
rect 1342 147 1345 177
rect 1185 122 1189 125
rect 1185 103 1189 118
rect 1201 115 1205 129
rect 1217 129 1221 133
rect 1217 122 1221 125
rect 1217 103 1221 118
rect 1342 115 1345 143
rect 1201 99 1205 100
rect 1217 95 1221 99
rect 1092 71 1095 81
rect 1099 41 1102 50
rect 1115 43 1118 56
rect 1128 28 1131 81
rect 1195 71 1198 81
rect 1135 56 1139 60
rect 1136 41 1139 50
rect 1091 14 1094 26
rect 1132 24 1133 28
rect 1142 14 1145 67
rect 1148 47 1151 52
rect 1157 41 1160 50
rect 1173 43 1176 56
rect 1194 41 1197 50
rect 1193 14 1196 24
rect 1201 0 1205 95
rect 1210 56 1213 88
rect 1224 71 1227 81
rect 1210 41 1213 50
rect 1231 41 1234 50
rect 1247 43 1250 56
rect 1260 28 1263 81
rect 1327 71 1330 81
rect 1267 56 1271 60
rect 1268 41 1271 50
rect 1223 14 1226 26
rect 1264 24 1265 28
rect 1274 14 1277 67
rect 1342 56 1345 103
rect 1280 47 1283 52
rect 1289 41 1292 50
rect 1305 43 1308 56
rect 1326 41 1329 50
rect 1342 48 1345 52
rect 1350 78 1356 214
rect 1342 41 1345 44
rect 1325 14 1328 24
rect 1350 0 1356 74
rect 1362 1902 1368 1973
rect 1362 1869 1368 1898
rect 1362 1816 1368 1865
rect 1362 1767 1368 1812
rect 1362 1684 1368 1763
rect 1362 1552 1368 1680
rect 1362 1420 1368 1548
rect 1362 1367 1368 1416
rect 1362 1257 1368 1363
rect 1362 1227 1368 1253
rect 1362 1171 1368 1223
rect 1362 1141 1368 1167
rect 1362 1001 1368 1137
rect 1362 922 1368 997
rect 1362 889 1368 918
rect 1362 836 1368 885
rect 1362 787 1368 832
rect 1362 704 1368 783
rect 1362 572 1368 700
rect 1362 440 1368 568
rect 1362 387 1368 436
rect 1362 277 1368 383
rect 1362 247 1368 273
rect 1362 191 1368 243
rect 1362 161 1368 187
rect 1362 21 1368 157
rect 1362 0 1368 17
rect 1374 1823 1380 1973
rect 1374 1809 1380 1819
rect 1374 1691 1380 1805
rect 1374 1677 1380 1687
rect 1374 1559 1380 1673
rect 1374 1545 1380 1555
rect 1374 1413 1380 1541
rect 1374 1339 1380 1409
rect 1374 843 1380 1335
rect 1374 829 1380 839
rect 1374 711 1380 825
rect 1374 697 1380 707
rect 1374 579 1380 693
rect 1374 565 1380 575
rect 1374 433 1380 561
rect 1374 359 1380 429
rect 1374 0 1380 355
rect 1386 1875 1392 1973
rect 1386 1743 1392 1871
rect 1386 1625 1392 1739
rect 1386 1611 1392 1621
rect 1386 1493 1392 1607
rect 1386 1479 1392 1489
rect 1386 1347 1392 1475
rect 1386 895 1392 1343
rect 1386 763 1392 891
rect 1386 645 1392 759
rect 1386 631 1392 641
rect 1386 513 1392 627
rect 1386 499 1392 509
rect 1386 367 1392 495
rect 1386 0 1392 363
rect 1398 1895 1404 1973
rect 1398 1862 1404 1891
rect 1398 1760 1404 1858
rect 1398 1361 1404 1756
rect 1398 1250 1404 1357
rect 1398 1220 1404 1246
rect 1398 1164 1404 1216
rect 1398 1134 1404 1160
rect 1398 994 1404 1130
rect 1398 915 1404 990
rect 1398 882 1404 911
rect 1398 780 1404 878
rect 1398 381 1404 776
rect 1398 270 1404 377
rect 1398 240 1404 266
rect 1398 184 1404 236
rect 1398 154 1404 180
rect 1398 14 1404 150
rect 1398 0 1404 10
rect 1410 1966 1416 1973
rect 1410 1933 1416 1962
rect 1432 1952 1435 1962
rect 1410 1831 1416 1929
rect 1439 1922 1442 1931
rect 1455 1924 1458 1937
rect 1468 1909 1471 1962
rect 1535 1952 1538 1962
rect 1564 1952 1567 1962
rect 1475 1937 1479 1941
rect 1476 1922 1479 1931
rect 1431 1895 1434 1907
rect 1472 1905 1473 1909
rect 1482 1895 1485 1948
rect 1488 1928 1491 1933
rect 1497 1922 1500 1931
rect 1513 1924 1516 1937
rect 1534 1922 1537 1931
rect 1550 1931 1553 1933
rect 1550 1928 1557 1931
rect 1550 1922 1553 1928
rect 1571 1922 1574 1931
rect 1587 1924 1590 1937
rect 1533 1895 1536 1905
rect 1550 1888 1553 1918
rect 1600 1909 1603 1962
rect 1667 1952 1670 1962
rect 1696 1952 1699 1962
rect 1607 1937 1611 1941
rect 1608 1922 1611 1931
rect 1563 1895 1566 1907
rect 1604 1905 1605 1909
rect 1614 1895 1617 1948
rect 1620 1928 1623 1933
rect 1629 1922 1632 1931
rect 1645 1924 1648 1937
rect 1666 1922 1669 1931
rect 1682 1931 1685 1933
rect 1682 1928 1689 1931
rect 1682 1922 1685 1928
rect 1703 1922 1706 1931
rect 1719 1924 1722 1937
rect 1665 1895 1668 1905
rect 1550 1885 1602 1888
rect 1430 1865 1433 1878
rect 1456 1868 1459 1871
rect 1463 1865 1466 1878
rect 1480 1865 1483 1878
rect 1410 1431 1416 1827
rect 1430 1816 1433 1831
rect 1444 1823 1447 1827
rect 1462 1816 1465 1831
rect 1481 1816 1484 1831
rect 1487 1830 1490 1871
rect 1503 1823 1506 1864
rect 1509 1831 1512 1871
rect 1528 1823 1531 1864
rect 1537 1865 1540 1878
rect 1553 1865 1556 1878
rect 1574 1868 1577 1871
rect 1581 1865 1584 1878
rect 1599 1874 1602 1885
rect 1682 1882 1685 1918
rect 1732 1909 1735 1962
rect 1799 1952 1802 1962
rect 1828 1952 1831 1962
rect 1739 1937 1743 1941
rect 1740 1922 1743 1931
rect 1695 1895 1698 1907
rect 1736 1905 1737 1909
rect 1746 1895 1749 1948
rect 1752 1928 1755 1933
rect 1761 1922 1764 1931
rect 1777 1924 1780 1937
rect 1798 1922 1801 1931
rect 1814 1931 1817 1933
rect 1814 1928 1821 1931
rect 1814 1922 1817 1928
rect 1835 1922 1838 1931
rect 1851 1924 1854 1937
rect 1797 1895 1800 1905
rect 1814 1888 1817 1910
rect 1864 1909 1867 1962
rect 1931 1952 1934 1962
rect 1871 1937 1875 1941
rect 1872 1922 1875 1931
rect 1827 1895 1830 1907
rect 1868 1905 1869 1909
rect 1878 1895 1881 1948
rect 1884 1928 1887 1933
rect 1893 1922 1896 1931
rect 1909 1924 1912 1937
rect 1930 1922 1933 1931
rect 1946 1931 1949 1933
rect 1946 1928 1950 1931
rect 1946 1922 1949 1928
rect 1946 1914 1949 1918
rect 1929 1895 1932 1905
rect 1680 1877 1685 1882
rect 1742 1884 1817 1888
rect 1599 1871 1644 1874
rect 1599 1861 1602 1871
rect 1617 1858 1637 1861
rect 1634 1839 1637 1858
rect 1537 1816 1540 1831
rect 1552 1816 1555 1831
rect 1559 1823 1563 1826
rect 1580 1816 1583 1831
rect 1430 1797 1433 1812
rect 1444 1801 1447 1805
rect 1462 1797 1465 1812
rect 1481 1797 1484 1812
rect 1430 1750 1433 1763
rect 1456 1757 1459 1760
rect 1430 1733 1433 1746
rect 1440 1743 1444 1753
rect 1463 1750 1466 1763
rect 1480 1750 1483 1763
rect 1487 1757 1490 1798
rect 1503 1764 1506 1805
rect 1509 1757 1512 1797
rect 1528 1764 1531 1805
rect 1537 1797 1540 1812
rect 1552 1797 1555 1812
rect 1559 1802 1563 1805
rect 1580 1797 1583 1812
rect 1537 1750 1540 1763
rect 1456 1736 1459 1739
rect 1463 1733 1466 1746
rect 1480 1733 1483 1746
rect 1430 1684 1433 1699
rect 1444 1691 1447 1695
rect 1462 1684 1465 1699
rect 1481 1684 1484 1699
rect 1487 1698 1490 1739
rect 1503 1691 1506 1732
rect 1509 1699 1512 1739
rect 1528 1691 1531 1732
rect 1537 1733 1540 1746
rect 1553 1750 1556 1763
rect 1574 1757 1577 1760
rect 1581 1750 1584 1763
rect 1634 1763 1637 1835
rect 1645 1799 1648 1871
rect 1680 1874 1683 1877
rect 1680 1871 1725 1874
rect 1680 1861 1683 1871
rect 1553 1733 1556 1746
rect 1574 1736 1577 1739
rect 1581 1733 1584 1746
rect 1634 1729 1637 1759
rect 1645 1743 1648 1795
rect 1652 1783 1656 1849
rect 1640 1739 1644 1742
rect 1633 1726 1637 1729
rect 1634 1707 1637 1726
rect 1537 1684 1540 1699
rect 1552 1684 1555 1699
rect 1559 1691 1563 1694
rect 1580 1684 1583 1699
rect 1430 1665 1433 1680
rect 1444 1669 1447 1673
rect 1462 1665 1465 1680
rect 1481 1665 1484 1680
rect 1430 1618 1433 1631
rect 1456 1625 1459 1628
rect 1430 1601 1433 1614
rect 1463 1618 1466 1631
rect 1480 1618 1483 1631
rect 1487 1625 1490 1666
rect 1503 1632 1506 1673
rect 1509 1625 1512 1665
rect 1528 1632 1531 1673
rect 1537 1665 1540 1680
rect 1552 1665 1555 1680
rect 1559 1670 1563 1673
rect 1580 1665 1583 1680
rect 1537 1618 1540 1631
rect 1456 1604 1459 1607
rect 1463 1601 1466 1614
rect 1480 1601 1483 1614
rect 1430 1552 1433 1567
rect 1444 1559 1447 1563
rect 1462 1552 1465 1567
rect 1481 1552 1484 1567
rect 1487 1566 1490 1607
rect 1503 1559 1506 1600
rect 1509 1567 1512 1607
rect 1528 1559 1531 1600
rect 1537 1601 1540 1614
rect 1553 1618 1556 1631
rect 1574 1625 1577 1628
rect 1581 1618 1584 1631
rect 1634 1632 1637 1703
rect 1645 1668 1648 1739
rect 1553 1601 1556 1614
rect 1574 1604 1577 1607
rect 1581 1601 1584 1614
rect 1634 1575 1637 1628
rect 1645 1611 1648 1664
rect 1652 1652 1656 1717
rect 1640 1607 1644 1610
rect 1683 1610 1686 1861
rect 1698 1858 1718 1861
rect 1715 1839 1718 1858
rect 1715 1763 1718 1835
rect 1726 1799 1729 1871
rect 1733 1783 1737 1849
rect 1742 1750 1745 1884
rect 1946 1881 1949 1910
rect 1770 1878 1877 1881
rect 1704 1746 1745 1750
rect 1704 1742 1707 1746
rect 1704 1739 1749 1742
rect 1704 1729 1707 1739
rect 1722 1726 1742 1729
rect 1704 1724 1707 1725
rect 1739 1707 1742 1726
rect 1739 1632 1742 1703
rect 1750 1668 1753 1739
rect 1757 1652 1761 1717
rect 1537 1552 1540 1567
rect 1552 1552 1555 1567
rect 1559 1559 1563 1562
rect 1580 1552 1583 1567
rect 1430 1533 1433 1548
rect 1444 1537 1447 1541
rect 1462 1533 1465 1548
rect 1481 1533 1484 1548
rect 1430 1486 1433 1499
rect 1456 1493 1459 1496
rect 1430 1469 1433 1482
rect 1463 1486 1466 1499
rect 1480 1486 1483 1499
rect 1487 1493 1490 1534
rect 1503 1500 1506 1541
rect 1509 1493 1512 1533
rect 1528 1500 1531 1541
rect 1537 1533 1540 1548
rect 1552 1533 1555 1548
rect 1559 1538 1563 1541
rect 1580 1533 1583 1548
rect 1537 1486 1540 1499
rect 1456 1472 1459 1475
rect 1463 1469 1466 1482
rect 1480 1469 1483 1482
rect 1410 1321 1416 1427
rect 1430 1420 1433 1435
rect 1444 1427 1447 1431
rect 1430 1401 1433 1416
rect 1453 1413 1457 1423
rect 1462 1420 1465 1435
rect 1481 1420 1484 1435
rect 1487 1434 1490 1475
rect 1503 1427 1506 1468
rect 1509 1435 1512 1475
rect 1528 1427 1531 1468
rect 1537 1469 1540 1482
rect 1553 1486 1556 1499
rect 1574 1493 1577 1496
rect 1581 1486 1584 1499
rect 1634 1497 1637 1571
rect 1645 1533 1648 1607
rect 1680 1607 1725 1610
rect 1680 1597 1683 1607
rect 1698 1594 1718 1597
rect 1553 1469 1556 1482
rect 1574 1472 1577 1475
rect 1581 1469 1584 1482
rect 1634 1443 1637 1493
rect 1645 1479 1648 1529
rect 1652 1517 1656 1585
rect 1715 1575 1718 1594
rect 1715 1497 1718 1571
rect 1726 1533 1729 1607
rect 1770 1610 1773 1878
rect 1881 1878 1949 1881
rect 1770 1607 1815 1610
rect 1770 1597 1773 1607
rect 1788 1594 1808 1597
rect 1733 1517 1737 1585
rect 1805 1575 1808 1594
rect 1805 1497 1808 1571
rect 1816 1533 1819 1607
rect 1823 1517 1827 1585
rect 1640 1475 1644 1478
rect 1537 1420 1540 1435
rect 1552 1420 1555 1435
rect 1559 1427 1563 1430
rect 1580 1420 1583 1435
rect 1444 1405 1447 1409
rect 1462 1401 1465 1416
rect 1481 1401 1484 1416
rect 1430 1354 1433 1367
rect 1456 1361 1459 1364
rect 1438 1347 1442 1357
rect 1463 1354 1466 1367
rect 1480 1354 1483 1367
rect 1487 1361 1490 1402
rect 1503 1368 1506 1409
rect 1509 1361 1512 1401
rect 1528 1368 1531 1409
rect 1537 1401 1540 1416
rect 1552 1401 1555 1416
rect 1559 1406 1563 1409
rect 1580 1401 1583 1416
rect 1537 1354 1540 1367
rect 1553 1354 1556 1367
rect 1574 1361 1577 1364
rect 1581 1354 1584 1367
rect 1634 1361 1637 1439
rect 1645 1397 1648 1475
rect 1652 1381 1656 1453
rect 1664 1354 1668 1367
rect 1673 1347 1676 1357
rect 1683 1340 1686 1409
rect 1705 1405 1708 1409
rect 1723 1401 1726 1416
rect 1742 1401 1745 1416
rect 1690 1354 1694 1367
rect 1717 1361 1720 1364
rect 1724 1354 1727 1367
rect 1741 1354 1744 1367
rect 1748 1361 1751 1402
rect 1764 1368 1767 1409
rect 1770 1361 1773 1401
rect 1789 1368 1792 1409
rect 1798 1401 1801 1416
rect 1813 1401 1816 1416
rect 1820 1406 1824 1409
rect 1841 1401 1844 1416
rect 1798 1354 1801 1367
rect 1814 1354 1817 1367
rect 1835 1361 1838 1364
rect 1842 1354 1845 1367
rect 1858 1348 1862 1584
rect 1851 1336 1852 1339
rect 1410 1291 1416 1317
rect 1410 1235 1416 1287
rect 1410 1205 1416 1231
rect 1716 1228 1720 1310
rect 1731 1307 1734 1317
rect 1738 1277 1741 1286
rect 1754 1279 1757 1292
rect 1767 1264 1770 1317
rect 1834 1307 1837 1317
rect 1774 1292 1778 1296
rect 1775 1277 1778 1286
rect 1730 1250 1733 1262
rect 1771 1260 1772 1264
rect 1781 1250 1784 1303
rect 1849 1292 1852 1336
rect 1787 1283 1790 1288
rect 1796 1277 1799 1286
rect 1812 1279 1815 1292
rect 1833 1277 1836 1286
rect 1849 1277 1852 1286
rect 1832 1250 1835 1260
rect 1849 1243 1852 1273
rect 1410 1065 1416 1201
rect 1724 1201 1727 1238
rect 1731 1221 1734 1231
rect 1738 1191 1741 1200
rect 1754 1193 1757 1206
rect 1767 1178 1770 1231
rect 1834 1221 1837 1231
rect 1774 1206 1778 1210
rect 1775 1191 1778 1200
rect 1730 1164 1733 1176
rect 1771 1174 1772 1178
rect 1781 1164 1784 1217
rect 1787 1197 1790 1202
rect 1796 1191 1799 1200
rect 1812 1193 1815 1206
rect 1833 1191 1836 1200
rect 1849 1201 1852 1202
rect 1870 1204 1874 1344
rect 1849 1196 1852 1197
rect 1832 1164 1835 1174
rect 1870 1102 1874 1184
rect 1410 986 1416 1061
rect 1410 953 1416 982
rect 1432 972 1435 982
rect 1410 851 1416 949
rect 1439 942 1442 951
rect 1455 944 1458 957
rect 1468 929 1471 982
rect 1535 972 1538 982
rect 1564 972 1567 982
rect 1475 957 1479 961
rect 1476 942 1479 951
rect 1431 915 1434 927
rect 1472 925 1473 929
rect 1482 915 1485 968
rect 1488 948 1491 953
rect 1497 942 1500 951
rect 1513 944 1516 957
rect 1534 942 1537 951
rect 1550 951 1553 953
rect 1550 948 1557 951
rect 1550 942 1553 948
rect 1571 942 1574 951
rect 1587 944 1590 957
rect 1533 915 1536 925
rect 1550 908 1553 938
rect 1600 929 1603 982
rect 1667 972 1670 982
rect 1696 972 1699 982
rect 1607 957 1611 961
rect 1608 942 1611 951
rect 1563 915 1566 927
rect 1604 925 1605 929
rect 1614 915 1617 968
rect 1620 948 1623 953
rect 1629 942 1632 951
rect 1645 944 1648 957
rect 1666 942 1669 951
rect 1682 951 1685 953
rect 1682 948 1689 951
rect 1682 942 1685 948
rect 1703 942 1706 951
rect 1719 944 1722 957
rect 1665 915 1668 925
rect 1550 905 1602 908
rect 1430 885 1433 898
rect 1456 888 1459 891
rect 1463 885 1466 898
rect 1480 885 1483 898
rect 1410 451 1416 847
rect 1430 836 1433 851
rect 1444 843 1447 847
rect 1462 836 1465 851
rect 1481 836 1484 851
rect 1487 850 1490 891
rect 1503 843 1506 884
rect 1509 851 1512 891
rect 1528 843 1531 884
rect 1537 885 1540 898
rect 1553 885 1556 898
rect 1574 888 1577 891
rect 1581 885 1584 898
rect 1599 894 1602 905
rect 1682 902 1685 938
rect 1732 929 1735 982
rect 1799 972 1802 982
rect 1828 972 1831 982
rect 1739 957 1743 961
rect 1740 942 1743 951
rect 1695 915 1698 927
rect 1736 925 1737 929
rect 1746 915 1749 968
rect 1752 948 1755 953
rect 1761 942 1764 951
rect 1777 944 1780 957
rect 1798 942 1801 951
rect 1814 951 1817 953
rect 1814 948 1821 951
rect 1814 942 1817 948
rect 1835 942 1838 951
rect 1851 944 1854 957
rect 1797 915 1800 925
rect 1814 908 1817 930
rect 1864 929 1867 982
rect 1931 972 1934 982
rect 1871 957 1875 961
rect 1872 942 1875 951
rect 1827 915 1830 927
rect 1868 925 1869 929
rect 1878 915 1881 968
rect 1884 948 1887 953
rect 1893 942 1896 951
rect 1909 944 1912 957
rect 1930 942 1933 951
rect 1946 951 1949 953
rect 1946 948 1950 951
rect 1946 942 1949 948
rect 1946 934 1949 938
rect 1929 915 1932 925
rect 1680 897 1685 902
rect 1742 904 1817 908
rect 1599 891 1644 894
rect 1599 881 1602 891
rect 1617 878 1637 881
rect 1634 859 1637 878
rect 1537 836 1540 851
rect 1552 836 1555 851
rect 1559 843 1563 846
rect 1580 836 1583 851
rect 1430 817 1433 832
rect 1444 821 1447 825
rect 1462 817 1465 832
rect 1481 817 1484 832
rect 1430 770 1433 783
rect 1456 777 1459 780
rect 1430 753 1433 766
rect 1440 763 1444 773
rect 1463 770 1466 783
rect 1480 770 1483 783
rect 1487 777 1490 818
rect 1503 784 1506 825
rect 1509 777 1512 817
rect 1528 784 1531 825
rect 1537 817 1540 832
rect 1552 817 1555 832
rect 1559 822 1563 825
rect 1580 817 1583 832
rect 1537 770 1540 783
rect 1456 756 1459 759
rect 1463 753 1466 766
rect 1480 753 1483 766
rect 1430 704 1433 719
rect 1444 711 1447 715
rect 1462 704 1465 719
rect 1481 704 1484 719
rect 1487 718 1490 759
rect 1503 711 1506 752
rect 1509 719 1512 759
rect 1528 711 1531 752
rect 1537 753 1540 766
rect 1553 770 1556 783
rect 1574 777 1577 780
rect 1581 770 1584 783
rect 1634 783 1637 855
rect 1645 819 1648 891
rect 1680 894 1683 897
rect 1680 891 1725 894
rect 1680 881 1683 891
rect 1553 753 1556 766
rect 1574 756 1577 759
rect 1581 753 1584 766
rect 1634 749 1637 779
rect 1645 763 1648 815
rect 1652 803 1656 869
rect 1640 759 1644 762
rect 1633 746 1637 749
rect 1634 727 1637 746
rect 1537 704 1540 719
rect 1552 704 1555 719
rect 1559 711 1563 714
rect 1580 704 1583 719
rect 1430 685 1433 700
rect 1444 689 1447 693
rect 1462 685 1465 700
rect 1481 685 1484 700
rect 1430 638 1433 651
rect 1456 645 1459 648
rect 1430 621 1433 634
rect 1463 638 1466 651
rect 1480 638 1483 651
rect 1487 645 1490 686
rect 1503 652 1506 693
rect 1509 645 1512 685
rect 1528 652 1531 693
rect 1537 685 1540 700
rect 1552 685 1555 700
rect 1559 690 1563 693
rect 1580 685 1583 700
rect 1537 638 1540 651
rect 1456 624 1459 627
rect 1463 621 1466 634
rect 1480 621 1483 634
rect 1430 572 1433 587
rect 1444 579 1447 583
rect 1462 572 1465 587
rect 1481 572 1484 587
rect 1487 586 1490 627
rect 1503 579 1506 620
rect 1509 587 1512 627
rect 1528 579 1531 620
rect 1537 621 1540 634
rect 1553 638 1556 651
rect 1574 645 1577 648
rect 1581 638 1584 651
rect 1634 652 1637 723
rect 1645 688 1648 759
rect 1553 621 1556 634
rect 1574 624 1577 627
rect 1581 621 1584 634
rect 1634 595 1637 648
rect 1645 631 1648 684
rect 1652 672 1656 737
rect 1640 627 1644 630
rect 1683 630 1686 881
rect 1698 878 1718 881
rect 1715 859 1718 878
rect 1715 783 1718 855
rect 1726 819 1729 891
rect 1733 803 1737 869
rect 1742 770 1745 904
rect 1946 901 1949 930
rect 1770 898 1877 901
rect 1704 766 1745 770
rect 1704 762 1707 766
rect 1704 759 1749 762
rect 1704 749 1707 759
rect 1722 746 1742 749
rect 1704 744 1707 745
rect 1739 727 1742 746
rect 1739 652 1742 723
rect 1750 688 1753 759
rect 1757 672 1761 737
rect 1537 572 1540 587
rect 1552 572 1555 587
rect 1559 579 1563 582
rect 1580 572 1583 587
rect 1430 553 1433 568
rect 1444 557 1447 561
rect 1462 553 1465 568
rect 1481 553 1484 568
rect 1430 506 1433 519
rect 1456 513 1459 516
rect 1430 489 1433 502
rect 1463 506 1466 519
rect 1480 506 1483 519
rect 1487 513 1490 554
rect 1503 520 1506 561
rect 1509 513 1512 553
rect 1528 520 1531 561
rect 1537 553 1540 568
rect 1552 553 1555 568
rect 1559 558 1563 561
rect 1580 553 1583 568
rect 1537 506 1540 519
rect 1456 492 1459 495
rect 1463 489 1466 502
rect 1480 489 1483 502
rect 1410 341 1416 447
rect 1430 440 1433 455
rect 1444 447 1447 451
rect 1430 421 1433 436
rect 1453 433 1457 443
rect 1462 440 1465 455
rect 1481 440 1484 455
rect 1487 454 1490 495
rect 1503 447 1506 488
rect 1509 455 1512 495
rect 1528 447 1531 488
rect 1537 489 1540 502
rect 1553 506 1556 519
rect 1574 513 1577 516
rect 1581 506 1584 519
rect 1634 517 1637 591
rect 1645 553 1648 627
rect 1680 627 1725 630
rect 1680 617 1683 627
rect 1698 614 1718 617
rect 1553 489 1556 502
rect 1574 492 1577 495
rect 1581 489 1584 502
rect 1634 463 1637 513
rect 1645 499 1648 549
rect 1652 537 1656 605
rect 1715 595 1718 614
rect 1715 517 1718 591
rect 1726 553 1729 627
rect 1770 630 1773 898
rect 1881 898 1949 901
rect 1770 627 1815 630
rect 1770 617 1773 627
rect 1788 614 1808 617
rect 1733 537 1737 605
rect 1805 595 1808 614
rect 1805 517 1808 591
rect 1816 553 1819 627
rect 1823 537 1827 605
rect 1640 495 1644 498
rect 1537 440 1540 455
rect 1552 440 1555 455
rect 1559 447 1563 450
rect 1580 440 1583 455
rect 1444 425 1447 429
rect 1462 421 1465 436
rect 1481 421 1484 436
rect 1430 374 1433 387
rect 1456 381 1459 384
rect 1438 367 1442 377
rect 1463 374 1466 387
rect 1480 374 1483 387
rect 1487 381 1490 422
rect 1503 388 1506 429
rect 1509 381 1512 421
rect 1528 388 1531 429
rect 1537 421 1540 436
rect 1552 421 1555 436
rect 1559 426 1563 429
rect 1580 421 1583 436
rect 1537 374 1540 387
rect 1553 374 1556 387
rect 1574 381 1577 384
rect 1581 374 1584 387
rect 1634 381 1637 459
rect 1645 417 1648 495
rect 1652 401 1656 473
rect 1664 374 1668 387
rect 1673 367 1676 377
rect 1683 360 1686 429
rect 1705 425 1708 429
rect 1723 421 1726 436
rect 1742 421 1745 436
rect 1690 374 1694 387
rect 1717 381 1720 384
rect 1724 374 1727 387
rect 1741 374 1744 387
rect 1748 381 1751 422
rect 1764 388 1767 429
rect 1770 381 1773 421
rect 1789 388 1792 429
rect 1798 421 1801 436
rect 1813 421 1816 436
rect 1820 426 1824 429
rect 1841 421 1844 436
rect 1798 374 1801 387
rect 1814 374 1817 387
rect 1835 381 1838 384
rect 1842 374 1845 387
rect 1858 368 1862 604
rect 1851 356 1852 359
rect 1410 311 1416 337
rect 1410 255 1416 307
rect 1410 225 1416 251
rect 1716 248 1720 330
rect 1731 327 1734 337
rect 1738 297 1741 306
rect 1754 299 1757 312
rect 1767 284 1770 337
rect 1834 327 1837 337
rect 1774 312 1778 316
rect 1775 297 1778 306
rect 1730 270 1733 282
rect 1771 280 1772 284
rect 1781 270 1784 323
rect 1849 312 1852 356
rect 1787 303 1790 308
rect 1796 297 1799 306
rect 1812 299 1815 312
rect 1833 297 1836 306
rect 1849 297 1852 306
rect 1832 270 1835 280
rect 1849 263 1852 293
rect 1410 85 1416 221
rect 1724 221 1727 258
rect 1731 241 1734 251
rect 1738 211 1741 220
rect 1754 213 1757 226
rect 1767 198 1770 251
rect 1834 241 1837 251
rect 1774 226 1778 230
rect 1775 211 1778 220
rect 1730 184 1733 196
rect 1771 194 1772 198
rect 1781 184 1784 237
rect 1787 217 1790 222
rect 1796 211 1799 220
rect 1812 213 1815 226
rect 1833 211 1836 220
rect 1849 221 1852 222
rect 1870 224 1874 364
rect 1849 216 1852 217
rect 1832 184 1835 194
rect 1870 122 1874 204
rect 1410 0 1416 81
<< m3contact >>
rect 20 1389 24 1393
rect 277 1892 281 1896
rect 276 1789 280 1793
rect 20 409 24 413
rect 409 1024 413 1028
rect 277 912 281 916
rect 276 809 280 813
rect 409 44 413 48
rect 488 1928 492 1932
rect 528 1845 533 1850
rect 539 1841 544 1846
rect 562 1850 567 1855
rect 586 1845 591 1850
rect 601 1849 606 1855
rect 631 1845 636 1850
rect 660 1844 665 1849
rect 615 1839 620 1844
rect 644 1839 648 1844
rect 686 1838 691 1843
rect 492 1785 497 1790
rect 528 1778 533 1783
rect 539 1782 544 1787
rect 562 1773 567 1778
rect 586 1778 591 1783
rect 615 1784 620 1789
rect 644 1784 648 1789
rect 601 1773 606 1779
rect 631 1778 636 1783
rect 660 1779 665 1784
rect 686 1779 691 1784
rect 491 1716 496 1721
rect 528 1713 533 1718
rect 539 1709 544 1714
rect 562 1718 567 1723
rect 586 1713 591 1718
rect 742 1844 747 1849
rect 601 1717 606 1723
rect 631 1713 636 1718
rect 660 1712 665 1717
rect 615 1707 620 1712
rect 644 1707 648 1712
rect 686 1706 691 1711
rect 492 1653 497 1658
rect 528 1646 533 1651
rect 539 1650 544 1655
rect 562 1641 567 1646
rect 586 1646 591 1651
rect 615 1652 620 1657
rect 644 1652 648 1657
rect 601 1641 606 1647
rect 631 1646 636 1651
rect 660 1647 665 1652
rect 685 1648 690 1653
rect 491 1584 496 1589
rect 528 1581 533 1586
rect 539 1577 544 1582
rect 562 1586 567 1591
rect 586 1581 591 1586
rect 601 1585 606 1591
rect 631 1581 636 1586
rect 660 1580 665 1585
rect 615 1575 620 1580
rect 644 1575 648 1580
rect 686 1574 691 1579
rect 742 1720 747 1725
rect 767 1838 772 1843
rect 766 1779 771 1784
rect 827 1844 832 1849
rect 791 1706 796 1711
rect 791 1648 796 1653
rect 492 1521 497 1526
rect 528 1514 533 1519
rect 539 1518 544 1523
rect 562 1509 567 1514
rect 586 1514 591 1519
rect 615 1520 620 1525
rect 644 1520 648 1525
rect 601 1509 606 1515
rect 631 1514 636 1519
rect 660 1515 665 1520
rect 686 1513 691 1518
rect 491 1452 496 1457
rect 528 1449 533 1454
rect 539 1445 544 1450
rect 562 1454 567 1459
rect 586 1449 591 1454
rect 601 1453 606 1459
rect 631 1449 636 1454
rect 660 1448 665 1453
rect 615 1443 620 1448
rect 644 1443 648 1448
rect 686 1442 691 1447
rect 742 1580 747 1585
rect 767 1574 772 1579
rect 766 1513 771 1518
rect 944 1877 948 1881
rect 849 1717 854 1722
rect 824 1589 829 1594
rect 858 1582 863 1587
rect 855 1509 860 1514
rect 492 1389 497 1394
rect 528 1382 533 1387
rect 539 1386 544 1391
rect 562 1377 567 1382
rect 586 1382 591 1387
rect 615 1388 620 1393
rect 644 1388 648 1393
rect 601 1377 606 1383
rect 631 1382 636 1387
rect 660 1383 665 1388
rect 685 1377 690 1382
rect 742 1456 747 1461
rect 730 1388 735 1393
rect 789 1382 794 1387
rect 800 1386 805 1391
rect 823 1377 828 1382
rect 847 1382 852 1387
rect 876 1388 881 1393
rect 905 1388 909 1393
rect 862 1377 867 1383
rect 892 1382 897 1387
rect 917 1388 922 1393
rect 953 1389 957 1393
rect 791 1279 795 1283
rect 1210 1892 1214 1896
rect 916 1197 920 1201
rect 488 948 492 952
rect 528 865 533 870
rect 539 861 544 866
rect 562 870 567 875
rect 586 865 591 870
rect 601 869 606 875
rect 631 865 636 870
rect 660 864 665 869
rect 615 859 620 864
rect 644 859 648 864
rect 686 858 691 863
rect 492 805 497 810
rect 528 798 533 803
rect 539 802 544 807
rect 562 793 567 798
rect 586 798 591 803
rect 615 804 620 809
rect 644 804 648 809
rect 601 793 606 799
rect 631 798 636 803
rect 660 799 665 804
rect 686 799 691 804
rect 491 736 496 741
rect 528 733 533 738
rect 539 729 544 734
rect 562 738 567 743
rect 586 733 591 738
rect 742 864 747 869
rect 601 737 606 743
rect 631 733 636 738
rect 660 732 665 737
rect 615 727 620 732
rect 644 727 648 732
rect 686 726 691 731
rect 492 673 497 678
rect 528 666 533 671
rect 539 670 544 675
rect 562 661 567 666
rect 586 666 591 671
rect 615 672 620 677
rect 644 672 648 677
rect 601 661 606 667
rect 631 666 636 671
rect 660 667 665 672
rect 685 668 690 673
rect 491 604 496 609
rect 528 601 533 606
rect 539 597 544 602
rect 562 606 567 611
rect 586 601 591 606
rect 601 605 606 611
rect 631 601 636 606
rect 660 600 665 605
rect 615 595 620 600
rect 644 595 648 600
rect 686 594 691 599
rect 742 740 747 745
rect 767 858 772 863
rect 766 799 771 804
rect 827 864 832 869
rect 791 726 796 731
rect 791 668 796 673
rect 492 541 497 546
rect 528 534 533 539
rect 539 538 544 543
rect 562 529 567 534
rect 586 534 591 539
rect 615 540 620 545
rect 644 540 648 545
rect 601 529 606 535
rect 631 534 636 539
rect 660 535 665 540
rect 686 533 691 538
rect 491 472 496 477
rect 528 469 533 474
rect 539 465 544 470
rect 562 474 567 479
rect 586 469 591 474
rect 601 473 606 479
rect 631 469 636 474
rect 660 468 665 473
rect 615 463 620 468
rect 644 463 648 468
rect 686 462 691 467
rect 742 600 747 605
rect 767 594 772 599
rect 766 533 771 538
rect 944 897 948 901
rect 1209 1789 1213 1793
rect 849 737 854 742
rect 824 609 829 614
rect 858 602 863 607
rect 855 529 860 534
rect 492 409 497 414
rect 528 402 533 407
rect 539 406 544 411
rect 562 397 567 402
rect 586 402 591 407
rect 615 408 620 413
rect 644 408 648 413
rect 601 397 606 403
rect 631 402 636 407
rect 660 403 665 408
rect 685 397 690 402
rect 742 476 747 481
rect 730 408 735 413
rect 789 402 794 407
rect 800 406 805 411
rect 823 397 828 402
rect 847 402 852 407
rect 876 408 881 413
rect 905 408 909 413
rect 862 397 867 403
rect 892 402 897 407
rect 917 408 922 413
rect 953 409 957 413
rect 791 299 795 303
rect 1342 1024 1346 1028
rect 1210 913 1214 917
rect 916 217 920 221
rect 1209 809 1213 813
rect 1342 44 1346 48
rect 1421 1928 1425 1932
rect 1461 1845 1466 1850
rect 1472 1841 1477 1846
rect 1495 1850 1500 1855
rect 1519 1845 1524 1850
rect 1534 1849 1539 1855
rect 1564 1845 1569 1850
rect 1593 1844 1598 1849
rect 1548 1839 1553 1844
rect 1577 1839 1581 1844
rect 1619 1838 1624 1843
rect 1425 1785 1430 1790
rect 1461 1778 1466 1783
rect 1472 1782 1477 1787
rect 1495 1773 1500 1778
rect 1519 1778 1524 1783
rect 1548 1784 1553 1789
rect 1577 1784 1581 1789
rect 1534 1773 1539 1779
rect 1564 1778 1569 1783
rect 1593 1779 1598 1784
rect 1619 1779 1624 1784
rect 1424 1716 1429 1721
rect 1461 1713 1466 1718
rect 1472 1709 1477 1714
rect 1495 1718 1500 1723
rect 1519 1713 1524 1718
rect 1675 1844 1680 1849
rect 1534 1717 1539 1723
rect 1564 1713 1569 1718
rect 1593 1712 1598 1717
rect 1548 1707 1553 1712
rect 1577 1707 1581 1712
rect 1619 1706 1624 1711
rect 1425 1653 1430 1658
rect 1461 1646 1466 1651
rect 1472 1650 1477 1655
rect 1495 1641 1500 1646
rect 1519 1646 1524 1651
rect 1548 1652 1553 1657
rect 1577 1652 1581 1657
rect 1534 1641 1539 1647
rect 1564 1646 1569 1651
rect 1593 1647 1598 1652
rect 1618 1648 1623 1653
rect 1424 1584 1429 1589
rect 1461 1581 1466 1586
rect 1472 1577 1477 1582
rect 1495 1586 1500 1591
rect 1519 1581 1524 1586
rect 1534 1585 1539 1591
rect 1564 1581 1569 1586
rect 1593 1580 1598 1585
rect 1548 1575 1553 1580
rect 1577 1575 1581 1580
rect 1619 1574 1624 1579
rect 1675 1720 1680 1725
rect 1700 1838 1705 1843
rect 1699 1779 1704 1784
rect 1760 1844 1765 1849
rect 1724 1706 1729 1711
rect 1724 1648 1729 1653
rect 1425 1521 1430 1526
rect 1461 1514 1466 1519
rect 1472 1518 1477 1523
rect 1495 1509 1500 1514
rect 1519 1514 1524 1519
rect 1548 1520 1553 1525
rect 1577 1520 1581 1525
rect 1534 1509 1539 1515
rect 1564 1514 1569 1519
rect 1593 1515 1598 1520
rect 1619 1513 1624 1518
rect 1424 1452 1429 1457
rect 1461 1449 1466 1454
rect 1472 1445 1477 1450
rect 1495 1454 1500 1459
rect 1519 1449 1524 1454
rect 1534 1453 1539 1459
rect 1564 1449 1569 1454
rect 1593 1448 1598 1453
rect 1548 1443 1553 1448
rect 1577 1443 1581 1448
rect 1619 1442 1624 1447
rect 1675 1580 1680 1585
rect 1700 1574 1705 1579
rect 1699 1513 1704 1518
rect 1877 1877 1881 1881
rect 1782 1717 1787 1722
rect 1757 1589 1762 1594
rect 1791 1582 1796 1587
rect 1788 1509 1793 1514
rect 1425 1389 1430 1394
rect 1461 1382 1466 1387
rect 1472 1386 1477 1391
rect 1495 1377 1500 1382
rect 1519 1382 1524 1387
rect 1548 1388 1553 1393
rect 1577 1388 1581 1393
rect 1534 1377 1539 1383
rect 1564 1382 1569 1387
rect 1593 1383 1598 1388
rect 1618 1377 1623 1382
rect 1675 1456 1680 1461
rect 1663 1388 1668 1393
rect 1722 1382 1727 1387
rect 1733 1386 1738 1391
rect 1756 1377 1761 1382
rect 1780 1382 1785 1387
rect 1809 1388 1814 1393
rect 1838 1388 1842 1393
rect 1795 1377 1800 1383
rect 1825 1382 1830 1387
rect 1850 1388 1855 1393
rect 1724 1279 1728 1283
rect 1849 1197 1853 1201
rect 1421 948 1425 952
rect 1461 865 1466 870
rect 1472 861 1477 866
rect 1495 870 1500 875
rect 1519 865 1524 870
rect 1534 869 1539 875
rect 1564 865 1569 870
rect 1593 864 1598 869
rect 1548 859 1553 864
rect 1577 859 1581 864
rect 1619 858 1624 863
rect 1425 805 1430 810
rect 1461 798 1466 803
rect 1472 802 1477 807
rect 1495 793 1500 798
rect 1519 798 1524 803
rect 1548 804 1553 809
rect 1577 804 1581 809
rect 1534 793 1539 799
rect 1564 798 1569 803
rect 1593 799 1598 804
rect 1619 799 1624 804
rect 1424 736 1429 741
rect 1461 733 1466 738
rect 1472 729 1477 734
rect 1495 738 1500 743
rect 1519 733 1524 738
rect 1675 864 1680 869
rect 1534 737 1539 743
rect 1564 733 1569 738
rect 1593 732 1598 737
rect 1548 727 1553 732
rect 1577 727 1581 732
rect 1619 726 1624 731
rect 1425 673 1430 678
rect 1461 666 1466 671
rect 1472 670 1477 675
rect 1495 661 1500 666
rect 1519 666 1524 671
rect 1548 672 1553 677
rect 1577 672 1581 677
rect 1534 661 1539 667
rect 1564 666 1569 671
rect 1593 667 1598 672
rect 1618 668 1623 673
rect 1424 604 1429 609
rect 1461 601 1466 606
rect 1472 597 1477 602
rect 1495 606 1500 611
rect 1519 601 1524 606
rect 1534 605 1539 611
rect 1564 601 1569 606
rect 1593 600 1598 605
rect 1548 595 1553 600
rect 1577 595 1581 600
rect 1619 594 1624 599
rect 1675 740 1680 745
rect 1700 858 1705 863
rect 1699 799 1704 804
rect 1760 864 1765 869
rect 1724 726 1729 731
rect 1724 668 1729 673
rect 1425 541 1430 546
rect 1461 534 1466 539
rect 1472 538 1477 543
rect 1495 529 1500 534
rect 1519 534 1524 539
rect 1548 540 1553 545
rect 1577 540 1581 545
rect 1534 529 1539 535
rect 1564 534 1569 539
rect 1593 535 1598 540
rect 1619 533 1624 538
rect 1424 472 1429 477
rect 1461 469 1466 474
rect 1472 465 1477 470
rect 1495 474 1500 479
rect 1519 469 1524 474
rect 1534 473 1539 479
rect 1564 469 1569 474
rect 1593 468 1598 473
rect 1548 463 1553 468
rect 1577 463 1581 468
rect 1619 462 1624 467
rect 1675 600 1680 605
rect 1700 594 1705 599
rect 1699 533 1704 538
rect 1877 897 1881 901
rect 1782 737 1787 742
rect 1757 609 1762 614
rect 1791 602 1796 607
rect 1788 529 1793 534
rect 1425 409 1430 414
rect 1461 402 1466 407
rect 1472 406 1477 411
rect 1495 397 1500 402
rect 1519 402 1524 407
rect 1548 408 1553 413
rect 1577 408 1581 413
rect 1534 397 1539 403
rect 1564 402 1569 407
rect 1593 403 1598 408
rect 1618 397 1623 402
rect 1675 476 1680 481
rect 1663 408 1668 413
rect 1722 402 1727 407
rect 1733 406 1738 411
rect 1756 397 1761 402
rect 1780 402 1785 407
rect 1809 408 1814 413
rect 1838 408 1842 413
rect 1795 397 1800 403
rect 1825 402 1830 407
rect 1850 408 1855 413
rect 1724 299 1728 303
rect 1849 217 1853 221
<< metal3 >>
rect 487 1932 493 1933
rect 487 1928 488 1932
rect 492 1928 493 1932
rect 487 1927 493 1928
rect 1420 1932 1426 1933
rect 1420 1928 1421 1932
rect 1425 1928 1426 1932
rect 1420 1927 1426 1928
rect 487 1897 492 1927
rect 1420 1897 1425 1927
rect 276 1896 492 1897
rect 276 1892 277 1896
rect 281 1892 492 1896
rect 1209 1896 1425 1897
rect 1209 1892 1210 1896
rect 1214 1892 1425 1896
rect 276 1891 282 1892
rect 1209 1891 1215 1892
rect 943 1881 949 1882
rect 943 1877 944 1881
rect 948 1877 949 1881
rect 943 1876 949 1877
rect 1876 1881 1882 1882
rect 1876 1877 1877 1881
rect 1881 1877 1882 1881
rect 1876 1876 1882 1877
rect 528 1855 568 1856
rect 528 1851 562 1855
rect 527 1850 534 1851
rect 527 1845 528 1850
rect 533 1845 534 1850
rect 561 1850 562 1851
rect 567 1850 568 1855
rect 600 1855 636 1860
rect 561 1849 568 1850
rect 585 1850 592 1851
rect 527 1844 534 1845
rect 538 1846 545 1847
rect 538 1841 539 1846
rect 544 1841 545 1846
rect 585 1845 586 1850
rect 591 1845 592 1850
rect 600 1849 601 1855
rect 606 1854 636 1855
rect 606 1849 607 1854
rect 631 1851 636 1854
rect 600 1848 607 1849
rect 630 1850 637 1851
rect 630 1845 631 1850
rect 636 1845 637 1850
rect 659 1849 666 1850
rect 585 1844 592 1845
rect 614 1844 621 1845
rect 630 1844 637 1845
rect 643 1844 649 1845
rect 586 1841 591 1844
rect 538 1836 591 1841
rect 614 1839 615 1844
rect 620 1839 621 1844
rect 643 1839 644 1844
rect 648 1839 649 1844
rect 614 1838 649 1839
rect 615 1834 649 1838
rect 659 1844 660 1849
rect 665 1844 666 1849
rect 741 1849 748 1850
rect 741 1844 742 1849
rect 747 1844 748 1849
rect 826 1849 833 1850
rect 826 1844 827 1849
rect 832 1844 833 1849
rect 659 1843 666 1844
rect 685 1843 692 1844
rect 741 1843 748 1844
rect 766 1843 773 1844
rect 826 1843 833 1844
rect 659 1838 686 1843
rect 691 1838 692 1843
rect 742 1838 767 1843
rect 772 1838 773 1843
rect 659 1817 664 1838
rect 685 1837 692 1838
rect 766 1837 773 1838
rect 823 1838 832 1843
rect 492 1811 664 1817
rect 275 1793 281 1794
rect 275 1789 276 1793
rect 280 1789 413 1793
rect 492 1791 497 1811
rect 275 1788 413 1789
rect 19 1393 25 1394
rect 19 1389 20 1393
rect 24 1389 25 1393
rect 19 1388 25 1389
rect 408 1029 413 1788
rect 491 1790 498 1791
rect 491 1785 492 1790
rect 497 1785 498 1790
rect 491 1784 498 1785
rect 538 1787 591 1792
rect 615 1790 649 1794
rect 527 1783 534 1784
rect 527 1778 528 1783
rect 533 1778 534 1783
rect 538 1782 539 1787
rect 544 1782 545 1787
rect 586 1784 591 1787
rect 614 1789 649 1790
rect 614 1784 615 1789
rect 620 1784 621 1789
rect 643 1784 644 1789
rect 648 1784 649 1789
rect 538 1781 545 1782
rect 585 1783 592 1784
rect 614 1783 621 1784
rect 630 1783 637 1784
rect 643 1783 649 1784
rect 659 1784 666 1785
rect 685 1784 692 1785
rect 765 1784 772 1785
rect 527 1777 534 1778
rect 561 1778 568 1779
rect 561 1777 562 1778
rect 528 1773 562 1777
rect 567 1773 568 1778
rect 585 1778 586 1783
rect 591 1778 592 1783
rect 585 1777 592 1778
rect 600 1779 607 1780
rect 528 1772 568 1773
rect 600 1773 601 1779
rect 606 1774 607 1779
rect 630 1778 631 1783
rect 636 1778 637 1783
rect 659 1779 660 1784
rect 665 1779 686 1784
rect 691 1779 692 1784
rect 659 1778 666 1779
rect 685 1778 692 1779
rect 742 1779 766 1784
rect 771 1779 772 1784
rect 630 1777 637 1778
rect 631 1774 636 1777
rect 606 1773 636 1774
rect 600 1768 636 1773
rect 660 1751 665 1778
rect 491 1745 665 1751
rect 491 1722 496 1745
rect 528 1723 568 1724
rect 490 1721 497 1722
rect 490 1716 491 1721
rect 496 1716 497 1721
rect 528 1719 562 1723
rect 490 1715 497 1716
rect 527 1718 534 1719
rect 527 1713 528 1718
rect 533 1713 534 1718
rect 561 1718 562 1719
rect 567 1718 568 1723
rect 600 1723 636 1728
rect 742 1726 747 1779
rect 765 1778 772 1779
rect 823 1750 828 1838
rect 785 1745 828 1750
rect 561 1717 568 1718
rect 585 1718 592 1719
rect 527 1712 534 1713
rect 538 1714 545 1715
rect 538 1709 539 1714
rect 544 1709 545 1714
rect 585 1713 586 1718
rect 591 1713 592 1718
rect 600 1717 601 1723
rect 606 1722 636 1723
rect 606 1717 607 1722
rect 631 1719 636 1722
rect 741 1725 748 1726
rect 741 1720 742 1725
rect 747 1720 748 1725
rect 741 1719 748 1720
rect 600 1716 607 1717
rect 630 1718 637 1719
rect 630 1713 631 1718
rect 636 1713 637 1718
rect 659 1717 666 1718
rect 585 1712 592 1713
rect 614 1712 621 1713
rect 630 1712 637 1713
rect 643 1712 649 1713
rect 586 1709 591 1712
rect 538 1704 591 1709
rect 614 1707 615 1712
rect 620 1707 621 1712
rect 643 1707 644 1712
rect 648 1707 649 1712
rect 614 1706 649 1707
rect 615 1702 649 1706
rect 659 1712 660 1717
rect 665 1712 666 1717
rect 785 1712 790 1745
rect 848 1722 855 1723
rect 848 1717 849 1722
rect 854 1717 855 1722
rect 848 1716 855 1717
rect 659 1711 666 1712
rect 685 1711 692 1712
rect 659 1706 686 1711
rect 691 1706 692 1711
rect 785 1711 797 1712
rect 785 1706 791 1711
rect 796 1706 797 1711
rect 659 1685 664 1706
rect 685 1705 692 1706
rect 790 1705 797 1706
rect 492 1679 664 1685
rect 492 1659 497 1679
rect 491 1658 498 1659
rect 491 1653 492 1658
rect 497 1653 498 1658
rect 491 1652 498 1653
rect 538 1655 591 1660
rect 615 1658 649 1662
rect 527 1651 534 1652
rect 527 1646 528 1651
rect 533 1646 534 1651
rect 538 1650 539 1655
rect 544 1650 545 1655
rect 586 1652 591 1655
rect 614 1657 649 1658
rect 614 1652 615 1657
rect 620 1652 621 1657
rect 643 1652 644 1657
rect 648 1652 649 1657
rect 684 1653 691 1654
rect 790 1653 797 1654
rect 538 1649 545 1650
rect 585 1651 592 1652
rect 614 1651 621 1652
rect 630 1651 637 1652
rect 643 1651 649 1652
rect 659 1652 685 1653
rect 527 1645 534 1646
rect 561 1646 568 1647
rect 561 1645 562 1646
rect 528 1641 562 1645
rect 567 1641 568 1646
rect 585 1646 586 1651
rect 591 1646 592 1651
rect 585 1645 592 1646
rect 600 1647 607 1648
rect 528 1640 568 1641
rect 600 1641 601 1647
rect 606 1642 607 1647
rect 630 1646 631 1651
rect 636 1646 637 1651
rect 630 1645 637 1646
rect 659 1647 660 1652
rect 665 1648 685 1652
rect 690 1648 691 1653
rect 665 1647 666 1648
rect 684 1647 691 1648
rect 786 1648 791 1653
rect 796 1648 797 1653
rect 786 1647 797 1648
rect 659 1646 666 1647
rect 631 1642 636 1645
rect 606 1641 636 1642
rect 600 1636 636 1641
rect 659 1619 664 1646
rect 491 1613 664 1619
rect 786 1619 791 1647
rect 786 1614 829 1619
rect 491 1590 496 1613
rect 528 1591 568 1592
rect 490 1589 497 1590
rect 490 1584 491 1589
rect 496 1584 497 1589
rect 528 1587 562 1591
rect 490 1583 497 1584
rect 527 1586 534 1587
rect 527 1581 528 1586
rect 533 1581 534 1586
rect 561 1586 562 1587
rect 567 1586 568 1591
rect 600 1591 636 1596
rect 824 1595 829 1614
rect 561 1585 568 1586
rect 585 1586 592 1587
rect 527 1580 534 1581
rect 538 1582 545 1583
rect 538 1577 539 1582
rect 544 1577 545 1582
rect 585 1581 586 1586
rect 591 1581 592 1586
rect 600 1585 601 1591
rect 606 1590 636 1591
rect 606 1585 607 1590
rect 631 1587 636 1590
rect 823 1594 830 1595
rect 823 1589 824 1594
rect 829 1589 830 1594
rect 823 1588 830 1589
rect 849 1587 854 1716
rect 857 1587 864 1588
rect 600 1584 607 1585
rect 630 1586 637 1587
rect 630 1581 631 1586
rect 636 1581 637 1586
rect 659 1585 666 1586
rect 585 1580 592 1581
rect 614 1580 621 1581
rect 630 1580 637 1581
rect 643 1580 649 1581
rect 586 1577 591 1580
rect 538 1572 591 1577
rect 614 1575 615 1580
rect 620 1575 621 1580
rect 643 1575 644 1580
rect 648 1575 649 1580
rect 614 1574 649 1575
rect 615 1570 649 1574
rect 659 1580 660 1585
rect 665 1580 666 1585
rect 741 1585 748 1586
rect 741 1580 742 1585
rect 747 1580 748 1585
rect 837 1582 858 1587
rect 863 1582 864 1587
rect 837 1581 849 1582
rect 857 1581 864 1582
rect 659 1579 666 1580
rect 685 1579 692 1580
rect 741 1579 748 1580
rect 766 1579 773 1580
rect 659 1574 686 1579
rect 691 1574 692 1579
rect 742 1574 767 1579
rect 772 1574 773 1579
rect 659 1553 664 1574
rect 685 1573 692 1574
rect 766 1573 773 1574
rect 837 1573 842 1581
rect 492 1547 664 1553
rect 804 1552 842 1573
rect 492 1527 497 1547
rect 491 1526 498 1527
rect 491 1521 492 1526
rect 497 1521 498 1526
rect 491 1520 498 1521
rect 538 1523 591 1528
rect 615 1526 649 1530
rect 527 1519 534 1520
rect 527 1514 528 1519
rect 533 1514 534 1519
rect 538 1518 539 1523
rect 544 1518 545 1523
rect 586 1520 591 1523
rect 614 1525 649 1526
rect 614 1520 615 1525
rect 620 1520 621 1525
rect 643 1520 644 1525
rect 648 1520 649 1525
rect 538 1517 545 1518
rect 585 1519 592 1520
rect 614 1519 621 1520
rect 630 1519 637 1520
rect 643 1519 649 1520
rect 659 1520 666 1521
rect 527 1513 534 1514
rect 561 1514 568 1515
rect 561 1513 562 1514
rect 528 1509 562 1513
rect 567 1509 568 1514
rect 585 1514 586 1519
rect 591 1514 592 1519
rect 585 1513 592 1514
rect 600 1515 607 1516
rect 528 1508 568 1509
rect 600 1509 601 1515
rect 606 1510 607 1515
rect 630 1514 631 1519
rect 636 1514 637 1519
rect 659 1515 660 1520
rect 665 1518 666 1520
rect 685 1518 692 1519
rect 765 1518 772 1519
rect 665 1515 686 1518
rect 659 1514 686 1515
rect 630 1513 637 1514
rect 660 1513 686 1514
rect 691 1513 692 1518
rect 631 1510 636 1513
rect 606 1509 636 1510
rect 600 1504 636 1509
rect 660 1487 665 1513
rect 685 1512 692 1513
rect 742 1513 766 1518
rect 771 1513 772 1518
rect 491 1481 665 1487
rect 491 1458 496 1481
rect 528 1459 568 1460
rect 490 1457 497 1458
rect 490 1452 491 1457
rect 496 1452 497 1457
rect 528 1455 562 1459
rect 490 1451 497 1452
rect 527 1454 534 1455
rect 527 1449 528 1454
rect 533 1449 534 1454
rect 561 1454 562 1455
rect 567 1454 568 1459
rect 600 1459 636 1464
rect 742 1462 747 1513
rect 765 1512 772 1513
rect 561 1453 568 1454
rect 585 1454 592 1455
rect 527 1448 534 1449
rect 538 1450 545 1451
rect 538 1445 539 1450
rect 544 1445 545 1450
rect 585 1449 586 1454
rect 591 1449 592 1454
rect 600 1453 601 1459
rect 606 1458 636 1459
rect 606 1453 607 1458
rect 631 1455 636 1458
rect 741 1461 748 1462
rect 741 1456 742 1461
rect 747 1456 748 1461
rect 741 1455 748 1456
rect 600 1452 607 1453
rect 630 1454 637 1455
rect 630 1449 631 1454
rect 636 1449 637 1454
rect 659 1453 666 1454
rect 585 1448 592 1449
rect 614 1448 621 1449
rect 630 1448 637 1449
rect 643 1448 649 1449
rect 586 1445 591 1448
rect 538 1440 591 1445
rect 614 1443 615 1448
rect 620 1443 621 1448
rect 643 1443 644 1448
rect 648 1443 649 1448
rect 614 1442 649 1443
rect 615 1438 649 1442
rect 659 1448 660 1453
rect 665 1448 666 1453
rect 659 1447 666 1448
rect 685 1447 692 1448
rect 659 1442 686 1447
rect 691 1442 692 1447
rect 804 1443 809 1552
rect 854 1514 861 1515
rect 854 1509 855 1514
rect 860 1509 861 1514
rect 854 1508 861 1509
rect 761 1442 809 1443
rect 659 1421 664 1442
rect 685 1441 692 1442
rect 492 1415 664 1421
rect 730 1437 809 1442
rect 855 1446 860 1508
rect 855 1440 922 1446
rect 492 1395 497 1415
rect 491 1394 498 1395
rect 491 1389 492 1394
rect 497 1389 498 1394
rect 491 1388 498 1389
rect 538 1391 591 1396
rect 615 1394 649 1398
rect 730 1394 735 1437
rect 527 1387 534 1388
rect 527 1382 528 1387
rect 533 1382 534 1387
rect 538 1386 539 1391
rect 544 1386 545 1391
rect 586 1388 591 1391
rect 614 1393 649 1394
rect 614 1388 615 1393
rect 620 1388 621 1393
rect 643 1388 644 1393
rect 648 1388 649 1393
rect 729 1393 736 1394
rect 538 1385 545 1386
rect 585 1387 592 1388
rect 614 1387 621 1388
rect 630 1387 637 1388
rect 643 1387 649 1388
rect 659 1388 666 1389
rect 527 1381 534 1382
rect 561 1382 568 1383
rect 561 1381 562 1382
rect 528 1377 562 1381
rect 567 1377 568 1382
rect 585 1382 586 1387
rect 591 1382 592 1387
rect 585 1381 592 1382
rect 600 1383 607 1384
rect 528 1376 568 1377
rect 600 1377 601 1383
rect 606 1378 607 1383
rect 630 1382 631 1387
rect 636 1382 637 1387
rect 659 1383 660 1388
rect 665 1383 666 1388
rect 729 1388 730 1393
rect 735 1388 736 1393
rect 799 1391 852 1396
rect 876 1394 910 1398
rect 917 1394 922 1440
rect 729 1387 736 1388
rect 788 1387 795 1388
rect 659 1382 666 1383
rect 684 1382 691 1383
rect 630 1381 637 1382
rect 631 1378 636 1381
rect 606 1377 636 1378
rect 600 1372 636 1377
rect 661 1377 685 1382
rect 690 1377 691 1382
rect 788 1382 789 1387
rect 794 1382 795 1387
rect 799 1386 800 1391
rect 805 1386 806 1391
rect 847 1388 852 1391
rect 875 1393 910 1394
rect 875 1388 876 1393
rect 881 1388 882 1393
rect 904 1388 905 1393
rect 909 1388 910 1393
rect 799 1385 806 1386
rect 846 1387 853 1388
rect 875 1387 882 1388
rect 891 1387 898 1388
rect 904 1387 910 1388
rect 916 1393 923 1394
rect 916 1388 917 1393
rect 922 1388 923 1393
rect 916 1387 923 1388
rect 788 1381 795 1382
rect 822 1382 829 1383
rect 822 1381 823 1382
rect 408 1028 414 1029
rect 408 1024 409 1028
rect 413 1024 414 1028
rect 408 1023 414 1024
rect 661 1011 666 1377
rect 684 1376 691 1377
rect 789 1377 823 1381
rect 828 1377 829 1382
rect 846 1382 847 1387
rect 852 1382 853 1387
rect 846 1381 853 1382
rect 861 1383 868 1384
rect 789 1376 829 1377
rect 861 1377 862 1383
rect 867 1378 868 1383
rect 891 1382 892 1387
rect 897 1382 898 1387
rect 891 1381 898 1382
rect 892 1378 897 1381
rect 867 1377 897 1378
rect 861 1372 897 1377
rect 944 1349 949 1876
rect 1461 1855 1501 1856
rect 1421 1853 1428 1854
rect 1411 1848 1428 1853
rect 1461 1851 1495 1855
rect 1208 1793 1214 1794
rect 1208 1789 1209 1793
rect 1213 1789 1346 1793
rect 1208 1788 1346 1789
rect 952 1393 958 1394
rect 952 1389 953 1393
rect 957 1389 958 1393
rect 952 1388 958 1389
rect 791 1344 949 1349
rect 791 1284 796 1344
rect 790 1283 796 1284
rect 790 1279 791 1283
rect 795 1279 796 1283
rect 790 1278 796 1279
rect 953 1221 958 1388
rect 916 1216 958 1221
rect 916 1202 921 1216
rect 915 1201 921 1202
rect 915 1197 916 1201
rect 920 1197 921 1201
rect 915 1196 921 1197
rect 1341 1029 1346 1788
rect 1341 1028 1347 1029
rect 1341 1024 1342 1028
rect 1346 1024 1347 1028
rect 1341 1023 1347 1024
rect 1411 1011 1416 1848
rect 1421 1847 1428 1848
rect 1460 1850 1467 1851
rect 1460 1845 1461 1850
rect 1466 1845 1467 1850
rect 1494 1850 1495 1851
rect 1500 1850 1501 1855
rect 1533 1855 1569 1860
rect 1494 1849 1501 1850
rect 1518 1850 1525 1851
rect 1460 1844 1467 1845
rect 1471 1846 1478 1847
rect 1471 1841 1472 1846
rect 1477 1841 1478 1846
rect 1518 1845 1519 1850
rect 1524 1845 1525 1850
rect 1533 1849 1534 1855
rect 1539 1854 1569 1855
rect 1539 1849 1540 1854
rect 1564 1851 1569 1854
rect 1533 1848 1540 1849
rect 1563 1850 1570 1851
rect 1563 1845 1564 1850
rect 1569 1845 1570 1850
rect 1592 1849 1599 1850
rect 1518 1844 1525 1845
rect 1547 1844 1554 1845
rect 1563 1844 1570 1845
rect 1576 1844 1582 1845
rect 1519 1841 1524 1844
rect 1471 1836 1524 1841
rect 1547 1839 1548 1844
rect 1553 1839 1554 1844
rect 1576 1839 1577 1844
rect 1581 1839 1582 1844
rect 1547 1838 1582 1839
rect 1548 1834 1582 1838
rect 1592 1844 1593 1849
rect 1598 1844 1599 1849
rect 1674 1849 1681 1850
rect 1674 1844 1675 1849
rect 1680 1844 1681 1849
rect 1759 1849 1766 1850
rect 1759 1844 1760 1849
rect 1765 1844 1766 1849
rect 1592 1843 1599 1844
rect 1618 1843 1625 1844
rect 1674 1843 1681 1844
rect 1699 1843 1706 1844
rect 1759 1843 1766 1844
rect 1592 1838 1619 1843
rect 1624 1838 1625 1843
rect 1675 1838 1700 1843
rect 1705 1838 1706 1843
rect 1592 1817 1597 1838
rect 1618 1837 1625 1838
rect 1699 1837 1706 1838
rect 1756 1838 1765 1843
rect 1425 1811 1597 1817
rect 1425 1791 1430 1811
rect 1424 1790 1431 1791
rect 1424 1785 1425 1790
rect 1430 1785 1431 1790
rect 1424 1784 1431 1785
rect 1471 1787 1524 1792
rect 1548 1790 1582 1794
rect 1460 1783 1467 1784
rect 1460 1778 1461 1783
rect 1466 1778 1467 1783
rect 1471 1782 1472 1787
rect 1477 1782 1478 1787
rect 1519 1784 1524 1787
rect 1547 1789 1582 1790
rect 1547 1784 1548 1789
rect 1553 1784 1554 1789
rect 1576 1784 1577 1789
rect 1581 1784 1582 1789
rect 1471 1781 1478 1782
rect 1518 1783 1525 1784
rect 1547 1783 1554 1784
rect 1563 1783 1570 1784
rect 1576 1783 1582 1784
rect 1592 1784 1599 1785
rect 1618 1784 1625 1785
rect 1698 1784 1705 1785
rect 1460 1777 1467 1778
rect 1494 1778 1501 1779
rect 1494 1777 1495 1778
rect 1461 1773 1495 1777
rect 1500 1773 1501 1778
rect 1518 1778 1519 1783
rect 1524 1778 1525 1783
rect 1518 1777 1525 1778
rect 1533 1779 1540 1780
rect 1461 1772 1501 1773
rect 1533 1773 1534 1779
rect 1539 1774 1540 1779
rect 1563 1778 1564 1783
rect 1569 1778 1570 1783
rect 1592 1779 1593 1784
rect 1598 1779 1619 1784
rect 1624 1779 1625 1784
rect 1592 1778 1599 1779
rect 1618 1778 1625 1779
rect 1675 1779 1699 1784
rect 1704 1779 1705 1784
rect 1563 1777 1570 1778
rect 1564 1774 1569 1777
rect 1539 1773 1569 1774
rect 1533 1768 1569 1773
rect 1593 1751 1598 1778
rect 1424 1745 1598 1751
rect 1424 1722 1429 1745
rect 1461 1723 1501 1724
rect 1423 1721 1430 1722
rect 1423 1716 1424 1721
rect 1429 1716 1430 1721
rect 1461 1719 1495 1723
rect 1423 1715 1430 1716
rect 1460 1718 1467 1719
rect 1460 1713 1461 1718
rect 1466 1713 1467 1718
rect 1494 1718 1495 1719
rect 1500 1718 1501 1723
rect 1533 1723 1569 1728
rect 1675 1726 1680 1779
rect 1698 1778 1705 1779
rect 1756 1750 1761 1838
rect 1718 1745 1761 1750
rect 1494 1717 1501 1718
rect 1518 1718 1525 1719
rect 1460 1712 1467 1713
rect 1471 1714 1478 1715
rect 1471 1709 1472 1714
rect 1477 1709 1478 1714
rect 1518 1713 1519 1718
rect 1524 1713 1525 1718
rect 1533 1717 1534 1723
rect 1539 1722 1569 1723
rect 1539 1717 1540 1722
rect 1564 1719 1569 1722
rect 1674 1725 1681 1726
rect 1674 1720 1675 1725
rect 1680 1720 1681 1725
rect 1674 1719 1681 1720
rect 1533 1716 1540 1717
rect 1563 1718 1570 1719
rect 1563 1713 1564 1718
rect 1569 1713 1570 1718
rect 1592 1717 1599 1718
rect 1518 1712 1525 1713
rect 1547 1712 1554 1713
rect 1563 1712 1570 1713
rect 1576 1712 1582 1713
rect 1519 1709 1524 1712
rect 1471 1704 1524 1709
rect 1547 1707 1548 1712
rect 1553 1707 1554 1712
rect 1576 1707 1577 1712
rect 1581 1707 1582 1712
rect 1547 1706 1582 1707
rect 1548 1702 1582 1706
rect 1592 1712 1593 1717
rect 1598 1712 1599 1717
rect 1718 1712 1723 1745
rect 1781 1722 1788 1723
rect 1781 1717 1782 1722
rect 1787 1717 1788 1722
rect 1781 1716 1788 1717
rect 1592 1711 1599 1712
rect 1618 1711 1625 1712
rect 1592 1706 1619 1711
rect 1624 1706 1625 1711
rect 1718 1711 1730 1712
rect 1718 1706 1724 1711
rect 1729 1706 1730 1711
rect 1592 1685 1597 1706
rect 1618 1705 1625 1706
rect 1723 1705 1730 1706
rect 1425 1679 1597 1685
rect 1425 1659 1430 1679
rect 1424 1658 1431 1659
rect 1424 1653 1425 1658
rect 1430 1653 1431 1658
rect 1424 1652 1431 1653
rect 1471 1655 1524 1660
rect 1548 1658 1582 1662
rect 1460 1651 1467 1652
rect 1460 1646 1461 1651
rect 1466 1646 1467 1651
rect 1471 1650 1472 1655
rect 1477 1650 1478 1655
rect 1519 1652 1524 1655
rect 1547 1657 1582 1658
rect 1547 1652 1548 1657
rect 1553 1652 1554 1657
rect 1576 1652 1577 1657
rect 1581 1652 1582 1657
rect 1617 1653 1624 1654
rect 1723 1653 1730 1654
rect 1471 1649 1478 1650
rect 1518 1651 1525 1652
rect 1547 1651 1554 1652
rect 1563 1651 1570 1652
rect 1576 1651 1582 1652
rect 1592 1652 1618 1653
rect 1460 1645 1467 1646
rect 1494 1646 1501 1647
rect 1494 1645 1495 1646
rect 1461 1641 1495 1645
rect 1500 1641 1501 1646
rect 1518 1646 1519 1651
rect 1524 1646 1525 1651
rect 1518 1645 1525 1646
rect 1533 1647 1540 1648
rect 1461 1640 1501 1641
rect 1533 1641 1534 1647
rect 1539 1642 1540 1647
rect 1563 1646 1564 1651
rect 1569 1646 1570 1651
rect 1563 1645 1570 1646
rect 1592 1647 1593 1652
rect 1598 1648 1618 1652
rect 1623 1648 1624 1653
rect 1598 1647 1599 1648
rect 1617 1647 1624 1648
rect 1719 1648 1724 1653
rect 1729 1648 1730 1653
rect 1719 1647 1730 1648
rect 1592 1646 1599 1647
rect 1564 1642 1569 1645
rect 1539 1641 1569 1642
rect 1533 1636 1569 1641
rect 1592 1619 1597 1646
rect 1424 1613 1597 1619
rect 1719 1619 1724 1647
rect 1719 1614 1762 1619
rect 1424 1590 1429 1613
rect 1461 1591 1501 1592
rect 1423 1589 1430 1590
rect 1423 1584 1424 1589
rect 1429 1584 1430 1589
rect 1461 1587 1495 1591
rect 1423 1583 1430 1584
rect 1460 1586 1467 1587
rect 1460 1581 1461 1586
rect 1466 1581 1467 1586
rect 1494 1586 1495 1587
rect 1500 1586 1501 1591
rect 1533 1591 1569 1596
rect 1757 1595 1762 1614
rect 1494 1585 1501 1586
rect 1518 1586 1525 1587
rect 1460 1580 1467 1581
rect 1471 1582 1478 1583
rect 1471 1577 1472 1582
rect 1477 1577 1478 1582
rect 1518 1581 1519 1586
rect 1524 1581 1525 1586
rect 1533 1585 1534 1591
rect 1539 1590 1569 1591
rect 1539 1585 1540 1590
rect 1564 1587 1569 1590
rect 1756 1594 1763 1595
rect 1756 1589 1757 1594
rect 1762 1589 1763 1594
rect 1756 1588 1763 1589
rect 1782 1587 1787 1716
rect 1790 1587 1797 1588
rect 1533 1584 1540 1585
rect 1563 1586 1570 1587
rect 1563 1581 1564 1586
rect 1569 1581 1570 1586
rect 1592 1585 1599 1586
rect 1518 1580 1525 1581
rect 1547 1580 1554 1581
rect 1563 1580 1570 1581
rect 1576 1580 1582 1581
rect 1519 1577 1524 1580
rect 1471 1572 1524 1577
rect 1547 1575 1548 1580
rect 1553 1575 1554 1580
rect 1576 1575 1577 1580
rect 1581 1575 1582 1580
rect 1547 1574 1582 1575
rect 1548 1570 1582 1574
rect 1592 1580 1593 1585
rect 1598 1580 1599 1585
rect 1674 1585 1681 1586
rect 1674 1580 1675 1585
rect 1680 1580 1681 1585
rect 1770 1582 1791 1587
rect 1796 1582 1797 1587
rect 1770 1581 1782 1582
rect 1790 1581 1797 1582
rect 1592 1579 1599 1580
rect 1618 1579 1625 1580
rect 1674 1579 1681 1580
rect 1699 1579 1706 1580
rect 1592 1574 1619 1579
rect 1624 1574 1625 1579
rect 1675 1574 1700 1579
rect 1705 1574 1706 1579
rect 1592 1553 1597 1574
rect 1618 1573 1625 1574
rect 1699 1573 1706 1574
rect 1770 1573 1775 1581
rect 1425 1547 1597 1553
rect 1737 1552 1775 1573
rect 1425 1527 1430 1547
rect 1424 1526 1431 1527
rect 1424 1521 1425 1526
rect 1430 1521 1431 1526
rect 1424 1520 1431 1521
rect 1471 1523 1524 1528
rect 1548 1526 1582 1530
rect 1460 1519 1467 1520
rect 1460 1514 1461 1519
rect 1466 1514 1467 1519
rect 1471 1518 1472 1523
rect 1477 1518 1478 1523
rect 1519 1520 1524 1523
rect 1547 1525 1582 1526
rect 1547 1520 1548 1525
rect 1553 1520 1554 1525
rect 1576 1520 1577 1525
rect 1581 1520 1582 1525
rect 1471 1517 1478 1518
rect 1518 1519 1525 1520
rect 1547 1519 1554 1520
rect 1563 1519 1570 1520
rect 1576 1519 1582 1520
rect 1592 1520 1599 1521
rect 1460 1513 1467 1514
rect 1494 1514 1501 1515
rect 1494 1513 1495 1514
rect 1461 1509 1495 1513
rect 1500 1509 1501 1514
rect 1518 1514 1519 1519
rect 1524 1514 1525 1519
rect 1518 1513 1525 1514
rect 1533 1515 1540 1516
rect 1461 1508 1501 1509
rect 1533 1509 1534 1515
rect 1539 1510 1540 1515
rect 1563 1514 1564 1519
rect 1569 1514 1570 1519
rect 1592 1515 1593 1520
rect 1598 1518 1599 1520
rect 1618 1518 1625 1519
rect 1698 1518 1705 1519
rect 1598 1515 1619 1518
rect 1592 1514 1619 1515
rect 1563 1513 1570 1514
rect 1593 1513 1619 1514
rect 1624 1513 1625 1518
rect 1564 1510 1569 1513
rect 1539 1509 1569 1510
rect 1533 1504 1569 1509
rect 1593 1487 1598 1513
rect 1618 1512 1625 1513
rect 1675 1513 1699 1518
rect 1704 1513 1705 1518
rect 1424 1481 1598 1487
rect 1424 1458 1429 1481
rect 1461 1459 1501 1460
rect 1423 1457 1430 1458
rect 1423 1452 1424 1457
rect 1429 1452 1430 1457
rect 1461 1455 1495 1459
rect 1423 1451 1430 1452
rect 1460 1454 1467 1455
rect 1460 1449 1461 1454
rect 1466 1449 1467 1454
rect 1494 1454 1495 1455
rect 1500 1454 1501 1459
rect 1533 1459 1569 1464
rect 1675 1462 1680 1513
rect 1698 1512 1705 1513
rect 1494 1453 1501 1454
rect 1518 1454 1525 1455
rect 1460 1448 1467 1449
rect 1471 1450 1478 1451
rect 1471 1445 1472 1450
rect 1477 1445 1478 1450
rect 1518 1449 1519 1454
rect 1524 1449 1525 1454
rect 1533 1453 1534 1459
rect 1539 1458 1569 1459
rect 1539 1453 1540 1458
rect 1564 1455 1569 1458
rect 1674 1461 1681 1462
rect 1674 1456 1675 1461
rect 1680 1456 1681 1461
rect 1674 1455 1681 1456
rect 1533 1452 1540 1453
rect 1563 1454 1570 1455
rect 1563 1449 1564 1454
rect 1569 1449 1570 1454
rect 1592 1453 1599 1454
rect 1518 1448 1525 1449
rect 1547 1448 1554 1449
rect 1563 1448 1570 1449
rect 1576 1448 1582 1449
rect 1519 1445 1524 1448
rect 1471 1440 1524 1445
rect 1547 1443 1548 1448
rect 1553 1443 1554 1448
rect 1576 1443 1577 1448
rect 1581 1443 1582 1448
rect 1547 1442 1582 1443
rect 1548 1438 1582 1442
rect 1592 1448 1593 1453
rect 1598 1448 1599 1453
rect 1592 1447 1599 1448
rect 1618 1447 1625 1448
rect 1592 1442 1619 1447
rect 1624 1442 1625 1447
rect 1737 1443 1742 1552
rect 1787 1514 1794 1515
rect 1787 1509 1788 1514
rect 1793 1509 1794 1514
rect 1787 1508 1794 1509
rect 1694 1442 1742 1443
rect 1592 1421 1597 1442
rect 1618 1441 1625 1442
rect 1425 1415 1597 1421
rect 1663 1437 1742 1442
rect 1788 1446 1793 1508
rect 1788 1440 1855 1446
rect 1425 1395 1430 1415
rect 1424 1394 1431 1395
rect 1424 1389 1425 1394
rect 1430 1389 1431 1394
rect 1424 1388 1431 1389
rect 1471 1391 1524 1396
rect 1548 1394 1582 1398
rect 1663 1394 1668 1437
rect 1460 1387 1467 1388
rect 1460 1382 1461 1387
rect 1466 1382 1467 1387
rect 1471 1386 1472 1391
rect 1477 1386 1478 1391
rect 1519 1388 1524 1391
rect 1547 1393 1582 1394
rect 1547 1388 1548 1393
rect 1553 1388 1554 1393
rect 1576 1388 1577 1393
rect 1581 1388 1582 1393
rect 1662 1393 1669 1394
rect 1471 1385 1478 1386
rect 1518 1387 1525 1388
rect 1547 1387 1554 1388
rect 1563 1387 1570 1388
rect 1576 1387 1582 1388
rect 1592 1388 1599 1389
rect 1460 1381 1467 1382
rect 1494 1382 1501 1383
rect 1494 1381 1495 1382
rect 1461 1377 1495 1381
rect 1500 1377 1501 1382
rect 1518 1382 1519 1387
rect 1524 1382 1525 1387
rect 1518 1381 1525 1382
rect 1533 1383 1540 1384
rect 1461 1376 1501 1377
rect 1533 1377 1534 1383
rect 1539 1378 1540 1383
rect 1563 1382 1564 1387
rect 1569 1382 1570 1387
rect 1592 1383 1593 1388
rect 1598 1383 1599 1388
rect 1662 1388 1663 1393
rect 1668 1388 1669 1393
rect 1732 1391 1785 1396
rect 1809 1394 1843 1398
rect 1850 1394 1855 1440
rect 1662 1387 1669 1388
rect 1721 1387 1728 1388
rect 1592 1382 1599 1383
rect 1617 1382 1624 1383
rect 1563 1381 1570 1382
rect 1564 1378 1569 1381
rect 1539 1377 1569 1378
rect 1533 1372 1569 1377
rect 1594 1377 1618 1382
rect 1623 1377 1624 1382
rect 1721 1382 1722 1387
rect 1727 1382 1728 1387
rect 1732 1386 1733 1391
rect 1738 1386 1739 1391
rect 1780 1388 1785 1391
rect 1808 1393 1843 1394
rect 1808 1388 1809 1393
rect 1814 1388 1815 1393
rect 1837 1388 1838 1393
rect 1842 1388 1843 1393
rect 1732 1385 1739 1386
rect 1779 1387 1786 1388
rect 1808 1387 1815 1388
rect 1824 1387 1831 1388
rect 1837 1387 1843 1388
rect 1849 1393 1856 1394
rect 1849 1388 1850 1393
rect 1855 1388 1856 1393
rect 1849 1387 1856 1388
rect 1721 1381 1728 1382
rect 1755 1382 1762 1383
rect 1755 1381 1756 1382
rect 1594 1248 1599 1377
rect 1617 1376 1624 1377
rect 1722 1377 1756 1381
rect 1761 1377 1762 1382
rect 1779 1382 1780 1387
rect 1785 1382 1786 1387
rect 1779 1381 1786 1382
rect 1794 1383 1801 1384
rect 1722 1376 1762 1377
rect 1794 1377 1795 1383
rect 1800 1378 1801 1383
rect 1824 1382 1825 1387
rect 1830 1382 1831 1387
rect 1824 1381 1831 1382
rect 1825 1378 1830 1381
rect 1800 1377 1830 1378
rect 1794 1372 1830 1377
rect 1877 1349 1882 1876
rect 1724 1344 1882 1349
rect 1724 1284 1729 1344
rect 1723 1283 1729 1284
rect 1723 1279 1724 1283
rect 1728 1279 1729 1283
rect 1723 1278 1729 1279
rect 1594 1242 1905 1248
rect 1848 1201 1854 1202
rect 1848 1197 1849 1201
rect 1853 1197 1854 1201
rect 1848 1196 1854 1197
rect 661 1005 1416 1011
rect 1849 992 1854 1196
rect 20 987 1854 992
rect 20 414 25 987
rect 414 952 493 953
rect 414 948 488 952
rect 492 948 493 952
rect 415 917 420 948
rect 487 947 493 948
rect 1420 952 1426 953
rect 1420 948 1421 952
rect 1425 948 1426 952
rect 1420 947 1426 948
rect 276 916 420 917
rect 276 912 277 916
rect 281 912 420 916
rect 1209 917 1215 918
rect 1420 917 1425 947
rect 276 911 282 912
rect 490 909 970 914
rect 1209 913 1210 917
rect 1214 913 1425 917
rect 1900 914 1905 1242
rect 1209 912 1425 913
rect 1563 909 1905 914
rect 490 874 495 909
rect 965 904 1591 909
rect 943 901 949 902
rect 943 897 944 901
rect 948 897 949 901
rect 943 896 949 897
rect 1876 901 1882 902
rect 1876 897 1877 901
rect 1881 897 1882 901
rect 1876 896 1882 897
rect 528 875 568 876
rect 489 867 496 874
rect 528 871 562 875
rect 527 870 534 871
rect 527 865 528 870
rect 533 865 534 870
rect 561 870 562 871
rect 567 870 568 875
rect 600 875 636 880
rect 561 869 568 870
rect 585 870 592 871
rect 527 864 534 865
rect 538 866 545 867
rect 538 861 539 866
rect 544 861 545 866
rect 585 865 586 870
rect 591 865 592 870
rect 600 869 601 875
rect 606 874 636 875
rect 606 869 607 874
rect 631 871 636 874
rect 600 868 607 869
rect 630 870 637 871
rect 630 865 631 870
rect 636 865 637 870
rect 659 869 666 870
rect 585 864 592 865
rect 614 864 621 865
rect 630 864 637 865
rect 643 864 649 865
rect 586 861 591 864
rect 538 856 591 861
rect 614 859 615 864
rect 620 859 621 864
rect 643 859 644 864
rect 648 859 649 864
rect 614 858 649 859
rect 615 854 649 858
rect 659 864 660 869
rect 665 864 666 869
rect 741 869 748 870
rect 741 864 742 869
rect 747 864 748 869
rect 826 869 833 870
rect 826 864 827 869
rect 832 864 833 869
rect 659 863 666 864
rect 685 863 692 864
rect 741 863 748 864
rect 766 863 773 864
rect 826 863 833 864
rect 659 858 686 863
rect 691 858 692 863
rect 742 858 767 863
rect 772 858 773 863
rect 659 837 664 858
rect 685 857 692 858
rect 766 857 773 858
rect 823 858 832 863
rect 492 831 664 837
rect 275 813 281 814
rect 275 809 276 813
rect 280 809 413 813
rect 492 811 497 831
rect 275 808 413 809
rect 19 413 25 414
rect 19 409 20 413
rect 24 409 25 413
rect 19 408 25 409
rect 408 49 413 808
rect 491 810 498 811
rect 491 805 492 810
rect 497 805 498 810
rect 491 804 498 805
rect 538 807 591 812
rect 615 810 649 814
rect 527 803 534 804
rect 527 798 528 803
rect 533 798 534 803
rect 538 802 539 807
rect 544 802 545 807
rect 586 804 591 807
rect 614 809 649 810
rect 614 804 615 809
rect 620 804 621 809
rect 643 804 644 809
rect 648 804 649 809
rect 538 801 545 802
rect 585 803 592 804
rect 614 803 621 804
rect 630 803 637 804
rect 643 803 649 804
rect 659 804 666 805
rect 685 804 692 805
rect 765 804 772 805
rect 527 797 534 798
rect 561 798 568 799
rect 561 797 562 798
rect 528 793 562 797
rect 567 793 568 798
rect 585 798 586 803
rect 591 798 592 803
rect 585 797 592 798
rect 600 799 607 800
rect 528 792 568 793
rect 600 793 601 799
rect 606 794 607 799
rect 630 798 631 803
rect 636 798 637 803
rect 659 799 660 804
rect 665 799 686 804
rect 691 799 692 804
rect 659 798 666 799
rect 685 798 692 799
rect 742 799 766 804
rect 771 799 772 804
rect 630 797 637 798
rect 631 794 636 797
rect 606 793 636 794
rect 600 788 636 793
rect 660 771 665 798
rect 491 765 665 771
rect 491 742 496 765
rect 528 743 568 744
rect 490 741 497 742
rect 490 736 491 741
rect 496 736 497 741
rect 528 739 562 743
rect 490 735 497 736
rect 527 738 534 739
rect 527 733 528 738
rect 533 733 534 738
rect 561 738 562 739
rect 567 738 568 743
rect 600 743 636 748
rect 742 746 747 799
rect 765 798 772 799
rect 823 770 828 858
rect 785 765 828 770
rect 561 737 568 738
rect 585 738 592 739
rect 527 732 534 733
rect 538 734 545 735
rect 538 729 539 734
rect 544 729 545 734
rect 585 733 586 738
rect 591 733 592 738
rect 600 737 601 743
rect 606 742 636 743
rect 606 737 607 742
rect 631 739 636 742
rect 741 745 748 746
rect 741 740 742 745
rect 747 740 748 745
rect 741 739 748 740
rect 600 736 607 737
rect 630 738 637 739
rect 630 733 631 738
rect 636 733 637 738
rect 659 737 666 738
rect 585 732 592 733
rect 614 732 621 733
rect 630 732 637 733
rect 643 732 649 733
rect 586 729 591 732
rect 538 724 591 729
rect 614 727 615 732
rect 620 727 621 732
rect 643 727 644 732
rect 648 727 649 732
rect 614 726 649 727
rect 615 722 649 726
rect 659 732 660 737
rect 665 732 666 737
rect 785 732 790 765
rect 848 742 855 743
rect 848 737 849 742
rect 854 737 855 742
rect 848 736 855 737
rect 659 731 666 732
rect 685 731 692 732
rect 659 726 686 731
rect 691 726 692 731
rect 785 731 797 732
rect 785 726 791 731
rect 796 726 797 731
rect 659 705 664 726
rect 685 725 692 726
rect 790 725 797 726
rect 492 699 664 705
rect 492 679 497 699
rect 491 678 498 679
rect 491 673 492 678
rect 497 673 498 678
rect 491 672 498 673
rect 538 675 591 680
rect 615 678 649 682
rect 527 671 534 672
rect 527 666 528 671
rect 533 666 534 671
rect 538 670 539 675
rect 544 670 545 675
rect 586 672 591 675
rect 614 677 649 678
rect 614 672 615 677
rect 620 672 621 677
rect 643 672 644 677
rect 648 672 649 677
rect 684 673 691 674
rect 790 673 797 674
rect 538 669 545 670
rect 585 671 592 672
rect 614 671 621 672
rect 630 671 637 672
rect 643 671 649 672
rect 659 672 685 673
rect 527 665 534 666
rect 561 666 568 667
rect 561 665 562 666
rect 528 661 562 665
rect 567 661 568 666
rect 585 666 586 671
rect 591 666 592 671
rect 585 665 592 666
rect 600 667 607 668
rect 528 660 568 661
rect 600 661 601 667
rect 606 662 607 667
rect 630 666 631 671
rect 636 666 637 671
rect 630 665 637 666
rect 659 667 660 672
rect 665 668 685 672
rect 690 668 691 673
rect 665 667 666 668
rect 684 667 691 668
rect 786 668 791 673
rect 796 668 797 673
rect 786 667 797 668
rect 659 666 666 667
rect 631 662 636 665
rect 606 661 636 662
rect 600 656 636 661
rect 659 639 664 666
rect 491 633 664 639
rect 786 639 791 667
rect 786 634 829 639
rect 491 610 496 633
rect 528 611 568 612
rect 490 609 497 610
rect 490 604 491 609
rect 496 604 497 609
rect 528 607 562 611
rect 490 603 497 604
rect 527 606 534 607
rect 527 601 528 606
rect 533 601 534 606
rect 561 606 562 607
rect 567 606 568 611
rect 600 611 636 616
rect 824 615 829 634
rect 561 605 568 606
rect 585 606 592 607
rect 527 600 534 601
rect 538 602 545 603
rect 538 597 539 602
rect 544 597 545 602
rect 585 601 586 606
rect 591 601 592 606
rect 600 605 601 611
rect 606 610 636 611
rect 606 605 607 610
rect 631 607 636 610
rect 823 614 830 615
rect 823 609 824 614
rect 829 609 830 614
rect 823 608 830 609
rect 849 607 854 736
rect 857 607 864 608
rect 600 604 607 605
rect 630 606 637 607
rect 630 601 631 606
rect 636 601 637 606
rect 659 605 666 606
rect 585 600 592 601
rect 614 600 621 601
rect 630 600 637 601
rect 643 600 649 601
rect 586 597 591 600
rect 538 592 591 597
rect 614 595 615 600
rect 620 595 621 600
rect 643 595 644 600
rect 648 595 649 600
rect 614 594 649 595
rect 615 590 649 594
rect 659 600 660 605
rect 665 600 666 605
rect 741 605 748 606
rect 741 600 742 605
rect 747 600 748 605
rect 837 602 858 607
rect 863 602 864 607
rect 837 601 849 602
rect 857 601 864 602
rect 659 599 666 600
rect 685 599 692 600
rect 741 599 748 600
rect 766 599 773 600
rect 659 594 686 599
rect 691 594 692 599
rect 742 594 767 599
rect 772 594 773 599
rect 659 573 664 594
rect 685 593 692 594
rect 766 593 773 594
rect 837 593 842 601
rect 492 567 664 573
rect 804 572 842 593
rect 492 547 497 567
rect 491 546 498 547
rect 491 541 492 546
rect 497 541 498 546
rect 491 540 498 541
rect 538 543 591 548
rect 615 546 649 550
rect 527 539 534 540
rect 527 534 528 539
rect 533 534 534 539
rect 538 538 539 543
rect 544 538 545 543
rect 586 540 591 543
rect 614 545 649 546
rect 614 540 615 545
rect 620 540 621 545
rect 643 540 644 545
rect 648 540 649 545
rect 538 537 545 538
rect 585 539 592 540
rect 614 539 621 540
rect 630 539 637 540
rect 643 539 649 540
rect 659 540 666 541
rect 527 533 534 534
rect 561 534 568 535
rect 561 533 562 534
rect 528 529 562 533
rect 567 529 568 534
rect 585 534 586 539
rect 591 534 592 539
rect 585 533 592 534
rect 600 535 607 536
rect 528 528 568 529
rect 600 529 601 535
rect 606 530 607 535
rect 630 534 631 539
rect 636 534 637 539
rect 659 535 660 540
rect 665 538 666 540
rect 685 538 692 539
rect 765 538 772 539
rect 665 535 686 538
rect 659 534 686 535
rect 630 533 637 534
rect 660 533 686 534
rect 691 533 692 538
rect 631 530 636 533
rect 606 529 636 530
rect 600 524 636 529
rect 660 507 665 533
rect 685 532 692 533
rect 742 533 766 538
rect 771 533 772 538
rect 491 501 665 507
rect 491 478 496 501
rect 528 479 568 480
rect 490 477 497 478
rect 490 472 491 477
rect 496 472 497 477
rect 528 475 562 479
rect 490 471 497 472
rect 527 474 534 475
rect 527 469 528 474
rect 533 469 534 474
rect 561 474 562 475
rect 567 474 568 479
rect 600 479 636 484
rect 742 482 747 533
rect 765 532 772 533
rect 561 473 568 474
rect 585 474 592 475
rect 527 468 534 469
rect 538 470 545 471
rect 538 465 539 470
rect 544 465 545 470
rect 585 469 586 474
rect 591 469 592 474
rect 600 473 601 479
rect 606 478 636 479
rect 606 473 607 478
rect 631 475 636 478
rect 741 481 748 482
rect 741 476 742 481
rect 747 476 748 481
rect 741 475 748 476
rect 600 472 607 473
rect 630 474 637 475
rect 630 469 631 474
rect 636 469 637 474
rect 659 473 666 474
rect 585 468 592 469
rect 614 468 621 469
rect 630 468 637 469
rect 643 468 649 469
rect 586 465 591 468
rect 538 460 591 465
rect 614 463 615 468
rect 620 463 621 468
rect 643 463 644 468
rect 648 463 649 468
rect 614 462 649 463
rect 615 458 649 462
rect 659 468 660 473
rect 665 468 666 473
rect 659 467 666 468
rect 685 467 692 468
rect 659 462 686 467
rect 691 462 692 467
rect 804 463 809 572
rect 854 534 861 535
rect 854 529 855 534
rect 860 529 861 534
rect 854 528 861 529
rect 761 462 809 463
rect 659 441 664 462
rect 685 461 692 462
rect 492 435 664 441
rect 730 457 809 462
rect 855 466 860 528
rect 855 460 922 466
rect 492 415 497 435
rect 491 414 498 415
rect 491 409 492 414
rect 497 409 498 414
rect 491 408 498 409
rect 538 411 591 416
rect 615 414 649 418
rect 730 414 735 457
rect 527 407 534 408
rect 527 402 528 407
rect 533 402 534 407
rect 538 406 539 411
rect 544 406 545 411
rect 586 408 591 411
rect 614 413 649 414
rect 614 408 615 413
rect 620 408 621 413
rect 643 408 644 413
rect 648 408 649 413
rect 729 413 736 414
rect 538 405 545 406
rect 585 407 592 408
rect 614 407 621 408
rect 630 407 637 408
rect 643 407 649 408
rect 659 408 666 409
rect 527 401 534 402
rect 561 402 568 403
rect 561 401 562 402
rect 528 397 562 401
rect 567 397 568 402
rect 585 402 586 407
rect 591 402 592 407
rect 585 401 592 402
rect 600 403 607 404
rect 528 396 568 397
rect 600 397 601 403
rect 606 398 607 403
rect 630 402 631 407
rect 636 402 637 407
rect 659 403 660 408
rect 665 403 666 408
rect 729 408 730 413
rect 735 408 736 413
rect 799 411 852 416
rect 876 414 910 418
rect 917 414 922 460
rect 729 407 736 408
rect 788 407 795 408
rect 659 402 666 403
rect 684 402 691 403
rect 630 401 637 402
rect 631 398 636 401
rect 606 397 636 398
rect 600 392 636 397
rect 661 397 685 402
rect 690 397 691 402
rect 788 402 789 407
rect 794 402 795 407
rect 799 406 800 411
rect 805 406 806 411
rect 847 408 852 411
rect 875 413 910 414
rect 875 408 876 413
rect 881 408 882 413
rect 904 408 905 413
rect 909 408 910 413
rect 799 405 806 406
rect 846 407 853 408
rect 875 407 882 408
rect 891 407 898 408
rect 904 407 910 408
rect 916 413 923 414
rect 916 408 917 413
rect 922 408 923 413
rect 916 407 923 408
rect 788 401 795 402
rect 822 402 829 403
rect 822 401 823 402
rect 408 48 414 49
rect 408 44 409 48
rect 413 44 414 48
rect 408 43 414 44
rect 661 37 666 397
rect 684 396 691 397
rect 789 397 823 401
rect 828 397 829 402
rect 846 402 847 407
rect 852 402 853 407
rect 846 401 853 402
rect 861 403 868 404
rect 789 396 829 397
rect 861 397 862 403
rect 867 398 868 403
rect 891 402 892 407
rect 897 402 898 407
rect 891 401 898 402
rect 892 398 897 401
rect 867 397 897 398
rect 861 392 897 397
rect 944 369 949 896
rect 1461 875 1501 876
rect 1422 873 1429 874
rect 1411 868 1429 873
rect 1461 871 1495 875
rect 1208 813 1214 814
rect 1208 809 1209 813
rect 1213 809 1346 813
rect 1208 808 1346 809
rect 952 413 958 414
rect 952 409 953 413
rect 957 409 958 413
rect 952 408 958 409
rect 791 364 949 369
rect 791 304 796 364
rect 790 303 796 304
rect 790 299 791 303
rect 795 299 796 303
rect 790 298 796 299
rect 953 241 958 408
rect 916 236 958 241
rect 916 222 921 236
rect 915 221 921 222
rect 915 217 916 221
rect 920 217 921 221
rect 915 216 921 217
rect 1341 49 1346 808
rect 1341 48 1347 49
rect 1341 44 1342 48
rect 1346 44 1347 48
rect 1341 43 1347 44
rect 1411 37 1416 868
rect 1422 867 1429 868
rect 1460 870 1467 871
rect 1460 865 1461 870
rect 1466 865 1467 870
rect 1494 870 1495 871
rect 1500 870 1501 875
rect 1533 875 1569 880
rect 1494 869 1501 870
rect 1518 870 1525 871
rect 1460 864 1467 865
rect 1471 866 1478 867
rect 1471 861 1472 866
rect 1477 861 1478 866
rect 1518 865 1519 870
rect 1524 865 1525 870
rect 1533 869 1534 875
rect 1539 874 1569 875
rect 1539 869 1540 874
rect 1564 871 1569 874
rect 1533 868 1540 869
rect 1563 870 1570 871
rect 1563 865 1564 870
rect 1569 865 1570 870
rect 1592 869 1599 870
rect 1518 864 1525 865
rect 1547 864 1554 865
rect 1563 864 1570 865
rect 1576 864 1582 865
rect 1519 861 1524 864
rect 1471 856 1524 861
rect 1547 859 1548 864
rect 1553 859 1554 864
rect 1576 859 1577 864
rect 1581 859 1582 864
rect 1547 858 1582 859
rect 1548 854 1582 858
rect 1592 864 1593 869
rect 1598 864 1599 869
rect 1674 869 1681 870
rect 1674 864 1675 869
rect 1680 864 1681 869
rect 1759 869 1766 870
rect 1759 864 1760 869
rect 1765 864 1766 869
rect 1592 863 1599 864
rect 1618 863 1625 864
rect 1674 863 1681 864
rect 1699 863 1706 864
rect 1759 863 1766 864
rect 1592 858 1619 863
rect 1624 858 1625 863
rect 1675 858 1700 863
rect 1705 858 1706 863
rect 1592 837 1597 858
rect 1618 857 1625 858
rect 1699 857 1706 858
rect 1756 858 1765 863
rect 1425 831 1597 837
rect 1425 811 1430 831
rect 1424 810 1431 811
rect 1424 805 1425 810
rect 1430 805 1431 810
rect 1424 804 1431 805
rect 1471 807 1524 812
rect 1548 810 1582 814
rect 1460 803 1467 804
rect 1460 798 1461 803
rect 1466 798 1467 803
rect 1471 802 1472 807
rect 1477 802 1478 807
rect 1519 804 1524 807
rect 1547 809 1582 810
rect 1547 804 1548 809
rect 1553 804 1554 809
rect 1576 804 1577 809
rect 1581 804 1582 809
rect 1471 801 1478 802
rect 1518 803 1525 804
rect 1547 803 1554 804
rect 1563 803 1570 804
rect 1576 803 1582 804
rect 1592 804 1599 805
rect 1618 804 1625 805
rect 1698 804 1705 805
rect 1460 797 1467 798
rect 1494 798 1501 799
rect 1494 797 1495 798
rect 1461 793 1495 797
rect 1500 793 1501 798
rect 1518 798 1519 803
rect 1524 798 1525 803
rect 1518 797 1525 798
rect 1533 799 1540 800
rect 1461 792 1501 793
rect 1533 793 1534 799
rect 1539 794 1540 799
rect 1563 798 1564 803
rect 1569 798 1570 803
rect 1592 799 1593 804
rect 1598 799 1619 804
rect 1624 799 1625 804
rect 1592 798 1599 799
rect 1618 798 1625 799
rect 1675 799 1699 804
rect 1704 799 1705 804
rect 1563 797 1570 798
rect 1564 794 1569 797
rect 1539 793 1569 794
rect 1533 788 1569 793
rect 1593 771 1598 798
rect 1424 765 1598 771
rect 1424 742 1429 765
rect 1461 743 1501 744
rect 1423 741 1430 742
rect 1423 736 1424 741
rect 1429 736 1430 741
rect 1461 739 1495 743
rect 1423 735 1430 736
rect 1460 738 1467 739
rect 1460 733 1461 738
rect 1466 733 1467 738
rect 1494 738 1495 739
rect 1500 738 1501 743
rect 1533 743 1569 748
rect 1675 746 1680 799
rect 1698 798 1705 799
rect 1756 770 1761 858
rect 1718 765 1761 770
rect 1494 737 1501 738
rect 1518 738 1525 739
rect 1460 732 1467 733
rect 1471 734 1478 735
rect 1471 729 1472 734
rect 1477 729 1478 734
rect 1518 733 1519 738
rect 1524 733 1525 738
rect 1533 737 1534 743
rect 1539 742 1569 743
rect 1539 737 1540 742
rect 1564 739 1569 742
rect 1674 745 1681 746
rect 1674 740 1675 745
rect 1680 740 1681 745
rect 1674 739 1681 740
rect 1533 736 1540 737
rect 1563 738 1570 739
rect 1563 733 1564 738
rect 1569 733 1570 738
rect 1592 737 1599 738
rect 1518 732 1525 733
rect 1547 732 1554 733
rect 1563 732 1570 733
rect 1576 732 1582 733
rect 1519 729 1524 732
rect 1471 724 1524 729
rect 1547 727 1548 732
rect 1553 727 1554 732
rect 1576 727 1577 732
rect 1581 727 1582 732
rect 1547 726 1582 727
rect 1548 722 1582 726
rect 1592 732 1593 737
rect 1598 732 1599 737
rect 1718 732 1723 765
rect 1781 742 1788 743
rect 1781 737 1782 742
rect 1787 737 1788 742
rect 1781 736 1788 737
rect 1592 731 1599 732
rect 1618 731 1625 732
rect 1592 726 1619 731
rect 1624 726 1625 731
rect 1718 731 1730 732
rect 1718 726 1724 731
rect 1729 726 1730 731
rect 1592 705 1597 726
rect 1618 725 1625 726
rect 1723 725 1730 726
rect 1425 699 1597 705
rect 1425 679 1430 699
rect 1424 678 1431 679
rect 1424 673 1425 678
rect 1430 673 1431 678
rect 1424 672 1431 673
rect 1471 675 1524 680
rect 1548 678 1582 682
rect 1460 671 1467 672
rect 1460 666 1461 671
rect 1466 666 1467 671
rect 1471 670 1472 675
rect 1477 670 1478 675
rect 1519 672 1524 675
rect 1547 677 1582 678
rect 1547 672 1548 677
rect 1553 672 1554 677
rect 1576 672 1577 677
rect 1581 672 1582 677
rect 1617 673 1624 674
rect 1723 673 1730 674
rect 1471 669 1478 670
rect 1518 671 1525 672
rect 1547 671 1554 672
rect 1563 671 1570 672
rect 1576 671 1582 672
rect 1592 672 1618 673
rect 1460 665 1467 666
rect 1494 666 1501 667
rect 1494 665 1495 666
rect 1461 661 1495 665
rect 1500 661 1501 666
rect 1518 666 1519 671
rect 1524 666 1525 671
rect 1518 665 1525 666
rect 1533 667 1540 668
rect 1461 660 1501 661
rect 1533 661 1534 667
rect 1539 662 1540 667
rect 1563 666 1564 671
rect 1569 666 1570 671
rect 1563 665 1570 666
rect 1592 667 1593 672
rect 1598 668 1618 672
rect 1623 668 1624 673
rect 1598 667 1599 668
rect 1617 667 1624 668
rect 1719 668 1724 673
rect 1729 668 1730 673
rect 1719 667 1730 668
rect 1592 666 1599 667
rect 1564 662 1569 665
rect 1539 661 1569 662
rect 1533 656 1569 661
rect 1592 639 1597 666
rect 1424 633 1597 639
rect 1719 639 1724 667
rect 1719 634 1762 639
rect 1424 610 1429 633
rect 1461 611 1501 612
rect 1423 609 1430 610
rect 1423 604 1424 609
rect 1429 604 1430 609
rect 1461 607 1495 611
rect 1423 603 1430 604
rect 1460 606 1467 607
rect 1460 601 1461 606
rect 1466 601 1467 606
rect 1494 606 1495 607
rect 1500 606 1501 611
rect 1533 611 1569 616
rect 1757 615 1762 634
rect 1494 605 1501 606
rect 1518 606 1525 607
rect 1460 600 1467 601
rect 1471 602 1478 603
rect 1471 597 1472 602
rect 1477 597 1478 602
rect 1518 601 1519 606
rect 1524 601 1525 606
rect 1533 605 1534 611
rect 1539 610 1569 611
rect 1539 605 1540 610
rect 1564 607 1569 610
rect 1756 614 1763 615
rect 1756 609 1757 614
rect 1762 609 1763 614
rect 1756 608 1763 609
rect 1782 607 1787 736
rect 1790 607 1797 608
rect 1533 604 1540 605
rect 1563 606 1570 607
rect 1563 601 1564 606
rect 1569 601 1570 606
rect 1592 605 1599 606
rect 1518 600 1525 601
rect 1547 600 1554 601
rect 1563 600 1570 601
rect 1576 600 1582 601
rect 1519 597 1524 600
rect 1471 592 1524 597
rect 1547 595 1548 600
rect 1553 595 1554 600
rect 1576 595 1577 600
rect 1581 595 1582 600
rect 1547 594 1582 595
rect 1548 590 1582 594
rect 1592 600 1593 605
rect 1598 600 1599 605
rect 1674 605 1681 606
rect 1674 600 1675 605
rect 1680 600 1681 605
rect 1770 602 1791 607
rect 1796 602 1797 607
rect 1770 601 1782 602
rect 1790 601 1797 602
rect 1592 599 1599 600
rect 1618 599 1625 600
rect 1674 599 1681 600
rect 1699 599 1706 600
rect 1592 594 1619 599
rect 1624 594 1625 599
rect 1675 594 1700 599
rect 1705 594 1706 599
rect 1592 573 1597 594
rect 1618 593 1625 594
rect 1699 593 1706 594
rect 1770 593 1775 601
rect 1425 567 1597 573
rect 1737 572 1775 593
rect 1425 547 1430 567
rect 1424 546 1431 547
rect 1424 541 1425 546
rect 1430 541 1431 546
rect 1424 540 1431 541
rect 1471 543 1524 548
rect 1548 546 1582 550
rect 1460 539 1467 540
rect 1460 534 1461 539
rect 1466 534 1467 539
rect 1471 538 1472 543
rect 1477 538 1478 543
rect 1519 540 1524 543
rect 1547 545 1582 546
rect 1547 540 1548 545
rect 1553 540 1554 545
rect 1576 540 1577 545
rect 1581 540 1582 545
rect 1471 537 1478 538
rect 1518 539 1525 540
rect 1547 539 1554 540
rect 1563 539 1570 540
rect 1576 539 1582 540
rect 1592 540 1599 541
rect 1460 533 1467 534
rect 1494 534 1501 535
rect 1494 533 1495 534
rect 1461 529 1495 533
rect 1500 529 1501 534
rect 1518 534 1519 539
rect 1524 534 1525 539
rect 1518 533 1525 534
rect 1533 535 1540 536
rect 1461 528 1501 529
rect 1533 529 1534 535
rect 1539 530 1540 535
rect 1563 534 1564 539
rect 1569 534 1570 539
rect 1592 535 1593 540
rect 1598 538 1599 540
rect 1618 538 1625 539
rect 1698 538 1705 539
rect 1598 535 1619 538
rect 1592 534 1619 535
rect 1563 533 1570 534
rect 1593 533 1619 534
rect 1624 533 1625 538
rect 1564 530 1569 533
rect 1539 529 1569 530
rect 1533 524 1569 529
rect 1593 507 1598 533
rect 1618 532 1625 533
rect 1675 533 1699 538
rect 1704 533 1705 538
rect 1424 501 1598 507
rect 1424 478 1429 501
rect 1461 479 1501 480
rect 1423 477 1430 478
rect 1423 472 1424 477
rect 1429 472 1430 477
rect 1461 475 1495 479
rect 1423 471 1430 472
rect 1460 474 1467 475
rect 1460 469 1461 474
rect 1466 469 1467 474
rect 1494 474 1495 475
rect 1500 474 1501 479
rect 1533 479 1569 484
rect 1675 482 1680 533
rect 1698 532 1705 533
rect 1494 473 1501 474
rect 1518 474 1525 475
rect 1460 468 1467 469
rect 1471 470 1478 471
rect 1471 465 1472 470
rect 1477 465 1478 470
rect 1518 469 1519 474
rect 1524 469 1525 474
rect 1533 473 1534 479
rect 1539 478 1569 479
rect 1539 473 1540 478
rect 1564 475 1569 478
rect 1674 481 1681 482
rect 1674 476 1675 481
rect 1680 476 1681 481
rect 1674 475 1681 476
rect 1533 472 1540 473
rect 1563 474 1570 475
rect 1563 469 1564 474
rect 1569 469 1570 474
rect 1592 473 1599 474
rect 1518 468 1525 469
rect 1547 468 1554 469
rect 1563 468 1570 469
rect 1576 468 1582 469
rect 1519 465 1524 468
rect 1471 460 1524 465
rect 1547 463 1548 468
rect 1553 463 1554 468
rect 1576 463 1577 468
rect 1581 463 1582 468
rect 1547 462 1582 463
rect 1548 458 1582 462
rect 1592 468 1593 473
rect 1598 468 1599 473
rect 1592 467 1599 468
rect 1618 467 1625 468
rect 1592 462 1619 467
rect 1624 462 1625 467
rect 1737 463 1742 572
rect 1787 534 1794 535
rect 1787 529 1788 534
rect 1793 529 1794 534
rect 1787 528 1794 529
rect 1694 462 1742 463
rect 1592 441 1597 462
rect 1618 461 1625 462
rect 1425 435 1597 441
rect 1663 457 1742 462
rect 1788 466 1793 528
rect 1788 460 1855 466
rect 1425 415 1430 435
rect 1424 414 1431 415
rect 1424 409 1425 414
rect 1430 409 1431 414
rect 1424 408 1431 409
rect 1471 411 1524 416
rect 1548 414 1582 418
rect 1663 414 1668 457
rect 1460 407 1467 408
rect 1460 402 1461 407
rect 1466 402 1467 407
rect 1471 406 1472 411
rect 1477 406 1478 411
rect 1519 408 1524 411
rect 1547 413 1582 414
rect 1547 408 1548 413
rect 1553 408 1554 413
rect 1576 408 1577 413
rect 1581 408 1582 413
rect 1662 413 1669 414
rect 1471 405 1478 406
rect 1518 407 1525 408
rect 1547 407 1554 408
rect 1563 407 1570 408
rect 1576 407 1582 408
rect 1592 408 1599 409
rect 1460 401 1467 402
rect 1494 402 1501 403
rect 1494 401 1495 402
rect 1461 397 1495 401
rect 1500 397 1501 402
rect 1518 402 1519 407
rect 1524 402 1525 407
rect 1518 401 1525 402
rect 1533 403 1540 404
rect 1461 396 1501 397
rect 1533 397 1534 403
rect 1539 398 1540 403
rect 1563 402 1564 407
rect 1569 402 1570 407
rect 1592 403 1593 408
rect 1598 403 1599 408
rect 1662 408 1663 413
rect 1668 408 1669 413
rect 1732 411 1785 416
rect 1809 414 1843 418
rect 1850 414 1855 460
rect 1662 407 1669 408
rect 1721 407 1728 408
rect 1592 402 1599 403
rect 1617 402 1624 403
rect 1563 401 1570 402
rect 1564 398 1569 401
rect 1539 397 1569 398
rect 1594 397 1618 402
rect 1623 397 1624 402
rect 1721 402 1722 407
rect 1727 402 1728 407
rect 1732 406 1733 411
rect 1738 406 1739 411
rect 1780 408 1785 411
rect 1808 413 1843 414
rect 1808 408 1809 413
rect 1814 408 1815 413
rect 1837 408 1838 413
rect 1842 408 1843 413
rect 1732 405 1739 406
rect 1779 407 1786 408
rect 1808 407 1815 408
rect 1824 407 1831 408
rect 1837 407 1843 408
rect 1849 413 1856 414
rect 1849 408 1850 413
rect 1855 408 1856 413
rect 1849 407 1856 408
rect 1721 401 1728 402
rect 1755 402 1762 403
rect 1755 401 1756 402
rect 1533 392 1569 397
rect 1617 396 1624 397
rect 1722 397 1756 401
rect 1761 397 1762 402
rect 1779 402 1780 407
rect 1785 402 1786 407
rect 1779 401 1786 402
rect 1794 403 1801 404
rect 1722 396 1762 397
rect 1794 397 1795 403
rect 1800 398 1801 403
rect 1824 402 1825 407
rect 1830 402 1831 407
rect 1824 401 1831 402
rect 1825 398 1830 401
rect 1800 397 1830 398
rect 1794 392 1830 397
rect 1877 369 1882 896
rect 1724 364 1882 369
rect 1895 413 1951 418
rect 1724 304 1729 364
rect 1723 303 1729 304
rect 1723 299 1724 303
rect 1728 299 1729 303
rect 1723 298 1729 299
rect 1895 241 1900 413
rect 1849 236 1900 241
rect 1849 222 1854 236
rect 1848 221 1854 222
rect 1848 217 1849 221
rect 1853 217 1854 221
rect 1848 216 1854 217
rect 661 32 1416 37
<< labels >>
rlabel metal2 1364 1971 1364 1971 1 GND!
rlabel metal2 1352 1971 1352 1971 1 Vdd!
rlabel metal2 1377 1970 1377 1970 4 f_clk_b
rlabel metal2 1389 1969 1389 1969 5 f_clk
rlabel metal2 1413 1970 1413 1970 5 p_clk
rlabel metal2 1401 1970 1401 1970 5 p_clk_b
rlabel metal2 431 1971 431 1971 1 GND!
rlabel metal2 419 1971 419 1971 1 Vdd!
rlabel metal2 444 1970 444 1970 4 f_clk_b
rlabel metal2 456 1969 456 1969 5 f_clk
rlabel metal2 480 1970 480 1970 5 p_clk
rlabel metal2 468 1970 468 1970 5 p_clk_b
rlabel metal2 153 1970 153 1970 1 in
rlabel metal1 1929 120 1929 120 1 out
rlabel m3contact 22 1391 22 1391 1 p_in
rlabel metal1 1280 1846 1280 1846 1 3
rlabel metal2 926 1361 926 1361 1 2
rlabel metal2 1860 1366 1860 1366 1 4
rlabel metal1 364 865 364 865 1 5
rlabel metal2 926 384 926 384 1 6
rlabel metal1 1274 865 1274 865 1 7
rlabel metal2 1859 380 1859 380 1 8
rlabel polysilicon 165 1840 165 1840 1 CB_1
rlabel polysilicon 931 1338 931 1338 1 CB_2
rlabel polysilicon 1074 1341 1074 1341 1 S_1
rlabel polysilicon 1098 1840 1098 1840 1 CB_3
rlabel polysilicon 1876 1194 1876 1194 1 CB_4
rlabel polysilicon 1211 1096 1211 1096 1 S_2
rlabel polysilicon 282 1080 282 1080 1 S_3
rlabel polysilicon 282 863 282 863 1 CB_5
rlabel polysilicon 931 358 931 358 1 CB_6
rlabel polysilicon 1074 354 1074 354 1 S_4
rlabel polysilicon 1098 854 1098 854 1 CB_7
rlabel polysilicon 1876 214 1876 214 1 CB_8
<< end >>
