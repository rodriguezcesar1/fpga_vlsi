magic
tech scmos
timestamp 1608351510
<< nwell >>
rect 1060 10033 1320 10293
rect 1369 10033 1629 10293
rect 1678 10033 1938 10293
rect 1987 10033 2247 10293
rect 2296 10033 2556 10293
rect 2605 10033 2865 10293
rect 2914 10033 3174 10293
rect 3223 10033 3483 10293
rect 3532 10033 3792 10293
rect 3841 10033 4101 10293
rect 86 9047 346 9307
rect 4826 9059 5086 9319
rect 86 8738 346 8998
rect 4826 8750 5086 9010
rect 86 8429 346 8689
rect 4826 8441 5086 8701
rect 86 8120 346 8380
rect 4826 8132 5086 8392
rect 86 7811 346 8071
rect 4826 7824 5086 8084
rect 86 7502 346 7762
rect 4826 7515 5086 7775
rect 86 7193 346 7453
rect 4826 7233 5086 7493
rect 86 6849 346 7109
rect 4826 6861 5086 7121
rect 86 6539 346 6799
rect 4826 6552 5086 6812
rect 86 6230 346 6490
rect 4826 6243 5086 6503
rect 86 5922 346 6182
rect 4826 5934 5086 6194
rect 86 5613 346 5873
rect 4826 5625 5086 5885
rect 86 5304 346 5564
rect 4826 5316 5086 5576
rect 86 4995 346 5255
rect 4826 5007 5086 5267
rect 1071 4021 1331 4281
rect 1380 4021 1640 4281
rect 1689 4021 1949 4281
rect 1998 4021 2258 4281
rect 2307 4021 2567 4281
rect 2616 4021 2876 4281
rect 2925 4021 3185 4281
rect 3234 4021 3494 4281
rect 3543 4021 3803 4281
rect 3852 4021 4112 4281
<< ntransistor >>
rect 1829 9824 1869 9826
rect 2138 9824 2178 9826
rect 2447 9824 2487 9826
rect 2756 9824 2796 9826
rect 3065 9824 3105 9826
rect 3992 9824 4032 9826
rect 1829 9816 1869 9818
rect 2138 9816 2178 9818
rect 2447 9816 2487 9818
rect 2756 9816 2796 9818
rect 3065 9816 3105 9818
rect 3992 9816 4032 9818
rect 1829 9808 1869 9810
rect 1829 9800 1869 9802
rect 1829 9792 1869 9794
rect 1829 9784 1869 9786
rect 2138 9808 2178 9810
rect 2138 9800 2178 9802
rect 2138 9792 2178 9794
rect 2138 9784 2178 9786
rect 2447 9808 2487 9810
rect 2447 9800 2487 9802
rect 2447 9792 2487 9794
rect 2447 9784 2487 9786
rect 2756 9808 2796 9810
rect 2756 9800 2796 9802
rect 2756 9792 2796 9794
rect 2756 9784 2796 9786
rect 3065 9808 3105 9810
rect 3065 9800 3105 9802
rect 3065 9792 3105 9794
rect 3065 9784 3105 9786
rect 3992 9808 4032 9810
rect 3992 9800 4032 9802
rect 3992 9792 4032 9794
rect 3992 9784 4032 9786
rect 428 6280 430 6339
rect 436 6280 438 6339
rect 444 6280 446 6339
rect 452 6280 454 6339
rect 469 6280 471 6339
rect 477 6280 479 6339
rect 485 6280 487 6339
rect 493 6280 495 6339
rect 512 6280 514 6339
rect 520 6280 522 6339
rect 528 6280 530 6339
rect 536 6280 538 6339
rect 551 6299 553 6339
rect 559 6299 561 6339
rect 567 6299 569 6339
rect 575 6299 577 6339
rect 583 6299 585 6339
rect 591 6299 593 6339
rect 2856 9299 2858 9303
rect 2861 9299 2863 9303
rect 2877 9299 2879 9303
rect 2893 9299 2895 9303
rect 2898 9299 2900 9303
rect 2919 9299 2921 9303
rect 2935 9299 2937 9303
rect 2951 9299 2953 9303
rect 2956 9299 2958 9303
rect 2972 9299 2974 9303
rect 2988 9299 2990 9303
rect 2993 9299 2995 9303
rect 3009 9299 3011 9303
rect 3025 9299 3027 9303
rect 3030 9299 3032 9303
rect 3051 9299 3053 9303
rect 3067 9299 3069 9303
rect 3083 9299 3085 9303
rect 3088 9299 3090 9303
rect 3104 9299 3106 9303
rect 3120 9299 3122 9303
rect 3125 9299 3127 9303
rect 3141 9299 3143 9303
rect 3157 9299 3159 9303
rect 3162 9299 3164 9303
rect 3183 9299 3185 9303
rect 3199 9299 3201 9303
rect 3215 9299 3217 9303
rect 3220 9299 3222 9303
rect 3236 9299 3238 9303
rect 3252 9299 3254 9303
rect 3257 9299 3259 9303
rect 3273 9299 3275 9303
rect 3289 9299 3291 9303
rect 3294 9299 3296 9303
rect 3315 9299 3317 9303
rect 3331 9299 3333 9303
rect 3347 9299 3349 9303
rect 3352 9299 3354 9303
rect 3368 9299 3370 9303
rect 3801 9299 3803 9303
rect 3806 9299 3808 9303
rect 3822 9299 3824 9303
rect 3838 9299 3840 9303
rect 3843 9299 3845 9303
rect 3864 9299 3866 9303
rect 3880 9299 3882 9303
rect 3896 9299 3898 9303
rect 3901 9299 3903 9303
rect 3917 9299 3919 9303
rect 3933 9299 3935 9303
rect 3938 9299 3940 9303
rect 3954 9299 3956 9303
rect 3970 9299 3972 9303
rect 3975 9299 3977 9303
rect 3996 9299 3998 9303
rect 4012 9299 4014 9303
rect 4028 9299 4030 9303
rect 4033 9299 4035 9303
rect 4049 9299 4051 9303
rect 4065 9299 4067 9303
rect 4070 9299 4072 9303
rect 4086 9299 4088 9303
rect 4102 9299 4104 9303
rect 4107 9299 4109 9303
rect 4128 9299 4130 9303
rect 4144 9299 4146 9303
rect 4160 9299 4162 9303
rect 4165 9299 4167 9303
rect 4181 9299 4183 9303
rect 4197 9299 4199 9303
rect 4202 9299 4204 9303
rect 4218 9299 4220 9303
rect 4234 9299 4236 9303
rect 4239 9299 4241 9303
rect 4260 9299 4262 9303
rect 4276 9299 4278 9303
rect 4292 9299 4294 9303
rect 4297 9299 4299 9303
rect 4313 9299 4315 9303
rect 2504 9266 2506 9270
rect 2509 9266 2511 9270
rect 2525 9266 2527 9270
rect 2541 9266 2543 9270
rect 2546 9266 2548 9270
rect 2567 9266 2569 9270
rect 2583 9266 2585 9270
rect 2599 9266 2601 9270
rect 2604 9266 2606 9270
rect 2620 9266 2622 9270
rect 3449 9266 3451 9270
rect 3454 9266 3456 9270
rect 3470 9266 3472 9270
rect 3486 9266 3488 9270
rect 3491 9266 3493 9270
rect 3512 9266 3514 9270
rect 3528 9266 3530 9270
rect 3544 9266 3546 9270
rect 3549 9266 3551 9270
rect 3565 9266 3567 9270
rect 2628 9229 2630 9233
rect 3035 9233 3037 9237
rect 3061 9229 3063 9233
rect 3066 9229 3068 9233
rect 3116 9233 3118 9237
rect 3142 9229 3144 9233
rect 3147 9229 3149 9233
rect 3089 9225 3091 9229
rect 2511 9220 2513 9224
rect 2861 9220 2863 9224
rect 2877 9220 2879 9224
rect 2893 9220 2895 9224
rect 2916 9220 2918 9224
rect 2921 9220 2923 9224
rect 2947 9220 2949 9224
rect 2968 9220 2970 9224
rect 2988 9220 2990 9224
rect 2993 9220 2995 9224
rect 3011 9220 3013 9224
rect 3170 9225 3172 9229
rect 3573 9229 3575 9233
rect 3980 9233 3982 9237
rect 4006 9229 4008 9233
rect 4011 9229 4013 9233
rect 4061 9233 4063 9237
rect 4087 9229 4089 9233
rect 4092 9229 4094 9233
rect 4034 9225 4036 9229
rect 3456 9220 3458 9224
rect 3806 9220 3808 9224
rect 3822 9220 3824 9224
rect 3838 9220 3840 9224
rect 3861 9220 3863 9224
rect 3866 9220 3868 9224
rect 3892 9220 3894 9224
rect 3913 9220 3915 9224
rect 3933 9220 3935 9224
rect 3938 9220 3940 9224
rect 3956 9220 3958 9224
rect 4115 9225 4117 9229
rect 2861 9174 2863 9178
rect 2877 9174 2879 9178
rect 2893 9174 2895 9178
rect 2916 9174 2918 9178
rect 2921 9174 2923 9178
rect 2947 9174 2949 9178
rect 2968 9174 2970 9178
rect 2988 9174 2990 9178
rect 2993 9174 2995 9178
rect 3011 9174 3013 9178
rect 2495 9164 2497 9168
rect 2511 9164 2513 9168
rect 2516 9164 2518 9168
rect 2532 9164 2534 9168
rect 2548 9164 2550 9168
rect 2569 9164 2571 9168
rect 2574 9164 2576 9168
rect 2590 9164 2592 9168
rect 2606 9164 2608 9168
rect 2611 9164 2613 9168
rect 3061 9173 3063 9177
rect 3066 9173 3068 9177
rect 3142 9173 3144 9177
rect 3147 9173 3149 9177
rect 3806 9174 3808 9178
rect 3822 9174 3824 9178
rect 3838 9174 3840 9178
rect 3861 9174 3863 9178
rect 3866 9174 3868 9178
rect 3892 9174 3894 9178
rect 3913 9174 3915 9178
rect 3933 9174 3935 9178
rect 3938 9174 3940 9178
rect 3956 9174 3958 9178
rect 3440 9164 3442 9168
rect 3456 9164 3458 9168
rect 3461 9164 3463 9168
rect 3477 9164 3479 9168
rect 3493 9164 3495 9168
rect 3514 9164 3516 9168
rect 3519 9164 3521 9168
rect 3535 9164 3537 9168
rect 3551 9164 3553 9168
rect 3556 9164 3558 9168
rect 4006 9173 4008 9177
rect 4011 9173 4013 9177
rect 4087 9173 4089 9177
rect 4092 9173 4094 9177
rect 3061 9097 3063 9101
rect 3066 9097 3068 9101
rect 3140 9101 3142 9105
rect 3166 9097 3168 9101
rect 3171 9097 3173 9101
rect 3089 9093 3091 9097
rect 2861 9088 2863 9092
rect 2877 9088 2879 9092
rect 2893 9088 2895 9092
rect 2916 9088 2918 9092
rect 2921 9088 2923 9092
rect 2947 9088 2949 9092
rect 2968 9088 2970 9092
rect 2988 9088 2990 9092
rect 2993 9088 2995 9092
rect 3011 9088 3013 9092
rect 3194 9093 3196 9097
rect 3371 9072 3373 9076
rect 3397 9068 3399 9072
rect 3402 9068 3404 9072
rect 3425 9064 3427 9068
rect 4006 9097 4008 9101
rect 4011 9097 4013 9101
rect 4085 9101 4087 9105
rect 4111 9097 4113 9101
rect 4116 9097 4118 9101
rect 4034 9093 4036 9097
rect 3806 9088 3808 9092
rect 3822 9088 3824 9092
rect 3838 9088 3840 9092
rect 3861 9088 3863 9092
rect 3866 9088 3868 9092
rect 3892 9088 3894 9092
rect 3913 9088 3915 9092
rect 3933 9088 3935 9092
rect 3938 9088 3940 9092
rect 3956 9088 3958 9092
rect 4139 9093 4141 9097
rect 2861 9042 2863 9046
rect 2877 9042 2879 9046
rect 2893 9042 2895 9046
rect 2916 9042 2918 9046
rect 2921 9042 2923 9046
rect 2947 9042 2949 9046
rect 2968 9042 2970 9046
rect 2988 9042 2990 9046
rect 2993 9042 2995 9046
rect 3011 9042 3013 9046
rect 3061 9042 3063 9046
rect 3066 9042 3068 9046
rect 3166 9042 3168 9046
rect 3171 9042 3173 9046
rect 3557 9033 3559 9045
rect 3610 9033 3612 9045
rect 3806 9042 3808 9046
rect 3822 9042 3824 9046
rect 3838 9042 3840 9046
rect 3861 9042 3863 9046
rect 3866 9042 3868 9046
rect 3892 9042 3894 9046
rect 3913 9042 3915 9046
rect 3933 9042 3935 9046
rect 3938 9042 3940 9046
rect 3956 9042 3958 9046
rect 4006 9042 4008 9046
rect 4011 9042 4013 9046
rect 4111 9042 4113 9046
rect 4116 9042 4118 9046
rect 3397 9008 3399 9012
rect 3402 9008 3404 9012
rect 3061 8965 3063 8969
rect 3066 8965 3068 8969
rect 3116 8969 3118 8973
rect 3142 8965 3144 8969
rect 3147 8965 3149 8969
rect 3206 8969 3208 8973
rect 3232 8965 3234 8969
rect 3237 8965 3239 8969
rect 3089 8961 3091 8965
rect 2861 8956 2863 8960
rect 2877 8956 2879 8960
rect 2893 8956 2895 8960
rect 2916 8956 2918 8960
rect 2921 8956 2923 8960
rect 2947 8956 2949 8960
rect 2968 8956 2970 8960
rect 2988 8956 2990 8960
rect 2993 8956 2995 8960
rect 3011 8956 3013 8960
rect 3170 8961 3172 8965
rect 3260 8961 3262 8965
rect 3349 8942 3351 8946
rect 3371 8942 3373 8946
rect 3397 8938 3399 8942
rect 3402 8938 3404 8942
rect 3425 8934 3427 8938
rect 4006 8965 4008 8969
rect 4011 8965 4013 8969
rect 4061 8969 4063 8973
rect 4087 8965 4089 8969
rect 4092 8965 4094 8969
rect 4151 8969 4153 8973
rect 4177 8965 4179 8969
rect 4182 8965 4184 8969
rect 4034 8961 4036 8965
rect 3806 8956 3808 8960
rect 3822 8956 3824 8960
rect 3838 8956 3840 8960
rect 3861 8956 3863 8960
rect 3866 8956 3868 8960
rect 3892 8956 3894 8960
rect 3913 8956 3915 8960
rect 3933 8956 3935 8960
rect 3938 8956 3940 8960
rect 3956 8956 3958 8960
rect 4115 8961 4117 8965
rect 4205 8961 4207 8965
rect 2861 8910 2863 8914
rect 2877 8910 2879 8914
rect 2893 8910 2895 8914
rect 2916 8910 2918 8914
rect 2921 8910 2923 8914
rect 2947 8910 2949 8914
rect 2968 8910 2970 8914
rect 2988 8910 2990 8914
rect 2993 8910 2995 8914
rect 3011 8910 3013 8914
rect 3061 8907 3063 8911
rect 3066 8907 3068 8911
rect 3142 8907 3144 8911
rect 3147 8907 3149 8911
rect 3232 8907 3234 8911
rect 3237 8907 3239 8911
rect 3463 8903 3465 8915
rect 3516 8903 3518 8915
rect 3806 8910 3808 8914
rect 3822 8910 3824 8914
rect 3838 8910 3840 8914
rect 3861 8910 3863 8914
rect 3866 8910 3868 8914
rect 3892 8910 3894 8914
rect 3913 8910 3915 8914
rect 3933 8910 3935 8914
rect 3938 8910 3940 8914
rect 3956 8910 3958 8914
rect 4006 8907 4008 8911
rect 4011 8907 4013 8911
rect 4087 8907 4089 8911
rect 4092 8907 4094 8911
rect 4177 8907 4179 8911
rect 4182 8907 4184 8911
rect 3397 8878 3399 8882
rect 3402 8878 3404 8882
rect 3061 8833 3063 8837
rect 3066 8833 3068 8837
rect 3089 8829 3091 8833
rect 2861 8824 2863 8828
rect 2877 8824 2879 8828
rect 2893 8824 2895 8828
rect 2916 8824 2918 8828
rect 2921 8824 2923 8828
rect 2947 8824 2949 8828
rect 2968 8824 2970 8828
rect 2988 8824 2990 8828
rect 2993 8824 2995 8828
rect 3011 8824 3013 8828
rect 4006 8833 4008 8837
rect 4011 8833 4013 8837
rect 4034 8829 4036 8833
rect 3806 8824 3808 8828
rect 3822 8824 3824 8828
rect 3838 8824 3840 8828
rect 3861 8824 3863 8828
rect 3866 8824 3868 8828
rect 3892 8824 3894 8828
rect 3913 8824 3915 8828
rect 3933 8824 3935 8828
rect 3938 8824 3940 8828
rect 3956 8824 3958 8828
rect 2861 8778 2863 8782
rect 2877 8778 2879 8782
rect 2893 8778 2895 8782
rect 2916 8778 2918 8782
rect 2921 8778 2923 8782
rect 2947 8778 2949 8782
rect 2968 8778 2970 8782
rect 2988 8778 2990 8782
rect 2993 8778 2995 8782
rect 3011 8778 3013 8782
rect 3095 8778 3097 8782
rect 3113 8778 3115 8782
rect 3138 8778 3140 8782
rect 3154 8778 3156 8782
rect 3177 8778 3179 8782
rect 3182 8778 3184 8782
rect 3208 8778 3210 8782
rect 3229 8778 3231 8782
rect 3249 8778 3251 8782
rect 3254 8778 3256 8782
rect 3272 8778 3274 8782
rect 2372 8764 2374 8768
rect 2377 8764 2379 8768
rect 2393 8764 2395 8768
rect 2409 8764 2411 8768
rect 2414 8764 2416 8768
rect 2435 8764 2437 8768
rect 2451 8764 2453 8768
rect 2467 8764 2469 8768
rect 2472 8764 2474 8768
rect 2488 8764 2490 8768
rect 2504 8764 2506 8768
rect 2509 8764 2511 8768
rect 2525 8764 2527 8768
rect 2541 8764 2543 8768
rect 2546 8764 2548 8768
rect 2567 8764 2569 8768
rect 2583 8764 2585 8768
rect 2599 8764 2601 8768
rect 2604 8764 2606 8768
rect 2620 8764 2622 8768
rect 2636 8764 2638 8768
rect 2641 8764 2643 8768
rect 2657 8764 2659 8768
rect 2673 8764 2675 8768
rect 2678 8764 2680 8768
rect 2699 8764 2701 8768
rect 2715 8764 2717 8768
rect 2731 8764 2733 8768
rect 2736 8764 2738 8768
rect 2752 8764 2754 8768
rect 3061 8771 3063 8775
rect 3066 8771 3068 8775
rect 3806 8778 3808 8782
rect 3822 8778 3824 8782
rect 3838 8778 3840 8782
rect 3861 8778 3863 8782
rect 3866 8778 3868 8782
rect 3892 8778 3894 8782
rect 3913 8778 3915 8782
rect 3933 8778 3935 8782
rect 3938 8778 3940 8782
rect 3956 8778 3958 8782
rect 4040 8778 4042 8782
rect 4058 8778 4060 8782
rect 4083 8778 4085 8782
rect 4099 8778 4101 8782
rect 4122 8778 4124 8782
rect 4127 8778 4129 8782
rect 4153 8778 4155 8782
rect 4174 8778 4176 8782
rect 4194 8778 4196 8782
rect 4199 8778 4201 8782
rect 4217 8778 4219 8782
rect 3317 8764 3319 8768
rect 3322 8764 3324 8768
rect 3338 8764 3340 8768
rect 3354 8764 3356 8768
rect 3359 8764 3361 8768
rect 3380 8764 3382 8768
rect 3396 8764 3398 8768
rect 3412 8764 3414 8768
rect 3417 8764 3419 8768
rect 3433 8764 3435 8768
rect 3449 8764 3451 8768
rect 3454 8764 3456 8768
rect 3470 8764 3472 8768
rect 3486 8764 3488 8768
rect 3491 8764 3493 8768
rect 3512 8764 3514 8768
rect 3528 8764 3530 8768
rect 3544 8764 3546 8768
rect 3549 8764 3551 8768
rect 3565 8764 3567 8768
rect 3581 8764 3583 8768
rect 3586 8764 3588 8768
rect 3602 8764 3604 8768
rect 3618 8764 3620 8768
rect 3623 8764 3625 8768
rect 3644 8764 3646 8768
rect 3660 8764 3662 8768
rect 3676 8764 3678 8768
rect 3681 8764 3683 8768
rect 3697 8764 3699 8768
rect 4006 8771 4008 8775
rect 4011 8771 4013 8775
rect 2487 8720 2489 8724
rect 2511 8720 2513 8724
rect 3284 8722 3288 8724
rect 3432 8720 3434 8724
rect 3456 8720 3458 8724
rect 4229 8722 4233 8724
rect 2507 8707 2509 8711
rect 3452 8707 3454 8711
rect 2498 8693 2502 8695
rect 3443 8693 3447 8695
rect 2487 8684 2489 8688
rect 2511 8684 2513 8688
rect 3432 8684 3434 8688
rect 3456 8684 3458 8688
rect 3155 8652 3157 8656
rect 3160 8652 3162 8656
rect 3176 8652 3178 8656
rect 3192 8652 3194 8656
rect 3197 8652 3199 8656
rect 3218 8652 3220 8656
rect 3234 8652 3236 8656
rect 3250 8652 3252 8656
rect 3255 8652 3257 8656
rect 3271 8652 3273 8656
rect 4100 8652 4102 8656
rect 4105 8652 4107 8656
rect 4121 8652 4123 8656
rect 4137 8652 4139 8656
rect 4142 8652 4144 8656
rect 4163 8652 4165 8656
rect 4179 8652 4181 8656
rect 4195 8652 4197 8656
rect 4200 8652 4202 8656
rect 4216 8652 4218 8656
rect 2372 8622 2374 8626
rect 2377 8622 2379 8626
rect 2393 8622 2395 8626
rect 2409 8622 2411 8626
rect 2414 8622 2416 8626
rect 2435 8622 2437 8626
rect 2451 8622 2453 8626
rect 2467 8622 2469 8626
rect 2472 8622 2474 8626
rect 2488 8622 2490 8626
rect 2504 8622 2506 8626
rect 2509 8622 2511 8626
rect 2525 8622 2527 8626
rect 2541 8622 2543 8626
rect 2546 8622 2548 8626
rect 2567 8622 2569 8626
rect 2583 8622 2585 8626
rect 2599 8622 2601 8626
rect 2604 8622 2606 8626
rect 2620 8622 2622 8626
rect 2636 8622 2638 8626
rect 2641 8622 2643 8626
rect 2657 8622 2659 8626
rect 2673 8622 2675 8626
rect 2678 8622 2680 8626
rect 2699 8622 2701 8626
rect 2715 8622 2717 8626
rect 2731 8622 2733 8626
rect 2736 8622 2738 8626
rect 2752 8622 2754 8626
rect 3317 8622 3319 8626
rect 3322 8622 3324 8626
rect 3338 8622 3340 8626
rect 3354 8622 3356 8626
rect 3359 8622 3361 8626
rect 3380 8622 3382 8626
rect 3396 8622 3398 8626
rect 3412 8622 3414 8626
rect 3417 8622 3419 8626
rect 3433 8622 3435 8626
rect 3449 8622 3451 8626
rect 3454 8622 3456 8626
rect 3470 8622 3472 8626
rect 3486 8622 3488 8626
rect 3491 8622 3493 8626
rect 3512 8622 3514 8626
rect 3528 8622 3530 8626
rect 3544 8622 3546 8626
rect 3549 8622 3551 8626
rect 3565 8622 3567 8626
rect 3581 8622 3583 8626
rect 3586 8622 3588 8626
rect 3602 8622 3604 8626
rect 3618 8622 3620 8626
rect 3623 8622 3625 8626
rect 3644 8622 3646 8626
rect 3660 8622 3662 8626
rect 3676 8622 3678 8626
rect 3681 8622 3683 8626
rect 3697 8622 3699 8626
rect 3296 8576 3300 8578
rect 4241 8576 4245 8578
rect 3155 8566 3157 8570
rect 3160 8566 3162 8570
rect 3176 8566 3178 8570
rect 3192 8566 3194 8570
rect 3197 8566 3199 8570
rect 3218 8566 3220 8570
rect 3234 8566 3236 8570
rect 3250 8566 3252 8570
rect 3255 8566 3257 8570
rect 3271 8566 3273 8570
rect 4100 8566 4102 8570
rect 4105 8566 4107 8570
rect 4121 8566 4123 8570
rect 4137 8566 4139 8570
rect 4142 8566 4144 8570
rect 4163 8566 4165 8570
rect 4179 8566 4181 8570
rect 4195 8566 4197 8570
rect 4200 8566 4202 8570
rect 4216 8566 4218 8570
rect 2372 8536 2374 8540
rect 2377 8536 2379 8540
rect 2393 8536 2395 8540
rect 2409 8536 2411 8540
rect 2414 8536 2416 8540
rect 2435 8536 2437 8540
rect 2451 8536 2453 8540
rect 2467 8536 2469 8540
rect 2472 8536 2474 8540
rect 2488 8536 2490 8540
rect 2504 8536 2506 8540
rect 2509 8536 2511 8540
rect 2525 8536 2527 8540
rect 2541 8536 2543 8540
rect 2546 8536 2548 8540
rect 2567 8536 2569 8540
rect 2583 8536 2585 8540
rect 2599 8536 2601 8540
rect 2604 8536 2606 8540
rect 2620 8536 2622 8540
rect 2636 8536 2638 8540
rect 2641 8536 2643 8540
rect 2657 8536 2659 8540
rect 2673 8536 2675 8540
rect 2678 8536 2680 8540
rect 2699 8536 2701 8540
rect 2715 8536 2717 8540
rect 2731 8536 2733 8540
rect 2736 8536 2738 8540
rect 2752 8536 2754 8540
rect 3317 8536 3319 8540
rect 3322 8536 3324 8540
rect 3338 8536 3340 8540
rect 3354 8536 3356 8540
rect 3359 8536 3361 8540
rect 3380 8536 3382 8540
rect 3396 8536 3398 8540
rect 3412 8536 3414 8540
rect 3417 8536 3419 8540
rect 3433 8536 3435 8540
rect 3449 8536 3451 8540
rect 3454 8536 3456 8540
rect 3470 8536 3472 8540
rect 3486 8536 3488 8540
rect 3491 8536 3493 8540
rect 3512 8536 3514 8540
rect 3528 8536 3530 8540
rect 3544 8536 3546 8540
rect 3549 8536 3551 8540
rect 3565 8536 3567 8540
rect 3581 8536 3583 8540
rect 3586 8536 3588 8540
rect 3602 8536 3604 8540
rect 3618 8536 3620 8540
rect 3623 8536 3625 8540
rect 3644 8536 3646 8540
rect 3660 8536 3662 8540
rect 3676 8536 3678 8540
rect 3681 8536 3683 8540
rect 3697 8536 3699 8540
rect 2604 8492 2606 8496
rect 2628 8492 2630 8496
rect 3549 8492 3551 8496
rect 3573 8492 3575 8496
rect 2624 8481 2626 8485
rect 3569 8481 3571 8485
rect 2615 8467 2619 8469
rect 3560 8467 3564 8469
rect 2604 8458 2606 8462
rect 2628 8458 2630 8462
rect 3549 8458 3551 8462
rect 3573 8458 3575 8462
rect 2372 8396 2374 8400
rect 2377 8396 2379 8400
rect 2393 8396 2395 8400
rect 2409 8396 2411 8400
rect 2414 8396 2416 8400
rect 2435 8396 2437 8400
rect 2451 8396 2453 8400
rect 2467 8396 2469 8400
rect 2472 8396 2474 8400
rect 2488 8396 2490 8400
rect 2504 8396 2506 8400
rect 2509 8396 2511 8400
rect 2525 8396 2527 8400
rect 2541 8396 2543 8400
rect 2546 8396 2548 8400
rect 2567 8396 2569 8400
rect 2583 8396 2585 8400
rect 2599 8396 2601 8400
rect 2604 8396 2606 8400
rect 2620 8396 2622 8400
rect 2636 8396 2638 8400
rect 2641 8396 2643 8400
rect 2657 8396 2659 8400
rect 2673 8396 2675 8400
rect 2678 8396 2680 8400
rect 2699 8396 2701 8400
rect 2715 8396 2717 8400
rect 2731 8396 2733 8400
rect 2736 8396 2738 8400
rect 2752 8396 2754 8400
rect 3317 8396 3319 8400
rect 3322 8396 3324 8400
rect 3338 8396 3340 8400
rect 3354 8396 3356 8400
rect 3359 8396 3361 8400
rect 3380 8396 3382 8400
rect 3396 8396 3398 8400
rect 3412 8396 3414 8400
rect 3417 8396 3419 8400
rect 3433 8396 3435 8400
rect 3449 8396 3451 8400
rect 3454 8396 3456 8400
rect 3470 8396 3472 8400
rect 3486 8396 3488 8400
rect 3491 8396 3493 8400
rect 3512 8396 3514 8400
rect 3528 8396 3530 8400
rect 3544 8396 3546 8400
rect 3549 8396 3551 8400
rect 3565 8396 3567 8400
rect 3581 8396 3583 8400
rect 3586 8396 3588 8400
rect 3602 8396 3604 8400
rect 3618 8396 3620 8400
rect 3623 8396 3625 8400
rect 3644 8396 3646 8400
rect 3660 8396 3662 8400
rect 3676 8396 3678 8400
rect 3681 8396 3683 8400
rect 3697 8396 3699 8400
rect 2856 8317 2858 8321
rect 2861 8317 2863 8321
rect 2877 8317 2879 8321
rect 2893 8317 2895 8321
rect 2898 8317 2900 8321
rect 2919 8317 2921 8321
rect 2935 8317 2937 8321
rect 2951 8317 2953 8321
rect 2956 8317 2958 8321
rect 2972 8317 2974 8321
rect 2988 8317 2990 8321
rect 2993 8317 2995 8321
rect 3009 8317 3011 8321
rect 3025 8317 3027 8321
rect 3030 8317 3032 8321
rect 3051 8317 3053 8321
rect 3067 8317 3069 8321
rect 3083 8317 3085 8321
rect 3088 8317 3090 8321
rect 3104 8317 3106 8321
rect 3120 8317 3122 8321
rect 3125 8317 3127 8321
rect 3141 8317 3143 8321
rect 3157 8317 3159 8321
rect 3162 8317 3164 8321
rect 3183 8317 3185 8321
rect 3199 8317 3201 8321
rect 3215 8317 3217 8321
rect 3220 8317 3222 8321
rect 3236 8317 3238 8321
rect 3252 8317 3254 8321
rect 3257 8317 3259 8321
rect 3273 8317 3275 8321
rect 3289 8317 3291 8321
rect 3294 8317 3296 8321
rect 3315 8317 3317 8321
rect 3331 8317 3333 8321
rect 3347 8317 3349 8321
rect 3352 8317 3354 8321
rect 3368 8317 3370 8321
rect 3801 8317 3803 8321
rect 3806 8317 3808 8321
rect 3822 8317 3824 8321
rect 3838 8317 3840 8321
rect 3843 8317 3845 8321
rect 3864 8317 3866 8321
rect 3880 8317 3882 8321
rect 3896 8317 3898 8321
rect 3901 8317 3903 8321
rect 3917 8317 3919 8321
rect 3933 8317 3935 8321
rect 3938 8317 3940 8321
rect 3954 8317 3956 8321
rect 3970 8317 3972 8321
rect 3975 8317 3977 8321
rect 3996 8317 3998 8321
rect 4012 8317 4014 8321
rect 4028 8317 4030 8321
rect 4033 8317 4035 8321
rect 4049 8317 4051 8321
rect 4065 8317 4067 8321
rect 4070 8317 4072 8321
rect 4086 8317 4088 8321
rect 4102 8317 4104 8321
rect 4107 8317 4109 8321
rect 4128 8317 4130 8321
rect 4144 8317 4146 8321
rect 4160 8317 4162 8321
rect 4165 8317 4167 8321
rect 4181 8317 4183 8321
rect 4197 8317 4199 8321
rect 4202 8317 4204 8321
rect 4218 8317 4220 8321
rect 4234 8317 4236 8321
rect 4239 8317 4241 8321
rect 4260 8317 4262 8321
rect 4276 8317 4278 8321
rect 4292 8317 4294 8321
rect 4297 8317 4299 8321
rect 4313 8317 4315 8321
rect 2504 8284 2506 8288
rect 2509 8284 2511 8288
rect 2525 8284 2527 8288
rect 2541 8284 2543 8288
rect 2546 8284 2548 8288
rect 2567 8284 2569 8288
rect 2583 8284 2585 8288
rect 2599 8284 2601 8288
rect 2604 8284 2606 8288
rect 2620 8284 2622 8288
rect 3449 8284 3451 8288
rect 3454 8284 3456 8288
rect 3470 8284 3472 8288
rect 3486 8284 3488 8288
rect 3491 8284 3493 8288
rect 3512 8284 3514 8288
rect 3528 8284 3530 8288
rect 3544 8284 3546 8288
rect 3549 8284 3551 8288
rect 3565 8284 3567 8288
rect 2628 8247 2630 8251
rect 3035 8251 3037 8255
rect 3061 8247 3063 8251
rect 3066 8247 3068 8251
rect 3116 8251 3118 8255
rect 3142 8247 3144 8251
rect 3147 8247 3149 8251
rect 3089 8243 3091 8247
rect 2511 8238 2513 8242
rect 2861 8238 2863 8242
rect 2877 8238 2879 8242
rect 2893 8238 2895 8242
rect 2916 8238 2918 8242
rect 2921 8238 2923 8242
rect 2947 8238 2949 8242
rect 2968 8238 2970 8242
rect 2988 8238 2990 8242
rect 2993 8238 2995 8242
rect 3011 8238 3013 8242
rect 3170 8243 3172 8247
rect 3573 8247 3575 8251
rect 3980 8251 3982 8255
rect 4006 8247 4008 8251
rect 4011 8247 4013 8251
rect 4061 8251 4063 8255
rect 4087 8247 4089 8251
rect 4092 8247 4094 8251
rect 4034 8243 4036 8247
rect 3456 8238 3458 8242
rect 3806 8238 3808 8242
rect 3822 8238 3824 8242
rect 3838 8238 3840 8242
rect 3861 8238 3863 8242
rect 3866 8238 3868 8242
rect 3892 8238 3894 8242
rect 3913 8238 3915 8242
rect 3933 8238 3935 8242
rect 3938 8238 3940 8242
rect 3956 8238 3958 8242
rect 4115 8243 4117 8247
rect 2861 8192 2863 8196
rect 2877 8192 2879 8196
rect 2893 8192 2895 8196
rect 2916 8192 2918 8196
rect 2921 8192 2923 8196
rect 2947 8192 2949 8196
rect 2968 8192 2970 8196
rect 2988 8192 2990 8196
rect 2993 8192 2995 8196
rect 3011 8192 3013 8196
rect 2495 8182 2497 8186
rect 2511 8182 2513 8186
rect 2516 8182 2518 8186
rect 2532 8182 2534 8186
rect 2548 8182 2550 8186
rect 2569 8182 2571 8186
rect 2574 8182 2576 8186
rect 2590 8182 2592 8186
rect 2606 8182 2608 8186
rect 2611 8182 2613 8186
rect 3061 8191 3063 8195
rect 3066 8191 3068 8195
rect 3142 8191 3144 8195
rect 3147 8191 3149 8195
rect 3806 8192 3808 8196
rect 3822 8192 3824 8196
rect 3838 8192 3840 8196
rect 3861 8192 3863 8196
rect 3866 8192 3868 8196
rect 3892 8192 3894 8196
rect 3913 8192 3915 8196
rect 3933 8192 3935 8196
rect 3938 8192 3940 8196
rect 3956 8192 3958 8196
rect 3440 8182 3442 8186
rect 3456 8182 3458 8186
rect 3461 8182 3463 8186
rect 3477 8182 3479 8186
rect 3493 8182 3495 8186
rect 3514 8182 3516 8186
rect 3519 8182 3521 8186
rect 3535 8182 3537 8186
rect 3551 8182 3553 8186
rect 3556 8182 3558 8186
rect 4006 8191 4008 8195
rect 4011 8191 4013 8195
rect 4087 8191 4089 8195
rect 4092 8191 4094 8195
rect 3061 8115 3063 8119
rect 3066 8115 3068 8119
rect 3140 8119 3142 8123
rect 3166 8115 3168 8119
rect 3171 8115 3173 8119
rect 3089 8111 3091 8115
rect 2861 8106 2863 8110
rect 2877 8106 2879 8110
rect 2893 8106 2895 8110
rect 2916 8106 2918 8110
rect 2921 8106 2923 8110
rect 2947 8106 2949 8110
rect 2968 8106 2970 8110
rect 2988 8106 2990 8110
rect 2993 8106 2995 8110
rect 3011 8106 3013 8110
rect 3194 8111 3196 8115
rect 4006 8115 4008 8119
rect 4011 8115 4013 8119
rect 4085 8119 4087 8123
rect 4111 8115 4113 8119
rect 4116 8115 4118 8119
rect 4034 8111 4036 8115
rect 3806 8106 3808 8110
rect 3822 8106 3824 8110
rect 3838 8106 3840 8110
rect 3861 8106 3863 8110
rect 3866 8106 3868 8110
rect 3892 8106 3894 8110
rect 3913 8106 3915 8110
rect 3933 8106 3935 8110
rect 3938 8106 3940 8110
rect 3956 8106 3958 8110
rect 4139 8111 4141 8115
rect 2861 8060 2863 8064
rect 2877 8060 2879 8064
rect 2893 8060 2895 8064
rect 2916 8060 2918 8064
rect 2921 8060 2923 8064
rect 2947 8060 2949 8064
rect 2968 8060 2970 8064
rect 2988 8060 2990 8064
rect 2993 8060 2995 8064
rect 3011 8060 3013 8064
rect 3061 8060 3063 8064
rect 3066 8060 3068 8064
rect 3166 8060 3168 8064
rect 3171 8060 3173 8064
rect 3806 8060 3808 8064
rect 3822 8060 3824 8064
rect 3838 8060 3840 8064
rect 3861 8060 3863 8064
rect 3866 8060 3868 8064
rect 3892 8060 3894 8064
rect 3913 8060 3915 8064
rect 3933 8060 3935 8064
rect 3938 8060 3940 8064
rect 3956 8060 3958 8064
rect 4006 8060 4008 8064
rect 4011 8060 4013 8064
rect 4111 8060 4113 8064
rect 4116 8060 4118 8064
rect 3061 7983 3063 7987
rect 3066 7983 3068 7987
rect 3116 7987 3118 7991
rect 3142 7983 3144 7987
rect 3147 7983 3149 7987
rect 3206 7987 3208 7991
rect 3232 7983 3234 7987
rect 3237 7983 3239 7987
rect 3089 7979 3091 7983
rect 2861 7974 2863 7978
rect 2877 7974 2879 7978
rect 2893 7974 2895 7978
rect 2916 7974 2918 7978
rect 2921 7974 2923 7978
rect 2947 7974 2949 7978
rect 2968 7974 2970 7978
rect 2988 7974 2990 7978
rect 2993 7974 2995 7978
rect 3011 7974 3013 7978
rect 3170 7979 3172 7983
rect 3260 7979 3262 7983
rect 4006 7983 4008 7987
rect 4011 7983 4013 7987
rect 4061 7987 4063 7991
rect 4087 7983 4089 7987
rect 4092 7983 4094 7987
rect 4151 7987 4153 7991
rect 4177 7983 4179 7987
rect 4182 7983 4184 7987
rect 4034 7979 4036 7983
rect 3806 7974 3808 7978
rect 3822 7974 3824 7978
rect 3838 7974 3840 7978
rect 3861 7974 3863 7978
rect 3866 7974 3868 7978
rect 3892 7974 3894 7978
rect 3913 7974 3915 7978
rect 3933 7974 3935 7978
rect 3938 7974 3940 7978
rect 3956 7974 3958 7978
rect 4115 7979 4117 7983
rect 4205 7979 4207 7983
rect 2861 7928 2863 7932
rect 2877 7928 2879 7932
rect 2893 7928 2895 7932
rect 2916 7928 2918 7932
rect 2921 7928 2923 7932
rect 2947 7928 2949 7932
rect 2968 7928 2970 7932
rect 2988 7928 2990 7932
rect 2993 7928 2995 7932
rect 3011 7928 3013 7932
rect 3061 7925 3063 7929
rect 3066 7925 3068 7929
rect 3142 7925 3144 7929
rect 3147 7925 3149 7929
rect 3232 7925 3234 7929
rect 3237 7925 3239 7929
rect 3806 7928 3808 7932
rect 3822 7928 3824 7932
rect 3838 7928 3840 7932
rect 3861 7928 3863 7932
rect 3866 7928 3868 7932
rect 3892 7928 3894 7932
rect 3913 7928 3915 7932
rect 3933 7928 3935 7932
rect 3938 7928 3940 7932
rect 3956 7928 3958 7932
rect 4006 7925 4008 7929
rect 4011 7925 4013 7929
rect 4087 7925 4089 7929
rect 4092 7925 4094 7929
rect 4177 7925 4179 7929
rect 4182 7925 4184 7929
rect 3061 7851 3063 7855
rect 3066 7851 3068 7855
rect 3089 7847 3091 7851
rect 2861 7842 2863 7846
rect 2877 7842 2879 7846
rect 2893 7842 2895 7846
rect 2916 7842 2918 7846
rect 2921 7842 2923 7846
rect 2947 7842 2949 7846
rect 2968 7842 2970 7846
rect 2988 7842 2990 7846
rect 2993 7842 2995 7846
rect 3011 7842 3013 7846
rect 4006 7851 4008 7855
rect 4011 7851 4013 7855
rect 4034 7847 4036 7851
rect 3806 7842 3808 7846
rect 3822 7842 3824 7846
rect 3838 7842 3840 7846
rect 3861 7842 3863 7846
rect 3866 7842 3868 7846
rect 3892 7842 3894 7846
rect 3913 7842 3915 7846
rect 3933 7842 3935 7846
rect 3938 7842 3940 7846
rect 3956 7842 3958 7846
rect 2861 7796 2863 7800
rect 2877 7796 2879 7800
rect 2893 7796 2895 7800
rect 2916 7796 2918 7800
rect 2921 7796 2923 7800
rect 2947 7796 2949 7800
rect 2968 7796 2970 7800
rect 2988 7796 2990 7800
rect 2993 7796 2995 7800
rect 3011 7796 3013 7800
rect 3095 7796 3097 7800
rect 3113 7796 3115 7800
rect 3138 7796 3140 7800
rect 3154 7796 3156 7800
rect 3177 7796 3179 7800
rect 3182 7796 3184 7800
rect 3208 7796 3210 7800
rect 3229 7796 3231 7800
rect 3249 7796 3251 7800
rect 3254 7796 3256 7800
rect 3272 7796 3274 7800
rect 2372 7782 2374 7786
rect 2377 7782 2379 7786
rect 2393 7782 2395 7786
rect 2409 7782 2411 7786
rect 2414 7782 2416 7786
rect 2435 7782 2437 7786
rect 2451 7782 2453 7786
rect 2467 7782 2469 7786
rect 2472 7782 2474 7786
rect 2488 7782 2490 7786
rect 2504 7782 2506 7786
rect 2509 7782 2511 7786
rect 2525 7782 2527 7786
rect 2541 7782 2543 7786
rect 2546 7782 2548 7786
rect 2567 7782 2569 7786
rect 2583 7782 2585 7786
rect 2599 7782 2601 7786
rect 2604 7782 2606 7786
rect 2620 7782 2622 7786
rect 2636 7782 2638 7786
rect 2641 7782 2643 7786
rect 2657 7782 2659 7786
rect 2673 7782 2675 7786
rect 2678 7782 2680 7786
rect 2699 7782 2701 7786
rect 2715 7782 2717 7786
rect 2731 7782 2733 7786
rect 2736 7782 2738 7786
rect 2752 7782 2754 7786
rect 3061 7789 3063 7793
rect 3066 7789 3068 7793
rect 3806 7796 3808 7800
rect 3822 7796 3824 7800
rect 3838 7796 3840 7800
rect 3861 7796 3863 7800
rect 3866 7796 3868 7800
rect 3892 7796 3894 7800
rect 3913 7796 3915 7800
rect 3933 7796 3935 7800
rect 3938 7796 3940 7800
rect 3956 7796 3958 7800
rect 4040 7796 4042 7800
rect 4058 7796 4060 7800
rect 4083 7796 4085 7800
rect 4099 7796 4101 7800
rect 4122 7796 4124 7800
rect 4127 7796 4129 7800
rect 4153 7796 4155 7800
rect 4174 7796 4176 7800
rect 4194 7796 4196 7800
rect 4199 7796 4201 7800
rect 4217 7796 4219 7800
rect 3317 7782 3319 7786
rect 3322 7782 3324 7786
rect 3338 7782 3340 7786
rect 3354 7782 3356 7786
rect 3359 7782 3361 7786
rect 3380 7782 3382 7786
rect 3396 7782 3398 7786
rect 3412 7782 3414 7786
rect 3417 7782 3419 7786
rect 3433 7782 3435 7786
rect 3449 7782 3451 7786
rect 3454 7782 3456 7786
rect 3470 7782 3472 7786
rect 3486 7782 3488 7786
rect 3491 7782 3493 7786
rect 3512 7782 3514 7786
rect 3528 7782 3530 7786
rect 3544 7782 3546 7786
rect 3549 7782 3551 7786
rect 3565 7782 3567 7786
rect 3581 7782 3583 7786
rect 3586 7782 3588 7786
rect 3602 7782 3604 7786
rect 3618 7782 3620 7786
rect 3623 7782 3625 7786
rect 3644 7782 3646 7786
rect 3660 7782 3662 7786
rect 3676 7782 3678 7786
rect 3681 7782 3683 7786
rect 3697 7782 3699 7786
rect 4006 7789 4008 7793
rect 4011 7789 4013 7793
rect 2487 7738 2489 7742
rect 2511 7738 2513 7742
rect 3284 7740 3288 7742
rect 3432 7738 3434 7742
rect 3456 7738 3458 7742
rect 4229 7740 4233 7742
rect 2507 7725 2509 7729
rect 3452 7725 3454 7729
rect 2498 7711 2502 7713
rect 3443 7711 3447 7713
rect 2487 7702 2489 7706
rect 2511 7702 2513 7706
rect 3432 7702 3434 7706
rect 3456 7702 3458 7706
rect 3155 7670 3157 7674
rect 3160 7670 3162 7674
rect 3176 7670 3178 7674
rect 3192 7670 3194 7674
rect 3197 7670 3199 7674
rect 3218 7670 3220 7674
rect 3234 7670 3236 7674
rect 3250 7670 3252 7674
rect 3255 7670 3257 7674
rect 3271 7670 3273 7674
rect 4100 7670 4102 7674
rect 4105 7670 4107 7674
rect 4121 7670 4123 7674
rect 4137 7670 4139 7674
rect 4142 7670 4144 7674
rect 4163 7670 4165 7674
rect 4179 7670 4181 7674
rect 4195 7670 4197 7674
rect 4200 7670 4202 7674
rect 4216 7670 4218 7674
rect 2372 7640 2374 7644
rect 2377 7640 2379 7644
rect 2393 7640 2395 7644
rect 2409 7640 2411 7644
rect 2414 7640 2416 7644
rect 2435 7640 2437 7644
rect 2451 7640 2453 7644
rect 2467 7640 2469 7644
rect 2472 7640 2474 7644
rect 2488 7640 2490 7644
rect 2504 7640 2506 7644
rect 2509 7640 2511 7644
rect 2525 7640 2527 7644
rect 2541 7640 2543 7644
rect 2546 7640 2548 7644
rect 2567 7640 2569 7644
rect 2583 7640 2585 7644
rect 2599 7640 2601 7644
rect 2604 7640 2606 7644
rect 2620 7640 2622 7644
rect 2636 7640 2638 7644
rect 2641 7640 2643 7644
rect 2657 7640 2659 7644
rect 2673 7640 2675 7644
rect 2678 7640 2680 7644
rect 2699 7640 2701 7644
rect 2715 7640 2717 7644
rect 2731 7640 2733 7644
rect 2736 7640 2738 7644
rect 2752 7640 2754 7644
rect 3317 7640 3319 7644
rect 3322 7640 3324 7644
rect 3338 7640 3340 7644
rect 3354 7640 3356 7644
rect 3359 7640 3361 7644
rect 3380 7640 3382 7644
rect 3396 7640 3398 7644
rect 3412 7640 3414 7644
rect 3417 7640 3419 7644
rect 3433 7640 3435 7644
rect 3449 7640 3451 7644
rect 3454 7640 3456 7644
rect 3470 7640 3472 7644
rect 3486 7640 3488 7644
rect 3491 7640 3493 7644
rect 3512 7640 3514 7644
rect 3528 7640 3530 7644
rect 3544 7640 3546 7644
rect 3549 7640 3551 7644
rect 3565 7640 3567 7644
rect 3581 7640 3583 7644
rect 3586 7640 3588 7644
rect 3602 7640 3604 7644
rect 3618 7640 3620 7644
rect 3623 7640 3625 7644
rect 3644 7640 3646 7644
rect 3660 7640 3662 7644
rect 3676 7640 3678 7644
rect 3681 7640 3683 7644
rect 3697 7640 3699 7644
rect 3296 7594 3300 7596
rect 4241 7594 4245 7596
rect 3155 7584 3157 7588
rect 3160 7584 3162 7588
rect 3176 7584 3178 7588
rect 3192 7584 3194 7588
rect 3197 7584 3199 7588
rect 3218 7584 3220 7588
rect 3234 7584 3236 7588
rect 3250 7584 3252 7588
rect 3255 7584 3257 7588
rect 3271 7584 3273 7588
rect 4100 7584 4102 7588
rect 4105 7584 4107 7588
rect 4121 7584 4123 7588
rect 4137 7584 4139 7588
rect 4142 7584 4144 7588
rect 4163 7584 4165 7588
rect 4179 7584 4181 7588
rect 4195 7584 4197 7588
rect 4200 7584 4202 7588
rect 4216 7584 4218 7588
rect 2372 7554 2374 7558
rect 2377 7554 2379 7558
rect 2393 7554 2395 7558
rect 2409 7554 2411 7558
rect 2414 7554 2416 7558
rect 2435 7554 2437 7558
rect 2451 7554 2453 7558
rect 2467 7554 2469 7558
rect 2472 7554 2474 7558
rect 2488 7554 2490 7558
rect 2504 7554 2506 7558
rect 2509 7554 2511 7558
rect 2525 7554 2527 7558
rect 2541 7554 2543 7558
rect 2546 7554 2548 7558
rect 2567 7554 2569 7558
rect 2583 7554 2585 7558
rect 2599 7554 2601 7558
rect 2604 7554 2606 7558
rect 2620 7554 2622 7558
rect 2636 7554 2638 7558
rect 2641 7554 2643 7558
rect 2657 7554 2659 7558
rect 2673 7554 2675 7558
rect 2678 7554 2680 7558
rect 2699 7554 2701 7558
rect 2715 7554 2717 7558
rect 2731 7554 2733 7558
rect 2736 7554 2738 7558
rect 2752 7554 2754 7558
rect 3317 7554 3319 7558
rect 3322 7554 3324 7558
rect 3338 7554 3340 7558
rect 3354 7554 3356 7558
rect 3359 7554 3361 7558
rect 3380 7554 3382 7558
rect 3396 7554 3398 7558
rect 3412 7554 3414 7558
rect 3417 7554 3419 7558
rect 3433 7554 3435 7558
rect 3449 7554 3451 7558
rect 3454 7554 3456 7558
rect 3470 7554 3472 7558
rect 3486 7554 3488 7558
rect 3491 7554 3493 7558
rect 3512 7554 3514 7558
rect 3528 7554 3530 7558
rect 3544 7554 3546 7558
rect 3549 7554 3551 7558
rect 3565 7554 3567 7558
rect 3581 7554 3583 7558
rect 3586 7554 3588 7558
rect 3602 7554 3604 7558
rect 3618 7554 3620 7558
rect 3623 7554 3625 7558
rect 3644 7554 3646 7558
rect 3660 7554 3662 7558
rect 3676 7554 3678 7558
rect 3681 7554 3683 7558
rect 3697 7554 3699 7558
rect 2604 7510 2606 7514
rect 2628 7510 2630 7514
rect 3549 7510 3551 7514
rect 3573 7510 3575 7514
rect 2624 7499 2626 7503
rect 3569 7499 3571 7503
rect 2615 7485 2619 7487
rect 3560 7485 3564 7487
rect 2604 7476 2606 7480
rect 2628 7476 2630 7480
rect 3549 7476 3551 7480
rect 3573 7476 3575 7480
rect 3836 7473 3844 7475
rect 2372 7414 2374 7418
rect 2377 7414 2379 7418
rect 2393 7414 2395 7418
rect 2409 7414 2411 7418
rect 2414 7414 2416 7418
rect 2435 7414 2437 7418
rect 2451 7414 2453 7418
rect 2467 7414 2469 7418
rect 2472 7414 2474 7418
rect 2488 7414 2490 7418
rect 2504 7414 2506 7418
rect 2509 7414 2511 7418
rect 2525 7414 2527 7418
rect 2541 7414 2543 7418
rect 2546 7414 2548 7418
rect 2567 7414 2569 7418
rect 2583 7414 2585 7418
rect 2599 7414 2601 7418
rect 2604 7414 2606 7418
rect 2620 7414 2622 7418
rect 2636 7414 2638 7418
rect 2641 7414 2643 7418
rect 2657 7414 2659 7418
rect 2673 7414 2675 7418
rect 2678 7414 2680 7418
rect 2699 7414 2701 7418
rect 2715 7414 2717 7418
rect 2731 7414 2733 7418
rect 2736 7414 2738 7418
rect 2752 7414 2754 7418
rect 3317 7414 3319 7418
rect 3322 7414 3324 7418
rect 3338 7414 3340 7418
rect 3354 7414 3356 7418
rect 3359 7414 3361 7418
rect 3380 7414 3382 7418
rect 3396 7414 3398 7418
rect 3412 7414 3414 7418
rect 3417 7414 3419 7418
rect 3433 7414 3435 7418
rect 3449 7414 3451 7418
rect 3454 7414 3456 7418
rect 3470 7414 3472 7418
rect 3486 7414 3488 7418
rect 3491 7414 3493 7418
rect 3512 7414 3514 7418
rect 3528 7414 3530 7418
rect 3544 7414 3546 7418
rect 3549 7414 3551 7418
rect 3565 7414 3567 7418
rect 3581 7414 3583 7418
rect 3586 7414 3588 7418
rect 3602 7414 3604 7418
rect 3618 7414 3620 7418
rect 3623 7414 3625 7418
rect 3644 7414 3646 7418
rect 3660 7414 3662 7418
rect 3676 7414 3678 7418
rect 3681 7414 3683 7418
rect 3697 7414 3699 7418
rect 1473 6896 1475 6900
rect 1489 6896 1491 6900
rect 1494 6896 1496 6900
rect 1510 6896 1512 6900
rect 1526 6896 1528 6900
rect 1547 6896 1549 6900
rect 1552 6896 1554 6900
rect 1568 6896 1570 6900
rect 1584 6896 1586 6900
rect 1589 6896 1591 6900
rect 1605 6896 1607 6900
rect 1621 6896 1623 6900
rect 1626 6896 1628 6900
rect 1642 6896 1644 6900
rect 1658 6896 1660 6900
rect 1679 6896 1681 6900
rect 1684 6896 1686 6900
rect 1700 6896 1702 6900
rect 1716 6896 1718 6900
rect 1721 6896 1723 6900
rect 1737 6896 1739 6900
rect 1753 6896 1755 6900
rect 1758 6896 1760 6900
rect 1774 6896 1776 6900
rect 1790 6896 1792 6900
rect 1811 6896 1813 6900
rect 1816 6896 1818 6900
rect 1832 6896 1834 6900
rect 1848 6896 1850 6900
rect 1853 6896 1855 6900
rect 2418 6896 2420 6900
rect 2434 6896 2436 6900
rect 2439 6896 2441 6900
rect 2455 6896 2457 6900
rect 2471 6896 2473 6900
rect 2492 6896 2494 6900
rect 2497 6896 2499 6900
rect 2513 6896 2515 6900
rect 2529 6896 2531 6900
rect 2534 6896 2536 6900
rect 2550 6896 2552 6900
rect 2566 6896 2568 6900
rect 2571 6896 2573 6900
rect 2587 6896 2589 6900
rect 2603 6896 2605 6900
rect 2624 6896 2626 6900
rect 2629 6896 2631 6900
rect 2645 6896 2647 6900
rect 2661 6896 2663 6900
rect 2666 6896 2668 6900
rect 2682 6896 2684 6900
rect 2698 6896 2700 6900
rect 2703 6896 2705 6900
rect 2719 6896 2721 6900
rect 2735 6896 2737 6900
rect 2756 6896 2758 6900
rect 2761 6896 2763 6900
rect 2777 6896 2779 6900
rect 2793 6896 2795 6900
rect 2798 6896 2800 6900
rect 1597 6834 1599 6838
rect 1621 6834 1623 6838
rect 2542 6834 2544 6838
rect 2566 6834 2568 6838
rect 1608 6827 1612 6829
rect 2553 6827 2557 6829
rect 1601 6811 1603 6815
rect 2546 6811 2548 6815
rect 1597 6800 1599 6804
rect 1621 6800 1623 6804
rect 2542 6800 2544 6804
rect 2566 6800 2568 6804
rect 1473 6756 1475 6760
rect 1489 6756 1491 6760
rect 1494 6756 1496 6760
rect 1510 6756 1512 6760
rect 1526 6756 1528 6760
rect 1547 6756 1549 6760
rect 1552 6756 1554 6760
rect 1568 6756 1570 6760
rect 1584 6756 1586 6760
rect 1589 6756 1591 6760
rect 1605 6756 1607 6760
rect 1621 6756 1623 6760
rect 1626 6756 1628 6760
rect 1642 6756 1644 6760
rect 1658 6756 1660 6760
rect 1679 6756 1681 6760
rect 1684 6756 1686 6760
rect 1700 6756 1702 6760
rect 1716 6756 1718 6760
rect 1721 6756 1723 6760
rect 1737 6756 1739 6760
rect 1753 6756 1755 6760
rect 1758 6756 1760 6760
rect 1774 6756 1776 6760
rect 1790 6756 1792 6760
rect 1811 6756 1813 6760
rect 1816 6756 1818 6760
rect 1832 6756 1834 6760
rect 1848 6756 1850 6760
rect 1853 6756 1855 6760
rect 2418 6756 2420 6760
rect 2434 6756 2436 6760
rect 2439 6756 2441 6760
rect 2455 6756 2457 6760
rect 2471 6756 2473 6760
rect 2492 6756 2494 6760
rect 2497 6756 2499 6760
rect 2513 6756 2515 6760
rect 2529 6756 2531 6760
rect 2534 6756 2536 6760
rect 2550 6756 2552 6760
rect 2566 6756 2568 6760
rect 2571 6756 2573 6760
rect 2587 6756 2589 6760
rect 2603 6756 2605 6760
rect 2624 6756 2626 6760
rect 2629 6756 2631 6760
rect 2645 6756 2647 6760
rect 2661 6756 2663 6760
rect 2666 6756 2668 6760
rect 2682 6756 2684 6760
rect 2698 6756 2700 6760
rect 2703 6756 2705 6760
rect 2719 6756 2721 6760
rect 2735 6756 2737 6760
rect 2756 6756 2758 6760
rect 2761 6756 2763 6760
rect 2777 6756 2779 6760
rect 2793 6756 2795 6760
rect 2798 6756 2800 6760
rect 954 6726 956 6730
rect 970 6726 972 6730
rect 975 6726 977 6730
rect 991 6726 993 6730
rect 1007 6726 1009 6730
rect 1028 6726 1030 6730
rect 1033 6726 1035 6730
rect 1049 6726 1051 6730
rect 1065 6726 1067 6730
rect 1070 6726 1072 6730
rect 1899 6726 1901 6730
rect 1915 6726 1917 6730
rect 1920 6726 1922 6730
rect 1936 6726 1938 6730
rect 1952 6726 1954 6730
rect 1973 6726 1975 6730
rect 1978 6726 1980 6730
rect 1994 6726 1996 6730
rect 2010 6726 2012 6730
rect 2015 6726 2017 6730
rect 927 6718 931 6720
rect 1872 6718 1876 6720
rect 1473 6670 1475 6674
rect 1489 6670 1491 6674
rect 1494 6670 1496 6674
rect 1510 6670 1512 6674
rect 1526 6670 1528 6674
rect 1547 6670 1549 6674
rect 1552 6670 1554 6674
rect 1568 6670 1570 6674
rect 1584 6670 1586 6674
rect 1589 6670 1591 6674
rect 1605 6670 1607 6674
rect 1621 6670 1623 6674
rect 1626 6670 1628 6674
rect 1642 6670 1644 6674
rect 1658 6670 1660 6674
rect 1679 6670 1681 6674
rect 1684 6670 1686 6674
rect 1700 6670 1702 6674
rect 1716 6670 1718 6674
rect 1721 6670 1723 6674
rect 1737 6670 1739 6674
rect 1753 6670 1755 6674
rect 1758 6670 1760 6674
rect 1774 6670 1776 6674
rect 1790 6670 1792 6674
rect 1811 6670 1813 6674
rect 1816 6670 1818 6674
rect 1832 6670 1834 6674
rect 1848 6670 1850 6674
rect 1853 6670 1855 6674
rect 2418 6670 2420 6674
rect 2434 6670 2436 6674
rect 2439 6670 2441 6674
rect 2455 6670 2457 6674
rect 2471 6670 2473 6674
rect 2492 6670 2494 6674
rect 2497 6670 2499 6674
rect 2513 6670 2515 6674
rect 2529 6670 2531 6674
rect 2534 6670 2536 6674
rect 2550 6670 2552 6674
rect 2566 6670 2568 6674
rect 2571 6670 2573 6674
rect 2587 6670 2589 6674
rect 2603 6670 2605 6674
rect 2624 6670 2626 6674
rect 2629 6670 2631 6674
rect 2645 6670 2647 6674
rect 2661 6670 2663 6674
rect 2666 6670 2668 6674
rect 2682 6670 2684 6674
rect 2698 6670 2700 6674
rect 2703 6670 2705 6674
rect 2719 6670 2721 6674
rect 2735 6670 2737 6674
rect 2756 6670 2758 6674
rect 2761 6670 2763 6674
rect 2777 6670 2779 6674
rect 2793 6670 2795 6674
rect 2798 6670 2800 6674
rect 954 6640 956 6644
rect 970 6640 972 6644
rect 975 6640 977 6644
rect 991 6640 993 6644
rect 1007 6640 1009 6644
rect 1028 6640 1030 6644
rect 1033 6640 1035 6644
rect 1049 6640 1051 6644
rect 1065 6640 1067 6644
rect 1070 6640 1072 6644
rect 1899 6640 1901 6644
rect 1915 6640 1917 6644
rect 1920 6640 1922 6644
rect 1936 6640 1938 6644
rect 1952 6640 1954 6644
rect 1973 6640 1975 6644
rect 1978 6640 1980 6644
rect 1994 6640 1996 6644
rect 2010 6640 2012 6644
rect 2015 6640 2017 6644
rect 1714 6608 1716 6612
rect 1738 6608 1740 6612
rect 2659 6608 2661 6612
rect 2683 6608 2685 6612
rect 1725 6601 1729 6603
rect 2670 6601 2674 6603
rect 1718 6585 1720 6589
rect 2663 6585 2665 6589
rect 939 6572 943 6574
rect 1714 6572 1716 6576
rect 1738 6572 1740 6576
rect 1884 6572 1888 6574
rect 2659 6572 2661 6576
rect 2683 6572 2685 6576
rect 1159 6521 1161 6525
rect 1164 6521 1166 6525
rect 1473 6528 1475 6532
rect 1489 6528 1491 6532
rect 1494 6528 1496 6532
rect 1510 6528 1512 6532
rect 1526 6528 1528 6532
rect 1547 6528 1549 6532
rect 1552 6528 1554 6532
rect 1568 6528 1570 6532
rect 1584 6528 1586 6532
rect 1589 6528 1591 6532
rect 1605 6528 1607 6532
rect 1621 6528 1623 6532
rect 1626 6528 1628 6532
rect 1642 6528 1644 6532
rect 1658 6528 1660 6532
rect 1679 6528 1681 6532
rect 1684 6528 1686 6532
rect 1700 6528 1702 6532
rect 1716 6528 1718 6532
rect 1721 6528 1723 6532
rect 1737 6528 1739 6532
rect 1753 6528 1755 6532
rect 1758 6528 1760 6532
rect 1774 6528 1776 6532
rect 1790 6528 1792 6532
rect 1811 6528 1813 6532
rect 1816 6528 1818 6532
rect 1832 6528 1834 6532
rect 1848 6528 1850 6532
rect 1853 6528 1855 6532
rect 953 6514 955 6518
rect 971 6514 973 6518
rect 976 6514 978 6518
rect 996 6514 998 6518
rect 1017 6514 1019 6518
rect 1043 6514 1045 6518
rect 1048 6514 1050 6518
rect 1071 6514 1073 6518
rect 1087 6514 1089 6518
rect 1112 6514 1114 6518
rect 1130 6514 1132 6518
rect 1214 6514 1216 6518
rect 1232 6514 1234 6518
rect 1237 6514 1239 6518
rect 1257 6514 1259 6518
rect 1278 6514 1280 6518
rect 1304 6514 1306 6518
rect 1309 6514 1311 6518
rect 1332 6514 1334 6518
rect 1348 6514 1350 6518
rect 1364 6514 1366 6518
rect 2104 6521 2106 6525
rect 2109 6521 2111 6525
rect 2418 6528 2420 6532
rect 2434 6528 2436 6532
rect 2439 6528 2441 6532
rect 2455 6528 2457 6532
rect 2471 6528 2473 6532
rect 2492 6528 2494 6532
rect 2497 6528 2499 6532
rect 2513 6528 2515 6532
rect 2529 6528 2531 6532
rect 2534 6528 2536 6532
rect 2550 6528 2552 6532
rect 2566 6528 2568 6532
rect 2571 6528 2573 6532
rect 2587 6528 2589 6532
rect 2603 6528 2605 6532
rect 2624 6528 2626 6532
rect 2629 6528 2631 6532
rect 2645 6528 2647 6532
rect 2661 6528 2663 6532
rect 2666 6528 2668 6532
rect 2682 6528 2684 6532
rect 2698 6528 2700 6532
rect 2703 6528 2705 6532
rect 2719 6528 2721 6532
rect 2735 6528 2737 6532
rect 2756 6528 2758 6532
rect 2761 6528 2763 6532
rect 2777 6528 2779 6532
rect 2793 6528 2795 6532
rect 2798 6528 2800 6532
rect 1898 6514 1900 6518
rect 1916 6514 1918 6518
rect 1921 6514 1923 6518
rect 1941 6514 1943 6518
rect 1962 6514 1964 6518
rect 1988 6514 1990 6518
rect 1993 6514 1995 6518
rect 2016 6514 2018 6518
rect 2032 6514 2034 6518
rect 2057 6514 2059 6518
rect 2075 6514 2077 6518
rect 2159 6514 2161 6518
rect 2177 6514 2179 6518
rect 2182 6514 2184 6518
rect 2202 6514 2204 6518
rect 2223 6514 2225 6518
rect 2249 6514 2251 6518
rect 2254 6514 2256 6518
rect 2277 6514 2279 6518
rect 2293 6514 2295 6518
rect 2309 6514 2311 6518
rect 1214 6468 1216 6472
rect 1232 6468 1234 6472
rect 1237 6468 1239 6472
rect 1257 6468 1259 6472
rect 1278 6468 1280 6472
rect 1304 6468 1306 6472
rect 1309 6468 1311 6472
rect 1332 6468 1334 6472
rect 1348 6468 1350 6472
rect 1364 6468 1366 6472
rect 1136 6463 1138 6467
rect 1159 6459 1161 6463
rect 1164 6459 1166 6463
rect 2159 6468 2161 6472
rect 2177 6468 2179 6472
rect 2182 6468 2184 6472
rect 2202 6468 2204 6472
rect 2223 6468 2225 6472
rect 2249 6468 2251 6472
rect 2254 6468 2256 6472
rect 2277 6468 2279 6472
rect 2293 6468 2295 6472
rect 2309 6468 2311 6472
rect 2081 6463 2083 6467
rect 2104 6459 2106 6463
rect 2109 6459 2111 6463
rect 988 6385 990 6389
rect 993 6385 995 6389
rect 1078 6385 1080 6389
rect 1083 6385 1085 6389
rect 1159 6385 1161 6389
rect 1164 6385 1166 6389
rect 1214 6382 1216 6386
rect 1232 6382 1234 6386
rect 1237 6382 1239 6386
rect 1257 6382 1259 6386
rect 1278 6382 1280 6386
rect 1304 6382 1306 6386
rect 1309 6382 1311 6386
rect 1332 6382 1334 6386
rect 1348 6382 1350 6386
rect 1364 6382 1366 6386
rect 1933 6385 1935 6389
rect 1938 6385 1940 6389
rect 2023 6385 2025 6389
rect 2028 6385 2030 6389
rect 2104 6385 2106 6389
rect 2109 6385 2111 6389
rect 2159 6382 2161 6386
rect 2177 6382 2179 6386
rect 2182 6382 2184 6386
rect 2202 6382 2204 6386
rect 2223 6382 2225 6386
rect 2249 6382 2251 6386
rect 2254 6382 2256 6386
rect 2277 6382 2279 6386
rect 2293 6382 2295 6386
rect 2309 6382 2311 6386
rect 965 6331 967 6335
rect 1055 6331 1057 6335
rect 1214 6336 1216 6340
rect 1232 6336 1234 6340
rect 1237 6336 1239 6340
rect 1257 6336 1259 6340
rect 1278 6336 1280 6340
rect 1304 6336 1306 6340
rect 1309 6336 1311 6340
rect 1332 6336 1334 6340
rect 1348 6336 1350 6340
rect 1364 6336 1366 6340
rect 1136 6331 1138 6335
rect 988 6327 990 6331
rect 993 6327 995 6331
rect 1019 6323 1021 6327
rect 1078 6327 1080 6331
rect 1083 6327 1085 6331
rect 1109 6323 1111 6327
rect 1159 6327 1161 6331
rect 1164 6327 1166 6331
rect 1910 6331 1912 6335
rect 2000 6331 2002 6335
rect 2159 6336 2161 6340
rect 2177 6336 2179 6340
rect 2182 6336 2184 6340
rect 2202 6336 2204 6340
rect 2223 6336 2225 6340
rect 2249 6336 2251 6340
rect 2254 6336 2256 6340
rect 2277 6336 2279 6340
rect 2293 6336 2295 6340
rect 2309 6336 2311 6340
rect 2081 6331 2083 6335
rect 1933 6327 1935 6331
rect 1938 6327 1940 6331
rect 1964 6323 1966 6327
rect 2023 6327 2025 6331
rect 2028 6327 2030 6331
rect 2054 6323 2056 6327
rect 2104 6327 2106 6331
rect 2109 6327 2111 6331
rect 1054 6250 1056 6254
rect 1059 6250 1061 6254
rect 1159 6250 1161 6254
rect 1164 6250 1166 6254
rect 1214 6250 1216 6254
rect 1232 6250 1234 6254
rect 1237 6250 1239 6254
rect 1257 6250 1259 6254
rect 1278 6250 1280 6254
rect 1304 6250 1306 6254
rect 1309 6250 1311 6254
rect 1332 6250 1334 6254
rect 1348 6250 1350 6254
rect 1364 6250 1366 6254
rect 1999 6250 2001 6254
rect 2004 6250 2006 6254
rect 2104 6250 2106 6254
rect 2109 6250 2111 6254
rect 2159 6250 2161 6254
rect 2177 6250 2179 6254
rect 2182 6250 2184 6254
rect 2202 6250 2204 6254
rect 2223 6250 2225 6254
rect 2249 6250 2251 6254
rect 2254 6250 2256 6254
rect 2277 6250 2279 6254
rect 2293 6250 2295 6254
rect 2309 6250 2311 6254
rect 1031 6199 1033 6203
rect 1214 6204 1216 6208
rect 1232 6204 1234 6208
rect 1237 6204 1239 6208
rect 1257 6204 1259 6208
rect 1278 6204 1280 6208
rect 1304 6204 1306 6208
rect 1309 6204 1311 6208
rect 1332 6204 1334 6208
rect 1348 6204 1350 6208
rect 1364 6204 1366 6208
rect 1136 6199 1138 6203
rect 1054 6195 1056 6199
rect 1059 6195 1061 6199
rect 1085 6191 1087 6195
rect 1159 6195 1161 6199
rect 1164 6195 1166 6199
rect 1976 6199 1978 6203
rect 2159 6204 2161 6208
rect 2177 6204 2179 6208
rect 2182 6204 2184 6208
rect 2202 6204 2204 6208
rect 2223 6204 2225 6208
rect 2249 6204 2251 6208
rect 2254 6204 2256 6208
rect 2277 6204 2279 6208
rect 2293 6204 2295 6208
rect 2309 6204 2311 6208
rect 2081 6199 2083 6203
rect 1999 6195 2001 6199
rect 2004 6195 2006 6199
rect 2030 6191 2032 6195
rect 2104 6195 2106 6199
rect 2109 6195 2111 6199
rect 1078 6119 1080 6123
rect 1083 6119 1085 6123
rect 1159 6119 1161 6123
rect 1164 6119 1166 6123
rect 1614 6128 1616 6132
rect 1619 6128 1621 6132
rect 1635 6128 1637 6132
rect 1651 6128 1653 6132
rect 1656 6128 1658 6132
rect 1677 6128 1679 6132
rect 1693 6128 1695 6132
rect 1709 6128 1711 6132
rect 1714 6128 1716 6132
rect 1730 6128 1732 6132
rect 1214 6118 1216 6122
rect 1232 6118 1234 6122
rect 1237 6118 1239 6122
rect 1257 6118 1259 6122
rect 1278 6118 1280 6122
rect 1304 6118 1306 6122
rect 1309 6118 1311 6122
rect 1332 6118 1334 6122
rect 1348 6118 1350 6122
rect 1364 6118 1366 6122
rect 2023 6119 2025 6123
rect 2028 6119 2030 6123
rect 2104 6119 2106 6123
rect 2109 6119 2111 6123
rect 2559 6128 2561 6132
rect 2564 6128 2566 6132
rect 2580 6128 2582 6132
rect 2596 6128 2598 6132
rect 2601 6128 2603 6132
rect 2622 6128 2624 6132
rect 2638 6128 2640 6132
rect 2654 6128 2656 6132
rect 2659 6128 2661 6132
rect 2675 6128 2677 6132
rect 2159 6118 2161 6122
rect 2177 6118 2179 6122
rect 2182 6118 2184 6122
rect 2202 6118 2204 6122
rect 2223 6118 2225 6122
rect 2249 6118 2251 6122
rect 2254 6118 2256 6122
rect 2277 6118 2279 6122
rect 2293 6118 2295 6122
rect 2309 6118 2311 6122
rect 1055 6067 1057 6071
rect 1214 6072 1216 6076
rect 1232 6072 1234 6076
rect 1237 6072 1239 6076
rect 1257 6072 1259 6076
rect 1278 6072 1280 6076
rect 1304 6072 1306 6076
rect 1309 6072 1311 6076
rect 1332 6072 1334 6076
rect 1348 6072 1350 6076
rect 1364 6072 1366 6076
rect 1714 6072 1716 6076
rect 1136 6067 1138 6071
rect 1078 6063 1080 6067
rect 1083 6063 1085 6067
rect 1109 6059 1111 6063
rect 1159 6063 1161 6067
rect 1164 6063 1166 6067
rect 1190 6059 1192 6063
rect 1597 6063 1599 6067
rect 2000 6067 2002 6071
rect 2159 6072 2161 6076
rect 2177 6072 2179 6076
rect 2182 6072 2184 6076
rect 2202 6072 2204 6076
rect 2223 6072 2225 6076
rect 2249 6072 2251 6076
rect 2254 6072 2256 6076
rect 2277 6072 2279 6076
rect 2293 6072 2295 6076
rect 2309 6072 2311 6076
rect 2659 6072 2661 6076
rect 2081 6067 2083 6071
rect 2023 6063 2025 6067
rect 2028 6063 2030 6067
rect 2054 6059 2056 6063
rect 2104 6063 2106 6067
rect 2109 6063 2111 6067
rect 2135 6059 2137 6063
rect 2542 6063 2544 6067
rect 1605 6026 1607 6030
rect 1621 6026 1623 6030
rect 1626 6026 1628 6030
rect 1642 6026 1644 6030
rect 1658 6026 1660 6030
rect 1679 6026 1681 6030
rect 1684 6026 1686 6030
rect 1700 6026 1702 6030
rect 1716 6026 1718 6030
rect 1721 6026 1723 6030
rect 2550 6026 2552 6030
rect 2566 6026 2568 6030
rect 2571 6026 2573 6030
rect 2587 6026 2589 6030
rect 2603 6026 2605 6030
rect 2624 6026 2626 6030
rect 2629 6026 2631 6030
rect 2645 6026 2647 6030
rect 2661 6026 2663 6030
rect 2666 6026 2668 6030
rect 857 5993 859 5997
rect 873 5993 875 5997
rect 878 5993 880 5997
rect 894 5993 896 5997
rect 910 5993 912 5997
rect 931 5993 933 5997
rect 936 5993 938 5997
rect 952 5993 954 5997
rect 968 5993 970 5997
rect 973 5993 975 5997
rect 989 5993 991 5997
rect 1005 5993 1007 5997
rect 1010 5993 1012 5997
rect 1026 5993 1028 5997
rect 1042 5993 1044 5997
rect 1063 5993 1065 5997
rect 1068 5993 1070 5997
rect 1084 5993 1086 5997
rect 1100 5993 1102 5997
rect 1105 5993 1107 5997
rect 1121 5993 1123 5997
rect 1137 5993 1139 5997
rect 1142 5993 1144 5997
rect 1158 5993 1160 5997
rect 1174 5993 1176 5997
rect 1195 5993 1197 5997
rect 1200 5993 1202 5997
rect 1216 5993 1218 5997
rect 1232 5993 1234 5997
rect 1237 5993 1239 5997
rect 1253 5993 1255 5997
rect 1269 5993 1271 5997
rect 1274 5993 1276 5997
rect 1290 5993 1292 5997
rect 1306 5993 1308 5997
rect 1327 5993 1329 5997
rect 1332 5993 1334 5997
rect 1348 5993 1350 5997
rect 1364 5993 1366 5997
rect 1369 5993 1371 5997
rect 1802 5993 1804 5997
rect 1818 5993 1820 5997
rect 1823 5993 1825 5997
rect 1839 5993 1841 5997
rect 1855 5993 1857 5997
rect 1876 5993 1878 5997
rect 1881 5993 1883 5997
rect 1897 5993 1899 5997
rect 1913 5993 1915 5997
rect 1918 5993 1920 5997
rect 1934 5993 1936 5997
rect 1950 5993 1952 5997
rect 1955 5993 1957 5997
rect 1971 5993 1973 5997
rect 1987 5993 1989 5997
rect 2008 5993 2010 5997
rect 2013 5993 2015 5997
rect 2029 5993 2031 5997
rect 2045 5993 2047 5997
rect 2050 5993 2052 5997
rect 2066 5993 2068 5997
rect 2082 5993 2084 5997
rect 2087 5993 2089 5997
rect 2103 5993 2105 5997
rect 2119 5993 2121 5997
rect 2140 5993 2142 5997
rect 2145 5993 2147 5997
rect 2161 5993 2163 5997
rect 2177 5993 2179 5997
rect 2182 5993 2184 5997
rect 2198 5993 2200 5997
rect 2214 5993 2216 5997
rect 2219 5993 2221 5997
rect 2235 5993 2237 5997
rect 2251 5993 2253 5997
rect 2272 5993 2274 5997
rect 2277 5993 2279 5997
rect 2293 5993 2295 5997
rect 2309 5993 2311 5997
rect 2314 5993 2316 5997
rect 1473 5914 1475 5918
rect 1489 5914 1491 5918
rect 1494 5914 1496 5918
rect 1510 5914 1512 5918
rect 1526 5914 1528 5918
rect 1547 5914 1549 5918
rect 1552 5914 1554 5918
rect 1568 5914 1570 5918
rect 1584 5914 1586 5918
rect 1589 5914 1591 5918
rect 1605 5914 1607 5918
rect 1621 5914 1623 5918
rect 1626 5914 1628 5918
rect 1642 5914 1644 5918
rect 1658 5914 1660 5918
rect 1679 5914 1681 5918
rect 1684 5914 1686 5918
rect 1700 5914 1702 5918
rect 1716 5914 1718 5918
rect 1721 5914 1723 5918
rect 1737 5914 1739 5918
rect 1753 5914 1755 5918
rect 1758 5914 1760 5918
rect 1774 5914 1776 5918
rect 1790 5914 1792 5918
rect 1811 5914 1813 5918
rect 1816 5914 1818 5918
rect 1832 5914 1834 5918
rect 1848 5914 1850 5918
rect 1853 5914 1855 5918
rect 2418 5914 2420 5918
rect 2434 5914 2436 5918
rect 2439 5914 2441 5918
rect 2455 5914 2457 5918
rect 2471 5914 2473 5918
rect 2492 5914 2494 5918
rect 2497 5914 2499 5918
rect 2513 5914 2515 5918
rect 2529 5914 2531 5918
rect 2534 5914 2536 5918
rect 2550 5914 2552 5918
rect 2566 5914 2568 5918
rect 2571 5914 2573 5918
rect 2587 5914 2589 5918
rect 2603 5914 2605 5918
rect 2624 5914 2626 5918
rect 2629 5914 2631 5918
rect 2645 5914 2647 5918
rect 2661 5914 2663 5918
rect 2666 5914 2668 5918
rect 2682 5914 2684 5918
rect 2698 5914 2700 5918
rect 2703 5914 2705 5918
rect 2719 5914 2721 5918
rect 2735 5914 2737 5918
rect 2756 5914 2758 5918
rect 2761 5914 2763 5918
rect 2777 5914 2779 5918
rect 2793 5914 2795 5918
rect 2798 5914 2800 5918
rect 1597 5852 1599 5856
rect 1621 5852 1623 5856
rect 2542 5852 2544 5856
rect 2566 5852 2568 5856
rect 1608 5845 1612 5847
rect 2553 5845 2557 5847
rect 1601 5829 1603 5833
rect 2546 5829 2548 5833
rect 1597 5818 1599 5822
rect 1621 5818 1623 5822
rect 2542 5818 2544 5822
rect 2566 5818 2568 5822
rect 1473 5774 1475 5778
rect 1489 5774 1491 5778
rect 1494 5774 1496 5778
rect 1510 5774 1512 5778
rect 1526 5774 1528 5778
rect 1547 5774 1549 5778
rect 1552 5774 1554 5778
rect 1568 5774 1570 5778
rect 1584 5774 1586 5778
rect 1589 5774 1591 5778
rect 1605 5774 1607 5778
rect 1621 5774 1623 5778
rect 1626 5774 1628 5778
rect 1642 5774 1644 5778
rect 1658 5774 1660 5778
rect 1679 5774 1681 5778
rect 1684 5774 1686 5778
rect 1700 5774 1702 5778
rect 1716 5774 1718 5778
rect 1721 5774 1723 5778
rect 1737 5774 1739 5778
rect 1753 5774 1755 5778
rect 1758 5774 1760 5778
rect 1774 5774 1776 5778
rect 1790 5774 1792 5778
rect 1811 5774 1813 5778
rect 1816 5774 1818 5778
rect 1832 5774 1834 5778
rect 1848 5774 1850 5778
rect 1853 5774 1855 5778
rect 2418 5774 2420 5778
rect 2434 5774 2436 5778
rect 2439 5774 2441 5778
rect 2455 5774 2457 5778
rect 2471 5774 2473 5778
rect 2492 5774 2494 5778
rect 2497 5774 2499 5778
rect 2513 5774 2515 5778
rect 2529 5774 2531 5778
rect 2534 5774 2536 5778
rect 2550 5774 2552 5778
rect 2566 5774 2568 5778
rect 2571 5774 2573 5778
rect 2587 5774 2589 5778
rect 2603 5774 2605 5778
rect 2624 5774 2626 5778
rect 2629 5774 2631 5778
rect 2645 5774 2647 5778
rect 2661 5774 2663 5778
rect 2666 5774 2668 5778
rect 2682 5774 2684 5778
rect 2698 5774 2700 5778
rect 2703 5774 2705 5778
rect 2719 5774 2721 5778
rect 2735 5774 2737 5778
rect 2756 5774 2758 5778
rect 2761 5774 2763 5778
rect 2777 5774 2779 5778
rect 2793 5774 2795 5778
rect 2798 5774 2800 5778
rect 954 5744 956 5748
rect 970 5744 972 5748
rect 975 5744 977 5748
rect 991 5744 993 5748
rect 1007 5744 1009 5748
rect 1028 5744 1030 5748
rect 1033 5744 1035 5748
rect 1049 5744 1051 5748
rect 1065 5744 1067 5748
rect 1070 5744 1072 5748
rect 1899 5744 1901 5748
rect 1915 5744 1917 5748
rect 1920 5744 1922 5748
rect 1936 5744 1938 5748
rect 1952 5744 1954 5748
rect 1973 5744 1975 5748
rect 1978 5744 1980 5748
rect 1994 5744 1996 5748
rect 2010 5744 2012 5748
rect 2015 5744 2017 5748
rect 927 5736 931 5738
rect 1872 5736 1876 5738
rect 1473 5688 1475 5692
rect 1489 5688 1491 5692
rect 1494 5688 1496 5692
rect 1510 5688 1512 5692
rect 1526 5688 1528 5692
rect 1547 5688 1549 5692
rect 1552 5688 1554 5692
rect 1568 5688 1570 5692
rect 1584 5688 1586 5692
rect 1589 5688 1591 5692
rect 1605 5688 1607 5692
rect 1621 5688 1623 5692
rect 1626 5688 1628 5692
rect 1642 5688 1644 5692
rect 1658 5688 1660 5692
rect 1679 5688 1681 5692
rect 1684 5688 1686 5692
rect 1700 5688 1702 5692
rect 1716 5688 1718 5692
rect 1721 5688 1723 5692
rect 1737 5688 1739 5692
rect 1753 5688 1755 5692
rect 1758 5688 1760 5692
rect 1774 5688 1776 5692
rect 1790 5688 1792 5692
rect 1811 5688 1813 5692
rect 1816 5688 1818 5692
rect 1832 5688 1834 5692
rect 1848 5688 1850 5692
rect 1853 5688 1855 5692
rect 2418 5688 2420 5692
rect 2434 5688 2436 5692
rect 2439 5688 2441 5692
rect 2455 5688 2457 5692
rect 2471 5688 2473 5692
rect 2492 5688 2494 5692
rect 2497 5688 2499 5692
rect 2513 5688 2515 5692
rect 2529 5688 2531 5692
rect 2534 5688 2536 5692
rect 2550 5688 2552 5692
rect 2566 5688 2568 5692
rect 2571 5688 2573 5692
rect 2587 5688 2589 5692
rect 2603 5688 2605 5692
rect 2624 5688 2626 5692
rect 2629 5688 2631 5692
rect 2645 5688 2647 5692
rect 2661 5688 2663 5692
rect 2666 5688 2668 5692
rect 2682 5688 2684 5692
rect 2698 5688 2700 5692
rect 2703 5688 2705 5692
rect 2719 5688 2721 5692
rect 2735 5688 2737 5692
rect 2756 5688 2758 5692
rect 2761 5688 2763 5692
rect 2777 5688 2779 5692
rect 2793 5688 2795 5692
rect 2798 5688 2800 5692
rect 954 5658 956 5662
rect 970 5658 972 5662
rect 975 5658 977 5662
rect 991 5658 993 5662
rect 1007 5658 1009 5662
rect 1028 5658 1030 5662
rect 1033 5658 1035 5662
rect 1049 5658 1051 5662
rect 1065 5658 1067 5662
rect 1070 5658 1072 5662
rect 1899 5658 1901 5662
rect 1915 5658 1917 5662
rect 1920 5658 1922 5662
rect 1936 5658 1938 5662
rect 1952 5658 1954 5662
rect 1973 5658 1975 5662
rect 1978 5658 1980 5662
rect 1994 5658 1996 5662
rect 2010 5658 2012 5662
rect 2015 5658 2017 5662
rect 1714 5626 1716 5630
rect 1738 5626 1740 5630
rect 2659 5626 2661 5630
rect 2683 5626 2685 5630
rect 1725 5619 1729 5621
rect 2670 5619 2674 5621
rect 1718 5603 1720 5607
rect 2663 5603 2665 5607
rect 939 5590 943 5592
rect 1714 5590 1716 5594
rect 1738 5590 1740 5594
rect 1884 5590 1888 5592
rect 2659 5590 2661 5594
rect 2683 5590 2685 5594
rect 1159 5539 1161 5543
rect 1164 5539 1166 5543
rect 1473 5546 1475 5550
rect 1489 5546 1491 5550
rect 1494 5546 1496 5550
rect 1510 5546 1512 5550
rect 1526 5546 1528 5550
rect 1547 5546 1549 5550
rect 1552 5546 1554 5550
rect 1568 5546 1570 5550
rect 1584 5546 1586 5550
rect 1589 5546 1591 5550
rect 1605 5546 1607 5550
rect 1621 5546 1623 5550
rect 1626 5546 1628 5550
rect 1642 5546 1644 5550
rect 1658 5546 1660 5550
rect 1679 5546 1681 5550
rect 1684 5546 1686 5550
rect 1700 5546 1702 5550
rect 1716 5546 1718 5550
rect 1721 5546 1723 5550
rect 1737 5546 1739 5550
rect 1753 5546 1755 5550
rect 1758 5546 1760 5550
rect 1774 5546 1776 5550
rect 1790 5546 1792 5550
rect 1811 5546 1813 5550
rect 1816 5546 1818 5550
rect 1832 5546 1834 5550
rect 1848 5546 1850 5550
rect 1853 5546 1855 5550
rect 953 5532 955 5536
rect 971 5532 973 5536
rect 976 5532 978 5536
rect 996 5532 998 5536
rect 1017 5532 1019 5536
rect 1043 5532 1045 5536
rect 1048 5532 1050 5536
rect 1071 5532 1073 5536
rect 1087 5532 1089 5536
rect 1112 5532 1114 5536
rect 1130 5532 1132 5536
rect 1214 5532 1216 5536
rect 1232 5532 1234 5536
rect 1237 5532 1239 5536
rect 1257 5532 1259 5536
rect 1278 5532 1280 5536
rect 1304 5532 1306 5536
rect 1309 5532 1311 5536
rect 1332 5532 1334 5536
rect 1348 5532 1350 5536
rect 1364 5532 1366 5536
rect 2104 5539 2106 5543
rect 2109 5539 2111 5543
rect 2418 5546 2420 5550
rect 2434 5546 2436 5550
rect 2439 5546 2441 5550
rect 2455 5546 2457 5550
rect 2471 5546 2473 5550
rect 2492 5546 2494 5550
rect 2497 5546 2499 5550
rect 2513 5546 2515 5550
rect 2529 5546 2531 5550
rect 2534 5546 2536 5550
rect 2550 5546 2552 5550
rect 2566 5546 2568 5550
rect 2571 5546 2573 5550
rect 2587 5546 2589 5550
rect 2603 5546 2605 5550
rect 2624 5546 2626 5550
rect 2629 5546 2631 5550
rect 2645 5546 2647 5550
rect 2661 5546 2663 5550
rect 2666 5546 2668 5550
rect 2682 5546 2684 5550
rect 2698 5546 2700 5550
rect 2703 5546 2705 5550
rect 2719 5546 2721 5550
rect 2735 5546 2737 5550
rect 2756 5546 2758 5550
rect 2761 5546 2763 5550
rect 2777 5546 2779 5550
rect 2793 5546 2795 5550
rect 2798 5546 2800 5550
rect 1898 5532 1900 5536
rect 1916 5532 1918 5536
rect 1921 5532 1923 5536
rect 1941 5532 1943 5536
rect 1962 5532 1964 5536
rect 1988 5532 1990 5536
rect 1993 5532 1995 5536
rect 2016 5532 2018 5536
rect 2032 5532 2034 5536
rect 2057 5532 2059 5536
rect 2075 5532 2077 5536
rect 2159 5532 2161 5536
rect 2177 5532 2179 5536
rect 2182 5532 2184 5536
rect 2202 5532 2204 5536
rect 2223 5532 2225 5536
rect 2249 5532 2251 5536
rect 2254 5532 2256 5536
rect 2277 5532 2279 5536
rect 2293 5532 2295 5536
rect 2309 5532 2311 5536
rect 1214 5486 1216 5490
rect 1232 5486 1234 5490
rect 1237 5486 1239 5490
rect 1257 5486 1259 5490
rect 1278 5486 1280 5490
rect 1304 5486 1306 5490
rect 1309 5486 1311 5490
rect 1332 5486 1334 5490
rect 1348 5486 1350 5490
rect 1364 5486 1366 5490
rect 1136 5481 1138 5485
rect 1159 5477 1161 5481
rect 1164 5477 1166 5481
rect 2159 5486 2161 5490
rect 2177 5486 2179 5490
rect 2182 5486 2184 5490
rect 2202 5486 2204 5490
rect 2223 5486 2225 5490
rect 2249 5486 2251 5490
rect 2254 5486 2256 5490
rect 2277 5486 2279 5490
rect 2293 5486 2295 5490
rect 2309 5486 2311 5490
rect 2081 5481 2083 5485
rect 2104 5477 2106 5481
rect 2109 5477 2111 5481
rect 1768 5432 1770 5436
rect 1773 5432 1775 5436
rect 988 5403 990 5407
rect 993 5403 995 5407
rect 1078 5403 1080 5407
rect 1083 5403 1085 5407
rect 1159 5403 1161 5407
rect 1164 5403 1166 5407
rect 1214 5400 1216 5404
rect 1232 5400 1234 5404
rect 1237 5400 1239 5404
rect 1257 5400 1259 5404
rect 1278 5400 1280 5404
rect 1304 5400 1306 5404
rect 1309 5400 1311 5404
rect 1332 5400 1334 5404
rect 1348 5400 1350 5404
rect 1364 5400 1366 5404
rect 1654 5399 1656 5411
rect 1707 5399 1709 5411
rect 1933 5403 1935 5407
rect 1938 5403 1940 5407
rect 2023 5403 2025 5407
rect 2028 5403 2030 5407
rect 2104 5403 2106 5407
rect 2109 5403 2111 5407
rect 2159 5400 2161 5404
rect 2177 5400 2179 5404
rect 2182 5400 2184 5404
rect 2202 5400 2204 5404
rect 2223 5400 2225 5404
rect 2249 5400 2251 5404
rect 2254 5400 2256 5404
rect 2277 5400 2279 5404
rect 2293 5400 2295 5404
rect 2309 5400 2311 5404
rect 965 5349 967 5353
rect 1055 5349 1057 5353
rect 1214 5354 1216 5358
rect 1232 5354 1234 5358
rect 1237 5354 1239 5358
rect 1257 5354 1259 5358
rect 1278 5354 1280 5358
rect 1304 5354 1306 5358
rect 1309 5354 1311 5358
rect 1332 5354 1334 5358
rect 1348 5354 1350 5358
rect 1364 5354 1366 5358
rect 1136 5349 1138 5353
rect 988 5345 990 5349
rect 993 5345 995 5349
rect 1019 5341 1021 5345
rect 1078 5345 1080 5349
rect 1083 5345 1085 5349
rect 1109 5341 1111 5345
rect 1159 5345 1161 5349
rect 1164 5345 1166 5349
rect 1745 5376 1747 5380
rect 1768 5372 1770 5376
rect 1773 5372 1775 5376
rect 1799 5368 1801 5372
rect 1821 5368 1823 5372
rect 1910 5349 1912 5353
rect 2000 5349 2002 5353
rect 2159 5354 2161 5358
rect 2177 5354 2179 5358
rect 2182 5354 2184 5358
rect 2202 5354 2204 5358
rect 2223 5354 2225 5358
rect 2249 5354 2251 5358
rect 2254 5354 2256 5358
rect 2277 5354 2279 5358
rect 2293 5354 2295 5358
rect 2309 5354 2311 5358
rect 2081 5349 2083 5353
rect 1933 5345 1935 5349
rect 1938 5345 1940 5349
rect 1964 5341 1966 5345
rect 2023 5345 2025 5349
rect 2028 5345 2030 5349
rect 2054 5341 2056 5345
rect 2104 5345 2106 5349
rect 2109 5345 2111 5349
rect 1768 5302 1770 5306
rect 1773 5302 1775 5306
rect 1054 5268 1056 5272
rect 1059 5268 1061 5272
rect 1159 5268 1161 5272
rect 1164 5268 1166 5272
rect 1214 5268 1216 5272
rect 1232 5268 1234 5272
rect 1237 5268 1239 5272
rect 1257 5268 1259 5272
rect 1278 5268 1280 5272
rect 1304 5268 1306 5272
rect 1309 5268 1311 5272
rect 1332 5268 1334 5272
rect 1348 5268 1350 5272
rect 1364 5268 1366 5272
rect 1560 5269 1562 5281
rect 1613 5269 1615 5281
rect 1999 5268 2001 5272
rect 2004 5268 2006 5272
rect 2104 5268 2106 5272
rect 2109 5268 2111 5272
rect 2159 5268 2161 5272
rect 2177 5268 2179 5272
rect 2182 5268 2184 5272
rect 2202 5268 2204 5272
rect 2223 5268 2225 5272
rect 2249 5268 2251 5272
rect 2254 5268 2256 5272
rect 2277 5268 2279 5272
rect 2293 5268 2295 5272
rect 2309 5268 2311 5272
rect 1031 5217 1033 5221
rect 1214 5222 1216 5226
rect 1232 5222 1234 5226
rect 1237 5222 1239 5226
rect 1257 5222 1259 5226
rect 1278 5222 1280 5226
rect 1304 5222 1306 5226
rect 1309 5222 1311 5226
rect 1332 5222 1334 5226
rect 1348 5222 1350 5226
rect 1364 5222 1366 5226
rect 1136 5217 1138 5221
rect 1054 5213 1056 5217
rect 1059 5213 1061 5217
rect 1085 5209 1087 5213
rect 1159 5213 1161 5217
rect 1164 5213 1166 5217
rect 1745 5246 1747 5250
rect 1768 5242 1770 5246
rect 1773 5242 1775 5246
rect 1799 5238 1801 5242
rect 1976 5217 1978 5221
rect 2159 5222 2161 5226
rect 2177 5222 2179 5226
rect 2182 5222 2184 5226
rect 2202 5222 2204 5226
rect 2223 5222 2225 5226
rect 2249 5222 2251 5226
rect 2254 5222 2256 5226
rect 2277 5222 2279 5226
rect 2293 5222 2295 5226
rect 2309 5222 2311 5226
rect 2081 5217 2083 5221
rect 1999 5213 2001 5217
rect 2004 5213 2006 5217
rect 2030 5209 2032 5213
rect 2104 5213 2106 5217
rect 2109 5213 2111 5217
rect 1078 5137 1080 5141
rect 1083 5137 1085 5141
rect 1159 5137 1161 5141
rect 1164 5137 1166 5141
rect 1614 5146 1616 5150
rect 1619 5146 1621 5150
rect 1635 5146 1637 5150
rect 1651 5146 1653 5150
rect 1656 5146 1658 5150
rect 1677 5146 1679 5150
rect 1693 5146 1695 5150
rect 1709 5146 1711 5150
rect 1714 5146 1716 5150
rect 1730 5146 1732 5150
rect 1214 5136 1216 5140
rect 1232 5136 1234 5140
rect 1237 5136 1239 5140
rect 1257 5136 1259 5140
rect 1278 5136 1280 5140
rect 1304 5136 1306 5140
rect 1309 5136 1311 5140
rect 1332 5136 1334 5140
rect 1348 5136 1350 5140
rect 1364 5136 1366 5140
rect 2023 5137 2025 5141
rect 2028 5137 2030 5141
rect 2104 5137 2106 5141
rect 2109 5137 2111 5141
rect 2559 5146 2561 5150
rect 2564 5146 2566 5150
rect 2580 5146 2582 5150
rect 2596 5146 2598 5150
rect 2601 5146 2603 5150
rect 2622 5146 2624 5150
rect 2638 5146 2640 5150
rect 2654 5146 2656 5150
rect 2659 5146 2661 5150
rect 2675 5146 2677 5150
rect 2159 5136 2161 5140
rect 2177 5136 2179 5140
rect 2182 5136 2184 5140
rect 2202 5136 2204 5140
rect 2223 5136 2225 5140
rect 2249 5136 2251 5140
rect 2254 5136 2256 5140
rect 2277 5136 2279 5140
rect 2293 5136 2295 5140
rect 2309 5136 2311 5140
rect 1055 5085 1057 5089
rect 1214 5090 1216 5094
rect 1232 5090 1234 5094
rect 1237 5090 1239 5094
rect 1257 5090 1259 5094
rect 1278 5090 1280 5094
rect 1304 5090 1306 5094
rect 1309 5090 1311 5094
rect 1332 5090 1334 5094
rect 1348 5090 1350 5094
rect 1364 5090 1366 5094
rect 1714 5090 1716 5094
rect 1136 5085 1138 5089
rect 1078 5081 1080 5085
rect 1083 5081 1085 5085
rect 1109 5077 1111 5081
rect 1159 5081 1161 5085
rect 1164 5081 1166 5085
rect 1190 5077 1192 5081
rect 1597 5081 1599 5085
rect 2000 5085 2002 5089
rect 2159 5090 2161 5094
rect 2177 5090 2179 5094
rect 2182 5090 2184 5094
rect 2202 5090 2204 5094
rect 2223 5090 2225 5094
rect 2249 5090 2251 5094
rect 2254 5090 2256 5094
rect 2277 5090 2279 5094
rect 2293 5090 2295 5094
rect 2309 5090 2311 5094
rect 2659 5090 2661 5094
rect 2081 5085 2083 5089
rect 2023 5081 2025 5085
rect 2028 5081 2030 5085
rect 2054 5077 2056 5081
rect 2104 5081 2106 5085
rect 2109 5081 2111 5085
rect 2135 5077 2137 5081
rect 2542 5081 2544 5085
rect 1605 5044 1607 5048
rect 1621 5044 1623 5048
rect 1626 5044 1628 5048
rect 1642 5044 1644 5048
rect 1658 5044 1660 5048
rect 1679 5044 1681 5048
rect 1684 5044 1686 5048
rect 1700 5044 1702 5048
rect 1716 5044 1718 5048
rect 1721 5044 1723 5048
rect 2550 5044 2552 5048
rect 2566 5044 2568 5048
rect 2571 5044 2573 5048
rect 2587 5044 2589 5048
rect 2603 5044 2605 5048
rect 2624 5044 2626 5048
rect 2629 5044 2631 5048
rect 2645 5044 2647 5048
rect 2661 5044 2663 5048
rect 2666 5044 2668 5048
rect 857 5011 859 5015
rect 873 5011 875 5015
rect 878 5011 880 5015
rect 894 5011 896 5015
rect 910 5011 912 5015
rect 931 5011 933 5015
rect 936 5011 938 5015
rect 952 5011 954 5015
rect 968 5011 970 5015
rect 973 5011 975 5015
rect 989 5011 991 5015
rect 1005 5011 1007 5015
rect 1010 5011 1012 5015
rect 1026 5011 1028 5015
rect 1042 5011 1044 5015
rect 1063 5011 1065 5015
rect 1068 5011 1070 5015
rect 1084 5011 1086 5015
rect 1100 5011 1102 5015
rect 1105 5011 1107 5015
rect 1121 5011 1123 5015
rect 1137 5011 1139 5015
rect 1142 5011 1144 5015
rect 1158 5011 1160 5015
rect 1174 5011 1176 5015
rect 1195 5011 1197 5015
rect 1200 5011 1202 5015
rect 1216 5011 1218 5015
rect 1232 5011 1234 5015
rect 1237 5011 1239 5015
rect 1253 5011 1255 5015
rect 1269 5011 1271 5015
rect 1274 5011 1276 5015
rect 1290 5011 1292 5015
rect 1306 5011 1308 5015
rect 1327 5011 1329 5015
rect 1332 5011 1334 5015
rect 1348 5011 1350 5015
rect 1364 5011 1366 5015
rect 1369 5011 1371 5015
rect 1802 5011 1804 5015
rect 1818 5011 1820 5015
rect 1823 5011 1825 5015
rect 1839 5011 1841 5015
rect 1855 5011 1857 5015
rect 1876 5011 1878 5015
rect 1881 5011 1883 5015
rect 1897 5011 1899 5015
rect 1913 5011 1915 5015
rect 1918 5011 1920 5015
rect 1934 5011 1936 5015
rect 1950 5011 1952 5015
rect 1955 5011 1957 5015
rect 1971 5011 1973 5015
rect 1987 5011 1989 5015
rect 2008 5011 2010 5015
rect 2013 5011 2015 5015
rect 2029 5011 2031 5015
rect 2045 5011 2047 5015
rect 2050 5011 2052 5015
rect 2066 5011 2068 5015
rect 2082 5011 2084 5015
rect 2087 5011 2089 5015
rect 2103 5011 2105 5015
rect 2119 5011 2121 5015
rect 2140 5011 2142 5015
rect 2145 5011 2147 5015
rect 2161 5011 2163 5015
rect 2177 5011 2179 5015
rect 2182 5011 2184 5015
rect 2198 5011 2200 5015
rect 2214 5011 2216 5015
rect 2219 5011 2221 5015
rect 2235 5011 2237 5015
rect 2251 5011 2253 5015
rect 2272 5011 2274 5015
rect 2277 5011 2279 5015
rect 2293 5011 2295 5015
rect 2309 5011 2311 5015
rect 2314 5011 2316 5015
rect 4579 7975 4581 8015
rect 4587 7975 4589 8015
rect 4595 7975 4597 8015
rect 4603 7975 4605 8015
rect 4611 7975 4613 8015
rect 4619 7975 4621 8015
rect 4634 7975 4636 8034
rect 4642 7975 4644 8034
rect 4650 7975 4652 8034
rect 4658 7975 4660 8034
rect 4677 7975 4679 8034
rect 4685 7975 4687 8034
rect 4693 7975 4695 8034
rect 4701 7975 4703 8034
rect 4718 7975 4720 8034
rect 4726 7975 4728 8034
rect 4734 7975 4736 8034
rect 4742 7975 4744 8034
rect 4577 7302 4579 7342
rect 4585 7302 4587 7342
rect 4593 7302 4595 7342
rect 4601 7302 4603 7342
rect 4609 7302 4611 7342
rect 4617 7302 4619 7342
rect 1140 4528 1180 4530
rect 1140 4520 1180 4522
rect 1140 4512 1180 4514
rect 1140 4504 1180 4506
rect 2067 4528 2107 4530
rect 2067 4520 2107 4522
rect 2067 4512 2107 4514
rect 2067 4504 2107 4506
rect 2376 4528 2416 4530
rect 2376 4520 2416 4522
rect 2376 4512 2416 4514
rect 2376 4504 2416 4506
rect 2685 4528 2725 4530
rect 2685 4520 2725 4522
rect 2685 4512 2725 4514
rect 2685 4504 2725 4506
rect 2994 4528 3034 4530
rect 2994 4520 3034 4522
rect 2994 4512 3034 4514
rect 2994 4504 3034 4506
rect 3303 4528 3343 4530
rect 3303 4520 3343 4522
rect 3303 4512 3343 4514
rect 3303 4504 3343 4506
rect 1140 4496 1180 4498
rect 2067 4496 2107 4498
rect 2376 4496 2416 4498
rect 2685 4496 2725 4498
rect 2994 4496 3034 4498
rect 3303 4496 3343 4498
rect 1140 4488 1180 4490
rect 2067 4488 2107 4490
rect 2376 4488 2416 4490
rect 2685 4488 2725 4490
rect 2994 4488 3034 4490
rect 3303 4488 3343 4490
<< ptransistor >>
rect 1743 9824 1799 9826
rect 2052 9824 2108 9826
rect 2361 9824 2417 9826
rect 2670 9824 2726 9826
rect 2979 9824 3035 9826
rect 3906 9824 3962 9826
rect 1743 9816 1799 9818
rect 2052 9816 2108 9818
rect 2361 9816 2417 9818
rect 2670 9816 2726 9818
rect 2979 9816 3035 9818
rect 3906 9816 3962 9818
rect 1743 9808 1799 9810
rect 1743 9800 1799 9802
rect 1743 9792 1799 9794
rect 1743 9784 1799 9786
rect 2052 9808 2108 9810
rect 2052 9800 2108 9802
rect 2052 9792 2108 9794
rect 2052 9784 2108 9786
rect 2361 9808 2417 9810
rect 2361 9800 2417 9802
rect 2361 9792 2417 9794
rect 2361 9784 2417 9786
rect 2670 9808 2726 9810
rect 2670 9800 2726 9802
rect 2670 9792 2726 9794
rect 2670 9784 2726 9786
rect 2979 9808 3035 9810
rect 2979 9800 3035 9802
rect 2979 9792 3035 9794
rect 2979 9784 3035 9786
rect 3906 9808 3962 9810
rect 3906 9800 3962 9802
rect 3906 9792 3962 9794
rect 3906 9784 3962 9786
rect 428 6369 430 6457
rect 436 6369 438 6457
rect 444 6369 446 6457
rect 452 6369 454 6457
rect 469 6369 471 6457
rect 477 6369 479 6457
rect 485 6369 487 6457
rect 493 6369 495 6457
rect 512 6369 514 6457
rect 520 6369 522 6457
rect 528 6369 530 6457
rect 536 6369 538 6457
rect 551 6369 553 6425
rect 559 6369 561 6425
rect 567 6369 569 6425
rect 575 6369 577 6425
rect 583 6369 585 6425
rect 591 6369 593 6425
rect 2856 9322 2858 9330
rect 2861 9322 2863 9330
rect 2877 9322 2879 9330
rect 2893 9322 2895 9330
rect 2898 9322 2900 9330
rect 2919 9322 2921 9330
rect 2935 9322 2937 9330
rect 2951 9322 2953 9330
rect 2956 9322 2958 9330
rect 2972 9322 2974 9330
rect 2988 9322 2990 9330
rect 2993 9322 2995 9330
rect 3009 9322 3011 9330
rect 3025 9322 3027 9330
rect 3030 9322 3032 9330
rect 3051 9322 3053 9330
rect 3067 9322 3069 9330
rect 3083 9322 3085 9330
rect 3088 9322 3090 9330
rect 3104 9322 3106 9330
rect 3120 9322 3122 9330
rect 3125 9322 3127 9330
rect 3141 9322 3143 9330
rect 3157 9322 3159 9330
rect 3162 9322 3164 9330
rect 3183 9322 3185 9330
rect 3199 9322 3201 9330
rect 3215 9322 3217 9330
rect 3220 9322 3222 9330
rect 3236 9322 3238 9330
rect 3252 9322 3254 9330
rect 3257 9322 3259 9330
rect 3273 9322 3275 9330
rect 3289 9322 3291 9330
rect 3294 9322 3296 9330
rect 3315 9322 3317 9330
rect 3331 9322 3333 9330
rect 3347 9322 3349 9330
rect 3352 9322 3354 9330
rect 3368 9322 3370 9330
rect 3801 9322 3803 9330
rect 3806 9322 3808 9330
rect 3822 9322 3824 9330
rect 3838 9322 3840 9330
rect 3843 9322 3845 9330
rect 3864 9322 3866 9330
rect 3880 9322 3882 9330
rect 3896 9322 3898 9330
rect 3901 9322 3903 9330
rect 3917 9322 3919 9330
rect 3933 9322 3935 9330
rect 3938 9322 3940 9330
rect 3954 9322 3956 9330
rect 3970 9322 3972 9330
rect 3975 9322 3977 9330
rect 3996 9322 3998 9330
rect 4012 9322 4014 9330
rect 4028 9322 4030 9330
rect 4033 9322 4035 9330
rect 4049 9322 4051 9330
rect 4065 9322 4067 9330
rect 4070 9322 4072 9330
rect 4086 9322 4088 9330
rect 4102 9322 4104 9330
rect 4107 9322 4109 9330
rect 4128 9322 4130 9330
rect 4144 9322 4146 9330
rect 4160 9322 4162 9330
rect 4165 9322 4167 9330
rect 4181 9322 4183 9330
rect 4197 9322 4199 9330
rect 4202 9322 4204 9330
rect 4218 9322 4220 9330
rect 4234 9322 4236 9330
rect 4239 9322 4241 9330
rect 4260 9322 4262 9330
rect 4276 9322 4278 9330
rect 4292 9322 4294 9330
rect 4297 9322 4299 9330
rect 4313 9322 4315 9330
rect 2504 9289 2506 9297
rect 2509 9289 2511 9297
rect 2525 9289 2527 9297
rect 2541 9289 2543 9297
rect 2546 9289 2548 9297
rect 2567 9289 2569 9297
rect 2583 9289 2585 9297
rect 2599 9289 2601 9297
rect 2604 9289 2606 9297
rect 2620 9289 2622 9297
rect 3449 9289 3451 9297
rect 3454 9289 3456 9297
rect 3470 9289 3472 9297
rect 3486 9289 3488 9297
rect 3491 9289 3493 9297
rect 3512 9289 3514 9297
rect 3528 9289 3530 9297
rect 3544 9289 3546 9297
rect 3549 9289 3551 9297
rect 3565 9289 3567 9297
rect 3035 9251 3037 9259
rect 2861 9238 2863 9246
rect 2877 9238 2879 9246
rect 2893 9238 2895 9246
rect 2916 9238 2918 9246
rect 2921 9238 2923 9246
rect 2947 9238 2949 9246
rect 2968 9238 2970 9246
rect 2988 9238 2990 9246
rect 2993 9238 2995 9246
rect 3011 9238 3013 9246
rect 3061 9245 3063 9253
rect 3066 9245 3068 9253
rect 3089 9251 3091 9259
rect 3116 9251 3118 9259
rect 3142 9245 3144 9253
rect 3147 9245 3149 9253
rect 3170 9251 3172 9259
rect 3980 9251 3982 9259
rect 3806 9238 3808 9246
rect 3822 9238 3824 9246
rect 3838 9238 3840 9246
rect 3861 9238 3863 9246
rect 3866 9238 3868 9246
rect 3892 9238 3894 9246
rect 3913 9238 3915 9246
rect 3933 9238 3935 9246
rect 3938 9238 3940 9246
rect 3956 9238 3958 9246
rect 4006 9245 4008 9253
rect 4011 9245 4013 9253
rect 4034 9251 4036 9259
rect 4061 9251 4063 9259
rect 4087 9245 4089 9253
rect 4092 9245 4094 9253
rect 4115 9251 4117 9259
rect 2495 9187 2497 9195
rect 2511 9187 2513 9195
rect 2516 9187 2518 9195
rect 2532 9187 2534 9195
rect 2548 9187 2550 9195
rect 2569 9187 2571 9195
rect 2574 9187 2576 9195
rect 2590 9187 2592 9195
rect 2606 9187 2608 9195
rect 2611 9187 2613 9195
rect 3440 9187 3442 9195
rect 3456 9187 3458 9195
rect 3461 9187 3463 9195
rect 3477 9187 3479 9195
rect 3493 9187 3495 9195
rect 3514 9187 3516 9195
rect 3519 9187 3521 9195
rect 3535 9187 3537 9195
rect 3551 9187 3553 9195
rect 3556 9187 3558 9195
rect 2861 9152 2863 9160
rect 2877 9152 2879 9160
rect 2893 9152 2895 9160
rect 2916 9152 2918 9160
rect 2921 9152 2923 9160
rect 2947 9152 2949 9160
rect 2968 9152 2970 9160
rect 2988 9152 2990 9160
rect 2993 9152 2995 9160
rect 3011 9152 3013 9160
rect 3061 9153 3063 9161
rect 3066 9153 3068 9161
rect 3142 9153 3144 9161
rect 3147 9153 3149 9161
rect 3806 9152 3808 9160
rect 3822 9152 3824 9160
rect 3838 9152 3840 9160
rect 3861 9152 3863 9160
rect 3866 9152 3868 9160
rect 3892 9152 3894 9160
rect 3913 9152 3915 9160
rect 3933 9152 3935 9160
rect 3938 9152 3940 9160
rect 3956 9152 3958 9160
rect 4006 9153 4008 9161
rect 4011 9153 4013 9161
rect 4087 9153 4089 9161
rect 4092 9153 4094 9161
rect 2861 9106 2863 9114
rect 2877 9106 2879 9114
rect 2893 9106 2895 9114
rect 2916 9106 2918 9114
rect 2921 9106 2923 9114
rect 2947 9106 2949 9114
rect 2968 9106 2970 9114
rect 2988 9106 2990 9114
rect 2993 9106 2995 9114
rect 3011 9106 3013 9114
rect 3061 9113 3063 9121
rect 3066 9113 3068 9121
rect 3089 9119 3091 9127
rect 3140 9119 3142 9127
rect 3166 9113 3168 9121
rect 3171 9113 3173 9121
rect 3194 9119 3196 9127
rect 3806 9106 3808 9114
rect 3822 9106 3824 9114
rect 3838 9106 3840 9114
rect 3861 9106 3863 9114
rect 3866 9106 3868 9114
rect 3892 9106 3894 9114
rect 3913 9106 3915 9114
rect 3933 9106 3935 9114
rect 3938 9106 3940 9114
rect 3956 9106 3958 9114
rect 4006 9113 4008 9121
rect 4011 9113 4013 9121
rect 4034 9119 4036 9127
rect 4085 9119 4087 9127
rect 3371 9090 3373 9098
rect 3397 9084 3399 9092
rect 3402 9084 3404 9092
rect 3425 9090 3427 9098
rect 3557 9065 3559 9095
rect 3610 9065 3612 9095
rect 4111 9113 4113 9121
rect 4116 9113 4118 9121
rect 4139 9119 4141 9127
rect 2861 9020 2863 9028
rect 2877 9020 2879 9028
rect 2893 9020 2895 9028
rect 2916 9020 2918 9028
rect 2921 9020 2923 9028
rect 2947 9020 2949 9028
rect 2968 9020 2970 9028
rect 2988 9020 2990 9028
rect 2993 9020 2995 9028
rect 3011 9020 3013 9028
rect 3061 9022 3063 9030
rect 3066 9022 3068 9030
rect 3166 9022 3168 9030
rect 3171 9022 3173 9030
rect 3806 9020 3808 9028
rect 3822 9020 3824 9028
rect 3838 9020 3840 9028
rect 3861 9020 3863 9028
rect 3866 9020 3868 9028
rect 3892 9020 3894 9028
rect 3913 9020 3915 9028
rect 3933 9020 3935 9028
rect 3938 9020 3940 9028
rect 3956 9020 3958 9028
rect 4006 9022 4008 9030
rect 4011 9022 4013 9030
rect 4111 9022 4113 9030
rect 4116 9022 4118 9030
rect 2861 8974 2863 8982
rect 2877 8974 2879 8982
rect 2893 8974 2895 8982
rect 2916 8974 2918 8982
rect 2921 8974 2923 8982
rect 2947 8974 2949 8982
rect 2968 8974 2970 8982
rect 2988 8974 2990 8982
rect 2993 8974 2995 8982
rect 3011 8974 3013 8982
rect 3061 8981 3063 8989
rect 3066 8981 3068 8989
rect 3089 8987 3091 8995
rect 3116 8987 3118 8995
rect 3142 8981 3144 8989
rect 3147 8981 3149 8989
rect 3170 8987 3172 8995
rect 3206 8987 3208 8995
rect 3232 8981 3234 8989
rect 3237 8981 3239 8989
rect 3260 8987 3262 8995
rect 3397 8988 3399 8996
rect 3402 8988 3404 8996
rect 3806 8974 3808 8982
rect 3822 8974 3824 8982
rect 3838 8974 3840 8982
rect 3861 8974 3863 8982
rect 3866 8974 3868 8982
rect 3892 8974 3894 8982
rect 3913 8974 3915 8982
rect 3933 8974 3935 8982
rect 3938 8974 3940 8982
rect 3956 8974 3958 8982
rect 4006 8981 4008 8989
rect 4011 8981 4013 8989
rect 4034 8987 4036 8995
rect 4061 8987 4063 8995
rect 3349 8960 3351 8968
rect 3371 8960 3373 8968
rect 3397 8954 3399 8962
rect 3402 8954 3404 8962
rect 3425 8960 3427 8968
rect 3463 8935 3465 8965
rect 3516 8935 3518 8965
rect 4087 8981 4089 8989
rect 4092 8981 4094 8989
rect 4115 8987 4117 8995
rect 4151 8987 4153 8995
rect 4177 8981 4179 8989
rect 4182 8981 4184 8989
rect 4205 8987 4207 8995
rect 2861 8888 2863 8896
rect 2877 8888 2879 8896
rect 2893 8888 2895 8896
rect 2916 8888 2918 8896
rect 2921 8888 2923 8896
rect 2947 8888 2949 8896
rect 2968 8888 2970 8896
rect 2988 8888 2990 8896
rect 2993 8888 2995 8896
rect 3011 8888 3013 8896
rect 3061 8887 3063 8895
rect 3066 8887 3068 8895
rect 3142 8887 3144 8895
rect 3147 8887 3149 8895
rect 3232 8887 3234 8895
rect 3237 8887 3239 8895
rect 3806 8888 3808 8896
rect 3822 8888 3824 8896
rect 3838 8888 3840 8896
rect 3861 8888 3863 8896
rect 3866 8888 3868 8896
rect 3892 8888 3894 8896
rect 3913 8888 3915 8896
rect 3933 8888 3935 8896
rect 3938 8888 3940 8896
rect 3956 8888 3958 8896
rect 4006 8887 4008 8895
rect 4011 8887 4013 8895
rect 4087 8887 4089 8895
rect 4092 8887 4094 8895
rect 4177 8887 4179 8895
rect 4182 8887 4184 8895
rect 2861 8842 2863 8850
rect 2877 8842 2879 8850
rect 2893 8842 2895 8850
rect 2916 8842 2918 8850
rect 2921 8842 2923 8850
rect 2947 8842 2949 8850
rect 2968 8842 2970 8850
rect 2988 8842 2990 8850
rect 2993 8842 2995 8850
rect 3011 8842 3013 8850
rect 3061 8849 3063 8857
rect 3066 8849 3068 8857
rect 3089 8855 3091 8863
rect 3397 8858 3399 8866
rect 3402 8858 3404 8866
rect 3806 8842 3808 8850
rect 3822 8842 3824 8850
rect 3838 8842 3840 8850
rect 3861 8842 3863 8850
rect 3866 8842 3868 8850
rect 3892 8842 3894 8850
rect 3913 8842 3915 8850
rect 3933 8842 3935 8850
rect 3938 8842 3940 8850
rect 3956 8842 3958 8850
rect 4006 8849 4008 8857
rect 4011 8849 4013 8857
rect 4034 8855 4036 8863
rect 2372 8787 2374 8795
rect 2377 8787 2379 8795
rect 2393 8787 2395 8795
rect 2409 8787 2411 8795
rect 2414 8787 2416 8795
rect 2435 8787 2437 8795
rect 2451 8787 2453 8795
rect 2467 8787 2469 8795
rect 2472 8787 2474 8795
rect 2488 8787 2490 8795
rect 2504 8787 2506 8795
rect 2509 8787 2511 8795
rect 2525 8787 2527 8795
rect 2541 8787 2543 8795
rect 2546 8787 2548 8795
rect 2567 8787 2569 8795
rect 2583 8787 2585 8795
rect 2599 8787 2601 8795
rect 2604 8787 2606 8795
rect 2620 8787 2622 8795
rect 2636 8787 2638 8795
rect 2641 8787 2643 8795
rect 2657 8787 2659 8795
rect 2673 8787 2675 8795
rect 2678 8787 2680 8795
rect 2699 8787 2701 8795
rect 2715 8787 2717 8795
rect 2731 8787 2733 8795
rect 2736 8787 2738 8795
rect 2752 8787 2754 8795
rect 3317 8787 3319 8795
rect 3322 8787 3324 8795
rect 3338 8787 3340 8795
rect 3354 8787 3356 8795
rect 3359 8787 3361 8795
rect 3380 8787 3382 8795
rect 3396 8787 3398 8795
rect 3412 8787 3414 8795
rect 3417 8787 3419 8795
rect 3433 8787 3435 8795
rect 3449 8787 3451 8795
rect 3454 8787 3456 8795
rect 3470 8787 3472 8795
rect 3486 8787 3488 8795
rect 3491 8787 3493 8795
rect 3512 8787 3514 8795
rect 3528 8787 3530 8795
rect 3544 8787 3546 8795
rect 3549 8787 3551 8795
rect 3565 8787 3567 8795
rect 3581 8787 3583 8795
rect 3586 8787 3588 8795
rect 3602 8787 3604 8795
rect 3618 8787 3620 8795
rect 3623 8787 3625 8795
rect 3644 8787 3646 8795
rect 3660 8787 3662 8795
rect 3676 8787 3678 8795
rect 3681 8787 3683 8795
rect 3697 8787 3699 8795
rect 2861 8756 2863 8764
rect 2877 8756 2879 8764
rect 2893 8756 2895 8764
rect 2916 8756 2918 8764
rect 2921 8756 2923 8764
rect 2947 8756 2949 8764
rect 2968 8756 2970 8764
rect 2988 8756 2990 8764
rect 2993 8756 2995 8764
rect 3011 8756 3013 8764
rect 3061 8751 3063 8759
rect 3066 8751 3068 8759
rect 3095 8756 3097 8764
rect 3113 8756 3115 8764
rect 3138 8756 3140 8764
rect 3154 8756 3156 8764
rect 3177 8756 3179 8764
rect 3182 8756 3184 8764
rect 3208 8756 3210 8764
rect 3229 8756 3231 8764
rect 3249 8756 3251 8764
rect 3254 8756 3256 8764
rect 3272 8756 3274 8764
rect 3806 8756 3808 8764
rect 3822 8756 3824 8764
rect 3838 8756 3840 8764
rect 3861 8756 3863 8764
rect 3866 8756 3868 8764
rect 3892 8756 3894 8764
rect 3913 8756 3915 8764
rect 3933 8756 3935 8764
rect 3938 8756 3940 8764
rect 3956 8756 3958 8764
rect 4006 8751 4008 8759
rect 4011 8751 4013 8759
rect 4040 8756 4042 8764
rect 4058 8756 4060 8764
rect 4083 8756 4085 8764
rect 4099 8756 4101 8764
rect 4122 8756 4124 8764
rect 4127 8756 4129 8764
rect 4153 8756 4155 8764
rect 4174 8756 4176 8764
rect 4194 8756 4196 8764
rect 4199 8756 4201 8764
rect 4217 8756 4219 8764
rect 3155 8675 3157 8683
rect 3160 8675 3162 8683
rect 3176 8675 3178 8683
rect 3192 8675 3194 8683
rect 3197 8675 3199 8683
rect 3218 8675 3220 8683
rect 3234 8675 3236 8683
rect 3250 8675 3252 8683
rect 3255 8675 3257 8683
rect 3271 8675 3273 8683
rect 4100 8675 4102 8683
rect 4105 8675 4107 8683
rect 4121 8675 4123 8683
rect 4137 8675 4139 8683
rect 4142 8675 4144 8683
rect 4163 8675 4165 8683
rect 4179 8675 4181 8683
rect 4195 8675 4197 8683
rect 4200 8675 4202 8683
rect 4216 8675 4218 8683
rect 2372 8645 2374 8653
rect 2377 8645 2379 8653
rect 2393 8645 2395 8653
rect 2409 8645 2411 8653
rect 2414 8645 2416 8653
rect 2435 8645 2437 8653
rect 2451 8645 2453 8653
rect 2467 8645 2469 8653
rect 2472 8645 2474 8653
rect 2488 8645 2490 8653
rect 2504 8645 2506 8653
rect 2509 8645 2511 8653
rect 2525 8645 2527 8653
rect 2541 8645 2543 8653
rect 2546 8645 2548 8653
rect 2567 8645 2569 8653
rect 2583 8645 2585 8653
rect 2599 8645 2601 8653
rect 2604 8645 2606 8653
rect 2620 8645 2622 8653
rect 2636 8645 2638 8653
rect 2641 8645 2643 8653
rect 2657 8645 2659 8653
rect 2673 8645 2675 8653
rect 2678 8645 2680 8653
rect 2699 8645 2701 8653
rect 2715 8645 2717 8653
rect 2731 8645 2733 8653
rect 2736 8645 2738 8653
rect 2752 8645 2754 8653
rect 3317 8645 3319 8653
rect 3322 8645 3324 8653
rect 3338 8645 3340 8653
rect 3354 8645 3356 8653
rect 3359 8645 3361 8653
rect 3380 8645 3382 8653
rect 3396 8645 3398 8653
rect 3412 8645 3414 8653
rect 3417 8645 3419 8653
rect 3433 8645 3435 8653
rect 3449 8645 3451 8653
rect 3454 8645 3456 8653
rect 3470 8645 3472 8653
rect 3486 8645 3488 8653
rect 3491 8645 3493 8653
rect 3512 8645 3514 8653
rect 3528 8645 3530 8653
rect 3544 8645 3546 8653
rect 3549 8645 3551 8653
rect 3565 8645 3567 8653
rect 3581 8645 3583 8653
rect 3586 8645 3588 8653
rect 3602 8645 3604 8653
rect 3618 8645 3620 8653
rect 3623 8645 3625 8653
rect 3644 8645 3646 8653
rect 3660 8645 3662 8653
rect 3676 8645 3678 8653
rect 3681 8645 3683 8653
rect 3697 8645 3699 8653
rect 3155 8589 3157 8597
rect 3160 8589 3162 8597
rect 3176 8589 3178 8597
rect 3192 8589 3194 8597
rect 3197 8589 3199 8597
rect 3218 8589 3220 8597
rect 3234 8589 3236 8597
rect 3250 8589 3252 8597
rect 3255 8589 3257 8597
rect 3271 8589 3273 8597
rect 4100 8589 4102 8597
rect 4105 8589 4107 8597
rect 4121 8589 4123 8597
rect 4137 8589 4139 8597
rect 4142 8589 4144 8597
rect 4163 8589 4165 8597
rect 4179 8589 4181 8597
rect 4195 8589 4197 8597
rect 4200 8589 4202 8597
rect 4216 8589 4218 8597
rect 2372 8559 2374 8567
rect 2377 8559 2379 8567
rect 2393 8559 2395 8567
rect 2409 8559 2411 8567
rect 2414 8559 2416 8567
rect 2435 8559 2437 8567
rect 2451 8559 2453 8567
rect 2467 8559 2469 8567
rect 2472 8559 2474 8567
rect 2488 8559 2490 8567
rect 2504 8559 2506 8567
rect 2509 8559 2511 8567
rect 2525 8559 2527 8567
rect 2541 8559 2543 8567
rect 2546 8559 2548 8567
rect 2567 8559 2569 8567
rect 2583 8559 2585 8567
rect 2599 8559 2601 8567
rect 2604 8559 2606 8567
rect 2620 8559 2622 8567
rect 2636 8559 2638 8567
rect 2641 8559 2643 8567
rect 2657 8559 2659 8567
rect 2673 8559 2675 8567
rect 2678 8559 2680 8567
rect 2699 8559 2701 8567
rect 2715 8559 2717 8567
rect 2731 8559 2733 8567
rect 2736 8559 2738 8567
rect 2752 8559 2754 8567
rect 3317 8559 3319 8567
rect 3322 8559 3324 8567
rect 3338 8559 3340 8567
rect 3354 8559 3356 8567
rect 3359 8559 3361 8567
rect 3380 8559 3382 8567
rect 3396 8559 3398 8567
rect 3412 8559 3414 8567
rect 3417 8559 3419 8567
rect 3433 8559 3435 8567
rect 3449 8559 3451 8567
rect 3454 8559 3456 8567
rect 3470 8559 3472 8567
rect 3486 8559 3488 8567
rect 3491 8559 3493 8567
rect 3512 8559 3514 8567
rect 3528 8559 3530 8567
rect 3544 8559 3546 8567
rect 3549 8559 3551 8567
rect 3565 8559 3567 8567
rect 3581 8559 3583 8567
rect 3586 8559 3588 8567
rect 3602 8559 3604 8567
rect 3618 8559 3620 8567
rect 3623 8559 3625 8567
rect 3644 8559 3646 8567
rect 3660 8559 3662 8567
rect 3676 8559 3678 8567
rect 3681 8559 3683 8567
rect 3697 8559 3699 8567
rect 2372 8419 2374 8427
rect 2377 8419 2379 8427
rect 2393 8419 2395 8427
rect 2409 8419 2411 8427
rect 2414 8419 2416 8427
rect 2435 8419 2437 8427
rect 2451 8419 2453 8427
rect 2467 8419 2469 8427
rect 2472 8419 2474 8427
rect 2488 8419 2490 8427
rect 2504 8419 2506 8427
rect 2509 8419 2511 8427
rect 2525 8419 2527 8427
rect 2541 8419 2543 8427
rect 2546 8419 2548 8427
rect 2567 8419 2569 8427
rect 2583 8419 2585 8427
rect 2599 8419 2601 8427
rect 2604 8419 2606 8427
rect 2620 8419 2622 8427
rect 2636 8419 2638 8427
rect 2641 8419 2643 8427
rect 2657 8419 2659 8427
rect 2673 8419 2675 8427
rect 2678 8419 2680 8427
rect 2699 8419 2701 8427
rect 2715 8419 2717 8427
rect 2731 8419 2733 8427
rect 2736 8419 2738 8427
rect 2752 8419 2754 8427
rect 3317 8419 3319 8427
rect 3322 8419 3324 8427
rect 3338 8419 3340 8427
rect 3354 8419 3356 8427
rect 3359 8419 3361 8427
rect 3380 8419 3382 8427
rect 3396 8419 3398 8427
rect 3412 8419 3414 8427
rect 3417 8419 3419 8427
rect 3433 8419 3435 8427
rect 3449 8419 3451 8427
rect 3454 8419 3456 8427
rect 3470 8419 3472 8427
rect 3486 8419 3488 8427
rect 3491 8419 3493 8427
rect 3512 8419 3514 8427
rect 3528 8419 3530 8427
rect 3544 8419 3546 8427
rect 3549 8419 3551 8427
rect 3565 8419 3567 8427
rect 3581 8419 3583 8427
rect 3586 8419 3588 8427
rect 3602 8419 3604 8427
rect 3618 8419 3620 8427
rect 3623 8419 3625 8427
rect 3644 8419 3646 8427
rect 3660 8419 3662 8427
rect 3676 8419 3678 8427
rect 3681 8419 3683 8427
rect 3697 8419 3699 8427
rect 2856 8340 2858 8348
rect 2861 8340 2863 8348
rect 2877 8340 2879 8348
rect 2893 8340 2895 8348
rect 2898 8340 2900 8348
rect 2919 8340 2921 8348
rect 2935 8340 2937 8348
rect 2951 8340 2953 8348
rect 2956 8340 2958 8348
rect 2972 8340 2974 8348
rect 2988 8340 2990 8348
rect 2993 8340 2995 8348
rect 3009 8340 3011 8348
rect 3025 8340 3027 8348
rect 3030 8340 3032 8348
rect 3051 8340 3053 8348
rect 3067 8340 3069 8348
rect 3083 8340 3085 8348
rect 3088 8340 3090 8348
rect 3104 8340 3106 8348
rect 3120 8340 3122 8348
rect 3125 8340 3127 8348
rect 3141 8340 3143 8348
rect 3157 8340 3159 8348
rect 3162 8340 3164 8348
rect 3183 8340 3185 8348
rect 3199 8340 3201 8348
rect 3215 8340 3217 8348
rect 3220 8340 3222 8348
rect 3236 8340 3238 8348
rect 3252 8340 3254 8348
rect 3257 8340 3259 8348
rect 3273 8340 3275 8348
rect 3289 8340 3291 8348
rect 3294 8340 3296 8348
rect 3315 8340 3317 8348
rect 3331 8340 3333 8348
rect 3347 8340 3349 8348
rect 3352 8340 3354 8348
rect 3368 8340 3370 8348
rect 3801 8340 3803 8348
rect 3806 8340 3808 8348
rect 3822 8340 3824 8348
rect 3838 8340 3840 8348
rect 3843 8340 3845 8348
rect 3864 8340 3866 8348
rect 3880 8340 3882 8348
rect 3896 8340 3898 8348
rect 3901 8340 3903 8348
rect 3917 8340 3919 8348
rect 3933 8340 3935 8348
rect 3938 8340 3940 8348
rect 3954 8340 3956 8348
rect 3970 8340 3972 8348
rect 3975 8340 3977 8348
rect 3996 8340 3998 8348
rect 4012 8340 4014 8348
rect 4028 8340 4030 8348
rect 4033 8340 4035 8348
rect 4049 8340 4051 8348
rect 4065 8340 4067 8348
rect 4070 8340 4072 8348
rect 4086 8340 4088 8348
rect 4102 8340 4104 8348
rect 4107 8340 4109 8348
rect 4128 8340 4130 8348
rect 4144 8340 4146 8348
rect 4160 8340 4162 8348
rect 4165 8340 4167 8348
rect 4181 8340 4183 8348
rect 4197 8340 4199 8348
rect 4202 8340 4204 8348
rect 4218 8340 4220 8348
rect 4234 8340 4236 8348
rect 4239 8340 4241 8348
rect 4260 8340 4262 8348
rect 4276 8340 4278 8348
rect 4292 8340 4294 8348
rect 4297 8340 4299 8348
rect 4313 8340 4315 8348
rect 2504 8307 2506 8315
rect 2509 8307 2511 8315
rect 2525 8307 2527 8315
rect 2541 8307 2543 8315
rect 2546 8307 2548 8315
rect 2567 8307 2569 8315
rect 2583 8307 2585 8315
rect 2599 8307 2601 8315
rect 2604 8307 2606 8315
rect 2620 8307 2622 8315
rect 3449 8307 3451 8315
rect 3454 8307 3456 8315
rect 3470 8307 3472 8315
rect 3486 8307 3488 8315
rect 3491 8307 3493 8315
rect 3512 8307 3514 8315
rect 3528 8307 3530 8315
rect 3544 8307 3546 8315
rect 3549 8307 3551 8315
rect 3565 8307 3567 8315
rect 3035 8269 3037 8277
rect 2861 8256 2863 8264
rect 2877 8256 2879 8264
rect 2893 8256 2895 8264
rect 2916 8256 2918 8264
rect 2921 8256 2923 8264
rect 2947 8256 2949 8264
rect 2968 8256 2970 8264
rect 2988 8256 2990 8264
rect 2993 8256 2995 8264
rect 3011 8256 3013 8264
rect 3061 8263 3063 8271
rect 3066 8263 3068 8271
rect 3089 8269 3091 8277
rect 3116 8269 3118 8277
rect 3142 8263 3144 8271
rect 3147 8263 3149 8271
rect 3170 8269 3172 8277
rect 3980 8269 3982 8277
rect 3806 8256 3808 8264
rect 3822 8256 3824 8264
rect 3838 8256 3840 8264
rect 3861 8256 3863 8264
rect 3866 8256 3868 8264
rect 3892 8256 3894 8264
rect 3913 8256 3915 8264
rect 3933 8256 3935 8264
rect 3938 8256 3940 8264
rect 3956 8256 3958 8264
rect 4006 8263 4008 8271
rect 4011 8263 4013 8271
rect 4034 8269 4036 8277
rect 4061 8269 4063 8277
rect 4087 8263 4089 8271
rect 4092 8263 4094 8271
rect 4115 8269 4117 8277
rect 2495 8205 2497 8213
rect 2511 8205 2513 8213
rect 2516 8205 2518 8213
rect 2532 8205 2534 8213
rect 2548 8205 2550 8213
rect 2569 8205 2571 8213
rect 2574 8205 2576 8213
rect 2590 8205 2592 8213
rect 2606 8205 2608 8213
rect 2611 8205 2613 8213
rect 3440 8205 3442 8213
rect 3456 8205 3458 8213
rect 3461 8205 3463 8213
rect 3477 8205 3479 8213
rect 3493 8205 3495 8213
rect 3514 8205 3516 8213
rect 3519 8205 3521 8213
rect 3535 8205 3537 8213
rect 3551 8205 3553 8213
rect 3556 8205 3558 8213
rect 2861 8170 2863 8178
rect 2877 8170 2879 8178
rect 2893 8170 2895 8178
rect 2916 8170 2918 8178
rect 2921 8170 2923 8178
rect 2947 8170 2949 8178
rect 2968 8170 2970 8178
rect 2988 8170 2990 8178
rect 2993 8170 2995 8178
rect 3011 8170 3013 8178
rect 3061 8171 3063 8179
rect 3066 8171 3068 8179
rect 3142 8171 3144 8179
rect 3147 8171 3149 8179
rect 3806 8170 3808 8178
rect 3822 8170 3824 8178
rect 3838 8170 3840 8178
rect 3861 8170 3863 8178
rect 3866 8170 3868 8178
rect 3892 8170 3894 8178
rect 3913 8170 3915 8178
rect 3933 8170 3935 8178
rect 3938 8170 3940 8178
rect 3956 8170 3958 8178
rect 4006 8171 4008 8179
rect 4011 8171 4013 8179
rect 4087 8171 4089 8179
rect 4092 8171 4094 8179
rect 2861 8124 2863 8132
rect 2877 8124 2879 8132
rect 2893 8124 2895 8132
rect 2916 8124 2918 8132
rect 2921 8124 2923 8132
rect 2947 8124 2949 8132
rect 2968 8124 2970 8132
rect 2988 8124 2990 8132
rect 2993 8124 2995 8132
rect 3011 8124 3013 8132
rect 3061 8131 3063 8139
rect 3066 8131 3068 8139
rect 3089 8137 3091 8145
rect 3140 8137 3142 8145
rect 3166 8131 3168 8139
rect 3171 8131 3173 8139
rect 3194 8137 3196 8145
rect 3806 8124 3808 8132
rect 3822 8124 3824 8132
rect 3838 8124 3840 8132
rect 3861 8124 3863 8132
rect 3866 8124 3868 8132
rect 3892 8124 3894 8132
rect 3913 8124 3915 8132
rect 3933 8124 3935 8132
rect 3938 8124 3940 8132
rect 3956 8124 3958 8132
rect 4006 8131 4008 8139
rect 4011 8131 4013 8139
rect 4034 8137 4036 8145
rect 4085 8137 4087 8145
rect 4111 8131 4113 8139
rect 4116 8131 4118 8139
rect 4139 8137 4141 8145
rect 2861 8038 2863 8046
rect 2877 8038 2879 8046
rect 2893 8038 2895 8046
rect 2916 8038 2918 8046
rect 2921 8038 2923 8046
rect 2947 8038 2949 8046
rect 2968 8038 2970 8046
rect 2988 8038 2990 8046
rect 2993 8038 2995 8046
rect 3011 8038 3013 8046
rect 3061 8040 3063 8048
rect 3066 8040 3068 8048
rect 3166 8040 3168 8048
rect 3171 8040 3173 8048
rect 3806 8038 3808 8046
rect 3822 8038 3824 8046
rect 3838 8038 3840 8046
rect 3861 8038 3863 8046
rect 3866 8038 3868 8046
rect 3892 8038 3894 8046
rect 3913 8038 3915 8046
rect 3933 8038 3935 8046
rect 3938 8038 3940 8046
rect 3956 8038 3958 8046
rect 4006 8040 4008 8048
rect 4011 8040 4013 8048
rect 4111 8040 4113 8048
rect 4116 8040 4118 8048
rect 2861 7992 2863 8000
rect 2877 7992 2879 8000
rect 2893 7992 2895 8000
rect 2916 7992 2918 8000
rect 2921 7992 2923 8000
rect 2947 7992 2949 8000
rect 2968 7992 2970 8000
rect 2988 7992 2990 8000
rect 2993 7992 2995 8000
rect 3011 7992 3013 8000
rect 3061 7999 3063 8007
rect 3066 7999 3068 8007
rect 3089 8005 3091 8013
rect 3116 8005 3118 8013
rect 3142 7999 3144 8007
rect 3147 7999 3149 8007
rect 3170 8005 3172 8013
rect 3206 8005 3208 8013
rect 3232 7999 3234 8007
rect 3237 7999 3239 8007
rect 3260 8005 3262 8013
rect 3806 7992 3808 8000
rect 3822 7992 3824 8000
rect 3838 7992 3840 8000
rect 3861 7992 3863 8000
rect 3866 7992 3868 8000
rect 3892 7992 3894 8000
rect 3913 7992 3915 8000
rect 3933 7992 3935 8000
rect 3938 7992 3940 8000
rect 3956 7992 3958 8000
rect 4006 7999 4008 8007
rect 4011 7999 4013 8007
rect 4034 8005 4036 8013
rect 4061 8005 4063 8013
rect 4087 7999 4089 8007
rect 4092 7999 4094 8007
rect 4115 8005 4117 8013
rect 4151 8005 4153 8013
rect 4177 7999 4179 8007
rect 4182 7999 4184 8007
rect 4205 8005 4207 8013
rect 2861 7906 2863 7914
rect 2877 7906 2879 7914
rect 2893 7906 2895 7914
rect 2916 7906 2918 7914
rect 2921 7906 2923 7914
rect 2947 7906 2949 7914
rect 2968 7906 2970 7914
rect 2988 7906 2990 7914
rect 2993 7906 2995 7914
rect 3011 7906 3013 7914
rect 3061 7905 3063 7913
rect 3066 7905 3068 7913
rect 3142 7905 3144 7913
rect 3147 7905 3149 7913
rect 3232 7905 3234 7913
rect 3237 7905 3239 7913
rect 3806 7906 3808 7914
rect 3822 7906 3824 7914
rect 3838 7906 3840 7914
rect 3861 7906 3863 7914
rect 3866 7906 3868 7914
rect 3892 7906 3894 7914
rect 3913 7906 3915 7914
rect 3933 7906 3935 7914
rect 3938 7906 3940 7914
rect 3956 7906 3958 7914
rect 4006 7905 4008 7913
rect 4011 7905 4013 7913
rect 4087 7905 4089 7913
rect 4092 7905 4094 7913
rect 4177 7905 4179 7913
rect 4182 7905 4184 7913
rect 2861 7860 2863 7868
rect 2877 7860 2879 7868
rect 2893 7860 2895 7868
rect 2916 7860 2918 7868
rect 2921 7860 2923 7868
rect 2947 7860 2949 7868
rect 2968 7860 2970 7868
rect 2988 7860 2990 7868
rect 2993 7860 2995 7868
rect 3011 7860 3013 7868
rect 3061 7867 3063 7875
rect 3066 7867 3068 7875
rect 3089 7873 3091 7881
rect 3806 7860 3808 7868
rect 3822 7860 3824 7868
rect 3838 7860 3840 7868
rect 3861 7860 3863 7868
rect 3866 7860 3868 7868
rect 3892 7860 3894 7868
rect 3913 7860 3915 7868
rect 3933 7860 3935 7868
rect 3938 7860 3940 7868
rect 3956 7860 3958 7868
rect 4006 7867 4008 7875
rect 4011 7867 4013 7875
rect 4034 7873 4036 7881
rect 2372 7805 2374 7813
rect 2377 7805 2379 7813
rect 2393 7805 2395 7813
rect 2409 7805 2411 7813
rect 2414 7805 2416 7813
rect 2435 7805 2437 7813
rect 2451 7805 2453 7813
rect 2467 7805 2469 7813
rect 2472 7805 2474 7813
rect 2488 7805 2490 7813
rect 2504 7805 2506 7813
rect 2509 7805 2511 7813
rect 2525 7805 2527 7813
rect 2541 7805 2543 7813
rect 2546 7805 2548 7813
rect 2567 7805 2569 7813
rect 2583 7805 2585 7813
rect 2599 7805 2601 7813
rect 2604 7805 2606 7813
rect 2620 7805 2622 7813
rect 2636 7805 2638 7813
rect 2641 7805 2643 7813
rect 2657 7805 2659 7813
rect 2673 7805 2675 7813
rect 2678 7805 2680 7813
rect 2699 7805 2701 7813
rect 2715 7805 2717 7813
rect 2731 7805 2733 7813
rect 2736 7805 2738 7813
rect 2752 7805 2754 7813
rect 3317 7805 3319 7813
rect 3322 7805 3324 7813
rect 3338 7805 3340 7813
rect 3354 7805 3356 7813
rect 3359 7805 3361 7813
rect 3380 7805 3382 7813
rect 3396 7805 3398 7813
rect 3412 7805 3414 7813
rect 3417 7805 3419 7813
rect 3433 7805 3435 7813
rect 3449 7805 3451 7813
rect 3454 7805 3456 7813
rect 3470 7805 3472 7813
rect 3486 7805 3488 7813
rect 3491 7805 3493 7813
rect 3512 7805 3514 7813
rect 3528 7805 3530 7813
rect 3544 7805 3546 7813
rect 3549 7805 3551 7813
rect 3565 7805 3567 7813
rect 3581 7805 3583 7813
rect 3586 7805 3588 7813
rect 3602 7805 3604 7813
rect 3618 7805 3620 7813
rect 3623 7805 3625 7813
rect 3644 7805 3646 7813
rect 3660 7805 3662 7813
rect 3676 7805 3678 7813
rect 3681 7805 3683 7813
rect 3697 7805 3699 7813
rect 2861 7774 2863 7782
rect 2877 7774 2879 7782
rect 2893 7774 2895 7782
rect 2916 7774 2918 7782
rect 2921 7774 2923 7782
rect 2947 7774 2949 7782
rect 2968 7774 2970 7782
rect 2988 7774 2990 7782
rect 2993 7774 2995 7782
rect 3011 7774 3013 7782
rect 3061 7769 3063 7777
rect 3066 7769 3068 7777
rect 3095 7774 3097 7782
rect 3113 7774 3115 7782
rect 3138 7774 3140 7782
rect 3154 7774 3156 7782
rect 3177 7774 3179 7782
rect 3182 7774 3184 7782
rect 3208 7774 3210 7782
rect 3229 7774 3231 7782
rect 3249 7774 3251 7782
rect 3254 7774 3256 7782
rect 3272 7774 3274 7782
rect 3806 7774 3808 7782
rect 3822 7774 3824 7782
rect 3838 7774 3840 7782
rect 3861 7774 3863 7782
rect 3866 7774 3868 7782
rect 3892 7774 3894 7782
rect 3913 7774 3915 7782
rect 3933 7774 3935 7782
rect 3938 7774 3940 7782
rect 3956 7774 3958 7782
rect 4006 7769 4008 7777
rect 4011 7769 4013 7777
rect 4040 7774 4042 7782
rect 4058 7774 4060 7782
rect 4083 7774 4085 7782
rect 4099 7774 4101 7782
rect 4122 7774 4124 7782
rect 4127 7774 4129 7782
rect 4153 7774 4155 7782
rect 4174 7774 4176 7782
rect 4194 7774 4196 7782
rect 4199 7774 4201 7782
rect 4217 7774 4219 7782
rect 3155 7693 3157 7701
rect 3160 7693 3162 7701
rect 3176 7693 3178 7701
rect 3192 7693 3194 7701
rect 3197 7693 3199 7701
rect 3218 7693 3220 7701
rect 3234 7693 3236 7701
rect 3250 7693 3252 7701
rect 3255 7693 3257 7701
rect 3271 7693 3273 7701
rect 4100 7693 4102 7701
rect 4105 7693 4107 7701
rect 4121 7693 4123 7701
rect 4137 7693 4139 7701
rect 4142 7693 4144 7701
rect 4163 7693 4165 7701
rect 4179 7693 4181 7701
rect 4195 7693 4197 7701
rect 4200 7693 4202 7701
rect 4216 7693 4218 7701
rect 2372 7663 2374 7671
rect 2377 7663 2379 7671
rect 2393 7663 2395 7671
rect 2409 7663 2411 7671
rect 2414 7663 2416 7671
rect 2435 7663 2437 7671
rect 2451 7663 2453 7671
rect 2467 7663 2469 7671
rect 2472 7663 2474 7671
rect 2488 7663 2490 7671
rect 2504 7663 2506 7671
rect 2509 7663 2511 7671
rect 2525 7663 2527 7671
rect 2541 7663 2543 7671
rect 2546 7663 2548 7671
rect 2567 7663 2569 7671
rect 2583 7663 2585 7671
rect 2599 7663 2601 7671
rect 2604 7663 2606 7671
rect 2620 7663 2622 7671
rect 2636 7663 2638 7671
rect 2641 7663 2643 7671
rect 2657 7663 2659 7671
rect 2673 7663 2675 7671
rect 2678 7663 2680 7671
rect 2699 7663 2701 7671
rect 2715 7663 2717 7671
rect 2731 7663 2733 7671
rect 2736 7663 2738 7671
rect 2752 7663 2754 7671
rect 3317 7663 3319 7671
rect 3322 7663 3324 7671
rect 3338 7663 3340 7671
rect 3354 7663 3356 7671
rect 3359 7663 3361 7671
rect 3380 7663 3382 7671
rect 3396 7663 3398 7671
rect 3412 7663 3414 7671
rect 3417 7663 3419 7671
rect 3433 7663 3435 7671
rect 3449 7663 3451 7671
rect 3454 7663 3456 7671
rect 3470 7663 3472 7671
rect 3486 7663 3488 7671
rect 3491 7663 3493 7671
rect 3512 7663 3514 7671
rect 3528 7663 3530 7671
rect 3544 7663 3546 7671
rect 3549 7663 3551 7671
rect 3565 7663 3567 7671
rect 3581 7663 3583 7671
rect 3586 7663 3588 7671
rect 3602 7663 3604 7671
rect 3618 7663 3620 7671
rect 3623 7663 3625 7671
rect 3644 7663 3646 7671
rect 3660 7663 3662 7671
rect 3676 7663 3678 7671
rect 3681 7663 3683 7671
rect 3697 7663 3699 7671
rect 3155 7607 3157 7615
rect 3160 7607 3162 7615
rect 3176 7607 3178 7615
rect 3192 7607 3194 7615
rect 3197 7607 3199 7615
rect 3218 7607 3220 7615
rect 3234 7607 3236 7615
rect 3250 7607 3252 7615
rect 3255 7607 3257 7615
rect 3271 7607 3273 7615
rect 4100 7607 4102 7615
rect 4105 7607 4107 7615
rect 4121 7607 4123 7615
rect 4137 7607 4139 7615
rect 4142 7607 4144 7615
rect 4163 7607 4165 7615
rect 4179 7607 4181 7615
rect 4195 7607 4197 7615
rect 4200 7607 4202 7615
rect 4216 7607 4218 7615
rect 2372 7577 2374 7585
rect 2377 7577 2379 7585
rect 2393 7577 2395 7585
rect 2409 7577 2411 7585
rect 2414 7577 2416 7585
rect 2435 7577 2437 7585
rect 2451 7577 2453 7585
rect 2467 7577 2469 7585
rect 2472 7577 2474 7585
rect 2488 7577 2490 7585
rect 2504 7577 2506 7585
rect 2509 7577 2511 7585
rect 2525 7577 2527 7585
rect 2541 7577 2543 7585
rect 2546 7577 2548 7585
rect 2567 7577 2569 7585
rect 2583 7577 2585 7585
rect 2599 7577 2601 7585
rect 2604 7577 2606 7585
rect 2620 7577 2622 7585
rect 2636 7577 2638 7585
rect 2641 7577 2643 7585
rect 2657 7577 2659 7585
rect 2673 7577 2675 7585
rect 2678 7577 2680 7585
rect 2699 7577 2701 7585
rect 2715 7577 2717 7585
rect 2731 7577 2733 7585
rect 2736 7577 2738 7585
rect 2752 7577 2754 7585
rect 3317 7577 3319 7585
rect 3322 7577 3324 7585
rect 3338 7577 3340 7585
rect 3354 7577 3356 7585
rect 3359 7577 3361 7585
rect 3380 7577 3382 7585
rect 3396 7577 3398 7585
rect 3412 7577 3414 7585
rect 3417 7577 3419 7585
rect 3433 7577 3435 7585
rect 3449 7577 3451 7585
rect 3454 7577 3456 7585
rect 3470 7577 3472 7585
rect 3486 7577 3488 7585
rect 3491 7577 3493 7585
rect 3512 7577 3514 7585
rect 3528 7577 3530 7585
rect 3544 7577 3546 7585
rect 3549 7577 3551 7585
rect 3565 7577 3567 7585
rect 3581 7577 3583 7585
rect 3586 7577 3588 7585
rect 3602 7577 3604 7585
rect 3618 7577 3620 7585
rect 3623 7577 3625 7585
rect 3644 7577 3646 7585
rect 3660 7577 3662 7585
rect 3676 7577 3678 7585
rect 3681 7577 3683 7585
rect 3697 7577 3699 7585
rect 2372 7437 2374 7445
rect 2377 7437 2379 7445
rect 2393 7437 2395 7445
rect 2409 7437 2411 7445
rect 2414 7437 2416 7445
rect 2435 7437 2437 7445
rect 2451 7437 2453 7445
rect 2467 7437 2469 7445
rect 2472 7437 2474 7445
rect 2488 7437 2490 7445
rect 2504 7437 2506 7445
rect 2509 7437 2511 7445
rect 2525 7437 2527 7445
rect 2541 7437 2543 7445
rect 2546 7437 2548 7445
rect 2567 7437 2569 7445
rect 2583 7437 2585 7445
rect 2599 7437 2601 7445
rect 2604 7437 2606 7445
rect 2620 7437 2622 7445
rect 2636 7437 2638 7445
rect 2641 7437 2643 7445
rect 2657 7437 2659 7445
rect 2673 7437 2675 7445
rect 2678 7437 2680 7445
rect 2699 7437 2701 7445
rect 2715 7437 2717 7445
rect 2731 7437 2733 7445
rect 2736 7437 2738 7445
rect 2752 7437 2754 7445
rect 3317 7437 3319 7445
rect 3322 7437 3324 7445
rect 3338 7437 3340 7445
rect 3354 7437 3356 7445
rect 3359 7437 3361 7445
rect 3380 7437 3382 7445
rect 3396 7437 3398 7445
rect 3412 7437 3414 7445
rect 3417 7437 3419 7445
rect 3433 7437 3435 7445
rect 3449 7437 3451 7445
rect 3454 7437 3456 7445
rect 3470 7437 3472 7445
rect 3486 7437 3488 7445
rect 3491 7437 3493 7445
rect 3512 7437 3514 7445
rect 3528 7437 3530 7445
rect 3544 7437 3546 7445
rect 3549 7437 3551 7445
rect 3565 7437 3567 7445
rect 3581 7437 3583 7445
rect 3586 7437 3588 7445
rect 3602 7437 3604 7445
rect 3618 7437 3620 7445
rect 3623 7437 3625 7445
rect 3644 7437 3646 7445
rect 3660 7437 3662 7445
rect 3676 7437 3678 7445
rect 3681 7437 3683 7445
rect 3697 7437 3699 7445
rect 1473 6869 1475 6877
rect 1489 6869 1491 6877
rect 1494 6869 1496 6877
rect 1510 6869 1512 6877
rect 1526 6869 1528 6877
rect 1547 6869 1549 6877
rect 1552 6869 1554 6877
rect 1568 6869 1570 6877
rect 1584 6869 1586 6877
rect 1589 6869 1591 6877
rect 1605 6869 1607 6877
rect 1621 6869 1623 6877
rect 1626 6869 1628 6877
rect 1642 6869 1644 6877
rect 1658 6869 1660 6877
rect 1679 6869 1681 6877
rect 1684 6869 1686 6877
rect 1700 6869 1702 6877
rect 1716 6869 1718 6877
rect 1721 6869 1723 6877
rect 1737 6869 1739 6877
rect 1753 6869 1755 6877
rect 1758 6869 1760 6877
rect 1774 6869 1776 6877
rect 1790 6869 1792 6877
rect 1811 6869 1813 6877
rect 1816 6869 1818 6877
rect 1832 6869 1834 6877
rect 1848 6869 1850 6877
rect 1853 6869 1855 6877
rect 2418 6869 2420 6877
rect 2434 6869 2436 6877
rect 2439 6869 2441 6877
rect 2455 6869 2457 6877
rect 2471 6869 2473 6877
rect 2492 6869 2494 6877
rect 2497 6869 2499 6877
rect 2513 6869 2515 6877
rect 2529 6869 2531 6877
rect 2534 6869 2536 6877
rect 2550 6869 2552 6877
rect 2566 6869 2568 6877
rect 2571 6869 2573 6877
rect 2587 6869 2589 6877
rect 2603 6869 2605 6877
rect 2624 6869 2626 6877
rect 2629 6869 2631 6877
rect 2645 6869 2647 6877
rect 2661 6869 2663 6877
rect 2666 6869 2668 6877
rect 2682 6869 2684 6877
rect 2698 6869 2700 6877
rect 2703 6869 2705 6877
rect 2719 6869 2721 6877
rect 2735 6869 2737 6877
rect 2756 6869 2758 6877
rect 2761 6869 2763 6877
rect 2777 6869 2779 6877
rect 2793 6869 2795 6877
rect 2798 6869 2800 6877
rect 1473 6729 1475 6737
rect 1489 6729 1491 6737
rect 1494 6729 1496 6737
rect 1510 6729 1512 6737
rect 1526 6729 1528 6737
rect 1547 6729 1549 6737
rect 1552 6729 1554 6737
rect 1568 6729 1570 6737
rect 1584 6729 1586 6737
rect 1589 6729 1591 6737
rect 1605 6729 1607 6737
rect 1621 6729 1623 6737
rect 1626 6729 1628 6737
rect 1642 6729 1644 6737
rect 1658 6729 1660 6737
rect 1679 6729 1681 6737
rect 1684 6729 1686 6737
rect 1700 6729 1702 6737
rect 1716 6729 1718 6737
rect 1721 6729 1723 6737
rect 1737 6729 1739 6737
rect 1753 6729 1755 6737
rect 1758 6729 1760 6737
rect 1774 6729 1776 6737
rect 1790 6729 1792 6737
rect 1811 6729 1813 6737
rect 1816 6729 1818 6737
rect 1832 6729 1834 6737
rect 1848 6729 1850 6737
rect 1853 6729 1855 6737
rect 2418 6729 2420 6737
rect 2434 6729 2436 6737
rect 2439 6729 2441 6737
rect 2455 6729 2457 6737
rect 2471 6729 2473 6737
rect 2492 6729 2494 6737
rect 2497 6729 2499 6737
rect 2513 6729 2515 6737
rect 2529 6729 2531 6737
rect 2534 6729 2536 6737
rect 2550 6729 2552 6737
rect 2566 6729 2568 6737
rect 2571 6729 2573 6737
rect 2587 6729 2589 6737
rect 2603 6729 2605 6737
rect 2624 6729 2626 6737
rect 2629 6729 2631 6737
rect 2645 6729 2647 6737
rect 2661 6729 2663 6737
rect 2666 6729 2668 6737
rect 2682 6729 2684 6737
rect 2698 6729 2700 6737
rect 2703 6729 2705 6737
rect 2719 6729 2721 6737
rect 2735 6729 2737 6737
rect 2756 6729 2758 6737
rect 2761 6729 2763 6737
rect 2777 6729 2779 6737
rect 2793 6729 2795 6737
rect 2798 6729 2800 6737
rect 954 6699 956 6707
rect 970 6699 972 6707
rect 975 6699 977 6707
rect 991 6699 993 6707
rect 1007 6699 1009 6707
rect 1028 6699 1030 6707
rect 1033 6699 1035 6707
rect 1049 6699 1051 6707
rect 1065 6699 1067 6707
rect 1070 6699 1072 6707
rect 1899 6699 1901 6707
rect 1915 6699 1917 6707
rect 1920 6699 1922 6707
rect 1936 6699 1938 6707
rect 1952 6699 1954 6707
rect 1973 6699 1975 6707
rect 1978 6699 1980 6707
rect 1994 6699 1996 6707
rect 2010 6699 2012 6707
rect 2015 6699 2017 6707
rect 1473 6643 1475 6651
rect 1489 6643 1491 6651
rect 1494 6643 1496 6651
rect 1510 6643 1512 6651
rect 1526 6643 1528 6651
rect 1547 6643 1549 6651
rect 1552 6643 1554 6651
rect 1568 6643 1570 6651
rect 1584 6643 1586 6651
rect 1589 6643 1591 6651
rect 1605 6643 1607 6651
rect 1621 6643 1623 6651
rect 1626 6643 1628 6651
rect 1642 6643 1644 6651
rect 1658 6643 1660 6651
rect 1679 6643 1681 6651
rect 1684 6643 1686 6651
rect 1700 6643 1702 6651
rect 1716 6643 1718 6651
rect 1721 6643 1723 6651
rect 1737 6643 1739 6651
rect 1753 6643 1755 6651
rect 1758 6643 1760 6651
rect 1774 6643 1776 6651
rect 1790 6643 1792 6651
rect 1811 6643 1813 6651
rect 1816 6643 1818 6651
rect 1832 6643 1834 6651
rect 1848 6643 1850 6651
rect 1853 6643 1855 6651
rect 2418 6643 2420 6651
rect 2434 6643 2436 6651
rect 2439 6643 2441 6651
rect 2455 6643 2457 6651
rect 2471 6643 2473 6651
rect 2492 6643 2494 6651
rect 2497 6643 2499 6651
rect 2513 6643 2515 6651
rect 2529 6643 2531 6651
rect 2534 6643 2536 6651
rect 2550 6643 2552 6651
rect 2566 6643 2568 6651
rect 2571 6643 2573 6651
rect 2587 6643 2589 6651
rect 2603 6643 2605 6651
rect 2624 6643 2626 6651
rect 2629 6643 2631 6651
rect 2645 6643 2647 6651
rect 2661 6643 2663 6651
rect 2666 6643 2668 6651
rect 2682 6643 2684 6651
rect 2698 6643 2700 6651
rect 2703 6643 2705 6651
rect 2719 6643 2721 6651
rect 2735 6643 2737 6651
rect 2756 6643 2758 6651
rect 2761 6643 2763 6651
rect 2777 6643 2779 6651
rect 2793 6643 2795 6651
rect 2798 6643 2800 6651
rect 954 6613 956 6621
rect 970 6613 972 6621
rect 975 6613 977 6621
rect 991 6613 993 6621
rect 1007 6613 1009 6621
rect 1028 6613 1030 6621
rect 1033 6613 1035 6621
rect 1049 6613 1051 6621
rect 1065 6613 1067 6621
rect 1070 6613 1072 6621
rect 1899 6613 1901 6621
rect 1915 6613 1917 6621
rect 1920 6613 1922 6621
rect 1936 6613 1938 6621
rect 1952 6613 1954 6621
rect 1973 6613 1975 6621
rect 1978 6613 1980 6621
rect 1994 6613 1996 6621
rect 2010 6613 2012 6621
rect 2015 6613 2017 6621
rect 953 6532 955 6540
rect 971 6532 973 6540
rect 976 6532 978 6540
rect 996 6532 998 6540
rect 1017 6532 1019 6540
rect 1043 6532 1045 6540
rect 1048 6532 1050 6540
rect 1071 6532 1073 6540
rect 1087 6532 1089 6540
rect 1112 6532 1114 6540
rect 1130 6532 1132 6540
rect 1159 6537 1161 6545
rect 1164 6537 1166 6545
rect 1214 6532 1216 6540
rect 1232 6532 1234 6540
rect 1237 6532 1239 6540
rect 1257 6532 1259 6540
rect 1278 6532 1280 6540
rect 1304 6532 1306 6540
rect 1309 6532 1311 6540
rect 1332 6532 1334 6540
rect 1348 6532 1350 6540
rect 1364 6532 1366 6540
rect 1898 6532 1900 6540
rect 1916 6532 1918 6540
rect 1921 6532 1923 6540
rect 1941 6532 1943 6540
rect 1962 6532 1964 6540
rect 1988 6532 1990 6540
rect 1993 6532 1995 6540
rect 2016 6532 2018 6540
rect 2032 6532 2034 6540
rect 2057 6532 2059 6540
rect 2075 6532 2077 6540
rect 2104 6537 2106 6545
rect 2109 6537 2111 6545
rect 2159 6532 2161 6540
rect 2177 6532 2179 6540
rect 2182 6532 2184 6540
rect 2202 6532 2204 6540
rect 2223 6532 2225 6540
rect 2249 6532 2251 6540
rect 2254 6532 2256 6540
rect 2277 6532 2279 6540
rect 2293 6532 2295 6540
rect 2309 6532 2311 6540
rect 1473 6501 1475 6509
rect 1489 6501 1491 6509
rect 1494 6501 1496 6509
rect 1510 6501 1512 6509
rect 1526 6501 1528 6509
rect 1547 6501 1549 6509
rect 1552 6501 1554 6509
rect 1568 6501 1570 6509
rect 1584 6501 1586 6509
rect 1589 6501 1591 6509
rect 1605 6501 1607 6509
rect 1621 6501 1623 6509
rect 1626 6501 1628 6509
rect 1642 6501 1644 6509
rect 1658 6501 1660 6509
rect 1679 6501 1681 6509
rect 1684 6501 1686 6509
rect 1700 6501 1702 6509
rect 1716 6501 1718 6509
rect 1721 6501 1723 6509
rect 1737 6501 1739 6509
rect 1753 6501 1755 6509
rect 1758 6501 1760 6509
rect 1774 6501 1776 6509
rect 1790 6501 1792 6509
rect 1811 6501 1813 6509
rect 1816 6501 1818 6509
rect 1832 6501 1834 6509
rect 1848 6501 1850 6509
rect 1853 6501 1855 6509
rect 2418 6501 2420 6509
rect 2434 6501 2436 6509
rect 2439 6501 2441 6509
rect 2455 6501 2457 6509
rect 2471 6501 2473 6509
rect 2492 6501 2494 6509
rect 2497 6501 2499 6509
rect 2513 6501 2515 6509
rect 2529 6501 2531 6509
rect 2534 6501 2536 6509
rect 2550 6501 2552 6509
rect 2566 6501 2568 6509
rect 2571 6501 2573 6509
rect 2587 6501 2589 6509
rect 2603 6501 2605 6509
rect 2624 6501 2626 6509
rect 2629 6501 2631 6509
rect 2645 6501 2647 6509
rect 2661 6501 2663 6509
rect 2666 6501 2668 6509
rect 2682 6501 2684 6509
rect 2698 6501 2700 6509
rect 2703 6501 2705 6509
rect 2719 6501 2721 6509
rect 2735 6501 2737 6509
rect 2756 6501 2758 6509
rect 2761 6501 2763 6509
rect 2777 6501 2779 6509
rect 2793 6501 2795 6509
rect 2798 6501 2800 6509
rect 1136 6433 1138 6441
rect 1159 6439 1161 6447
rect 1164 6439 1166 6447
rect 1214 6446 1216 6454
rect 1232 6446 1234 6454
rect 1237 6446 1239 6454
rect 1257 6446 1259 6454
rect 1278 6446 1280 6454
rect 1304 6446 1306 6454
rect 1309 6446 1311 6454
rect 1332 6446 1334 6454
rect 1348 6446 1350 6454
rect 1364 6446 1366 6454
rect 2081 6433 2083 6441
rect 2104 6439 2106 6447
rect 2109 6439 2111 6447
rect 2159 6446 2161 6454
rect 2177 6446 2179 6454
rect 2182 6446 2184 6454
rect 2202 6446 2204 6454
rect 2223 6446 2225 6454
rect 2249 6446 2251 6454
rect 2254 6446 2256 6454
rect 2277 6446 2279 6454
rect 2293 6446 2295 6454
rect 2309 6446 2311 6454
rect 988 6401 990 6409
rect 993 6401 995 6409
rect 1078 6401 1080 6409
rect 1083 6401 1085 6409
rect 1159 6401 1161 6409
rect 1164 6401 1166 6409
rect 1214 6400 1216 6408
rect 1232 6400 1234 6408
rect 1237 6400 1239 6408
rect 1257 6400 1259 6408
rect 1278 6400 1280 6408
rect 1304 6400 1306 6408
rect 1309 6400 1311 6408
rect 1332 6400 1334 6408
rect 1348 6400 1350 6408
rect 1364 6400 1366 6408
rect 1933 6401 1935 6409
rect 1938 6401 1940 6409
rect 2023 6401 2025 6409
rect 2028 6401 2030 6409
rect 2104 6401 2106 6409
rect 2109 6401 2111 6409
rect 2159 6400 2161 6408
rect 2177 6400 2179 6408
rect 2182 6400 2184 6408
rect 2202 6400 2204 6408
rect 2223 6400 2225 6408
rect 2249 6400 2251 6408
rect 2254 6400 2256 6408
rect 2277 6400 2279 6408
rect 2293 6400 2295 6408
rect 2309 6400 2311 6408
rect 965 6301 967 6309
rect 988 6307 990 6315
rect 993 6307 995 6315
rect 1019 6301 1021 6309
rect 1055 6301 1057 6309
rect 1078 6307 1080 6315
rect 1083 6307 1085 6315
rect 1109 6301 1111 6309
rect 1136 6301 1138 6309
rect 1159 6307 1161 6315
rect 1164 6307 1166 6315
rect 1214 6314 1216 6322
rect 1232 6314 1234 6322
rect 1237 6314 1239 6322
rect 1257 6314 1259 6322
rect 1278 6314 1280 6322
rect 1304 6314 1306 6322
rect 1309 6314 1311 6322
rect 1332 6314 1334 6322
rect 1348 6314 1350 6322
rect 1364 6314 1366 6322
rect 1910 6301 1912 6309
rect 1933 6307 1935 6315
rect 1938 6307 1940 6315
rect 1964 6301 1966 6309
rect 2000 6301 2002 6309
rect 2023 6307 2025 6315
rect 2028 6307 2030 6315
rect 2054 6301 2056 6309
rect 2081 6301 2083 6309
rect 2104 6307 2106 6315
rect 2109 6307 2111 6315
rect 2159 6314 2161 6322
rect 2177 6314 2179 6322
rect 2182 6314 2184 6322
rect 2202 6314 2204 6322
rect 2223 6314 2225 6322
rect 2249 6314 2251 6322
rect 2254 6314 2256 6322
rect 2277 6314 2279 6322
rect 2293 6314 2295 6322
rect 2309 6314 2311 6322
rect 1054 6266 1056 6274
rect 1059 6266 1061 6274
rect 1159 6266 1161 6274
rect 1164 6266 1166 6274
rect 1214 6268 1216 6276
rect 1232 6268 1234 6276
rect 1237 6268 1239 6276
rect 1257 6268 1259 6276
rect 1278 6268 1280 6276
rect 1304 6268 1306 6276
rect 1309 6268 1311 6276
rect 1332 6268 1334 6276
rect 1348 6268 1350 6276
rect 1364 6268 1366 6276
rect 1999 6266 2001 6274
rect 2004 6266 2006 6274
rect 2104 6266 2106 6274
rect 2109 6266 2111 6274
rect 2159 6268 2161 6276
rect 2177 6268 2179 6276
rect 2182 6268 2184 6276
rect 2202 6268 2204 6276
rect 2223 6268 2225 6276
rect 2249 6268 2251 6276
rect 2254 6268 2256 6276
rect 2277 6268 2279 6276
rect 2293 6268 2295 6276
rect 2309 6268 2311 6276
rect 1031 6169 1033 6177
rect 1054 6175 1056 6183
rect 1059 6175 1061 6183
rect 1085 6169 1087 6177
rect 1136 6169 1138 6177
rect 1159 6175 1161 6183
rect 1164 6175 1166 6183
rect 1214 6182 1216 6190
rect 1232 6182 1234 6190
rect 1237 6182 1239 6190
rect 1257 6182 1259 6190
rect 1278 6182 1280 6190
rect 1304 6182 1306 6190
rect 1309 6182 1311 6190
rect 1332 6182 1334 6190
rect 1348 6182 1350 6190
rect 1364 6182 1366 6190
rect 1976 6169 1978 6177
rect 1999 6175 2001 6183
rect 2004 6175 2006 6183
rect 2030 6169 2032 6177
rect 2081 6169 2083 6177
rect 2104 6175 2106 6183
rect 2109 6175 2111 6183
rect 2159 6182 2161 6190
rect 2177 6182 2179 6190
rect 2182 6182 2184 6190
rect 2202 6182 2204 6190
rect 2223 6182 2225 6190
rect 2249 6182 2251 6190
rect 2254 6182 2256 6190
rect 2277 6182 2279 6190
rect 2293 6182 2295 6190
rect 2309 6182 2311 6190
rect 1078 6135 1080 6143
rect 1083 6135 1085 6143
rect 1159 6135 1161 6143
rect 1164 6135 1166 6143
rect 1214 6136 1216 6144
rect 1232 6136 1234 6144
rect 1237 6136 1239 6144
rect 1257 6136 1259 6144
rect 1278 6136 1280 6144
rect 1304 6136 1306 6144
rect 1309 6136 1311 6144
rect 1332 6136 1334 6144
rect 1348 6136 1350 6144
rect 1364 6136 1366 6144
rect 2023 6135 2025 6143
rect 2028 6135 2030 6143
rect 2104 6135 2106 6143
rect 2109 6135 2111 6143
rect 2159 6136 2161 6144
rect 2177 6136 2179 6144
rect 2182 6136 2184 6144
rect 2202 6136 2204 6144
rect 2223 6136 2225 6144
rect 2249 6136 2251 6144
rect 2254 6136 2256 6144
rect 2277 6136 2279 6144
rect 2293 6136 2295 6144
rect 2309 6136 2311 6144
rect 1614 6101 1616 6109
rect 1619 6101 1621 6109
rect 1635 6101 1637 6109
rect 1651 6101 1653 6109
rect 1656 6101 1658 6109
rect 1677 6101 1679 6109
rect 1693 6101 1695 6109
rect 1709 6101 1711 6109
rect 1714 6101 1716 6109
rect 1730 6101 1732 6109
rect 2559 6101 2561 6109
rect 2564 6101 2566 6109
rect 2580 6101 2582 6109
rect 2596 6101 2598 6109
rect 2601 6101 2603 6109
rect 2622 6101 2624 6109
rect 2638 6101 2640 6109
rect 2654 6101 2656 6109
rect 2659 6101 2661 6109
rect 2675 6101 2677 6109
rect 1055 6037 1057 6045
rect 1078 6043 1080 6051
rect 1083 6043 1085 6051
rect 1109 6037 1111 6045
rect 1136 6037 1138 6045
rect 1159 6043 1161 6051
rect 1164 6043 1166 6051
rect 1214 6050 1216 6058
rect 1232 6050 1234 6058
rect 1237 6050 1239 6058
rect 1257 6050 1259 6058
rect 1278 6050 1280 6058
rect 1304 6050 1306 6058
rect 1309 6050 1311 6058
rect 1332 6050 1334 6058
rect 1348 6050 1350 6058
rect 1364 6050 1366 6058
rect 1190 6037 1192 6045
rect 2000 6037 2002 6045
rect 2023 6043 2025 6051
rect 2028 6043 2030 6051
rect 2054 6037 2056 6045
rect 2081 6037 2083 6045
rect 2104 6043 2106 6051
rect 2109 6043 2111 6051
rect 2159 6050 2161 6058
rect 2177 6050 2179 6058
rect 2182 6050 2184 6058
rect 2202 6050 2204 6058
rect 2223 6050 2225 6058
rect 2249 6050 2251 6058
rect 2254 6050 2256 6058
rect 2277 6050 2279 6058
rect 2293 6050 2295 6058
rect 2309 6050 2311 6058
rect 2135 6037 2137 6045
rect 1605 5999 1607 6007
rect 1621 5999 1623 6007
rect 1626 5999 1628 6007
rect 1642 5999 1644 6007
rect 1658 5999 1660 6007
rect 1679 5999 1681 6007
rect 1684 5999 1686 6007
rect 1700 5999 1702 6007
rect 1716 5999 1718 6007
rect 1721 5999 1723 6007
rect 2550 5999 2552 6007
rect 2566 5999 2568 6007
rect 2571 5999 2573 6007
rect 2587 5999 2589 6007
rect 2603 5999 2605 6007
rect 2624 5999 2626 6007
rect 2629 5999 2631 6007
rect 2645 5999 2647 6007
rect 2661 5999 2663 6007
rect 2666 5999 2668 6007
rect 857 5966 859 5974
rect 873 5966 875 5974
rect 878 5966 880 5974
rect 894 5966 896 5974
rect 910 5966 912 5974
rect 931 5966 933 5974
rect 936 5966 938 5974
rect 952 5966 954 5974
rect 968 5966 970 5974
rect 973 5966 975 5974
rect 989 5966 991 5974
rect 1005 5966 1007 5974
rect 1010 5966 1012 5974
rect 1026 5966 1028 5974
rect 1042 5966 1044 5974
rect 1063 5966 1065 5974
rect 1068 5966 1070 5974
rect 1084 5966 1086 5974
rect 1100 5966 1102 5974
rect 1105 5966 1107 5974
rect 1121 5966 1123 5974
rect 1137 5966 1139 5974
rect 1142 5966 1144 5974
rect 1158 5966 1160 5974
rect 1174 5966 1176 5974
rect 1195 5966 1197 5974
rect 1200 5966 1202 5974
rect 1216 5966 1218 5974
rect 1232 5966 1234 5974
rect 1237 5966 1239 5974
rect 1253 5966 1255 5974
rect 1269 5966 1271 5974
rect 1274 5966 1276 5974
rect 1290 5966 1292 5974
rect 1306 5966 1308 5974
rect 1327 5966 1329 5974
rect 1332 5966 1334 5974
rect 1348 5966 1350 5974
rect 1364 5966 1366 5974
rect 1369 5966 1371 5974
rect 1802 5966 1804 5974
rect 1818 5966 1820 5974
rect 1823 5966 1825 5974
rect 1839 5966 1841 5974
rect 1855 5966 1857 5974
rect 1876 5966 1878 5974
rect 1881 5966 1883 5974
rect 1897 5966 1899 5974
rect 1913 5966 1915 5974
rect 1918 5966 1920 5974
rect 1934 5966 1936 5974
rect 1950 5966 1952 5974
rect 1955 5966 1957 5974
rect 1971 5966 1973 5974
rect 1987 5966 1989 5974
rect 2008 5966 2010 5974
rect 2013 5966 2015 5974
rect 2029 5966 2031 5974
rect 2045 5966 2047 5974
rect 2050 5966 2052 5974
rect 2066 5966 2068 5974
rect 2082 5966 2084 5974
rect 2087 5966 2089 5974
rect 2103 5966 2105 5974
rect 2119 5966 2121 5974
rect 2140 5966 2142 5974
rect 2145 5966 2147 5974
rect 2161 5966 2163 5974
rect 2177 5966 2179 5974
rect 2182 5966 2184 5974
rect 2198 5966 2200 5974
rect 2214 5966 2216 5974
rect 2219 5966 2221 5974
rect 2235 5966 2237 5974
rect 2251 5966 2253 5974
rect 2272 5966 2274 5974
rect 2277 5966 2279 5974
rect 2293 5966 2295 5974
rect 2309 5966 2311 5974
rect 2314 5966 2316 5974
rect 1473 5887 1475 5895
rect 1489 5887 1491 5895
rect 1494 5887 1496 5895
rect 1510 5887 1512 5895
rect 1526 5887 1528 5895
rect 1547 5887 1549 5895
rect 1552 5887 1554 5895
rect 1568 5887 1570 5895
rect 1584 5887 1586 5895
rect 1589 5887 1591 5895
rect 1605 5887 1607 5895
rect 1621 5887 1623 5895
rect 1626 5887 1628 5895
rect 1642 5887 1644 5895
rect 1658 5887 1660 5895
rect 1679 5887 1681 5895
rect 1684 5887 1686 5895
rect 1700 5887 1702 5895
rect 1716 5887 1718 5895
rect 1721 5887 1723 5895
rect 1737 5887 1739 5895
rect 1753 5887 1755 5895
rect 1758 5887 1760 5895
rect 1774 5887 1776 5895
rect 1790 5887 1792 5895
rect 1811 5887 1813 5895
rect 1816 5887 1818 5895
rect 1832 5887 1834 5895
rect 1848 5887 1850 5895
rect 1853 5887 1855 5895
rect 2418 5887 2420 5895
rect 2434 5887 2436 5895
rect 2439 5887 2441 5895
rect 2455 5887 2457 5895
rect 2471 5887 2473 5895
rect 2492 5887 2494 5895
rect 2497 5887 2499 5895
rect 2513 5887 2515 5895
rect 2529 5887 2531 5895
rect 2534 5887 2536 5895
rect 2550 5887 2552 5895
rect 2566 5887 2568 5895
rect 2571 5887 2573 5895
rect 2587 5887 2589 5895
rect 2603 5887 2605 5895
rect 2624 5887 2626 5895
rect 2629 5887 2631 5895
rect 2645 5887 2647 5895
rect 2661 5887 2663 5895
rect 2666 5887 2668 5895
rect 2682 5887 2684 5895
rect 2698 5887 2700 5895
rect 2703 5887 2705 5895
rect 2719 5887 2721 5895
rect 2735 5887 2737 5895
rect 2756 5887 2758 5895
rect 2761 5887 2763 5895
rect 2777 5887 2779 5895
rect 2793 5887 2795 5895
rect 2798 5887 2800 5895
rect 1473 5747 1475 5755
rect 1489 5747 1491 5755
rect 1494 5747 1496 5755
rect 1510 5747 1512 5755
rect 1526 5747 1528 5755
rect 1547 5747 1549 5755
rect 1552 5747 1554 5755
rect 1568 5747 1570 5755
rect 1584 5747 1586 5755
rect 1589 5747 1591 5755
rect 1605 5747 1607 5755
rect 1621 5747 1623 5755
rect 1626 5747 1628 5755
rect 1642 5747 1644 5755
rect 1658 5747 1660 5755
rect 1679 5747 1681 5755
rect 1684 5747 1686 5755
rect 1700 5747 1702 5755
rect 1716 5747 1718 5755
rect 1721 5747 1723 5755
rect 1737 5747 1739 5755
rect 1753 5747 1755 5755
rect 1758 5747 1760 5755
rect 1774 5747 1776 5755
rect 1790 5747 1792 5755
rect 1811 5747 1813 5755
rect 1816 5747 1818 5755
rect 1832 5747 1834 5755
rect 1848 5747 1850 5755
rect 1853 5747 1855 5755
rect 2418 5747 2420 5755
rect 2434 5747 2436 5755
rect 2439 5747 2441 5755
rect 2455 5747 2457 5755
rect 2471 5747 2473 5755
rect 2492 5747 2494 5755
rect 2497 5747 2499 5755
rect 2513 5747 2515 5755
rect 2529 5747 2531 5755
rect 2534 5747 2536 5755
rect 2550 5747 2552 5755
rect 2566 5747 2568 5755
rect 2571 5747 2573 5755
rect 2587 5747 2589 5755
rect 2603 5747 2605 5755
rect 2624 5747 2626 5755
rect 2629 5747 2631 5755
rect 2645 5747 2647 5755
rect 2661 5747 2663 5755
rect 2666 5747 2668 5755
rect 2682 5747 2684 5755
rect 2698 5747 2700 5755
rect 2703 5747 2705 5755
rect 2719 5747 2721 5755
rect 2735 5747 2737 5755
rect 2756 5747 2758 5755
rect 2761 5747 2763 5755
rect 2777 5747 2779 5755
rect 2793 5747 2795 5755
rect 2798 5747 2800 5755
rect 954 5717 956 5725
rect 970 5717 972 5725
rect 975 5717 977 5725
rect 991 5717 993 5725
rect 1007 5717 1009 5725
rect 1028 5717 1030 5725
rect 1033 5717 1035 5725
rect 1049 5717 1051 5725
rect 1065 5717 1067 5725
rect 1070 5717 1072 5725
rect 1899 5717 1901 5725
rect 1915 5717 1917 5725
rect 1920 5717 1922 5725
rect 1936 5717 1938 5725
rect 1952 5717 1954 5725
rect 1973 5717 1975 5725
rect 1978 5717 1980 5725
rect 1994 5717 1996 5725
rect 2010 5717 2012 5725
rect 2015 5717 2017 5725
rect 1473 5661 1475 5669
rect 1489 5661 1491 5669
rect 1494 5661 1496 5669
rect 1510 5661 1512 5669
rect 1526 5661 1528 5669
rect 1547 5661 1549 5669
rect 1552 5661 1554 5669
rect 1568 5661 1570 5669
rect 1584 5661 1586 5669
rect 1589 5661 1591 5669
rect 1605 5661 1607 5669
rect 1621 5661 1623 5669
rect 1626 5661 1628 5669
rect 1642 5661 1644 5669
rect 1658 5661 1660 5669
rect 1679 5661 1681 5669
rect 1684 5661 1686 5669
rect 1700 5661 1702 5669
rect 1716 5661 1718 5669
rect 1721 5661 1723 5669
rect 1737 5661 1739 5669
rect 1753 5661 1755 5669
rect 1758 5661 1760 5669
rect 1774 5661 1776 5669
rect 1790 5661 1792 5669
rect 1811 5661 1813 5669
rect 1816 5661 1818 5669
rect 1832 5661 1834 5669
rect 1848 5661 1850 5669
rect 1853 5661 1855 5669
rect 2418 5661 2420 5669
rect 2434 5661 2436 5669
rect 2439 5661 2441 5669
rect 2455 5661 2457 5669
rect 2471 5661 2473 5669
rect 2492 5661 2494 5669
rect 2497 5661 2499 5669
rect 2513 5661 2515 5669
rect 2529 5661 2531 5669
rect 2534 5661 2536 5669
rect 2550 5661 2552 5669
rect 2566 5661 2568 5669
rect 2571 5661 2573 5669
rect 2587 5661 2589 5669
rect 2603 5661 2605 5669
rect 2624 5661 2626 5669
rect 2629 5661 2631 5669
rect 2645 5661 2647 5669
rect 2661 5661 2663 5669
rect 2666 5661 2668 5669
rect 2682 5661 2684 5669
rect 2698 5661 2700 5669
rect 2703 5661 2705 5669
rect 2719 5661 2721 5669
rect 2735 5661 2737 5669
rect 2756 5661 2758 5669
rect 2761 5661 2763 5669
rect 2777 5661 2779 5669
rect 2793 5661 2795 5669
rect 2798 5661 2800 5669
rect 954 5631 956 5639
rect 970 5631 972 5639
rect 975 5631 977 5639
rect 991 5631 993 5639
rect 1007 5631 1009 5639
rect 1028 5631 1030 5639
rect 1033 5631 1035 5639
rect 1049 5631 1051 5639
rect 1065 5631 1067 5639
rect 1070 5631 1072 5639
rect 1899 5631 1901 5639
rect 1915 5631 1917 5639
rect 1920 5631 1922 5639
rect 1936 5631 1938 5639
rect 1952 5631 1954 5639
rect 1973 5631 1975 5639
rect 1978 5631 1980 5639
rect 1994 5631 1996 5639
rect 2010 5631 2012 5639
rect 2015 5631 2017 5639
rect 953 5550 955 5558
rect 971 5550 973 5558
rect 976 5550 978 5558
rect 996 5550 998 5558
rect 1017 5550 1019 5558
rect 1043 5550 1045 5558
rect 1048 5550 1050 5558
rect 1071 5550 1073 5558
rect 1087 5550 1089 5558
rect 1112 5550 1114 5558
rect 1130 5550 1132 5558
rect 1159 5555 1161 5563
rect 1164 5555 1166 5563
rect 1214 5550 1216 5558
rect 1232 5550 1234 5558
rect 1237 5550 1239 5558
rect 1257 5550 1259 5558
rect 1278 5550 1280 5558
rect 1304 5550 1306 5558
rect 1309 5550 1311 5558
rect 1332 5550 1334 5558
rect 1348 5550 1350 5558
rect 1364 5550 1366 5558
rect 1898 5550 1900 5558
rect 1916 5550 1918 5558
rect 1921 5550 1923 5558
rect 1941 5550 1943 5558
rect 1962 5550 1964 5558
rect 1988 5550 1990 5558
rect 1993 5550 1995 5558
rect 2016 5550 2018 5558
rect 2032 5550 2034 5558
rect 2057 5550 2059 5558
rect 2075 5550 2077 5558
rect 2104 5555 2106 5563
rect 2109 5555 2111 5563
rect 2159 5550 2161 5558
rect 2177 5550 2179 5558
rect 2182 5550 2184 5558
rect 2202 5550 2204 5558
rect 2223 5550 2225 5558
rect 2249 5550 2251 5558
rect 2254 5550 2256 5558
rect 2277 5550 2279 5558
rect 2293 5550 2295 5558
rect 2309 5550 2311 5558
rect 1473 5519 1475 5527
rect 1489 5519 1491 5527
rect 1494 5519 1496 5527
rect 1510 5519 1512 5527
rect 1526 5519 1528 5527
rect 1547 5519 1549 5527
rect 1552 5519 1554 5527
rect 1568 5519 1570 5527
rect 1584 5519 1586 5527
rect 1589 5519 1591 5527
rect 1605 5519 1607 5527
rect 1621 5519 1623 5527
rect 1626 5519 1628 5527
rect 1642 5519 1644 5527
rect 1658 5519 1660 5527
rect 1679 5519 1681 5527
rect 1684 5519 1686 5527
rect 1700 5519 1702 5527
rect 1716 5519 1718 5527
rect 1721 5519 1723 5527
rect 1737 5519 1739 5527
rect 1753 5519 1755 5527
rect 1758 5519 1760 5527
rect 1774 5519 1776 5527
rect 1790 5519 1792 5527
rect 1811 5519 1813 5527
rect 1816 5519 1818 5527
rect 1832 5519 1834 5527
rect 1848 5519 1850 5527
rect 1853 5519 1855 5527
rect 2418 5519 2420 5527
rect 2434 5519 2436 5527
rect 2439 5519 2441 5527
rect 2455 5519 2457 5527
rect 2471 5519 2473 5527
rect 2492 5519 2494 5527
rect 2497 5519 2499 5527
rect 2513 5519 2515 5527
rect 2529 5519 2531 5527
rect 2534 5519 2536 5527
rect 2550 5519 2552 5527
rect 2566 5519 2568 5527
rect 2571 5519 2573 5527
rect 2587 5519 2589 5527
rect 2603 5519 2605 5527
rect 2624 5519 2626 5527
rect 2629 5519 2631 5527
rect 2645 5519 2647 5527
rect 2661 5519 2663 5527
rect 2666 5519 2668 5527
rect 2682 5519 2684 5527
rect 2698 5519 2700 5527
rect 2703 5519 2705 5527
rect 2719 5519 2721 5527
rect 2735 5519 2737 5527
rect 2756 5519 2758 5527
rect 2761 5519 2763 5527
rect 2777 5519 2779 5527
rect 2793 5519 2795 5527
rect 2798 5519 2800 5527
rect 1136 5451 1138 5459
rect 1159 5457 1161 5465
rect 1164 5457 1166 5465
rect 1214 5464 1216 5472
rect 1232 5464 1234 5472
rect 1237 5464 1239 5472
rect 1257 5464 1259 5472
rect 1278 5464 1280 5472
rect 1304 5464 1306 5472
rect 1309 5464 1311 5472
rect 1332 5464 1334 5472
rect 1348 5464 1350 5472
rect 1364 5464 1366 5472
rect 1768 5448 1770 5456
rect 1773 5448 1775 5456
rect 2081 5451 2083 5459
rect 2104 5457 2106 5465
rect 2109 5457 2111 5465
rect 2159 5464 2161 5472
rect 2177 5464 2179 5472
rect 2182 5464 2184 5472
rect 2202 5464 2204 5472
rect 2223 5464 2225 5472
rect 2249 5464 2251 5472
rect 2254 5464 2256 5472
rect 2277 5464 2279 5472
rect 2293 5464 2295 5472
rect 2309 5464 2311 5472
rect 988 5419 990 5427
rect 993 5419 995 5427
rect 1078 5419 1080 5427
rect 1083 5419 1085 5427
rect 1159 5419 1161 5427
rect 1164 5419 1166 5427
rect 1214 5418 1216 5426
rect 1232 5418 1234 5426
rect 1237 5418 1239 5426
rect 1257 5418 1259 5426
rect 1278 5418 1280 5426
rect 1304 5418 1306 5426
rect 1309 5418 1311 5426
rect 1332 5418 1334 5426
rect 1348 5418 1350 5426
rect 1364 5418 1366 5426
rect 1933 5419 1935 5427
rect 1938 5419 1940 5427
rect 2023 5419 2025 5427
rect 2028 5419 2030 5427
rect 2104 5419 2106 5427
rect 2109 5419 2111 5427
rect 2159 5418 2161 5426
rect 2177 5418 2179 5426
rect 2182 5418 2184 5426
rect 2202 5418 2204 5426
rect 2223 5418 2225 5426
rect 2249 5418 2251 5426
rect 2254 5418 2256 5426
rect 2277 5418 2279 5426
rect 2293 5418 2295 5426
rect 2309 5418 2311 5426
rect 965 5319 967 5327
rect 988 5325 990 5333
rect 993 5325 995 5333
rect 1019 5319 1021 5327
rect 1055 5319 1057 5327
rect 1078 5325 1080 5333
rect 1083 5325 1085 5333
rect 1654 5349 1656 5379
rect 1707 5349 1709 5379
rect 1745 5346 1747 5354
rect 1768 5352 1770 5360
rect 1773 5352 1775 5360
rect 1799 5346 1801 5354
rect 1821 5346 1823 5354
rect 1109 5319 1111 5327
rect 1136 5319 1138 5327
rect 1159 5325 1161 5333
rect 1164 5325 1166 5333
rect 1214 5332 1216 5340
rect 1232 5332 1234 5340
rect 1237 5332 1239 5340
rect 1257 5332 1259 5340
rect 1278 5332 1280 5340
rect 1304 5332 1306 5340
rect 1309 5332 1311 5340
rect 1332 5332 1334 5340
rect 1348 5332 1350 5340
rect 1364 5332 1366 5340
rect 1768 5318 1770 5326
rect 1773 5318 1775 5326
rect 1910 5319 1912 5327
rect 1933 5325 1935 5333
rect 1938 5325 1940 5333
rect 1964 5319 1966 5327
rect 2000 5319 2002 5327
rect 2023 5325 2025 5333
rect 2028 5325 2030 5333
rect 2054 5319 2056 5327
rect 2081 5319 2083 5327
rect 2104 5325 2106 5333
rect 2109 5325 2111 5333
rect 2159 5332 2161 5340
rect 2177 5332 2179 5340
rect 2182 5332 2184 5340
rect 2202 5332 2204 5340
rect 2223 5332 2225 5340
rect 2249 5332 2251 5340
rect 2254 5332 2256 5340
rect 2277 5332 2279 5340
rect 2293 5332 2295 5340
rect 2309 5332 2311 5340
rect 1054 5284 1056 5292
rect 1059 5284 1061 5292
rect 1159 5284 1161 5292
rect 1164 5284 1166 5292
rect 1214 5286 1216 5294
rect 1232 5286 1234 5294
rect 1237 5286 1239 5294
rect 1257 5286 1259 5294
rect 1278 5286 1280 5294
rect 1304 5286 1306 5294
rect 1309 5286 1311 5294
rect 1332 5286 1334 5294
rect 1348 5286 1350 5294
rect 1364 5286 1366 5294
rect 1999 5284 2001 5292
rect 2004 5284 2006 5292
rect 2104 5284 2106 5292
rect 2109 5284 2111 5292
rect 2159 5286 2161 5294
rect 2177 5286 2179 5294
rect 2182 5286 2184 5294
rect 2202 5286 2204 5294
rect 2223 5286 2225 5294
rect 2249 5286 2251 5294
rect 2254 5286 2256 5294
rect 2277 5286 2279 5294
rect 2293 5286 2295 5294
rect 2309 5286 2311 5294
rect 1031 5187 1033 5195
rect 1054 5193 1056 5201
rect 1059 5193 1061 5201
rect 1560 5219 1562 5249
rect 1613 5219 1615 5249
rect 1745 5216 1747 5224
rect 1768 5222 1770 5230
rect 1773 5222 1775 5230
rect 1799 5216 1801 5224
rect 1085 5187 1087 5195
rect 1136 5187 1138 5195
rect 1159 5193 1161 5201
rect 1164 5193 1166 5201
rect 1214 5200 1216 5208
rect 1232 5200 1234 5208
rect 1237 5200 1239 5208
rect 1257 5200 1259 5208
rect 1278 5200 1280 5208
rect 1304 5200 1306 5208
rect 1309 5200 1311 5208
rect 1332 5200 1334 5208
rect 1348 5200 1350 5208
rect 1364 5200 1366 5208
rect 1976 5187 1978 5195
rect 1999 5193 2001 5201
rect 2004 5193 2006 5201
rect 2030 5187 2032 5195
rect 2081 5187 2083 5195
rect 2104 5193 2106 5201
rect 2109 5193 2111 5201
rect 2159 5200 2161 5208
rect 2177 5200 2179 5208
rect 2182 5200 2184 5208
rect 2202 5200 2204 5208
rect 2223 5200 2225 5208
rect 2249 5200 2251 5208
rect 2254 5200 2256 5208
rect 2277 5200 2279 5208
rect 2293 5200 2295 5208
rect 2309 5200 2311 5208
rect 1078 5153 1080 5161
rect 1083 5153 1085 5161
rect 1159 5153 1161 5161
rect 1164 5153 1166 5161
rect 1214 5154 1216 5162
rect 1232 5154 1234 5162
rect 1237 5154 1239 5162
rect 1257 5154 1259 5162
rect 1278 5154 1280 5162
rect 1304 5154 1306 5162
rect 1309 5154 1311 5162
rect 1332 5154 1334 5162
rect 1348 5154 1350 5162
rect 1364 5154 1366 5162
rect 2023 5153 2025 5161
rect 2028 5153 2030 5161
rect 2104 5153 2106 5161
rect 2109 5153 2111 5161
rect 2159 5154 2161 5162
rect 2177 5154 2179 5162
rect 2182 5154 2184 5162
rect 2202 5154 2204 5162
rect 2223 5154 2225 5162
rect 2249 5154 2251 5162
rect 2254 5154 2256 5162
rect 2277 5154 2279 5162
rect 2293 5154 2295 5162
rect 2309 5154 2311 5162
rect 1614 5119 1616 5127
rect 1619 5119 1621 5127
rect 1635 5119 1637 5127
rect 1651 5119 1653 5127
rect 1656 5119 1658 5127
rect 1677 5119 1679 5127
rect 1693 5119 1695 5127
rect 1709 5119 1711 5127
rect 1714 5119 1716 5127
rect 1730 5119 1732 5127
rect 2559 5119 2561 5127
rect 2564 5119 2566 5127
rect 2580 5119 2582 5127
rect 2596 5119 2598 5127
rect 2601 5119 2603 5127
rect 2622 5119 2624 5127
rect 2638 5119 2640 5127
rect 2654 5119 2656 5127
rect 2659 5119 2661 5127
rect 2675 5119 2677 5127
rect 1055 5055 1057 5063
rect 1078 5061 1080 5069
rect 1083 5061 1085 5069
rect 1109 5055 1111 5063
rect 1136 5055 1138 5063
rect 1159 5061 1161 5069
rect 1164 5061 1166 5069
rect 1214 5068 1216 5076
rect 1232 5068 1234 5076
rect 1237 5068 1239 5076
rect 1257 5068 1259 5076
rect 1278 5068 1280 5076
rect 1304 5068 1306 5076
rect 1309 5068 1311 5076
rect 1332 5068 1334 5076
rect 1348 5068 1350 5076
rect 1364 5068 1366 5076
rect 1190 5055 1192 5063
rect 2000 5055 2002 5063
rect 2023 5061 2025 5069
rect 2028 5061 2030 5069
rect 2054 5055 2056 5063
rect 2081 5055 2083 5063
rect 2104 5061 2106 5069
rect 2109 5061 2111 5069
rect 2159 5068 2161 5076
rect 2177 5068 2179 5076
rect 2182 5068 2184 5076
rect 2202 5068 2204 5076
rect 2223 5068 2225 5076
rect 2249 5068 2251 5076
rect 2254 5068 2256 5076
rect 2277 5068 2279 5076
rect 2293 5068 2295 5076
rect 2309 5068 2311 5076
rect 2135 5055 2137 5063
rect 1605 5017 1607 5025
rect 1621 5017 1623 5025
rect 1626 5017 1628 5025
rect 1642 5017 1644 5025
rect 1658 5017 1660 5025
rect 1679 5017 1681 5025
rect 1684 5017 1686 5025
rect 1700 5017 1702 5025
rect 1716 5017 1718 5025
rect 1721 5017 1723 5025
rect 2550 5017 2552 5025
rect 2566 5017 2568 5025
rect 2571 5017 2573 5025
rect 2587 5017 2589 5025
rect 2603 5017 2605 5025
rect 2624 5017 2626 5025
rect 2629 5017 2631 5025
rect 2645 5017 2647 5025
rect 2661 5017 2663 5025
rect 2666 5017 2668 5025
rect 857 4984 859 4992
rect 873 4984 875 4992
rect 878 4984 880 4992
rect 894 4984 896 4992
rect 910 4984 912 4992
rect 931 4984 933 4992
rect 936 4984 938 4992
rect 952 4984 954 4992
rect 968 4984 970 4992
rect 973 4984 975 4992
rect 989 4984 991 4992
rect 1005 4984 1007 4992
rect 1010 4984 1012 4992
rect 1026 4984 1028 4992
rect 1042 4984 1044 4992
rect 1063 4984 1065 4992
rect 1068 4984 1070 4992
rect 1084 4984 1086 4992
rect 1100 4984 1102 4992
rect 1105 4984 1107 4992
rect 1121 4984 1123 4992
rect 1137 4984 1139 4992
rect 1142 4984 1144 4992
rect 1158 4984 1160 4992
rect 1174 4984 1176 4992
rect 1195 4984 1197 4992
rect 1200 4984 1202 4992
rect 1216 4984 1218 4992
rect 1232 4984 1234 4992
rect 1237 4984 1239 4992
rect 1253 4984 1255 4992
rect 1269 4984 1271 4992
rect 1274 4984 1276 4992
rect 1290 4984 1292 4992
rect 1306 4984 1308 4992
rect 1327 4984 1329 4992
rect 1332 4984 1334 4992
rect 1348 4984 1350 4992
rect 1364 4984 1366 4992
rect 1369 4984 1371 4992
rect 1802 4984 1804 4992
rect 1818 4984 1820 4992
rect 1823 4984 1825 4992
rect 1839 4984 1841 4992
rect 1855 4984 1857 4992
rect 1876 4984 1878 4992
rect 1881 4984 1883 4992
rect 1897 4984 1899 4992
rect 1913 4984 1915 4992
rect 1918 4984 1920 4992
rect 1934 4984 1936 4992
rect 1950 4984 1952 4992
rect 1955 4984 1957 4992
rect 1971 4984 1973 4992
rect 1987 4984 1989 4992
rect 2008 4984 2010 4992
rect 2013 4984 2015 4992
rect 2029 4984 2031 4992
rect 2045 4984 2047 4992
rect 2050 4984 2052 4992
rect 2066 4984 2068 4992
rect 2082 4984 2084 4992
rect 2087 4984 2089 4992
rect 2103 4984 2105 4992
rect 2119 4984 2121 4992
rect 2140 4984 2142 4992
rect 2145 4984 2147 4992
rect 2161 4984 2163 4992
rect 2177 4984 2179 4992
rect 2182 4984 2184 4992
rect 2198 4984 2200 4992
rect 2214 4984 2216 4992
rect 2219 4984 2221 4992
rect 2235 4984 2237 4992
rect 2251 4984 2253 4992
rect 2272 4984 2274 4992
rect 2277 4984 2279 4992
rect 2293 4984 2295 4992
rect 2309 4984 2311 4992
rect 2314 4984 2316 4992
rect 4579 7889 4581 7945
rect 4587 7889 4589 7945
rect 4595 7889 4597 7945
rect 4603 7889 4605 7945
rect 4611 7889 4613 7945
rect 4619 7889 4621 7945
rect 4634 7857 4636 7945
rect 4642 7857 4644 7945
rect 4650 7857 4652 7945
rect 4658 7857 4660 7945
rect 4677 7857 4679 7945
rect 4685 7857 4687 7945
rect 4693 7857 4695 7945
rect 4701 7857 4703 7945
rect 4718 7857 4720 7945
rect 4726 7857 4728 7945
rect 4734 7857 4736 7945
rect 4742 7857 4744 7945
rect 4577 7372 4579 7428
rect 4585 7372 4587 7428
rect 4593 7372 4595 7428
rect 4601 7372 4603 7428
rect 4609 7372 4611 7428
rect 4617 7372 4619 7428
rect 1210 4528 1266 4530
rect 1210 4520 1266 4522
rect 1210 4512 1266 4514
rect 1210 4504 1266 4506
rect 2137 4528 2193 4530
rect 2137 4520 2193 4522
rect 2137 4512 2193 4514
rect 2137 4504 2193 4506
rect 2446 4528 2502 4530
rect 2446 4520 2502 4522
rect 2446 4512 2502 4514
rect 2446 4504 2502 4506
rect 2755 4528 2811 4530
rect 2755 4520 2811 4522
rect 2755 4512 2811 4514
rect 2755 4504 2811 4506
rect 3064 4528 3120 4530
rect 3064 4520 3120 4522
rect 3064 4512 3120 4514
rect 3064 4504 3120 4506
rect 3373 4528 3429 4530
rect 3373 4520 3429 4522
rect 3373 4512 3429 4514
rect 3373 4504 3429 4506
rect 1210 4496 1266 4498
rect 2137 4496 2193 4498
rect 2446 4496 2502 4498
rect 2755 4496 2811 4498
rect 3064 4496 3120 4498
rect 3373 4496 3429 4498
rect 1210 4488 1266 4490
rect 2137 4488 2193 4490
rect 2446 4488 2502 4490
rect 2755 4488 2811 4490
rect 3064 4488 3120 4490
rect 3373 4488 3429 4490
<< ndiffusion >>
rect 1397 9949 1402 9953
rect 1406 9949 1412 9953
rect 1416 9949 1422 9953
rect 1426 9949 1432 9953
rect 1436 9949 1441 9953
rect 1397 9948 1441 9949
rect 1401 9944 1407 9948
rect 1411 9944 1417 9948
rect 1421 9944 1427 9948
rect 1431 9944 1437 9948
rect 1397 9943 1441 9944
rect 1397 9939 1402 9943
rect 1406 9939 1412 9943
rect 1416 9939 1422 9943
rect 1426 9939 1432 9943
rect 1436 9939 1441 9943
rect 1397 9938 1441 9939
rect 1401 9934 1407 9938
rect 1411 9934 1417 9938
rect 1421 9934 1427 9938
rect 1431 9934 1437 9938
rect 1397 9933 1441 9934
rect 1397 9929 1402 9933
rect 1406 9929 1412 9933
rect 1416 9929 1422 9933
rect 1426 9929 1432 9933
rect 1436 9929 1441 9933
rect 1397 9928 1441 9929
rect 1401 9924 1407 9928
rect 1411 9924 1417 9928
rect 1421 9924 1427 9928
rect 1431 9924 1437 9928
rect 1397 9923 1441 9924
rect 1397 9919 1402 9923
rect 1406 9919 1412 9923
rect 1416 9919 1422 9923
rect 1426 9919 1432 9923
rect 1436 9919 1441 9923
rect 1397 9918 1441 9919
rect 1401 9914 1407 9918
rect 1411 9914 1417 9918
rect 1421 9914 1427 9918
rect 1431 9914 1437 9918
rect 1397 9913 1441 9914
rect 1397 9909 1402 9913
rect 1406 9909 1412 9913
rect 1416 9909 1422 9913
rect 1426 9909 1432 9913
rect 1436 9909 1441 9913
rect 1397 9908 1441 9909
rect 1401 9904 1407 9908
rect 1411 9904 1417 9908
rect 1421 9904 1427 9908
rect 1431 9904 1437 9908
rect 1397 9903 1441 9904
rect 1397 9899 1402 9903
rect 1406 9899 1412 9903
rect 1416 9899 1422 9903
rect 1426 9899 1432 9903
rect 1436 9899 1441 9903
rect 1397 9898 1441 9899
rect 1401 9894 1407 9898
rect 1411 9894 1417 9898
rect 1421 9894 1427 9898
rect 1431 9894 1437 9898
rect 1397 9893 1441 9894
rect 1397 9889 1402 9893
rect 1406 9889 1412 9893
rect 1416 9889 1422 9893
rect 1426 9889 1432 9893
rect 1436 9889 1441 9893
rect 1397 9888 1441 9889
rect 1401 9884 1407 9888
rect 1411 9884 1417 9888
rect 1421 9884 1427 9888
rect 1431 9884 1437 9888
rect 1397 9883 1441 9884
rect 1397 9879 1402 9883
rect 1406 9879 1412 9883
rect 1416 9879 1422 9883
rect 1426 9879 1432 9883
rect 1436 9879 1441 9883
rect 1397 9878 1441 9879
rect 1401 9874 1407 9878
rect 1411 9874 1417 9878
rect 1421 9874 1427 9878
rect 1431 9874 1437 9878
rect 1397 9873 1441 9874
rect 1397 9869 1402 9873
rect 1406 9869 1412 9873
rect 1416 9869 1422 9873
rect 1426 9869 1432 9873
rect 1436 9869 1441 9873
rect 1397 9868 1441 9869
rect 1401 9864 1407 9868
rect 1411 9864 1417 9868
rect 1421 9864 1427 9868
rect 1431 9864 1437 9868
rect 1706 9949 1711 9953
rect 1715 9949 1721 9953
rect 1725 9949 1731 9953
rect 1735 9949 1741 9953
rect 1745 9949 1750 9953
rect 1706 9948 1750 9949
rect 1710 9944 1716 9948
rect 1720 9944 1726 9948
rect 1730 9944 1736 9948
rect 1740 9944 1746 9948
rect 1706 9943 1750 9944
rect 1706 9939 1711 9943
rect 1715 9939 1721 9943
rect 1725 9939 1731 9943
rect 1735 9939 1741 9943
rect 1745 9939 1750 9943
rect 1706 9938 1750 9939
rect 1710 9934 1716 9938
rect 1720 9934 1726 9938
rect 1730 9934 1736 9938
rect 1740 9934 1746 9938
rect 1706 9933 1750 9934
rect 1706 9929 1711 9933
rect 1715 9929 1721 9933
rect 1725 9929 1731 9933
rect 1735 9929 1741 9933
rect 1745 9929 1750 9933
rect 1706 9928 1750 9929
rect 1710 9924 1716 9928
rect 1720 9924 1726 9928
rect 1730 9924 1736 9928
rect 1740 9924 1746 9928
rect 1706 9923 1750 9924
rect 1706 9919 1711 9923
rect 1715 9919 1721 9923
rect 1725 9919 1731 9923
rect 1735 9919 1741 9923
rect 1745 9919 1750 9923
rect 1706 9918 1750 9919
rect 1710 9914 1716 9918
rect 1720 9914 1726 9918
rect 1730 9914 1736 9918
rect 1740 9914 1746 9918
rect 1706 9913 1750 9914
rect 1706 9909 1711 9913
rect 1715 9909 1721 9913
rect 1725 9909 1731 9913
rect 1735 9909 1741 9913
rect 1745 9909 1750 9913
rect 1706 9908 1750 9909
rect 1710 9904 1716 9908
rect 1720 9904 1726 9908
rect 1730 9904 1736 9908
rect 1740 9904 1746 9908
rect 1706 9903 1750 9904
rect 1706 9899 1711 9903
rect 1715 9899 1721 9903
rect 1725 9899 1731 9903
rect 1735 9899 1741 9903
rect 1745 9899 1750 9903
rect 1706 9898 1750 9899
rect 1710 9894 1716 9898
rect 1720 9894 1726 9898
rect 1730 9894 1736 9898
rect 1740 9894 1746 9898
rect 1706 9893 1750 9894
rect 1706 9889 1711 9893
rect 1715 9889 1721 9893
rect 1725 9889 1731 9893
rect 1735 9889 1741 9893
rect 1745 9889 1750 9893
rect 1706 9888 1750 9889
rect 1710 9884 1716 9888
rect 1720 9884 1726 9888
rect 1730 9884 1736 9888
rect 1740 9884 1746 9888
rect 1706 9883 1750 9884
rect 1706 9879 1711 9883
rect 1715 9879 1721 9883
rect 1725 9879 1731 9883
rect 1735 9879 1741 9883
rect 1745 9879 1750 9883
rect 1706 9878 1750 9879
rect 1710 9874 1716 9878
rect 1720 9874 1726 9878
rect 1730 9874 1736 9878
rect 1740 9874 1746 9878
rect 1706 9873 1750 9874
rect 1706 9869 1711 9873
rect 1715 9869 1721 9873
rect 1725 9869 1731 9873
rect 1735 9869 1741 9873
rect 1745 9869 1750 9873
rect 1706 9868 1750 9869
rect 1710 9864 1716 9868
rect 1720 9864 1726 9868
rect 1730 9864 1736 9868
rect 1740 9864 1746 9868
rect 2015 9949 2020 9953
rect 2024 9949 2030 9953
rect 2034 9949 2040 9953
rect 2044 9949 2050 9953
rect 2054 9949 2059 9953
rect 2015 9948 2059 9949
rect 2019 9944 2025 9948
rect 2029 9944 2035 9948
rect 2039 9944 2045 9948
rect 2049 9944 2055 9948
rect 2015 9943 2059 9944
rect 2015 9939 2020 9943
rect 2024 9939 2030 9943
rect 2034 9939 2040 9943
rect 2044 9939 2050 9943
rect 2054 9939 2059 9943
rect 2015 9938 2059 9939
rect 2019 9934 2025 9938
rect 2029 9934 2035 9938
rect 2039 9934 2045 9938
rect 2049 9934 2055 9938
rect 2015 9933 2059 9934
rect 2015 9929 2020 9933
rect 2024 9929 2030 9933
rect 2034 9929 2040 9933
rect 2044 9929 2050 9933
rect 2054 9929 2059 9933
rect 2015 9928 2059 9929
rect 2019 9924 2025 9928
rect 2029 9924 2035 9928
rect 2039 9924 2045 9928
rect 2049 9924 2055 9928
rect 2015 9923 2059 9924
rect 2015 9919 2020 9923
rect 2024 9919 2030 9923
rect 2034 9919 2040 9923
rect 2044 9919 2050 9923
rect 2054 9919 2059 9923
rect 2015 9918 2059 9919
rect 2019 9914 2025 9918
rect 2029 9914 2035 9918
rect 2039 9914 2045 9918
rect 2049 9914 2055 9918
rect 2015 9913 2059 9914
rect 2015 9909 2020 9913
rect 2024 9909 2030 9913
rect 2034 9909 2040 9913
rect 2044 9909 2050 9913
rect 2054 9909 2059 9913
rect 2015 9908 2059 9909
rect 2019 9904 2025 9908
rect 2029 9904 2035 9908
rect 2039 9904 2045 9908
rect 2049 9904 2055 9908
rect 2015 9903 2059 9904
rect 2015 9899 2020 9903
rect 2024 9899 2030 9903
rect 2034 9899 2040 9903
rect 2044 9899 2050 9903
rect 2054 9899 2059 9903
rect 2015 9898 2059 9899
rect 2019 9894 2025 9898
rect 2029 9894 2035 9898
rect 2039 9894 2045 9898
rect 2049 9894 2055 9898
rect 2015 9893 2059 9894
rect 2015 9889 2020 9893
rect 2024 9889 2030 9893
rect 2034 9889 2040 9893
rect 2044 9889 2050 9893
rect 2054 9889 2059 9893
rect 2015 9888 2059 9889
rect 2019 9884 2025 9888
rect 2029 9884 2035 9888
rect 2039 9884 2045 9888
rect 2049 9884 2055 9888
rect 2015 9883 2059 9884
rect 2015 9879 2020 9883
rect 2024 9879 2030 9883
rect 2034 9879 2040 9883
rect 2044 9879 2050 9883
rect 2054 9879 2059 9883
rect 2015 9878 2059 9879
rect 2019 9874 2025 9878
rect 2029 9874 2035 9878
rect 2039 9874 2045 9878
rect 2049 9874 2055 9878
rect 2015 9873 2059 9874
rect 2015 9869 2020 9873
rect 2024 9869 2030 9873
rect 2034 9869 2040 9873
rect 2044 9869 2050 9873
rect 2054 9869 2059 9873
rect 2015 9868 2059 9869
rect 2019 9864 2025 9868
rect 2029 9864 2035 9868
rect 2039 9864 2045 9868
rect 2049 9864 2055 9868
rect 2324 9949 2329 9953
rect 2333 9949 2339 9953
rect 2343 9949 2349 9953
rect 2353 9949 2359 9953
rect 2363 9949 2368 9953
rect 2324 9948 2368 9949
rect 2328 9944 2334 9948
rect 2338 9944 2344 9948
rect 2348 9944 2354 9948
rect 2358 9944 2364 9948
rect 2324 9943 2368 9944
rect 2324 9939 2329 9943
rect 2333 9939 2339 9943
rect 2343 9939 2349 9943
rect 2353 9939 2359 9943
rect 2363 9939 2368 9943
rect 2324 9938 2368 9939
rect 2328 9934 2334 9938
rect 2338 9934 2344 9938
rect 2348 9934 2354 9938
rect 2358 9934 2364 9938
rect 2324 9933 2368 9934
rect 2324 9929 2329 9933
rect 2333 9929 2339 9933
rect 2343 9929 2349 9933
rect 2353 9929 2359 9933
rect 2363 9929 2368 9933
rect 2324 9928 2368 9929
rect 2328 9924 2334 9928
rect 2338 9924 2344 9928
rect 2348 9924 2354 9928
rect 2358 9924 2364 9928
rect 2324 9923 2368 9924
rect 2324 9919 2329 9923
rect 2333 9919 2339 9923
rect 2343 9919 2349 9923
rect 2353 9919 2359 9923
rect 2363 9919 2368 9923
rect 2324 9918 2368 9919
rect 2328 9914 2334 9918
rect 2338 9914 2344 9918
rect 2348 9914 2354 9918
rect 2358 9914 2364 9918
rect 2324 9913 2368 9914
rect 2324 9909 2329 9913
rect 2333 9909 2339 9913
rect 2343 9909 2349 9913
rect 2353 9909 2359 9913
rect 2363 9909 2368 9913
rect 2324 9908 2368 9909
rect 2328 9904 2334 9908
rect 2338 9904 2344 9908
rect 2348 9904 2354 9908
rect 2358 9904 2364 9908
rect 2324 9903 2368 9904
rect 2324 9899 2329 9903
rect 2333 9899 2339 9903
rect 2343 9899 2349 9903
rect 2353 9899 2359 9903
rect 2363 9899 2368 9903
rect 2324 9898 2368 9899
rect 2328 9894 2334 9898
rect 2338 9894 2344 9898
rect 2348 9894 2354 9898
rect 2358 9894 2364 9898
rect 2324 9893 2368 9894
rect 2324 9889 2329 9893
rect 2333 9889 2339 9893
rect 2343 9889 2349 9893
rect 2353 9889 2359 9893
rect 2363 9889 2368 9893
rect 2324 9888 2368 9889
rect 2328 9884 2334 9888
rect 2338 9884 2344 9888
rect 2348 9884 2354 9888
rect 2358 9884 2364 9888
rect 2324 9883 2368 9884
rect 2324 9879 2329 9883
rect 2333 9879 2339 9883
rect 2343 9879 2349 9883
rect 2353 9879 2359 9883
rect 2363 9879 2368 9883
rect 2324 9878 2368 9879
rect 2328 9874 2334 9878
rect 2338 9874 2344 9878
rect 2348 9874 2354 9878
rect 2358 9874 2364 9878
rect 2324 9873 2368 9874
rect 2324 9869 2329 9873
rect 2333 9869 2339 9873
rect 2343 9869 2349 9873
rect 2353 9869 2359 9873
rect 2363 9869 2368 9873
rect 2324 9868 2368 9869
rect 2328 9864 2334 9868
rect 2338 9864 2344 9868
rect 2348 9864 2354 9868
rect 2358 9864 2364 9868
rect 2633 9949 2638 9953
rect 2642 9949 2648 9953
rect 2652 9949 2658 9953
rect 2662 9949 2668 9953
rect 2672 9949 2677 9953
rect 2633 9948 2677 9949
rect 2637 9944 2643 9948
rect 2647 9944 2653 9948
rect 2657 9944 2663 9948
rect 2667 9944 2673 9948
rect 2633 9943 2677 9944
rect 2633 9939 2638 9943
rect 2642 9939 2648 9943
rect 2652 9939 2658 9943
rect 2662 9939 2668 9943
rect 2672 9939 2677 9943
rect 2633 9938 2677 9939
rect 2637 9934 2643 9938
rect 2647 9934 2653 9938
rect 2657 9934 2663 9938
rect 2667 9934 2673 9938
rect 2633 9933 2677 9934
rect 2633 9929 2638 9933
rect 2642 9929 2648 9933
rect 2652 9929 2658 9933
rect 2662 9929 2668 9933
rect 2672 9929 2677 9933
rect 2633 9928 2677 9929
rect 2637 9924 2643 9928
rect 2647 9924 2653 9928
rect 2657 9924 2663 9928
rect 2667 9924 2673 9928
rect 2633 9923 2677 9924
rect 2633 9919 2638 9923
rect 2642 9919 2648 9923
rect 2652 9919 2658 9923
rect 2662 9919 2668 9923
rect 2672 9919 2677 9923
rect 2633 9918 2677 9919
rect 2637 9914 2643 9918
rect 2647 9914 2653 9918
rect 2657 9914 2663 9918
rect 2667 9914 2673 9918
rect 2633 9913 2677 9914
rect 2633 9909 2638 9913
rect 2642 9909 2648 9913
rect 2652 9909 2658 9913
rect 2662 9909 2668 9913
rect 2672 9909 2677 9913
rect 2633 9908 2677 9909
rect 2637 9904 2643 9908
rect 2647 9904 2653 9908
rect 2657 9904 2663 9908
rect 2667 9904 2673 9908
rect 2633 9903 2677 9904
rect 2633 9899 2638 9903
rect 2642 9899 2648 9903
rect 2652 9899 2658 9903
rect 2662 9899 2668 9903
rect 2672 9899 2677 9903
rect 2633 9898 2677 9899
rect 2637 9894 2643 9898
rect 2647 9894 2653 9898
rect 2657 9894 2663 9898
rect 2667 9894 2673 9898
rect 2633 9893 2677 9894
rect 2633 9889 2638 9893
rect 2642 9889 2648 9893
rect 2652 9889 2658 9893
rect 2662 9889 2668 9893
rect 2672 9889 2677 9893
rect 2633 9888 2677 9889
rect 2637 9884 2643 9888
rect 2647 9884 2653 9888
rect 2657 9884 2663 9888
rect 2667 9884 2673 9888
rect 2633 9883 2677 9884
rect 2633 9879 2638 9883
rect 2642 9879 2648 9883
rect 2652 9879 2658 9883
rect 2662 9879 2668 9883
rect 2672 9879 2677 9883
rect 2633 9878 2677 9879
rect 2637 9874 2643 9878
rect 2647 9874 2653 9878
rect 2657 9874 2663 9878
rect 2667 9874 2673 9878
rect 2633 9873 2677 9874
rect 2633 9869 2638 9873
rect 2642 9869 2648 9873
rect 2652 9869 2658 9873
rect 2662 9869 2668 9873
rect 2672 9869 2677 9873
rect 2633 9868 2677 9869
rect 2637 9864 2643 9868
rect 2647 9864 2653 9868
rect 2657 9864 2663 9868
rect 2667 9864 2673 9868
rect 2942 9949 2947 9953
rect 2951 9949 2957 9953
rect 2961 9949 2967 9953
rect 2971 9949 2977 9953
rect 2981 9949 2986 9953
rect 2942 9948 2986 9949
rect 2946 9944 2952 9948
rect 2956 9944 2962 9948
rect 2966 9944 2972 9948
rect 2976 9944 2982 9948
rect 2942 9943 2986 9944
rect 2942 9939 2947 9943
rect 2951 9939 2957 9943
rect 2961 9939 2967 9943
rect 2971 9939 2977 9943
rect 2981 9939 2986 9943
rect 2942 9938 2986 9939
rect 2946 9934 2952 9938
rect 2956 9934 2962 9938
rect 2966 9934 2972 9938
rect 2976 9934 2982 9938
rect 2942 9933 2986 9934
rect 2942 9929 2947 9933
rect 2951 9929 2957 9933
rect 2961 9929 2967 9933
rect 2971 9929 2977 9933
rect 2981 9929 2986 9933
rect 2942 9928 2986 9929
rect 2946 9924 2952 9928
rect 2956 9924 2962 9928
rect 2966 9924 2972 9928
rect 2976 9924 2982 9928
rect 2942 9923 2986 9924
rect 2942 9919 2947 9923
rect 2951 9919 2957 9923
rect 2961 9919 2967 9923
rect 2971 9919 2977 9923
rect 2981 9919 2986 9923
rect 2942 9918 2986 9919
rect 2946 9914 2952 9918
rect 2956 9914 2962 9918
rect 2966 9914 2972 9918
rect 2976 9914 2982 9918
rect 2942 9913 2986 9914
rect 2942 9909 2947 9913
rect 2951 9909 2957 9913
rect 2961 9909 2967 9913
rect 2971 9909 2977 9913
rect 2981 9909 2986 9913
rect 2942 9908 2986 9909
rect 2946 9904 2952 9908
rect 2956 9904 2962 9908
rect 2966 9904 2972 9908
rect 2976 9904 2982 9908
rect 2942 9903 2986 9904
rect 2942 9899 2947 9903
rect 2951 9899 2957 9903
rect 2961 9899 2967 9903
rect 2971 9899 2977 9903
rect 2981 9899 2986 9903
rect 2942 9898 2986 9899
rect 2946 9894 2952 9898
rect 2956 9894 2962 9898
rect 2966 9894 2972 9898
rect 2976 9894 2982 9898
rect 2942 9893 2986 9894
rect 2942 9889 2947 9893
rect 2951 9889 2957 9893
rect 2961 9889 2967 9893
rect 2971 9889 2977 9893
rect 2981 9889 2986 9893
rect 2942 9888 2986 9889
rect 2946 9884 2952 9888
rect 2956 9884 2962 9888
rect 2966 9884 2972 9888
rect 2976 9884 2982 9888
rect 2942 9883 2986 9884
rect 2942 9879 2947 9883
rect 2951 9879 2957 9883
rect 2961 9879 2967 9883
rect 2971 9879 2977 9883
rect 2981 9879 2986 9883
rect 2942 9878 2986 9879
rect 2946 9874 2952 9878
rect 2956 9874 2962 9878
rect 2966 9874 2972 9878
rect 2976 9874 2982 9878
rect 2942 9873 2986 9874
rect 2942 9869 2947 9873
rect 2951 9869 2957 9873
rect 2961 9869 2967 9873
rect 2971 9869 2977 9873
rect 2981 9869 2986 9873
rect 2942 9868 2986 9869
rect 2946 9864 2952 9868
rect 2956 9864 2962 9868
rect 2966 9864 2972 9868
rect 2976 9864 2982 9868
rect 3251 9949 3256 9953
rect 3260 9949 3266 9953
rect 3270 9949 3276 9953
rect 3280 9949 3286 9953
rect 3290 9949 3295 9953
rect 3251 9948 3295 9949
rect 3255 9944 3261 9948
rect 3265 9944 3271 9948
rect 3275 9944 3281 9948
rect 3285 9944 3291 9948
rect 3251 9943 3295 9944
rect 3251 9939 3256 9943
rect 3260 9939 3266 9943
rect 3270 9939 3276 9943
rect 3280 9939 3286 9943
rect 3290 9939 3295 9943
rect 3251 9938 3295 9939
rect 3255 9934 3261 9938
rect 3265 9934 3271 9938
rect 3275 9934 3281 9938
rect 3285 9934 3291 9938
rect 3251 9933 3295 9934
rect 3251 9929 3256 9933
rect 3260 9929 3266 9933
rect 3270 9929 3276 9933
rect 3280 9929 3286 9933
rect 3290 9929 3295 9933
rect 3251 9928 3295 9929
rect 3255 9924 3261 9928
rect 3265 9924 3271 9928
rect 3275 9924 3281 9928
rect 3285 9924 3291 9928
rect 3251 9923 3295 9924
rect 3251 9919 3256 9923
rect 3260 9919 3266 9923
rect 3270 9919 3276 9923
rect 3280 9919 3286 9923
rect 3290 9919 3295 9923
rect 3251 9918 3295 9919
rect 3255 9914 3261 9918
rect 3265 9914 3271 9918
rect 3275 9914 3281 9918
rect 3285 9914 3291 9918
rect 3251 9913 3295 9914
rect 3251 9909 3256 9913
rect 3260 9909 3266 9913
rect 3270 9909 3276 9913
rect 3280 9909 3286 9913
rect 3290 9909 3295 9913
rect 3251 9908 3295 9909
rect 3255 9904 3261 9908
rect 3265 9904 3271 9908
rect 3275 9904 3281 9908
rect 3285 9904 3291 9908
rect 3251 9903 3295 9904
rect 3251 9899 3256 9903
rect 3260 9899 3266 9903
rect 3270 9899 3276 9903
rect 3280 9899 3286 9903
rect 3290 9899 3295 9903
rect 3251 9898 3295 9899
rect 3255 9894 3261 9898
rect 3265 9894 3271 9898
rect 3275 9894 3281 9898
rect 3285 9894 3291 9898
rect 3251 9893 3295 9894
rect 3251 9889 3256 9893
rect 3260 9889 3266 9893
rect 3270 9889 3276 9893
rect 3280 9889 3286 9893
rect 3290 9889 3295 9893
rect 3251 9888 3295 9889
rect 3255 9884 3261 9888
rect 3265 9884 3271 9888
rect 3275 9884 3281 9888
rect 3285 9884 3291 9888
rect 3251 9883 3295 9884
rect 3251 9879 3256 9883
rect 3260 9879 3266 9883
rect 3270 9879 3276 9883
rect 3280 9879 3286 9883
rect 3290 9879 3295 9883
rect 3251 9878 3295 9879
rect 3255 9874 3261 9878
rect 3265 9874 3271 9878
rect 3275 9874 3281 9878
rect 3285 9874 3291 9878
rect 3251 9873 3295 9874
rect 3251 9869 3256 9873
rect 3260 9869 3266 9873
rect 3270 9869 3276 9873
rect 3280 9869 3286 9873
rect 3290 9869 3295 9873
rect 3251 9868 3295 9869
rect 3255 9864 3261 9868
rect 3265 9864 3271 9868
rect 3275 9864 3281 9868
rect 3285 9864 3291 9868
rect 3560 9949 3565 9953
rect 3569 9949 3575 9953
rect 3579 9949 3585 9953
rect 3589 9949 3595 9953
rect 3599 9949 3604 9953
rect 3560 9948 3604 9949
rect 3564 9944 3570 9948
rect 3574 9944 3580 9948
rect 3584 9944 3590 9948
rect 3594 9944 3600 9948
rect 3560 9943 3604 9944
rect 3560 9939 3565 9943
rect 3569 9939 3575 9943
rect 3579 9939 3585 9943
rect 3589 9939 3595 9943
rect 3599 9939 3604 9943
rect 3560 9938 3604 9939
rect 3564 9934 3570 9938
rect 3574 9934 3580 9938
rect 3584 9934 3590 9938
rect 3594 9934 3600 9938
rect 3560 9933 3604 9934
rect 3560 9929 3565 9933
rect 3569 9929 3575 9933
rect 3579 9929 3585 9933
rect 3589 9929 3595 9933
rect 3599 9929 3604 9933
rect 3560 9928 3604 9929
rect 3564 9924 3570 9928
rect 3574 9924 3580 9928
rect 3584 9924 3590 9928
rect 3594 9924 3600 9928
rect 3560 9923 3604 9924
rect 3560 9919 3565 9923
rect 3569 9919 3575 9923
rect 3579 9919 3585 9923
rect 3589 9919 3595 9923
rect 3599 9919 3604 9923
rect 3560 9918 3604 9919
rect 3564 9914 3570 9918
rect 3574 9914 3580 9918
rect 3584 9914 3590 9918
rect 3594 9914 3600 9918
rect 3560 9913 3604 9914
rect 3560 9909 3565 9913
rect 3569 9909 3575 9913
rect 3579 9909 3585 9913
rect 3589 9909 3595 9913
rect 3599 9909 3604 9913
rect 3560 9908 3604 9909
rect 3564 9904 3570 9908
rect 3574 9904 3580 9908
rect 3584 9904 3590 9908
rect 3594 9904 3600 9908
rect 3560 9903 3604 9904
rect 3560 9899 3565 9903
rect 3569 9899 3575 9903
rect 3579 9899 3585 9903
rect 3589 9899 3595 9903
rect 3599 9899 3604 9903
rect 3560 9898 3604 9899
rect 3564 9894 3570 9898
rect 3574 9894 3580 9898
rect 3584 9894 3590 9898
rect 3594 9894 3600 9898
rect 3560 9893 3604 9894
rect 3560 9889 3565 9893
rect 3569 9889 3575 9893
rect 3579 9889 3585 9893
rect 3589 9889 3595 9893
rect 3599 9889 3604 9893
rect 3560 9888 3604 9889
rect 3564 9884 3570 9888
rect 3574 9884 3580 9888
rect 3584 9884 3590 9888
rect 3594 9884 3600 9888
rect 3560 9883 3604 9884
rect 3560 9879 3565 9883
rect 3569 9879 3575 9883
rect 3579 9879 3585 9883
rect 3589 9879 3595 9883
rect 3599 9879 3604 9883
rect 3560 9878 3604 9879
rect 3564 9874 3570 9878
rect 3574 9874 3580 9878
rect 3584 9874 3590 9878
rect 3594 9874 3600 9878
rect 3560 9873 3604 9874
rect 3560 9869 3565 9873
rect 3569 9869 3575 9873
rect 3579 9869 3585 9873
rect 3589 9869 3595 9873
rect 3599 9869 3604 9873
rect 3560 9868 3604 9869
rect 3564 9864 3570 9868
rect 3574 9864 3580 9868
rect 3584 9864 3590 9868
rect 3594 9864 3600 9868
rect 3869 9949 3874 9953
rect 3878 9949 3884 9953
rect 3888 9949 3894 9953
rect 3898 9949 3904 9953
rect 3908 9949 3913 9953
rect 3869 9948 3913 9949
rect 3873 9944 3879 9948
rect 3883 9944 3889 9948
rect 3893 9944 3899 9948
rect 3903 9944 3909 9948
rect 3869 9943 3913 9944
rect 3869 9939 3874 9943
rect 3878 9939 3884 9943
rect 3888 9939 3894 9943
rect 3898 9939 3904 9943
rect 3908 9939 3913 9943
rect 3869 9938 3913 9939
rect 3873 9934 3879 9938
rect 3883 9934 3889 9938
rect 3893 9934 3899 9938
rect 3903 9934 3909 9938
rect 3869 9933 3913 9934
rect 3869 9929 3874 9933
rect 3878 9929 3884 9933
rect 3888 9929 3894 9933
rect 3898 9929 3904 9933
rect 3908 9929 3913 9933
rect 3869 9928 3913 9929
rect 3873 9924 3879 9928
rect 3883 9924 3889 9928
rect 3893 9924 3899 9928
rect 3903 9924 3909 9928
rect 3869 9923 3913 9924
rect 3869 9919 3874 9923
rect 3878 9919 3884 9923
rect 3888 9919 3894 9923
rect 3898 9919 3904 9923
rect 3908 9919 3913 9923
rect 3869 9918 3913 9919
rect 3873 9914 3879 9918
rect 3883 9914 3889 9918
rect 3893 9914 3899 9918
rect 3903 9914 3909 9918
rect 3869 9913 3913 9914
rect 3869 9909 3874 9913
rect 3878 9909 3884 9913
rect 3888 9909 3894 9913
rect 3898 9909 3904 9913
rect 3908 9909 3913 9913
rect 3869 9908 3913 9909
rect 3873 9904 3879 9908
rect 3883 9904 3889 9908
rect 3893 9904 3899 9908
rect 3903 9904 3909 9908
rect 3869 9903 3913 9904
rect 3869 9899 3874 9903
rect 3878 9899 3884 9903
rect 3888 9899 3894 9903
rect 3898 9899 3904 9903
rect 3908 9899 3913 9903
rect 3869 9898 3913 9899
rect 3873 9894 3879 9898
rect 3883 9894 3889 9898
rect 3893 9894 3899 9898
rect 3903 9894 3909 9898
rect 3869 9893 3913 9894
rect 3869 9889 3874 9893
rect 3878 9889 3884 9893
rect 3888 9889 3894 9893
rect 3898 9889 3904 9893
rect 3908 9889 3913 9893
rect 3869 9888 3913 9889
rect 3873 9884 3879 9888
rect 3883 9884 3889 9888
rect 3893 9884 3899 9888
rect 3903 9884 3909 9888
rect 3869 9883 3913 9884
rect 3869 9879 3874 9883
rect 3878 9879 3884 9883
rect 3888 9879 3894 9883
rect 3898 9879 3904 9883
rect 3908 9879 3913 9883
rect 3869 9878 3913 9879
rect 3873 9874 3879 9878
rect 3883 9874 3889 9878
rect 3893 9874 3899 9878
rect 3903 9874 3909 9878
rect 3869 9873 3913 9874
rect 3869 9869 3874 9873
rect 3878 9869 3884 9873
rect 3888 9869 3894 9873
rect 3898 9869 3904 9873
rect 3908 9869 3913 9873
rect 3869 9868 3913 9869
rect 3873 9864 3879 9868
rect 3883 9864 3889 9868
rect 3893 9864 3899 9868
rect 3903 9864 3909 9868
rect 1836 9827 1840 9831
rect 1829 9826 1869 9827
rect 2145 9827 2149 9831
rect 2138 9826 2178 9827
rect 2454 9827 2458 9831
rect 2447 9826 2487 9827
rect 2763 9827 2767 9831
rect 2756 9826 2796 9827
rect 3072 9827 3076 9831
rect 3065 9826 3105 9827
rect 3999 9827 4003 9831
rect 3992 9826 4032 9827
rect 1829 9823 1869 9824
rect 1829 9818 1869 9819
rect 2138 9823 2178 9824
rect 2138 9818 2178 9819
rect 2447 9823 2487 9824
rect 2447 9818 2487 9819
rect 2756 9823 2796 9824
rect 2756 9818 2796 9819
rect 3065 9823 3105 9824
rect 3065 9818 3105 9819
rect 3992 9823 4032 9824
rect 3992 9818 4032 9819
rect 1829 9815 1869 9816
rect 1836 9811 1840 9815
rect 1829 9810 1869 9811
rect 2138 9815 2178 9816
rect 1829 9807 1869 9808
rect 1829 9802 1869 9803
rect 1829 9799 1869 9800
rect 1836 9795 1840 9799
rect 1829 9794 1869 9795
rect 1829 9791 1869 9792
rect 1829 9786 1869 9787
rect 2145 9811 2149 9815
rect 2138 9810 2178 9811
rect 2447 9815 2487 9816
rect 2138 9807 2178 9808
rect 2138 9802 2178 9803
rect 2138 9799 2178 9800
rect 2145 9795 2149 9799
rect 2138 9794 2178 9795
rect 2138 9791 2178 9792
rect 2138 9786 2178 9787
rect 2454 9811 2458 9815
rect 2447 9810 2487 9811
rect 2756 9815 2796 9816
rect 2447 9807 2487 9808
rect 2447 9802 2487 9803
rect 2447 9799 2487 9800
rect 2454 9795 2458 9799
rect 2447 9794 2487 9795
rect 2447 9791 2487 9792
rect 2447 9786 2487 9787
rect 2763 9811 2767 9815
rect 2756 9810 2796 9811
rect 3065 9815 3105 9816
rect 2756 9807 2796 9808
rect 2756 9802 2796 9803
rect 2756 9799 2796 9800
rect 2763 9795 2767 9799
rect 2756 9794 2796 9795
rect 2756 9791 2796 9792
rect 2756 9786 2796 9787
rect 3072 9811 3076 9815
rect 3065 9810 3105 9811
rect 3992 9815 4032 9816
rect 3065 9807 3105 9808
rect 3065 9802 3105 9803
rect 3065 9799 3105 9800
rect 3072 9795 3076 9799
rect 3065 9794 3105 9795
rect 3065 9791 3105 9792
rect 3065 9786 3105 9787
rect 3999 9811 4003 9815
rect 3992 9810 4032 9811
rect 3992 9807 4032 9808
rect 3992 9802 4032 9803
rect 3992 9799 4032 9800
rect 3999 9795 4003 9799
rect 3992 9794 4032 9795
rect 3992 9791 4032 9792
rect 3992 9786 4032 9787
rect 1829 9783 1869 9784
rect 1836 9779 1840 9783
rect 2138 9783 2178 9784
rect 2145 9779 2149 9783
rect 2447 9783 2487 9784
rect 2454 9779 2458 9783
rect 2756 9783 2796 9784
rect 2763 9779 2767 9783
rect 3065 9783 3105 9784
rect 3072 9779 3076 9783
rect 3992 9783 4032 9784
rect 3999 9779 4003 9783
rect 422 6332 423 6339
rect 427 6332 428 6339
rect 422 6328 428 6332
rect 422 6280 423 6328
rect 427 6280 428 6328
rect 430 6280 431 6339
rect 435 6280 436 6339
rect 438 6328 444 6339
rect 438 6280 439 6328
rect 443 6280 444 6328
rect 446 6280 447 6339
rect 451 6280 452 6339
rect 454 6280 459 6339
rect 463 6332 464 6339
rect 468 6332 469 6339
rect 463 6328 469 6332
rect 463 6280 464 6328
rect 468 6280 469 6328
rect 471 6280 472 6339
rect 476 6280 477 6339
rect 479 6328 485 6339
rect 479 6280 480 6328
rect 484 6280 485 6328
rect 487 6280 488 6339
rect 492 6280 493 6339
rect 495 6280 502 6339
rect 506 6332 507 6339
rect 511 6332 512 6339
rect 506 6328 512 6332
rect 506 6280 507 6328
rect 511 6280 512 6328
rect 514 6280 515 6339
rect 519 6280 520 6339
rect 522 6332 523 6339
rect 527 6332 528 6339
rect 522 6328 528 6332
rect 522 6280 523 6328
rect 527 6280 528 6328
rect 530 6280 531 6339
rect 535 6280 536 6339
rect 538 6280 541 6339
rect 545 6332 546 6339
rect 550 6332 551 6339
rect 545 6328 551 6332
rect 545 6299 546 6328
rect 550 6299 551 6328
rect 553 6299 554 6339
rect 558 6299 559 6339
rect 561 6332 562 6339
rect 566 6332 567 6339
rect 561 6328 567 6332
rect 561 6299 562 6328
rect 566 6299 567 6328
rect 569 6299 570 6339
rect 574 6299 575 6339
rect 577 6332 578 6339
rect 582 6332 583 6339
rect 577 6328 583 6332
rect 577 6299 578 6328
rect 582 6299 583 6328
rect 585 6299 586 6339
rect 590 6299 591 6339
rect 593 6332 594 6339
rect 593 6328 598 6332
rect 593 6299 594 6328
rect 2855 9299 2856 9303
rect 2858 9299 2861 9303
rect 2863 9299 2864 9303
rect 2876 9299 2877 9303
rect 2879 9299 2880 9303
rect 2892 9299 2893 9303
rect 2895 9299 2898 9303
rect 2900 9299 2901 9303
rect 2918 9299 2919 9303
rect 2921 9299 2922 9303
rect 2934 9299 2935 9303
rect 2937 9299 2938 9303
rect 2950 9299 2951 9303
rect 2953 9299 2956 9303
rect 2958 9299 2959 9303
rect 2971 9299 2972 9303
rect 2974 9299 2975 9303
rect 2987 9299 2988 9303
rect 2990 9299 2993 9303
rect 2995 9299 2996 9303
rect 3008 9299 3009 9303
rect 3011 9299 3012 9303
rect 3024 9299 3025 9303
rect 3027 9299 3030 9303
rect 3032 9299 3033 9303
rect 3050 9299 3051 9303
rect 3053 9299 3054 9303
rect 3066 9299 3067 9303
rect 3069 9299 3070 9303
rect 3082 9299 3083 9303
rect 3085 9299 3088 9303
rect 3090 9299 3091 9303
rect 3103 9299 3104 9303
rect 3106 9299 3107 9303
rect 3119 9299 3120 9303
rect 3122 9299 3125 9303
rect 3127 9299 3128 9303
rect 3140 9299 3141 9303
rect 3143 9299 3144 9303
rect 3156 9299 3157 9303
rect 3159 9299 3162 9303
rect 3164 9299 3165 9303
rect 3182 9299 3183 9303
rect 3185 9299 3186 9303
rect 3198 9299 3199 9303
rect 3201 9299 3202 9303
rect 3214 9299 3215 9303
rect 3217 9299 3220 9303
rect 3222 9299 3223 9303
rect 3235 9299 3236 9303
rect 3238 9299 3239 9303
rect 3251 9299 3252 9303
rect 3254 9299 3257 9303
rect 3259 9299 3260 9303
rect 3272 9299 3273 9303
rect 3275 9299 3276 9303
rect 3288 9299 3289 9303
rect 3291 9299 3294 9303
rect 3296 9299 3297 9303
rect 3314 9299 3315 9303
rect 3317 9299 3318 9303
rect 3330 9299 3331 9303
rect 3333 9299 3334 9303
rect 3346 9299 3347 9303
rect 3349 9299 3352 9303
rect 3354 9299 3355 9303
rect 3367 9299 3368 9303
rect 3370 9299 3371 9303
rect 3800 9299 3801 9303
rect 3803 9299 3806 9303
rect 3808 9299 3809 9303
rect 3821 9299 3822 9303
rect 3824 9299 3825 9303
rect 3837 9299 3838 9303
rect 3840 9299 3843 9303
rect 3845 9299 3846 9303
rect 3863 9299 3864 9303
rect 3866 9299 3867 9303
rect 3879 9299 3880 9303
rect 3882 9299 3883 9303
rect 3895 9299 3896 9303
rect 3898 9299 3901 9303
rect 3903 9299 3904 9303
rect 3916 9299 3917 9303
rect 3919 9299 3920 9303
rect 3932 9299 3933 9303
rect 3935 9299 3938 9303
rect 3940 9299 3941 9303
rect 3953 9299 3954 9303
rect 3956 9299 3957 9303
rect 3969 9299 3970 9303
rect 3972 9299 3975 9303
rect 3977 9299 3978 9303
rect 3995 9299 3996 9303
rect 3998 9299 3999 9303
rect 4011 9299 4012 9303
rect 4014 9299 4015 9303
rect 4027 9299 4028 9303
rect 4030 9299 4033 9303
rect 4035 9299 4036 9303
rect 4048 9299 4049 9303
rect 4051 9299 4052 9303
rect 4064 9299 4065 9303
rect 4067 9299 4070 9303
rect 4072 9299 4073 9303
rect 4085 9299 4086 9303
rect 4088 9299 4089 9303
rect 4101 9299 4102 9303
rect 4104 9299 4107 9303
rect 4109 9299 4110 9303
rect 4127 9299 4128 9303
rect 4130 9299 4131 9303
rect 4143 9299 4144 9303
rect 4146 9299 4147 9303
rect 4159 9299 4160 9303
rect 4162 9299 4165 9303
rect 4167 9299 4168 9303
rect 4180 9299 4181 9303
rect 4183 9299 4184 9303
rect 4196 9299 4197 9303
rect 4199 9299 4202 9303
rect 4204 9299 4205 9303
rect 4217 9299 4218 9303
rect 4220 9299 4221 9303
rect 4233 9299 4234 9303
rect 4236 9299 4239 9303
rect 4241 9299 4242 9303
rect 4259 9299 4260 9303
rect 4262 9299 4263 9303
rect 4275 9299 4276 9303
rect 4278 9299 4279 9303
rect 4291 9299 4292 9303
rect 4294 9299 4297 9303
rect 4299 9299 4300 9303
rect 4312 9299 4313 9303
rect 4315 9299 4316 9303
rect 2503 9266 2504 9270
rect 2506 9266 2509 9270
rect 2511 9266 2512 9270
rect 2524 9266 2525 9270
rect 2527 9266 2528 9270
rect 2540 9266 2541 9270
rect 2543 9266 2546 9270
rect 2548 9266 2549 9270
rect 2566 9266 2567 9270
rect 2569 9266 2570 9270
rect 2582 9266 2583 9270
rect 2585 9266 2586 9270
rect 2598 9266 2599 9270
rect 2601 9266 2604 9270
rect 2606 9266 2607 9270
rect 2619 9266 2620 9270
rect 2622 9266 2623 9270
rect 3448 9266 3449 9270
rect 3451 9266 3454 9270
rect 3456 9266 3457 9270
rect 3469 9266 3470 9270
rect 3472 9266 3473 9270
rect 3485 9266 3486 9270
rect 3488 9266 3491 9270
rect 3493 9266 3494 9270
rect 3511 9266 3512 9270
rect 3514 9266 3515 9270
rect 3527 9266 3528 9270
rect 3530 9266 3531 9270
rect 3543 9266 3544 9270
rect 3546 9266 3549 9270
rect 3551 9266 3552 9270
rect 3564 9266 3565 9270
rect 3567 9266 3568 9270
rect 2627 9229 2628 9233
rect 2630 9229 2631 9233
rect 3034 9233 3035 9237
rect 3037 9233 3038 9237
rect 3058 9229 3061 9233
rect 3063 9229 3066 9233
rect 3068 9229 3069 9233
rect 3115 9233 3116 9237
rect 3118 9233 3119 9237
rect 3139 9229 3142 9233
rect 3144 9229 3147 9233
rect 3149 9229 3150 9233
rect 3088 9225 3089 9229
rect 3091 9225 3092 9229
rect 2510 9220 2511 9224
rect 2513 9220 2514 9224
rect 2860 9220 2861 9224
rect 2863 9220 2864 9224
rect 2876 9220 2877 9224
rect 2879 9220 2880 9224
rect 2892 9220 2893 9224
rect 2895 9220 2896 9224
rect 2911 9220 2916 9224
rect 2918 9220 2921 9224
rect 2923 9220 2924 9224
rect 2945 9220 2947 9224
rect 2949 9220 2950 9224
rect 2967 9220 2968 9224
rect 2970 9220 2971 9224
rect 2983 9220 2988 9224
rect 2990 9220 2993 9224
rect 2995 9220 2996 9224
rect 3010 9220 3011 9224
rect 3013 9220 3014 9224
rect 3169 9225 3170 9229
rect 3172 9225 3173 9229
rect 3572 9229 3573 9233
rect 3575 9229 3576 9233
rect 3979 9233 3980 9237
rect 3982 9233 3983 9237
rect 4003 9229 4006 9233
rect 4008 9229 4011 9233
rect 4013 9229 4014 9233
rect 4060 9233 4061 9237
rect 4063 9233 4064 9237
rect 4084 9229 4087 9233
rect 4089 9229 4092 9233
rect 4094 9229 4095 9233
rect 4033 9225 4034 9229
rect 4036 9225 4037 9229
rect 3455 9220 3456 9224
rect 3458 9220 3459 9224
rect 3805 9220 3806 9224
rect 3808 9220 3809 9224
rect 3821 9220 3822 9224
rect 3824 9220 3825 9224
rect 3837 9220 3838 9224
rect 3840 9220 3841 9224
rect 3856 9220 3861 9224
rect 3863 9220 3866 9224
rect 3868 9220 3869 9224
rect 3890 9220 3892 9224
rect 3894 9220 3895 9224
rect 3912 9220 3913 9224
rect 3915 9220 3916 9224
rect 3928 9220 3933 9224
rect 3935 9220 3938 9224
rect 3940 9220 3941 9224
rect 3955 9220 3956 9224
rect 3958 9220 3959 9224
rect 4114 9225 4115 9229
rect 4117 9225 4118 9229
rect 2860 9174 2861 9178
rect 2863 9174 2864 9178
rect 2876 9174 2877 9178
rect 2879 9174 2880 9178
rect 2892 9174 2893 9178
rect 2895 9174 2896 9178
rect 2911 9174 2916 9178
rect 2918 9174 2921 9178
rect 2923 9174 2924 9178
rect 2945 9174 2947 9178
rect 2949 9174 2950 9178
rect 2967 9174 2968 9178
rect 2970 9174 2971 9178
rect 2983 9174 2988 9178
rect 2990 9174 2993 9178
rect 2995 9174 2996 9178
rect 3010 9174 3011 9178
rect 3013 9174 3014 9178
rect 2494 9164 2495 9168
rect 2497 9164 2498 9168
rect 2510 9164 2511 9168
rect 2513 9164 2516 9168
rect 2518 9164 2519 9168
rect 2531 9164 2532 9168
rect 2534 9164 2535 9168
rect 2547 9164 2548 9168
rect 2550 9164 2551 9168
rect 2568 9164 2569 9168
rect 2571 9164 2574 9168
rect 2576 9164 2577 9168
rect 2589 9164 2590 9168
rect 2592 9164 2593 9168
rect 2605 9164 2606 9168
rect 2608 9164 2611 9168
rect 2613 9164 2614 9168
rect 3058 9173 3061 9177
rect 3063 9173 3066 9177
rect 3068 9173 3069 9177
rect 3139 9173 3142 9177
rect 3144 9173 3147 9177
rect 3149 9173 3150 9177
rect 3805 9174 3806 9178
rect 3808 9174 3809 9178
rect 3821 9174 3822 9178
rect 3824 9174 3825 9178
rect 3837 9174 3838 9178
rect 3840 9174 3841 9178
rect 3856 9174 3861 9178
rect 3863 9174 3866 9178
rect 3868 9174 3869 9178
rect 3890 9174 3892 9178
rect 3894 9174 3895 9178
rect 3912 9174 3913 9178
rect 3915 9174 3916 9178
rect 3928 9174 3933 9178
rect 3935 9174 3938 9178
rect 3940 9174 3941 9178
rect 3955 9174 3956 9178
rect 3958 9174 3959 9178
rect 3439 9164 3440 9168
rect 3442 9164 3443 9168
rect 3455 9164 3456 9168
rect 3458 9164 3461 9168
rect 3463 9164 3464 9168
rect 3476 9164 3477 9168
rect 3479 9164 3480 9168
rect 3492 9164 3493 9168
rect 3495 9164 3496 9168
rect 3513 9164 3514 9168
rect 3516 9164 3519 9168
rect 3521 9164 3522 9168
rect 3534 9164 3535 9168
rect 3537 9164 3538 9168
rect 3550 9164 3551 9168
rect 3553 9164 3556 9168
rect 3558 9164 3559 9168
rect 4003 9173 4006 9177
rect 4008 9173 4011 9177
rect 4013 9173 4014 9177
rect 4084 9173 4087 9177
rect 4089 9173 4092 9177
rect 4094 9173 4095 9177
rect 3058 9097 3061 9101
rect 3063 9097 3066 9101
rect 3068 9097 3069 9101
rect 3139 9101 3140 9105
rect 3142 9101 3143 9105
rect 3163 9097 3166 9101
rect 3168 9097 3171 9101
rect 3173 9097 3174 9101
rect 3088 9093 3089 9097
rect 3091 9093 3092 9097
rect 2860 9088 2861 9092
rect 2863 9088 2864 9092
rect 2876 9088 2877 9092
rect 2879 9088 2880 9092
rect 2892 9088 2893 9092
rect 2895 9088 2896 9092
rect 2911 9088 2916 9092
rect 2918 9088 2921 9092
rect 2923 9088 2924 9092
rect 2945 9088 2947 9092
rect 2949 9088 2950 9092
rect 2967 9088 2968 9092
rect 2970 9088 2971 9092
rect 2983 9088 2988 9092
rect 2990 9088 2993 9092
rect 2995 9088 2996 9092
rect 3010 9088 3011 9092
rect 3013 9088 3014 9092
rect 3193 9093 3194 9097
rect 3196 9093 3197 9097
rect 3370 9072 3371 9076
rect 3373 9072 3374 9076
rect 3394 9068 3397 9072
rect 3399 9068 3402 9072
rect 3404 9068 3405 9072
rect 3424 9064 3425 9068
rect 3427 9064 3428 9068
rect 4003 9097 4006 9101
rect 4008 9097 4011 9101
rect 4013 9097 4014 9101
rect 4084 9101 4085 9105
rect 4087 9101 4088 9105
rect 4108 9097 4111 9101
rect 4113 9097 4116 9101
rect 4118 9097 4119 9101
rect 4033 9093 4034 9097
rect 4036 9093 4037 9097
rect 3805 9088 3806 9092
rect 3808 9088 3809 9092
rect 3821 9088 3822 9092
rect 3824 9088 3825 9092
rect 3837 9088 3838 9092
rect 3840 9088 3841 9092
rect 3856 9088 3861 9092
rect 3863 9088 3866 9092
rect 3868 9088 3869 9092
rect 3890 9088 3892 9092
rect 3894 9088 3895 9092
rect 3912 9088 3913 9092
rect 3915 9088 3916 9092
rect 3928 9088 3933 9092
rect 3935 9088 3938 9092
rect 3940 9088 3941 9092
rect 3955 9088 3956 9092
rect 3958 9088 3959 9092
rect 4138 9093 4139 9097
rect 4141 9093 4142 9097
rect 2860 9042 2861 9046
rect 2863 9042 2864 9046
rect 2876 9042 2877 9046
rect 2879 9042 2880 9046
rect 2892 9042 2893 9046
rect 2895 9042 2896 9046
rect 2911 9042 2916 9046
rect 2918 9042 2921 9046
rect 2923 9042 2924 9046
rect 2945 9042 2947 9046
rect 2949 9042 2950 9046
rect 2967 9042 2968 9046
rect 2970 9042 2971 9046
rect 2983 9042 2988 9046
rect 2990 9042 2993 9046
rect 2995 9042 2996 9046
rect 3010 9042 3011 9046
rect 3013 9042 3014 9046
rect 3058 9042 3061 9046
rect 3063 9042 3066 9046
rect 3068 9042 3069 9046
rect 3163 9042 3166 9046
rect 3168 9042 3171 9046
rect 3173 9042 3174 9046
rect 3556 9033 3557 9045
rect 3559 9033 3560 9045
rect 3609 9033 3610 9045
rect 3612 9033 3613 9045
rect 3805 9042 3806 9046
rect 3808 9042 3809 9046
rect 3821 9042 3822 9046
rect 3824 9042 3825 9046
rect 3837 9042 3838 9046
rect 3840 9042 3841 9046
rect 3856 9042 3861 9046
rect 3863 9042 3866 9046
rect 3868 9042 3869 9046
rect 3890 9042 3892 9046
rect 3894 9042 3895 9046
rect 3912 9042 3913 9046
rect 3915 9042 3916 9046
rect 3928 9042 3933 9046
rect 3935 9042 3938 9046
rect 3940 9042 3941 9046
rect 3955 9042 3956 9046
rect 3958 9042 3959 9046
rect 4003 9042 4006 9046
rect 4008 9042 4011 9046
rect 4013 9042 4014 9046
rect 4108 9042 4111 9046
rect 4113 9042 4116 9046
rect 4118 9042 4119 9046
rect 3394 9008 3397 9012
rect 3399 9008 3402 9012
rect 3404 9008 3405 9012
rect 3058 8965 3061 8969
rect 3063 8965 3066 8969
rect 3068 8965 3069 8969
rect 3115 8969 3116 8973
rect 3118 8969 3119 8973
rect 3139 8965 3142 8969
rect 3144 8965 3147 8969
rect 3149 8965 3150 8969
rect 3205 8969 3206 8973
rect 3208 8969 3209 8973
rect 3229 8965 3232 8969
rect 3234 8965 3237 8969
rect 3239 8965 3240 8969
rect 3088 8961 3089 8965
rect 3091 8961 3092 8965
rect 2860 8956 2861 8960
rect 2863 8956 2864 8960
rect 2876 8956 2877 8960
rect 2879 8956 2880 8960
rect 2892 8956 2893 8960
rect 2895 8956 2896 8960
rect 2911 8956 2916 8960
rect 2918 8956 2921 8960
rect 2923 8956 2924 8960
rect 2945 8956 2947 8960
rect 2949 8956 2950 8960
rect 2967 8956 2968 8960
rect 2970 8956 2971 8960
rect 2983 8956 2988 8960
rect 2990 8956 2993 8960
rect 2995 8956 2996 8960
rect 3010 8956 3011 8960
rect 3013 8956 3014 8960
rect 3169 8961 3170 8965
rect 3172 8961 3173 8965
rect 3259 8961 3260 8965
rect 3262 8961 3263 8965
rect 3348 8942 3349 8946
rect 3351 8942 3352 8946
rect 3370 8942 3371 8946
rect 3373 8942 3374 8946
rect 3394 8938 3397 8942
rect 3399 8938 3402 8942
rect 3404 8938 3405 8942
rect 3424 8934 3425 8938
rect 3427 8934 3428 8938
rect 4003 8965 4006 8969
rect 4008 8965 4011 8969
rect 4013 8965 4014 8969
rect 4060 8969 4061 8973
rect 4063 8969 4064 8973
rect 4084 8965 4087 8969
rect 4089 8965 4092 8969
rect 4094 8965 4095 8969
rect 4150 8969 4151 8973
rect 4153 8969 4154 8973
rect 4174 8965 4177 8969
rect 4179 8965 4182 8969
rect 4184 8965 4185 8969
rect 4033 8961 4034 8965
rect 4036 8961 4037 8965
rect 3805 8956 3806 8960
rect 3808 8956 3809 8960
rect 3821 8956 3822 8960
rect 3824 8956 3825 8960
rect 3837 8956 3838 8960
rect 3840 8956 3841 8960
rect 3856 8956 3861 8960
rect 3863 8956 3866 8960
rect 3868 8956 3869 8960
rect 3890 8956 3892 8960
rect 3894 8956 3895 8960
rect 3912 8956 3913 8960
rect 3915 8956 3916 8960
rect 3928 8956 3933 8960
rect 3935 8956 3938 8960
rect 3940 8956 3941 8960
rect 3955 8956 3956 8960
rect 3958 8956 3959 8960
rect 4114 8961 4115 8965
rect 4117 8961 4118 8965
rect 4204 8961 4205 8965
rect 4207 8961 4208 8965
rect 2860 8910 2861 8914
rect 2863 8910 2864 8914
rect 2876 8910 2877 8914
rect 2879 8910 2880 8914
rect 2892 8910 2893 8914
rect 2895 8910 2896 8914
rect 2911 8910 2916 8914
rect 2918 8910 2921 8914
rect 2923 8910 2924 8914
rect 2945 8910 2947 8914
rect 2949 8910 2950 8914
rect 2967 8910 2968 8914
rect 2970 8910 2971 8914
rect 2983 8910 2988 8914
rect 2990 8910 2993 8914
rect 2995 8910 2996 8914
rect 3010 8910 3011 8914
rect 3013 8910 3014 8914
rect 3058 8907 3061 8911
rect 3063 8907 3066 8911
rect 3068 8907 3069 8911
rect 3139 8907 3142 8911
rect 3144 8907 3147 8911
rect 3149 8907 3150 8911
rect 3229 8907 3232 8911
rect 3234 8907 3237 8911
rect 3239 8907 3240 8911
rect 3462 8903 3463 8915
rect 3465 8903 3466 8915
rect 3515 8903 3516 8915
rect 3518 8903 3519 8915
rect 3805 8910 3806 8914
rect 3808 8910 3809 8914
rect 3821 8910 3822 8914
rect 3824 8910 3825 8914
rect 3837 8910 3838 8914
rect 3840 8910 3841 8914
rect 3856 8910 3861 8914
rect 3863 8910 3866 8914
rect 3868 8910 3869 8914
rect 3890 8910 3892 8914
rect 3894 8910 3895 8914
rect 3912 8910 3913 8914
rect 3915 8910 3916 8914
rect 3928 8910 3933 8914
rect 3935 8910 3938 8914
rect 3940 8910 3941 8914
rect 3955 8910 3956 8914
rect 3958 8910 3959 8914
rect 4003 8907 4006 8911
rect 4008 8907 4011 8911
rect 4013 8907 4014 8911
rect 4084 8907 4087 8911
rect 4089 8907 4092 8911
rect 4094 8907 4095 8911
rect 4174 8907 4177 8911
rect 4179 8907 4182 8911
rect 4184 8907 4185 8911
rect 3394 8878 3397 8882
rect 3399 8878 3402 8882
rect 3404 8878 3405 8882
rect 3058 8833 3061 8837
rect 3063 8833 3066 8837
rect 3068 8833 3069 8837
rect 3088 8829 3089 8833
rect 3091 8829 3092 8833
rect 2860 8824 2861 8828
rect 2863 8824 2864 8828
rect 2876 8824 2877 8828
rect 2879 8824 2880 8828
rect 2892 8824 2893 8828
rect 2895 8824 2896 8828
rect 2911 8824 2916 8828
rect 2918 8824 2921 8828
rect 2923 8824 2924 8828
rect 2945 8824 2947 8828
rect 2949 8824 2950 8828
rect 2967 8824 2968 8828
rect 2970 8824 2971 8828
rect 2983 8824 2988 8828
rect 2990 8824 2993 8828
rect 2995 8824 2996 8828
rect 3010 8824 3011 8828
rect 3013 8824 3014 8828
rect 4003 8833 4006 8837
rect 4008 8833 4011 8837
rect 4013 8833 4014 8837
rect 4033 8829 4034 8833
rect 4036 8829 4037 8833
rect 3805 8824 3806 8828
rect 3808 8824 3809 8828
rect 3821 8824 3822 8828
rect 3824 8824 3825 8828
rect 3837 8824 3838 8828
rect 3840 8824 3841 8828
rect 3856 8824 3861 8828
rect 3863 8824 3866 8828
rect 3868 8824 3869 8828
rect 3890 8824 3892 8828
rect 3894 8824 3895 8828
rect 3912 8824 3913 8828
rect 3915 8824 3916 8828
rect 3928 8824 3933 8828
rect 3935 8824 3938 8828
rect 3940 8824 3941 8828
rect 3955 8824 3956 8828
rect 3958 8824 3959 8828
rect 2860 8778 2861 8782
rect 2863 8778 2864 8782
rect 2876 8778 2877 8782
rect 2879 8778 2880 8782
rect 2892 8778 2893 8782
rect 2895 8778 2896 8782
rect 2911 8778 2916 8782
rect 2918 8778 2921 8782
rect 2923 8778 2924 8782
rect 2945 8778 2947 8782
rect 2949 8778 2950 8782
rect 2967 8778 2968 8782
rect 2970 8778 2971 8782
rect 2983 8778 2988 8782
rect 2990 8778 2993 8782
rect 2995 8778 2996 8782
rect 3010 8778 3011 8782
rect 3013 8778 3014 8782
rect 3094 8778 3095 8782
rect 3097 8778 3098 8782
rect 3102 8778 3108 8782
rect 3112 8778 3113 8782
rect 3115 8778 3116 8782
rect 3137 8778 3138 8782
rect 3140 8778 3141 8782
rect 3153 8778 3154 8782
rect 3156 8778 3157 8782
rect 3172 8778 3177 8782
rect 3179 8778 3182 8782
rect 3184 8778 3185 8782
rect 3206 8778 3208 8782
rect 3210 8778 3211 8782
rect 3228 8778 3229 8782
rect 3231 8778 3232 8782
rect 3244 8778 3249 8782
rect 3251 8778 3254 8782
rect 3256 8778 3257 8782
rect 3271 8778 3272 8782
rect 3274 8778 3275 8782
rect 2371 8764 2372 8768
rect 2374 8764 2377 8768
rect 2379 8764 2380 8768
rect 2392 8764 2393 8768
rect 2395 8764 2396 8768
rect 2408 8764 2409 8768
rect 2411 8764 2414 8768
rect 2416 8764 2417 8768
rect 2434 8764 2435 8768
rect 2437 8764 2438 8768
rect 2450 8764 2451 8768
rect 2453 8764 2454 8768
rect 2466 8764 2467 8768
rect 2469 8764 2472 8768
rect 2474 8764 2475 8768
rect 2487 8764 2488 8768
rect 2490 8764 2491 8768
rect 2503 8764 2504 8768
rect 2506 8764 2509 8768
rect 2511 8764 2512 8768
rect 2524 8764 2525 8768
rect 2527 8764 2528 8768
rect 2540 8764 2541 8768
rect 2543 8764 2546 8768
rect 2548 8764 2549 8768
rect 2566 8764 2567 8768
rect 2569 8764 2570 8768
rect 2582 8764 2583 8768
rect 2585 8764 2586 8768
rect 2598 8764 2599 8768
rect 2601 8764 2604 8768
rect 2606 8764 2607 8768
rect 2619 8764 2620 8768
rect 2622 8764 2623 8768
rect 2635 8764 2636 8768
rect 2638 8764 2641 8768
rect 2643 8764 2644 8768
rect 2656 8764 2657 8768
rect 2659 8764 2660 8768
rect 2672 8764 2673 8768
rect 2675 8764 2678 8768
rect 2680 8764 2681 8768
rect 2698 8764 2699 8768
rect 2701 8764 2702 8768
rect 2714 8764 2715 8768
rect 2717 8764 2718 8768
rect 2730 8764 2731 8768
rect 2733 8764 2736 8768
rect 2738 8764 2739 8768
rect 2751 8764 2752 8768
rect 2754 8764 2755 8768
rect 3058 8771 3061 8775
rect 3063 8771 3066 8775
rect 3068 8771 3069 8775
rect 3805 8778 3806 8782
rect 3808 8778 3809 8782
rect 3821 8778 3822 8782
rect 3824 8778 3825 8782
rect 3837 8778 3838 8782
rect 3840 8778 3841 8782
rect 3856 8778 3861 8782
rect 3863 8778 3866 8782
rect 3868 8778 3869 8782
rect 3890 8778 3892 8782
rect 3894 8778 3895 8782
rect 3912 8778 3913 8782
rect 3915 8778 3916 8782
rect 3928 8778 3933 8782
rect 3935 8778 3938 8782
rect 3940 8778 3941 8782
rect 3955 8778 3956 8782
rect 3958 8778 3959 8782
rect 4039 8778 4040 8782
rect 4042 8778 4043 8782
rect 4047 8778 4053 8782
rect 4057 8778 4058 8782
rect 4060 8778 4061 8782
rect 4082 8778 4083 8782
rect 4085 8778 4086 8782
rect 4098 8778 4099 8782
rect 4101 8778 4102 8782
rect 4117 8778 4122 8782
rect 4124 8778 4127 8782
rect 4129 8778 4130 8782
rect 4151 8778 4153 8782
rect 4155 8778 4156 8782
rect 4173 8778 4174 8782
rect 4176 8778 4177 8782
rect 4189 8778 4194 8782
rect 4196 8778 4199 8782
rect 4201 8778 4202 8782
rect 4216 8778 4217 8782
rect 4219 8778 4220 8782
rect 3316 8764 3317 8768
rect 3319 8764 3322 8768
rect 3324 8764 3325 8768
rect 3337 8764 3338 8768
rect 3340 8764 3341 8768
rect 3353 8764 3354 8768
rect 3356 8764 3359 8768
rect 3361 8764 3362 8768
rect 3379 8764 3380 8768
rect 3382 8764 3383 8768
rect 3395 8764 3396 8768
rect 3398 8764 3399 8768
rect 3411 8764 3412 8768
rect 3414 8764 3417 8768
rect 3419 8764 3420 8768
rect 3432 8764 3433 8768
rect 3435 8764 3436 8768
rect 3448 8764 3449 8768
rect 3451 8764 3454 8768
rect 3456 8764 3457 8768
rect 3469 8764 3470 8768
rect 3472 8764 3473 8768
rect 3485 8764 3486 8768
rect 3488 8764 3491 8768
rect 3493 8764 3494 8768
rect 3511 8764 3512 8768
rect 3514 8764 3515 8768
rect 3527 8764 3528 8768
rect 3530 8764 3531 8768
rect 3543 8764 3544 8768
rect 3546 8764 3549 8768
rect 3551 8764 3552 8768
rect 3564 8764 3565 8768
rect 3567 8764 3568 8768
rect 3580 8764 3581 8768
rect 3583 8764 3586 8768
rect 3588 8764 3589 8768
rect 3601 8764 3602 8768
rect 3604 8764 3605 8768
rect 3617 8764 3618 8768
rect 3620 8764 3623 8768
rect 3625 8764 3626 8768
rect 3643 8764 3644 8768
rect 3646 8764 3647 8768
rect 3659 8764 3660 8768
rect 3662 8764 3663 8768
rect 3675 8764 3676 8768
rect 3678 8764 3681 8768
rect 3683 8764 3684 8768
rect 3696 8764 3697 8768
rect 3699 8764 3700 8768
rect 4003 8771 4006 8775
rect 4008 8771 4011 8775
rect 4013 8771 4014 8775
rect 2486 8720 2487 8724
rect 2489 8720 2490 8724
rect 2510 8720 2511 8724
rect 2513 8720 2514 8724
rect 3284 8724 3288 8725
rect 3284 8721 3288 8722
rect 3431 8720 3432 8724
rect 3434 8720 3435 8724
rect 3455 8720 3456 8724
rect 3458 8720 3459 8724
rect 4229 8724 4233 8725
rect 4229 8721 4233 8722
rect 2506 8707 2507 8711
rect 2509 8707 2510 8711
rect 3451 8707 3452 8711
rect 3454 8707 3455 8711
rect 2498 8695 2502 8696
rect 2498 8692 2502 8693
rect 3443 8695 3447 8696
rect 3443 8692 3447 8693
rect 2486 8684 2487 8688
rect 2489 8684 2490 8688
rect 2510 8684 2511 8688
rect 2513 8684 2514 8688
rect 3431 8684 3432 8688
rect 3434 8684 3435 8688
rect 3455 8684 3456 8688
rect 3458 8684 3459 8688
rect 3154 8652 3155 8656
rect 3157 8652 3160 8656
rect 3162 8652 3163 8656
rect 3175 8652 3176 8656
rect 3178 8652 3179 8656
rect 3191 8652 3192 8656
rect 3194 8652 3197 8656
rect 3199 8652 3200 8656
rect 3217 8652 3218 8656
rect 3220 8652 3221 8656
rect 3233 8652 3234 8656
rect 3236 8652 3237 8656
rect 3249 8652 3250 8656
rect 3252 8652 3255 8656
rect 3257 8652 3258 8656
rect 3270 8652 3271 8656
rect 3273 8652 3274 8656
rect 4099 8652 4100 8656
rect 4102 8652 4105 8656
rect 4107 8652 4108 8656
rect 4120 8652 4121 8656
rect 4123 8652 4124 8656
rect 4136 8652 4137 8656
rect 4139 8652 4142 8656
rect 4144 8652 4145 8656
rect 4162 8652 4163 8656
rect 4165 8652 4166 8656
rect 4178 8652 4179 8656
rect 4181 8652 4182 8656
rect 4194 8652 4195 8656
rect 4197 8652 4200 8656
rect 4202 8652 4203 8656
rect 4215 8652 4216 8656
rect 4218 8652 4219 8656
rect 2371 8622 2372 8626
rect 2374 8622 2377 8626
rect 2379 8622 2380 8626
rect 2392 8622 2393 8626
rect 2395 8622 2396 8626
rect 2408 8622 2409 8626
rect 2411 8622 2414 8626
rect 2416 8622 2417 8626
rect 2434 8622 2435 8626
rect 2437 8622 2438 8626
rect 2450 8622 2451 8626
rect 2453 8622 2454 8626
rect 2466 8622 2467 8626
rect 2469 8622 2472 8626
rect 2474 8622 2475 8626
rect 2487 8622 2488 8626
rect 2490 8622 2491 8626
rect 2503 8622 2504 8626
rect 2506 8622 2509 8626
rect 2511 8622 2512 8626
rect 2524 8622 2525 8626
rect 2527 8622 2528 8626
rect 2540 8622 2541 8626
rect 2543 8622 2546 8626
rect 2548 8622 2549 8626
rect 2566 8622 2567 8626
rect 2569 8622 2570 8626
rect 2582 8622 2583 8626
rect 2585 8622 2586 8626
rect 2598 8622 2599 8626
rect 2601 8622 2604 8626
rect 2606 8622 2607 8626
rect 2619 8622 2620 8626
rect 2622 8622 2623 8626
rect 2635 8622 2636 8626
rect 2638 8622 2641 8626
rect 2643 8622 2644 8626
rect 2656 8622 2657 8626
rect 2659 8622 2660 8626
rect 2672 8622 2673 8626
rect 2675 8622 2678 8626
rect 2680 8622 2681 8626
rect 2698 8622 2699 8626
rect 2701 8622 2702 8626
rect 2714 8622 2715 8626
rect 2717 8622 2718 8626
rect 2730 8622 2731 8626
rect 2733 8622 2736 8626
rect 2738 8622 2739 8626
rect 2751 8622 2752 8626
rect 2754 8622 2755 8626
rect 3316 8622 3317 8626
rect 3319 8622 3322 8626
rect 3324 8622 3325 8626
rect 3337 8622 3338 8626
rect 3340 8622 3341 8626
rect 3353 8622 3354 8626
rect 3356 8622 3359 8626
rect 3361 8622 3362 8626
rect 3379 8622 3380 8626
rect 3382 8622 3383 8626
rect 3395 8622 3396 8626
rect 3398 8622 3399 8626
rect 3411 8622 3412 8626
rect 3414 8622 3417 8626
rect 3419 8622 3420 8626
rect 3432 8622 3433 8626
rect 3435 8622 3436 8626
rect 3448 8622 3449 8626
rect 3451 8622 3454 8626
rect 3456 8622 3457 8626
rect 3469 8622 3470 8626
rect 3472 8622 3473 8626
rect 3485 8622 3486 8626
rect 3488 8622 3491 8626
rect 3493 8622 3494 8626
rect 3511 8622 3512 8626
rect 3514 8622 3515 8626
rect 3527 8622 3528 8626
rect 3530 8622 3531 8626
rect 3543 8622 3544 8626
rect 3546 8622 3549 8626
rect 3551 8622 3552 8626
rect 3564 8622 3565 8626
rect 3567 8622 3568 8626
rect 3580 8622 3581 8626
rect 3583 8622 3586 8626
rect 3588 8622 3589 8626
rect 3601 8622 3602 8626
rect 3604 8622 3605 8626
rect 3617 8622 3618 8626
rect 3620 8622 3623 8626
rect 3625 8622 3626 8626
rect 3643 8622 3644 8626
rect 3646 8622 3647 8626
rect 3659 8622 3660 8626
rect 3662 8622 3663 8626
rect 3675 8622 3676 8626
rect 3678 8622 3681 8626
rect 3683 8622 3684 8626
rect 3696 8622 3697 8626
rect 3699 8622 3700 8626
rect 3296 8578 3300 8579
rect 3296 8575 3300 8576
rect 4241 8578 4245 8579
rect 4241 8575 4245 8576
rect 3154 8566 3155 8570
rect 3157 8566 3160 8570
rect 3162 8566 3163 8570
rect 3175 8566 3176 8570
rect 3178 8566 3179 8570
rect 3191 8566 3192 8570
rect 3194 8566 3197 8570
rect 3199 8566 3200 8570
rect 3217 8566 3218 8570
rect 3220 8566 3221 8570
rect 3233 8566 3234 8570
rect 3236 8566 3237 8570
rect 3249 8566 3250 8570
rect 3252 8566 3255 8570
rect 3257 8566 3258 8570
rect 3270 8566 3271 8570
rect 3273 8566 3274 8570
rect 4099 8566 4100 8570
rect 4102 8566 4105 8570
rect 4107 8566 4108 8570
rect 4120 8566 4121 8570
rect 4123 8566 4124 8570
rect 4136 8566 4137 8570
rect 4139 8566 4142 8570
rect 4144 8566 4145 8570
rect 4162 8566 4163 8570
rect 4165 8566 4166 8570
rect 4178 8566 4179 8570
rect 4181 8566 4182 8570
rect 4194 8566 4195 8570
rect 4197 8566 4200 8570
rect 4202 8566 4203 8570
rect 4215 8566 4216 8570
rect 4218 8566 4219 8570
rect 2371 8536 2372 8540
rect 2374 8536 2377 8540
rect 2379 8536 2380 8540
rect 2392 8536 2393 8540
rect 2395 8536 2396 8540
rect 2408 8536 2409 8540
rect 2411 8536 2414 8540
rect 2416 8536 2417 8540
rect 2434 8536 2435 8540
rect 2437 8536 2438 8540
rect 2450 8536 2451 8540
rect 2453 8536 2454 8540
rect 2466 8536 2467 8540
rect 2469 8536 2472 8540
rect 2474 8536 2475 8540
rect 2487 8536 2488 8540
rect 2490 8536 2491 8540
rect 2503 8536 2504 8540
rect 2506 8536 2509 8540
rect 2511 8536 2512 8540
rect 2524 8536 2525 8540
rect 2527 8536 2528 8540
rect 2540 8536 2541 8540
rect 2543 8536 2546 8540
rect 2548 8536 2549 8540
rect 2566 8536 2567 8540
rect 2569 8536 2570 8540
rect 2582 8536 2583 8540
rect 2585 8536 2586 8540
rect 2598 8536 2599 8540
rect 2601 8536 2604 8540
rect 2606 8536 2607 8540
rect 2619 8536 2620 8540
rect 2622 8536 2623 8540
rect 2635 8536 2636 8540
rect 2638 8536 2641 8540
rect 2643 8536 2644 8540
rect 2656 8536 2657 8540
rect 2659 8536 2660 8540
rect 2672 8536 2673 8540
rect 2675 8536 2678 8540
rect 2680 8536 2681 8540
rect 2698 8536 2699 8540
rect 2701 8536 2702 8540
rect 2714 8536 2715 8540
rect 2717 8536 2718 8540
rect 2730 8536 2731 8540
rect 2733 8536 2736 8540
rect 2738 8536 2739 8540
rect 2751 8536 2752 8540
rect 2754 8536 2755 8540
rect 3316 8536 3317 8540
rect 3319 8536 3322 8540
rect 3324 8536 3325 8540
rect 3337 8536 3338 8540
rect 3340 8536 3341 8540
rect 3353 8536 3354 8540
rect 3356 8536 3359 8540
rect 3361 8536 3362 8540
rect 3379 8536 3380 8540
rect 3382 8536 3383 8540
rect 3395 8536 3396 8540
rect 3398 8536 3399 8540
rect 3411 8536 3412 8540
rect 3414 8536 3417 8540
rect 3419 8536 3420 8540
rect 3432 8536 3433 8540
rect 3435 8536 3436 8540
rect 3448 8536 3449 8540
rect 3451 8536 3454 8540
rect 3456 8536 3457 8540
rect 3469 8536 3470 8540
rect 3472 8536 3473 8540
rect 3485 8536 3486 8540
rect 3488 8536 3491 8540
rect 3493 8536 3494 8540
rect 3511 8536 3512 8540
rect 3514 8536 3515 8540
rect 3527 8536 3528 8540
rect 3530 8536 3531 8540
rect 3543 8536 3544 8540
rect 3546 8536 3549 8540
rect 3551 8536 3552 8540
rect 3564 8536 3565 8540
rect 3567 8536 3568 8540
rect 3580 8536 3581 8540
rect 3583 8536 3586 8540
rect 3588 8536 3589 8540
rect 3601 8536 3602 8540
rect 3604 8536 3605 8540
rect 3617 8536 3618 8540
rect 3620 8536 3623 8540
rect 3625 8536 3626 8540
rect 3643 8536 3644 8540
rect 3646 8536 3647 8540
rect 3659 8536 3660 8540
rect 3662 8536 3663 8540
rect 3675 8536 3676 8540
rect 3678 8536 3681 8540
rect 3683 8536 3684 8540
rect 3696 8536 3697 8540
rect 3699 8536 3700 8540
rect 2603 8492 2604 8496
rect 2606 8492 2607 8496
rect 2627 8492 2628 8496
rect 2630 8492 2631 8496
rect 3548 8492 3549 8496
rect 3551 8492 3552 8496
rect 3572 8492 3573 8496
rect 3575 8492 3576 8496
rect 2623 8481 2624 8485
rect 2626 8481 2627 8485
rect 3568 8481 3569 8485
rect 3571 8481 3572 8485
rect 2615 8469 2619 8470
rect 2615 8466 2619 8467
rect 3560 8469 3564 8470
rect 3560 8466 3564 8467
rect 2603 8458 2604 8462
rect 2606 8458 2607 8462
rect 2627 8458 2628 8462
rect 2630 8458 2631 8462
rect 3548 8458 3549 8462
rect 3551 8458 3552 8462
rect 3572 8458 3573 8462
rect 3575 8458 3576 8462
rect 2371 8396 2372 8400
rect 2374 8396 2377 8400
rect 2379 8396 2380 8400
rect 2392 8396 2393 8400
rect 2395 8396 2396 8400
rect 2408 8396 2409 8400
rect 2411 8396 2414 8400
rect 2416 8396 2417 8400
rect 2434 8396 2435 8400
rect 2437 8396 2438 8400
rect 2450 8396 2451 8400
rect 2453 8396 2454 8400
rect 2466 8396 2467 8400
rect 2469 8396 2472 8400
rect 2474 8396 2475 8400
rect 2487 8396 2488 8400
rect 2490 8396 2491 8400
rect 2503 8396 2504 8400
rect 2506 8396 2509 8400
rect 2511 8396 2512 8400
rect 2524 8396 2525 8400
rect 2527 8396 2528 8400
rect 2540 8396 2541 8400
rect 2543 8396 2546 8400
rect 2548 8396 2549 8400
rect 2566 8396 2567 8400
rect 2569 8396 2570 8400
rect 2582 8396 2583 8400
rect 2585 8396 2586 8400
rect 2598 8396 2599 8400
rect 2601 8396 2604 8400
rect 2606 8396 2607 8400
rect 2619 8396 2620 8400
rect 2622 8396 2623 8400
rect 2635 8396 2636 8400
rect 2638 8396 2641 8400
rect 2643 8396 2644 8400
rect 2656 8396 2657 8400
rect 2659 8396 2660 8400
rect 2672 8396 2673 8400
rect 2675 8396 2678 8400
rect 2680 8396 2681 8400
rect 2698 8396 2699 8400
rect 2701 8396 2702 8400
rect 2714 8396 2715 8400
rect 2717 8396 2718 8400
rect 2730 8396 2731 8400
rect 2733 8396 2736 8400
rect 2738 8396 2739 8400
rect 2751 8396 2752 8400
rect 2754 8396 2755 8400
rect 3316 8396 3317 8400
rect 3319 8396 3322 8400
rect 3324 8396 3325 8400
rect 3337 8396 3338 8400
rect 3340 8396 3341 8400
rect 3353 8396 3354 8400
rect 3356 8396 3359 8400
rect 3361 8396 3362 8400
rect 3379 8396 3380 8400
rect 3382 8396 3383 8400
rect 3395 8396 3396 8400
rect 3398 8396 3399 8400
rect 3411 8396 3412 8400
rect 3414 8396 3417 8400
rect 3419 8396 3420 8400
rect 3432 8396 3433 8400
rect 3435 8396 3436 8400
rect 3448 8396 3449 8400
rect 3451 8396 3454 8400
rect 3456 8396 3457 8400
rect 3469 8396 3470 8400
rect 3472 8396 3473 8400
rect 3485 8396 3486 8400
rect 3488 8396 3491 8400
rect 3493 8396 3494 8400
rect 3511 8396 3512 8400
rect 3514 8396 3515 8400
rect 3527 8396 3528 8400
rect 3530 8396 3531 8400
rect 3543 8396 3544 8400
rect 3546 8396 3549 8400
rect 3551 8396 3552 8400
rect 3564 8396 3565 8400
rect 3567 8396 3568 8400
rect 3580 8396 3581 8400
rect 3583 8396 3586 8400
rect 3588 8396 3589 8400
rect 3601 8396 3602 8400
rect 3604 8396 3605 8400
rect 3617 8396 3618 8400
rect 3620 8396 3623 8400
rect 3625 8396 3626 8400
rect 3643 8396 3644 8400
rect 3646 8396 3647 8400
rect 3659 8396 3660 8400
rect 3662 8396 3663 8400
rect 3675 8396 3676 8400
rect 3678 8396 3681 8400
rect 3683 8396 3684 8400
rect 3696 8396 3697 8400
rect 3699 8396 3700 8400
rect 2855 8317 2856 8321
rect 2858 8317 2861 8321
rect 2863 8317 2864 8321
rect 2876 8317 2877 8321
rect 2879 8317 2880 8321
rect 2892 8317 2893 8321
rect 2895 8317 2898 8321
rect 2900 8317 2901 8321
rect 2918 8317 2919 8321
rect 2921 8317 2922 8321
rect 2934 8317 2935 8321
rect 2937 8317 2938 8321
rect 2950 8317 2951 8321
rect 2953 8317 2956 8321
rect 2958 8317 2959 8321
rect 2971 8317 2972 8321
rect 2974 8317 2975 8321
rect 2987 8317 2988 8321
rect 2990 8317 2993 8321
rect 2995 8317 2996 8321
rect 3008 8317 3009 8321
rect 3011 8317 3012 8321
rect 3024 8317 3025 8321
rect 3027 8317 3030 8321
rect 3032 8317 3033 8321
rect 3050 8317 3051 8321
rect 3053 8317 3054 8321
rect 3066 8317 3067 8321
rect 3069 8317 3070 8321
rect 3082 8317 3083 8321
rect 3085 8317 3088 8321
rect 3090 8317 3091 8321
rect 3103 8317 3104 8321
rect 3106 8317 3107 8321
rect 3119 8317 3120 8321
rect 3122 8317 3125 8321
rect 3127 8317 3128 8321
rect 3140 8317 3141 8321
rect 3143 8317 3144 8321
rect 3156 8317 3157 8321
rect 3159 8317 3162 8321
rect 3164 8317 3165 8321
rect 3182 8317 3183 8321
rect 3185 8317 3186 8321
rect 3198 8317 3199 8321
rect 3201 8317 3202 8321
rect 3214 8317 3215 8321
rect 3217 8317 3220 8321
rect 3222 8317 3223 8321
rect 3235 8317 3236 8321
rect 3238 8317 3239 8321
rect 3251 8317 3252 8321
rect 3254 8317 3257 8321
rect 3259 8317 3260 8321
rect 3272 8317 3273 8321
rect 3275 8317 3276 8321
rect 3288 8317 3289 8321
rect 3291 8317 3294 8321
rect 3296 8317 3297 8321
rect 3314 8317 3315 8321
rect 3317 8317 3318 8321
rect 3330 8317 3331 8321
rect 3333 8317 3334 8321
rect 3346 8317 3347 8321
rect 3349 8317 3352 8321
rect 3354 8317 3355 8321
rect 3367 8317 3368 8321
rect 3370 8317 3371 8321
rect 3800 8317 3801 8321
rect 3803 8317 3806 8321
rect 3808 8317 3809 8321
rect 3821 8317 3822 8321
rect 3824 8317 3825 8321
rect 3837 8317 3838 8321
rect 3840 8317 3843 8321
rect 3845 8317 3846 8321
rect 3863 8317 3864 8321
rect 3866 8317 3867 8321
rect 3879 8317 3880 8321
rect 3882 8317 3883 8321
rect 3895 8317 3896 8321
rect 3898 8317 3901 8321
rect 3903 8317 3904 8321
rect 3916 8317 3917 8321
rect 3919 8317 3920 8321
rect 3932 8317 3933 8321
rect 3935 8317 3938 8321
rect 3940 8317 3941 8321
rect 3953 8317 3954 8321
rect 3956 8317 3957 8321
rect 3969 8317 3970 8321
rect 3972 8317 3975 8321
rect 3977 8317 3978 8321
rect 3995 8317 3996 8321
rect 3998 8317 3999 8321
rect 4011 8317 4012 8321
rect 4014 8317 4015 8321
rect 4027 8317 4028 8321
rect 4030 8317 4033 8321
rect 4035 8317 4036 8321
rect 4048 8317 4049 8321
rect 4051 8317 4052 8321
rect 4064 8317 4065 8321
rect 4067 8317 4070 8321
rect 4072 8317 4073 8321
rect 4085 8317 4086 8321
rect 4088 8317 4089 8321
rect 4101 8317 4102 8321
rect 4104 8317 4107 8321
rect 4109 8317 4110 8321
rect 4127 8317 4128 8321
rect 4130 8317 4131 8321
rect 4143 8317 4144 8321
rect 4146 8317 4147 8321
rect 4159 8317 4160 8321
rect 4162 8317 4165 8321
rect 4167 8317 4168 8321
rect 4180 8317 4181 8321
rect 4183 8317 4184 8321
rect 4196 8317 4197 8321
rect 4199 8317 4202 8321
rect 4204 8317 4205 8321
rect 4217 8317 4218 8321
rect 4220 8317 4221 8321
rect 4233 8317 4234 8321
rect 4236 8317 4239 8321
rect 4241 8317 4242 8321
rect 4259 8317 4260 8321
rect 4262 8317 4263 8321
rect 4275 8317 4276 8321
rect 4278 8317 4279 8321
rect 4291 8317 4292 8321
rect 4294 8317 4297 8321
rect 4299 8317 4300 8321
rect 4312 8317 4313 8321
rect 4315 8317 4316 8321
rect 2503 8284 2504 8288
rect 2506 8284 2509 8288
rect 2511 8284 2512 8288
rect 2524 8284 2525 8288
rect 2527 8284 2528 8288
rect 2540 8284 2541 8288
rect 2543 8284 2546 8288
rect 2548 8284 2549 8288
rect 2566 8284 2567 8288
rect 2569 8284 2570 8288
rect 2582 8284 2583 8288
rect 2585 8284 2586 8288
rect 2598 8284 2599 8288
rect 2601 8284 2604 8288
rect 2606 8284 2607 8288
rect 2619 8284 2620 8288
rect 2622 8284 2623 8288
rect 3448 8284 3449 8288
rect 3451 8284 3454 8288
rect 3456 8284 3457 8288
rect 3469 8284 3470 8288
rect 3472 8284 3473 8288
rect 3485 8284 3486 8288
rect 3488 8284 3491 8288
rect 3493 8284 3494 8288
rect 3511 8284 3512 8288
rect 3514 8284 3515 8288
rect 3527 8284 3528 8288
rect 3530 8284 3531 8288
rect 3543 8284 3544 8288
rect 3546 8284 3549 8288
rect 3551 8284 3552 8288
rect 3564 8284 3565 8288
rect 3567 8284 3568 8288
rect 2627 8247 2628 8251
rect 2630 8247 2631 8251
rect 3034 8251 3035 8255
rect 3037 8251 3038 8255
rect 3058 8247 3061 8251
rect 3063 8247 3066 8251
rect 3068 8247 3069 8251
rect 3115 8251 3116 8255
rect 3118 8251 3119 8255
rect 3139 8247 3142 8251
rect 3144 8247 3147 8251
rect 3149 8247 3150 8251
rect 3088 8243 3089 8247
rect 3091 8243 3092 8247
rect 2510 8238 2511 8242
rect 2513 8238 2514 8242
rect 2860 8238 2861 8242
rect 2863 8238 2864 8242
rect 2876 8238 2877 8242
rect 2879 8238 2880 8242
rect 2892 8238 2893 8242
rect 2895 8238 2896 8242
rect 2911 8238 2916 8242
rect 2918 8238 2921 8242
rect 2923 8238 2924 8242
rect 2945 8238 2947 8242
rect 2949 8238 2950 8242
rect 2967 8238 2968 8242
rect 2970 8238 2971 8242
rect 2983 8238 2988 8242
rect 2990 8238 2993 8242
rect 2995 8238 2996 8242
rect 3010 8238 3011 8242
rect 3013 8238 3014 8242
rect 3169 8243 3170 8247
rect 3172 8243 3173 8247
rect 3572 8247 3573 8251
rect 3575 8247 3576 8251
rect 3979 8251 3980 8255
rect 3982 8251 3983 8255
rect 4003 8247 4006 8251
rect 4008 8247 4011 8251
rect 4013 8247 4014 8251
rect 4060 8251 4061 8255
rect 4063 8251 4064 8255
rect 4084 8247 4087 8251
rect 4089 8247 4092 8251
rect 4094 8247 4095 8251
rect 4033 8243 4034 8247
rect 4036 8243 4037 8247
rect 3455 8238 3456 8242
rect 3458 8238 3459 8242
rect 3805 8238 3806 8242
rect 3808 8238 3809 8242
rect 3821 8238 3822 8242
rect 3824 8238 3825 8242
rect 3837 8238 3838 8242
rect 3840 8238 3841 8242
rect 3856 8238 3861 8242
rect 3863 8238 3866 8242
rect 3868 8238 3869 8242
rect 3890 8238 3892 8242
rect 3894 8238 3895 8242
rect 3912 8238 3913 8242
rect 3915 8238 3916 8242
rect 3928 8238 3933 8242
rect 3935 8238 3938 8242
rect 3940 8238 3941 8242
rect 3955 8238 3956 8242
rect 3958 8238 3959 8242
rect 4114 8243 4115 8247
rect 4117 8243 4118 8247
rect 2860 8192 2861 8196
rect 2863 8192 2864 8196
rect 2876 8192 2877 8196
rect 2879 8192 2880 8196
rect 2892 8192 2893 8196
rect 2895 8192 2896 8196
rect 2911 8192 2916 8196
rect 2918 8192 2921 8196
rect 2923 8192 2924 8196
rect 2945 8192 2947 8196
rect 2949 8192 2950 8196
rect 2967 8192 2968 8196
rect 2970 8192 2971 8196
rect 2983 8192 2988 8196
rect 2990 8192 2993 8196
rect 2995 8192 2996 8196
rect 3010 8192 3011 8196
rect 3013 8192 3014 8196
rect 2494 8182 2495 8186
rect 2497 8182 2498 8186
rect 2510 8182 2511 8186
rect 2513 8182 2516 8186
rect 2518 8182 2519 8186
rect 2531 8182 2532 8186
rect 2534 8182 2535 8186
rect 2547 8182 2548 8186
rect 2550 8182 2551 8186
rect 2568 8182 2569 8186
rect 2571 8182 2574 8186
rect 2576 8182 2577 8186
rect 2589 8182 2590 8186
rect 2592 8182 2593 8186
rect 2605 8182 2606 8186
rect 2608 8182 2611 8186
rect 2613 8182 2614 8186
rect 3058 8191 3061 8195
rect 3063 8191 3066 8195
rect 3068 8191 3069 8195
rect 3139 8191 3142 8195
rect 3144 8191 3147 8195
rect 3149 8191 3150 8195
rect 3805 8192 3806 8196
rect 3808 8192 3809 8196
rect 3821 8192 3822 8196
rect 3824 8192 3825 8196
rect 3837 8192 3838 8196
rect 3840 8192 3841 8196
rect 3856 8192 3861 8196
rect 3863 8192 3866 8196
rect 3868 8192 3869 8196
rect 3890 8192 3892 8196
rect 3894 8192 3895 8196
rect 3912 8192 3913 8196
rect 3915 8192 3916 8196
rect 3928 8192 3933 8196
rect 3935 8192 3938 8196
rect 3940 8192 3941 8196
rect 3955 8192 3956 8196
rect 3958 8192 3959 8196
rect 3439 8182 3440 8186
rect 3442 8182 3443 8186
rect 3455 8182 3456 8186
rect 3458 8182 3461 8186
rect 3463 8182 3464 8186
rect 3476 8182 3477 8186
rect 3479 8182 3480 8186
rect 3492 8182 3493 8186
rect 3495 8182 3496 8186
rect 3513 8182 3514 8186
rect 3516 8182 3519 8186
rect 3521 8182 3522 8186
rect 3534 8182 3535 8186
rect 3537 8182 3538 8186
rect 3550 8182 3551 8186
rect 3553 8182 3556 8186
rect 3558 8182 3559 8186
rect 4003 8191 4006 8195
rect 4008 8191 4011 8195
rect 4013 8191 4014 8195
rect 4084 8191 4087 8195
rect 4089 8191 4092 8195
rect 4094 8191 4095 8195
rect 3058 8115 3061 8119
rect 3063 8115 3066 8119
rect 3068 8115 3069 8119
rect 3139 8119 3140 8123
rect 3142 8119 3143 8123
rect 3163 8115 3166 8119
rect 3168 8115 3171 8119
rect 3173 8115 3174 8119
rect 3088 8111 3089 8115
rect 3091 8111 3092 8115
rect 2860 8106 2861 8110
rect 2863 8106 2864 8110
rect 2876 8106 2877 8110
rect 2879 8106 2880 8110
rect 2892 8106 2893 8110
rect 2895 8106 2896 8110
rect 2911 8106 2916 8110
rect 2918 8106 2921 8110
rect 2923 8106 2924 8110
rect 2945 8106 2947 8110
rect 2949 8106 2950 8110
rect 2967 8106 2968 8110
rect 2970 8106 2971 8110
rect 2983 8106 2988 8110
rect 2990 8106 2993 8110
rect 2995 8106 2996 8110
rect 3010 8106 3011 8110
rect 3013 8106 3014 8110
rect 3193 8111 3194 8115
rect 3196 8111 3197 8115
rect 4003 8115 4006 8119
rect 4008 8115 4011 8119
rect 4013 8115 4014 8119
rect 4084 8119 4085 8123
rect 4087 8119 4088 8123
rect 4108 8115 4111 8119
rect 4113 8115 4116 8119
rect 4118 8115 4119 8119
rect 4033 8111 4034 8115
rect 4036 8111 4037 8115
rect 3805 8106 3806 8110
rect 3808 8106 3809 8110
rect 3821 8106 3822 8110
rect 3824 8106 3825 8110
rect 3837 8106 3838 8110
rect 3840 8106 3841 8110
rect 3856 8106 3861 8110
rect 3863 8106 3866 8110
rect 3868 8106 3869 8110
rect 3890 8106 3892 8110
rect 3894 8106 3895 8110
rect 3912 8106 3913 8110
rect 3915 8106 3916 8110
rect 3928 8106 3933 8110
rect 3935 8106 3938 8110
rect 3940 8106 3941 8110
rect 3955 8106 3956 8110
rect 3958 8106 3959 8110
rect 4138 8111 4139 8115
rect 4141 8111 4142 8115
rect 2860 8060 2861 8064
rect 2863 8060 2864 8064
rect 2876 8060 2877 8064
rect 2879 8060 2880 8064
rect 2892 8060 2893 8064
rect 2895 8060 2896 8064
rect 2911 8060 2916 8064
rect 2918 8060 2921 8064
rect 2923 8060 2924 8064
rect 2945 8060 2947 8064
rect 2949 8060 2950 8064
rect 2967 8060 2968 8064
rect 2970 8060 2971 8064
rect 2983 8060 2988 8064
rect 2990 8060 2993 8064
rect 2995 8060 2996 8064
rect 3010 8060 3011 8064
rect 3013 8060 3014 8064
rect 3058 8060 3061 8064
rect 3063 8060 3066 8064
rect 3068 8060 3069 8064
rect 3163 8060 3166 8064
rect 3168 8060 3171 8064
rect 3173 8060 3174 8064
rect 3805 8060 3806 8064
rect 3808 8060 3809 8064
rect 3821 8060 3822 8064
rect 3824 8060 3825 8064
rect 3837 8060 3838 8064
rect 3840 8060 3841 8064
rect 3856 8060 3861 8064
rect 3863 8060 3866 8064
rect 3868 8060 3869 8064
rect 3890 8060 3892 8064
rect 3894 8060 3895 8064
rect 3912 8060 3913 8064
rect 3915 8060 3916 8064
rect 3928 8060 3933 8064
rect 3935 8060 3938 8064
rect 3940 8060 3941 8064
rect 3955 8060 3956 8064
rect 3958 8060 3959 8064
rect 4003 8060 4006 8064
rect 4008 8060 4011 8064
rect 4013 8060 4014 8064
rect 4108 8060 4111 8064
rect 4113 8060 4116 8064
rect 4118 8060 4119 8064
rect 3058 7983 3061 7987
rect 3063 7983 3066 7987
rect 3068 7983 3069 7987
rect 3115 7987 3116 7991
rect 3118 7987 3119 7991
rect 3139 7983 3142 7987
rect 3144 7983 3147 7987
rect 3149 7983 3150 7987
rect 3205 7987 3206 7991
rect 3208 7987 3209 7991
rect 3229 7983 3232 7987
rect 3234 7983 3237 7987
rect 3239 7983 3240 7987
rect 3088 7979 3089 7983
rect 3091 7979 3092 7983
rect 2860 7974 2861 7978
rect 2863 7974 2864 7978
rect 2876 7974 2877 7978
rect 2879 7974 2880 7978
rect 2892 7974 2893 7978
rect 2895 7974 2896 7978
rect 2911 7974 2916 7978
rect 2918 7974 2921 7978
rect 2923 7974 2924 7978
rect 2945 7974 2947 7978
rect 2949 7974 2950 7978
rect 2967 7974 2968 7978
rect 2970 7974 2971 7978
rect 2983 7974 2988 7978
rect 2990 7974 2993 7978
rect 2995 7974 2996 7978
rect 3010 7974 3011 7978
rect 3013 7974 3014 7978
rect 3169 7979 3170 7983
rect 3172 7979 3173 7983
rect 3259 7979 3260 7983
rect 3262 7979 3263 7983
rect 4003 7983 4006 7987
rect 4008 7983 4011 7987
rect 4013 7983 4014 7987
rect 4060 7987 4061 7991
rect 4063 7987 4064 7991
rect 4084 7983 4087 7987
rect 4089 7983 4092 7987
rect 4094 7983 4095 7987
rect 4150 7987 4151 7991
rect 4153 7987 4154 7991
rect 4174 7983 4177 7987
rect 4179 7983 4182 7987
rect 4184 7983 4185 7987
rect 4033 7979 4034 7983
rect 4036 7979 4037 7983
rect 3805 7974 3806 7978
rect 3808 7974 3809 7978
rect 3821 7974 3822 7978
rect 3824 7974 3825 7978
rect 3837 7974 3838 7978
rect 3840 7974 3841 7978
rect 3856 7974 3861 7978
rect 3863 7974 3866 7978
rect 3868 7974 3869 7978
rect 3890 7974 3892 7978
rect 3894 7974 3895 7978
rect 3912 7974 3913 7978
rect 3915 7974 3916 7978
rect 3928 7974 3933 7978
rect 3935 7974 3938 7978
rect 3940 7974 3941 7978
rect 3955 7974 3956 7978
rect 3958 7974 3959 7978
rect 4114 7979 4115 7983
rect 4117 7979 4118 7983
rect 4204 7979 4205 7983
rect 4207 7979 4208 7983
rect 2860 7928 2861 7932
rect 2863 7928 2864 7932
rect 2876 7928 2877 7932
rect 2879 7928 2880 7932
rect 2892 7928 2893 7932
rect 2895 7928 2896 7932
rect 2911 7928 2916 7932
rect 2918 7928 2921 7932
rect 2923 7928 2924 7932
rect 2945 7928 2947 7932
rect 2949 7928 2950 7932
rect 2967 7928 2968 7932
rect 2970 7928 2971 7932
rect 2983 7928 2988 7932
rect 2990 7928 2993 7932
rect 2995 7928 2996 7932
rect 3010 7928 3011 7932
rect 3013 7928 3014 7932
rect 3058 7925 3061 7929
rect 3063 7925 3066 7929
rect 3068 7925 3069 7929
rect 3139 7925 3142 7929
rect 3144 7925 3147 7929
rect 3149 7925 3150 7929
rect 3229 7925 3232 7929
rect 3234 7925 3237 7929
rect 3239 7925 3240 7929
rect 3805 7928 3806 7932
rect 3808 7928 3809 7932
rect 3821 7928 3822 7932
rect 3824 7928 3825 7932
rect 3837 7928 3838 7932
rect 3840 7928 3841 7932
rect 3856 7928 3861 7932
rect 3863 7928 3866 7932
rect 3868 7928 3869 7932
rect 3890 7928 3892 7932
rect 3894 7928 3895 7932
rect 3912 7928 3913 7932
rect 3915 7928 3916 7932
rect 3928 7928 3933 7932
rect 3935 7928 3938 7932
rect 3940 7928 3941 7932
rect 3955 7928 3956 7932
rect 3958 7928 3959 7932
rect 4003 7925 4006 7929
rect 4008 7925 4011 7929
rect 4013 7925 4014 7929
rect 4084 7925 4087 7929
rect 4089 7925 4092 7929
rect 4094 7925 4095 7929
rect 4174 7925 4177 7929
rect 4179 7925 4182 7929
rect 4184 7925 4185 7929
rect 3058 7851 3061 7855
rect 3063 7851 3066 7855
rect 3068 7851 3069 7855
rect 3088 7847 3089 7851
rect 3091 7847 3092 7851
rect 2860 7842 2861 7846
rect 2863 7842 2864 7846
rect 2876 7842 2877 7846
rect 2879 7842 2880 7846
rect 2892 7842 2893 7846
rect 2895 7842 2896 7846
rect 2911 7842 2916 7846
rect 2918 7842 2921 7846
rect 2923 7842 2924 7846
rect 2945 7842 2947 7846
rect 2949 7842 2950 7846
rect 2967 7842 2968 7846
rect 2970 7842 2971 7846
rect 2983 7842 2988 7846
rect 2990 7842 2993 7846
rect 2995 7842 2996 7846
rect 3010 7842 3011 7846
rect 3013 7842 3014 7846
rect 4003 7851 4006 7855
rect 4008 7851 4011 7855
rect 4013 7851 4014 7855
rect 4033 7847 4034 7851
rect 4036 7847 4037 7851
rect 3805 7842 3806 7846
rect 3808 7842 3809 7846
rect 3821 7842 3822 7846
rect 3824 7842 3825 7846
rect 3837 7842 3838 7846
rect 3840 7842 3841 7846
rect 3856 7842 3861 7846
rect 3863 7842 3866 7846
rect 3868 7842 3869 7846
rect 3890 7842 3892 7846
rect 3894 7842 3895 7846
rect 3912 7842 3913 7846
rect 3915 7842 3916 7846
rect 3928 7842 3933 7846
rect 3935 7842 3938 7846
rect 3940 7842 3941 7846
rect 3955 7842 3956 7846
rect 3958 7842 3959 7846
rect 2860 7796 2861 7800
rect 2863 7796 2864 7800
rect 2876 7796 2877 7800
rect 2879 7796 2880 7800
rect 2892 7796 2893 7800
rect 2895 7796 2896 7800
rect 2911 7796 2916 7800
rect 2918 7796 2921 7800
rect 2923 7796 2924 7800
rect 2945 7796 2947 7800
rect 2949 7796 2950 7800
rect 2967 7796 2968 7800
rect 2970 7796 2971 7800
rect 2983 7796 2988 7800
rect 2990 7796 2993 7800
rect 2995 7796 2996 7800
rect 3010 7796 3011 7800
rect 3013 7796 3014 7800
rect 3094 7796 3095 7800
rect 3097 7796 3098 7800
rect 3102 7796 3108 7800
rect 3112 7796 3113 7800
rect 3115 7796 3116 7800
rect 3137 7796 3138 7800
rect 3140 7796 3141 7800
rect 3153 7796 3154 7800
rect 3156 7796 3157 7800
rect 3172 7796 3177 7800
rect 3179 7796 3182 7800
rect 3184 7796 3185 7800
rect 3206 7796 3208 7800
rect 3210 7796 3211 7800
rect 3228 7796 3229 7800
rect 3231 7796 3232 7800
rect 3244 7796 3249 7800
rect 3251 7796 3254 7800
rect 3256 7796 3257 7800
rect 3271 7796 3272 7800
rect 3274 7796 3275 7800
rect 2371 7782 2372 7786
rect 2374 7782 2377 7786
rect 2379 7782 2380 7786
rect 2392 7782 2393 7786
rect 2395 7782 2396 7786
rect 2408 7782 2409 7786
rect 2411 7782 2414 7786
rect 2416 7782 2417 7786
rect 2434 7782 2435 7786
rect 2437 7782 2438 7786
rect 2450 7782 2451 7786
rect 2453 7782 2454 7786
rect 2466 7782 2467 7786
rect 2469 7782 2472 7786
rect 2474 7782 2475 7786
rect 2487 7782 2488 7786
rect 2490 7782 2491 7786
rect 2503 7782 2504 7786
rect 2506 7782 2509 7786
rect 2511 7782 2512 7786
rect 2524 7782 2525 7786
rect 2527 7782 2528 7786
rect 2540 7782 2541 7786
rect 2543 7782 2546 7786
rect 2548 7782 2549 7786
rect 2566 7782 2567 7786
rect 2569 7782 2570 7786
rect 2582 7782 2583 7786
rect 2585 7782 2586 7786
rect 2598 7782 2599 7786
rect 2601 7782 2604 7786
rect 2606 7782 2607 7786
rect 2619 7782 2620 7786
rect 2622 7782 2623 7786
rect 2635 7782 2636 7786
rect 2638 7782 2641 7786
rect 2643 7782 2644 7786
rect 2656 7782 2657 7786
rect 2659 7782 2660 7786
rect 2672 7782 2673 7786
rect 2675 7782 2678 7786
rect 2680 7782 2681 7786
rect 2698 7782 2699 7786
rect 2701 7782 2702 7786
rect 2714 7782 2715 7786
rect 2717 7782 2718 7786
rect 2730 7782 2731 7786
rect 2733 7782 2736 7786
rect 2738 7782 2739 7786
rect 2751 7782 2752 7786
rect 2754 7782 2755 7786
rect 3058 7789 3061 7793
rect 3063 7789 3066 7793
rect 3068 7789 3069 7793
rect 3805 7796 3806 7800
rect 3808 7796 3809 7800
rect 3821 7796 3822 7800
rect 3824 7796 3825 7800
rect 3837 7796 3838 7800
rect 3840 7796 3841 7800
rect 3856 7796 3861 7800
rect 3863 7796 3866 7800
rect 3868 7796 3869 7800
rect 3890 7796 3892 7800
rect 3894 7796 3895 7800
rect 3912 7796 3913 7800
rect 3915 7796 3916 7800
rect 3928 7796 3933 7800
rect 3935 7796 3938 7800
rect 3940 7796 3941 7800
rect 3955 7796 3956 7800
rect 3958 7796 3959 7800
rect 4039 7796 4040 7800
rect 4042 7796 4043 7800
rect 4047 7796 4053 7800
rect 4057 7796 4058 7800
rect 4060 7796 4061 7800
rect 4082 7796 4083 7800
rect 4085 7796 4086 7800
rect 4098 7796 4099 7800
rect 4101 7796 4102 7800
rect 4117 7796 4122 7800
rect 4124 7796 4127 7800
rect 4129 7796 4130 7800
rect 4151 7796 4153 7800
rect 4155 7796 4156 7800
rect 4173 7796 4174 7800
rect 4176 7796 4177 7800
rect 4189 7796 4194 7800
rect 4196 7796 4199 7800
rect 4201 7796 4202 7800
rect 4216 7796 4217 7800
rect 4219 7796 4220 7800
rect 3316 7782 3317 7786
rect 3319 7782 3322 7786
rect 3324 7782 3325 7786
rect 3337 7782 3338 7786
rect 3340 7782 3341 7786
rect 3353 7782 3354 7786
rect 3356 7782 3359 7786
rect 3361 7782 3362 7786
rect 3379 7782 3380 7786
rect 3382 7782 3383 7786
rect 3395 7782 3396 7786
rect 3398 7782 3399 7786
rect 3411 7782 3412 7786
rect 3414 7782 3417 7786
rect 3419 7782 3420 7786
rect 3432 7782 3433 7786
rect 3435 7782 3436 7786
rect 3448 7782 3449 7786
rect 3451 7782 3454 7786
rect 3456 7782 3457 7786
rect 3469 7782 3470 7786
rect 3472 7782 3473 7786
rect 3485 7782 3486 7786
rect 3488 7782 3491 7786
rect 3493 7782 3494 7786
rect 3511 7782 3512 7786
rect 3514 7782 3515 7786
rect 3527 7782 3528 7786
rect 3530 7782 3531 7786
rect 3543 7782 3544 7786
rect 3546 7782 3549 7786
rect 3551 7782 3552 7786
rect 3564 7782 3565 7786
rect 3567 7782 3568 7786
rect 3580 7782 3581 7786
rect 3583 7782 3586 7786
rect 3588 7782 3589 7786
rect 3601 7782 3602 7786
rect 3604 7782 3605 7786
rect 3617 7782 3618 7786
rect 3620 7782 3623 7786
rect 3625 7782 3626 7786
rect 3643 7782 3644 7786
rect 3646 7782 3647 7786
rect 3659 7782 3660 7786
rect 3662 7782 3663 7786
rect 3675 7782 3676 7786
rect 3678 7782 3681 7786
rect 3683 7782 3684 7786
rect 3696 7782 3697 7786
rect 3699 7782 3700 7786
rect 4003 7789 4006 7793
rect 4008 7789 4011 7793
rect 4013 7789 4014 7793
rect 2486 7738 2487 7742
rect 2489 7738 2490 7742
rect 2510 7738 2511 7742
rect 2513 7738 2514 7742
rect 3284 7742 3288 7743
rect 3284 7739 3288 7740
rect 3431 7738 3432 7742
rect 3434 7738 3435 7742
rect 3455 7738 3456 7742
rect 3458 7738 3459 7742
rect 4229 7742 4233 7743
rect 4229 7739 4233 7740
rect 2506 7725 2507 7729
rect 2509 7725 2510 7729
rect 3451 7725 3452 7729
rect 3454 7725 3455 7729
rect 2498 7713 2502 7714
rect 2498 7710 2502 7711
rect 3443 7713 3447 7714
rect 3443 7710 3447 7711
rect 2486 7702 2487 7706
rect 2489 7702 2490 7706
rect 2510 7702 2511 7706
rect 2513 7702 2514 7706
rect 3431 7702 3432 7706
rect 3434 7702 3435 7706
rect 3455 7702 3456 7706
rect 3458 7702 3459 7706
rect 3154 7670 3155 7674
rect 3157 7670 3160 7674
rect 3162 7670 3163 7674
rect 3175 7670 3176 7674
rect 3178 7670 3179 7674
rect 3191 7670 3192 7674
rect 3194 7670 3197 7674
rect 3199 7670 3200 7674
rect 3217 7670 3218 7674
rect 3220 7670 3221 7674
rect 3233 7670 3234 7674
rect 3236 7670 3237 7674
rect 3249 7670 3250 7674
rect 3252 7670 3255 7674
rect 3257 7670 3258 7674
rect 3270 7670 3271 7674
rect 3273 7670 3274 7674
rect 4099 7670 4100 7674
rect 4102 7670 4105 7674
rect 4107 7670 4108 7674
rect 4120 7670 4121 7674
rect 4123 7670 4124 7674
rect 4136 7670 4137 7674
rect 4139 7670 4142 7674
rect 4144 7670 4145 7674
rect 4162 7670 4163 7674
rect 4165 7670 4166 7674
rect 4178 7670 4179 7674
rect 4181 7670 4182 7674
rect 4194 7670 4195 7674
rect 4197 7670 4200 7674
rect 4202 7670 4203 7674
rect 4215 7670 4216 7674
rect 4218 7670 4219 7674
rect 2371 7640 2372 7644
rect 2374 7640 2377 7644
rect 2379 7640 2380 7644
rect 2392 7640 2393 7644
rect 2395 7640 2396 7644
rect 2408 7640 2409 7644
rect 2411 7640 2414 7644
rect 2416 7640 2417 7644
rect 2434 7640 2435 7644
rect 2437 7640 2438 7644
rect 2450 7640 2451 7644
rect 2453 7640 2454 7644
rect 2466 7640 2467 7644
rect 2469 7640 2472 7644
rect 2474 7640 2475 7644
rect 2487 7640 2488 7644
rect 2490 7640 2491 7644
rect 2503 7640 2504 7644
rect 2506 7640 2509 7644
rect 2511 7640 2512 7644
rect 2524 7640 2525 7644
rect 2527 7640 2528 7644
rect 2540 7640 2541 7644
rect 2543 7640 2546 7644
rect 2548 7640 2549 7644
rect 2566 7640 2567 7644
rect 2569 7640 2570 7644
rect 2582 7640 2583 7644
rect 2585 7640 2586 7644
rect 2598 7640 2599 7644
rect 2601 7640 2604 7644
rect 2606 7640 2607 7644
rect 2619 7640 2620 7644
rect 2622 7640 2623 7644
rect 2635 7640 2636 7644
rect 2638 7640 2641 7644
rect 2643 7640 2644 7644
rect 2656 7640 2657 7644
rect 2659 7640 2660 7644
rect 2672 7640 2673 7644
rect 2675 7640 2678 7644
rect 2680 7640 2681 7644
rect 2698 7640 2699 7644
rect 2701 7640 2702 7644
rect 2714 7640 2715 7644
rect 2717 7640 2718 7644
rect 2730 7640 2731 7644
rect 2733 7640 2736 7644
rect 2738 7640 2739 7644
rect 2751 7640 2752 7644
rect 2754 7640 2755 7644
rect 3316 7640 3317 7644
rect 3319 7640 3322 7644
rect 3324 7640 3325 7644
rect 3337 7640 3338 7644
rect 3340 7640 3341 7644
rect 3353 7640 3354 7644
rect 3356 7640 3359 7644
rect 3361 7640 3362 7644
rect 3379 7640 3380 7644
rect 3382 7640 3383 7644
rect 3395 7640 3396 7644
rect 3398 7640 3399 7644
rect 3411 7640 3412 7644
rect 3414 7640 3417 7644
rect 3419 7640 3420 7644
rect 3432 7640 3433 7644
rect 3435 7640 3436 7644
rect 3448 7640 3449 7644
rect 3451 7640 3454 7644
rect 3456 7640 3457 7644
rect 3469 7640 3470 7644
rect 3472 7640 3473 7644
rect 3485 7640 3486 7644
rect 3488 7640 3491 7644
rect 3493 7640 3494 7644
rect 3511 7640 3512 7644
rect 3514 7640 3515 7644
rect 3527 7640 3528 7644
rect 3530 7640 3531 7644
rect 3543 7640 3544 7644
rect 3546 7640 3549 7644
rect 3551 7640 3552 7644
rect 3564 7640 3565 7644
rect 3567 7640 3568 7644
rect 3580 7640 3581 7644
rect 3583 7640 3586 7644
rect 3588 7640 3589 7644
rect 3601 7640 3602 7644
rect 3604 7640 3605 7644
rect 3617 7640 3618 7644
rect 3620 7640 3623 7644
rect 3625 7640 3626 7644
rect 3643 7640 3644 7644
rect 3646 7640 3647 7644
rect 3659 7640 3660 7644
rect 3662 7640 3663 7644
rect 3675 7640 3676 7644
rect 3678 7640 3681 7644
rect 3683 7640 3684 7644
rect 3696 7640 3697 7644
rect 3699 7640 3700 7644
rect 3296 7596 3300 7597
rect 3296 7593 3300 7594
rect 4241 7596 4245 7597
rect 4241 7593 4245 7594
rect 3154 7584 3155 7588
rect 3157 7584 3160 7588
rect 3162 7584 3163 7588
rect 3175 7584 3176 7588
rect 3178 7584 3179 7588
rect 3191 7584 3192 7588
rect 3194 7584 3197 7588
rect 3199 7584 3200 7588
rect 3217 7584 3218 7588
rect 3220 7584 3221 7588
rect 3233 7584 3234 7588
rect 3236 7584 3237 7588
rect 3249 7584 3250 7588
rect 3252 7584 3255 7588
rect 3257 7584 3258 7588
rect 3270 7584 3271 7588
rect 3273 7584 3274 7588
rect 4099 7584 4100 7588
rect 4102 7584 4105 7588
rect 4107 7584 4108 7588
rect 4120 7584 4121 7588
rect 4123 7584 4124 7588
rect 4136 7584 4137 7588
rect 4139 7584 4142 7588
rect 4144 7584 4145 7588
rect 4162 7584 4163 7588
rect 4165 7584 4166 7588
rect 4178 7584 4179 7588
rect 4181 7584 4182 7588
rect 4194 7584 4195 7588
rect 4197 7584 4200 7588
rect 4202 7584 4203 7588
rect 4215 7584 4216 7588
rect 4218 7584 4219 7588
rect 2371 7554 2372 7558
rect 2374 7554 2377 7558
rect 2379 7554 2380 7558
rect 2392 7554 2393 7558
rect 2395 7554 2396 7558
rect 2408 7554 2409 7558
rect 2411 7554 2414 7558
rect 2416 7554 2417 7558
rect 2434 7554 2435 7558
rect 2437 7554 2438 7558
rect 2450 7554 2451 7558
rect 2453 7554 2454 7558
rect 2466 7554 2467 7558
rect 2469 7554 2472 7558
rect 2474 7554 2475 7558
rect 2487 7554 2488 7558
rect 2490 7554 2491 7558
rect 2503 7554 2504 7558
rect 2506 7554 2509 7558
rect 2511 7554 2512 7558
rect 2524 7554 2525 7558
rect 2527 7554 2528 7558
rect 2540 7554 2541 7558
rect 2543 7554 2546 7558
rect 2548 7554 2549 7558
rect 2566 7554 2567 7558
rect 2569 7554 2570 7558
rect 2582 7554 2583 7558
rect 2585 7554 2586 7558
rect 2598 7554 2599 7558
rect 2601 7554 2604 7558
rect 2606 7554 2607 7558
rect 2619 7554 2620 7558
rect 2622 7554 2623 7558
rect 2635 7554 2636 7558
rect 2638 7554 2641 7558
rect 2643 7554 2644 7558
rect 2656 7554 2657 7558
rect 2659 7554 2660 7558
rect 2672 7554 2673 7558
rect 2675 7554 2678 7558
rect 2680 7554 2681 7558
rect 2698 7554 2699 7558
rect 2701 7554 2702 7558
rect 2714 7554 2715 7558
rect 2717 7554 2718 7558
rect 2730 7554 2731 7558
rect 2733 7554 2736 7558
rect 2738 7554 2739 7558
rect 2751 7554 2752 7558
rect 2754 7554 2755 7558
rect 3316 7554 3317 7558
rect 3319 7554 3322 7558
rect 3324 7554 3325 7558
rect 3337 7554 3338 7558
rect 3340 7554 3341 7558
rect 3353 7554 3354 7558
rect 3356 7554 3359 7558
rect 3361 7554 3362 7558
rect 3379 7554 3380 7558
rect 3382 7554 3383 7558
rect 3395 7554 3396 7558
rect 3398 7554 3399 7558
rect 3411 7554 3412 7558
rect 3414 7554 3417 7558
rect 3419 7554 3420 7558
rect 3432 7554 3433 7558
rect 3435 7554 3436 7558
rect 3448 7554 3449 7558
rect 3451 7554 3454 7558
rect 3456 7554 3457 7558
rect 3469 7554 3470 7558
rect 3472 7554 3473 7558
rect 3485 7554 3486 7558
rect 3488 7554 3491 7558
rect 3493 7554 3494 7558
rect 3511 7554 3512 7558
rect 3514 7554 3515 7558
rect 3527 7554 3528 7558
rect 3530 7554 3531 7558
rect 3543 7554 3544 7558
rect 3546 7554 3549 7558
rect 3551 7554 3552 7558
rect 3564 7554 3565 7558
rect 3567 7554 3568 7558
rect 3580 7554 3581 7558
rect 3583 7554 3586 7558
rect 3588 7554 3589 7558
rect 3601 7554 3602 7558
rect 3604 7554 3605 7558
rect 3617 7554 3618 7558
rect 3620 7554 3623 7558
rect 3625 7554 3626 7558
rect 3643 7554 3644 7558
rect 3646 7554 3647 7558
rect 3659 7554 3660 7558
rect 3662 7554 3663 7558
rect 3675 7554 3676 7558
rect 3678 7554 3681 7558
rect 3683 7554 3684 7558
rect 3696 7554 3697 7558
rect 3699 7554 3700 7558
rect 2603 7510 2604 7514
rect 2606 7510 2607 7514
rect 2627 7510 2628 7514
rect 2630 7510 2631 7514
rect 3548 7510 3549 7514
rect 3551 7510 3552 7514
rect 3572 7510 3573 7514
rect 3575 7510 3576 7514
rect 2623 7499 2624 7503
rect 2626 7499 2627 7503
rect 3568 7499 3569 7503
rect 3571 7499 3572 7503
rect 2615 7487 2619 7488
rect 2615 7484 2619 7485
rect 3560 7487 3564 7488
rect 3560 7484 3564 7485
rect 2603 7476 2604 7480
rect 2606 7476 2607 7480
rect 2627 7476 2628 7480
rect 2630 7476 2631 7480
rect 3548 7476 3549 7480
rect 3551 7476 3552 7480
rect 3572 7476 3573 7480
rect 3575 7476 3576 7480
rect 3836 7475 3844 7476
rect 3836 7472 3844 7473
rect 2371 7414 2372 7418
rect 2374 7414 2377 7418
rect 2379 7414 2380 7418
rect 2392 7414 2393 7418
rect 2395 7414 2396 7418
rect 2408 7414 2409 7418
rect 2411 7414 2414 7418
rect 2416 7414 2417 7418
rect 2434 7414 2435 7418
rect 2437 7414 2438 7418
rect 2450 7414 2451 7418
rect 2453 7414 2454 7418
rect 2466 7414 2467 7418
rect 2469 7414 2472 7418
rect 2474 7414 2475 7418
rect 2487 7414 2488 7418
rect 2490 7414 2491 7418
rect 2503 7414 2504 7418
rect 2506 7414 2509 7418
rect 2511 7414 2512 7418
rect 2524 7414 2525 7418
rect 2527 7414 2528 7418
rect 2540 7414 2541 7418
rect 2543 7414 2546 7418
rect 2548 7414 2549 7418
rect 2566 7414 2567 7418
rect 2569 7414 2570 7418
rect 2582 7414 2583 7418
rect 2585 7414 2586 7418
rect 2598 7414 2599 7418
rect 2601 7414 2604 7418
rect 2606 7414 2607 7418
rect 2619 7414 2620 7418
rect 2622 7414 2623 7418
rect 2635 7414 2636 7418
rect 2638 7414 2641 7418
rect 2643 7414 2644 7418
rect 2656 7414 2657 7418
rect 2659 7414 2660 7418
rect 2672 7414 2673 7418
rect 2675 7414 2678 7418
rect 2680 7414 2681 7418
rect 2698 7414 2699 7418
rect 2701 7414 2702 7418
rect 2714 7414 2715 7418
rect 2717 7414 2718 7418
rect 2730 7414 2731 7418
rect 2733 7414 2736 7418
rect 2738 7414 2739 7418
rect 2751 7414 2752 7418
rect 2754 7414 2755 7418
rect 3316 7414 3317 7418
rect 3319 7414 3322 7418
rect 3324 7414 3325 7418
rect 3337 7414 3338 7418
rect 3340 7414 3341 7418
rect 3353 7414 3354 7418
rect 3356 7414 3359 7418
rect 3361 7414 3362 7418
rect 3379 7414 3380 7418
rect 3382 7414 3383 7418
rect 3395 7414 3396 7418
rect 3398 7414 3399 7418
rect 3411 7414 3412 7418
rect 3414 7414 3417 7418
rect 3419 7414 3420 7418
rect 3432 7414 3433 7418
rect 3435 7414 3436 7418
rect 3448 7414 3449 7418
rect 3451 7414 3454 7418
rect 3456 7414 3457 7418
rect 3469 7414 3470 7418
rect 3472 7414 3473 7418
rect 3485 7414 3486 7418
rect 3488 7414 3491 7418
rect 3493 7414 3494 7418
rect 3511 7414 3512 7418
rect 3514 7414 3515 7418
rect 3527 7414 3528 7418
rect 3530 7414 3531 7418
rect 3543 7414 3544 7418
rect 3546 7414 3549 7418
rect 3551 7414 3552 7418
rect 3564 7414 3565 7418
rect 3567 7414 3568 7418
rect 3580 7414 3581 7418
rect 3583 7414 3586 7418
rect 3588 7414 3589 7418
rect 3601 7414 3602 7418
rect 3604 7414 3605 7418
rect 3617 7414 3618 7418
rect 3620 7414 3623 7418
rect 3625 7414 3626 7418
rect 3643 7414 3644 7418
rect 3646 7414 3647 7418
rect 3659 7414 3660 7418
rect 3662 7414 3663 7418
rect 3675 7414 3676 7418
rect 3678 7414 3681 7418
rect 3683 7414 3684 7418
rect 3696 7414 3697 7418
rect 3699 7414 3700 7418
rect 1472 6896 1473 6900
rect 1475 6896 1476 6900
rect 1488 6896 1489 6900
rect 1491 6896 1494 6900
rect 1496 6896 1497 6900
rect 1509 6896 1510 6900
rect 1512 6896 1513 6900
rect 1525 6896 1526 6900
rect 1528 6896 1529 6900
rect 1546 6896 1547 6900
rect 1549 6896 1552 6900
rect 1554 6896 1555 6900
rect 1567 6896 1568 6900
rect 1570 6896 1571 6900
rect 1583 6896 1584 6900
rect 1586 6896 1589 6900
rect 1591 6896 1592 6900
rect 1604 6896 1605 6900
rect 1607 6896 1608 6900
rect 1620 6896 1621 6900
rect 1623 6896 1626 6900
rect 1628 6896 1629 6900
rect 1641 6896 1642 6900
rect 1644 6896 1645 6900
rect 1657 6896 1658 6900
rect 1660 6896 1661 6900
rect 1678 6896 1679 6900
rect 1681 6896 1684 6900
rect 1686 6896 1687 6900
rect 1699 6896 1700 6900
rect 1702 6896 1703 6900
rect 1715 6896 1716 6900
rect 1718 6896 1721 6900
rect 1723 6896 1724 6900
rect 1736 6896 1737 6900
rect 1739 6896 1740 6900
rect 1752 6896 1753 6900
rect 1755 6896 1758 6900
rect 1760 6896 1761 6900
rect 1773 6896 1774 6900
rect 1776 6896 1777 6900
rect 1789 6896 1790 6900
rect 1792 6896 1793 6900
rect 1810 6896 1811 6900
rect 1813 6896 1816 6900
rect 1818 6896 1819 6900
rect 1831 6896 1832 6900
rect 1834 6896 1835 6900
rect 1847 6896 1848 6900
rect 1850 6896 1853 6900
rect 1855 6896 1856 6900
rect 2417 6896 2418 6900
rect 2420 6896 2421 6900
rect 2433 6896 2434 6900
rect 2436 6896 2439 6900
rect 2441 6896 2442 6900
rect 2454 6896 2455 6900
rect 2457 6896 2458 6900
rect 2470 6896 2471 6900
rect 2473 6896 2474 6900
rect 2491 6896 2492 6900
rect 2494 6896 2497 6900
rect 2499 6896 2500 6900
rect 2512 6896 2513 6900
rect 2515 6896 2516 6900
rect 2528 6896 2529 6900
rect 2531 6896 2534 6900
rect 2536 6896 2537 6900
rect 2549 6896 2550 6900
rect 2552 6896 2553 6900
rect 2565 6896 2566 6900
rect 2568 6896 2571 6900
rect 2573 6896 2574 6900
rect 2586 6896 2587 6900
rect 2589 6896 2590 6900
rect 2602 6896 2603 6900
rect 2605 6896 2606 6900
rect 2623 6896 2624 6900
rect 2626 6896 2629 6900
rect 2631 6896 2632 6900
rect 2644 6896 2645 6900
rect 2647 6896 2648 6900
rect 2660 6896 2661 6900
rect 2663 6896 2666 6900
rect 2668 6896 2669 6900
rect 2681 6896 2682 6900
rect 2684 6896 2685 6900
rect 2697 6896 2698 6900
rect 2700 6896 2703 6900
rect 2705 6896 2706 6900
rect 2718 6896 2719 6900
rect 2721 6896 2722 6900
rect 2734 6896 2735 6900
rect 2737 6896 2738 6900
rect 2755 6896 2756 6900
rect 2758 6896 2761 6900
rect 2763 6896 2764 6900
rect 2776 6896 2777 6900
rect 2779 6896 2780 6900
rect 2792 6896 2793 6900
rect 2795 6896 2798 6900
rect 2800 6896 2801 6900
rect 1596 6834 1597 6838
rect 1599 6834 1600 6838
rect 1620 6834 1621 6838
rect 1623 6834 1624 6838
rect 2541 6834 2542 6838
rect 2544 6834 2545 6838
rect 2565 6834 2566 6838
rect 2568 6834 2569 6838
rect 1608 6829 1612 6830
rect 1608 6826 1612 6827
rect 2553 6829 2557 6830
rect 2553 6826 2557 6827
rect 1600 6811 1601 6815
rect 1603 6811 1604 6815
rect 2545 6811 2546 6815
rect 2548 6811 2549 6815
rect 1596 6800 1597 6804
rect 1599 6800 1600 6804
rect 1620 6800 1621 6804
rect 1623 6800 1624 6804
rect 2541 6800 2542 6804
rect 2544 6800 2545 6804
rect 2565 6800 2566 6804
rect 2568 6800 2569 6804
rect 1472 6756 1473 6760
rect 1475 6756 1476 6760
rect 1488 6756 1489 6760
rect 1491 6756 1494 6760
rect 1496 6756 1497 6760
rect 1509 6756 1510 6760
rect 1512 6756 1513 6760
rect 1525 6756 1526 6760
rect 1528 6756 1529 6760
rect 1546 6756 1547 6760
rect 1549 6756 1552 6760
rect 1554 6756 1555 6760
rect 1567 6756 1568 6760
rect 1570 6756 1571 6760
rect 1583 6756 1584 6760
rect 1586 6756 1589 6760
rect 1591 6756 1592 6760
rect 1604 6756 1605 6760
rect 1607 6756 1608 6760
rect 1620 6756 1621 6760
rect 1623 6756 1626 6760
rect 1628 6756 1629 6760
rect 1641 6756 1642 6760
rect 1644 6756 1645 6760
rect 1657 6756 1658 6760
rect 1660 6756 1661 6760
rect 1678 6756 1679 6760
rect 1681 6756 1684 6760
rect 1686 6756 1687 6760
rect 1699 6756 1700 6760
rect 1702 6756 1703 6760
rect 1715 6756 1716 6760
rect 1718 6756 1721 6760
rect 1723 6756 1724 6760
rect 1736 6756 1737 6760
rect 1739 6756 1740 6760
rect 1752 6756 1753 6760
rect 1755 6756 1758 6760
rect 1760 6756 1761 6760
rect 1773 6756 1774 6760
rect 1776 6756 1777 6760
rect 1789 6756 1790 6760
rect 1792 6756 1793 6760
rect 1810 6756 1811 6760
rect 1813 6756 1816 6760
rect 1818 6756 1819 6760
rect 1831 6756 1832 6760
rect 1834 6756 1835 6760
rect 1847 6756 1848 6760
rect 1850 6756 1853 6760
rect 1855 6756 1856 6760
rect 2417 6756 2418 6760
rect 2420 6756 2421 6760
rect 2433 6756 2434 6760
rect 2436 6756 2439 6760
rect 2441 6756 2442 6760
rect 2454 6756 2455 6760
rect 2457 6756 2458 6760
rect 2470 6756 2471 6760
rect 2473 6756 2474 6760
rect 2491 6756 2492 6760
rect 2494 6756 2497 6760
rect 2499 6756 2500 6760
rect 2512 6756 2513 6760
rect 2515 6756 2516 6760
rect 2528 6756 2529 6760
rect 2531 6756 2534 6760
rect 2536 6756 2537 6760
rect 2549 6756 2550 6760
rect 2552 6756 2553 6760
rect 2565 6756 2566 6760
rect 2568 6756 2571 6760
rect 2573 6756 2574 6760
rect 2586 6756 2587 6760
rect 2589 6756 2590 6760
rect 2602 6756 2603 6760
rect 2605 6756 2606 6760
rect 2623 6756 2624 6760
rect 2626 6756 2629 6760
rect 2631 6756 2632 6760
rect 2644 6756 2645 6760
rect 2647 6756 2648 6760
rect 2660 6756 2661 6760
rect 2663 6756 2666 6760
rect 2668 6756 2669 6760
rect 2681 6756 2682 6760
rect 2684 6756 2685 6760
rect 2697 6756 2698 6760
rect 2700 6756 2703 6760
rect 2705 6756 2706 6760
rect 2718 6756 2719 6760
rect 2721 6756 2722 6760
rect 2734 6756 2735 6760
rect 2737 6756 2738 6760
rect 2755 6756 2756 6760
rect 2758 6756 2761 6760
rect 2763 6756 2764 6760
rect 2776 6756 2777 6760
rect 2779 6756 2780 6760
rect 2792 6756 2793 6760
rect 2795 6756 2798 6760
rect 2800 6756 2801 6760
rect 953 6726 954 6730
rect 956 6726 957 6730
rect 969 6726 970 6730
rect 972 6726 975 6730
rect 977 6726 978 6730
rect 990 6726 991 6730
rect 993 6726 994 6730
rect 1006 6726 1007 6730
rect 1009 6726 1010 6730
rect 1027 6726 1028 6730
rect 1030 6726 1033 6730
rect 1035 6726 1036 6730
rect 1048 6726 1049 6730
rect 1051 6726 1052 6730
rect 1064 6726 1065 6730
rect 1067 6726 1070 6730
rect 1072 6726 1073 6730
rect 1898 6726 1899 6730
rect 1901 6726 1902 6730
rect 1914 6726 1915 6730
rect 1917 6726 1920 6730
rect 1922 6726 1923 6730
rect 1935 6726 1936 6730
rect 1938 6726 1939 6730
rect 1951 6726 1952 6730
rect 1954 6726 1955 6730
rect 1972 6726 1973 6730
rect 1975 6726 1978 6730
rect 1980 6726 1981 6730
rect 1993 6726 1994 6730
rect 1996 6726 1997 6730
rect 2009 6726 2010 6730
rect 2012 6726 2015 6730
rect 2017 6726 2018 6730
rect 927 6720 931 6721
rect 927 6717 931 6718
rect 1872 6720 1876 6721
rect 1872 6717 1876 6718
rect 1472 6670 1473 6674
rect 1475 6670 1476 6674
rect 1488 6670 1489 6674
rect 1491 6670 1494 6674
rect 1496 6670 1497 6674
rect 1509 6670 1510 6674
rect 1512 6670 1513 6674
rect 1525 6670 1526 6674
rect 1528 6670 1529 6674
rect 1546 6670 1547 6674
rect 1549 6670 1552 6674
rect 1554 6670 1555 6674
rect 1567 6670 1568 6674
rect 1570 6670 1571 6674
rect 1583 6670 1584 6674
rect 1586 6670 1589 6674
rect 1591 6670 1592 6674
rect 1604 6670 1605 6674
rect 1607 6670 1608 6674
rect 1620 6670 1621 6674
rect 1623 6670 1626 6674
rect 1628 6670 1629 6674
rect 1641 6670 1642 6674
rect 1644 6670 1645 6674
rect 1657 6670 1658 6674
rect 1660 6670 1661 6674
rect 1678 6670 1679 6674
rect 1681 6670 1684 6674
rect 1686 6670 1687 6674
rect 1699 6670 1700 6674
rect 1702 6670 1703 6674
rect 1715 6670 1716 6674
rect 1718 6670 1721 6674
rect 1723 6670 1724 6674
rect 1736 6670 1737 6674
rect 1739 6670 1740 6674
rect 1752 6670 1753 6674
rect 1755 6670 1758 6674
rect 1760 6670 1761 6674
rect 1773 6670 1774 6674
rect 1776 6670 1777 6674
rect 1789 6670 1790 6674
rect 1792 6670 1793 6674
rect 1810 6670 1811 6674
rect 1813 6670 1816 6674
rect 1818 6670 1819 6674
rect 1831 6670 1832 6674
rect 1834 6670 1835 6674
rect 1847 6670 1848 6674
rect 1850 6670 1853 6674
rect 1855 6670 1856 6674
rect 2417 6670 2418 6674
rect 2420 6670 2421 6674
rect 2433 6670 2434 6674
rect 2436 6670 2439 6674
rect 2441 6670 2442 6674
rect 2454 6670 2455 6674
rect 2457 6670 2458 6674
rect 2470 6670 2471 6674
rect 2473 6670 2474 6674
rect 2491 6670 2492 6674
rect 2494 6670 2497 6674
rect 2499 6670 2500 6674
rect 2512 6670 2513 6674
rect 2515 6670 2516 6674
rect 2528 6670 2529 6674
rect 2531 6670 2534 6674
rect 2536 6670 2537 6674
rect 2549 6670 2550 6674
rect 2552 6670 2553 6674
rect 2565 6670 2566 6674
rect 2568 6670 2571 6674
rect 2573 6670 2574 6674
rect 2586 6670 2587 6674
rect 2589 6670 2590 6674
rect 2602 6670 2603 6674
rect 2605 6670 2606 6674
rect 2623 6670 2624 6674
rect 2626 6670 2629 6674
rect 2631 6670 2632 6674
rect 2644 6670 2645 6674
rect 2647 6670 2648 6674
rect 2660 6670 2661 6674
rect 2663 6670 2666 6674
rect 2668 6670 2669 6674
rect 2681 6670 2682 6674
rect 2684 6670 2685 6674
rect 2697 6670 2698 6674
rect 2700 6670 2703 6674
rect 2705 6670 2706 6674
rect 2718 6670 2719 6674
rect 2721 6670 2722 6674
rect 2734 6670 2735 6674
rect 2737 6670 2738 6674
rect 2755 6670 2756 6674
rect 2758 6670 2761 6674
rect 2763 6670 2764 6674
rect 2776 6670 2777 6674
rect 2779 6670 2780 6674
rect 2792 6670 2793 6674
rect 2795 6670 2798 6674
rect 2800 6670 2801 6674
rect 953 6640 954 6644
rect 956 6640 957 6644
rect 969 6640 970 6644
rect 972 6640 975 6644
rect 977 6640 978 6644
rect 990 6640 991 6644
rect 993 6640 994 6644
rect 1006 6640 1007 6644
rect 1009 6640 1010 6644
rect 1027 6640 1028 6644
rect 1030 6640 1033 6644
rect 1035 6640 1036 6644
rect 1048 6640 1049 6644
rect 1051 6640 1052 6644
rect 1064 6640 1065 6644
rect 1067 6640 1070 6644
rect 1072 6640 1073 6644
rect 1898 6640 1899 6644
rect 1901 6640 1902 6644
rect 1914 6640 1915 6644
rect 1917 6640 1920 6644
rect 1922 6640 1923 6644
rect 1935 6640 1936 6644
rect 1938 6640 1939 6644
rect 1951 6640 1952 6644
rect 1954 6640 1955 6644
rect 1972 6640 1973 6644
rect 1975 6640 1978 6644
rect 1980 6640 1981 6644
rect 1993 6640 1994 6644
rect 1996 6640 1997 6644
rect 2009 6640 2010 6644
rect 2012 6640 2015 6644
rect 2017 6640 2018 6644
rect 1713 6608 1714 6612
rect 1716 6608 1717 6612
rect 1737 6608 1738 6612
rect 1740 6608 1741 6612
rect 2658 6608 2659 6612
rect 2661 6608 2662 6612
rect 2682 6608 2683 6612
rect 2685 6608 2686 6612
rect 1725 6603 1729 6604
rect 1725 6600 1729 6601
rect 2670 6603 2674 6604
rect 2670 6600 2674 6601
rect 1717 6585 1718 6589
rect 1720 6585 1721 6589
rect 2662 6585 2663 6589
rect 2665 6585 2666 6589
rect 939 6574 943 6575
rect 939 6571 943 6572
rect 1713 6572 1714 6576
rect 1716 6572 1717 6576
rect 1737 6572 1738 6576
rect 1740 6572 1741 6576
rect 1884 6574 1888 6575
rect 1884 6571 1888 6572
rect 2658 6572 2659 6576
rect 2661 6572 2662 6576
rect 2682 6572 2683 6576
rect 2685 6572 2686 6576
rect 1158 6521 1159 6525
rect 1161 6521 1164 6525
rect 1166 6521 1169 6525
rect 1472 6528 1473 6532
rect 1475 6528 1476 6532
rect 1488 6528 1489 6532
rect 1491 6528 1494 6532
rect 1496 6528 1497 6532
rect 1509 6528 1510 6532
rect 1512 6528 1513 6532
rect 1525 6528 1526 6532
rect 1528 6528 1529 6532
rect 1546 6528 1547 6532
rect 1549 6528 1552 6532
rect 1554 6528 1555 6532
rect 1567 6528 1568 6532
rect 1570 6528 1571 6532
rect 1583 6528 1584 6532
rect 1586 6528 1589 6532
rect 1591 6528 1592 6532
rect 1604 6528 1605 6532
rect 1607 6528 1608 6532
rect 1620 6528 1621 6532
rect 1623 6528 1626 6532
rect 1628 6528 1629 6532
rect 1641 6528 1642 6532
rect 1644 6528 1645 6532
rect 1657 6528 1658 6532
rect 1660 6528 1661 6532
rect 1678 6528 1679 6532
rect 1681 6528 1684 6532
rect 1686 6528 1687 6532
rect 1699 6528 1700 6532
rect 1702 6528 1703 6532
rect 1715 6528 1716 6532
rect 1718 6528 1721 6532
rect 1723 6528 1724 6532
rect 1736 6528 1737 6532
rect 1739 6528 1740 6532
rect 1752 6528 1753 6532
rect 1755 6528 1758 6532
rect 1760 6528 1761 6532
rect 1773 6528 1774 6532
rect 1776 6528 1777 6532
rect 1789 6528 1790 6532
rect 1792 6528 1793 6532
rect 1810 6528 1811 6532
rect 1813 6528 1816 6532
rect 1818 6528 1819 6532
rect 1831 6528 1832 6532
rect 1834 6528 1835 6532
rect 1847 6528 1848 6532
rect 1850 6528 1853 6532
rect 1855 6528 1856 6532
rect 952 6514 953 6518
rect 955 6514 956 6518
rect 970 6514 971 6518
rect 973 6514 976 6518
rect 978 6514 983 6518
rect 995 6514 996 6518
rect 998 6514 999 6518
rect 1016 6514 1017 6518
rect 1019 6514 1021 6518
rect 1042 6514 1043 6518
rect 1045 6514 1048 6518
rect 1050 6514 1055 6518
rect 1070 6514 1071 6518
rect 1073 6514 1074 6518
rect 1086 6514 1087 6518
rect 1089 6514 1090 6518
rect 1111 6514 1112 6518
rect 1114 6514 1115 6518
rect 1119 6514 1125 6518
rect 1129 6514 1130 6518
rect 1132 6514 1133 6518
rect 1213 6514 1214 6518
rect 1216 6514 1217 6518
rect 1231 6514 1232 6518
rect 1234 6514 1237 6518
rect 1239 6514 1244 6518
rect 1256 6514 1257 6518
rect 1259 6514 1260 6518
rect 1277 6514 1278 6518
rect 1280 6514 1282 6518
rect 1303 6514 1304 6518
rect 1306 6514 1309 6518
rect 1311 6514 1316 6518
rect 1331 6514 1332 6518
rect 1334 6514 1335 6518
rect 1347 6514 1348 6518
rect 1350 6514 1351 6518
rect 1363 6514 1364 6518
rect 1366 6514 1367 6518
rect 2103 6521 2104 6525
rect 2106 6521 2109 6525
rect 2111 6521 2114 6525
rect 2417 6528 2418 6532
rect 2420 6528 2421 6532
rect 2433 6528 2434 6532
rect 2436 6528 2439 6532
rect 2441 6528 2442 6532
rect 2454 6528 2455 6532
rect 2457 6528 2458 6532
rect 2470 6528 2471 6532
rect 2473 6528 2474 6532
rect 2491 6528 2492 6532
rect 2494 6528 2497 6532
rect 2499 6528 2500 6532
rect 2512 6528 2513 6532
rect 2515 6528 2516 6532
rect 2528 6528 2529 6532
rect 2531 6528 2534 6532
rect 2536 6528 2537 6532
rect 2549 6528 2550 6532
rect 2552 6528 2553 6532
rect 2565 6528 2566 6532
rect 2568 6528 2571 6532
rect 2573 6528 2574 6532
rect 2586 6528 2587 6532
rect 2589 6528 2590 6532
rect 2602 6528 2603 6532
rect 2605 6528 2606 6532
rect 2623 6528 2624 6532
rect 2626 6528 2629 6532
rect 2631 6528 2632 6532
rect 2644 6528 2645 6532
rect 2647 6528 2648 6532
rect 2660 6528 2661 6532
rect 2663 6528 2666 6532
rect 2668 6528 2669 6532
rect 2681 6528 2682 6532
rect 2684 6528 2685 6532
rect 2697 6528 2698 6532
rect 2700 6528 2703 6532
rect 2705 6528 2706 6532
rect 2718 6528 2719 6532
rect 2721 6528 2722 6532
rect 2734 6528 2735 6532
rect 2737 6528 2738 6532
rect 2755 6528 2756 6532
rect 2758 6528 2761 6532
rect 2763 6528 2764 6532
rect 2776 6528 2777 6532
rect 2779 6528 2780 6532
rect 2792 6528 2793 6532
rect 2795 6528 2798 6532
rect 2800 6528 2801 6532
rect 1897 6514 1898 6518
rect 1900 6514 1901 6518
rect 1915 6514 1916 6518
rect 1918 6514 1921 6518
rect 1923 6514 1928 6518
rect 1940 6514 1941 6518
rect 1943 6514 1944 6518
rect 1961 6514 1962 6518
rect 1964 6514 1966 6518
rect 1987 6514 1988 6518
rect 1990 6514 1993 6518
rect 1995 6514 2000 6518
rect 2015 6514 2016 6518
rect 2018 6514 2019 6518
rect 2031 6514 2032 6518
rect 2034 6514 2035 6518
rect 2056 6514 2057 6518
rect 2059 6514 2060 6518
rect 2064 6514 2070 6518
rect 2074 6514 2075 6518
rect 2077 6514 2078 6518
rect 2158 6514 2159 6518
rect 2161 6514 2162 6518
rect 2176 6514 2177 6518
rect 2179 6514 2182 6518
rect 2184 6514 2189 6518
rect 2201 6514 2202 6518
rect 2204 6514 2205 6518
rect 2222 6514 2223 6518
rect 2225 6514 2227 6518
rect 2248 6514 2249 6518
rect 2251 6514 2254 6518
rect 2256 6514 2261 6518
rect 2276 6514 2277 6518
rect 2279 6514 2280 6518
rect 2292 6514 2293 6518
rect 2295 6514 2296 6518
rect 2308 6514 2309 6518
rect 2311 6514 2312 6518
rect 1213 6468 1214 6472
rect 1216 6468 1217 6472
rect 1231 6468 1232 6472
rect 1234 6468 1237 6472
rect 1239 6468 1244 6472
rect 1256 6468 1257 6472
rect 1259 6468 1260 6472
rect 1277 6468 1278 6472
rect 1280 6468 1282 6472
rect 1303 6468 1304 6472
rect 1306 6468 1309 6472
rect 1311 6468 1316 6472
rect 1331 6468 1332 6472
rect 1334 6468 1335 6472
rect 1347 6468 1348 6472
rect 1350 6468 1351 6472
rect 1363 6468 1364 6472
rect 1366 6468 1367 6472
rect 1135 6463 1136 6467
rect 1138 6463 1139 6467
rect 1158 6459 1159 6463
rect 1161 6459 1164 6463
rect 1166 6459 1169 6463
rect 2158 6468 2159 6472
rect 2161 6468 2162 6472
rect 2176 6468 2177 6472
rect 2179 6468 2182 6472
rect 2184 6468 2189 6472
rect 2201 6468 2202 6472
rect 2204 6468 2205 6472
rect 2222 6468 2223 6472
rect 2225 6468 2227 6472
rect 2248 6468 2249 6472
rect 2251 6468 2254 6472
rect 2256 6468 2261 6472
rect 2276 6468 2277 6472
rect 2279 6468 2280 6472
rect 2292 6468 2293 6472
rect 2295 6468 2296 6472
rect 2308 6468 2309 6472
rect 2311 6468 2312 6472
rect 2080 6463 2081 6467
rect 2083 6463 2084 6467
rect 2103 6459 2104 6463
rect 2106 6459 2109 6463
rect 2111 6459 2114 6463
rect 987 6385 988 6389
rect 990 6385 993 6389
rect 995 6385 998 6389
rect 1077 6385 1078 6389
rect 1080 6385 1083 6389
rect 1085 6385 1088 6389
rect 1158 6385 1159 6389
rect 1161 6385 1164 6389
rect 1166 6385 1169 6389
rect 1213 6382 1214 6386
rect 1216 6382 1217 6386
rect 1231 6382 1232 6386
rect 1234 6382 1237 6386
rect 1239 6382 1244 6386
rect 1256 6382 1257 6386
rect 1259 6382 1260 6386
rect 1277 6382 1278 6386
rect 1280 6382 1282 6386
rect 1303 6382 1304 6386
rect 1306 6382 1309 6386
rect 1311 6382 1316 6386
rect 1331 6382 1332 6386
rect 1334 6382 1335 6386
rect 1347 6382 1348 6386
rect 1350 6382 1351 6386
rect 1363 6382 1364 6386
rect 1366 6382 1367 6386
rect 1932 6385 1933 6389
rect 1935 6385 1938 6389
rect 1940 6385 1943 6389
rect 2022 6385 2023 6389
rect 2025 6385 2028 6389
rect 2030 6385 2033 6389
rect 2103 6385 2104 6389
rect 2106 6385 2109 6389
rect 2111 6385 2114 6389
rect 2158 6382 2159 6386
rect 2161 6382 2162 6386
rect 2176 6382 2177 6386
rect 2179 6382 2182 6386
rect 2184 6382 2189 6386
rect 2201 6382 2202 6386
rect 2204 6382 2205 6386
rect 2222 6382 2223 6386
rect 2225 6382 2227 6386
rect 2248 6382 2249 6386
rect 2251 6382 2254 6386
rect 2256 6382 2261 6386
rect 2276 6382 2277 6386
rect 2279 6382 2280 6386
rect 2292 6382 2293 6386
rect 2295 6382 2296 6386
rect 2308 6382 2309 6386
rect 2311 6382 2312 6386
rect 964 6331 965 6335
rect 967 6331 968 6335
rect 1054 6331 1055 6335
rect 1057 6331 1058 6335
rect 1213 6336 1214 6340
rect 1216 6336 1217 6340
rect 1231 6336 1232 6340
rect 1234 6336 1237 6340
rect 1239 6336 1244 6340
rect 1256 6336 1257 6340
rect 1259 6336 1260 6340
rect 1277 6336 1278 6340
rect 1280 6336 1282 6340
rect 1303 6336 1304 6340
rect 1306 6336 1309 6340
rect 1311 6336 1316 6340
rect 1331 6336 1332 6340
rect 1334 6336 1335 6340
rect 1347 6336 1348 6340
rect 1350 6336 1351 6340
rect 1363 6336 1364 6340
rect 1366 6336 1367 6340
rect 1135 6331 1136 6335
rect 1138 6331 1139 6335
rect 987 6327 988 6331
rect 990 6327 993 6331
rect 995 6327 998 6331
rect 1018 6323 1019 6327
rect 1021 6323 1022 6327
rect 1077 6327 1078 6331
rect 1080 6327 1083 6331
rect 1085 6327 1088 6331
rect 1108 6323 1109 6327
rect 1111 6323 1112 6327
rect 1158 6327 1159 6331
rect 1161 6327 1164 6331
rect 1166 6327 1169 6331
rect 1909 6331 1910 6335
rect 1912 6331 1913 6335
rect 1999 6331 2000 6335
rect 2002 6331 2003 6335
rect 2158 6336 2159 6340
rect 2161 6336 2162 6340
rect 2176 6336 2177 6340
rect 2179 6336 2182 6340
rect 2184 6336 2189 6340
rect 2201 6336 2202 6340
rect 2204 6336 2205 6340
rect 2222 6336 2223 6340
rect 2225 6336 2227 6340
rect 2248 6336 2249 6340
rect 2251 6336 2254 6340
rect 2256 6336 2261 6340
rect 2276 6336 2277 6340
rect 2279 6336 2280 6340
rect 2292 6336 2293 6340
rect 2295 6336 2296 6340
rect 2308 6336 2309 6340
rect 2311 6336 2312 6340
rect 2080 6331 2081 6335
rect 2083 6331 2084 6335
rect 1932 6327 1933 6331
rect 1935 6327 1938 6331
rect 1940 6327 1943 6331
rect 1963 6323 1964 6327
rect 1966 6323 1967 6327
rect 2022 6327 2023 6331
rect 2025 6327 2028 6331
rect 2030 6327 2033 6331
rect 2053 6323 2054 6327
rect 2056 6323 2057 6327
rect 2103 6327 2104 6331
rect 2106 6327 2109 6331
rect 2111 6327 2114 6331
rect 1053 6250 1054 6254
rect 1056 6250 1059 6254
rect 1061 6250 1064 6254
rect 1158 6250 1159 6254
rect 1161 6250 1164 6254
rect 1166 6250 1169 6254
rect 1213 6250 1214 6254
rect 1216 6250 1217 6254
rect 1231 6250 1232 6254
rect 1234 6250 1237 6254
rect 1239 6250 1244 6254
rect 1256 6250 1257 6254
rect 1259 6250 1260 6254
rect 1277 6250 1278 6254
rect 1280 6250 1282 6254
rect 1303 6250 1304 6254
rect 1306 6250 1309 6254
rect 1311 6250 1316 6254
rect 1331 6250 1332 6254
rect 1334 6250 1335 6254
rect 1347 6250 1348 6254
rect 1350 6250 1351 6254
rect 1363 6250 1364 6254
rect 1366 6250 1367 6254
rect 1998 6250 1999 6254
rect 2001 6250 2004 6254
rect 2006 6250 2009 6254
rect 2103 6250 2104 6254
rect 2106 6250 2109 6254
rect 2111 6250 2114 6254
rect 2158 6250 2159 6254
rect 2161 6250 2162 6254
rect 2176 6250 2177 6254
rect 2179 6250 2182 6254
rect 2184 6250 2189 6254
rect 2201 6250 2202 6254
rect 2204 6250 2205 6254
rect 2222 6250 2223 6254
rect 2225 6250 2227 6254
rect 2248 6250 2249 6254
rect 2251 6250 2254 6254
rect 2256 6250 2261 6254
rect 2276 6250 2277 6254
rect 2279 6250 2280 6254
rect 2292 6250 2293 6254
rect 2295 6250 2296 6254
rect 2308 6250 2309 6254
rect 2311 6250 2312 6254
rect 1030 6199 1031 6203
rect 1033 6199 1034 6203
rect 1213 6204 1214 6208
rect 1216 6204 1217 6208
rect 1231 6204 1232 6208
rect 1234 6204 1237 6208
rect 1239 6204 1244 6208
rect 1256 6204 1257 6208
rect 1259 6204 1260 6208
rect 1277 6204 1278 6208
rect 1280 6204 1282 6208
rect 1303 6204 1304 6208
rect 1306 6204 1309 6208
rect 1311 6204 1316 6208
rect 1331 6204 1332 6208
rect 1334 6204 1335 6208
rect 1347 6204 1348 6208
rect 1350 6204 1351 6208
rect 1363 6204 1364 6208
rect 1366 6204 1367 6208
rect 1135 6199 1136 6203
rect 1138 6199 1139 6203
rect 1053 6195 1054 6199
rect 1056 6195 1059 6199
rect 1061 6195 1064 6199
rect 1084 6191 1085 6195
rect 1087 6191 1088 6195
rect 1158 6195 1159 6199
rect 1161 6195 1164 6199
rect 1166 6195 1169 6199
rect 1975 6199 1976 6203
rect 1978 6199 1979 6203
rect 2158 6204 2159 6208
rect 2161 6204 2162 6208
rect 2176 6204 2177 6208
rect 2179 6204 2182 6208
rect 2184 6204 2189 6208
rect 2201 6204 2202 6208
rect 2204 6204 2205 6208
rect 2222 6204 2223 6208
rect 2225 6204 2227 6208
rect 2248 6204 2249 6208
rect 2251 6204 2254 6208
rect 2256 6204 2261 6208
rect 2276 6204 2277 6208
rect 2279 6204 2280 6208
rect 2292 6204 2293 6208
rect 2295 6204 2296 6208
rect 2308 6204 2309 6208
rect 2311 6204 2312 6208
rect 2080 6199 2081 6203
rect 2083 6199 2084 6203
rect 1998 6195 1999 6199
rect 2001 6195 2004 6199
rect 2006 6195 2009 6199
rect 2029 6191 2030 6195
rect 2032 6191 2033 6195
rect 2103 6195 2104 6199
rect 2106 6195 2109 6199
rect 2111 6195 2114 6199
rect 1077 6119 1078 6123
rect 1080 6119 1083 6123
rect 1085 6119 1088 6123
rect 1158 6119 1159 6123
rect 1161 6119 1164 6123
rect 1166 6119 1169 6123
rect 1613 6128 1614 6132
rect 1616 6128 1619 6132
rect 1621 6128 1622 6132
rect 1634 6128 1635 6132
rect 1637 6128 1638 6132
rect 1650 6128 1651 6132
rect 1653 6128 1656 6132
rect 1658 6128 1659 6132
rect 1676 6128 1677 6132
rect 1679 6128 1680 6132
rect 1692 6128 1693 6132
rect 1695 6128 1696 6132
rect 1708 6128 1709 6132
rect 1711 6128 1714 6132
rect 1716 6128 1717 6132
rect 1729 6128 1730 6132
rect 1732 6128 1733 6132
rect 1213 6118 1214 6122
rect 1216 6118 1217 6122
rect 1231 6118 1232 6122
rect 1234 6118 1237 6122
rect 1239 6118 1244 6122
rect 1256 6118 1257 6122
rect 1259 6118 1260 6122
rect 1277 6118 1278 6122
rect 1280 6118 1282 6122
rect 1303 6118 1304 6122
rect 1306 6118 1309 6122
rect 1311 6118 1316 6122
rect 1331 6118 1332 6122
rect 1334 6118 1335 6122
rect 1347 6118 1348 6122
rect 1350 6118 1351 6122
rect 1363 6118 1364 6122
rect 1366 6118 1367 6122
rect 2022 6119 2023 6123
rect 2025 6119 2028 6123
rect 2030 6119 2033 6123
rect 2103 6119 2104 6123
rect 2106 6119 2109 6123
rect 2111 6119 2114 6123
rect 2558 6128 2559 6132
rect 2561 6128 2564 6132
rect 2566 6128 2567 6132
rect 2579 6128 2580 6132
rect 2582 6128 2583 6132
rect 2595 6128 2596 6132
rect 2598 6128 2601 6132
rect 2603 6128 2604 6132
rect 2621 6128 2622 6132
rect 2624 6128 2625 6132
rect 2637 6128 2638 6132
rect 2640 6128 2641 6132
rect 2653 6128 2654 6132
rect 2656 6128 2659 6132
rect 2661 6128 2662 6132
rect 2674 6128 2675 6132
rect 2677 6128 2678 6132
rect 2158 6118 2159 6122
rect 2161 6118 2162 6122
rect 2176 6118 2177 6122
rect 2179 6118 2182 6122
rect 2184 6118 2189 6122
rect 2201 6118 2202 6122
rect 2204 6118 2205 6122
rect 2222 6118 2223 6122
rect 2225 6118 2227 6122
rect 2248 6118 2249 6122
rect 2251 6118 2254 6122
rect 2256 6118 2261 6122
rect 2276 6118 2277 6122
rect 2279 6118 2280 6122
rect 2292 6118 2293 6122
rect 2295 6118 2296 6122
rect 2308 6118 2309 6122
rect 2311 6118 2312 6122
rect 1054 6067 1055 6071
rect 1057 6067 1058 6071
rect 1213 6072 1214 6076
rect 1216 6072 1217 6076
rect 1231 6072 1232 6076
rect 1234 6072 1237 6076
rect 1239 6072 1244 6076
rect 1256 6072 1257 6076
rect 1259 6072 1260 6076
rect 1277 6072 1278 6076
rect 1280 6072 1282 6076
rect 1303 6072 1304 6076
rect 1306 6072 1309 6076
rect 1311 6072 1316 6076
rect 1331 6072 1332 6076
rect 1334 6072 1335 6076
rect 1347 6072 1348 6076
rect 1350 6072 1351 6076
rect 1363 6072 1364 6076
rect 1366 6072 1367 6076
rect 1713 6072 1714 6076
rect 1716 6072 1717 6076
rect 1135 6067 1136 6071
rect 1138 6067 1139 6071
rect 1077 6063 1078 6067
rect 1080 6063 1083 6067
rect 1085 6063 1088 6067
rect 1108 6059 1109 6063
rect 1111 6059 1112 6063
rect 1158 6063 1159 6067
rect 1161 6063 1164 6067
rect 1166 6063 1169 6067
rect 1189 6059 1190 6063
rect 1192 6059 1193 6063
rect 1596 6063 1597 6067
rect 1599 6063 1600 6067
rect 1999 6067 2000 6071
rect 2002 6067 2003 6071
rect 2158 6072 2159 6076
rect 2161 6072 2162 6076
rect 2176 6072 2177 6076
rect 2179 6072 2182 6076
rect 2184 6072 2189 6076
rect 2201 6072 2202 6076
rect 2204 6072 2205 6076
rect 2222 6072 2223 6076
rect 2225 6072 2227 6076
rect 2248 6072 2249 6076
rect 2251 6072 2254 6076
rect 2256 6072 2261 6076
rect 2276 6072 2277 6076
rect 2279 6072 2280 6076
rect 2292 6072 2293 6076
rect 2295 6072 2296 6076
rect 2308 6072 2309 6076
rect 2311 6072 2312 6076
rect 2658 6072 2659 6076
rect 2661 6072 2662 6076
rect 2080 6067 2081 6071
rect 2083 6067 2084 6071
rect 2022 6063 2023 6067
rect 2025 6063 2028 6067
rect 2030 6063 2033 6067
rect 2053 6059 2054 6063
rect 2056 6059 2057 6063
rect 2103 6063 2104 6067
rect 2106 6063 2109 6067
rect 2111 6063 2114 6067
rect 2134 6059 2135 6063
rect 2137 6059 2138 6063
rect 2541 6063 2542 6067
rect 2544 6063 2545 6067
rect 1604 6026 1605 6030
rect 1607 6026 1608 6030
rect 1620 6026 1621 6030
rect 1623 6026 1626 6030
rect 1628 6026 1629 6030
rect 1641 6026 1642 6030
rect 1644 6026 1645 6030
rect 1657 6026 1658 6030
rect 1660 6026 1661 6030
rect 1678 6026 1679 6030
rect 1681 6026 1684 6030
rect 1686 6026 1687 6030
rect 1699 6026 1700 6030
rect 1702 6026 1703 6030
rect 1715 6026 1716 6030
rect 1718 6026 1721 6030
rect 1723 6026 1724 6030
rect 2549 6026 2550 6030
rect 2552 6026 2553 6030
rect 2565 6026 2566 6030
rect 2568 6026 2571 6030
rect 2573 6026 2574 6030
rect 2586 6026 2587 6030
rect 2589 6026 2590 6030
rect 2602 6026 2603 6030
rect 2605 6026 2606 6030
rect 2623 6026 2624 6030
rect 2626 6026 2629 6030
rect 2631 6026 2632 6030
rect 2644 6026 2645 6030
rect 2647 6026 2648 6030
rect 2660 6026 2661 6030
rect 2663 6026 2666 6030
rect 2668 6026 2669 6030
rect 856 5993 857 5997
rect 859 5993 860 5997
rect 872 5993 873 5997
rect 875 5993 878 5997
rect 880 5993 881 5997
rect 893 5993 894 5997
rect 896 5993 897 5997
rect 909 5993 910 5997
rect 912 5993 913 5997
rect 930 5993 931 5997
rect 933 5993 936 5997
rect 938 5993 939 5997
rect 951 5993 952 5997
rect 954 5993 955 5997
rect 967 5993 968 5997
rect 970 5993 973 5997
rect 975 5993 976 5997
rect 988 5993 989 5997
rect 991 5993 992 5997
rect 1004 5993 1005 5997
rect 1007 5993 1010 5997
rect 1012 5993 1013 5997
rect 1025 5993 1026 5997
rect 1028 5993 1029 5997
rect 1041 5993 1042 5997
rect 1044 5993 1045 5997
rect 1062 5993 1063 5997
rect 1065 5993 1068 5997
rect 1070 5993 1071 5997
rect 1083 5993 1084 5997
rect 1086 5993 1087 5997
rect 1099 5993 1100 5997
rect 1102 5993 1105 5997
rect 1107 5993 1108 5997
rect 1120 5993 1121 5997
rect 1123 5993 1124 5997
rect 1136 5993 1137 5997
rect 1139 5993 1142 5997
rect 1144 5993 1145 5997
rect 1157 5993 1158 5997
rect 1160 5993 1161 5997
rect 1173 5993 1174 5997
rect 1176 5993 1177 5997
rect 1194 5993 1195 5997
rect 1197 5993 1200 5997
rect 1202 5993 1203 5997
rect 1215 5993 1216 5997
rect 1218 5993 1219 5997
rect 1231 5993 1232 5997
rect 1234 5993 1237 5997
rect 1239 5993 1240 5997
rect 1252 5993 1253 5997
rect 1255 5993 1256 5997
rect 1268 5993 1269 5997
rect 1271 5993 1274 5997
rect 1276 5993 1277 5997
rect 1289 5993 1290 5997
rect 1292 5993 1293 5997
rect 1305 5993 1306 5997
rect 1308 5993 1309 5997
rect 1326 5993 1327 5997
rect 1329 5993 1332 5997
rect 1334 5993 1335 5997
rect 1347 5993 1348 5997
rect 1350 5993 1351 5997
rect 1363 5993 1364 5997
rect 1366 5993 1369 5997
rect 1371 5993 1372 5997
rect 1801 5993 1802 5997
rect 1804 5993 1805 5997
rect 1817 5993 1818 5997
rect 1820 5993 1823 5997
rect 1825 5993 1826 5997
rect 1838 5993 1839 5997
rect 1841 5993 1842 5997
rect 1854 5993 1855 5997
rect 1857 5993 1858 5997
rect 1875 5993 1876 5997
rect 1878 5993 1881 5997
rect 1883 5993 1884 5997
rect 1896 5993 1897 5997
rect 1899 5993 1900 5997
rect 1912 5993 1913 5997
rect 1915 5993 1918 5997
rect 1920 5993 1921 5997
rect 1933 5993 1934 5997
rect 1936 5993 1937 5997
rect 1949 5993 1950 5997
rect 1952 5993 1955 5997
rect 1957 5993 1958 5997
rect 1970 5993 1971 5997
rect 1973 5993 1974 5997
rect 1986 5993 1987 5997
rect 1989 5993 1990 5997
rect 2007 5993 2008 5997
rect 2010 5993 2013 5997
rect 2015 5993 2016 5997
rect 2028 5993 2029 5997
rect 2031 5993 2032 5997
rect 2044 5993 2045 5997
rect 2047 5993 2050 5997
rect 2052 5993 2053 5997
rect 2065 5993 2066 5997
rect 2068 5993 2069 5997
rect 2081 5993 2082 5997
rect 2084 5993 2087 5997
rect 2089 5993 2090 5997
rect 2102 5993 2103 5997
rect 2105 5993 2106 5997
rect 2118 5993 2119 5997
rect 2121 5993 2122 5997
rect 2139 5993 2140 5997
rect 2142 5993 2145 5997
rect 2147 5993 2148 5997
rect 2160 5993 2161 5997
rect 2163 5993 2164 5997
rect 2176 5993 2177 5997
rect 2179 5993 2182 5997
rect 2184 5993 2185 5997
rect 2197 5993 2198 5997
rect 2200 5993 2201 5997
rect 2213 5993 2214 5997
rect 2216 5993 2219 5997
rect 2221 5993 2222 5997
rect 2234 5993 2235 5997
rect 2237 5993 2238 5997
rect 2250 5993 2251 5997
rect 2253 5993 2254 5997
rect 2271 5993 2272 5997
rect 2274 5993 2277 5997
rect 2279 5993 2280 5997
rect 2292 5993 2293 5997
rect 2295 5993 2296 5997
rect 2308 5993 2309 5997
rect 2311 5993 2314 5997
rect 2316 5993 2317 5997
rect 1472 5914 1473 5918
rect 1475 5914 1476 5918
rect 1488 5914 1489 5918
rect 1491 5914 1494 5918
rect 1496 5914 1497 5918
rect 1509 5914 1510 5918
rect 1512 5914 1513 5918
rect 1525 5914 1526 5918
rect 1528 5914 1529 5918
rect 1546 5914 1547 5918
rect 1549 5914 1552 5918
rect 1554 5914 1555 5918
rect 1567 5914 1568 5918
rect 1570 5914 1571 5918
rect 1583 5914 1584 5918
rect 1586 5914 1589 5918
rect 1591 5914 1592 5918
rect 1604 5914 1605 5918
rect 1607 5914 1608 5918
rect 1620 5914 1621 5918
rect 1623 5914 1626 5918
rect 1628 5914 1629 5918
rect 1641 5914 1642 5918
rect 1644 5914 1645 5918
rect 1657 5914 1658 5918
rect 1660 5914 1661 5918
rect 1678 5914 1679 5918
rect 1681 5914 1684 5918
rect 1686 5914 1687 5918
rect 1699 5914 1700 5918
rect 1702 5914 1703 5918
rect 1715 5914 1716 5918
rect 1718 5914 1721 5918
rect 1723 5914 1724 5918
rect 1736 5914 1737 5918
rect 1739 5914 1740 5918
rect 1752 5914 1753 5918
rect 1755 5914 1758 5918
rect 1760 5914 1761 5918
rect 1773 5914 1774 5918
rect 1776 5914 1777 5918
rect 1789 5914 1790 5918
rect 1792 5914 1793 5918
rect 1810 5914 1811 5918
rect 1813 5914 1816 5918
rect 1818 5914 1819 5918
rect 1831 5914 1832 5918
rect 1834 5914 1835 5918
rect 1847 5914 1848 5918
rect 1850 5914 1853 5918
rect 1855 5914 1856 5918
rect 2417 5914 2418 5918
rect 2420 5914 2421 5918
rect 2433 5914 2434 5918
rect 2436 5914 2439 5918
rect 2441 5914 2442 5918
rect 2454 5914 2455 5918
rect 2457 5914 2458 5918
rect 2470 5914 2471 5918
rect 2473 5914 2474 5918
rect 2491 5914 2492 5918
rect 2494 5914 2497 5918
rect 2499 5914 2500 5918
rect 2512 5914 2513 5918
rect 2515 5914 2516 5918
rect 2528 5914 2529 5918
rect 2531 5914 2534 5918
rect 2536 5914 2537 5918
rect 2549 5914 2550 5918
rect 2552 5914 2553 5918
rect 2565 5914 2566 5918
rect 2568 5914 2571 5918
rect 2573 5914 2574 5918
rect 2586 5914 2587 5918
rect 2589 5914 2590 5918
rect 2602 5914 2603 5918
rect 2605 5914 2606 5918
rect 2623 5914 2624 5918
rect 2626 5914 2629 5918
rect 2631 5914 2632 5918
rect 2644 5914 2645 5918
rect 2647 5914 2648 5918
rect 2660 5914 2661 5918
rect 2663 5914 2666 5918
rect 2668 5914 2669 5918
rect 2681 5914 2682 5918
rect 2684 5914 2685 5918
rect 2697 5914 2698 5918
rect 2700 5914 2703 5918
rect 2705 5914 2706 5918
rect 2718 5914 2719 5918
rect 2721 5914 2722 5918
rect 2734 5914 2735 5918
rect 2737 5914 2738 5918
rect 2755 5914 2756 5918
rect 2758 5914 2761 5918
rect 2763 5914 2764 5918
rect 2776 5914 2777 5918
rect 2779 5914 2780 5918
rect 2792 5914 2793 5918
rect 2795 5914 2798 5918
rect 2800 5914 2801 5918
rect 1596 5852 1597 5856
rect 1599 5852 1600 5856
rect 1620 5852 1621 5856
rect 1623 5852 1624 5856
rect 2541 5852 2542 5856
rect 2544 5852 2545 5856
rect 2565 5852 2566 5856
rect 2568 5852 2569 5856
rect 1608 5847 1612 5848
rect 1608 5844 1612 5845
rect 2553 5847 2557 5848
rect 2553 5844 2557 5845
rect 1600 5829 1601 5833
rect 1603 5829 1604 5833
rect 2545 5829 2546 5833
rect 2548 5829 2549 5833
rect 1596 5818 1597 5822
rect 1599 5818 1600 5822
rect 1620 5818 1621 5822
rect 1623 5818 1624 5822
rect 2541 5818 2542 5822
rect 2544 5818 2545 5822
rect 2565 5818 2566 5822
rect 2568 5818 2569 5822
rect 1472 5774 1473 5778
rect 1475 5774 1476 5778
rect 1488 5774 1489 5778
rect 1491 5774 1494 5778
rect 1496 5774 1497 5778
rect 1509 5774 1510 5778
rect 1512 5774 1513 5778
rect 1525 5774 1526 5778
rect 1528 5774 1529 5778
rect 1546 5774 1547 5778
rect 1549 5774 1552 5778
rect 1554 5774 1555 5778
rect 1567 5774 1568 5778
rect 1570 5774 1571 5778
rect 1583 5774 1584 5778
rect 1586 5774 1589 5778
rect 1591 5774 1592 5778
rect 1604 5774 1605 5778
rect 1607 5774 1608 5778
rect 1620 5774 1621 5778
rect 1623 5774 1626 5778
rect 1628 5774 1629 5778
rect 1641 5774 1642 5778
rect 1644 5774 1645 5778
rect 1657 5774 1658 5778
rect 1660 5774 1661 5778
rect 1678 5774 1679 5778
rect 1681 5774 1684 5778
rect 1686 5774 1687 5778
rect 1699 5774 1700 5778
rect 1702 5774 1703 5778
rect 1715 5774 1716 5778
rect 1718 5774 1721 5778
rect 1723 5774 1724 5778
rect 1736 5774 1737 5778
rect 1739 5774 1740 5778
rect 1752 5774 1753 5778
rect 1755 5774 1758 5778
rect 1760 5774 1761 5778
rect 1773 5774 1774 5778
rect 1776 5774 1777 5778
rect 1789 5774 1790 5778
rect 1792 5774 1793 5778
rect 1810 5774 1811 5778
rect 1813 5774 1816 5778
rect 1818 5774 1819 5778
rect 1831 5774 1832 5778
rect 1834 5774 1835 5778
rect 1847 5774 1848 5778
rect 1850 5774 1853 5778
rect 1855 5774 1856 5778
rect 2417 5774 2418 5778
rect 2420 5774 2421 5778
rect 2433 5774 2434 5778
rect 2436 5774 2439 5778
rect 2441 5774 2442 5778
rect 2454 5774 2455 5778
rect 2457 5774 2458 5778
rect 2470 5774 2471 5778
rect 2473 5774 2474 5778
rect 2491 5774 2492 5778
rect 2494 5774 2497 5778
rect 2499 5774 2500 5778
rect 2512 5774 2513 5778
rect 2515 5774 2516 5778
rect 2528 5774 2529 5778
rect 2531 5774 2534 5778
rect 2536 5774 2537 5778
rect 2549 5774 2550 5778
rect 2552 5774 2553 5778
rect 2565 5774 2566 5778
rect 2568 5774 2571 5778
rect 2573 5774 2574 5778
rect 2586 5774 2587 5778
rect 2589 5774 2590 5778
rect 2602 5774 2603 5778
rect 2605 5774 2606 5778
rect 2623 5774 2624 5778
rect 2626 5774 2629 5778
rect 2631 5774 2632 5778
rect 2644 5774 2645 5778
rect 2647 5774 2648 5778
rect 2660 5774 2661 5778
rect 2663 5774 2666 5778
rect 2668 5774 2669 5778
rect 2681 5774 2682 5778
rect 2684 5774 2685 5778
rect 2697 5774 2698 5778
rect 2700 5774 2703 5778
rect 2705 5774 2706 5778
rect 2718 5774 2719 5778
rect 2721 5774 2722 5778
rect 2734 5774 2735 5778
rect 2737 5774 2738 5778
rect 2755 5774 2756 5778
rect 2758 5774 2761 5778
rect 2763 5774 2764 5778
rect 2776 5774 2777 5778
rect 2779 5774 2780 5778
rect 2792 5774 2793 5778
rect 2795 5774 2798 5778
rect 2800 5774 2801 5778
rect 953 5744 954 5748
rect 956 5744 957 5748
rect 969 5744 970 5748
rect 972 5744 975 5748
rect 977 5744 978 5748
rect 990 5744 991 5748
rect 993 5744 994 5748
rect 1006 5744 1007 5748
rect 1009 5744 1010 5748
rect 1027 5744 1028 5748
rect 1030 5744 1033 5748
rect 1035 5744 1036 5748
rect 1048 5744 1049 5748
rect 1051 5744 1052 5748
rect 1064 5744 1065 5748
rect 1067 5744 1070 5748
rect 1072 5744 1073 5748
rect 1898 5744 1899 5748
rect 1901 5744 1902 5748
rect 1914 5744 1915 5748
rect 1917 5744 1920 5748
rect 1922 5744 1923 5748
rect 1935 5744 1936 5748
rect 1938 5744 1939 5748
rect 1951 5744 1952 5748
rect 1954 5744 1955 5748
rect 1972 5744 1973 5748
rect 1975 5744 1978 5748
rect 1980 5744 1981 5748
rect 1993 5744 1994 5748
rect 1996 5744 1997 5748
rect 2009 5744 2010 5748
rect 2012 5744 2015 5748
rect 2017 5744 2018 5748
rect 927 5738 931 5739
rect 927 5735 931 5736
rect 1872 5738 1876 5739
rect 1872 5735 1876 5736
rect 1472 5688 1473 5692
rect 1475 5688 1476 5692
rect 1488 5688 1489 5692
rect 1491 5688 1494 5692
rect 1496 5688 1497 5692
rect 1509 5688 1510 5692
rect 1512 5688 1513 5692
rect 1525 5688 1526 5692
rect 1528 5688 1529 5692
rect 1546 5688 1547 5692
rect 1549 5688 1552 5692
rect 1554 5688 1555 5692
rect 1567 5688 1568 5692
rect 1570 5688 1571 5692
rect 1583 5688 1584 5692
rect 1586 5688 1589 5692
rect 1591 5688 1592 5692
rect 1604 5688 1605 5692
rect 1607 5688 1608 5692
rect 1620 5688 1621 5692
rect 1623 5688 1626 5692
rect 1628 5688 1629 5692
rect 1641 5688 1642 5692
rect 1644 5688 1645 5692
rect 1657 5688 1658 5692
rect 1660 5688 1661 5692
rect 1678 5688 1679 5692
rect 1681 5688 1684 5692
rect 1686 5688 1687 5692
rect 1699 5688 1700 5692
rect 1702 5688 1703 5692
rect 1715 5688 1716 5692
rect 1718 5688 1721 5692
rect 1723 5688 1724 5692
rect 1736 5688 1737 5692
rect 1739 5688 1740 5692
rect 1752 5688 1753 5692
rect 1755 5688 1758 5692
rect 1760 5688 1761 5692
rect 1773 5688 1774 5692
rect 1776 5688 1777 5692
rect 1789 5688 1790 5692
rect 1792 5688 1793 5692
rect 1810 5688 1811 5692
rect 1813 5688 1816 5692
rect 1818 5688 1819 5692
rect 1831 5688 1832 5692
rect 1834 5688 1835 5692
rect 1847 5688 1848 5692
rect 1850 5688 1853 5692
rect 1855 5688 1856 5692
rect 2417 5688 2418 5692
rect 2420 5688 2421 5692
rect 2433 5688 2434 5692
rect 2436 5688 2439 5692
rect 2441 5688 2442 5692
rect 2454 5688 2455 5692
rect 2457 5688 2458 5692
rect 2470 5688 2471 5692
rect 2473 5688 2474 5692
rect 2491 5688 2492 5692
rect 2494 5688 2497 5692
rect 2499 5688 2500 5692
rect 2512 5688 2513 5692
rect 2515 5688 2516 5692
rect 2528 5688 2529 5692
rect 2531 5688 2534 5692
rect 2536 5688 2537 5692
rect 2549 5688 2550 5692
rect 2552 5688 2553 5692
rect 2565 5688 2566 5692
rect 2568 5688 2571 5692
rect 2573 5688 2574 5692
rect 2586 5688 2587 5692
rect 2589 5688 2590 5692
rect 2602 5688 2603 5692
rect 2605 5688 2606 5692
rect 2623 5688 2624 5692
rect 2626 5688 2629 5692
rect 2631 5688 2632 5692
rect 2644 5688 2645 5692
rect 2647 5688 2648 5692
rect 2660 5688 2661 5692
rect 2663 5688 2666 5692
rect 2668 5688 2669 5692
rect 2681 5688 2682 5692
rect 2684 5688 2685 5692
rect 2697 5688 2698 5692
rect 2700 5688 2703 5692
rect 2705 5688 2706 5692
rect 2718 5688 2719 5692
rect 2721 5688 2722 5692
rect 2734 5688 2735 5692
rect 2737 5688 2738 5692
rect 2755 5688 2756 5692
rect 2758 5688 2761 5692
rect 2763 5688 2764 5692
rect 2776 5688 2777 5692
rect 2779 5688 2780 5692
rect 2792 5688 2793 5692
rect 2795 5688 2798 5692
rect 2800 5688 2801 5692
rect 953 5658 954 5662
rect 956 5658 957 5662
rect 969 5658 970 5662
rect 972 5658 975 5662
rect 977 5658 978 5662
rect 990 5658 991 5662
rect 993 5658 994 5662
rect 1006 5658 1007 5662
rect 1009 5658 1010 5662
rect 1027 5658 1028 5662
rect 1030 5658 1033 5662
rect 1035 5658 1036 5662
rect 1048 5658 1049 5662
rect 1051 5658 1052 5662
rect 1064 5658 1065 5662
rect 1067 5658 1070 5662
rect 1072 5658 1073 5662
rect 1898 5658 1899 5662
rect 1901 5658 1902 5662
rect 1914 5658 1915 5662
rect 1917 5658 1920 5662
rect 1922 5658 1923 5662
rect 1935 5658 1936 5662
rect 1938 5658 1939 5662
rect 1951 5658 1952 5662
rect 1954 5658 1955 5662
rect 1972 5658 1973 5662
rect 1975 5658 1978 5662
rect 1980 5658 1981 5662
rect 1993 5658 1994 5662
rect 1996 5658 1997 5662
rect 2009 5658 2010 5662
rect 2012 5658 2015 5662
rect 2017 5658 2018 5662
rect 1713 5626 1714 5630
rect 1716 5626 1717 5630
rect 1737 5626 1738 5630
rect 1740 5626 1741 5630
rect 2658 5626 2659 5630
rect 2661 5626 2662 5630
rect 2682 5626 2683 5630
rect 2685 5626 2686 5630
rect 1725 5621 1729 5622
rect 1725 5618 1729 5619
rect 2670 5621 2674 5622
rect 2670 5618 2674 5619
rect 1717 5603 1718 5607
rect 1720 5603 1721 5607
rect 2662 5603 2663 5607
rect 2665 5603 2666 5607
rect 939 5592 943 5593
rect 939 5589 943 5590
rect 1713 5590 1714 5594
rect 1716 5590 1717 5594
rect 1737 5590 1738 5594
rect 1740 5590 1741 5594
rect 1884 5592 1888 5593
rect 1884 5589 1888 5590
rect 2658 5590 2659 5594
rect 2661 5590 2662 5594
rect 2682 5590 2683 5594
rect 2685 5590 2686 5594
rect 1158 5539 1159 5543
rect 1161 5539 1164 5543
rect 1166 5539 1169 5543
rect 1472 5546 1473 5550
rect 1475 5546 1476 5550
rect 1488 5546 1489 5550
rect 1491 5546 1494 5550
rect 1496 5546 1497 5550
rect 1509 5546 1510 5550
rect 1512 5546 1513 5550
rect 1525 5546 1526 5550
rect 1528 5546 1529 5550
rect 1546 5546 1547 5550
rect 1549 5546 1552 5550
rect 1554 5546 1555 5550
rect 1567 5546 1568 5550
rect 1570 5546 1571 5550
rect 1583 5546 1584 5550
rect 1586 5546 1589 5550
rect 1591 5546 1592 5550
rect 1604 5546 1605 5550
rect 1607 5546 1608 5550
rect 1620 5546 1621 5550
rect 1623 5546 1626 5550
rect 1628 5546 1629 5550
rect 1641 5546 1642 5550
rect 1644 5546 1645 5550
rect 1657 5546 1658 5550
rect 1660 5546 1661 5550
rect 1678 5546 1679 5550
rect 1681 5546 1684 5550
rect 1686 5546 1687 5550
rect 1699 5546 1700 5550
rect 1702 5546 1703 5550
rect 1715 5546 1716 5550
rect 1718 5546 1721 5550
rect 1723 5546 1724 5550
rect 1736 5546 1737 5550
rect 1739 5546 1740 5550
rect 1752 5546 1753 5550
rect 1755 5546 1758 5550
rect 1760 5546 1761 5550
rect 1773 5546 1774 5550
rect 1776 5546 1777 5550
rect 1789 5546 1790 5550
rect 1792 5546 1793 5550
rect 1810 5546 1811 5550
rect 1813 5546 1816 5550
rect 1818 5546 1819 5550
rect 1831 5546 1832 5550
rect 1834 5546 1835 5550
rect 1847 5546 1848 5550
rect 1850 5546 1853 5550
rect 1855 5546 1856 5550
rect 952 5532 953 5536
rect 955 5532 956 5536
rect 970 5532 971 5536
rect 973 5532 976 5536
rect 978 5532 983 5536
rect 995 5532 996 5536
rect 998 5532 999 5536
rect 1016 5532 1017 5536
rect 1019 5532 1021 5536
rect 1042 5532 1043 5536
rect 1045 5532 1048 5536
rect 1050 5532 1055 5536
rect 1070 5532 1071 5536
rect 1073 5532 1074 5536
rect 1086 5532 1087 5536
rect 1089 5532 1090 5536
rect 1111 5532 1112 5536
rect 1114 5532 1115 5536
rect 1119 5532 1125 5536
rect 1129 5532 1130 5536
rect 1132 5532 1133 5536
rect 1213 5532 1214 5536
rect 1216 5532 1217 5536
rect 1231 5532 1232 5536
rect 1234 5532 1237 5536
rect 1239 5532 1244 5536
rect 1256 5532 1257 5536
rect 1259 5532 1260 5536
rect 1277 5532 1278 5536
rect 1280 5532 1282 5536
rect 1303 5532 1304 5536
rect 1306 5532 1309 5536
rect 1311 5532 1316 5536
rect 1331 5532 1332 5536
rect 1334 5532 1335 5536
rect 1347 5532 1348 5536
rect 1350 5532 1351 5536
rect 1363 5532 1364 5536
rect 1366 5532 1367 5536
rect 2103 5539 2104 5543
rect 2106 5539 2109 5543
rect 2111 5539 2114 5543
rect 2417 5546 2418 5550
rect 2420 5546 2421 5550
rect 2433 5546 2434 5550
rect 2436 5546 2439 5550
rect 2441 5546 2442 5550
rect 2454 5546 2455 5550
rect 2457 5546 2458 5550
rect 2470 5546 2471 5550
rect 2473 5546 2474 5550
rect 2491 5546 2492 5550
rect 2494 5546 2497 5550
rect 2499 5546 2500 5550
rect 2512 5546 2513 5550
rect 2515 5546 2516 5550
rect 2528 5546 2529 5550
rect 2531 5546 2534 5550
rect 2536 5546 2537 5550
rect 2549 5546 2550 5550
rect 2552 5546 2553 5550
rect 2565 5546 2566 5550
rect 2568 5546 2571 5550
rect 2573 5546 2574 5550
rect 2586 5546 2587 5550
rect 2589 5546 2590 5550
rect 2602 5546 2603 5550
rect 2605 5546 2606 5550
rect 2623 5546 2624 5550
rect 2626 5546 2629 5550
rect 2631 5546 2632 5550
rect 2644 5546 2645 5550
rect 2647 5546 2648 5550
rect 2660 5546 2661 5550
rect 2663 5546 2666 5550
rect 2668 5546 2669 5550
rect 2681 5546 2682 5550
rect 2684 5546 2685 5550
rect 2697 5546 2698 5550
rect 2700 5546 2703 5550
rect 2705 5546 2706 5550
rect 2718 5546 2719 5550
rect 2721 5546 2722 5550
rect 2734 5546 2735 5550
rect 2737 5546 2738 5550
rect 2755 5546 2756 5550
rect 2758 5546 2761 5550
rect 2763 5546 2764 5550
rect 2776 5546 2777 5550
rect 2779 5546 2780 5550
rect 2792 5546 2793 5550
rect 2795 5546 2798 5550
rect 2800 5546 2801 5550
rect 1897 5532 1898 5536
rect 1900 5532 1901 5536
rect 1915 5532 1916 5536
rect 1918 5532 1921 5536
rect 1923 5532 1928 5536
rect 1940 5532 1941 5536
rect 1943 5532 1944 5536
rect 1961 5532 1962 5536
rect 1964 5532 1966 5536
rect 1987 5532 1988 5536
rect 1990 5532 1993 5536
rect 1995 5532 2000 5536
rect 2015 5532 2016 5536
rect 2018 5532 2019 5536
rect 2031 5532 2032 5536
rect 2034 5532 2035 5536
rect 2056 5532 2057 5536
rect 2059 5532 2060 5536
rect 2064 5532 2070 5536
rect 2074 5532 2075 5536
rect 2077 5532 2078 5536
rect 2158 5532 2159 5536
rect 2161 5532 2162 5536
rect 2176 5532 2177 5536
rect 2179 5532 2182 5536
rect 2184 5532 2189 5536
rect 2201 5532 2202 5536
rect 2204 5532 2205 5536
rect 2222 5532 2223 5536
rect 2225 5532 2227 5536
rect 2248 5532 2249 5536
rect 2251 5532 2254 5536
rect 2256 5532 2261 5536
rect 2276 5532 2277 5536
rect 2279 5532 2280 5536
rect 2292 5532 2293 5536
rect 2295 5532 2296 5536
rect 2308 5532 2309 5536
rect 2311 5532 2312 5536
rect 1213 5486 1214 5490
rect 1216 5486 1217 5490
rect 1231 5486 1232 5490
rect 1234 5486 1237 5490
rect 1239 5486 1244 5490
rect 1256 5486 1257 5490
rect 1259 5486 1260 5490
rect 1277 5486 1278 5490
rect 1280 5486 1282 5490
rect 1303 5486 1304 5490
rect 1306 5486 1309 5490
rect 1311 5486 1316 5490
rect 1331 5486 1332 5490
rect 1334 5486 1335 5490
rect 1347 5486 1348 5490
rect 1350 5486 1351 5490
rect 1363 5486 1364 5490
rect 1366 5486 1367 5490
rect 1135 5481 1136 5485
rect 1138 5481 1139 5485
rect 1158 5477 1159 5481
rect 1161 5477 1164 5481
rect 1166 5477 1169 5481
rect 2158 5486 2159 5490
rect 2161 5486 2162 5490
rect 2176 5486 2177 5490
rect 2179 5486 2182 5490
rect 2184 5486 2189 5490
rect 2201 5486 2202 5490
rect 2204 5486 2205 5490
rect 2222 5486 2223 5490
rect 2225 5486 2227 5490
rect 2248 5486 2249 5490
rect 2251 5486 2254 5490
rect 2256 5486 2261 5490
rect 2276 5486 2277 5490
rect 2279 5486 2280 5490
rect 2292 5486 2293 5490
rect 2295 5486 2296 5490
rect 2308 5486 2309 5490
rect 2311 5486 2312 5490
rect 2080 5481 2081 5485
rect 2083 5481 2084 5485
rect 2103 5477 2104 5481
rect 2106 5477 2109 5481
rect 2111 5477 2114 5481
rect 1767 5432 1768 5436
rect 1770 5432 1773 5436
rect 1775 5432 1778 5436
rect 987 5403 988 5407
rect 990 5403 993 5407
rect 995 5403 998 5407
rect 1077 5403 1078 5407
rect 1080 5403 1083 5407
rect 1085 5403 1088 5407
rect 1158 5403 1159 5407
rect 1161 5403 1164 5407
rect 1166 5403 1169 5407
rect 1213 5400 1214 5404
rect 1216 5400 1217 5404
rect 1231 5400 1232 5404
rect 1234 5400 1237 5404
rect 1239 5400 1244 5404
rect 1256 5400 1257 5404
rect 1259 5400 1260 5404
rect 1277 5400 1278 5404
rect 1280 5400 1282 5404
rect 1303 5400 1304 5404
rect 1306 5400 1309 5404
rect 1311 5400 1316 5404
rect 1331 5400 1332 5404
rect 1334 5400 1335 5404
rect 1347 5400 1348 5404
rect 1350 5400 1351 5404
rect 1363 5400 1364 5404
rect 1366 5400 1367 5404
rect 1653 5399 1654 5411
rect 1656 5399 1657 5411
rect 1706 5399 1707 5411
rect 1709 5399 1710 5411
rect 1932 5403 1933 5407
rect 1935 5403 1938 5407
rect 1940 5403 1943 5407
rect 2022 5403 2023 5407
rect 2025 5403 2028 5407
rect 2030 5403 2033 5407
rect 2103 5403 2104 5407
rect 2106 5403 2109 5407
rect 2111 5403 2114 5407
rect 2158 5400 2159 5404
rect 2161 5400 2162 5404
rect 2176 5400 2177 5404
rect 2179 5400 2182 5404
rect 2184 5400 2189 5404
rect 2201 5400 2202 5404
rect 2204 5400 2205 5404
rect 2222 5400 2223 5404
rect 2225 5400 2227 5404
rect 2248 5400 2249 5404
rect 2251 5400 2254 5404
rect 2256 5400 2261 5404
rect 2276 5400 2277 5404
rect 2279 5400 2280 5404
rect 2292 5400 2293 5404
rect 2295 5400 2296 5404
rect 2308 5400 2309 5404
rect 2311 5400 2312 5404
rect 964 5349 965 5353
rect 967 5349 968 5353
rect 1054 5349 1055 5353
rect 1057 5349 1058 5353
rect 1213 5354 1214 5358
rect 1216 5354 1217 5358
rect 1231 5354 1232 5358
rect 1234 5354 1237 5358
rect 1239 5354 1244 5358
rect 1256 5354 1257 5358
rect 1259 5354 1260 5358
rect 1277 5354 1278 5358
rect 1280 5354 1282 5358
rect 1303 5354 1304 5358
rect 1306 5354 1309 5358
rect 1311 5354 1316 5358
rect 1331 5354 1332 5358
rect 1334 5354 1335 5358
rect 1347 5354 1348 5358
rect 1350 5354 1351 5358
rect 1363 5354 1364 5358
rect 1366 5354 1367 5358
rect 1135 5349 1136 5353
rect 1138 5349 1139 5353
rect 987 5345 988 5349
rect 990 5345 993 5349
rect 995 5345 998 5349
rect 1018 5341 1019 5345
rect 1021 5341 1022 5345
rect 1077 5345 1078 5349
rect 1080 5345 1083 5349
rect 1085 5345 1088 5349
rect 1108 5341 1109 5345
rect 1111 5341 1112 5345
rect 1158 5345 1159 5349
rect 1161 5345 1164 5349
rect 1166 5345 1169 5349
rect 1744 5376 1745 5380
rect 1747 5376 1748 5380
rect 1767 5372 1768 5376
rect 1770 5372 1773 5376
rect 1775 5372 1778 5376
rect 1798 5368 1799 5372
rect 1801 5368 1802 5372
rect 1820 5368 1821 5372
rect 1823 5368 1824 5372
rect 1909 5349 1910 5353
rect 1912 5349 1913 5353
rect 1999 5349 2000 5353
rect 2002 5349 2003 5353
rect 2158 5354 2159 5358
rect 2161 5354 2162 5358
rect 2176 5354 2177 5358
rect 2179 5354 2182 5358
rect 2184 5354 2189 5358
rect 2201 5354 2202 5358
rect 2204 5354 2205 5358
rect 2222 5354 2223 5358
rect 2225 5354 2227 5358
rect 2248 5354 2249 5358
rect 2251 5354 2254 5358
rect 2256 5354 2261 5358
rect 2276 5354 2277 5358
rect 2279 5354 2280 5358
rect 2292 5354 2293 5358
rect 2295 5354 2296 5358
rect 2308 5354 2309 5358
rect 2311 5354 2312 5358
rect 2080 5349 2081 5353
rect 2083 5349 2084 5353
rect 1932 5345 1933 5349
rect 1935 5345 1938 5349
rect 1940 5345 1943 5349
rect 1963 5341 1964 5345
rect 1966 5341 1967 5345
rect 2022 5345 2023 5349
rect 2025 5345 2028 5349
rect 2030 5345 2033 5349
rect 2053 5341 2054 5345
rect 2056 5341 2057 5345
rect 2103 5345 2104 5349
rect 2106 5345 2109 5349
rect 2111 5345 2114 5349
rect 1767 5302 1768 5306
rect 1770 5302 1773 5306
rect 1775 5302 1778 5306
rect 1053 5268 1054 5272
rect 1056 5268 1059 5272
rect 1061 5268 1064 5272
rect 1158 5268 1159 5272
rect 1161 5268 1164 5272
rect 1166 5268 1169 5272
rect 1213 5268 1214 5272
rect 1216 5268 1217 5272
rect 1231 5268 1232 5272
rect 1234 5268 1237 5272
rect 1239 5268 1244 5272
rect 1256 5268 1257 5272
rect 1259 5268 1260 5272
rect 1277 5268 1278 5272
rect 1280 5268 1282 5272
rect 1303 5268 1304 5272
rect 1306 5268 1309 5272
rect 1311 5268 1316 5272
rect 1331 5268 1332 5272
rect 1334 5268 1335 5272
rect 1347 5268 1348 5272
rect 1350 5268 1351 5272
rect 1363 5268 1364 5272
rect 1366 5268 1367 5272
rect 1559 5269 1560 5281
rect 1562 5269 1563 5281
rect 1612 5269 1613 5281
rect 1615 5269 1616 5281
rect 1998 5268 1999 5272
rect 2001 5268 2004 5272
rect 2006 5268 2009 5272
rect 2103 5268 2104 5272
rect 2106 5268 2109 5272
rect 2111 5268 2114 5272
rect 2158 5268 2159 5272
rect 2161 5268 2162 5272
rect 2176 5268 2177 5272
rect 2179 5268 2182 5272
rect 2184 5268 2189 5272
rect 2201 5268 2202 5272
rect 2204 5268 2205 5272
rect 2222 5268 2223 5272
rect 2225 5268 2227 5272
rect 2248 5268 2249 5272
rect 2251 5268 2254 5272
rect 2256 5268 2261 5272
rect 2276 5268 2277 5272
rect 2279 5268 2280 5272
rect 2292 5268 2293 5272
rect 2295 5268 2296 5272
rect 2308 5268 2309 5272
rect 2311 5268 2312 5272
rect 1030 5217 1031 5221
rect 1033 5217 1034 5221
rect 1213 5222 1214 5226
rect 1216 5222 1217 5226
rect 1231 5222 1232 5226
rect 1234 5222 1237 5226
rect 1239 5222 1244 5226
rect 1256 5222 1257 5226
rect 1259 5222 1260 5226
rect 1277 5222 1278 5226
rect 1280 5222 1282 5226
rect 1303 5222 1304 5226
rect 1306 5222 1309 5226
rect 1311 5222 1316 5226
rect 1331 5222 1332 5226
rect 1334 5222 1335 5226
rect 1347 5222 1348 5226
rect 1350 5222 1351 5226
rect 1363 5222 1364 5226
rect 1366 5222 1367 5226
rect 1135 5217 1136 5221
rect 1138 5217 1139 5221
rect 1053 5213 1054 5217
rect 1056 5213 1059 5217
rect 1061 5213 1064 5217
rect 1084 5209 1085 5213
rect 1087 5209 1088 5213
rect 1158 5213 1159 5217
rect 1161 5213 1164 5217
rect 1166 5213 1169 5217
rect 1744 5246 1745 5250
rect 1747 5246 1748 5250
rect 1767 5242 1768 5246
rect 1770 5242 1773 5246
rect 1775 5242 1778 5246
rect 1798 5238 1799 5242
rect 1801 5238 1802 5242
rect 1975 5217 1976 5221
rect 1978 5217 1979 5221
rect 2158 5222 2159 5226
rect 2161 5222 2162 5226
rect 2176 5222 2177 5226
rect 2179 5222 2182 5226
rect 2184 5222 2189 5226
rect 2201 5222 2202 5226
rect 2204 5222 2205 5226
rect 2222 5222 2223 5226
rect 2225 5222 2227 5226
rect 2248 5222 2249 5226
rect 2251 5222 2254 5226
rect 2256 5222 2261 5226
rect 2276 5222 2277 5226
rect 2279 5222 2280 5226
rect 2292 5222 2293 5226
rect 2295 5222 2296 5226
rect 2308 5222 2309 5226
rect 2311 5222 2312 5226
rect 2080 5217 2081 5221
rect 2083 5217 2084 5221
rect 1998 5213 1999 5217
rect 2001 5213 2004 5217
rect 2006 5213 2009 5217
rect 2029 5209 2030 5213
rect 2032 5209 2033 5213
rect 2103 5213 2104 5217
rect 2106 5213 2109 5217
rect 2111 5213 2114 5217
rect 1077 5137 1078 5141
rect 1080 5137 1083 5141
rect 1085 5137 1088 5141
rect 1158 5137 1159 5141
rect 1161 5137 1164 5141
rect 1166 5137 1169 5141
rect 1613 5146 1614 5150
rect 1616 5146 1619 5150
rect 1621 5146 1622 5150
rect 1634 5146 1635 5150
rect 1637 5146 1638 5150
rect 1650 5146 1651 5150
rect 1653 5146 1656 5150
rect 1658 5146 1659 5150
rect 1676 5146 1677 5150
rect 1679 5146 1680 5150
rect 1692 5146 1693 5150
rect 1695 5146 1696 5150
rect 1708 5146 1709 5150
rect 1711 5146 1714 5150
rect 1716 5146 1717 5150
rect 1729 5146 1730 5150
rect 1732 5146 1733 5150
rect 1213 5136 1214 5140
rect 1216 5136 1217 5140
rect 1231 5136 1232 5140
rect 1234 5136 1237 5140
rect 1239 5136 1244 5140
rect 1256 5136 1257 5140
rect 1259 5136 1260 5140
rect 1277 5136 1278 5140
rect 1280 5136 1282 5140
rect 1303 5136 1304 5140
rect 1306 5136 1309 5140
rect 1311 5136 1316 5140
rect 1331 5136 1332 5140
rect 1334 5136 1335 5140
rect 1347 5136 1348 5140
rect 1350 5136 1351 5140
rect 1363 5136 1364 5140
rect 1366 5136 1367 5140
rect 2022 5137 2023 5141
rect 2025 5137 2028 5141
rect 2030 5137 2033 5141
rect 2103 5137 2104 5141
rect 2106 5137 2109 5141
rect 2111 5137 2114 5141
rect 2558 5146 2559 5150
rect 2561 5146 2564 5150
rect 2566 5146 2567 5150
rect 2579 5146 2580 5150
rect 2582 5146 2583 5150
rect 2595 5146 2596 5150
rect 2598 5146 2601 5150
rect 2603 5146 2604 5150
rect 2621 5146 2622 5150
rect 2624 5146 2625 5150
rect 2637 5146 2638 5150
rect 2640 5146 2641 5150
rect 2653 5146 2654 5150
rect 2656 5146 2659 5150
rect 2661 5146 2662 5150
rect 2674 5146 2675 5150
rect 2677 5146 2678 5150
rect 2158 5136 2159 5140
rect 2161 5136 2162 5140
rect 2176 5136 2177 5140
rect 2179 5136 2182 5140
rect 2184 5136 2189 5140
rect 2201 5136 2202 5140
rect 2204 5136 2205 5140
rect 2222 5136 2223 5140
rect 2225 5136 2227 5140
rect 2248 5136 2249 5140
rect 2251 5136 2254 5140
rect 2256 5136 2261 5140
rect 2276 5136 2277 5140
rect 2279 5136 2280 5140
rect 2292 5136 2293 5140
rect 2295 5136 2296 5140
rect 2308 5136 2309 5140
rect 2311 5136 2312 5140
rect 1054 5085 1055 5089
rect 1057 5085 1058 5089
rect 1213 5090 1214 5094
rect 1216 5090 1217 5094
rect 1231 5090 1232 5094
rect 1234 5090 1237 5094
rect 1239 5090 1244 5094
rect 1256 5090 1257 5094
rect 1259 5090 1260 5094
rect 1277 5090 1278 5094
rect 1280 5090 1282 5094
rect 1303 5090 1304 5094
rect 1306 5090 1309 5094
rect 1311 5090 1316 5094
rect 1331 5090 1332 5094
rect 1334 5090 1335 5094
rect 1347 5090 1348 5094
rect 1350 5090 1351 5094
rect 1363 5090 1364 5094
rect 1366 5090 1367 5094
rect 1713 5090 1714 5094
rect 1716 5090 1717 5094
rect 1135 5085 1136 5089
rect 1138 5085 1139 5089
rect 1077 5081 1078 5085
rect 1080 5081 1083 5085
rect 1085 5081 1088 5085
rect 1108 5077 1109 5081
rect 1111 5077 1112 5081
rect 1158 5081 1159 5085
rect 1161 5081 1164 5085
rect 1166 5081 1169 5085
rect 1189 5077 1190 5081
rect 1192 5077 1193 5081
rect 1596 5081 1597 5085
rect 1599 5081 1600 5085
rect 1999 5085 2000 5089
rect 2002 5085 2003 5089
rect 2158 5090 2159 5094
rect 2161 5090 2162 5094
rect 2176 5090 2177 5094
rect 2179 5090 2182 5094
rect 2184 5090 2189 5094
rect 2201 5090 2202 5094
rect 2204 5090 2205 5094
rect 2222 5090 2223 5094
rect 2225 5090 2227 5094
rect 2248 5090 2249 5094
rect 2251 5090 2254 5094
rect 2256 5090 2261 5094
rect 2276 5090 2277 5094
rect 2279 5090 2280 5094
rect 2292 5090 2293 5094
rect 2295 5090 2296 5094
rect 2308 5090 2309 5094
rect 2311 5090 2312 5094
rect 2658 5090 2659 5094
rect 2661 5090 2662 5094
rect 2080 5085 2081 5089
rect 2083 5085 2084 5089
rect 2022 5081 2023 5085
rect 2025 5081 2028 5085
rect 2030 5081 2033 5085
rect 2053 5077 2054 5081
rect 2056 5077 2057 5081
rect 2103 5081 2104 5085
rect 2106 5081 2109 5085
rect 2111 5081 2114 5085
rect 2134 5077 2135 5081
rect 2137 5077 2138 5081
rect 2541 5081 2542 5085
rect 2544 5081 2545 5085
rect 1604 5044 1605 5048
rect 1607 5044 1608 5048
rect 1620 5044 1621 5048
rect 1623 5044 1626 5048
rect 1628 5044 1629 5048
rect 1641 5044 1642 5048
rect 1644 5044 1645 5048
rect 1657 5044 1658 5048
rect 1660 5044 1661 5048
rect 1678 5044 1679 5048
rect 1681 5044 1684 5048
rect 1686 5044 1687 5048
rect 1699 5044 1700 5048
rect 1702 5044 1703 5048
rect 1715 5044 1716 5048
rect 1718 5044 1721 5048
rect 1723 5044 1724 5048
rect 2549 5044 2550 5048
rect 2552 5044 2553 5048
rect 2565 5044 2566 5048
rect 2568 5044 2571 5048
rect 2573 5044 2574 5048
rect 2586 5044 2587 5048
rect 2589 5044 2590 5048
rect 2602 5044 2603 5048
rect 2605 5044 2606 5048
rect 2623 5044 2624 5048
rect 2626 5044 2629 5048
rect 2631 5044 2632 5048
rect 2644 5044 2645 5048
rect 2647 5044 2648 5048
rect 2660 5044 2661 5048
rect 2663 5044 2666 5048
rect 2668 5044 2669 5048
rect 856 5011 857 5015
rect 859 5011 860 5015
rect 872 5011 873 5015
rect 875 5011 878 5015
rect 880 5011 881 5015
rect 893 5011 894 5015
rect 896 5011 897 5015
rect 909 5011 910 5015
rect 912 5011 913 5015
rect 930 5011 931 5015
rect 933 5011 936 5015
rect 938 5011 939 5015
rect 951 5011 952 5015
rect 954 5011 955 5015
rect 967 5011 968 5015
rect 970 5011 973 5015
rect 975 5011 976 5015
rect 988 5011 989 5015
rect 991 5011 992 5015
rect 1004 5011 1005 5015
rect 1007 5011 1010 5015
rect 1012 5011 1013 5015
rect 1025 5011 1026 5015
rect 1028 5011 1029 5015
rect 1041 5011 1042 5015
rect 1044 5011 1045 5015
rect 1062 5011 1063 5015
rect 1065 5011 1068 5015
rect 1070 5011 1071 5015
rect 1083 5011 1084 5015
rect 1086 5011 1087 5015
rect 1099 5011 1100 5015
rect 1102 5011 1105 5015
rect 1107 5011 1108 5015
rect 1120 5011 1121 5015
rect 1123 5011 1124 5015
rect 1136 5011 1137 5015
rect 1139 5011 1142 5015
rect 1144 5011 1145 5015
rect 1157 5011 1158 5015
rect 1160 5011 1161 5015
rect 1173 5011 1174 5015
rect 1176 5011 1177 5015
rect 1194 5011 1195 5015
rect 1197 5011 1200 5015
rect 1202 5011 1203 5015
rect 1215 5011 1216 5015
rect 1218 5011 1219 5015
rect 1231 5011 1232 5015
rect 1234 5011 1237 5015
rect 1239 5011 1240 5015
rect 1252 5011 1253 5015
rect 1255 5011 1256 5015
rect 1268 5011 1269 5015
rect 1271 5011 1274 5015
rect 1276 5011 1277 5015
rect 1289 5011 1290 5015
rect 1292 5011 1293 5015
rect 1305 5011 1306 5015
rect 1308 5011 1309 5015
rect 1326 5011 1327 5015
rect 1329 5011 1332 5015
rect 1334 5011 1335 5015
rect 1347 5011 1348 5015
rect 1350 5011 1351 5015
rect 1363 5011 1364 5015
rect 1366 5011 1369 5015
rect 1371 5011 1372 5015
rect 1801 5011 1802 5015
rect 1804 5011 1805 5015
rect 1817 5011 1818 5015
rect 1820 5011 1823 5015
rect 1825 5011 1826 5015
rect 1838 5011 1839 5015
rect 1841 5011 1842 5015
rect 1854 5011 1855 5015
rect 1857 5011 1858 5015
rect 1875 5011 1876 5015
rect 1878 5011 1881 5015
rect 1883 5011 1884 5015
rect 1896 5011 1897 5015
rect 1899 5011 1900 5015
rect 1912 5011 1913 5015
rect 1915 5011 1918 5015
rect 1920 5011 1921 5015
rect 1933 5011 1934 5015
rect 1936 5011 1937 5015
rect 1949 5011 1950 5015
rect 1952 5011 1955 5015
rect 1957 5011 1958 5015
rect 1970 5011 1971 5015
rect 1973 5011 1974 5015
rect 1986 5011 1987 5015
rect 1989 5011 1990 5015
rect 2007 5011 2008 5015
rect 2010 5011 2013 5015
rect 2015 5011 2016 5015
rect 2028 5011 2029 5015
rect 2031 5011 2032 5015
rect 2044 5011 2045 5015
rect 2047 5011 2050 5015
rect 2052 5011 2053 5015
rect 2065 5011 2066 5015
rect 2068 5011 2069 5015
rect 2081 5011 2082 5015
rect 2084 5011 2087 5015
rect 2089 5011 2090 5015
rect 2102 5011 2103 5015
rect 2105 5011 2106 5015
rect 2118 5011 2119 5015
rect 2121 5011 2122 5015
rect 2139 5011 2140 5015
rect 2142 5011 2145 5015
rect 2147 5011 2148 5015
rect 2160 5011 2161 5015
rect 2163 5011 2164 5015
rect 2176 5011 2177 5015
rect 2179 5011 2182 5015
rect 2184 5011 2185 5015
rect 2197 5011 2198 5015
rect 2200 5011 2201 5015
rect 2213 5011 2214 5015
rect 2216 5011 2219 5015
rect 2221 5011 2222 5015
rect 2234 5011 2235 5015
rect 2237 5011 2238 5015
rect 2250 5011 2251 5015
rect 2253 5011 2254 5015
rect 2271 5011 2272 5015
rect 2274 5011 2277 5015
rect 2279 5011 2280 5015
rect 2292 5011 2293 5015
rect 2295 5011 2296 5015
rect 2308 5011 2309 5015
rect 2311 5011 2314 5015
rect 2316 5011 2317 5015
rect 4578 7986 4579 8015
rect 4574 7982 4579 7986
rect 4578 7975 4579 7982
rect 4581 7975 4582 8015
rect 4586 7975 4587 8015
rect 4589 7986 4590 8015
rect 4594 7986 4595 8015
rect 4589 7982 4595 7986
rect 4589 7975 4590 7982
rect 4594 7975 4595 7982
rect 4597 7975 4598 8015
rect 4602 7975 4603 8015
rect 4605 7986 4606 8015
rect 4610 7986 4611 8015
rect 4605 7982 4611 7986
rect 4605 7975 4606 7982
rect 4610 7975 4611 7982
rect 4613 7975 4614 8015
rect 4618 7975 4619 8015
rect 4621 7986 4622 8015
rect 4626 7986 4627 8015
rect 4621 7982 4627 7986
rect 4621 7975 4622 7982
rect 4626 7975 4627 7982
rect 4631 7975 4634 8034
rect 4636 7975 4637 8034
rect 4641 7975 4642 8034
rect 4644 7986 4645 8034
rect 4649 7986 4650 8034
rect 4644 7982 4650 7986
rect 4644 7975 4645 7982
rect 4649 7975 4650 7982
rect 4652 7975 4653 8034
rect 4657 7975 4658 8034
rect 4660 7986 4661 8034
rect 4665 7986 4666 8034
rect 4660 7982 4666 7986
rect 4660 7975 4661 7982
rect 4665 7975 4666 7982
rect 4670 7975 4677 8034
rect 4679 7975 4680 8034
rect 4684 7975 4685 8034
rect 4687 7986 4688 8034
rect 4692 7986 4693 8034
rect 4687 7975 4693 7986
rect 4695 7975 4696 8034
rect 4700 7975 4701 8034
rect 4703 7986 4704 8034
rect 4708 7986 4709 8034
rect 4703 7982 4709 7986
rect 4703 7975 4704 7982
rect 4708 7975 4709 7982
rect 4713 7975 4718 8034
rect 4720 7975 4721 8034
rect 4725 7975 4726 8034
rect 4728 7986 4729 8034
rect 4733 7986 4734 8034
rect 4728 7975 4734 7986
rect 4736 7975 4737 8034
rect 4741 7975 4742 8034
rect 4744 7986 4745 8034
rect 4749 7986 4750 8034
rect 4744 7982 4750 7986
rect 4744 7975 4745 7982
rect 4749 7975 4750 7982
rect 4661 7461 4667 7465
rect 4671 7461 4677 7465
rect 4681 7461 4687 7465
rect 4691 7461 4697 7465
rect 4701 7461 4707 7465
rect 4711 7461 4717 7465
rect 4721 7461 4727 7465
rect 4731 7461 4737 7465
rect 4741 7461 4746 7465
rect 4657 7460 4746 7461
rect 4657 7456 4662 7460
rect 4666 7456 4672 7460
rect 4676 7456 4682 7460
rect 4686 7456 4692 7460
rect 4696 7456 4702 7460
rect 4706 7456 4712 7460
rect 4716 7456 4722 7460
rect 4726 7456 4732 7460
rect 4736 7456 4742 7460
rect 4657 7455 4746 7456
rect 4661 7451 4667 7455
rect 4671 7451 4677 7455
rect 4681 7451 4687 7455
rect 4691 7451 4697 7455
rect 4701 7451 4707 7455
rect 4711 7451 4717 7455
rect 4721 7451 4727 7455
rect 4731 7451 4737 7455
rect 4741 7451 4746 7455
rect 4657 7450 4746 7451
rect 4657 7446 4662 7450
rect 4666 7446 4672 7450
rect 4676 7446 4682 7450
rect 4686 7446 4692 7450
rect 4696 7446 4702 7450
rect 4706 7446 4712 7450
rect 4716 7446 4722 7450
rect 4726 7446 4732 7450
rect 4736 7446 4742 7450
rect 4657 7445 4746 7446
rect 4661 7441 4667 7445
rect 4671 7441 4677 7445
rect 4681 7441 4687 7445
rect 4691 7441 4697 7445
rect 4701 7441 4707 7445
rect 4711 7441 4717 7445
rect 4721 7441 4727 7445
rect 4731 7441 4737 7445
rect 4741 7441 4746 7445
rect 4657 7440 4746 7441
rect 4657 7436 4662 7440
rect 4666 7436 4672 7440
rect 4676 7436 4682 7440
rect 4686 7436 4692 7440
rect 4696 7436 4702 7440
rect 4706 7436 4712 7440
rect 4716 7436 4722 7440
rect 4726 7436 4732 7440
rect 4736 7436 4742 7440
rect 4657 7435 4746 7436
rect 4661 7431 4667 7435
rect 4671 7431 4677 7435
rect 4681 7431 4687 7435
rect 4691 7431 4697 7435
rect 4701 7431 4707 7435
rect 4711 7431 4717 7435
rect 4721 7431 4727 7435
rect 4731 7431 4737 7435
rect 4741 7431 4746 7435
rect 4657 7430 4746 7431
rect 4657 7426 4662 7430
rect 4666 7426 4672 7430
rect 4676 7426 4682 7430
rect 4686 7426 4692 7430
rect 4696 7426 4702 7430
rect 4706 7426 4712 7430
rect 4716 7426 4722 7430
rect 4726 7426 4732 7430
rect 4736 7426 4742 7430
rect 4657 7425 4746 7426
rect 4661 7421 4667 7425
rect 4671 7421 4677 7425
rect 4681 7421 4687 7425
rect 4691 7421 4697 7425
rect 4701 7421 4707 7425
rect 4711 7421 4717 7425
rect 4721 7421 4727 7425
rect 4731 7421 4737 7425
rect 4741 7421 4746 7425
rect 4576 7335 4577 7342
rect 4572 7331 4577 7335
rect 4576 7302 4577 7331
rect 4579 7302 4580 7342
rect 4584 7302 4585 7342
rect 4587 7335 4588 7342
rect 4592 7335 4593 7342
rect 4587 7331 4593 7335
rect 4587 7302 4588 7331
rect 4592 7302 4593 7331
rect 4595 7302 4596 7342
rect 4600 7302 4601 7342
rect 4603 7335 4604 7342
rect 4608 7335 4609 7342
rect 4603 7331 4609 7335
rect 4603 7302 4604 7331
rect 4608 7302 4609 7331
rect 4611 7302 4612 7342
rect 4616 7302 4617 7342
rect 4619 7335 4620 7342
rect 4619 7331 4624 7335
rect 4619 7302 4620 7331
rect 1169 4531 1173 4535
rect 1140 4530 1180 4531
rect 2096 4531 2100 4535
rect 2067 4530 2107 4531
rect 2405 4531 2409 4535
rect 2376 4530 2416 4531
rect 2714 4531 2718 4535
rect 2685 4530 2725 4531
rect 3023 4531 3027 4535
rect 2994 4530 3034 4531
rect 3332 4531 3336 4535
rect 3303 4530 3343 4531
rect 1140 4527 1180 4528
rect 1140 4522 1180 4523
rect 1140 4519 1180 4520
rect 1169 4515 1173 4519
rect 1140 4514 1180 4515
rect 1140 4511 1180 4512
rect 1140 4506 1180 4507
rect 1140 4503 1180 4504
rect 1169 4499 1173 4503
rect 2067 4527 2107 4528
rect 2067 4522 2107 4523
rect 2067 4519 2107 4520
rect 2096 4515 2100 4519
rect 2067 4514 2107 4515
rect 2067 4511 2107 4512
rect 2067 4506 2107 4507
rect 1140 4498 1180 4499
rect 2067 4503 2107 4504
rect 2096 4499 2100 4503
rect 2376 4527 2416 4528
rect 2376 4522 2416 4523
rect 2376 4519 2416 4520
rect 2405 4515 2409 4519
rect 2376 4514 2416 4515
rect 2376 4511 2416 4512
rect 2376 4506 2416 4507
rect 2067 4498 2107 4499
rect 2376 4503 2416 4504
rect 2405 4499 2409 4503
rect 2685 4527 2725 4528
rect 2685 4522 2725 4523
rect 2685 4519 2725 4520
rect 2714 4515 2718 4519
rect 2685 4514 2725 4515
rect 2685 4511 2725 4512
rect 2685 4506 2725 4507
rect 2376 4498 2416 4499
rect 2685 4503 2725 4504
rect 2714 4499 2718 4503
rect 2994 4527 3034 4528
rect 2994 4522 3034 4523
rect 2994 4519 3034 4520
rect 3023 4515 3027 4519
rect 2994 4514 3034 4515
rect 2994 4511 3034 4512
rect 2994 4506 3034 4507
rect 2685 4498 2725 4499
rect 2994 4503 3034 4504
rect 3023 4499 3027 4503
rect 3303 4527 3343 4528
rect 3303 4522 3343 4523
rect 3303 4519 3343 4520
rect 3332 4515 3336 4519
rect 3303 4514 3343 4515
rect 3303 4511 3343 4512
rect 3303 4506 3343 4507
rect 2994 4498 3034 4499
rect 3303 4503 3343 4504
rect 3332 4499 3336 4503
rect 3303 4498 3343 4499
rect 1140 4495 1180 4496
rect 1140 4490 1180 4491
rect 2067 4495 2107 4496
rect 2067 4490 2107 4491
rect 2376 4495 2416 4496
rect 2376 4490 2416 4491
rect 2685 4495 2725 4496
rect 2685 4490 2725 4491
rect 2994 4495 3034 4496
rect 2994 4490 3034 4491
rect 3303 4495 3343 4496
rect 3303 4490 3343 4491
rect 1140 4487 1180 4488
rect 1169 4483 1173 4487
rect 2067 4487 2107 4488
rect 2096 4483 2100 4487
rect 2376 4487 2416 4488
rect 2405 4483 2409 4487
rect 2685 4487 2725 4488
rect 2714 4483 2718 4487
rect 2994 4487 3034 4488
rect 3023 4483 3027 4487
rect 3303 4487 3343 4488
rect 3332 4483 3336 4487
rect 1263 4446 1269 4450
rect 1273 4446 1279 4450
rect 1283 4446 1289 4450
rect 1293 4446 1299 4450
rect 1259 4445 1303 4446
rect 1259 4441 1264 4445
rect 1268 4441 1274 4445
rect 1278 4441 1284 4445
rect 1288 4441 1294 4445
rect 1298 4441 1303 4445
rect 1259 4440 1303 4441
rect 1263 4436 1269 4440
rect 1273 4436 1279 4440
rect 1283 4436 1289 4440
rect 1293 4436 1299 4440
rect 1259 4435 1303 4436
rect 1259 4431 1264 4435
rect 1268 4431 1274 4435
rect 1278 4431 1284 4435
rect 1288 4431 1294 4435
rect 1298 4431 1303 4435
rect 1259 4430 1303 4431
rect 1263 4426 1269 4430
rect 1273 4426 1279 4430
rect 1283 4426 1289 4430
rect 1293 4426 1299 4430
rect 1259 4425 1303 4426
rect 1259 4421 1264 4425
rect 1268 4421 1274 4425
rect 1278 4421 1284 4425
rect 1288 4421 1294 4425
rect 1298 4421 1303 4425
rect 1259 4420 1303 4421
rect 1263 4416 1269 4420
rect 1273 4416 1279 4420
rect 1283 4416 1289 4420
rect 1293 4416 1299 4420
rect 1259 4415 1303 4416
rect 1259 4411 1264 4415
rect 1268 4411 1274 4415
rect 1278 4411 1284 4415
rect 1288 4411 1294 4415
rect 1298 4411 1303 4415
rect 1259 4410 1303 4411
rect 1263 4406 1269 4410
rect 1273 4406 1279 4410
rect 1283 4406 1289 4410
rect 1293 4406 1299 4410
rect 1259 4405 1303 4406
rect 1259 4401 1264 4405
rect 1268 4401 1274 4405
rect 1278 4401 1284 4405
rect 1288 4401 1294 4405
rect 1298 4401 1303 4405
rect 1259 4400 1303 4401
rect 1263 4396 1269 4400
rect 1273 4396 1279 4400
rect 1283 4396 1289 4400
rect 1293 4396 1299 4400
rect 1259 4395 1303 4396
rect 1259 4391 1264 4395
rect 1268 4391 1274 4395
rect 1278 4391 1284 4395
rect 1288 4391 1294 4395
rect 1298 4391 1303 4395
rect 1259 4390 1303 4391
rect 1263 4386 1269 4390
rect 1273 4386 1279 4390
rect 1283 4386 1289 4390
rect 1293 4386 1299 4390
rect 1259 4385 1303 4386
rect 1259 4381 1264 4385
rect 1268 4381 1274 4385
rect 1278 4381 1284 4385
rect 1288 4381 1294 4385
rect 1298 4381 1303 4385
rect 1259 4380 1303 4381
rect 1263 4376 1269 4380
rect 1273 4376 1279 4380
rect 1283 4376 1289 4380
rect 1293 4376 1299 4380
rect 1259 4375 1303 4376
rect 1259 4371 1264 4375
rect 1268 4371 1274 4375
rect 1278 4371 1284 4375
rect 1288 4371 1294 4375
rect 1298 4371 1303 4375
rect 1259 4370 1303 4371
rect 1263 4366 1269 4370
rect 1273 4366 1279 4370
rect 1283 4366 1289 4370
rect 1293 4366 1299 4370
rect 1259 4365 1303 4366
rect 1259 4361 1264 4365
rect 1268 4361 1274 4365
rect 1278 4361 1284 4365
rect 1288 4361 1294 4365
rect 1298 4361 1303 4365
rect 1572 4446 1578 4450
rect 1582 4446 1588 4450
rect 1592 4446 1598 4450
rect 1602 4446 1608 4450
rect 1568 4445 1612 4446
rect 1568 4441 1573 4445
rect 1577 4441 1583 4445
rect 1587 4441 1593 4445
rect 1597 4441 1603 4445
rect 1607 4441 1612 4445
rect 1568 4440 1612 4441
rect 1572 4436 1578 4440
rect 1582 4436 1588 4440
rect 1592 4436 1598 4440
rect 1602 4436 1608 4440
rect 1568 4435 1612 4436
rect 1568 4431 1573 4435
rect 1577 4431 1583 4435
rect 1587 4431 1593 4435
rect 1597 4431 1603 4435
rect 1607 4431 1612 4435
rect 1568 4430 1612 4431
rect 1572 4426 1578 4430
rect 1582 4426 1588 4430
rect 1592 4426 1598 4430
rect 1602 4426 1608 4430
rect 1568 4425 1612 4426
rect 1568 4421 1573 4425
rect 1577 4421 1583 4425
rect 1587 4421 1593 4425
rect 1597 4421 1603 4425
rect 1607 4421 1612 4425
rect 1568 4420 1612 4421
rect 1572 4416 1578 4420
rect 1582 4416 1588 4420
rect 1592 4416 1598 4420
rect 1602 4416 1608 4420
rect 1568 4415 1612 4416
rect 1568 4411 1573 4415
rect 1577 4411 1583 4415
rect 1587 4411 1593 4415
rect 1597 4411 1603 4415
rect 1607 4411 1612 4415
rect 1568 4410 1612 4411
rect 1572 4406 1578 4410
rect 1582 4406 1588 4410
rect 1592 4406 1598 4410
rect 1602 4406 1608 4410
rect 1568 4405 1612 4406
rect 1568 4401 1573 4405
rect 1577 4401 1583 4405
rect 1587 4401 1593 4405
rect 1597 4401 1603 4405
rect 1607 4401 1612 4405
rect 1568 4400 1612 4401
rect 1572 4396 1578 4400
rect 1582 4396 1588 4400
rect 1592 4396 1598 4400
rect 1602 4396 1608 4400
rect 1568 4395 1612 4396
rect 1568 4391 1573 4395
rect 1577 4391 1583 4395
rect 1587 4391 1593 4395
rect 1597 4391 1603 4395
rect 1607 4391 1612 4395
rect 1568 4390 1612 4391
rect 1572 4386 1578 4390
rect 1582 4386 1588 4390
rect 1592 4386 1598 4390
rect 1602 4386 1608 4390
rect 1568 4385 1612 4386
rect 1568 4381 1573 4385
rect 1577 4381 1583 4385
rect 1587 4381 1593 4385
rect 1597 4381 1603 4385
rect 1607 4381 1612 4385
rect 1568 4380 1612 4381
rect 1572 4376 1578 4380
rect 1582 4376 1588 4380
rect 1592 4376 1598 4380
rect 1602 4376 1608 4380
rect 1568 4375 1612 4376
rect 1568 4371 1573 4375
rect 1577 4371 1583 4375
rect 1587 4371 1593 4375
rect 1597 4371 1603 4375
rect 1607 4371 1612 4375
rect 1568 4370 1612 4371
rect 1572 4366 1578 4370
rect 1582 4366 1588 4370
rect 1592 4366 1598 4370
rect 1602 4366 1608 4370
rect 1568 4365 1612 4366
rect 1568 4361 1573 4365
rect 1577 4361 1583 4365
rect 1587 4361 1593 4365
rect 1597 4361 1603 4365
rect 1607 4361 1612 4365
rect 1881 4446 1887 4450
rect 1891 4446 1897 4450
rect 1901 4446 1907 4450
rect 1911 4446 1917 4450
rect 1877 4445 1921 4446
rect 1877 4441 1882 4445
rect 1886 4441 1892 4445
rect 1896 4441 1902 4445
rect 1906 4441 1912 4445
rect 1916 4441 1921 4445
rect 1877 4440 1921 4441
rect 1881 4436 1887 4440
rect 1891 4436 1897 4440
rect 1901 4436 1907 4440
rect 1911 4436 1917 4440
rect 1877 4435 1921 4436
rect 1877 4431 1882 4435
rect 1886 4431 1892 4435
rect 1896 4431 1902 4435
rect 1906 4431 1912 4435
rect 1916 4431 1921 4435
rect 1877 4430 1921 4431
rect 1881 4426 1887 4430
rect 1891 4426 1897 4430
rect 1901 4426 1907 4430
rect 1911 4426 1917 4430
rect 1877 4425 1921 4426
rect 1877 4421 1882 4425
rect 1886 4421 1892 4425
rect 1896 4421 1902 4425
rect 1906 4421 1912 4425
rect 1916 4421 1921 4425
rect 1877 4420 1921 4421
rect 1881 4416 1887 4420
rect 1891 4416 1897 4420
rect 1901 4416 1907 4420
rect 1911 4416 1917 4420
rect 1877 4415 1921 4416
rect 1877 4411 1882 4415
rect 1886 4411 1892 4415
rect 1896 4411 1902 4415
rect 1906 4411 1912 4415
rect 1916 4411 1921 4415
rect 1877 4410 1921 4411
rect 1881 4406 1887 4410
rect 1891 4406 1897 4410
rect 1901 4406 1907 4410
rect 1911 4406 1917 4410
rect 1877 4405 1921 4406
rect 1877 4401 1882 4405
rect 1886 4401 1892 4405
rect 1896 4401 1902 4405
rect 1906 4401 1912 4405
rect 1916 4401 1921 4405
rect 1877 4400 1921 4401
rect 1881 4396 1887 4400
rect 1891 4396 1897 4400
rect 1901 4396 1907 4400
rect 1911 4396 1917 4400
rect 1877 4395 1921 4396
rect 1877 4391 1882 4395
rect 1886 4391 1892 4395
rect 1896 4391 1902 4395
rect 1906 4391 1912 4395
rect 1916 4391 1921 4395
rect 1877 4390 1921 4391
rect 1881 4386 1887 4390
rect 1891 4386 1897 4390
rect 1901 4386 1907 4390
rect 1911 4386 1917 4390
rect 1877 4385 1921 4386
rect 1877 4381 1882 4385
rect 1886 4381 1892 4385
rect 1896 4381 1902 4385
rect 1906 4381 1912 4385
rect 1916 4381 1921 4385
rect 1877 4380 1921 4381
rect 1881 4376 1887 4380
rect 1891 4376 1897 4380
rect 1901 4376 1907 4380
rect 1911 4376 1917 4380
rect 1877 4375 1921 4376
rect 1877 4371 1882 4375
rect 1886 4371 1892 4375
rect 1896 4371 1902 4375
rect 1906 4371 1912 4375
rect 1916 4371 1921 4375
rect 1877 4370 1921 4371
rect 1881 4366 1887 4370
rect 1891 4366 1897 4370
rect 1901 4366 1907 4370
rect 1911 4366 1917 4370
rect 1877 4365 1921 4366
rect 1877 4361 1882 4365
rect 1886 4361 1892 4365
rect 1896 4361 1902 4365
rect 1906 4361 1912 4365
rect 1916 4361 1921 4365
rect 2190 4446 2196 4450
rect 2200 4446 2206 4450
rect 2210 4446 2216 4450
rect 2220 4446 2226 4450
rect 2186 4445 2230 4446
rect 2186 4441 2191 4445
rect 2195 4441 2201 4445
rect 2205 4441 2211 4445
rect 2215 4441 2221 4445
rect 2225 4441 2230 4445
rect 2186 4440 2230 4441
rect 2190 4436 2196 4440
rect 2200 4436 2206 4440
rect 2210 4436 2216 4440
rect 2220 4436 2226 4440
rect 2186 4435 2230 4436
rect 2186 4431 2191 4435
rect 2195 4431 2201 4435
rect 2205 4431 2211 4435
rect 2215 4431 2221 4435
rect 2225 4431 2230 4435
rect 2186 4430 2230 4431
rect 2190 4426 2196 4430
rect 2200 4426 2206 4430
rect 2210 4426 2216 4430
rect 2220 4426 2226 4430
rect 2186 4425 2230 4426
rect 2186 4421 2191 4425
rect 2195 4421 2201 4425
rect 2205 4421 2211 4425
rect 2215 4421 2221 4425
rect 2225 4421 2230 4425
rect 2186 4420 2230 4421
rect 2190 4416 2196 4420
rect 2200 4416 2206 4420
rect 2210 4416 2216 4420
rect 2220 4416 2226 4420
rect 2186 4415 2230 4416
rect 2186 4411 2191 4415
rect 2195 4411 2201 4415
rect 2205 4411 2211 4415
rect 2215 4411 2221 4415
rect 2225 4411 2230 4415
rect 2186 4410 2230 4411
rect 2190 4406 2196 4410
rect 2200 4406 2206 4410
rect 2210 4406 2216 4410
rect 2220 4406 2226 4410
rect 2186 4405 2230 4406
rect 2186 4401 2191 4405
rect 2195 4401 2201 4405
rect 2205 4401 2211 4405
rect 2215 4401 2221 4405
rect 2225 4401 2230 4405
rect 2186 4400 2230 4401
rect 2190 4396 2196 4400
rect 2200 4396 2206 4400
rect 2210 4396 2216 4400
rect 2220 4396 2226 4400
rect 2186 4395 2230 4396
rect 2186 4391 2191 4395
rect 2195 4391 2201 4395
rect 2205 4391 2211 4395
rect 2215 4391 2221 4395
rect 2225 4391 2230 4395
rect 2186 4390 2230 4391
rect 2190 4386 2196 4390
rect 2200 4386 2206 4390
rect 2210 4386 2216 4390
rect 2220 4386 2226 4390
rect 2186 4385 2230 4386
rect 2186 4381 2191 4385
rect 2195 4381 2201 4385
rect 2205 4381 2211 4385
rect 2215 4381 2221 4385
rect 2225 4381 2230 4385
rect 2186 4380 2230 4381
rect 2190 4376 2196 4380
rect 2200 4376 2206 4380
rect 2210 4376 2216 4380
rect 2220 4376 2226 4380
rect 2186 4375 2230 4376
rect 2186 4371 2191 4375
rect 2195 4371 2201 4375
rect 2205 4371 2211 4375
rect 2215 4371 2221 4375
rect 2225 4371 2230 4375
rect 2186 4370 2230 4371
rect 2190 4366 2196 4370
rect 2200 4366 2206 4370
rect 2210 4366 2216 4370
rect 2220 4366 2226 4370
rect 2186 4365 2230 4366
rect 2186 4361 2191 4365
rect 2195 4361 2201 4365
rect 2205 4361 2211 4365
rect 2215 4361 2221 4365
rect 2225 4361 2230 4365
rect 2499 4446 2505 4450
rect 2509 4446 2515 4450
rect 2519 4446 2525 4450
rect 2529 4446 2535 4450
rect 2495 4445 2539 4446
rect 2495 4441 2500 4445
rect 2504 4441 2510 4445
rect 2514 4441 2520 4445
rect 2524 4441 2530 4445
rect 2534 4441 2539 4445
rect 2495 4440 2539 4441
rect 2499 4436 2505 4440
rect 2509 4436 2515 4440
rect 2519 4436 2525 4440
rect 2529 4436 2535 4440
rect 2495 4435 2539 4436
rect 2495 4431 2500 4435
rect 2504 4431 2510 4435
rect 2514 4431 2520 4435
rect 2524 4431 2530 4435
rect 2534 4431 2539 4435
rect 2495 4430 2539 4431
rect 2499 4426 2505 4430
rect 2509 4426 2515 4430
rect 2519 4426 2525 4430
rect 2529 4426 2535 4430
rect 2495 4425 2539 4426
rect 2495 4421 2500 4425
rect 2504 4421 2510 4425
rect 2514 4421 2520 4425
rect 2524 4421 2530 4425
rect 2534 4421 2539 4425
rect 2495 4420 2539 4421
rect 2499 4416 2505 4420
rect 2509 4416 2515 4420
rect 2519 4416 2525 4420
rect 2529 4416 2535 4420
rect 2495 4415 2539 4416
rect 2495 4411 2500 4415
rect 2504 4411 2510 4415
rect 2514 4411 2520 4415
rect 2524 4411 2530 4415
rect 2534 4411 2539 4415
rect 2495 4410 2539 4411
rect 2499 4406 2505 4410
rect 2509 4406 2515 4410
rect 2519 4406 2525 4410
rect 2529 4406 2535 4410
rect 2495 4405 2539 4406
rect 2495 4401 2500 4405
rect 2504 4401 2510 4405
rect 2514 4401 2520 4405
rect 2524 4401 2530 4405
rect 2534 4401 2539 4405
rect 2495 4400 2539 4401
rect 2499 4396 2505 4400
rect 2509 4396 2515 4400
rect 2519 4396 2525 4400
rect 2529 4396 2535 4400
rect 2495 4395 2539 4396
rect 2495 4391 2500 4395
rect 2504 4391 2510 4395
rect 2514 4391 2520 4395
rect 2524 4391 2530 4395
rect 2534 4391 2539 4395
rect 2495 4390 2539 4391
rect 2499 4386 2505 4390
rect 2509 4386 2515 4390
rect 2519 4386 2525 4390
rect 2529 4386 2535 4390
rect 2495 4385 2539 4386
rect 2495 4381 2500 4385
rect 2504 4381 2510 4385
rect 2514 4381 2520 4385
rect 2524 4381 2530 4385
rect 2534 4381 2539 4385
rect 2495 4380 2539 4381
rect 2499 4376 2505 4380
rect 2509 4376 2515 4380
rect 2519 4376 2525 4380
rect 2529 4376 2535 4380
rect 2495 4375 2539 4376
rect 2495 4371 2500 4375
rect 2504 4371 2510 4375
rect 2514 4371 2520 4375
rect 2524 4371 2530 4375
rect 2534 4371 2539 4375
rect 2495 4370 2539 4371
rect 2499 4366 2505 4370
rect 2509 4366 2515 4370
rect 2519 4366 2525 4370
rect 2529 4366 2535 4370
rect 2495 4365 2539 4366
rect 2495 4361 2500 4365
rect 2504 4361 2510 4365
rect 2514 4361 2520 4365
rect 2524 4361 2530 4365
rect 2534 4361 2539 4365
rect 2808 4446 2814 4450
rect 2818 4446 2824 4450
rect 2828 4446 2834 4450
rect 2838 4446 2844 4450
rect 2804 4445 2848 4446
rect 2804 4441 2809 4445
rect 2813 4441 2819 4445
rect 2823 4441 2829 4445
rect 2833 4441 2839 4445
rect 2843 4441 2848 4445
rect 2804 4440 2848 4441
rect 2808 4436 2814 4440
rect 2818 4436 2824 4440
rect 2828 4436 2834 4440
rect 2838 4436 2844 4440
rect 2804 4435 2848 4436
rect 2804 4431 2809 4435
rect 2813 4431 2819 4435
rect 2823 4431 2829 4435
rect 2833 4431 2839 4435
rect 2843 4431 2848 4435
rect 2804 4430 2848 4431
rect 2808 4426 2814 4430
rect 2818 4426 2824 4430
rect 2828 4426 2834 4430
rect 2838 4426 2844 4430
rect 2804 4425 2848 4426
rect 2804 4421 2809 4425
rect 2813 4421 2819 4425
rect 2823 4421 2829 4425
rect 2833 4421 2839 4425
rect 2843 4421 2848 4425
rect 2804 4420 2848 4421
rect 2808 4416 2814 4420
rect 2818 4416 2824 4420
rect 2828 4416 2834 4420
rect 2838 4416 2844 4420
rect 2804 4415 2848 4416
rect 2804 4411 2809 4415
rect 2813 4411 2819 4415
rect 2823 4411 2829 4415
rect 2833 4411 2839 4415
rect 2843 4411 2848 4415
rect 2804 4410 2848 4411
rect 2808 4406 2814 4410
rect 2818 4406 2824 4410
rect 2828 4406 2834 4410
rect 2838 4406 2844 4410
rect 2804 4405 2848 4406
rect 2804 4401 2809 4405
rect 2813 4401 2819 4405
rect 2823 4401 2829 4405
rect 2833 4401 2839 4405
rect 2843 4401 2848 4405
rect 2804 4400 2848 4401
rect 2808 4396 2814 4400
rect 2818 4396 2824 4400
rect 2828 4396 2834 4400
rect 2838 4396 2844 4400
rect 2804 4395 2848 4396
rect 2804 4391 2809 4395
rect 2813 4391 2819 4395
rect 2823 4391 2829 4395
rect 2833 4391 2839 4395
rect 2843 4391 2848 4395
rect 2804 4390 2848 4391
rect 2808 4386 2814 4390
rect 2818 4386 2824 4390
rect 2828 4386 2834 4390
rect 2838 4386 2844 4390
rect 2804 4385 2848 4386
rect 2804 4381 2809 4385
rect 2813 4381 2819 4385
rect 2823 4381 2829 4385
rect 2833 4381 2839 4385
rect 2843 4381 2848 4385
rect 2804 4380 2848 4381
rect 2808 4376 2814 4380
rect 2818 4376 2824 4380
rect 2828 4376 2834 4380
rect 2838 4376 2844 4380
rect 2804 4375 2848 4376
rect 2804 4371 2809 4375
rect 2813 4371 2819 4375
rect 2823 4371 2829 4375
rect 2833 4371 2839 4375
rect 2843 4371 2848 4375
rect 2804 4370 2848 4371
rect 2808 4366 2814 4370
rect 2818 4366 2824 4370
rect 2828 4366 2834 4370
rect 2838 4366 2844 4370
rect 2804 4365 2848 4366
rect 2804 4361 2809 4365
rect 2813 4361 2819 4365
rect 2823 4361 2829 4365
rect 2833 4361 2839 4365
rect 2843 4361 2848 4365
rect 3117 4446 3123 4450
rect 3127 4446 3133 4450
rect 3137 4446 3143 4450
rect 3147 4446 3153 4450
rect 3113 4445 3157 4446
rect 3113 4441 3118 4445
rect 3122 4441 3128 4445
rect 3132 4441 3138 4445
rect 3142 4441 3148 4445
rect 3152 4441 3157 4445
rect 3113 4440 3157 4441
rect 3117 4436 3123 4440
rect 3127 4436 3133 4440
rect 3137 4436 3143 4440
rect 3147 4436 3153 4440
rect 3113 4435 3157 4436
rect 3113 4431 3118 4435
rect 3122 4431 3128 4435
rect 3132 4431 3138 4435
rect 3142 4431 3148 4435
rect 3152 4431 3157 4435
rect 3113 4430 3157 4431
rect 3117 4426 3123 4430
rect 3127 4426 3133 4430
rect 3137 4426 3143 4430
rect 3147 4426 3153 4430
rect 3113 4425 3157 4426
rect 3113 4421 3118 4425
rect 3122 4421 3128 4425
rect 3132 4421 3138 4425
rect 3142 4421 3148 4425
rect 3152 4421 3157 4425
rect 3113 4420 3157 4421
rect 3117 4416 3123 4420
rect 3127 4416 3133 4420
rect 3137 4416 3143 4420
rect 3147 4416 3153 4420
rect 3113 4415 3157 4416
rect 3113 4411 3118 4415
rect 3122 4411 3128 4415
rect 3132 4411 3138 4415
rect 3142 4411 3148 4415
rect 3152 4411 3157 4415
rect 3113 4410 3157 4411
rect 3117 4406 3123 4410
rect 3127 4406 3133 4410
rect 3137 4406 3143 4410
rect 3147 4406 3153 4410
rect 3113 4405 3157 4406
rect 3113 4401 3118 4405
rect 3122 4401 3128 4405
rect 3132 4401 3138 4405
rect 3142 4401 3148 4405
rect 3152 4401 3157 4405
rect 3113 4400 3157 4401
rect 3117 4396 3123 4400
rect 3127 4396 3133 4400
rect 3137 4396 3143 4400
rect 3147 4396 3153 4400
rect 3113 4395 3157 4396
rect 3113 4391 3118 4395
rect 3122 4391 3128 4395
rect 3132 4391 3138 4395
rect 3142 4391 3148 4395
rect 3152 4391 3157 4395
rect 3113 4390 3157 4391
rect 3117 4386 3123 4390
rect 3127 4386 3133 4390
rect 3137 4386 3143 4390
rect 3147 4386 3153 4390
rect 3113 4385 3157 4386
rect 3113 4381 3118 4385
rect 3122 4381 3128 4385
rect 3132 4381 3138 4385
rect 3142 4381 3148 4385
rect 3152 4381 3157 4385
rect 3113 4380 3157 4381
rect 3117 4376 3123 4380
rect 3127 4376 3133 4380
rect 3137 4376 3143 4380
rect 3147 4376 3153 4380
rect 3113 4375 3157 4376
rect 3113 4371 3118 4375
rect 3122 4371 3128 4375
rect 3132 4371 3138 4375
rect 3142 4371 3148 4375
rect 3152 4371 3157 4375
rect 3113 4370 3157 4371
rect 3117 4366 3123 4370
rect 3127 4366 3133 4370
rect 3137 4366 3143 4370
rect 3147 4366 3153 4370
rect 3113 4365 3157 4366
rect 3113 4361 3118 4365
rect 3122 4361 3128 4365
rect 3132 4361 3138 4365
rect 3142 4361 3148 4365
rect 3152 4361 3157 4365
rect 3426 4446 3432 4450
rect 3436 4446 3442 4450
rect 3446 4446 3452 4450
rect 3456 4446 3462 4450
rect 3422 4445 3466 4446
rect 3422 4441 3427 4445
rect 3431 4441 3437 4445
rect 3441 4441 3447 4445
rect 3451 4441 3457 4445
rect 3461 4441 3466 4445
rect 3422 4440 3466 4441
rect 3426 4436 3432 4440
rect 3436 4436 3442 4440
rect 3446 4436 3452 4440
rect 3456 4436 3462 4440
rect 3422 4435 3466 4436
rect 3422 4431 3427 4435
rect 3431 4431 3437 4435
rect 3441 4431 3447 4435
rect 3451 4431 3457 4435
rect 3461 4431 3466 4435
rect 3422 4430 3466 4431
rect 3426 4426 3432 4430
rect 3436 4426 3442 4430
rect 3446 4426 3452 4430
rect 3456 4426 3462 4430
rect 3422 4425 3466 4426
rect 3422 4421 3427 4425
rect 3431 4421 3437 4425
rect 3441 4421 3447 4425
rect 3451 4421 3457 4425
rect 3461 4421 3466 4425
rect 3422 4420 3466 4421
rect 3426 4416 3432 4420
rect 3436 4416 3442 4420
rect 3446 4416 3452 4420
rect 3456 4416 3462 4420
rect 3422 4415 3466 4416
rect 3422 4411 3427 4415
rect 3431 4411 3437 4415
rect 3441 4411 3447 4415
rect 3451 4411 3457 4415
rect 3461 4411 3466 4415
rect 3422 4410 3466 4411
rect 3426 4406 3432 4410
rect 3436 4406 3442 4410
rect 3446 4406 3452 4410
rect 3456 4406 3462 4410
rect 3422 4405 3466 4406
rect 3422 4401 3427 4405
rect 3431 4401 3437 4405
rect 3441 4401 3447 4405
rect 3451 4401 3457 4405
rect 3461 4401 3466 4405
rect 3422 4400 3466 4401
rect 3426 4396 3432 4400
rect 3436 4396 3442 4400
rect 3446 4396 3452 4400
rect 3456 4396 3462 4400
rect 3422 4395 3466 4396
rect 3422 4391 3427 4395
rect 3431 4391 3437 4395
rect 3441 4391 3447 4395
rect 3451 4391 3457 4395
rect 3461 4391 3466 4395
rect 3422 4390 3466 4391
rect 3426 4386 3432 4390
rect 3436 4386 3442 4390
rect 3446 4386 3452 4390
rect 3456 4386 3462 4390
rect 3422 4385 3466 4386
rect 3422 4381 3427 4385
rect 3431 4381 3437 4385
rect 3441 4381 3447 4385
rect 3451 4381 3457 4385
rect 3461 4381 3466 4385
rect 3422 4380 3466 4381
rect 3426 4376 3432 4380
rect 3436 4376 3442 4380
rect 3446 4376 3452 4380
rect 3456 4376 3462 4380
rect 3422 4375 3466 4376
rect 3422 4371 3427 4375
rect 3431 4371 3437 4375
rect 3441 4371 3447 4375
rect 3451 4371 3457 4375
rect 3461 4371 3466 4375
rect 3422 4370 3466 4371
rect 3426 4366 3432 4370
rect 3436 4366 3442 4370
rect 3446 4366 3452 4370
rect 3456 4366 3462 4370
rect 3422 4365 3466 4366
rect 3422 4361 3427 4365
rect 3431 4361 3437 4365
rect 3441 4361 3447 4365
rect 3451 4361 3457 4365
rect 3461 4361 3466 4365
rect 3735 4446 3741 4450
rect 3745 4446 3751 4450
rect 3755 4446 3761 4450
rect 3765 4446 3771 4450
rect 3731 4445 3775 4446
rect 3731 4441 3736 4445
rect 3740 4441 3746 4445
rect 3750 4441 3756 4445
rect 3760 4441 3766 4445
rect 3770 4441 3775 4445
rect 3731 4440 3775 4441
rect 3735 4436 3741 4440
rect 3745 4436 3751 4440
rect 3755 4436 3761 4440
rect 3765 4436 3771 4440
rect 3731 4435 3775 4436
rect 3731 4431 3736 4435
rect 3740 4431 3746 4435
rect 3750 4431 3756 4435
rect 3760 4431 3766 4435
rect 3770 4431 3775 4435
rect 3731 4430 3775 4431
rect 3735 4426 3741 4430
rect 3745 4426 3751 4430
rect 3755 4426 3761 4430
rect 3765 4426 3771 4430
rect 3731 4425 3775 4426
rect 3731 4421 3736 4425
rect 3740 4421 3746 4425
rect 3750 4421 3756 4425
rect 3760 4421 3766 4425
rect 3770 4421 3775 4425
rect 3731 4420 3775 4421
rect 3735 4416 3741 4420
rect 3745 4416 3751 4420
rect 3755 4416 3761 4420
rect 3765 4416 3771 4420
rect 3731 4415 3775 4416
rect 3731 4411 3736 4415
rect 3740 4411 3746 4415
rect 3750 4411 3756 4415
rect 3760 4411 3766 4415
rect 3770 4411 3775 4415
rect 3731 4410 3775 4411
rect 3735 4406 3741 4410
rect 3745 4406 3751 4410
rect 3755 4406 3761 4410
rect 3765 4406 3771 4410
rect 3731 4405 3775 4406
rect 3731 4401 3736 4405
rect 3740 4401 3746 4405
rect 3750 4401 3756 4405
rect 3760 4401 3766 4405
rect 3770 4401 3775 4405
rect 3731 4400 3775 4401
rect 3735 4396 3741 4400
rect 3745 4396 3751 4400
rect 3755 4396 3761 4400
rect 3765 4396 3771 4400
rect 3731 4395 3775 4396
rect 3731 4391 3736 4395
rect 3740 4391 3746 4395
rect 3750 4391 3756 4395
rect 3760 4391 3766 4395
rect 3770 4391 3775 4395
rect 3731 4390 3775 4391
rect 3735 4386 3741 4390
rect 3745 4386 3751 4390
rect 3755 4386 3761 4390
rect 3765 4386 3771 4390
rect 3731 4385 3775 4386
rect 3731 4381 3736 4385
rect 3740 4381 3746 4385
rect 3750 4381 3756 4385
rect 3760 4381 3766 4385
rect 3770 4381 3775 4385
rect 3731 4380 3775 4381
rect 3735 4376 3741 4380
rect 3745 4376 3751 4380
rect 3755 4376 3761 4380
rect 3765 4376 3771 4380
rect 3731 4375 3775 4376
rect 3731 4371 3736 4375
rect 3740 4371 3746 4375
rect 3750 4371 3756 4375
rect 3760 4371 3766 4375
rect 3770 4371 3775 4375
rect 3731 4370 3775 4371
rect 3735 4366 3741 4370
rect 3745 4366 3751 4370
rect 3755 4366 3761 4370
rect 3765 4366 3771 4370
rect 3731 4365 3775 4366
rect 3731 4361 3736 4365
rect 3740 4361 3746 4365
rect 3750 4361 3756 4365
rect 3760 4361 3766 4365
rect 3770 4361 3775 4365
<< pdiffusion >>
rect 1556 9949 1562 9953
rect 1566 9949 1572 9953
rect 1576 9949 1582 9953
rect 1586 9949 1592 9953
rect 1596 9949 1601 9953
rect 1556 9948 1601 9949
rect 1556 9944 1557 9948
rect 1561 9944 1567 9948
rect 1571 9944 1577 9948
rect 1581 9944 1587 9948
rect 1591 9944 1597 9948
rect 1556 9943 1601 9944
rect 1556 9939 1562 9943
rect 1566 9939 1572 9943
rect 1576 9939 1582 9943
rect 1586 9939 1592 9943
rect 1596 9939 1601 9943
rect 1556 9938 1601 9939
rect 1556 9934 1557 9938
rect 1561 9934 1567 9938
rect 1571 9934 1577 9938
rect 1581 9934 1587 9938
rect 1591 9934 1597 9938
rect 1556 9933 1601 9934
rect 1556 9929 1562 9933
rect 1566 9929 1572 9933
rect 1576 9929 1582 9933
rect 1586 9929 1592 9933
rect 1596 9929 1601 9933
rect 1556 9928 1601 9929
rect 1556 9924 1557 9928
rect 1561 9924 1567 9928
rect 1571 9924 1577 9928
rect 1581 9924 1587 9928
rect 1591 9924 1597 9928
rect 1556 9923 1601 9924
rect 1556 9919 1562 9923
rect 1566 9919 1572 9923
rect 1576 9919 1582 9923
rect 1586 9919 1592 9923
rect 1596 9919 1601 9923
rect 1556 9918 1601 9919
rect 1556 9914 1557 9918
rect 1561 9914 1567 9918
rect 1571 9914 1577 9918
rect 1581 9914 1587 9918
rect 1591 9914 1597 9918
rect 1556 9913 1601 9914
rect 1556 9909 1562 9913
rect 1566 9909 1572 9913
rect 1576 9909 1582 9913
rect 1586 9909 1592 9913
rect 1596 9909 1601 9913
rect 1556 9908 1601 9909
rect 1556 9904 1557 9908
rect 1561 9904 1567 9908
rect 1571 9904 1577 9908
rect 1581 9904 1587 9908
rect 1591 9904 1597 9908
rect 1556 9903 1601 9904
rect 1556 9899 1562 9903
rect 1566 9899 1572 9903
rect 1576 9899 1582 9903
rect 1586 9899 1592 9903
rect 1596 9899 1601 9903
rect 1556 9898 1601 9899
rect 1556 9894 1557 9898
rect 1561 9894 1567 9898
rect 1571 9894 1577 9898
rect 1581 9894 1587 9898
rect 1591 9894 1597 9898
rect 1556 9893 1601 9894
rect 1556 9889 1562 9893
rect 1566 9889 1572 9893
rect 1576 9889 1582 9893
rect 1586 9889 1592 9893
rect 1596 9889 1601 9893
rect 1556 9888 1601 9889
rect 1556 9884 1557 9888
rect 1561 9884 1567 9888
rect 1571 9884 1577 9888
rect 1581 9884 1587 9888
rect 1591 9884 1597 9888
rect 1556 9883 1601 9884
rect 1556 9879 1562 9883
rect 1566 9879 1572 9883
rect 1576 9879 1582 9883
rect 1586 9879 1592 9883
rect 1596 9879 1601 9883
rect 1556 9878 1601 9879
rect 1556 9874 1557 9878
rect 1561 9874 1567 9878
rect 1571 9874 1577 9878
rect 1581 9874 1587 9878
rect 1591 9874 1597 9878
rect 1556 9873 1601 9874
rect 1556 9869 1562 9873
rect 1566 9869 1572 9873
rect 1576 9869 1582 9873
rect 1586 9869 1592 9873
rect 1596 9869 1601 9873
rect 1556 9868 1601 9869
rect 1556 9864 1557 9868
rect 1561 9864 1567 9868
rect 1571 9864 1577 9868
rect 1581 9864 1587 9868
rect 1591 9864 1597 9868
rect 1865 9949 1871 9953
rect 1875 9949 1881 9953
rect 1885 9949 1891 9953
rect 1895 9949 1901 9953
rect 1905 9949 1910 9953
rect 1865 9948 1910 9949
rect 1865 9944 1866 9948
rect 1870 9944 1876 9948
rect 1880 9944 1886 9948
rect 1890 9944 1896 9948
rect 1900 9944 1906 9948
rect 1865 9943 1910 9944
rect 1865 9939 1871 9943
rect 1875 9939 1881 9943
rect 1885 9939 1891 9943
rect 1895 9939 1901 9943
rect 1905 9939 1910 9943
rect 1865 9938 1910 9939
rect 1865 9934 1866 9938
rect 1870 9934 1876 9938
rect 1880 9934 1886 9938
rect 1890 9934 1896 9938
rect 1900 9934 1906 9938
rect 1865 9933 1910 9934
rect 1865 9929 1871 9933
rect 1875 9929 1881 9933
rect 1885 9929 1891 9933
rect 1895 9929 1901 9933
rect 1905 9929 1910 9933
rect 1865 9928 1910 9929
rect 1865 9924 1866 9928
rect 1870 9924 1876 9928
rect 1880 9924 1886 9928
rect 1890 9924 1896 9928
rect 1900 9924 1906 9928
rect 1865 9923 1910 9924
rect 1865 9919 1871 9923
rect 1875 9919 1881 9923
rect 1885 9919 1891 9923
rect 1895 9919 1901 9923
rect 1905 9919 1910 9923
rect 1865 9918 1910 9919
rect 1865 9914 1866 9918
rect 1870 9914 1876 9918
rect 1880 9914 1886 9918
rect 1890 9914 1896 9918
rect 1900 9914 1906 9918
rect 1865 9913 1910 9914
rect 1865 9909 1871 9913
rect 1875 9909 1881 9913
rect 1885 9909 1891 9913
rect 1895 9909 1901 9913
rect 1905 9909 1910 9913
rect 1865 9908 1910 9909
rect 1865 9904 1866 9908
rect 1870 9904 1876 9908
rect 1880 9904 1886 9908
rect 1890 9904 1896 9908
rect 1900 9904 1906 9908
rect 1865 9903 1910 9904
rect 1865 9899 1871 9903
rect 1875 9899 1881 9903
rect 1885 9899 1891 9903
rect 1895 9899 1901 9903
rect 1905 9899 1910 9903
rect 1865 9898 1910 9899
rect 1865 9894 1866 9898
rect 1870 9894 1876 9898
rect 1880 9894 1886 9898
rect 1890 9894 1896 9898
rect 1900 9894 1906 9898
rect 1865 9893 1910 9894
rect 1865 9889 1871 9893
rect 1875 9889 1881 9893
rect 1885 9889 1891 9893
rect 1895 9889 1901 9893
rect 1905 9889 1910 9893
rect 1865 9888 1910 9889
rect 1865 9884 1866 9888
rect 1870 9884 1876 9888
rect 1880 9884 1886 9888
rect 1890 9884 1896 9888
rect 1900 9884 1906 9888
rect 1865 9883 1910 9884
rect 1865 9879 1871 9883
rect 1875 9879 1881 9883
rect 1885 9879 1891 9883
rect 1895 9879 1901 9883
rect 1905 9879 1910 9883
rect 1865 9878 1910 9879
rect 1865 9874 1866 9878
rect 1870 9874 1876 9878
rect 1880 9874 1886 9878
rect 1890 9874 1896 9878
rect 1900 9874 1906 9878
rect 1865 9873 1910 9874
rect 1865 9869 1871 9873
rect 1875 9869 1881 9873
rect 1885 9869 1891 9873
rect 1895 9869 1901 9873
rect 1905 9869 1910 9873
rect 1865 9868 1910 9869
rect 1865 9864 1866 9868
rect 1870 9864 1876 9868
rect 1880 9864 1886 9868
rect 1890 9864 1896 9868
rect 1900 9864 1906 9868
rect 2174 9949 2180 9953
rect 2184 9949 2190 9953
rect 2194 9949 2200 9953
rect 2204 9949 2210 9953
rect 2214 9949 2219 9953
rect 2174 9948 2219 9949
rect 2174 9944 2175 9948
rect 2179 9944 2185 9948
rect 2189 9944 2195 9948
rect 2199 9944 2205 9948
rect 2209 9944 2215 9948
rect 2174 9943 2219 9944
rect 2174 9939 2180 9943
rect 2184 9939 2190 9943
rect 2194 9939 2200 9943
rect 2204 9939 2210 9943
rect 2214 9939 2219 9943
rect 2174 9938 2219 9939
rect 2174 9934 2175 9938
rect 2179 9934 2185 9938
rect 2189 9934 2195 9938
rect 2199 9934 2205 9938
rect 2209 9934 2215 9938
rect 2174 9933 2219 9934
rect 2174 9929 2180 9933
rect 2184 9929 2190 9933
rect 2194 9929 2200 9933
rect 2204 9929 2210 9933
rect 2214 9929 2219 9933
rect 2174 9928 2219 9929
rect 2174 9924 2175 9928
rect 2179 9924 2185 9928
rect 2189 9924 2195 9928
rect 2199 9924 2205 9928
rect 2209 9924 2215 9928
rect 2174 9923 2219 9924
rect 2174 9919 2180 9923
rect 2184 9919 2190 9923
rect 2194 9919 2200 9923
rect 2204 9919 2210 9923
rect 2214 9919 2219 9923
rect 2174 9918 2219 9919
rect 2174 9914 2175 9918
rect 2179 9914 2185 9918
rect 2189 9914 2195 9918
rect 2199 9914 2205 9918
rect 2209 9914 2215 9918
rect 2174 9913 2219 9914
rect 2174 9909 2180 9913
rect 2184 9909 2190 9913
rect 2194 9909 2200 9913
rect 2204 9909 2210 9913
rect 2214 9909 2219 9913
rect 2174 9908 2219 9909
rect 2174 9904 2175 9908
rect 2179 9904 2185 9908
rect 2189 9904 2195 9908
rect 2199 9904 2205 9908
rect 2209 9904 2215 9908
rect 2174 9903 2219 9904
rect 2174 9899 2180 9903
rect 2184 9899 2190 9903
rect 2194 9899 2200 9903
rect 2204 9899 2210 9903
rect 2214 9899 2219 9903
rect 2174 9898 2219 9899
rect 2174 9894 2175 9898
rect 2179 9894 2185 9898
rect 2189 9894 2195 9898
rect 2199 9894 2205 9898
rect 2209 9894 2215 9898
rect 2174 9893 2219 9894
rect 2174 9889 2180 9893
rect 2184 9889 2190 9893
rect 2194 9889 2200 9893
rect 2204 9889 2210 9893
rect 2214 9889 2219 9893
rect 2174 9888 2219 9889
rect 2174 9884 2175 9888
rect 2179 9884 2185 9888
rect 2189 9884 2195 9888
rect 2199 9884 2205 9888
rect 2209 9884 2215 9888
rect 2174 9883 2219 9884
rect 2174 9879 2180 9883
rect 2184 9879 2190 9883
rect 2194 9879 2200 9883
rect 2204 9879 2210 9883
rect 2214 9879 2219 9883
rect 2174 9878 2219 9879
rect 2174 9874 2175 9878
rect 2179 9874 2185 9878
rect 2189 9874 2195 9878
rect 2199 9874 2205 9878
rect 2209 9874 2215 9878
rect 2174 9873 2219 9874
rect 2174 9869 2180 9873
rect 2184 9869 2190 9873
rect 2194 9869 2200 9873
rect 2204 9869 2210 9873
rect 2214 9869 2219 9873
rect 2174 9868 2219 9869
rect 2174 9864 2175 9868
rect 2179 9864 2185 9868
rect 2189 9864 2195 9868
rect 2199 9864 2205 9868
rect 2209 9864 2215 9868
rect 2483 9949 2489 9953
rect 2493 9949 2499 9953
rect 2503 9949 2509 9953
rect 2513 9949 2519 9953
rect 2523 9949 2528 9953
rect 2483 9948 2528 9949
rect 2483 9944 2484 9948
rect 2488 9944 2494 9948
rect 2498 9944 2504 9948
rect 2508 9944 2514 9948
rect 2518 9944 2524 9948
rect 2483 9943 2528 9944
rect 2483 9939 2489 9943
rect 2493 9939 2499 9943
rect 2503 9939 2509 9943
rect 2513 9939 2519 9943
rect 2523 9939 2528 9943
rect 2483 9938 2528 9939
rect 2483 9934 2484 9938
rect 2488 9934 2494 9938
rect 2498 9934 2504 9938
rect 2508 9934 2514 9938
rect 2518 9934 2524 9938
rect 2483 9933 2528 9934
rect 2483 9929 2489 9933
rect 2493 9929 2499 9933
rect 2503 9929 2509 9933
rect 2513 9929 2519 9933
rect 2523 9929 2528 9933
rect 2483 9928 2528 9929
rect 2483 9924 2484 9928
rect 2488 9924 2494 9928
rect 2498 9924 2504 9928
rect 2508 9924 2514 9928
rect 2518 9924 2524 9928
rect 2483 9923 2528 9924
rect 2483 9919 2489 9923
rect 2493 9919 2499 9923
rect 2503 9919 2509 9923
rect 2513 9919 2519 9923
rect 2523 9919 2528 9923
rect 2483 9918 2528 9919
rect 2483 9914 2484 9918
rect 2488 9914 2494 9918
rect 2498 9914 2504 9918
rect 2508 9914 2514 9918
rect 2518 9914 2524 9918
rect 2483 9913 2528 9914
rect 2483 9909 2489 9913
rect 2493 9909 2499 9913
rect 2503 9909 2509 9913
rect 2513 9909 2519 9913
rect 2523 9909 2528 9913
rect 2483 9908 2528 9909
rect 2483 9904 2484 9908
rect 2488 9904 2494 9908
rect 2498 9904 2504 9908
rect 2508 9904 2514 9908
rect 2518 9904 2524 9908
rect 2483 9903 2528 9904
rect 2483 9899 2489 9903
rect 2493 9899 2499 9903
rect 2503 9899 2509 9903
rect 2513 9899 2519 9903
rect 2523 9899 2528 9903
rect 2483 9898 2528 9899
rect 2483 9894 2484 9898
rect 2488 9894 2494 9898
rect 2498 9894 2504 9898
rect 2508 9894 2514 9898
rect 2518 9894 2524 9898
rect 2483 9893 2528 9894
rect 2483 9889 2489 9893
rect 2493 9889 2499 9893
rect 2503 9889 2509 9893
rect 2513 9889 2519 9893
rect 2523 9889 2528 9893
rect 2483 9888 2528 9889
rect 2483 9884 2484 9888
rect 2488 9884 2494 9888
rect 2498 9884 2504 9888
rect 2508 9884 2514 9888
rect 2518 9884 2524 9888
rect 2483 9883 2528 9884
rect 2483 9879 2489 9883
rect 2493 9879 2499 9883
rect 2503 9879 2509 9883
rect 2513 9879 2519 9883
rect 2523 9879 2528 9883
rect 2483 9878 2528 9879
rect 2483 9874 2484 9878
rect 2488 9874 2494 9878
rect 2498 9874 2504 9878
rect 2508 9874 2514 9878
rect 2518 9874 2524 9878
rect 2483 9873 2528 9874
rect 2483 9869 2489 9873
rect 2493 9869 2499 9873
rect 2503 9869 2509 9873
rect 2513 9869 2519 9873
rect 2523 9869 2528 9873
rect 2483 9868 2528 9869
rect 2483 9864 2484 9868
rect 2488 9864 2494 9868
rect 2498 9864 2504 9868
rect 2508 9864 2514 9868
rect 2518 9864 2524 9868
rect 2792 9949 2798 9953
rect 2802 9949 2808 9953
rect 2812 9949 2818 9953
rect 2822 9949 2828 9953
rect 2832 9949 2837 9953
rect 2792 9948 2837 9949
rect 2792 9944 2793 9948
rect 2797 9944 2803 9948
rect 2807 9944 2813 9948
rect 2817 9944 2823 9948
rect 2827 9944 2833 9948
rect 2792 9943 2837 9944
rect 2792 9939 2798 9943
rect 2802 9939 2808 9943
rect 2812 9939 2818 9943
rect 2822 9939 2828 9943
rect 2832 9939 2837 9943
rect 2792 9938 2837 9939
rect 2792 9934 2793 9938
rect 2797 9934 2803 9938
rect 2807 9934 2813 9938
rect 2817 9934 2823 9938
rect 2827 9934 2833 9938
rect 2792 9933 2837 9934
rect 2792 9929 2798 9933
rect 2802 9929 2808 9933
rect 2812 9929 2818 9933
rect 2822 9929 2828 9933
rect 2832 9929 2837 9933
rect 2792 9928 2837 9929
rect 2792 9924 2793 9928
rect 2797 9924 2803 9928
rect 2807 9924 2813 9928
rect 2817 9924 2823 9928
rect 2827 9924 2833 9928
rect 2792 9923 2837 9924
rect 2792 9919 2798 9923
rect 2802 9919 2808 9923
rect 2812 9919 2818 9923
rect 2822 9919 2828 9923
rect 2832 9919 2837 9923
rect 2792 9918 2837 9919
rect 2792 9914 2793 9918
rect 2797 9914 2803 9918
rect 2807 9914 2813 9918
rect 2817 9914 2823 9918
rect 2827 9914 2833 9918
rect 2792 9913 2837 9914
rect 2792 9909 2798 9913
rect 2802 9909 2808 9913
rect 2812 9909 2818 9913
rect 2822 9909 2828 9913
rect 2832 9909 2837 9913
rect 2792 9908 2837 9909
rect 2792 9904 2793 9908
rect 2797 9904 2803 9908
rect 2807 9904 2813 9908
rect 2817 9904 2823 9908
rect 2827 9904 2833 9908
rect 2792 9903 2837 9904
rect 2792 9899 2798 9903
rect 2802 9899 2808 9903
rect 2812 9899 2818 9903
rect 2822 9899 2828 9903
rect 2832 9899 2837 9903
rect 2792 9898 2837 9899
rect 2792 9894 2793 9898
rect 2797 9894 2803 9898
rect 2807 9894 2813 9898
rect 2817 9894 2823 9898
rect 2827 9894 2833 9898
rect 2792 9893 2837 9894
rect 2792 9889 2798 9893
rect 2802 9889 2808 9893
rect 2812 9889 2818 9893
rect 2822 9889 2828 9893
rect 2832 9889 2837 9893
rect 2792 9888 2837 9889
rect 2792 9884 2793 9888
rect 2797 9884 2803 9888
rect 2807 9884 2813 9888
rect 2817 9884 2823 9888
rect 2827 9884 2833 9888
rect 2792 9883 2837 9884
rect 2792 9879 2798 9883
rect 2802 9879 2808 9883
rect 2812 9879 2818 9883
rect 2822 9879 2828 9883
rect 2832 9879 2837 9883
rect 2792 9878 2837 9879
rect 2792 9874 2793 9878
rect 2797 9874 2803 9878
rect 2807 9874 2813 9878
rect 2817 9874 2823 9878
rect 2827 9874 2833 9878
rect 2792 9873 2837 9874
rect 2792 9869 2798 9873
rect 2802 9869 2808 9873
rect 2812 9869 2818 9873
rect 2822 9869 2828 9873
rect 2832 9869 2837 9873
rect 2792 9868 2837 9869
rect 2792 9864 2793 9868
rect 2797 9864 2803 9868
rect 2807 9864 2813 9868
rect 2817 9864 2823 9868
rect 2827 9864 2833 9868
rect 3101 9949 3107 9953
rect 3111 9949 3117 9953
rect 3121 9949 3127 9953
rect 3131 9949 3137 9953
rect 3141 9949 3146 9953
rect 3101 9948 3146 9949
rect 3101 9944 3102 9948
rect 3106 9944 3112 9948
rect 3116 9944 3122 9948
rect 3126 9944 3132 9948
rect 3136 9944 3142 9948
rect 3101 9943 3146 9944
rect 3101 9939 3107 9943
rect 3111 9939 3117 9943
rect 3121 9939 3127 9943
rect 3131 9939 3137 9943
rect 3141 9939 3146 9943
rect 3101 9938 3146 9939
rect 3101 9934 3102 9938
rect 3106 9934 3112 9938
rect 3116 9934 3122 9938
rect 3126 9934 3132 9938
rect 3136 9934 3142 9938
rect 3101 9933 3146 9934
rect 3101 9929 3107 9933
rect 3111 9929 3117 9933
rect 3121 9929 3127 9933
rect 3131 9929 3137 9933
rect 3141 9929 3146 9933
rect 3101 9928 3146 9929
rect 3101 9924 3102 9928
rect 3106 9924 3112 9928
rect 3116 9924 3122 9928
rect 3126 9924 3132 9928
rect 3136 9924 3142 9928
rect 3101 9923 3146 9924
rect 3101 9919 3107 9923
rect 3111 9919 3117 9923
rect 3121 9919 3127 9923
rect 3131 9919 3137 9923
rect 3141 9919 3146 9923
rect 3101 9918 3146 9919
rect 3101 9914 3102 9918
rect 3106 9914 3112 9918
rect 3116 9914 3122 9918
rect 3126 9914 3132 9918
rect 3136 9914 3142 9918
rect 3101 9913 3146 9914
rect 3101 9909 3107 9913
rect 3111 9909 3117 9913
rect 3121 9909 3127 9913
rect 3131 9909 3137 9913
rect 3141 9909 3146 9913
rect 3101 9908 3146 9909
rect 3101 9904 3102 9908
rect 3106 9904 3112 9908
rect 3116 9904 3122 9908
rect 3126 9904 3132 9908
rect 3136 9904 3142 9908
rect 3101 9903 3146 9904
rect 3101 9899 3107 9903
rect 3111 9899 3117 9903
rect 3121 9899 3127 9903
rect 3131 9899 3137 9903
rect 3141 9899 3146 9903
rect 3101 9898 3146 9899
rect 3101 9894 3102 9898
rect 3106 9894 3112 9898
rect 3116 9894 3122 9898
rect 3126 9894 3132 9898
rect 3136 9894 3142 9898
rect 3101 9893 3146 9894
rect 3101 9889 3107 9893
rect 3111 9889 3117 9893
rect 3121 9889 3127 9893
rect 3131 9889 3137 9893
rect 3141 9889 3146 9893
rect 3101 9888 3146 9889
rect 3101 9884 3102 9888
rect 3106 9884 3112 9888
rect 3116 9884 3122 9888
rect 3126 9884 3132 9888
rect 3136 9884 3142 9888
rect 3101 9883 3146 9884
rect 3101 9879 3107 9883
rect 3111 9879 3117 9883
rect 3121 9879 3127 9883
rect 3131 9879 3137 9883
rect 3141 9879 3146 9883
rect 3101 9878 3146 9879
rect 3101 9874 3102 9878
rect 3106 9874 3112 9878
rect 3116 9874 3122 9878
rect 3126 9874 3132 9878
rect 3136 9874 3142 9878
rect 3101 9873 3146 9874
rect 3101 9869 3107 9873
rect 3111 9869 3117 9873
rect 3121 9869 3127 9873
rect 3131 9869 3137 9873
rect 3141 9869 3146 9873
rect 3101 9868 3146 9869
rect 3101 9864 3102 9868
rect 3106 9864 3112 9868
rect 3116 9864 3122 9868
rect 3126 9864 3132 9868
rect 3136 9864 3142 9868
rect 3410 9949 3416 9953
rect 3420 9949 3426 9953
rect 3430 9949 3436 9953
rect 3440 9949 3446 9953
rect 3450 9949 3455 9953
rect 3410 9948 3455 9949
rect 3410 9944 3411 9948
rect 3415 9944 3421 9948
rect 3425 9944 3431 9948
rect 3435 9944 3441 9948
rect 3445 9944 3451 9948
rect 3410 9943 3455 9944
rect 3410 9939 3416 9943
rect 3420 9939 3426 9943
rect 3430 9939 3436 9943
rect 3440 9939 3446 9943
rect 3450 9939 3455 9943
rect 3410 9938 3455 9939
rect 3410 9934 3411 9938
rect 3415 9934 3421 9938
rect 3425 9934 3431 9938
rect 3435 9934 3441 9938
rect 3445 9934 3451 9938
rect 3410 9933 3455 9934
rect 3410 9929 3416 9933
rect 3420 9929 3426 9933
rect 3430 9929 3436 9933
rect 3440 9929 3446 9933
rect 3450 9929 3455 9933
rect 3410 9928 3455 9929
rect 3410 9924 3411 9928
rect 3415 9924 3421 9928
rect 3425 9924 3431 9928
rect 3435 9924 3441 9928
rect 3445 9924 3451 9928
rect 3410 9923 3455 9924
rect 3410 9919 3416 9923
rect 3420 9919 3426 9923
rect 3430 9919 3436 9923
rect 3440 9919 3446 9923
rect 3450 9919 3455 9923
rect 3410 9918 3455 9919
rect 3410 9914 3411 9918
rect 3415 9914 3421 9918
rect 3425 9914 3431 9918
rect 3435 9914 3441 9918
rect 3445 9914 3451 9918
rect 3410 9913 3455 9914
rect 3410 9909 3416 9913
rect 3420 9909 3426 9913
rect 3430 9909 3436 9913
rect 3440 9909 3446 9913
rect 3450 9909 3455 9913
rect 3410 9908 3455 9909
rect 3410 9904 3411 9908
rect 3415 9904 3421 9908
rect 3425 9904 3431 9908
rect 3435 9904 3441 9908
rect 3445 9904 3451 9908
rect 3410 9903 3455 9904
rect 3410 9899 3416 9903
rect 3420 9899 3426 9903
rect 3430 9899 3436 9903
rect 3440 9899 3446 9903
rect 3450 9899 3455 9903
rect 3410 9898 3455 9899
rect 3410 9894 3411 9898
rect 3415 9894 3421 9898
rect 3425 9894 3431 9898
rect 3435 9894 3441 9898
rect 3445 9894 3451 9898
rect 3410 9893 3455 9894
rect 3410 9889 3416 9893
rect 3420 9889 3426 9893
rect 3430 9889 3436 9893
rect 3440 9889 3446 9893
rect 3450 9889 3455 9893
rect 3410 9888 3455 9889
rect 3410 9884 3411 9888
rect 3415 9884 3421 9888
rect 3425 9884 3431 9888
rect 3435 9884 3441 9888
rect 3445 9884 3451 9888
rect 3410 9883 3455 9884
rect 3410 9879 3416 9883
rect 3420 9879 3426 9883
rect 3430 9879 3436 9883
rect 3440 9879 3446 9883
rect 3450 9879 3455 9883
rect 3410 9878 3455 9879
rect 3410 9874 3411 9878
rect 3415 9874 3421 9878
rect 3425 9874 3431 9878
rect 3435 9874 3441 9878
rect 3445 9874 3451 9878
rect 3410 9873 3455 9874
rect 3410 9869 3416 9873
rect 3420 9869 3426 9873
rect 3430 9869 3436 9873
rect 3440 9869 3446 9873
rect 3450 9869 3455 9873
rect 3410 9868 3455 9869
rect 3410 9864 3411 9868
rect 3415 9864 3421 9868
rect 3425 9864 3431 9868
rect 3435 9864 3441 9868
rect 3445 9864 3451 9868
rect 3719 9949 3725 9953
rect 3729 9949 3735 9953
rect 3739 9949 3745 9953
rect 3749 9949 3755 9953
rect 3759 9949 3764 9953
rect 3719 9948 3764 9949
rect 3719 9944 3720 9948
rect 3724 9944 3730 9948
rect 3734 9944 3740 9948
rect 3744 9944 3750 9948
rect 3754 9944 3760 9948
rect 3719 9943 3764 9944
rect 3719 9939 3725 9943
rect 3729 9939 3735 9943
rect 3739 9939 3745 9943
rect 3749 9939 3755 9943
rect 3759 9939 3764 9943
rect 3719 9938 3764 9939
rect 3719 9934 3720 9938
rect 3724 9934 3730 9938
rect 3734 9934 3740 9938
rect 3744 9934 3750 9938
rect 3754 9934 3760 9938
rect 3719 9933 3764 9934
rect 3719 9929 3725 9933
rect 3729 9929 3735 9933
rect 3739 9929 3745 9933
rect 3749 9929 3755 9933
rect 3759 9929 3764 9933
rect 3719 9928 3764 9929
rect 3719 9924 3720 9928
rect 3724 9924 3730 9928
rect 3734 9924 3740 9928
rect 3744 9924 3750 9928
rect 3754 9924 3760 9928
rect 3719 9923 3764 9924
rect 3719 9919 3725 9923
rect 3729 9919 3735 9923
rect 3739 9919 3745 9923
rect 3749 9919 3755 9923
rect 3759 9919 3764 9923
rect 3719 9918 3764 9919
rect 3719 9914 3720 9918
rect 3724 9914 3730 9918
rect 3734 9914 3740 9918
rect 3744 9914 3750 9918
rect 3754 9914 3760 9918
rect 3719 9913 3764 9914
rect 3719 9909 3725 9913
rect 3729 9909 3735 9913
rect 3739 9909 3745 9913
rect 3749 9909 3755 9913
rect 3759 9909 3764 9913
rect 3719 9908 3764 9909
rect 3719 9904 3720 9908
rect 3724 9904 3730 9908
rect 3734 9904 3740 9908
rect 3744 9904 3750 9908
rect 3754 9904 3760 9908
rect 3719 9903 3764 9904
rect 3719 9899 3725 9903
rect 3729 9899 3735 9903
rect 3739 9899 3745 9903
rect 3749 9899 3755 9903
rect 3759 9899 3764 9903
rect 3719 9898 3764 9899
rect 3719 9894 3720 9898
rect 3724 9894 3730 9898
rect 3734 9894 3740 9898
rect 3744 9894 3750 9898
rect 3754 9894 3760 9898
rect 3719 9893 3764 9894
rect 3719 9889 3725 9893
rect 3729 9889 3735 9893
rect 3739 9889 3745 9893
rect 3749 9889 3755 9893
rect 3759 9889 3764 9893
rect 3719 9888 3764 9889
rect 3719 9884 3720 9888
rect 3724 9884 3730 9888
rect 3734 9884 3740 9888
rect 3744 9884 3750 9888
rect 3754 9884 3760 9888
rect 3719 9883 3764 9884
rect 3719 9879 3725 9883
rect 3729 9879 3735 9883
rect 3739 9879 3745 9883
rect 3749 9879 3755 9883
rect 3759 9879 3764 9883
rect 3719 9878 3764 9879
rect 3719 9874 3720 9878
rect 3724 9874 3730 9878
rect 3734 9874 3740 9878
rect 3744 9874 3750 9878
rect 3754 9874 3760 9878
rect 3719 9873 3764 9874
rect 3719 9869 3725 9873
rect 3729 9869 3735 9873
rect 3739 9869 3745 9873
rect 3749 9869 3755 9873
rect 3759 9869 3764 9873
rect 3719 9868 3764 9869
rect 3719 9864 3720 9868
rect 3724 9864 3730 9868
rect 3734 9864 3740 9868
rect 3744 9864 3750 9868
rect 3754 9864 3760 9868
rect 4028 9949 4034 9953
rect 4038 9949 4044 9953
rect 4048 9949 4054 9953
rect 4058 9949 4064 9953
rect 4068 9949 4073 9953
rect 4028 9948 4073 9949
rect 4028 9944 4029 9948
rect 4033 9944 4039 9948
rect 4043 9944 4049 9948
rect 4053 9944 4059 9948
rect 4063 9944 4069 9948
rect 4028 9943 4073 9944
rect 4028 9939 4034 9943
rect 4038 9939 4044 9943
rect 4048 9939 4054 9943
rect 4058 9939 4064 9943
rect 4068 9939 4073 9943
rect 4028 9938 4073 9939
rect 4028 9934 4029 9938
rect 4033 9934 4039 9938
rect 4043 9934 4049 9938
rect 4053 9934 4059 9938
rect 4063 9934 4069 9938
rect 4028 9933 4073 9934
rect 4028 9929 4034 9933
rect 4038 9929 4044 9933
rect 4048 9929 4054 9933
rect 4058 9929 4064 9933
rect 4068 9929 4073 9933
rect 4028 9928 4073 9929
rect 4028 9924 4029 9928
rect 4033 9924 4039 9928
rect 4043 9924 4049 9928
rect 4053 9924 4059 9928
rect 4063 9924 4069 9928
rect 4028 9923 4073 9924
rect 4028 9919 4034 9923
rect 4038 9919 4044 9923
rect 4048 9919 4054 9923
rect 4058 9919 4064 9923
rect 4068 9919 4073 9923
rect 4028 9918 4073 9919
rect 4028 9914 4029 9918
rect 4033 9914 4039 9918
rect 4043 9914 4049 9918
rect 4053 9914 4059 9918
rect 4063 9914 4069 9918
rect 4028 9913 4073 9914
rect 4028 9909 4034 9913
rect 4038 9909 4044 9913
rect 4048 9909 4054 9913
rect 4058 9909 4064 9913
rect 4068 9909 4073 9913
rect 4028 9908 4073 9909
rect 4028 9904 4029 9908
rect 4033 9904 4039 9908
rect 4043 9904 4049 9908
rect 4053 9904 4059 9908
rect 4063 9904 4069 9908
rect 4028 9903 4073 9904
rect 4028 9899 4034 9903
rect 4038 9899 4044 9903
rect 4048 9899 4054 9903
rect 4058 9899 4064 9903
rect 4068 9899 4073 9903
rect 4028 9898 4073 9899
rect 4028 9894 4029 9898
rect 4033 9894 4039 9898
rect 4043 9894 4049 9898
rect 4053 9894 4059 9898
rect 4063 9894 4069 9898
rect 4028 9893 4073 9894
rect 4028 9889 4034 9893
rect 4038 9889 4044 9893
rect 4048 9889 4054 9893
rect 4058 9889 4064 9893
rect 4068 9889 4073 9893
rect 4028 9888 4073 9889
rect 4028 9884 4029 9888
rect 4033 9884 4039 9888
rect 4043 9884 4049 9888
rect 4053 9884 4059 9888
rect 4063 9884 4069 9888
rect 4028 9883 4073 9884
rect 4028 9879 4034 9883
rect 4038 9879 4044 9883
rect 4048 9879 4054 9883
rect 4058 9879 4064 9883
rect 4068 9879 4073 9883
rect 4028 9878 4073 9879
rect 4028 9874 4029 9878
rect 4033 9874 4039 9878
rect 4043 9874 4049 9878
rect 4053 9874 4059 9878
rect 4063 9874 4069 9878
rect 4028 9873 4073 9874
rect 4028 9869 4034 9873
rect 4038 9869 4044 9873
rect 4048 9869 4054 9873
rect 4058 9869 4064 9873
rect 4068 9869 4073 9873
rect 4028 9868 4073 9869
rect 4028 9864 4029 9868
rect 4033 9864 4039 9868
rect 4043 9864 4049 9868
rect 4053 9864 4059 9868
rect 4063 9864 4069 9868
rect 1778 9827 1782 9831
rect 1743 9826 1799 9827
rect 2087 9827 2091 9831
rect 2052 9826 2108 9827
rect 2396 9827 2400 9831
rect 2361 9826 2417 9827
rect 2705 9827 2709 9831
rect 2670 9826 2726 9827
rect 3014 9827 3018 9831
rect 2979 9826 3035 9827
rect 3941 9827 3945 9831
rect 3906 9826 3962 9827
rect 1743 9823 1799 9824
rect 1743 9818 1799 9819
rect 2052 9823 2108 9824
rect 2052 9818 2108 9819
rect 2361 9823 2417 9824
rect 2361 9818 2417 9819
rect 2670 9823 2726 9824
rect 2670 9818 2726 9819
rect 2979 9823 3035 9824
rect 2979 9818 3035 9819
rect 3906 9823 3962 9824
rect 3906 9818 3962 9819
rect 1743 9815 1799 9816
rect 1778 9811 1782 9815
rect 1743 9810 1799 9811
rect 2052 9815 2108 9816
rect 2087 9811 2091 9815
rect 2052 9810 2108 9811
rect 1743 9807 1799 9808
rect 1743 9802 1799 9803
rect 1743 9799 1799 9800
rect 1778 9795 1782 9799
rect 1743 9794 1799 9795
rect 1743 9791 1799 9792
rect 1743 9786 1799 9787
rect 2361 9815 2417 9816
rect 2396 9811 2400 9815
rect 2361 9810 2417 9811
rect 2052 9807 2108 9808
rect 2052 9802 2108 9803
rect 2052 9799 2108 9800
rect 2087 9795 2091 9799
rect 2052 9794 2108 9795
rect 2052 9791 2108 9792
rect 2052 9786 2108 9787
rect 2670 9815 2726 9816
rect 2705 9811 2709 9815
rect 2670 9810 2726 9811
rect 2361 9807 2417 9808
rect 2361 9802 2417 9803
rect 2361 9799 2417 9800
rect 2396 9795 2400 9799
rect 2361 9794 2417 9795
rect 2361 9791 2417 9792
rect 2361 9786 2417 9787
rect 2979 9815 3035 9816
rect 3014 9811 3018 9815
rect 2979 9810 3035 9811
rect 2670 9807 2726 9808
rect 2670 9802 2726 9803
rect 2670 9799 2726 9800
rect 2705 9795 2709 9799
rect 2670 9794 2726 9795
rect 2670 9791 2726 9792
rect 2670 9786 2726 9787
rect 3906 9815 3962 9816
rect 3941 9811 3945 9815
rect 3906 9810 3962 9811
rect 2979 9807 3035 9808
rect 2979 9802 3035 9803
rect 2979 9799 3035 9800
rect 3014 9795 3018 9799
rect 2979 9794 3035 9795
rect 2979 9791 3035 9792
rect 2979 9786 3035 9787
rect 3906 9807 3962 9808
rect 3906 9802 3962 9803
rect 3906 9799 3962 9800
rect 3941 9795 3945 9799
rect 3906 9794 3962 9795
rect 3906 9791 3962 9792
rect 3906 9786 3962 9787
rect 1743 9783 1799 9784
rect 1778 9779 1782 9783
rect 2052 9783 2108 9784
rect 2087 9779 2091 9783
rect 2361 9783 2417 9784
rect 2396 9779 2400 9783
rect 2670 9783 2726 9784
rect 2705 9779 2709 9783
rect 2979 9783 3035 9784
rect 3014 9779 3018 9783
rect 3906 9783 3962 9784
rect 3941 9779 3945 9783
rect 422 6390 423 6457
rect 427 6390 428 6457
rect 422 6386 428 6390
rect 422 6369 423 6386
rect 427 6369 428 6386
rect 430 6369 431 6457
rect 435 6369 436 6457
rect 438 6390 439 6457
rect 443 6390 444 6457
rect 438 6386 444 6390
rect 438 6378 439 6386
rect 443 6378 444 6386
rect 438 6369 444 6378
rect 446 6369 447 6457
rect 451 6369 452 6457
rect 454 6369 459 6457
rect 463 6390 464 6457
rect 468 6390 469 6457
rect 463 6386 469 6390
rect 463 6369 464 6386
rect 468 6369 469 6386
rect 471 6369 472 6457
rect 476 6369 477 6457
rect 479 6390 480 6457
rect 484 6390 485 6457
rect 479 6386 485 6390
rect 479 6378 480 6386
rect 484 6378 485 6386
rect 479 6369 485 6378
rect 487 6369 488 6457
rect 492 6369 493 6457
rect 495 6369 498 6457
rect 506 6390 507 6457
rect 511 6390 512 6457
rect 506 6386 512 6390
rect 506 6369 507 6386
rect 511 6369 512 6386
rect 514 6369 515 6457
rect 519 6369 520 6457
rect 522 6390 523 6457
rect 527 6390 528 6457
rect 522 6386 528 6390
rect 522 6378 523 6386
rect 527 6378 528 6386
rect 522 6369 528 6378
rect 530 6369 531 6457
rect 535 6369 536 6457
rect 538 6369 541 6457
rect 545 6390 546 6425
rect 550 6390 551 6425
rect 545 6386 551 6390
rect 545 6369 546 6386
rect 550 6369 551 6386
rect 553 6369 554 6425
rect 558 6369 559 6425
rect 561 6390 562 6425
rect 566 6390 567 6425
rect 561 6386 567 6390
rect 561 6369 562 6386
rect 566 6369 567 6386
rect 569 6369 570 6425
rect 574 6369 575 6425
rect 577 6390 578 6425
rect 582 6390 583 6425
rect 577 6386 583 6390
rect 577 6369 578 6386
rect 582 6369 583 6386
rect 585 6369 586 6425
rect 590 6369 591 6425
rect 593 6390 594 6425
rect 593 6386 598 6390
rect 593 6369 594 6386
rect 2855 9322 2856 9330
rect 2858 9322 2861 9330
rect 2863 9322 2864 9330
rect 2876 9322 2877 9330
rect 2879 9326 2880 9330
rect 2879 9322 2884 9326
rect 2892 9322 2893 9330
rect 2895 9322 2898 9330
rect 2900 9322 2901 9330
rect 2918 9322 2919 9330
rect 2921 9322 2922 9330
rect 2934 9322 2935 9330
rect 2937 9326 2938 9330
rect 2937 9322 2942 9326
rect 2950 9322 2951 9330
rect 2953 9322 2956 9330
rect 2958 9322 2959 9330
rect 2971 9322 2972 9330
rect 2974 9322 2975 9330
rect 2987 9322 2988 9330
rect 2990 9322 2993 9330
rect 2995 9322 2996 9330
rect 3008 9322 3009 9330
rect 3011 9326 3012 9330
rect 3011 9322 3016 9326
rect 3024 9322 3025 9330
rect 3027 9322 3030 9330
rect 3032 9322 3033 9330
rect 3050 9322 3051 9330
rect 3053 9322 3054 9330
rect 3066 9322 3067 9330
rect 3069 9326 3070 9330
rect 3069 9322 3074 9326
rect 3082 9322 3083 9330
rect 3085 9322 3088 9330
rect 3090 9322 3091 9330
rect 3103 9322 3104 9330
rect 3106 9322 3107 9330
rect 3119 9322 3120 9330
rect 3122 9322 3125 9330
rect 3127 9322 3128 9330
rect 3140 9322 3141 9330
rect 3143 9326 3144 9330
rect 3143 9322 3148 9326
rect 3156 9322 3157 9330
rect 3159 9322 3162 9330
rect 3164 9322 3165 9330
rect 3182 9322 3183 9330
rect 3185 9322 3186 9330
rect 3198 9322 3199 9330
rect 3201 9326 3202 9330
rect 3201 9322 3206 9326
rect 3214 9322 3215 9330
rect 3217 9322 3220 9330
rect 3222 9322 3223 9330
rect 3235 9322 3236 9330
rect 3238 9322 3239 9330
rect 3251 9322 3252 9330
rect 3254 9322 3257 9330
rect 3259 9322 3260 9330
rect 3272 9322 3273 9330
rect 3275 9326 3276 9330
rect 3275 9322 3280 9326
rect 3288 9322 3289 9330
rect 3291 9322 3294 9330
rect 3296 9322 3297 9330
rect 3314 9322 3315 9330
rect 3317 9322 3318 9330
rect 3330 9322 3331 9330
rect 3333 9326 3334 9330
rect 3333 9322 3338 9326
rect 3346 9322 3347 9330
rect 3349 9322 3352 9330
rect 3354 9322 3355 9330
rect 3367 9322 3368 9330
rect 3370 9322 3371 9330
rect 3800 9322 3801 9330
rect 3803 9322 3806 9330
rect 3808 9322 3809 9330
rect 3821 9322 3822 9330
rect 3824 9326 3825 9330
rect 3824 9322 3829 9326
rect 3837 9322 3838 9330
rect 3840 9322 3843 9330
rect 3845 9322 3846 9330
rect 3863 9322 3864 9330
rect 3866 9322 3867 9330
rect 3879 9322 3880 9330
rect 3882 9326 3883 9330
rect 3882 9322 3887 9326
rect 3895 9322 3896 9330
rect 3898 9322 3901 9330
rect 3903 9322 3904 9330
rect 3916 9322 3917 9330
rect 3919 9322 3920 9330
rect 3932 9322 3933 9330
rect 3935 9322 3938 9330
rect 3940 9322 3941 9330
rect 3953 9322 3954 9330
rect 3956 9326 3957 9330
rect 3956 9322 3961 9326
rect 3969 9322 3970 9330
rect 3972 9322 3975 9330
rect 3977 9322 3978 9330
rect 3995 9322 3996 9330
rect 3998 9322 3999 9330
rect 4011 9322 4012 9330
rect 4014 9326 4015 9330
rect 4014 9322 4019 9326
rect 4027 9322 4028 9330
rect 4030 9322 4033 9330
rect 4035 9322 4036 9330
rect 4048 9322 4049 9330
rect 4051 9322 4052 9330
rect 4064 9322 4065 9330
rect 4067 9322 4070 9330
rect 4072 9322 4073 9330
rect 4085 9322 4086 9330
rect 4088 9326 4089 9330
rect 4088 9322 4093 9326
rect 4101 9322 4102 9330
rect 4104 9322 4107 9330
rect 4109 9322 4110 9330
rect 4127 9322 4128 9330
rect 4130 9322 4131 9330
rect 4143 9322 4144 9330
rect 4146 9326 4147 9330
rect 4146 9322 4151 9326
rect 4159 9322 4160 9330
rect 4162 9322 4165 9330
rect 4167 9322 4168 9330
rect 4180 9322 4181 9330
rect 4183 9322 4184 9330
rect 4196 9322 4197 9330
rect 4199 9322 4202 9330
rect 4204 9322 4205 9330
rect 4217 9322 4218 9330
rect 4220 9326 4221 9330
rect 4220 9322 4225 9326
rect 4233 9322 4234 9330
rect 4236 9322 4239 9330
rect 4241 9322 4242 9330
rect 4259 9322 4260 9330
rect 4262 9322 4263 9330
rect 4275 9322 4276 9330
rect 4278 9326 4279 9330
rect 4278 9322 4283 9326
rect 4291 9322 4292 9330
rect 4294 9322 4297 9330
rect 4299 9322 4300 9330
rect 4312 9322 4313 9330
rect 4315 9322 4316 9330
rect 2503 9289 2504 9297
rect 2506 9289 2509 9297
rect 2511 9289 2512 9297
rect 2524 9289 2525 9297
rect 2527 9293 2528 9297
rect 2527 9289 2532 9293
rect 2540 9289 2541 9297
rect 2543 9289 2546 9297
rect 2548 9289 2549 9297
rect 2566 9289 2567 9297
rect 2569 9289 2570 9297
rect 2582 9289 2583 9297
rect 2585 9293 2586 9297
rect 2585 9289 2590 9293
rect 2598 9289 2599 9297
rect 2601 9289 2604 9297
rect 2606 9289 2607 9297
rect 2619 9289 2620 9297
rect 2622 9289 2623 9297
rect 3448 9289 3449 9297
rect 3451 9289 3454 9297
rect 3456 9289 3457 9297
rect 3469 9289 3470 9297
rect 3472 9293 3473 9297
rect 3472 9289 3477 9293
rect 3485 9289 3486 9297
rect 3488 9289 3491 9297
rect 3493 9289 3494 9297
rect 3511 9289 3512 9297
rect 3514 9289 3515 9297
rect 3527 9289 3528 9297
rect 3530 9293 3531 9297
rect 3530 9289 3535 9293
rect 3543 9289 3544 9297
rect 3546 9289 3549 9297
rect 3551 9289 3552 9297
rect 3564 9289 3565 9297
rect 3567 9289 3568 9297
rect 3034 9251 3035 9259
rect 3037 9251 3038 9259
rect 2860 9238 2861 9246
rect 2863 9238 2864 9246
rect 2876 9238 2877 9246
rect 2879 9238 2880 9246
rect 2892 9238 2893 9246
rect 2895 9238 2896 9246
rect 2911 9238 2916 9246
rect 2918 9238 2921 9246
rect 2923 9238 2924 9246
rect 2945 9238 2947 9246
rect 2949 9238 2950 9246
rect 2967 9238 2968 9246
rect 2970 9238 2971 9246
rect 2983 9238 2988 9246
rect 2990 9238 2993 9246
rect 2995 9238 2996 9246
rect 3010 9238 3011 9246
rect 3013 9238 3014 9246
rect 3058 9245 3061 9253
rect 3063 9245 3066 9253
rect 3068 9245 3069 9253
rect 3088 9251 3089 9259
rect 3091 9251 3092 9259
rect 3115 9251 3116 9259
rect 3118 9251 3119 9259
rect 3139 9245 3142 9253
rect 3144 9245 3147 9253
rect 3149 9245 3150 9253
rect 3169 9251 3170 9259
rect 3172 9251 3173 9259
rect 3979 9251 3980 9259
rect 3982 9251 3983 9259
rect 3805 9238 3806 9246
rect 3808 9238 3809 9246
rect 3821 9238 3822 9246
rect 3824 9238 3825 9246
rect 3837 9238 3838 9246
rect 3840 9238 3841 9246
rect 3856 9238 3861 9246
rect 3863 9238 3866 9246
rect 3868 9238 3869 9246
rect 3890 9238 3892 9246
rect 3894 9238 3895 9246
rect 3912 9238 3913 9246
rect 3915 9238 3916 9246
rect 3928 9238 3933 9246
rect 3935 9238 3938 9246
rect 3940 9238 3941 9246
rect 3955 9238 3956 9246
rect 3958 9238 3959 9246
rect 4003 9245 4006 9253
rect 4008 9245 4011 9253
rect 4013 9245 4014 9253
rect 4033 9251 4034 9259
rect 4036 9251 4037 9259
rect 4060 9251 4061 9259
rect 4063 9251 4064 9259
rect 4084 9245 4087 9253
rect 4089 9245 4092 9253
rect 4094 9245 4095 9253
rect 4114 9251 4115 9259
rect 4117 9251 4118 9259
rect 2494 9187 2495 9195
rect 2497 9187 2498 9195
rect 2510 9187 2511 9195
rect 2513 9187 2516 9195
rect 2518 9187 2519 9195
rect 2531 9191 2532 9195
rect 2527 9187 2532 9191
rect 2534 9187 2535 9195
rect 2547 9187 2548 9195
rect 2550 9187 2551 9195
rect 2568 9187 2569 9195
rect 2571 9187 2574 9195
rect 2576 9187 2577 9195
rect 2589 9191 2590 9195
rect 2585 9187 2590 9191
rect 2592 9187 2593 9195
rect 2605 9187 2606 9195
rect 2608 9187 2611 9195
rect 2613 9187 2614 9195
rect 3439 9187 3440 9195
rect 3442 9187 3443 9195
rect 3455 9187 3456 9195
rect 3458 9187 3461 9195
rect 3463 9187 3464 9195
rect 3476 9191 3477 9195
rect 3472 9187 3477 9191
rect 3479 9187 3480 9195
rect 3492 9187 3493 9195
rect 3495 9187 3496 9195
rect 3513 9187 3514 9195
rect 3516 9187 3519 9195
rect 3521 9187 3522 9195
rect 3534 9191 3535 9195
rect 3530 9187 3535 9191
rect 3537 9187 3538 9195
rect 3550 9187 3551 9195
rect 3553 9187 3556 9195
rect 3558 9187 3559 9195
rect 2860 9152 2861 9160
rect 2863 9152 2864 9160
rect 2876 9152 2877 9160
rect 2879 9152 2880 9160
rect 2892 9152 2893 9160
rect 2895 9152 2896 9160
rect 2911 9152 2916 9160
rect 2918 9152 2921 9160
rect 2923 9152 2924 9160
rect 2945 9152 2947 9160
rect 2949 9152 2950 9160
rect 2967 9152 2968 9160
rect 2970 9152 2971 9160
rect 2983 9152 2988 9160
rect 2990 9152 2993 9160
rect 2995 9152 2996 9160
rect 3010 9152 3011 9160
rect 3013 9152 3014 9160
rect 3058 9153 3061 9161
rect 3063 9153 3066 9161
rect 3068 9153 3069 9161
rect 3139 9153 3142 9161
rect 3144 9153 3147 9161
rect 3149 9153 3150 9161
rect 3805 9152 3806 9160
rect 3808 9152 3809 9160
rect 3821 9152 3822 9160
rect 3824 9152 3825 9160
rect 3837 9152 3838 9160
rect 3840 9152 3841 9160
rect 3856 9152 3861 9160
rect 3863 9152 3866 9160
rect 3868 9152 3869 9160
rect 3890 9152 3892 9160
rect 3894 9152 3895 9160
rect 3912 9152 3913 9160
rect 3915 9152 3916 9160
rect 3928 9152 3933 9160
rect 3935 9152 3938 9160
rect 3940 9152 3941 9160
rect 3955 9152 3956 9160
rect 3958 9152 3959 9160
rect 4003 9153 4006 9161
rect 4008 9153 4011 9161
rect 4013 9153 4014 9161
rect 4084 9153 4087 9161
rect 4089 9153 4092 9161
rect 4094 9153 4095 9161
rect 2860 9106 2861 9114
rect 2863 9106 2864 9114
rect 2876 9106 2877 9114
rect 2879 9106 2880 9114
rect 2892 9106 2893 9114
rect 2895 9106 2896 9114
rect 2911 9106 2916 9114
rect 2918 9106 2921 9114
rect 2923 9106 2924 9114
rect 2945 9106 2947 9114
rect 2949 9106 2950 9114
rect 2967 9106 2968 9114
rect 2970 9106 2971 9114
rect 2983 9106 2988 9114
rect 2990 9106 2993 9114
rect 2995 9106 2996 9114
rect 3010 9106 3011 9114
rect 3013 9106 3014 9114
rect 3058 9113 3061 9121
rect 3063 9113 3066 9121
rect 3068 9113 3069 9121
rect 3088 9119 3089 9127
rect 3091 9119 3092 9127
rect 3139 9119 3140 9127
rect 3142 9119 3143 9127
rect 3163 9113 3166 9121
rect 3168 9113 3171 9121
rect 3173 9113 3174 9121
rect 3193 9119 3194 9127
rect 3196 9119 3197 9127
rect 3805 9106 3806 9114
rect 3808 9106 3809 9114
rect 3821 9106 3822 9114
rect 3824 9106 3825 9114
rect 3837 9106 3838 9114
rect 3840 9106 3841 9114
rect 3856 9106 3861 9114
rect 3863 9106 3866 9114
rect 3868 9106 3869 9114
rect 3890 9106 3892 9114
rect 3894 9106 3895 9114
rect 3912 9106 3913 9114
rect 3915 9106 3916 9114
rect 3928 9106 3933 9114
rect 3935 9106 3938 9114
rect 3940 9106 3941 9114
rect 3955 9106 3956 9114
rect 3958 9106 3959 9114
rect 4003 9113 4006 9121
rect 4008 9113 4011 9121
rect 4013 9113 4014 9121
rect 4033 9119 4034 9127
rect 4036 9119 4037 9127
rect 4084 9119 4085 9127
rect 4087 9119 4088 9127
rect 3370 9090 3371 9098
rect 3373 9090 3374 9098
rect 3394 9084 3397 9092
rect 3399 9084 3402 9092
rect 3404 9084 3405 9092
rect 3424 9090 3425 9098
rect 3427 9090 3428 9098
rect 3556 9065 3557 9095
rect 3559 9065 3560 9095
rect 3609 9065 3610 9095
rect 3612 9065 3613 9095
rect 4108 9113 4111 9121
rect 4113 9113 4116 9121
rect 4118 9113 4119 9121
rect 4138 9119 4139 9127
rect 4141 9119 4142 9127
rect 2860 9020 2861 9028
rect 2863 9020 2864 9028
rect 2876 9020 2877 9028
rect 2879 9020 2880 9028
rect 2892 9020 2893 9028
rect 2895 9020 2896 9028
rect 2911 9020 2916 9028
rect 2918 9020 2921 9028
rect 2923 9020 2924 9028
rect 2945 9020 2947 9028
rect 2949 9020 2950 9028
rect 2967 9020 2968 9028
rect 2970 9020 2971 9028
rect 2983 9020 2988 9028
rect 2990 9020 2993 9028
rect 2995 9020 2996 9028
rect 3010 9020 3011 9028
rect 3013 9020 3014 9028
rect 3058 9022 3061 9030
rect 3063 9022 3066 9030
rect 3068 9022 3069 9030
rect 3163 9022 3166 9030
rect 3168 9022 3171 9030
rect 3173 9022 3174 9030
rect 3805 9020 3806 9028
rect 3808 9020 3809 9028
rect 3821 9020 3822 9028
rect 3824 9020 3825 9028
rect 3837 9020 3838 9028
rect 3840 9020 3841 9028
rect 3856 9020 3861 9028
rect 3863 9020 3866 9028
rect 3868 9020 3869 9028
rect 3890 9020 3892 9028
rect 3894 9020 3895 9028
rect 3912 9020 3913 9028
rect 3915 9020 3916 9028
rect 3928 9020 3933 9028
rect 3935 9020 3938 9028
rect 3940 9020 3941 9028
rect 3955 9020 3956 9028
rect 3958 9020 3959 9028
rect 4003 9022 4006 9030
rect 4008 9022 4011 9030
rect 4013 9022 4014 9030
rect 4108 9022 4111 9030
rect 4113 9022 4116 9030
rect 4118 9022 4119 9030
rect 2860 8974 2861 8982
rect 2863 8974 2864 8982
rect 2876 8974 2877 8982
rect 2879 8974 2880 8982
rect 2892 8974 2893 8982
rect 2895 8974 2896 8982
rect 2911 8974 2916 8982
rect 2918 8974 2921 8982
rect 2923 8974 2924 8982
rect 2945 8974 2947 8982
rect 2949 8974 2950 8982
rect 2967 8974 2968 8982
rect 2970 8974 2971 8982
rect 2983 8974 2988 8982
rect 2990 8974 2993 8982
rect 2995 8974 2996 8982
rect 3010 8974 3011 8982
rect 3013 8974 3014 8982
rect 3058 8981 3061 8989
rect 3063 8981 3066 8989
rect 3068 8981 3069 8989
rect 3088 8987 3089 8995
rect 3091 8987 3092 8995
rect 3115 8987 3116 8995
rect 3118 8987 3119 8995
rect 3139 8981 3142 8989
rect 3144 8981 3147 8989
rect 3149 8981 3150 8989
rect 3169 8987 3170 8995
rect 3172 8987 3173 8995
rect 3205 8987 3206 8995
rect 3208 8987 3209 8995
rect 3229 8981 3232 8989
rect 3234 8981 3237 8989
rect 3239 8981 3240 8989
rect 3259 8987 3260 8995
rect 3262 8987 3263 8995
rect 3394 8988 3397 8996
rect 3399 8988 3402 8996
rect 3404 8988 3405 8996
rect 3805 8974 3806 8982
rect 3808 8974 3809 8982
rect 3821 8974 3822 8982
rect 3824 8974 3825 8982
rect 3837 8974 3838 8982
rect 3840 8974 3841 8982
rect 3856 8974 3861 8982
rect 3863 8974 3866 8982
rect 3868 8974 3869 8982
rect 3890 8974 3892 8982
rect 3894 8974 3895 8982
rect 3912 8974 3913 8982
rect 3915 8974 3916 8982
rect 3928 8974 3933 8982
rect 3935 8974 3938 8982
rect 3940 8974 3941 8982
rect 3955 8974 3956 8982
rect 3958 8974 3959 8982
rect 4003 8981 4006 8989
rect 4008 8981 4011 8989
rect 4013 8981 4014 8989
rect 4033 8987 4034 8995
rect 4036 8987 4037 8995
rect 4060 8987 4061 8995
rect 4063 8987 4064 8995
rect 3348 8960 3349 8968
rect 3351 8960 3352 8968
rect 3370 8960 3371 8968
rect 3373 8960 3374 8968
rect 3394 8954 3397 8962
rect 3399 8954 3402 8962
rect 3404 8954 3405 8962
rect 3424 8960 3425 8968
rect 3427 8960 3428 8968
rect 3462 8935 3463 8965
rect 3465 8935 3466 8965
rect 3515 8935 3516 8965
rect 3518 8935 3519 8965
rect 4084 8981 4087 8989
rect 4089 8981 4092 8989
rect 4094 8981 4095 8989
rect 4114 8987 4115 8995
rect 4117 8987 4118 8995
rect 4150 8987 4151 8995
rect 4153 8987 4154 8995
rect 4174 8981 4177 8989
rect 4179 8981 4182 8989
rect 4184 8981 4185 8989
rect 4204 8987 4205 8995
rect 4207 8987 4208 8995
rect 2860 8888 2861 8896
rect 2863 8888 2864 8896
rect 2876 8888 2877 8896
rect 2879 8888 2880 8896
rect 2892 8888 2893 8896
rect 2895 8888 2896 8896
rect 2911 8888 2916 8896
rect 2918 8888 2921 8896
rect 2923 8888 2924 8896
rect 2945 8888 2947 8896
rect 2949 8888 2950 8896
rect 2967 8888 2968 8896
rect 2970 8888 2971 8896
rect 2983 8888 2988 8896
rect 2990 8888 2993 8896
rect 2995 8888 2996 8896
rect 3010 8888 3011 8896
rect 3013 8888 3014 8896
rect 3058 8887 3061 8895
rect 3063 8887 3066 8895
rect 3068 8887 3069 8895
rect 3139 8887 3142 8895
rect 3144 8887 3147 8895
rect 3149 8887 3150 8895
rect 3229 8887 3232 8895
rect 3234 8887 3237 8895
rect 3239 8887 3240 8895
rect 3805 8888 3806 8896
rect 3808 8888 3809 8896
rect 3821 8888 3822 8896
rect 3824 8888 3825 8896
rect 3837 8888 3838 8896
rect 3840 8888 3841 8896
rect 3856 8888 3861 8896
rect 3863 8888 3866 8896
rect 3868 8888 3869 8896
rect 3890 8888 3892 8896
rect 3894 8888 3895 8896
rect 3912 8888 3913 8896
rect 3915 8888 3916 8896
rect 3928 8888 3933 8896
rect 3935 8888 3938 8896
rect 3940 8888 3941 8896
rect 3955 8888 3956 8896
rect 3958 8888 3959 8896
rect 4003 8887 4006 8895
rect 4008 8887 4011 8895
rect 4013 8887 4014 8895
rect 4084 8887 4087 8895
rect 4089 8887 4092 8895
rect 4094 8887 4095 8895
rect 4174 8887 4177 8895
rect 4179 8887 4182 8895
rect 4184 8887 4185 8895
rect 2860 8842 2861 8850
rect 2863 8842 2864 8850
rect 2876 8842 2877 8850
rect 2879 8842 2880 8850
rect 2892 8842 2893 8850
rect 2895 8842 2896 8850
rect 2911 8842 2916 8850
rect 2918 8842 2921 8850
rect 2923 8842 2924 8850
rect 2945 8842 2947 8850
rect 2949 8842 2950 8850
rect 2967 8842 2968 8850
rect 2970 8842 2971 8850
rect 2983 8842 2988 8850
rect 2990 8842 2993 8850
rect 2995 8842 2996 8850
rect 3010 8842 3011 8850
rect 3013 8842 3014 8850
rect 3058 8849 3061 8857
rect 3063 8849 3066 8857
rect 3068 8849 3069 8857
rect 3088 8855 3089 8863
rect 3091 8855 3092 8863
rect 3394 8858 3397 8866
rect 3399 8858 3402 8866
rect 3404 8858 3405 8866
rect 3805 8842 3806 8850
rect 3808 8842 3809 8850
rect 3821 8842 3822 8850
rect 3824 8842 3825 8850
rect 3837 8842 3838 8850
rect 3840 8842 3841 8850
rect 3856 8842 3861 8850
rect 3863 8842 3866 8850
rect 3868 8842 3869 8850
rect 3890 8842 3892 8850
rect 3894 8842 3895 8850
rect 3912 8842 3913 8850
rect 3915 8842 3916 8850
rect 3928 8842 3933 8850
rect 3935 8842 3938 8850
rect 3940 8842 3941 8850
rect 3955 8842 3956 8850
rect 3958 8842 3959 8850
rect 4003 8849 4006 8857
rect 4008 8849 4011 8857
rect 4013 8849 4014 8857
rect 4033 8855 4034 8863
rect 4036 8855 4037 8863
rect 2371 8787 2372 8795
rect 2374 8787 2377 8795
rect 2379 8787 2380 8795
rect 2392 8787 2393 8795
rect 2395 8791 2396 8795
rect 2395 8787 2400 8791
rect 2408 8787 2409 8795
rect 2411 8787 2414 8795
rect 2416 8787 2417 8795
rect 2434 8787 2435 8795
rect 2437 8787 2438 8795
rect 2450 8787 2451 8795
rect 2453 8791 2454 8795
rect 2453 8787 2458 8791
rect 2466 8787 2467 8795
rect 2469 8787 2472 8795
rect 2474 8787 2475 8795
rect 2487 8787 2488 8795
rect 2490 8787 2491 8795
rect 2503 8787 2504 8795
rect 2506 8787 2509 8795
rect 2511 8787 2512 8795
rect 2524 8787 2525 8795
rect 2527 8791 2528 8795
rect 2527 8787 2532 8791
rect 2540 8787 2541 8795
rect 2543 8787 2546 8795
rect 2548 8787 2549 8795
rect 2566 8787 2567 8795
rect 2569 8787 2570 8795
rect 2582 8787 2583 8795
rect 2585 8791 2586 8795
rect 2585 8787 2590 8791
rect 2598 8787 2599 8795
rect 2601 8787 2604 8795
rect 2606 8787 2607 8795
rect 2619 8787 2620 8795
rect 2622 8787 2623 8795
rect 2635 8787 2636 8795
rect 2638 8787 2641 8795
rect 2643 8787 2644 8795
rect 2656 8787 2657 8795
rect 2659 8791 2660 8795
rect 2659 8787 2664 8791
rect 2672 8787 2673 8795
rect 2675 8787 2678 8795
rect 2680 8787 2681 8795
rect 2698 8787 2699 8795
rect 2701 8787 2702 8795
rect 2714 8787 2715 8795
rect 2717 8791 2718 8795
rect 2717 8787 2722 8791
rect 2730 8787 2731 8795
rect 2733 8787 2736 8795
rect 2738 8787 2739 8795
rect 2751 8787 2752 8795
rect 2754 8787 2755 8795
rect 3316 8787 3317 8795
rect 3319 8787 3322 8795
rect 3324 8787 3325 8795
rect 3337 8787 3338 8795
rect 3340 8791 3341 8795
rect 3340 8787 3345 8791
rect 3353 8787 3354 8795
rect 3356 8787 3359 8795
rect 3361 8787 3362 8795
rect 3379 8787 3380 8795
rect 3382 8787 3383 8795
rect 3395 8787 3396 8795
rect 3398 8791 3399 8795
rect 3398 8787 3403 8791
rect 3411 8787 3412 8795
rect 3414 8787 3417 8795
rect 3419 8787 3420 8795
rect 3432 8787 3433 8795
rect 3435 8787 3436 8795
rect 3448 8787 3449 8795
rect 3451 8787 3454 8795
rect 3456 8787 3457 8795
rect 3469 8787 3470 8795
rect 3472 8791 3473 8795
rect 3472 8787 3477 8791
rect 3485 8787 3486 8795
rect 3488 8787 3491 8795
rect 3493 8787 3494 8795
rect 3511 8787 3512 8795
rect 3514 8787 3515 8795
rect 3527 8787 3528 8795
rect 3530 8791 3531 8795
rect 3530 8787 3535 8791
rect 3543 8787 3544 8795
rect 3546 8787 3549 8795
rect 3551 8787 3552 8795
rect 3564 8787 3565 8795
rect 3567 8787 3568 8795
rect 3580 8787 3581 8795
rect 3583 8787 3586 8795
rect 3588 8787 3589 8795
rect 3601 8787 3602 8795
rect 3604 8791 3605 8795
rect 3604 8787 3609 8791
rect 3617 8787 3618 8795
rect 3620 8787 3623 8795
rect 3625 8787 3626 8795
rect 3643 8787 3644 8795
rect 3646 8787 3647 8795
rect 3659 8787 3660 8795
rect 3662 8791 3663 8795
rect 3662 8787 3667 8791
rect 3675 8787 3676 8795
rect 3678 8787 3681 8795
rect 3683 8787 3684 8795
rect 3696 8787 3697 8795
rect 3699 8787 3700 8795
rect 2860 8756 2861 8764
rect 2863 8756 2864 8764
rect 2876 8756 2877 8764
rect 2879 8756 2880 8764
rect 2892 8756 2893 8764
rect 2895 8756 2896 8764
rect 2911 8756 2916 8764
rect 2918 8756 2921 8764
rect 2923 8756 2924 8764
rect 2945 8756 2947 8764
rect 2949 8756 2950 8764
rect 2967 8756 2968 8764
rect 2970 8756 2971 8764
rect 2983 8756 2988 8764
rect 2990 8756 2993 8764
rect 2995 8756 2996 8764
rect 3010 8756 3011 8764
rect 3013 8756 3014 8764
rect 3058 8751 3061 8759
rect 3063 8751 3066 8759
rect 3068 8751 3069 8759
rect 3094 8756 3095 8764
rect 3097 8756 3098 8764
rect 3102 8756 3108 8764
rect 3112 8756 3113 8764
rect 3115 8756 3116 8764
rect 3137 8756 3138 8764
rect 3140 8756 3141 8764
rect 3153 8756 3154 8764
rect 3156 8756 3157 8764
rect 3172 8756 3177 8764
rect 3179 8756 3182 8764
rect 3184 8756 3185 8764
rect 3206 8756 3208 8764
rect 3210 8756 3211 8764
rect 3228 8756 3229 8764
rect 3231 8756 3232 8764
rect 3244 8756 3249 8764
rect 3251 8756 3254 8764
rect 3256 8756 3257 8764
rect 3271 8756 3272 8764
rect 3274 8756 3275 8764
rect 3805 8756 3806 8764
rect 3808 8756 3809 8764
rect 3821 8756 3822 8764
rect 3824 8756 3825 8764
rect 3837 8756 3838 8764
rect 3840 8756 3841 8764
rect 3856 8756 3861 8764
rect 3863 8756 3866 8764
rect 3868 8756 3869 8764
rect 3890 8756 3892 8764
rect 3894 8756 3895 8764
rect 3912 8756 3913 8764
rect 3915 8756 3916 8764
rect 3928 8756 3933 8764
rect 3935 8756 3938 8764
rect 3940 8756 3941 8764
rect 3955 8756 3956 8764
rect 3958 8756 3959 8764
rect 4003 8751 4006 8759
rect 4008 8751 4011 8759
rect 4013 8751 4014 8759
rect 4039 8756 4040 8764
rect 4042 8756 4043 8764
rect 4047 8756 4053 8764
rect 4057 8756 4058 8764
rect 4060 8756 4061 8764
rect 4082 8756 4083 8764
rect 4085 8756 4086 8764
rect 4098 8756 4099 8764
rect 4101 8756 4102 8764
rect 4117 8756 4122 8764
rect 4124 8756 4127 8764
rect 4129 8756 4130 8764
rect 4151 8756 4153 8764
rect 4155 8756 4156 8764
rect 4173 8756 4174 8764
rect 4176 8756 4177 8764
rect 4189 8756 4194 8764
rect 4196 8756 4199 8764
rect 4201 8756 4202 8764
rect 4216 8756 4217 8764
rect 4219 8756 4220 8764
rect 3154 8675 3155 8683
rect 3157 8675 3160 8683
rect 3162 8675 3163 8683
rect 3175 8675 3176 8683
rect 3178 8679 3179 8683
rect 3178 8675 3183 8679
rect 3191 8675 3192 8683
rect 3194 8675 3197 8683
rect 3199 8675 3200 8683
rect 3217 8675 3218 8683
rect 3220 8675 3221 8683
rect 3233 8675 3234 8683
rect 3236 8679 3237 8683
rect 3236 8675 3241 8679
rect 3249 8675 3250 8683
rect 3252 8675 3255 8683
rect 3257 8675 3258 8683
rect 3270 8675 3271 8683
rect 3273 8675 3274 8683
rect 4099 8675 4100 8683
rect 4102 8675 4105 8683
rect 4107 8675 4108 8683
rect 4120 8675 4121 8683
rect 4123 8679 4124 8683
rect 4123 8675 4128 8679
rect 4136 8675 4137 8683
rect 4139 8675 4142 8683
rect 4144 8675 4145 8683
rect 4162 8675 4163 8683
rect 4165 8675 4166 8683
rect 4178 8675 4179 8683
rect 4181 8679 4182 8683
rect 4181 8675 4186 8679
rect 4194 8675 4195 8683
rect 4197 8675 4200 8683
rect 4202 8675 4203 8683
rect 4215 8675 4216 8683
rect 4218 8675 4219 8683
rect 2371 8645 2372 8653
rect 2374 8645 2377 8653
rect 2379 8645 2380 8653
rect 2392 8645 2393 8653
rect 2395 8649 2396 8653
rect 2395 8645 2400 8649
rect 2408 8645 2409 8653
rect 2411 8645 2414 8653
rect 2416 8645 2417 8653
rect 2434 8645 2435 8653
rect 2437 8645 2438 8653
rect 2450 8645 2451 8653
rect 2453 8649 2454 8653
rect 2453 8645 2458 8649
rect 2466 8645 2467 8653
rect 2469 8645 2472 8653
rect 2474 8645 2475 8653
rect 2487 8645 2488 8653
rect 2490 8645 2491 8653
rect 2503 8645 2504 8653
rect 2506 8645 2509 8653
rect 2511 8645 2512 8653
rect 2524 8645 2525 8653
rect 2527 8649 2528 8653
rect 2527 8645 2532 8649
rect 2540 8645 2541 8653
rect 2543 8645 2546 8653
rect 2548 8645 2549 8653
rect 2566 8645 2567 8653
rect 2569 8645 2570 8653
rect 2582 8645 2583 8653
rect 2585 8649 2586 8653
rect 2585 8645 2590 8649
rect 2598 8645 2599 8653
rect 2601 8645 2604 8653
rect 2606 8645 2607 8653
rect 2619 8645 2620 8653
rect 2622 8645 2623 8653
rect 2635 8645 2636 8653
rect 2638 8645 2641 8653
rect 2643 8645 2644 8653
rect 2656 8645 2657 8653
rect 2659 8649 2660 8653
rect 2659 8645 2664 8649
rect 2672 8645 2673 8653
rect 2675 8645 2678 8653
rect 2680 8645 2681 8653
rect 2698 8645 2699 8653
rect 2701 8645 2702 8653
rect 2714 8645 2715 8653
rect 2717 8649 2718 8653
rect 2717 8645 2722 8649
rect 2730 8645 2731 8653
rect 2733 8645 2736 8653
rect 2738 8645 2739 8653
rect 2751 8645 2752 8653
rect 2754 8645 2755 8653
rect 3316 8645 3317 8653
rect 3319 8645 3322 8653
rect 3324 8645 3325 8653
rect 3337 8645 3338 8653
rect 3340 8649 3341 8653
rect 3340 8645 3345 8649
rect 3353 8645 3354 8653
rect 3356 8645 3359 8653
rect 3361 8645 3362 8653
rect 3379 8645 3380 8653
rect 3382 8645 3383 8653
rect 3395 8645 3396 8653
rect 3398 8649 3399 8653
rect 3398 8645 3403 8649
rect 3411 8645 3412 8653
rect 3414 8645 3417 8653
rect 3419 8645 3420 8653
rect 3432 8645 3433 8653
rect 3435 8645 3436 8653
rect 3448 8645 3449 8653
rect 3451 8645 3454 8653
rect 3456 8645 3457 8653
rect 3469 8645 3470 8653
rect 3472 8649 3473 8653
rect 3472 8645 3477 8649
rect 3485 8645 3486 8653
rect 3488 8645 3491 8653
rect 3493 8645 3494 8653
rect 3511 8645 3512 8653
rect 3514 8645 3515 8653
rect 3527 8645 3528 8653
rect 3530 8649 3531 8653
rect 3530 8645 3535 8649
rect 3543 8645 3544 8653
rect 3546 8645 3549 8653
rect 3551 8645 3552 8653
rect 3564 8645 3565 8653
rect 3567 8645 3568 8653
rect 3580 8645 3581 8653
rect 3583 8645 3586 8653
rect 3588 8645 3589 8653
rect 3601 8645 3602 8653
rect 3604 8649 3605 8653
rect 3604 8645 3609 8649
rect 3617 8645 3618 8653
rect 3620 8645 3623 8653
rect 3625 8645 3626 8653
rect 3643 8645 3644 8653
rect 3646 8645 3647 8653
rect 3659 8645 3660 8653
rect 3662 8649 3663 8653
rect 3662 8645 3667 8649
rect 3675 8645 3676 8653
rect 3678 8645 3681 8653
rect 3683 8645 3684 8653
rect 3696 8645 3697 8653
rect 3699 8645 3700 8653
rect 3154 8589 3155 8597
rect 3157 8589 3160 8597
rect 3162 8589 3163 8597
rect 3175 8589 3176 8597
rect 3178 8593 3179 8597
rect 3178 8589 3183 8593
rect 3191 8589 3192 8597
rect 3194 8589 3197 8597
rect 3199 8589 3200 8597
rect 3217 8589 3218 8597
rect 3220 8589 3221 8597
rect 3233 8589 3234 8597
rect 3236 8593 3237 8597
rect 3236 8589 3241 8593
rect 3249 8589 3250 8597
rect 3252 8589 3255 8597
rect 3257 8589 3258 8597
rect 3270 8589 3271 8597
rect 3273 8589 3274 8597
rect 4099 8589 4100 8597
rect 4102 8589 4105 8597
rect 4107 8589 4108 8597
rect 4120 8589 4121 8597
rect 4123 8593 4124 8597
rect 4123 8589 4128 8593
rect 4136 8589 4137 8597
rect 4139 8589 4142 8597
rect 4144 8589 4145 8597
rect 4162 8589 4163 8597
rect 4165 8589 4166 8597
rect 4178 8589 4179 8597
rect 4181 8593 4182 8597
rect 4181 8589 4186 8593
rect 4194 8589 4195 8597
rect 4197 8589 4200 8597
rect 4202 8589 4203 8597
rect 4215 8589 4216 8597
rect 4218 8589 4219 8597
rect 2371 8559 2372 8567
rect 2374 8559 2377 8567
rect 2379 8559 2380 8567
rect 2392 8559 2393 8567
rect 2395 8563 2396 8567
rect 2395 8559 2400 8563
rect 2408 8559 2409 8567
rect 2411 8559 2414 8567
rect 2416 8559 2417 8567
rect 2434 8559 2435 8567
rect 2437 8559 2438 8567
rect 2450 8559 2451 8567
rect 2453 8563 2454 8567
rect 2453 8559 2458 8563
rect 2466 8559 2467 8567
rect 2469 8559 2472 8567
rect 2474 8559 2475 8567
rect 2487 8559 2488 8567
rect 2490 8559 2491 8567
rect 2503 8559 2504 8567
rect 2506 8559 2509 8567
rect 2511 8559 2512 8567
rect 2524 8559 2525 8567
rect 2527 8563 2528 8567
rect 2527 8559 2532 8563
rect 2540 8559 2541 8567
rect 2543 8559 2546 8567
rect 2548 8559 2549 8567
rect 2566 8559 2567 8567
rect 2569 8559 2570 8567
rect 2582 8559 2583 8567
rect 2585 8563 2586 8567
rect 2585 8559 2590 8563
rect 2598 8559 2599 8567
rect 2601 8559 2604 8567
rect 2606 8559 2607 8567
rect 2619 8559 2620 8567
rect 2622 8559 2623 8567
rect 2635 8559 2636 8567
rect 2638 8559 2641 8567
rect 2643 8559 2644 8567
rect 2656 8559 2657 8567
rect 2659 8563 2660 8567
rect 2659 8559 2664 8563
rect 2672 8559 2673 8567
rect 2675 8559 2678 8567
rect 2680 8559 2681 8567
rect 2698 8559 2699 8567
rect 2701 8559 2702 8567
rect 2714 8559 2715 8567
rect 2717 8563 2718 8567
rect 2717 8559 2722 8563
rect 2730 8559 2731 8567
rect 2733 8559 2736 8567
rect 2738 8559 2739 8567
rect 2751 8559 2752 8567
rect 2754 8559 2755 8567
rect 3316 8559 3317 8567
rect 3319 8559 3322 8567
rect 3324 8559 3325 8567
rect 3337 8559 3338 8567
rect 3340 8563 3341 8567
rect 3340 8559 3345 8563
rect 3353 8559 3354 8567
rect 3356 8559 3359 8567
rect 3361 8559 3362 8567
rect 3379 8559 3380 8567
rect 3382 8559 3383 8567
rect 3395 8559 3396 8567
rect 3398 8563 3399 8567
rect 3398 8559 3403 8563
rect 3411 8559 3412 8567
rect 3414 8559 3417 8567
rect 3419 8559 3420 8567
rect 3432 8559 3433 8567
rect 3435 8559 3436 8567
rect 3448 8559 3449 8567
rect 3451 8559 3454 8567
rect 3456 8559 3457 8567
rect 3469 8559 3470 8567
rect 3472 8563 3473 8567
rect 3472 8559 3477 8563
rect 3485 8559 3486 8567
rect 3488 8559 3491 8567
rect 3493 8559 3494 8567
rect 3511 8559 3512 8567
rect 3514 8559 3515 8567
rect 3527 8559 3528 8567
rect 3530 8563 3531 8567
rect 3530 8559 3535 8563
rect 3543 8559 3544 8567
rect 3546 8559 3549 8567
rect 3551 8559 3552 8567
rect 3564 8559 3565 8567
rect 3567 8559 3568 8567
rect 3580 8559 3581 8567
rect 3583 8559 3586 8567
rect 3588 8559 3589 8567
rect 3601 8559 3602 8567
rect 3604 8563 3605 8567
rect 3604 8559 3609 8563
rect 3617 8559 3618 8567
rect 3620 8559 3623 8567
rect 3625 8559 3626 8567
rect 3643 8559 3644 8567
rect 3646 8559 3647 8567
rect 3659 8559 3660 8567
rect 3662 8563 3663 8567
rect 3662 8559 3667 8563
rect 3675 8559 3676 8567
rect 3678 8559 3681 8567
rect 3683 8559 3684 8567
rect 3696 8559 3697 8567
rect 3699 8559 3700 8567
rect 2371 8419 2372 8427
rect 2374 8419 2377 8427
rect 2379 8419 2380 8427
rect 2392 8419 2393 8427
rect 2395 8423 2396 8427
rect 2395 8419 2400 8423
rect 2408 8419 2409 8427
rect 2411 8419 2414 8427
rect 2416 8419 2417 8427
rect 2434 8419 2435 8427
rect 2437 8419 2438 8427
rect 2450 8419 2451 8427
rect 2453 8423 2454 8427
rect 2453 8419 2458 8423
rect 2466 8419 2467 8427
rect 2469 8419 2472 8427
rect 2474 8419 2475 8427
rect 2487 8419 2488 8427
rect 2490 8419 2491 8427
rect 2503 8419 2504 8427
rect 2506 8419 2509 8427
rect 2511 8419 2512 8427
rect 2524 8419 2525 8427
rect 2527 8423 2528 8427
rect 2527 8419 2532 8423
rect 2540 8419 2541 8427
rect 2543 8419 2546 8427
rect 2548 8419 2549 8427
rect 2566 8419 2567 8427
rect 2569 8419 2570 8427
rect 2582 8419 2583 8427
rect 2585 8423 2586 8427
rect 2585 8419 2590 8423
rect 2598 8419 2599 8427
rect 2601 8419 2604 8427
rect 2606 8419 2607 8427
rect 2619 8419 2620 8427
rect 2622 8419 2623 8427
rect 2635 8419 2636 8427
rect 2638 8419 2641 8427
rect 2643 8419 2644 8427
rect 2656 8419 2657 8427
rect 2659 8423 2660 8427
rect 2659 8419 2664 8423
rect 2672 8419 2673 8427
rect 2675 8419 2678 8427
rect 2680 8419 2681 8427
rect 2698 8419 2699 8427
rect 2701 8419 2702 8427
rect 2714 8419 2715 8427
rect 2717 8423 2718 8427
rect 2717 8419 2722 8423
rect 2730 8419 2731 8427
rect 2733 8419 2736 8427
rect 2738 8419 2739 8427
rect 2751 8419 2752 8427
rect 2754 8419 2755 8427
rect 3316 8419 3317 8427
rect 3319 8419 3322 8427
rect 3324 8419 3325 8427
rect 3337 8419 3338 8427
rect 3340 8423 3341 8427
rect 3340 8419 3345 8423
rect 3353 8419 3354 8427
rect 3356 8419 3359 8427
rect 3361 8419 3362 8427
rect 3379 8419 3380 8427
rect 3382 8419 3383 8427
rect 3395 8419 3396 8427
rect 3398 8423 3399 8427
rect 3398 8419 3403 8423
rect 3411 8419 3412 8427
rect 3414 8419 3417 8427
rect 3419 8419 3420 8427
rect 3432 8419 3433 8427
rect 3435 8419 3436 8427
rect 3448 8419 3449 8427
rect 3451 8419 3454 8427
rect 3456 8419 3457 8427
rect 3469 8419 3470 8427
rect 3472 8423 3473 8427
rect 3472 8419 3477 8423
rect 3485 8419 3486 8427
rect 3488 8419 3491 8427
rect 3493 8419 3494 8427
rect 3511 8419 3512 8427
rect 3514 8419 3515 8427
rect 3527 8419 3528 8427
rect 3530 8423 3531 8427
rect 3530 8419 3535 8423
rect 3543 8419 3544 8427
rect 3546 8419 3549 8427
rect 3551 8419 3552 8427
rect 3564 8419 3565 8427
rect 3567 8419 3568 8427
rect 3580 8419 3581 8427
rect 3583 8419 3586 8427
rect 3588 8419 3589 8427
rect 3601 8419 3602 8427
rect 3604 8423 3605 8427
rect 3604 8419 3609 8423
rect 3617 8419 3618 8427
rect 3620 8419 3623 8427
rect 3625 8419 3626 8427
rect 3643 8419 3644 8427
rect 3646 8419 3647 8427
rect 3659 8419 3660 8427
rect 3662 8423 3663 8427
rect 3662 8419 3667 8423
rect 3675 8419 3676 8427
rect 3678 8419 3681 8427
rect 3683 8419 3684 8427
rect 3696 8419 3697 8427
rect 3699 8419 3700 8427
rect 2855 8340 2856 8348
rect 2858 8340 2861 8348
rect 2863 8340 2864 8348
rect 2876 8340 2877 8348
rect 2879 8344 2880 8348
rect 2879 8340 2884 8344
rect 2892 8340 2893 8348
rect 2895 8340 2898 8348
rect 2900 8340 2901 8348
rect 2918 8340 2919 8348
rect 2921 8340 2922 8348
rect 2934 8340 2935 8348
rect 2937 8344 2938 8348
rect 2937 8340 2942 8344
rect 2950 8340 2951 8348
rect 2953 8340 2956 8348
rect 2958 8340 2959 8348
rect 2971 8340 2972 8348
rect 2974 8340 2975 8348
rect 2987 8340 2988 8348
rect 2990 8340 2993 8348
rect 2995 8340 2996 8348
rect 3008 8340 3009 8348
rect 3011 8344 3012 8348
rect 3011 8340 3016 8344
rect 3024 8340 3025 8348
rect 3027 8340 3030 8348
rect 3032 8340 3033 8348
rect 3050 8340 3051 8348
rect 3053 8340 3054 8348
rect 3066 8340 3067 8348
rect 3069 8344 3070 8348
rect 3069 8340 3074 8344
rect 3082 8340 3083 8348
rect 3085 8340 3088 8348
rect 3090 8340 3091 8348
rect 3103 8340 3104 8348
rect 3106 8340 3107 8348
rect 3119 8340 3120 8348
rect 3122 8340 3125 8348
rect 3127 8340 3128 8348
rect 3140 8340 3141 8348
rect 3143 8344 3144 8348
rect 3143 8340 3148 8344
rect 3156 8340 3157 8348
rect 3159 8340 3162 8348
rect 3164 8340 3165 8348
rect 3182 8340 3183 8348
rect 3185 8340 3186 8348
rect 3198 8340 3199 8348
rect 3201 8344 3202 8348
rect 3201 8340 3206 8344
rect 3214 8340 3215 8348
rect 3217 8340 3220 8348
rect 3222 8340 3223 8348
rect 3235 8340 3236 8348
rect 3238 8340 3239 8348
rect 3251 8340 3252 8348
rect 3254 8340 3257 8348
rect 3259 8340 3260 8348
rect 3272 8340 3273 8348
rect 3275 8344 3276 8348
rect 3275 8340 3280 8344
rect 3288 8340 3289 8348
rect 3291 8340 3294 8348
rect 3296 8340 3297 8348
rect 3314 8340 3315 8348
rect 3317 8340 3318 8348
rect 3330 8340 3331 8348
rect 3333 8344 3334 8348
rect 3333 8340 3338 8344
rect 3346 8340 3347 8348
rect 3349 8340 3352 8348
rect 3354 8340 3355 8348
rect 3367 8340 3368 8348
rect 3370 8340 3371 8348
rect 3800 8340 3801 8348
rect 3803 8340 3806 8348
rect 3808 8340 3809 8348
rect 3821 8340 3822 8348
rect 3824 8344 3825 8348
rect 3824 8340 3829 8344
rect 3837 8340 3838 8348
rect 3840 8340 3843 8348
rect 3845 8340 3846 8348
rect 3863 8340 3864 8348
rect 3866 8340 3867 8348
rect 3879 8340 3880 8348
rect 3882 8344 3883 8348
rect 3882 8340 3887 8344
rect 3895 8340 3896 8348
rect 3898 8340 3901 8348
rect 3903 8340 3904 8348
rect 3916 8340 3917 8348
rect 3919 8340 3920 8348
rect 3932 8340 3933 8348
rect 3935 8340 3938 8348
rect 3940 8340 3941 8348
rect 3953 8340 3954 8348
rect 3956 8344 3957 8348
rect 3956 8340 3961 8344
rect 3969 8340 3970 8348
rect 3972 8340 3975 8348
rect 3977 8340 3978 8348
rect 3995 8340 3996 8348
rect 3998 8340 3999 8348
rect 4011 8340 4012 8348
rect 4014 8344 4015 8348
rect 4014 8340 4019 8344
rect 4027 8340 4028 8348
rect 4030 8340 4033 8348
rect 4035 8340 4036 8348
rect 4048 8340 4049 8348
rect 4051 8340 4052 8348
rect 4064 8340 4065 8348
rect 4067 8340 4070 8348
rect 4072 8340 4073 8348
rect 4085 8340 4086 8348
rect 4088 8344 4089 8348
rect 4088 8340 4093 8344
rect 4101 8340 4102 8348
rect 4104 8340 4107 8348
rect 4109 8340 4110 8348
rect 4127 8340 4128 8348
rect 4130 8340 4131 8348
rect 4143 8340 4144 8348
rect 4146 8344 4147 8348
rect 4146 8340 4151 8344
rect 4159 8340 4160 8348
rect 4162 8340 4165 8348
rect 4167 8340 4168 8348
rect 4180 8340 4181 8348
rect 4183 8340 4184 8348
rect 4196 8340 4197 8348
rect 4199 8340 4202 8348
rect 4204 8340 4205 8348
rect 4217 8340 4218 8348
rect 4220 8344 4221 8348
rect 4220 8340 4225 8344
rect 4233 8340 4234 8348
rect 4236 8340 4239 8348
rect 4241 8340 4242 8348
rect 4259 8340 4260 8348
rect 4262 8340 4263 8348
rect 4275 8340 4276 8348
rect 4278 8344 4279 8348
rect 4278 8340 4283 8344
rect 4291 8340 4292 8348
rect 4294 8340 4297 8348
rect 4299 8340 4300 8348
rect 4312 8340 4313 8348
rect 4315 8340 4316 8348
rect 2503 8307 2504 8315
rect 2506 8307 2509 8315
rect 2511 8307 2512 8315
rect 2524 8307 2525 8315
rect 2527 8311 2528 8315
rect 2527 8307 2532 8311
rect 2540 8307 2541 8315
rect 2543 8307 2546 8315
rect 2548 8307 2549 8315
rect 2566 8307 2567 8315
rect 2569 8307 2570 8315
rect 2582 8307 2583 8315
rect 2585 8311 2586 8315
rect 2585 8307 2590 8311
rect 2598 8307 2599 8315
rect 2601 8307 2604 8315
rect 2606 8307 2607 8315
rect 2619 8307 2620 8315
rect 2622 8307 2623 8315
rect 3448 8307 3449 8315
rect 3451 8307 3454 8315
rect 3456 8307 3457 8315
rect 3469 8307 3470 8315
rect 3472 8311 3473 8315
rect 3472 8307 3477 8311
rect 3485 8307 3486 8315
rect 3488 8307 3491 8315
rect 3493 8307 3494 8315
rect 3511 8307 3512 8315
rect 3514 8307 3515 8315
rect 3527 8307 3528 8315
rect 3530 8311 3531 8315
rect 3530 8307 3535 8311
rect 3543 8307 3544 8315
rect 3546 8307 3549 8315
rect 3551 8307 3552 8315
rect 3564 8307 3565 8315
rect 3567 8307 3568 8315
rect 3034 8269 3035 8277
rect 3037 8269 3038 8277
rect 2860 8256 2861 8264
rect 2863 8256 2864 8264
rect 2876 8256 2877 8264
rect 2879 8256 2880 8264
rect 2892 8256 2893 8264
rect 2895 8256 2896 8264
rect 2911 8256 2916 8264
rect 2918 8256 2921 8264
rect 2923 8256 2924 8264
rect 2945 8256 2947 8264
rect 2949 8256 2950 8264
rect 2967 8256 2968 8264
rect 2970 8256 2971 8264
rect 2983 8256 2988 8264
rect 2990 8256 2993 8264
rect 2995 8256 2996 8264
rect 3010 8256 3011 8264
rect 3013 8256 3014 8264
rect 3058 8263 3061 8271
rect 3063 8263 3066 8271
rect 3068 8263 3069 8271
rect 3088 8269 3089 8277
rect 3091 8269 3092 8277
rect 3115 8269 3116 8277
rect 3118 8269 3119 8277
rect 3139 8263 3142 8271
rect 3144 8263 3147 8271
rect 3149 8263 3150 8271
rect 3169 8269 3170 8277
rect 3172 8269 3173 8277
rect 3979 8269 3980 8277
rect 3982 8269 3983 8277
rect 3805 8256 3806 8264
rect 3808 8256 3809 8264
rect 3821 8256 3822 8264
rect 3824 8256 3825 8264
rect 3837 8256 3838 8264
rect 3840 8256 3841 8264
rect 3856 8256 3861 8264
rect 3863 8256 3866 8264
rect 3868 8256 3869 8264
rect 3890 8256 3892 8264
rect 3894 8256 3895 8264
rect 3912 8256 3913 8264
rect 3915 8256 3916 8264
rect 3928 8256 3933 8264
rect 3935 8256 3938 8264
rect 3940 8256 3941 8264
rect 3955 8256 3956 8264
rect 3958 8256 3959 8264
rect 4003 8263 4006 8271
rect 4008 8263 4011 8271
rect 4013 8263 4014 8271
rect 4033 8269 4034 8277
rect 4036 8269 4037 8277
rect 4060 8269 4061 8277
rect 4063 8269 4064 8277
rect 4084 8263 4087 8271
rect 4089 8263 4092 8271
rect 4094 8263 4095 8271
rect 4114 8269 4115 8277
rect 4117 8269 4118 8277
rect 2494 8205 2495 8213
rect 2497 8205 2498 8213
rect 2510 8205 2511 8213
rect 2513 8205 2516 8213
rect 2518 8205 2519 8213
rect 2531 8209 2532 8213
rect 2527 8205 2532 8209
rect 2534 8205 2535 8213
rect 2547 8205 2548 8213
rect 2550 8205 2551 8213
rect 2568 8205 2569 8213
rect 2571 8205 2574 8213
rect 2576 8205 2577 8213
rect 2589 8209 2590 8213
rect 2585 8205 2590 8209
rect 2592 8205 2593 8213
rect 2605 8205 2606 8213
rect 2608 8205 2611 8213
rect 2613 8205 2614 8213
rect 3439 8205 3440 8213
rect 3442 8205 3443 8213
rect 3455 8205 3456 8213
rect 3458 8205 3461 8213
rect 3463 8205 3464 8213
rect 3476 8209 3477 8213
rect 3472 8205 3477 8209
rect 3479 8205 3480 8213
rect 3492 8205 3493 8213
rect 3495 8205 3496 8213
rect 3513 8205 3514 8213
rect 3516 8205 3519 8213
rect 3521 8205 3522 8213
rect 3534 8209 3535 8213
rect 3530 8205 3535 8209
rect 3537 8205 3538 8213
rect 3550 8205 3551 8213
rect 3553 8205 3556 8213
rect 3558 8205 3559 8213
rect 2860 8170 2861 8178
rect 2863 8170 2864 8178
rect 2876 8170 2877 8178
rect 2879 8170 2880 8178
rect 2892 8170 2893 8178
rect 2895 8170 2896 8178
rect 2911 8170 2916 8178
rect 2918 8170 2921 8178
rect 2923 8170 2924 8178
rect 2945 8170 2947 8178
rect 2949 8170 2950 8178
rect 2967 8170 2968 8178
rect 2970 8170 2971 8178
rect 2983 8170 2988 8178
rect 2990 8170 2993 8178
rect 2995 8170 2996 8178
rect 3010 8170 3011 8178
rect 3013 8170 3014 8178
rect 3058 8171 3061 8179
rect 3063 8171 3066 8179
rect 3068 8171 3069 8179
rect 3139 8171 3142 8179
rect 3144 8171 3147 8179
rect 3149 8171 3150 8179
rect 3805 8170 3806 8178
rect 3808 8170 3809 8178
rect 3821 8170 3822 8178
rect 3824 8170 3825 8178
rect 3837 8170 3838 8178
rect 3840 8170 3841 8178
rect 3856 8170 3861 8178
rect 3863 8170 3866 8178
rect 3868 8170 3869 8178
rect 3890 8170 3892 8178
rect 3894 8170 3895 8178
rect 3912 8170 3913 8178
rect 3915 8170 3916 8178
rect 3928 8170 3933 8178
rect 3935 8170 3938 8178
rect 3940 8170 3941 8178
rect 3955 8170 3956 8178
rect 3958 8170 3959 8178
rect 4003 8171 4006 8179
rect 4008 8171 4011 8179
rect 4013 8171 4014 8179
rect 4084 8171 4087 8179
rect 4089 8171 4092 8179
rect 4094 8171 4095 8179
rect 2860 8124 2861 8132
rect 2863 8124 2864 8132
rect 2876 8124 2877 8132
rect 2879 8124 2880 8132
rect 2892 8124 2893 8132
rect 2895 8124 2896 8132
rect 2911 8124 2916 8132
rect 2918 8124 2921 8132
rect 2923 8124 2924 8132
rect 2945 8124 2947 8132
rect 2949 8124 2950 8132
rect 2967 8124 2968 8132
rect 2970 8124 2971 8132
rect 2983 8124 2988 8132
rect 2990 8124 2993 8132
rect 2995 8124 2996 8132
rect 3010 8124 3011 8132
rect 3013 8124 3014 8132
rect 3058 8131 3061 8139
rect 3063 8131 3066 8139
rect 3068 8131 3069 8139
rect 3088 8137 3089 8145
rect 3091 8137 3092 8145
rect 3139 8137 3140 8145
rect 3142 8137 3143 8145
rect 3163 8131 3166 8139
rect 3168 8131 3171 8139
rect 3173 8131 3174 8139
rect 3193 8137 3194 8145
rect 3196 8137 3197 8145
rect 3805 8124 3806 8132
rect 3808 8124 3809 8132
rect 3821 8124 3822 8132
rect 3824 8124 3825 8132
rect 3837 8124 3838 8132
rect 3840 8124 3841 8132
rect 3856 8124 3861 8132
rect 3863 8124 3866 8132
rect 3868 8124 3869 8132
rect 3890 8124 3892 8132
rect 3894 8124 3895 8132
rect 3912 8124 3913 8132
rect 3915 8124 3916 8132
rect 3928 8124 3933 8132
rect 3935 8124 3938 8132
rect 3940 8124 3941 8132
rect 3955 8124 3956 8132
rect 3958 8124 3959 8132
rect 4003 8131 4006 8139
rect 4008 8131 4011 8139
rect 4013 8131 4014 8139
rect 4033 8137 4034 8145
rect 4036 8137 4037 8145
rect 4084 8137 4085 8145
rect 4087 8137 4088 8145
rect 4108 8131 4111 8139
rect 4113 8131 4116 8139
rect 4118 8131 4119 8139
rect 4138 8137 4139 8145
rect 4141 8137 4142 8145
rect 2860 8038 2861 8046
rect 2863 8038 2864 8046
rect 2876 8038 2877 8046
rect 2879 8038 2880 8046
rect 2892 8038 2893 8046
rect 2895 8038 2896 8046
rect 2911 8038 2916 8046
rect 2918 8038 2921 8046
rect 2923 8038 2924 8046
rect 2945 8038 2947 8046
rect 2949 8038 2950 8046
rect 2967 8038 2968 8046
rect 2970 8038 2971 8046
rect 2983 8038 2988 8046
rect 2990 8038 2993 8046
rect 2995 8038 2996 8046
rect 3010 8038 3011 8046
rect 3013 8038 3014 8046
rect 3058 8040 3061 8048
rect 3063 8040 3066 8048
rect 3068 8040 3069 8048
rect 3163 8040 3166 8048
rect 3168 8040 3171 8048
rect 3173 8040 3174 8048
rect 3805 8038 3806 8046
rect 3808 8038 3809 8046
rect 3821 8038 3822 8046
rect 3824 8038 3825 8046
rect 3837 8038 3838 8046
rect 3840 8038 3841 8046
rect 3856 8038 3861 8046
rect 3863 8038 3866 8046
rect 3868 8038 3869 8046
rect 3890 8038 3892 8046
rect 3894 8038 3895 8046
rect 3912 8038 3913 8046
rect 3915 8038 3916 8046
rect 3928 8038 3933 8046
rect 3935 8038 3938 8046
rect 3940 8038 3941 8046
rect 3955 8038 3956 8046
rect 3958 8038 3959 8046
rect 4003 8040 4006 8048
rect 4008 8040 4011 8048
rect 4013 8040 4014 8048
rect 4108 8040 4111 8048
rect 4113 8040 4116 8048
rect 4118 8040 4119 8048
rect 2860 7992 2861 8000
rect 2863 7992 2864 8000
rect 2876 7992 2877 8000
rect 2879 7992 2880 8000
rect 2892 7992 2893 8000
rect 2895 7992 2896 8000
rect 2911 7992 2916 8000
rect 2918 7992 2921 8000
rect 2923 7992 2924 8000
rect 2945 7992 2947 8000
rect 2949 7992 2950 8000
rect 2967 7992 2968 8000
rect 2970 7992 2971 8000
rect 2983 7992 2988 8000
rect 2990 7992 2993 8000
rect 2995 7992 2996 8000
rect 3010 7992 3011 8000
rect 3013 7992 3014 8000
rect 3058 7999 3061 8007
rect 3063 7999 3066 8007
rect 3068 7999 3069 8007
rect 3088 8005 3089 8013
rect 3091 8005 3092 8013
rect 3115 8005 3116 8013
rect 3118 8005 3119 8013
rect 3139 7999 3142 8007
rect 3144 7999 3147 8007
rect 3149 7999 3150 8007
rect 3169 8005 3170 8013
rect 3172 8005 3173 8013
rect 3205 8005 3206 8013
rect 3208 8005 3209 8013
rect 3229 7999 3232 8007
rect 3234 7999 3237 8007
rect 3239 7999 3240 8007
rect 3259 8005 3260 8013
rect 3262 8005 3263 8013
rect 3805 7992 3806 8000
rect 3808 7992 3809 8000
rect 3821 7992 3822 8000
rect 3824 7992 3825 8000
rect 3837 7992 3838 8000
rect 3840 7992 3841 8000
rect 3856 7992 3861 8000
rect 3863 7992 3866 8000
rect 3868 7992 3869 8000
rect 3890 7992 3892 8000
rect 3894 7992 3895 8000
rect 3912 7992 3913 8000
rect 3915 7992 3916 8000
rect 3928 7992 3933 8000
rect 3935 7992 3938 8000
rect 3940 7992 3941 8000
rect 3955 7992 3956 8000
rect 3958 7992 3959 8000
rect 4003 7999 4006 8007
rect 4008 7999 4011 8007
rect 4013 7999 4014 8007
rect 4033 8005 4034 8013
rect 4036 8005 4037 8013
rect 4060 8005 4061 8013
rect 4063 8005 4064 8013
rect 4084 7999 4087 8007
rect 4089 7999 4092 8007
rect 4094 7999 4095 8007
rect 4114 8005 4115 8013
rect 4117 8005 4118 8013
rect 4150 8005 4151 8013
rect 4153 8005 4154 8013
rect 4174 7999 4177 8007
rect 4179 7999 4182 8007
rect 4184 7999 4185 8007
rect 4204 8005 4205 8013
rect 4207 8005 4208 8013
rect 2860 7906 2861 7914
rect 2863 7906 2864 7914
rect 2876 7906 2877 7914
rect 2879 7906 2880 7914
rect 2892 7906 2893 7914
rect 2895 7906 2896 7914
rect 2911 7906 2916 7914
rect 2918 7906 2921 7914
rect 2923 7906 2924 7914
rect 2945 7906 2947 7914
rect 2949 7906 2950 7914
rect 2967 7906 2968 7914
rect 2970 7906 2971 7914
rect 2983 7906 2988 7914
rect 2990 7906 2993 7914
rect 2995 7906 2996 7914
rect 3010 7906 3011 7914
rect 3013 7906 3014 7914
rect 3058 7905 3061 7913
rect 3063 7905 3066 7913
rect 3068 7905 3069 7913
rect 3139 7905 3142 7913
rect 3144 7905 3147 7913
rect 3149 7905 3150 7913
rect 3229 7905 3232 7913
rect 3234 7905 3237 7913
rect 3239 7905 3240 7913
rect 3805 7906 3806 7914
rect 3808 7906 3809 7914
rect 3821 7906 3822 7914
rect 3824 7906 3825 7914
rect 3837 7906 3838 7914
rect 3840 7906 3841 7914
rect 3856 7906 3861 7914
rect 3863 7906 3866 7914
rect 3868 7906 3869 7914
rect 3890 7906 3892 7914
rect 3894 7906 3895 7914
rect 3912 7906 3913 7914
rect 3915 7906 3916 7914
rect 3928 7906 3933 7914
rect 3935 7906 3938 7914
rect 3940 7906 3941 7914
rect 3955 7906 3956 7914
rect 3958 7906 3959 7914
rect 4003 7905 4006 7913
rect 4008 7905 4011 7913
rect 4013 7905 4014 7913
rect 4084 7905 4087 7913
rect 4089 7905 4092 7913
rect 4094 7905 4095 7913
rect 4174 7905 4177 7913
rect 4179 7905 4182 7913
rect 4184 7905 4185 7913
rect 2860 7860 2861 7868
rect 2863 7860 2864 7868
rect 2876 7860 2877 7868
rect 2879 7860 2880 7868
rect 2892 7860 2893 7868
rect 2895 7860 2896 7868
rect 2911 7860 2916 7868
rect 2918 7860 2921 7868
rect 2923 7860 2924 7868
rect 2945 7860 2947 7868
rect 2949 7860 2950 7868
rect 2967 7860 2968 7868
rect 2970 7860 2971 7868
rect 2983 7860 2988 7868
rect 2990 7860 2993 7868
rect 2995 7860 2996 7868
rect 3010 7860 3011 7868
rect 3013 7860 3014 7868
rect 3058 7867 3061 7875
rect 3063 7867 3066 7875
rect 3068 7867 3069 7875
rect 3088 7873 3089 7881
rect 3091 7873 3092 7881
rect 3805 7860 3806 7868
rect 3808 7860 3809 7868
rect 3821 7860 3822 7868
rect 3824 7860 3825 7868
rect 3837 7860 3838 7868
rect 3840 7860 3841 7868
rect 3856 7860 3861 7868
rect 3863 7860 3866 7868
rect 3868 7860 3869 7868
rect 3890 7860 3892 7868
rect 3894 7860 3895 7868
rect 3912 7860 3913 7868
rect 3915 7860 3916 7868
rect 3928 7860 3933 7868
rect 3935 7860 3938 7868
rect 3940 7860 3941 7868
rect 3955 7860 3956 7868
rect 3958 7860 3959 7868
rect 4003 7867 4006 7875
rect 4008 7867 4011 7875
rect 4013 7867 4014 7875
rect 4033 7873 4034 7881
rect 4036 7873 4037 7881
rect 2371 7805 2372 7813
rect 2374 7805 2377 7813
rect 2379 7805 2380 7813
rect 2392 7805 2393 7813
rect 2395 7809 2396 7813
rect 2395 7805 2400 7809
rect 2408 7805 2409 7813
rect 2411 7805 2414 7813
rect 2416 7805 2417 7813
rect 2434 7805 2435 7813
rect 2437 7805 2438 7813
rect 2450 7805 2451 7813
rect 2453 7809 2454 7813
rect 2453 7805 2458 7809
rect 2466 7805 2467 7813
rect 2469 7805 2472 7813
rect 2474 7805 2475 7813
rect 2487 7805 2488 7813
rect 2490 7805 2491 7813
rect 2503 7805 2504 7813
rect 2506 7805 2509 7813
rect 2511 7805 2512 7813
rect 2524 7805 2525 7813
rect 2527 7809 2528 7813
rect 2527 7805 2532 7809
rect 2540 7805 2541 7813
rect 2543 7805 2546 7813
rect 2548 7805 2549 7813
rect 2566 7805 2567 7813
rect 2569 7805 2570 7813
rect 2582 7805 2583 7813
rect 2585 7809 2586 7813
rect 2585 7805 2590 7809
rect 2598 7805 2599 7813
rect 2601 7805 2604 7813
rect 2606 7805 2607 7813
rect 2619 7805 2620 7813
rect 2622 7805 2623 7813
rect 2635 7805 2636 7813
rect 2638 7805 2641 7813
rect 2643 7805 2644 7813
rect 2656 7805 2657 7813
rect 2659 7809 2660 7813
rect 2659 7805 2664 7809
rect 2672 7805 2673 7813
rect 2675 7805 2678 7813
rect 2680 7805 2681 7813
rect 2698 7805 2699 7813
rect 2701 7805 2702 7813
rect 2714 7805 2715 7813
rect 2717 7809 2718 7813
rect 2717 7805 2722 7809
rect 2730 7805 2731 7813
rect 2733 7805 2736 7813
rect 2738 7805 2739 7813
rect 2751 7805 2752 7813
rect 2754 7805 2755 7813
rect 3316 7805 3317 7813
rect 3319 7805 3322 7813
rect 3324 7805 3325 7813
rect 3337 7805 3338 7813
rect 3340 7809 3341 7813
rect 3340 7805 3345 7809
rect 3353 7805 3354 7813
rect 3356 7805 3359 7813
rect 3361 7805 3362 7813
rect 3379 7805 3380 7813
rect 3382 7805 3383 7813
rect 3395 7805 3396 7813
rect 3398 7809 3399 7813
rect 3398 7805 3403 7809
rect 3411 7805 3412 7813
rect 3414 7805 3417 7813
rect 3419 7805 3420 7813
rect 3432 7805 3433 7813
rect 3435 7805 3436 7813
rect 3448 7805 3449 7813
rect 3451 7805 3454 7813
rect 3456 7805 3457 7813
rect 3469 7805 3470 7813
rect 3472 7809 3473 7813
rect 3472 7805 3477 7809
rect 3485 7805 3486 7813
rect 3488 7805 3491 7813
rect 3493 7805 3494 7813
rect 3511 7805 3512 7813
rect 3514 7805 3515 7813
rect 3527 7805 3528 7813
rect 3530 7809 3531 7813
rect 3530 7805 3535 7809
rect 3543 7805 3544 7813
rect 3546 7805 3549 7813
rect 3551 7805 3552 7813
rect 3564 7805 3565 7813
rect 3567 7805 3568 7813
rect 3580 7805 3581 7813
rect 3583 7805 3586 7813
rect 3588 7805 3589 7813
rect 3601 7805 3602 7813
rect 3604 7809 3605 7813
rect 3604 7805 3609 7809
rect 3617 7805 3618 7813
rect 3620 7805 3623 7813
rect 3625 7805 3626 7813
rect 3643 7805 3644 7813
rect 3646 7805 3647 7813
rect 3659 7805 3660 7813
rect 3662 7809 3663 7813
rect 3662 7805 3667 7809
rect 3675 7805 3676 7813
rect 3678 7805 3681 7813
rect 3683 7805 3684 7813
rect 3696 7805 3697 7813
rect 3699 7805 3700 7813
rect 2860 7774 2861 7782
rect 2863 7774 2864 7782
rect 2876 7774 2877 7782
rect 2879 7774 2880 7782
rect 2892 7774 2893 7782
rect 2895 7774 2896 7782
rect 2911 7774 2916 7782
rect 2918 7774 2921 7782
rect 2923 7774 2924 7782
rect 2945 7774 2947 7782
rect 2949 7774 2950 7782
rect 2967 7774 2968 7782
rect 2970 7774 2971 7782
rect 2983 7774 2988 7782
rect 2990 7774 2993 7782
rect 2995 7774 2996 7782
rect 3010 7774 3011 7782
rect 3013 7774 3014 7782
rect 3058 7769 3061 7777
rect 3063 7769 3066 7777
rect 3068 7769 3069 7777
rect 3094 7774 3095 7782
rect 3097 7774 3098 7782
rect 3102 7774 3108 7782
rect 3112 7774 3113 7782
rect 3115 7774 3116 7782
rect 3137 7774 3138 7782
rect 3140 7774 3141 7782
rect 3153 7774 3154 7782
rect 3156 7774 3157 7782
rect 3172 7774 3177 7782
rect 3179 7774 3182 7782
rect 3184 7774 3185 7782
rect 3206 7774 3208 7782
rect 3210 7774 3211 7782
rect 3228 7774 3229 7782
rect 3231 7774 3232 7782
rect 3244 7774 3249 7782
rect 3251 7774 3254 7782
rect 3256 7774 3257 7782
rect 3271 7774 3272 7782
rect 3274 7774 3275 7782
rect 3805 7774 3806 7782
rect 3808 7774 3809 7782
rect 3821 7774 3822 7782
rect 3824 7774 3825 7782
rect 3837 7774 3838 7782
rect 3840 7774 3841 7782
rect 3856 7774 3861 7782
rect 3863 7774 3866 7782
rect 3868 7774 3869 7782
rect 3890 7774 3892 7782
rect 3894 7774 3895 7782
rect 3912 7774 3913 7782
rect 3915 7774 3916 7782
rect 3928 7774 3933 7782
rect 3935 7774 3938 7782
rect 3940 7774 3941 7782
rect 3955 7774 3956 7782
rect 3958 7774 3959 7782
rect 4003 7769 4006 7777
rect 4008 7769 4011 7777
rect 4013 7769 4014 7777
rect 4039 7774 4040 7782
rect 4042 7774 4043 7782
rect 4047 7774 4053 7782
rect 4057 7774 4058 7782
rect 4060 7774 4061 7782
rect 4082 7774 4083 7782
rect 4085 7774 4086 7782
rect 4098 7774 4099 7782
rect 4101 7774 4102 7782
rect 4117 7774 4122 7782
rect 4124 7774 4127 7782
rect 4129 7774 4130 7782
rect 4151 7774 4153 7782
rect 4155 7774 4156 7782
rect 4173 7774 4174 7782
rect 4176 7774 4177 7782
rect 4189 7774 4194 7782
rect 4196 7774 4199 7782
rect 4201 7774 4202 7782
rect 4216 7774 4217 7782
rect 4219 7774 4220 7782
rect 3154 7693 3155 7701
rect 3157 7693 3160 7701
rect 3162 7693 3163 7701
rect 3175 7693 3176 7701
rect 3178 7697 3179 7701
rect 3178 7693 3183 7697
rect 3191 7693 3192 7701
rect 3194 7693 3197 7701
rect 3199 7693 3200 7701
rect 3217 7693 3218 7701
rect 3220 7693 3221 7701
rect 3233 7693 3234 7701
rect 3236 7697 3237 7701
rect 3236 7693 3241 7697
rect 3249 7693 3250 7701
rect 3252 7693 3255 7701
rect 3257 7693 3258 7701
rect 3270 7693 3271 7701
rect 3273 7693 3274 7701
rect 4099 7693 4100 7701
rect 4102 7693 4105 7701
rect 4107 7693 4108 7701
rect 4120 7693 4121 7701
rect 4123 7697 4124 7701
rect 4123 7693 4128 7697
rect 4136 7693 4137 7701
rect 4139 7693 4142 7701
rect 4144 7693 4145 7701
rect 4162 7693 4163 7701
rect 4165 7693 4166 7701
rect 4178 7693 4179 7701
rect 4181 7697 4182 7701
rect 4181 7693 4186 7697
rect 4194 7693 4195 7701
rect 4197 7693 4200 7701
rect 4202 7693 4203 7701
rect 4215 7693 4216 7701
rect 4218 7693 4219 7701
rect 2371 7663 2372 7671
rect 2374 7663 2377 7671
rect 2379 7663 2380 7671
rect 2392 7663 2393 7671
rect 2395 7667 2396 7671
rect 2395 7663 2400 7667
rect 2408 7663 2409 7671
rect 2411 7663 2414 7671
rect 2416 7663 2417 7671
rect 2434 7663 2435 7671
rect 2437 7663 2438 7671
rect 2450 7663 2451 7671
rect 2453 7667 2454 7671
rect 2453 7663 2458 7667
rect 2466 7663 2467 7671
rect 2469 7663 2472 7671
rect 2474 7663 2475 7671
rect 2487 7663 2488 7671
rect 2490 7663 2491 7671
rect 2503 7663 2504 7671
rect 2506 7663 2509 7671
rect 2511 7663 2512 7671
rect 2524 7663 2525 7671
rect 2527 7667 2528 7671
rect 2527 7663 2532 7667
rect 2540 7663 2541 7671
rect 2543 7663 2546 7671
rect 2548 7663 2549 7671
rect 2566 7663 2567 7671
rect 2569 7663 2570 7671
rect 2582 7663 2583 7671
rect 2585 7667 2586 7671
rect 2585 7663 2590 7667
rect 2598 7663 2599 7671
rect 2601 7663 2604 7671
rect 2606 7663 2607 7671
rect 2619 7663 2620 7671
rect 2622 7663 2623 7671
rect 2635 7663 2636 7671
rect 2638 7663 2641 7671
rect 2643 7663 2644 7671
rect 2656 7663 2657 7671
rect 2659 7667 2660 7671
rect 2659 7663 2664 7667
rect 2672 7663 2673 7671
rect 2675 7663 2678 7671
rect 2680 7663 2681 7671
rect 2698 7663 2699 7671
rect 2701 7663 2702 7671
rect 2714 7663 2715 7671
rect 2717 7667 2718 7671
rect 2717 7663 2722 7667
rect 2730 7663 2731 7671
rect 2733 7663 2736 7671
rect 2738 7663 2739 7671
rect 2751 7663 2752 7671
rect 2754 7663 2755 7671
rect 3316 7663 3317 7671
rect 3319 7663 3322 7671
rect 3324 7663 3325 7671
rect 3337 7663 3338 7671
rect 3340 7667 3341 7671
rect 3340 7663 3345 7667
rect 3353 7663 3354 7671
rect 3356 7663 3359 7671
rect 3361 7663 3362 7671
rect 3379 7663 3380 7671
rect 3382 7663 3383 7671
rect 3395 7663 3396 7671
rect 3398 7667 3399 7671
rect 3398 7663 3403 7667
rect 3411 7663 3412 7671
rect 3414 7663 3417 7671
rect 3419 7663 3420 7671
rect 3432 7663 3433 7671
rect 3435 7663 3436 7671
rect 3448 7663 3449 7671
rect 3451 7663 3454 7671
rect 3456 7663 3457 7671
rect 3469 7663 3470 7671
rect 3472 7667 3473 7671
rect 3472 7663 3477 7667
rect 3485 7663 3486 7671
rect 3488 7663 3491 7671
rect 3493 7663 3494 7671
rect 3511 7663 3512 7671
rect 3514 7663 3515 7671
rect 3527 7663 3528 7671
rect 3530 7667 3531 7671
rect 3530 7663 3535 7667
rect 3543 7663 3544 7671
rect 3546 7663 3549 7671
rect 3551 7663 3552 7671
rect 3564 7663 3565 7671
rect 3567 7663 3568 7671
rect 3580 7663 3581 7671
rect 3583 7663 3586 7671
rect 3588 7663 3589 7671
rect 3601 7663 3602 7671
rect 3604 7667 3605 7671
rect 3604 7663 3609 7667
rect 3617 7663 3618 7671
rect 3620 7663 3623 7671
rect 3625 7663 3626 7671
rect 3643 7663 3644 7671
rect 3646 7663 3647 7671
rect 3659 7663 3660 7671
rect 3662 7667 3663 7671
rect 3662 7663 3667 7667
rect 3675 7663 3676 7671
rect 3678 7663 3681 7671
rect 3683 7663 3684 7671
rect 3696 7663 3697 7671
rect 3699 7663 3700 7671
rect 3154 7607 3155 7615
rect 3157 7607 3160 7615
rect 3162 7607 3163 7615
rect 3175 7607 3176 7615
rect 3178 7611 3179 7615
rect 3178 7607 3183 7611
rect 3191 7607 3192 7615
rect 3194 7607 3197 7615
rect 3199 7607 3200 7615
rect 3217 7607 3218 7615
rect 3220 7607 3221 7615
rect 3233 7607 3234 7615
rect 3236 7611 3237 7615
rect 3236 7607 3241 7611
rect 3249 7607 3250 7615
rect 3252 7607 3255 7615
rect 3257 7607 3258 7615
rect 3270 7607 3271 7615
rect 3273 7607 3274 7615
rect 4099 7607 4100 7615
rect 4102 7607 4105 7615
rect 4107 7607 4108 7615
rect 4120 7607 4121 7615
rect 4123 7611 4124 7615
rect 4123 7607 4128 7611
rect 4136 7607 4137 7615
rect 4139 7607 4142 7615
rect 4144 7607 4145 7615
rect 4162 7607 4163 7615
rect 4165 7607 4166 7615
rect 4178 7607 4179 7615
rect 4181 7611 4182 7615
rect 4181 7607 4186 7611
rect 4194 7607 4195 7615
rect 4197 7607 4200 7615
rect 4202 7607 4203 7615
rect 4215 7607 4216 7615
rect 4218 7607 4219 7615
rect 2371 7577 2372 7585
rect 2374 7577 2377 7585
rect 2379 7577 2380 7585
rect 2392 7577 2393 7585
rect 2395 7581 2396 7585
rect 2395 7577 2400 7581
rect 2408 7577 2409 7585
rect 2411 7577 2414 7585
rect 2416 7577 2417 7585
rect 2434 7577 2435 7585
rect 2437 7577 2438 7585
rect 2450 7577 2451 7585
rect 2453 7581 2454 7585
rect 2453 7577 2458 7581
rect 2466 7577 2467 7585
rect 2469 7577 2472 7585
rect 2474 7577 2475 7585
rect 2487 7577 2488 7585
rect 2490 7577 2491 7585
rect 2503 7577 2504 7585
rect 2506 7577 2509 7585
rect 2511 7577 2512 7585
rect 2524 7577 2525 7585
rect 2527 7581 2528 7585
rect 2527 7577 2532 7581
rect 2540 7577 2541 7585
rect 2543 7577 2546 7585
rect 2548 7577 2549 7585
rect 2566 7577 2567 7585
rect 2569 7577 2570 7585
rect 2582 7577 2583 7585
rect 2585 7581 2586 7585
rect 2585 7577 2590 7581
rect 2598 7577 2599 7585
rect 2601 7577 2604 7585
rect 2606 7577 2607 7585
rect 2619 7577 2620 7585
rect 2622 7577 2623 7585
rect 2635 7577 2636 7585
rect 2638 7577 2641 7585
rect 2643 7577 2644 7585
rect 2656 7577 2657 7585
rect 2659 7581 2660 7585
rect 2659 7577 2664 7581
rect 2672 7577 2673 7585
rect 2675 7577 2678 7585
rect 2680 7577 2681 7585
rect 2698 7577 2699 7585
rect 2701 7577 2702 7585
rect 2714 7577 2715 7585
rect 2717 7581 2718 7585
rect 2717 7577 2722 7581
rect 2730 7577 2731 7585
rect 2733 7577 2736 7585
rect 2738 7577 2739 7585
rect 2751 7577 2752 7585
rect 2754 7577 2755 7585
rect 3316 7577 3317 7585
rect 3319 7577 3322 7585
rect 3324 7577 3325 7585
rect 3337 7577 3338 7585
rect 3340 7581 3341 7585
rect 3340 7577 3345 7581
rect 3353 7577 3354 7585
rect 3356 7577 3359 7585
rect 3361 7577 3362 7585
rect 3379 7577 3380 7585
rect 3382 7577 3383 7585
rect 3395 7577 3396 7585
rect 3398 7581 3399 7585
rect 3398 7577 3403 7581
rect 3411 7577 3412 7585
rect 3414 7577 3417 7585
rect 3419 7577 3420 7585
rect 3432 7577 3433 7585
rect 3435 7577 3436 7585
rect 3448 7577 3449 7585
rect 3451 7577 3454 7585
rect 3456 7577 3457 7585
rect 3469 7577 3470 7585
rect 3472 7581 3473 7585
rect 3472 7577 3477 7581
rect 3485 7577 3486 7585
rect 3488 7577 3491 7585
rect 3493 7577 3494 7585
rect 3511 7577 3512 7585
rect 3514 7577 3515 7585
rect 3527 7577 3528 7585
rect 3530 7581 3531 7585
rect 3530 7577 3535 7581
rect 3543 7577 3544 7585
rect 3546 7577 3549 7585
rect 3551 7577 3552 7585
rect 3564 7577 3565 7585
rect 3567 7577 3568 7585
rect 3580 7577 3581 7585
rect 3583 7577 3586 7585
rect 3588 7577 3589 7585
rect 3601 7577 3602 7585
rect 3604 7581 3605 7585
rect 3604 7577 3609 7581
rect 3617 7577 3618 7585
rect 3620 7577 3623 7585
rect 3625 7577 3626 7585
rect 3643 7577 3644 7585
rect 3646 7577 3647 7585
rect 3659 7577 3660 7585
rect 3662 7581 3663 7585
rect 3662 7577 3667 7581
rect 3675 7577 3676 7585
rect 3678 7577 3681 7585
rect 3683 7577 3684 7585
rect 3696 7577 3697 7585
rect 3699 7577 3700 7585
rect 2371 7437 2372 7445
rect 2374 7437 2377 7445
rect 2379 7437 2380 7445
rect 2392 7437 2393 7445
rect 2395 7441 2396 7445
rect 2395 7437 2400 7441
rect 2408 7437 2409 7445
rect 2411 7437 2414 7445
rect 2416 7437 2417 7445
rect 2434 7437 2435 7445
rect 2437 7437 2438 7445
rect 2450 7437 2451 7445
rect 2453 7441 2454 7445
rect 2453 7437 2458 7441
rect 2466 7437 2467 7445
rect 2469 7437 2472 7445
rect 2474 7437 2475 7445
rect 2487 7437 2488 7445
rect 2490 7437 2491 7445
rect 2503 7437 2504 7445
rect 2506 7437 2509 7445
rect 2511 7437 2512 7445
rect 2524 7437 2525 7445
rect 2527 7441 2528 7445
rect 2527 7437 2532 7441
rect 2540 7437 2541 7445
rect 2543 7437 2546 7445
rect 2548 7437 2549 7445
rect 2566 7437 2567 7445
rect 2569 7437 2570 7445
rect 2582 7437 2583 7445
rect 2585 7441 2586 7445
rect 2585 7437 2590 7441
rect 2598 7437 2599 7445
rect 2601 7437 2604 7445
rect 2606 7437 2607 7445
rect 2619 7437 2620 7445
rect 2622 7437 2623 7445
rect 2635 7437 2636 7445
rect 2638 7437 2641 7445
rect 2643 7437 2644 7445
rect 2656 7437 2657 7445
rect 2659 7441 2660 7445
rect 2659 7437 2664 7441
rect 2672 7437 2673 7445
rect 2675 7437 2678 7445
rect 2680 7437 2681 7445
rect 2698 7437 2699 7445
rect 2701 7437 2702 7445
rect 2714 7437 2715 7445
rect 2717 7441 2718 7445
rect 2717 7437 2722 7441
rect 2730 7437 2731 7445
rect 2733 7437 2736 7445
rect 2738 7437 2739 7445
rect 2751 7437 2752 7445
rect 2754 7437 2755 7445
rect 3316 7437 3317 7445
rect 3319 7437 3322 7445
rect 3324 7437 3325 7445
rect 3337 7437 3338 7445
rect 3340 7441 3341 7445
rect 3340 7437 3345 7441
rect 3353 7437 3354 7445
rect 3356 7437 3359 7445
rect 3361 7437 3362 7445
rect 3379 7437 3380 7445
rect 3382 7437 3383 7445
rect 3395 7437 3396 7445
rect 3398 7441 3399 7445
rect 3398 7437 3403 7441
rect 3411 7437 3412 7445
rect 3414 7437 3417 7445
rect 3419 7437 3420 7445
rect 3432 7437 3433 7445
rect 3435 7437 3436 7445
rect 3448 7437 3449 7445
rect 3451 7437 3454 7445
rect 3456 7437 3457 7445
rect 3469 7437 3470 7445
rect 3472 7441 3473 7445
rect 3472 7437 3477 7441
rect 3485 7437 3486 7445
rect 3488 7437 3491 7445
rect 3493 7437 3494 7445
rect 3511 7437 3512 7445
rect 3514 7437 3515 7445
rect 3527 7437 3528 7445
rect 3530 7441 3531 7445
rect 3530 7437 3535 7441
rect 3543 7437 3544 7445
rect 3546 7437 3549 7445
rect 3551 7437 3552 7445
rect 3564 7437 3565 7445
rect 3567 7437 3568 7445
rect 3580 7437 3581 7445
rect 3583 7437 3586 7445
rect 3588 7437 3589 7445
rect 3601 7437 3602 7445
rect 3604 7441 3605 7445
rect 3604 7437 3609 7441
rect 3617 7437 3618 7445
rect 3620 7437 3623 7445
rect 3625 7437 3626 7445
rect 3643 7437 3644 7445
rect 3646 7437 3647 7445
rect 3659 7437 3660 7445
rect 3662 7441 3663 7445
rect 3662 7437 3667 7441
rect 3675 7437 3676 7445
rect 3678 7437 3681 7445
rect 3683 7437 3684 7445
rect 3696 7437 3697 7445
rect 3699 7437 3700 7445
rect 1472 6869 1473 6877
rect 1475 6869 1476 6877
rect 1488 6869 1489 6877
rect 1491 6869 1494 6877
rect 1496 6869 1497 6877
rect 1505 6873 1510 6877
rect 1509 6869 1510 6873
rect 1512 6869 1513 6877
rect 1525 6869 1526 6877
rect 1528 6869 1529 6877
rect 1546 6869 1547 6877
rect 1549 6869 1552 6877
rect 1554 6869 1555 6877
rect 1563 6873 1568 6877
rect 1567 6869 1568 6873
rect 1570 6869 1571 6877
rect 1583 6869 1584 6877
rect 1586 6869 1589 6877
rect 1591 6869 1592 6877
rect 1604 6869 1605 6877
rect 1607 6869 1608 6877
rect 1620 6869 1621 6877
rect 1623 6869 1626 6877
rect 1628 6869 1629 6877
rect 1637 6873 1642 6877
rect 1641 6869 1642 6873
rect 1644 6869 1645 6877
rect 1657 6869 1658 6877
rect 1660 6869 1661 6877
rect 1678 6869 1679 6877
rect 1681 6869 1684 6877
rect 1686 6869 1687 6877
rect 1695 6873 1700 6877
rect 1699 6869 1700 6873
rect 1702 6869 1703 6877
rect 1715 6869 1716 6877
rect 1718 6869 1721 6877
rect 1723 6869 1724 6877
rect 1736 6869 1737 6877
rect 1739 6869 1740 6877
rect 1752 6869 1753 6877
rect 1755 6869 1758 6877
rect 1760 6869 1761 6877
rect 1769 6873 1774 6877
rect 1773 6869 1774 6873
rect 1776 6869 1777 6877
rect 1789 6869 1790 6877
rect 1792 6869 1793 6877
rect 1810 6869 1811 6877
rect 1813 6869 1816 6877
rect 1818 6869 1819 6877
rect 1827 6873 1832 6877
rect 1831 6869 1832 6873
rect 1834 6869 1835 6877
rect 1847 6869 1848 6877
rect 1850 6869 1853 6877
rect 1855 6869 1856 6877
rect 2417 6869 2418 6877
rect 2420 6869 2421 6877
rect 2433 6869 2434 6877
rect 2436 6869 2439 6877
rect 2441 6869 2442 6877
rect 2450 6873 2455 6877
rect 2454 6869 2455 6873
rect 2457 6869 2458 6877
rect 2470 6869 2471 6877
rect 2473 6869 2474 6877
rect 2491 6869 2492 6877
rect 2494 6869 2497 6877
rect 2499 6869 2500 6877
rect 2508 6873 2513 6877
rect 2512 6869 2513 6873
rect 2515 6869 2516 6877
rect 2528 6869 2529 6877
rect 2531 6869 2534 6877
rect 2536 6869 2537 6877
rect 2549 6869 2550 6877
rect 2552 6869 2553 6877
rect 2565 6869 2566 6877
rect 2568 6869 2571 6877
rect 2573 6869 2574 6877
rect 2582 6873 2587 6877
rect 2586 6869 2587 6873
rect 2589 6869 2590 6877
rect 2602 6869 2603 6877
rect 2605 6869 2606 6877
rect 2623 6869 2624 6877
rect 2626 6869 2629 6877
rect 2631 6869 2632 6877
rect 2640 6873 2645 6877
rect 2644 6869 2645 6873
rect 2647 6869 2648 6877
rect 2660 6869 2661 6877
rect 2663 6869 2666 6877
rect 2668 6869 2669 6877
rect 2681 6869 2682 6877
rect 2684 6869 2685 6877
rect 2697 6869 2698 6877
rect 2700 6869 2703 6877
rect 2705 6869 2706 6877
rect 2714 6873 2719 6877
rect 2718 6869 2719 6873
rect 2721 6869 2722 6877
rect 2734 6869 2735 6877
rect 2737 6869 2738 6877
rect 2755 6869 2756 6877
rect 2758 6869 2761 6877
rect 2763 6869 2764 6877
rect 2772 6873 2777 6877
rect 2776 6869 2777 6873
rect 2779 6869 2780 6877
rect 2792 6869 2793 6877
rect 2795 6869 2798 6877
rect 2800 6869 2801 6877
rect 1472 6729 1473 6737
rect 1475 6729 1476 6737
rect 1488 6729 1489 6737
rect 1491 6729 1494 6737
rect 1496 6729 1497 6737
rect 1505 6733 1510 6737
rect 1509 6729 1510 6733
rect 1512 6729 1513 6737
rect 1525 6729 1526 6737
rect 1528 6729 1529 6737
rect 1546 6729 1547 6737
rect 1549 6729 1552 6737
rect 1554 6729 1555 6737
rect 1563 6733 1568 6737
rect 1567 6729 1568 6733
rect 1570 6729 1571 6737
rect 1583 6729 1584 6737
rect 1586 6729 1589 6737
rect 1591 6729 1592 6737
rect 1604 6729 1605 6737
rect 1607 6729 1608 6737
rect 1620 6729 1621 6737
rect 1623 6729 1626 6737
rect 1628 6729 1629 6737
rect 1637 6733 1642 6737
rect 1641 6729 1642 6733
rect 1644 6729 1645 6737
rect 1657 6729 1658 6737
rect 1660 6729 1661 6737
rect 1678 6729 1679 6737
rect 1681 6729 1684 6737
rect 1686 6729 1687 6737
rect 1695 6733 1700 6737
rect 1699 6729 1700 6733
rect 1702 6729 1703 6737
rect 1715 6729 1716 6737
rect 1718 6729 1721 6737
rect 1723 6729 1724 6737
rect 1736 6729 1737 6737
rect 1739 6729 1740 6737
rect 1752 6729 1753 6737
rect 1755 6729 1758 6737
rect 1760 6729 1761 6737
rect 1769 6733 1774 6737
rect 1773 6729 1774 6733
rect 1776 6729 1777 6737
rect 1789 6729 1790 6737
rect 1792 6729 1793 6737
rect 1810 6729 1811 6737
rect 1813 6729 1816 6737
rect 1818 6729 1819 6737
rect 1827 6733 1832 6737
rect 1831 6729 1832 6733
rect 1834 6729 1835 6737
rect 1847 6729 1848 6737
rect 1850 6729 1853 6737
rect 1855 6729 1856 6737
rect 2417 6729 2418 6737
rect 2420 6729 2421 6737
rect 2433 6729 2434 6737
rect 2436 6729 2439 6737
rect 2441 6729 2442 6737
rect 2450 6733 2455 6737
rect 2454 6729 2455 6733
rect 2457 6729 2458 6737
rect 2470 6729 2471 6737
rect 2473 6729 2474 6737
rect 2491 6729 2492 6737
rect 2494 6729 2497 6737
rect 2499 6729 2500 6737
rect 2508 6733 2513 6737
rect 2512 6729 2513 6733
rect 2515 6729 2516 6737
rect 2528 6729 2529 6737
rect 2531 6729 2534 6737
rect 2536 6729 2537 6737
rect 2549 6729 2550 6737
rect 2552 6729 2553 6737
rect 2565 6729 2566 6737
rect 2568 6729 2571 6737
rect 2573 6729 2574 6737
rect 2582 6733 2587 6737
rect 2586 6729 2587 6733
rect 2589 6729 2590 6737
rect 2602 6729 2603 6737
rect 2605 6729 2606 6737
rect 2623 6729 2624 6737
rect 2626 6729 2629 6737
rect 2631 6729 2632 6737
rect 2640 6733 2645 6737
rect 2644 6729 2645 6733
rect 2647 6729 2648 6737
rect 2660 6729 2661 6737
rect 2663 6729 2666 6737
rect 2668 6729 2669 6737
rect 2681 6729 2682 6737
rect 2684 6729 2685 6737
rect 2697 6729 2698 6737
rect 2700 6729 2703 6737
rect 2705 6729 2706 6737
rect 2714 6733 2719 6737
rect 2718 6729 2719 6733
rect 2721 6729 2722 6737
rect 2734 6729 2735 6737
rect 2737 6729 2738 6737
rect 2755 6729 2756 6737
rect 2758 6729 2761 6737
rect 2763 6729 2764 6737
rect 2772 6733 2777 6737
rect 2776 6729 2777 6733
rect 2779 6729 2780 6737
rect 2792 6729 2793 6737
rect 2795 6729 2798 6737
rect 2800 6729 2801 6737
rect 953 6699 954 6707
rect 956 6699 957 6707
rect 969 6699 970 6707
rect 972 6699 975 6707
rect 977 6699 978 6707
rect 986 6703 991 6707
rect 990 6699 991 6703
rect 993 6699 994 6707
rect 1006 6699 1007 6707
rect 1009 6699 1010 6707
rect 1027 6699 1028 6707
rect 1030 6699 1033 6707
rect 1035 6699 1036 6707
rect 1044 6703 1049 6707
rect 1048 6699 1049 6703
rect 1051 6699 1052 6707
rect 1064 6699 1065 6707
rect 1067 6699 1070 6707
rect 1072 6699 1073 6707
rect 1898 6699 1899 6707
rect 1901 6699 1902 6707
rect 1914 6699 1915 6707
rect 1917 6699 1920 6707
rect 1922 6699 1923 6707
rect 1931 6703 1936 6707
rect 1935 6699 1936 6703
rect 1938 6699 1939 6707
rect 1951 6699 1952 6707
rect 1954 6699 1955 6707
rect 1972 6699 1973 6707
rect 1975 6699 1978 6707
rect 1980 6699 1981 6707
rect 1989 6703 1994 6707
rect 1993 6699 1994 6703
rect 1996 6699 1997 6707
rect 2009 6699 2010 6707
rect 2012 6699 2015 6707
rect 2017 6699 2018 6707
rect 1472 6643 1473 6651
rect 1475 6643 1476 6651
rect 1488 6643 1489 6651
rect 1491 6643 1494 6651
rect 1496 6643 1497 6651
rect 1505 6647 1510 6651
rect 1509 6643 1510 6647
rect 1512 6643 1513 6651
rect 1525 6643 1526 6651
rect 1528 6643 1529 6651
rect 1546 6643 1547 6651
rect 1549 6643 1552 6651
rect 1554 6643 1555 6651
rect 1563 6647 1568 6651
rect 1567 6643 1568 6647
rect 1570 6643 1571 6651
rect 1583 6643 1584 6651
rect 1586 6643 1589 6651
rect 1591 6643 1592 6651
rect 1604 6643 1605 6651
rect 1607 6643 1608 6651
rect 1620 6643 1621 6651
rect 1623 6643 1626 6651
rect 1628 6643 1629 6651
rect 1637 6647 1642 6651
rect 1641 6643 1642 6647
rect 1644 6643 1645 6651
rect 1657 6643 1658 6651
rect 1660 6643 1661 6651
rect 1678 6643 1679 6651
rect 1681 6643 1684 6651
rect 1686 6643 1687 6651
rect 1695 6647 1700 6651
rect 1699 6643 1700 6647
rect 1702 6643 1703 6651
rect 1715 6643 1716 6651
rect 1718 6643 1721 6651
rect 1723 6643 1724 6651
rect 1736 6643 1737 6651
rect 1739 6643 1740 6651
rect 1752 6643 1753 6651
rect 1755 6643 1758 6651
rect 1760 6643 1761 6651
rect 1769 6647 1774 6651
rect 1773 6643 1774 6647
rect 1776 6643 1777 6651
rect 1789 6643 1790 6651
rect 1792 6643 1793 6651
rect 1810 6643 1811 6651
rect 1813 6643 1816 6651
rect 1818 6643 1819 6651
rect 1827 6647 1832 6651
rect 1831 6643 1832 6647
rect 1834 6643 1835 6651
rect 1847 6643 1848 6651
rect 1850 6643 1853 6651
rect 1855 6643 1856 6651
rect 2417 6643 2418 6651
rect 2420 6643 2421 6651
rect 2433 6643 2434 6651
rect 2436 6643 2439 6651
rect 2441 6643 2442 6651
rect 2450 6647 2455 6651
rect 2454 6643 2455 6647
rect 2457 6643 2458 6651
rect 2470 6643 2471 6651
rect 2473 6643 2474 6651
rect 2491 6643 2492 6651
rect 2494 6643 2497 6651
rect 2499 6643 2500 6651
rect 2508 6647 2513 6651
rect 2512 6643 2513 6647
rect 2515 6643 2516 6651
rect 2528 6643 2529 6651
rect 2531 6643 2534 6651
rect 2536 6643 2537 6651
rect 2549 6643 2550 6651
rect 2552 6643 2553 6651
rect 2565 6643 2566 6651
rect 2568 6643 2571 6651
rect 2573 6643 2574 6651
rect 2582 6647 2587 6651
rect 2586 6643 2587 6647
rect 2589 6643 2590 6651
rect 2602 6643 2603 6651
rect 2605 6643 2606 6651
rect 2623 6643 2624 6651
rect 2626 6643 2629 6651
rect 2631 6643 2632 6651
rect 2640 6647 2645 6651
rect 2644 6643 2645 6647
rect 2647 6643 2648 6651
rect 2660 6643 2661 6651
rect 2663 6643 2666 6651
rect 2668 6643 2669 6651
rect 2681 6643 2682 6651
rect 2684 6643 2685 6651
rect 2697 6643 2698 6651
rect 2700 6643 2703 6651
rect 2705 6643 2706 6651
rect 2714 6647 2719 6651
rect 2718 6643 2719 6647
rect 2721 6643 2722 6651
rect 2734 6643 2735 6651
rect 2737 6643 2738 6651
rect 2755 6643 2756 6651
rect 2758 6643 2761 6651
rect 2763 6643 2764 6651
rect 2772 6647 2777 6651
rect 2776 6643 2777 6647
rect 2779 6643 2780 6651
rect 2792 6643 2793 6651
rect 2795 6643 2798 6651
rect 2800 6643 2801 6651
rect 953 6613 954 6621
rect 956 6613 957 6621
rect 969 6613 970 6621
rect 972 6613 975 6621
rect 977 6613 978 6621
rect 986 6617 991 6621
rect 990 6613 991 6617
rect 993 6613 994 6621
rect 1006 6613 1007 6621
rect 1009 6613 1010 6621
rect 1027 6613 1028 6621
rect 1030 6613 1033 6621
rect 1035 6613 1036 6621
rect 1044 6617 1049 6621
rect 1048 6613 1049 6617
rect 1051 6613 1052 6621
rect 1064 6613 1065 6621
rect 1067 6613 1070 6621
rect 1072 6613 1073 6621
rect 1898 6613 1899 6621
rect 1901 6613 1902 6621
rect 1914 6613 1915 6621
rect 1917 6613 1920 6621
rect 1922 6613 1923 6621
rect 1931 6617 1936 6621
rect 1935 6613 1936 6617
rect 1938 6613 1939 6621
rect 1951 6613 1952 6621
rect 1954 6613 1955 6621
rect 1972 6613 1973 6621
rect 1975 6613 1978 6621
rect 1980 6613 1981 6621
rect 1989 6617 1994 6621
rect 1993 6613 1994 6617
rect 1996 6613 1997 6621
rect 2009 6613 2010 6621
rect 2012 6613 2015 6621
rect 2017 6613 2018 6621
rect 952 6532 953 6540
rect 955 6532 956 6540
rect 970 6532 971 6540
rect 973 6532 976 6540
rect 978 6532 983 6540
rect 995 6532 996 6540
rect 998 6532 999 6540
rect 1016 6532 1017 6540
rect 1019 6532 1021 6540
rect 1042 6532 1043 6540
rect 1045 6532 1048 6540
rect 1050 6532 1055 6540
rect 1070 6532 1071 6540
rect 1073 6532 1074 6540
rect 1086 6532 1087 6540
rect 1089 6532 1090 6540
rect 1111 6532 1112 6540
rect 1114 6532 1115 6540
rect 1119 6532 1125 6540
rect 1129 6532 1130 6540
rect 1132 6532 1133 6540
rect 1158 6537 1159 6545
rect 1161 6537 1164 6545
rect 1166 6537 1169 6545
rect 1213 6532 1214 6540
rect 1216 6532 1217 6540
rect 1231 6532 1232 6540
rect 1234 6532 1237 6540
rect 1239 6532 1244 6540
rect 1256 6532 1257 6540
rect 1259 6532 1260 6540
rect 1277 6532 1278 6540
rect 1280 6532 1282 6540
rect 1303 6532 1304 6540
rect 1306 6532 1309 6540
rect 1311 6532 1316 6540
rect 1331 6532 1332 6540
rect 1334 6532 1335 6540
rect 1347 6532 1348 6540
rect 1350 6532 1351 6540
rect 1363 6532 1364 6540
rect 1366 6532 1367 6540
rect 1897 6532 1898 6540
rect 1900 6532 1901 6540
rect 1915 6532 1916 6540
rect 1918 6532 1921 6540
rect 1923 6532 1928 6540
rect 1940 6532 1941 6540
rect 1943 6532 1944 6540
rect 1961 6532 1962 6540
rect 1964 6532 1966 6540
rect 1987 6532 1988 6540
rect 1990 6532 1993 6540
rect 1995 6532 2000 6540
rect 2015 6532 2016 6540
rect 2018 6532 2019 6540
rect 2031 6532 2032 6540
rect 2034 6532 2035 6540
rect 2056 6532 2057 6540
rect 2059 6532 2060 6540
rect 2064 6532 2070 6540
rect 2074 6532 2075 6540
rect 2077 6532 2078 6540
rect 2103 6537 2104 6545
rect 2106 6537 2109 6545
rect 2111 6537 2114 6545
rect 2158 6532 2159 6540
rect 2161 6532 2162 6540
rect 2176 6532 2177 6540
rect 2179 6532 2182 6540
rect 2184 6532 2189 6540
rect 2201 6532 2202 6540
rect 2204 6532 2205 6540
rect 2222 6532 2223 6540
rect 2225 6532 2227 6540
rect 2248 6532 2249 6540
rect 2251 6532 2254 6540
rect 2256 6532 2261 6540
rect 2276 6532 2277 6540
rect 2279 6532 2280 6540
rect 2292 6532 2293 6540
rect 2295 6532 2296 6540
rect 2308 6532 2309 6540
rect 2311 6532 2312 6540
rect 1472 6501 1473 6509
rect 1475 6501 1476 6509
rect 1488 6501 1489 6509
rect 1491 6501 1494 6509
rect 1496 6501 1497 6509
rect 1505 6505 1510 6509
rect 1509 6501 1510 6505
rect 1512 6501 1513 6509
rect 1525 6501 1526 6509
rect 1528 6501 1529 6509
rect 1546 6501 1547 6509
rect 1549 6501 1552 6509
rect 1554 6501 1555 6509
rect 1563 6505 1568 6509
rect 1567 6501 1568 6505
rect 1570 6501 1571 6509
rect 1583 6501 1584 6509
rect 1586 6501 1589 6509
rect 1591 6501 1592 6509
rect 1604 6501 1605 6509
rect 1607 6501 1608 6509
rect 1620 6501 1621 6509
rect 1623 6501 1626 6509
rect 1628 6501 1629 6509
rect 1637 6505 1642 6509
rect 1641 6501 1642 6505
rect 1644 6501 1645 6509
rect 1657 6501 1658 6509
rect 1660 6501 1661 6509
rect 1678 6501 1679 6509
rect 1681 6501 1684 6509
rect 1686 6501 1687 6509
rect 1695 6505 1700 6509
rect 1699 6501 1700 6505
rect 1702 6501 1703 6509
rect 1715 6501 1716 6509
rect 1718 6501 1721 6509
rect 1723 6501 1724 6509
rect 1736 6501 1737 6509
rect 1739 6501 1740 6509
rect 1752 6501 1753 6509
rect 1755 6501 1758 6509
rect 1760 6501 1761 6509
rect 1769 6505 1774 6509
rect 1773 6501 1774 6505
rect 1776 6501 1777 6509
rect 1789 6501 1790 6509
rect 1792 6501 1793 6509
rect 1810 6501 1811 6509
rect 1813 6501 1816 6509
rect 1818 6501 1819 6509
rect 1827 6505 1832 6509
rect 1831 6501 1832 6505
rect 1834 6501 1835 6509
rect 1847 6501 1848 6509
rect 1850 6501 1853 6509
rect 1855 6501 1856 6509
rect 2417 6501 2418 6509
rect 2420 6501 2421 6509
rect 2433 6501 2434 6509
rect 2436 6501 2439 6509
rect 2441 6501 2442 6509
rect 2450 6505 2455 6509
rect 2454 6501 2455 6505
rect 2457 6501 2458 6509
rect 2470 6501 2471 6509
rect 2473 6501 2474 6509
rect 2491 6501 2492 6509
rect 2494 6501 2497 6509
rect 2499 6501 2500 6509
rect 2508 6505 2513 6509
rect 2512 6501 2513 6505
rect 2515 6501 2516 6509
rect 2528 6501 2529 6509
rect 2531 6501 2534 6509
rect 2536 6501 2537 6509
rect 2549 6501 2550 6509
rect 2552 6501 2553 6509
rect 2565 6501 2566 6509
rect 2568 6501 2571 6509
rect 2573 6501 2574 6509
rect 2582 6505 2587 6509
rect 2586 6501 2587 6505
rect 2589 6501 2590 6509
rect 2602 6501 2603 6509
rect 2605 6501 2606 6509
rect 2623 6501 2624 6509
rect 2626 6501 2629 6509
rect 2631 6501 2632 6509
rect 2640 6505 2645 6509
rect 2644 6501 2645 6505
rect 2647 6501 2648 6509
rect 2660 6501 2661 6509
rect 2663 6501 2666 6509
rect 2668 6501 2669 6509
rect 2681 6501 2682 6509
rect 2684 6501 2685 6509
rect 2697 6501 2698 6509
rect 2700 6501 2703 6509
rect 2705 6501 2706 6509
rect 2714 6505 2719 6509
rect 2718 6501 2719 6505
rect 2721 6501 2722 6509
rect 2734 6501 2735 6509
rect 2737 6501 2738 6509
rect 2755 6501 2756 6509
rect 2758 6501 2761 6509
rect 2763 6501 2764 6509
rect 2772 6505 2777 6509
rect 2776 6501 2777 6505
rect 2779 6501 2780 6509
rect 2792 6501 2793 6509
rect 2795 6501 2798 6509
rect 2800 6501 2801 6509
rect 1135 6433 1136 6441
rect 1138 6433 1139 6441
rect 1158 6439 1159 6447
rect 1161 6439 1164 6447
rect 1166 6439 1169 6447
rect 1213 6446 1214 6454
rect 1216 6446 1217 6454
rect 1231 6446 1232 6454
rect 1234 6446 1237 6454
rect 1239 6446 1244 6454
rect 1256 6446 1257 6454
rect 1259 6446 1260 6454
rect 1277 6446 1278 6454
rect 1280 6446 1282 6454
rect 1303 6446 1304 6454
rect 1306 6446 1309 6454
rect 1311 6446 1316 6454
rect 1331 6446 1332 6454
rect 1334 6446 1335 6454
rect 1347 6446 1348 6454
rect 1350 6446 1351 6454
rect 1363 6446 1364 6454
rect 1366 6446 1367 6454
rect 2080 6433 2081 6441
rect 2083 6433 2084 6441
rect 2103 6439 2104 6447
rect 2106 6439 2109 6447
rect 2111 6439 2114 6447
rect 2158 6446 2159 6454
rect 2161 6446 2162 6454
rect 2176 6446 2177 6454
rect 2179 6446 2182 6454
rect 2184 6446 2189 6454
rect 2201 6446 2202 6454
rect 2204 6446 2205 6454
rect 2222 6446 2223 6454
rect 2225 6446 2227 6454
rect 2248 6446 2249 6454
rect 2251 6446 2254 6454
rect 2256 6446 2261 6454
rect 2276 6446 2277 6454
rect 2279 6446 2280 6454
rect 2292 6446 2293 6454
rect 2295 6446 2296 6454
rect 2308 6446 2309 6454
rect 2311 6446 2312 6454
rect 987 6401 988 6409
rect 990 6401 993 6409
rect 995 6401 998 6409
rect 1077 6401 1078 6409
rect 1080 6401 1083 6409
rect 1085 6401 1088 6409
rect 1158 6401 1159 6409
rect 1161 6401 1164 6409
rect 1166 6401 1169 6409
rect 1213 6400 1214 6408
rect 1216 6400 1217 6408
rect 1231 6400 1232 6408
rect 1234 6400 1237 6408
rect 1239 6400 1244 6408
rect 1256 6400 1257 6408
rect 1259 6400 1260 6408
rect 1277 6400 1278 6408
rect 1280 6400 1282 6408
rect 1303 6400 1304 6408
rect 1306 6400 1309 6408
rect 1311 6400 1316 6408
rect 1331 6400 1332 6408
rect 1334 6400 1335 6408
rect 1347 6400 1348 6408
rect 1350 6400 1351 6408
rect 1363 6400 1364 6408
rect 1366 6400 1367 6408
rect 1932 6401 1933 6409
rect 1935 6401 1938 6409
rect 1940 6401 1943 6409
rect 2022 6401 2023 6409
rect 2025 6401 2028 6409
rect 2030 6401 2033 6409
rect 2103 6401 2104 6409
rect 2106 6401 2109 6409
rect 2111 6401 2114 6409
rect 2158 6400 2159 6408
rect 2161 6400 2162 6408
rect 2176 6400 2177 6408
rect 2179 6400 2182 6408
rect 2184 6400 2189 6408
rect 2201 6400 2202 6408
rect 2204 6400 2205 6408
rect 2222 6400 2223 6408
rect 2225 6400 2227 6408
rect 2248 6400 2249 6408
rect 2251 6400 2254 6408
rect 2256 6400 2261 6408
rect 2276 6400 2277 6408
rect 2279 6400 2280 6408
rect 2292 6400 2293 6408
rect 2295 6400 2296 6408
rect 2308 6400 2309 6408
rect 2311 6400 2312 6408
rect 964 6301 965 6309
rect 967 6301 968 6309
rect 987 6307 988 6315
rect 990 6307 993 6315
rect 995 6307 998 6315
rect 1018 6301 1019 6309
rect 1021 6301 1022 6309
rect 1054 6301 1055 6309
rect 1057 6301 1058 6309
rect 1077 6307 1078 6315
rect 1080 6307 1083 6315
rect 1085 6307 1088 6315
rect 1108 6301 1109 6309
rect 1111 6301 1112 6309
rect 1135 6301 1136 6309
rect 1138 6301 1139 6309
rect 1158 6307 1159 6315
rect 1161 6307 1164 6315
rect 1166 6307 1169 6315
rect 1213 6314 1214 6322
rect 1216 6314 1217 6322
rect 1231 6314 1232 6322
rect 1234 6314 1237 6322
rect 1239 6314 1244 6322
rect 1256 6314 1257 6322
rect 1259 6314 1260 6322
rect 1277 6314 1278 6322
rect 1280 6314 1282 6322
rect 1303 6314 1304 6322
rect 1306 6314 1309 6322
rect 1311 6314 1316 6322
rect 1331 6314 1332 6322
rect 1334 6314 1335 6322
rect 1347 6314 1348 6322
rect 1350 6314 1351 6322
rect 1363 6314 1364 6322
rect 1366 6314 1367 6322
rect 1909 6301 1910 6309
rect 1912 6301 1913 6309
rect 1932 6307 1933 6315
rect 1935 6307 1938 6315
rect 1940 6307 1943 6315
rect 1963 6301 1964 6309
rect 1966 6301 1967 6309
rect 1999 6301 2000 6309
rect 2002 6301 2003 6309
rect 2022 6307 2023 6315
rect 2025 6307 2028 6315
rect 2030 6307 2033 6315
rect 2053 6301 2054 6309
rect 2056 6301 2057 6309
rect 2080 6301 2081 6309
rect 2083 6301 2084 6309
rect 2103 6307 2104 6315
rect 2106 6307 2109 6315
rect 2111 6307 2114 6315
rect 2158 6314 2159 6322
rect 2161 6314 2162 6322
rect 2176 6314 2177 6322
rect 2179 6314 2182 6322
rect 2184 6314 2189 6322
rect 2201 6314 2202 6322
rect 2204 6314 2205 6322
rect 2222 6314 2223 6322
rect 2225 6314 2227 6322
rect 2248 6314 2249 6322
rect 2251 6314 2254 6322
rect 2256 6314 2261 6322
rect 2276 6314 2277 6322
rect 2279 6314 2280 6322
rect 2292 6314 2293 6322
rect 2295 6314 2296 6322
rect 2308 6314 2309 6322
rect 2311 6314 2312 6322
rect 1053 6266 1054 6274
rect 1056 6266 1059 6274
rect 1061 6266 1064 6274
rect 1158 6266 1159 6274
rect 1161 6266 1164 6274
rect 1166 6266 1169 6274
rect 1213 6268 1214 6276
rect 1216 6268 1217 6276
rect 1231 6268 1232 6276
rect 1234 6268 1237 6276
rect 1239 6268 1244 6276
rect 1256 6268 1257 6276
rect 1259 6268 1260 6276
rect 1277 6268 1278 6276
rect 1280 6268 1282 6276
rect 1303 6268 1304 6276
rect 1306 6268 1309 6276
rect 1311 6268 1316 6276
rect 1331 6268 1332 6276
rect 1334 6268 1335 6276
rect 1347 6268 1348 6276
rect 1350 6268 1351 6276
rect 1363 6268 1364 6276
rect 1366 6268 1367 6276
rect 1998 6266 1999 6274
rect 2001 6266 2004 6274
rect 2006 6266 2009 6274
rect 2103 6266 2104 6274
rect 2106 6266 2109 6274
rect 2111 6266 2114 6274
rect 2158 6268 2159 6276
rect 2161 6268 2162 6276
rect 2176 6268 2177 6276
rect 2179 6268 2182 6276
rect 2184 6268 2189 6276
rect 2201 6268 2202 6276
rect 2204 6268 2205 6276
rect 2222 6268 2223 6276
rect 2225 6268 2227 6276
rect 2248 6268 2249 6276
rect 2251 6268 2254 6276
rect 2256 6268 2261 6276
rect 2276 6268 2277 6276
rect 2279 6268 2280 6276
rect 2292 6268 2293 6276
rect 2295 6268 2296 6276
rect 2308 6268 2309 6276
rect 2311 6268 2312 6276
rect 1030 6169 1031 6177
rect 1033 6169 1034 6177
rect 1053 6175 1054 6183
rect 1056 6175 1059 6183
rect 1061 6175 1064 6183
rect 1084 6169 1085 6177
rect 1087 6169 1088 6177
rect 1135 6169 1136 6177
rect 1138 6169 1139 6177
rect 1158 6175 1159 6183
rect 1161 6175 1164 6183
rect 1166 6175 1169 6183
rect 1213 6182 1214 6190
rect 1216 6182 1217 6190
rect 1231 6182 1232 6190
rect 1234 6182 1237 6190
rect 1239 6182 1244 6190
rect 1256 6182 1257 6190
rect 1259 6182 1260 6190
rect 1277 6182 1278 6190
rect 1280 6182 1282 6190
rect 1303 6182 1304 6190
rect 1306 6182 1309 6190
rect 1311 6182 1316 6190
rect 1331 6182 1332 6190
rect 1334 6182 1335 6190
rect 1347 6182 1348 6190
rect 1350 6182 1351 6190
rect 1363 6182 1364 6190
rect 1366 6182 1367 6190
rect 1975 6169 1976 6177
rect 1978 6169 1979 6177
rect 1998 6175 1999 6183
rect 2001 6175 2004 6183
rect 2006 6175 2009 6183
rect 2029 6169 2030 6177
rect 2032 6169 2033 6177
rect 2080 6169 2081 6177
rect 2083 6169 2084 6177
rect 2103 6175 2104 6183
rect 2106 6175 2109 6183
rect 2111 6175 2114 6183
rect 2158 6182 2159 6190
rect 2161 6182 2162 6190
rect 2176 6182 2177 6190
rect 2179 6182 2182 6190
rect 2184 6182 2189 6190
rect 2201 6182 2202 6190
rect 2204 6182 2205 6190
rect 2222 6182 2223 6190
rect 2225 6182 2227 6190
rect 2248 6182 2249 6190
rect 2251 6182 2254 6190
rect 2256 6182 2261 6190
rect 2276 6182 2277 6190
rect 2279 6182 2280 6190
rect 2292 6182 2293 6190
rect 2295 6182 2296 6190
rect 2308 6182 2309 6190
rect 2311 6182 2312 6190
rect 1077 6135 1078 6143
rect 1080 6135 1083 6143
rect 1085 6135 1088 6143
rect 1158 6135 1159 6143
rect 1161 6135 1164 6143
rect 1166 6135 1169 6143
rect 1213 6136 1214 6144
rect 1216 6136 1217 6144
rect 1231 6136 1232 6144
rect 1234 6136 1237 6144
rect 1239 6136 1244 6144
rect 1256 6136 1257 6144
rect 1259 6136 1260 6144
rect 1277 6136 1278 6144
rect 1280 6136 1282 6144
rect 1303 6136 1304 6144
rect 1306 6136 1309 6144
rect 1311 6136 1316 6144
rect 1331 6136 1332 6144
rect 1334 6136 1335 6144
rect 1347 6136 1348 6144
rect 1350 6136 1351 6144
rect 1363 6136 1364 6144
rect 1366 6136 1367 6144
rect 2022 6135 2023 6143
rect 2025 6135 2028 6143
rect 2030 6135 2033 6143
rect 2103 6135 2104 6143
rect 2106 6135 2109 6143
rect 2111 6135 2114 6143
rect 2158 6136 2159 6144
rect 2161 6136 2162 6144
rect 2176 6136 2177 6144
rect 2179 6136 2182 6144
rect 2184 6136 2189 6144
rect 2201 6136 2202 6144
rect 2204 6136 2205 6144
rect 2222 6136 2223 6144
rect 2225 6136 2227 6144
rect 2248 6136 2249 6144
rect 2251 6136 2254 6144
rect 2256 6136 2261 6144
rect 2276 6136 2277 6144
rect 2279 6136 2280 6144
rect 2292 6136 2293 6144
rect 2295 6136 2296 6144
rect 2308 6136 2309 6144
rect 2311 6136 2312 6144
rect 1613 6101 1614 6109
rect 1616 6101 1619 6109
rect 1621 6101 1622 6109
rect 1634 6101 1635 6109
rect 1637 6105 1642 6109
rect 1637 6101 1638 6105
rect 1650 6101 1651 6109
rect 1653 6101 1656 6109
rect 1658 6101 1659 6109
rect 1676 6101 1677 6109
rect 1679 6101 1680 6109
rect 1692 6101 1693 6109
rect 1695 6105 1700 6109
rect 1695 6101 1696 6105
rect 1708 6101 1709 6109
rect 1711 6101 1714 6109
rect 1716 6101 1717 6109
rect 1729 6101 1730 6109
rect 1732 6101 1733 6109
rect 2558 6101 2559 6109
rect 2561 6101 2564 6109
rect 2566 6101 2567 6109
rect 2579 6101 2580 6109
rect 2582 6105 2587 6109
rect 2582 6101 2583 6105
rect 2595 6101 2596 6109
rect 2598 6101 2601 6109
rect 2603 6101 2604 6109
rect 2621 6101 2622 6109
rect 2624 6101 2625 6109
rect 2637 6101 2638 6109
rect 2640 6105 2645 6109
rect 2640 6101 2641 6105
rect 2653 6101 2654 6109
rect 2656 6101 2659 6109
rect 2661 6101 2662 6109
rect 2674 6101 2675 6109
rect 2677 6101 2678 6109
rect 1054 6037 1055 6045
rect 1057 6037 1058 6045
rect 1077 6043 1078 6051
rect 1080 6043 1083 6051
rect 1085 6043 1088 6051
rect 1108 6037 1109 6045
rect 1111 6037 1112 6045
rect 1135 6037 1136 6045
rect 1138 6037 1139 6045
rect 1158 6043 1159 6051
rect 1161 6043 1164 6051
rect 1166 6043 1169 6051
rect 1213 6050 1214 6058
rect 1216 6050 1217 6058
rect 1231 6050 1232 6058
rect 1234 6050 1237 6058
rect 1239 6050 1244 6058
rect 1256 6050 1257 6058
rect 1259 6050 1260 6058
rect 1277 6050 1278 6058
rect 1280 6050 1282 6058
rect 1303 6050 1304 6058
rect 1306 6050 1309 6058
rect 1311 6050 1316 6058
rect 1331 6050 1332 6058
rect 1334 6050 1335 6058
rect 1347 6050 1348 6058
rect 1350 6050 1351 6058
rect 1363 6050 1364 6058
rect 1366 6050 1367 6058
rect 1189 6037 1190 6045
rect 1192 6037 1193 6045
rect 1999 6037 2000 6045
rect 2002 6037 2003 6045
rect 2022 6043 2023 6051
rect 2025 6043 2028 6051
rect 2030 6043 2033 6051
rect 2053 6037 2054 6045
rect 2056 6037 2057 6045
rect 2080 6037 2081 6045
rect 2083 6037 2084 6045
rect 2103 6043 2104 6051
rect 2106 6043 2109 6051
rect 2111 6043 2114 6051
rect 2158 6050 2159 6058
rect 2161 6050 2162 6058
rect 2176 6050 2177 6058
rect 2179 6050 2182 6058
rect 2184 6050 2189 6058
rect 2201 6050 2202 6058
rect 2204 6050 2205 6058
rect 2222 6050 2223 6058
rect 2225 6050 2227 6058
rect 2248 6050 2249 6058
rect 2251 6050 2254 6058
rect 2256 6050 2261 6058
rect 2276 6050 2277 6058
rect 2279 6050 2280 6058
rect 2292 6050 2293 6058
rect 2295 6050 2296 6058
rect 2308 6050 2309 6058
rect 2311 6050 2312 6058
rect 2134 6037 2135 6045
rect 2137 6037 2138 6045
rect 1604 5999 1605 6007
rect 1607 5999 1608 6007
rect 1620 5999 1621 6007
rect 1623 5999 1626 6007
rect 1628 5999 1629 6007
rect 1637 6003 1642 6007
rect 1641 5999 1642 6003
rect 1644 5999 1645 6007
rect 1657 5999 1658 6007
rect 1660 5999 1661 6007
rect 1678 5999 1679 6007
rect 1681 5999 1684 6007
rect 1686 5999 1687 6007
rect 1695 6003 1700 6007
rect 1699 5999 1700 6003
rect 1702 5999 1703 6007
rect 1715 5999 1716 6007
rect 1718 5999 1721 6007
rect 1723 5999 1724 6007
rect 2549 5999 2550 6007
rect 2552 5999 2553 6007
rect 2565 5999 2566 6007
rect 2568 5999 2571 6007
rect 2573 5999 2574 6007
rect 2582 6003 2587 6007
rect 2586 5999 2587 6003
rect 2589 5999 2590 6007
rect 2602 5999 2603 6007
rect 2605 5999 2606 6007
rect 2623 5999 2624 6007
rect 2626 5999 2629 6007
rect 2631 5999 2632 6007
rect 2640 6003 2645 6007
rect 2644 5999 2645 6003
rect 2647 5999 2648 6007
rect 2660 5999 2661 6007
rect 2663 5999 2666 6007
rect 2668 5999 2669 6007
rect 856 5966 857 5974
rect 859 5966 860 5974
rect 872 5966 873 5974
rect 875 5966 878 5974
rect 880 5966 881 5974
rect 889 5970 894 5974
rect 893 5966 894 5970
rect 896 5966 897 5974
rect 909 5966 910 5974
rect 912 5966 913 5974
rect 930 5966 931 5974
rect 933 5966 936 5974
rect 938 5966 939 5974
rect 947 5970 952 5974
rect 951 5966 952 5970
rect 954 5966 955 5974
rect 967 5966 968 5974
rect 970 5966 973 5974
rect 975 5966 976 5974
rect 988 5966 989 5974
rect 991 5966 992 5974
rect 1004 5966 1005 5974
rect 1007 5966 1010 5974
rect 1012 5966 1013 5974
rect 1021 5970 1026 5974
rect 1025 5966 1026 5970
rect 1028 5966 1029 5974
rect 1041 5966 1042 5974
rect 1044 5966 1045 5974
rect 1062 5966 1063 5974
rect 1065 5966 1068 5974
rect 1070 5966 1071 5974
rect 1079 5970 1084 5974
rect 1083 5966 1084 5970
rect 1086 5966 1087 5974
rect 1099 5966 1100 5974
rect 1102 5966 1105 5974
rect 1107 5966 1108 5974
rect 1120 5966 1121 5974
rect 1123 5966 1124 5974
rect 1136 5966 1137 5974
rect 1139 5966 1142 5974
rect 1144 5966 1145 5974
rect 1153 5970 1158 5974
rect 1157 5966 1158 5970
rect 1160 5966 1161 5974
rect 1173 5966 1174 5974
rect 1176 5966 1177 5974
rect 1194 5966 1195 5974
rect 1197 5966 1200 5974
rect 1202 5966 1203 5974
rect 1211 5970 1216 5974
rect 1215 5966 1216 5970
rect 1218 5966 1219 5974
rect 1231 5966 1232 5974
rect 1234 5966 1237 5974
rect 1239 5966 1240 5974
rect 1252 5966 1253 5974
rect 1255 5966 1256 5974
rect 1268 5966 1269 5974
rect 1271 5966 1274 5974
rect 1276 5966 1277 5974
rect 1285 5970 1290 5974
rect 1289 5966 1290 5970
rect 1292 5966 1293 5974
rect 1305 5966 1306 5974
rect 1308 5966 1309 5974
rect 1326 5966 1327 5974
rect 1329 5966 1332 5974
rect 1334 5966 1335 5974
rect 1343 5970 1348 5974
rect 1347 5966 1348 5970
rect 1350 5966 1351 5974
rect 1363 5966 1364 5974
rect 1366 5966 1369 5974
rect 1371 5966 1372 5974
rect 1801 5966 1802 5974
rect 1804 5966 1805 5974
rect 1817 5966 1818 5974
rect 1820 5966 1823 5974
rect 1825 5966 1826 5974
rect 1834 5970 1839 5974
rect 1838 5966 1839 5970
rect 1841 5966 1842 5974
rect 1854 5966 1855 5974
rect 1857 5966 1858 5974
rect 1875 5966 1876 5974
rect 1878 5966 1881 5974
rect 1883 5966 1884 5974
rect 1892 5970 1897 5974
rect 1896 5966 1897 5970
rect 1899 5966 1900 5974
rect 1912 5966 1913 5974
rect 1915 5966 1918 5974
rect 1920 5966 1921 5974
rect 1933 5966 1934 5974
rect 1936 5966 1937 5974
rect 1949 5966 1950 5974
rect 1952 5966 1955 5974
rect 1957 5966 1958 5974
rect 1966 5970 1971 5974
rect 1970 5966 1971 5970
rect 1973 5966 1974 5974
rect 1986 5966 1987 5974
rect 1989 5966 1990 5974
rect 2007 5966 2008 5974
rect 2010 5966 2013 5974
rect 2015 5966 2016 5974
rect 2024 5970 2029 5974
rect 2028 5966 2029 5970
rect 2031 5966 2032 5974
rect 2044 5966 2045 5974
rect 2047 5966 2050 5974
rect 2052 5966 2053 5974
rect 2065 5966 2066 5974
rect 2068 5966 2069 5974
rect 2081 5966 2082 5974
rect 2084 5966 2087 5974
rect 2089 5966 2090 5974
rect 2098 5970 2103 5974
rect 2102 5966 2103 5970
rect 2105 5966 2106 5974
rect 2118 5966 2119 5974
rect 2121 5966 2122 5974
rect 2139 5966 2140 5974
rect 2142 5966 2145 5974
rect 2147 5966 2148 5974
rect 2156 5970 2161 5974
rect 2160 5966 2161 5970
rect 2163 5966 2164 5974
rect 2176 5966 2177 5974
rect 2179 5966 2182 5974
rect 2184 5966 2185 5974
rect 2197 5966 2198 5974
rect 2200 5966 2201 5974
rect 2213 5966 2214 5974
rect 2216 5966 2219 5974
rect 2221 5966 2222 5974
rect 2230 5970 2235 5974
rect 2234 5966 2235 5970
rect 2237 5966 2238 5974
rect 2250 5966 2251 5974
rect 2253 5966 2254 5974
rect 2271 5966 2272 5974
rect 2274 5966 2277 5974
rect 2279 5966 2280 5974
rect 2288 5970 2293 5974
rect 2292 5966 2293 5970
rect 2295 5966 2296 5974
rect 2308 5966 2309 5974
rect 2311 5966 2314 5974
rect 2316 5966 2317 5974
rect 1472 5887 1473 5895
rect 1475 5887 1476 5895
rect 1488 5887 1489 5895
rect 1491 5887 1494 5895
rect 1496 5887 1497 5895
rect 1505 5891 1510 5895
rect 1509 5887 1510 5891
rect 1512 5887 1513 5895
rect 1525 5887 1526 5895
rect 1528 5887 1529 5895
rect 1546 5887 1547 5895
rect 1549 5887 1552 5895
rect 1554 5887 1555 5895
rect 1563 5891 1568 5895
rect 1567 5887 1568 5891
rect 1570 5887 1571 5895
rect 1583 5887 1584 5895
rect 1586 5887 1589 5895
rect 1591 5887 1592 5895
rect 1604 5887 1605 5895
rect 1607 5887 1608 5895
rect 1620 5887 1621 5895
rect 1623 5887 1626 5895
rect 1628 5887 1629 5895
rect 1637 5891 1642 5895
rect 1641 5887 1642 5891
rect 1644 5887 1645 5895
rect 1657 5887 1658 5895
rect 1660 5887 1661 5895
rect 1678 5887 1679 5895
rect 1681 5887 1684 5895
rect 1686 5887 1687 5895
rect 1695 5891 1700 5895
rect 1699 5887 1700 5891
rect 1702 5887 1703 5895
rect 1715 5887 1716 5895
rect 1718 5887 1721 5895
rect 1723 5887 1724 5895
rect 1736 5887 1737 5895
rect 1739 5887 1740 5895
rect 1752 5887 1753 5895
rect 1755 5887 1758 5895
rect 1760 5887 1761 5895
rect 1769 5891 1774 5895
rect 1773 5887 1774 5891
rect 1776 5887 1777 5895
rect 1789 5887 1790 5895
rect 1792 5887 1793 5895
rect 1810 5887 1811 5895
rect 1813 5887 1816 5895
rect 1818 5887 1819 5895
rect 1827 5891 1832 5895
rect 1831 5887 1832 5891
rect 1834 5887 1835 5895
rect 1847 5887 1848 5895
rect 1850 5887 1853 5895
rect 1855 5887 1856 5895
rect 2417 5887 2418 5895
rect 2420 5887 2421 5895
rect 2433 5887 2434 5895
rect 2436 5887 2439 5895
rect 2441 5887 2442 5895
rect 2450 5891 2455 5895
rect 2454 5887 2455 5891
rect 2457 5887 2458 5895
rect 2470 5887 2471 5895
rect 2473 5887 2474 5895
rect 2491 5887 2492 5895
rect 2494 5887 2497 5895
rect 2499 5887 2500 5895
rect 2508 5891 2513 5895
rect 2512 5887 2513 5891
rect 2515 5887 2516 5895
rect 2528 5887 2529 5895
rect 2531 5887 2534 5895
rect 2536 5887 2537 5895
rect 2549 5887 2550 5895
rect 2552 5887 2553 5895
rect 2565 5887 2566 5895
rect 2568 5887 2571 5895
rect 2573 5887 2574 5895
rect 2582 5891 2587 5895
rect 2586 5887 2587 5891
rect 2589 5887 2590 5895
rect 2602 5887 2603 5895
rect 2605 5887 2606 5895
rect 2623 5887 2624 5895
rect 2626 5887 2629 5895
rect 2631 5887 2632 5895
rect 2640 5891 2645 5895
rect 2644 5887 2645 5891
rect 2647 5887 2648 5895
rect 2660 5887 2661 5895
rect 2663 5887 2666 5895
rect 2668 5887 2669 5895
rect 2681 5887 2682 5895
rect 2684 5887 2685 5895
rect 2697 5887 2698 5895
rect 2700 5887 2703 5895
rect 2705 5887 2706 5895
rect 2714 5891 2719 5895
rect 2718 5887 2719 5891
rect 2721 5887 2722 5895
rect 2734 5887 2735 5895
rect 2737 5887 2738 5895
rect 2755 5887 2756 5895
rect 2758 5887 2761 5895
rect 2763 5887 2764 5895
rect 2772 5891 2777 5895
rect 2776 5887 2777 5891
rect 2779 5887 2780 5895
rect 2792 5887 2793 5895
rect 2795 5887 2798 5895
rect 2800 5887 2801 5895
rect 1472 5747 1473 5755
rect 1475 5747 1476 5755
rect 1488 5747 1489 5755
rect 1491 5747 1494 5755
rect 1496 5747 1497 5755
rect 1505 5751 1510 5755
rect 1509 5747 1510 5751
rect 1512 5747 1513 5755
rect 1525 5747 1526 5755
rect 1528 5747 1529 5755
rect 1546 5747 1547 5755
rect 1549 5747 1552 5755
rect 1554 5747 1555 5755
rect 1563 5751 1568 5755
rect 1567 5747 1568 5751
rect 1570 5747 1571 5755
rect 1583 5747 1584 5755
rect 1586 5747 1589 5755
rect 1591 5747 1592 5755
rect 1604 5747 1605 5755
rect 1607 5747 1608 5755
rect 1620 5747 1621 5755
rect 1623 5747 1626 5755
rect 1628 5747 1629 5755
rect 1637 5751 1642 5755
rect 1641 5747 1642 5751
rect 1644 5747 1645 5755
rect 1657 5747 1658 5755
rect 1660 5747 1661 5755
rect 1678 5747 1679 5755
rect 1681 5747 1684 5755
rect 1686 5747 1687 5755
rect 1695 5751 1700 5755
rect 1699 5747 1700 5751
rect 1702 5747 1703 5755
rect 1715 5747 1716 5755
rect 1718 5747 1721 5755
rect 1723 5747 1724 5755
rect 1736 5747 1737 5755
rect 1739 5747 1740 5755
rect 1752 5747 1753 5755
rect 1755 5747 1758 5755
rect 1760 5747 1761 5755
rect 1769 5751 1774 5755
rect 1773 5747 1774 5751
rect 1776 5747 1777 5755
rect 1789 5747 1790 5755
rect 1792 5747 1793 5755
rect 1810 5747 1811 5755
rect 1813 5747 1816 5755
rect 1818 5747 1819 5755
rect 1827 5751 1832 5755
rect 1831 5747 1832 5751
rect 1834 5747 1835 5755
rect 1847 5747 1848 5755
rect 1850 5747 1853 5755
rect 1855 5747 1856 5755
rect 2417 5747 2418 5755
rect 2420 5747 2421 5755
rect 2433 5747 2434 5755
rect 2436 5747 2439 5755
rect 2441 5747 2442 5755
rect 2450 5751 2455 5755
rect 2454 5747 2455 5751
rect 2457 5747 2458 5755
rect 2470 5747 2471 5755
rect 2473 5747 2474 5755
rect 2491 5747 2492 5755
rect 2494 5747 2497 5755
rect 2499 5747 2500 5755
rect 2508 5751 2513 5755
rect 2512 5747 2513 5751
rect 2515 5747 2516 5755
rect 2528 5747 2529 5755
rect 2531 5747 2534 5755
rect 2536 5747 2537 5755
rect 2549 5747 2550 5755
rect 2552 5747 2553 5755
rect 2565 5747 2566 5755
rect 2568 5747 2571 5755
rect 2573 5747 2574 5755
rect 2582 5751 2587 5755
rect 2586 5747 2587 5751
rect 2589 5747 2590 5755
rect 2602 5747 2603 5755
rect 2605 5747 2606 5755
rect 2623 5747 2624 5755
rect 2626 5747 2629 5755
rect 2631 5747 2632 5755
rect 2640 5751 2645 5755
rect 2644 5747 2645 5751
rect 2647 5747 2648 5755
rect 2660 5747 2661 5755
rect 2663 5747 2666 5755
rect 2668 5747 2669 5755
rect 2681 5747 2682 5755
rect 2684 5747 2685 5755
rect 2697 5747 2698 5755
rect 2700 5747 2703 5755
rect 2705 5747 2706 5755
rect 2714 5751 2719 5755
rect 2718 5747 2719 5751
rect 2721 5747 2722 5755
rect 2734 5747 2735 5755
rect 2737 5747 2738 5755
rect 2755 5747 2756 5755
rect 2758 5747 2761 5755
rect 2763 5747 2764 5755
rect 2772 5751 2777 5755
rect 2776 5747 2777 5751
rect 2779 5747 2780 5755
rect 2792 5747 2793 5755
rect 2795 5747 2798 5755
rect 2800 5747 2801 5755
rect 953 5717 954 5725
rect 956 5717 957 5725
rect 969 5717 970 5725
rect 972 5717 975 5725
rect 977 5717 978 5725
rect 986 5721 991 5725
rect 990 5717 991 5721
rect 993 5717 994 5725
rect 1006 5717 1007 5725
rect 1009 5717 1010 5725
rect 1027 5717 1028 5725
rect 1030 5717 1033 5725
rect 1035 5717 1036 5725
rect 1044 5721 1049 5725
rect 1048 5717 1049 5721
rect 1051 5717 1052 5725
rect 1064 5717 1065 5725
rect 1067 5717 1070 5725
rect 1072 5717 1073 5725
rect 1898 5717 1899 5725
rect 1901 5717 1902 5725
rect 1914 5717 1915 5725
rect 1917 5717 1920 5725
rect 1922 5717 1923 5725
rect 1931 5721 1936 5725
rect 1935 5717 1936 5721
rect 1938 5717 1939 5725
rect 1951 5717 1952 5725
rect 1954 5717 1955 5725
rect 1972 5717 1973 5725
rect 1975 5717 1978 5725
rect 1980 5717 1981 5725
rect 1989 5721 1994 5725
rect 1993 5717 1994 5721
rect 1996 5717 1997 5725
rect 2009 5717 2010 5725
rect 2012 5717 2015 5725
rect 2017 5717 2018 5725
rect 1472 5661 1473 5669
rect 1475 5661 1476 5669
rect 1488 5661 1489 5669
rect 1491 5661 1494 5669
rect 1496 5661 1497 5669
rect 1505 5665 1510 5669
rect 1509 5661 1510 5665
rect 1512 5661 1513 5669
rect 1525 5661 1526 5669
rect 1528 5661 1529 5669
rect 1546 5661 1547 5669
rect 1549 5661 1552 5669
rect 1554 5661 1555 5669
rect 1563 5665 1568 5669
rect 1567 5661 1568 5665
rect 1570 5661 1571 5669
rect 1583 5661 1584 5669
rect 1586 5661 1589 5669
rect 1591 5661 1592 5669
rect 1604 5661 1605 5669
rect 1607 5661 1608 5669
rect 1620 5661 1621 5669
rect 1623 5661 1626 5669
rect 1628 5661 1629 5669
rect 1637 5665 1642 5669
rect 1641 5661 1642 5665
rect 1644 5661 1645 5669
rect 1657 5661 1658 5669
rect 1660 5661 1661 5669
rect 1678 5661 1679 5669
rect 1681 5661 1684 5669
rect 1686 5661 1687 5669
rect 1695 5665 1700 5669
rect 1699 5661 1700 5665
rect 1702 5661 1703 5669
rect 1715 5661 1716 5669
rect 1718 5661 1721 5669
rect 1723 5661 1724 5669
rect 1736 5661 1737 5669
rect 1739 5661 1740 5669
rect 1752 5661 1753 5669
rect 1755 5661 1758 5669
rect 1760 5661 1761 5669
rect 1769 5665 1774 5669
rect 1773 5661 1774 5665
rect 1776 5661 1777 5669
rect 1789 5661 1790 5669
rect 1792 5661 1793 5669
rect 1810 5661 1811 5669
rect 1813 5661 1816 5669
rect 1818 5661 1819 5669
rect 1827 5665 1832 5669
rect 1831 5661 1832 5665
rect 1834 5661 1835 5669
rect 1847 5661 1848 5669
rect 1850 5661 1853 5669
rect 1855 5661 1856 5669
rect 2417 5661 2418 5669
rect 2420 5661 2421 5669
rect 2433 5661 2434 5669
rect 2436 5661 2439 5669
rect 2441 5661 2442 5669
rect 2450 5665 2455 5669
rect 2454 5661 2455 5665
rect 2457 5661 2458 5669
rect 2470 5661 2471 5669
rect 2473 5661 2474 5669
rect 2491 5661 2492 5669
rect 2494 5661 2497 5669
rect 2499 5661 2500 5669
rect 2508 5665 2513 5669
rect 2512 5661 2513 5665
rect 2515 5661 2516 5669
rect 2528 5661 2529 5669
rect 2531 5661 2534 5669
rect 2536 5661 2537 5669
rect 2549 5661 2550 5669
rect 2552 5661 2553 5669
rect 2565 5661 2566 5669
rect 2568 5661 2571 5669
rect 2573 5661 2574 5669
rect 2582 5665 2587 5669
rect 2586 5661 2587 5665
rect 2589 5661 2590 5669
rect 2602 5661 2603 5669
rect 2605 5661 2606 5669
rect 2623 5661 2624 5669
rect 2626 5661 2629 5669
rect 2631 5661 2632 5669
rect 2640 5665 2645 5669
rect 2644 5661 2645 5665
rect 2647 5661 2648 5669
rect 2660 5661 2661 5669
rect 2663 5661 2666 5669
rect 2668 5661 2669 5669
rect 2681 5661 2682 5669
rect 2684 5661 2685 5669
rect 2697 5661 2698 5669
rect 2700 5661 2703 5669
rect 2705 5661 2706 5669
rect 2714 5665 2719 5669
rect 2718 5661 2719 5665
rect 2721 5661 2722 5669
rect 2734 5661 2735 5669
rect 2737 5661 2738 5669
rect 2755 5661 2756 5669
rect 2758 5661 2761 5669
rect 2763 5661 2764 5669
rect 2772 5665 2777 5669
rect 2776 5661 2777 5665
rect 2779 5661 2780 5669
rect 2792 5661 2793 5669
rect 2795 5661 2798 5669
rect 2800 5661 2801 5669
rect 953 5631 954 5639
rect 956 5631 957 5639
rect 969 5631 970 5639
rect 972 5631 975 5639
rect 977 5631 978 5639
rect 986 5635 991 5639
rect 990 5631 991 5635
rect 993 5631 994 5639
rect 1006 5631 1007 5639
rect 1009 5631 1010 5639
rect 1027 5631 1028 5639
rect 1030 5631 1033 5639
rect 1035 5631 1036 5639
rect 1044 5635 1049 5639
rect 1048 5631 1049 5635
rect 1051 5631 1052 5639
rect 1064 5631 1065 5639
rect 1067 5631 1070 5639
rect 1072 5631 1073 5639
rect 1898 5631 1899 5639
rect 1901 5631 1902 5639
rect 1914 5631 1915 5639
rect 1917 5631 1920 5639
rect 1922 5631 1923 5639
rect 1931 5635 1936 5639
rect 1935 5631 1936 5635
rect 1938 5631 1939 5639
rect 1951 5631 1952 5639
rect 1954 5631 1955 5639
rect 1972 5631 1973 5639
rect 1975 5631 1978 5639
rect 1980 5631 1981 5639
rect 1989 5635 1994 5639
rect 1993 5631 1994 5635
rect 1996 5631 1997 5639
rect 2009 5631 2010 5639
rect 2012 5631 2015 5639
rect 2017 5631 2018 5639
rect 952 5550 953 5558
rect 955 5550 956 5558
rect 970 5550 971 5558
rect 973 5550 976 5558
rect 978 5550 983 5558
rect 995 5550 996 5558
rect 998 5550 999 5558
rect 1016 5550 1017 5558
rect 1019 5550 1021 5558
rect 1042 5550 1043 5558
rect 1045 5550 1048 5558
rect 1050 5550 1055 5558
rect 1070 5550 1071 5558
rect 1073 5550 1074 5558
rect 1086 5550 1087 5558
rect 1089 5550 1090 5558
rect 1111 5550 1112 5558
rect 1114 5550 1115 5558
rect 1119 5550 1125 5558
rect 1129 5550 1130 5558
rect 1132 5550 1133 5558
rect 1158 5555 1159 5563
rect 1161 5555 1164 5563
rect 1166 5555 1169 5563
rect 1213 5550 1214 5558
rect 1216 5550 1217 5558
rect 1231 5550 1232 5558
rect 1234 5550 1237 5558
rect 1239 5550 1244 5558
rect 1256 5550 1257 5558
rect 1259 5550 1260 5558
rect 1277 5550 1278 5558
rect 1280 5550 1282 5558
rect 1303 5550 1304 5558
rect 1306 5550 1309 5558
rect 1311 5550 1316 5558
rect 1331 5550 1332 5558
rect 1334 5550 1335 5558
rect 1347 5550 1348 5558
rect 1350 5550 1351 5558
rect 1363 5550 1364 5558
rect 1366 5550 1367 5558
rect 1897 5550 1898 5558
rect 1900 5550 1901 5558
rect 1915 5550 1916 5558
rect 1918 5550 1921 5558
rect 1923 5550 1928 5558
rect 1940 5550 1941 5558
rect 1943 5550 1944 5558
rect 1961 5550 1962 5558
rect 1964 5550 1966 5558
rect 1987 5550 1988 5558
rect 1990 5550 1993 5558
rect 1995 5550 2000 5558
rect 2015 5550 2016 5558
rect 2018 5550 2019 5558
rect 2031 5550 2032 5558
rect 2034 5550 2035 5558
rect 2056 5550 2057 5558
rect 2059 5550 2060 5558
rect 2064 5550 2070 5558
rect 2074 5550 2075 5558
rect 2077 5550 2078 5558
rect 2103 5555 2104 5563
rect 2106 5555 2109 5563
rect 2111 5555 2114 5563
rect 2158 5550 2159 5558
rect 2161 5550 2162 5558
rect 2176 5550 2177 5558
rect 2179 5550 2182 5558
rect 2184 5550 2189 5558
rect 2201 5550 2202 5558
rect 2204 5550 2205 5558
rect 2222 5550 2223 5558
rect 2225 5550 2227 5558
rect 2248 5550 2249 5558
rect 2251 5550 2254 5558
rect 2256 5550 2261 5558
rect 2276 5550 2277 5558
rect 2279 5550 2280 5558
rect 2292 5550 2293 5558
rect 2295 5550 2296 5558
rect 2308 5550 2309 5558
rect 2311 5550 2312 5558
rect 1472 5519 1473 5527
rect 1475 5519 1476 5527
rect 1488 5519 1489 5527
rect 1491 5519 1494 5527
rect 1496 5519 1497 5527
rect 1505 5523 1510 5527
rect 1509 5519 1510 5523
rect 1512 5519 1513 5527
rect 1525 5519 1526 5527
rect 1528 5519 1529 5527
rect 1546 5519 1547 5527
rect 1549 5519 1552 5527
rect 1554 5519 1555 5527
rect 1563 5523 1568 5527
rect 1567 5519 1568 5523
rect 1570 5519 1571 5527
rect 1583 5519 1584 5527
rect 1586 5519 1589 5527
rect 1591 5519 1592 5527
rect 1604 5519 1605 5527
rect 1607 5519 1608 5527
rect 1620 5519 1621 5527
rect 1623 5519 1626 5527
rect 1628 5519 1629 5527
rect 1637 5523 1642 5527
rect 1641 5519 1642 5523
rect 1644 5519 1645 5527
rect 1657 5519 1658 5527
rect 1660 5519 1661 5527
rect 1678 5519 1679 5527
rect 1681 5519 1684 5527
rect 1686 5519 1687 5527
rect 1695 5523 1700 5527
rect 1699 5519 1700 5523
rect 1702 5519 1703 5527
rect 1715 5519 1716 5527
rect 1718 5519 1721 5527
rect 1723 5519 1724 5527
rect 1736 5519 1737 5527
rect 1739 5519 1740 5527
rect 1752 5519 1753 5527
rect 1755 5519 1758 5527
rect 1760 5519 1761 5527
rect 1769 5523 1774 5527
rect 1773 5519 1774 5523
rect 1776 5519 1777 5527
rect 1789 5519 1790 5527
rect 1792 5519 1793 5527
rect 1810 5519 1811 5527
rect 1813 5519 1816 5527
rect 1818 5519 1819 5527
rect 1827 5523 1832 5527
rect 1831 5519 1832 5523
rect 1834 5519 1835 5527
rect 1847 5519 1848 5527
rect 1850 5519 1853 5527
rect 1855 5519 1856 5527
rect 2417 5519 2418 5527
rect 2420 5519 2421 5527
rect 2433 5519 2434 5527
rect 2436 5519 2439 5527
rect 2441 5519 2442 5527
rect 2450 5523 2455 5527
rect 2454 5519 2455 5523
rect 2457 5519 2458 5527
rect 2470 5519 2471 5527
rect 2473 5519 2474 5527
rect 2491 5519 2492 5527
rect 2494 5519 2497 5527
rect 2499 5519 2500 5527
rect 2508 5523 2513 5527
rect 2512 5519 2513 5523
rect 2515 5519 2516 5527
rect 2528 5519 2529 5527
rect 2531 5519 2534 5527
rect 2536 5519 2537 5527
rect 2549 5519 2550 5527
rect 2552 5519 2553 5527
rect 2565 5519 2566 5527
rect 2568 5519 2571 5527
rect 2573 5519 2574 5527
rect 2582 5523 2587 5527
rect 2586 5519 2587 5523
rect 2589 5519 2590 5527
rect 2602 5519 2603 5527
rect 2605 5519 2606 5527
rect 2623 5519 2624 5527
rect 2626 5519 2629 5527
rect 2631 5519 2632 5527
rect 2640 5523 2645 5527
rect 2644 5519 2645 5523
rect 2647 5519 2648 5527
rect 2660 5519 2661 5527
rect 2663 5519 2666 5527
rect 2668 5519 2669 5527
rect 2681 5519 2682 5527
rect 2684 5519 2685 5527
rect 2697 5519 2698 5527
rect 2700 5519 2703 5527
rect 2705 5519 2706 5527
rect 2714 5523 2719 5527
rect 2718 5519 2719 5523
rect 2721 5519 2722 5527
rect 2734 5519 2735 5527
rect 2737 5519 2738 5527
rect 2755 5519 2756 5527
rect 2758 5519 2761 5527
rect 2763 5519 2764 5527
rect 2772 5523 2777 5527
rect 2776 5519 2777 5523
rect 2779 5519 2780 5527
rect 2792 5519 2793 5527
rect 2795 5519 2798 5527
rect 2800 5519 2801 5527
rect 1135 5451 1136 5459
rect 1138 5451 1139 5459
rect 1158 5457 1159 5465
rect 1161 5457 1164 5465
rect 1166 5457 1169 5465
rect 1213 5464 1214 5472
rect 1216 5464 1217 5472
rect 1231 5464 1232 5472
rect 1234 5464 1237 5472
rect 1239 5464 1244 5472
rect 1256 5464 1257 5472
rect 1259 5464 1260 5472
rect 1277 5464 1278 5472
rect 1280 5464 1282 5472
rect 1303 5464 1304 5472
rect 1306 5464 1309 5472
rect 1311 5464 1316 5472
rect 1331 5464 1332 5472
rect 1334 5464 1335 5472
rect 1347 5464 1348 5472
rect 1350 5464 1351 5472
rect 1363 5464 1364 5472
rect 1366 5464 1367 5472
rect 1767 5448 1768 5456
rect 1770 5448 1773 5456
rect 1775 5448 1778 5456
rect 2080 5451 2081 5459
rect 2083 5451 2084 5459
rect 2103 5457 2104 5465
rect 2106 5457 2109 5465
rect 2111 5457 2114 5465
rect 2158 5464 2159 5472
rect 2161 5464 2162 5472
rect 2176 5464 2177 5472
rect 2179 5464 2182 5472
rect 2184 5464 2189 5472
rect 2201 5464 2202 5472
rect 2204 5464 2205 5472
rect 2222 5464 2223 5472
rect 2225 5464 2227 5472
rect 2248 5464 2249 5472
rect 2251 5464 2254 5472
rect 2256 5464 2261 5472
rect 2276 5464 2277 5472
rect 2279 5464 2280 5472
rect 2292 5464 2293 5472
rect 2295 5464 2296 5472
rect 2308 5464 2309 5472
rect 2311 5464 2312 5472
rect 987 5419 988 5427
rect 990 5419 993 5427
rect 995 5419 998 5427
rect 1077 5419 1078 5427
rect 1080 5419 1083 5427
rect 1085 5419 1088 5427
rect 1158 5419 1159 5427
rect 1161 5419 1164 5427
rect 1166 5419 1169 5427
rect 1213 5418 1214 5426
rect 1216 5418 1217 5426
rect 1231 5418 1232 5426
rect 1234 5418 1237 5426
rect 1239 5418 1244 5426
rect 1256 5418 1257 5426
rect 1259 5418 1260 5426
rect 1277 5418 1278 5426
rect 1280 5418 1282 5426
rect 1303 5418 1304 5426
rect 1306 5418 1309 5426
rect 1311 5418 1316 5426
rect 1331 5418 1332 5426
rect 1334 5418 1335 5426
rect 1347 5418 1348 5426
rect 1350 5418 1351 5426
rect 1363 5418 1364 5426
rect 1366 5418 1367 5426
rect 1932 5419 1933 5427
rect 1935 5419 1938 5427
rect 1940 5419 1943 5427
rect 2022 5419 2023 5427
rect 2025 5419 2028 5427
rect 2030 5419 2033 5427
rect 2103 5419 2104 5427
rect 2106 5419 2109 5427
rect 2111 5419 2114 5427
rect 2158 5418 2159 5426
rect 2161 5418 2162 5426
rect 2176 5418 2177 5426
rect 2179 5418 2182 5426
rect 2184 5418 2189 5426
rect 2201 5418 2202 5426
rect 2204 5418 2205 5426
rect 2222 5418 2223 5426
rect 2225 5418 2227 5426
rect 2248 5418 2249 5426
rect 2251 5418 2254 5426
rect 2256 5418 2261 5426
rect 2276 5418 2277 5426
rect 2279 5418 2280 5426
rect 2292 5418 2293 5426
rect 2295 5418 2296 5426
rect 2308 5418 2309 5426
rect 2311 5418 2312 5426
rect 964 5319 965 5327
rect 967 5319 968 5327
rect 987 5325 988 5333
rect 990 5325 993 5333
rect 995 5325 998 5333
rect 1018 5319 1019 5327
rect 1021 5319 1022 5327
rect 1054 5319 1055 5327
rect 1057 5319 1058 5327
rect 1077 5325 1078 5333
rect 1080 5325 1083 5333
rect 1085 5325 1088 5333
rect 1653 5349 1654 5379
rect 1656 5349 1657 5379
rect 1706 5349 1707 5379
rect 1709 5349 1710 5379
rect 1744 5346 1745 5354
rect 1747 5346 1748 5354
rect 1767 5352 1768 5360
rect 1770 5352 1773 5360
rect 1775 5352 1778 5360
rect 1798 5346 1799 5354
rect 1801 5346 1802 5354
rect 1820 5346 1821 5354
rect 1823 5346 1824 5354
rect 1108 5319 1109 5327
rect 1111 5319 1112 5327
rect 1135 5319 1136 5327
rect 1138 5319 1139 5327
rect 1158 5325 1159 5333
rect 1161 5325 1164 5333
rect 1166 5325 1169 5333
rect 1213 5332 1214 5340
rect 1216 5332 1217 5340
rect 1231 5332 1232 5340
rect 1234 5332 1237 5340
rect 1239 5332 1244 5340
rect 1256 5332 1257 5340
rect 1259 5332 1260 5340
rect 1277 5332 1278 5340
rect 1280 5332 1282 5340
rect 1303 5332 1304 5340
rect 1306 5332 1309 5340
rect 1311 5332 1316 5340
rect 1331 5332 1332 5340
rect 1334 5332 1335 5340
rect 1347 5332 1348 5340
rect 1350 5332 1351 5340
rect 1363 5332 1364 5340
rect 1366 5332 1367 5340
rect 1767 5318 1768 5326
rect 1770 5318 1773 5326
rect 1775 5318 1778 5326
rect 1909 5319 1910 5327
rect 1912 5319 1913 5327
rect 1932 5325 1933 5333
rect 1935 5325 1938 5333
rect 1940 5325 1943 5333
rect 1963 5319 1964 5327
rect 1966 5319 1967 5327
rect 1999 5319 2000 5327
rect 2002 5319 2003 5327
rect 2022 5325 2023 5333
rect 2025 5325 2028 5333
rect 2030 5325 2033 5333
rect 2053 5319 2054 5327
rect 2056 5319 2057 5327
rect 2080 5319 2081 5327
rect 2083 5319 2084 5327
rect 2103 5325 2104 5333
rect 2106 5325 2109 5333
rect 2111 5325 2114 5333
rect 2158 5332 2159 5340
rect 2161 5332 2162 5340
rect 2176 5332 2177 5340
rect 2179 5332 2182 5340
rect 2184 5332 2189 5340
rect 2201 5332 2202 5340
rect 2204 5332 2205 5340
rect 2222 5332 2223 5340
rect 2225 5332 2227 5340
rect 2248 5332 2249 5340
rect 2251 5332 2254 5340
rect 2256 5332 2261 5340
rect 2276 5332 2277 5340
rect 2279 5332 2280 5340
rect 2292 5332 2293 5340
rect 2295 5332 2296 5340
rect 2308 5332 2309 5340
rect 2311 5332 2312 5340
rect 1053 5284 1054 5292
rect 1056 5284 1059 5292
rect 1061 5284 1064 5292
rect 1158 5284 1159 5292
rect 1161 5284 1164 5292
rect 1166 5284 1169 5292
rect 1213 5286 1214 5294
rect 1216 5286 1217 5294
rect 1231 5286 1232 5294
rect 1234 5286 1237 5294
rect 1239 5286 1244 5294
rect 1256 5286 1257 5294
rect 1259 5286 1260 5294
rect 1277 5286 1278 5294
rect 1280 5286 1282 5294
rect 1303 5286 1304 5294
rect 1306 5286 1309 5294
rect 1311 5286 1316 5294
rect 1331 5286 1332 5294
rect 1334 5286 1335 5294
rect 1347 5286 1348 5294
rect 1350 5286 1351 5294
rect 1363 5286 1364 5294
rect 1366 5286 1367 5294
rect 1998 5284 1999 5292
rect 2001 5284 2004 5292
rect 2006 5284 2009 5292
rect 2103 5284 2104 5292
rect 2106 5284 2109 5292
rect 2111 5284 2114 5292
rect 2158 5286 2159 5294
rect 2161 5286 2162 5294
rect 2176 5286 2177 5294
rect 2179 5286 2182 5294
rect 2184 5286 2189 5294
rect 2201 5286 2202 5294
rect 2204 5286 2205 5294
rect 2222 5286 2223 5294
rect 2225 5286 2227 5294
rect 2248 5286 2249 5294
rect 2251 5286 2254 5294
rect 2256 5286 2261 5294
rect 2276 5286 2277 5294
rect 2279 5286 2280 5294
rect 2292 5286 2293 5294
rect 2295 5286 2296 5294
rect 2308 5286 2309 5294
rect 2311 5286 2312 5294
rect 1030 5187 1031 5195
rect 1033 5187 1034 5195
rect 1053 5193 1054 5201
rect 1056 5193 1059 5201
rect 1061 5193 1064 5201
rect 1559 5219 1560 5249
rect 1562 5219 1563 5249
rect 1612 5219 1613 5249
rect 1615 5219 1616 5249
rect 1744 5216 1745 5224
rect 1747 5216 1748 5224
rect 1767 5222 1768 5230
rect 1770 5222 1773 5230
rect 1775 5222 1778 5230
rect 1798 5216 1799 5224
rect 1801 5216 1802 5224
rect 1084 5187 1085 5195
rect 1087 5187 1088 5195
rect 1135 5187 1136 5195
rect 1138 5187 1139 5195
rect 1158 5193 1159 5201
rect 1161 5193 1164 5201
rect 1166 5193 1169 5201
rect 1213 5200 1214 5208
rect 1216 5200 1217 5208
rect 1231 5200 1232 5208
rect 1234 5200 1237 5208
rect 1239 5200 1244 5208
rect 1256 5200 1257 5208
rect 1259 5200 1260 5208
rect 1277 5200 1278 5208
rect 1280 5200 1282 5208
rect 1303 5200 1304 5208
rect 1306 5200 1309 5208
rect 1311 5200 1316 5208
rect 1331 5200 1332 5208
rect 1334 5200 1335 5208
rect 1347 5200 1348 5208
rect 1350 5200 1351 5208
rect 1363 5200 1364 5208
rect 1366 5200 1367 5208
rect 1975 5187 1976 5195
rect 1978 5187 1979 5195
rect 1998 5193 1999 5201
rect 2001 5193 2004 5201
rect 2006 5193 2009 5201
rect 2029 5187 2030 5195
rect 2032 5187 2033 5195
rect 2080 5187 2081 5195
rect 2083 5187 2084 5195
rect 2103 5193 2104 5201
rect 2106 5193 2109 5201
rect 2111 5193 2114 5201
rect 2158 5200 2159 5208
rect 2161 5200 2162 5208
rect 2176 5200 2177 5208
rect 2179 5200 2182 5208
rect 2184 5200 2189 5208
rect 2201 5200 2202 5208
rect 2204 5200 2205 5208
rect 2222 5200 2223 5208
rect 2225 5200 2227 5208
rect 2248 5200 2249 5208
rect 2251 5200 2254 5208
rect 2256 5200 2261 5208
rect 2276 5200 2277 5208
rect 2279 5200 2280 5208
rect 2292 5200 2293 5208
rect 2295 5200 2296 5208
rect 2308 5200 2309 5208
rect 2311 5200 2312 5208
rect 1077 5153 1078 5161
rect 1080 5153 1083 5161
rect 1085 5153 1088 5161
rect 1158 5153 1159 5161
rect 1161 5153 1164 5161
rect 1166 5153 1169 5161
rect 1213 5154 1214 5162
rect 1216 5154 1217 5162
rect 1231 5154 1232 5162
rect 1234 5154 1237 5162
rect 1239 5154 1244 5162
rect 1256 5154 1257 5162
rect 1259 5154 1260 5162
rect 1277 5154 1278 5162
rect 1280 5154 1282 5162
rect 1303 5154 1304 5162
rect 1306 5154 1309 5162
rect 1311 5154 1316 5162
rect 1331 5154 1332 5162
rect 1334 5154 1335 5162
rect 1347 5154 1348 5162
rect 1350 5154 1351 5162
rect 1363 5154 1364 5162
rect 1366 5154 1367 5162
rect 2022 5153 2023 5161
rect 2025 5153 2028 5161
rect 2030 5153 2033 5161
rect 2103 5153 2104 5161
rect 2106 5153 2109 5161
rect 2111 5153 2114 5161
rect 2158 5154 2159 5162
rect 2161 5154 2162 5162
rect 2176 5154 2177 5162
rect 2179 5154 2182 5162
rect 2184 5154 2189 5162
rect 2201 5154 2202 5162
rect 2204 5154 2205 5162
rect 2222 5154 2223 5162
rect 2225 5154 2227 5162
rect 2248 5154 2249 5162
rect 2251 5154 2254 5162
rect 2256 5154 2261 5162
rect 2276 5154 2277 5162
rect 2279 5154 2280 5162
rect 2292 5154 2293 5162
rect 2295 5154 2296 5162
rect 2308 5154 2309 5162
rect 2311 5154 2312 5162
rect 1613 5119 1614 5127
rect 1616 5119 1619 5127
rect 1621 5119 1622 5127
rect 1634 5119 1635 5127
rect 1637 5123 1642 5127
rect 1637 5119 1638 5123
rect 1650 5119 1651 5127
rect 1653 5119 1656 5127
rect 1658 5119 1659 5127
rect 1676 5119 1677 5127
rect 1679 5119 1680 5127
rect 1692 5119 1693 5127
rect 1695 5123 1700 5127
rect 1695 5119 1696 5123
rect 1708 5119 1709 5127
rect 1711 5119 1714 5127
rect 1716 5119 1717 5127
rect 1729 5119 1730 5127
rect 1732 5119 1733 5127
rect 2558 5119 2559 5127
rect 2561 5119 2564 5127
rect 2566 5119 2567 5127
rect 2579 5119 2580 5127
rect 2582 5123 2587 5127
rect 2582 5119 2583 5123
rect 2595 5119 2596 5127
rect 2598 5119 2601 5127
rect 2603 5119 2604 5127
rect 2621 5119 2622 5127
rect 2624 5119 2625 5127
rect 2637 5119 2638 5127
rect 2640 5123 2645 5127
rect 2640 5119 2641 5123
rect 2653 5119 2654 5127
rect 2656 5119 2659 5127
rect 2661 5119 2662 5127
rect 2674 5119 2675 5127
rect 2677 5119 2678 5127
rect 1054 5055 1055 5063
rect 1057 5055 1058 5063
rect 1077 5061 1078 5069
rect 1080 5061 1083 5069
rect 1085 5061 1088 5069
rect 1108 5055 1109 5063
rect 1111 5055 1112 5063
rect 1135 5055 1136 5063
rect 1138 5055 1139 5063
rect 1158 5061 1159 5069
rect 1161 5061 1164 5069
rect 1166 5061 1169 5069
rect 1213 5068 1214 5076
rect 1216 5068 1217 5076
rect 1231 5068 1232 5076
rect 1234 5068 1237 5076
rect 1239 5068 1244 5076
rect 1256 5068 1257 5076
rect 1259 5068 1260 5076
rect 1277 5068 1278 5076
rect 1280 5068 1282 5076
rect 1303 5068 1304 5076
rect 1306 5068 1309 5076
rect 1311 5068 1316 5076
rect 1331 5068 1332 5076
rect 1334 5068 1335 5076
rect 1347 5068 1348 5076
rect 1350 5068 1351 5076
rect 1363 5068 1364 5076
rect 1366 5068 1367 5076
rect 1189 5055 1190 5063
rect 1192 5055 1193 5063
rect 1999 5055 2000 5063
rect 2002 5055 2003 5063
rect 2022 5061 2023 5069
rect 2025 5061 2028 5069
rect 2030 5061 2033 5069
rect 2053 5055 2054 5063
rect 2056 5055 2057 5063
rect 2080 5055 2081 5063
rect 2083 5055 2084 5063
rect 2103 5061 2104 5069
rect 2106 5061 2109 5069
rect 2111 5061 2114 5069
rect 2158 5068 2159 5076
rect 2161 5068 2162 5076
rect 2176 5068 2177 5076
rect 2179 5068 2182 5076
rect 2184 5068 2189 5076
rect 2201 5068 2202 5076
rect 2204 5068 2205 5076
rect 2222 5068 2223 5076
rect 2225 5068 2227 5076
rect 2248 5068 2249 5076
rect 2251 5068 2254 5076
rect 2256 5068 2261 5076
rect 2276 5068 2277 5076
rect 2279 5068 2280 5076
rect 2292 5068 2293 5076
rect 2295 5068 2296 5076
rect 2308 5068 2309 5076
rect 2311 5068 2312 5076
rect 2134 5055 2135 5063
rect 2137 5055 2138 5063
rect 1604 5017 1605 5025
rect 1607 5017 1608 5025
rect 1620 5017 1621 5025
rect 1623 5017 1626 5025
rect 1628 5017 1629 5025
rect 1637 5021 1642 5025
rect 1641 5017 1642 5021
rect 1644 5017 1645 5025
rect 1657 5017 1658 5025
rect 1660 5017 1661 5025
rect 1678 5017 1679 5025
rect 1681 5017 1684 5025
rect 1686 5017 1687 5025
rect 1695 5021 1700 5025
rect 1699 5017 1700 5021
rect 1702 5017 1703 5025
rect 1715 5017 1716 5025
rect 1718 5017 1721 5025
rect 1723 5017 1724 5025
rect 2549 5017 2550 5025
rect 2552 5017 2553 5025
rect 2565 5017 2566 5025
rect 2568 5017 2571 5025
rect 2573 5017 2574 5025
rect 2582 5021 2587 5025
rect 2586 5017 2587 5021
rect 2589 5017 2590 5025
rect 2602 5017 2603 5025
rect 2605 5017 2606 5025
rect 2623 5017 2624 5025
rect 2626 5017 2629 5025
rect 2631 5017 2632 5025
rect 2640 5021 2645 5025
rect 2644 5017 2645 5021
rect 2647 5017 2648 5025
rect 2660 5017 2661 5025
rect 2663 5017 2666 5025
rect 2668 5017 2669 5025
rect 856 4984 857 4992
rect 859 4984 860 4992
rect 872 4984 873 4992
rect 875 4984 878 4992
rect 880 4984 881 4992
rect 889 4988 894 4992
rect 893 4984 894 4988
rect 896 4984 897 4992
rect 909 4984 910 4992
rect 912 4984 913 4992
rect 930 4984 931 4992
rect 933 4984 936 4992
rect 938 4984 939 4992
rect 947 4988 952 4992
rect 951 4984 952 4988
rect 954 4984 955 4992
rect 967 4984 968 4992
rect 970 4984 973 4992
rect 975 4984 976 4992
rect 988 4984 989 4992
rect 991 4984 992 4992
rect 1004 4984 1005 4992
rect 1007 4984 1010 4992
rect 1012 4984 1013 4992
rect 1021 4988 1026 4992
rect 1025 4984 1026 4988
rect 1028 4984 1029 4992
rect 1041 4984 1042 4992
rect 1044 4984 1045 4992
rect 1062 4984 1063 4992
rect 1065 4984 1068 4992
rect 1070 4984 1071 4992
rect 1079 4988 1084 4992
rect 1083 4984 1084 4988
rect 1086 4984 1087 4992
rect 1099 4984 1100 4992
rect 1102 4984 1105 4992
rect 1107 4984 1108 4992
rect 1120 4984 1121 4992
rect 1123 4984 1124 4992
rect 1136 4984 1137 4992
rect 1139 4984 1142 4992
rect 1144 4984 1145 4992
rect 1153 4988 1158 4992
rect 1157 4984 1158 4988
rect 1160 4984 1161 4992
rect 1173 4984 1174 4992
rect 1176 4984 1177 4992
rect 1194 4984 1195 4992
rect 1197 4984 1200 4992
rect 1202 4984 1203 4992
rect 1211 4988 1216 4992
rect 1215 4984 1216 4988
rect 1218 4984 1219 4992
rect 1231 4984 1232 4992
rect 1234 4984 1237 4992
rect 1239 4984 1240 4992
rect 1252 4984 1253 4992
rect 1255 4984 1256 4992
rect 1268 4984 1269 4992
rect 1271 4984 1274 4992
rect 1276 4984 1277 4992
rect 1285 4988 1290 4992
rect 1289 4984 1290 4988
rect 1292 4984 1293 4992
rect 1305 4984 1306 4992
rect 1308 4984 1309 4992
rect 1326 4984 1327 4992
rect 1329 4984 1332 4992
rect 1334 4984 1335 4992
rect 1343 4988 1348 4992
rect 1347 4984 1348 4988
rect 1350 4984 1351 4992
rect 1363 4984 1364 4992
rect 1366 4984 1369 4992
rect 1371 4984 1372 4992
rect 1801 4984 1802 4992
rect 1804 4984 1805 4992
rect 1817 4984 1818 4992
rect 1820 4984 1823 4992
rect 1825 4984 1826 4992
rect 1834 4988 1839 4992
rect 1838 4984 1839 4988
rect 1841 4984 1842 4992
rect 1854 4984 1855 4992
rect 1857 4984 1858 4992
rect 1875 4984 1876 4992
rect 1878 4984 1881 4992
rect 1883 4984 1884 4992
rect 1892 4988 1897 4992
rect 1896 4984 1897 4988
rect 1899 4984 1900 4992
rect 1912 4984 1913 4992
rect 1915 4984 1918 4992
rect 1920 4984 1921 4992
rect 1933 4984 1934 4992
rect 1936 4984 1937 4992
rect 1949 4984 1950 4992
rect 1952 4984 1955 4992
rect 1957 4984 1958 4992
rect 1966 4988 1971 4992
rect 1970 4984 1971 4988
rect 1973 4984 1974 4992
rect 1986 4984 1987 4992
rect 1989 4984 1990 4992
rect 2007 4984 2008 4992
rect 2010 4984 2013 4992
rect 2015 4984 2016 4992
rect 2024 4988 2029 4992
rect 2028 4984 2029 4988
rect 2031 4984 2032 4992
rect 2044 4984 2045 4992
rect 2047 4984 2050 4992
rect 2052 4984 2053 4992
rect 2065 4984 2066 4992
rect 2068 4984 2069 4992
rect 2081 4984 2082 4992
rect 2084 4984 2087 4992
rect 2089 4984 2090 4992
rect 2098 4988 2103 4992
rect 2102 4984 2103 4988
rect 2105 4984 2106 4992
rect 2118 4984 2119 4992
rect 2121 4984 2122 4992
rect 2139 4984 2140 4992
rect 2142 4984 2145 4992
rect 2147 4984 2148 4992
rect 2156 4988 2161 4992
rect 2160 4984 2161 4988
rect 2163 4984 2164 4992
rect 2176 4984 2177 4992
rect 2179 4984 2182 4992
rect 2184 4984 2185 4992
rect 2197 4984 2198 4992
rect 2200 4984 2201 4992
rect 2213 4984 2214 4992
rect 2216 4984 2219 4992
rect 2221 4984 2222 4992
rect 2230 4988 2235 4992
rect 2234 4984 2235 4988
rect 2237 4984 2238 4992
rect 2250 4984 2251 4992
rect 2253 4984 2254 4992
rect 2271 4984 2272 4992
rect 2274 4984 2277 4992
rect 2279 4984 2280 4992
rect 2288 4988 2293 4992
rect 2292 4984 2293 4988
rect 2295 4984 2296 4992
rect 2308 4984 2309 4992
rect 2311 4984 2314 4992
rect 2316 4984 2317 4992
rect 4578 7928 4579 7945
rect 4574 7924 4579 7928
rect 4578 7889 4579 7924
rect 4581 7889 4582 7945
rect 4586 7889 4587 7945
rect 4589 7928 4590 7945
rect 4594 7928 4595 7945
rect 4589 7924 4595 7928
rect 4589 7889 4590 7924
rect 4594 7889 4595 7924
rect 4597 7889 4598 7945
rect 4602 7889 4603 7945
rect 4605 7928 4606 7945
rect 4610 7928 4611 7945
rect 4605 7924 4611 7928
rect 4605 7889 4606 7924
rect 4610 7889 4611 7924
rect 4613 7889 4614 7945
rect 4618 7889 4619 7945
rect 4621 7928 4622 7945
rect 4626 7928 4627 7945
rect 4621 7924 4627 7928
rect 4621 7889 4622 7924
rect 4626 7889 4627 7924
rect 4631 7857 4634 7945
rect 4636 7857 4637 7945
rect 4641 7857 4642 7945
rect 4644 7936 4650 7945
rect 4644 7928 4645 7936
rect 4649 7928 4650 7936
rect 4644 7924 4650 7928
rect 4644 7857 4645 7924
rect 4649 7857 4650 7924
rect 4652 7857 4653 7945
rect 4657 7857 4658 7945
rect 4660 7928 4661 7945
rect 4665 7928 4666 7945
rect 4660 7924 4666 7928
rect 4660 7857 4661 7924
rect 4665 7857 4666 7924
rect 4674 7857 4677 7945
rect 4679 7857 4680 7945
rect 4684 7857 4685 7945
rect 4687 7936 4693 7945
rect 4687 7928 4688 7936
rect 4692 7928 4693 7936
rect 4687 7924 4693 7928
rect 4687 7857 4688 7924
rect 4692 7857 4693 7924
rect 4695 7857 4696 7945
rect 4700 7857 4701 7945
rect 4703 7928 4704 7945
rect 4708 7928 4709 7945
rect 4703 7924 4709 7928
rect 4703 7857 4704 7924
rect 4708 7857 4709 7924
rect 4713 7857 4718 7945
rect 4720 7857 4721 7945
rect 4725 7857 4726 7945
rect 4728 7936 4734 7945
rect 4728 7928 4729 7936
rect 4733 7928 4734 7936
rect 4728 7924 4734 7928
rect 4728 7857 4729 7924
rect 4733 7857 4734 7924
rect 4736 7857 4737 7945
rect 4741 7857 4742 7945
rect 4744 7928 4745 7945
rect 4749 7928 4750 7945
rect 4744 7924 4750 7928
rect 4744 7857 4745 7924
rect 4749 7857 4750 7924
rect 4576 7393 4577 7428
rect 4572 7389 4577 7393
rect 4576 7372 4577 7389
rect 4579 7372 4580 7428
rect 4584 7372 4585 7428
rect 4587 7393 4588 7428
rect 4592 7393 4593 7428
rect 4587 7389 4593 7393
rect 4587 7372 4588 7389
rect 4592 7372 4593 7389
rect 4595 7372 4596 7428
rect 4600 7372 4601 7428
rect 4603 7393 4604 7428
rect 4608 7393 4609 7428
rect 4603 7389 4609 7393
rect 4603 7372 4604 7389
rect 4608 7372 4609 7389
rect 4611 7372 4612 7428
rect 4616 7372 4617 7428
rect 4619 7393 4620 7428
rect 4619 7389 4624 7393
rect 4619 7372 4620 7389
rect 4657 7305 4746 7306
rect 4661 7301 4667 7305
rect 4671 7301 4677 7305
rect 4681 7301 4687 7305
rect 4691 7301 4697 7305
rect 4701 7301 4707 7305
rect 4711 7301 4717 7305
rect 4721 7301 4727 7305
rect 4731 7301 4737 7305
rect 4741 7301 4746 7305
rect 4657 7300 4746 7301
rect 4657 7296 4662 7300
rect 4666 7296 4672 7300
rect 4676 7296 4682 7300
rect 4686 7296 4692 7300
rect 4696 7296 4702 7300
rect 4706 7296 4712 7300
rect 4716 7296 4722 7300
rect 4726 7296 4732 7300
rect 4736 7296 4742 7300
rect 4657 7295 4746 7296
rect 4661 7291 4667 7295
rect 4671 7291 4677 7295
rect 4681 7291 4687 7295
rect 4691 7291 4697 7295
rect 4701 7291 4707 7295
rect 4711 7291 4717 7295
rect 4721 7291 4727 7295
rect 4731 7291 4737 7295
rect 4741 7291 4746 7295
rect 4657 7290 4746 7291
rect 4657 7286 4662 7290
rect 4666 7286 4672 7290
rect 4676 7286 4682 7290
rect 4686 7286 4692 7290
rect 4696 7286 4702 7290
rect 4706 7286 4712 7290
rect 4716 7286 4722 7290
rect 4726 7286 4732 7290
rect 4736 7286 4742 7290
rect 4657 7285 4746 7286
rect 4661 7281 4667 7285
rect 4671 7281 4677 7285
rect 4681 7281 4687 7285
rect 4691 7281 4697 7285
rect 4701 7281 4707 7285
rect 4711 7281 4717 7285
rect 4721 7281 4727 7285
rect 4731 7281 4737 7285
rect 4741 7281 4746 7285
rect 4657 7280 4746 7281
rect 4657 7276 4662 7280
rect 4666 7276 4672 7280
rect 4676 7276 4682 7280
rect 4686 7276 4692 7280
rect 4696 7276 4702 7280
rect 4706 7276 4712 7280
rect 4716 7276 4722 7280
rect 4726 7276 4732 7280
rect 4736 7276 4742 7280
rect 4657 7275 4746 7276
rect 4661 7271 4667 7275
rect 4671 7271 4677 7275
rect 4681 7271 4687 7275
rect 4691 7271 4697 7275
rect 4701 7271 4707 7275
rect 4711 7271 4717 7275
rect 4721 7271 4727 7275
rect 4731 7271 4737 7275
rect 4741 7271 4746 7275
rect 4657 7270 4746 7271
rect 4657 7266 4662 7270
rect 4666 7266 4672 7270
rect 4676 7266 4682 7270
rect 4686 7266 4692 7270
rect 4696 7266 4702 7270
rect 4706 7266 4712 7270
rect 4716 7266 4722 7270
rect 4726 7266 4732 7270
rect 4736 7266 4742 7270
rect 4657 7265 4746 7266
rect 4661 7261 4667 7265
rect 4671 7261 4677 7265
rect 4681 7261 4687 7265
rect 4691 7261 4697 7265
rect 4701 7261 4707 7265
rect 4711 7261 4717 7265
rect 4721 7261 4727 7265
rect 4731 7261 4737 7265
rect 4741 7261 4746 7265
rect 1227 4531 1231 4535
rect 1210 4530 1266 4531
rect 2154 4531 2158 4535
rect 2137 4530 2193 4531
rect 2463 4531 2467 4535
rect 2446 4530 2502 4531
rect 2772 4531 2776 4535
rect 2755 4530 2811 4531
rect 3081 4531 3085 4535
rect 3064 4530 3120 4531
rect 3390 4531 3394 4535
rect 3373 4530 3429 4531
rect 1210 4527 1266 4528
rect 1210 4522 1266 4523
rect 1210 4519 1266 4520
rect 1227 4515 1231 4519
rect 1210 4514 1266 4515
rect 1210 4511 1266 4512
rect 1210 4506 1266 4507
rect 2137 4527 2193 4528
rect 2137 4522 2193 4523
rect 2137 4519 2193 4520
rect 2154 4515 2158 4519
rect 2137 4514 2193 4515
rect 2137 4511 2193 4512
rect 2137 4506 2193 4507
rect 1210 4503 1266 4504
rect 1227 4499 1231 4503
rect 1210 4498 1266 4499
rect 2446 4527 2502 4528
rect 2446 4522 2502 4523
rect 2446 4519 2502 4520
rect 2463 4515 2467 4519
rect 2446 4514 2502 4515
rect 2446 4511 2502 4512
rect 2446 4506 2502 4507
rect 2137 4503 2193 4504
rect 2154 4499 2158 4503
rect 2137 4498 2193 4499
rect 2755 4527 2811 4528
rect 2755 4522 2811 4523
rect 2755 4519 2811 4520
rect 2772 4515 2776 4519
rect 2755 4514 2811 4515
rect 2755 4511 2811 4512
rect 2755 4506 2811 4507
rect 2446 4503 2502 4504
rect 2463 4499 2467 4503
rect 2446 4498 2502 4499
rect 3064 4527 3120 4528
rect 3064 4522 3120 4523
rect 3064 4519 3120 4520
rect 3081 4515 3085 4519
rect 3064 4514 3120 4515
rect 3064 4511 3120 4512
rect 3064 4506 3120 4507
rect 2755 4503 2811 4504
rect 2772 4499 2776 4503
rect 2755 4498 2811 4499
rect 3373 4527 3429 4528
rect 3373 4522 3429 4523
rect 3373 4519 3429 4520
rect 3390 4515 3394 4519
rect 3373 4514 3429 4515
rect 3373 4511 3429 4512
rect 3373 4506 3429 4507
rect 3064 4503 3120 4504
rect 3081 4499 3085 4503
rect 3064 4498 3120 4499
rect 3373 4503 3429 4504
rect 3390 4499 3394 4503
rect 3373 4498 3429 4499
rect 1210 4495 1266 4496
rect 1210 4490 1266 4491
rect 2137 4495 2193 4496
rect 2137 4490 2193 4491
rect 2446 4495 2502 4496
rect 2446 4490 2502 4491
rect 2755 4495 2811 4496
rect 2755 4490 2811 4491
rect 3064 4495 3120 4496
rect 3064 4490 3120 4491
rect 3373 4495 3429 4496
rect 3373 4490 3429 4491
rect 1210 4487 1266 4488
rect 1227 4483 1231 4487
rect 2137 4487 2193 4488
rect 2154 4483 2158 4487
rect 2446 4487 2502 4488
rect 2463 4483 2467 4487
rect 2755 4487 2811 4488
rect 2772 4483 2776 4487
rect 3064 4487 3120 4488
rect 3081 4483 3085 4487
rect 3373 4487 3429 4488
rect 3390 4483 3394 4487
rect 1103 4446 1109 4450
rect 1113 4446 1119 4450
rect 1123 4446 1129 4450
rect 1133 4446 1139 4450
rect 1143 4446 1144 4450
rect 1099 4445 1144 4446
rect 1099 4441 1104 4445
rect 1108 4441 1114 4445
rect 1118 4441 1124 4445
rect 1128 4441 1134 4445
rect 1138 4441 1144 4445
rect 1099 4440 1144 4441
rect 1103 4436 1109 4440
rect 1113 4436 1119 4440
rect 1123 4436 1129 4440
rect 1133 4436 1139 4440
rect 1143 4436 1144 4440
rect 1099 4435 1144 4436
rect 1099 4431 1104 4435
rect 1108 4431 1114 4435
rect 1118 4431 1124 4435
rect 1128 4431 1134 4435
rect 1138 4431 1144 4435
rect 1099 4430 1144 4431
rect 1103 4426 1109 4430
rect 1113 4426 1119 4430
rect 1123 4426 1129 4430
rect 1133 4426 1139 4430
rect 1143 4426 1144 4430
rect 1099 4425 1144 4426
rect 1099 4421 1104 4425
rect 1108 4421 1114 4425
rect 1118 4421 1124 4425
rect 1128 4421 1134 4425
rect 1138 4421 1144 4425
rect 1099 4420 1144 4421
rect 1103 4416 1109 4420
rect 1113 4416 1119 4420
rect 1123 4416 1129 4420
rect 1133 4416 1139 4420
rect 1143 4416 1144 4420
rect 1099 4415 1144 4416
rect 1099 4411 1104 4415
rect 1108 4411 1114 4415
rect 1118 4411 1124 4415
rect 1128 4411 1134 4415
rect 1138 4411 1144 4415
rect 1099 4410 1144 4411
rect 1103 4406 1109 4410
rect 1113 4406 1119 4410
rect 1123 4406 1129 4410
rect 1133 4406 1139 4410
rect 1143 4406 1144 4410
rect 1099 4405 1144 4406
rect 1099 4401 1104 4405
rect 1108 4401 1114 4405
rect 1118 4401 1124 4405
rect 1128 4401 1134 4405
rect 1138 4401 1144 4405
rect 1099 4400 1144 4401
rect 1103 4396 1109 4400
rect 1113 4396 1119 4400
rect 1123 4396 1129 4400
rect 1133 4396 1139 4400
rect 1143 4396 1144 4400
rect 1099 4395 1144 4396
rect 1099 4391 1104 4395
rect 1108 4391 1114 4395
rect 1118 4391 1124 4395
rect 1128 4391 1134 4395
rect 1138 4391 1144 4395
rect 1099 4390 1144 4391
rect 1103 4386 1109 4390
rect 1113 4386 1119 4390
rect 1123 4386 1129 4390
rect 1133 4386 1139 4390
rect 1143 4386 1144 4390
rect 1099 4385 1144 4386
rect 1099 4381 1104 4385
rect 1108 4381 1114 4385
rect 1118 4381 1124 4385
rect 1128 4381 1134 4385
rect 1138 4381 1144 4385
rect 1099 4380 1144 4381
rect 1103 4376 1109 4380
rect 1113 4376 1119 4380
rect 1123 4376 1129 4380
rect 1133 4376 1139 4380
rect 1143 4376 1144 4380
rect 1099 4375 1144 4376
rect 1099 4371 1104 4375
rect 1108 4371 1114 4375
rect 1118 4371 1124 4375
rect 1128 4371 1134 4375
rect 1138 4371 1144 4375
rect 1099 4370 1144 4371
rect 1103 4366 1109 4370
rect 1113 4366 1119 4370
rect 1123 4366 1129 4370
rect 1133 4366 1139 4370
rect 1143 4366 1144 4370
rect 1099 4365 1144 4366
rect 1099 4361 1104 4365
rect 1108 4361 1114 4365
rect 1118 4361 1124 4365
rect 1128 4361 1134 4365
rect 1138 4361 1144 4365
rect 1412 4446 1418 4450
rect 1422 4446 1428 4450
rect 1432 4446 1438 4450
rect 1442 4446 1448 4450
rect 1452 4446 1453 4450
rect 1408 4445 1453 4446
rect 1408 4441 1413 4445
rect 1417 4441 1423 4445
rect 1427 4441 1433 4445
rect 1437 4441 1443 4445
rect 1447 4441 1453 4445
rect 1408 4440 1453 4441
rect 1412 4436 1418 4440
rect 1422 4436 1428 4440
rect 1432 4436 1438 4440
rect 1442 4436 1448 4440
rect 1452 4436 1453 4440
rect 1408 4435 1453 4436
rect 1408 4431 1413 4435
rect 1417 4431 1423 4435
rect 1427 4431 1433 4435
rect 1437 4431 1443 4435
rect 1447 4431 1453 4435
rect 1408 4430 1453 4431
rect 1412 4426 1418 4430
rect 1422 4426 1428 4430
rect 1432 4426 1438 4430
rect 1442 4426 1448 4430
rect 1452 4426 1453 4430
rect 1408 4425 1453 4426
rect 1408 4421 1413 4425
rect 1417 4421 1423 4425
rect 1427 4421 1433 4425
rect 1437 4421 1443 4425
rect 1447 4421 1453 4425
rect 1408 4420 1453 4421
rect 1412 4416 1418 4420
rect 1422 4416 1428 4420
rect 1432 4416 1438 4420
rect 1442 4416 1448 4420
rect 1452 4416 1453 4420
rect 1408 4415 1453 4416
rect 1408 4411 1413 4415
rect 1417 4411 1423 4415
rect 1427 4411 1433 4415
rect 1437 4411 1443 4415
rect 1447 4411 1453 4415
rect 1408 4410 1453 4411
rect 1412 4406 1418 4410
rect 1422 4406 1428 4410
rect 1432 4406 1438 4410
rect 1442 4406 1448 4410
rect 1452 4406 1453 4410
rect 1408 4405 1453 4406
rect 1408 4401 1413 4405
rect 1417 4401 1423 4405
rect 1427 4401 1433 4405
rect 1437 4401 1443 4405
rect 1447 4401 1453 4405
rect 1408 4400 1453 4401
rect 1412 4396 1418 4400
rect 1422 4396 1428 4400
rect 1432 4396 1438 4400
rect 1442 4396 1448 4400
rect 1452 4396 1453 4400
rect 1408 4395 1453 4396
rect 1408 4391 1413 4395
rect 1417 4391 1423 4395
rect 1427 4391 1433 4395
rect 1437 4391 1443 4395
rect 1447 4391 1453 4395
rect 1408 4390 1453 4391
rect 1412 4386 1418 4390
rect 1422 4386 1428 4390
rect 1432 4386 1438 4390
rect 1442 4386 1448 4390
rect 1452 4386 1453 4390
rect 1408 4385 1453 4386
rect 1408 4381 1413 4385
rect 1417 4381 1423 4385
rect 1427 4381 1433 4385
rect 1437 4381 1443 4385
rect 1447 4381 1453 4385
rect 1408 4380 1453 4381
rect 1412 4376 1418 4380
rect 1422 4376 1428 4380
rect 1432 4376 1438 4380
rect 1442 4376 1448 4380
rect 1452 4376 1453 4380
rect 1408 4375 1453 4376
rect 1408 4371 1413 4375
rect 1417 4371 1423 4375
rect 1427 4371 1433 4375
rect 1437 4371 1443 4375
rect 1447 4371 1453 4375
rect 1408 4370 1453 4371
rect 1412 4366 1418 4370
rect 1422 4366 1428 4370
rect 1432 4366 1438 4370
rect 1442 4366 1448 4370
rect 1452 4366 1453 4370
rect 1408 4365 1453 4366
rect 1408 4361 1413 4365
rect 1417 4361 1423 4365
rect 1427 4361 1433 4365
rect 1437 4361 1443 4365
rect 1447 4361 1453 4365
rect 1721 4446 1727 4450
rect 1731 4446 1737 4450
rect 1741 4446 1747 4450
rect 1751 4446 1757 4450
rect 1761 4446 1762 4450
rect 1717 4445 1762 4446
rect 1717 4441 1722 4445
rect 1726 4441 1732 4445
rect 1736 4441 1742 4445
rect 1746 4441 1752 4445
rect 1756 4441 1762 4445
rect 1717 4440 1762 4441
rect 1721 4436 1727 4440
rect 1731 4436 1737 4440
rect 1741 4436 1747 4440
rect 1751 4436 1757 4440
rect 1761 4436 1762 4440
rect 1717 4435 1762 4436
rect 1717 4431 1722 4435
rect 1726 4431 1732 4435
rect 1736 4431 1742 4435
rect 1746 4431 1752 4435
rect 1756 4431 1762 4435
rect 1717 4430 1762 4431
rect 1721 4426 1727 4430
rect 1731 4426 1737 4430
rect 1741 4426 1747 4430
rect 1751 4426 1757 4430
rect 1761 4426 1762 4430
rect 1717 4425 1762 4426
rect 1717 4421 1722 4425
rect 1726 4421 1732 4425
rect 1736 4421 1742 4425
rect 1746 4421 1752 4425
rect 1756 4421 1762 4425
rect 1717 4420 1762 4421
rect 1721 4416 1727 4420
rect 1731 4416 1737 4420
rect 1741 4416 1747 4420
rect 1751 4416 1757 4420
rect 1761 4416 1762 4420
rect 1717 4415 1762 4416
rect 1717 4411 1722 4415
rect 1726 4411 1732 4415
rect 1736 4411 1742 4415
rect 1746 4411 1752 4415
rect 1756 4411 1762 4415
rect 1717 4410 1762 4411
rect 1721 4406 1727 4410
rect 1731 4406 1737 4410
rect 1741 4406 1747 4410
rect 1751 4406 1757 4410
rect 1761 4406 1762 4410
rect 1717 4405 1762 4406
rect 1717 4401 1722 4405
rect 1726 4401 1732 4405
rect 1736 4401 1742 4405
rect 1746 4401 1752 4405
rect 1756 4401 1762 4405
rect 1717 4400 1762 4401
rect 1721 4396 1727 4400
rect 1731 4396 1737 4400
rect 1741 4396 1747 4400
rect 1751 4396 1757 4400
rect 1761 4396 1762 4400
rect 1717 4395 1762 4396
rect 1717 4391 1722 4395
rect 1726 4391 1732 4395
rect 1736 4391 1742 4395
rect 1746 4391 1752 4395
rect 1756 4391 1762 4395
rect 1717 4390 1762 4391
rect 1721 4386 1727 4390
rect 1731 4386 1737 4390
rect 1741 4386 1747 4390
rect 1751 4386 1757 4390
rect 1761 4386 1762 4390
rect 1717 4385 1762 4386
rect 1717 4381 1722 4385
rect 1726 4381 1732 4385
rect 1736 4381 1742 4385
rect 1746 4381 1752 4385
rect 1756 4381 1762 4385
rect 1717 4380 1762 4381
rect 1721 4376 1727 4380
rect 1731 4376 1737 4380
rect 1741 4376 1747 4380
rect 1751 4376 1757 4380
rect 1761 4376 1762 4380
rect 1717 4375 1762 4376
rect 1717 4371 1722 4375
rect 1726 4371 1732 4375
rect 1736 4371 1742 4375
rect 1746 4371 1752 4375
rect 1756 4371 1762 4375
rect 1717 4370 1762 4371
rect 1721 4366 1727 4370
rect 1731 4366 1737 4370
rect 1741 4366 1747 4370
rect 1751 4366 1757 4370
rect 1761 4366 1762 4370
rect 1717 4365 1762 4366
rect 1717 4361 1722 4365
rect 1726 4361 1732 4365
rect 1736 4361 1742 4365
rect 1746 4361 1752 4365
rect 1756 4361 1762 4365
rect 2030 4446 2036 4450
rect 2040 4446 2046 4450
rect 2050 4446 2056 4450
rect 2060 4446 2066 4450
rect 2070 4446 2071 4450
rect 2026 4445 2071 4446
rect 2026 4441 2031 4445
rect 2035 4441 2041 4445
rect 2045 4441 2051 4445
rect 2055 4441 2061 4445
rect 2065 4441 2071 4445
rect 2026 4440 2071 4441
rect 2030 4436 2036 4440
rect 2040 4436 2046 4440
rect 2050 4436 2056 4440
rect 2060 4436 2066 4440
rect 2070 4436 2071 4440
rect 2026 4435 2071 4436
rect 2026 4431 2031 4435
rect 2035 4431 2041 4435
rect 2045 4431 2051 4435
rect 2055 4431 2061 4435
rect 2065 4431 2071 4435
rect 2026 4430 2071 4431
rect 2030 4426 2036 4430
rect 2040 4426 2046 4430
rect 2050 4426 2056 4430
rect 2060 4426 2066 4430
rect 2070 4426 2071 4430
rect 2026 4425 2071 4426
rect 2026 4421 2031 4425
rect 2035 4421 2041 4425
rect 2045 4421 2051 4425
rect 2055 4421 2061 4425
rect 2065 4421 2071 4425
rect 2026 4420 2071 4421
rect 2030 4416 2036 4420
rect 2040 4416 2046 4420
rect 2050 4416 2056 4420
rect 2060 4416 2066 4420
rect 2070 4416 2071 4420
rect 2026 4415 2071 4416
rect 2026 4411 2031 4415
rect 2035 4411 2041 4415
rect 2045 4411 2051 4415
rect 2055 4411 2061 4415
rect 2065 4411 2071 4415
rect 2026 4410 2071 4411
rect 2030 4406 2036 4410
rect 2040 4406 2046 4410
rect 2050 4406 2056 4410
rect 2060 4406 2066 4410
rect 2070 4406 2071 4410
rect 2026 4405 2071 4406
rect 2026 4401 2031 4405
rect 2035 4401 2041 4405
rect 2045 4401 2051 4405
rect 2055 4401 2061 4405
rect 2065 4401 2071 4405
rect 2026 4400 2071 4401
rect 2030 4396 2036 4400
rect 2040 4396 2046 4400
rect 2050 4396 2056 4400
rect 2060 4396 2066 4400
rect 2070 4396 2071 4400
rect 2026 4395 2071 4396
rect 2026 4391 2031 4395
rect 2035 4391 2041 4395
rect 2045 4391 2051 4395
rect 2055 4391 2061 4395
rect 2065 4391 2071 4395
rect 2026 4390 2071 4391
rect 2030 4386 2036 4390
rect 2040 4386 2046 4390
rect 2050 4386 2056 4390
rect 2060 4386 2066 4390
rect 2070 4386 2071 4390
rect 2026 4385 2071 4386
rect 2026 4381 2031 4385
rect 2035 4381 2041 4385
rect 2045 4381 2051 4385
rect 2055 4381 2061 4385
rect 2065 4381 2071 4385
rect 2026 4380 2071 4381
rect 2030 4376 2036 4380
rect 2040 4376 2046 4380
rect 2050 4376 2056 4380
rect 2060 4376 2066 4380
rect 2070 4376 2071 4380
rect 2026 4375 2071 4376
rect 2026 4371 2031 4375
rect 2035 4371 2041 4375
rect 2045 4371 2051 4375
rect 2055 4371 2061 4375
rect 2065 4371 2071 4375
rect 2026 4370 2071 4371
rect 2030 4366 2036 4370
rect 2040 4366 2046 4370
rect 2050 4366 2056 4370
rect 2060 4366 2066 4370
rect 2070 4366 2071 4370
rect 2026 4365 2071 4366
rect 2026 4361 2031 4365
rect 2035 4361 2041 4365
rect 2045 4361 2051 4365
rect 2055 4361 2061 4365
rect 2065 4361 2071 4365
rect 2339 4446 2345 4450
rect 2349 4446 2355 4450
rect 2359 4446 2365 4450
rect 2369 4446 2375 4450
rect 2379 4446 2380 4450
rect 2335 4445 2380 4446
rect 2335 4441 2340 4445
rect 2344 4441 2350 4445
rect 2354 4441 2360 4445
rect 2364 4441 2370 4445
rect 2374 4441 2380 4445
rect 2335 4440 2380 4441
rect 2339 4436 2345 4440
rect 2349 4436 2355 4440
rect 2359 4436 2365 4440
rect 2369 4436 2375 4440
rect 2379 4436 2380 4440
rect 2335 4435 2380 4436
rect 2335 4431 2340 4435
rect 2344 4431 2350 4435
rect 2354 4431 2360 4435
rect 2364 4431 2370 4435
rect 2374 4431 2380 4435
rect 2335 4430 2380 4431
rect 2339 4426 2345 4430
rect 2349 4426 2355 4430
rect 2359 4426 2365 4430
rect 2369 4426 2375 4430
rect 2379 4426 2380 4430
rect 2335 4425 2380 4426
rect 2335 4421 2340 4425
rect 2344 4421 2350 4425
rect 2354 4421 2360 4425
rect 2364 4421 2370 4425
rect 2374 4421 2380 4425
rect 2335 4420 2380 4421
rect 2339 4416 2345 4420
rect 2349 4416 2355 4420
rect 2359 4416 2365 4420
rect 2369 4416 2375 4420
rect 2379 4416 2380 4420
rect 2335 4415 2380 4416
rect 2335 4411 2340 4415
rect 2344 4411 2350 4415
rect 2354 4411 2360 4415
rect 2364 4411 2370 4415
rect 2374 4411 2380 4415
rect 2335 4410 2380 4411
rect 2339 4406 2345 4410
rect 2349 4406 2355 4410
rect 2359 4406 2365 4410
rect 2369 4406 2375 4410
rect 2379 4406 2380 4410
rect 2335 4405 2380 4406
rect 2335 4401 2340 4405
rect 2344 4401 2350 4405
rect 2354 4401 2360 4405
rect 2364 4401 2370 4405
rect 2374 4401 2380 4405
rect 2335 4400 2380 4401
rect 2339 4396 2345 4400
rect 2349 4396 2355 4400
rect 2359 4396 2365 4400
rect 2369 4396 2375 4400
rect 2379 4396 2380 4400
rect 2335 4395 2380 4396
rect 2335 4391 2340 4395
rect 2344 4391 2350 4395
rect 2354 4391 2360 4395
rect 2364 4391 2370 4395
rect 2374 4391 2380 4395
rect 2335 4390 2380 4391
rect 2339 4386 2345 4390
rect 2349 4386 2355 4390
rect 2359 4386 2365 4390
rect 2369 4386 2375 4390
rect 2379 4386 2380 4390
rect 2335 4385 2380 4386
rect 2335 4381 2340 4385
rect 2344 4381 2350 4385
rect 2354 4381 2360 4385
rect 2364 4381 2370 4385
rect 2374 4381 2380 4385
rect 2335 4380 2380 4381
rect 2339 4376 2345 4380
rect 2349 4376 2355 4380
rect 2359 4376 2365 4380
rect 2369 4376 2375 4380
rect 2379 4376 2380 4380
rect 2335 4375 2380 4376
rect 2335 4371 2340 4375
rect 2344 4371 2350 4375
rect 2354 4371 2360 4375
rect 2364 4371 2370 4375
rect 2374 4371 2380 4375
rect 2335 4370 2380 4371
rect 2339 4366 2345 4370
rect 2349 4366 2355 4370
rect 2359 4366 2365 4370
rect 2369 4366 2375 4370
rect 2379 4366 2380 4370
rect 2335 4365 2380 4366
rect 2335 4361 2340 4365
rect 2344 4361 2350 4365
rect 2354 4361 2360 4365
rect 2364 4361 2370 4365
rect 2374 4361 2380 4365
rect 2648 4446 2654 4450
rect 2658 4446 2664 4450
rect 2668 4446 2674 4450
rect 2678 4446 2684 4450
rect 2688 4446 2689 4450
rect 2644 4445 2689 4446
rect 2644 4441 2649 4445
rect 2653 4441 2659 4445
rect 2663 4441 2669 4445
rect 2673 4441 2679 4445
rect 2683 4441 2689 4445
rect 2644 4440 2689 4441
rect 2648 4436 2654 4440
rect 2658 4436 2664 4440
rect 2668 4436 2674 4440
rect 2678 4436 2684 4440
rect 2688 4436 2689 4440
rect 2644 4435 2689 4436
rect 2644 4431 2649 4435
rect 2653 4431 2659 4435
rect 2663 4431 2669 4435
rect 2673 4431 2679 4435
rect 2683 4431 2689 4435
rect 2644 4430 2689 4431
rect 2648 4426 2654 4430
rect 2658 4426 2664 4430
rect 2668 4426 2674 4430
rect 2678 4426 2684 4430
rect 2688 4426 2689 4430
rect 2644 4425 2689 4426
rect 2644 4421 2649 4425
rect 2653 4421 2659 4425
rect 2663 4421 2669 4425
rect 2673 4421 2679 4425
rect 2683 4421 2689 4425
rect 2644 4420 2689 4421
rect 2648 4416 2654 4420
rect 2658 4416 2664 4420
rect 2668 4416 2674 4420
rect 2678 4416 2684 4420
rect 2688 4416 2689 4420
rect 2644 4415 2689 4416
rect 2644 4411 2649 4415
rect 2653 4411 2659 4415
rect 2663 4411 2669 4415
rect 2673 4411 2679 4415
rect 2683 4411 2689 4415
rect 2644 4410 2689 4411
rect 2648 4406 2654 4410
rect 2658 4406 2664 4410
rect 2668 4406 2674 4410
rect 2678 4406 2684 4410
rect 2688 4406 2689 4410
rect 2644 4405 2689 4406
rect 2644 4401 2649 4405
rect 2653 4401 2659 4405
rect 2663 4401 2669 4405
rect 2673 4401 2679 4405
rect 2683 4401 2689 4405
rect 2644 4400 2689 4401
rect 2648 4396 2654 4400
rect 2658 4396 2664 4400
rect 2668 4396 2674 4400
rect 2678 4396 2684 4400
rect 2688 4396 2689 4400
rect 2644 4395 2689 4396
rect 2644 4391 2649 4395
rect 2653 4391 2659 4395
rect 2663 4391 2669 4395
rect 2673 4391 2679 4395
rect 2683 4391 2689 4395
rect 2644 4390 2689 4391
rect 2648 4386 2654 4390
rect 2658 4386 2664 4390
rect 2668 4386 2674 4390
rect 2678 4386 2684 4390
rect 2688 4386 2689 4390
rect 2644 4385 2689 4386
rect 2644 4381 2649 4385
rect 2653 4381 2659 4385
rect 2663 4381 2669 4385
rect 2673 4381 2679 4385
rect 2683 4381 2689 4385
rect 2644 4380 2689 4381
rect 2648 4376 2654 4380
rect 2658 4376 2664 4380
rect 2668 4376 2674 4380
rect 2678 4376 2684 4380
rect 2688 4376 2689 4380
rect 2644 4375 2689 4376
rect 2644 4371 2649 4375
rect 2653 4371 2659 4375
rect 2663 4371 2669 4375
rect 2673 4371 2679 4375
rect 2683 4371 2689 4375
rect 2644 4370 2689 4371
rect 2648 4366 2654 4370
rect 2658 4366 2664 4370
rect 2668 4366 2674 4370
rect 2678 4366 2684 4370
rect 2688 4366 2689 4370
rect 2644 4365 2689 4366
rect 2644 4361 2649 4365
rect 2653 4361 2659 4365
rect 2663 4361 2669 4365
rect 2673 4361 2679 4365
rect 2683 4361 2689 4365
rect 2957 4446 2963 4450
rect 2967 4446 2973 4450
rect 2977 4446 2983 4450
rect 2987 4446 2993 4450
rect 2997 4446 2998 4450
rect 2953 4445 2998 4446
rect 2953 4441 2958 4445
rect 2962 4441 2968 4445
rect 2972 4441 2978 4445
rect 2982 4441 2988 4445
rect 2992 4441 2998 4445
rect 2953 4440 2998 4441
rect 2957 4436 2963 4440
rect 2967 4436 2973 4440
rect 2977 4436 2983 4440
rect 2987 4436 2993 4440
rect 2997 4436 2998 4440
rect 2953 4435 2998 4436
rect 2953 4431 2958 4435
rect 2962 4431 2968 4435
rect 2972 4431 2978 4435
rect 2982 4431 2988 4435
rect 2992 4431 2998 4435
rect 2953 4430 2998 4431
rect 2957 4426 2963 4430
rect 2967 4426 2973 4430
rect 2977 4426 2983 4430
rect 2987 4426 2993 4430
rect 2997 4426 2998 4430
rect 2953 4425 2998 4426
rect 2953 4421 2958 4425
rect 2962 4421 2968 4425
rect 2972 4421 2978 4425
rect 2982 4421 2988 4425
rect 2992 4421 2998 4425
rect 2953 4420 2998 4421
rect 2957 4416 2963 4420
rect 2967 4416 2973 4420
rect 2977 4416 2983 4420
rect 2987 4416 2993 4420
rect 2997 4416 2998 4420
rect 2953 4415 2998 4416
rect 2953 4411 2958 4415
rect 2962 4411 2968 4415
rect 2972 4411 2978 4415
rect 2982 4411 2988 4415
rect 2992 4411 2998 4415
rect 2953 4410 2998 4411
rect 2957 4406 2963 4410
rect 2967 4406 2973 4410
rect 2977 4406 2983 4410
rect 2987 4406 2993 4410
rect 2997 4406 2998 4410
rect 2953 4405 2998 4406
rect 2953 4401 2958 4405
rect 2962 4401 2968 4405
rect 2972 4401 2978 4405
rect 2982 4401 2988 4405
rect 2992 4401 2998 4405
rect 2953 4400 2998 4401
rect 2957 4396 2963 4400
rect 2967 4396 2973 4400
rect 2977 4396 2983 4400
rect 2987 4396 2993 4400
rect 2997 4396 2998 4400
rect 2953 4395 2998 4396
rect 2953 4391 2958 4395
rect 2962 4391 2968 4395
rect 2972 4391 2978 4395
rect 2982 4391 2988 4395
rect 2992 4391 2998 4395
rect 2953 4390 2998 4391
rect 2957 4386 2963 4390
rect 2967 4386 2973 4390
rect 2977 4386 2983 4390
rect 2987 4386 2993 4390
rect 2997 4386 2998 4390
rect 2953 4385 2998 4386
rect 2953 4381 2958 4385
rect 2962 4381 2968 4385
rect 2972 4381 2978 4385
rect 2982 4381 2988 4385
rect 2992 4381 2998 4385
rect 2953 4380 2998 4381
rect 2957 4376 2963 4380
rect 2967 4376 2973 4380
rect 2977 4376 2983 4380
rect 2987 4376 2993 4380
rect 2997 4376 2998 4380
rect 2953 4375 2998 4376
rect 2953 4371 2958 4375
rect 2962 4371 2968 4375
rect 2972 4371 2978 4375
rect 2982 4371 2988 4375
rect 2992 4371 2998 4375
rect 2953 4370 2998 4371
rect 2957 4366 2963 4370
rect 2967 4366 2973 4370
rect 2977 4366 2983 4370
rect 2987 4366 2993 4370
rect 2997 4366 2998 4370
rect 2953 4365 2998 4366
rect 2953 4361 2958 4365
rect 2962 4361 2968 4365
rect 2972 4361 2978 4365
rect 2982 4361 2988 4365
rect 2992 4361 2998 4365
rect 3266 4446 3272 4450
rect 3276 4446 3282 4450
rect 3286 4446 3292 4450
rect 3296 4446 3302 4450
rect 3306 4446 3307 4450
rect 3262 4445 3307 4446
rect 3262 4441 3267 4445
rect 3271 4441 3277 4445
rect 3281 4441 3287 4445
rect 3291 4441 3297 4445
rect 3301 4441 3307 4445
rect 3262 4440 3307 4441
rect 3266 4436 3272 4440
rect 3276 4436 3282 4440
rect 3286 4436 3292 4440
rect 3296 4436 3302 4440
rect 3306 4436 3307 4440
rect 3262 4435 3307 4436
rect 3262 4431 3267 4435
rect 3271 4431 3277 4435
rect 3281 4431 3287 4435
rect 3291 4431 3297 4435
rect 3301 4431 3307 4435
rect 3262 4430 3307 4431
rect 3266 4426 3272 4430
rect 3276 4426 3282 4430
rect 3286 4426 3292 4430
rect 3296 4426 3302 4430
rect 3306 4426 3307 4430
rect 3262 4425 3307 4426
rect 3262 4421 3267 4425
rect 3271 4421 3277 4425
rect 3281 4421 3287 4425
rect 3291 4421 3297 4425
rect 3301 4421 3307 4425
rect 3262 4420 3307 4421
rect 3266 4416 3272 4420
rect 3276 4416 3282 4420
rect 3286 4416 3292 4420
rect 3296 4416 3302 4420
rect 3306 4416 3307 4420
rect 3262 4415 3307 4416
rect 3262 4411 3267 4415
rect 3271 4411 3277 4415
rect 3281 4411 3287 4415
rect 3291 4411 3297 4415
rect 3301 4411 3307 4415
rect 3262 4410 3307 4411
rect 3266 4406 3272 4410
rect 3276 4406 3282 4410
rect 3286 4406 3292 4410
rect 3296 4406 3302 4410
rect 3306 4406 3307 4410
rect 3262 4405 3307 4406
rect 3262 4401 3267 4405
rect 3271 4401 3277 4405
rect 3281 4401 3287 4405
rect 3291 4401 3297 4405
rect 3301 4401 3307 4405
rect 3262 4400 3307 4401
rect 3266 4396 3272 4400
rect 3276 4396 3282 4400
rect 3286 4396 3292 4400
rect 3296 4396 3302 4400
rect 3306 4396 3307 4400
rect 3262 4395 3307 4396
rect 3262 4391 3267 4395
rect 3271 4391 3277 4395
rect 3281 4391 3287 4395
rect 3291 4391 3297 4395
rect 3301 4391 3307 4395
rect 3262 4390 3307 4391
rect 3266 4386 3272 4390
rect 3276 4386 3282 4390
rect 3286 4386 3292 4390
rect 3296 4386 3302 4390
rect 3306 4386 3307 4390
rect 3262 4385 3307 4386
rect 3262 4381 3267 4385
rect 3271 4381 3277 4385
rect 3281 4381 3287 4385
rect 3291 4381 3297 4385
rect 3301 4381 3307 4385
rect 3262 4380 3307 4381
rect 3266 4376 3272 4380
rect 3276 4376 3282 4380
rect 3286 4376 3292 4380
rect 3296 4376 3302 4380
rect 3306 4376 3307 4380
rect 3262 4375 3307 4376
rect 3262 4371 3267 4375
rect 3271 4371 3277 4375
rect 3281 4371 3287 4375
rect 3291 4371 3297 4375
rect 3301 4371 3307 4375
rect 3262 4370 3307 4371
rect 3266 4366 3272 4370
rect 3276 4366 3282 4370
rect 3286 4366 3292 4370
rect 3296 4366 3302 4370
rect 3306 4366 3307 4370
rect 3262 4365 3307 4366
rect 3262 4361 3267 4365
rect 3271 4361 3277 4365
rect 3281 4361 3287 4365
rect 3291 4361 3297 4365
rect 3301 4361 3307 4365
rect 3575 4446 3581 4450
rect 3585 4446 3591 4450
rect 3595 4446 3601 4450
rect 3605 4446 3611 4450
rect 3615 4446 3616 4450
rect 3571 4445 3616 4446
rect 3571 4441 3576 4445
rect 3580 4441 3586 4445
rect 3590 4441 3596 4445
rect 3600 4441 3606 4445
rect 3610 4441 3616 4445
rect 3571 4440 3616 4441
rect 3575 4436 3581 4440
rect 3585 4436 3591 4440
rect 3595 4436 3601 4440
rect 3605 4436 3611 4440
rect 3615 4436 3616 4440
rect 3571 4435 3616 4436
rect 3571 4431 3576 4435
rect 3580 4431 3586 4435
rect 3590 4431 3596 4435
rect 3600 4431 3606 4435
rect 3610 4431 3616 4435
rect 3571 4430 3616 4431
rect 3575 4426 3581 4430
rect 3585 4426 3591 4430
rect 3595 4426 3601 4430
rect 3605 4426 3611 4430
rect 3615 4426 3616 4430
rect 3571 4425 3616 4426
rect 3571 4421 3576 4425
rect 3580 4421 3586 4425
rect 3590 4421 3596 4425
rect 3600 4421 3606 4425
rect 3610 4421 3616 4425
rect 3571 4420 3616 4421
rect 3575 4416 3581 4420
rect 3585 4416 3591 4420
rect 3595 4416 3601 4420
rect 3605 4416 3611 4420
rect 3615 4416 3616 4420
rect 3571 4415 3616 4416
rect 3571 4411 3576 4415
rect 3580 4411 3586 4415
rect 3590 4411 3596 4415
rect 3600 4411 3606 4415
rect 3610 4411 3616 4415
rect 3571 4410 3616 4411
rect 3575 4406 3581 4410
rect 3585 4406 3591 4410
rect 3595 4406 3601 4410
rect 3605 4406 3611 4410
rect 3615 4406 3616 4410
rect 3571 4405 3616 4406
rect 3571 4401 3576 4405
rect 3580 4401 3586 4405
rect 3590 4401 3596 4405
rect 3600 4401 3606 4405
rect 3610 4401 3616 4405
rect 3571 4400 3616 4401
rect 3575 4396 3581 4400
rect 3585 4396 3591 4400
rect 3595 4396 3601 4400
rect 3605 4396 3611 4400
rect 3615 4396 3616 4400
rect 3571 4395 3616 4396
rect 3571 4391 3576 4395
rect 3580 4391 3586 4395
rect 3590 4391 3596 4395
rect 3600 4391 3606 4395
rect 3610 4391 3616 4395
rect 3571 4390 3616 4391
rect 3575 4386 3581 4390
rect 3585 4386 3591 4390
rect 3595 4386 3601 4390
rect 3605 4386 3611 4390
rect 3615 4386 3616 4390
rect 3571 4385 3616 4386
rect 3571 4381 3576 4385
rect 3580 4381 3586 4385
rect 3590 4381 3596 4385
rect 3600 4381 3606 4385
rect 3610 4381 3616 4385
rect 3571 4380 3616 4381
rect 3575 4376 3581 4380
rect 3585 4376 3591 4380
rect 3595 4376 3601 4380
rect 3605 4376 3611 4380
rect 3615 4376 3616 4380
rect 3571 4375 3616 4376
rect 3571 4371 3576 4375
rect 3580 4371 3586 4375
rect 3590 4371 3596 4375
rect 3600 4371 3606 4375
rect 3610 4371 3616 4375
rect 3571 4370 3616 4371
rect 3575 4366 3581 4370
rect 3585 4366 3591 4370
rect 3595 4366 3601 4370
rect 3605 4366 3611 4370
rect 3615 4366 3616 4370
rect 3571 4365 3616 4366
rect 3571 4361 3576 4365
rect 3580 4361 3586 4365
rect 3590 4361 3596 4365
rect 3600 4361 3606 4365
rect 3610 4361 3616 4365
<< ndcontact >>
rect 1402 9949 1406 9953
rect 1412 9949 1416 9953
rect 1422 9949 1426 9953
rect 1432 9949 1436 9953
rect 1397 9944 1401 9948
rect 1407 9944 1411 9948
rect 1417 9944 1421 9948
rect 1427 9944 1431 9948
rect 1437 9944 1441 9948
rect 1402 9939 1406 9943
rect 1412 9939 1416 9943
rect 1422 9939 1426 9943
rect 1432 9939 1436 9943
rect 1397 9934 1401 9938
rect 1407 9934 1411 9938
rect 1417 9934 1421 9938
rect 1427 9934 1431 9938
rect 1437 9934 1441 9938
rect 1402 9929 1406 9933
rect 1412 9929 1416 9933
rect 1422 9929 1426 9933
rect 1432 9929 1436 9933
rect 1397 9924 1401 9928
rect 1407 9924 1411 9928
rect 1417 9924 1421 9928
rect 1427 9924 1431 9928
rect 1437 9924 1441 9928
rect 1402 9919 1406 9923
rect 1412 9919 1416 9923
rect 1422 9919 1426 9923
rect 1432 9919 1436 9923
rect 1397 9914 1401 9918
rect 1407 9914 1411 9918
rect 1417 9914 1421 9918
rect 1427 9914 1431 9918
rect 1437 9914 1441 9918
rect 1402 9909 1406 9913
rect 1412 9909 1416 9913
rect 1422 9909 1426 9913
rect 1432 9909 1436 9913
rect 1397 9904 1401 9908
rect 1407 9904 1411 9908
rect 1417 9904 1421 9908
rect 1427 9904 1431 9908
rect 1437 9904 1441 9908
rect 1402 9899 1406 9903
rect 1412 9899 1416 9903
rect 1422 9899 1426 9903
rect 1432 9899 1436 9903
rect 1397 9894 1401 9898
rect 1407 9894 1411 9898
rect 1417 9894 1421 9898
rect 1427 9894 1431 9898
rect 1437 9894 1441 9898
rect 1402 9889 1406 9893
rect 1412 9889 1416 9893
rect 1422 9889 1426 9893
rect 1432 9889 1436 9893
rect 1397 9884 1401 9888
rect 1407 9884 1411 9888
rect 1417 9884 1421 9888
rect 1427 9884 1431 9888
rect 1437 9884 1441 9888
rect 1402 9879 1406 9883
rect 1412 9879 1416 9883
rect 1422 9879 1426 9883
rect 1432 9879 1436 9883
rect 1397 9874 1401 9878
rect 1407 9874 1411 9878
rect 1417 9874 1421 9878
rect 1427 9874 1431 9878
rect 1437 9874 1441 9878
rect 1402 9869 1406 9873
rect 1412 9869 1416 9873
rect 1422 9869 1426 9873
rect 1432 9869 1436 9873
rect 1397 9864 1401 9868
rect 1407 9864 1411 9868
rect 1417 9864 1421 9868
rect 1427 9864 1431 9868
rect 1437 9864 1441 9868
rect 1711 9949 1715 9953
rect 1721 9949 1725 9953
rect 1731 9949 1735 9953
rect 1741 9949 1745 9953
rect 1706 9944 1710 9948
rect 1716 9944 1720 9948
rect 1726 9944 1730 9948
rect 1736 9944 1740 9948
rect 1746 9944 1750 9948
rect 1711 9939 1715 9943
rect 1721 9939 1725 9943
rect 1731 9939 1735 9943
rect 1741 9939 1745 9943
rect 1706 9934 1710 9938
rect 1716 9934 1720 9938
rect 1726 9934 1730 9938
rect 1736 9934 1740 9938
rect 1746 9934 1750 9938
rect 1711 9929 1715 9933
rect 1721 9929 1725 9933
rect 1731 9929 1735 9933
rect 1741 9929 1745 9933
rect 1706 9924 1710 9928
rect 1716 9924 1720 9928
rect 1726 9924 1730 9928
rect 1736 9924 1740 9928
rect 1746 9924 1750 9928
rect 1711 9919 1715 9923
rect 1721 9919 1725 9923
rect 1731 9919 1735 9923
rect 1741 9919 1745 9923
rect 1706 9914 1710 9918
rect 1716 9914 1720 9918
rect 1726 9914 1730 9918
rect 1736 9914 1740 9918
rect 1746 9914 1750 9918
rect 1711 9909 1715 9913
rect 1721 9909 1725 9913
rect 1731 9909 1735 9913
rect 1741 9909 1745 9913
rect 1706 9904 1710 9908
rect 1716 9904 1720 9908
rect 1726 9904 1730 9908
rect 1736 9904 1740 9908
rect 1746 9904 1750 9908
rect 1711 9899 1715 9903
rect 1721 9899 1725 9903
rect 1731 9899 1735 9903
rect 1741 9899 1745 9903
rect 1706 9894 1710 9898
rect 1716 9894 1720 9898
rect 1726 9894 1730 9898
rect 1736 9894 1740 9898
rect 1746 9894 1750 9898
rect 1711 9889 1715 9893
rect 1721 9889 1725 9893
rect 1731 9889 1735 9893
rect 1741 9889 1745 9893
rect 1706 9884 1710 9888
rect 1716 9884 1720 9888
rect 1726 9884 1730 9888
rect 1736 9884 1740 9888
rect 1746 9884 1750 9888
rect 1711 9879 1715 9883
rect 1721 9879 1725 9883
rect 1731 9879 1735 9883
rect 1741 9879 1745 9883
rect 1706 9874 1710 9878
rect 1716 9874 1720 9878
rect 1726 9874 1730 9878
rect 1736 9874 1740 9878
rect 1746 9874 1750 9878
rect 1711 9869 1715 9873
rect 1721 9869 1725 9873
rect 1731 9869 1735 9873
rect 1741 9869 1745 9873
rect 1706 9864 1710 9868
rect 1716 9864 1720 9868
rect 1726 9864 1730 9868
rect 1736 9864 1740 9868
rect 1746 9864 1750 9868
rect 2020 9949 2024 9953
rect 2030 9949 2034 9953
rect 2040 9949 2044 9953
rect 2050 9949 2054 9953
rect 2015 9944 2019 9948
rect 2025 9944 2029 9948
rect 2035 9944 2039 9948
rect 2045 9944 2049 9948
rect 2055 9944 2059 9948
rect 2020 9939 2024 9943
rect 2030 9939 2034 9943
rect 2040 9939 2044 9943
rect 2050 9939 2054 9943
rect 2015 9934 2019 9938
rect 2025 9934 2029 9938
rect 2035 9934 2039 9938
rect 2045 9934 2049 9938
rect 2055 9934 2059 9938
rect 2020 9929 2024 9933
rect 2030 9929 2034 9933
rect 2040 9929 2044 9933
rect 2050 9929 2054 9933
rect 2015 9924 2019 9928
rect 2025 9924 2029 9928
rect 2035 9924 2039 9928
rect 2045 9924 2049 9928
rect 2055 9924 2059 9928
rect 2020 9919 2024 9923
rect 2030 9919 2034 9923
rect 2040 9919 2044 9923
rect 2050 9919 2054 9923
rect 2015 9914 2019 9918
rect 2025 9914 2029 9918
rect 2035 9914 2039 9918
rect 2045 9914 2049 9918
rect 2055 9914 2059 9918
rect 2020 9909 2024 9913
rect 2030 9909 2034 9913
rect 2040 9909 2044 9913
rect 2050 9909 2054 9913
rect 2015 9904 2019 9908
rect 2025 9904 2029 9908
rect 2035 9904 2039 9908
rect 2045 9904 2049 9908
rect 2055 9904 2059 9908
rect 2020 9899 2024 9903
rect 2030 9899 2034 9903
rect 2040 9899 2044 9903
rect 2050 9899 2054 9903
rect 2015 9894 2019 9898
rect 2025 9894 2029 9898
rect 2035 9894 2039 9898
rect 2045 9894 2049 9898
rect 2055 9894 2059 9898
rect 2020 9889 2024 9893
rect 2030 9889 2034 9893
rect 2040 9889 2044 9893
rect 2050 9889 2054 9893
rect 2015 9884 2019 9888
rect 2025 9884 2029 9888
rect 2035 9884 2039 9888
rect 2045 9884 2049 9888
rect 2055 9884 2059 9888
rect 2020 9879 2024 9883
rect 2030 9879 2034 9883
rect 2040 9879 2044 9883
rect 2050 9879 2054 9883
rect 2015 9874 2019 9878
rect 2025 9874 2029 9878
rect 2035 9874 2039 9878
rect 2045 9874 2049 9878
rect 2055 9874 2059 9878
rect 2020 9869 2024 9873
rect 2030 9869 2034 9873
rect 2040 9869 2044 9873
rect 2050 9869 2054 9873
rect 2015 9864 2019 9868
rect 2025 9864 2029 9868
rect 2035 9864 2039 9868
rect 2045 9864 2049 9868
rect 2055 9864 2059 9868
rect 2329 9949 2333 9953
rect 2339 9949 2343 9953
rect 2349 9949 2353 9953
rect 2359 9949 2363 9953
rect 2324 9944 2328 9948
rect 2334 9944 2338 9948
rect 2344 9944 2348 9948
rect 2354 9944 2358 9948
rect 2364 9944 2368 9948
rect 2329 9939 2333 9943
rect 2339 9939 2343 9943
rect 2349 9939 2353 9943
rect 2359 9939 2363 9943
rect 2324 9934 2328 9938
rect 2334 9934 2338 9938
rect 2344 9934 2348 9938
rect 2354 9934 2358 9938
rect 2364 9934 2368 9938
rect 2329 9929 2333 9933
rect 2339 9929 2343 9933
rect 2349 9929 2353 9933
rect 2359 9929 2363 9933
rect 2324 9924 2328 9928
rect 2334 9924 2338 9928
rect 2344 9924 2348 9928
rect 2354 9924 2358 9928
rect 2364 9924 2368 9928
rect 2329 9919 2333 9923
rect 2339 9919 2343 9923
rect 2349 9919 2353 9923
rect 2359 9919 2363 9923
rect 2324 9914 2328 9918
rect 2334 9914 2338 9918
rect 2344 9914 2348 9918
rect 2354 9914 2358 9918
rect 2364 9914 2368 9918
rect 2329 9909 2333 9913
rect 2339 9909 2343 9913
rect 2349 9909 2353 9913
rect 2359 9909 2363 9913
rect 2324 9904 2328 9908
rect 2334 9904 2338 9908
rect 2344 9904 2348 9908
rect 2354 9904 2358 9908
rect 2364 9904 2368 9908
rect 2329 9899 2333 9903
rect 2339 9899 2343 9903
rect 2349 9899 2353 9903
rect 2359 9899 2363 9903
rect 2324 9894 2328 9898
rect 2334 9894 2338 9898
rect 2344 9894 2348 9898
rect 2354 9894 2358 9898
rect 2364 9894 2368 9898
rect 2329 9889 2333 9893
rect 2339 9889 2343 9893
rect 2349 9889 2353 9893
rect 2359 9889 2363 9893
rect 2324 9884 2328 9888
rect 2334 9884 2338 9888
rect 2344 9884 2348 9888
rect 2354 9884 2358 9888
rect 2364 9884 2368 9888
rect 2329 9879 2333 9883
rect 2339 9879 2343 9883
rect 2349 9879 2353 9883
rect 2359 9879 2363 9883
rect 2324 9874 2328 9878
rect 2334 9874 2338 9878
rect 2344 9874 2348 9878
rect 2354 9874 2358 9878
rect 2364 9874 2368 9878
rect 2329 9869 2333 9873
rect 2339 9869 2343 9873
rect 2349 9869 2353 9873
rect 2359 9869 2363 9873
rect 2324 9864 2328 9868
rect 2334 9864 2338 9868
rect 2344 9864 2348 9868
rect 2354 9864 2358 9868
rect 2364 9864 2368 9868
rect 2638 9949 2642 9953
rect 2648 9949 2652 9953
rect 2658 9949 2662 9953
rect 2668 9949 2672 9953
rect 2633 9944 2637 9948
rect 2643 9944 2647 9948
rect 2653 9944 2657 9948
rect 2663 9944 2667 9948
rect 2673 9944 2677 9948
rect 2638 9939 2642 9943
rect 2648 9939 2652 9943
rect 2658 9939 2662 9943
rect 2668 9939 2672 9943
rect 2633 9934 2637 9938
rect 2643 9934 2647 9938
rect 2653 9934 2657 9938
rect 2663 9934 2667 9938
rect 2673 9934 2677 9938
rect 2638 9929 2642 9933
rect 2648 9929 2652 9933
rect 2658 9929 2662 9933
rect 2668 9929 2672 9933
rect 2633 9924 2637 9928
rect 2643 9924 2647 9928
rect 2653 9924 2657 9928
rect 2663 9924 2667 9928
rect 2673 9924 2677 9928
rect 2638 9919 2642 9923
rect 2648 9919 2652 9923
rect 2658 9919 2662 9923
rect 2668 9919 2672 9923
rect 2633 9914 2637 9918
rect 2643 9914 2647 9918
rect 2653 9914 2657 9918
rect 2663 9914 2667 9918
rect 2673 9914 2677 9918
rect 2638 9909 2642 9913
rect 2648 9909 2652 9913
rect 2658 9909 2662 9913
rect 2668 9909 2672 9913
rect 2633 9904 2637 9908
rect 2643 9904 2647 9908
rect 2653 9904 2657 9908
rect 2663 9904 2667 9908
rect 2673 9904 2677 9908
rect 2638 9899 2642 9903
rect 2648 9899 2652 9903
rect 2658 9899 2662 9903
rect 2668 9899 2672 9903
rect 2633 9894 2637 9898
rect 2643 9894 2647 9898
rect 2653 9894 2657 9898
rect 2663 9894 2667 9898
rect 2673 9894 2677 9898
rect 2638 9889 2642 9893
rect 2648 9889 2652 9893
rect 2658 9889 2662 9893
rect 2668 9889 2672 9893
rect 2633 9884 2637 9888
rect 2643 9884 2647 9888
rect 2653 9884 2657 9888
rect 2663 9884 2667 9888
rect 2673 9884 2677 9888
rect 2638 9879 2642 9883
rect 2648 9879 2652 9883
rect 2658 9879 2662 9883
rect 2668 9879 2672 9883
rect 2633 9874 2637 9878
rect 2643 9874 2647 9878
rect 2653 9874 2657 9878
rect 2663 9874 2667 9878
rect 2673 9874 2677 9878
rect 2638 9869 2642 9873
rect 2648 9869 2652 9873
rect 2658 9869 2662 9873
rect 2668 9869 2672 9873
rect 2633 9864 2637 9868
rect 2643 9864 2647 9868
rect 2653 9864 2657 9868
rect 2663 9864 2667 9868
rect 2673 9864 2677 9868
rect 2947 9949 2951 9953
rect 2957 9949 2961 9953
rect 2967 9949 2971 9953
rect 2977 9949 2981 9953
rect 2942 9944 2946 9948
rect 2952 9944 2956 9948
rect 2962 9944 2966 9948
rect 2972 9944 2976 9948
rect 2982 9944 2986 9948
rect 2947 9939 2951 9943
rect 2957 9939 2961 9943
rect 2967 9939 2971 9943
rect 2977 9939 2981 9943
rect 2942 9934 2946 9938
rect 2952 9934 2956 9938
rect 2962 9934 2966 9938
rect 2972 9934 2976 9938
rect 2982 9934 2986 9938
rect 2947 9929 2951 9933
rect 2957 9929 2961 9933
rect 2967 9929 2971 9933
rect 2977 9929 2981 9933
rect 2942 9924 2946 9928
rect 2952 9924 2956 9928
rect 2962 9924 2966 9928
rect 2972 9924 2976 9928
rect 2982 9924 2986 9928
rect 2947 9919 2951 9923
rect 2957 9919 2961 9923
rect 2967 9919 2971 9923
rect 2977 9919 2981 9923
rect 2942 9914 2946 9918
rect 2952 9914 2956 9918
rect 2962 9914 2966 9918
rect 2972 9914 2976 9918
rect 2982 9914 2986 9918
rect 2947 9909 2951 9913
rect 2957 9909 2961 9913
rect 2967 9909 2971 9913
rect 2977 9909 2981 9913
rect 2942 9904 2946 9908
rect 2952 9904 2956 9908
rect 2962 9904 2966 9908
rect 2972 9904 2976 9908
rect 2982 9904 2986 9908
rect 2947 9899 2951 9903
rect 2957 9899 2961 9903
rect 2967 9899 2971 9903
rect 2977 9899 2981 9903
rect 2942 9894 2946 9898
rect 2952 9894 2956 9898
rect 2962 9894 2966 9898
rect 2972 9894 2976 9898
rect 2982 9894 2986 9898
rect 2947 9889 2951 9893
rect 2957 9889 2961 9893
rect 2967 9889 2971 9893
rect 2977 9889 2981 9893
rect 2942 9884 2946 9888
rect 2952 9884 2956 9888
rect 2962 9884 2966 9888
rect 2972 9884 2976 9888
rect 2982 9884 2986 9888
rect 2947 9879 2951 9883
rect 2957 9879 2961 9883
rect 2967 9879 2971 9883
rect 2977 9879 2981 9883
rect 2942 9874 2946 9878
rect 2952 9874 2956 9878
rect 2962 9874 2966 9878
rect 2972 9874 2976 9878
rect 2982 9874 2986 9878
rect 2947 9869 2951 9873
rect 2957 9869 2961 9873
rect 2967 9869 2971 9873
rect 2977 9869 2981 9873
rect 2942 9864 2946 9868
rect 2952 9864 2956 9868
rect 2962 9864 2966 9868
rect 2972 9864 2976 9868
rect 2982 9864 2986 9868
rect 3256 9949 3260 9953
rect 3266 9949 3270 9953
rect 3276 9949 3280 9953
rect 3286 9949 3290 9953
rect 3251 9944 3255 9948
rect 3261 9944 3265 9948
rect 3271 9944 3275 9948
rect 3281 9944 3285 9948
rect 3291 9944 3295 9948
rect 3256 9939 3260 9943
rect 3266 9939 3270 9943
rect 3276 9939 3280 9943
rect 3286 9939 3290 9943
rect 3251 9934 3255 9938
rect 3261 9934 3265 9938
rect 3271 9934 3275 9938
rect 3281 9934 3285 9938
rect 3291 9934 3295 9938
rect 3256 9929 3260 9933
rect 3266 9929 3270 9933
rect 3276 9929 3280 9933
rect 3286 9929 3290 9933
rect 3251 9924 3255 9928
rect 3261 9924 3265 9928
rect 3271 9924 3275 9928
rect 3281 9924 3285 9928
rect 3291 9924 3295 9928
rect 3256 9919 3260 9923
rect 3266 9919 3270 9923
rect 3276 9919 3280 9923
rect 3286 9919 3290 9923
rect 3251 9914 3255 9918
rect 3261 9914 3265 9918
rect 3271 9914 3275 9918
rect 3281 9914 3285 9918
rect 3291 9914 3295 9918
rect 3256 9909 3260 9913
rect 3266 9909 3270 9913
rect 3276 9909 3280 9913
rect 3286 9909 3290 9913
rect 3251 9904 3255 9908
rect 3261 9904 3265 9908
rect 3271 9904 3275 9908
rect 3281 9904 3285 9908
rect 3291 9904 3295 9908
rect 3256 9899 3260 9903
rect 3266 9899 3270 9903
rect 3276 9899 3280 9903
rect 3286 9899 3290 9903
rect 3251 9894 3255 9898
rect 3261 9894 3265 9898
rect 3271 9894 3275 9898
rect 3281 9894 3285 9898
rect 3291 9894 3295 9898
rect 3256 9889 3260 9893
rect 3266 9889 3270 9893
rect 3276 9889 3280 9893
rect 3286 9889 3290 9893
rect 3251 9884 3255 9888
rect 3261 9884 3265 9888
rect 3271 9884 3275 9888
rect 3281 9884 3285 9888
rect 3291 9884 3295 9888
rect 3256 9879 3260 9883
rect 3266 9879 3270 9883
rect 3276 9879 3280 9883
rect 3286 9879 3290 9883
rect 3251 9874 3255 9878
rect 3261 9874 3265 9878
rect 3271 9874 3275 9878
rect 3281 9874 3285 9878
rect 3291 9874 3295 9878
rect 3256 9869 3260 9873
rect 3266 9869 3270 9873
rect 3276 9869 3280 9873
rect 3286 9869 3290 9873
rect 3251 9864 3255 9868
rect 3261 9864 3265 9868
rect 3271 9864 3275 9868
rect 3281 9864 3285 9868
rect 3291 9864 3295 9868
rect 3565 9949 3569 9953
rect 3575 9949 3579 9953
rect 3585 9949 3589 9953
rect 3595 9949 3599 9953
rect 3560 9944 3564 9948
rect 3570 9944 3574 9948
rect 3580 9944 3584 9948
rect 3590 9944 3594 9948
rect 3600 9944 3604 9948
rect 3565 9939 3569 9943
rect 3575 9939 3579 9943
rect 3585 9939 3589 9943
rect 3595 9939 3599 9943
rect 3560 9934 3564 9938
rect 3570 9934 3574 9938
rect 3580 9934 3584 9938
rect 3590 9934 3594 9938
rect 3600 9934 3604 9938
rect 3565 9929 3569 9933
rect 3575 9929 3579 9933
rect 3585 9929 3589 9933
rect 3595 9929 3599 9933
rect 3560 9924 3564 9928
rect 3570 9924 3574 9928
rect 3580 9924 3584 9928
rect 3590 9924 3594 9928
rect 3600 9924 3604 9928
rect 3565 9919 3569 9923
rect 3575 9919 3579 9923
rect 3585 9919 3589 9923
rect 3595 9919 3599 9923
rect 3560 9914 3564 9918
rect 3570 9914 3574 9918
rect 3580 9914 3584 9918
rect 3590 9914 3594 9918
rect 3600 9914 3604 9918
rect 3565 9909 3569 9913
rect 3575 9909 3579 9913
rect 3585 9909 3589 9913
rect 3595 9909 3599 9913
rect 3560 9904 3564 9908
rect 3570 9904 3574 9908
rect 3580 9904 3584 9908
rect 3590 9904 3594 9908
rect 3600 9904 3604 9908
rect 3565 9899 3569 9903
rect 3575 9899 3579 9903
rect 3585 9899 3589 9903
rect 3595 9899 3599 9903
rect 3560 9894 3564 9898
rect 3570 9894 3574 9898
rect 3580 9894 3584 9898
rect 3590 9894 3594 9898
rect 3600 9894 3604 9898
rect 3565 9889 3569 9893
rect 3575 9889 3579 9893
rect 3585 9889 3589 9893
rect 3595 9889 3599 9893
rect 3560 9884 3564 9888
rect 3570 9884 3574 9888
rect 3580 9884 3584 9888
rect 3590 9884 3594 9888
rect 3600 9884 3604 9888
rect 3565 9879 3569 9883
rect 3575 9879 3579 9883
rect 3585 9879 3589 9883
rect 3595 9879 3599 9883
rect 3560 9874 3564 9878
rect 3570 9874 3574 9878
rect 3580 9874 3584 9878
rect 3590 9874 3594 9878
rect 3600 9874 3604 9878
rect 3565 9869 3569 9873
rect 3575 9869 3579 9873
rect 3585 9869 3589 9873
rect 3595 9869 3599 9873
rect 3560 9864 3564 9868
rect 3570 9864 3574 9868
rect 3580 9864 3584 9868
rect 3590 9864 3594 9868
rect 3600 9864 3604 9868
rect 3874 9949 3878 9953
rect 3884 9949 3888 9953
rect 3894 9949 3898 9953
rect 3904 9949 3908 9953
rect 3869 9944 3873 9948
rect 3879 9944 3883 9948
rect 3889 9944 3893 9948
rect 3899 9944 3903 9948
rect 3909 9944 3913 9948
rect 3874 9939 3878 9943
rect 3884 9939 3888 9943
rect 3894 9939 3898 9943
rect 3904 9939 3908 9943
rect 3869 9934 3873 9938
rect 3879 9934 3883 9938
rect 3889 9934 3893 9938
rect 3899 9934 3903 9938
rect 3909 9934 3913 9938
rect 3874 9929 3878 9933
rect 3884 9929 3888 9933
rect 3894 9929 3898 9933
rect 3904 9929 3908 9933
rect 3869 9924 3873 9928
rect 3879 9924 3883 9928
rect 3889 9924 3893 9928
rect 3899 9924 3903 9928
rect 3909 9924 3913 9928
rect 3874 9919 3878 9923
rect 3884 9919 3888 9923
rect 3894 9919 3898 9923
rect 3904 9919 3908 9923
rect 3869 9914 3873 9918
rect 3879 9914 3883 9918
rect 3889 9914 3893 9918
rect 3899 9914 3903 9918
rect 3909 9914 3913 9918
rect 3874 9909 3878 9913
rect 3884 9909 3888 9913
rect 3894 9909 3898 9913
rect 3904 9909 3908 9913
rect 3869 9904 3873 9908
rect 3879 9904 3883 9908
rect 3889 9904 3893 9908
rect 3899 9904 3903 9908
rect 3909 9904 3913 9908
rect 3874 9899 3878 9903
rect 3884 9899 3888 9903
rect 3894 9899 3898 9903
rect 3904 9899 3908 9903
rect 3869 9894 3873 9898
rect 3879 9894 3883 9898
rect 3889 9894 3893 9898
rect 3899 9894 3903 9898
rect 3909 9894 3913 9898
rect 3874 9889 3878 9893
rect 3884 9889 3888 9893
rect 3894 9889 3898 9893
rect 3904 9889 3908 9893
rect 3869 9884 3873 9888
rect 3879 9884 3883 9888
rect 3889 9884 3893 9888
rect 3899 9884 3903 9888
rect 3909 9884 3913 9888
rect 3874 9879 3878 9883
rect 3884 9879 3888 9883
rect 3894 9879 3898 9883
rect 3904 9879 3908 9883
rect 3869 9874 3873 9878
rect 3879 9874 3883 9878
rect 3889 9874 3893 9878
rect 3899 9874 3903 9878
rect 3909 9874 3913 9878
rect 3874 9869 3878 9873
rect 3884 9869 3888 9873
rect 3894 9869 3898 9873
rect 3904 9869 3908 9873
rect 3869 9864 3873 9868
rect 3879 9864 3883 9868
rect 3889 9864 3893 9868
rect 3899 9864 3903 9868
rect 3909 9864 3913 9868
rect 1829 9827 1836 9831
rect 1840 9827 1869 9831
rect 2138 9827 2145 9831
rect 2149 9827 2178 9831
rect 2447 9827 2454 9831
rect 2458 9827 2487 9831
rect 2756 9827 2763 9831
rect 2767 9827 2796 9831
rect 3065 9827 3072 9831
rect 3076 9827 3105 9831
rect 3992 9827 3999 9831
rect 4003 9827 4032 9831
rect 1829 9819 1869 9823
rect 2138 9819 2178 9823
rect 2447 9819 2487 9823
rect 2756 9819 2796 9823
rect 3065 9819 3105 9823
rect 3992 9819 4032 9823
rect 1829 9811 1836 9815
rect 1840 9811 1869 9815
rect 1829 9803 1869 9807
rect 1829 9795 1836 9799
rect 1840 9795 1869 9799
rect 1829 9787 1869 9791
rect 2138 9811 2145 9815
rect 2149 9811 2178 9815
rect 2138 9803 2178 9807
rect 2138 9795 2145 9799
rect 2149 9795 2178 9799
rect 2138 9787 2178 9791
rect 2447 9811 2454 9815
rect 2458 9811 2487 9815
rect 2447 9803 2487 9807
rect 2447 9795 2454 9799
rect 2458 9795 2487 9799
rect 2447 9787 2487 9791
rect 2756 9811 2763 9815
rect 2767 9811 2796 9815
rect 2756 9803 2796 9807
rect 2756 9795 2763 9799
rect 2767 9795 2796 9799
rect 2756 9787 2796 9791
rect 3065 9811 3072 9815
rect 3076 9811 3105 9815
rect 3065 9803 3105 9807
rect 3065 9795 3072 9799
rect 3076 9795 3105 9799
rect 3065 9787 3105 9791
rect 3992 9811 3999 9815
rect 4003 9811 4032 9815
rect 3992 9803 4032 9807
rect 3992 9795 3999 9799
rect 4003 9795 4032 9799
rect 3992 9787 4032 9791
rect 1829 9779 1836 9783
rect 1840 9779 1869 9783
rect 2138 9779 2145 9783
rect 2149 9779 2178 9783
rect 2447 9779 2454 9783
rect 2458 9779 2487 9783
rect 2756 9779 2763 9783
rect 2767 9779 2796 9783
rect 3065 9779 3072 9783
rect 3076 9779 3105 9783
rect 3992 9779 3999 9783
rect 4003 9779 4032 9783
rect 423 6332 427 6339
rect 423 6280 427 6328
rect 431 6280 435 6339
rect 439 6280 443 6328
rect 447 6280 451 6339
rect 464 6332 468 6339
rect 464 6280 468 6328
rect 472 6280 476 6339
rect 480 6280 484 6328
rect 488 6280 492 6339
rect 507 6332 511 6339
rect 507 6280 511 6328
rect 515 6280 519 6339
rect 523 6332 527 6339
rect 523 6280 527 6328
rect 531 6280 535 6339
rect 546 6332 550 6339
rect 546 6299 550 6328
rect 554 6299 558 6339
rect 562 6332 566 6339
rect 562 6299 566 6328
rect 570 6299 574 6339
rect 578 6332 582 6339
rect 578 6299 582 6328
rect 586 6299 590 6339
rect 594 6332 598 6339
rect 594 6299 598 6328
rect 2851 9299 2855 9303
rect 2864 9299 2868 9303
rect 2872 9299 2876 9303
rect 2880 9299 2884 9303
rect 2888 9299 2892 9303
rect 2901 9299 2905 9303
rect 2914 9299 2918 9303
rect 2922 9299 2926 9303
rect 2930 9299 2934 9303
rect 2938 9299 2942 9303
rect 2946 9299 2950 9303
rect 2959 9299 2963 9303
rect 2967 9299 2971 9303
rect 2975 9299 2979 9303
rect 2983 9299 2987 9303
rect 2996 9299 3000 9303
rect 3004 9299 3008 9303
rect 3012 9299 3016 9303
rect 3020 9299 3024 9303
rect 3033 9299 3037 9303
rect 3046 9299 3050 9303
rect 3054 9299 3058 9303
rect 3062 9299 3066 9303
rect 3070 9299 3074 9303
rect 3078 9299 3082 9303
rect 3091 9299 3095 9303
rect 3099 9299 3103 9303
rect 3107 9299 3111 9303
rect 3115 9299 3119 9303
rect 3128 9299 3132 9303
rect 3136 9299 3140 9303
rect 3144 9299 3148 9303
rect 3152 9299 3156 9303
rect 3165 9299 3169 9303
rect 3178 9299 3182 9303
rect 3186 9299 3190 9303
rect 3194 9299 3198 9303
rect 3202 9299 3206 9303
rect 3210 9299 3214 9303
rect 3223 9299 3227 9303
rect 3231 9299 3235 9303
rect 3239 9299 3243 9303
rect 3247 9299 3251 9303
rect 3260 9299 3264 9303
rect 3268 9299 3272 9303
rect 3276 9299 3280 9303
rect 3284 9299 3288 9303
rect 3297 9299 3301 9303
rect 3310 9299 3314 9303
rect 3318 9299 3322 9303
rect 3326 9299 3330 9303
rect 3334 9299 3338 9303
rect 3342 9299 3346 9303
rect 3355 9299 3359 9303
rect 3363 9299 3367 9303
rect 3371 9299 3375 9303
rect 3796 9299 3800 9303
rect 3809 9299 3813 9303
rect 3817 9299 3821 9303
rect 3825 9299 3829 9303
rect 3833 9299 3837 9303
rect 3846 9299 3850 9303
rect 3859 9299 3863 9303
rect 3867 9299 3871 9303
rect 3875 9299 3879 9303
rect 3883 9299 3887 9303
rect 3891 9299 3895 9303
rect 3904 9299 3908 9303
rect 3912 9299 3916 9303
rect 3920 9299 3924 9303
rect 3928 9299 3932 9303
rect 3941 9299 3945 9303
rect 3949 9299 3953 9303
rect 3957 9299 3961 9303
rect 3965 9299 3969 9303
rect 3978 9299 3982 9303
rect 3991 9299 3995 9303
rect 3999 9299 4003 9303
rect 4007 9299 4011 9303
rect 4015 9299 4019 9303
rect 4023 9299 4027 9303
rect 4036 9299 4040 9303
rect 4044 9299 4048 9303
rect 4052 9299 4056 9303
rect 4060 9299 4064 9303
rect 4073 9299 4077 9303
rect 4081 9299 4085 9303
rect 4089 9299 4093 9303
rect 4097 9299 4101 9303
rect 4110 9299 4114 9303
rect 4123 9299 4127 9303
rect 4131 9299 4135 9303
rect 4139 9299 4143 9303
rect 4147 9299 4151 9303
rect 4155 9299 4159 9303
rect 4168 9299 4172 9303
rect 4176 9299 4180 9303
rect 4184 9299 4188 9303
rect 4192 9299 4196 9303
rect 4205 9299 4209 9303
rect 4213 9299 4217 9303
rect 4221 9299 4225 9303
rect 4229 9299 4233 9303
rect 4242 9299 4246 9303
rect 4255 9299 4259 9303
rect 4263 9299 4267 9303
rect 4271 9299 4275 9303
rect 4279 9299 4283 9303
rect 4287 9299 4291 9303
rect 4300 9299 4304 9303
rect 4308 9299 4312 9303
rect 4316 9299 4320 9303
rect 2499 9266 2503 9270
rect 2512 9266 2516 9270
rect 2520 9266 2524 9270
rect 2528 9266 2532 9270
rect 2536 9266 2540 9270
rect 2549 9266 2553 9270
rect 2562 9266 2566 9270
rect 2570 9266 2574 9270
rect 2578 9266 2582 9270
rect 2586 9266 2590 9270
rect 2594 9266 2598 9270
rect 2607 9266 2611 9270
rect 2615 9266 2619 9270
rect 2623 9266 2627 9270
rect 3444 9266 3448 9270
rect 3457 9266 3461 9270
rect 3465 9266 3469 9270
rect 3473 9266 3477 9270
rect 3481 9266 3485 9270
rect 3494 9266 3498 9270
rect 3507 9266 3511 9270
rect 3515 9266 3519 9270
rect 3523 9266 3527 9270
rect 3531 9266 3535 9270
rect 3539 9266 3543 9270
rect 3552 9266 3556 9270
rect 3560 9266 3564 9270
rect 3568 9266 3572 9270
rect 2623 9229 2627 9233
rect 2631 9229 2635 9233
rect 3030 9233 3034 9237
rect 3038 9233 3042 9237
rect 3054 9229 3058 9233
rect 3069 9229 3073 9233
rect 3111 9233 3115 9237
rect 3119 9233 3123 9237
rect 3135 9229 3139 9233
rect 3150 9229 3154 9233
rect 3084 9225 3088 9229
rect 3092 9225 3096 9229
rect 2506 9220 2510 9224
rect 2514 9220 2518 9224
rect 2856 9220 2860 9224
rect 2864 9220 2868 9224
rect 2872 9220 2876 9224
rect 2880 9220 2884 9224
rect 2888 9220 2892 9224
rect 2896 9220 2900 9224
rect 2907 9220 2911 9224
rect 2924 9220 2928 9224
rect 2941 9220 2945 9224
rect 2950 9220 2954 9224
rect 2963 9220 2967 9224
rect 2971 9220 2975 9224
rect 2979 9220 2983 9224
rect 2996 9220 3000 9224
rect 3006 9220 3010 9224
rect 3014 9220 3018 9224
rect 3165 9225 3169 9229
rect 3173 9225 3177 9229
rect 3568 9229 3572 9233
rect 3576 9229 3580 9233
rect 3975 9233 3979 9237
rect 3983 9233 3987 9237
rect 3999 9229 4003 9233
rect 4014 9229 4018 9233
rect 4056 9233 4060 9237
rect 4064 9233 4068 9237
rect 4080 9229 4084 9233
rect 4095 9229 4099 9233
rect 4029 9225 4033 9229
rect 4037 9225 4041 9229
rect 3451 9220 3455 9224
rect 3459 9220 3463 9224
rect 3801 9220 3805 9224
rect 3809 9220 3813 9224
rect 3817 9220 3821 9224
rect 3825 9220 3829 9224
rect 3833 9220 3837 9224
rect 3841 9220 3845 9224
rect 3852 9220 3856 9224
rect 3869 9220 3873 9224
rect 3886 9220 3890 9224
rect 3895 9220 3899 9224
rect 3908 9220 3912 9224
rect 3916 9220 3920 9224
rect 3924 9220 3928 9224
rect 3941 9220 3945 9224
rect 3951 9220 3955 9224
rect 3959 9220 3963 9224
rect 4110 9225 4114 9229
rect 4118 9225 4122 9229
rect 2856 9174 2860 9178
rect 2864 9174 2868 9178
rect 2872 9174 2876 9178
rect 2880 9174 2884 9178
rect 2888 9174 2892 9178
rect 2896 9174 2900 9178
rect 2907 9174 2911 9178
rect 2924 9174 2928 9178
rect 2941 9174 2945 9178
rect 2950 9174 2954 9178
rect 2963 9174 2967 9178
rect 2971 9174 2975 9178
rect 2979 9174 2983 9178
rect 2996 9174 3000 9178
rect 3006 9174 3010 9178
rect 3014 9174 3018 9178
rect 2490 9164 2494 9168
rect 2498 9164 2502 9168
rect 2506 9164 2510 9168
rect 2519 9164 2523 9168
rect 2527 9164 2531 9168
rect 2535 9164 2539 9168
rect 2543 9164 2547 9168
rect 2551 9164 2555 9168
rect 2564 9164 2568 9168
rect 2577 9164 2581 9168
rect 2585 9164 2589 9168
rect 2593 9164 2597 9168
rect 2601 9164 2605 9168
rect 2614 9164 2618 9168
rect 3054 9173 3058 9177
rect 3069 9173 3073 9177
rect 3135 9173 3139 9177
rect 3150 9173 3154 9177
rect 3801 9174 3805 9178
rect 3809 9174 3813 9178
rect 3817 9174 3821 9178
rect 3825 9174 3829 9178
rect 3833 9174 3837 9178
rect 3841 9174 3845 9178
rect 3852 9174 3856 9178
rect 3869 9174 3873 9178
rect 3886 9174 3890 9178
rect 3895 9174 3899 9178
rect 3908 9174 3912 9178
rect 3916 9174 3920 9178
rect 3924 9174 3928 9178
rect 3941 9174 3945 9178
rect 3951 9174 3955 9178
rect 3959 9174 3963 9178
rect 3435 9164 3439 9168
rect 3443 9164 3447 9168
rect 3451 9164 3455 9168
rect 3464 9164 3468 9168
rect 3472 9164 3476 9168
rect 3480 9164 3484 9168
rect 3488 9164 3492 9168
rect 3496 9164 3500 9168
rect 3509 9164 3513 9168
rect 3522 9164 3526 9168
rect 3530 9164 3534 9168
rect 3538 9164 3542 9168
rect 3546 9164 3550 9168
rect 3559 9164 3563 9168
rect 3999 9173 4003 9177
rect 4014 9173 4018 9177
rect 4080 9173 4084 9177
rect 4095 9173 4099 9177
rect 3054 9097 3058 9101
rect 3069 9097 3073 9101
rect 3135 9101 3139 9105
rect 3143 9101 3147 9105
rect 3159 9097 3163 9101
rect 3174 9097 3178 9101
rect 3084 9093 3088 9097
rect 3092 9093 3096 9097
rect 2856 9088 2860 9092
rect 2864 9088 2868 9092
rect 2872 9088 2876 9092
rect 2880 9088 2884 9092
rect 2888 9088 2892 9092
rect 2896 9088 2900 9092
rect 2907 9088 2911 9092
rect 2924 9088 2928 9092
rect 2941 9088 2945 9092
rect 2950 9088 2954 9092
rect 2963 9088 2967 9092
rect 2971 9088 2975 9092
rect 2979 9088 2983 9092
rect 2996 9088 3000 9092
rect 3006 9088 3010 9092
rect 3014 9088 3018 9092
rect 3189 9093 3193 9097
rect 3197 9093 3201 9097
rect 3366 9072 3370 9076
rect 3374 9072 3378 9076
rect 3390 9068 3394 9072
rect 3405 9068 3409 9072
rect 3420 9064 3424 9068
rect 3428 9064 3432 9068
rect 3999 9097 4003 9101
rect 4014 9097 4018 9101
rect 4080 9101 4084 9105
rect 4088 9101 4092 9105
rect 4104 9097 4108 9101
rect 4119 9097 4123 9101
rect 4029 9093 4033 9097
rect 4037 9093 4041 9097
rect 3801 9088 3805 9092
rect 3809 9088 3813 9092
rect 3817 9088 3821 9092
rect 3825 9088 3829 9092
rect 3833 9088 3837 9092
rect 3841 9088 3845 9092
rect 3852 9088 3856 9092
rect 3869 9088 3873 9092
rect 3886 9088 3890 9092
rect 3895 9088 3899 9092
rect 3908 9088 3912 9092
rect 3916 9088 3920 9092
rect 3924 9088 3928 9092
rect 3941 9088 3945 9092
rect 3951 9088 3955 9092
rect 3959 9088 3963 9092
rect 4134 9093 4138 9097
rect 4142 9093 4146 9097
rect 2856 9042 2860 9046
rect 2864 9042 2868 9046
rect 2872 9042 2876 9046
rect 2880 9042 2884 9046
rect 2888 9042 2892 9046
rect 2896 9042 2900 9046
rect 2907 9042 2911 9046
rect 2924 9042 2928 9046
rect 2941 9042 2945 9046
rect 2950 9042 2954 9046
rect 2963 9042 2967 9046
rect 2971 9042 2975 9046
rect 2979 9042 2983 9046
rect 2996 9042 3000 9046
rect 3006 9042 3010 9046
rect 3014 9042 3018 9046
rect 3054 9042 3058 9046
rect 3069 9042 3073 9046
rect 3159 9042 3163 9046
rect 3174 9042 3178 9046
rect 3540 9033 3556 9045
rect 3560 9033 3576 9045
rect 3593 9033 3609 9045
rect 3613 9033 3629 9045
rect 3801 9042 3805 9046
rect 3809 9042 3813 9046
rect 3817 9042 3821 9046
rect 3825 9042 3829 9046
rect 3833 9042 3837 9046
rect 3841 9042 3845 9046
rect 3852 9042 3856 9046
rect 3869 9042 3873 9046
rect 3886 9042 3890 9046
rect 3895 9042 3899 9046
rect 3908 9042 3912 9046
rect 3916 9042 3920 9046
rect 3924 9042 3928 9046
rect 3941 9042 3945 9046
rect 3951 9042 3955 9046
rect 3959 9042 3963 9046
rect 3999 9042 4003 9046
rect 4014 9042 4018 9046
rect 4104 9042 4108 9046
rect 4119 9042 4123 9046
rect 3390 9008 3394 9012
rect 3405 9008 3409 9012
rect 3054 8965 3058 8969
rect 3069 8965 3073 8969
rect 3111 8969 3115 8973
rect 3119 8969 3123 8973
rect 3135 8965 3139 8969
rect 3150 8965 3154 8969
rect 3201 8969 3205 8973
rect 3209 8969 3213 8973
rect 3225 8965 3229 8969
rect 3240 8965 3244 8969
rect 3084 8961 3088 8965
rect 3092 8961 3096 8965
rect 2856 8956 2860 8960
rect 2864 8956 2868 8960
rect 2872 8956 2876 8960
rect 2880 8956 2884 8960
rect 2888 8956 2892 8960
rect 2896 8956 2900 8960
rect 2907 8956 2911 8960
rect 2924 8956 2928 8960
rect 2941 8956 2945 8960
rect 2950 8956 2954 8960
rect 2963 8956 2967 8960
rect 2971 8956 2975 8960
rect 2979 8956 2983 8960
rect 2996 8956 3000 8960
rect 3006 8956 3010 8960
rect 3014 8956 3018 8960
rect 3165 8961 3169 8965
rect 3173 8961 3177 8965
rect 3255 8961 3259 8965
rect 3263 8961 3267 8965
rect 3344 8942 3348 8946
rect 3352 8942 3356 8946
rect 3366 8942 3370 8946
rect 3374 8942 3378 8946
rect 3390 8938 3394 8942
rect 3405 8938 3409 8942
rect 3420 8934 3424 8938
rect 3428 8934 3432 8938
rect 3999 8965 4003 8969
rect 4014 8965 4018 8969
rect 4056 8969 4060 8973
rect 4064 8969 4068 8973
rect 4080 8965 4084 8969
rect 4095 8965 4099 8969
rect 4146 8969 4150 8973
rect 4154 8969 4158 8973
rect 4170 8965 4174 8969
rect 4185 8965 4189 8969
rect 4029 8961 4033 8965
rect 4037 8961 4041 8965
rect 3801 8956 3805 8960
rect 3809 8956 3813 8960
rect 3817 8956 3821 8960
rect 3825 8956 3829 8960
rect 3833 8956 3837 8960
rect 3841 8956 3845 8960
rect 3852 8956 3856 8960
rect 3869 8956 3873 8960
rect 3886 8956 3890 8960
rect 3895 8956 3899 8960
rect 3908 8956 3912 8960
rect 3916 8956 3920 8960
rect 3924 8956 3928 8960
rect 3941 8956 3945 8960
rect 3951 8956 3955 8960
rect 3959 8956 3963 8960
rect 4110 8961 4114 8965
rect 4118 8961 4122 8965
rect 4200 8961 4204 8965
rect 4208 8961 4212 8965
rect 2856 8910 2860 8914
rect 2864 8910 2868 8914
rect 2872 8910 2876 8914
rect 2880 8910 2884 8914
rect 2888 8910 2892 8914
rect 2896 8910 2900 8914
rect 2907 8910 2911 8914
rect 2924 8910 2928 8914
rect 2941 8910 2945 8914
rect 2950 8910 2954 8914
rect 2963 8910 2967 8914
rect 2971 8910 2975 8914
rect 2979 8910 2983 8914
rect 2996 8910 3000 8914
rect 3006 8910 3010 8914
rect 3014 8910 3018 8914
rect 3054 8907 3058 8911
rect 3069 8907 3073 8911
rect 3135 8907 3139 8911
rect 3150 8907 3154 8911
rect 3225 8907 3229 8911
rect 3240 8907 3244 8911
rect 3446 8903 3462 8915
rect 3466 8903 3482 8915
rect 3499 8903 3515 8915
rect 3519 8903 3535 8915
rect 3801 8910 3805 8914
rect 3809 8910 3813 8914
rect 3817 8910 3821 8914
rect 3825 8910 3829 8914
rect 3833 8910 3837 8914
rect 3841 8910 3845 8914
rect 3852 8910 3856 8914
rect 3869 8910 3873 8914
rect 3886 8910 3890 8914
rect 3895 8910 3899 8914
rect 3908 8910 3912 8914
rect 3916 8910 3920 8914
rect 3924 8910 3928 8914
rect 3941 8910 3945 8914
rect 3951 8910 3955 8914
rect 3959 8910 3963 8914
rect 3999 8907 4003 8911
rect 4014 8907 4018 8911
rect 4080 8907 4084 8911
rect 4095 8907 4099 8911
rect 4170 8907 4174 8911
rect 4185 8907 4189 8911
rect 3390 8878 3394 8882
rect 3405 8878 3409 8882
rect 3054 8833 3058 8837
rect 3069 8833 3073 8837
rect 3084 8829 3088 8833
rect 3092 8829 3096 8833
rect 2856 8824 2860 8828
rect 2864 8824 2868 8828
rect 2872 8824 2876 8828
rect 2880 8824 2884 8828
rect 2888 8824 2892 8828
rect 2896 8824 2900 8828
rect 2907 8824 2911 8828
rect 2924 8824 2928 8828
rect 2941 8824 2945 8828
rect 2950 8824 2954 8828
rect 2963 8824 2967 8828
rect 2971 8824 2975 8828
rect 2979 8824 2983 8828
rect 2996 8824 3000 8828
rect 3006 8824 3010 8828
rect 3014 8824 3018 8828
rect 3999 8833 4003 8837
rect 4014 8833 4018 8837
rect 4029 8829 4033 8833
rect 4037 8829 4041 8833
rect 3801 8824 3805 8828
rect 3809 8824 3813 8828
rect 3817 8824 3821 8828
rect 3825 8824 3829 8828
rect 3833 8824 3837 8828
rect 3841 8824 3845 8828
rect 3852 8824 3856 8828
rect 3869 8824 3873 8828
rect 3886 8824 3890 8828
rect 3895 8824 3899 8828
rect 3908 8824 3912 8828
rect 3916 8824 3920 8828
rect 3924 8824 3928 8828
rect 3941 8824 3945 8828
rect 3951 8824 3955 8828
rect 3959 8824 3963 8828
rect 2856 8778 2860 8782
rect 2864 8778 2868 8782
rect 2872 8778 2876 8782
rect 2880 8778 2884 8782
rect 2888 8778 2892 8782
rect 2896 8778 2900 8782
rect 2907 8778 2911 8782
rect 2924 8778 2928 8782
rect 2941 8778 2945 8782
rect 2950 8778 2954 8782
rect 2963 8778 2967 8782
rect 2971 8778 2975 8782
rect 2979 8778 2983 8782
rect 2996 8778 3000 8782
rect 3006 8778 3010 8782
rect 3014 8778 3018 8782
rect 3090 8778 3094 8782
rect 3098 8778 3102 8782
rect 3108 8778 3112 8782
rect 3116 8778 3120 8782
rect 3125 8778 3129 8782
rect 3133 8778 3137 8782
rect 3141 8778 3145 8782
rect 3149 8778 3153 8782
rect 3157 8778 3161 8782
rect 3168 8778 3172 8782
rect 3185 8778 3189 8782
rect 3202 8778 3206 8782
rect 3211 8778 3215 8782
rect 3224 8778 3228 8782
rect 3232 8778 3236 8782
rect 3240 8778 3244 8782
rect 3257 8778 3261 8782
rect 3267 8778 3271 8782
rect 3275 8778 3279 8782
rect 2367 8764 2371 8768
rect 2380 8764 2384 8768
rect 2388 8764 2392 8768
rect 2396 8764 2400 8768
rect 2404 8764 2408 8768
rect 2417 8764 2421 8768
rect 2430 8764 2434 8768
rect 2438 8764 2442 8768
rect 2446 8764 2450 8768
rect 2454 8764 2458 8768
rect 2462 8764 2466 8768
rect 2475 8764 2479 8768
rect 2483 8764 2487 8768
rect 2491 8764 2495 8768
rect 2499 8764 2503 8768
rect 2512 8764 2516 8768
rect 2520 8764 2524 8768
rect 2528 8764 2532 8768
rect 2536 8764 2540 8768
rect 2549 8764 2553 8768
rect 2562 8764 2566 8768
rect 2570 8764 2574 8768
rect 2578 8764 2582 8768
rect 2586 8764 2590 8768
rect 2594 8764 2598 8768
rect 2607 8764 2611 8768
rect 2615 8764 2619 8768
rect 2623 8764 2627 8768
rect 2631 8764 2635 8768
rect 2644 8764 2648 8768
rect 2652 8764 2656 8768
rect 2660 8764 2664 8768
rect 2668 8764 2672 8768
rect 2681 8764 2685 8768
rect 2694 8764 2698 8768
rect 2702 8764 2706 8768
rect 2710 8764 2714 8768
rect 2718 8764 2722 8768
rect 2726 8764 2730 8768
rect 2739 8764 2743 8768
rect 2747 8764 2751 8768
rect 2755 8764 2759 8768
rect 3054 8771 3058 8775
rect 3069 8771 3073 8775
rect 3801 8778 3805 8782
rect 3809 8778 3813 8782
rect 3817 8778 3821 8782
rect 3825 8778 3829 8782
rect 3833 8778 3837 8782
rect 3841 8778 3845 8782
rect 3852 8778 3856 8782
rect 3869 8778 3873 8782
rect 3886 8778 3890 8782
rect 3895 8778 3899 8782
rect 3908 8778 3912 8782
rect 3916 8778 3920 8782
rect 3924 8778 3928 8782
rect 3941 8778 3945 8782
rect 3951 8778 3955 8782
rect 3959 8778 3963 8782
rect 4035 8778 4039 8782
rect 4043 8778 4047 8782
rect 4053 8778 4057 8782
rect 4061 8778 4065 8782
rect 4070 8778 4074 8782
rect 4078 8778 4082 8782
rect 4086 8778 4090 8782
rect 4094 8778 4098 8782
rect 4102 8778 4106 8782
rect 4113 8778 4117 8782
rect 4130 8778 4134 8782
rect 4147 8778 4151 8782
rect 4156 8778 4160 8782
rect 4169 8778 4173 8782
rect 4177 8778 4181 8782
rect 4185 8778 4189 8782
rect 4202 8778 4206 8782
rect 4212 8778 4216 8782
rect 4220 8778 4224 8782
rect 3312 8764 3316 8768
rect 3325 8764 3329 8768
rect 3333 8764 3337 8768
rect 3341 8764 3345 8768
rect 3349 8764 3353 8768
rect 3362 8764 3366 8768
rect 3375 8764 3379 8768
rect 3383 8764 3387 8768
rect 3391 8764 3395 8768
rect 3399 8764 3403 8768
rect 3407 8764 3411 8768
rect 3420 8764 3424 8768
rect 3428 8764 3432 8768
rect 3436 8764 3440 8768
rect 3444 8764 3448 8768
rect 3457 8764 3461 8768
rect 3465 8764 3469 8768
rect 3473 8764 3477 8768
rect 3481 8764 3485 8768
rect 3494 8764 3498 8768
rect 3507 8764 3511 8768
rect 3515 8764 3519 8768
rect 3523 8764 3527 8768
rect 3531 8764 3535 8768
rect 3539 8764 3543 8768
rect 3552 8764 3556 8768
rect 3560 8764 3564 8768
rect 3568 8764 3572 8768
rect 3576 8764 3580 8768
rect 3589 8764 3593 8768
rect 3597 8764 3601 8768
rect 3605 8764 3609 8768
rect 3613 8764 3617 8768
rect 3626 8764 3630 8768
rect 3639 8764 3643 8768
rect 3647 8764 3651 8768
rect 3655 8764 3659 8768
rect 3663 8764 3667 8768
rect 3671 8764 3675 8768
rect 3684 8764 3688 8768
rect 3692 8764 3696 8768
rect 3700 8764 3704 8768
rect 3999 8771 4003 8775
rect 4014 8771 4018 8775
rect 2482 8720 2486 8724
rect 2490 8720 2494 8724
rect 2506 8720 2510 8724
rect 2514 8720 2518 8724
rect 3284 8725 3288 8729
rect 3284 8716 3288 8721
rect 3427 8720 3431 8724
rect 3435 8720 3439 8724
rect 3451 8720 3455 8724
rect 3459 8720 3463 8724
rect 4229 8725 4233 8729
rect 4229 8716 4233 8721
rect 2502 8707 2506 8711
rect 2510 8707 2514 8711
rect 3447 8707 3451 8711
rect 3455 8707 3459 8711
rect 2498 8696 2502 8700
rect 3443 8696 3447 8700
rect 2498 8688 2502 8692
rect 2482 8684 2486 8688
rect 2490 8684 2494 8688
rect 2506 8684 2510 8688
rect 2514 8684 2518 8688
rect 3443 8688 3447 8692
rect 3427 8684 3431 8688
rect 3435 8684 3439 8688
rect 3451 8684 3455 8688
rect 3459 8684 3463 8688
rect 3150 8652 3154 8656
rect 3163 8652 3167 8656
rect 3171 8652 3175 8656
rect 3179 8652 3183 8656
rect 3187 8652 3191 8656
rect 3200 8652 3204 8656
rect 3213 8652 3217 8656
rect 3221 8652 3225 8656
rect 3229 8652 3233 8656
rect 3237 8652 3241 8656
rect 3245 8652 3249 8656
rect 3258 8652 3262 8656
rect 3266 8652 3270 8656
rect 3274 8652 3278 8656
rect 4095 8652 4099 8656
rect 4108 8652 4112 8656
rect 4116 8652 4120 8656
rect 4124 8652 4128 8656
rect 4132 8652 4136 8656
rect 4145 8652 4149 8656
rect 4158 8652 4162 8656
rect 4166 8652 4170 8656
rect 4174 8652 4178 8656
rect 4182 8652 4186 8656
rect 4190 8652 4194 8656
rect 4203 8652 4207 8656
rect 4211 8652 4215 8656
rect 4219 8652 4223 8656
rect 2367 8622 2371 8626
rect 2380 8622 2384 8626
rect 2388 8622 2392 8626
rect 2396 8622 2400 8626
rect 2404 8622 2408 8626
rect 2417 8622 2421 8626
rect 2430 8622 2434 8626
rect 2438 8622 2442 8626
rect 2446 8622 2450 8626
rect 2454 8622 2458 8626
rect 2462 8622 2466 8626
rect 2475 8622 2479 8626
rect 2483 8622 2487 8626
rect 2491 8622 2495 8626
rect 2499 8622 2503 8626
rect 2512 8622 2516 8626
rect 2520 8622 2524 8626
rect 2528 8622 2532 8626
rect 2536 8622 2540 8626
rect 2549 8622 2553 8626
rect 2562 8622 2566 8626
rect 2570 8622 2574 8626
rect 2578 8622 2582 8626
rect 2586 8622 2590 8626
rect 2594 8622 2598 8626
rect 2607 8622 2611 8626
rect 2615 8622 2619 8626
rect 2623 8622 2627 8626
rect 2631 8622 2635 8626
rect 2644 8622 2648 8626
rect 2652 8622 2656 8626
rect 2660 8622 2664 8626
rect 2668 8622 2672 8626
rect 2681 8622 2685 8626
rect 2694 8622 2698 8626
rect 2702 8622 2706 8626
rect 2710 8622 2714 8626
rect 2718 8622 2722 8626
rect 2726 8622 2730 8626
rect 2739 8622 2743 8626
rect 2747 8622 2751 8626
rect 2755 8622 2759 8626
rect 3312 8622 3316 8626
rect 3325 8622 3329 8626
rect 3333 8622 3337 8626
rect 3341 8622 3345 8626
rect 3349 8622 3353 8626
rect 3362 8622 3366 8626
rect 3375 8622 3379 8626
rect 3383 8622 3387 8626
rect 3391 8622 3395 8626
rect 3399 8622 3403 8626
rect 3407 8622 3411 8626
rect 3420 8622 3424 8626
rect 3428 8622 3432 8626
rect 3436 8622 3440 8626
rect 3444 8622 3448 8626
rect 3457 8622 3461 8626
rect 3465 8622 3469 8626
rect 3473 8622 3477 8626
rect 3481 8622 3485 8626
rect 3494 8622 3498 8626
rect 3507 8622 3511 8626
rect 3515 8622 3519 8626
rect 3523 8622 3527 8626
rect 3531 8622 3535 8626
rect 3539 8622 3543 8626
rect 3552 8622 3556 8626
rect 3560 8622 3564 8626
rect 3568 8622 3572 8626
rect 3576 8622 3580 8626
rect 3589 8622 3593 8626
rect 3597 8622 3601 8626
rect 3605 8622 3609 8626
rect 3613 8622 3617 8626
rect 3626 8622 3630 8626
rect 3639 8622 3643 8626
rect 3647 8622 3651 8626
rect 3655 8622 3659 8626
rect 3663 8622 3667 8626
rect 3671 8622 3675 8626
rect 3684 8622 3688 8626
rect 3692 8622 3696 8626
rect 3700 8622 3704 8626
rect 3296 8579 3300 8583
rect 3296 8571 3300 8575
rect 4241 8579 4245 8583
rect 4241 8571 4245 8575
rect 3150 8566 3154 8570
rect 3163 8566 3167 8570
rect 3171 8566 3175 8570
rect 3179 8566 3183 8570
rect 3187 8566 3191 8570
rect 3200 8566 3204 8570
rect 3213 8566 3217 8570
rect 3221 8566 3225 8570
rect 3229 8566 3233 8570
rect 3237 8566 3241 8570
rect 3245 8566 3249 8570
rect 3258 8566 3262 8570
rect 3266 8566 3270 8570
rect 3274 8566 3278 8570
rect 4095 8566 4099 8570
rect 4108 8566 4112 8570
rect 4116 8566 4120 8570
rect 4124 8566 4128 8570
rect 4132 8566 4136 8570
rect 4145 8566 4149 8570
rect 4158 8566 4162 8570
rect 4166 8566 4170 8570
rect 4174 8566 4178 8570
rect 4182 8566 4186 8570
rect 4190 8566 4194 8570
rect 4203 8566 4207 8570
rect 4211 8566 4215 8570
rect 4219 8566 4223 8570
rect 2367 8536 2371 8540
rect 2380 8536 2384 8540
rect 2388 8536 2392 8540
rect 2396 8536 2400 8540
rect 2404 8536 2408 8540
rect 2417 8536 2421 8540
rect 2430 8536 2434 8540
rect 2438 8536 2442 8540
rect 2446 8536 2450 8540
rect 2454 8536 2458 8540
rect 2462 8536 2466 8540
rect 2475 8536 2479 8540
rect 2483 8536 2487 8540
rect 2491 8536 2495 8540
rect 2499 8536 2503 8540
rect 2512 8536 2516 8540
rect 2520 8536 2524 8540
rect 2528 8536 2532 8540
rect 2536 8536 2540 8540
rect 2549 8536 2553 8540
rect 2562 8536 2566 8540
rect 2570 8536 2574 8540
rect 2578 8536 2582 8540
rect 2586 8536 2590 8540
rect 2594 8536 2598 8540
rect 2607 8536 2611 8540
rect 2615 8536 2619 8540
rect 2623 8536 2627 8540
rect 2631 8536 2635 8540
rect 2644 8536 2648 8540
rect 2652 8536 2656 8540
rect 2660 8536 2664 8540
rect 2668 8536 2672 8540
rect 2681 8536 2685 8540
rect 2694 8536 2698 8540
rect 2702 8536 2706 8540
rect 2710 8536 2714 8540
rect 2718 8536 2722 8540
rect 2726 8536 2730 8540
rect 2739 8536 2743 8540
rect 2747 8536 2751 8540
rect 2755 8536 2759 8540
rect 3312 8536 3316 8540
rect 3325 8536 3329 8540
rect 3333 8536 3337 8540
rect 3341 8536 3345 8540
rect 3349 8536 3353 8540
rect 3362 8536 3366 8540
rect 3375 8536 3379 8540
rect 3383 8536 3387 8540
rect 3391 8536 3395 8540
rect 3399 8536 3403 8540
rect 3407 8536 3411 8540
rect 3420 8536 3424 8540
rect 3428 8536 3432 8540
rect 3436 8536 3440 8540
rect 3444 8536 3448 8540
rect 3457 8536 3461 8540
rect 3465 8536 3469 8540
rect 3473 8536 3477 8540
rect 3481 8536 3485 8540
rect 3494 8536 3498 8540
rect 3507 8536 3511 8540
rect 3515 8536 3519 8540
rect 3523 8536 3527 8540
rect 3531 8536 3535 8540
rect 3539 8536 3543 8540
rect 3552 8536 3556 8540
rect 3560 8536 3564 8540
rect 3568 8536 3572 8540
rect 3576 8536 3580 8540
rect 3589 8536 3593 8540
rect 3597 8536 3601 8540
rect 3605 8536 3609 8540
rect 3613 8536 3617 8540
rect 3626 8536 3630 8540
rect 3639 8536 3643 8540
rect 3647 8536 3651 8540
rect 3655 8536 3659 8540
rect 3663 8536 3667 8540
rect 3671 8536 3675 8540
rect 3684 8536 3688 8540
rect 3692 8536 3696 8540
rect 3700 8536 3704 8540
rect 2599 8492 2603 8496
rect 2607 8492 2611 8496
rect 2623 8492 2627 8496
rect 2631 8492 2635 8496
rect 3544 8492 3548 8496
rect 3552 8492 3556 8496
rect 3568 8492 3572 8496
rect 3576 8492 3580 8496
rect 2619 8481 2623 8485
rect 2627 8481 2631 8485
rect 3564 8481 3568 8485
rect 3572 8481 3576 8485
rect 2615 8470 2619 8474
rect 3560 8470 3564 8474
rect 2615 8462 2619 8466
rect 3560 8462 3564 8466
rect 2599 8458 2603 8462
rect 2607 8458 2611 8462
rect 2623 8458 2627 8462
rect 2631 8458 2635 8462
rect 3544 8458 3548 8462
rect 3552 8458 3556 8462
rect 3568 8458 3572 8462
rect 3576 8458 3580 8462
rect 2367 8396 2371 8400
rect 2380 8396 2384 8400
rect 2388 8396 2392 8400
rect 2396 8396 2400 8400
rect 2404 8396 2408 8400
rect 2417 8396 2421 8400
rect 2430 8396 2434 8400
rect 2438 8396 2442 8400
rect 2446 8396 2450 8400
rect 2454 8396 2458 8400
rect 2462 8396 2466 8400
rect 2475 8396 2479 8400
rect 2483 8396 2487 8400
rect 2491 8396 2495 8400
rect 2499 8396 2503 8400
rect 2512 8396 2516 8400
rect 2520 8396 2524 8400
rect 2528 8396 2532 8400
rect 2536 8396 2540 8400
rect 2549 8396 2553 8400
rect 2562 8396 2566 8400
rect 2570 8396 2574 8400
rect 2578 8396 2582 8400
rect 2586 8396 2590 8400
rect 2594 8396 2598 8400
rect 2607 8396 2611 8400
rect 2615 8396 2619 8400
rect 2623 8396 2627 8400
rect 2631 8396 2635 8400
rect 2644 8396 2648 8400
rect 2652 8396 2656 8400
rect 2660 8396 2664 8400
rect 2668 8396 2672 8400
rect 2681 8396 2685 8400
rect 2694 8396 2698 8400
rect 2702 8396 2706 8400
rect 2710 8396 2714 8400
rect 2718 8396 2722 8400
rect 2726 8396 2730 8400
rect 2739 8396 2743 8400
rect 2747 8396 2751 8400
rect 2755 8396 2759 8400
rect 3312 8396 3316 8400
rect 3325 8396 3329 8400
rect 3333 8396 3337 8400
rect 3341 8396 3345 8400
rect 3349 8396 3353 8400
rect 3362 8396 3366 8400
rect 3375 8396 3379 8400
rect 3383 8396 3387 8400
rect 3391 8396 3395 8400
rect 3399 8396 3403 8400
rect 3407 8396 3411 8400
rect 3420 8396 3424 8400
rect 3428 8396 3432 8400
rect 3436 8396 3440 8400
rect 3444 8396 3448 8400
rect 3457 8396 3461 8400
rect 3465 8396 3469 8400
rect 3473 8396 3477 8400
rect 3481 8396 3485 8400
rect 3494 8396 3498 8400
rect 3507 8396 3511 8400
rect 3515 8396 3519 8400
rect 3523 8396 3527 8400
rect 3531 8396 3535 8400
rect 3539 8396 3543 8400
rect 3552 8396 3556 8400
rect 3560 8396 3564 8400
rect 3568 8396 3572 8400
rect 3576 8396 3580 8400
rect 3589 8396 3593 8400
rect 3597 8396 3601 8400
rect 3605 8396 3609 8400
rect 3613 8396 3617 8400
rect 3626 8396 3630 8400
rect 3639 8396 3643 8400
rect 3647 8396 3651 8400
rect 3655 8396 3659 8400
rect 3663 8396 3667 8400
rect 3671 8396 3675 8400
rect 3684 8396 3688 8400
rect 3692 8396 3696 8400
rect 3700 8396 3704 8400
rect 2851 8317 2855 8321
rect 2864 8317 2868 8321
rect 2872 8317 2876 8321
rect 2880 8317 2884 8321
rect 2888 8317 2892 8321
rect 2901 8317 2905 8321
rect 2914 8317 2918 8321
rect 2922 8317 2926 8321
rect 2930 8317 2934 8321
rect 2938 8317 2942 8321
rect 2946 8317 2950 8321
rect 2959 8317 2963 8321
rect 2967 8317 2971 8321
rect 2975 8317 2979 8321
rect 2983 8317 2987 8321
rect 2996 8317 3000 8321
rect 3004 8317 3008 8321
rect 3012 8317 3016 8321
rect 3020 8317 3024 8321
rect 3033 8317 3037 8321
rect 3046 8317 3050 8321
rect 3054 8317 3058 8321
rect 3062 8317 3066 8321
rect 3070 8317 3074 8321
rect 3078 8317 3082 8321
rect 3091 8317 3095 8321
rect 3099 8317 3103 8321
rect 3107 8317 3111 8321
rect 3115 8317 3119 8321
rect 3128 8317 3132 8321
rect 3136 8317 3140 8321
rect 3144 8317 3148 8321
rect 3152 8317 3156 8321
rect 3165 8317 3169 8321
rect 3178 8317 3182 8321
rect 3186 8317 3190 8321
rect 3194 8317 3198 8321
rect 3202 8317 3206 8321
rect 3210 8317 3214 8321
rect 3223 8317 3227 8321
rect 3231 8317 3235 8321
rect 3239 8317 3243 8321
rect 3247 8317 3251 8321
rect 3260 8317 3264 8321
rect 3268 8317 3272 8321
rect 3276 8317 3280 8321
rect 3284 8317 3288 8321
rect 3297 8317 3301 8321
rect 3310 8317 3314 8321
rect 3318 8317 3322 8321
rect 3326 8317 3330 8321
rect 3334 8317 3338 8321
rect 3342 8317 3346 8321
rect 3355 8317 3359 8321
rect 3363 8317 3367 8321
rect 3371 8317 3375 8321
rect 3796 8317 3800 8321
rect 3809 8317 3813 8321
rect 3817 8317 3821 8321
rect 3825 8317 3829 8321
rect 3833 8317 3837 8321
rect 3846 8317 3850 8321
rect 3859 8317 3863 8321
rect 3867 8317 3871 8321
rect 3875 8317 3879 8321
rect 3883 8317 3887 8321
rect 3891 8317 3895 8321
rect 3904 8317 3908 8321
rect 3912 8317 3916 8321
rect 3920 8317 3924 8321
rect 3928 8317 3932 8321
rect 3941 8317 3945 8321
rect 3949 8317 3953 8321
rect 3957 8317 3961 8321
rect 3965 8317 3969 8321
rect 3978 8317 3982 8321
rect 3991 8317 3995 8321
rect 3999 8317 4003 8321
rect 4007 8317 4011 8321
rect 4015 8317 4019 8321
rect 4023 8317 4027 8321
rect 4036 8317 4040 8321
rect 4044 8317 4048 8321
rect 4052 8317 4056 8321
rect 4060 8317 4064 8321
rect 4073 8317 4077 8321
rect 4081 8317 4085 8321
rect 4089 8317 4093 8321
rect 4097 8317 4101 8321
rect 4110 8317 4114 8321
rect 4123 8317 4127 8321
rect 4131 8317 4135 8321
rect 4139 8317 4143 8321
rect 4147 8317 4151 8321
rect 4155 8317 4159 8321
rect 4168 8317 4172 8321
rect 4176 8317 4180 8321
rect 4184 8317 4188 8321
rect 4192 8317 4196 8321
rect 4205 8317 4209 8321
rect 4213 8317 4217 8321
rect 4221 8317 4225 8321
rect 4229 8317 4233 8321
rect 4242 8317 4246 8321
rect 4255 8317 4259 8321
rect 4263 8317 4267 8321
rect 4271 8317 4275 8321
rect 4279 8317 4283 8321
rect 4287 8317 4291 8321
rect 4300 8317 4304 8321
rect 4308 8317 4312 8321
rect 4316 8317 4320 8321
rect 2499 8284 2503 8288
rect 2512 8284 2516 8288
rect 2520 8284 2524 8288
rect 2528 8284 2532 8288
rect 2536 8284 2540 8288
rect 2549 8284 2553 8288
rect 2562 8284 2566 8288
rect 2570 8284 2574 8288
rect 2578 8284 2582 8288
rect 2586 8284 2590 8288
rect 2594 8284 2598 8288
rect 2607 8284 2611 8288
rect 2615 8284 2619 8288
rect 2623 8284 2627 8288
rect 3444 8284 3448 8288
rect 3457 8284 3461 8288
rect 3465 8284 3469 8288
rect 3473 8284 3477 8288
rect 3481 8284 3485 8288
rect 3494 8284 3498 8288
rect 3507 8284 3511 8288
rect 3515 8284 3519 8288
rect 3523 8284 3527 8288
rect 3531 8284 3535 8288
rect 3539 8284 3543 8288
rect 3552 8284 3556 8288
rect 3560 8284 3564 8288
rect 3568 8284 3572 8288
rect 2623 8247 2627 8251
rect 2631 8247 2635 8251
rect 3030 8251 3034 8255
rect 3038 8251 3042 8255
rect 3054 8247 3058 8251
rect 3069 8247 3073 8251
rect 3111 8251 3115 8255
rect 3119 8251 3123 8255
rect 3135 8247 3139 8251
rect 3150 8247 3154 8251
rect 3084 8243 3088 8247
rect 3092 8243 3096 8247
rect 2506 8238 2510 8242
rect 2514 8238 2518 8242
rect 2856 8238 2860 8242
rect 2864 8238 2868 8242
rect 2872 8238 2876 8242
rect 2880 8238 2884 8242
rect 2888 8238 2892 8242
rect 2896 8238 2900 8242
rect 2907 8238 2911 8242
rect 2924 8238 2928 8242
rect 2941 8238 2945 8242
rect 2950 8238 2954 8242
rect 2963 8238 2967 8242
rect 2971 8238 2975 8242
rect 2979 8238 2983 8242
rect 2996 8238 3000 8242
rect 3006 8238 3010 8242
rect 3014 8238 3018 8242
rect 3165 8243 3169 8247
rect 3173 8243 3177 8247
rect 3568 8247 3572 8251
rect 3576 8247 3580 8251
rect 3975 8251 3979 8255
rect 3983 8251 3987 8255
rect 3999 8247 4003 8251
rect 4014 8247 4018 8251
rect 4056 8251 4060 8255
rect 4064 8251 4068 8255
rect 4080 8247 4084 8251
rect 4095 8247 4099 8251
rect 4029 8243 4033 8247
rect 4037 8243 4041 8247
rect 3451 8238 3455 8242
rect 3459 8238 3463 8242
rect 3801 8238 3805 8242
rect 3809 8238 3813 8242
rect 3817 8238 3821 8242
rect 3825 8238 3829 8242
rect 3833 8238 3837 8242
rect 3841 8238 3845 8242
rect 3852 8238 3856 8242
rect 3869 8238 3873 8242
rect 3886 8238 3890 8242
rect 3895 8238 3899 8242
rect 3908 8238 3912 8242
rect 3916 8238 3920 8242
rect 3924 8238 3928 8242
rect 3941 8238 3945 8242
rect 3951 8238 3955 8242
rect 3959 8238 3963 8242
rect 4110 8243 4114 8247
rect 4118 8243 4122 8247
rect 2856 8192 2860 8196
rect 2864 8192 2868 8196
rect 2872 8192 2876 8196
rect 2880 8192 2884 8196
rect 2888 8192 2892 8196
rect 2896 8192 2900 8196
rect 2907 8192 2911 8196
rect 2924 8192 2928 8196
rect 2941 8192 2945 8196
rect 2950 8192 2954 8196
rect 2963 8192 2967 8196
rect 2971 8192 2975 8196
rect 2979 8192 2983 8196
rect 2996 8192 3000 8196
rect 3006 8192 3010 8196
rect 3014 8192 3018 8196
rect 2490 8182 2494 8186
rect 2498 8182 2502 8186
rect 2506 8182 2510 8186
rect 2519 8182 2523 8186
rect 2527 8182 2531 8186
rect 2535 8182 2539 8186
rect 2543 8182 2547 8186
rect 2551 8182 2555 8186
rect 2564 8182 2568 8186
rect 2577 8182 2581 8186
rect 2585 8182 2589 8186
rect 2593 8182 2597 8186
rect 2601 8182 2605 8186
rect 2614 8182 2618 8186
rect 3054 8191 3058 8195
rect 3069 8191 3073 8195
rect 3135 8191 3139 8195
rect 3150 8191 3154 8195
rect 3801 8192 3805 8196
rect 3809 8192 3813 8196
rect 3817 8192 3821 8196
rect 3825 8192 3829 8196
rect 3833 8192 3837 8196
rect 3841 8192 3845 8196
rect 3852 8192 3856 8196
rect 3869 8192 3873 8196
rect 3886 8192 3890 8196
rect 3895 8192 3899 8196
rect 3908 8192 3912 8196
rect 3916 8192 3920 8196
rect 3924 8192 3928 8196
rect 3941 8192 3945 8196
rect 3951 8192 3955 8196
rect 3959 8192 3963 8196
rect 3435 8182 3439 8186
rect 3443 8182 3447 8186
rect 3451 8182 3455 8186
rect 3464 8182 3468 8186
rect 3472 8182 3476 8186
rect 3480 8182 3484 8186
rect 3488 8182 3492 8186
rect 3496 8182 3500 8186
rect 3509 8182 3513 8186
rect 3522 8182 3526 8186
rect 3530 8182 3534 8186
rect 3538 8182 3542 8186
rect 3546 8182 3550 8186
rect 3559 8182 3563 8186
rect 3999 8191 4003 8195
rect 4014 8191 4018 8195
rect 4080 8191 4084 8195
rect 4095 8191 4099 8195
rect 3054 8115 3058 8119
rect 3069 8115 3073 8119
rect 3135 8119 3139 8123
rect 3143 8119 3147 8123
rect 3159 8115 3163 8119
rect 3174 8115 3178 8119
rect 3084 8111 3088 8115
rect 3092 8111 3096 8115
rect 2856 8106 2860 8110
rect 2864 8106 2868 8110
rect 2872 8106 2876 8110
rect 2880 8106 2884 8110
rect 2888 8106 2892 8110
rect 2896 8106 2900 8110
rect 2907 8106 2911 8110
rect 2924 8106 2928 8110
rect 2941 8106 2945 8110
rect 2950 8106 2954 8110
rect 2963 8106 2967 8110
rect 2971 8106 2975 8110
rect 2979 8106 2983 8110
rect 2996 8106 3000 8110
rect 3006 8106 3010 8110
rect 3014 8106 3018 8110
rect 3189 8111 3193 8115
rect 3197 8111 3201 8115
rect 3999 8115 4003 8119
rect 4014 8115 4018 8119
rect 4080 8119 4084 8123
rect 4088 8119 4092 8123
rect 4104 8115 4108 8119
rect 4119 8115 4123 8119
rect 4029 8111 4033 8115
rect 4037 8111 4041 8115
rect 3801 8106 3805 8110
rect 3809 8106 3813 8110
rect 3817 8106 3821 8110
rect 3825 8106 3829 8110
rect 3833 8106 3837 8110
rect 3841 8106 3845 8110
rect 3852 8106 3856 8110
rect 3869 8106 3873 8110
rect 3886 8106 3890 8110
rect 3895 8106 3899 8110
rect 3908 8106 3912 8110
rect 3916 8106 3920 8110
rect 3924 8106 3928 8110
rect 3941 8106 3945 8110
rect 3951 8106 3955 8110
rect 3959 8106 3963 8110
rect 4134 8111 4138 8115
rect 4142 8111 4146 8115
rect 2856 8060 2860 8064
rect 2864 8060 2868 8064
rect 2872 8060 2876 8064
rect 2880 8060 2884 8064
rect 2888 8060 2892 8064
rect 2896 8060 2900 8064
rect 2907 8060 2911 8064
rect 2924 8060 2928 8064
rect 2941 8060 2945 8064
rect 2950 8060 2954 8064
rect 2963 8060 2967 8064
rect 2971 8060 2975 8064
rect 2979 8060 2983 8064
rect 2996 8060 3000 8064
rect 3006 8060 3010 8064
rect 3014 8060 3018 8064
rect 3054 8060 3058 8064
rect 3069 8060 3073 8064
rect 3159 8060 3163 8064
rect 3174 8060 3178 8064
rect 3801 8060 3805 8064
rect 3809 8060 3813 8064
rect 3817 8060 3821 8064
rect 3825 8060 3829 8064
rect 3833 8060 3837 8064
rect 3841 8060 3845 8064
rect 3852 8060 3856 8064
rect 3869 8060 3873 8064
rect 3886 8060 3890 8064
rect 3895 8060 3899 8064
rect 3908 8060 3912 8064
rect 3916 8060 3920 8064
rect 3924 8060 3928 8064
rect 3941 8060 3945 8064
rect 3951 8060 3955 8064
rect 3959 8060 3963 8064
rect 3999 8060 4003 8064
rect 4014 8060 4018 8064
rect 4104 8060 4108 8064
rect 4119 8060 4123 8064
rect 3054 7983 3058 7987
rect 3069 7983 3073 7987
rect 3111 7987 3115 7991
rect 3119 7987 3123 7991
rect 3135 7983 3139 7987
rect 3150 7983 3154 7987
rect 3201 7987 3205 7991
rect 3209 7987 3213 7991
rect 3225 7983 3229 7987
rect 3240 7983 3244 7987
rect 3084 7979 3088 7983
rect 3092 7979 3096 7983
rect 2856 7974 2860 7978
rect 2864 7974 2868 7978
rect 2872 7974 2876 7978
rect 2880 7974 2884 7978
rect 2888 7974 2892 7978
rect 2896 7974 2900 7978
rect 2907 7974 2911 7978
rect 2924 7974 2928 7978
rect 2941 7974 2945 7978
rect 2950 7974 2954 7978
rect 2963 7974 2967 7978
rect 2971 7974 2975 7978
rect 2979 7974 2983 7978
rect 2996 7974 3000 7978
rect 3006 7974 3010 7978
rect 3014 7974 3018 7978
rect 3165 7979 3169 7983
rect 3173 7979 3177 7983
rect 3255 7979 3259 7983
rect 3263 7979 3267 7983
rect 3999 7983 4003 7987
rect 4014 7983 4018 7987
rect 4056 7987 4060 7991
rect 4064 7987 4068 7991
rect 4080 7983 4084 7987
rect 4095 7983 4099 7987
rect 4146 7987 4150 7991
rect 4154 7987 4158 7991
rect 4170 7983 4174 7987
rect 4185 7983 4189 7987
rect 4029 7979 4033 7983
rect 4037 7979 4041 7983
rect 3801 7974 3805 7978
rect 3809 7974 3813 7978
rect 3817 7974 3821 7978
rect 3825 7974 3829 7978
rect 3833 7974 3837 7978
rect 3841 7974 3845 7978
rect 3852 7974 3856 7978
rect 3869 7974 3873 7978
rect 3886 7974 3890 7978
rect 3895 7974 3899 7978
rect 3908 7974 3912 7978
rect 3916 7974 3920 7978
rect 3924 7974 3928 7978
rect 3941 7974 3945 7978
rect 3951 7974 3955 7978
rect 3959 7974 3963 7978
rect 4110 7979 4114 7983
rect 4118 7979 4122 7983
rect 4200 7979 4204 7983
rect 4208 7979 4212 7983
rect 2856 7928 2860 7932
rect 2864 7928 2868 7932
rect 2872 7928 2876 7932
rect 2880 7928 2884 7932
rect 2888 7928 2892 7932
rect 2896 7928 2900 7932
rect 2907 7928 2911 7932
rect 2924 7928 2928 7932
rect 2941 7928 2945 7932
rect 2950 7928 2954 7932
rect 2963 7928 2967 7932
rect 2971 7928 2975 7932
rect 2979 7928 2983 7932
rect 2996 7928 3000 7932
rect 3006 7928 3010 7932
rect 3014 7928 3018 7932
rect 3054 7925 3058 7929
rect 3069 7925 3073 7929
rect 3135 7925 3139 7929
rect 3150 7925 3154 7929
rect 3225 7925 3229 7929
rect 3240 7925 3244 7929
rect 3801 7928 3805 7932
rect 3809 7928 3813 7932
rect 3817 7928 3821 7932
rect 3825 7928 3829 7932
rect 3833 7928 3837 7932
rect 3841 7928 3845 7932
rect 3852 7928 3856 7932
rect 3869 7928 3873 7932
rect 3886 7928 3890 7932
rect 3895 7928 3899 7932
rect 3908 7928 3912 7932
rect 3916 7928 3920 7932
rect 3924 7928 3928 7932
rect 3941 7928 3945 7932
rect 3951 7928 3955 7932
rect 3959 7928 3963 7932
rect 3999 7925 4003 7929
rect 4014 7925 4018 7929
rect 4080 7925 4084 7929
rect 4095 7925 4099 7929
rect 4170 7925 4174 7929
rect 4185 7925 4189 7929
rect 3054 7851 3058 7855
rect 3069 7851 3073 7855
rect 3084 7847 3088 7851
rect 3092 7847 3096 7851
rect 2856 7842 2860 7846
rect 2864 7842 2868 7846
rect 2872 7842 2876 7846
rect 2880 7842 2884 7846
rect 2888 7842 2892 7846
rect 2896 7842 2900 7846
rect 2907 7842 2911 7846
rect 2924 7842 2928 7846
rect 2941 7842 2945 7846
rect 2950 7842 2954 7846
rect 2963 7842 2967 7846
rect 2971 7842 2975 7846
rect 2979 7842 2983 7846
rect 2996 7842 3000 7846
rect 3006 7842 3010 7846
rect 3014 7842 3018 7846
rect 3999 7851 4003 7855
rect 4014 7851 4018 7855
rect 4029 7847 4033 7851
rect 4037 7847 4041 7851
rect 3801 7842 3805 7846
rect 3809 7842 3813 7846
rect 3817 7842 3821 7846
rect 3825 7842 3829 7846
rect 3833 7842 3837 7846
rect 3841 7842 3845 7846
rect 3852 7842 3856 7846
rect 3869 7842 3873 7846
rect 3886 7842 3890 7846
rect 3895 7842 3899 7846
rect 3908 7842 3912 7846
rect 3916 7842 3920 7846
rect 3924 7842 3928 7846
rect 3941 7842 3945 7846
rect 3951 7842 3955 7846
rect 3959 7842 3963 7846
rect 2856 7796 2860 7800
rect 2864 7796 2868 7800
rect 2872 7796 2876 7800
rect 2880 7796 2884 7800
rect 2888 7796 2892 7800
rect 2896 7796 2900 7800
rect 2907 7796 2911 7800
rect 2924 7796 2928 7800
rect 2941 7796 2945 7800
rect 2950 7796 2954 7800
rect 2963 7796 2967 7800
rect 2971 7796 2975 7800
rect 2979 7796 2983 7800
rect 2996 7796 3000 7800
rect 3006 7796 3010 7800
rect 3014 7796 3018 7800
rect 3090 7796 3094 7800
rect 3098 7796 3102 7800
rect 3108 7796 3112 7800
rect 3116 7796 3120 7800
rect 3125 7796 3129 7800
rect 3133 7796 3137 7800
rect 3141 7796 3145 7800
rect 3149 7796 3153 7800
rect 3157 7796 3161 7800
rect 3168 7796 3172 7800
rect 3185 7796 3189 7800
rect 3202 7796 3206 7800
rect 3211 7796 3215 7800
rect 3224 7796 3228 7800
rect 3232 7796 3236 7800
rect 3240 7796 3244 7800
rect 3257 7796 3261 7800
rect 3267 7796 3271 7800
rect 3275 7796 3279 7800
rect 2367 7782 2371 7786
rect 2380 7782 2384 7786
rect 2388 7782 2392 7786
rect 2396 7782 2400 7786
rect 2404 7782 2408 7786
rect 2417 7782 2421 7786
rect 2430 7782 2434 7786
rect 2438 7782 2442 7786
rect 2446 7782 2450 7786
rect 2454 7782 2458 7786
rect 2462 7782 2466 7786
rect 2475 7782 2479 7786
rect 2483 7782 2487 7786
rect 2491 7782 2495 7786
rect 2499 7782 2503 7786
rect 2512 7782 2516 7786
rect 2520 7782 2524 7786
rect 2528 7782 2532 7786
rect 2536 7782 2540 7786
rect 2549 7782 2553 7786
rect 2562 7782 2566 7786
rect 2570 7782 2574 7786
rect 2578 7782 2582 7786
rect 2586 7782 2590 7786
rect 2594 7782 2598 7786
rect 2607 7782 2611 7786
rect 2615 7782 2619 7786
rect 2623 7782 2627 7786
rect 2631 7782 2635 7786
rect 2644 7782 2648 7786
rect 2652 7782 2656 7786
rect 2660 7782 2664 7786
rect 2668 7782 2672 7786
rect 2681 7782 2685 7786
rect 2694 7782 2698 7786
rect 2702 7782 2706 7786
rect 2710 7782 2714 7786
rect 2718 7782 2722 7786
rect 2726 7782 2730 7786
rect 2739 7782 2743 7786
rect 2747 7782 2751 7786
rect 2755 7782 2759 7786
rect 3054 7789 3058 7793
rect 3069 7789 3073 7793
rect 3801 7796 3805 7800
rect 3809 7796 3813 7800
rect 3817 7796 3821 7800
rect 3825 7796 3829 7800
rect 3833 7796 3837 7800
rect 3841 7796 3845 7800
rect 3852 7796 3856 7800
rect 3869 7796 3873 7800
rect 3886 7796 3890 7800
rect 3895 7796 3899 7800
rect 3908 7796 3912 7800
rect 3916 7796 3920 7800
rect 3924 7796 3928 7800
rect 3941 7796 3945 7800
rect 3951 7796 3955 7800
rect 3959 7796 3963 7800
rect 4035 7796 4039 7800
rect 4043 7796 4047 7800
rect 4053 7796 4057 7800
rect 4061 7796 4065 7800
rect 4070 7796 4074 7800
rect 4078 7796 4082 7800
rect 4086 7796 4090 7800
rect 4094 7796 4098 7800
rect 4102 7796 4106 7800
rect 4113 7796 4117 7800
rect 4130 7796 4134 7800
rect 4147 7796 4151 7800
rect 4156 7796 4160 7800
rect 4169 7796 4173 7800
rect 4177 7796 4181 7800
rect 4185 7796 4189 7800
rect 4202 7796 4206 7800
rect 4212 7796 4216 7800
rect 4220 7796 4224 7800
rect 3312 7782 3316 7786
rect 3325 7782 3329 7786
rect 3333 7782 3337 7786
rect 3341 7782 3345 7786
rect 3349 7782 3353 7786
rect 3362 7782 3366 7786
rect 3375 7782 3379 7786
rect 3383 7782 3387 7786
rect 3391 7782 3395 7786
rect 3399 7782 3403 7786
rect 3407 7782 3411 7786
rect 3420 7782 3424 7786
rect 3428 7782 3432 7786
rect 3436 7782 3440 7786
rect 3444 7782 3448 7786
rect 3457 7782 3461 7786
rect 3465 7782 3469 7786
rect 3473 7782 3477 7786
rect 3481 7782 3485 7786
rect 3494 7782 3498 7786
rect 3507 7782 3511 7786
rect 3515 7782 3519 7786
rect 3523 7782 3527 7786
rect 3531 7782 3535 7786
rect 3539 7782 3543 7786
rect 3552 7782 3556 7786
rect 3560 7782 3564 7786
rect 3568 7782 3572 7786
rect 3576 7782 3580 7786
rect 3589 7782 3593 7786
rect 3597 7782 3601 7786
rect 3605 7782 3609 7786
rect 3613 7782 3617 7786
rect 3626 7782 3630 7786
rect 3639 7782 3643 7786
rect 3647 7782 3651 7786
rect 3655 7782 3659 7786
rect 3663 7782 3667 7786
rect 3671 7782 3675 7786
rect 3684 7782 3688 7786
rect 3692 7782 3696 7786
rect 3700 7782 3704 7786
rect 3999 7789 4003 7793
rect 4014 7789 4018 7793
rect 2482 7738 2486 7742
rect 2490 7738 2494 7742
rect 2506 7738 2510 7742
rect 2514 7738 2518 7742
rect 3284 7743 3288 7747
rect 3284 7735 3288 7739
rect 3427 7738 3431 7742
rect 3435 7738 3439 7742
rect 3451 7738 3455 7742
rect 3459 7738 3463 7742
rect 4229 7743 4233 7747
rect 4229 7735 4233 7739
rect 2502 7725 2506 7729
rect 2510 7725 2514 7729
rect 3447 7725 3451 7729
rect 3455 7725 3459 7729
rect 2498 7714 2502 7718
rect 3443 7714 3447 7718
rect 2498 7706 2502 7710
rect 2482 7702 2486 7706
rect 2490 7702 2494 7706
rect 2506 7702 2510 7706
rect 2514 7702 2518 7706
rect 3443 7706 3447 7710
rect 3427 7702 3431 7706
rect 3435 7702 3439 7706
rect 3451 7702 3455 7706
rect 3459 7702 3463 7706
rect 3150 7670 3154 7674
rect 3163 7670 3167 7674
rect 3171 7670 3175 7674
rect 3179 7670 3183 7674
rect 3187 7670 3191 7674
rect 3200 7670 3204 7674
rect 3213 7670 3217 7674
rect 3221 7670 3225 7674
rect 3229 7670 3233 7674
rect 3237 7670 3241 7674
rect 3245 7670 3249 7674
rect 3258 7670 3262 7674
rect 3266 7670 3270 7674
rect 3274 7670 3278 7674
rect 4095 7670 4099 7674
rect 4108 7670 4112 7674
rect 4116 7670 4120 7674
rect 4124 7670 4128 7674
rect 4132 7670 4136 7674
rect 4145 7670 4149 7674
rect 4158 7670 4162 7674
rect 4166 7670 4170 7674
rect 4174 7670 4178 7674
rect 4182 7670 4186 7674
rect 4190 7670 4194 7674
rect 4203 7670 4207 7674
rect 4211 7670 4215 7674
rect 4219 7670 4223 7674
rect 2367 7640 2371 7644
rect 2380 7640 2384 7644
rect 2388 7640 2392 7644
rect 2396 7640 2400 7644
rect 2404 7640 2408 7644
rect 2417 7640 2421 7644
rect 2430 7640 2434 7644
rect 2438 7640 2442 7644
rect 2446 7640 2450 7644
rect 2454 7640 2458 7644
rect 2462 7640 2466 7644
rect 2475 7640 2479 7644
rect 2483 7640 2487 7644
rect 2491 7640 2495 7644
rect 2499 7640 2503 7644
rect 2512 7640 2516 7644
rect 2520 7640 2524 7644
rect 2528 7640 2532 7644
rect 2536 7640 2540 7644
rect 2549 7640 2553 7644
rect 2562 7640 2566 7644
rect 2570 7640 2574 7644
rect 2578 7640 2582 7644
rect 2586 7640 2590 7644
rect 2594 7640 2598 7644
rect 2607 7640 2611 7644
rect 2615 7640 2619 7644
rect 2623 7640 2627 7644
rect 2631 7640 2635 7644
rect 2644 7640 2648 7644
rect 2652 7640 2656 7644
rect 2660 7640 2664 7644
rect 2668 7640 2672 7644
rect 2681 7640 2685 7644
rect 2694 7640 2698 7644
rect 2702 7640 2706 7644
rect 2710 7640 2714 7644
rect 2718 7640 2722 7644
rect 2726 7640 2730 7644
rect 2739 7640 2743 7644
rect 2747 7640 2751 7644
rect 2755 7640 2759 7644
rect 3312 7640 3316 7644
rect 3325 7640 3329 7644
rect 3333 7640 3337 7644
rect 3341 7640 3345 7644
rect 3349 7640 3353 7644
rect 3362 7640 3366 7644
rect 3375 7640 3379 7644
rect 3383 7640 3387 7644
rect 3391 7640 3395 7644
rect 3399 7640 3403 7644
rect 3407 7640 3411 7644
rect 3420 7640 3424 7644
rect 3428 7640 3432 7644
rect 3436 7640 3440 7644
rect 3444 7640 3448 7644
rect 3457 7640 3461 7644
rect 3465 7640 3469 7644
rect 3473 7640 3477 7644
rect 3481 7640 3485 7644
rect 3494 7640 3498 7644
rect 3507 7640 3511 7644
rect 3515 7640 3519 7644
rect 3523 7640 3527 7644
rect 3531 7640 3535 7644
rect 3539 7640 3543 7644
rect 3552 7640 3556 7644
rect 3560 7640 3564 7644
rect 3568 7640 3572 7644
rect 3576 7640 3580 7644
rect 3589 7640 3593 7644
rect 3597 7640 3601 7644
rect 3605 7640 3609 7644
rect 3613 7640 3617 7644
rect 3626 7640 3630 7644
rect 3639 7640 3643 7644
rect 3647 7640 3651 7644
rect 3655 7640 3659 7644
rect 3663 7640 3667 7644
rect 3671 7640 3675 7644
rect 3684 7640 3688 7644
rect 3692 7640 3696 7644
rect 3700 7640 3704 7644
rect 3296 7597 3300 7601
rect 3296 7589 3300 7593
rect 4241 7597 4245 7601
rect 4241 7589 4245 7593
rect 3150 7584 3154 7588
rect 3163 7584 3167 7588
rect 3171 7584 3175 7588
rect 3179 7584 3183 7588
rect 3187 7584 3191 7588
rect 3200 7584 3204 7588
rect 3213 7584 3217 7588
rect 3221 7584 3225 7588
rect 3229 7584 3233 7588
rect 3237 7584 3241 7588
rect 3245 7584 3249 7588
rect 3258 7584 3262 7588
rect 3266 7584 3270 7588
rect 3274 7584 3278 7588
rect 4095 7584 4099 7588
rect 4108 7584 4112 7588
rect 4116 7584 4120 7588
rect 4124 7584 4128 7588
rect 4132 7584 4136 7588
rect 4145 7584 4149 7588
rect 4158 7584 4162 7588
rect 4166 7584 4170 7588
rect 4174 7584 4178 7588
rect 4182 7584 4186 7588
rect 4190 7584 4194 7588
rect 4203 7584 4207 7588
rect 4211 7584 4215 7588
rect 4219 7584 4223 7588
rect 2367 7554 2371 7558
rect 2380 7554 2384 7558
rect 2388 7554 2392 7558
rect 2396 7554 2400 7558
rect 2404 7554 2408 7558
rect 2417 7554 2421 7558
rect 2430 7554 2434 7558
rect 2438 7554 2442 7558
rect 2446 7554 2450 7558
rect 2454 7554 2458 7558
rect 2462 7554 2466 7558
rect 2475 7554 2479 7558
rect 2483 7554 2487 7558
rect 2491 7554 2495 7558
rect 2499 7554 2503 7558
rect 2512 7554 2516 7558
rect 2520 7554 2524 7558
rect 2528 7554 2532 7558
rect 2536 7554 2540 7558
rect 2549 7554 2553 7558
rect 2562 7554 2566 7558
rect 2570 7554 2574 7558
rect 2578 7554 2582 7558
rect 2586 7554 2590 7558
rect 2594 7554 2598 7558
rect 2607 7554 2611 7558
rect 2615 7554 2619 7558
rect 2623 7554 2627 7558
rect 2631 7554 2635 7558
rect 2644 7554 2648 7558
rect 2652 7554 2656 7558
rect 2660 7554 2664 7558
rect 2668 7554 2672 7558
rect 2681 7554 2685 7558
rect 2694 7554 2698 7558
rect 2702 7554 2706 7558
rect 2710 7554 2714 7558
rect 2718 7554 2722 7558
rect 2726 7554 2730 7558
rect 2739 7554 2743 7558
rect 2747 7554 2751 7558
rect 2755 7554 2759 7558
rect 3312 7554 3316 7558
rect 3325 7554 3329 7558
rect 3333 7554 3337 7558
rect 3341 7554 3345 7558
rect 3349 7554 3353 7558
rect 3362 7554 3366 7558
rect 3375 7554 3379 7558
rect 3383 7554 3387 7558
rect 3391 7554 3395 7558
rect 3399 7554 3403 7558
rect 3407 7554 3411 7558
rect 3420 7554 3424 7558
rect 3428 7554 3432 7558
rect 3436 7554 3440 7558
rect 3444 7554 3448 7558
rect 3457 7554 3461 7558
rect 3465 7554 3469 7558
rect 3473 7554 3477 7558
rect 3481 7554 3485 7558
rect 3494 7554 3498 7558
rect 3507 7554 3511 7558
rect 3515 7554 3519 7558
rect 3523 7554 3527 7558
rect 3531 7554 3535 7558
rect 3539 7554 3543 7558
rect 3552 7554 3556 7558
rect 3560 7554 3564 7558
rect 3568 7554 3572 7558
rect 3576 7554 3580 7558
rect 3589 7554 3593 7558
rect 3597 7554 3601 7558
rect 3605 7554 3609 7558
rect 3613 7554 3617 7558
rect 3626 7554 3630 7558
rect 3639 7554 3643 7558
rect 3647 7554 3651 7558
rect 3655 7554 3659 7558
rect 3663 7554 3667 7558
rect 3671 7554 3675 7558
rect 3684 7554 3688 7558
rect 3692 7554 3696 7558
rect 3700 7554 3704 7558
rect 2599 7510 2603 7514
rect 2607 7510 2611 7514
rect 2623 7510 2627 7514
rect 2631 7510 2635 7514
rect 3544 7510 3548 7514
rect 3552 7510 3556 7514
rect 3568 7510 3572 7514
rect 3576 7510 3580 7514
rect 2619 7499 2623 7503
rect 2627 7499 2631 7503
rect 3564 7499 3568 7503
rect 3572 7499 3576 7503
rect 2615 7488 2619 7492
rect 3560 7488 3564 7492
rect 2615 7480 2619 7484
rect 3560 7480 3564 7484
rect 2599 7476 2603 7480
rect 2607 7476 2611 7480
rect 2623 7476 2627 7480
rect 2631 7476 2635 7480
rect 3544 7476 3548 7480
rect 3552 7476 3556 7480
rect 3568 7476 3572 7480
rect 3576 7476 3580 7480
rect 3836 7476 3844 7480
rect 3836 7468 3844 7472
rect 2367 7414 2371 7418
rect 2380 7414 2384 7418
rect 2388 7414 2392 7418
rect 2396 7414 2400 7418
rect 2404 7414 2408 7418
rect 2417 7414 2421 7418
rect 2430 7414 2434 7418
rect 2438 7414 2442 7418
rect 2446 7414 2450 7418
rect 2454 7414 2458 7418
rect 2462 7414 2466 7418
rect 2475 7414 2479 7418
rect 2483 7414 2487 7418
rect 2491 7414 2495 7418
rect 2499 7414 2503 7418
rect 2512 7414 2516 7418
rect 2520 7414 2524 7418
rect 2528 7414 2532 7418
rect 2536 7414 2540 7418
rect 2549 7414 2553 7418
rect 2562 7414 2566 7418
rect 2570 7414 2574 7418
rect 2578 7414 2582 7418
rect 2586 7414 2590 7418
rect 2594 7414 2598 7418
rect 2607 7414 2611 7418
rect 2615 7414 2619 7418
rect 2623 7414 2627 7418
rect 2631 7414 2635 7418
rect 2644 7414 2648 7418
rect 2652 7414 2656 7418
rect 2660 7414 2664 7418
rect 2668 7414 2672 7418
rect 2681 7414 2685 7418
rect 2694 7414 2698 7418
rect 2702 7414 2706 7418
rect 2710 7414 2714 7418
rect 2718 7414 2722 7418
rect 2726 7414 2730 7418
rect 2739 7414 2743 7418
rect 2747 7414 2751 7418
rect 2755 7414 2759 7418
rect 3312 7414 3316 7418
rect 3325 7414 3329 7418
rect 3333 7414 3337 7418
rect 3341 7414 3345 7418
rect 3349 7414 3353 7418
rect 3362 7414 3366 7418
rect 3375 7414 3379 7418
rect 3383 7414 3387 7418
rect 3391 7414 3395 7418
rect 3399 7414 3403 7418
rect 3407 7414 3411 7418
rect 3420 7414 3424 7418
rect 3428 7414 3432 7418
rect 3436 7414 3440 7418
rect 3444 7414 3448 7418
rect 3457 7414 3461 7418
rect 3465 7414 3469 7418
rect 3473 7414 3477 7418
rect 3481 7414 3485 7418
rect 3494 7414 3498 7418
rect 3507 7414 3511 7418
rect 3515 7414 3519 7418
rect 3523 7414 3527 7418
rect 3531 7414 3535 7418
rect 3539 7414 3543 7418
rect 3552 7414 3556 7418
rect 3560 7414 3564 7418
rect 3568 7414 3572 7418
rect 3576 7414 3580 7418
rect 3589 7414 3593 7418
rect 3597 7414 3601 7418
rect 3605 7414 3609 7418
rect 3613 7414 3617 7418
rect 3626 7414 3630 7418
rect 3639 7414 3643 7418
rect 3647 7414 3651 7418
rect 3655 7414 3659 7418
rect 3663 7414 3667 7418
rect 3671 7414 3675 7418
rect 3684 7414 3688 7418
rect 3692 7414 3696 7418
rect 3700 7414 3704 7418
rect 1468 6896 1472 6900
rect 1476 6896 1480 6900
rect 1484 6896 1488 6900
rect 1497 6896 1501 6900
rect 1505 6896 1509 6900
rect 1513 6896 1517 6900
rect 1521 6896 1525 6900
rect 1529 6896 1533 6900
rect 1542 6896 1546 6900
rect 1555 6896 1559 6900
rect 1563 6896 1567 6900
rect 1571 6896 1575 6900
rect 1579 6896 1583 6900
rect 1592 6896 1596 6900
rect 1600 6896 1604 6900
rect 1608 6896 1612 6900
rect 1616 6896 1620 6900
rect 1629 6896 1633 6900
rect 1637 6896 1641 6900
rect 1645 6896 1649 6900
rect 1653 6896 1657 6900
rect 1661 6896 1665 6900
rect 1674 6896 1678 6900
rect 1687 6896 1691 6900
rect 1695 6896 1699 6900
rect 1703 6896 1707 6900
rect 1711 6896 1715 6900
rect 1724 6896 1728 6900
rect 1732 6896 1736 6900
rect 1740 6896 1744 6900
rect 1748 6896 1752 6900
rect 1761 6896 1765 6900
rect 1769 6896 1773 6900
rect 1777 6896 1781 6900
rect 1785 6896 1789 6900
rect 1793 6896 1797 6900
rect 1806 6896 1810 6900
rect 1819 6896 1823 6900
rect 1827 6896 1831 6900
rect 1835 6896 1839 6900
rect 1843 6896 1847 6900
rect 1856 6896 1860 6900
rect 2413 6896 2417 6900
rect 2421 6896 2425 6900
rect 2429 6896 2433 6900
rect 2442 6896 2446 6900
rect 2450 6896 2454 6900
rect 2458 6896 2462 6900
rect 2466 6896 2470 6900
rect 2474 6896 2478 6900
rect 2487 6896 2491 6900
rect 2500 6896 2504 6900
rect 2508 6896 2512 6900
rect 2516 6896 2520 6900
rect 2524 6896 2528 6900
rect 2537 6896 2541 6900
rect 2545 6896 2549 6900
rect 2553 6896 2557 6900
rect 2561 6896 2565 6900
rect 2574 6896 2578 6900
rect 2582 6896 2586 6900
rect 2590 6896 2594 6900
rect 2598 6896 2602 6900
rect 2606 6896 2610 6900
rect 2619 6896 2623 6900
rect 2632 6896 2636 6900
rect 2640 6896 2644 6900
rect 2648 6896 2652 6900
rect 2656 6896 2660 6900
rect 2669 6896 2673 6900
rect 2677 6896 2681 6900
rect 2685 6896 2689 6900
rect 2693 6896 2697 6900
rect 2706 6896 2710 6900
rect 2714 6896 2718 6900
rect 2722 6896 2726 6900
rect 2730 6896 2734 6900
rect 2738 6896 2742 6900
rect 2751 6896 2755 6900
rect 2764 6896 2768 6900
rect 2772 6896 2776 6900
rect 2780 6896 2784 6900
rect 2788 6896 2792 6900
rect 2801 6896 2805 6900
rect 1592 6834 1596 6838
rect 1600 6834 1604 6838
rect 1616 6834 1620 6838
rect 1624 6834 1628 6838
rect 2537 6834 2541 6838
rect 2545 6834 2549 6838
rect 2561 6834 2565 6838
rect 2569 6834 2573 6838
rect 1608 6830 1612 6834
rect 2553 6830 2557 6834
rect 1608 6822 1612 6826
rect 2553 6822 2557 6826
rect 1596 6811 1600 6815
rect 1604 6811 1608 6815
rect 2541 6811 2545 6815
rect 2549 6811 2553 6815
rect 1592 6800 1596 6804
rect 1600 6800 1604 6804
rect 1616 6800 1620 6804
rect 1624 6800 1628 6804
rect 2537 6800 2541 6804
rect 2545 6800 2549 6804
rect 2561 6800 2565 6804
rect 2569 6800 2573 6804
rect 1468 6756 1472 6760
rect 1476 6756 1480 6760
rect 1484 6756 1488 6760
rect 1497 6756 1501 6760
rect 1505 6756 1509 6760
rect 1513 6756 1517 6760
rect 1521 6756 1525 6760
rect 1529 6756 1533 6760
rect 1542 6756 1546 6760
rect 1555 6756 1559 6760
rect 1563 6756 1567 6760
rect 1571 6756 1575 6760
rect 1579 6756 1583 6760
rect 1592 6756 1596 6760
rect 1600 6756 1604 6760
rect 1608 6756 1612 6760
rect 1616 6756 1620 6760
rect 1629 6756 1633 6760
rect 1637 6756 1641 6760
rect 1645 6756 1649 6760
rect 1653 6756 1657 6760
rect 1661 6756 1665 6760
rect 1674 6756 1678 6760
rect 1687 6756 1691 6760
rect 1695 6756 1699 6760
rect 1703 6756 1707 6760
rect 1711 6756 1715 6760
rect 1724 6756 1728 6760
rect 1732 6756 1736 6760
rect 1740 6756 1744 6760
rect 1748 6756 1752 6760
rect 1761 6756 1765 6760
rect 1769 6756 1773 6760
rect 1777 6756 1781 6760
rect 1785 6756 1789 6760
rect 1793 6756 1797 6760
rect 1806 6756 1810 6760
rect 1819 6756 1823 6760
rect 1827 6756 1831 6760
rect 1835 6756 1839 6760
rect 1843 6756 1847 6760
rect 1856 6756 1860 6760
rect 2413 6756 2417 6760
rect 2421 6756 2425 6760
rect 2429 6756 2433 6760
rect 2442 6756 2446 6760
rect 2450 6756 2454 6760
rect 2458 6756 2462 6760
rect 2466 6756 2470 6760
rect 2474 6756 2478 6760
rect 2487 6756 2491 6760
rect 2500 6756 2504 6760
rect 2508 6756 2512 6760
rect 2516 6756 2520 6760
rect 2524 6756 2528 6760
rect 2537 6756 2541 6760
rect 2545 6756 2549 6760
rect 2553 6756 2557 6760
rect 2561 6756 2565 6760
rect 2574 6756 2578 6760
rect 2582 6756 2586 6760
rect 2590 6756 2594 6760
rect 2598 6756 2602 6760
rect 2606 6756 2610 6760
rect 2619 6756 2623 6760
rect 2632 6756 2636 6760
rect 2640 6756 2644 6760
rect 2648 6756 2652 6760
rect 2656 6756 2660 6760
rect 2669 6756 2673 6760
rect 2677 6756 2681 6760
rect 2685 6756 2689 6760
rect 2693 6756 2697 6760
rect 2706 6756 2710 6760
rect 2714 6756 2718 6760
rect 2722 6756 2726 6760
rect 2730 6756 2734 6760
rect 2738 6756 2742 6760
rect 2751 6756 2755 6760
rect 2764 6756 2768 6760
rect 2772 6756 2776 6760
rect 2780 6756 2784 6760
rect 2788 6756 2792 6760
rect 2801 6756 2805 6760
rect 949 6726 953 6730
rect 957 6726 961 6730
rect 965 6726 969 6730
rect 978 6726 982 6730
rect 986 6726 990 6730
rect 994 6726 998 6730
rect 1002 6726 1006 6730
rect 1010 6726 1014 6730
rect 1023 6726 1027 6730
rect 1036 6726 1040 6730
rect 1044 6726 1048 6730
rect 1052 6726 1056 6730
rect 1060 6726 1064 6730
rect 1073 6726 1077 6730
rect 1894 6726 1898 6730
rect 1902 6726 1906 6730
rect 1910 6726 1914 6730
rect 1923 6726 1927 6730
rect 1931 6726 1935 6730
rect 1939 6726 1943 6730
rect 1947 6726 1951 6730
rect 1955 6726 1959 6730
rect 1968 6726 1972 6730
rect 1981 6726 1985 6730
rect 1989 6726 1993 6730
rect 1997 6726 2001 6730
rect 2005 6726 2009 6730
rect 2018 6726 2022 6730
rect 927 6721 931 6725
rect 927 6713 931 6717
rect 1872 6721 1876 6725
rect 1872 6713 1876 6717
rect 1468 6670 1472 6674
rect 1476 6670 1480 6674
rect 1484 6670 1488 6674
rect 1497 6670 1501 6674
rect 1505 6670 1509 6674
rect 1513 6670 1517 6674
rect 1521 6670 1525 6674
rect 1529 6670 1533 6674
rect 1542 6670 1546 6674
rect 1555 6670 1559 6674
rect 1563 6670 1567 6674
rect 1571 6670 1575 6674
rect 1579 6670 1583 6674
rect 1592 6670 1596 6674
rect 1600 6670 1604 6674
rect 1608 6670 1612 6674
rect 1616 6670 1620 6674
rect 1629 6670 1633 6674
rect 1637 6670 1641 6674
rect 1645 6670 1649 6674
rect 1653 6670 1657 6674
rect 1661 6670 1665 6674
rect 1674 6670 1678 6674
rect 1687 6670 1691 6674
rect 1695 6670 1699 6674
rect 1703 6670 1707 6674
rect 1711 6670 1715 6674
rect 1724 6670 1728 6674
rect 1732 6670 1736 6674
rect 1740 6670 1744 6674
rect 1748 6670 1752 6674
rect 1761 6670 1765 6674
rect 1769 6670 1773 6674
rect 1777 6670 1781 6674
rect 1785 6670 1789 6674
rect 1793 6670 1797 6674
rect 1806 6670 1810 6674
rect 1819 6670 1823 6674
rect 1827 6670 1831 6674
rect 1835 6670 1839 6674
rect 1843 6670 1847 6674
rect 1856 6670 1860 6674
rect 2413 6670 2417 6674
rect 2421 6670 2425 6674
rect 2429 6670 2433 6674
rect 2442 6670 2446 6674
rect 2450 6670 2454 6674
rect 2458 6670 2462 6674
rect 2466 6670 2470 6674
rect 2474 6670 2478 6674
rect 2487 6670 2491 6674
rect 2500 6670 2504 6674
rect 2508 6670 2512 6674
rect 2516 6670 2520 6674
rect 2524 6670 2528 6674
rect 2537 6670 2541 6674
rect 2545 6670 2549 6674
rect 2553 6670 2557 6674
rect 2561 6670 2565 6674
rect 2574 6670 2578 6674
rect 2582 6670 2586 6674
rect 2590 6670 2594 6674
rect 2598 6670 2602 6674
rect 2606 6670 2610 6674
rect 2619 6670 2623 6674
rect 2632 6670 2636 6674
rect 2640 6670 2644 6674
rect 2648 6670 2652 6674
rect 2656 6670 2660 6674
rect 2669 6670 2673 6674
rect 2677 6670 2681 6674
rect 2685 6670 2689 6674
rect 2693 6670 2697 6674
rect 2706 6670 2710 6674
rect 2714 6670 2718 6674
rect 2722 6670 2726 6674
rect 2730 6670 2734 6674
rect 2738 6670 2742 6674
rect 2751 6670 2755 6674
rect 2764 6670 2768 6674
rect 2772 6670 2776 6674
rect 2780 6670 2784 6674
rect 2788 6670 2792 6674
rect 2801 6670 2805 6674
rect 949 6640 953 6644
rect 957 6640 961 6644
rect 965 6640 969 6644
rect 978 6640 982 6644
rect 986 6640 990 6644
rect 994 6640 998 6644
rect 1002 6640 1006 6644
rect 1010 6640 1014 6644
rect 1023 6640 1027 6644
rect 1036 6640 1040 6644
rect 1044 6640 1048 6644
rect 1052 6640 1056 6644
rect 1060 6640 1064 6644
rect 1073 6640 1077 6644
rect 1894 6640 1898 6644
rect 1902 6640 1906 6644
rect 1910 6640 1914 6644
rect 1923 6640 1927 6644
rect 1931 6640 1935 6644
rect 1939 6640 1943 6644
rect 1947 6640 1951 6644
rect 1955 6640 1959 6644
rect 1968 6640 1972 6644
rect 1981 6640 1985 6644
rect 1989 6640 1993 6644
rect 1997 6640 2001 6644
rect 2005 6640 2009 6644
rect 2018 6640 2022 6644
rect 1709 6608 1713 6612
rect 1717 6608 1721 6612
rect 1733 6608 1737 6612
rect 1741 6608 1745 6612
rect 1725 6604 1729 6608
rect 2654 6608 2658 6612
rect 2662 6608 2666 6612
rect 2678 6608 2682 6612
rect 2686 6608 2690 6612
rect 2670 6604 2674 6608
rect 1725 6596 1729 6600
rect 2670 6596 2674 6600
rect 1713 6585 1717 6589
rect 1721 6585 1725 6589
rect 2658 6585 2662 6589
rect 2666 6585 2670 6589
rect 939 6575 943 6579
rect 939 6567 943 6571
rect 1709 6572 1713 6576
rect 1717 6572 1721 6576
rect 1733 6572 1737 6576
rect 1741 6572 1745 6576
rect 1884 6575 1888 6579
rect 1884 6567 1888 6571
rect 2654 6572 2658 6576
rect 2662 6572 2666 6576
rect 2678 6572 2682 6576
rect 2686 6572 2690 6576
rect 1154 6521 1158 6525
rect 1169 6521 1173 6525
rect 1468 6528 1472 6532
rect 1476 6528 1480 6532
rect 1484 6528 1488 6532
rect 1497 6528 1501 6532
rect 1505 6528 1509 6532
rect 1513 6528 1517 6532
rect 1521 6528 1525 6532
rect 1529 6528 1533 6532
rect 1542 6528 1546 6532
rect 1555 6528 1559 6532
rect 1563 6528 1567 6532
rect 1571 6528 1575 6532
rect 1579 6528 1583 6532
rect 1592 6528 1596 6532
rect 1600 6528 1604 6532
rect 1608 6528 1612 6532
rect 1616 6528 1620 6532
rect 1629 6528 1633 6532
rect 1637 6528 1641 6532
rect 1645 6528 1649 6532
rect 1653 6528 1657 6532
rect 1661 6528 1665 6532
rect 1674 6528 1678 6532
rect 1687 6528 1691 6532
rect 1695 6528 1699 6532
rect 1703 6528 1707 6532
rect 1711 6528 1715 6532
rect 1724 6528 1728 6532
rect 1732 6528 1736 6532
rect 1740 6528 1744 6532
rect 1748 6528 1752 6532
rect 1761 6528 1765 6532
rect 1769 6528 1773 6532
rect 1777 6528 1781 6532
rect 1785 6528 1789 6532
rect 1793 6528 1797 6532
rect 1806 6528 1810 6532
rect 1819 6528 1823 6532
rect 1827 6528 1831 6532
rect 1835 6528 1839 6532
rect 1843 6528 1847 6532
rect 1856 6528 1860 6532
rect 948 6514 952 6518
rect 956 6514 960 6518
rect 966 6514 970 6518
rect 983 6514 987 6518
rect 991 6514 995 6518
rect 999 6514 1003 6518
rect 1012 6514 1016 6518
rect 1021 6514 1025 6518
rect 1038 6514 1042 6518
rect 1055 6514 1059 6518
rect 1066 6514 1070 6518
rect 1074 6514 1078 6518
rect 1082 6514 1086 6518
rect 1090 6514 1094 6518
rect 1098 6514 1102 6518
rect 1107 6514 1111 6518
rect 1115 6514 1119 6518
rect 1125 6514 1129 6518
rect 1133 6514 1137 6518
rect 1209 6514 1213 6518
rect 1217 6514 1221 6518
rect 1227 6514 1231 6518
rect 1244 6514 1248 6518
rect 1252 6514 1256 6518
rect 1260 6514 1264 6518
rect 1273 6514 1277 6518
rect 1282 6514 1286 6518
rect 1299 6514 1303 6518
rect 1316 6514 1320 6518
rect 1327 6514 1331 6518
rect 1335 6514 1339 6518
rect 1343 6514 1347 6518
rect 1351 6514 1355 6518
rect 1359 6514 1363 6518
rect 1367 6514 1371 6518
rect 2099 6521 2103 6525
rect 2114 6521 2118 6525
rect 2413 6528 2417 6532
rect 2421 6528 2425 6532
rect 2429 6528 2433 6532
rect 2442 6528 2446 6532
rect 2450 6528 2454 6532
rect 2458 6528 2462 6532
rect 2466 6528 2470 6532
rect 2474 6528 2478 6532
rect 2487 6528 2491 6532
rect 2500 6528 2504 6532
rect 2508 6528 2512 6532
rect 2516 6528 2520 6532
rect 2524 6528 2528 6532
rect 2537 6528 2541 6532
rect 2545 6528 2549 6532
rect 2553 6528 2557 6532
rect 2561 6528 2565 6532
rect 2574 6528 2578 6532
rect 2582 6528 2586 6532
rect 2590 6528 2594 6532
rect 2598 6528 2602 6532
rect 2606 6528 2610 6532
rect 2619 6528 2623 6532
rect 2632 6528 2636 6532
rect 2640 6528 2644 6532
rect 2648 6528 2652 6532
rect 2656 6528 2660 6532
rect 2669 6528 2673 6532
rect 2677 6528 2681 6532
rect 2685 6528 2689 6532
rect 2693 6528 2697 6532
rect 2706 6528 2710 6532
rect 2714 6528 2718 6532
rect 2722 6528 2726 6532
rect 2730 6528 2734 6532
rect 2738 6528 2742 6532
rect 2751 6528 2755 6532
rect 2764 6528 2768 6532
rect 2772 6528 2776 6532
rect 2780 6528 2784 6532
rect 2788 6528 2792 6532
rect 2801 6528 2805 6532
rect 1893 6514 1897 6518
rect 1901 6514 1905 6518
rect 1911 6514 1915 6518
rect 1928 6514 1932 6518
rect 1936 6514 1940 6518
rect 1944 6514 1948 6518
rect 1957 6514 1961 6518
rect 1966 6514 1970 6518
rect 1983 6514 1987 6518
rect 2000 6514 2004 6518
rect 2011 6514 2015 6518
rect 2019 6514 2023 6518
rect 2027 6514 2031 6518
rect 2035 6514 2039 6518
rect 2043 6514 2047 6518
rect 2052 6514 2056 6518
rect 2060 6514 2064 6518
rect 2070 6514 2074 6518
rect 2078 6514 2082 6518
rect 2154 6514 2158 6518
rect 2162 6514 2166 6518
rect 2172 6514 2176 6518
rect 2189 6514 2193 6518
rect 2197 6514 2201 6518
rect 2205 6514 2209 6518
rect 2218 6514 2222 6518
rect 2227 6514 2231 6518
rect 2244 6514 2248 6518
rect 2261 6514 2265 6518
rect 2272 6514 2276 6518
rect 2280 6514 2284 6518
rect 2288 6514 2292 6518
rect 2296 6514 2300 6518
rect 2304 6514 2308 6518
rect 2312 6514 2316 6518
rect 1209 6468 1213 6472
rect 1217 6468 1221 6472
rect 1227 6468 1231 6472
rect 1244 6468 1248 6472
rect 1252 6468 1256 6472
rect 1260 6468 1264 6472
rect 1273 6468 1277 6472
rect 1282 6468 1286 6472
rect 1299 6468 1303 6472
rect 1316 6468 1320 6472
rect 1327 6468 1331 6472
rect 1335 6468 1339 6472
rect 1343 6468 1347 6472
rect 1351 6468 1355 6472
rect 1359 6468 1363 6472
rect 1367 6468 1371 6472
rect 1131 6463 1135 6467
rect 1139 6463 1143 6467
rect 1154 6459 1158 6463
rect 1169 6459 1173 6463
rect 2154 6468 2158 6472
rect 2162 6468 2166 6472
rect 2172 6468 2176 6472
rect 2189 6468 2193 6472
rect 2197 6468 2201 6472
rect 2205 6468 2209 6472
rect 2218 6468 2222 6472
rect 2227 6468 2231 6472
rect 2244 6468 2248 6472
rect 2261 6468 2265 6472
rect 2272 6468 2276 6472
rect 2280 6468 2284 6472
rect 2288 6468 2292 6472
rect 2296 6468 2300 6472
rect 2304 6468 2308 6472
rect 2312 6468 2316 6472
rect 2076 6463 2080 6467
rect 2084 6463 2088 6467
rect 2099 6459 2103 6463
rect 2114 6459 2118 6463
rect 983 6385 987 6389
rect 998 6385 1002 6389
rect 1073 6385 1077 6389
rect 1088 6385 1092 6389
rect 1154 6385 1158 6389
rect 1169 6385 1173 6389
rect 1209 6382 1213 6386
rect 1217 6382 1221 6386
rect 1227 6382 1231 6386
rect 1244 6382 1248 6386
rect 1252 6382 1256 6386
rect 1260 6382 1264 6386
rect 1273 6382 1277 6386
rect 1282 6382 1286 6386
rect 1299 6382 1303 6386
rect 1316 6382 1320 6386
rect 1327 6382 1331 6386
rect 1335 6382 1339 6386
rect 1343 6382 1347 6386
rect 1351 6382 1355 6386
rect 1359 6382 1363 6386
rect 1367 6382 1371 6386
rect 1928 6385 1932 6389
rect 1943 6385 1947 6389
rect 2018 6385 2022 6389
rect 2033 6385 2037 6389
rect 2099 6385 2103 6389
rect 2114 6385 2118 6389
rect 2154 6382 2158 6386
rect 2162 6382 2166 6386
rect 2172 6382 2176 6386
rect 2189 6382 2193 6386
rect 2197 6382 2201 6386
rect 2205 6382 2209 6386
rect 2218 6382 2222 6386
rect 2227 6382 2231 6386
rect 2244 6382 2248 6386
rect 2261 6382 2265 6386
rect 2272 6382 2276 6386
rect 2280 6382 2284 6386
rect 2288 6382 2292 6386
rect 2296 6382 2300 6386
rect 2304 6382 2308 6386
rect 2312 6382 2316 6386
rect 960 6331 964 6335
rect 968 6331 972 6335
rect 1050 6331 1054 6335
rect 1058 6331 1062 6335
rect 1209 6336 1213 6340
rect 1217 6336 1221 6340
rect 1227 6336 1231 6340
rect 1244 6336 1248 6340
rect 1252 6336 1256 6340
rect 1260 6336 1264 6340
rect 1273 6336 1277 6340
rect 1282 6336 1286 6340
rect 1299 6336 1303 6340
rect 1316 6336 1320 6340
rect 1327 6336 1331 6340
rect 1335 6336 1339 6340
rect 1343 6336 1347 6340
rect 1351 6336 1355 6340
rect 1359 6336 1363 6340
rect 1367 6336 1371 6340
rect 1131 6331 1135 6335
rect 1139 6331 1143 6335
rect 983 6327 987 6331
rect 998 6327 1002 6331
rect 1014 6323 1018 6327
rect 1022 6323 1026 6327
rect 1073 6327 1077 6331
rect 1088 6327 1092 6331
rect 1104 6323 1108 6327
rect 1112 6323 1116 6327
rect 1154 6327 1158 6331
rect 1169 6327 1173 6331
rect 1905 6331 1909 6335
rect 1913 6331 1917 6335
rect 1995 6331 1999 6335
rect 2003 6331 2007 6335
rect 2154 6336 2158 6340
rect 2162 6336 2166 6340
rect 2172 6336 2176 6340
rect 2189 6336 2193 6340
rect 2197 6336 2201 6340
rect 2205 6336 2209 6340
rect 2218 6336 2222 6340
rect 2227 6336 2231 6340
rect 2244 6336 2248 6340
rect 2261 6336 2265 6340
rect 2272 6336 2276 6340
rect 2280 6336 2284 6340
rect 2288 6336 2292 6340
rect 2296 6336 2300 6340
rect 2304 6336 2308 6340
rect 2312 6336 2316 6340
rect 2076 6331 2080 6335
rect 2084 6331 2088 6335
rect 1928 6327 1932 6331
rect 1943 6327 1947 6331
rect 1959 6323 1963 6327
rect 1967 6323 1971 6327
rect 2018 6327 2022 6331
rect 2033 6327 2037 6331
rect 2049 6323 2053 6327
rect 2057 6323 2061 6327
rect 2099 6327 2103 6331
rect 2114 6327 2118 6331
rect 1049 6250 1053 6254
rect 1064 6250 1068 6254
rect 1154 6250 1158 6254
rect 1169 6250 1173 6254
rect 1209 6250 1213 6254
rect 1217 6250 1221 6254
rect 1227 6250 1231 6254
rect 1244 6250 1248 6254
rect 1252 6250 1256 6254
rect 1260 6250 1264 6254
rect 1273 6250 1277 6254
rect 1282 6250 1286 6254
rect 1299 6250 1303 6254
rect 1316 6250 1320 6254
rect 1327 6250 1331 6254
rect 1335 6250 1339 6254
rect 1343 6250 1347 6254
rect 1351 6250 1355 6254
rect 1359 6250 1363 6254
rect 1367 6250 1371 6254
rect 1994 6250 1998 6254
rect 2009 6250 2013 6254
rect 2099 6250 2103 6254
rect 2114 6250 2118 6254
rect 2154 6250 2158 6254
rect 2162 6250 2166 6254
rect 2172 6250 2176 6254
rect 2189 6250 2193 6254
rect 2197 6250 2201 6254
rect 2205 6250 2209 6254
rect 2218 6250 2222 6254
rect 2227 6250 2231 6254
rect 2244 6250 2248 6254
rect 2261 6250 2265 6254
rect 2272 6250 2276 6254
rect 2280 6250 2284 6254
rect 2288 6250 2292 6254
rect 2296 6250 2300 6254
rect 2304 6250 2308 6254
rect 2312 6250 2316 6254
rect 1026 6199 1030 6203
rect 1034 6199 1038 6203
rect 1209 6204 1213 6208
rect 1217 6204 1221 6208
rect 1227 6204 1231 6208
rect 1244 6204 1248 6208
rect 1252 6204 1256 6208
rect 1260 6204 1264 6208
rect 1273 6204 1277 6208
rect 1282 6204 1286 6208
rect 1299 6204 1303 6208
rect 1316 6204 1320 6208
rect 1327 6204 1331 6208
rect 1335 6204 1339 6208
rect 1343 6204 1347 6208
rect 1351 6204 1355 6208
rect 1359 6204 1363 6208
rect 1367 6204 1371 6208
rect 1131 6199 1135 6203
rect 1139 6199 1143 6203
rect 1049 6195 1053 6199
rect 1064 6195 1068 6199
rect 1080 6191 1084 6195
rect 1088 6191 1092 6195
rect 1154 6195 1158 6199
rect 1169 6195 1173 6199
rect 1971 6199 1975 6203
rect 1979 6199 1983 6203
rect 2154 6204 2158 6208
rect 2162 6204 2166 6208
rect 2172 6204 2176 6208
rect 2189 6204 2193 6208
rect 2197 6204 2201 6208
rect 2205 6204 2209 6208
rect 2218 6204 2222 6208
rect 2227 6204 2231 6208
rect 2244 6204 2248 6208
rect 2261 6204 2265 6208
rect 2272 6204 2276 6208
rect 2280 6204 2284 6208
rect 2288 6204 2292 6208
rect 2296 6204 2300 6208
rect 2304 6204 2308 6208
rect 2312 6204 2316 6208
rect 2076 6199 2080 6203
rect 2084 6199 2088 6203
rect 1994 6195 1998 6199
rect 2009 6195 2013 6199
rect 2025 6191 2029 6195
rect 2033 6191 2037 6195
rect 2099 6195 2103 6199
rect 2114 6195 2118 6199
rect 1073 6119 1077 6123
rect 1088 6119 1092 6123
rect 1154 6119 1158 6123
rect 1169 6119 1173 6123
rect 1609 6128 1613 6132
rect 1622 6128 1626 6132
rect 1630 6128 1634 6132
rect 1638 6128 1642 6132
rect 1646 6128 1650 6132
rect 1659 6128 1663 6132
rect 1672 6128 1676 6132
rect 1680 6128 1684 6132
rect 1688 6128 1692 6132
rect 1696 6128 1700 6132
rect 1704 6128 1708 6132
rect 1717 6128 1721 6132
rect 1725 6128 1729 6132
rect 1733 6128 1737 6132
rect 1209 6118 1213 6122
rect 1217 6118 1221 6122
rect 1227 6118 1231 6122
rect 1244 6118 1248 6122
rect 1252 6118 1256 6122
rect 1260 6118 1264 6122
rect 1273 6118 1277 6122
rect 1282 6118 1286 6122
rect 1299 6118 1303 6122
rect 1316 6118 1320 6122
rect 1327 6118 1331 6122
rect 1335 6118 1339 6122
rect 1343 6118 1347 6122
rect 1351 6118 1355 6122
rect 1359 6118 1363 6122
rect 1367 6118 1371 6122
rect 2018 6119 2022 6123
rect 2033 6119 2037 6123
rect 2099 6119 2103 6123
rect 2114 6119 2118 6123
rect 2554 6128 2558 6132
rect 2567 6128 2571 6132
rect 2575 6128 2579 6132
rect 2583 6128 2587 6132
rect 2591 6128 2595 6132
rect 2604 6128 2608 6132
rect 2617 6128 2621 6132
rect 2625 6128 2629 6132
rect 2633 6128 2637 6132
rect 2641 6128 2645 6132
rect 2649 6128 2653 6132
rect 2662 6128 2666 6132
rect 2670 6128 2674 6132
rect 2678 6128 2682 6132
rect 2154 6118 2158 6122
rect 2162 6118 2166 6122
rect 2172 6118 2176 6122
rect 2189 6118 2193 6122
rect 2197 6118 2201 6122
rect 2205 6118 2209 6122
rect 2218 6118 2222 6122
rect 2227 6118 2231 6122
rect 2244 6118 2248 6122
rect 2261 6118 2265 6122
rect 2272 6118 2276 6122
rect 2280 6118 2284 6122
rect 2288 6118 2292 6122
rect 2296 6118 2300 6122
rect 2304 6118 2308 6122
rect 2312 6118 2316 6122
rect 1050 6067 1054 6071
rect 1058 6067 1062 6071
rect 1209 6072 1213 6076
rect 1217 6072 1221 6076
rect 1227 6072 1231 6076
rect 1244 6072 1248 6076
rect 1252 6072 1256 6076
rect 1260 6072 1264 6076
rect 1273 6072 1277 6076
rect 1282 6072 1286 6076
rect 1299 6072 1303 6076
rect 1316 6072 1320 6076
rect 1327 6072 1331 6076
rect 1335 6072 1339 6076
rect 1343 6072 1347 6076
rect 1351 6072 1355 6076
rect 1359 6072 1363 6076
rect 1367 6072 1371 6076
rect 1709 6072 1713 6076
rect 1717 6072 1721 6076
rect 1131 6067 1135 6071
rect 1139 6067 1143 6071
rect 1073 6063 1077 6067
rect 1088 6063 1092 6067
rect 1104 6059 1108 6063
rect 1112 6059 1116 6063
rect 1154 6063 1158 6067
rect 1169 6063 1173 6067
rect 1185 6059 1189 6063
rect 1193 6059 1197 6063
rect 1592 6063 1596 6067
rect 1600 6063 1604 6067
rect 1995 6067 1999 6071
rect 2003 6067 2007 6071
rect 2154 6072 2158 6076
rect 2162 6072 2166 6076
rect 2172 6072 2176 6076
rect 2189 6072 2193 6076
rect 2197 6072 2201 6076
rect 2205 6072 2209 6076
rect 2218 6072 2222 6076
rect 2227 6072 2231 6076
rect 2244 6072 2248 6076
rect 2261 6072 2265 6076
rect 2272 6072 2276 6076
rect 2280 6072 2284 6076
rect 2288 6072 2292 6076
rect 2296 6072 2300 6076
rect 2304 6072 2308 6076
rect 2312 6072 2316 6076
rect 2654 6072 2658 6076
rect 2662 6072 2666 6076
rect 2076 6067 2080 6071
rect 2084 6067 2088 6071
rect 2018 6063 2022 6067
rect 2033 6063 2037 6067
rect 2049 6059 2053 6063
rect 2057 6059 2061 6063
rect 2099 6063 2103 6067
rect 2114 6063 2118 6067
rect 2130 6059 2134 6063
rect 2138 6059 2142 6063
rect 2537 6063 2541 6067
rect 2545 6063 2549 6067
rect 1600 6026 1604 6030
rect 1608 6026 1612 6030
rect 1616 6026 1620 6030
rect 1629 6026 1633 6030
rect 1637 6026 1641 6030
rect 1645 6026 1649 6030
rect 1653 6026 1657 6030
rect 1661 6026 1665 6030
rect 1674 6026 1678 6030
rect 1687 6026 1691 6030
rect 1695 6026 1699 6030
rect 1703 6026 1707 6030
rect 1711 6026 1715 6030
rect 1724 6026 1728 6030
rect 2545 6026 2549 6030
rect 2553 6026 2557 6030
rect 2561 6026 2565 6030
rect 2574 6026 2578 6030
rect 2582 6026 2586 6030
rect 2590 6026 2594 6030
rect 2598 6026 2602 6030
rect 2606 6026 2610 6030
rect 2619 6026 2623 6030
rect 2632 6026 2636 6030
rect 2640 6026 2644 6030
rect 2648 6026 2652 6030
rect 2656 6026 2660 6030
rect 2669 6026 2673 6030
rect 852 5993 856 5997
rect 860 5993 864 5997
rect 868 5993 872 5997
rect 881 5993 885 5997
rect 889 5993 893 5997
rect 897 5993 901 5997
rect 905 5993 909 5997
rect 913 5993 917 5997
rect 926 5993 930 5997
rect 939 5993 943 5997
rect 947 5993 951 5997
rect 955 5993 959 5997
rect 963 5993 967 5997
rect 976 5993 980 5997
rect 984 5993 988 5997
rect 992 5993 996 5997
rect 1000 5993 1004 5997
rect 1013 5993 1017 5997
rect 1021 5993 1025 5997
rect 1029 5993 1033 5997
rect 1037 5993 1041 5997
rect 1045 5993 1049 5997
rect 1058 5993 1062 5997
rect 1071 5993 1075 5997
rect 1079 5993 1083 5997
rect 1087 5993 1091 5997
rect 1095 5993 1099 5997
rect 1108 5993 1112 5997
rect 1116 5993 1120 5997
rect 1124 5993 1128 5997
rect 1132 5993 1136 5997
rect 1145 5993 1149 5997
rect 1153 5993 1157 5997
rect 1161 5993 1165 5997
rect 1169 5993 1173 5997
rect 1177 5993 1181 5997
rect 1190 5993 1194 5997
rect 1203 5993 1207 5997
rect 1211 5993 1215 5997
rect 1219 5993 1223 5997
rect 1227 5993 1231 5997
rect 1240 5993 1244 5997
rect 1248 5993 1252 5997
rect 1256 5993 1260 5997
rect 1264 5993 1268 5997
rect 1277 5993 1281 5997
rect 1285 5993 1289 5997
rect 1293 5993 1297 5997
rect 1301 5993 1305 5997
rect 1309 5993 1313 5997
rect 1322 5993 1326 5997
rect 1335 5993 1339 5997
rect 1343 5993 1347 5997
rect 1351 5993 1355 5997
rect 1359 5993 1363 5997
rect 1372 5993 1376 5997
rect 1797 5993 1801 5997
rect 1805 5993 1809 5997
rect 1813 5993 1817 5997
rect 1826 5993 1830 5997
rect 1834 5993 1838 5997
rect 1842 5993 1846 5997
rect 1850 5993 1854 5997
rect 1858 5993 1862 5997
rect 1871 5993 1875 5997
rect 1884 5993 1888 5997
rect 1892 5993 1896 5997
rect 1900 5993 1904 5997
rect 1908 5993 1912 5997
rect 1921 5993 1925 5997
rect 1929 5993 1933 5997
rect 1937 5993 1941 5997
rect 1945 5993 1949 5997
rect 1958 5993 1962 5997
rect 1966 5993 1970 5997
rect 1974 5993 1978 5997
rect 1982 5993 1986 5997
rect 1990 5993 1994 5997
rect 2003 5993 2007 5997
rect 2016 5993 2020 5997
rect 2024 5993 2028 5997
rect 2032 5993 2036 5997
rect 2040 5993 2044 5997
rect 2053 5993 2057 5997
rect 2061 5993 2065 5997
rect 2069 5993 2073 5997
rect 2077 5993 2081 5997
rect 2090 5993 2094 5997
rect 2098 5993 2102 5997
rect 2106 5993 2110 5997
rect 2114 5993 2118 5997
rect 2122 5993 2126 5997
rect 2135 5993 2139 5997
rect 2148 5993 2152 5997
rect 2156 5993 2160 5997
rect 2164 5993 2168 5997
rect 2172 5993 2176 5997
rect 2185 5993 2189 5997
rect 2193 5993 2197 5997
rect 2201 5993 2205 5997
rect 2209 5993 2213 5997
rect 2222 5993 2226 5997
rect 2230 5993 2234 5997
rect 2238 5993 2242 5997
rect 2246 5993 2250 5997
rect 2254 5993 2258 5997
rect 2267 5993 2271 5997
rect 2280 5993 2284 5997
rect 2288 5993 2292 5997
rect 2296 5993 2300 5997
rect 2304 5993 2308 5997
rect 2317 5993 2321 5997
rect 1468 5914 1472 5918
rect 1476 5914 1480 5918
rect 1484 5914 1488 5918
rect 1497 5914 1501 5918
rect 1505 5914 1509 5918
rect 1513 5914 1517 5918
rect 1521 5914 1525 5918
rect 1529 5914 1533 5918
rect 1542 5914 1546 5918
rect 1555 5914 1559 5918
rect 1563 5914 1567 5918
rect 1571 5914 1575 5918
rect 1579 5914 1583 5918
rect 1592 5914 1596 5918
rect 1600 5914 1604 5918
rect 1608 5914 1612 5918
rect 1616 5914 1620 5918
rect 1629 5914 1633 5918
rect 1637 5914 1641 5918
rect 1645 5914 1649 5918
rect 1653 5914 1657 5918
rect 1661 5914 1665 5918
rect 1674 5914 1678 5918
rect 1687 5914 1691 5918
rect 1695 5914 1699 5918
rect 1703 5914 1707 5918
rect 1711 5914 1715 5918
rect 1724 5914 1728 5918
rect 1732 5914 1736 5918
rect 1740 5914 1744 5918
rect 1748 5914 1752 5918
rect 1761 5914 1765 5918
rect 1769 5914 1773 5918
rect 1777 5914 1781 5918
rect 1785 5914 1789 5918
rect 1793 5914 1797 5918
rect 1806 5914 1810 5918
rect 1819 5914 1823 5918
rect 1827 5914 1831 5918
rect 1835 5914 1839 5918
rect 1843 5914 1847 5918
rect 1856 5914 1860 5918
rect 2413 5914 2417 5918
rect 2421 5914 2425 5918
rect 2429 5914 2433 5918
rect 2442 5914 2446 5918
rect 2450 5914 2454 5918
rect 2458 5914 2462 5918
rect 2466 5914 2470 5918
rect 2474 5914 2478 5918
rect 2487 5914 2491 5918
rect 2500 5914 2504 5918
rect 2508 5914 2512 5918
rect 2516 5914 2520 5918
rect 2524 5914 2528 5918
rect 2537 5914 2541 5918
rect 2545 5914 2549 5918
rect 2553 5914 2557 5918
rect 2561 5914 2565 5918
rect 2574 5914 2578 5918
rect 2582 5914 2586 5918
rect 2590 5914 2594 5918
rect 2598 5914 2602 5918
rect 2606 5914 2610 5918
rect 2619 5914 2623 5918
rect 2632 5914 2636 5918
rect 2640 5914 2644 5918
rect 2648 5914 2652 5918
rect 2656 5914 2660 5918
rect 2669 5914 2673 5918
rect 2677 5914 2681 5918
rect 2685 5914 2689 5918
rect 2693 5914 2697 5918
rect 2706 5914 2710 5918
rect 2714 5914 2718 5918
rect 2722 5914 2726 5918
rect 2730 5914 2734 5918
rect 2738 5914 2742 5918
rect 2751 5914 2755 5918
rect 2764 5914 2768 5918
rect 2772 5914 2776 5918
rect 2780 5914 2784 5918
rect 2788 5914 2792 5918
rect 2801 5914 2805 5918
rect 1592 5852 1596 5856
rect 1600 5852 1604 5856
rect 1616 5852 1620 5856
rect 1624 5852 1628 5856
rect 2537 5852 2541 5856
rect 2545 5852 2549 5856
rect 2561 5852 2565 5856
rect 2569 5852 2573 5856
rect 1608 5848 1612 5852
rect 2553 5848 2557 5852
rect 1608 5840 1612 5844
rect 2553 5840 2557 5844
rect 1596 5829 1600 5833
rect 1604 5829 1608 5833
rect 2541 5829 2545 5833
rect 2549 5829 2553 5833
rect 1592 5818 1596 5822
rect 1600 5818 1604 5822
rect 1616 5818 1620 5822
rect 1624 5818 1628 5822
rect 2537 5818 2541 5822
rect 2545 5818 2549 5822
rect 2561 5818 2565 5822
rect 2569 5818 2573 5822
rect 1468 5774 1472 5778
rect 1476 5774 1480 5778
rect 1484 5774 1488 5778
rect 1497 5774 1501 5778
rect 1505 5774 1509 5778
rect 1513 5774 1517 5778
rect 1521 5774 1525 5778
rect 1529 5774 1533 5778
rect 1542 5774 1546 5778
rect 1555 5774 1559 5778
rect 1563 5774 1567 5778
rect 1571 5774 1575 5778
rect 1579 5774 1583 5778
rect 1592 5774 1596 5778
rect 1600 5774 1604 5778
rect 1608 5774 1612 5778
rect 1616 5774 1620 5778
rect 1629 5774 1633 5778
rect 1637 5774 1641 5778
rect 1645 5774 1649 5778
rect 1653 5774 1657 5778
rect 1661 5774 1665 5778
rect 1674 5774 1678 5778
rect 1687 5774 1691 5778
rect 1695 5774 1699 5778
rect 1703 5774 1707 5778
rect 1711 5774 1715 5778
rect 1724 5774 1728 5778
rect 1732 5774 1736 5778
rect 1740 5774 1744 5778
rect 1748 5774 1752 5778
rect 1761 5774 1765 5778
rect 1769 5774 1773 5778
rect 1777 5774 1781 5778
rect 1785 5774 1789 5778
rect 1793 5774 1797 5778
rect 1806 5774 1810 5778
rect 1819 5774 1823 5778
rect 1827 5774 1831 5778
rect 1835 5774 1839 5778
rect 1843 5774 1847 5778
rect 1856 5774 1860 5778
rect 2413 5774 2417 5778
rect 2421 5774 2425 5778
rect 2429 5774 2433 5778
rect 2442 5774 2446 5778
rect 2450 5774 2454 5778
rect 2458 5774 2462 5778
rect 2466 5774 2470 5778
rect 2474 5774 2478 5778
rect 2487 5774 2491 5778
rect 2500 5774 2504 5778
rect 2508 5774 2512 5778
rect 2516 5774 2520 5778
rect 2524 5774 2528 5778
rect 2537 5774 2541 5778
rect 2545 5774 2549 5778
rect 2553 5774 2557 5778
rect 2561 5774 2565 5778
rect 2574 5774 2578 5778
rect 2582 5774 2586 5778
rect 2590 5774 2594 5778
rect 2598 5774 2602 5778
rect 2606 5774 2610 5778
rect 2619 5774 2623 5778
rect 2632 5774 2636 5778
rect 2640 5774 2644 5778
rect 2648 5774 2652 5778
rect 2656 5774 2660 5778
rect 2669 5774 2673 5778
rect 2677 5774 2681 5778
rect 2685 5774 2689 5778
rect 2693 5774 2697 5778
rect 2706 5774 2710 5778
rect 2714 5774 2718 5778
rect 2722 5774 2726 5778
rect 2730 5774 2734 5778
rect 2738 5774 2742 5778
rect 2751 5774 2755 5778
rect 2764 5774 2768 5778
rect 2772 5774 2776 5778
rect 2780 5774 2784 5778
rect 2788 5774 2792 5778
rect 2801 5774 2805 5778
rect 949 5744 953 5748
rect 957 5744 961 5748
rect 965 5744 969 5748
rect 978 5744 982 5748
rect 986 5744 990 5748
rect 994 5744 998 5748
rect 1002 5744 1006 5748
rect 1010 5744 1014 5748
rect 1023 5744 1027 5748
rect 1036 5744 1040 5748
rect 1044 5744 1048 5748
rect 1052 5744 1056 5748
rect 1060 5744 1064 5748
rect 1073 5744 1077 5748
rect 1894 5744 1898 5748
rect 1902 5744 1906 5748
rect 1910 5744 1914 5748
rect 1923 5744 1927 5748
rect 1931 5744 1935 5748
rect 1939 5744 1943 5748
rect 1947 5744 1951 5748
rect 1955 5744 1959 5748
rect 1968 5744 1972 5748
rect 1981 5744 1985 5748
rect 1989 5744 1993 5748
rect 1997 5744 2001 5748
rect 2005 5744 2009 5748
rect 2018 5744 2022 5748
rect 927 5739 931 5743
rect 927 5731 931 5735
rect 1872 5739 1876 5743
rect 1872 5731 1876 5735
rect 1468 5688 1472 5692
rect 1476 5688 1480 5692
rect 1484 5688 1488 5692
rect 1497 5688 1501 5692
rect 1505 5688 1509 5692
rect 1513 5688 1517 5692
rect 1521 5688 1525 5692
rect 1529 5688 1533 5692
rect 1542 5688 1546 5692
rect 1555 5688 1559 5692
rect 1563 5688 1567 5692
rect 1571 5688 1575 5692
rect 1579 5688 1583 5692
rect 1592 5688 1596 5692
rect 1600 5688 1604 5692
rect 1608 5688 1612 5692
rect 1616 5688 1620 5692
rect 1629 5688 1633 5692
rect 1637 5688 1641 5692
rect 1645 5688 1649 5692
rect 1653 5688 1657 5692
rect 1661 5688 1665 5692
rect 1674 5688 1678 5692
rect 1687 5688 1691 5692
rect 1695 5688 1699 5692
rect 1703 5688 1707 5692
rect 1711 5688 1715 5692
rect 1724 5688 1728 5692
rect 1732 5688 1736 5692
rect 1740 5688 1744 5692
rect 1748 5688 1752 5692
rect 1761 5688 1765 5692
rect 1769 5688 1773 5692
rect 1777 5688 1781 5692
rect 1785 5688 1789 5692
rect 1793 5688 1797 5692
rect 1806 5688 1810 5692
rect 1819 5688 1823 5692
rect 1827 5688 1831 5692
rect 1835 5688 1839 5692
rect 1843 5688 1847 5692
rect 1856 5688 1860 5692
rect 2413 5688 2417 5692
rect 2421 5688 2425 5692
rect 2429 5688 2433 5692
rect 2442 5688 2446 5692
rect 2450 5688 2454 5692
rect 2458 5688 2462 5692
rect 2466 5688 2470 5692
rect 2474 5688 2478 5692
rect 2487 5688 2491 5692
rect 2500 5688 2504 5692
rect 2508 5688 2512 5692
rect 2516 5688 2520 5692
rect 2524 5688 2528 5692
rect 2537 5688 2541 5692
rect 2545 5688 2549 5692
rect 2553 5688 2557 5692
rect 2561 5688 2565 5692
rect 2574 5688 2578 5692
rect 2582 5688 2586 5692
rect 2590 5688 2594 5692
rect 2598 5688 2602 5692
rect 2606 5688 2610 5692
rect 2619 5688 2623 5692
rect 2632 5688 2636 5692
rect 2640 5688 2644 5692
rect 2648 5688 2652 5692
rect 2656 5688 2660 5692
rect 2669 5688 2673 5692
rect 2677 5688 2681 5692
rect 2685 5688 2689 5692
rect 2693 5688 2697 5692
rect 2706 5688 2710 5692
rect 2714 5688 2718 5692
rect 2722 5688 2726 5692
rect 2730 5688 2734 5692
rect 2738 5688 2742 5692
rect 2751 5688 2755 5692
rect 2764 5688 2768 5692
rect 2772 5688 2776 5692
rect 2780 5688 2784 5692
rect 2788 5688 2792 5692
rect 2801 5688 2805 5692
rect 949 5658 953 5662
rect 957 5658 961 5662
rect 965 5658 969 5662
rect 978 5658 982 5662
rect 986 5658 990 5662
rect 994 5658 998 5662
rect 1002 5658 1006 5662
rect 1010 5658 1014 5662
rect 1023 5658 1027 5662
rect 1036 5658 1040 5662
rect 1044 5658 1048 5662
rect 1052 5658 1056 5662
rect 1060 5658 1064 5662
rect 1073 5658 1077 5662
rect 1894 5658 1898 5662
rect 1902 5658 1906 5662
rect 1910 5658 1914 5662
rect 1923 5658 1927 5662
rect 1931 5658 1935 5662
rect 1939 5658 1943 5662
rect 1947 5658 1951 5662
rect 1955 5658 1959 5662
rect 1968 5658 1972 5662
rect 1981 5658 1985 5662
rect 1989 5658 1993 5662
rect 1997 5658 2001 5662
rect 2005 5658 2009 5662
rect 2018 5658 2022 5662
rect 1709 5626 1713 5630
rect 1717 5626 1721 5630
rect 1733 5626 1737 5630
rect 1741 5626 1745 5630
rect 1725 5622 1729 5626
rect 2654 5626 2658 5630
rect 2662 5626 2666 5630
rect 2678 5626 2682 5630
rect 2686 5626 2690 5630
rect 2670 5622 2674 5626
rect 1725 5614 1729 5618
rect 2670 5614 2674 5618
rect 1713 5603 1717 5607
rect 1721 5603 1725 5607
rect 2658 5603 2662 5607
rect 2666 5603 2670 5607
rect 939 5593 943 5598
rect 939 5585 943 5589
rect 1709 5590 1713 5594
rect 1717 5590 1721 5594
rect 1733 5590 1737 5594
rect 1741 5590 1745 5594
rect 1884 5593 1888 5598
rect 1884 5585 1888 5589
rect 2654 5590 2658 5594
rect 2662 5590 2666 5594
rect 2678 5590 2682 5594
rect 2686 5590 2690 5594
rect 1154 5539 1158 5543
rect 1169 5539 1173 5543
rect 1468 5546 1472 5550
rect 1476 5546 1480 5550
rect 1484 5546 1488 5550
rect 1497 5546 1501 5550
rect 1505 5546 1509 5550
rect 1513 5546 1517 5550
rect 1521 5546 1525 5550
rect 1529 5546 1533 5550
rect 1542 5546 1546 5550
rect 1555 5546 1559 5550
rect 1563 5546 1567 5550
rect 1571 5546 1575 5550
rect 1579 5546 1583 5550
rect 1592 5546 1596 5550
rect 1600 5546 1604 5550
rect 1608 5546 1612 5550
rect 1616 5546 1620 5550
rect 1629 5546 1633 5550
rect 1637 5546 1641 5550
rect 1645 5546 1649 5550
rect 1653 5546 1657 5550
rect 1661 5546 1665 5550
rect 1674 5546 1678 5550
rect 1687 5546 1691 5550
rect 1695 5546 1699 5550
rect 1703 5546 1707 5550
rect 1711 5546 1715 5550
rect 1724 5546 1728 5550
rect 1732 5546 1736 5550
rect 1740 5546 1744 5550
rect 1748 5546 1752 5550
rect 1761 5546 1765 5550
rect 1769 5546 1773 5550
rect 1777 5546 1781 5550
rect 1785 5546 1789 5550
rect 1793 5546 1797 5550
rect 1806 5546 1810 5550
rect 1819 5546 1823 5550
rect 1827 5546 1831 5550
rect 1835 5546 1839 5550
rect 1843 5546 1847 5550
rect 1856 5546 1860 5550
rect 948 5532 952 5536
rect 956 5532 960 5536
rect 966 5532 970 5536
rect 983 5532 987 5536
rect 991 5532 995 5536
rect 999 5532 1003 5536
rect 1012 5532 1016 5536
rect 1021 5532 1025 5536
rect 1038 5532 1042 5536
rect 1055 5532 1059 5536
rect 1066 5532 1070 5536
rect 1074 5532 1078 5536
rect 1082 5532 1086 5536
rect 1090 5532 1094 5536
rect 1098 5532 1102 5536
rect 1107 5532 1111 5536
rect 1115 5532 1119 5536
rect 1125 5532 1129 5536
rect 1133 5532 1137 5536
rect 1209 5532 1213 5536
rect 1217 5532 1221 5536
rect 1227 5532 1231 5536
rect 1244 5532 1248 5536
rect 1252 5532 1256 5536
rect 1260 5532 1264 5536
rect 1273 5532 1277 5536
rect 1282 5532 1286 5536
rect 1299 5532 1303 5536
rect 1316 5532 1320 5536
rect 1327 5532 1331 5536
rect 1335 5532 1339 5536
rect 1343 5532 1347 5536
rect 1351 5532 1355 5536
rect 1359 5532 1363 5536
rect 1367 5532 1371 5536
rect 2099 5539 2103 5543
rect 2114 5539 2118 5543
rect 2413 5546 2417 5550
rect 2421 5546 2425 5550
rect 2429 5546 2433 5550
rect 2442 5546 2446 5550
rect 2450 5546 2454 5550
rect 2458 5546 2462 5550
rect 2466 5546 2470 5550
rect 2474 5546 2478 5550
rect 2487 5546 2491 5550
rect 2500 5546 2504 5550
rect 2508 5546 2512 5550
rect 2516 5546 2520 5550
rect 2524 5546 2528 5550
rect 2537 5546 2541 5550
rect 2545 5546 2549 5550
rect 2553 5546 2557 5550
rect 2561 5546 2565 5550
rect 2574 5546 2578 5550
rect 2582 5546 2586 5550
rect 2590 5546 2594 5550
rect 2598 5546 2602 5550
rect 2606 5546 2610 5550
rect 2619 5546 2623 5550
rect 2632 5546 2636 5550
rect 2640 5546 2644 5550
rect 2648 5546 2652 5550
rect 2656 5546 2660 5550
rect 2669 5546 2673 5550
rect 2677 5546 2681 5550
rect 2685 5546 2689 5550
rect 2693 5546 2697 5550
rect 2706 5546 2710 5550
rect 2714 5546 2718 5550
rect 2722 5546 2726 5550
rect 2730 5546 2734 5550
rect 2738 5546 2742 5550
rect 2751 5546 2755 5550
rect 2764 5546 2768 5550
rect 2772 5546 2776 5550
rect 2780 5546 2784 5550
rect 2788 5546 2792 5550
rect 2801 5546 2805 5550
rect 1893 5532 1897 5536
rect 1901 5532 1905 5536
rect 1911 5532 1915 5536
rect 1928 5532 1932 5536
rect 1936 5532 1940 5536
rect 1944 5532 1948 5536
rect 1957 5532 1961 5536
rect 1966 5532 1970 5536
rect 1983 5532 1987 5536
rect 2000 5532 2004 5536
rect 2011 5532 2015 5536
rect 2019 5532 2023 5536
rect 2027 5532 2031 5536
rect 2035 5532 2039 5536
rect 2043 5532 2047 5536
rect 2052 5532 2056 5536
rect 2060 5532 2064 5536
rect 2070 5532 2074 5536
rect 2078 5532 2082 5536
rect 2154 5532 2158 5536
rect 2162 5532 2166 5536
rect 2172 5532 2176 5536
rect 2189 5532 2193 5536
rect 2197 5532 2201 5536
rect 2205 5532 2209 5536
rect 2218 5532 2222 5536
rect 2227 5532 2231 5536
rect 2244 5532 2248 5536
rect 2261 5532 2265 5536
rect 2272 5532 2276 5536
rect 2280 5532 2284 5536
rect 2288 5532 2292 5536
rect 2296 5532 2300 5536
rect 2304 5532 2308 5536
rect 2312 5532 2316 5536
rect 1209 5486 1213 5490
rect 1217 5486 1221 5490
rect 1227 5486 1231 5490
rect 1244 5486 1248 5490
rect 1252 5486 1256 5490
rect 1260 5486 1264 5490
rect 1273 5486 1277 5490
rect 1282 5486 1286 5490
rect 1299 5486 1303 5490
rect 1316 5486 1320 5490
rect 1327 5486 1331 5490
rect 1335 5486 1339 5490
rect 1343 5486 1347 5490
rect 1351 5486 1355 5490
rect 1359 5486 1363 5490
rect 1367 5486 1371 5490
rect 1131 5481 1135 5485
rect 1139 5481 1143 5485
rect 1154 5477 1158 5481
rect 1169 5477 1173 5481
rect 2154 5486 2158 5490
rect 2162 5486 2166 5490
rect 2172 5486 2176 5490
rect 2189 5486 2193 5490
rect 2197 5486 2201 5490
rect 2205 5486 2209 5490
rect 2218 5486 2222 5490
rect 2227 5486 2231 5490
rect 2244 5486 2248 5490
rect 2261 5486 2265 5490
rect 2272 5486 2276 5490
rect 2280 5486 2284 5490
rect 2288 5486 2292 5490
rect 2296 5486 2300 5490
rect 2304 5486 2308 5490
rect 2312 5486 2316 5490
rect 2076 5481 2080 5485
rect 2084 5481 2088 5485
rect 2099 5477 2103 5481
rect 2114 5477 2118 5481
rect 1763 5432 1767 5436
rect 1778 5432 1782 5436
rect 983 5403 987 5407
rect 998 5403 1002 5407
rect 1073 5403 1077 5407
rect 1088 5403 1092 5407
rect 1154 5403 1158 5407
rect 1169 5403 1173 5407
rect 1209 5400 1213 5404
rect 1217 5400 1221 5404
rect 1227 5400 1231 5404
rect 1244 5400 1248 5404
rect 1252 5400 1256 5404
rect 1260 5400 1264 5404
rect 1273 5400 1277 5404
rect 1282 5400 1286 5404
rect 1299 5400 1303 5404
rect 1316 5400 1320 5404
rect 1327 5400 1331 5404
rect 1335 5400 1339 5404
rect 1343 5400 1347 5404
rect 1351 5400 1355 5404
rect 1359 5400 1363 5404
rect 1367 5400 1371 5404
rect 1637 5399 1653 5411
rect 1657 5399 1673 5411
rect 1690 5399 1706 5411
rect 1710 5399 1726 5411
rect 1928 5403 1932 5407
rect 1943 5403 1947 5407
rect 2018 5403 2022 5407
rect 2033 5403 2037 5407
rect 2099 5403 2103 5407
rect 2114 5403 2118 5407
rect 2154 5400 2158 5404
rect 2162 5400 2166 5404
rect 2172 5400 2176 5404
rect 2189 5400 2193 5404
rect 2197 5400 2201 5404
rect 2205 5400 2209 5404
rect 2218 5400 2222 5404
rect 2227 5400 2231 5404
rect 2244 5400 2248 5404
rect 2261 5400 2265 5404
rect 2272 5400 2276 5404
rect 2280 5400 2284 5404
rect 2288 5400 2292 5404
rect 2296 5400 2300 5404
rect 2304 5400 2308 5404
rect 2312 5400 2316 5404
rect 960 5349 964 5353
rect 968 5349 972 5353
rect 1050 5349 1054 5353
rect 1058 5349 1062 5353
rect 1209 5354 1213 5358
rect 1217 5354 1221 5358
rect 1227 5354 1231 5358
rect 1244 5354 1248 5358
rect 1252 5354 1256 5358
rect 1260 5354 1264 5358
rect 1273 5354 1277 5358
rect 1282 5354 1286 5358
rect 1299 5354 1303 5358
rect 1316 5354 1320 5358
rect 1327 5354 1331 5358
rect 1335 5354 1339 5358
rect 1343 5354 1347 5358
rect 1351 5354 1355 5358
rect 1359 5354 1363 5358
rect 1367 5354 1371 5358
rect 1131 5349 1135 5353
rect 1139 5349 1143 5353
rect 983 5345 987 5349
rect 998 5345 1002 5349
rect 1014 5341 1018 5345
rect 1022 5341 1026 5345
rect 1073 5345 1077 5349
rect 1088 5345 1092 5349
rect 1104 5341 1108 5345
rect 1112 5341 1116 5345
rect 1154 5345 1158 5349
rect 1169 5345 1173 5349
rect 1740 5376 1744 5380
rect 1748 5376 1752 5380
rect 1763 5372 1767 5376
rect 1778 5372 1782 5376
rect 1794 5368 1798 5372
rect 1802 5368 1806 5372
rect 1816 5368 1820 5372
rect 1824 5368 1828 5372
rect 1905 5349 1909 5353
rect 1913 5349 1917 5353
rect 1995 5349 1999 5353
rect 2003 5349 2007 5353
rect 2154 5354 2158 5358
rect 2162 5354 2166 5358
rect 2172 5354 2176 5358
rect 2189 5354 2193 5358
rect 2197 5354 2201 5358
rect 2205 5354 2209 5358
rect 2218 5354 2222 5358
rect 2227 5354 2231 5358
rect 2244 5354 2248 5358
rect 2261 5354 2265 5358
rect 2272 5354 2276 5358
rect 2280 5354 2284 5358
rect 2288 5354 2292 5358
rect 2296 5354 2300 5358
rect 2304 5354 2308 5358
rect 2312 5354 2316 5358
rect 2076 5349 2080 5353
rect 2084 5349 2088 5353
rect 1928 5345 1932 5349
rect 1943 5345 1947 5349
rect 1959 5341 1963 5345
rect 1967 5341 1971 5345
rect 2018 5345 2022 5349
rect 2033 5345 2037 5349
rect 2049 5341 2053 5345
rect 2057 5341 2061 5345
rect 2099 5345 2103 5349
rect 2114 5345 2118 5349
rect 1763 5302 1767 5306
rect 1778 5302 1782 5306
rect 1049 5268 1053 5272
rect 1064 5268 1068 5272
rect 1154 5268 1158 5272
rect 1169 5268 1173 5272
rect 1209 5268 1213 5272
rect 1217 5268 1221 5272
rect 1227 5268 1231 5272
rect 1244 5268 1248 5272
rect 1252 5268 1256 5272
rect 1260 5268 1264 5272
rect 1273 5268 1277 5272
rect 1282 5268 1286 5272
rect 1299 5268 1303 5272
rect 1316 5268 1320 5272
rect 1327 5268 1331 5272
rect 1335 5268 1339 5272
rect 1343 5268 1347 5272
rect 1351 5268 1355 5272
rect 1359 5268 1363 5272
rect 1367 5268 1371 5272
rect 1543 5269 1559 5281
rect 1563 5269 1579 5281
rect 1596 5269 1612 5281
rect 1616 5269 1632 5281
rect 1994 5268 1998 5272
rect 2009 5268 2013 5272
rect 2099 5268 2103 5272
rect 2114 5268 2118 5272
rect 2154 5268 2158 5272
rect 2162 5268 2166 5272
rect 2172 5268 2176 5272
rect 2189 5268 2193 5272
rect 2197 5268 2201 5272
rect 2205 5268 2209 5272
rect 2218 5268 2222 5272
rect 2227 5268 2231 5272
rect 2244 5268 2248 5272
rect 2261 5268 2265 5272
rect 2272 5268 2276 5272
rect 2280 5268 2284 5272
rect 2288 5268 2292 5272
rect 2296 5268 2300 5272
rect 2304 5268 2308 5272
rect 2312 5268 2316 5272
rect 1026 5217 1030 5221
rect 1034 5217 1038 5221
rect 1209 5222 1213 5226
rect 1217 5222 1221 5226
rect 1227 5222 1231 5226
rect 1244 5222 1248 5226
rect 1252 5222 1256 5226
rect 1260 5222 1264 5226
rect 1273 5222 1277 5226
rect 1282 5222 1286 5226
rect 1299 5222 1303 5226
rect 1316 5222 1320 5226
rect 1327 5222 1331 5226
rect 1335 5222 1339 5226
rect 1343 5222 1347 5226
rect 1351 5222 1355 5226
rect 1359 5222 1363 5226
rect 1367 5222 1371 5226
rect 1131 5217 1135 5221
rect 1139 5217 1143 5221
rect 1049 5213 1053 5217
rect 1064 5213 1068 5217
rect 1080 5209 1084 5213
rect 1088 5209 1092 5213
rect 1154 5213 1158 5217
rect 1169 5213 1173 5217
rect 1740 5246 1744 5250
rect 1748 5246 1752 5250
rect 1763 5242 1767 5246
rect 1778 5242 1782 5246
rect 1794 5238 1798 5242
rect 1802 5238 1806 5242
rect 1971 5217 1975 5221
rect 1979 5217 1983 5221
rect 2154 5222 2158 5226
rect 2162 5222 2166 5226
rect 2172 5222 2176 5226
rect 2189 5222 2193 5226
rect 2197 5222 2201 5226
rect 2205 5222 2209 5226
rect 2218 5222 2222 5226
rect 2227 5222 2231 5226
rect 2244 5222 2248 5226
rect 2261 5222 2265 5226
rect 2272 5222 2276 5226
rect 2280 5222 2284 5226
rect 2288 5222 2292 5226
rect 2296 5222 2300 5226
rect 2304 5222 2308 5226
rect 2312 5222 2316 5226
rect 2076 5217 2080 5221
rect 2084 5217 2088 5221
rect 1994 5213 1998 5217
rect 2009 5213 2013 5217
rect 2025 5209 2029 5213
rect 2033 5209 2037 5213
rect 2099 5213 2103 5217
rect 2114 5213 2118 5217
rect 1073 5137 1077 5141
rect 1088 5137 1092 5141
rect 1154 5137 1158 5141
rect 1169 5137 1173 5141
rect 1609 5146 1613 5150
rect 1622 5146 1626 5150
rect 1630 5146 1634 5150
rect 1638 5146 1642 5150
rect 1646 5146 1650 5150
rect 1659 5146 1663 5150
rect 1672 5146 1676 5150
rect 1680 5146 1684 5150
rect 1688 5146 1692 5150
rect 1696 5146 1700 5150
rect 1704 5146 1708 5150
rect 1717 5146 1721 5150
rect 1725 5146 1729 5150
rect 1733 5146 1737 5150
rect 1209 5136 1213 5140
rect 1217 5136 1221 5140
rect 1227 5136 1231 5140
rect 1244 5136 1248 5140
rect 1252 5136 1256 5140
rect 1260 5136 1264 5140
rect 1273 5136 1277 5140
rect 1282 5136 1286 5140
rect 1299 5136 1303 5140
rect 1316 5136 1320 5140
rect 1327 5136 1331 5140
rect 1335 5136 1339 5140
rect 1343 5136 1347 5140
rect 1351 5136 1355 5140
rect 1359 5136 1363 5140
rect 1367 5136 1371 5140
rect 2018 5137 2022 5141
rect 2033 5137 2037 5141
rect 2099 5137 2103 5141
rect 2114 5137 2118 5141
rect 2554 5146 2558 5150
rect 2567 5146 2571 5150
rect 2575 5146 2579 5150
rect 2583 5146 2587 5150
rect 2591 5146 2595 5150
rect 2604 5146 2608 5150
rect 2617 5146 2621 5150
rect 2625 5146 2629 5150
rect 2633 5146 2637 5150
rect 2641 5146 2645 5150
rect 2649 5146 2653 5150
rect 2662 5146 2666 5150
rect 2670 5146 2674 5150
rect 2678 5146 2682 5150
rect 2154 5136 2158 5140
rect 2162 5136 2166 5140
rect 2172 5136 2176 5140
rect 2189 5136 2193 5140
rect 2197 5136 2201 5140
rect 2205 5136 2209 5140
rect 2218 5136 2222 5140
rect 2227 5136 2231 5140
rect 2244 5136 2248 5140
rect 2261 5136 2265 5140
rect 2272 5136 2276 5140
rect 2280 5136 2284 5140
rect 2288 5136 2292 5140
rect 2296 5136 2300 5140
rect 2304 5136 2308 5140
rect 2312 5136 2316 5140
rect 1050 5085 1054 5089
rect 1058 5085 1062 5089
rect 1209 5090 1213 5094
rect 1217 5090 1221 5094
rect 1227 5090 1231 5094
rect 1244 5090 1248 5094
rect 1252 5090 1256 5094
rect 1260 5090 1264 5094
rect 1273 5090 1277 5094
rect 1282 5090 1286 5094
rect 1299 5090 1303 5094
rect 1316 5090 1320 5094
rect 1327 5090 1331 5094
rect 1335 5090 1339 5094
rect 1343 5090 1347 5094
rect 1351 5090 1355 5094
rect 1359 5090 1363 5094
rect 1367 5090 1371 5094
rect 1709 5090 1713 5094
rect 1717 5090 1721 5094
rect 1131 5085 1135 5089
rect 1139 5085 1143 5089
rect 1073 5081 1077 5085
rect 1088 5081 1092 5085
rect 1104 5077 1108 5081
rect 1112 5077 1116 5081
rect 1154 5081 1158 5085
rect 1169 5081 1173 5085
rect 1185 5077 1189 5081
rect 1193 5077 1197 5081
rect 1592 5081 1596 5085
rect 1600 5081 1604 5085
rect 1995 5085 1999 5089
rect 2003 5085 2007 5089
rect 2154 5090 2158 5094
rect 2162 5090 2166 5094
rect 2172 5090 2176 5094
rect 2189 5090 2193 5094
rect 2197 5090 2201 5094
rect 2205 5090 2209 5094
rect 2218 5090 2222 5094
rect 2227 5090 2231 5094
rect 2244 5090 2248 5094
rect 2261 5090 2265 5094
rect 2272 5090 2276 5094
rect 2280 5090 2284 5094
rect 2288 5090 2292 5094
rect 2296 5090 2300 5094
rect 2304 5090 2308 5094
rect 2312 5090 2316 5094
rect 2654 5090 2658 5094
rect 2662 5090 2666 5094
rect 2076 5085 2080 5089
rect 2084 5085 2088 5089
rect 2018 5081 2022 5085
rect 2033 5081 2037 5085
rect 2049 5077 2053 5081
rect 2057 5077 2061 5081
rect 2099 5081 2103 5085
rect 2114 5081 2118 5085
rect 2130 5077 2134 5081
rect 2138 5077 2142 5081
rect 2537 5081 2541 5085
rect 2545 5081 2549 5085
rect 1600 5044 1604 5048
rect 1608 5044 1612 5048
rect 1616 5044 1620 5048
rect 1629 5044 1633 5048
rect 1637 5044 1641 5048
rect 1645 5044 1649 5048
rect 1653 5044 1657 5048
rect 1661 5044 1665 5048
rect 1674 5044 1678 5048
rect 1687 5044 1691 5048
rect 1695 5044 1699 5048
rect 1703 5044 1707 5048
rect 1711 5044 1715 5048
rect 1724 5044 1728 5048
rect 2545 5044 2549 5048
rect 2553 5044 2557 5048
rect 2561 5044 2565 5048
rect 2574 5044 2578 5048
rect 2582 5044 2586 5048
rect 2590 5044 2594 5048
rect 2598 5044 2602 5048
rect 2606 5044 2610 5048
rect 2619 5044 2623 5048
rect 2632 5044 2636 5048
rect 2640 5044 2644 5048
rect 2648 5044 2652 5048
rect 2656 5044 2660 5048
rect 2669 5044 2673 5048
rect 852 5011 856 5015
rect 860 5011 864 5015
rect 868 5011 872 5015
rect 881 5011 885 5015
rect 889 5011 893 5015
rect 897 5011 901 5015
rect 905 5011 909 5015
rect 913 5011 917 5015
rect 926 5011 930 5015
rect 939 5011 943 5015
rect 947 5011 951 5015
rect 955 5011 959 5015
rect 963 5011 967 5015
rect 976 5011 980 5015
rect 984 5011 988 5015
rect 992 5011 996 5015
rect 1000 5011 1004 5015
rect 1013 5011 1017 5015
rect 1021 5011 1025 5015
rect 1029 5011 1033 5015
rect 1037 5011 1041 5015
rect 1045 5011 1049 5015
rect 1058 5011 1062 5015
rect 1071 5011 1075 5015
rect 1079 5011 1083 5015
rect 1087 5011 1091 5015
rect 1095 5011 1099 5015
rect 1108 5011 1112 5015
rect 1116 5011 1120 5015
rect 1124 5011 1128 5015
rect 1132 5011 1136 5015
rect 1145 5011 1149 5015
rect 1153 5011 1157 5015
rect 1161 5011 1165 5015
rect 1169 5011 1173 5015
rect 1177 5011 1181 5015
rect 1190 5011 1194 5015
rect 1203 5011 1207 5015
rect 1211 5011 1215 5015
rect 1219 5011 1223 5015
rect 1227 5011 1231 5015
rect 1240 5011 1244 5015
rect 1248 5011 1252 5015
rect 1256 5011 1260 5015
rect 1264 5011 1268 5015
rect 1277 5011 1281 5015
rect 1285 5011 1289 5015
rect 1293 5011 1297 5015
rect 1301 5011 1305 5015
rect 1309 5011 1313 5015
rect 1322 5011 1326 5015
rect 1335 5011 1339 5015
rect 1343 5011 1347 5015
rect 1351 5011 1355 5015
rect 1359 5011 1363 5015
rect 1372 5011 1376 5015
rect 1797 5011 1801 5015
rect 1805 5011 1809 5015
rect 1813 5011 1817 5015
rect 1826 5011 1830 5015
rect 1834 5011 1838 5015
rect 1842 5011 1846 5015
rect 1850 5011 1854 5015
rect 1858 5011 1862 5015
rect 1871 5011 1875 5015
rect 1884 5011 1888 5015
rect 1892 5011 1896 5015
rect 1900 5011 1904 5015
rect 1908 5011 1912 5015
rect 1921 5011 1925 5015
rect 1929 5011 1933 5015
rect 1937 5011 1941 5015
rect 1945 5011 1949 5015
rect 1958 5011 1962 5015
rect 1966 5011 1970 5015
rect 1974 5011 1978 5015
rect 1982 5011 1986 5015
rect 1990 5011 1994 5015
rect 2003 5011 2007 5015
rect 2016 5011 2020 5015
rect 2024 5011 2028 5015
rect 2032 5011 2036 5015
rect 2040 5011 2044 5015
rect 2053 5011 2057 5015
rect 2061 5011 2065 5015
rect 2069 5011 2073 5015
rect 2077 5011 2081 5015
rect 2090 5011 2094 5015
rect 2098 5011 2102 5015
rect 2106 5011 2110 5015
rect 2114 5011 2118 5015
rect 2122 5011 2126 5015
rect 2135 5011 2139 5015
rect 2148 5011 2152 5015
rect 2156 5011 2160 5015
rect 2164 5011 2168 5015
rect 2172 5011 2176 5015
rect 2185 5011 2189 5015
rect 2193 5011 2197 5015
rect 2201 5011 2205 5015
rect 2209 5011 2213 5015
rect 2222 5011 2226 5015
rect 2230 5011 2234 5015
rect 2238 5011 2242 5015
rect 2246 5011 2250 5015
rect 2254 5011 2258 5015
rect 2267 5011 2271 5015
rect 2280 5011 2284 5015
rect 2288 5011 2292 5015
rect 2296 5011 2300 5015
rect 2304 5011 2308 5015
rect 2317 5011 2321 5015
rect 4574 7986 4578 8015
rect 4574 7975 4578 7982
rect 4582 7975 4586 8015
rect 4590 7986 4594 8015
rect 4590 7975 4594 7982
rect 4598 7975 4602 8015
rect 4606 7986 4610 8015
rect 4606 7975 4610 7982
rect 4614 7975 4618 8015
rect 4622 7986 4626 8015
rect 4622 7975 4626 7982
rect 4637 7975 4641 8034
rect 4645 7986 4649 8034
rect 4645 7975 4649 7982
rect 4653 7975 4657 8034
rect 4661 7986 4665 8034
rect 4661 7975 4665 7982
rect 4680 7975 4684 8034
rect 4688 7986 4692 8034
rect 4696 7975 4700 8034
rect 4704 7986 4708 8034
rect 4704 7975 4708 7982
rect 4721 7975 4725 8034
rect 4729 7986 4733 8034
rect 4737 7975 4741 8034
rect 4745 7986 4749 8034
rect 4745 7975 4749 7982
rect 4657 7461 4661 7465
rect 4667 7461 4671 7465
rect 4677 7461 4681 7465
rect 4687 7461 4691 7465
rect 4697 7461 4701 7465
rect 4707 7461 4711 7465
rect 4717 7461 4721 7465
rect 4727 7461 4731 7465
rect 4737 7461 4741 7465
rect 4662 7456 4666 7460
rect 4672 7456 4676 7460
rect 4682 7456 4686 7460
rect 4692 7456 4696 7460
rect 4702 7456 4706 7460
rect 4712 7456 4716 7460
rect 4722 7456 4726 7460
rect 4732 7456 4736 7460
rect 4742 7456 4746 7460
rect 4657 7451 4661 7455
rect 4667 7451 4671 7455
rect 4677 7451 4681 7455
rect 4687 7451 4691 7455
rect 4697 7451 4701 7455
rect 4707 7451 4711 7455
rect 4717 7451 4721 7455
rect 4727 7451 4731 7455
rect 4737 7451 4741 7455
rect 4662 7446 4666 7450
rect 4672 7446 4676 7450
rect 4682 7446 4686 7450
rect 4692 7446 4696 7450
rect 4702 7446 4706 7450
rect 4712 7446 4716 7450
rect 4722 7446 4726 7450
rect 4732 7446 4736 7450
rect 4742 7446 4746 7450
rect 4657 7441 4661 7445
rect 4667 7441 4671 7445
rect 4677 7441 4681 7445
rect 4687 7441 4691 7445
rect 4697 7441 4701 7445
rect 4707 7441 4711 7445
rect 4717 7441 4721 7445
rect 4727 7441 4731 7445
rect 4737 7441 4741 7445
rect 4662 7436 4666 7440
rect 4672 7436 4676 7440
rect 4682 7436 4686 7440
rect 4692 7436 4696 7440
rect 4702 7436 4706 7440
rect 4712 7436 4716 7440
rect 4722 7436 4726 7440
rect 4732 7436 4736 7440
rect 4742 7436 4746 7440
rect 4657 7431 4661 7435
rect 4667 7431 4671 7435
rect 4677 7431 4681 7435
rect 4687 7431 4691 7435
rect 4697 7431 4701 7435
rect 4707 7431 4711 7435
rect 4717 7431 4721 7435
rect 4727 7431 4731 7435
rect 4737 7431 4741 7435
rect 4662 7426 4666 7430
rect 4672 7426 4676 7430
rect 4682 7426 4686 7430
rect 4692 7426 4696 7430
rect 4702 7426 4706 7430
rect 4712 7426 4716 7430
rect 4722 7426 4726 7430
rect 4732 7426 4736 7430
rect 4742 7426 4746 7430
rect 4657 7421 4661 7425
rect 4667 7421 4671 7425
rect 4677 7421 4681 7425
rect 4687 7421 4691 7425
rect 4697 7421 4701 7425
rect 4707 7421 4711 7425
rect 4717 7421 4721 7425
rect 4727 7421 4731 7425
rect 4737 7421 4741 7425
rect 4572 7335 4576 7342
rect 4572 7302 4576 7331
rect 4580 7302 4584 7342
rect 4588 7335 4592 7342
rect 4588 7302 4592 7331
rect 4596 7302 4600 7342
rect 4604 7335 4608 7342
rect 4604 7302 4608 7331
rect 4612 7302 4616 7342
rect 4620 7335 4624 7342
rect 4620 7302 4624 7331
rect 1140 4531 1169 4535
rect 1173 4531 1180 4535
rect 2067 4531 2096 4535
rect 2100 4531 2107 4535
rect 2376 4531 2405 4535
rect 2409 4531 2416 4535
rect 2685 4531 2714 4535
rect 2718 4531 2725 4535
rect 2994 4531 3023 4535
rect 3027 4531 3034 4535
rect 3303 4531 3332 4535
rect 3336 4531 3343 4535
rect 1140 4523 1180 4527
rect 1140 4515 1169 4519
rect 1173 4515 1180 4519
rect 1140 4507 1180 4511
rect 1140 4499 1169 4503
rect 1173 4499 1180 4503
rect 2067 4523 2107 4527
rect 2067 4515 2096 4519
rect 2100 4515 2107 4519
rect 2067 4507 2107 4511
rect 2067 4499 2096 4503
rect 2100 4499 2107 4503
rect 2376 4523 2416 4527
rect 2376 4515 2405 4519
rect 2409 4515 2416 4519
rect 2376 4507 2416 4511
rect 2376 4499 2405 4503
rect 2409 4499 2416 4503
rect 2685 4523 2725 4527
rect 2685 4515 2714 4519
rect 2718 4515 2725 4519
rect 2685 4507 2725 4511
rect 2685 4499 2714 4503
rect 2718 4499 2725 4503
rect 2994 4523 3034 4527
rect 2994 4515 3023 4519
rect 3027 4515 3034 4519
rect 2994 4507 3034 4511
rect 2994 4499 3023 4503
rect 3027 4499 3034 4503
rect 3303 4523 3343 4527
rect 3303 4515 3332 4519
rect 3336 4515 3343 4519
rect 3303 4507 3343 4511
rect 3303 4499 3332 4503
rect 3336 4499 3343 4503
rect 1140 4491 1180 4495
rect 2067 4491 2107 4495
rect 2376 4491 2416 4495
rect 2685 4491 2725 4495
rect 2994 4491 3034 4495
rect 3303 4491 3343 4495
rect 1140 4483 1169 4487
rect 1173 4483 1180 4487
rect 2067 4483 2096 4487
rect 2100 4483 2107 4487
rect 2376 4483 2405 4487
rect 2409 4483 2416 4487
rect 2685 4483 2714 4487
rect 2718 4483 2725 4487
rect 2994 4483 3023 4487
rect 3027 4483 3034 4487
rect 3303 4483 3332 4487
rect 3336 4483 3343 4487
rect 1259 4446 1263 4450
rect 1269 4446 1273 4450
rect 1279 4446 1283 4450
rect 1289 4446 1293 4450
rect 1299 4446 1303 4450
rect 1264 4441 1268 4445
rect 1274 4441 1278 4445
rect 1284 4441 1288 4445
rect 1294 4441 1298 4445
rect 1259 4436 1263 4440
rect 1269 4436 1273 4440
rect 1279 4436 1283 4440
rect 1289 4436 1293 4440
rect 1299 4436 1303 4440
rect 1264 4431 1268 4435
rect 1274 4431 1278 4435
rect 1284 4431 1288 4435
rect 1294 4431 1298 4435
rect 1259 4426 1263 4430
rect 1269 4426 1273 4430
rect 1279 4426 1283 4430
rect 1289 4426 1293 4430
rect 1299 4426 1303 4430
rect 1264 4421 1268 4425
rect 1274 4421 1278 4425
rect 1284 4421 1288 4425
rect 1294 4421 1298 4425
rect 1259 4416 1263 4420
rect 1269 4416 1273 4420
rect 1279 4416 1283 4420
rect 1289 4416 1293 4420
rect 1299 4416 1303 4420
rect 1264 4411 1268 4415
rect 1274 4411 1278 4415
rect 1284 4411 1288 4415
rect 1294 4411 1298 4415
rect 1259 4406 1263 4410
rect 1269 4406 1273 4410
rect 1279 4406 1283 4410
rect 1289 4406 1293 4410
rect 1299 4406 1303 4410
rect 1264 4401 1268 4405
rect 1274 4401 1278 4405
rect 1284 4401 1288 4405
rect 1294 4401 1298 4405
rect 1259 4396 1263 4400
rect 1269 4396 1273 4400
rect 1279 4396 1283 4400
rect 1289 4396 1293 4400
rect 1299 4396 1303 4400
rect 1264 4391 1268 4395
rect 1274 4391 1278 4395
rect 1284 4391 1288 4395
rect 1294 4391 1298 4395
rect 1259 4386 1263 4390
rect 1269 4386 1273 4390
rect 1279 4386 1283 4390
rect 1289 4386 1293 4390
rect 1299 4386 1303 4390
rect 1264 4381 1268 4385
rect 1274 4381 1278 4385
rect 1284 4381 1288 4385
rect 1294 4381 1298 4385
rect 1259 4376 1263 4380
rect 1269 4376 1273 4380
rect 1279 4376 1283 4380
rect 1289 4376 1293 4380
rect 1299 4376 1303 4380
rect 1264 4371 1268 4375
rect 1274 4371 1278 4375
rect 1284 4371 1288 4375
rect 1294 4371 1298 4375
rect 1259 4366 1263 4370
rect 1269 4366 1273 4370
rect 1279 4366 1283 4370
rect 1289 4366 1293 4370
rect 1299 4366 1303 4370
rect 1264 4361 1268 4365
rect 1274 4361 1278 4365
rect 1284 4361 1288 4365
rect 1294 4361 1298 4365
rect 1568 4446 1572 4450
rect 1578 4446 1582 4450
rect 1588 4446 1592 4450
rect 1598 4446 1602 4450
rect 1608 4446 1612 4450
rect 1573 4441 1577 4445
rect 1583 4441 1587 4445
rect 1593 4441 1597 4445
rect 1603 4441 1607 4445
rect 1568 4436 1572 4440
rect 1578 4436 1582 4440
rect 1588 4436 1592 4440
rect 1598 4436 1602 4440
rect 1608 4436 1612 4440
rect 1573 4431 1577 4435
rect 1583 4431 1587 4435
rect 1593 4431 1597 4435
rect 1603 4431 1607 4435
rect 1568 4426 1572 4430
rect 1578 4426 1582 4430
rect 1588 4426 1592 4430
rect 1598 4426 1602 4430
rect 1608 4426 1612 4430
rect 1573 4421 1577 4425
rect 1583 4421 1587 4425
rect 1593 4421 1597 4425
rect 1603 4421 1607 4425
rect 1568 4416 1572 4420
rect 1578 4416 1582 4420
rect 1588 4416 1592 4420
rect 1598 4416 1602 4420
rect 1608 4416 1612 4420
rect 1573 4411 1577 4415
rect 1583 4411 1587 4415
rect 1593 4411 1597 4415
rect 1603 4411 1607 4415
rect 1568 4406 1572 4410
rect 1578 4406 1582 4410
rect 1588 4406 1592 4410
rect 1598 4406 1602 4410
rect 1608 4406 1612 4410
rect 1573 4401 1577 4405
rect 1583 4401 1587 4405
rect 1593 4401 1597 4405
rect 1603 4401 1607 4405
rect 1568 4396 1572 4400
rect 1578 4396 1582 4400
rect 1588 4396 1592 4400
rect 1598 4396 1602 4400
rect 1608 4396 1612 4400
rect 1573 4391 1577 4395
rect 1583 4391 1587 4395
rect 1593 4391 1597 4395
rect 1603 4391 1607 4395
rect 1568 4386 1572 4390
rect 1578 4386 1582 4390
rect 1588 4386 1592 4390
rect 1598 4386 1602 4390
rect 1608 4386 1612 4390
rect 1573 4381 1577 4385
rect 1583 4381 1587 4385
rect 1593 4381 1597 4385
rect 1603 4381 1607 4385
rect 1568 4376 1572 4380
rect 1578 4376 1582 4380
rect 1588 4376 1592 4380
rect 1598 4376 1602 4380
rect 1608 4376 1612 4380
rect 1573 4371 1577 4375
rect 1583 4371 1587 4375
rect 1593 4371 1597 4375
rect 1603 4371 1607 4375
rect 1568 4366 1572 4370
rect 1578 4366 1582 4370
rect 1588 4366 1592 4370
rect 1598 4366 1602 4370
rect 1608 4366 1612 4370
rect 1573 4361 1577 4365
rect 1583 4361 1587 4365
rect 1593 4361 1597 4365
rect 1603 4361 1607 4365
rect 1877 4446 1881 4450
rect 1887 4446 1891 4450
rect 1897 4446 1901 4450
rect 1907 4446 1911 4450
rect 1917 4446 1921 4450
rect 1882 4441 1886 4445
rect 1892 4441 1896 4445
rect 1902 4441 1906 4445
rect 1912 4441 1916 4445
rect 1877 4436 1881 4440
rect 1887 4436 1891 4440
rect 1897 4436 1901 4440
rect 1907 4436 1911 4440
rect 1917 4436 1921 4440
rect 1882 4431 1886 4435
rect 1892 4431 1896 4435
rect 1902 4431 1906 4435
rect 1912 4431 1916 4435
rect 1877 4426 1881 4430
rect 1887 4426 1891 4430
rect 1897 4426 1901 4430
rect 1907 4426 1911 4430
rect 1917 4426 1921 4430
rect 1882 4421 1886 4425
rect 1892 4421 1896 4425
rect 1902 4421 1906 4425
rect 1912 4421 1916 4425
rect 1877 4416 1881 4420
rect 1887 4416 1891 4420
rect 1897 4416 1901 4420
rect 1907 4416 1911 4420
rect 1917 4416 1921 4420
rect 1882 4411 1886 4415
rect 1892 4411 1896 4415
rect 1902 4411 1906 4415
rect 1912 4411 1916 4415
rect 1877 4406 1881 4410
rect 1887 4406 1891 4410
rect 1897 4406 1901 4410
rect 1907 4406 1911 4410
rect 1917 4406 1921 4410
rect 1882 4401 1886 4405
rect 1892 4401 1896 4405
rect 1902 4401 1906 4405
rect 1912 4401 1916 4405
rect 1877 4396 1881 4400
rect 1887 4396 1891 4400
rect 1897 4396 1901 4400
rect 1907 4396 1911 4400
rect 1917 4396 1921 4400
rect 1882 4391 1886 4395
rect 1892 4391 1896 4395
rect 1902 4391 1906 4395
rect 1912 4391 1916 4395
rect 1877 4386 1881 4390
rect 1887 4386 1891 4390
rect 1897 4386 1901 4390
rect 1907 4386 1911 4390
rect 1917 4386 1921 4390
rect 1882 4381 1886 4385
rect 1892 4381 1896 4385
rect 1902 4381 1906 4385
rect 1912 4381 1916 4385
rect 1877 4376 1881 4380
rect 1887 4376 1891 4380
rect 1897 4376 1901 4380
rect 1907 4376 1911 4380
rect 1917 4376 1921 4380
rect 1882 4371 1886 4375
rect 1892 4371 1896 4375
rect 1902 4371 1906 4375
rect 1912 4371 1916 4375
rect 1877 4366 1881 4370
rect 1887 4366 1891 4370
rect 1897 4366 1901 4370
rect 1907 4366 1911 4370
rect 1917 4366 1921 4370
rect 1882 4361 1886 4365
rect 1892 4361 1896 4365
rect 1902 4361 1906 4365
rect 1912 4361 1916 4365
rect 2186 4446 2190 4450
rect 2196 4446 2200 4450
rect 2206 4446 2210 4450
rect 2216 4446 2220 4450
rect 2226 4446 2230 4450
rect 2191 4441 2195 4445
rect 2201 4441 2205 4445
rect 2211 4441 2215 4445
rect 2221 4441 2225 4445
rect 2186 4436 2190 4440
rect 2196 4436 2200 4440
rect 2206 4436 2210 4440
rect 2216 4436 2220 4440
rect 2226 4436 2230 4440
rect 2191 4431 2195 4435
rect 2201 4431 2205 4435
rect 2211 4431 2215 4435
rect 2221 4431 2225 4435
rect 2186 4426 2190 4430
rect 2196 4426 2200 4430
rect 2206 4426 2210 4430
rect 2216 4426 2220 4430
rect 2226 4426 2230 4430
rect 2191 4421 2195 4425
rect 2201 4421 2205 4425
rect 2211 4421 2215 4425
rect 2221 4421 2225 4425
rect 2186 4416 2190 4420
rect 2196 4416 2200 4420
rect 2206 4416 2210 4420
rect 2216 4416 2220 4420
rect 2226 4416 2230 4420
rect 2191 4411 2195 4415
rect 2201 4411 2205 4415
rect 2211 4411 2215 4415
rect 2221 4411 2225 4415
rect 2186 4406 2190 4410
rect 2196 4406 2200 4410
rect 2206 4406 2210 4410
rect 2216 4406 2220 4410
rect 2226 4406 2230 4410
rect 2191 4401 2195 4405
rect 2201 4401 2205 4405
rect 2211 4401 2215 4405
rect 2221 4401 2225 4405
rect 2186 4396 2190 4400
rect 2196 4396 2200 4400
rect 2206 4396 2210 4400
rect 2216 4396 2220 4400
rect 2226 4396 2230 4400
rect 2191 4391 2195 4395
rect 2201 4391 2205 4395
rect 2211 4391 2215 4395
rect 2221 4391 2225 4395
rect 2186 4386 2190 4390
rect 2196 4386 2200 4390
rect 2206 4386 2210 4390
rect 2216 4386 2220 4390
rect 2226 4386 2230 4390
rect 2191 4381 2195 4385
rect 2201 4381 2205 4385
rect 2211 4381 2215 4385
rect 2221 4381 2225 4385
rect 2186 4376 2190 4380
rect 2196 4376 2200 4380
rect 2206 4376 2210 4380
rect 2216 4376 2220 4380
rect 2226 4376 2230 4380
rect 2191 4371 2195 4375
rect 2201 4371 2205 4375
rect 2211 4371 2215 4375
rect 2221 4371 2225 4375
rect 2186 4366 2190 4370
rect 2196 4366 2200 4370
rect 2206 4366 2210 4370
rect 2216 4366 2220 4370
rect 2226 4366 2230 4370
rect 2191 4361 2195 4365
rect 2201 4361 2205 4365
rect 2211 4361 2215 4365
rect 2221 4361 2225 4365
rect 2495 4446 2499 4450
rect 2505 4446 2509 4450
rect 2515 4446 2519 4450
rect 2525 4446 2529 4450
rect 2535 4446 2539 4450
rect 2500 4441 2504 4445
rect 2510 4441 2514 4445
rect 2520 4441 2524 4445
rect 2530 4441 2534 4445
rect 2495 4436 2499 4440
rect 2505 4436 2509 4440
rect 2515 4436 2519 4440
rect 2525 4436 2529 4440
rect 2535 4436 2539 4440
rect 2500 4431 2504 4435
rect 2510 4431 2514 4435
rect 2520 4431 2524 4435
rect 2530 4431 2534 4435
rect 2495 4426 2499 4430
rect 2505 4426 2509 4430
rect 2515 4426 2519 4430
rect 2525 4426 2529 4430
rect 2535 4426 2539 4430
rect 2500 4421 2504 4425
rect 2510 4421 2514 4425
rect 2520 4421 2524 4425
rect 2530 4421 2534 4425
rect 2495 4416 2499 4420
rect 2505 4416 2509 4420
rect 2515 4416 2519 4420
rect 2525 4416 2529 4420
rect 2535 4416 2539 4420
rect 2500 4411 2504 4415
rect 2510 4411 2514 4415
rect 2520 4411 2524 4415
rect 2530 4411 2534 4415
rect 2495 4406 2499 4410
rect 2505 4406 2509 4410
rect 2515 4406 2519 4410
rect 2525 4406 2529 4410
rect 2535 4406 2539 4410
rect 2500 4401 2504 4405
rect 2510 4401 2514 4405
rect 2520 4401 2524 4405
rect 2530 4401 2534 4405
rect 2495 4396 2499 4400
rect 2505 4396 2509 4400
rect 2515 4396 2519 4400
rect 2525 4396 2529 4400
rect 2535 4396 2539 4400
rect 2500 4391 2504 4395
rect 2510 4391 2514 4395
rect 2520 4391 2524 4395
rect 2530 4391 2534 4395
rect 2495 4386 2499 4390
rect 2505 4386 2509 4390
rect 2515 4386 2519 4390
rect 2525 4386 2529 4390
rect 2535 4386 2539 4390
rect 2500 4381 2504 4385
rect 2510 4381 2514 4385
rect 2520 4381 2524 4385
rect 2530 4381 2534 4385
rect 2495 4376 2499 4380
rect 2505 4376 2509 4380
rect 2515 4376 2519 4380
rect 2525 4376 2529 4380
rect 2535 4376 2539 4380
rect 2500 4371 2504 4375
rect 2510 4371 2514 4375
rect 2520 4371 2524 4375
rect 2530 4371 2534 4375
rect 2495 4366 2499 4370
rect 2505 4366 2509 4370
rect 2515 4366 2519 4370
rect 2525 4366 2529 4370
rect 2535 4366 2539 4370
rect 2500 4361 2504 4365
rect 2510 4361 2514 4365
rect 2520 4361 2524 4365
rect 2530 4361 2534 4365
rect 2804 4446 2808 4450
rect 2814 4446 2818 4450
rect 2824 4446 2828 4450
rect 2834 4446 2838 4450
rect 2844 4446 2848 4450
rect 2809 4441 2813 4445
rect 2819 4441 2823 4445
rect 2829 4441 2833 4445
rect 2839 4441 2843 4445
rect 2804 4436 2808 4440
rect 2814 4436 2818 4440
rect 2824 4436 2828 4440
rect 2834 4436 2838 4440
rect 2844 4436 2848 4440
rect 2809 4431 2813 4435
rect 2819 4431 2823 4435
rect 2829 4431 2833 4435
rect 2839 4431 2843 4435
rect 2804 4426 2808 4430
rect 2814 4426 2818 4430
rect 2824 4426 2828 4430
rect 2834 4426 2838 4430
rect 2844 4426 2848 4430
rect 2809 4421 2813 4425
rect 2819 4421 2823 4425
rect 2829 4421 2833 4425
rect 2839 4421 2843 4425
rect 2804 4416 2808 4420
rect 2814 4416 2818 4420
rect 2824 4416 2828 4420
rect 2834 4416 2838 4420
rect 2844 4416 2848 4420
rect 2809 4411 2813 4415
rect 2819 4411 2823 4415
rect 2829 4411 2833 4415
rect 2839 4411 2843 4415
rect 2804 4406 2808 4410
rect 2814 4406 2818 4410
rect 2824 4406 2828 4410
rect 2834 4406 2838 4410
rect 2844 4406 2848 4410
rect 2809 4401 2813 4405
rect 2819 4401 2823 4405
rect 2829 4401 2833 4405
rect 2839 4401 2843 4405
rect 2804 4396 2808 4400
rect 2814 4396 2818 4400
rect 2824 4396 2828 4400
rect 2834 4396 2838 4400
rect 2844 4396 2848 4400
rect 2809 4391 2813 4395
rect 2819 4391 2823 4395
rect 2829 4391 2833 4395
rect 2839 4391 2843 4395
rect 2804 4386 2808 4390
rect 2814 4386 2818 4390
rect 2824 4386 2828 4390
rect 2834 4386 2838 4390
rect 2844 4386 2848 4390
rect 2809 4381 2813 4385
rect 2819 4381 2823 4385
rect 2829 4381 2833 4385
rect 2839 4381 2843 4385
rect 2804 4376 2808 4380
rect 2814 4376 2818 4380
rect 2824 4376 2828 4380
rect 2834 4376 2838 4380
rect 2844 4376 2848 4380
rect 2809 4371 2813 4375
rect 2819 4371 2823 4375
rect 2829 4371 2833 4375
rect 2839 4371 2843 4375
rect 2804 4366 2808 4370
rect 2814 4366 2818 4370
rect 2824 4366 2828 4370
rect 2834 4366 2838 4370
rect 2844 4366 2848 4370
rect 2809 4361 2813 4365
rect 2819 4361 2823 4365
rect 2829 4361 2833 4365
rect 2839 4361 2843 4365
rect 3113 4446 3117 4450
rect 3123 4446 3127 4450
rect 3133 4446 3137 4450
rect 3143 4446 3147 4450
rect 3153 4446 3157 4450
rect 3118 4441 3122 4445
rect 3128 4441 3132 4445
rect 3138 4441 3142 4445
rect 3148 4441 3152 4445
rect 3113 4436 3117 4440
rect 3123 4436 3127 4440
rect 3133 4436 3137 4440
rect 3143 4436 3147 4440
rect 3153 4436 3157 4440
rect 3118 4431 3122 4435
rect 3128 4431 3132 4435
rect 3138 4431 3142 4435
rect 3148 4431 3152 4435
rect 3113 4426 3117 4430
rect 3123 4426 3127 4430
rect 3133 4426 3137 4430
rect 3143 4426 3147 4430
rect 3153 4426 3157 4430
rect 3118 4421 3122 4425
rect 3128 4421 3132 4425
rect 3138 4421 3142 4425
rect 3148 4421 3152 4425
rect 3113 4416 3117 4420
rect 3123 4416 3127 4420
rect 3133 4416 3137 4420
rect 3143 4416 3147 4420
rect 3153 4416 3157 4420
rect 3118 4411 3122 4415
rect 3128 4411 3132 4415
rect 3138 4411 3142 4415
rect 3148 4411 3152 4415
rect 3113 4406 3117 4410
rect 3123 4406 3127 4410
rect 3133 4406 3137 4410
rect 3143 4406 3147 4410
rect 3153 4406 3157 4410
rect 3118 4401 3122 4405
rect 3128 4401 3132 4405
rect 3138 4401 3142 4405
rect 3148 4401 3152 4405
rect 3113 4396 3117 4400
rect 3123 4396 3127 4400
rect 3133 4396 3137 4400
rect 3143 4396 3147 4400
rect 3153 4396 3157 4400
rect 3118 4391 3122 4395
rect 3128 4391 3132 4395
rect 3138 4391 3142 4395
rect 3148 4391 3152 4395
rect 3113 4386 3117 4390
rect 3123 4386 3127 4390
rect 3133 4386 3137 4390
rect 3143 4386 3147 4390
rect 3153 4386 3157 4390
rect 3118 4381 3122 4385
rect 3128 4381 3132 4385
rect 3138 4381 3142 4385
rect 3148 4381 3152 4385
rect 3113 4376 3117 4380
rect 3123 4376 3127 4380
rect 3133 4376 3137 4380
rect 3143 4376 3147 4380
rect 3153 4376 3157 4380
rect 3118 4371 3122 4375
rect 3128 4371 3132 4375
rect 3138 4371 3142 4375
rect 3148 4371 3152 4375
rect 3113 4366 3117 4370
rect 3123 4366 3127 4370
rect 3133 4366 3137 4370
rect 3143 4366 3147 4370
rect 3153 4366 3157 4370
rect 3118 4361 3122 4365
rect 3128 4361 3132 4365
rect 3138 4361 3142 4365
rect 3148 4361 3152 4365
rect 3422 4446 3426 4450
rect 3432 4446 3436 4450
rect 3442 4446 3446 4450
rect 3452 4446 3456 4450
rect 3462 4446 3466 4450
rect 3427 4441 3431 4445
rect 3437 4441 3441 4445
rect 3447 4441 3451 4445
rect 3457 4441 3461 4445
rect 3422 4436 3426 4440
rect 3432 4436 3436 4440
rect 3442 4436 3446 4440
rect 3452 4436 3456 4440
rect 3462 4436 3466 4440
rect 3427 4431 3431 4435
rect 3437 4431 3441 4435
rect 3447 4431 3451 4435
rect 3457 4431 3461 4435
rect 3422 4426 3426 4430
rect 3432 4426 3436 4430
rect 3442 4426 3446 4430
rect 3452 4426 3456 4430
rect 3462 4426 3466 4430
rect 3427 4421 3431 4425
rect 3437 4421 3441 4425
rect 3447 4421 3451 4425
rect 3457 4421 3461 4425
rect 3422 4416 3426 4420
rect 3432 4416 3436 4420
rect 3442 4416 3446 4420
rect 3452 4416 3456 4420
rect 3462 4416 3466 4420
rect 3427 4411 3431 4415
rect 3437 4411 3441 4415
rect 3447 4411 3451 4415
rect 3457 4411 3461 4415
rect 3422 4406 3426 4410
rect 3432 4406 3436 4410
rect 3442 4406 3446 4410
rect 3452 4406 3456 4410
rect 3462 4406 3466 4410
rect 3427 4401 3431 4405
rect 3437 4401 3441 4405
rect 3447 4401 3451 4405
rect 3457 4401 3461 4405
rect 3422 4396 3426 4400
rect 3432 4396 3436 4400
rect 3442 4396 3446 4400
rect 3452 4396 3456 4400
rect 3462 4396 3466 4400
rect 3427 4391 3431 4395
rect 3437 4391 3441 4395
rect 3447 4391 3451 4395
rect 3457 4391 3461 4395
rect 3422 4386 3426 4390
rect 3432 4386 3436 4390
rect 3442 4386 3446 4390
rect 3452 4386 3456 4390
rect 3462 4386 3466 4390
rect 3427 4381 3431 4385
rect 3437 4381 3441 4385
rect 3447 4381 3451 4385
rect 3457 4381 3461 4385
rect 3422 4376 3426 4380
rect 3432 4376 3436 4380
rect 3442 4376 3446 4380
rect 3452 4376 3456 4380
rect 3462 4376 3466 4380
rect 3427 4371 3431 4375
rect 3437 4371 3441 4375
rect 3447 4371 3451 4375
rect 3457 4371 3461 4375
rect 3422 4366 3426 4370
rect 3432 4366 3436 4370
rect 3442 4366 3446 4370
rect 3452 4366 3456 4370
rect 3462 4366 3466 4370
rect 3427 4361 3431 4365
rect 3437 4361 3441 4365
rect 3447 4361 3451 4365
rect 3457 4361 3461 4365
rect 3731 4446 3735 4450
rect 3741 4446 3745 4450
rect 3751 4446 3755 4450
rect 3761 4446 3765 4450
rect 3771 4446 3775 4450
rect 3736 4441 3740 4445
rect 3746 4441 3750 4445
rect 3756 4441 3760 4445
rect 3766 4441 3770 4445
rect 3731 4436 3735 4440
rect 3741 4436 3745 4440
rect 3751 4436 3755 4440
rect 3761 4436 3765 4440
rect 3771 4436 3775 4440
rect 3736 4431 3740 4435
rect 3746 4431 3750 4435
rect 3756 4431 3760 4435
rect 3766 4431 3770 4435
rect 3731 4426 3735 4430
rect 3741 4426 3745 4430
rect 3751 4426 3755 4430
rect 3761 4426 3765 4430
rect 3771 4426 3775 4430
rect 3736 4421 3740 4425
rect 3746 4421 3750 4425
rect 3756 4421 3760 4425
rect 3766 4421 3770 4425
rect 3731 4416 3735 4420
rect 3741 4416 3745 4420
rect 3751 4416 3755 4420
rect 3761 4416 3765 4420
rect 3771 4416 3775 4420
rect 3736 4411 3740 4415
rect 3746 4411 3750 4415
rect 3756 4411 3760 4415
rect 3766 4411 3770 4415
rect 3731 4406 3735 4410
rect 3741 4406 3745 4410
rect 3751 4406 3755 4410
rect 3761 4406 3765 4410
rect 3771 4406 3775 4410
rect 3736 4401 3740 4405
rect 3746 4401 3750 4405
rect 3756 4401 3760 4405
rect 3766 4401 3770 4405
rect 3731 4396 3735 4400
rect 3741 4396 3745 4400
rect 3751 4396 3755 4400
rect 3761 4396 3765 4400
rect 3771 4396 3775 4400
rect 3736 4391 3740 4395
rect 3746 4391 3750 4395
rect 3756 4391 3760 4395
rect 3766 4391 3770 4395
rect 3731 4386 3735 4390
rect 3741 4386 3745 4390
rect 3751 4386 3755 4390
rect 3761 4386 3765 4390
rect 3771 4386 3775 4390
rect 3736 4381 3740 4385
rect 3746 4381 3750 4385
rect 3756 4381 3760 4385
rect 3766 4381 3770 4385
rect 3731 4376 3735 4380
rect 3741 4376 3745 4380
rect 3751 4376 3755 4380
rect 3761 4376 3765 4380
rect 3771 4376 3775 4380
rect 3736 4371 3740 4375
rect 3746 4371 3750 4375
rect 3756 4371 3760 4375
rect 3766 4371 3770 4375
rect 3731 4366 3735 4370
rect 3741 4366 3745 4370
rect 3751 4366 3755 4370
rect 3761 4366 3765 4370
rect 3771 4366 3775 4370
rect 3736 4361 3740 4365
rect 3746 4361 3750 4365
rect 3756 4361 3760 4365
rect 3766 4361 3770 4365
<< pdcontact >>
rect 1562 9949 1566 9953
rect 1572 9949 1576 9953
rect 1582 9949 1586 9953
rect 1592 9949 1596 9953
rect 1557 9944 1561 9948
rect 1567 9944 1571 9948
rect 1577 9944 1581 9948
rect 1587 9944 1591 9948
rect 1597 9944 1601 9948
rect 1562 9939 1566 9943
rect 1572 9939 1576 9943
rect 1582 9939 1586 9943
rect 1592 9939 1596 9943
rect 1557 9934 1561 9938
rect 1567 9934 1571 9938
rect 1577 9934 1581 9938
rect 1587 9934 1591 9938
rect 1597 9934 1601 9938
rect 1562 9929 1566 9933
rect 1572 9929 1576 9933
rect 1582 9929 1586 9933
rect 1592 9929 1596 9933
rect 1557 9924 1561 9928
rect 1567 9924 1571 9928
rect 1577 9924 1581 9928
rect 1587 9924 1591 9928
rect 1597 9924 1601 9928
rect 1562 9919 1566 9923
rect 1572 9919 1576 9923
rect 1582 9919 1586 9923
rect 1592 9919 1596 9923
rect 1557 9914 1561 9918
rect 1567 9914 1571 9918
rect 1577 9914 1581 9918
rect 1587 9914 1591 9918
rect 1597 9914 1601 9918
rect 1562 9909 1566 9913
rect 1572 9909 1576 9913
rect 1582 9909 1586 9913
rect 1592 9909 1596 9913
rect 1557 9904 1561 9908
rect 1567 9904 1571 9908
rect 1577 9904 1581 9908
rect 1587 9904 1591 9908
rect 1597 9904 1601 9908
rect 1562 9899 1566 9903
rect 1572 9899 1576 9903
rect 1582 9899 1586 9903
rect 1592 9899 1596 9903
rect 1557 9894 1561 9898
rect 1567 9894 1571 9898
rect 1577 9894 1581 9898
rect 1587 9894 1591 9898
rect 1597 9894 1601 9898
rect 1562 9889 1566 9893
rect 1572 9889 1576 9893
rect 1582 9889 1586 9893
rect 1592 9889 1596 9893
rect 1557 9884 1561 9888
rect 1567 9884 1571 9888
rect 1577 9884 1581 9888
rect 1587 9884 1591 9888
rect 1597 9884 1601 9888
rect 1562 9879 1566 9883
rect 1572 9879 1576 9883
rect 1582 9879 1586 9883
rect 1592 9879 1596 9883
rect 1557 9874 1561 9878
rect 1567 9874 1571 9878
rect 1577 9874 1581 9878
rect 1587 9874 1591 9878
rect 1597 9874 1601 9878
rect 1562 9869 1566 9873
rect 1572 9869 1576 9873
rect 1582 9869 1586 9873
rect 1592 9869 1596 9873
rect 1557 9864 1561 9868
rect 1567 9864 1571 9868
rect 1577 9864 1581 9868
rect 1587 9864 1591 9868
rect 1597 9864 1601 9868
rect 1871 9949 1875 9953
rect 1881 9949 1885 9953
rect 1891 9949 1895 9953
rect 1901 9949 1905 9953
rect 1866 9944 1870 9948
rect 1876 9944 1880 9948
rect 1886 9944 1890 9948
rect 1896 9944 1900 9948
rect 1906 9944 1910 9948
rect 1871 9939 1875 9943
rect 1881 9939 1885 9943
rect 1891 9939 1895 9943
rect 1901 9939 1905 9943
rect 1866 9934 1870 9938
rect 1876 9934 1880 9938
rect 1886 9934 1890 9938
rect 1896 9934 1900 9938
rect 1906 9934 1910 9938
rect 1871 9929 1875 9933
rect 1881 9929 1885 9933
rect 1891 9929 1895 9933
rect 1901 9929 1905 9933
rect 1866 9924 1870 9928
rect 1876 9924 1880 9928
rect 1886 9924 1890 9928
rect 1896 9924 1900 9928
rect 1906 9924 1910 9928
rect 1871 9919 1875 9923
rect 1881 9919 1885 9923
rect 1891 9919 1895 9923
rect 1901 9919 1905 9923
rect 1866 9914 1870 9918
rect 1876 9914 1880 9918
rect 1886 9914 1890 9918
rect 1896 9914 1900 9918
rect 1906 9914 1910 9918
rect 1871 9909 1875 9913
rect 1881 9909 1885 9913
rect 1891 9909 1895 9913
rect 1901 9909 1905 9913
rect 1866 9904 1870 9908
rect 1876 9904 1880 9908
rect 1886 9904 1890 9908
rect 1896 9904 1900 9908
rect 1906 9904 1910 9908
rect 1871 9899 1875 9903
rect 1881 9899 1885 9903
rect 1891 9899 1895 9903
rect 1901 9899 1905 9903
rect 1866 9894 1870 9898
rect 1876 9894 1880 9898
rect 1886 9894 1890 9898
rect 1896 9894 1900 9898
rect 1906 9894 1910 9898
rect 1871 9889 1875 9893
rect 1881 9889 1885 9893
rect 1891 9889 1895 9893
rect 1901 9889 1905 9893
rect 1866 9884 1870 9888
rect 1876 9884 1880 9888
rect 1886 9884 1890 9888
rect 1896 9884 1900 9888
rect 1906 9884 1910 9888
rect 1871 9879 1875 9883
rect 1881 9879 1885 9883
rect 1891 9879 1895 9883
rect 1901 9879 1905 9883
rect 1866 9874 1870 9878
rect 1876 9874 1880 9878
rect 1886 9874 1890 9878
rect 1896 9874 1900 9878
rect 1906 9874 1910 9878
rect 1871 9869 1875 9873
rect 1881 9869 1885 9873
rect 1891 9869 1895 9873
rect 1901 9869 1905 9873
rect 1866 9864 1870 9868
rect 1876 9864 1880 9868
rect 1886 9864 1890 9868
rect 1896 9864 1900 9868
rect 1906 9864 1910 9868
rect 2180 9949 2184 9953
rect 2190 9949 2194 9953
rect 2200 9949 2204 9953
rect 2210 9949 2214 9953
rect 2175 9944 2179 9948
rect 2185 9944 2189 9948
rect 2195 9944 2199 9948
rect 2205 9944 2209 9948
rect 2215 9944 2219 9948
rect 2180 9939 2184 9943
rect 2190 9939 2194 9943
rect 2200 9939 2204 9943
rect 2210 9939 2214 9943
rect 2175 9934 2179 9938
rect 2185 9934 2189 9938
rect 2195 9934 2199 9938
rect 2205 9934 2209 9938
rect 2215 9934 2219 9938
rect 2180 9929 2184 9933
rect 2190 9929 2194 9933
rect 2200 9929 2204 9933
rect 2210 9929 2214 9933
rect 2175 9924 2179 9928
rect 2185 9924 2189 9928
rect 2195 9924 2199 9928
rect 2205 9924 2209 9928
rect 2215 9924 2219 9928
rect 2180 9919 2184 9923
rect 2190 9919 2194 9923
rect 2200 9919 2204 9923
rect 2210 9919 2214 9923
rect 2175 9914 2179 9918
rect 2185 9914 2189 9918
rect 2195 9914 2199 9918
rect 2205 9914 2209 9918
rect 2215 9914 2219 9918
rect 2180 9909 2184 9913
rect 2190 9909 2194 9913
rect 2200 9909 2204 9913
rect 2210 9909 2214 9913
rect 2175 9904 2179 9908
rect 2185 9904 2189 9908
rect 2195 9904 2199 9908
rect 2205 9904 2209 9908
rect 2215 9904 2219 9908
rect 2180 9899 2184 9903
rect 2190 9899 2194 9903
rect 2200 9899 2204 9903
rect 2210 9899 2214 9903
rect 2175 9894 2179 9898
rect 2185 9894 2189 9898
rect 2195 9894 2199 9898
rect 2205 9894 2209 9898
rect 2215 9894 2219 9898
rect 2180 9889 2184 9893
rect 2190 9889 2194 9893
rect 2200 9889 2204 9893
rect 2210 9889 2214 9893
rect 2175 9884 2179 9888
rect 2185 9884 2189 9888
rect 2195 9884 2199 9888
rect 2205 9884 2209 9888
rect 2215 9884 2219 9888
rect 2180 9879 2184 9883
rect 2190 9879 2194 9883
rect 2200 9879 2204 9883
rect 2210 9879 2214 9883
rect 2175 9874 2179 9878
rect 2185 9874 2189 9878
rect 2195 9874 2199 9878
rect 2205 9874 2209 9878
rect 2215 9874 2219 9878
rect 2180 9869 2184 9873
rect 2190 9869 2194 9873
rect 2200 9869 2204 9873
rect 2210 9869 2214 9873
rect 2175 9864 2179 9868
rect 2185 9864 2189 9868
rect 2195 9864 2199 9868
rect 2205 9864 2209 9868
rect 2215 9864 2219 9868
rect 2489 9949 2493 9953
rect 2499 9949 2503 9953
rect 2509 9949 2513 9953
rect 2519 9949 2523 9953
rect 2484 9944 2488 9948
rect 2494 9944 2498 9948
rect 2504 9944 2508 9948
rect 2514 9944 2518 9948
rect 2524 9944 2528 9948
rect 2489 9939 2493 9943
rect 2499 9939 2503 9943
rect 2509 9939 2513 9943
rect 2519 9939 2523 9943
rect 2484 9934 2488 9938
rect 2494 9934 2498 9938
rect 2504 9934 2508 9938
rect 2514 9934 2518 9938
rect 2524 9934 2528 9938
rect 2489 9929 2493 9933
rect 2499 9929 2503 9933
rect 2509 9929 2513 9933
rect 2519 9929 2523 9933
rect 2484 9924 2488 9928
rect 2494 9924 2498 9928
rect 2504 9924 2508 9928
rect 2514 9924 2518 9928
rect 2524 9924 2528 9928
rect 2489 9919 2493 9923
rect 2499 9919 2503 9923
rect 2509 9919 2513 9923
rect 2519 9919 2523 9923
rect 2484 9914 2488 9918
rect 2494 9914 2498 9918
rect 2504 9914 2508 9918
rect 2514 9914 2518 9918
rect 2524 9914 2528 9918
rect 2489 9909 2493 9913
rect 2499 9909 2503 9913
rect 2509 9909 2513 9913
rect 2519 9909 2523 9913
rect 2484 9904 2488 9908
rect 2494 9904 2498 9908
rect 2504 9904 2508 9908
rect 2514 9904 2518 9908
rect 2524 9904 2528 9908
rect 2489 9899 2493 9903
rect 2499 9899 2503 9903
rect 2509 9899 2513 9903
rect 2519 9899 2523 9903
rect 2484 9894 2488 9898
rect 2494 9894 2498 9898
rect 2504 9894 2508 9898
rect 2514 9894 2518 9898
rect 2524 9894 2528 9898
rect 2489 9889 2493 9893
rect 2499 9889 2503 9893
rect 2509 9889 2513 9893
rect 2519 9889 2523 9893
rect 2484 9884 2488 9888
rect 2494 9884 2498 9888
rect 2504 9884 2508 9888
rect 2514 9884 2518 9888
rect 2524 9884 2528 9888
rect 2489 9879 2493 9883
rect 2499 9879 2503 9883
rect 2509 9879 2513 9883
rect 2519 9879 2523 9883
rect 2484 9874 2488 9878
rect 2494 9874 2498 9878
rect 2504 9874 2508 9878
rect 2514 9874 2518 9878
rect 2524 9874 2528 9878
rect 2489 9869 2493 9873
rect 2499 9869 2503 9873
rect 2509 9869 2513 9873
rect 2519 9869 2523 9873
rect 2484 9864 2488 9868
rect 2494 9864 2498 9868
rect 2504 9864 2508 9868
rect 2514 9864 2518 9868
rect 2524 9864 2528 9868
rect 2798 9949 2802 9953
rect 2808 9949 2812 9953
rect 2818 9949 2822 9953
rect 2828 9949 2832 9953
rect 2793 9944 2797 9948
rect 2803 9944 2807 9948
rect 2813 9944 2817 9948
rect 2823 9944 2827 9948
rect 2833 9944 2837 9948
rect 2798 9939 2802 9943
rect 2808 9939 2812 9943
rect 2818 9939 2822 9943
rect 2828 9939 2832 9943
rect 2793 9934 2797 9938
rect 2803 9934 2807 9938
rect 2813 9934 2817 9938
rect 2823 9934 2827 9938
rect 2833 9934 2837 9938
rect 2798 9929 2802 9933
rect 2808 9929 2812 9933
rect 2818 9929 2822 9933
rect 2828 9929 2832 9933
rect 2793 9924 2797 9928
rect 2803 9924 2807 9928
rect 2813 9924 2817 9928
rect 2823 9924 2827 9928
rect 2833 9924 2837 9928
rect 2798 9919 2802 9923
rect 2808 9919 2812 9923
rect 2818 9919 2822 9923
rect 2828 9919 2832 9923
rect 2793 9914 2797 9918
rect 2803 9914 2807 9918
rect 2813 9914 2817 9918
rect 2823 9914 2827 9918
rect 2833 9914 2837 9918
rect 2798 9909 2802 9913
rect 2808 9909 2812 9913
rect 2818 9909 2822 9913
rect 2828 9909 2832 9913
rect 2793 9904 2797 9908
rect 2803 9904 2807 9908
rect 2813 9904 2817 9908
rect 2823 9904 2827 9908
rect 2833 9904 2837 9908
rect 2798 9899 2802 9903
rect 2808 9899 2812 9903
rect 2818 9899 2822 9903
rect 2828 9899 2832 9903
rect 2793 9894 2797 9898
rect 2803 9894 2807 9898
rect 2813 9894 2817 9898
rect 2823 9894 2827 9898
rect 2833 9894 2837 9898
rect 2798 9889 2802 9893
rect 2808 9889 2812 9893
rect 2818 9889 2822 9893
rect 2828 9889 2832 9893
rect 2793 9884 2797 9888
rect 2803 9884 2807 9888
rect 2813 9884 2817 9888
rect 2823 9884 2827 9888
rect 2833 9884 2837 9888
rect 2798 9879 2802 9883
rect 2808 9879 2812 9883
rect 2818 9879 2822 9883
rect 2828 9879 2832 9883
rect 2793 9874 2797 9878
rect 2803 9874 2807 9878
rect 2813 9874 2817 9878
rect 2823 9874 2827 9878
rect 2833 9874 2837 9878
rect 2798 9869 2802 9873
rect 2808 9869 2812 9873
rect 2818 9869 2822 9873
rect 2828 9869 2832 9873
rect 2793 9864 2797 9868
rect 2803 9864 2807 9868
rect 2813 9864 2817 9868
rect 2823 9864 2827 9868
rect 2833 9864 2837 9868
rect 3107 9949 3111 9953
rect 3117 9949 3121 9953
rect 3127 9949 3131 9953
rect 3137 9949 3141 9953
rect 3102 9944 3106 9948
rect 3112 9944 3116 9948
rect 3122 9944 3126 9948
rect 3132 9944 3136 9948
rect 3142 9944 3146 9948
rect 3107 9939 3111 9943
rect 3117 9939 3121 9943
rect 3127 9939 3131 9943
rect 3137 9939 3141 9943
rect 3102 9934 3106 9938
rect 3112 9934 3116 9938
rect 3122 9934 3126 9938
rect 3132 9934 3136 9938
rect 3142 9934 3146 9938
rect 3107 9929 3111 9933
rect 3117 9929 3121 9933
rect 3127 9929 3131 9933
rect 3137 9929 3141 9933
rect 3102 9924 3106 9928
rect 3112 9924 3116 9928
rect 3122 9924 3126 9928
rect 3132 9924 3136 9928
rect 3142 9924 3146 9928
rect 3107 9919 3111 9923
rect 3117 9919 3121 9923
rect 3127 9919 3131 9923
rect 3137 9919 3141 9923
rect 3102 9914 3106 9918
rect 3112 9914 3116 9918
rect 3122 9914 3126 9918
rect 3132 9914 3136 9918
rect 3142 9914 3146 9918
rect 3107 9909 3111 9913
rect 3117 9909 3121 9913
rect 3127 9909 3131 9913
rect 3137 9909 3141 9913
rect 3102 9904 3106 9908
rect 3112 9904 3116 9908
rect 3122 9904 3126 9908
rect 3132 9904 3136 9908
rect 3142 9904 3146 9908
rect 3107 9899 3111 9903
rect 3117 9899 3121 9903
rect 3127 9899 3131 9903
rect 3137 9899 3141 9903
rect 3102 9894 3106 9898
rect 3112 9894 3116 9898
rect 3122 9894 3126 9898
rect 3132 9894 3136 9898
rect 3142 9894 3146 9898
rect 3107 9889 3111 9893
rect 3117 9889 3121 9893
rect 3127 9889 3131 9893
rect 3137 9889 3141 9893
rect 3102 9884 3106 9888
rect 3112 9884 3116 9888
rect 3122 9884 3126 9888
rect 3132 9884 3136 9888
rect 3142 9884 3146 9888
rect 3107 9879 3111 9883
rect 3117 9879 3121 9883
rect 3127 9879 3131 9883
rect 3137 9879 3141 9883
rect 3102 9874 3106 9878
rect 3112 9874 3116 9878
rect 3122 9874 3126 9878
rect 3132 9874 3136 9878
rect 3142 9874 3146 9878
rect 3107 9869 3111 9873
rect 3117 9869 3121 9873
rect 3127 9869 3131 9873
rect 3137 9869 3141 9873
rect 3102 9864 3106 9868
rect 3112 9864 3116 9868
rect 3122 9864 3126 9868
rect 3132 9864 3136 9868
rect 3142 9864 3146 9868
rect 3416 9949 3420 9953
rect 3426 9949 3430 9953
rect 3436 9949 3440 9953
rect 3446 9949 3450 9953
rect 3411 9944 3415 9948
rect 3421 9944 3425 9948
rect 3431 9944 3435 9948
rect 3441 9944 3445 9948
rect 3451 9944 3455 9948
rect 3416 9939 3420 9943
rect 3426 9939 3430 9943
rect 3436 9939 3440 9943
rect 3446 9939 3450 9943
rect 3411 9934 3415 9938
rect 3421 9934 3425 9938
rect 3431 9934 3435 9938
rect 3441 9934 3445 9938
rect 3451 9934 3455 9938
rect 3416 9929 3420 9933
rect 3426 9929 3430 9933
rect 3436 9929 3440 9933
rect 3446 9929 3450 9933
rect 3411 9924 3415 9928
rect 3421 9924 3425 9928
rect 3431 9924 3435 9928
rect 3441 9924 3445 9928
rect 3451 9924 3455 9928
rect 3416 9919 3420 9923
rect 3426 9919 3430 9923
rect 3436 9919 3440 9923
rect 3446 9919 3450 9923
rect 3411 9914 3415 9918
rect 3421 9914 3425 9918
rect 3431 9914 3435 9918
rect 3441 9914 3445 9918
rect 3451 9914 3455 9918
rect 3416 9909 3420 9913
rect 3426 9909 3430 9913
rect 3436 9909 3440 9913
rect 3446 9909 3450 9913
rect 3411 9904 3415 9908
rect 3421 9904 3425 9908
rect 3431 9904 3435 9908
rect 3441 9904 3445 9908
rect 3451 9904 3455 9908
rect 3416 9899 3420 9903
rect 3426 9899 3430 9903
rect 3436 9899 3440 9903
rect 3446 9899 3450 9903
rect 3411 9894 3415 9898
rect 3421 9894 3425 9898
rect 3431 9894 3435 9898
rect 3441 9894 3445 9898
rect 3451 9894 3455 9898
rect 3416 9889 3420 9893
rect 3426 9889 3430 9893
rect 3436 9889 3440 9893
rect 3446 9889 3450 9893
rect 3411 9884 3415 9888
rect 3421 9884 3425 9888
rect 3431 9884 3435 9888
rect 3441 9884 3445 9888
rect 3451 9884 3455 9888
rect 3416 9879 3420 9883
rect 3426 9879 3430 9883
rect 3436 9879 3440 9883
rect 3446 9879 3450 9883
rect 3411 9874 3415 9878
rect 3421 9874 3425 9878
rect 3431 9874 3435 9878
rect 3441 9874 3445 9878
rect 3451 9874 3455 9878
rect 3416 9869 3420 9873
rect 3426 9869 3430 9873
rect 3436 9869 3440 9873
rect 3446 9869 3450 9873
rect 3411 9864 3415 9868
rect 3421 9864 3425 9868
rect 3431 9864 3435 9868
rect 3441 9864 3445 9868
rect 3451 9864 3455 9868
rect 3725 9949 3729 9953
rect 3735 9949 3739 9953
rect 3745 9949 3749 9953
rect 3755 9949 3759 9953
rect 3720 9944 3724 9948
rect 3730 9944 3734 9948
rect 3740 9944 3744 9948
rect 3750 9944 3754 9948
rect 3760 9944 3764 9948
rect 3725 9939 3729 9943
rect 3735 9939 3739 9943
rect 3745 9939 3749 9943
rect 3755 9939 3759 9943
rect 3720 9934 3724 9938
rect 3730 9934 3734 9938
rect 3740 9934 3744 9938
rect 3750 9934 3754 9938
rect 3760 9934 3764 9938
rect 3725 9929 3729 9933
rect 3735 9929 3739 9933
rect 3745 9929 3749 9933
rect 3755 9929 3759 9933
rect 3720 9924 3724 9928
rect 3730 9924 3734 9928
rect 3740 9924 3744 9928
rect 3750 9924 3754 9928
rect 3760 9924 3764 9928
rect 3725 9919 3729 9923
rect 3735 9919 3739 9923
rect 3745 9919 3749 9923
rect 3755 9919 3759 9923
rect 3720 9914 3724 9918
rect 3730 9914 3734 9918
rect 3740 9914 3744 9918
rect 3750 9914 3754 9918
rect 3760 9914 3764 9918
rect 3725 9909 3729 9913
rect 3735 9909 3739 9913
rect 3745 9909 3749 9913
rect 3755 9909 3759 9913
rect 3720 9904 3724 9908
rect 3730 9904 3734 9908
rect 3740 9904 3744 9908
rect 3750 9904 3754 9908
rect 3760 9904 3764 9908
rect 3725 9899 3729 9903
rect 3735 9899 3739 9903
rect 3745 9899 3749 9903
rect 3755 9899 3759 9903
rect 3720 9894 3724 9898
rect 3730 9894 3734 9898
rect 3740 9894 3744 9898
rect 3750 9894 3754 9898
rect 3760 9894 3764 9898
rect 3725 9889 3729 9893
rect 3735 9889 3739 9893
rect 3745 9889 3749 9893
rect 3755 9889 3759 9893
rect 3720 9884 3724 9888
rect 3730 9884 3734 9888
rect 3740 9884 3744 9888
rect 3750 9884 3754 9888
rect 3760 9884 3764 9888
rect 3725 9879 3729 9883
rect 3735 9879 3739 9883
rect 3745 9879 3749 9883
rect 3755 9879 3759 9883
rect 3720 9874 3724 9878
rect 3730 9874 3734 9878
rect 3740 9874 3744 9878
rect 3750 9874 3754 9878
rect 3760 9874 3764 9878
rect 3725 9869 3729 9873
rect 3735 9869 3739 9873
rect 3745 9869 3749 9873
rect 3755 9869 3759 9873
rect 3720 9864 3724 9868
rect 3730 9864 3734 9868
rect 3740 9864 3744 9868
rect 3750 9864 3754 9868
rect 3760 9864 3764 9868
rect 4034 9949 4038 9953
rect 4044 9949 4048 9953
rect 4054 9949 4058 9953
rect 4064 9949 4068 9953
rect 4029 9944 4033 9948
rect 4039 9944 4043 9948
rect 4049 9944 4053 9948
rect 4059 9944 4063 9948
rect 4069 9944 4073 9948
rect 4034 9939 4038 9943
rect 4044 9939 4048 9943
rect 4054 9939 4058 9943
rect 4064 9939 4068 9943
rect 4029 9934 4033 9938
rect 4039 9934 4043 9938
rect 4049 9934 4053 9938
rect 4059 9934 4063 9938
rect 4069 9934 4073 9938
rect 4034 9929 4038 9933
rect 4044 9929 4048 9933
rect 4054 9929 4058 9933
rect 4064 9929 4068 9933
rect 4029 9924 4033 9928
rect 4039 9924 4043 9928
rect 4049 9924 4053 9928
rect 4059 9924 4063 9928
rect 4069 9924 4073 9928
rect 4034 9919 4038 9923
rect 4044 9919 4048 9923
rect 4054 9919 4058 9923
rect 4064 9919 4068 9923
rect 4029 9914 4033 9918
rect 4039 9914 4043 9918
rect 4049 9914 4053 9918
rect 4059 9914 4063 9918
rect 4069 9914 4073 9918
rect 4034 9909 4038 9913
rect 4044 9909 4048 9913
rect 4054 9909 4058 9913
rect 4064 9909 4068 9913
rect 4029 9904 4033 9908
rect 4039 9904 4043 9908
rect 4049 9904 4053 9908
rect 4059 9904 4063 9908
rect 4069 9904 4073 9908
rect 4034 9899 4038 9903
rect 4044 9899 4048 9903
rect 4054 9899 4058 9903
rect 4064 9899 4068 9903
rect 4029 9894 4033 9898
rect 4039 9894 4043 9898
rect 4049 9894 4053 9898
rect 4059 9894 4063 9898
rect 4069 9894 4073 9898
rect 4034 9889 4038 9893
rect 4044 9889 4048 9893
rect 4054 9889 4058 9893
rect 4064 9889 4068 9893
rect 4029 9884 4033 9888
rect 4039 9884 4043 9888
rect 4049 9884 4053 9888
rect 4059 9884 4063 9888
rect 4069 9884 4073 9888
rect 4034 9879 4038 9883
rect 4044 9879 4048 9883
rect 4054 9879 4058 9883
rect 4064 9879 4068 9883
rect 4029 9874 4033 9878
rect 4039 9874 4043 9878
rect 4049 9874 4053 9878
rect 4059 9874 4063 9878
rect 4069 9874 4073 9878
rect 4034 9869 4038 9873
rect 4044 9869 4048 9873
rect 4054 9869 4058 9873
rect 4064 9869 4068 9873
rect 4029 9864 4033 9868
rect 4039 9864 4043 9868
rect 4049 9864 4053 9868
rect 4059 9864 4063 9868
rect 4069 9864 4073 9868
rect 1743 9827 1778 9831
rect 1782 9827 1799 9831
rect 2052 9827 2087 9831
rect 2091 9827 2108 9831
rect 2361 9827 2396 9831
rect 2400 9827 2417 9831
rect 2670 9827 2705 9831
rect 2709 9827 2726 9831
rect 2979 9827 3014 9831
rect 3018 9827 3035 9831
rect 3906 9827 3941 9831
rect 3945 9827 3962 9831
rect 1743 9819 1799 9823
rect 2052 9819 2108 9823
rect 2361 9819 2417 9823
rect 2670 9819 2726 9823
rect 2979 9819 3035 9823
rect 3906 9819 3962 9823
rect 1743 9811 1778 9815
rect 1782 9811 1799 9815
rect 2052 9811 2087 9815
rect 2091 9811 2108 9815
rect 1743 9803 1799 9807
rect 1743 9795 1778 9799
rect 1782 9795 1799 9799
rect 1743 9787 1799 9791
rect 2361 9811 2396 9815
rect 2400 9811 2417 9815
rect 2052 9803 2108 9807
rect 2052 9795 2087 9799
rect 2091 9795 2108 9799
rect 2052 9787 2108 9791
rect 2670 9811 2705 9815
rect 2709 9811 2726 9815
rect 2361 9803 2417 9807
rect 2361 9795 2396 9799
rect 2400 9795 2417 9799
rect 2361 9787 2417 9791
rect 2979 9811 3014 9815
rect 3018 9811 3035 9815
rect 2670 9803 2726 9807
rect 2670 9795 2705 9799
rect 2709 9795 2726 9799
rect 2670 9787 2726 9791
rect 3906 9811 3941 9815
rect 3945 9811 3962 9815
rect 2979 9803 3035 9807
rect 2979 9795 3014 9799
rect 3018 9795 3035 9799
rect 2979 9787 3035 9791
rect 3906 9803 3962 9807
rect 3906 9795 3941 9799
rect 3945 9795 3962 9799
rect 3906 9787 3962 9791
rect 1743 9779 1778 9783
rect 1782 9779 1799 9783
rect 2052 9779 2087 9783
rect 2091 9779 2108 9783
rect 2361 9779 2396 9783
rect 2400 9779 2417 9783
rect 2670 9779 2705 9783
rect 2709 9779 2726 9783
rect 2979 9779 3014 9783
rect 3018 9779 3035 9783
rect 3906 9779 3941 9783
rect 3945 9779 3962 9783
rect 423 6390 427 6457
rect 423 6369 427 6386
rect 431 6369 435 6457
rect 439 6390 443 6457
rect 439 6378 443 6386
rect 447 6369 451 6457
rect 464 6390 468 6457
rect 464 6369 468 6386
rect 472 6369 476 6457
rect 480 6390 484 6457
rect 480 6378 484 6386
rect 488 6369 492 6457
rect 507 6390 511 6457
rect 507 6369 511 6386
rect 515 6369 519 6457
rect 523 6390 527 6457
rect 523 6378 527 6386
rect 531 6369 535 6457
rect 546 6390 550 6425
rect 546 6369 550 6386
rect 554 6369 558 6425
rect 562 6390 566 6425
rect 562 6369 566 6386
rect 570 6369 574 6425
rect 578 6390 582 6425
rect 578 6369 582 6386
rect 586 6369 590 6425
rect 594 6390 598 6425
rect 594 6369 598 6386
rect 2851 9322 2855 9330
rect 2864 9322 2868 9330
rect 2872 9322 2876 9330
rect 2880 9326 2884 9330
rect 2888 9322 2892 9330
rect 2901 9322 2905 9330
rect 2914 9322 2918 9330
rect 2922 9322 2926 9330
rect 2930 9322 2934 9330
rect 2938 9326 2942 9330
rect 2946 9322 2950 9330
rect 2959 9322 2963 9330
rect 2967 9322 2971 9330
rect 2975 9322 2979 9330
rect 2983 9322 2987 9330
rect 2996 9322 3000 9330
rect 3004 9322 3008 9330
rect 3012 9326 3016 9330
rect 3020 9322 3024 9330
rect 3033 9322 3037 9330
rect 3046 9322 3050 9330
rect 3054 9322 3058 9330
rect 3062 9322 3066 9330
rect 3070 9326 3074 9330
rect 3078 9322 3082 9330
rect 3091 9322 3095 9330
rect 3099 9322 3103 9330
rect 3107 9322 3111 9330
rect 3115 9322 3119 9330
rect 3128 9322 3132 9330
rect 3136 9322 3140 9330
rect 3144 9326 3148 9330
rect 3152 9322 3156 9330
rect 3165 9322 3169 9330
rect 3178 9322 3182 9330
rect 3186 9322 3190 9330
rect 3194 9322 3198 9330
rect 3202 9326 3206 9330
rect 3210 9322 3214 9330
rect 3223 9322 3227 9330
rect 3231 9322 3235 9330
rect 3239 9322 3243 9330
rect 3247 9322 3251 9330
rect 3260 9322 3264 9330
rect 3268 9322 3272 9330
rect 3276 9326 3280 9330
rect 3284 9322 3288 9330
rect 3297 9322 3301 9330
rect 3310 9322 3314 9330
rect 3318 9322 3322 9330
rect 3326 9322 3330 9330
rect 3334 9326 3338 9330
rect 3342 9322 3346 9330
rect 3355 9322 3359 9330
rect 3363 9322 3367 9330
rect 3371 9322 3375 9330
rect 3796 9322 3800 9330
rect 3809 9322 3813 9330
rect 3817 9322 3821 9330
rect 3825 9326 3829 9330
rect 3833 9322 3837 9330
rect 3846 9322 3850 9330
rect 3859 9322 3863 9330
rect 3867 9322 3871 9330
rect 3875 9322 3879 9330
rect 3883 9326 3887 9330
rect 3891 9322 3895 9330
rect 3904 9322 3908 9330
rect 3912 9322 3916 9330
rect 3920 9322 3924 9330
rect 3928 9322 3932 9330
rect 3941 9322 3945 9330
rect 3949 9322 3953 9330
rect 3957 9326 3961 9330
rect 3965 9322 3969 9330
rect 3978 9322 3982 9330
rect 3991 9322 3995 9330
rect 3999 9322 4003 9330
rect 4007 9322 4011 9330
rect 4015 9326 4019 9330
rect 4023 9322 4027 9330
rect 4036 9322 4040 9330
rect 4044 9322 4048 9330
rect 4052 9322 4056 9330
rect 4060 9322 4064 9330
rect 4073 9322 4077 9330
rect 4081 9322 4085 9330
rect 4089 9326 4093 9330
rect 4097 9322 4101 9330
rect 4110 9322 4114 9330
rect 4123 9322 4127 9330
rect 4131 9322 4135 9330
rect 4139 9322 4143 9330
rect 4147 9326 4151 9330
rect 4155 9322 4159 9330
rect 4168 9322 4172 9330
rect 4176 9322 4180 9330
rect 4184 9322 4188 9330
rect 4192 9322 4196 9330
rect 4205 9322 4209 9330
rect 4213 9322 4217 9330
rect 4221 9326 4225 9330
rect 4229 9322 4233 9330
rect 4242 9322 4246 9330
rect 4255 9322 4259 9330
rect 4263 9322 4267 9330
rect 4271 9322 4275 9330
rect 4279 9326 4283 9330
rect 4287 9322 4291 9330
rect 4300 9322 4304 9330
rect 4308 9322 4312 9330
rect 4316 9322 4320 9330
rect 2499 9289 2503 9297
rect 2512 9289 2516 9297
rect 2520 9289 2524 9297
rect 2528 9293 2532 9297
rect 2536 9289 2540 9297
rect 2549 9289 2553 9297
rect 2562 9289 2566 9297
rect 2570 9289 2574 9297
rect 2578 9289 2582 9297
rect 2586 9293 2590 9297
rect 2594 9289 2598 9297
rect 2607 9289 2611 9297
rect 2615 9289 2619 9297
rect 2623 9289 2627 9297
rect 3444 9289 3448 9297
rect 3457 9289 3461 9297
rect 3465 9289 3469 9297
rect 3473 9293 3477 9297
rect 3481 9289 3485 9297
rect 3494 9289 3498 9297
rect 3507 9289 3511 9297
rect 3515 9289 3519 9297
rect 3523 9289 3527 9297
rect 3531 9293 3535 9297
rect 3539 9289 3543 9297
rect 3552 9289 3556 9297
rect 3560 9289 3564 9297
rect 3568 9289 3572 9297
rect 3030 9251 3034 9259
rect 3038 9251 3042 9259
rect 2856 9238 2860 9246
rect 2864 9238 2868 9246
rect 2872 9238 2876 9246
rect 2880 9238 2884 9246
rect 2888 9238 2892 9246
rect 2896 9238 2900 9246
rect 2907 9238 2911 9246
rect 2924 9238 2928 9246
rect 2941 9238 2945 9246
rect 2950 9238 2954 9246
rect 2963 9238 2967 9246
rect 2971 9238 2975 9246
rect 2979 9238 2983 9246
rect 2996 9238 3000 9246
rect 3006 9238 3010 9246
rect 3014 9238 3018 9246
rect 3054 9245 3058 9253
rect 3069 9245 3073 9253
rect 3084 9251 3088 9259
rect 3092 9251 3096 9259
rect 3111 9251 3115 9259
rect 3119 9251 3123 9259
rect 3135 9245 3139 9253
rect 3150 9245 3154 9253
rect 3165 9251 3169 9259
rect 3173 9251 3177 9259
rect 3975 9251 3979 9259
rect 3983 9251 3987 9259
rect 3801 9238 3805 9246
rect 3809 9238 3813 9246
rect 3817 9238 3821 9246
rect 3825 9238 3829 9246
rect 3833 9238 3837 9246
rect 3841 9238 3845 9246
rect 3852 9238 3856 9246
rect 3869 9238 3873 9246
rect 3886 9238 3890 9246
rect 3895 9238 3899 9246
rect 3908 9238 3912 9246
rect 3916 9238 3920 9246
rect 3924 9238 3928 9246
rect 3941 9238 3945 9246
rect 3951 9238 3955 9246
rect 3959 9238 3963 9246
rect 3999 9245 4003 9253
rect 4014 9245 4018 9253
rect 4029 9251 4033 9259
rect 4037 9251 4041 9259
rect 4056 9251 4060 9259
rect 4064 9251 4068 9259
rect 4080 9245 4084 9253
rect 4095 9245 4099 9253
rect 4110 9251 4114 9259
rect 4118 9251 4122 9259
rect 2490 9187 2494 9195
rect 2498 9187 2502 9195
rect 2506 9187 2510 9195
rect 2519 9187 2523 9195
rect 2527 9191 2531 9195
rect 2535 9187 2539 9195
rect 2543 9187 2547 9195
rect 2551 9187 2555 9195
rect 2564 9187 2568 9195
rect 2577 9187 2581 9195
rect 2585 9191 2589 9195
rect 2593 9187 2597 9195
rect 2601 9187 2605 9195
rect 2614 9187 2618 9195
rect 3435 9187 3439 9195
rect 3443 9187 3447 9195
rect 3451 9187 3455 9195
rect 3464 9187 3468 9195
rect 3472 9191 3476 9195
rect 3480 9187 3484 9195
rect 3488 9187 3492 9195
rect 3496 9187 3500 9195
rect 3509 9187 3513 9195
rect 3522 9187 3526 9195
rect 3530 9191 3534 9195
rect 3538 9187 3542 9195
rect 3546 9187 3550 9195
rect 3559 9187 3563 9195
rect 2856 9152 2860 9160
rect 2864 9152 2868 9160
rect 2872 9152 2876 9160
rect 2880 9152 2884 9160
rect 2888 9152 2892 9160
rect 2896 9152 2900 9160
rect 2907 9152 2911 9160
rect 2924 9152 2928 9160
rect 2941 9152 2945 9160
rect 2950 9152 2954 9160
rect 2963 9152 2967 9160
rect 2971 9152 2975 9160
rect 2979 9152 2983 9160
rect 2996 9152 3000 9160
rect 3006 9152 3010 9160
rect 3014 9152 3018 9160
rect 3054 9153 3058 9161
rect 3069 9153 3073 9161
rect 3135 9153 3139 9161
rect 3150 9153 3154 9161
rect 3801 9152 3805 9160
rect 3809 9152 3813 9160
rect 3817 9152 3821 9160
rect 3825 9152 3829 9160
rect 3833 9152 3837 9160
rect 3841 9152 3845 9160
rect 3852 9152 3856 9160
rect 3869 9152 3873 9160
rect 3886 9152 3890 9160
rect 3895 9152 3899 9160
rect 3908 9152 3912 9160
rect 3916 9152 3920 9160
rect 3924 9152 3928 9160
rect 3941 9152 3945 9160
rect 3951 9152 3955 9160
rect 3959 9152 3963 9160
rect 3999 9153 4003 9161
rect 4014 9153 4018 9161
rect 4080 9153 4084 9161
rect 4095 9153 4099 9161
rect 2856 9106 2860 9114
rect 2864 9106 2868 9114
rect 2872 9106 2876 9114
rect 2880 9106 2884 9114
rect 2888 9106 2892 9114
rect 2896 9106 2900 9114
rect 2907 9106 2911 9114
rect 2924 9106 2928 9114
rect 2941 9106 2945 9114
rect 2950 9106 2954 9114
rect 2963 9106 2967 9114
rect 2971 9106 2975 9114
rect 2979 9106 2983 9114
rect 2996 9106 3000 9114
rect 3006 9106 3010 9114
rect 3014 9106 3018 9114
rect 3054 9113 3058 9121
rect 3069 9113 3073 9121
rect 3084 9119 3088 9127
rect 3092 9119 3096 9127
rect 3135 9119 3139 9127
rect 3143 9119 3147 9127
rect 3159 9113 3163 9121
rect 3174 9113 3178 9121
rect 3189 9119 3193 9127
rect 3197 9119 3201 9127
rect 3801 9106 3805 9114
rect 3809 9106 3813 9114
rect 3817 9106 3821 9114
rect 3825 9106 3829 9114
rect 3833 9106 3837 9114
rect 3841 9106 3845 9114
rect 3852 9106 3856 9114
rect 3869 9106 3873 9114
rect 3886 9106 3890 9114
rect 3895 9106 3899 9114
rect 3908 9106 3912 9114
rect 3916 9106 3920 9114
rect 3924 9106 3928 9114
rect 3941 9106 3945 9114
rect 3951 9106 3955 9114
rect 3959 9106 3963 9114
rect 3999 9113 4003 9121
rect 4014 9113 4018 9121
rect 4029 9119 4033 9127
rect 4037 9119 4041 9127
rect 4080 9119 4084 9127
rect 4088 9119 4092 9127
rect 3366 9090 3370 9098
rect 3374 9090 3378 9098
rect 3390 9084 3394 9092
rect 3405 9084 3409 9092
rect 3420 9090 3424 9098
rect 3428 9090 3432 9098
rect 3540 9065 3556 9095
rect 3560 9065 3576 9095
rect 3593 9065 3609 9095
rect 3613 9065 3629 9095
rect 4104 9113 4108 9121
rect 4119 9113 4123 9121
rect 4134 9119 4138 9127
rect 4142 9119 4146 9127
rect 2856 9020 2860 9028
rect 2864 9020 2868 9028
rect 2872 9020 2876 9028
rect 2880 9020 2884 9028
rect 2888 9020 2892 9028
rect 2896 9020 2900 9028
rect 2907 9020 2911 9028
rect 2924 9020 2928 9028
rect 2941 9020 2945 9028
rect 2950 9020 2954 9028
rect 2963 9020 2967 9028
rect 2971 9020 2975 9028
rect 2979 9020 2983 9028
rect 2996 9020 3000 9028
rect 3006 9020 3010 9028
rect 3014 9020 3018 9028
rect 3054 9022 3058 9030
rect 3069 9022 3073 9030
rect 3159 9022 3163 9030
rect 3174 9022 3178 9030
rect 3801 9020 3805 9028
rect 3809 9020 3813 9028
rect 3817 9020 3821 9028
rect 3825 9020 3829 9028
rect 3833 9020 3837 9028
rect 3841 9020 3845 9028
rect 3852 9020 3856 9028
rect 3869 9020 3873 9028
rect 3886 9020 3890 9028
rect 3895 9020 3899 9028
rect 3908 9020 3912 9028
rect 3916 9020 3920 9028
rect 3924 9020 3928 9028
rect 3941 9020 3945 9028
rect 3951 9020 3955 9028
rect 3959 9020 3963 9028
rect 3999 9022 4003 9030
rect 4014 9022 4018 9030
rect 4104 9022 4108 9030
rect 4119 9022 4123 9030
rect 2856 8974 2860 8982
rect 2864 8974 2868 8982
rect 2872 8974 2876 8982
rect 2880 8974 2884 8982
rect 2888 8974 2892 8982
rect 2896 8974 2900 8982
rect 2907 8974 2911 8982
rect 2924 8974 2928 8982
rect 2941 8974 2945 8982
rect 2950 8974 2954 8982
rect 2963 8974 2967 8982
rect 2971 8974 2975 8982
rect 2979 8974 2983 8982
rect 2996 8974 3000 8982
rect 3006 8974 3010 8982
rect 3014 8974 3018 8982
rect 3054 8981 3058 8989
rect 3069 8981 3073 8989
rect 3084 8987 3088 8995
rect 3092 8987 3096 8995
rect 3111 8987 3115 8995
rect 3119 8987 3123 8995
rect 3135 8981 3139 8989
rect 3150 8981 3154 8989
rect 3165 8987 3169 8995
rect 3173 8987 3177 8995
rect 3201 8987 3205 8995
rect 3209 8987 3213 8995
rect 3225 8981 3229 8989
rect 3240 8981 3244 8989
rect 3255 8987 3259 8995
rect 3263 8987 3267 8995
rect 3390 8988 3394 8996
rect 3405 8988 3409 8996
rect 3801 8974 3805 8982
rect 3809 8974 3813 8982
rect 3817 8974 3821 8982
rect 3825 8974 3829 8982
rect 3833 8974 3837 8982
rect 3841 8974 3845 8982
rect 3852 8974 3856 8982
rect 3869 8974 3873 8982
rect 3886 8974 3890 8982
rect 3895 8974 3899 8982
rect 3908 8974 3912 8982
rect 3916 8974 3920 8982
rect 3924 8974 3928 8982
rect 3941 8974 3945 8982
rect 3951 8974 3955 8982
rect 3959 8974 3963 8982
rect 3999 8981 4003 8989
rect 4014 8981 4018 8989
rect 4029 8987 4033 8995
rect 4037 8987 4041 8995
rect 4056 8987 4060 8995
rect 4064 8987 4068 8995
rect 3344 8960 3348 8968
rect 3352 8960 3356 8968
rect 3366 8960 3370 8968
rect 3374 8960 3378 8968
rect 3390 8954 3394 8962
rect 3405 8954 3409 8962
rect 3420 8960 3424 8968
rect 3428 8960 3432 8968
rect 3446 8935 3462 8965
rect 3466 8935 3482 8965
rect 3499 8935 3515 8965
rect 3519 8935 3535 8965
rect 4080 8981 4084 8989
rect 4095 8981 4099 8989
rect 4110 8987 4114 8995
rect 4118 8987 4122 8995
rect 4146 8987 4150 8995
rect 4154 8987 4158 8995
rect 4170 8981 4174 8989
rect 4185 8981 4189 8989
rect 4200 8987 4204 8995
rect 4208 8987 4212 8995
rect 2856 8888 2860 8896
rect 2864 8888 2868 8896
rect 2872 8888 2876 8896
rect 2880 8888 2884 8896
rect 2888 8888 2892 8896
rect 2896 8888 2900 8896
rect 2907 8888 2911 8896
rect 2924 8888 2928 8896
rect 2941 8888 2945 8896
rect 2950 8888 2954 8896
rect 2963 8888 2967 8896
rect 2971 8888 2975 8896
rect 2979 8888 2983 8896
rect 2996 8888 3000 8896
rect 3006 8888 3010 8896
rect 3014 8888 3018 8896
rect 3054 8887 3058 8895
rect 3069 8887 3073 8895
rect 3135 8887 3139 8895
rect 3150 8887 3154 8895
rect 3225 8887 3229 8895
rect 3240 8887 3244 8895
rect 3801 8888 3805 8896
rect 3809 8888 3813 8896
rect 3817 8888 3821 8896
rect 3825 8888 3829 8896
rect 3833 8888 3837 8896
rect 3841 8888 3845 8896
rect 3852 8888 3856 8896
rect 3869 8888 3873 8896
rect 3886 8888 3890 8896
rect 3895 8888 3899 8896
rect 3908 8888 3912 8896
rect 3916 8888 3920 8896
rect 3924 8888 3928 8896
rect 3941 8888 3945 8896
rect 3951 8888 3955 8896
rect 3959 8888 3963 8896
rect 3999 8887 4003 8895
rect 4014 8887 4018 8895
rect 4080 8887 4084 8895
rect 4095 8887 4099 8895
rect 4170 8887 4174 8895
rect 4185 8887 4189 8895
rect 2856 8842 2860 8850
rect 2864 8842 2868 8850
rect 2872 8842 2876 8850
rect 2880 8842 2884 8850
rect 2888 8842 2892 8850
rect 2896 8842 2900 8850
rect 2907 8842 2911 8850
rect 2924 8842 2928 8850
rect 2941 8842 2945 8850
rect 2950 8842 2954 8850
rect 2963 8842 2967 8850
rect 2971 8842 2975 8850
rect 2979 8842 2983 8850
rect 2996 8842 3000 8850
rect 3006 8842 3010 8850
rect 3014 8842 3018 8850
rect 3054 8849 3058 8857
rect 3069 8849 3073 8857
rect 3084 8855 3088 8863
rect 3092 8855 3096 8863
rect 3390 8858 3394 8866
rect 3405 8858 3409 8866
rect 3801 8842 3805 8850
rect 3809 8842 3813 8850
rect 3817 8842 3821 8850
rect 3825 8842 3829 8850
rect 3833 8842 3837 8850
rect 3841 8842 3845 8850
rect 3852 8842 3856 8850
rect 3869 8842 3873 8850
rect 3886 8842 3890 8850
rect 3895 8842 3899 8850
rect 3908 8842 3912 8850
rect 3916 8842 3920 8850
rect 3924 8842 3928 8850
rect 3941 8842 3945 8850
rect 3951 8842 3955 8850
rect 3959 8842 3963 8850
rect 3999 8849 4003 8857
rect 4014 8849 4018 8857
rect 4029 8855 4033 8863
rect 4037 8855 4041 8863
rect 2367 8787 2371 8795
rect 2380 8787 2384 8795
rect 2388 8787 2392 8795
rect 2396 8791 2400 8795
rect 2404 8787 2408 8795
rect 2417 8787 2421 8795
rect 2430 8787 2434 8795
rect 2438 8787 2442 8795
rect 2446 8787 2450 8795
rect 2454 8791 2458 8795
rect 2462 8787 2466 8795
rect 2475 8787 2479 8795
rect 2483 8787 2487 8795
rect 2491 8787 2495 8795
rect 2499 8787 2503 8795
rect 2512 8787 2516 8795
rect 2520 8787 2524 8795
rect 2528 8791 2532 8795
rect 2536 8787 2540 8795
rect 2549 8787 2553 8795
rect 2562 8787 2566 8795
rect 2570 8787 2574 8795
rect 2578 8787 2582 8795
rect 2586 8791 2590 8795
rect 2594 8787 2598 8795
rect 2607 8787 2611 8795
rect 2615 8787 2619 8795
rect 2623 8787 2627 8795
rect 2631 8787 2635 8795
rect 2644 8787 2648 8795
rect 2652 8787 2656 8795
rect 2660 8791 2664 8795
rect 2668 8787 2672 8795
rect 2681 8787 2685 8795
rect 2694 8787 2698 8795
rect 2702 8787 2706 8795
rect 2710 8787 2714 8795
rect 2718 8791 2722 8795
rect 2726 8787 2730 8795
rect 2739 8787 2743 8795
rect 2747 8787 2751 8795
rect 2755 8787 2759 8795
rect 3312 8787 3316 8795
rect 3325 8787 3329 8795
rect 3333 8787 3337 8795
rect 3341 8791 3345 8795
rect 3349 8787 3353 8795
rect 3362 8787 3366 8795
rect 3375 8787 3379 8795
rect 3383 8787 3387 8795
rect 3391 8787 3395 8795
rect 3399 8791 3403 8795
rect 3407 8787 3411 8795
rect 3420 8787 3424 8795
rect 3428 8787 3432 8795
rect 3436 8787 3440 8795
rect 3444 8787 3448 8795
rect 3457 8787 3461 8795
rect 3465 8787 3469 8795
rect 3473 8791 3477 8795
rect 3481 8787 3485 8795
rect 3494 8787 3498 8795
rect 3507 8787 3511 8795
rect 3515 8787 3519 8795
rect 3523 8787 3527 8795
rect 3531 8791 3535 8795
rect 3539 8787 3543 8795
rect 3552 8787 3556 8795
rect 3560 8787 3564 8795
rect 3568 8787 3572 8795
rect 3576 8787 3580 8795
rect 3589 8787 3593 8795
rect 3597 8787 3601 8795
rect 3605 8791 3609 8795
rect 3613 8787 3617 8795
rect 3626 8787 3630 8795
rect 3639 8787 3643 8795
rect 3647 8787 3651 8795
rect 3655 8787 3659 8795
rect 3663 8791 3667 8795
rect 3671 8787 3675 8795
rect 3684 8787 3688 8795
rect 3692 8787 3696 8795
rect 3700 8787 3704 8795
rect 2856 8756 2860 8764
rect 2864 8756 2868 8764
rect 2872 8756 2876 8764
rect 2880 8756 2884 8764
rect 2888 8756 2892 8764
rect 2896 8756 2900 8764
rect 2907 8756 2911 8764
rect 2924 8756 2928 8764
rect 2941 8756 2945 8764
rect 2950 8756 2954 8764
rect 2963 8756 2967 8764
rect 2971 8756 2975 8764
rect 2979 8756 2983 8764
rect 2996 8756 3000 8764
rect 3006 8756 3010 8764
rect 3014 8756 3018 8764
rect 3054 8751 3058 8759
rect 3069 8751 3073 8759
rect 3090 8756 3094 8764
rect 3098 8756 3102 8764
rect 3108 8756 3112 8764
rect 3116 8756 3120 8764
rect 3125 8756 3129 8764
rect 3133 8756 3137 8764
rect 3141 8756 3145 8764
rect 3149 8756 3153 8764
rect 3157 8756 3161 8764
rect 3168 8756 3172 8764
rect 3185 8756 3189 8764
rect 3202 8756 3206 8764
rect 3211 8756 3215 8764
rect 3224 8756 3228 8764
rect 3232 8756 3236 8764
rect 3240 8756 3244 8764
rect 3257 8756 3261 8764
rect 3267 8756 3271 8764
rect 3275 8756 3279 8764
rect 3801 8756 3805 8764
rect 3809 8756 3813 8764
rect 3817 8756 3821 8764
rect 3825 8756 3829 8764
rect 3833 8756 3837 8764
rect 3841 8756 3845 8764
rect 3852 8756 3856 8764
rect 3869 8756 3873 8764
rect 3886 8756 3890 8764
rect 3895 8756 3899 8764
rect 3908 8756 3912 8764
rect 3916 8756 3920 8764
rect 3924 8756 3928 8764
rect 3941 8756 3945 8764
rect 3951 8756 3955 8764
rect 3959 8756 3963 8764
rect 3999 8751 4003 8759
rect 4014 8751 4018 8759
rect 4035 8756 4039 8764
rect 4043 8756 4047 8764
rect 4053 8756 4057 8764
rect 4061 8756 4065 8764
rect 4070 8756 4074 8764
rect 4078 8756 4082 8764
rect 4086 8756 4090 8764
rect 4094 8756 4098 8764
rect 4102 8756 4106 8764
rect 4113 8756 4117 8764
rect 4130 8756 4134 8764
rect 4147 8756 4151 8764
rect 4156 8756 4160 8764
rect 4169 8756 4173 8764
rect 4177 8756 4181 8764
rect 4185 8756 4189 8764
rect 4202 8756 4206 8764
rect 4212 8756 4216 8764
rect 4220 8756 4224 8764
rect 3150 8675 3154 8683
rect 3163 8675 3167 8683
rect 3171 8675 3175 8683
rect 3179 8679 3183 8683
rect 3187 8675 3191 8683
rect 3200 8675 3204 8683
rect 3213 8675 3217 8683
rect 3221 8675 3225 8683
rect 3229 8675 3233 8683
rect 3237 8679 3241 8683
rect 3245 8675 3249 8683
rect 3258 8675 3262 8683
rect 3266 8675 3270 8683
rect 3274 8675 3278 8683
rect 4095 8675 4099 8683
rect 4108 8675 4112 8683
rect 4116 8675 4120 8683
rect 4124 8679 4128 8683
rect 4132 8675 4136 8683
rect 4145 8675 4149 8683
rect 4158 8675 4162 8683
rect 4166 8675 4170 8683
rect 4174 8675 4178 8683
rect 4182 8679 4186 8683
rect 4190 8675 4194 8683
rect 4203 8675 4207 8683
rect 4211 8675 4215 8683
rect 4219 8675 4223 8683
rect 2367 8645 2371 8653
rect 2380 8645 2384 8653
rect 2388 8645 2392 8653
rect 2396 8649 2400 8653
rect 2404 8645 2408 8653
rect 2417 8645 2421 8653
rect 2430 8645 2434 8653
rect 2438 8645 2442 8653
rect 2446 8645 2450 8653
rect 2454 8649 2458 8653
rect 2462 8645 2466 8653
rect 2475 8645 2479 8653
rect 2483 8645 2487 8653
rect 2491 8645 2495 8653
rect 2499 8645 2503 8653
rect 2512 8645 2516 8653
rect 2520 8645 2524 8653
rect 2528 8649 2532 8653
rect 2536 8645 2540 8653
rect 2549 8645 2553 8653
rect 2562 8645 2566 8653
rect 2570 8645 2574 8653
rect 2578 8645 2582 8653
rect 2586 8649 2590 8653
rect 2594 8645 2598 8653
rect 2607 8645 2611 8653
rect 2615 8645 2619 8653
rect 2623 8645 2627 8653
rect 2631 8645 2635 8653
rect 2644 8645 2648 8653
rect 2652 8645 2656 8653
rect 2660 8649 2664 8653
rect 2668 8645 2672 8653
rect 2681 8645 2685 8653
rect 2694 8645 2698 8653
rect 2702 8645 2706 8653
rect 2710 8645 2714 8653
rect 2718 8649 2722 8653
rect 2726 8645 2730 8653
rect 2739 8645 2743 8653
rect 2747 8645 2751 8653
rect 2755 8645 2759 8653
rect 3312 8645 3316 8653
rect 3325 8645 3329 8653
rect 3333 8645 3337 8653
rect 3341 8649 3345 8653
rect 3349 8645 3353 8653
rect 3362 8645 3366 8653
rect 3375 8645 3379 8653
rect 3383 8645 3387 8653
rect 3391 8645 3395 8653
rect 3399 8649 3403 8653
rect 3407 8645 3411 8653
rect 3420 8645 3424 8653
rect 3428 8645 3432 8653
rect 3436 8645 3440 8653
rect 3444 8645 3448 8653
rect 3457 8645 3461 8653
rect 3465 8645 3469 8653
rect 3473 8649 3477 8653
rect 3481 8645 3485 8653
rect 3494 8645 3498 8653
rect 3507 8645 3511 8653
rect 3515 8645 3519 8653
rect 3523 8645 3527 8653
rect 3531 8649 3535 8653
rect 3539 8645 3543 8653
rect 3552 8645 3556 8653
rect 3560 8645 3564 8653
rect 3568 8645 3572 8653
rect 3576 8645 3580 8653
rect 3589 8645 3593 8653
rect 3597 8645 3601 8653
rect 3605 8649 3609 8653
rect 3613 8645 3617 8653
rect 3626 8645 3630 8653
rect 3639 8645 3643 8653
rect 3647 8645 3651 8653
rect 3655 8645 3659 8653
rect 3663 8649 3667 8653
rect 3671 8645 3675 8653
rect 3684 8645 3688 8653
rect 3692 8645 3696 8653
rect 3700 8645 3704 8653
rect 3150 8589 3154 8597
rect 3163 8589 3167 8597
rect 3171 8589 3175 8597
rect 3179 8593 3183 8597
rect 3187 8589 3191 8597
rect 3200 8589 3204 8597
rect 3213 8589 3217 8597
rect 3221 8589 3225 8597
rect 3229 8589 3233 8597
rect 3237 8593 3241 8597
rect 3245 8589 3249 8597
rect 3258 8589 3262 8597
rect 3266 8589 3270 8597
rect 3274 8589 3278 8597
rect 4095 8589 4099 8597
rect 4108 8589 4112 8597
rect 4116 8589 4120 8597
rect 4124 8593 4128 8597
rect 4132 8589 4136 8597
rect 4145 8589 4149 8597
rect 4158 8589 4162 8597
rect 4166 8589 4170 8597
rect 4174 8589 4178 8597
rect 4182 8593 4186 8597
rect 4190 8589 4194 8597
rect 4203 8589 4207 8597
rect 4211 8589 4215 8597
rect 4219 8589 4223 8597
rect 2367 8559 2371 8567
rect 2380 8559 2384 8567
rect 2388 8559 2392 8567
rect 2396 8563 2400 8567
rect 2404 8559 2408 8567
rect 2417 8559 2421 8567
rect 2430 8559 2434 8567
rect 2438 8559 2442 8567
rect 2446 8559 2450 8567
rect 2454 8563 2458 8567
rect 2462 8559 2466 8567
rect 2475 8559 2479 8567
rect 2483 8559 2487 8567
rect 2491 8559 2495 8567
rect 2499 8559 2503 8567
rect 2512 8559 2516 8567
rect 2520 8559 2524 8567
rect 2528 8563 2532 8567
rect 2536 8559 2540 8567
rect 2549 8559 2553 8567
rect 2562 8559 2566 8567
rect 2570 8559 2574 8567
rect 2578 8559 2582 8567
rect 2586 8563 2590 8567
rect 2594 8559 2598 8567
rect 2607 8559 2611 8567
rect 2615 8559 2619 8567
rect 2623 8559 2627 8567
rect 2631 8559 2635 8567
rect 2644 8559 2648 8567
rect 2652 8559 2656 8567
rect 2660 8563 2664 8567
rect 2668 8559 2672 8567
rect 2681 8559 2685 8567
rect 2694 8559 2698 8567
rect 2702 8559 2706 8567
rect 2710 8559 2714 8567
rect 2718 8563 2722 8567
rect 2726 8559 2730 8567
rect 2739 8559 2743 8567
rect 2747 8559 2751 8567
rect 2755 8559 2759 8567
rect 3312 8559 3316 8567
rect 3325 8559 3329 8567
rect 3333 8559 3337 8567
rect 3341 8563 3345 8567
rect 3349 8559 3353 8567
rect 3362 8559 3366 8567
rect 3375 8559 3379 8567
rect 3383 8559 3387 8567
rect 3391 8559 3395 8567
rect 3399 8563 3403 8567
rect 3407 8559 3411 8567
rect 3420 8559 3424 8567
rect 3428 8559 3432 8567
rect 3436 8559 3440 8567
rect 3444 8559 3448 8567
rect 3457 8559 3461 8567
rect 3465 8559 3469 8567
rect 3473 8563 3477 8567
rect 3481 8559 3485 8567
rect 3494 8559 3498 8567
rect 3507 8559 3511 8567
rect 3515 8559 3519 8567
rect 3523 8559 3527 8567
rect 3531 8563 3535 8567
rect 3539 8559 3543 8567
rect 3552 8559 3556 8567
rect 3560 8559 3564 8567
rect 3568 8559 3572 8567
rect 3576 8559 3580 8567
rect 3589 8559 3593 8567
rect 3597 8559 3601 8567
rect 3605 8563 3609 8567
rect 3613 8559 3617 8567
rect 3626 8559 3630 8567
rect 3639 8559 3643 8567
rect 3647 8559 3651 8567
rect 3655 8559 3659 8567
rect 3663 8563 3667 8567
rect 3671 8559 3675 8567
rect 3684 8559 3688 8567
rect 3692 8559 3696 8567
rect 3700 8559 3704 8567
rect 2367 8419 2371 8427
rect 2380 8419 2384 8427
rect 2388 8419 2392 8427
rect 2396 8423 2400 8427
rect 2404 8419 2408 8427
rect 2417 8419 2421 8427
rect 2430 8419 2434 8427
rect 2438 8419 2442 8427
rect 2446 8419 2450 8427
rect 2454 8423 2458 8427
rect 2462 8419 2466 8427
rect 2475 8419 2479 8427
rect 2483 8419 2487 8427
rect 2491 8419 2495 8427
rect 2499 8419 2503 8427
rect 2512 8419 2516 8427
rect 2520 8419 2524 8427
rect 2528 8423 2532 8427
rect 2536 8419 2540 8427
rect 2549 8419 2553 8427
rect 2562 8419 2566 8427
rect 2570 8419 2574 8427
rect 2578 8419 2582 8427
rect 2586 8423 2590 8427
rect 2594 8419 2598 8427
rect 2607 8419 2611 8427
rect 2615 8419 2619 8427
rect 2623 8419 2627 8427
rect 2631 8419 2635 8427
rect 2644 8419 2648 8427
rect 2652 8419 2656 8427
rect 2660 8423 2664 8427
rect 2668 8419 2672 8427
rect 2681 8419 2685 8427
rect 2694 8419 2698 8427
rect 2702 8419 2706 8427
rect 2710 8419 2714 8427
rect 2718 8423 2722 8427
rect 2726 8419 2730 8427
rect 2739 8419 2743 8427
rect 2747 8419 2751 8427
rect 2755 8419 2759 8427
rect 3312 8419 3316 8427
rect 3325 8419 3329 8427
rect 3333 8419 3337 8427
rect 3341 8423 3345 8427
rect 3349 8419 3353 8427
rect 3362 8419 3366 8427
rect 3375 8419 3379 8427
rect 3383 8419 3387 8427
rect 3391 8419 3395 8427
rect 3399 8423 3403 8427
rect 3407 8419 3411 8427
rect 3420 8419 3424 8427
rect 3428 8419 3432 8427
rect 3436 8419 3440 8427
rect 3444 8419 3448 8427
rect 3457 8419 3461 8427
rect 3465 8419 3469 8427
rect 3473 8423 3477 8427
rect 3481 8419 3485 8427
rect 3494 8419 3498 8427
rect 3507 8419 3511 8427
rect 3515 8419 3519 8427
rect 3523 8419 3527 8427
rect 3531 8423 3535 8427
rect 3539 8419 3543 8427
rect 3552 8419 3556 8427
rect 3560 8419 3564 8427
rect 3568 8419 3572 8427
rect 3576 8419 3580 8427
rect 3589 8419 3593 8427
rect 3597 8419 3601 8427
rect 3605 8423 3609 8427
rect 3613 8419 3617 8427
rect 3626 8419 3630 8427
rect 3639 8419 3643 8427
rect 3647 8419 3651 8427
rect 3655 8419 3659 8427
rect 3663 8423 3667 8427
rect 3671 8419 3675 8427
rect 3684 8419 3688 8427
rect 3692 8419 3696 8427
rect 3700 8419 3704 8427
rect 2851 8340 2855 8348
rect 2864 8340 2868 8348
rect 2872 8340 2876 8348
rect 2880 8344 2884 8348
rect 2888 8340 2892 8348
rect 2901 8340 2905 8348
rect 2914 8340 2918 8348
rect 2922 8340 2926 8348
rect 2930 8340 2934 8348
rect 2938 8344 2942 8348
rect 2946 8340 2950 8348
rect 2959 8340 2963 8348
rect 2967 8340 2971 8348
rect 2975 8340 2979 8348
rect 2983 8340 2987 8348
rect 2996 8340 3000 8348
rect 3004 8340 3008 8348
rect 3012 8344 3016 8348
rect 3020 8340 3024 8348
rect 3033 8340 3037 8348
rect 3046 8340 3050 8348
rect 3054 8340 3058 8348
rect 3062 8340 3066 8348
rect 3070 8344 3074 8348
rect 3078 8340 3082 8348
rect 3091 8340 3095 8348
rect 3099 8340 3103 8348
rect 3107 8340 3111 8348
rect 3115 8340 3119 8348
rect 3128 8340 3132 8348
rect 3136 8340 3140 8348
rect 3144 8344 3148 8348
rect 3152 8340 3156 8348
rect 3165 8340 3169 8348
rect 3178 8340 3182 8348
rect 3186 8340 3190 8348
rect 3194 8340 3198 8348
rect 3202 8344 3206 8348
rect 3210 8340 3214 8348
rect 3223 8340 3227 8348
rect 3231 8340 3235 8348
rect 3239 8340 3243 8348
rect 3247 8340 3251 8348
rect 3260 8340 3264 8348
rect 3268 8340 3272 8348
rect 3276 8344 3280 8348
rect 3284 8340 3288 8348
rect 3297 8340 3301 8348
rect 3310 8340 3314 8348
rect 3318 8340 3322 8348
rect 3326 8340 3330 8348
rect 3334 8344 3338 8348
rect 3342 8340 3346 8348
rect 3355 8340 3359 8348
rect 3363 8340 3367 8348
rect 3371 8340 3375 8348
rect 3796 8340 3800 8348
rect 3809 8340 3813 8348
rect 3817 8340 3821 8348
rect 3825 8344 3829 8348
rect 3833 8340 3837 8348
rect 3846 8340 3850 8348
rect 3859 8340 3863 8348
rect 3867 8340 3871 8348
rect 3875 8340 3879 8348
rect 3883 8344 3887 8348
rect 3891 8340 3895 8348
rect 3904 8340 3908 8348
rect 3912 8340 3916 8348
rect 3920 8340 3924 8348
rect 3928 8340 3932 8348
rect 3941 8340 3945 8348
rect 3949 8340 3953 8348
rect 3957 8344 3961 8348
rect 3965 8340 3969 8348
rect 3978 8340 3982 8348
rect 3991 8340 3995 8348
rect 3999 8340 4003 8348
rect 4007 8340 4011 8348
rect 4015 8344 4019 8348
rect 4023 8340 4027 8348
rect 4036 8340 4040 8348
rect 4044 8340 4048 8348
rect 4052 8340 4056 8348
rect 4060 8340 4064 8348
rect 4073 8340 4077 8348
rect 4081 8340 4085 8348
rect 4089 8344 4093 8348
rect 4097 8340 4101 8348
rect 4110 8340 4114 8348
rect 4123 8340 4127 8348
rect 4131 8340 4135 8348
rect 4139 8340 4143 8348
rect 4147 8344 4151 8348
rect 4155 8340 4159 8348
rect 4168 8340 4172 8348
rect 4176 8340 4180 8348
rect 4184 8340 4188 8348
rect 4192 8340 4196 8348
rect 4205 8340 4209 8348
rect 4213 8340 4217 8348
rect 4221 8344 4225 8348
rect 4229 8340 4233 8348
rect 4242 8340 4246 8348
rect 4255 8340 4259 8348
rect 4263 8340 4267 8348
rect 4271 8340 4275 8348
rect 4279 8344 4283 8348
rect 4287 8340 4291 8348
rect 4300 8340 4304 8348
rect 4308 8340 4312 8348
rect 4316 8340 4320 8348
rect 2499 8307 2503 8315
rect 2512 8307 2516 8315
rect 2520 8307 2524 8315
rect 2528 8311 2532 8315
rect 2536 8307 2540 8315
rect 2549 8307 2553 8315
rect 2562 8307 2566 8315
rect 2570 8307 2574 8315
rect 2578 8307 2582 8315
rect 2586 8311 2590 8315
rect 2594 8307 2598 8315
rect 2607 8307 2611 8315
rect 2615 8307 2619 8315
rect 2623 8307 2627 8315
rect 3444 8307 3448 8315
rect 3457 8307 3461 8315
rect 3465 8307 3469 8315
rect 3473 8311 3477 8315
rect 3481 8307 3485 8315
rect 3494 8307 3498 8315
rect 3507 8307 3511 8315
rect 3515 8307 3519 8315
rect 3523 8307 3527 8315
rect 3531 8311 3535 8315
rect 3539 8307 3543 8315
rect 3552 8307 3556 8315
rect 3560 8307 3564 8315
rect 3568 8307 3572 8315
rect 3030 8269 3034 8277
rect 3038 8269 3042 8277
rect 2856 8256 2860 8264
rect 2864 8256 2868 8264
rect 2872 8256 2876 8264
rect 2880 8256 2884 8264
rect 2888 8256 2892 8264
rect 2896 8256 2900 8264
rect 2907 8256 2911 8264
rect 2924 8256 2928 8264
rect 2941 8256 2945 8264
rect 2950 8256 2954 8264
rect 2963 8256 2967 8264
rect 2971 8256 2975 8264
rect 2979 8256 2983 8264
rect 2996 8256 3000 8264
rect 3006 8256 3010 8264
rect 3014 8256 3018 8264
rect 3054 8263 3058 8271
rect 3069 8263 3073 8271
rect 3084 8269 3088 8277
rect 3092 8269 3096 8277
rect 3111 8269 3115 8277
rect 3119 8269 3123 8277
rect 3135 8263 3139 8271
rect 3150 8263 3154 8271
rect 3165 8269 3169 8277
rect 3173 8269 3177 8277
rect 3975 8269 3979 8277
rect 3983 8269 3987 8277
rect 3801 8256 3805 8264
rect 3809 8256 3813 8264
rect 3817 8256 3821 8264
rect 3825 8256 3829 8264
rect 3833 8256 3837 8264
rect 3841 8256 3845 8264
rect 3852 8256 3856 8264
rect 3869 8256 3873 8264
rect 3886 8256 3890 8264
rect 3895 8256 3899 8264
rect 3908 8256 3912 8264
rect 3916 8256 3920 8264
rect 3924 8256 3928 8264
rect 3941 8256 3945 8264
rect 3951 8256 3955 8264
rect 3959 8256 3963 8264
rect 3999 8263 4003 8271
rect 4014 8263 4018 8271
rect 4029 8269 4033 8277
rect 4037 8269 4041 8277
rect 4056 8269 4060 8277
rect 4064 8269 4068 8277
rect 4080 8263 4084 8271
rect 4095 8263 4099 8271
rect 4110 8269 4114 8277
rect 4118 8269 4122 8277
rect 2490 8205 2494 8213
rect 2498 8205 2502 8213
rect 2506 8205 2510 8213
rect 2519 8205 2523 8213
rect 2527 8209 2531 8213
rect 2535 8205 2539 8213
rect 2543 8205 2547 8213
rect 2551 8205 2555 8213
rect 2564 8205 2568 8213
rect 2577 8205 2581 8213
rect 2585 8209 2589 8213
rect 2593 8205 2597 8213
rect 2601 8205 2605 8213
rect 2614 8205 2618 8213
rect 3435 8205 3439 8213
rect 3443 8205 3447 8213
rect 3451 8205 3455 8213
rect 3464 8205 3468 8213
rect 3472 8209 3476 8213
rect 3480 8205 3484 8213
rect 3488 8205 3492 8213
rect 3496 8205 3500 8213
rect 3509 8205 3513 8213
rect 3522 8205 3526 8213
rect 3530 8209 3534 8213
rect 3538 8205 3542 8213
rect 3546 8205 3550 8213
rect 3559 8205 3563 8213
rect 2856 8170 2860 8178
rect 2864 8170 2868 8178
rect 2872 8170 2876 8178
rect 2880 8170 2884 8178
rect 2888 8170 2892 8178
rect 2896 8170 2900 8178
rect 2907 8170 2911 8178
rect 2924 8170 2928 8178
rect 2941 8170 2945 8178
rect 2950 8170 2954 8178
rect 2963 8170 2967 8178
rect 2971 8170 2975 8178
rect 2979 8170 2983 8178
rect 2996 8170 3000 8178
rect 3006 8170 3010 8178
rect 3014 8170 3018 8178
rect 3054 8171 3058 8179
rect 3069 8171 3073 8179
rect 3135 8171 3139 8179
rect 3150 8171 3154 8179
rect 3801 8170 3805 8178
rect 3809 8170 3813 8178
rect 3817 8170 3821 8178
rect 3825 8170 3829 8178
rect 3833 8170 3837 8178
rect 3841 8170 3845 8178
rect 3852 8170 3856 8178
rect 3869 8170 3873 8178
rect 3886 8170 3890 8178
rect 3895 8170 3899 8178
rect 3908 8170 3912 8178
rect 3916 8170 3920 8178
rect 3924 8170 3928 8178
rect 3941 8170 3945 8178
rect 3951 8170 3955 8178
rect 3959 8170 3963 8178
rect 3999 8171 4003 8179
rect 4014 8171 4018 8179
rect 4080 8171 4084 8179
rect 4095 8171 4099 8179
rect 2856 8124 2860 8132
rect 2864 8124 2868 8132
rect 2872 8124 2876 8132
rect 2880 8124 2884 8132
rect 2888 8124 2892 8132
rect 2896 8124 2900 8132
rect 2907 8124 2911 8132
rect 2924 8124 2928 8132
rect 2941 8124 2945 8132
rect 2950 8124 2954 8132
rect 2963 8124 2967 8132
rect 2971 8124 2975 8132
rect 2979 8124 2983 8132
rect 2996 8124 3000 8132
rect 3006 8124 3010 8132
rect 3014 8124 3018 8132
rect 3054 8131 3058 8139
rect 3069 8131 3073 8139
rect 3084 8137 3088 8145
rect 3092 8137 3096 8145
rect 3135 8137 3139 8145
rect 3143 8137 3147 8145
rect 3159 8131 3163 8139
rect 3174 8131 3178 8139
rect 3189 8137 3193 8145
rect 3197 8137 3201 8145
rect 3801 8124 3805 8132
rect 3809 8124 3813 8132
rect 3817 8124 3821 8132
rect 3825 8124 3829 8132
rect 3833 8124 3837 8132
rect 3841 8124 3845 8132
rect 3852 8124 3856 8132
rect 3869 8124 3873 8132
rect 3886 8124 3890 8132
rect 3895 8124 3899 8132
rect 3908 8124 3912 8132
rect 3916 8124 3920 8132
rect 3924 8124 3928 8132
rect 3941 8124 3945 8132
rect 3951 8124 3955 8132
rect 3959 8124 3963 8132
rect 3999 8131 4003 8139
rect 4014 8131 4018 8139
rect 4029 8137 4033 8145
rect 4037 8137 4041 8145
rect 4080 8137 4084 8145
rect 4088 8137 4092 8145
rect 4104 8131 4108 8139
rect 4119 8131 4123 8139
rect 4134 8137 4138 8145
rect 4142 8137 4146 8145
rect 2856 8038 2860 8046
rect 2864 8038 2868 8046
rect 2872 8038 2876 8046
rect 2880 8038 2884 8046
rect 2888 8038 2892 8046
rect 2896 8038 2900 8046
rect 2907 8038 2911 8046
rect 2924 8038 2928 8046
rect 2941 8038 2945 8046
rect 2950 8038 2954 8046
rect 2963 8038 2967 8046
rect 2971 8038 2975 8046
rect 2979 8038 2983 8046
rect 2996 8038 3000 8046
rect 3006 8038 3010 8046
rect 3014 8038 3018 8046
rect 3054 8040 3058 8048
rect 3069 8040 3073 8048
rect 3159 8040 3163 8048
rect 3174 8040 3178 8048
rect 3801 8038 3805 8046
rect 3809 8038 3813 8046
rect 3817 8038 3821 8046
rect 3825 8038 3829 8046
rect 3833 8038 3837 8046
rect 3841 8038 3845 8046
rect 3852 8038 3856 8046
rect 3869 8038 3873 8046
rect 3886 8038 3890 8046
rect 3895 8038 3899 8046
rect 3908 8038 3912 8046
rect 3916 8038 3920 8046
rect 3924 8038 3928 8046
rect 3941 8038 3945 8046
rect 3951 8038 3955 8046
rect 3959 8038 3963 8046
rect 3999 8040 4003 8048
rect 4014 8040 4018 8048
rect 4104 8040 4108 8048
rect 4119 8040 4123 8048
rect 2856 7992 2860 8000
rect 2864 7992 2868 8000
rect 2872 7992 2876 8000
rect 2880 7992 2884 8000
rect 2888 7992 2892 8000
rect 2896 7992 2900 8000
rect 2907 7992 2911 8000
rect 2924 7992 2928 8000
rect 2941 7992 2945 8000
rect 2950 7992 2954 8000
rect 2963 7992 2967 8000
rect 2971 7992 2975 8000
rect 2979 7992 2983 8000
rect 2996 7992 3000 8000
rect 3006 7992 3010 8000
rect 3014 7992 3018 8000
rect 3054 7999 3058 8007
rect 3069 7999 3073 8007
rect 3084 8005 3088 8013
rect 3092 8005 3096 8013
rect 3111 8005 3115 8013
rect 3119 8005 3123 8013
rect 3135 7999 3139 8007
rect 3150 7999 3154 8007
rect 3165 8005 3169 8013
rect 3173 8005 3177 8013
rect 3201 8005 3205 8013
rect 3209 8005 3213 8013
rect 3225 7999 3229 8007
rect 3240 7999 3244 8007
rect 3255 8005 3259 8013
rect 3263 8005 3267 8013
rect 3801 7992 3805 8000
rect 3809 7992 3813 8000
rect 3817 7992 3821 8000
rect 3825 7992 3829 8000
rect 3833 7992 3837 8000
rect 3841 7992 3845 8000
rect 3852 7992 3856 8000
rect 3869 7992 3873 8000
rect 3886 7992 3890 8000
rect 3895 7992 3899 8000
rect 3908 7992 3912 8000
rect 3916 7992 3920 8000
rect 3924 7992 3928 8000
rect 3941 7992 3945 8000
rect 3951 7992 3955 8000
rect 3959 7992 3963 8000
rect 3999 7999 4003 8007
rect 4014 7999 4018 8007
rect 4029 8005 4033 8013
rect 4037 8005 4041 8013
rect 4056 8005 4060 8013
rect 4064 8005 4068 8013
rect 4080 7999 4084 8007
rect 4095 7999 4099 8007
rect 4110 8005 4114 8013
rect 4118 8005 4122 8013
rect 4146 8005 4150 8013
rect 4154 8005 4158 8013
rect 4170 7999 4174 8007
rect 4185 7999 4189 8007
rect 4200 8005 4204 8013
rect 4208 8005 4212 8013
rect 2856 7906 2860 7914
rect 2864 7906 2868 7914
rect 2872 7906 2876 7914
rect 2880 7906 2884 7914
rect 2888 7906 2892 7914
rect 2896 7906 2900 7914
rect 2907 7906 2911 7914
rect 2924 7906 2928 7914
rect 2941 7906 2945 7914
rect 2950 7906 2954 7914
rect 2963 7906 2967 7914
rect 2971 7906 2975 7914
rect 2979 7906 2983 7914
rect 2996 7906 3000 7914
rect 3006 7906 3010 7914
rect 3014 7906 3018 7914
rect 3054 7905 3058 7913
rect 3069 7905 3073 7913
rect 3135 7905 3139 7913
rect 3150 7905 3154 7913
rect 3225 7905 3229 7913
rect 3240 7905 3244 7913
rect 3801 7906 3805 7914
rect 3809 7906 3813 7914
rect 3817 7906 3821 7914
rect 3825 7906 3829 7914
rect 3833 7906 3837 7914
rect 3841 7906 3845 7914
rect 3852 7906 3856 7914
rect 3869 7906 3873 7914
rect 3886 7906 3890 7914
rect 3895 7906 3899 7914
rect 3908 7906 3912 7914
rect 3916 7906 3920 7914
rect 3924 7906 3928 7914
rect 3941 7906 3945 7914
rect 3951 7906 3955 7914
rect 3959 7906 3963 7914
rect 3999 7905 4003 7913
rect 4014 7905 4018 7913
rect 4080 7905 4084 7913
rect 4095 7905 4099 7913
rect 4170 7905 4174 7913
rect 4185 7905 4189 7913
rect 2856 7860 2860 7868
rect 2864 7860 2868 7868
rect 2872 7860 2876 7868
rect 2880 7860 2884 7868
rect 2888 7860 2892 7868
rect 2896 7860 2900 7868
rect 2907 7860 2911 7868
rect 2924 7860 2928 7868
rect 2941 7860 2945 7868
rect 2950 7860 2954 7868
rect 2963 7860 2967 7868
rect 2971 7860 2975 7868
rect 2979 7860 2983 7868
rect 2996 7860 3000 7868
rect 3006 7860 3010 7868
rect 3014 7860 3018 7868
rect 3054 7867 3058 7875
rect 3069 7867 3073 7875
rect 3084 7873 3088 7881
rect 3092 7873 3096 7881
rect 3801 7860 3805 7868
rect 3809 7860 3813 7868
rect 3817 7860 3821 7868
rect 3825 7860 3829 7868
rect 3833 7860 3837 7868
rect 3841 7860 3845 7868
rect 3852 7860 3856 7868
rect 3869 7860 3873 7868
rect 3886 7860 3890 7868
rect 3895 7860 3899 7868
rect 3908 7860 3912 7868
rect 3916 7860 3920 7868
rect 3924 7860 3928 7868
rect 3941 7860 3945 7868
rect 3951 7860 3955 7868
rect 3959 7860 3963 7868
rect 3999 7867 4003 7875
rect 4014 7867 4018 7875
rect 4029 7873 4033 7881
rect 4037 7873 4041 7881
rect 2367 7805 2371 7813
rect 2380 7805 2384 7813
rect 2388 7805 2392 7813
rect 2396 7809 2400 7813
rect 2404 7805 2408 7813
rect 2417 7805 2421 7813
rect 2430 7805 2434 7813
rect 2438 7805 2442 7813
rect 2446 7805 2450 7813
rect 2454 7809 2458 7813
rect 2462 7805 2466 7813
rect 2475 7805 2479 7813
rect 2483 7805 2487 7813
rect 2491 7805 2495 7813
rect 2499 7805 2503 7813
rect 2512 7805 2516 7813
rect 2520 7805 2524 7813
rect 2528 7809 2532 7813
rect 2536 7805 2540 7813
rect 2549 7805 2553 7813
rect 2562 7805 2566 7813
rect 2570 7805 2574 7813
rect 2578 7805 2582 7813
rect 2586 7809 2590 7813
rect 2594 7805 2598 7813
rect 2607 7805 2611 7813
rect 2615 7805 2619 7813
rect 2623 7805 2627 7813
rect 2631 7805 2635 7813
rect 2644 7805 2648 7813
rect 2652 7805 2656 7813
rect 2660 7809 2664 7813
rect 2668 7805 2672 7813
rect 2681 7805 2685 7813
rect 2694 7805 2698 7813
rect 2702 7805 2706 7813
rect 2710 7805 2714 7813
rect 2718 7809 2722 7813
rect 2726 7805 2730 7813
rect 2739 7805 2743 7813
rect 2747 7805 2751 7813
rect 2755 7805 2759 7813
rect 3312 7805 3316 7813
rect 3325 7805 3329 7813
rect 3333 7805 3337 7813
rect 3341 7809 3345 7813
rect 3349 7805 3353 7813
rect 3362 7805 3366 7813
rect 3375 7805 3379 7813
rect 3383 7805 3387 7813
rect 3391 7805 3395 7813
rect 3399 7809 3403 7813
rect 3407 7805 3411 7813
rect 3420 7805 3424 7813
rect 3428 7805 3432 7813
rect 3436 7805 3440 7813
rect 3444 7805 3448 7813
rect 3457 7805 3461 7813
rect 3465 7805 3469 7813
rect 3473 7809 3477 7813
rect 3481 7805 3485 7813
rect 3494 7805 3498 7813
rect 3507 7805 3511 7813
rect 3515 7805 3519 7813
rect 3523 7805 3527 7813
rect 3531 7809 3535 7813
rect 3539 7805 3543 7813
rect 3552 7805 3556 7813
rect 3560 7805 3564 7813
rect 3568 7805 3572 7813
rect 3576 7805 3580 7813
rect 3589 7805 3593 7813
rect 3597 7805 3601 7813
rect 3605 7809 3609 7813
rect 3613 7805 3617 7813
rect 3626 7805 3630 7813
rect 3639 7805 3643 7813
rect 3647 7805 3651 7813
rect 3655 7805 3659 7813
rect 3663 7809 3667 7813
rect 3671 7805 3675 7813
rect 3684 7805 3688 7813
rect 3692 7805 3696 7813
rect 3700 7805 3704 7813
rect 2856 7774 2860 7782
rect 2864 7774 2868 7782
rect 2872 7774 2876 7782
rect 2880 7774 2884 7782
rect 2888 7774 2892 7782
rect 2896 7774 2900 7782
rect 2907 7774 2911 7782
rect 2924 7774 2928 7782
rect 2941 7774 2945 7782
rect 2950 7774 2954 7782
rect 2963 7774 2967 7782
rect 2971 7774 2975 7782
rect 2979 7774 2983 7782
rect 2996 7774 3000 7782
rect 3006 7774 3010 7782
rect 3014 7774 3018 7782
rect 3054 7769 3058 7777
rect 3069 7769 3073 7777
rect 3090 7774 3094 7782
rect 3098 7774 3102 7782
rect 3108 7774 3112 7782
rect 3116 7774 3120 7782
rect 3125 7774 3129 7782
rect 3133 7774 3137 7782
rect 3141 7774 3145 7782
rect 3149 7774 3153 7782
rect 3157 7774 3161 7782
rect 3168 7774 3172 7782
rect 3185 7774 3189 7782
rect 3202 7774 3206 7782
rect 3211 7774 3215 7782
rect 3224 7774 3228 7782
rect 3232 7774 3236 7782
rect 3240 7774 3244 7782
rect 3257 7774 3261 7782
rect 3267 7774 3271 7782
rect 3275 7774 3279 7782
rect 3801 7774 3805 7782
rect 3809 7774 3813 7782
rect 3817 7774 3821 7782
rect 3825 7774 3829 7782
rect 3833 7774 3837 7782
rect 3841 7774 3845 7782
rect 3852 7774 3856 7782
rect 3869 7774 3873 7782
rect 3886 7774 3890 7782
rect 3895 7774 3899 7782
rect 3908 7774 3912 7782
rect 3916 7774 3920 7782
rect 3924 7774 3928 7782
rect 3941 7774 3945 7782
rect 3951 7774 3955 7782
rect 3959 7774 3963 7782
rect 3999 7769 4003 7777
rect 4014 7769 4018 7777
rect 4035 7774 4039 7782
rect 4043 7774 4047 7782
rect 4053 7774 4057 7782
rect 4061 7774 4065 7782
rect 4070 7774 4074 7782
rect 4078 7774 4082 7782
rect 4086 7774 4090 7782
rect 4094 7774 4098 7782
rect 4102 7774 4106 7782
rect 4113 7774 4117 7782
rect 4130 7774 4134 7782
rect 4147 7774 4151 7782
rect 4156 7774 4160 7782
rect 4169 7774 4173 7782
rect 4177 7774 4181 7782
rect 4185 7774 4189 7782
rect 4202 7774 4206 7782
rect 4212 7774 4216 7782
rect 4220 7774 4224 7782
rect 3150 7693 3154 7701
rect 3163 7693 3167 7701
rect 3171 7693 3175 7701
rect 3179 7697 3183 7701
rect 3187 7693 3191 7701
rect 3200 7693 3204 7701
rect 3213 7693 3217 7701
rect 3221 7693 3225 7701
rect 3229 7693 3233 7701
rect 3237 7697 3241 7701
rect 3245 7693 3249 7701
rect 3258 7693 3262 7701
rect 3266 7693 3270 7701
rect 3274 7693 3278 7701
rect 4095 7693 4099 7701
rect 4108 7693 4112 7701
rect 4116 7693 4120 7701
rect 4124 7697 4128 7701
rect 4132 7693 4136 7701
rect 4145 7693 4149 7701
rect 4158 7693 4162 7701
rect 4166 7693 4170 7701
rect 4174 7693 4178 7701
rect 4182 7697 4186 7701
rect 4190 7693 4194 7701
rect 4203 7693 4207 7701
rect 4211 7693 4215 7701
rect 4219 7693 4223 7701
rect 2367 7663 2371 7671
rect 2380 7663 2384 7671
rect 2388 7663 2392 7671
rect 2396 7667 2400 7671
rect 2404 7663 2408 7671
rect 2417 7663 2421 7671
rect 2430 7663 2434 7671
rect 2438 7663 2442 7671
rect 2446 7663 2450 7671
rect 2454 7667 2458 7671
rect 2462 7663 2466 7671
rect 2475 7663 2479 7671
rect 2483 7663 2487 7671
rect 2491 7663 2495 7671
rect 2499 7663 2503 7671
rect 2512 7663 2516 7671
rect 2520 7663 2524 7671
rect 2528 7667 2532 7671
rect 2536 7663 2540 7671
rect 2549 7663 2553 7671
rect 2562 7663 2566 7671
rect 2570 7663 2574 7671
rect 2578 7663 2582 7671
rect 2586 7667 2590 7671
rect 2594 7663 2598 7671
rect 2607 7663 2611 7671
rect 2615 7663 2619 7671
rect 2623 7663 2627 7671
rect 2631 7663 2635 7671
rect 2644 7663 2648 7671
rect 2652 7663 2656 7671
rect 2660 7667 2664 7671
rect 2668 7663 2672 7671
rect 2681 7663 2685 7671
rect 2694 7663 2698 7671
rect 2702 7663 2706 7671
rect 2710 7663 2714 7671
rect 2718 7667 2722 7671
rect 2726 7663 2730 7671
rect 2739 7663 2743 7671
rect 2747 7663 2751 7671
rect 2755 7663 2759 7671
rect 3312 7663 3316 7671
rect 3325 7663 3329 7671
rect 3333 7663 3337 7671
rect 3341 7667 3345 7671
rect 3349 7663 3353 7671
rect 3362 7663 3366 7671
rect 3375 7663 3379 7671
rect 3383 7663 3387 7671
rect 3391 7663 3395 7671
rect 3399 7667 3403 7671
rect 3407 7663 3411 7671
rect 3420 7663 3424 7671
rect 3428 7663 3432 7671
rect 3436 7663 3440 7671
rect 3444 7663 3448 7671
rect 3457 7663 3461 7671
rect 3465 7663 3469 7671
rect 3473 7667 3477 7671
rect 3481 7663 3485 7671
rect 3494 7663 3498 7671
rect 3507 7663 3511 7671
rect 3515 7663 3519 7671
rect 3523 7663 3527 7671
rect 3531 7667 3535 7671
rect 3539 7663 3543 7671
rect 3552 7663 3556 7671
rect 3560 7663 3564 7671
rect 3568 7663 3572 7671
rect 3576 7663 3580 7671
rect 3589 7663 3593 7671
rect 3597 7663 3601 7671
rect 3605 7667 3609 7671
rect 3613 7663 3617 7671
rect 3626 7663 3630 7671
rect 3639 7663 3643 7671
rect 3647 7663 3651 7671
rect 3655 7663 3659 7671
rect 3663 7667 3667 7671
rect 3671 7663 3675 7671
rect 3684 7663 3688 7671
rect 3692 7663 3696 7671
rect 3700 7663 3704 7671
rect 3150 7607 3154 7615
rect 3163 7607 3167 7615
rect 3171 7607 3175 7615
rect 3179 7611 3183 7615
rect 3187 7607 3191 7615
rect 3200 7607 3204 7615
rect 3213 7607 3217 7615
rect 3221 7607 3225 7615
rect 3229 7607 3233 7615
rect 3237 7611 3241 7615
rect 3245 7607 3249 7615
rect 3258 7607 3262 7615
rect 3266 7607 3270 7615
rect 3274 7607 3278 7615
rect 4095 7607 4099 7615
rect 4108 7607 4112 7615
rect 4116 7607 4120 7615
rect 4124 7611 4128 7615
rect 4132 7607 4136 7615
rect 4145 7607 4149 7615
rect 4158 7607 4162 7615
rect 4166 7607 4170 7615
rect 4174 7607 4178 7615
rect 4182 7611 4186 7615
rect 4190 7607 4194 7615
rect 4203 7607 4207 7615
rect 4211 7607 4215 7615
rect 4219 7607 4223 7615
rect 2367 7577 2371 7585
rect 2380 7577 2384 7585
rect 2388 7577 2392 7585
rect 2396 7581 2400 7585
rect 2404 7577 2408 7585
rect 2417 7577 2421 7585
rect 2430 7577 2434 7585
rect 2438 7577 2442 7585
rect 2446 7577 2450 7585
rect 2454 7581 2458 7585
rect 2462 7577 2466 7585
rect 2475 7577 2479 7585
rect 2483 7577 2487 7585
rect 2491 7577 2495 7585
rect 2499 7577 2503 7585
rect 2512 7577 2516 7585
rect 2520 7577 2524 7585
rect 2528 7581 2532 7585
rect 2536 7577 2540 7585
rect 2549 7577 2553 7585
rect 2562 7577 2566 7585
rect 2570 7577 2574 7585
rect 2578 7577 2582 7585
rect 2586 7581 2590 7585
rect 2594 7577 2598 7585
rect 2607 7577 2611 7585
rect 2615 7577 2619 7585
rect 2623 7577 2627 7585
rect 2631 7577 2635 7585
rect 2644 7577 2648 7585
rect 2652 7577 2656 7585
rect 2660 7581 2664 7585
rect 2668 7577 2672 7585
rect 2681 7577 2685 7585
rect 2694 7577 2698 7585
rect 2702 7577 2706 7585
rect 2710 7577 2714 7585
rect 2718 7581 2722 7585
rect 2726 7577 2730 7585
rect 2739 7577 2743 7585
rect 2747 7577 2751 7585
rect 2755 7577 2759 7585
rect 3312 7577 3316 7585
rect 3325 7577 3329 7585
rect 3333 7577 3337 7585
rect 3341 7581 3345 7585
rect 3349 7577 3353 7585
rect 3362 7577 3366 7585
rect 3375 7577 3379 7585
rect 3383 7577 3387 7585
rect 3391 7577 3395 7585
rect 3399 7581 3403 7585
rect 3407 7577 3411 7585
rect 3420 7577 3424 7585
rect 3428 7577 3432 7585
rect 3436 7577 3440 7585
rect 3444 7577 3448 7585
rect 3457 7577 3461 7585
rect 3465 7577 3469 7585
rect 3473 7581 3477 7585
rect 3481 7577 3485 7585
rect 3494 7577 3498 7585
rect 3507 7577 3511 7585
rect 3515 7577 3519 7585
rect 3523 7577 3527 7585
rect 3531 7581 3535 7585
rect 3539 7577 3543 7585
rect 3552 7577 3556 7585
rect 3560 7577 3564 7585
rect 3568 7577 3572 7585
rect 3576 7577 3580 7585
rect 3589 7577 3593 7585
rect 3597 7577 3601 7585
rect 3605 7581 3609 7585
rect 3613 7577 3617 7585
rect 3626 7577 3630 7585
rect 3639 7577 3643 7585
rect 3647 7577 3651 7585
rect 3655 7577 3659 7585
rect 3663 7581 3667 7585
rect 3671 7577 3675 7585
rect 3684 7577 3688 7585
rect 3692 7577 3696 7585
rect 3700 7577 3704 7585
rect 2367 7437 2371 7445
rect 2380 7437 2384 7445
rect 2388 7437 2392 7445
rect 2396 7441 2400 7445
rect 2404 7437 2408 7445
rect 2417 7437 2421 7445
rect 2430 7437 2434 7445
rect 2438 7437 2442 7445
rect 2446 7437 2450 7445
rect 2454 7441 2458 7445
rect 2462 7437 2466 7445
rect 2475 7437 2479 7445
rect 2483 7437 2487 7445
rect 2491 7437 2495 7445
rect 2499 7437 2503 7445
rect 2512 7437 2516 7445
rect 2520 7437 2524 7445
rect 2528 7441 2532 7445
rect 2536 7437 2540 7445
rect 2549 7437 2553 7445
rect 2562 7437 2566 7445
rect 2570 7437 2574 7445
rect 2578 7437 2582 7445
rect 2586 7441 2590 7445
rect 2594 7437 2598 7445
rect 2607 7437 2611 7445
rect 2615 7437 2619 7445
rect 2623 7437 2627 7445
rect 2631 7437 2635 7445
rect 2644 7437 2648 7445
rect 2652 7437 2656 7445
rect 2660 7441 2664 7445
rect 2668 7437 2672 7445
rect 2681 7437 2685 7445
rect 2694 7437 2698 7445
rect 2702 7437 2706 7445
rect 2710 7437 2714 7445
rect 2718 7441 2722 7445
rect 2726 7437 2730 7445
rect 2739 7437 2743 7445
rect 2747 7437 2751 7445
rect 2755 7437 2759 7445
rect 3312 7437 3316 7445
rect 3325 7437 3329 7445
rect 3333 7437 3337 7445
rect 3341 7441 3345 7445
rect 3349 7437 3353 7445
rect 3362 7437 3366 7445
rect 3375 7437 3379 7445
rect 3383 7437 3387 7445
rect 3391 7437 3395 7445
rect 3399 7441 3403 7445
rect 3407 7437 3411 7445
rect 3420 7437 3424 7445
rect 3428 7437 3432 7445
rect 3436 7437 3440 7445
rect 3444 7437 3448 7445
rect 3457 7437 3461 7445
rect 3465 7437 3469 7445
rect 3473 7441 3477 7445
rect 3481 7437 3485 7445
rect 3494 7437 3498 7445
rect 3507 7437 3511 7445
rect 3515 7437 3519 7445
rect 3523 7437 3527 7445
rect 3531 7441 3535 7445
rect 3539 7437 3543 7445
rect 3552 7437 3556 7445
rect 3560 7437 3564 7445
rect 3568 7437 3572 7445
rect 3576 7437 3580 7445
rect 3589 7437 3593 7445
rect 3597 7437 3601 7445
rect 3605 7441 3609 7445
rect 3613 7437 3617 7445
rect 3626 7437 3630 7445
rect 3639 7437 3643 7445
rect 3647 7437 3651 7445
rect 3655 7437 3659 7445
rect 3663 7441 3667 7445
rect 3671 7437 3675 7445
rect 3684 7437 3688 7445
rect 3692 7437 3696 7445
rect 3700 7437 3704 7445
rect 1468 6869 1472 6877
rect 1476 6869 1480 6877
rect 1484 6869 1488 6877
rect 1497 6869 1501 6877
rect 1505 6869 1509 6873
rect 1513 6869 1517 6877
rect 1521 6869 1525 6877
rect 1529 6869 1533 6877
rect 1542 6869 1546 6877
rect 1555 6869 1559 6877
rect 1563 6869 1567 6873
rect 1571 6869 1575 6877
rect 1579 6869 1583 6877
rect 1592 6869 1596 6877
rect 1600 6869 1604 6877
rect 1608 6869 1612 6877
rect 1616 6869 1620 6877
rect 1629 6869 1633 6877
rect 1637 6869 1641 6873
rect 1645 6869 1649 6877
rect 1653 6869 1657 6877
rect 1661 6869 1665 6877
rect 1674 6869 1678 6877
rect 1687 6869 1691 6877
rect 1695 6869 1699 6873
rect 1703 6869 1707 6877
rect 1711 6869 1715 6877
rect 1724 6869 1728 6877
rect 1732 6869 1736 6877
rect 1740 6869 1744 6877
rect 1748 6869 1752 6877
rect 1761 6869 1765 6877
rect 1769 6869 1773 6873
rect 1777 6869 1781 6877
rect 1785 6869 1789 6877
rect 1793 6869 1797 6877
rect 1806 6869 1810 6877
rect 1819 6869 1823 6877
rect 1827 6869 1831 6873
rect 1835 6869 1839 6877
rect 1843 6869 1847 6877
rect 1856 6869 1860 6877
rect 2413 6869 2417 6877
rect 2421 6869 2425 6877
rect 2429 6869 2433 6877
rect 2442 6869 2446 6877
rect 2450 6869 2454 6873
rect 2458 6869 2462 6877
rect 2466 6869 2470 6877
rect 2474 6869 2478 6877
rect 2487 6869 2491 6877
rect 2500 6869 2504 6877
rect 2508 6869 2512 6873
rect 2516 6869 2520 6877
rect 2524 6869 2528 6877
rect 2537 6869 2541 6877
rect 2545 6869 2549 6877
rect 2553 6869 2557 6877
rect 2561 6869 2565 6877
rect 2574 6869 2578 6877
rect 2582 6869 2586 6873
rect 2590 6869 2594 6877
rect 2598 6869 2602 6877
rect 2606 6869 2610 6877
rect 2619 6869 2623 6877
rect 2632 6869 2636 6877
rect 2640 6869 2644 6873
rect 2648 6869 2652 6877
rect 2656 6869 2660 6877
rect 2669 6869 2673 6877
rect 2677 6869 2681 6877
rect 2685 6869 2689 6877
rect 2693 6869 2697 6877
rect 2706 6869 2710 6877
rect 2714 6869 2718 6873
rect 2722 6869 2726 6877
rect 2730 6869 2734 6877
rect 2738 6869 2742 6877
rect 2751 6869 2755 6877
rect 2764 6869 2768 6877
rect 2772 6869 2776 6873
rect 2780 6869 2784 6877
rect 2788 6869 2792 6877
rect 2801 6869 2805 6877
rect 1468 6729 1472 6737
rect 1476 6729 1480 6737
rect 1484 6729 1488 6737
rect 1497 6729 1501 6737
rect 1505 6729 1509 6733
rect 1513 6729 1517 6737
rect 1521 6729 1525 6737
rect 1529 6729 1533 6737
rect 1542 6729 1546 6737
rect 1555 6729 1559 6737
rect 1563 6729 1567 6733
rect 1571 6729 1575 6737
rect 1579 6729 1583 6737
rect 1592 6729 1596 6737
rect 1600 6729 1604 6737
rect 1608 6729 1612 6737
rect 1616 6729 1620 6737
rect 1629 6729 1633 6737
rect 1637 6729 1641 6733
rect 1645 6729 1649 6737
rect 1653 6729 1657 6737
rect 1661 6729 1665 6737
rect 1674 6729 1678 6737
rect 1687 6729 1691 6737
rect 1695 6729 1699 6733
rect 1703 6729 1707 6737
rect 1711 6729 1715 6737
rect 1724 6729 1728 6737
rect 1732 6729 1736 6737
rect 1740 6729 1744 6737
rect 1748 6729 1752 6737
rect 1761 6729 1765 6737
rect 1769 6729 1773 6733
rect 1777 6729 1781 6737
rect 1785 6729 1789 6737
rect 1793 6729 1797 6737
rect 1806 6729 1810 6737
rect 1819 6729 1823 6737
rect 1827 6729 1831 6733
rect 1835 6729 1839 6737
rect 1843 6729 1847 6737
rect 1856 6729 1860 6737
rect 2413 6729 2417 6737
rect 2421 6729 2425 6737
rect 2429 6729 2433 6737
rect 2442 6729 2446 6737
rect 2450 6729 2454 6733
rect 2458 6729 2462 6737
rect 2466 6729 2470 6737
rect 2474 6729 2478 6737
rect 2487 6729 2491 6737
rect 2500 6729 2504 6737
rect 2508 6729 2512 6733
rect 2516 6729 2520 6737
rect 2524 6729 2528 6737
rect 2537 6729 2541 6737
rect 2545 6729 2549 6737
rect 2553 6729 2557 6737
rect 2561 6729 2565 6737
rect 2574 6729 2578 6737
rect 2582 6729 2586 6733
rect 2590 6729 2594 6737
rect 2598 6729 2602 6737
rect 2606 6729 2610 6737
rect 2619 6729 2623 6737
rect 2632 6729 2636 6737
rect 2640 6729 2644 6733
rect 2648 6729 2652 6737
rect 2656 6729 2660 6737
rect 2669 6729 2673 6737
rect 2677 6729 2681 6737
rect 2685 6729 2689 6737
rect 2693 6729 2697 6737
rect 2706 6729 2710 6737
rect 2714 6729 2718 6733
rect 2722 6729 2726 6737
rect 2730 6729 2734 6737
rect 2738 6729 2742 6737
rect 2751 6729 2755 6737
rect 2764 6729 2768 6737
rect 2772 6729 2776 6733
rect 2780 6729 2784 6737
rect 2788 6729 2792 6737
rect 2801 6729 2805 6737
rect 949 6699 953 6707
rect 957 6699 961 6707
rect 965 6699 969 6707
rect 978 6699 982 6707
rect 986 6699 990 6703
rect 994 6699 998 6707
rect 1002 6699 1006 6707
rect 1010 6699 1014 6707
rect 1023 6699 1027 6707
rect 1036 6699 1040 6707
rect 1044 6699 1048 6703
rect 1052 6699 1056 6707
rect 1060 6699 1064 6707
rect 1073 6699 1077 6707
rect 1894 6699 1898 6707
rect 1902 6699 1906 6707
rect 1910 6699 1914 6707
rect 1923 6699 1927 6707
rect 1931 6699 1935 6703
rect 1939 6699 1943 6707
rect 1947 6699 1951 6707
rect 1955 6699 1959 6707
rect 1968 6699 1972 6707
rect 1981 6699 1985 6707
rect 1989 6699 1993 6703
rect 1997 6699 2001 6707
rect 2005 6699 2009 6707
rect 2018 6699 2022 6707
rect 1468 6643 1472 6651
rect 1476 6643 1480 6651
rect 1484 6643 1488 6651
rect 1497 6643 1501 6651
rect 1505 6643 1509 6647
rect 1513 6643 1517 6651
rect 1521 6643 1525 6651
rect 1529 6643 1533 6651
rect 1542 6643 1546 6651
rect 1555 6643 1559 6651
rect 1563 6643 1567 6647
rect 1571 6643 1575 6651
rect 1579 6643 1583 6651
rect 1592 6643 1596 6651
rect 1600 6643 1604 6651
rect 1608 6643 1612 6651
rect 1616 6643 1620 6651
rect 1629 6643 1633 6651
rect 1637 6643 1641 6647
rect 1645 6643 1649 6651
rect 1653 6643 1657 6651
rect 1661 6643 1665 6651
rect 1674 6643 1678 6651
rect 1687 6643 1691 6651
rect 1695 6643 1699 6647
rect 1703 6643 1707 6651
rect 1711 6643 1715 6651
rect 1724 6643 1728 6651
rect 1732 6643 1736 6651
rect 1740 6643 1744 6651
rect 1748 6643 1752 6651
rect 1761 6643 1765 6651
rect 1769 6643 1773 6647
rect 1777 6643 1781 6651
rect 1785 6643 1789 6651
rect 1793 6643 1797 6651
rect 1806 6643 1810 6651
rect 1819 6643 1823 6651
rect 1827 6643 1831 6647
rect 1835 6643 1839 6651
rect 1843 6643 1847 6651
rect 1856 6643 1860 6651
rect 2413 6643 2417 6651
rect 2421 6643 2425 6651
rect 2429 6643 2433 6651
rect 2442 6643 2446 6651
rect 2450 6643 2454 6647
rect 2458 6643 2462 6651
rect 2466 6643 2470 6651
rect 2474 6643 2478 6651
rect 2487 6643 2491 6651
rect 2500 6643 2504 6651
rect 2508 6643 2512 6647
rect 2516 6643 2520 6651
rect 2524 6643 2528 6651
rect 2537 6643 2541 6651
rect 2545 6643 2549 6651
rect 2553 6643 2557 6651
rect 2561 6643 2565 6651
rect 2574 6643 2578 6651
rect 2582 6643 2586 6647
rect 2590 6643 2594 6651
rect 2598 6643 2602 6651
rect 2606 6643 2610 6651
rect 2619 6643 2623 6651
rect 2632 6643 2636 6651
rect 2640 6643 2644 6647
rect 2648 6643 2652 6651
rect 2656 6643 2660 6651
rect 2669 6643 2673 6651
rect 2677 6643 2681 6651
rect 2685 6643 2689 6651
rect 2693 6643 2697 6651
rect 2706 6643 2710 6651
rect 2714 6643 2718 6647
rect 2722 6643 2726 6651
rect 2730 6643 2734 6651
rect 2738 6643 2742 6651
rect 2751 6643 2755 6651
rect 2764 6643 2768 6651
rect 2772 6643 2776 6647
rect 2780 6643 2784 6651
rect 2788 6643 2792 6651
rect 2801 6643 2805 6651
rect 949 6613 953 6621
rect 957 6613 961 6621
rect 965 6613 969 6621
rect 978 6613 982 6621
rect 986 6613 990 6617
rect 994 6613 998 6621
rect 1002 6613 1006 6621
rect 1010 6613 1014 6621
rect 1023 6613 1027 6621
rect 1036 6613 1040 6621
rect 1044 6613 1048 6617
rect 1052 6613 1056 6621
rect 1060 6613 1064 6621
rect 1073 6613 1077 6621
rect 1894 6613 1898 6621
rect 1902 6613 1906 6621
rect 1910 6613 1914 6621
rect 1923 6613 1927 6621
rect 1931 6613 1935 6617
rect 1939 6613 1943 6621
rect 1947 6613 1951 6621
rect 1955 6613 1959 6621
rect 1968 6613 1972 6621
rect 1981 6613 1985 6621
rect 1989 6613 1993 6617
rect 1997 6613 2001 6621
rect 2005 6613 2009 6621
rect 2018 6613 2022 6621
rect 948 6532 952 6540
rect 956 6532 960 6540
rect 966 6532 970 6540
rect 983 6532 987 6540
rect 991 6532 995 6540
rect 999 6532 1003 6540
rect 1012 6532 1016 6540
rect 1021 6532 1025 6540
rect 1038 6532 1042 6540
rect 1055 6532 1059 6540
rect 1066 6532 1070 6540
rect 1074 6532 1078 6540
rect 1082 6532 1086 6540
rect 1090 6532 1094 6540
rect 1098 6532 1102 6540
rect 1107 6532 1111 6540
rect 1115 6532 1119 6540
rect 1125 6532 1129 6540
rect 1133 6532 1137 6540
rect 1154 6537 1158 6545
rect 1169 6537 1173 6545
rect 1209 6532 1213 6540
rect 1217 6532 1221 6540
rect 1227 6532 1231 6540
rect 1244 6532 1248 6540
rect 1252 6532 1256 6540
rect 1260 6532 1264 6540
rect 1273 6532 1277 6540
rect 1282 6532 1286 6540
rect 1299 6532 1303 6540
rect 1316 6532 1320 6540
rect 1327 6532 1331 6540
rect 1335 6532 1339 6540
rect 1343 6532 1347 6540
rect 1351 6532 1355 6540
rect 1359 6532 1363 6540
rect 1367 6532 1371 6540
rect 1893 6532 1897 6540
rect 1901 6532 1905 6540
rect 1911 6532 1915 6540
rect 1928 6532 1932 6540
rect 1936 6532 1940 6540
rect 1944 6532 1948 6540
rect 1957 6532 1961 6540
rect 1966 6532 1970 6540
rect 1983 6532 1987 6540
rect 2000 6532 2004 6540
rect 2011 6532 2015 6540
rect 2019 6532 2023 6540
rect 2027 6532 2031 6540
rect 2035 6532 2039 6540
rect 2043 6532 2047 6540
rect 2052 6532 2056 6540
rect 2060 6532 2064 6540
rect 2070 6532 2074 6540
rect 2078 6532 2082 6540
rect 2099 6537 2103 6545
rect 2114 6537 2118 6545
rect 2154 6532 2158 6540
rect 2162 6532 2166 6540
rect 2172 6532 2176 6540
rect 2189 6532 2193 6540
rect 2197 6532 2201 6540
rect 2205 6532 2209 6540
rect 2218 6532 2222 6540
rect 2227 6532 2231 6540
rect 2244 6532 2248 6540
rect 2261 6532 2265 6540
rect 2272 6532 2276 6540
rect 2280 6532 2284 6540
rect 2288 6532 2292 6540
rect 2296 6532 2300 6540
rect 2304 6532 2308 6540
rect 2312 6532 2316 6540
rect 1468 6501 1472 6509
rect 1476 6501 1480 6509
rect 1484 6501 1488 6509
rect 1497 6501 1501 6509
rect 1505 6501 1509 6505
rect 1513 6501 1517 6509
rect 1521 6501 1525 6509
rect 1529 6501 1533 6509
rect 1542 6501 1546 6509
rect 1555 6501 1559 6509
rect 1563 6501 1567 6505
rect 1571 6501 1575 6509
rect 1579 6501 1583 6509
rect 1592 6501 1596 6509
rect 1600 6501 1604 6509
rect 1608 6501 1612 6509
rect 1616 6501 1620 6509
rect 1629 6501 1633 6509
rect 1637 6501 1641 6505
rect 1645 6501 1649 6509
rect 1653 6501 1657 6509
rect 1661 6501 1665 6509
rect 1674 6501 1678 6509
rect 1687 6501 1691 6509
rect 1695 6501 1699 6505
rect 1703 6501 1707 6509
rect 1711 6501 1715 6509
rect 1724 6501 1728 6509
rect 1732 6501 1736 6509
rect 1740 6501 1744 6509
rect 1748 6501 1752 6509
rect 1761 6501 1765 6509
rect 1769 6501 1773 6505
rect 1777 6501 1781 6509
rect 1785 6501 1789 6509
rect 1793 6501 1797 6509
rect 1806 6501 1810 6509
rect 1819 6501 1823 6509
rect 1827 6501 1831 6505
rect 1835 6501 1839 6509
rect 1843 6501 1847 6509
rect 1856 6501 1860 6509
rect 2413 6501 2417 6509
rect 2421 6501 2425 6509
rect 2429 6501 2433 6509
rect 2442 6501 2446 6509
rect 2450 6501 2454 6505
rect 2458 6501 2462 6509
rect 2466 6501 2470 6509
rect 2474 6501 2478 6509
rect 2487 6501 2491 6509
rect 2500 6501 2504 6509
rect 2508 6501 2512 6505
rect 2516 6501 2520 6509
rect 2524 6501 2528 6509
rect 2537 6501 2541 6509
rect 2545 6501 2549 6509
rect 2553 6501 2557 6509
rect 2561 6501 2565 6509
rect 2574 6501 2578 6509
rect 2582 6501 2586 6505
rect 2590 6501 2594 6509
rect 2598 6501 2602 6509
rect 2606 6501 2610 6509
rect 2619 6501 2623 6509
rect 2632 6501 2636 6509
rect 2640 6501 2644 6505
rect 2648 6501 2652 6509
rect 2656 6501 2660 6509
rect 2669 6501 2673 6509
rect 2677 6501 2681 6509
rect 2685 6501 2689 6509
rect 2693 6501 2697 6509
rect 2706 6501 2710 6509
rect 2714 6501 2718 6505
rect 2722 6501 2726 6509
rect 2730 6501 2734 6509
rect 2738 6501 2742 6509
rect 2751 6501 2755 6509
rect 2764 6501 2768 6509
rect 2772 6501 2776 6505
rect 2780 6501 2784 6509
rect 2788 6501 2792 6509
rect 2801 6501 2805 6509
rect 1131 6433 1135 6441
rect 1139 6433 1143 6441
rect 1154 6439 1158 6447
rect 1169 6439 1173 6447
rect 1209 6446 1213 6454
rect 1217 6446 1221 6454
rect 1227 6446 1231 6454
rect 1244 6446 1248 6454
rect 1252 6446 1256 6454
rect 1260 6446 1264 6454
rect 1273 6446 1277 6454
rect 1282 6446 1286 6454
rect 1299 6446 1303 6454
rect 1316 6446 1320 6454
rect 1327 6446 1331 6454
rect 1335 6446 1339 6454
rect 1343 6446 1347 6454
rect 1351 6446 1355 6454
rect 1359 6446 1363 6454
rect 1367 6446 1371 6454
rect 2076 6433 2080 6441
rect 2084 6433 2088 6441
rect 2099 6439 2103 6447
rect 2114 6439 2118 6447
rect 2154 6446 2158 6454
rect 2162 6446 2166 6454
rect 2172 6446 2176 6454
rect 2189 6446 2193 6454
rect 2197 6446 2201 6454
rect 2205 6446 2209 6454
rect 2218 6446 2222 6454
rect 2227 6446 2231 6454
rect 2244 6446 2248 6454
rect 2261 6446 2265 6454
rect 2272 6446 2276 6454
rect 2280 6446 2284 6454
rect 2288 6446 2292 6454
rect 2296 6446 2300 6454
rect 2304 6446 2308 6454
rect 2312 6446 2316 6454
rect 983 6401 987 6409
rect 998 6401 1002 6409
rect 1073 6401 1077 6409
rect 1088 6401 1092 6409
rect 1154 6401 1158 6409
rect 1169 6401 1173 6409
rect 1209 6400 1213 6408
rect 1217 6400 1221 6408
rect 1227 6400 1231 6408
rect 1244 6400 1248 6408
rect 1252 6400 1256 6408
rect 1260 6400 1264 6408
rect 1273 6400 1277 6408
rect 1282 6400 1286 6408
rect 1299 6400 1303 6408
rect 1316 6400 1320 6408
rect 1327 6400 1331 6408
rect 1335 6400 1339 6408
rect 1343 6400 1347 6408
rect 1351 6400 1355 6408
rect 1359 6400 1363 6408
rect 1367 6400 1371 6408
rect 1928 6401 1932 6409
rect 1943 6401 1947 6409
rect 2018 6401 2022 6409
rect 2033 6401 2037 6409
rect 2099 6401 2103 6409
rect 2114 6401 2118 6409
rect 2154 6400 2158 6408
rect 2162 6400 2166 6408
rect 2172 6400 2176 6408
rect 2189 6400 2193 6408
rect 2197 6400 2201 6408
rect 2205 6400 2209 6408
rect 2218 6400 2222 6408
rect 2227 6400 2231 6408
rect 2244 6400 2248 6408
rect 2261 6400 2265 6408
rect 2272 6400 2276 6408
rect 2280 6400 2284 6408
rect 2288 6400 2292 6408
rect 2296 6400 2300 6408
rect 2304 6400 2308 6408
rect 2312 6400 2316 6408
rect 960 6301 964 6309
rect 968 6301 972 6309
rect 983 6307 987 6315
rect 998 6307 1002 6315
rect 1014 6301 1018 6309
rect 1022 6301 1026 6309
rect 1050 6301 1054 6309
rect 1058 6301 1062 6309
rect 1073 6307 1077 6315
rect 1088 6307 1092 6315
rect 1104 6301 1108 6309
rect 1112 6301 1116 6309
rect 1131 6301 1135 6309
rect 1139 6301 1143 6309
rect 1154 6307 1158 6315
rect 1169 6307 1173 6315
rect 1209 6314 1213 6322
rect 1217 6314 1221 6322
rect 1227 6314 1231 6322
rect 1244 6314 1248 6322
rect 1252 6314 1256 6322
rect 1260 6314 1264 6322
rect 1273 6314 1277 6322
rect 1282 6314 1286 6322
rect 1299 6314 1303 6322
rect 1316 6314 1320 6322
rect 1327 6314 1331 6322
rect 1335 6314 1339 6322
rect 1343 6314 1347 6322
rect 1351 6314 1355 6322
rect 1359 6314 1363 6322
rect 1367 6314 1371 6322
rect 1905 6301 1909 6309
rect 1913 6301 1917 6309
rect 1928 6307 1932 6315
rect 1943 6307 1947 6315
rect 1959 6301 1963 6309
rect 1967 6301 1971 6309
rect 1995 6301 1999 6309
rect 2003 6301 2007 6309
rect 2018 6307 2022 6315
rect 2033 6307 2037 6315
rect 2049 6301 2053 6309
rect 2057 6301 2061 6309
rect 2076 6301 2080 6309
rect 2084 6301 2088 6309
rect 2099 6307 2103 6315
rect 2114 6307 2118 6315
rect 2154 6314 2158 6322
rect 2162 6314 2166 6322
rect 2172 6314 2176 6322
rect 2189 6314 2193 6322
rect 2197 6314 2201 6322
rect 2205 6314 2209 6322
rect 2218 6314 2222 6322
rect 2227 6314 2231 6322
rect 2244 6314 2248 6322
rect 2261 6314 2265 6322
rect 2272 6314 2276 6322
rect 2280 6314 2284 6322
rect 2288 6314 2292 6322
rect 2296 6314 2300 6322
rect 2304 6314 2308 6322
rect 2312 6314 2316 6322
rect 1049 6266 1053 6274
rect 1064 6266 1068 6274
rect 1154 6266 1158 6274
rect 1169 6266 1173 6274
rect 1209 6268 1213 6276
rect 1217 6268 1221 6276
rect 1227 6268 1231 6276
rect 1244 6268 1248 6276
rect 1252 6268 1256 6276
rect 1260 6268 1264 6276
rect 1273 6268 1277 6276
rect 1282 6268 1286 6276
rect 1299 6268 1303 6276
rect 1316 6268 1320 6276
rect 1327 6268 1331 6276
rect 1335 6268 1339 6276
rect 1343 6268 1347 6276
rect 1351 6268 1355 6276
rect 1359 6268 1363 6276
rect 1367 6268 1371 6276
rect 1994 6266 1998 6274
rect 2009 6266 2013 6274
rect 2099 6266 2103 6274
rect 2114 6266 2118 6274
rect 2154 6268 2158 6276
rect 2162 6268 2166 6276
rect 2172 6268 2176 6276
rect 2189 6268 2193 6276
rect 2197 6268 2201 6276
rect 2205 6268 2209 6276
rect 2218 6268 2222 6276
rect 2227 6268 2231 6276
rect 2244 6268 2248 6276
rect 2261 6268 2265 6276
rect 2272 6268 2276 6276
rect 2280 6268 2284 6276
rect 2288 6268 2292 6276
rect 2296 6268 2300 6276
rect 2304 6268 2308 6276
rect 2312 6268 2316 6276
rect 1026 6169 1030 6177
rect 1034 6169 1038 6177
rect 1049 6175 1053 6183
rect 1064 6175 1068 6183
rect 1080 6169 1084 6177
rect 1088 6169 1092 6177
rect 1131 6169 1135 6177
rect 1139 6169 1143 6177
rect 1154 6175 1158 6183
rect 1169 6175 1173 6183
rect 1209 6182 1213 6190
rect 1217 6182 1221 6190
rect 1227 6182 1231 6190
rect 1244 6182 1248 6190
rect 1252 6182 1256 6190
rect 1260 6182 1264 6190
rect 1273 6182 1277 6190
rect 1282 6182 1286 6190
rect 1299 6182 1303 6190
rect 1316 6182 1320 6190
rect 1327 6182 1331 6190
rect 1335 6182 1339 6190
rect 1343 6182 1347 6190
rect 1351 6182 1355 6190
rect 1359 6182 1363 6190
rect 1367 6182 1371 6190
rect 1971 6169 1975 6177
rect 1979 6169 1983 6177
rect 1994 6175 1998 6183
rect 2009 6175 2013 6183
rect 2025 6169 2029 6177
rect 2033 6169 2037 6177
rect 2076 6169 2080 6177
rect 2084 6169 2088 6177
rect 2099 6175 2103 6183
rect 2114 6175 2118 6183
rect 2154 6182 2158 6190
rect 2162 6182 2166 6190
rect 2172 6182 2176 6190
rect 2189 6182 2193 6190
rect 2197 6182 2201 6190
rect 2205 6182 2209 6190
rect 2218 6182 2222 6190
rect 2227 6182 2231 6190
rect 2244 6182 2248 6190
rect 2261 6182 2265 6190
rect 2272 6182 2276 6190
rect 2280 6182 2284 6190
rect 2288 6182 2292 6190
rect 2296 6182 2300 6190
rect 2304 6182 2308 6190
rect 2312 6182 2316 6190
rect 1073 6135 1077 6143
rect 1088 6135 1092 6143
rect 1154 6135 1158 6143
rect 1169 6135 1173 6143
rect 1209 6136 1213 6144
rect 1217 6136 1221 6144
rect 1227 6136 1231 6144
rect 1244 6136 1248 6144
rect 1252 6136 1256 6144
rect 1260 6136 1264 6144
rect 1273 6136 1277 6144
rect 1282 6136 1286 6144
rect 1299 6136 1303 6144
rect 1316 6136 1320 6144
rect 1327 6136 1331 6144
rect 1335 6136 1339 6144
rect 1343 6136 1347 6144
rect 1351 6136 1355 6144
rect 1359 6136 1363 6144
rect 1367 6136 1371 6144
rect 2018 6135 2022 6143
rect 2033 6135 2037 6143
rect 2099 6135 2103 6143
rect 2114 6135 2118 6143
rect 2154 6136 2158 6144
rect 2162 6136 2166 6144
rect 2172 6136 2176 6144
rect 2189 6136 2193 6144
rect 2197 6136 2201 6144
rect 2205 6136 2209 6144
rect 2218 6136 2222 6144
rect 2227 6136 2231 6144
rect 2244 6136 2248 6144
rect 2261 6136 2265 6144
rect 2272 6136 2276 6144
rect 2280 6136 2284 6144
rect 2288 6136 2292 6144
rect 2296 6136 2300 6144
rect 2304 6136 2308 6144
rect 2312 6136 2316 6144
rect 1609 6101 1613 6109
rect 1622 6101 1626 6109
rect 1630 6101 1634 6109
rect 1638 6101 1642 6105
rect 1646 6101 1650 6109
rect 1659 6101 1663 6109
rect 1672 6101 1676 6109
rect 1680 6101 1684 6109
rect 1688 6101 1692 6109
rect 1696 6101 1700 6105
rect 1704 6101 1708 6109
rect 1717 6101 1721 6109
rect 1725 6101 1729 6109
rect 1733 6101 1737 6109
rect 2554 6101 2558 6109
rect 2567 6101 2571 6109
rect 2575 6101 2579 6109
rect 2583 6101 2587 6105
rect 2591 6101 2595 6109
rect 2604 6101 2608 6109
rect 2617 6101 2621 6109
rect 2625 6101 2629 6109
rect 2633 6101 2637 6109
rect 2641 6101 2645 6105
rect 2649 6101 2653 6109
rect 2662 6101 2666 6109
rect 2670 6101 2674 6109
rect 2678 6101 2682 6109
rect 1050 6037 1054 6045
rect 1058 6037 1062 6045
rect 1073 6043 1077 6051
rect 1088 6043 1092 6051
rect 1104 6037 1108 6045
rect 1112 6037 1116 6045
rect 1131 6037 1135 6045
rect 1139 6037 1143 6045
rect 1154 6043 1158 6051
rect 1169 6043 1173 6051
rect 1209 6050 1213 6058
rect 1217 6050 1221 6058
rect 1227 6050 1231 6058
rect 1244 6050 1248 6058
rect 1252 6050 1256 6058
rect 1260 6050 1264 6058
rect 1273 6050 1277 6058
rect 1282 6050 1286 6058
rect 1299 6050 1303 6058
rect 1316 6050 1320 6058
rect 1327 6050 1331 6058
rect 1335 6050 1339 6058
rect 1343 6050 1347 6058
rect 1351 6050 1355 6058
rect 1359 6050 1363 6058
rect 1367 6050 1371 6058
rect 1185 6037 1189 6045
rect 1193 6037 1197 6045
rect 1995 6037 1999 6045
rect 2003 6037 2007 6045
rect 2018 6043 2022 6051
rect 2033 6043 2037 6051
rect 2049 6037 2053 6045
rect 2057 6037 2061 6045
rect 2076 6037 2080 6045
rect 2084 6037 2088 6045
rect 2099 6043 2103 6051
rect 2114 6043 2118 6051
rect 2154 6050 2158 6058
rect 2162 6050 2166 6058
rect 2172 6050 2176 6058
rect 2189 6050 2193 6058
rect 2197 6050 2201 6058
rect 2205 6050 2209 6058
rect 2218 6050 2222 6058
rect 2227 6050 2231 6058
rect 2244 6050 2248 6058
rect 2261 6050 2265 6058
rect 2272 6050 2276 6058
rect 2280 6050 2284 6058
rect 2288 6050 2292 6058
rect 2296 6050 2300 6058
rect 2304 6050 2308 6058
rect 2312 6050 2316 6058
rect 2130 6037 2134 6045
rect 2138 6037 2142 6045
rect 1600 5999 1604 6007
rect 1608 5999 1612 6007
rect 1616 5999 1620 6007
rect 1629 5999 1633 6007
rect 1637 5999 1641 6003
rect 1645 5999 1649 6007
rect 1653 5999 1657 6007
rect 1661 5999 1665 6007
rect 1674 5999 1678 6007
rect 1687 5999 1691 6007
rect 1695 5999 1699 6003
rect 1703 5999 1707 6007
rect 1711 5999 1715 6007
rect 1724 5999 1728 6007
rect 2545 5999 2549 6007
rect 2553 5999 2557 6007
rect 2561 5999 2565 6007
rect 2574 5999 2578 6007
rect 2582 5999 2586 6003
rect 2590 5999 2594 6007
rect 2598 5999 2602 6007
rect 2606 5999 2610 6007
rect 2619 5999 2623 6007
rect 2632 5999 2636 6007
rect 2640 5999 2644 6003
rect 2648 5999 2652 6007
rect 2656 5999 2660 6007
rect 2669 5999 2673 6007
rect 852 5966 856 5974
rect 860 5966 864 5974
rect 868 5966 872 5974
rect 881 5966 885 5974
rect 889 5966 893 5970
rect 897 5966 901 5974
rect 905 5966 909 5974
rect 913 5966 917 5974
rect 926 5966 930 5974
rect 939 5966 943 5974
rect 947 5966 951 5970
rect 955 5966 959 5974
rect 963 5966 967 5974
rect 976 5966 980 5974
rect 984 5966 988 5974
rect 992 5966 996 5974
rect 1000 5966 1004 5974
rect 1013 5966 1017 5974
rect 1021 5966 1025 5970
rect 1029 5966 1033 5974
rect 1037 5966 1041 5974
rect 1045 5966 1049 5974
rect 1058 5966 1062 5974
rect 1071 5966 1075 5974
rect 1079 5966 1083 5970
rect 1087 5966 1091 5974
rect 1095 5966 1099 5974
rect 1108 5966 1112 5974
rect 1116 5966 1120 5974
rect 1124 5966 1128 5974
rect 1132 5966 1136 5974
rect 1145 5966 1149 5974
rect 1153 5966 1157 5970
rect 1161 5966 1165 5974
rect 1169 5966 1173 5974
rect 1177 5966 1181 5974
rect 1190 5966 1194 5974
rect 1203 5966 1207 5974
rect 1211 5966 1215 5970
rect 1219 5966 1223 5974
rect 1227 5966 1231 5974
rect 1240 5966 1244 5974
rect 1248 5966 1252 5974
rect 1256 5966 1260 5974
rect 1264 5966 1268 5974
rect 1277 5966 1281 5974
rect 1285 5966 1289 5970
rect 1293 5966 1297 5974
rect 1301 5966 1305 5974
rect 1309 5966 1313 5974
rect 1322 5966 1326 5974
rect 1335 5966 1339 5974
rect 1343 5966 1347 5970
rect 1351 5966 1355 5974
rect 1359 5966 1363 5974
rect 1372 5966 1376 5974
rect 1797 5966 1801 5974
rect 1805 5966 1809 5974
rect 1813 5966 1817 5974
rect 1826 5966 1830 5974
rect 1834 5966 1838 5970
rect 1842 5966 1846 5974
rect 1850 5966 1854 5974
rect 1858 5966 1862 5974
rect 1871 5966 1875 5974
rect 1884 5966 1888 5974
rect 1892 5966 1896 5970
rect 1900 5966 1904 5974
rect 1908 5966 1912 5974
rect 1921 5966 1925 5974
rect 1929 5966 1933 5974
rect 1937 5966 1941 5974
rect 1945 5966 1949 5974
rect 1958 5966 1962 5974
rect 1966 5966 1970 5970
rect 1974 5966 1978 5974
rect 1982 5966 1986 5974
rect 1990 5966 1994 5974
rect 2003 5966 2007 5974
rect 2016 5966 2020 5974
rect 2024 5966 2028 5970
rect 2032 5966 2036 5974
rect 2040 5966 2044 5974
rect 2053 5966 2057 5974
rect 2061 5966 2065 5974
rect 2069 5966 2073 5974
rect 2077 5966 2081 5974
rect 2090 5966 2094 5974
rect 2098 5966 2102 5970
rect 2106 5966 2110 5974
rect 2114 5966 2118 5974
rect 2122 5966 2126 5974
rect 2135 5966 2139 5974
rect 2148 5966 2152 5974
rect 2156 5966 2160 5970
rect 2164 5966 2168 5974
rect 2172 5966 2176 5974
rect 2185 5966 2189 5974
rect 2193 5966 2197 5974
rect 2201 5966 2205 5974
rect 2209 5966 2213 5974
rect 2222 5966 2226 5974
rect 2230 5966 2234 5970
rect 2238 5966 2242 5974
rect 2246 5966 2250 5974
rect 2254 5966 2258 5974
rect 2267 5966 2271 5974
rect 2280 5966 2284 5974
rect 2288 5966 2292 5970
rect 2296 5966 2300 5974
rect 2304 5966 2308 5974
rect 2317 5966 2321 5974
rect 1468 5887 1472 5895
rect 1476 5887 1480 5895
rect 1484 5887 1488 5895
rect 1497 5887 1501 5895
rect 1505 5887 1509 5891
rect 1513 5887 1517 5895
rect 1521 5887 1525 5895
rect 1529 5887 1533 5895
rect 1542 5887 1546 5895
rect 1555 5887 1559 5895
rect 1563 5887 1567 5891
rect 1571 5887 1575 5895
rect 1579 5887 1583 5895
rect 1592 5887 1596 5895
rect 1600 5887 1604 5895
rect 1608 5887 1612 5895
rect 1616 5887 1620 5895
rect 1629 5887 1633 5895
rect 1637 5887 1641 5891
rect 1645 5887 1649 5895
rect 1653 5887 1657 5895
rect 1661 5887 1665 5895
rect 1674 5887 1678 5895
rect 1687 5887 1691 5895
rect 1695 5887 1699 5891
rect 1703 5887 1707 5895
rect 1711 5887 1715 5895
rect 1724 5887 1728 5895
rect 1732 5887 1736 5895
rect 1740 5887 1744 5895
rect 1748 5887 1752 5895
rect 1761 5887 1765 5895
rect 1769 5887 1773 5891
rect 1777 5887 1781 5895
rect 1785 5887 1789 5895
rect 1793 5887 1797 5895
rect 1806 5887 1810 5895
rect 1819 5887 1823 5895
rect 1827 5887 1831 5891
rect 1835 5887 1839 5895
rect 1843 5887 1847 5895
rect 1856 5887 1860 5895
rect 2413 5887 2417 5895
rect 2421 5887 2425 5895
rect 2429 5887 2433 5895
rect 2442 5887 2446 5895
rect 2450 5887 2454 5891
rect 2458 5887 2462 5895
rect 2466 5887 2470 5895
rect 2474 5887 2478 5895
rect 2487 5887 2491 5895
rect 2500 5887 2504 5895
rect 2508 5887 2512 5891
rect 2516 5887 2520 5895
rect 2524 5887 2528 5895
rect 2537 5887 2541 5895
rect 2545 5887 2549 5895
rect 2553 5887 2557 5895
rect 2561 5887 2565 5895
rect 2574 5887 2578 5895
rect 2582 5887 2586 5891
rect 2590 5887 2594 5895
rect 2598 5887 2602 5895
rect 2606 5887 2610 5895
rect 2619 5887 2623 5895
rect 2632 5887 2636 5895
rect 2640 5887 2644 5891
rect 2648 5887 2652 5895
rect 2656 5887 2660 5895
rect 2669 5887 2673 5895
rect 2677 5887 2681 5895
rect 2685 5887 2689 5895
rect 2693 5887 2697 5895
rect 2706 5887 2710 5895
rect 2714 5887 2718 5891
rect 2722 5887 2726 5895
rect 2730 5887 2734 5895
rect 2738 5887 2742 5895
rect 2751 5887 2755 5895
rect 2764 5887 2768 5895
rect 2772 5887 2776 5891
rect 2780 5887 2784 5895
rect 2788 5887 2792 5895
rect 2801 5887 2805 5895
rect 1468 5747 1472 5755
rect 1476 5747 1480 5755
rect 1484 5747 1488 5755
rect 1497 5747 1501 5755
rect 1505 5747 1509 5751
rect 1513 5747 1517 5755
rect 1521 5747 1525 5755
rect 1529 5747 1533 5755
rect 1542 5747 1546 5755
rect 1555 5747 1559 5755
rect 1563 5747 1567 5751
rect 1571 5747 1575 5755
rect 1579 5747 1583 5755
rect 1592 5747 1596 5755
rect 1600 5747 1604 5755
rect 1608 5747 1612 5755
rect 1616 5747 1620 5755
rect 1629 5747 1633 5755
rect 1637 5747 1641 5751
rect 1645 5747 1649 5755
rect 1653 5747 1657 5755
rect 1661 5747 1665 5755
rect 1674 5747 1678 5755
rect 1687 5747 1691 5755
rect 1695 5747 1699 5751
rect 1703 5747 1707 5755
rect 1711 5747 1715 5755
rect 1724 5747 1728 5755
rect 1732 5747 1736 5755
rect 1740 5747 1744 5755
rect 1748 5747 1752 5755
rect 1761 5747 1765 5755
rect 1769 5747 1773 5751
rect 1777 5747 1781 5755
rect 1785 5747 1789 5755
rect 1793 5747 1797 5755
rect 1806 5747 1810 5755
rect 1819 5747 1823 5755
rect 1827 5747 1831 5751
rect 1835 5747 1839 5755
rect 1843 5747 1847 5755
rect 1856 5747 1860 5755
rect 2413 5747 2417 5755
rect 2421 5747 2425 5755
rect 2429 5747 2433 5755
rect 2442 5747 2446 5755
rect 2450 5747 2454 5751
rect 2458 5747 2462 5755
rect 2466 5747 2470 5755
rect 2474 5747 2478 5755
rect 2487 5747 2491 5755
rect 2500 5747 2504 5755
rect 2508 5747 2512 5751
rect 2516 5747 2520 5755
rect 2524 5747 2528 5755
rect 2537 5747 2541 5755
rect 2545 5747 2549 5755
rect 2553 5747 2557 5755
rect 2561 5747 2565 5755
rect 2574 5747 2578 5755
rect 2582 5747 2586 5751
rect 2590 5747 2594 5755
rect 2598 5747 2602 5755
rect 2606 5747 2610 5755
rect 2619 5747 2623 5755
rect 2632 5747 2636 5755
rect 2640 5747 2644 5751
rect 2648 5747 2652 5755
rect 2656 5747 2660 5755
rect 2669 5747 2673 5755
rect 2677 5747 2681 5755
rect 2685 5747 2689 5755
rect 2693 5747 2697 5755
rect 2706 5747 2710 5755
rect 2714 5747 2718 5751
rect 2722 5747 2726 5755
rect 2730 5747 2734 5755
rect 2738 5747 2742 5755
rect 2751 5747 2755 5755
rect 2764 5747 2768 5755
rect 2772 5747 2776 5751
rect 2780 5747 2784 5755
rect 2788 5747 2792 5755
rect 2801 5747 2805 5755
rect 949 5717 953 5725
rect 957 5717 961 5725
rect 965 5717 969 5725
rect 978 5717 982 5725
rect 986 5717 990 5721
rect 994 5717 998 5725
rect 1002 5717 1006 5725
rect 1010 5717 1014 5725
rect 1023 5717 1027 5725
rect 1036 5717 1040 5725
rect 1044 5717 1048 5721
rect 1052 5717 1056 5725
rect 1060 5717 1064 5725
rect 1073 5717 1077 5725
rect 1894 5717 1898 5725
rect 1902 5717 1906 5725
rect 1910 5717 1914 5725
rect 1923 5717 1927 5725
rect 1931 5717 1935 5721
rect 1939 5717 1943 5725
rect 1947 5717 1951 5725
rect 1955 5717 1959 5725
rect 1968 5717 1972 5725
rect 1981 5717 1985 5725
rect 1989 5717 1993 5721
rect 1997 5717 2001 5725
rect 2005 5717 2009 5725
rect 2018 5717 2022 5725
rect 1468 5661 1472 5669
rect 1476 5661 1480 5669
rect 1484 5661 1488 5669
rect 1497 5661 1501 5669
rect 1505 5661 1509 5665
rect 1513 5661 1517 5669
rect 1521 5661 1525 5669
rect 1529 5661 1533 5669
rect 1542 5661 1546 5669
rect 1555 5661 1559 5669
rect 1563 5661 1567 5665
rect 1571 5661 1575 5669
rect 1579 5661 1583 5669
rect 1592 5661 1596 5669
rect 1600 5661 1604 5669
rect 1608 5661 1612 5669
rect 1616 5661 1620 5669
rect 1629 5661 1633 5669
rect 1637 5661 1641 5665
rect 1645 5661 1649 5669
rect 1653 5661 1657 5669
rect 1661 5661 1665 5669
rect 1674 5661 1678 5669
rect 1687 5661 1691 5669
rect 1695 5661 1699 5665
rect 1703 5661 1707 5669
rect 1711 5661 1715 5669
rect 1724 5661 1728 5669
rect 1732 5661 1736 5669
rect 1740 5661 1744 5669
rect 1748 5661 1752 5669
rect 1761 5661 1765 5669
rect 1769 5661 1773 5665
rect 1777 5661 1781 5669
rect 1785 5661 1789 5669
rect 1793 5661 1797 5669
rect 1806 5661 1810 5669
rect 1819 5661 1823 5669
rect 1827 5661 1831 5665
rect 1835 5661 1839 5669
rect 1843 5661 1847 5669
rect 1856 5661 1860 5669
rect 2413 5661 2417 5669
rect 2421 5661 2425 5669
rect 2429 5661 2433 5669
rect 2442 5661 2446 5669
rect 2450 5661 2454 5665
rect 2458 5661 2462 5669
rect 2466 5661 2470 5669
rect 2474 5661 2478 5669
rect 2487 5661 2491 5669
rect 2500 5661 2504 5669
rect 2508 5661 2512 5665
rect 2516 5661 2520 5669
rect 2524 5661 2528 5669
rect 2537 5661 2541 5669
rect 2545 5661 2549 5669
rect 2553 5661 2557 5669
rect 2561 5661 2565 5669
rect 2574 5661 2578 5669
rect 2582 5661 2586 5665
rect 2590 5661 2594 5669
rect 2598 5661 2602 5669
rect 2606 5661 2610 5669
rect 2619 5661 2623 5669
rect 2632 5661 2636 5669
rect 2640 5661 2644 5665
rect 2648 5661 2652 5669
rect 2656 5661 2660 5669
rect 2669 5661 2673 5669
rect 2677 5661 2681 5669
rect 2685 5661 2689 5669
rect 2693 5661 2697 5669
rect 2706 5661 2710 5669
rect 2714 5661 2718 5665
rect 2722 5661 2726 5669
rect 2730 5661 2734 5669
rect 2738 5661 2742 5669
rect 2751 5661 2755 5669
rect 2764 5661 2768 5669
rect 2772 5661 2776 5665
rect 2780 5661 2784 5669
rect 2788 5661 2792 5669
rect 2801 5661 2805 5669
rect 949 5631 953 5639
rect 957 5631 961 5639
rect 965 5631 969 5639
rect 978 5631 982 5639
rect 986 5631 990 5635
rect 994 5631 998 5639
rect 1002 5631 1006 5639
rect 1010 5631 1014 5639
rect 1023 5631 1027 5639
rect 1036 5631 1040 5639
rect 1044 5631 1048 5635
rect 1052 5631 1056 5639
rect 1060 5631 1064 5639
rect 1073 5631 1077 5639
rect 1894 5631 1898 5639
rect 1902 5631 1906 5639
rect 1910 5631 1914 5639
rect 1923 5631 1927 5639
rect 1931 5631 1935 5635
rect 1939 5631 1943 5639
rect 1947 5631 1951 5639
rect 1955 5631 1959 5639
rect 1968 5631 1972 5639
rect 1981 5631 1985 5639
rect 1989 5631 1993 5635
rect 1997 5631 2001 5639
rect 2005 5631 2009 5639
rect 2018 5631 2022 5639
rect 948 5550 952 5558
rect 956 5550 960 5558
rect 966 5550 970 5558
rect 983 5550 987 5558
rect 991 5550 995 5558
rect 999 5550 1003 5558
rect 1012 5550 1016 5558
rect 1021 5550 1025 5558
rect 1038 5550 1042 5558
rect 1055 5550 1059 5558
rect 1066 5550 1070 5558
rect 1074 5550 1078 5558
rect 1082 5550 1086 5558
rect 1090 5550 1094 5558
rect 1098 5550 1102 5558
rect 1107 5550 1111 5558
rect 1115 5550 1119 5558
rect 1125 5550 1129 5558
rect 1133 5550 1137 5558
rect 1154 5555 1158 5563
rect 1169 5555 1173 5563
rect 1209 5550 1213 5558
rect 1217 5550 1221 5558
rect 1227 5550 1231 5558
rect 1244 5550 1248 5558
rect 1252 5550 1256 5558
rect 1260 5550 1264 5558
rect 1273 5550 1277 5558
rect 1282 5550 1286 5558
rect 1299 5550 1303 5558
rect 1316 5550 1320 5558
rect 1327 5550 1331 5558
rect 1335 5550 1339 5558
rect 1343 5550 1347 5558
rect 1351 5550 1355 5558
rect 1359 5550 1363 5558
rect 1367 5550 1371 5558
rect 1893 5550 1897 5558
rect 1901 5550 1905 5558
rect 1911 5550 1915 5558
rect 1928 5550 1932 5558
rect 1936 5550 1940 5558
rect 1944 5550 1948 5558
rect 1957 5550 1961 5558
rect 1966 5550 1970 5558
rect 1983 5550 1987 5558
rect 2000 5550 2004 5558
rect 2011 5550 2015 5558
rect 2019 5550 2023 5558
rect 2027 5550 2031 5558
rect 2035 5550 2039 5558
rect 2043 5550 2047 5558
rect 2052 5550 2056 5558
rect 2060 5550 2064 5558
rect 2070 5550 2074 5558
rect 2078 5550 2082 5558
rect 2099 5555 2103 5563
rect 2114 5555 2118 5563
rect 2154 5550 2158 5558
rect 2162 5550 2166 5558
rect 2172 5550 2176 5558
rect 2189 5550 2193 5558
rect 2197 5550 2201 5558
rect 2205 5550 2209 5558
rect 2218 5550 2222 5558
rect 2227 5550 2231 5558
rect 2244 5550 2248 5558
rect 2261 5550 2265 5558
rect 2272 5550 2276 5558
rect 2280 5550 2284 5558
rect 2288 5550 2292 5558
rect 2296 5550 2300 5558
rect 2304 5550 2308 5558
rect 2312 5550 2316 5558
rect 1468 5519 1472 5527
rect 1476 5519 1480 5527
rect 1484 5519 1488 5527
rect 1497 5519 1501 5527
rect 1505 5519 1509 5523
rect 1513 5519 1517 5527
rect 1521 5519 1525 5527
rect 1529 5519 1533 5527
rect 1542 5519 1546 5527
rect 1555 5519 1559 5527
rect 1563 5519 1567 5523
rect 1571 5519 1575 5527
rect 1579 5519 1583 5527
rect 1592 5519 1596 5527
rect 1600 5519 1604 5527
rect 1608 5519 1612 5527
rect 1616 5519 1620 5527
rect 1629 5519 1633 5527
rect 1637 5519 1641 5523
rect 1645 5519 1649 5527
rect 1653 5519 1657 5527
rect 1661 5519 1665 5527
rect 1674 5519 1678 5527
rect 1687 5519 1691 5527
rect 1695 5519 1699 5523
rect 1703 5519 1707 5527
rect 1711 5519 1715 5527
rect 1724 5519 1728 5527
rect 1732 5519 1736 5527
rect 1740 5519 1744 5527
rect 1748 5519 1752 5527
rect 1761 5519 1765 5527
rect 1769 5519 1773 5523
rect 1777 5519 1781 5527
rect 1785 5519 1789 5527
rect 1793 5519 1797 5527
rect 1806 5519 1810 5527
rect 1819 5519 1823 5527
rect 1827 5519 1831 5523
rect 1835 5519 1839 5527
rect 1843 5519 1847 5527
rect 1856 5519 1860 5527
rect 2413 5519 2417 5527
rect 2421 5519 2425 5527
rect 2429 5519 2433 5527
rect 2442 5519 2446 5527
rect 2450 5519 2454 5523
rect 2458 5519 2462 5527
rect 2466 5519 2470 5527
rect 2474 5519 2478 5527
rect 2487 5519 2491 5527
rect 2500 5519 2504 5527
rect 2508 5519 2512 5523
rect 2516 5519 2520 5527
rect 2524 5519 2528 5527
rect 2537 5519 2541 5527
rect 2545 5519 2549 5527
rect 2553 5519 2557 5527
rect 2561 5519 2565 5527
rect 2574 5519 2578 5527
rect 2582 5519 2586 5523
rect 2590 5519 2594 5527
rect 2598 5519 2602 5527
rect 2606 5519 2610 5527
rect 2619 5519 2623 5527
rect 2632 5519 2636 5527
rect 2640 5519 2644 5523
rect 2648 5519 2652 5527
rect 2656 5519 2660 5527
rect 2669 5519 2673 5527
rect 2677 5519 2681 5527
rect 2685 5519 2689 5527
rect 2693 5519 2697 5527
rect 2706 5519 2710 5527
rect 2714 5519 2718 5523
rect 2722 5519 2726 5527
rect 2730 5519 2734 5527
rect 2738 5519 2742 5527
rect 2751 5519 2755 5527
rect 2764 5519 2768 5527
rect 2772 5519 2776 5523
rect 2780 5519 2784 5527
rect 2788 5519 2792 5527
rect 2801 5519 2805 5527
rect 1131 5451 1135 5459
rect 1139 5451 1143 5459
rect 1154 5457 1158 5465
rect 1169 5457 1173 5465
rect 1209 5464 1213 5472
rect 1217 5464 1221 5472
rect 1227 5464 1231 5472
rect 1244 5464 1248 5472
rect 1252 5464 1256 5472
rect 1260 5464 1264 5472
rect 1273 5464 1277 5472
rect 1282 5464 1286 5472
rect 1299 5464 1303 5472
rect 1316 5464 1320 5472
rect 1327 5464 1331 5472
rect 1335 5464 1339 5472
rect 1343 5464 1347 5472
rect 1351 5464 1355 5472
rect 1359 5464 1363 5472
rect 1367 5464 1371 5472
rect 1763 5448 1767 5456
rect 1778 5448 1782 5456
rect 2076 5451 2080 5459
rect 2084 5451 2088 5459
rect 2099 5457 2103 5465
rect 2114 5457 2118 5465
rect 2154 5464 2158 5472
rect 2162 5464 2166 5472
rect 2172 5464 2176 5472
rect 2189 5464 2193 5472
rect 2197 5464 2201 5472
rect 2205 5464 2209 5472
rect 2218 5464 2222 5472
rect 2227 5464 2231 5472
rect 2244 5464 2248 5472
rect 2261 5464 2265 5472
rect 2272 5464 2276 5472
rect 2280 5464 2284 5472
rect 2288 5464 2292 5472
rect 2296 5464 2300 5472
rect 2304 5464 2308 5472
rect 2312 5464 2316 5472
rect 983 5419 987 5427
rect 998 5419 1002 5427
rect 1073 5419 1077 5427
rect 1088 5419 1092 5427
rect 1154 5419 1158 5427
rect 1169 5419 1173 5427
rect 1209 5418 1213 5426
rect 1217 5418 1221 5426
rect 1227 5418 1231 5426
rect 1244 5418 1248 5426
rect 1252 5418 1256 5426
rect 1260 5418 1264 5426
rect 1273 5418 1277 5426
rect 1282 5418 1286 5426
rect 1299 5418 1303 5426
rect 1316 5418 1320 5426
rect 1327 5418 1331 5426
rect 1335 5418 1339 5426
rect 1343 5418 1347 5426
rect 1351 5418 1355 5426
rect 1359 5418 1363 5426
rect 1367 5418 1371 5426
rect 1928 5419 1932 5427
rect 1943 5419 1947 5427
rect 2018 5419 2022 5427
rect 2033 5419 2037 5427
rect 2099 5419 2103 5427
rect 2114 5419 2118 5427
rect 2154 5418 2158 5426
rect 2162 5418 2166 5426
rect 2172 5418 2176 5426
rect 2189 5418 2193 5426
rect 2197 5418 2201 5426
rect 2205 5418 2209 5426
rect 2218 5418 2222 5426
rect 2227 5418 2231 5426
rect 2244 5418 2248 5426
rect 2261 5418 2265 5426
rect 2272 5418 2276 5426
rect 2280 5418 2284 5426
rect 2288 5418 2292 5426
rect 2296 5418 2300 5426
rect 2304 5418 2308 5426
rect 2312 5418 2316 5426
rect 960 5319 964 5327
rect 968 5319 972 5327
rect 983 5325 987 5333
rect 998 5325 1002 5333
rect 1014 5319 1018 5327
rect 1022 5319 1026 5327
rect 1050 5319 1054 5327
rect 1058 5319 1062 5327
rect 1073 5325 1077 5333
rect 1088 5325 1092 5333
rect 1637 5349 1653 5379
rect 1657 5349 1673 5379
rect 1690 5349 1706 5379
rect 1710 5349 1726 5379
rect 1740 5346 1744 5354
rect 1748 5346 1752 5354
rect 1763 5352 1767 5360
rect 1778 5352 1782 5360
rect 1794 5346 1798 5354
rect 1802 5346 1806 5354
rect 1816 5346 1820 5354
rect 1824 5346 1828 5354
rect 1104 5319 1108 5327
rect 1112 5319 1116 5327
rect 1131 5319 1135 5327
rect 1139 5319 1143 5327
rect 1154 5325 1158 5333
rect 1169 5325 1173 5333
rect 1209 5332 1213 5340
rect 1217 5332 1221 5340
rect 1227 5332 1231 5340
rect 1244 5332 1248 5340
rect 1252 5332 1256 5340
rect 1260 5332 1264 5340
rect 1273 5332 1277 5340
rect 1282 5332 1286 5340
rect 1299 5332 1303 5340
rect 1316 5332 1320 5340
rect 1327 5332 1331 5340
rect 1335 5332 1339 5340
rect 1343 5332 1347 5340
rect 1351 5332 1355 5340
rect 1359 5332 1363 5340
rect 1367 5332 1371 5340
rect 1763 5318 1767 5326
rect 1778 5318 1782 5326
rect 1905 5319 1909 5327
rect 1913 5319 1917 5327
rect 1928 5325 1932 5333
rect 1943 5325 1947 5333
rect 1959 5319 1963 5327
rect 1967 5319 1971 5327
rect 1995 5319 1999 5327
rect 2003 5319 2007 5327
rect 2018 5325 2022 5333
rect 2033 5325 2037 5333
rect 2049 5319 2053 5327
rect 2057 5319 2061 5327
rect 2076 5319 2080 5327
rect 2084 5319 2088 5327
rect 2099 5325 2103 5333
rect 2114 5325 2118 5333
rect 2154 5332 2158 5340
rect 2162 5332 2166 5340
rect 2172 5332 2176 5340
rect 2189 5332 2193 5340
rect 2197 5332 2201 5340
rect 2205 5332 2209 5340
rect 2218 5332 2222 5340
rect 2227 5332 2231 5340
rect 2244 5332 2248 5340
rect 2261 5332 2265 5340
rect 2272 5332 2276 5340
rect 2280 5332 2284 5340
rect 2288 5332 2292 5340
rect 2296 5332 2300 5340
rect 2304 5332 2308 5340
rect 2312 5332 2316 5340
rect 1049 5284 1053 5292
rect 1064 5284 1068 5292
rect 1154 5284 1158 5292
rect 1169 5284 1173 5292
rect 1209 5286 1213 5294
rect 1217 5286 1221 5294
rect 1227 5286 1231 5294
rect 1244 5286 1248 5294
rect 1252 5286 1256 5294
rect 1260 5286 1264 5294
rect 1273 5286 1277 5294
rect 1282 5286 1286 5294
rect 1299 5286 1303 5294
rect 1316 5286 1320 5294
rect 1327 5286 1331 5294
rect 1335 5286 1339 5294
rect 1343 5286 1347 5294
rect 1351 5286 1355 5294
rect 1359 5286 1363 5294
rect 1367 5286 1371 5294
rect 1994 5284 1998 5292
rect 2009 5284 2013 5292
rect 2099 5284 2103 5292
rect 2114 5284 2118 5292
rect 2154 5286 2158 5294
rect 2162 5286 2166 5294
rect 2172 5286 2176 5294
rect 2189 5286 2193 5294
rect 2197 5286 2201 5294
rect 2205 5286 2209 5294
rect 2218 5286 2222 5294
rect 2227 5286 2231 5294
rect 2244 5286 2248 5294
rect 2261 5286 2265 5294
rect 2272 5286 2276 5294
rect 2280 5286 2284 5294
rect 2288 5286 2292 5294
rect 2296 5286 2300 5294
rect 2304 5286 2308 5294
rect 2312 5286 2316 5294
rect 1026 5187 1030 5195
rect 1034 5187 1038 5195
rect 1049 5193 1053 5201
rect 1064 5193 1068 5201
rect 1543 5219 1559 5249
rect 1563 5219 1579 5249
rect 1596 5219 1612 5249
rect 1616 5219 1632 5249
rect 1740 5216 1744 5224
rect 1748 5216 1752 5224
rect 1763 5222 1767 5230
rect 1778 5222 1782 5230
rect 1794 5216 1798 5224
rect 1802 5216 1806 5224
rect 1080 5187 1084 5195
rect 1088 5187 1092 5195
rect 1131 5187 1135 5195
rect 1139 5187 1143 5195
rect 1154 5193 1158 5201
rect 1169 5193 1173 5201
rect 1209 5200 1213 5208
rect 1217 5200 1221 5208
rect 1227 5200 1231 5208
rect 1244 5200 1248 5208
rect 1252 5200 1256 5208
rect 1260 5200 1264 5208
rect 1273 5200 1277 5208
rect 1282 5200 1286 5208
rect 1299 5200 1303 5208
rect 1316 5200 1320 5208
rect 1327 5200 1331 5208
rect 1335 5200 1339 5208
rect 1343 5200 1347 5208
rect 1351 5200 1355 5208
rect 1359 5200 1363 5208
rect 1367 5200 1371 5208
rect 1971 5187 1975 5195
rect 1979 5187 1983 5195
rect 1994 5193 1998 5201
rect 2009 5193 2013 5201
rect 2025 5187 2029 5195
rect 2033 5187 2037 5195
rect 2076 5187 2080 5195
rect 2084 5187 2088 5195
rect 2099 5193 2103 5201
rect 2114 5193 2118 5201
rect 2154 5200 2158 5208
rect 2162 5200 2166 5208
rect 2172 5200 2176 5208
rect 2189 5200 2193 5208
rect 2197 5200 2201 5208
rect 2205 5200 2209 5208
rect 2218 5200 2222 5208
rect 2227 5200 2231 5208
rect 2244 5200 2248 5208
rect 2261 5200 2265 5208
rect 2272 5200 2276 5208
rect 2280 5200 2284 5208
rect 2288 5200 2292 5208
rect 2296 5200 2300 5208
rect 2304 5200 2308 5208
rect 2312 5200 2316 5208
rect 1073 5153 1077 5161
rect 1088 5153 1092 5161
rect 1154 5153 1158 5161
rect 1169 5153 1173 5161
rect 1209 5154 1213 5162
rect 1217 5154 1221 5162
rect 1227 5154 1231 5162
rect 1244 5154 1248 5162
rect 1252 5154 1256 5162
rect 1260 5154 1264 5162
rect 1273 5154 1277 5162
rect 1282 5154 1286 5162
rect 1299 5154 1303 5162
rect 1316 5154 1320 5162
rect 1327 5154 1331 5162
rect 1335 5154 1339 5162
rect 1343 5154 1347 5162
rect 1351 5154 1355 5162
rect 1359 5154 1363 5162
rect 1367 5154 1371 5162
rect 2018 5153 2022 5161
rect 2033 5153 2037 5161
rect 2099 5153 2103 5161
rect 2114 5153 2118 5161
rect 2154 5154 2158 5162
rect 2162 5154 2166 5162
rect 2172 5154 2176 5162
rect 2189 5154 2193 5162
rect 2197 5154 2201 5162
rect 2205 5154 2209 5162
rect 2218 5154 2222 5162
rect 2227 5154 2231 5162
rect 2244 5154 2248 5162
rect 2261 5154 2265 5162
rect 2272 5154 2276 5162
rect 2280 5154 2284 5162
rect 2288 5154 2292 5162
rect 2296 5154 2300 5162
rect 2304 5154 2308 5162
rect 2312 5154 2316 5162
rect 1609 5119 1613 5127
rect 1622 5119 1626 5127
rect 1630 5119 1634 5127
rect 1638 5119 1642 5123
rect 1646 5119 1650 5127
rect 1659 5119 1663 5127
rect 1672 5119 1676 5127
rect 1680 5119 1684 5127
rect 1688 5119 1692 5127
rect 1696 5119 1700 5123
rect 1704 5119 1708 5127
rect 1717 5119 1721 5127
rect 1725 5119 1729 5127
rect 1733 5119 1737 5127
rect 2554 5119 2558 5127
rect 2567 5119 2571 5127
rect 2575 5119 2579 5127
rect 2583 5119 2587 5123
rect 2591 5119 2595 5127
rect 2604 5119 2608 5127
rect 2617 5119 2621 5127
rect 2625 5119 2629 5127
rect 2633 5119 2637 5127
rect 2641 5119 2645 5123
rect 2649 5119 2653 5127
rect 2662 5119 2666 5127
rect 2670 5119 2674 5127
rect 2678 5119 2682 5127
rect 1050 5055 1054 5063
rect 1058 5055 1062 5063
rect 1073 5061 1077 5069
rect 1088 5061 1092 5069
rect 1104 5055 1108 5063
rect 1112 5055 1116 5063
rect 1131 5055 1135 5063
rect 1139 5055 1143 5063
rect 1154 5061 1158 5069
rect 1169 5061 1173 5069
rect 1209 5068 1213 5076
rect 1217 5068 1221 5076
rect 1227 5068 1231 5076
rect 1244 5068 1248 5076
rect 1252 5068 1256 5076
rect 1260 5068 1264 5076
rect 1273 5068 1277 5076
rect 1282 5068 1286 5076
rect 1299 5068 1303 5076
rect 1316 5068 1320 5076
rect 1327 5068 1331 5076
rect 1335 5068 1339 5076
rect 1343 5068 1347 5076
rect 1351 5068 1355 5076
rect 1359 5068 1363 5076
rect 1367 5068 1371 5076
rect 1185 5055 1189 5063
rect 1193 5055 1197 5063
rect 1995 5055 1999 5063
rect 2003 5055 2007 5063
rect 2018 5061 2022 5069
rect 2033 5061 2037 5069
rect 2049 5055 2053 5063
rect 2057 5055 2061 5063
rect 2076 5055 2080 5063
rect 2084 5055 2088 5063
rect 2099 5061 2103 5069
rect 2114 5061 2118 5069
rect 2154 5068 2158 5076
rect 2162 5068 2166 5076
rect 2172 5068 2176 5076
rect 2189 5068 2193 5076
rect 2197 5068 2201 5076
rect 2205 5068 2209 5076
rect 2218 5068 2222 5076
rect 2227 5068 2231 5076
rect 2244 5068 2248 5076
rect 2261 5068 2265 5076
rect 2272 5068 2276 5076
rect 2280 5068 2284 5076
rect 2288 5068 2292 5076
rect 2296 5068 2300 5076
rect 2304 5068 2308 5076
rect 2312 5068 2316 5076
rect 2130 5055 2134 5063
rect 2138 5055 2142 5063
rect 1600 5017 1604 5025
rect 1608 5017 1612 5025
rect 1616 5017 1620 5025
rect 1629 5017 1633 5025
rect 1637 5017 1641 5021
rect 1645 5017 1649 5025
rect 1653 5017 1657 5025
rect 1661 5017 1665 5025
rect 1674 5017 1678 5025
rect 1687 5017 1691 5025
rect 1695 5017 1699 5021
rect 1703 5017 1707 5025
rect 1711 5017 1715 5025
rect 1724 5017 1728 5025
rect 2545 5017 2549 5025
rect 2553 5017 2557 5025
rect 2561 5017 2565 5025
rect 2574 5017 2578 5025
rect 2582 5017 2586 5021
rect 2590 5017 2594 5025
rect 2598 5017 2602 5025
rect 2606 5017 2610 5025
rect 2619 5017 2623 5025
rect 2632 5017 2636 5025
rect 2640 5017 2644 5021
rect 2648 5017 2652 5025
rect 2656 5017 2660 5025
rect 2669 5017 2673 5025
rect 852 4984 856 4992
rect 860 4984 864 4992
rect 868 4984 872 4992
rect 881 4984 885 4992
rect 889 4984 893 4988
rect 897 4984 901 4992
rect 905 4984 909 4992
rect 913 4984 917 4992
rect 926 4984 930 4992
rect 939 4984 943 4992
rect 947 4984 951 4988
rect 955 4984 959 4992
rect 963 4984 967 4992
rect 976 4984 980 4992
rect 984 4984 988 4992
rect 992 4984 996 4992
rect 1000 4984 1004 4992
rect 1013 4984 1017 4992
rect 1021 4984 1025 4988
rect 1029 4984 1033 4992
rect 1037 4984 1041 4992
rect 1045 4984 1049 4992
rect 1058 4984 1062 4992
rect 1071 4984 1075 4992
rect 1079 4984 1083 4988
rect 1087 4984 1091 4992
rect 1095 4984 1099 4992
rect 1108 4984 1112 4992
rect 1116 4984 1120 4992
rect 1124 4984 1128 4992
rect 1132 4984 1136 4992
rect 1145 4984 1149 4992
rect 1153 4984 1157 4988
rect 1161 4984 1165 4992
rect 1169 4984 1173 4992
rect 1177 4984 1181 4992
rect 1190 4984 1194 4992
rect 1203 4984 1207 4992
rect 1211 4984 1215 4988
rect 1219 4984 1223 4992
rect 1227 4984 1231 4992
rect 1240 4984 1244 4992
rect 1248 4984 1252 4992
rect 1256 4984 1260 4992
rect 1264 4984 1268 4992
rect 1277 4984 1281 4992
rect 1285 4984 1289 4988
rect 1293 4984 1297 4992
rect 1301 4984 1305 4992
rect 1309 4984 1313 4992
rect 1322 4984 1326 4992
rect 1335 4984 1339 4992
rect 1343 4984 1347 4988
rect 1351 4984 1355 4992
rect 1359 4984 1363 4992
rect 1372 4984 1376 4992
rect 1797 4984 1801 4992
rect 1805 4984 1809 4992
rect 1813 4984 1817 4992
rect 1826 4984 1830 4992
rect 1834 4984 1838 4988
rect 1842 4984 1846 4992
rect 1850 4984 1854 4992
rect 1858 4984 1862 4992
rect 1871 4984 1875 4992
rect 1884 4984 1888 4992
rect 1892 4984 1896 4988
rect 1900 4984 1904 4992
rect 1908 4984 1912 4992
rect 1921 4984 1925 4992
rect 1929 4984 1933 4992
rect 1937 4984 1941 4992
rect 1945 4984 1949 4992
rect 1958 4984 1962 4992
rect 1966 4984 1970 4988
rect 1974 4984 1978 4992
rect 1982 4984 1986 4992
rect 1990 4984 1994 4992
rect 2003 4984 2007 4992
rect 2016 4984 2020 4992
rect 2024 4984 2028 4988
rect 2032 4984 2036 4992
rect 2040 4984 2044 4992
rect 2053 4984 2057 4992
rect 2061 4984 2065 4992
rect 2069 4984 2073 4992
rect 2077 4984 2081 4992
rect 2090 4984 2094 4992
rect 2098 4984 2102 4988
rect 2106 4984 2110 4992
rect 2114 4984 2118 4992
rect 2122 4984 2126 4992
rect 2135 4984 2139 4992
rect 2148 4984 2152 4992
rect 2156 4984 2160 4988
rect 2164 4984 2168 4992
rect 2172 4984 2176 4992
rect 2185 4984 2189 4992
rect 2193 4984 2197 4992
rect 2201 4984 2205 4992
rect 2209 4984 2213 4992
rect 2222 4984 2226 4992
rect 2230 4984 2234 4988
rect 2238 4984 2242 4992
rect 2246 4984 2250 4992
rect 2254 4984 2258 4992
rect 2267 4984 2271 4992
rect 2280 4984 2284 4992
rect 2288 4984 2292 4988
rect 2296 4984 2300 4992
rect 2304 4984 2308 4992
rect 2317 4984 2321 4992
rect 4574 7928 4578 7945
rect 4574 7889 4578 7924
rect 4582 7889 4586 7945
rect 4590 7928 4594 7945
rect 4590 7889 4594 7924
rect 4598 7889 4602 7945
rect 4606 7928 4610 7945
rect 4606 7889 4610 7924
rect 4614 7889 4618 7945
rect 4622 7928 4626 7945
rect 4622 7889 4626 7924
rect 4637 7857 4641 7945
rect 4645 7928 4649 7936
rect 4645 7857 4649 7924
rect 4653 7857 4657 7945
rect 4661 7928 4665 7945
rect 4661 7857 4665 7924
rect 4680 7857 4684 7945
rect 4688 7928 4692 7936
rect 4688 7857 4692 7924
rect 4696 7857 4700 7945
rect 4704 7928 4708 7945
rect 4704 7857 4708 7924
rect 4721 7857 4725 7945
rect 4729 7928 4733 7936
rect 4729 7857 4733 7924
rect 4737 7857 4741 7945
rect 4745 7928 4749 7945
rect 4745 7857 4749 7924
rect 4572 7393 4576 7428
rect 4572 7372 4576 7389
rect 4580 7372 4584 7428
rect 4588 7393 4592 7428
rect 4588 7372 4592 7389
rect 4596 7372 4600 7428
rect 4604 7393 4608 7428
rect 4604 7372 4608 7389
rect 4612 7372 4616 7428
rect 4620 7393 4624 7428
rect 4620 7372 4624 7389
rect 4657 7301 4661 7305
rect 4667 7301 4671 7305
rect 4677 7301 4681 7305
rect 4687 7301 4691 7305
rect 4697 7301 4701 7305
rect 4707 7301 4711 7305
rect 4717 7301 4721 7305
rect 4727 7301 4731 7305
rect 4737 7301 4741 7305
rect 4662 7296 4666 7300
rect 4672 7296 4676 7300
rect 4682 7296 4686 7300
rect 4692 7296 4696 7300
rect 4702 7296 4706 7300
rect 4712 7296 4716 7300
rect 4722 7296 4726 7300
rect 4732 7296 4736 7300
rect 4742 7296 4746 7300
rect 4657 7291 4661 7295
rect 4667 7291 4671 7295
rect 4677 7291 4681 7295
rect 4687 7291 4691 7295
rect 4697 7291 4701 7295
rect 4707 7291 4711 7295
rect 4717 7291 4721 7295
rect 4727 7291 4731 7295
rect 4737 7291 4741 7295
rect 4662 7286 4666 7290
rect 4672 7286 4676 7290
rect 4682 7286 4686 7290
rect 4692 7286 4696 7290
rect 4702 7286 4706 7290
rect 4712 7286 4716 7290
rect 4722 7286 4726 7290
rect 4732 7286 4736 7290
rect 4742 7286 4746 7290
rect 4657 7281 4661 7285
rect 4667 7281 4671 7285
rect 4677 7281 4681 7285
rect 4687 7281 4691 7285
rect 4697 7281 4701 7285
rect 4707 7281 4711 7285
rect 4717 7281 4721 7285
rect 4727 7281 4731 7285
rect 4737 7281 4741 7285
rect 4662 7276 4666 7280
rect 4672 7276 4676 7280
rect 4682 7276 4686 7280
rect 4692 7276 4696 7280
rect 4702 7276 4706 7280
rect 4712 7276 4716 7280
rect 4722 7276 4726 7280
rect 4732 7276 4736 7280
rect 4742 7276 4746 7280
rect 4657 7271 4661 7275
rect 4667 7271 4671 7275
rect 4677 7271 4681 7275
rect 4687 7271 4691 7275
rect 4697 7271 4701 7275
rect 4707 7271 4711 7275
rect 4717 7271 4721 7275
rect 4727 7271 4731 7275
rect 4737 7271 4741 7275
rect 4662 7266 4666 7270
rect 4672 7266 4676 7270
rect 4682 7266 4686 7270
rect 4692 7266 4696 7270
rect 4702 7266 4706 7270
rect 4712 7266 4716 7270
rect 4722 7266 4726 7270
rect 4732 7266 4736 7270
rect 4742 7266 4746 7270
rect 4657 7261 4661 7265
rect 4667 7261 4671 7265
rect 4677 7261 4681 7265
rect 4687 7261 4691 7265
rect 4697 7261 4701 7265
rect 4707 7261 4711 7265
rect 4717 7261 4721 7265
rect 4727 7261 4731 7265
rect 4737 7261 4741 7265
rect 1210 4531 1227 4535
rect 1231 4531 1266 4535
rect 2137 4531 2154 4535
rect 2158 4531 2193 4535
rect 2446 4531 2463 4535
rect 2467 4531 2502 4535
rect 2755 4531 2772 4535
rect 2776 4531 2811 4535
rect 3064 4531 3081 4535
rect 3085 4531 3120 4535
rect 3373 4531 3390 4535
rect 3394 4531 3429 4535
rect 1210 4523 1266 4527
rect 1210 4515 1227 4519
rect 1231 4515 1266 4519
rect 1210 4507 1266 4511
rect 2137 4523 2193 4527
rect 2137 4515 2154 4519
rect 2158 4515 2193 4519
rect 2137 4507 2193 4511
rect 1210 4499 1227 4503
rect 1231 4499 1266 4503
rect 2446 4523 2502 4527
rect 2446 4515 2463 4519
rect 2467 4515 2502 4519
rect 2446 4507 2502 4511
rect 2137 4499 2154 4503
rect 2158 4499 2193 4503
rect 2755 4523 2811 4527
rect 2755 4515 2772 4519
rect 2776 4515 2811 4519
rect 2755 4507 2811 4511
rect 2446 4499 2463 4503
rect 2467 4499 2502 4503
rect 3064 4523 3120 4527
rect 3064 4515 3081 4519
rect 3085 4515 3120 4519
rect 3064 4507 3120 4511
rect 2755 4499 2772 4503
rect 2776 4499 2811 4503
rect 3373 4523 3429 4527
rect 3373 4515 3390 4519
rect 3394 4515 3429 4519
rect 3373 4507 3429 4511
rect 3064 4499 3081 4503
rect 3085 4499 3120 4503
rect 3373 4499 3390 4503
rect 3394 4499 3429 4503
rect 1210 4491 1266 4495
rect 2137 4491 2193 4495
rect 2446 4491 2502 4495
rect 2755 4491 2811 4495
rect 3064 4491 3120 4495
rect 3373 4491 3429 4495
rect 1210 4483 1227 4487
rect 1231 4483 1266 4487
rect 2137 4483 2154 4487
rect 2158 4483 2193 4487
rect 2446 4483 2463 4487
rect 2467 4483 2502 4487
rect 2755 4483 2772 4487
rect 2776 4483 2811 4487
rect 3064 4483 3081 4487
rect 3085 4483 3120 4487
rect 3373 4483 3390 4487
rect 3394 4483 3429 4487
rect 1099 4446 1103 4450
rect 1109 4446 1113 4450
rect 1119 4446 1123 4450
rect 1129 4446 1133 4450
rect 1139 4446 1143 4450
rect 1104 4441 1108 4445
rect 1114 4441 1118 4445
rect 1124 4441 1128 4445
rect 1134 4441 1138 4445
rect 1099 4436 1103 4440
rect 1109 4436 1113 4440
rect 1119 4436 1123 4440
rect 1129 4436 1133 4440
rect 1139 4436 1143 4440
rect 1104 4431 1108 4435
rect 1114 4431 1118 4435
rect 1124 4431 1128 4435
rect 1134 4431 1138 4435
rect 1099 4426 1103 4430
rect 1109 4426 1113 4430
rect 1119 4426 1123 4430
rect 1129 4426 1133 4430
rect 1139 4426 1143 4430
rect 1104 4421 1108 4425
rect 1114 4421 1118 4425
rect 1124 4421 1128 4425
rect 1134 4421 1138 4425
rect 1099 4416 1103 4420
rect 1109 4416 1113 4420
rect 1119 4416 1123 4420
rect 1129 4416 1133 4420
rect 1139 4416 1143 4420
rect 1104 4411 1108 4415
rect 1114 4411 1118 4415
rect 1124 4411 1128 4415
rect 1134 4411 1138 4415
rect 1099 4406 1103 4410
rect 1109 4406 1113 4410
rect 1119 4406 1123 4410
rect 1129 4406 1133 4410
rect 1139 4406 1143 4410
rect 1104 4401 1108 4405
rect 1114 4401 1118 4405
rect 1124 4401 1128 4405
rect 1134 4401 1138 4405
rect 1099 4396 1103 4400
rect 1109 4396 1113 4400
rect 1119 4396 1123 4400
rect 1129 4396 1133 4400
rect 1139 4396 1143 4400
rect 1104 4391 1108 4395
rect 1114 4391 1118 4395
rect 1124 4391 1128 4395
rect 1134 4391 1138 4395
rect 1099 4386 1103 4390
rect 1109 4386 1113 4390
rect 1119 4386 1123 4390
rect 1129 4386 1133 4390
rect 1139 4386 1143 4390
rect 1104 4381 1108 4385
rect 1114 4381 1118 4385
rect 1124 4381 1128 4385
rect 1134 4381 1138 4385
rect 1099 4376 1103 4380
rect 1109 4376 1113 4380
rect 1119 4376 1123 4380
rect 1129 4376 1133 4380
rect 1139 4376 1143 4380
rect 1104 4371 1108 4375
rect 1114 4371 1118 4375
rect 1124 4371 1128 4375
rect 1134 4371 1138 4375
rect 1099 4366 1103 4370
rect 1109 4366 1113 4370
rect 1119 4366 1123 4370
rect 1129 4366 1133 4370
rect 1139 4366 1143 4370
rect 1104 4361 1108 4365
rect 1114 4361 1118 4365
rect 1124 4361 1128 4365
rect 1134 4361 1138 4365
rect 1408 4446 1412 4450
rect 1418 4446 1422 4450
rect 1428 4446 1432 4450
rect 1438 4446 1442 4450
rect 1448 4446 1452 4450
rect 1413 4441 1417 4445
rect 1423 4441 1427 4445
rect 1433 4441 1437 4445
rect 1443 4441 1447 4445
rect 1408 4436 1412 4440
rect 1418 4436 1422 4440
rect 1428 4436 1432 4440
rect 1438 4436 1442 4440
rect 1448 4436 1452 4440
rect 1413 4431 1417 4435
rect 1423 4431 1427 4435
rect 1433 4431 1437 4435
rect 1443 4431 1447 4435
rect 1408 4426 1412 4430
rect 1418 4426 1422 4430
rect 1428 4426 1432 4430
rect 1438 4426 1442 4430
rect 1448 4426 1452 4430
rect 1413 4421 1417 4425
rect 1423 4421 1427 4425
rect 1433 4421 1437 4425
rect 1443 4421 1447 4425
rect 1408 4416 1412 4420
rect 1418 4416 1422 4420
rect 1428 4416 1432 4420
rect 1438 4416 1442 4420
rect 1448 4416 1452 4420
rect 1413 4411 1417 4415
rect 1423 4411 1427 4415
rect 1433 4411 1437 4415
rect 1443 4411 1447 4415
rect 1408 4406 1412 4410
rect 1418 4406 1422 4410
rect 1428 4406 1432 4410
rect 1438 4406 1442 4410
rect 1448 4406 1452 4410
rect 1413 4401 1417 4405
rect 1423 4401 1427 4405
rect 1433 4401 1437 4405
rect 1443 4401 1447 4405
rect 1408 4396 1412 4400
rect 1418 4396 1422 4400
rect 1428 4396 1432 4400
rect 1438 4396 1442 4400
rect 1448 4396 1452 4400
rect 1413 4391 1417 4395
rect 1423 4391 1427 4395
rect 1433 4391 1437 4395
rect 1443 4391 1447 4395
rect 1408 4386 1412 4390
rect 1418 4386 1422 4390
rect 1428 4386 1432 4390
rect 1438 4386 1442 4390
rect 1448 4386 1452 4390
rect 1413 4381 1417 4385
rect 1423 4381 1427 4385
rect 1433 4381 1437 4385
rect 1443 4381 1447 4385
rect 1408 4376 1412 4380
rect 1418 4376 1422 4380
rect 1428 4376 1432 4380
rect 1438 4376 1442 4380
rect 1448 4376 1452 4380
rect 1413 4371 1417 4375
rect 1423 4371 1427 4375
rect 1433 4371 1437 4375
rect 1443 4371 1447 4375
rect 1408 4366 1412 4370
rect 1418 4366 1422 4370
rect 1428 4366 1432 4370
rect 1438 4366 1442 4370
rect 1448 4366 1452 4370
rect 1413 4361 1417 4365
rect 1423 4361 1427 4365
rect 1433 4361 1437 4365
rect 1443 4361 1447 4365
rect 1717 4446 1721 4450
rect 1727 4446 1731 4450
rect 1737 4446 1741 4450
rect 1747 4446 1751 4450
rect 1757 4446 1761 4450
rect 1722 4441 1726 4445
rect 1732 4441 1736 4445
rect 1742 4441 1746 4445
rect 1752 4441 1756 4445
rect 1717 4436 1721 4440
rect 1727 4436 1731 4440
rect 1737 4436 1741 4440
rect 1747 4436 1751 4440
rect 1757 4436 1761 4440
rect 1722 4431 1726 4435
rect 1732 4431 1736 4435
rect 1742 4431 1746 4435
rect 1752 4431 1756 4435
rect 1717 4426 1721 4430
rect 1727 4426 1731 4430
rect 1737 4426 1741 4430
rect 1747 4426 1751 4430
rect 1757 4426 1761 4430
rect 1722 4421 1726 4425
rect 1732 4421 1736 4425
rect 1742 4421 1746 4425
rect 1752 4421 1756 4425
rect 1717 4416 1721 4420
rect 1727 4416 1731 4420
rect 1737 4416 1741 4420
rect 1747 4416 1751 4420
rect 1757 4416 1761 4420
rect 1722 4411 1726 4415
rect 1732 4411 1736 4415
rect 1742 4411 1746 4415
rect 1752 4411 1756 4415
rect 1717 4406 1721 4410
rect 1727 4406 1731 4410
rect 1737 4406 1741 4410
rect 1747 4406 1751 4410
rect 1757 4406 1761 4410
rect 1722 4401 1726 4405
rect 1732 4401 1736 4405
rect 1742 4401 1746 4405
rect 1752 4401 1756 4405
rect 1717 4396 1721 4400
rect 1727 4396 1731 4400
rect 1737 4396 1741 4400
rect 1747 4396 1751 4400
rect 1757 4396 1761 4400
rect 1722 4391 1726 4395
rect 1732 4391 1736 4395
rect 1742 4391 1746 4395
rect 1752 4391 1756 4395
rect 1717 4386 1721 4390
rect 1727 4386 1731 4390
rect 1737 4386 1741 4390
rect 1747 4386 1751 4390
rect 1757 4386 1761 4390
rect 1722 4381 1726 4385
rect 1732 4381 1736 4385
rect 1742 4381 1746 4385
rect 1752 4381 1756 4385
rect 1717 4376 1721 4380
rect 1727 4376 1731 4380
rect 1737 4376 1741 4380
rect 1747 4376 1751 4380
rect 1757 4376 1761 4380
rect 1722 4371 1726 4375
rect 1732 4371 1736 4375
rect 1742 4371 1746 4375
rect 1752 4371 1756 4375
rect 1717 4366 1721 4370
rect 1727 4366 1731 4370
rect 1737 4366 1741 4370
rect 1747 4366 1751 4370
rect 1757 4366 1761 4370
rect 1722 4361 1726 4365
rect 1732 4361 1736 4365
rect 1742 4361 1746 4365
rect 1752 4361 1756 4365
rect 2026 4446 2030 4450
rect 2036 4446 2040 4450
rect 2046 4446 2050 4450
rect 2056 4446 2060 4450
rect 2066 4446 2070 4450
rect 2031 4441 2035 4445
rect 2041 4441 2045 4445
rect 2051 4441 2055 4445
rect 2061 4441 2065 4445
rect 2026 4436 2030 4440
rect 2036 4436 2040 4440
rect 2046 4436 2050 4440
rect 2056 4436 2060 4440
rect 2066 4436 2070 4440
rect 2031 4431 2035 4435
rect 2041 4431 2045 4435
rect 2051 4431 2055 4435
rect 2061 4431 2065 4435
rect 2026 4426 2030 4430
rect 2036 4426 2040 4430
rect 2046 4426 2050 4430
rect 2056 4426 2060 4430
rect 2066 4426 2070 4430
rect 2031 4421 2035 4425
rect 2041 4421 2045 4425
rect 2051 4421 2055 4425
rect 2061 4421 2065 4425
rect 2026 4416 2030 4420
rect 2036 4416 2040 4420
rect 2046 4416 2050 4420
rect 2056 4416 2060 4420
rect 2066 4416 2070 4420
rect 2031 4411 2035 4415
rect 2041 4411 2045 4415
rect 2051 4411 2055 4415
rect 2061 4411 2065 4415
rect 2026 4406 2030 4410
rect 2036 4406 2040 4410
rect 2046 4406 2050 4410
rect 2056 4406 2060 4410
rect 2066 4406 2070 4410
rect 2031 4401 2035 4405
rect 2041 4401 2045 4405
rect 2051 4401 2055 4405
rect 2061 4401 2065 4405
rect 2026 4396 2030 4400
rect 2036 4396 2040 4400
rect 2046 4396 2050 4400
rect 2056 4396 2060 4400
rect 2066 4396 2070 4400
rect 2031 4391 2035 4395
rect 2041 4391 2045 4395
rect 2051 4391 2055 4395
rect 2061 4391 2065 4395
rect 2026 4386 2030 4390
rect 2036 4386 2040 4390
rect 2046 4386 2050 4390
rect 2056 4386 2060 4390
rect 2066 4386 2070 4390
rect 2031 4381 2035 4385
rect 2041 4381 2045 4385
rect 2051 4381 2055 4385
rect 2061 4381 2065 4385
rect 2026 4376 2030 4380
rect 2036 4376 2040 4380
rect 2046 4376 2050 4380
rect 2056 4376 2060 4380
rect 2066 4376 2070 4380
rect 2031 4371 2035 4375
rect 2041 4371 2045 4375
rect 2051 4371 2055 4375
rect 2061 4371 2065 4375
rect 2026 4366 2030 4370
rect 2036 4366 2040 4370
rect 2046 4366 2050 4370
rect 2056 4366 2060 4370
rect 2066 4366 2070 4370
rect 2031 4361 2035 4365
rect 2041 4361 2045 4365
rect 2051 4361 2055 4365
rect 2061 4361 2065 4365
rect 2335 4446 2339 4450
rect 2345 4446 2349 4450
rect 2355 4446 2359 4450
rect 2365 4446 2369 4450
rect 2375 4446 2379 4450
rect 2340 4441 2344 4445
rect 2350 4441 2354 4445
rect 2360 4441 2364 4445
rect 2370 4441 2374 4445
rect 2335 4436 2339 4440
rect 2345 4436 2349 4440
rect 2355 4436 2359 4440
rect 2365 4436 2369 4440
rect 2375 4436 2379 4440
rect 2340 4431 2344 4435
rect 2350 4431 2354 4435
rect 2360 4431 2364 4435
rect 2370 4431 2374 4435
rect 2335 4426 2339 4430
rect 2345 4426 2349 4430
rect 2355 4426 2359 4430
rect 2365 4426 2369 4430
rect 2375 4426 2379 4430
rect 2340 4421 2344 4425
rect 2350 4421 2354 4425
rect 2360 4421 2364 4425
rect 2370 4421 2374 4425
rect 2335 4416 2339 4420
rect 2345 4416 2349 4420
rect 2355 4416 2359 4420
rect 2365 4416 2369 4420
rect 2375 4416 2379 4420
rect 2340 4411 2344 4415
rect 2350 4411 2354 4415
rect 2360 4411 2364 4415
rect 2370 4411 2374 4415
rect 2335 4406 2339 4410
rect 2345 4406 2349 4410
rect 2355 4406 2359 4410
rect 2365 4406 2369 4410
rect 2375 4406 2379 4410
rect 2340 4401 2344 4405
rect 2350 4401 2354 4405
rect 2360 4401 2364 4405
rect 2370 4401 2374 4405
rect 2335 4396 2339 4400
rect 2345 4396 2349 4400
rect 2355 4396 2359 4400
rect 2365 4396 2369 4400
rect 2375 4396 2379 4400
rect 2340 4391 2344 4395
rect 2350 4391 2354 4395
rect 2360 4391 2364 4395
rect 2370 4391 2374 4395
rect 2335 4386 2339 4390
rect 2345 4386 2349 4390
rect 2355 4386 2359 4390
rect 2365 4386 2369 4390
rect 2375 4386 2379 4390
rect 2340 4381 2344 4385
rect 2350 4381 2354 4385
rect 2360 4381 2364 4385
rect 2370 4381 2374 4385
rect 2335 4376 2339 4380
rect 2345 4376 2349 4380
rect 2355 4376 2359 4380
rect 2365 4376 2369 4380
rect 2375 4376 2379 4380
rect 2340 4371 2344 4375
rect 2350 4371 2354 4375
rect 2360 4371 2364 4375
rect 2370 4371 2374 4375
rect 2335 4366 2339 4370
rect 2345 4366 2349 4370
rect 2355 4366 2359 4370
rect 2365 4366 2369 4370
rect 2375 4366 2379 4370
rect 2340 4361 2344 4365
rect 2350 4361 2354 4365
rect 2360 4361 2364 4365
rect 2370 4361 2374 4365
rect 2644 4446 2648 4450
rect 2654 4446 2658 4450
rect 2664 4446 2668 4450
rect 2674 4446 2678 4450
rect 2684 4446 2688 4450
rect 2649 4441 2653 4445
rect 2659 4441 2663 4445
rect 2669 4441 2673 4445
rect 2679 4441 2683 4445
rect 2644 4436 2648 4440
rect 2654 4436 2658 4440
rect 2664 4436 2668 4440
rect 2674 4436 2678 4440
rect 2684 4436 2688 4440
rect 2649 4431 2653 4435
rect 2659 4431 2663 4435
rect 2669 4431 2673 4435
rect 2679 4431 2683 4435
rect 2644 4426 2648 4430
rect 2654 4426 2658 4430
rect 2664 4426 2668 4430
rect 2674 4426 2678 4430
rect 2684 4426 2688 4430
rect 2649 4421 2653 4425
rect 2659 4421 2663 4425
rect 2669 4421 2673 4425
rect 2679 4421 2683 4425
rect 2644 4416 2648 4420
rect 2654 4416 2658 4420
rect 2664 4416 2668 4420
rect 2674 4416 2678 4420
rect 2684 4416 2688 4420
rect 2649 4411 2653 4415
rect 2659 4411 2663 4415
rect 2669 4411 2673 4415
rect 2679 4411 2683 4415
rect 2644 4406 2648 4410
rect 2654 4406 2658 4410
rect 2664 4406 2668 4410
rect 2674 4406 2678 4410
rect 2684 4406 2688 4410
rect 2649 4401 2653 4405
rect 2659 4401 2663 4405
rect 2669 4401 2673 4405
rect 2679 4401 2683 4405
rect 2644 4396 2648 4400
rect 2654 4396 2658 4400
rect 2664 4396 2668 4400
rect 2674 4396 2678 4400
rect 2684 4396 2688 4400
rect 2649 4391 2653 4395
rect 2659 4391 2663 4395
rect 2669 4391 2673 4395
rect 2679 4391 2683 4395
rect 2644 4386 2648 4390
rect 2654 4386 2658 4390
rect 2664 4386 2668 4390
rect 2674 4386 2678 4390
rect 2684 4386 2688 4390
rect 2649 4381 2653 4385
rect 2659 4381 2663 4385
rect 2669 4381 2673 4385
rect 2679 4381 2683 4385
rect 2644 4376 2648 4380
rect 2654 4376 2658 4380
rect 2664 4376 2668 4380
rect 2674 4376 2678 4380
rect 2684 4376 2688 4380
rect 2649 4371 2653 4375
rect 2659 4371 2663 4375
rect 2669 4371 2673 4375
rect 2679 4371 2683 4375
rect 2644 4366 2648 4370
rect 2654 4366 2658 4370
rect 2664 4366 2668 4370
rect 2674 4366 2678 4370
rect 2684 4366 2688 4370
rect 2649 4361 2653 4365
rect 2659 4361 2663 4365
rect 2669 4361 2673 4365
rect 2679 4361 2683 4365
rect 2953 4446 2957 4450
rect 2963 4446 2967 4450
rect 2973 4446 2977 4450
rect 2983 4446 2987 4450
rect 2993 4446 2997 4450
rect 2958 4441 2962 4445
rect 2968 4441 2972 4445
rect 2978 4441 2982 4445
rect 2988 4441 2992 4445
rect 2953 4436 2957 4440
rect 2963 4436 2967 4440
rect 2973 4436 2977 4440
rect 2983 4436 2987 4440
rect 2993 4436 2997 4440
rect 2958 4431 2962 4435
rect 2968 4431 2972 4435
rect 2978 4431 2982 4435
rect 2988 4431 2992 4435
rect 2953 4426 2957 4430
rect 2963 4426 2967 4430
rect 2973 4426 2977 4430
rect 2983 4426 2987 4430
rect 2993 4426 2997 4430
rect 2958 4421 2962 4425
rect 2968 4421 2972 4425
rect 2978 4421 2982 4425
rect 2988 4421 2992 4425
rect 2953 4416 2957 4420
rect 2963 4416 2967 4420
rect 2973 4416 2977 4420
rect 2983 4416 2987 4420
rect 2993 4416 2997 4420
rect 2958 4411 2962 4415
rect 2968 4411 2972 4415
rect 2978 4411 2982 4415
rect 2988 4411 2992 4415
rect 2953 4406 2957 4410
rect 2963 4406 2967 4410
rect 2973 4406 2977 4410
rect 2983 4406 2987 4410
rect 2993 4406 2997 4410
rect 2958 4401 2962 4405
rect 2968 4401 2972 4405
rect 2978 4401 2982 4405
rect 2988 4401 2992 4405
rect 2953 4396 2957 4400
rect 2963 4396 2967 4400
rect 2973 4396 2977 4400
rect 2983 4396 2987 4400
rect 2993 4396 2997 4400
rect 2958 4391 2962 4395
rect 2968 4391 2972 4395
rect 2978 4391 2982 4395
rect 2988 4391 2992 4395
rect 2953 4386 2957 4390
rect 2963 4386 2967 4390
rect 2973 4386 2977 4390
rect 2983 4386 2987 4390
rect 2993 4386 2997 4390
rect 2958 4381 2962 4385
rect 2968 4381 2972 4385
rect 2978 4381 2982 4385
rect 2988 4381 2992 4385
rect 2953 4376 2957 4380
rect 2963 4376 2967 4380
rect 2973 4376 2977 4380
rect 2983 4376 2987 4380
rect 2993 4376 2997 4380
rect 2958 4371 2962 4375
rect 2968 4371 2972 4375
rect 2978 4371 2982 4375
rect 2988 4371 2992 4375
rect 2953 4366 2957 4370
rect 2963 4366 2967 4370
rect 2973 4366 2977 4370
rect 2983 4366 2987 4370
rect 2993 4366 2997 4370
rect 2958 4361 2962 4365
rect 2968 4361 2972 4365
rect 2978 4361 2982 4365
rect 2988 4361 2992 4365
rect 3262 4446 3266 4450
rect 3272 4446 3276 4450
rect 3282 4446 3286 4450
rect 3292 4446 3296 4450
rect 3302 4446 3306 4450
rect 3267 4441 3271 4445
rect 3277 4441 3281 4445
rect 3287 4441 3291 4445
rect 3297 4441 3301 4445
rect 3262 4436 3266 4440
rect 3272 4436 3276 4440
rect 3282 4436 3286 4440
rect 3292 4436 3296 4440
rect 3302 4436 3306 4440
rect 3267 4431 3271 4435
rect 3277 4431 3281 4435
rect 3287 4431 3291 4435
rect 3297 4431 3301 4435
rect 3262 4426 3266 4430
rect 3272 4426 3276 4430
rect 3282 4426 3286 4430
rect 3292 4426 3296 4430
rect 3302 4426 3306 4430
rect 3267 4421 3271 4425
rect 3277 4421 3281 4425
rect 3287 4421 3291 4425
rect 3297 4421 3301 4425
rect 3262 4416 3266 4420
rect 3272 4416 3276 4420
rect 3282 4416 3286 4420
rect 3292 4416 3296 4420
rect 3302 4416 3306 4420
rect 3267 4411 3271 4415
rect 3277 4411 3281 4415
rect 3287 4411 3291 4415
rect 3297 4411 3301 4415
rect 3262 4406 3266 4410
rect 3272 4406 3276 4410
rect 3282 4406 3286 4410
rect 3292 4406 3296 4410
rect 3302 4406 3306 4410
rect 3267 4401 3271 4405
rect 3277 4401 3281 4405
rect 3287 4401 3291 4405
rect 3297 4401 3301 4405
rect 3262 4396 3266 4400
rect 3272 4396 3276 4400
rect 3282 4396 3286 4400
rect 3292 4396 3296 4400
rect 3302 4396 3306 4400
rect 3267 4391 3271 4395
rect 3277 4391 3281 4395
rect 3287 4391 3291 4395
rect 3297 4391 3301 4395
rect 3262 4386 3266 4390
rect 3272 4386 3276 4390
rect 3282 4386 3286 4390
rect 3292 4386 3296 4390
rect 3302 4386 3306 4390
rect 3267 4381 3271 4385
rect 3277 4381 3281 4385
rect 3287 4381 3291 4385
rect 3297 4381 3301 4385
rect 3262 4376 3266 4380
rect 3272 4376 3276 4380
rect 3282 4376 3286 4380
rect 3292 4376 3296 4380
rect 3302 4376 3306 4380
rect 3267 4371 3271 4375
rect 3277 4371 3281 4375
rect 3287 4371 3291 4375
rect 3297 4371 3301 4375
rect 3262 4366 3266 4370
rect 3272 4366 3276 4370
rect 3282 4366 3286 4370
rect 3292 4366 3296 4370
rect 3302 4366 3306 4370
rect 3267 4361 3271 4365
rect 3277 4361 3281 4365
rect 3287 4361 3291 4365
rect 3297 4361 3301 4365
rect 3571 4446 3575 4450
rect 3581 4446 3585 4450
rect 3591 4446 3595 4450
rect 3601 4446 3605 4450
rect 3611 4446 3615 4450
rect 3576 4441 3580 4445
rect 3586 4441 3590 4445
rect 3596 4441 3600 4445
rect 3606 4441 3610 4445
rect 3571 4436 3575 4440
rect 3581 4436 3585 4440
rect 3591 4436 3595 4440
rect 3601 4436 3605 4440
rect 3611 4436 3615 4440
rect 3576 4431 3580 4435
rect 3586 4431 3590 4435
rect 3596 4431 3600 4435
rect 3606 4431 3610 4435
rect 3571 4426 3575 4430
rect 3581 4426 3585 4430
rect 3591 4426 3595 4430
rect 3601 4426 3605 4430
rect 3611 4426 3615 4430
rect 3576 4421 3580 4425
rect 3586 4421 3590 4425
rect 3596 4421 3600 4425
rect 3606 4421 3610 4425
rect 3571 4416 3575 4420
rect 3581 4416 3585 4420
rect 3591 4416 3595 4420
rect 3601 4416 3605 4420
rect 3611 4416 3615 4420
rect 3576 4411 3580 4415
rect 3586 4411 3590 4415
rect 3596 4411 3600 4415
rect 3606 4411 3610 4415
rect 3571 4406 3575 4410
rect 3581 4406 3585 4410
rect 3591 4406 3595 4410
rect 3601 4406 3605 4410
rect 3611 4406 3615 4410
rect 3576 4401 3580 4405
rect 3586 4401 3590 4405
rect 3596 4401 3600 4405
rect 3606 4401 3610 4405
rect 3571 4396 3575 4400
rect 3581 4396 3585 4400
rect 3591 4396 3595 4400
rect 3601 4396 3605 4400
rect 3611 4396 3615 4400
rect 3576 4391 3580 4395
rect 3586 4391 3590 4395
rect 3596 4391 3600 4395
rect 3606 4391 3610 4395
rect 3571 4386 3575 4390
rect 3581 4386 3585 4390
rect 3591 4386 3595 4390
rect 3601 4386 3605 4390
rect 3611 4386 3615 4390
rect 3576 4381 3580 4385
rect 3586 4381 3590 4385
rect 3596 4381 3600 4385
rect 3606 4381 3610 4385
rect 3571 4376 3575 4380
rect 3581 4376 3585 4380
rect 3591 4376 3595 4380
rect 3601 4376 3605 4380
rect 3611 4376 3615 4380
rect 3576 4371 3580 4375
rect 3586 4371 3590 4375
rect 3596 4371 3600 4375
rect 3606 4371 3610 4375
rect 3571 4366 3575 4370
rect 3581 4366 3585 4370
rect 3591 4366 3595 4370
rect 3601 4366 3605 4370
rect 3611 4366 3615 4370
rect 3576 4361 3580 4365
rect 3586 4361 3590 4365
rect 3596 4361 3600 4365
rect 3606 4361 3610 4365
<< psubstratepdiff >>
rect 1383 9965 1455 9967
rect 1383 9961 1385 9965
rect 1389 9961 1392 9965
rect 1396 9961 1397 9965
rect 1401 9961 1402 9965
rect 1406 9961 1407 9965
rect 1411 9961 1412 9965
rect 1416 9961 1417 9965
rect 1421 9961 1422 9965
rect 1426 9961 1427 9965
rect 1431 9961 1432 9965
rect 1436 9961 1437 9965
rect 1441 9961 1442 9965
rect 1446 9961 1449 9965
rect 1453 9961 1455 9965
rect 1383 9959 1455 9961
rect 1383 9958 1391 9959
rect 1383 9954 1385 9958
rect 1389 9954 1391 9958
rect 1383 9953 1391 9954
rect 1447 9958 1455 9959
rect 1447 9954 1449 9958
rect 1453 9954 1455 9958
rect 1447 9953 1455 9954
rect 1383 9949 1385 9953
rect 1389 9949 1391 9953
rect 1383 9948 1391 9949
rect 1383 9944 1385 9948
rect 1389 9944 1391 9948
rect 1383 9943 1391 9944
rect 1383 9939 1385 9943
rect 1389 9939 1391 9943
rect 1383 9938 1391 9939
rect 1383 9934 1385 9938
rect 1389 9934 1391 9938
rect 1383 9933 1391 9934
rect 1383 9929 1385 9933
rect 1389 9929 1391 9933
rect 1383 9928 1391 9929
rect 1383 9924 1385 9928
rect 1389 9924 1391 9928
rect 1383 9923 1391 9924
rect 1383 9919 1385 9923
rect 1389 9919 1391 9923
rect 1383 9918 1391 9919
rect 1383 9914 1385 9918
rect 1389 9914 1391 9918
rect 1383 9913 1391 9914
rect 1383 9909 1385 9913
rect 1389 9909 1391 9913
rect 1383 9908 1391 9909
rect 1383 9904 1385 9908
rect 1389 9904 1391 9908
rect 1383 9903 1391 9904
rect 1383 9899 1385 9903
rect 1389 9899 1391 9903
rect 1383 9898 1391 9899
rect 1383 9894 1385 9898
rect 1389 9894 1391 9898
rect 1383 9893 1391 9894
rect 1383 9889 1385 9893
rect 1389 9889 1391 9893
rect 1383 9888 1391 9889
rect 1383 9884 1385 9888
rect 1389 9884 1391 9888
rect 1383 9883 1391 9884
rect 1383 9879 1385 9883
rect 1389 9879 1391 9883
rect 1383 9878 1391 9879
rect 1383 9874 1385 9878
rect 1389 9874 1391 9878
rect 1383 9873 1391 9874
rect 1383 9869 1385 9873
rect 1389 9869 1391 9873
rect 1383 9868 1391 9869
rect 1383 9864 1385 9868
rect 1389 9864 1391 9868
rect 1447 9949 1449 9953
rect 1453 9949 1455 9953
rect 1447 9948 1455 9949
rect 1447 9944 1449 9948
rect 1453 9944 1455 9948
rect 1447 9943 1455 9944
rect 1447 9939 1449 9943
rect 1453 9939 1455 9943
rect 1447 9938 1455 9939
rect 1447 9934 1449 9938
rect 1453 9934 1455 9938
rect 1447 9933 1455 9934
rect 1447 9929 1449 9933
rect 1453 9929 1455 9933
rect 1447 9928 1455 9929
rect 1447 9924 1449 9928
rect 1453 9924 1455 9928
rect 1447 9923 1455 9924
rect 1447 9919 1449 9923
rect 1453 9919 1455 9923
rect 1447 9918 1455 9919
rect 1447 9914 1449 9918
rect 1453 9914 1455 9918
rect 1447 9913 1455 9914
rect 1447 9909 1449 9913
rect 1453 9909 1455 9913
rect 1447 9908 1455 9909
rect 1447 9904 1449 9908
rect 1453 9904 1455 9908
rect 1447 9903 1455 9904
rect 1447 9899 1449 9903
rect 1453 9899 1455 9903
rect 1447 9898 1455 9899
rect 1447 9894 1449 9898
rect 1453 9894 1455 9898
rect 1447 9893 1455 9894
rect 1447 9889 1449 9893
rect 1453 9889 1455 9893
rect 1447 9888 1455 9889
rect 1447 9884 1449 9888
rect 1453 9884 1455 9888
rect 1447 9883 1455 9884
rect 1447 9879 1449 9883
rect 1453 9879 1455 9883
rect 1447 9878 1455 9879
rect 1447 9874 1449 9878
rect 1453 9874 1455 9878
rect 1447 9873 1455 9874
rect 1447 9869 1449 9873
rect 1453 9869 1455 9873
rect 1447 9868 1455 9869
rect 1447 9864 1449 9868
rect 1453 9864 1455 9868
rect 1383 9863 1391 9864
rect 1383 9859 1385 9863
rect 1389 9859 1391 9863
rect 1383 9858 1391 9859
rect 1447 9863 1455 9864
rect 1447 9859 1449 9863
rect 1453 9859 1455 9863
rect 1447 9858 1455 9859
rect 1383 9856 1455 9858
rect 1383 9852 1385 9856
rect 1389 9852 1392 9856
rect 1396 9852 1397 9856
rect 1401 9852 1402 9856
rect 1406 9852 1407 9856
rect 1411 9852 1412 9856
rect 1416 9852 1417 9856
rect 1421 9852 1422 9856
rect 1426 9852 1427 9856
rect 1431 9852 1432 9856
rect 1436 9852 1437 9856
rect 1441 9852 1442 9856
rect 1446 9852 1449 9856
rect 1453 9852 1455 9856
rect 1383 9850 1455 9852
rect 1531 9978 1627 9979
rect 1531 9974 1532 9978
rect 1536 9974 1537 9978
rect 1541 9974 1542 9978
rect 1546 9974 1547 9978
rect 1551 9974 1552 9978
rect 1556 9974 1557 9978
rect 1561 9974 1562 9978
rect 1566 9974 1567 9978
rect 1571 9974 1572 9978
rect 1576 9974 1577 9978
rect 1581 9974 1582 9978
rect 1586 9974 1587 9978
rect 1591 9974 1592 9978
rect 1596 9974 1597 9978
rect 1601 9974 1602 9978
rect 1606 9974 1607 9978
rect 1611 9974 1612 9978
rect 1616 9974 1617 9978
rect 1621 9974 1622 9978
rect 1626 9974 1627 9978
rect 1531 9973 1627 9974
rect 1531 9969 1532 9973
rect 1536 9969 1537 9973
rect 1531 9968 1537 9969
rect 1531 9964 1532 9968
rect 1536 9964 1537 9968
rect 1621 9969 1622 9973
rect 1626 9969 1627 9973
rect 1621 9968 1627 9969
rect 1531 9963 1537 9964
rect 1531 9959 1532 9963
rect 1536 9959 1537 9963
rect 1531 9958 1537 9959
rect 1531 9954 1532 9958
rect 1536 9954 1537 9958
rect 1531 9953 1537 9954
rect 1531 9949 1532 9953
rect 1536 9949 1537 9953
rect 1531 9948 1537 9949
rect 1531 9944 1532 9948
rect 1536 9944 1537 9948
rect 1531 9943 1537 9944
rect 1531 9939 1532 9943
rect 1536 9939 1537 9943
rect 1531 9938 1537 9939
rect 1531 9934 1532 9938
rect 1536 9934 1537 9938
rect 1531 9933 1537 9934
rect 1531 9929 1532 9933
rect 1536 9929 1537 9933
rect 1531 9928 1537 9929
rect 1531 9924 1532 9928
rect 1536 9924 1537 9928
rect 1531 9923 1537 9924
rect 1531 9919 1532 9923
rect 1536 9919 1537 9923
rect 1531 9918 1537 9919
rect 1531 9914 1532 9918
rect 1536 9914 1537 9918
rect 1531 9913 1537 9914
rect 1531 9909 1532 9913
rect 1536 9909 1537 9913
rect 1531 9908 1537 9909
rect 1531 9904 1532 9908
rect 1536 9904 1537 9908
rect 1531 9903 1537 9904
rect 1531 9899 1532 9903
rect 1536 9899 1537 9903
rect 1531 9898 1537 9899
rect 1531 9894 1532 9898
rect 1536 9894 1537 9898
rect 1531 9893 1537 9894
rect 1531 9889 1532 9893
rect 1536 9889 1537 9893
rect 1531 9888 1537 9889
rect 1531 9884 1532 9888
rect 1536 9884 1537 9888
rect 1531 9883 1537 9884
rect 1531 9879 1532 9883
rect 1536 9879 1537 9883
rect 1531 9878 1537 9879
rect 1531 9874 1532 9878
rect 1536 9874 1537 9878
rect 1531 9873 1537 9874
rect 1531 9869 1532 9873
rect 1536 9869 1537 9873
rect 1531 9868 1537 9869
rect 1531 9864 1532 9868
rect 1536 9864 1537 9868
rect 1531 9863 1537 9864
rect 1531 9859 1532 9863
rect 1536 9859 1537 9863
rect 1531 9858 1537 9859
rect 1531 9854 1532 9858
rect 1536 9854 1537 9858
rect 1531 9853 1537 9854
rect 1531 9849 1532 9853
rect 1536 9849 1537 9853
rect 1621 9964 1622 9968
rect 1626 9964 1627 9968
rect 1621 9963 1627 9964
rect 1621 9959 1622 9963
rect 1626 9959 1627 9963
rect 1621 9958 1627 9959
rect 1621 9954 1622 9958
rect 1626 9954 1627 9958
rect 1621 9953 1627 9954
rect 1621 9949 1622 9953
rect 1626 9949 1627 9953
rect 1621 9948 1627 9949
rect 1621 9944 1622 9948
rect 1626 9944 1627 9948
rect 1621 9943 1627 9944
rect 1621 9939 1622 9943
rect 1626 9939 1627 9943
rect 1621 9938 1627 9939
rect 1621 9934 1622 9938
rect 1626 9934 1627 9938
rect 1621 9933 1627 9934
rect 1621 9929 1622 9933
rect 1626 9929 1627 9933
rect 1621 9928 1627 9929
rect 1621 9924 1622 9928
rect 1626 9924 1627 9928
rect 1621 9923 1627 9924
rect 1621 9919 1622 9923
rect 1626 9919 1627 9923
rect 1621 9918 1627 9919
rect 1621 9914 1622 9918
rect 1626 9914 1627 9918
rect 1621 9913 1627 9914
rect 1621 9909 1622 9913
rect 1626 9909 1627 9913
rect 1621 9908 1627 9909
rect 1621 9904 1622 9908
rect 1626 9904 1627 9908
rect 1621 9903 1627 9904
rect 1621 9899 1622 9903
rect 1626 9899 1627 9903
rect 1621 9898 1627 9899
rect 1621 9894 1622 9898
rect 1626 9894 1627 9898
rect 1621 9893 1627 9894
rect 1621 9889 1622 9893
rect 1626 9889 1627 9893
rect 1621 9888 1627 9889
rect 1621 9884 1622 9888
rect 1626 9884 1627 9888
rect 1621 9883 1627 9884
rect 1621 9879 1622 9883
rect 1626 9879 1627 9883
rect 1621 9878 1627 9879
rect 1621 9874 1622 9878
rect 1626 9874 1627 9878
rect 1621 9873 1627 9874
rect 1621 9869 1622 9873
rect 1626 9869 1627 9873
rect 1621 9868 1627 9869
rect 1621 9864 1622 9868
rect 1626 9864 1627 9868
rect 1621 9863 1627 9864
rect 1621 9859 1622 9863
rect 1626 9859 1627 9863
rect 1621 9858 1627 9859
rect 1621 9854 1622 9858
rect 1626 9854 1627 9858
rect 1621 9853 1627 9854
rect 1531 9848 1537 9849
rect 1531 9844 1532 9848
rect 1536 9844 1537 9848
rect 1621 9849 1622 9853
rect 1626 9849 1627 9853
rect 1621 9848 1627 9849
rect 1621 9844 1622 9848
rect 1626 9844 1627 9848
rect 1531 9843 1627 9844
rect 1531 9839 1532 9843
rect 1536 9839 1537 9843
rect 1541 9839 1542 9843
rect 1546 9839 1547 9843
rect 1551 9839 1552 9843
rect 1556 9839 1557 9843
rect 1561 9839 1562 9843
rect 1566 9839 1567 9843
rect 1571 9839 1572 9843
rect 1576 9839 1577 9843
rect 1581 9839 1582 9843
rect 1586 9839 1587 9843
rect 1591 9839 1592 9843
rect 1596 9839 1597 9843
rect 1601 9839 1602 9843
rect 1606 9839 1607 9843
rect 1611 9839 1612 9843
rect 1616 9839 1617 9843
rect 1621 9839 1622 9843
rect 1626 9839 1627 9843
rect 1531 9838 1627 9839
rect 1692 9965 1764 9967
rect 1692 9961 1694 9965
rect 1698 9961 1701 9965
rect 1705 9961 1706 9965
rect 1710 9961 1711 9965
rect 1715 9961 1716 9965
rect 1720 9961 1721 9965
rect 1725 9961 1726 9965
rect 1730 9961 1731 9965
rect 1735 9961 1736 9965
rect 1740 9961 1741 9965
rect 1745 9961 1746 9965
rect 1750 9961 1751 9965
rect 1755 9961 1758 9965
rect 1762 9961 1764 9965
rect 1692 9959 1764 9961
rect 1692 9958 1700 9959
rect 1692 9954 1694 9958
rect 1698 9954 1700 9958
rect 1692 9953 1700 9954
rect 1756 9958 1764 9959
rect 1756 9954 1758 9958
rect 1762 9954 1764 9958
rect 1756 9953 1764 9954
rect 1692 9949 1694 9953
rect 1698 9949 1700 9953
rect 1692 9948 1700 9949
rect 1692 9944 1694 9948
rect 1698 9944 1700 9948
rect 1692 9943 1700 9944
rect 1692 9939 1694 9943
rect 1698 9939 1700 9943
rect 1692 9938 1700 9939
rect 1692 9934 1694 9938
rect 1698 9934 1700 9938
rect 1692 9933 1700 9934
rect 1692 9929 1694 9933
rect 1698 9929 1700 9933
rect 1692 9928 1700 9929
rect 1692 9924 1694 9928
rect 1698 9924 1700 9928
rect 1692 9923 1700 9924
rect 1692 9919 1694 9923
rect 1698 9919 1700 9923
rect 1692 9918 1700 9919
rect 1692 9914 1694 9918
rect 1698 9914 1700 9918
rect 1692 9913 1700 9914
rect 1692 9909 1694 9913
rect 1698 9909 1700 9913
rect 1692 9908 1700 9909
rect 1692 9904 1694 9908
rect 1698 9904 1700 9908
rect 1692 9903 1700 9904
rect 1692 9899 1694 9903
rect 1698 9899 1700 9903
rect 1692 9898 1700 9899
rect 1692 9894 1694 9898
rect 1698 9894 1700 9898
rect 1692 9893 1700 9894
rect 1692 9889 1694 9893
rect 1698 9889 1700 9893
rect 1692 9888 1700 9889
rect 1692 9884 1694 9888
rect 1698 9884 1700 9888
rect 1692 9883 1700 9884
rect 1692 9879 1694 9883
rect 1698 9879 1700 9883
rect 1692 9878 1700 9879
rect 1692 9874 1694 9878
rect 1698 9874 1700 9878
rect 1692 9873 1700 9874
rect 1692 9869 1694 9873
rect 1698 9869 1700 9873
rect 1692 9868 1700 9869
rect 1692 9864 1694 9868
rect 1698 9864 1700 9868
rect 1756 9949 1758 9953
rect 1762 9949 1764 9953
rect 1756 9948 1764 9949
rect 1756 9944 1758 9948
rect 1762 9944 1764 9948
rect 1756 9943 1764 9944
rect 1756 9939 1758 9943
rect 1762 9939 1764 9943
rect 1756 9938 1764 9939
rect 1756 9934 1758 9938
rect 1762 9934 1764 9938
rect 1756 9933 1764 9934
rect 1756 9929 1758 9933
rect 1762 9929 1764 9933
rect 1756 9928 1764 9929
rect 1756 9924 1758 9928
rect 1762 9924 1764 9928
rect 1756 9923 1764 9924
rect 1756 9919 1758 9923
rect 1762 9919 1764 9923
rect 1756 9918 1764 9919
rect 1756 9914 1758 9918
rect 1762 9914 1764 9918
rect 1756 9913 1764 9914
rect 1756 9909 1758 9913
rect 1762 9909 1764 9913
rect 1756 9908 1764 9909
rect 1756 9904 1758 9908
rect 1762 9904 1764 9908
rect 1756 9903 1764 9904
rect 1756 9899 1758 9903
rect 1762 9899 1764 9903
rect 1756 9898 1764 9899
rect 1756 9894 1758 9898
rect 1762 9894 1764 9898
rect 1756 9893 1764 9894
rect 1756 9889 1758 9893
rect 1762 9889 1764 9893
rect 1756 9888 1764 9889
rect 1756 9884 1758 9888
rect 1762 9884 1764 9888
rect 1756 9883 1764 9884
rect 1756 9879 1758 9883
rect 1762 9879 1764 9883
rect 1756 9878 1764 9879
rect 1756 9874 1758 9878
rect 1762 9874 1764 9878
rect 1756 9873 1764 9874
rect 1756 9869 1758 9873
rect 1762 9869 1764 9873
rect 1756 9868 1764 9869
rect 1756 9864 1758 9868
rect 1762 9864 1764 9868
rect 1692 9863 1700 9864
rect 1692 9859 1694 9863
rect 1698 9859 1700 9863
rect 1692 9858 1700 9859
rect 1756 9863 1764 9864
rect 1756 9859 1758 9863
rect 1762 9859 1764 9863
rect 1756 9858 1764 9859
rect 1692 9856 1764 9858
rect 1692 9852 1694 9856
rect 1698 9852 1701 9856
rect 1705 9852 1706 9856
rect 1710 9852 1711 9856
rect 1715 9852 1716 9856
rect 1720 9852 1721 9856
rect 1725 9852 1726 9856
rect 1730 9852 1731 9856
rect 1735 9852 1736 9856
rect 1740 9852 1741 9856
rect 1745 9852 1746 9856
rect 1750 9852 1751 9856
rect 1755 9852 1758 9856
rect 1762 9852 1764 9856
rect 1692 9850 1764 9852
rect 1840 9978 1936 9979
rect 1840 9974 1841 9978
rect 1845 9974 1846 9978
rect 1850 9974 1851 9978
rect 1855 9974 1856 9978
rect 1860 9974 1861 9978
rect 1865 9974 1866 9978
rect 1870 9974 1871 9978
rect 1875 9974 1876 9978
rect 1880 9974 1881 9978
rect 1885 9974 1886 9978
rect 1890 9974 1891 9978
rect 1895 9974 1896 9978
rect 1900 9974 1901 9978
rect 1905 9974 1906 9978
rect 1910 9974 1911 9978
rect 1915 9974 1916 9978
rect 1920 9974 1921 9978
rect 1925 9974 1926 9978
rect 1930 9974 1931 9978
rect 1935 9974 1936 9978
rect 1840 9973 1936 9974
rect 1840 9969 1841 9973
rect 1845 9969 1846 9973
rect 1840 9968 1846 9969
rect 1840 9964 1841 9968
rect 1845 9964 1846 9968
rect 1930 9969 1931 9973
rect 1935 9969 1936 9973
rect 1930 9968 1936 9969
rect 1840 9963 1846 9964
rect 1840 9959 1841 9963
rect 1845 9959 1846 9963
rect 1840 9958 1846 9959
rect 1840 9954 1841 9958
rect 1845 9954 1846 9958
rect 1840 9953 1846 9954
rect 1840 9949 1841 9953
rect 1845 9949 1846 9953
rect 1840 9948 1846 9949
rect 1840 9944 1841 9948
rect 1845 9944 1846 9948
rect 1840 9943 1846 9944
rect 1840 9939 1841 9943
rect 1845 9939 1846 9943
rect 1840 9938 1846 9939
rect 1840 9934 1841 9938
rect 1845 9934 1846 9938
rect 1840 9933 1846 9934
rect 1840 9929 1841 9933
rect 1845 9929 1846 9933
rect 1840 9928 1846 9929
rect 1840 9924 1841 9928
rect 1845 9924 1846 9928
rect 1840 9923 1846 9924
rect 1840 9919 1841 9923
rect 1845 9919 1846 9923
rect 1840 9918 1846 9919
rect 1840 9914 1841 9918
rect 1845 9914 1846 9918
rect 1840 9913 1846 9914
rect 1840 9909 1841 9913
rect 1845 9909 1846 9913
rect 1840 9908 1846 9909
rect 1840 9904 1841 9908
rect 1845 9904 1846 9908
rect 1840 9903 1846 9904
rect 1840 9899 1841 9903
rect 1845 9899 1846 9903
rect 1840 9898 1846 9899
rect 1840 9894 1841 9898
rect 1845 9894 1846 9898
rect 1840 9893 1846 9894
rect 1840 9889 1841 9893
rect 1845 9889 1846 9893
rect 1840 9888 1846 9889
rect 1840 9884 1841 9888
rect 1845 9884 1846 9888
rect 1840 9883 1846 9884
rect 1840 9879 1841 9883
rect 1845 9879 1846 9883
rect 1840 9878 1846 9879
rect 1840 9874 1841 9878
rect 1845 9874 1846 9878
rect 1840 9873 1846 9874
rect 1840 9869 1841 9873
rect 1845 9869 1846 9873
rect 1840 9868 1846 9869
rect 1840 9864 1841 9868
rect 1845 9864 1846 9868
rect 1840 9863 1846 9864
rect 1840 9859 1841 9863
rect 1845 9859 1846 9863
rect 1840 9858 1846 9859
rect 1840 9854 1841 9858
rect 1845 9854 1846 9858
rect 1840 9853 1846 9854
rect 1840 9849 1841 9853
rect 1845 9849 1846 9853
rect 1930 9964 1931 9968
rect 1935 9964 1936 9968
rect 1930 9963 1936 9964
rect 1930 9959 1931 9963
rect 1935 9959 1936 9963
rect 1930 9958 1936 9959
rect 1930 9954 1931 9958
rect 1935 9954 1936 9958
rect 1930 9953 1936 9954
rect 1930 9949 1931 9953
rect 1935 9949 1936 9953
rect 1930 9948 1936 9949
rect 1930 9944 1931 9948
rect 1935 9944 1936 9948
rect 1930 9943 1936 9944
rect 1930 9939 1931 9943
rect 1935 9939 1936 9943
rect 1930 9938 1936 9939
rect 1930 9934 1931 9938
rect 1935 9934 1936 9938
rect 1930 9933 1936 9934
rect 1930 9929 1931 9933
rect 1935 9929 1936 9933
rect 1930 9928 1936 9929
rect 1930 9924 1931 9928
rect 1935 9924 1936 9928
rect 1930 9923 1936 9924
rect 1930 9919 1931 9923
rect 1935 9919 1936 9923
rect 1930 9918 1936 9919
rect 1930 9914 1931 9918
rect 1935 9914 1936 9918
rect 1930 9913 1936 9914
rect 1930 9909 1931 9913
rect 1935 9909 1936 9913
rect 1930 9908 1936 9909
rect 1930 9904 1931 9908
rect 1935 9904 1936 9908
rect 1930 9903 1936 9904
rect 1930 9899 1931 9903
rect 1935 9899 1936 9903
rect 1930 9898 1936 9899
rect 1930 9894 1931 9898
rect 1935 9894 1936 9898
rect 1930 9893 1936 9894
rect 1930 9889 1931 9893
rect 1935 9889 1936 9893
rect 1930 9888 1936 9889
rect 1930 9884 1931 9888
rect 1935 9884 1936 9888
rect 1930 9883 1936 9884
rect 1930 9879 1931 9883
rect 1935 9879 1936 9883
rect 1930 9878 1936 9879
rect 1930 9874 1931 9878
rect 1935 9874 1936 9878
rect 1930 9873 1936 9874
rect 1930 9869 1931 9873
rect 1935 9869 1936 9873
rect 1930 9868 1936 9869
rect 1930 9864 1931 9868
rect 1935 9864 1936 9868
rect 1930 9863 1936 9864
rect 1930 9859 1931 9863
rect 1935 9859 1936 9863
rect 1930 9858 1936 9859
rect 1930 9854 1931 9858
rect 1935 9854 1936 9858
rect 1930 9853 1936 9854
rect 1840 9848 1846 9849
rect 1840 9844 1841 9848
rect 1845 9844 1846 9848
rect 1930 9849 1931 9853
rect 1935 9849 1936 9853
rect 1930 9848 1936 9849
rect 1930 9844 1931 9848
rect 1935 9844 1936 9848
rect 1840 9843 1936 9844
rect 1840 9839 1841 9843
rect 1845 9839 1846 9843
rect 1850 9839 1851 9843
rect 1855 9839 1856 9843
rect 1860 9839 1861 9843
rect 1865 9839 1866 9843
rect 1870 9839 1871 9843
rect 1875 9839 1876 9843
rect 1880 9839 1881 9843
rect 1885 9839 1886 9843
rect 1890 9839 1891 9843
rect 1895 9839 1896 9843
rect 1900 9839 1901 9843
rect 1905 9839 1906 9843
rect 1910 9839 1911 9843
rect 1915 9839 1916 9843
rect 1920 9839 1921 9843
rect 1925 9839 1926 9843
rect 1930 9839 1931 9843
rect 1935 9839 1936 9843
rect 1840 9838 1936 9839
rect 2001 9965 2073 9967
rect 2001 9961 2003 9965
rect 2007 9961 2010 9965
rect 2014 9961 2015 9965
rect 2019 9961 2020 9965
rect 2024 9961 2025 9965
rect 2029 9961 2030 9965
rect 2034 9961 2035 9965
rect 2039 9961 2040 9965
rect 2044 9961 2045 9965
rect 2049 9961 2050 9965
rect 2054 9961 2055 9965
rect 2059 9961 2060 9965
rect 2064 9961 2067 9965
rect 2071 9961 2073 9965
rect 2001 9959 2073 9961
rect 2001 9958 2009 9959
rect 2001 9954 2003 9958
rect 2007 9954 2009 9958
rect 2001 9953 2009 9954
rect 2065 9958 2073 9959
rect 2065 9954 2067 9958
rect 2071 9954 2073 9958
rect 2065 9953 2073 9954
rect 2001 9949 2003 9953
rect 2007 9949 2009 9953
rect 2001 9948 2009 9949
rect 2001 9944 2003 9948
rect 2007 9944 2009 9948
rect 2001 9943 2009 9944
rect 2001 9939 2003 9943
rect 2007 9939 2009 9943
rect 2001 9938 2009 9939
rect 2001 9934 2003 9938
rect 2007 9934 2009 9938
rect 2001 9933 2009 9934
rect 2001 9929 2003 9933
rect 2007 9929 2009 9933
rect 2001 9928 2009 9929
rect 2001 9924 2003 9928
rect 2007 9924 2009 9928
rect 2001 9923 2009 9924
rect 2001 9919 2003 9923
rect 2007 9919 2009 9923
rect 2001 9918 2009 9919
rect 2001 9914 2003 9918
rect 2007 9914 2009 9918
rect 2001 9913 2009 9914
rect 2001 9909 2003 9913
rect 2007 9909 2009 9913
rect 2001 9908 2009 9909
rect 2001 9904 2003 9908
rect 2007 9904 2009 9908
rect 2001 9903 2009 9904
rect 2001 9899 2003 9903
rect 2007 9899 2009 9903
rect 2001 9898 2009 9899
rect 2001 9894 2003 9898
rect 2007 9894 2009 9898
rect 2001 9893 2009 9894
rect 2001 9889 2003 9893
rect 2007 9889 2009 9893
rect 2001 9888 2009 9889
rect 2001 9884 2003 9888
rect 2007 9884 2009 9888
rect 2001 9883 2009 9884
rect 2001 9879 2003 9883
rect 2007 9879 2009 9883
rect 2001 9878 2009 9879
rect 2001 9874 2003 9878
rect 2007 9874 2009 9878
rect 2001 9873 2009 9874
rect 2001 9869 2003 9873
rect 2007 9869 2009 9873
rect 2001 9868 2009 9869
rect 2001 9864 2003 9868
rect 2007 9864 2009 9868
rect 2065 9949 2067 9953
rect 2071 9949 2073 9953
rect 2065 9948 2073 9949
rect 2065 9944 2067 9948
rect 2071 9944 2073 9948
rect 2065 9943 2073 9944
rect 2065 9939 2067 9943
rect 2071 9939 2073 9943
rect 2065 9938 2073 9939
rect 2065 9934 2067 9938
rect 2071 9934 2073 9938
rect 2065 9933 2073 9934
rect 2065 9929 2067 9933
rect 2071 9929 2073 9933
rect 2065 9928 2073 9929
rect 2065 9924 2067 9928
rect 2071 9924 2073 9928
rect 2065 9923 2073 9924
rect 2065 9919 2067 9923
rect 2071 9919 2073 9923
rect 2065 9918 2073 9919
rect 2065 9914 2067 9918
rect 2071 9914 2073 9918
rect 2065 9913 2073 9914
rect 2065 9909 2067 9913
rect 2071 9909 2073 9913
rect 2065 9908 2073 9909
rect 2065 9904 2067 9908
rect 2071 9904 2073 9908
rect 2065 9903 2073 9904
rect 2065 9899 2067 9903
rect 2071 9899 2073 9903
rect 2065 9898 2073 9899
rect 2065 9894 2067 9898
rect 2071 9894 2073 9898
rect 2065 9893 2073 9894
rect 2065 9889 2067 9893
rect 2071 9889 2073 9893
rect 2065 9888 2073 9889
rect 2065 9884 2067 9888
rect 2071 9884 2073 9888
rect 2065 9883 2073 9884
rect 2065 9879 2067 9883
rect 2071 9879 2073 9883
rect 2065 9878 2073 9879
rect 2065 9874 2067 9878
rect 2071 9874 2073 9878
rect 2065 9873 2073 9874
rect 2065 9869 2067 9873
rect 2071 9869 2073 9873
rect 2065 9868 2073 9869
rect 2065 9864 2067 9868
rect 2071 9864 2073 9868
rect 2001 9863 2009 9864
rect 2001 9859 2003 9863
rect 2007 9859 2009 9863
rect 2001 9858 2009 9859
rect 2065 9863 2073 9864
rect 2065 9859 2067 9863
rect 2071 9859 2073 9863
rect 2065 9858 2073 9859
rect 2001 9856 2073 9858
rect 2001 9852 2003 9856
rect 2007 9852 2010 9856
rect 2014 9852 2015 9856
rect 2019 9852 2020 9856
rect 2024 9852 2025 9856
rect 2029 9852 2030 9856
rect 2034 9852 2035 9856
rect 2039 9852 2040 9856
rect 2044 9852 2045 9856
rect 2049 9852 2050 9856
rect 2054 9852 2055 9856
rect 2059 9852 2060 9856
rect 2064 9852 2067 9856
rect 2071 9852 2073 9856
rect 2001 9850 2073 9852
rect 2149 9978 2245 9979
rect 2149 9974 2150 9978
rect 2154 9974 2155 9978
rect 2159 9974 2160 9978
rect 2164 9974 2165 9978
rect 2169 9974 2170 9978
rect 2174 9974 2175 9978
rect 2179 9974 2180 9978
rect 2184 9974 2185 9978
rect 2189 9974 2190 9978
rect 2194 9974 2195 9978
rect 2199 9974 2200 9978
rect 2204 9974 2205 9978
rect 2209 9974 2210 9978
rect 2214 9974 2215 9978
rect 2219 9974 2220 9978
rect 2224 9974 2225 9978
rect 2229 9974 2230 9978
rect 2234 9974 2235 9978
rect 2239 9974 2240 9978
rect 2244 9974 2245 9978
rect 2149 9973 2245 9974
rect 2149 9969 2150 9973
rect 2154 9969 2155 9973
rect 2149 9968 2155 9969
rect 2149 9964 2150 9968
rect 2154 9964 2155 9968
rect 2239 9969 2240 9973
rect 2244 9969 2245 9973
rect 2239 9968 2245 9969
rect 2149 9963 2155 9964
rect 2149 9959 2150 9963
rect 2154 9959 2155 9963
rect 2149 9958 2155 9959
rect 2149 9954 2150 9958
rect 2154 9954 2155 9958
rect 2149 9953 2155 9954
rect 2149 9949 2150 9953
rect 2154 9949 2155 9953
rect 2149 9948 2155 9949
rect 2149 9944 2150 9948
rect 2154 9944 2155 9948
rect 2149 9943 2155 9944
rect 2149 9939 2150 9943
rect 2154 9939 2155 9943
rect 2149 9938 2155 9939
rect 2149 9934 2150 9938
rect 2154 9934 2155 9938
rect 2149 9933 2155 9934
rect 2149 9929 2150 9933
rect 2154 9929 2155 9933
rect 2149 9928 2155 9929
rect 2149 9924 2150 9928
rect 2154 9924 2155 9928
rect 2149 9923 2155 9924
rect 2149 9919 2150 9923
rect 2154 9919 2155 9923
rect 2149 9918 2155 9919
rect 2149 9914 2150 9918
rect 2154 9914 2155 9918
rect 2149 9913 2155 9914
rect 2149 9909 2150 9913
rect 2154 9909 2155 9913
rect 2149 9908 2155 9909
rect 2149 9904 2150 9908
rect 2154 9904 2155 9908
rect 2149 9903 2155 9904
rect 2149 9899 2150 9903
rect 2154 9899 2155 9903
rect 2149 9898 2155 9899
rect 2149 9894 2150 9898
rect 2154 9894 2155 9898
rect 2149 9893 2155 9894
rect 2149 9889 2150 9893
rect 2154 9889 2155 9893
rect 2149 9888 2155 9889
rect 2149 9884 2150 9888
rect 2154 9884 2155 9888
rect 2149 9883 2155 9884
rect 2149 9879 2150 9883
rect 2154 9879 2155 9883
rect 2149 9878 2155 9879
rect 2149 9874 2150 9878
rect 2154 9874 2155 9878
rect 2149 9873 2155 9874
rect 2149 9869 2150 9873
rect 2154 9869 2155 9873
rect 2149 9868 2155 9869
rect 2149 9864 2150 9868
rect 2154 9864 2155 9868
rect 2149 9863 2155 9864
rect 2149 9859 2150 9863
rect 2154 9859 2155 9863
rect 2149 9858 2155 9859
rect 2149 9854 2150 9858
rect 2154 9854 2155 9858
rect 2149 9853 2155 9854
rect 2149 9849 2150 9853
rect 2154 9849 2155 9853
rect 2239 9964 2240 9968
rect 2244 9964 2245 9968
rect 2239 9963 2245 9964
rect 2239 9959 2240 9963
rect 2244 9959 2245 9963
rect 2239 9958 2245 9959
rect 2239 9954 2240 9958
rect 2244 9954 2245 9958
rect 2239 9953 2245 9954
rect 2239 9949 2240 9953
rect 2244 9949 2245 9953
rect 2239 9948 2245 9949
rect 2239 9944 2240 9948
rect 2244 9944 2245 9948
rect 2239 9943 2245 9944
rect 2239 9939 2240 9943
rect 2244 9939 2245 9943
rect 2239 9938 2245 9939
rect 2239 9934 2240 9938
rect 2244 9934 2245 9938
rect 2239 9933 2245 9934
rect 2239 9929 2240 9933
rect 2244 9929 2245 9933
rect 2239 9928 2245 9929
rect 2239 9924 2240 9928
rect 2244 9924 2245 9928
rect 2239 9923 2245 9924
rect 2239 9919 2240 9923
rect 2244 9919 2245 9923
rect 2239 9918 2245 9919
rect 2239 9914 2240 9918
rect 2244 9914 2245 9918
rect 2239 9913 2245 9914
rect 2239 9909 2240 9913
rect 2244 9909 2245 9913
rect 2239 9908 2245 9909
rect 2239 9904 2240 9908
rect 2244 9904 2245 9908
rect 2239 9903 2245 9904
rect 2239 9899 2240 9903
rect 2244 9899 2245 9903
rect 2239 9898 2245 9899
rect 2239 9894 2240 9898
rect 2244 9894 2245 9898
rect 2239 9893 2245 9894
rect 2239 9889 2240 9893
rect 2244 9889 2245 9893
rect 2239 9888 2245 9889
rect 2239 9884 2240 9888
rect 2244 9884 2245 9888
rect 2239 9883 2245 9884
rect 2239 9879 2240 9883
rect 2244 9879 2245 9883
rect 2239 9878 2245 9879
rect 2239 9874 2240 9878
rect 2244 9874 2245 9878
rect 2239 9873 2245 9874
rect 2239 9869 2240 9873
rect 2244 9869 2245 9873
rect 2239 9868 2245 9869
rect 2239 9864 2240 9868
rect 2244 9864 2245 9868
rect 2239 9863 2245 9864
rect 2239 9859 2240 9863
rect 2244 9859 2245 9863
rect 2239 9858 2245 9859
rect 2239 9854 2240 9858
rect 2244 9854 2245 9858
rect 2239 9853 2245 9854
rect 2149 9848 2155 9849
rect 2149 9844 2150 9848
rect 2154 9844 2155 9848
rect 2239 9849 2240 9853
rect 2244 9849 2245 9853
rect 2239 9848 2245 9849
rect 2239 9844 2240 9848
rect 2244 9844 2245 9848
rect 2149 9843 2245 9844
rect 2149 9839 2150 9843
rect 2154 9839 2155 9843
rect 2159 9839 2160 9843
rect 2164 9839 2165 9843
rect 2169 9839 2170 9843
rect 2174 9839 2175 9843
rect 2179 9839 2180 9843
rect 2184 9839 2185 9843
rect 2189 9839 2190 9843
rect 2194 9839 2195 9843
rect 2199 9839 2200 9843
rect 2204 9839 2205 9843
rect 2209 9839 2210 9843
rect 2214 9839 2215 9843
rect 2219 9839 2220 9843
rect 2224 9839 2225 9843
rect 2229 9839 2230 9843
rect 2234 9839 2235 9843
rect 2239 9839 2240 9843
rect 2244 9839 2245 9843
rect 2149 9838 2245 9839
rect 2310 9965 2382 9967
rect 2310 9961 2312 9965
rect 2316 9961 2319 9965
rect 2323 9961 2324 9965
rect 2328 9961 2329 9965
rect 2333 9961 2334 9965
rect 2338 9961 2339 9965
rect 2343 9961 2344 9965
rect 2348 9961 2349 9965
rect 2353 9961 2354 9965
rect 2358 9961 2359 9965
rect 2363 9961 2364 9965
rect 2368 9961 2369 9965
rect 2373 9961 2376 9965
rect 2380 9961 2382 9965
rect 2310 9959 2382 9961
rect 2310 9958 2318 9959
rect 2310 9954 2312 9958
rect 2316 9954 2318 9958
rect 2310 9953 2318 9954
rect 2374 9958 2382 9959
rect 2374 9954 2376 9958
rect 2380 9954 2382 9958
rect 2374 9953 2382 9954
rect 2310 9949 2312 9953
rect 2316 9949 2318 9953
rect 2310 9948 2318 9949
rect 2310 9944 2312 9948
rect 2316 9944 2318 9948
rect 2310 9943 2318 9944
rect 2310 9939 2312 9943
rect 2316 9939 2318 9943
rect 2310 9938 2318 9939
rect 2310 9934 2312 9938
rect 2316 9934 2318 9938
rect 2310 9933 2318 9934
rect 2310 9929 2312 9933
rect 2316 9929 2318 9933
rect 2310 9928 2318 9929
rect 2310 9924 2312 9928
rect 2316 9924 2318 9928
rect 2310 9923 2318 9924
rect 2310 9919 2312 9923
rect 2316 9919 2318 9923
rect 2310 9918 2318 9919
rect 2310 9914 2312 9918
rect 2316 9914 2318 9918
rect 2310 9913 2318 9914
rect 2310 9909 2312 9913
rect 2316 9909 2318 9913
rect 2310 9908 2318 9909
rect 2310 9904 2312 9908
rect 2316 9904 2318 9908
rect 2310 9903 2318 9904
rect 2310 9899 2312 9903
rect 2316 9899 2318 9903
rect 2310 9898 2318 9899
rect 2310 9894 2312 9898
rect 2316 9894 2318 9898
rect 2310 9893 2318 9894
rect 2310 9889 2312 9893
rect 2316 9889 2318 9893
rect 2310 9888 2318 9889
rect 2310 9884 2312 9888
rect 2316 9884 2318 9888
rect 2310 9883 2318 9884
rect 2310 9879 2312 9883
rect 2316 9879 2318 9883
rect 2310 9878 2318 9879
rect 2310 9874 2312 9878
rect 2316 9874 2318 9878
rect 2310 9873 2318 9874
rect 2310 9869 2312 9873
rect 2316 9869 2318 9873
rect 2310 9868 2318 9869
rect 2310 9864 2312 9868
rect 2316 9864 2318 9868
rect 2374 9949 2376 9953
rect 2380 9949 2382 9953
rect 2374 9948 2382 9949
rect 2374 9944 2376 9948
rect 2380 9944 2382 9948
rect 2374 9943 2382 9944
rect 2374 9939 2376 9943
rect 2380 9939 2382 9943
rect 2374 9938 2382 9939
rect 2374 9934 2376 9938
rect 2380 9934 2382 9938
rect 2374 9933 2382 9934
rect 2374 9929 2376 9933
rect 2380 9929 2382 9933
rect 2374 9928 2382 9929
rect 2374 9924 2376 9928
rect 2380 9924 2382 9928
rect 2374 9923 2382 9924
rect 2374 9919 2376 9923
rect 2380 9919 2382 9923
rect 2374 9918 2382 9919
rect 2374 9914 2376 9918
rect 2380 9914 2382 9918
rect 2374 9913 2382 9914
rect 2374 9909 2376 9913
rect 2380 9909 2382 9913
rect 2374 9908 2382 9909
rect 2374 9904 2376 9908
rect 2380 9904 2382 9908
rect 2374 9903 2382 9904
rect 2374 9899 2376 9903
rect 2380 9899 2382 9903
rect 2374 9898 2382 9899
rect 2374 9894 2376 9898
rect 2380 9894 2382 9898
rect 2374 9893 2382 9894
rect 2374 9889 2376 9893
rect 2380 9889 2382 9893
rect 2374 9888 2382 9889
rect 2374 9884 2376 9888
rect 2380 9884 2382 9888
rect 2374 9883 2382 9884
rect 2374 9879 2376 9883
rect 2380 9879 2382 9883
rect 2374 9878 2382 9879
rect 2374 9874 2376 9878
rect 2380 9874 2382 9878
rect 2374 9873 2382 9874
rect 2374 9869 2376 9873
rect 2380 9869 2382 9873
rect 2374 9868 2382 9869
rect 2374 9864 2376 9868
rect 2380 9864 2382 9868
rect 2310 9863 2318 9864
rect 2310 9859 2312 9863
rect 2316 9859 2318 9863
rect 2310 9858 2318 9859
rect 2374 9863 2382 9864
rect 2374 9859 2376 9863
rect 2380 9859 2382 9863
rect 2374 9858 2382 9859
rect 2310 9856 2382 9858
rect 2310 9852 2312 9856
rect 2316 9852 2319 9856
rect 2323 9852 2324 9856
rect 2328 9852 2329 9856
rect 2333 9852 2334 9856
rect 2338 9852 2339 9856
rect 2343 9852 2344 9856
rect 2348 9852 2349 9856
rect 2353 9852 2354 9856
rect 2358 9852 2359 9856
rect 2363 9852 2364 9856
rect 2368 9852 2369 9856
rect 2373 9852 2376 9856
rect 2380 9852 2382 9856
rect 2310 9850 2382 9852
rect 2458 9978 2554 9979
rect 2458 9974 2459 9978
rect 2463 9974 2464 9978
rect 2468 9974 2469 9978
rect 2473 9974 2474 9978
rect 2478 9974 2479 9978
rect 2483 9974 2484 9978
rect 2488 9974 2489 9978
rect 2493 9974 2494 9978
rect 2498 9974 2499 9978
rect 2503 9974 2504 9978
rect 2508 9974 2509 9978
rect 2513 9974 2514 9978
rect 2518 9974 2519 9978
rect 2523 9974 2524 9978
rect 2528 9974 2529 9978
rect 2533 9974 2534 9978
rect 2538 9974 2539 9978
rect 2543 9974 2544 9978
rect 2548 9974 2549 9978
rect 2553 9974 2554 9978
rect 2458 9973 2554 9974
rect 2458 9969 2459 9973
rect 2463 9969 2464 9973
rect 2458 9968 2464 9969
rect 2458 9964 2459 9968
rect 2463 9964 2464 9968
rect 2548 9969 2549 9973
rect 2553 9969 2554 9973
rect 2548 9968 2554 9969
rect 2458 9963 2464 9964
rect 2458 9959 2459 9963
rect 2463 9959 2464 9963
rect 2458 9958 2464 9959
rect 2458 9954 2459 9958
rect 2463 9954 2464 9958
rect 2458 9953 2464 9954
rect 2458 9949 2459 9953
rect 2463 9949 2464 9953
rect 2458 9948 2464 9949
rect 2458 9944 2459 9948
rect 2463 9944 2464 9948
rect 2458 9943 2464 9944
rect 2458 9939 2459 9943
rect 2463 9939 2464 9943
rect 2458 9938 2464 9939
rect 2458 9934 2459 9938
rect 2463 9934 2464 9938
rect 2458 9933 2464 9934
rect 2458 9929 2459 9933
rect 2463 9929 2464 9933
rect 2458 9928 2464 9929
rect 2458 9924 2459 9928
rect 2463 9924 2464 9928
rect 2458 9923 2464 9924
rect 2458 9919 2459 9923
rect 2463 9919 2464 9923
rect 2458 9918 2464 9919
rect 2458 9914 2459 9918
rect 2463 9914 2464 9918
rect 2458 9913 2464 9914
rect 2458 9909 2459 9913
rect 2463 9909 2464 9913
rect 2458 9908 2464 9909
rect 2458 9904 2459 9908
rect 2463 9904 2464 9908
rect 2458 9903 2464 9904
rect 2458 9899 2459 9903
rect 2463 9899 2464 9903
rect 2458 9898 2464 9899
rect 2458 9894 2459 9898
rect 2463 9894 2464 9898
rect 2458 9893 2464 9894
rect 2458 9889 2459 9893
rect 2463 9889 2464 9893
rect 2458 9888 2464 9889
rect 2458 9884 2459 9888
rect 2463 9884 2464 9888
rect 2458 9883 2464 9884
rect 2458 9879 2459 9883
rect 2463 9879 2464 9883
rect 2458 9878 2464 9879
rect 2458 9874 2459 9878
rect 2463 9874 2464 9878
rect 2458 9873 2464 9874
rect 2458 9869 2459 9873
rect 2463 9869 2464 9873
rect 2458 9868 2464 9869
rect 2458 9864 2459 9868
rect 2463 9864 2464 9868
rect 2458 9863 2464 9864
rect 2458 9859 2459 9863
rect 2463 9859 2464 9863
rect 2458 9858 2464 9859
rect 2458 9854 2459 9858
rect 2463 9854 2464 9858
rect 2458 9853 2464 9854
rect 2458 9849 2459 9853
rect 2463 9849 2464 9853
rect 2548 9964 2549 9968
rect 2553 9964 2554 9968
rect 2548 9963 2554 9964
rect 2548 9959 2549 9963
rect 2553 9959 2554 9963
rect 2548 9958 2554 9959
rect 2548 9954 2549 9958
rect 2553 9954 2554 9958
rect 2548 9953 2554 9954
rect 2548 9949 2549 9953
rect 2553 9949 2554 9953
rect 2548 9948 2554 9949
rect 2548 9944 2549 9948
rect 2553 9944 2554 9948
rect 2548 9943 2554 9944
rect 2548 9939 2549 9943
rect 2553 9939 2554 9943
rect 2548 9938 2554 9939
rect 2548 9934 2549 9938
rect 2553 9934 2554 9938
rect 2548 9933 2554 9934
rect 2548 9929 2549 9933
rect 2553 9929 2554 9933
rect 2548 9928 2554 9929
rect 2548 9924 2549 9928
rect 2553 9924 2554 9928
rect 2548 9923 2554 9924
rect 2548 9919 2549 9923
rect 2553 9919 2554 9923
rect 2548 9918 2554 9919
rect 2548 9914 2549 9918
rect 2553 9914 2554 9918
rect 2548 9913 2554 9914
rect 2548 9909 2549 9913
rect 2553 9909 2554 9913
rect 2548 9908 2554 9909
rect 2548 9904 2549 9908
rect 2553 9904 2554 9908
rect 2548 9903 2554 9904
rect 2548 9899 2549 9903
rect 2553 9899 2554 9903
rect 2548 9898 2554 9899
rect 2548 9894 2549 9898
rect 2553 9894 2554 9898
rect 2548 9893 2554 9894
rect 2548 9889 2549 9893
rect 2553 9889 2554 9893
rect 2548 9888 2554 9889
rect 2548 9884 2549 9888
rect 2553 9884 2554 9888
rect 2548 9883 2554 9884
rect 2548 9879 2549 9883
rect 2553 9879 2554 9883
rect 2548 9878 2554 9879
rect 2548 9874 2549 9878
rect 2553 9874 2554 9878
rect 2548 9873 2554 9874
rect 2548 9869 2549 9873
rect 2553 9869 2554 9873
rect 2548 9868 2554 9869
rect 2548 9864 2549 9868
rect 2553 9864 2554 9868
rect 2548 9863 2554 9864
rect 2548 9859 2549 9863
rect 2553 9859 2554 9863
rect 2548 9858 2554 9859
rect 2548 9854 2549 9858
rect 2553 9854 2554 9858
rect 2548 9853 2554 9854
rect 2458 9848 2464 9849
rect 2458 9844 2459 9848
rect 2463 9844 2464 9848
rect 2548 9849 2549 9853
rect 2553 9849 2554 9853
rect 2548 9848 2554 9849
rect 2548 9844 2549 9848
rect 2553 9844 2554 9848
rect 2458 9843 2554 9844
rect 2458 9839 2459 9843
rect 2463 9839 2464 9843
rect 2468 9839 2469 9843
rect 2473 9839 2474 9843
rect 2478 9839 2479 9843
rect 2483 9839 2484 9843
rect 2488 9839 2489 9843
rect 2493 9839 2494 9843
rect 2498 9839 2499 9843
rect 2503 9839 2504 9843
rect 2508 9839 2509 9843
rect 2513 9839 2514 9843
rect 2518 9839 2519 9843
rect 2523 9839 2524 9843
rect 2528 9839 2529 9843
rect 2533 9839 2534 9843
rect 2538 9839 2539 9843
rect 2543 9839 2544 9843
rect 2548 9839 2549 9843
rect 2553 9839 2554 9843
rect 2458 9838 2554 9839
rect 2619 9965 2691 9967
rect 2619 9961 2621 9965
rect 2625 9961 2628 9965
rect 2632 9961 2633 9965
rect 2637 9961 2638 9965
rect 2642 9961 2643 9965
rect 2647 9961 2648 9965
rect 2652 9961 2653 9965
rect 2657 9961 2658 9965
rect 2662 9961 2663 9965
rect 2667 9961 2668 9965
rect 2672 9961 2673 9965
rect 2677 9961 2678 9965
rect 2682 9961 2685 9965
rect 2689 9961 2691 9965
rect 2619 9959 2691 9961
rect 2619 9958 2627 9959
rect 2619 9954 2621 9958
rect 2625 9954 2627 9958
rect 2619 9953 2627 9954
rect 2683 9958 2691 9959
rect 2683 9954 2685 9958
rect 2689 9954 2691 9958
rect 2683 9953 2691 9954
rect 2619 9949 2621 9953
rect 2625 9949 2627 9953
rect 2619 9948 2627 9949
rect 2619 9944 2621 9948
rect 2625 9944 2627 9948
rect 2619 9943 2627 9944
rect 2619 9939 2621 9943
rect 2625 9939 2627 9943
rect 2619 9938 2627 9939
rect 2619 9934 2621 9938
rect 2625 9934 2627 9938
rect 2619 9933 2627 9934
rect 2619 9929 2621 9933
rect 2625 9929 2627 9933
rect 2619 9928 2627 9929
rect 2619 9924 2621 9928
rect 2625 9924 2627 9928
rect 2619 9923 2627 9924
rect 2619 9919 2621 9923
rect 2625 9919 2627 9923
rect 2619 9918 2627 9919
rect 2619 9914 2621 9918
rect 2625 9914 2627 9918
rect 2619 9913 2627 9914
rect 2619 9909 2621 9913
rect 2625 9909 2627 9913
rect 2619 9908 2627 9909
rect 2619 9904 2621 9908
rect 2625 9904 2627 9908
rect 2619 9903 2627 9904
rect 2619 9899 2621 9903
rect 2625 9899 2627 9903
rect 2619 9898 2627 9899
rect 2619 9894 2621 9898
rect 2625 9894 2627 9898
rect 2619 9893 2627 9894
rect 2619 9889 2621 9893
rect 2625 9889 2627 9893
rect 2619 9888 2627 9889
rect 2619 9884 2621 9888
rect 2625 9884 2627 9888
rect 2619 9883 2627 9884
rect 2619 9879 2621 9883
rect 2625 9879 2627 9883
rect 2619 9878 2627 9879
rect 2619 9874 2621 9878
rect 2625 9874 2627 9878
rect 2619 9873 2627 9874
rect 2619 9869 2621 9873
rect 2625 9869 2627 9873
rect 2619 9868 2627 9869
rect 2619 9864 2621 9868
rect 2625 9864 2627 9868
rect 2683 9949 2685 9953
rect 2689 9949 2691 9953
rect 2683 9948 2691 9949
rect 2683 9944 2685 9948
rect 2689 9944 2691 9948
rect 2683 9943 2691 9944
rect 2683 9939 2685 9943
rect 2689 9939 2691 9943
rect 2683 9938 2691 9939
rect 2683 9934 2685 9938
rect 2689 9934 2691 9938
rect 2683 9933 2691 9934
rect 2683 9929 2685 9933
rect 2689 9929 2691 9933
rect 2683 9928 2691 9929
rect 2683 9924 2685 9928
rect 2689 9924 2691 9928
rect 2683 9923 2691 9924
rect 2683 9919 2685 9923
rect 2689 9919 2691 9923
rect 2683 9918 2691 9919
rect 2683 9914 2685 9918
rect 2689 9914 2691 9918
rect 2683 9913 2691 9914
rect 2683 9909 2685 9913
rect 2689 9909 2691 9913
rect 2683 9908 2691 9909
rect 2683 9904 2685 9908
rect 2689 9904 2691 9908
rect 2683 9903 2691 9904
rect 2683 9899 2685 9903
rect 2689 9899 2691 9903
rect 2683 9898 2691 9899
rect 2683 9894 2685 9898
rect 2689 9894 2691 9898
rect 2683 9893 2691 9894
rect 2683 9889 2685 9893
rect 2689 9889 2691 9893
rect 2683 9888 2691 9889
rect 2683 9884 2685 9888
rect 2689 9884 2691 9888
rect 2683 9883 2691 9884
rect 2683 9879 2685 9883
rect 2689 9879 2691 9883
rect 2683 9878 2691 9879
rect 2683 9874 2685 9878
rect 2689 9874 2691 9878
rect 2683 9873 2691 9874
rect 2683 9869 2685 9873
rect 2689 9869 2691 9873
rect 2683 9868 2691 9869
rect 2683 9864 2685 9868
rect 2689 9864 2691 9868
rect 2619 9863 2627 9864
rect 2619 9859 2621 9863
rect 2625 9859 2627 9863
rect 2619 9858 2627 9859
rect 2683 9863 2691 9864
rect 2683 9859 2685 9863
rect 2689 9859 2691 9863
rect 2683 9858 2691 9859
rect 2619 9856 2691 9858
rect 2619 9852 2621 9856
rect 2625 9852 2628 9856
rect 2632 9852 2633 9856
rect 2637 9852 2638 9856
rect 2642 9852 2643 9856
rect 2647 9852 2648 9856
rect 2652 9852 2653 9856
rect 2657 9852 2658 9856
rect 2662 9852 2663 9856
rect 2667 9852 2668 9856
rect 2672 9852 2673 9856
rect 2677 9852 2678 9856
rect 2682 9852 2685 9856
rect 2689 9852 2691 9856
rect 2619 9850 2691 9852
rect 2767 9978 2863 9979
rect 2767 9974 2768 9978
rect 2772 9974 2773 9978
rect 2777 9974 2778 9978
rect 2782 9974 2783 9978
rect 2787 9974 2788 9978
rect 2792 9974 2793 9978
rect 2797 9974 2798 9978
rect 2802 9974 2803 9978
rect 2807 9974 2808 9978
rect 2812 9974 2813 9978
rect 2817 9974 2818 9978
rect 2822 9974 2823 9978
rect 2827 9974 2828 9978
rect 2832 9974 2833 9978
rect 2837 9974 2838 9978
rect 2842 9974 2843 9978
rect 2847 9974 2848 9978
rect 2852 9974 2853 9978
rect 2857 9974 2858 9978
rect 2862 9974 2863 9978
rect 2767 9973 2863 9974
rect 2767 9969 2768 9973
rect 2772 9969 2773 9973
rect 2767 9968 2773 9969
rect 2767 9964 2768 9968
rect 2772 9964 2773 9968
rect 2857 9969 2858 9973
rect 2862 9969 2863 9973
rect 2857 9968 2863 9969
rect 2767 9963 2773 9964
rect 2767 9959 2768 9963
rect 2772 9959 2773 9963
rect 2767 9958 2773 9959
rect 2767 9954 2768 9958
rect 2772 9954 2773 9958
rect 2767 9953 2773 9954
rect 2767 9949 2768 9953
rect 2772 9949 2773 9953
rect 2767 9948 2773 9949
rect 2767 9944 2768 9948
rect 2772 9944 2773 9948
rect 2767 9943 2773 9944
rect 2767 9939 2768 9943
rect 2772 9939 2773 9943
rect 2767 9938 2773 9939
rect 2767 9934 2768 9938
rect 2772 9934 2773 9938
rect 2767 9933 2773 9934
rect 2767 9929 2768 9933
rect 2772 9929 2773 9933
rect 2767 9928 2773 9929
rect 2767 9924 2768 9928
rect 2772 9924 2773 9928
rect 2767 9923 2773 9924
rect 2767 9919 2768 9923
rect 2772 9919 2773 9923
rect 2767 9918 2773 9919
rect 2767 9914 2768 9918
rect 2772 9914 2773 9918
rect 2767 9913 2773 9914
rect 2767 9909 2768 9913
rect 2772 9909 2773 9913
rect 2767 9908 2773 9909
rect 2767 9904 2768 9908
rect 2772 9904 2773 9908
rect 2767 9903 2773 9904
rect 2767 9899 2768 9903
rect 2772 9899 2773 9903
rect 2767 9898 2773 9899
rect 2767 9894 2768 9898
rect 2772 9894 2773 9898
rect 2767 9893 2773 9894
rect 2767 9889 2768 9893
rect 2772 9889 2773 9893
rect 2767 9888 2773 9889
rect 2767 9884 2768 9888
rect 2772 9884 2773 9888
rect 2767 9883 2773 9884
rect 2767 9879 2768 9883
rect 2772 9879 2773 9883
rect 2767 9878 2773 9879
rect 2767 9874 2768 9878
rect 2772 9874 2773 9878
rect 2767 9873 2773 9874
rect 2767 9869 2768 9873
rect 2772 9869 2773 9873
rect 2767 9868 2773 9869
rect 2767 9864 2768 9868
rect 2772 9864 2773 9868
rect 2767 9863 2773 9864
rect 2767 9859 2768 9863
rect 2772 9859 2773 9863
rect 2767 9858 2773 9859
rect 2767 9854 2768 9858
rect 2772 9854 2773 9858
rect 2767 9853 2773 9854
rect 2767 9849 2768 9853
rect 2772 9849 2773 9853
rect 2857 9964 2858 9968
rect 2862 9964 2863 9968
rect 2857 9963 2863 9964
rect 2857 9959 2858 9963
rect 2862 9959 2863 9963
rect 2857 9958 2863 9959
rect 2857 9954 2858 9958
rect 2862 9954 2863 9958
rect 2857 9953 2863 9954
rect 2857 9949 2858 9953
rect 2862 9949 2863 9953
rect 2857 9948 2863 9949
rect 2857 9944 2858 9948
rect 2862 9944 2863 9948
rect 2857 9943 2863 9944
rect 2857 9939 2858 9943
rect 2862 9939 2863 9943
rect 2857 9938 2863 9939
rect 2857 9934 2858 9938
rect 2862 9934 2863 9938
rect 2857 9933 2863 9934
rect 2857 9929 2858 9933
rect 2862 9929 2863 9933
rect 2857 9928 2863 9929
rect 2857 9924 2858 9928
rect 2862 9924 2863 9928
rect 2857 9923 2863 9924
rect 2857 9919 2858 9923
rect 2862 9919 2863 9923
rect 2857 9918 2863 9919
rect 2857 9914 2858 9918
rect 2862 9914 2863 9918
rect 2857 9913 2863 9914
rect 2857 9909 2858 9913
rect 2862 9909 2863 9913
rect 2857 9908 2863 9909
rect 2857 9904 2858 9908
rect 2862 9904 2863 9908
rect 2857 9903 2863 9904
rect 2857 9899 2858 9903
rect 2862 9899 2863 9903
rect 2857 9898 2863 9899
rect 2857 9894 2858 9898
rect 2862 9894 2863 9898
rect 2857 9893 2863 9894
rect 2857 9889 2858 9893
rect 2862 9889 2863 9893
rect 2857 9888 2863 9889
rect 2857 9884 2858 9888
rect 2862 9884 2863 9888
rect 2857 9883 2863 9884
rect 2857 9879 2858 9883
rect 2862 9879 2863 9883
rect 2857 9878 2863 9879
rect 2857 9874 2858 9878
rect 2862 9874 2863 9878
rect 2857 9873 2863 9874
rect 2857 9869 2858 9873
rect 2862 9869 2863 9873
rect 2857 9868 2863 9869
rect 2857 9864 2858 9868
rect 2862 9864 2863 9868
rect 2857 9863 2863 9864
rect 2857 9859 2858 9863
rect 2862 9859 2863 9863
rect 2857 9858 2863 9859
rect 2857 9854 2858 9858
rect 2862 9854 2863 9858
rect 2857 9853 2863 9854
rect 2767 9848 2773 9849
rect 2767 9844 2768 9848
rect 2772 9844 2773 9848
rect 2857 9849 2858 9853
rect 2862 9849 2863 9853
rect 2857 9848 2863 9849
rect 2857 9844 2858 9848
rect 2862 9844 2863 9848
rect 2767 9843 2863 9844
rect 2767 9839 2768 9843
rect 2772 9839 2773 9843
rect 2777 9839 2778 9843
rect 2782 9839 2783 9843
rect 2787 9839 2788 9843
rect 2792 9839 2793 9843
rect 2797 9839 2798 9843
rect 2802 9839 2803 9843
rect 2807 9839 2808 9843
rect 2812 9839 2813 9843
rect 2817 9839 2818 9843
rect 2822 9839 2823 9843
rect 2827 9839 2828 9843
rect 2832 9839 2833 9843
rect 2837 9839 2838 9843
rect 2842 9839 2843 9843
rect 2847 9839 2848 9843
rect 2852 9839 2853 9843
rect 2857 9839 2858 9843
rect 2862 9839 2863 9843
rect 2767 9838 2863 9839
rect 2928 9965 3000 9967
rect 2928 9961 2930 9965
rect 2934 9961 2937 9965
rect 2941 9961 2942 9965
rect 2946 9961 2947 9965
rect 2951 9961 2952 9965
rect 2956 9961 2957 9965
rect 2961 9961 2962 9965
rect 2966 9961 2967 9965
rect 2971 9961 2972 9965
rect 2976 9961 2977 9965
rect 2981 9961 2982 9965
rect 2986 9961 2987 9965
rect 2991 9961 2994 9965
rect 2998 9961 3000 9965
rect 2928 9959 3000 9961
rect 2928 9958 2936 9959
rect 2928 9954 2930 9958
rect 2934 9954 2936 9958
rect 2928 9953 2936 9954
rect 2992 9958 3000 9959
rect 2992 9954 2994 9958
rect 2998 9954 3000 9958
rect 2992 9953 3000 9954
rect 2928 9949 2930 9953
rect 2934 9949 2936 9953
rect 2928 9948 2936 9949
rect 2928 9944 2930 9948
rect 2934 9944 2936 9948
rect 2928 9943 2936 9944
rect 2928 9939 2930 9943
rect 2934 9939 2936 9943
rect 2928 9938 2936 9939
rect 2928 9934 2930 9938
rect 2934 9934 2936 9938
rect 2928 9933 2936 9934
rect 2928 9929 2930 9933
rect 2934 9929 2936 9933
rect 2928 9928 2936 9929
rect 2928 9924 2930 9928
rect 2934 9924 2936 9928
rect 2928 9923 2936 9924
rect 2928 9919 2930 9923
rect 2934 9919 2936 9923
rect 2928 9918 2936 9919
rect 2928 9914 2930 9918
rect 2934 9914 2936 9918
rect 2928 9913 2936 9914
rect 2928 9909 2930 9913
rect 2934 9909 2936 9913
rect 2928 9908 2936 9909
rect 2928 9904 2930 9908
rect 2934 9904 2936 9908
rect 2928 9903 2936 9904
rect 2928 9899 2930 9903
rect 2934 9899 2936 9903
rect 2928 9898 2936 9899
rect 2928 9894 2930 9898
rect 2934 9894 2936 9898
rect 2928 9893 2936 9894
rect 2928 9889 2930 9893
rect 2934 9889 2936 9893
rect 2928 9888 2936 9889
rect 2928 9884 2930 9888
rect 2934 9884 2936 9888
rect 2928 9883 2936 9884
rect 2928 9879 2930 9883
rect 2934 9879 2936 9883
rect 2928 9878 2936 9879
rect 2928 9874 2930 9878
rect 2934 9874 2936 9878
rect 2928 9873 2936 9874
rect 2928 9869 2930 9873
rect 2934 9869 2936 9873
rect 2928 9868 2936 9869
rect 2928 9864 2930 9868
rect 2934 9864 2936 9868
rect 2992 9949 2994 9953
rect 2998 9949 3000 9953
rect 2992 9948 3000 9949
rect 2992 9944 2994 9948
rect 2998 9944 3000 9948
rect 2992 9943 3000 9944
rect 2992 9939 2994 9943
rect 2998 9939 3000 9943
rect 2992 9938 3000 9939
rect 2992 9934 2994 9938
rect 2998 9934 3000 9938
rect 2992 9933 3000 9934
rect 2992 9929 2994 9933
rect 2998 9929 3000 9933
rect 2992 9928 3000 9929
rect 2992 9924 2994 9928
rect 2998 9924 3000 9928
rect 2992 9923 3000 9924
rect 2992 9919 2994 9923
rect 2998 9919 3000 9923
rect 2992 9918 3000 9919
rect 2992 9914 2994 9918
rect 2998 9914 3000 9918
rect 2992 9913 3000 9914
rect 2992 9909 2994 9913
rect 2998 9909 3000 9913
rect 2992 9908 3000 9909
rect 2992 9904 2994 9908
rect 2998 9904 3000 9908
rect 2992 9903 3000 9904
rect 2992 9899 2994 9903
rect 2998 9899 3000 9903
rect 2992 9898 3000 9899
rect 2992 9894 2994 9898
rect 2998 9894 3000 9898
rect 2992 9893 3000 9894
rect 2992 9889 2994 9893
rect 2998 9889 3000 9893
rect 2992 9888 3000 9889
rect 2992 9884 2994 9888
rect 2998 9884 3000 9888
rect 2992 9883 3000 9884
rect 2992 9879 2994 9883
rect 2998 9879 3000 9883
rect 2992 9878 3000 9879
rect 2992 9874 2994 9878
rect 2998 9874 3000 9878
rect 2992 9873 3000 9874
rect 2992 9869 2994 9873
rect 2998 9869 3000 9873
rect 2992 9868 3000 9869
rect 2992 9864 2994 9868
rect 2998 9864 3000 9868
rect 2928 9863 2936 9864
rect 2928 9859 2930 9863
rect 2934 9859 2936 9863
rect 2928 9858 2936 9859
rect 2992 9863 3000 9864
rect 2992 9859 2994 9863
rect 2998 9859 3000 9863
rect 2992 9858 3000 9859
rect 2928 9856 3000 9858
rect 2928 9852 2930 9856
rect 2934 9852 2937 9856
rect 2941 9852 2942 9856
rect 2946 9852 2947 9856
rect 2951 9852 2952 9856
rect 2956 9852 2957 9856
rect 2961 9852 2962 9856
rect 2966 9852 2967 9856
rect 2971 9852 2972 9856
rect 2976 9852 2977 9856
rect 2981 9852 2982 9856
rect 2986 9852 2987 9856
rect 2991 9852 2994 9856
rect 2998 9852 3000 9856
rect 2928 9850 3000 9852
rect 3076 9978 3172 9979
rect 3076 9974 3077 9978
rect 3081 9974 3082 9978
rect 3086 9974 3087 9978
rect 3091 9974 3092 9978
rect 3096 9974 3097 9978
rect 3101 9974 3102 9978
rect 3106 9974 3107 9978
rect 3111 9974 3112 9978
rect 3116 9974 3117 9978
rect 3121 9974 3122 9978
rect 3126 9974 3127 9978
rect 3131 9974 3132 9978
rect 3136 9974 3137 9978
rect 3141 9974 3142 9978
rect 3146 9974 3147 9978
rect 3151 9974 3152 9978
rect 3156 9974 3157 9978
rect 3161 9974 3162 9978
rect 3166 9974 3167 9978
rect 3171 9974 3172 9978
rect 3076 9973 3172 9974
rect 3076 9969 3077 9973
rect 3081 9969 3082 9973
rect 3076 9968 3082 9969
rect 3076 9964 3077 9968
rect 3081 9964 3082 9968
rect 3166 9969 3167 9973
rect 3171 9969 3172 9973
rect 3166 9968 3172 9969
rect 3076 9963 3082 9964
rect 3076 9959 3077 9963
rect 3081 9959 3082 9963
rect 3076 9958 3082 9959
rect 3076 9954 3077 9958
rect 3081 9954 3082 9958
rect 3076 9953 3082 9954
rect 3076 9949 3077 9953
rect 3081 9949 3082 9953
rect 3076 9948 3082 9949
rect 3076 9944 3077 9948
rect 3081 9944 3082 9948
rect 3076 9943 3082 9944
rect 3076 9939 3077 9943
rect 3081 9939 3082 9943
rect 3076 9938 3082 9939
rect 3076 9934 3077 9938
rect 3081 9934 3082 9938
rect 3076 9933 3082 9934
rect 3076 9929 3077 9933
rect 3081 9929 3082 9933
rect 3076 9928 3082 9929
rect 3076 9924 3077 9928
rect 3081 9924 3082 9928
rect 3076 9923 3082 9924
rect 3076 9919 3077 9923
rect 3081 9919 3082 9923
rect 3076 9918 3082 9919
rect 3076 9914 3077 9918
rect 3081 9914 3082 9918
rect 3076 9913 3082 9914
rect 3076 9909 3077 9913
rect 3081 9909 3082 9913
rect 3076 9908 3082 9909
rect 3076 9904 3077 9908
rect 3081 9904 3082 9908
rect 3076 9903 3082 9904
rect 3076 9899 3077 9903
rect 3081 9899 3082 9903
rect 3076 9898 3082 9899
rect 3076 9894 3077 9898
rect 3081 9894 3082 9898
rect 3076 9893 3082 9894
rect 3076 9889 3077 9893
rect 3081 9889 3082 9893
rect 3076 9888 3082 9889
rect 3076 9884 3077 9888
rect 3081 9884 3082 9888
rect 3076 9883 3082 9884
rect 3076 9879 3077 9883
rect 3081 9879 3082 9883
rect 3076 9878 3082 9879
rect 3076 9874 3077 9878
rect 3081 9874 3082 9878
rect 3076 9873 3082 9874
rect 3076 9869 3077 9873
rect 3081 9869 3082 9873
rect 3076 9868 3082 9869
rect 3076 9864 3077 9868
rect 3081 9864 3082 9868
rect 3076 9863 3082 9864
rect 3076 9859 3077 9863
rect 3081 9859 3082 9863
rect 3076 9858 3082 9859
rect 3076 9854 3077 9858
rect 3081 9854 3082 9858
rect 3076 9853 3082 9854
rect 3076 9849 3077 9853
rect 3081 9849 3082 9853
rect 3166 9964 3167 9968
rect 3171 9964 3172 9968
rect 3166 9963 3172 9964
rect 3166 9959 3167 9963
rect 3171 9959 3172 9963
rect 3166 9958 3172 9959
rect 3166 9954 3167 9958
rect 3171 9954 3172 9958
rect 3166 9953 3172 9954
rect 3166 9949 3167 9953
rect 3171 9949 3172 9953
rect 3166 9948 3172 9949
rect 3166 9944 3167 9948
rect 3171 9944 3172 9948
rect 3166 9943 3172 9944
rect 3166 9939 3167 9943
rect 3171 9939 3172 9943
rect 3166 9938 3172 9939
rect 3166 9934 3167 9938
rect 3171 9934 3172 9938
rect 3166 9933 3172 9934
rect 3166 9929 3167 9933
rect 3171 9929 3172 9933
rect 3166 9928 3172 9929
rect 3166 9924 3167 9928
rect 3171 9924 3172 9928
rect 3166 9923 3172 9924
rect 3166 9919 3167 9923
rect 3171 9919 3172 9923
rect 3166 9918 3172 9919
rect 3166 9914 3167 9918
rect 3171 9914 3172 9918
rect 3166 9913 3172 9914
rect 3166 9909 3167 9913
rect 3171 9909 3172 9913
rect 3166 9908 3172 9909
rect 3166 9904 3167 9908
rect 3171 9904 3172 9908
rect 3166 9903 3172 9904
rect 3166 9899 3167 9903
rect 3171 9899 3172 9903
rect 3166 9898 3172 9899
rect 3166 9894 3167 9898
rect 3171 9894 3172 9898
rect 3166 9893 3172 9894
rect 3166 9889 3167 9893
rect 3171 9889 3172 9893
rect 3166 9888 3172 9889
rect 3166 9884 3167 9888
rect 3171 9884 3172 9888
rect 3166 9883 3172 9884
rect 3166 9879 3167 9883
rect 3171 9879 3172 9883
rect 3166 9878 3172 9879
rect 3166 9874 3167 9878
rect 3171 9874 3172 9878
rect 3166 9873 3172 9874
rect 3166 9869 3167 9873
rect 3171 9869 3172 9873
rect 3166 9868 3172 9869
rect 3166 9864 3167 9868
rect 3171 9864 3172 9868
rect 3166 9863 3172 9864
rect 3166 9859 3167 9863
rect 3171 9859 3172 9863
rect 3166 9858 3172 9859
rect 3166 9854 3167 9858
rect 3171 9854 3172 9858
rect 3166 9853 3172 9854
rect 3076 9848 3082 9849
rect 3076 9844 3077 9848
rect 3081 9844 3082 9848
rect 3166 9849 3167 9853
rect 3171 9849 3172 9853
rect 3166 9848 3172 9849
rect 3166 9844 3167 9848
rect 3171 9844 3172 9848
rect 3076 9843 3172 9844
rect 3076 9839 3077 9843
rect 3081 9839 3082 9843
rect 3086 9839 3087 9843
rect 3091 9839 3092 9843
rect 3096 9839 3097 9843
rect 3101 9839 3102 9843
rect 3106 9839 3107 9843
rect 3111 9839 3112 9843
rect 3116 9839 3117 9843
rect 3121 9839 3122 9843
rect 3126 9839 3127 9843
rect 3131 9839 3132 9843
rect 3136 9839 3137 9843
rect 3141 9839 3142 9843
rect 3146 9839 3147 9843
rect 3151 9839 3152 9843
rect 3156 9839 3157 9843
rect 3161 9839 3162 9843
rect 3166 9839 3167 9843
rect 3171 9839 3172 9843
rect 3076 9838 3172 9839
rect 3237 9965 3309 9967
rect 3237 9961 3239 9965
rect 3243 9961 3246 9965
rect 3250 9961 3251 9965
rect 3255 9961 3256 9965
rect 3260 9961 3261 9965
rect 3265 9961 3266 9965
rect 3270 9961 3271 9965
rect 3275 9961 3276 9965
rect 3280 9961 3281 9965
rect 3285 9961 3286 9965
rect 3290 9961 3291 9965
rect 3295 9961 3296 9965
rect 3300 9961 3303 9965
rect 3307 9961 3309 9965
rect 3237 9959 3309 9961
rect 3237 9958 3245 9959
rect 3237 9954 3239 9958
rect 3243 9954 3245 9958
rect 3237 9953 3245 9954
rect 3301 9958 3309 9959
rect 3301 9954 3303 9958
rect 3307 9954 3309 9958
rect 3301 9953 3309 9954
rect 3237 9949 3239 9953
rect 3243 9949 3245 9953
rect 3237 9948 3245 9949
rect 3237 9944 3239 9948
rect 3243 9944 3245 9948
rect 3237 9943 3245 9944
rect 3237 9939 3239 9943
rect 3243 9939 3245 9943
rect 3237 9938 3245 9939
rect 3237 9934 3239 9938
rect 3243 9934 3245 9938
rect 3237 9933 3245 9934
rect 3237 9929 3239 9933
rect 3243 9929 3245 9933
rect 3237 9928 3245 9929
rect 3237 9924 3239 9928
rect 3243 9924 3245 9928
rect 3237 9923 3245 9924
rect 3237 9919 3239 9923
rect 3243 9919 3245 9923
rect 3237 9918 3245 9919
rect 3237 9914 3239 9918
rect 3243 9914 3245 9918
rect 3237 9913 3245 9914
rect 3237 9909 3239 9913
rect 3243 9909 3245 9913
rect 3237 9908 3245 9909
rect 3237 9904 3239 9908
rect 3243 9904 3245 9908
rect 3237 9903 3245 9904
rect 3237 9899 3239 9903
rect 3243 9899 3245 9903
rect 3237 9898 3245 9899
rect 3237 9894 3239 9898
rect 3243 9894 3245 9898
rect 3237 9893 3245 9894
rect 3237 9889 3239 9893
rect 3243 9889 3245 9893
rect 3237 9888 3245 9889
rect 3237 9884 3239 9888
rect 3243 9884 3245 9888
rect 3237 9883 3245 9884
rect 3237 9879 3239 9883
rect 3243 9879 3245 9883
rect 3237 9878 3245 9879
rect 3237 9874 3239 9878
rect 3243 9874 3245 9878
rect 3237 9873 3245 9874
rect 3237 9869 3239 9873
rect 3243 9869 3245 9873
rect 3237 9868 3245 9869
rect 3237 9864 3239 9868
rect 3243 9864 3245 9868
rect 3301 9949 3303 9953
rect 3307 9949 3309 9953
rect 3301 9948 3309 9949
rect 3301 9944 3303 9948
rect 3307 9944 3309 9948
rect 3301 9943 3309 9944
rect 3301 9939 3303 9943
rect 3307 9939 3309 9943
rect 3301 9938 3309 9939
rect 3301 9934 3303 9938
rect 3307 9934 3309 9938
rect 3301 9933 3309 9934
rect 3301 9929 3303 9933
rect 3307 9929 3309 9933
rect 3301 9928 3309 9929
rect 3301 9924 3303 9928
rect 3307 9924 3309 9928
rect 3301 9923 3309 9924
rect 3301 9919 3303 9923
rect 3307 9919 3309 9923
rect 3301 9918 3309 9919
rect 3301 9914 3303 9918
rect 3307 9914 3309 9918
rect 3301 9913 3309 9914
rect 3301 9909 3303 9913
rect 3307 9909 3309 9913
rect 3301 9908 3309 9909
rect 3301 9904 3303 9908
rect 3307 9904 3309 9908
rect 3301 9903 3309 9904
rect 3301 9899 3303 9903
rect 3307 9899 3309 9903
rect 3301 9898 3309 9899
rect 3301 9894 3303 9898
rect 3307 9894 3309 9898
rect 3301 9893 3309 9894
rect 3301 9889 3303 9893
rect 3307 9889 3309 9893
rect 3301 9888 3309 9889
rect 3301 9884 3303 9888
rect 3307 9884 3309 9888
rect 3301 9883 3309 9884
rect 3301 9879 3303 9883
rect 3307 9879 3309 9883
rect 3301 9878 3309 9879
rect 3301 9874 3303 9878
rect 3307 9874 3309 9878
rect 3301 9873 3309 9874
rect 3301 9869 3303 9873
rect 3307 9869 3309 9873
rect 3301 9868 3309 9869
rect 3301 9864 3303 9868
rect 3307 9864 3309 9868
rect 3237 9863 3245 9864
rect 3237 9859 3239 9863
rect 3243 9859 3245 9863
rect 3237 9858 3245 9859
rect 3301 9863 3309 9864
rect 3301 9859 3303 9863
rect 3307 9859 3309 9863
rect 3301 9858 3309 9859
rect 3237 9856 3309 9858
rect 3237 9852 3239 9856
rect 3243 9852 3246 9856
rect 3250 9852 3251 9856
rect 3255 9852 3256 9856
rect 3260 9852 3261 9856
rect 3265 9852 3266 9856
rect 3270 9852 3271 9856
rect 3275 9852 3276 9856
rect 3280 9852 3281 9856
rect 3285 9852 3286 9856
rect 3290 9852 3291 9856
rect 3295 9852 3296 9856
rect 3300 9852 3303 9856
rect 3307 9852 3309 9856
rect 3237 9850 3309 9852
rect 3385 9978 3481 9979
rect 3385 9974 3386 9978
rect 3390 9974 3391 9978
rect 3395 9974 3396 9978
rect 3400 9974 3401 9978
rect 3405 9974 3406 9978
rect 3410 9974 3411 9978
rect 3415 9974 3416 9978
rect 3420 9974 3421 9978
rect 3425 9974 3426 9978
rect 3430 9974 3431 9978
rect 3435 9974 3436 9978
rect 3440 9974 3441 9978
rect 3445 9974 3446 9978
rect 3450 9974 3451 9978
rect 3455 9974 3456 9978
rect 3460 9974 3461 9978
rect 3465 9974 3466 9978
rect 3470 9974 3471 9978
rect 3475 9974 3476 9978
rect 3480 9974 3481 9978
rect 3385 9973 3481 9974
rect 3385 9969 3386 9973
rect 3390 9969 3391 9973
rect 3385 9968 3391 9969
rect 3385 9964 3386 9968
rect 3390 9964 3391 9968
rect 3475 9969 3476 9973
rect 3480 9969 3481 9973
rect 3475 9968 3481 9969
rect 3385 9963 3391 9964
rect 3385 9959 3386 9963
rect 3390 9959 3391 9963
rect 3385 9958 3391 9959
rect 3385 9954 3386 9958
rect 3390 9954 3391 9958
rect 3385 9953 3391 9954
rect 3385 9949 3386 9953
rect 3390 9949 3391 9953
rect 3385 9948 3391 9949
rect 3385 9944 3386 9948
rect 3390 9944 3391 9948
rect 3385 9943 3391 9944
rect 3385 9939 3386 9943
rect 3390 9939 3391 9943
rect 3385 9938 3391 9939
rect 3385 9934 3386 9938
rect 3390 9934 3391 9938
rect 3385 9933 3391 9934
rect 3385 9929 3386 9933
rect 3390 9929 3391 9933
rect 3385 9928 3391 9929
rect 3385 9924 3386 9928
rect 3390 9924 3391 9928
rect 3385 9923 3391 9924
rect 3385 9919 3386 9923
rect 3390 9919 3391 9923
rect 3385 9918 3391 9919
rect 3385 9914 3386 9918
rect 3390 9914 3391 9918
rect 3385 9913 3391 9914
rect 3385 9909 3386 9913
rect 3390 9909 3391 9913
rect 3385 9908 3391 9909
rect 3385 9904 3386 9908
rect 3390 9904 3391 9908
rect 3385 9903 3391 9904
rect 3385 9899 3386 9903
rect 3390 9899 3391 9903
rect 3385 9898 3391 9899
rect 3385 9894 3386 9898
rect 3390 9894 3391 9898
rect 3385 9893 3391 9894
rect 3385 9889 3386 9893
rect 3390 9889 3391 9893
rect 3385 9888 3391 9889
rect 3385 9884 3386 9888
rect 3390 9884 3391 9888
rect 3385 9883 3391 9884
rect 3385 9879 3386 9883
rect 3390 9879 3391 9883
rect 3385 9878 3391 9879
rect 3385 9874 3386 9878
rect 3390 9874 3391 9878
rect 3385 9873 3391 9874
rect 3385 9869 3386 9873
rect 3390 9869 3391 9873
rect 3385 9868 3391 9869
rect 3385 9864 3386 9868
rect 3390 9864 3391 9868
rect 3385 9863 3391 9864
rect 3385 9859 3386 9863
rect 3390 9859 3391 9863
rect 3385 9858 3391 9859
rect 3385 9854 3386 9858
rect 3390 9854 3391 9858
rect 3385 9853 3391 9854
rect 3385 9849 3386 9853
rect 3390 9849 3391 9853
rect 3475 9964 3476 9968
rect 3480 9964 3481 9968
rect 3475 9963 3481 9964
rect 3475 9959 3476 9963
rect 3480 9959 3481 9963
rect 3475 9958 3481 9959
rect 3475 9954 3476 9958
rect 3480 9954 3481 9958
rect 3475 9953 3481 9954
rect 3475 9949 3476 9953
rect 3480 9949 3481 9953
rect 3475 9948 3481 9949
rect 3475 9944 3476 9948
rect 3480 9944 3481 9948
rect 3475 9943 3481 9944
rect 3475 9939 3476 9943
rect 3480 9939 3481 9943
rect 3475 9938 3481 9939
rect 3475 9934 3476 9938
rect 3480 9934 3481 9938
rect 3475 9933 3481 9934
rect 3475 9929 3476 9933
rect 3480 9929 3481 9933
rect 3475 9928 3481 9929
rect 3475 9924 3476 9928
rect 3480 9924 3481 9928
rect 3475 9923 3481 9924
rect 3475 9919 3476 9923
rect 3480 9919 3481 9923
rect 3475 9918 3481 9919
rect 3475 9914 3476 9918
rect 3480 9914 3481 9918
rect 3475 9913 3481 9914
rect 3475 9909 3476 9913
rect 3480 9909 3481 9913
rect 3475 9908 3481 9909
rect 3475 9904 3476 9908
rect 3480 9904 3481 9908
rect 3475 9903 3481 9904
rect 3475 9899 3476 9903
rect 3480 9899 3481 9903
rect 3475 9898 3481 9899
rect 3475 9894 3476 9898
rect 3480 9894 3481 9898
rect 3475 9893 3481 9894
rect 3475 9889 3476 9893
rect 3480 9889 3481 9893
rect 3475 9888 3481 9889
rect 3475 9884 3476 9888
rect 3480 9884 3481 9888
rect 3475 9883 3481 9884
rect 3475 9879 3476 9883
rect 3480 9879 3481 9883
rect 3475 9878 3481 9879
rect 3475 9874 3476 9878
rect 3480 9874 3481 9878
rect 3475 9873 3481 9874
rect 3475 9869 3476 9873
rect 3480 9869 3481 9873
rect 3475 9868 3481 9869
rect 3475 9864 3476 9868
rect 3480 9864 3481 9868
rect 3475 9863 3481 9864
rect 3475 9859 3476 9863
rect 3480 9859 3481 9863
rect 3475 9858 3481 9859
rect 3475 9854 3476 9858
rect 3480 9854 3481 9858
rect 3475 9853 3481 9854
rect 3385 9848 3391 9849
rect 3385 9844 3386 9848
rect 3390 9844 3391 9848
rect 3475 9849 3476 9853
rect 3480 9849 3481 9853
rect 3475 9848 3481 9849
rect 3475 9844 3476 9848
rect 3480 9844 3481 9848
rect 3385 9843 3481 9844
rect 3385 9839 3386 9843
rect 3390 9839 3391 9843
rect 3395 9839 3396 9843
rect 3400 9839 3401 9843
rect 3405 9839 3406 9843
rect 3410 9839 3411 9843
rect 3415 9839 3416 9843
rect 3420 9839 3421 9843
rect 3425 9839 3426 9843
rect 3430 9839 3431 9843
rect 3435 9839 3436 9843
rect 3440 9839 3441 9843
rect 3445 9839 3446 9843
rect 3450 9839 3451 9843
rect 3455 9839 3456 9843
rect 3460 9839 3461 9843
rect 3465 9839 3466 9843
rect 3470 9839 3471 9843
rect 3475 9839 3476 9843
rect 3480 9839 3481 9843
rect 3385 9838 3481 9839
rect 3546 9965 3618 9967
rect 3546 9961 3548 9965
rect 3552 9961 3555 9965
rect 3559 9961 3560 9965
rect 3564 9961 3565 9965
rect 3569 9961 3570 9965
rect 3574 9961 3575 9965
rect 3579 9961 3580 9965
rect 3584 9961 3585 9965
rect 3589 9961 3590 9965
rect 3594 9961 3595 9965
rect 3599 9961 3600 9965
rect 3604 9961 3605 9965
rect 3609 9961 3612 9965
rect 3616 9961 3618 9965
rect 3546 9959 3618 9961
rect 3546 9958 3554 9959
rect 3546 9954 3548 9958
rect 3552 9954 3554 9958
rect 3546 9953 3554 9954
rect 3610 9958 3618 9959
rect 3610 9954 3612 9958
rect 3616 9954 3618 9958
rect 3610 9953 3618 9954
rect 3546 9949 3548 9953
rect 3552 9949 3554 9953
rect 3546 9948 3554 9949
rect 3546 9944 3548 9948
rect 3552 9944 3554 9948
rect 3546 9943 3554 9944
rect 3546 9939 3548 9943
rect 3552 9939 3554 9943
rect 3546 9938 3554 9939
rect 3546 9934 3548 9938
rect 3552 9934 3554 9938
rect 3546 9933 3554 9934
rect 3546 9929 3548 9933
rect 3552 9929 3554 9933
rect 3546 9928 3554 9929
rect 3546 9924 3548 9928
rect 3552 9924 3554 9928
rect 3546 9923 3554 9924
rect 3546 9919 3548 9923
rect 3552 9919 3554 9923
rect 3546 9918 3554 9919
rect 3546 9914 3548 9918
rect 3552 9914 3554 9918
rect 3546 9913 3554 9914
rect 3546 9909 3548 9913
rect 3552 9909 3554 9913
rect 3546 9908 3554 9909
rect 3546 9904 3548 9908
rect 3552 9904 3554 9908
rect 3546 9903 3554 9904
rect 3546 9899 3548 9903
rect 3552 9899 3554 9903
rect 3546 9898 3554 9899
rect 3546 9894 3548 9898
rect 3552 9894 3554 9898
rect 3546 9893 3554 9894
rect 3546 9889 3548 9893
rect 3552 9889 3554 9893
rect 3546 9888 3554 9889
rect 3546 9884 3548 9888
rect 3552 9884 3554 9888
rect 3546 9883 3554 9884
rect 3546 9879 3548 9883
rect 3552 9879 3554 9883
rect 3546 9878 3554 9879
rect 3546 9874 3548 9878
rect 3552 9874 3554 9878
rect 3546 9873 3554 9874
rect 3546 9869 3548 9873
rect 3552 9869 3554 9873
rect 3546 9868 3554 9869
rect 3546 9864 3548 9868
rect 3552 9864 3554 9868
rect 3610 9949 3612 9953
rect 3616 9949 3618 9953
rect 3610 9948 3618 9949
rect 3610 9944 3612 9948
rect 3616 9944 3618 9948
rect 3610 9943 3618 9944
rect 3610 9939 3612 9943
rect 3616 9939 3618 9943
rect 3610 9938 3618 9939
rect 3610 9934 3612 9938
rect 3616 9934 3618 9938
rect 3610 9933 3618 9934
rect 3610 9929 3612 9933
rect 3616 9929 3618 9933
rect 3610 9928 3618 9929
rect 3610 9924 3612 9928
rect 3616 9924 3618 9928
rect 3610 9923 3618 9924
rect 3610 9919 3612 9923
rect 3616 9919 3618 9923
rect 3610 9918 3618 9919
rect 3610 9914 3612 9918
rect 3616 9914 3618 9918
rect 3610 9913 3618 9914
rect 3610 9909 3612 9913
rect 3616 9909 3618 9913
rect 3610 9908 3618 9909
rect 3610 9904 3612 9908
rect 3616 9904 3618 9908
rect 3610 9903 3618 9904
rect 3610 9899 3612 9903
rect 3616 9899 3618 9903
rect 3610 9898 3618 9899
rect 3610 9894 3612 9898
rect 3616 9894 3618 9898
rect 3610 9893 3618 9894
rect 3610 9889 3612 9893
rect 3616 9889 3618 9893
rect 3610 9888 3618 9889
rect 3610 9884 3612 9888
rect 3616 9884 3618 9888
rect 3610 9883 3618 9884
rect 3610 9879 3612 9883
rect 3616 9879 3618 9883
rect 3610 9878 3618 9879
rect 3610 9874 3612 9878
rect 3616 9874 3618 9878
rect 3610 9873 3618 9874
rect 3610 9869 3612 9873
rect 3616 9869 3618 9873
rect 3610 9868 3618 9869
rect 3610 9864 3612 9868
rect 3616 9864 3618 9868
rect 3546 9863 3554 9864
rect 3546 9859 3548 9863
rect 3552 9859 3554 9863
rect 3546 9858 3554 9859
rect 3610 9863 3618 9864
rect 3610 9859 3612 9863
rect 3616 9859 3618 9863
rect 3610 9858 3618 9859
rect 3546 9856 3618 9858
rect 3546 9852 3548 9856
rect 3552 9852 3555 9856
rect 3559 9852 3560 9856
rect 3564 9852 3565 9856
rect 3569 9852 3570 9856
rect 3574 9852 3575 9856
rect 3579 9852 3580 9856
rect 3584 9852 3585 9856
rect 3589 9852 3590 9856
rect 3594 9852 3595 9856
rect 3599 9852 3600 9856
rect 3604 9852 3605 9856
rect 3609 9852 3612 9856
rect 3616 9852 3618 9856
rect 3546 9850 3618 9852
rect 3694 9978 3790 9979
rect 3694 9974 3695 9978
rect 3699 9974 3700 9978
rect 3704 9974 3705 9978
rect 3709 9974 3710 9978
rect 3714 9974 3715 9978
rect 3719 9974 3720 9978
rect 3724 9974 3725 9978
rect 3729 9974 3730 9978
rect 3734 9974 3735 9978
rect 3739 9974 3740 9978
rect 3744 9974 3745 9978
rect 3749 9974 3750 9978
rect 3754 9974 3755 9978
rect 3759 9974 3760 9978
rect 3764 9974 3765 9978
rect 3769 9974 3770 9978
rect 3774 9974 3775 9978
rect 3779 9974 3780 9978
rect 3784 9974 3785 9978
rect 3789 9974 3790 9978
rect 3694 9973 3790 9974
rect 3694 9969 3695 9973
rect 3699 9969 3700 9973
rect 3694 9968 3700 9969
rect 3694 9964 3695 9968
rect 3699 9964 3700 9968
rect 3784 9969 3785 9973
rect 3789 9969 3790 9973
rect 3784 9968 3790 9969
rect 3694 9963 3700 9964
rect 3694 9959 3695 9963
rect 3699 9959 3700 9963
rect 3694 9958 3700 9959
rect 3694 9954 3695 9958
rect 3699 9954 3700 9958
rect 3694 9953 3700 9954
rect 3694 9949 3695 9953
rect 3699 9949 3700 9953
rect 3694 9948 3700 9949
rect 3694 9944 3695 9948
rect 3699 9944 3700 9948
rect 3694 9943 3700 9944
rect 3694 9939 3695 9943
rect 3699 9939 3700 9943
rect 3694 9938 3700 9939
rect 3694 9934 3695 9938
rect 3699 9934 3700 9938
rect 3694 9933 3700 9934
rect 3694 9929 3695 9933
rect 3699 9929 3700 9933
rect 3694 9928 3700 9929
rect 3694 9924 3695 9928
rect 3699 9924 3700 9928
rect 3694 9923 3700 9924
rect 3694 9919 3695 9923
rect 3699 9919 3700 9923
rect 3694 9918 3700 9919
rect 3694 9914 3695 9918
rect 3699 9914 3700 9918
rect 3694 9913 3700 9914
rect 3694 9909 3695 9913
rect 3699 9909 3700 9913
rect 3694 9908 3700 9909
rect 3694 9904 3695 9908
rect 3699 9904 3700 9908
rect 3694 9903 3700 9904
rect 3694 9899 3695 9903
rect 3699 9899 3700 9903
rect 3694 9898 3700 9899
rect 3694 9894 3695 9898
rect 3699 9894 3700 9898
rect 3694 9893 3700 9894
rect 3694 9889 3695 9893
rect 3699 9889 3700 9893
rect 3694 9888 3700 9889
rect 3694 9884 3695 9888
rect 3699 9884 3700 9888
rect 3694 9883 3700 9884
rect 3694 9879 3695 9883
rect 3699 9879 3700 9883
rect 3694 9878 3700 9879
rect 3694 9874 3695 9878
rect 3699 9874 3700 9878
rect 3694 9873 3700 9874
rect 3694 9869 3695 9873
rect 3699 9869 3700 9873
rect 3694 9868 3700 9869
rect 3694 9864 3695 9868
rect 3699 9864 3700 9868
rect 3694 9863 3700 9864
rect 3694 9859 3695 9863
rect 3699 9859 3700 9863
rect 3694 9858 3700 9859
rect 3694 9854 3695 9858
rect 3699 9854 3700 9858
rect 3694 9853 3700 9854
rect 3694 9849 3695 9853
rect 3699 9849 3700 9853
rect 3784 9964 3785 9968
rect 3789 9964 3790 9968
rect 3784 9963 3790 9964
rect 3784 9959 3785 9963
rect 3789 9959 3790 9963
rect 3784 9958 3790 9959
rect 3784 9954 3785 9958
rect 3789 9954 3790 9958
rect 3784 9953 3790 9954
rect 3784 9949 3785 9953
rect 3789 9949 3790 9953
rect 3784 9948 3790 9949
rect 3784 9944 3785 9948
rect 3789 9944 3790 9948
rect 3784 9943 3790 9944
rect 3784 9939 3785 9943
rect 3789 9939 3790 9943
rect 3784 9938 3790 9939
rect 3784 9934 3785 9938
rect 3789 9934 3790 9938
rect 3784 9933 3790 9934
rect 3784 9929 3785 9933
rect 3789 9929 3790 9933
rect 3784 9928 3790 9929
rect 3784 9924 3785 9928
rect 3789 9924 3790 9928
rect 3784 9923 3790 9924
rect 3784 9919 3785 9923
rect 3789 9919 3790 9923
rect 3784 9918 3790 9919
rect 3784 9914 3785 9918
rect 3789 9914 3790 9918
rect 3784 9913 3790 9914
rect 3784 9909 3785 9913
rect 3789 9909 3790 9913
rect 3784 9908 3790 9909
rect 3784 9904 3785 9908
rect 3789 9904 3790 9908
rect 3784 9903 3790 9904
rect 3784 9899 3785 9903
rect 3789 9899 3790 9903
rect 3784 9898 3790 9899
rect 3784 9894 3785 9898
rect 3789 9894 3790 9898
rect 3784 9893 3790 9894
rect 3784 9889 3785 9893
rect 3789 9889 3790 9893
rect 3784 9888 3790 9889
rect 3784 9884 3785 9888
rect 3789 9884 3790 9888
rect 3784 9883 3790 9884
rect 3784 9879 3785 9883
rect 3789 9879 3790 9883
rect 3784 9878 3790 9879
rect 3784 9874 3785 9878
rect 3789 9874 3790 9878
rect 3784 9873 3790 9874
rect 3784 9869 3785 9873
rect 3789 9869 3790 9873
rect 3784 9868 3790 9869
rect 3784 9864 3785 9868
rect 3789 9864 3790 9868
rect 3784 9863 3790 9864
rect 3784 9859 3785 9863
rect 3789 9859 3790 9863
rect 3784 9858 3790 9859
rect 3784 9854 3785 9858
rect 3789 9854 3790 9858
rect 3784 9853 3790 9854
rect 3694 9848 3700 9849
rect 3694 9844 3695 9848
rect 3699 9844 3700 9848
rect 3784 9849 3785 9853
rect 3789 9849 3790 9853
rect 3784 9848 3790 9849
rect 3784 9844 3785 9848
rect 3789 9844 3790 9848
rect 3694 9843 3790 9844
rect 3694 9839 3695 9843
rect 3699 9839 3700 9843
rect 3704 9839 3705 9843
rect 3709 9839 3710 9843
rect 3714 9839 3715 9843
rect 3719 9839 3720 9843
rect 3724 9839 3725 9843
rect 3729 9839 3730 9843
rect 3734 9839 3735 9843
rect 3739 9839 3740 9843
rect 3744 9839 3745 9843
rect 3749 9839 3750 9843
rect 3754 9839 3755 9843
rect 3759 9839 3760 9843
rect 3764 9839 3765 9843
rect 3769 9839 3770 9843
rect 3774 9839 3775 9843
rect 3779 9839 3780 9843
rect 3784 9839 3785 9843
rect 3789 9839 3790 9843
rect 3694 9838 3790 9839
rect 3855 9965 3927 9967
rect 3855 9961 3857 9965
rect 3861 9961 3864 9965
rect 3868 9961 3869 9965
rect 3873 9961 3874 9965
rect 3878 9961 3879 9965
rect 3883 9961 3884 9965
rect 3888 9961 3889 9965
rect 3893 9961 3894 9965
rect 3898 9961 3899 9965
rect 3903 9961 3904 9965
rect 3908 9961 3909 9965
rect 3913 9961 3914 9965
rect 3918 9961 3921 9965
rect 3925 9961 3927 9965
rect 3855 9959 3927 9961
rect 3855 9958 3863 9959
rect 3855 9954 3857 9958
rect 3861 9954 3863 9958
rect 3855 9953 3863 9954
rect 3919 9958 3927 9959
rect 3919 9954 3921 9958
rect 3925 9954 3927 9958
rect 3919 9953 3927 9954
rect 3855 9949 3857 9953
rect 3861 9949 3863 9953
rect 3855 9948 3863 9949
rect 3855 9944 3857 9948
rect 3861 9944 3863 9948
rect 3855 9943 3863 9944
rect 3855 9939 3857 9943
rect 3861 9939 3863 9943
rect 3855 9938 3863 9939
rect 3855 9934 3857 9938
rect 3861 9934 3863 9938
rect 3855 9933 3863 9934
rect 3855 9929 3857 9933
rect 3861 9929 3863 9933
rect 3855 9928 3863 9929
rect 3855 9924 3857 9928
rect 3861 9924 3863 9928
rect 3855 9923 3863 9924
rect 3855 9919 3857 9923
rect 3861 9919 3863 9923
rect 3855 9918 3863 9919
rect 3855 9914 3857 9918
rect 3861 9914 3863 9918
rect 3855 9913 3863 9914
rect 3855 9909 3857 9913
rect 3861 9909 3863 9913
rect 3855 9908 3863 9909
rect 3855 9904 3857 9908
rect 3861 9904 3863 9908
rect 3855 9903 3863 9904
rect 3855 9899 3857 9903
rect 3861 9899 3863 9903
rect 3855 9898 3863 9899
rect 3855 9894 3857 9898
rect 3861 9894 3863 9898
rect 3855 9893 3863 9894
rect 3855 9889 3857 9893
rect 3861 9889 3863 9893
rect 3855 9888 3863 9889
rect 3855 9884 3857 9888
rect 3861 9884 3863 9888
rect 3855 9883 3863 9884
rect 3855 9879 3857 9883
rect 3861 9879 3863 9883
rect 3855 9878 3863 9879
rect 3855 9874 3857 9878
rect 3861 9874 3863 9878
rect 3855 9873 3863 9874
rect 3855 9869 3857 9873
rect 3861 9869 3863 9873
rect 3855 9868 3863 9869
rect 3855 9864 3857 9868
rect 3861 9864 3863 9868
rect 3919 9949 3921 9953
rect 3925 9949 3927 9953
rect 3919 9948 3927 9949
rect 3919 9944 3921 9948
rect 3925 9944 3927 9948
rect 3919 9943 3927 9944
rect 3919 9939 3921 9943
rect 3925 9939 3927 9943
rect 3919 9938 3927 9939
rect 3919 9934 3921 9938
rect 3925 9934 3927 9938
rect 3919 9933 3927 9934
rect 3919 9929 3921 9933
rect 3925 9929 3927 9933
rect 3919 9928 3927 9929
rect 3919 9924 3921 9928
rect 3925 9924 3927 9928
rect 3919 9923 3927 9924
rect 3919 9919 3921 9923
rect 3925 9919 3927 9923
rect 3919 9918 3927 9919
rect 3919 9914 3921 9918
rect 3925 9914 3927 9918
rect 3919 9913 3927 9914
rect 3919 9909 3921 9913
rect 3925 9909 3927 9913
rect 3919 9908 3927 9909
rect 3919 9904 3921 9908
rect 3925 9904 3927 9908
rect 3919 9903 3927 9904
rect 3919 9899 3921 9903
rect 3925 9899 3927 9903
rect 3919 9898 3927 9899
rect 3919 9894 3921 9898
rect 3925 9894 3927 9898
rect 3919 9893 3927 9894
rect 3919 9889 3921 9893
rect 3925 9889 3927 9893
rect 3919 9888 3927 9889
rect 3919 9884 3921 9888
rect 3925 9884 3927 9888
rect 3919 9883 3927 9884
rect 3919 9879 3921 9883
rect 3925 9879 3927 9883
rect 3919 9878 3927 9879
rect 3919 9874 3921 9878
rect 3925 9874 3927 9878
rect 3919 9873 3927 9874
rect 3919 9869 3921 9873
rect 3925 9869 3927 9873
rect 3919 9868 3927 9869
rect 3919 9864 3921 9868
rect 3925 9864 3927 9868
rect 3855 9863 3863 9864
rect 3855 9859 3857 9863
rect 3861 9859 3863 9863
rect 3855 9858 3863 9859
rect 3919 9863 3927 9864
rect 3919 9859 3921 9863
rect 3925 9859 3927 9863
rect 3919 9858 3927 9859
rect 3855 9856 3927 9858
rect 3855 9852 3857 9856
rect 3861 9852 3864 9856
rect 3868 9852 3869 9856
rect 3873 9852 3874 9856
rect 3878 9852 3879 9856
rect 3883 9852 3884 9856
rect 3888 9852 3889 9856
rect 3893 9852 3894 9856
rect 3898 9852 3899 9856
rect 3903 9852 3904 9856
rect 3908 9852 3909 9856
rect 3913 9852 3914 9856
rect 3918 9852 3921 9856
rect 3925 9852 3927 9856
rect 3855 9850 3927 9852
rect 4003 9978 4099 9979
rect 4003 9974 4004 9978
rect 4008 9974 4009 9978
rect 4013 9974 4014 9978
rect 4018 9974 4019 9978
rect 4023 9974 4024 9978
rect 4028 9974 4029 9978
rect 4033 9974 4034 9978
rect 4038 9974 4039 9978
rect 4043 9974 4044 9978
rect 4048 9974 4049 9978
rect 4053 9974 4054 9978
rect 4058 9974 4059 9978
rect 4063 9974 4064 9978
rect 4068 9974 4069 9978
rect 4073 9974 4074 9978
rect 4078 9974 4079 9978
rect 4083 9974 4084 9978
rect 4088 9974 4089 9978
rect 4093 9974 4094 9978
rect 4098 9974 4099 9978
rect 4003 9973 4099 9974
rect 4003 9969 4004 9973
rect 4008 9969 4009 9973
rect 4003 9968 4009 9969
rect 4003 9964 4004 9968
rect 4008 9964 4009 9968
rect 4093 9969 4094 9973
rect 4098 9969 4099 9973
rect 4093 9968 4099 9969
rect 4003 9963 4009 9964
rect 4003 9959 4004 9963
rect 4008 9959 4009 9963
rect 4003 9958 4009 9959
rect 4003 9954 4004 9958
rect 4008 9954 4009 9958
rect 4003 9953 4009 9954
rect 4003 9949 4004 9953
rect 4008 9949 4009 9953
rect 4003 9948 4009 9949
rect 4003 9944 4004 9948
rect 4008 9944 4009 9948
rect 4003 9943 4009 9944
rect 4003 9939 4004 9943
rect 4008 9939 4009 9943
rect 4003 9938 4009 9939
rect 4003 9934 4004 9938
rect 4008 9934 4009 9938
rect 4003 9933 4009 9934
rect 4003 9929 4004 9933
rect 4008 9929 4009 9933
rect 4003 9928 4009 9929
rect 4003 9924 4004 9928
rect 4008 9924 4009 9928
rect 4003 9923 4009 9924
rect 4003 9919 4004 9923
rect 4008 9919 4009 9923
rect 4003 9918 4009 9919
rect 4003 9914 4004 9918
rect 4008 9914 4009 9918
rect 4003 9913 4009 9914
rect 4003 9909 4004 9913
rect 4008 9909 4009 9913
rect 4003 9908 4009 9909
rect 4003 9904 4004 9908
rect 4008 9904 4009 9908
rect 4003 9903 4009 9904
rect 4003 9899 4004 9903
rect 4008 9899 4009 9903
rect 4003 9898 4009 9899
rect 4003 9894 4004 9898
rect 4008 9894 4009 9898
rect 4003 9893 4009 9894
rect 4003 9889 4004 9893
rect 4008 9889 4009 9893
rect 4003 9888 4009 9889
rect 4003 9884 4004 9888
rect 4008 9884 4009 9888
rect 4003 9883 4009 9884
rect 4003 9879 4004 9883
rect 4008 9879 4009 9883
rect 4003 9878 4009 9879
rect 4003 9874 4004 9878
rect 4008 9874 4009 9878
rect 4003 9873 4009 9874
rect 4003 9869 4004 9873
rect 4008 9869 4009 9873
rect 4003 9868 4009 9869
rect 4003 9864 4004 9868
rect 4008 9864 4009 9868
rect 4003 9863 4009 9864
rect 4003 9859 4004 9863
rect 4008 9859 4009 9863
rect 4003 9858 4009 9859
rect 4003 9854 4004 9858
rect 4008 9854 4009 9858
rect 4003 9853 4009 9854
rect 4003 9849 4004 9853
rect 4008 9849 4009 9853
rect 4093 9964 4094 9968
rect 4098 9964 4099 9968
rect 4093 9963 4099 9964
rect 4093 9959 4094 9963
rect 4098 9959 4099 9963
rect 4093 9958 4099 9959
rect 4093 9954 4094 9958
rect 4098 9954 4099 9958
rect 4093 9953 4099 9954
rect 4093 9949 4094 9953
rect 4098 9949 4099 9953
rect 4093 9948 4099 9949
rect 4093 9944 4094 9948
rect 4098 9944 4099 9948
rect 4093 9943 4099 9944
rect 4093 9939 4094 9943
rect 4098 9939 4099 9943
rect 4093 9938 4099 9939
rect 4093 9934 4094 9938
rect 4098 9934 4099 9938
rect 4093 9933 4099 9934
rect 4093 9929 4094 9933
rect 4098 9929 4099 9933
rect 4093 9928 4099 9929
rect 4093 9924 4094 9928
rect 4098 9924 4099 9928
rect 4093 9923 4099 9924
rect 4093 9919 4094 9923
rect 4098 9919 4099 9923
rect 4093 9918 4099 9919
rect 4093 9914 4094 9918
rect 4098 9914 4099 9918
rect 4093 9913 4099 9914
rect 4093 9909 4094 9913
rect 4098 9909 4099 9913
rect 4093 9908 4099 9909
rect 4093 9904 4094 9908
rect 4098 9904 4099 9908
rect 4093 9903 4099 9904
rect 4093 9899 4094 9903
rect 4098 9899 4099 9903
rect 4093 9898 4099 9899
rect 4093 9894 4094 9898
rect 4098 9894 4099 9898
rect 4093 9893 4099 9894
rect 4093 9889 4094 9893
rect 4098 9889 4099 9893
rect 4093 9888 4099 9889
rect 4093 9884 4094 9888
rect 4098 9884 4099 9888
rect 4093 9883 4099 9884
rect 4093 9879 4094 9883
rect 4098 9879 4099 9883
rect 4093 9878 4099 9879
rect 4093 9874 4094 9878
rect 4098 9874 4099 9878
rect 4093 9873 4099 9874
rect 4093 9869 4094 9873
rect 4098 9869 4099 9873
rect 4093 9868 4099 9869
rect 4093 9864 4094 9868
rect 4098 9864 4099 9868
rect 4093 9863 4099 9864
rect 4093 9859 4094 9863
rect 4098 9859 4099 9863
rect 4093 9858 4099 9859
rect 4093 9854 4094 9858
rect 4098 9854 4099 9858
rect 4093 9853 4099 9854
rect 4003 9848 4009 9849
rect 4003 9844 4004 9848
rect 4008 9844 4009 9848
rect 4093 9849 4094 9853
rect 4098 9849 4099 9853
rect 4093 9848 4099 9849
rect 4093 9844 4094 9848
rect 4098 9844 4099 9848
rect 4003 9843 4099 9844
rect 4003 9839 4004 9843
rect 4008 9839 4009 9843
rect 4013 9839 4014 9843
rect 4018 9839 4019 9843
rect 4023 9839 4024 9843
rect 4028 9839 4029 9843
rect 4033 9839 4034 9843
rect 4038 9839 4039 9843
rect 4043 9839 4044 9843
rect 4048 9839 4049 9843
rect 4053 9839 4054 9843
rect 4058 9839 4059 9843
rect 4063 9839 4064 9843
rect 4068 9839 4069 9843
rect 4073 9839 4074 9843
rect 4078 9839 4079 9843
rect 4083 9839 4084 9843
rect 4088 9839 4089 9843
rect 4093 9839 4094 9843
rect 4098 9839 4099 9843
rect 4003 9838 4099 9839
rect 655 9720 4517 9724
rect 655 9716 802 9720
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 821 9716 831 9720
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 850 9716 860 9720
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 879 9716 889 9720
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 908 9716 918 9720
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 937 9716 1319 9720
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1338 9716 1628 9720
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1647 9716 1937 9720
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1956 9716 2246 9720
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2265 9716 2555 9720
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2574 9716 2864 9720
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2883 9716 3173 9720
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3192 9716 3482 9720
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3501 9716 3791 9720
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3810 9716 4100 9720
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4119 9716 4292 9720
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4311 9716 4318 9720
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4337 9716 4344 9720
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4363 9716 4370 9720
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4389 9716 4396 9720
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4415 9716 4517 9720
rect 655 9710 4517 9716
rect 655 9706 802 9710
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 821 9706 831 9710
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 850 9706 860 9710
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 879 9706 889 9710
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 908 9706 918 9710
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 937 9706 1319 9710
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1338 9706 1628 9710
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1647 9706 1937 9710
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1956 9706 2246 9710
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2265 9706 2555 9710
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2574 9706 2864 9710
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2883 9706 3173 9710
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3192 9706 3482 9710
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3501 9706 3791 9710
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3810 9706 4100 9710
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4119 9706 4292 9710
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4311 9706 4318 9710
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4337 9706 4344 9710
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4363 9706 4370 9710
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4389 9706 4396 9710
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4415 9706 4517 9710
rect 655 9700 4517 9706
rect 655 9696 802 9700
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 821 9696 831 9700
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 850 9696 860 9700
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 879 9696 889 9700
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 908 9696 918 9700
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 937 9696 1319 9700
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1338 9696 1628 9700
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1647 9696 1937 9700
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1956 9696 2246 9700
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2265 9696 2555 9700
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2574 9696 2864 9700
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2883 9696 3173 9700
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3192 9696 3482 9700
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3501 9696 3791 9700
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3810 9696 4100 9700
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4119 9696 4292 9700
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4311 9696 4318 9700
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4337 9696 4344 9700
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4363 9696 4370 9700
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4389 9696 4396 9700
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4415 9696 4517 9700
rect 655 9690 4517 9696
rect 655 9686 802 9690
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 821 9686 831 9690
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 850 9686 860 9690
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 879 9686 889 9690
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 908 9686 918 9690
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 937 9686 1319 9690
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1338 9686 1628 9690
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1647 9686 1937 9690
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 1956 9686 2246 9690
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2265 9686 2555 9690
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2574 9686 2864 9690
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 2883 9686 3173 9690
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3192 9686 3482 9690
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 3501 9686 3791 9690
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 3810 9686 4100 9690
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4119 9686 4292 9690
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4311 9686 4318 9690
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4337 9686 4344 9690
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4363 9686 4370 9690
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4389 9686 4396 9690
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 4415 9686 4517 9690
rect 655 9684 4517 9686
rect 655 9622 695 9684
rect 655 9618 659 9622
rect 663 9618 669 9622
rect 673 9618 679 9622
rect 683 9618 689 9622
rect 693 9618 695 9622
rect 655 9617 695 9618
rect 655 9613 659 9617
rect 663 9613 669 9617
rect 673 9613 679 9617
rect 683 9613 689 9617
rect 693 9613 695 9617
rect 655 9612 695 9613
rect 655 9608 659 9612
rect 663 9608 669 9612
rect 673 9608 679 9612
rect 683 9608 689 9612
rect 693 9608 695 9612
rect 655 9607 695 9608
rect 655 9603 659 9607
rect 663 9603 669 9607
rect 673 9603 679 9607
rect 683 9603 689 9607
rect 693 9603 695 9607
rect 655 9596 695 9603
rect 655 9592 659 9596
rect 663 9592 669 9596
rect 673 9592 679 9596
rect 683 9592 689 9596
rect 693 9592 695 9596
rect 655 9591 695 9592
rect 655 9587 659 9591
rect 663 9587 669 9591
rect 673 9587 679 9591
rect 683 9587 689 9591
rect 693 9587 695 9591
rect 655 9586 695 9587
rect 655 9582 659 9586
rect 663 9582 669 9586
rect 673 9582 679 9586
rect 683 9582 689 9586
rect 693 9582 695 9586
rect 655 9581 695 9582
rect 655 9577 659 9581
rect 663 9577 669 9581
rect 673 9577 679 9581
rect 683 9577 689 9581
rect 693 9577 695 9581
rect 655 9570 695 9577
rect 655 9566 659 9570
rect 663 9566 669 9570
rect 673 9566 679 9570
rect 683 9566 689 9570
rect 693 9566 695 9570
rect 655 9565 695 9566
rect 655 9561 659 9565
rect 663 9561 669 9565
rect 673 9561 679 9565
rect 683 9561 689 9565
rect 693 9561 695 9565
rect 655 9560 695 9561
rect 655 9556 659 9560
rect 663 9556 669 9560
rect 673 9556 679 9560
rect 683 9556 689 9560
rect 693 9556 695 9560
rect 655 9555 695 9556
rect 655 9551 659 9555
rect 663 9551 669 9555
rect 673 9551 679 9555
rect 683 9551 689 9555
rect 693 9551 695 9555
rect 655 9544 695 9551
rect 655 9540 659 9544
rect 663 9540 669 9544
rect 673 9540 679 9544
rect 683 9540 689 9544
rect 693 9540 695 9544
rect 655 9539 695 9540
rect 655 9535 659 9539
rect 663 9535 669 9539
rect 673 9535 679 9539
rect 683 9535 689 9539
rect 693 9535 695 9539
rect 655 9534 695 9535
rect 655 9530 659 9534
rect 663 9530 669 9534
rect 673 9530 679 9534
rect 683 9530 689 9534
rect 693 9530 695 9534
rect 655 9529 695 9530
rect 655 9525 659 9529
rect 663 9525 669 9529
rect 673 9525 679 9529
rect 683 9525 689 9529
rect 693 9525 695 9529
rect 655 9518 695 9525
rect 655 9514 659 9518
rect 663 9514 669 9518
rect 673 9514 679 9518
rect 683 9514 689 9518
rect 693 9514 695 9518
rect 655 9513 695 9514
rect 655 9509 659 9513
rect 663 9509 669 9513
rect 673 9509 679 9513
rect 683 9509 689 9513
rect 693 9509 695 9513
rect 655 9508 695 9509
rect 655 9504 659 9508
rect 663 9504 669 9508
rect 673 9504 679 9508
rect 683 9504 689 9508
rect 693 9504 695 9508
rect 655 9503 695 9504
rect 655 9499 659 9503
rect 663 9499 669 9503
rect 673 9499 679 9503
rect 683 9499 689 9503
rect 693 9499 695 9503
rect 655 9325 695 9499
rect 4477 9577 4517 9684
rect 4477 9573 4479 9577
rect 4483 9573 4489 9577
rect 4493 9573 4499 9577
rect 4503 9573 4509 9577
rect 4513 9573 4517 9577
rect 4477 9572 4517 9573
rect 4477 9568 4479 9572
rect 4483 9568 4489 9572
rect 4493 9568 4499 9572
rect 4503 9568 4509 9572
rect 4513 9568 4517 9572
rect 4477 9567 4517 9568
rect 4477 9563 4479 9567
rect 4483 9563 4489 9567
rect 4493 9563 4499 9567
rect 4503 9563 4509 9567
rect 4513 9563 4517 9567
rect 4477 9562 4517 9563
rect 4477 9558 4479 9562
rect 4483 9558 4489 9562
rect 4493 9558 4499 9562
rect 4503 9558 4509 9562
rect 4513 9558 4517 9562
rect 4477 9548 4517 9558
rect 4477 9544 4479 9548
rect 4483 9544 4489 9548
rect 4493 9544 4499 9548
rect 4503 9544 4509 9548
rect 4513 9544 4517 9548
rect 4477 9543 4517 9544
rect 4477 9539 4479 9543
rect 4483 9539 4489 9543
rect 4493 9539 4499 9543
rect 4503 9539 4509 9543
rect 4513 9539 4517 9543
rect 4477 9538 4517 9539
rect 4477 9534 4479 9538
rect 4483 9534 4489 9538
rect 4493 9534 4499 9538
rect 4503 9534 4509 9538
rect 4513 9534 4517 9538
rect 4477 9533 4517 9534
rect 4477 9529 4479 9533
rect 4483 9529 4489 9533
rect 4493 9529 4499 9533
rect 4503 9529 4509 9533
rect 4513 9529 4517 9533
rect 4477 9519 4517 9529
rect 4477 9515 4479 9519
rect 4483 9515 4489 9519
rect 4493 9515 4499 9519
rect 4503 9515 4509 9519
rect 4513 9515 4517 9519
rect 4477 9514 4517 9515
rect 4477 9510 4479 9514
rect 4483 9510 4489 9514
rect 4493 9510 4499 9514
rect 4503 9510 4509 9514
rect 4513 9510 4517 9514
rect 4477 9509 4517 9510
rect 4477 9505 4479 9509
rect 4483 9505 4489 9509
rect 4493 9505 4499 9509
rect 4503 9505 4509 9509
rect 4513 9505 4517 9509
rect 4477 9504 4517 9505
rect 4477 9500 4479 9504
rect 4483 9500 4489 9504
rect 4493 9500 4499 9504
rect 4503 9500 4509 9504
rect 4513 9500 4517 9504
rect 4477 9490 4517 9500
rect 4477 9486 4479 9490
rect 4483 9486 4489 9490
rect 4493 9486 4499 9490
rect 4503 9486 4509 9490
rect 4513 9486 4517 9490
rect 4477 9485 4517 9486
rect 4477 9481 4479 9485
rect 4483 9481 4489 9485
rect 4493 9481 4499 9485
rect 4503 9481 4509 9485
rect 4513 9481 4517 9485
rect 4477 9480 4517 9481
rect 4477 9476 4479 9480
rect 4483 9476 4489 9480
rect 4493 9476 4499 9480
rect 4503 9476 4509 9480
rect 4513 9476 4517 9480
rect 4477 9475 4517 9476
rect 4477 9471 4479 9475
rect 4483 9471 4489 9475
rect 4493 9471 4499 9475
rect 4503 9471 4509 9475
rect 4513 9471 4517 9475
rect 4477 9461 4517 9471
rect 4477 9457 4479 9461
rect 4483 9457 4489 9461
rect 4493 9457 4499 9461
rect 4503 9457 4509 9461
rect 4513 9457 4517 9461
rect 4477 9456 4517 9457
rect 4477 9452 4479 9456
rect 4483 9452 4489 9456
rect 4493 9452 4499 9456
rect 4503 9452 4509 9456
rect 4513 9452 4517 9456
rect 4477 9451 4517 9452
rect 4477 9447 4479 9451
rect 4483 9447 4489 9451
rect 4493 9447 4499 9451
rect 4503 9447 4509 9451
rect 4513 9447 4517 9451
rect 4477 9446 4517 9447
rect 4477 9442 4479 9446
rect 4483 9442 4489 9446
rect 4493 9442 4499 9446
rect 4503 9442 4509 9446
rect 4513 9442 4517 9446
rect 655 9321 659 9325
rect 663 9321 669 9325
rect 673 9321 679 9325
rect 683 9321 689 9325
rect 693 9321 695 9325
rect 655 9320 695 9321
rect 655 9316 659 9320
rect 663 9316 669 9320
rect 673 9316 679 9320
rect 683 9316 689 9320
rect 693 9316 695 9320
rect 655 9315 695 9316
rect 655 9311 659 9315
rect 663 9311 669 9315
rect 673 9311 679 9315
rect 683 9311 689 9315
rect 693 9311 695 9315
rect 655 9310 695 9311
rect 655 9306 659 9310
rect 663 9306 669 9310
rect 673 9306 679 9310
rect 683 9306 689 9310
rect 693 9306 695 9310
rect 655 9016 695 9306
rect 4477 9060 4517 9442
rect 4477 9056 4479 9060
rect 4483 9056 4489 9060
rect 4493 9056 4499 9060
rect 4503 9056 4509 9060
rect 4513 9056 4517 9060
rect 4477 9055 4517 9056
rect 4477 9051 4479 9055
rect 4483 9051 4489 9055
rect 4493 9051 4499 9055
rect 4503 9051 4509 9055
rect 4513 9051 4517 9055
rect 4477 9050 4517 9051
rect 4477 9046 4479 9050
rect 4483 9046 4489 9050
rect 4493 9046 4499 9050
rect 4503 9046 4509 9050
rect 4513 9046 4517 9050
rect 4477 9045 4517 9046
rect 4477 9041 4479 9045
rect 4483 9041 4489 9045
rect 4493 9041 4499 9045
rect 4503 9041 4509 9045
rect 4513 9041 4517 9045
rect 655 9012 659 9016
rect 663 9012 669 9016
rect 673 9012 679 9016
rect 683 9012 689 9016
rect 693 9012 695 9016
rect 655 9011 695 9012
rect 655 9007 659 9011
rect 663 9007 669 9011
rect 673 9007 679 9011
rect 683 9007 689 9011
rect 693 9007 695 9011
rect 655 9006 695 9007
rect 655 9002 659 9006
rect 663 9002 669 9006
rect 673 9002 679 9006
rect 683 9002 689 9006
rect 693 9002 695 9006
rect 655 9001 695 9002
rect 655 8997 659 9001
rect 663 8997 669 9001
rect 673 8997 679 9001
rect 683 8997 689 9001
rect 693 8997 695 9001
rect 655 8707 695 8997
rect 4477 8751 4517 9041
rect 4477 8747 4479 8751
rect 4483 8747 4489 8751
rect 4493 8747 4499 8751
rect 4503 8747 4509 8751
rect 4513 8747 4517 8751
rect 4477 8746 4517 8747
rect 4477 8742 4479 8746
rect 4483 8742 4489 8746
rect 4493 8742 4499 8746
rect 4503 8742 4509 8746
rect 4513 8742 4517 8746
rect 4477 8741 4517 8742
rect 4477 8737 4479 8741
rect 4483 8737 4489 8741
rect 4493 8737 4499 8741
rect 4503 8737 4509 8741
rect 4513 8737 4517 8741
rect 4477 8736 4517 8737
rect 4477 8732 4479 8736
rect 4483 8732 4489 8736
rect 4493 8732 4499 8736
rect 4503 8732 4509 8736
rect 4513 8732 4517 8736
rect 655 8703 659 8707
rect 663 8703 669 8707
rect 673 8703 679 8707
rect 683 8703 689 8707
rect 693 8703 695 8707
rect 655 8702 695 8703
rect 655 8698 659 8702
rect 663 8698 669 8702
rect 673 8698 679 8702
rect 683 8698 689 8702
rect 693 8698 695 8702
rect 655 8697 695 8698
rect 655 8693 659 8697
rect 663 8693 669 8697
rect 673 8693 679 8697
rect 683 8693 689 8697
rect 693 8693 695 8697
rect 655 8692 695 8693
rect 655 8688 659 8692
rect 663 8688 669 8692
rect 673 8688 679 8692
rect 683 8688 689 8692
rect 693 8688 695 8692
rect 655 8398 695 8688
rect 4477 8442 4517 8732
rect 4477 8438 4479 8442
rect 4483 8438 4489 8442
rect 4493 8438 4499 8442
rect 4503 8438 4509 8442
rect 4513 8438 4517 8442
rect 4477 8437 4517 8438
rect 4477 8433 4479 8437
rect 4483 8433 4489 8437
rect 4493 8433 4499 8437
rect 4503 8433 4509 8437
rect 4513 8433 4517 8437
rect 4477 8432 4517 8433
rect 4477 8428 4479 8432
rect 4483 8428 4489 8432
rect 4493 8428 4499 8432
rect 4503 8428 4509 8432
rect 4513 8428 4517 8432
rect 4477 8427 4517 8428
rect 4477 8423 4479 8427
rect 4483 8423 4489 8427
rect 4493 8423 4499 8427
rect 4503 8423 4509 8427
rect 4513 8423 4517 8427
rect 655 8394 659 8398
rect 663 8394 669 8398
rect 673 8394 679 8398
rect 683 8394 689 8398
rect 693 8394 695 8398
rect 655 8393 695 8394
rect 655 8389 659 8393
rect 663 8389 669 8393
rect 673 8389 679 8393
rect 683 8389 689 8393
rect 693 8389 695 8393
rect 655 8388 695 8389
rect 655 8384 659 8388
rect 663 8384 669 8388
rect 673 8384 679 8388
rect 683 8384 689 8388
rect 693 8384 695 8388
rect 655 8383 695 8384
rect 655 8379 659 8383
rect 663 8379 669 8383
rect 673 8379 679 8383
rect 683 8379 689 8383
rect 693 8379 695 8383
rect 655 8089 695 8379
rect 4477 8133 4517 8423
rect 4477 8129 4479 8133
rect 4483 8129 4489 8133
rect 4493 8129 4499 8133
rect 4503 8129 4509 8133
rect 4513 8129 4517 8133
rect 4477 8128 4517 8129
rect 4477 8124 4479 8128
rect 4483 8124 4489 8128
rect 4493 8124 4499 8128
rect 4503 8124 4509 8128
rect 4513 8124 4517 8128
rect 4477 8123 4517 8124
rect 4477 8119 4479 8123
rect 4483 8119 4489 8123
rect 4493 8119 4499 8123
rect 4503 8119 4509 8123
rect 4513 8119 4517 8123
rect 4477 8118 4517 8119
rect 4477 8114 4479 8118
rect 4483 8114 4489 8118
rect 4493 8114 4499 8118
rect 4503 8114 4509 8118
rect 4513 8114 4517 8118
rect 4477 8102 4517 8114
rect 4477 8098 4479 8102
rect 4483 8098 4489 8102
rect 4493 8098 4499 8102
rect 4503 8098 4509 8102
rect 4513 8098 4517 8102
rect 4477 8097 4517 8098
rect 655 8085 659 8089
rect 663 8085 669 8089
rect 673 8085 679 8089
rect 683 8085 689 8089
rect 693 8085 695 8089
rect 4477 8093 4479 8097
rect 4483 8093 4489 8097
rect 4493 8093 4499 8097
rect 4503 8093 4509 8097
rect 4513 8093 4517 8097
rect 4477 8092 4517 8093
rect 4477 8088 4479 8092
rect 4483 8088 4489 8092
rect 4493 8088 4499 8092
rect 4503 8088 4509 8092
rect 4513 8088 4517 8092
rect 4477 8087 4517 8088
rect 655 8084 695 8085
rect 655 8080 659 8084
rect 663 8080 669 8084
rect 673 8080 679 8084
rect 683 8080 689 8084
rect 693 8080 695 8084
rect 4477 8083 4479 8087
rect 4483 8083 4489 8087
rect 4493 8083 4499 8087
rect 4503 8083 4509 8087
rect 4513 8083 4517 8087
rect 655 8079 695 8080
rect 655 8075 659 8079
rect 663 8075 669 8079
rect 673 8075 679 8079
rect 683 8075 689 8079
rect 693 8075 695 8079
rect 655 8074 695 8075
rect 655 8070 659 8074
rect 663 8070 669 8074
rect 673 8070 679 8074
rect 683 8070 689 8074
rect 693 8070 695 8074
rect 655 7780 695 8070
rect 655 7776 659 7780
rect 663 7776 669 7780
rect 673 7776 679 7780
rect 683 7776 689 7780
rect 693 7776 695 7780
rect 655 7775 695 7776
rect 655 7771 659 7775
rect 663 7771 669 7775
rect 673 7771 679 7775
rect 683 7771 689 7775
rect 693 7771 695 7775
rect 655 7770 695 7771
rect 655 7766 659 7770
rect 663 7766 669 7770
rect 673 7766 679 7770
rect 683 7766 689 7770
rect 693 7766 695 7770
rect 655 7765 695 7766
rect 655 7761 659 7765
rect 663 7761 669 7765
rect 673 7761 679 7765
rect 683 7761 689 7765
rect 693 7761 695 7765
rect 655 7471 695 7761
rect 4477 7793 4517 8083
rect 4477 7789 4479 7793
rect 4483 7789 4489 7793
rect 4493 7789 4499 7793
rect 4503 7789 4509 7793
rect 4513 7789 4517 7793
rect 4477 7788 4517 7789
rect 4477 7784 4479 7788
rect 4483 7784 4489 7788
rect 4493 7784 4499 7788
rect 4503 7784 4509 7788
rect 4513 7784 4517 7788
rect 4477 7783 4517 7784
rect 4477 7779 4479 7783
rect 4483 7779 4489 7783
rect 4493 7779 4499 7783
rect 4503 7779 4509 7783
rect 4513 7779 4517 7783
rect 4477 7778 4517 7779
rect 4477 7774 4479 7778
rect 4483 7774 4489 7778
rect 4493 7774 4499 7778
rect 4503 7774 4509 7778
rect 4513 7774 4517 7778
rect 655 7467 659 7471
rect 663 7467 669 7471
rect 673 7467 679 7471
rect 683 7467 689 7471
rect 693 7467 695 7471
rect 655 7466 695 7467
rect 655 7462 659 7466
rect 663 7462 669 7466
rect 673 7462 679 7466
rect 683 7462 689 7466
rect 693 7462 695 7466
rect 655 7461 695 7462
rect 655 7457 659 7461
rect 663 7457 669 7461
rect 673 7457 679 7461
rect 683 7457 689 7461
rect 693 7457 695 7461
rect 655 7456 695 7457
rect 655 7452 659 7456
rect 663 7452 669 7456
rect 673 7452 679 7456
rect 683 7452 689 7456
rect 693 7452 695 7456
rect 655 7162 695 7452
rect 655 7158 659 7162
rect 663 7158 669 7162
rect 673 7158 679 7162
rect 683 7158 689 7162
rect 693 7158 695 7162
rect 655 7127 695 7158
rect 655 7123 659 7127
rect 663 7123 669 7127
rect 673 7123 679 7127
rect 683 7123 689 7127
rect 693 7123 695 7127
rect 655 7122 695 7123
rect 655 7118 659 7122
rect 663 7118 669 7122
rect 673 7118 679 7122
rect 683 7118 689 7122
rect 693 7118 695 7122
rect 655 7117 695 7118
rect 655 7113 659 7117
rect 663 7113 669 7117
rect 673 7113 679 7117
rect 683 7113 689 7117
rect 693 7113 695 7117
rect 655 7112 695 7113
rect 655 7108 659 7112
rect 663 7108 669 7112
rect 673 7108 679 7112
rect 683 7108 689 7112
rect 693 7108 695 7112
rect 655 6540 695 7108
rect 4477 7234 4517 7774
rect 4477 7230 4479 7234
rect 4483 7230 4489 7234
rect 4493 7230 4499 7234
rect 4503 7230 4509 7234
rect 4513 7230 4517 7234
rect 4477 7229 4517 7230
rect 4477 7225 4479 7229
rect 4483 7225 4489 7229
rect 4493 7225 4499 7229
rect 4503 7225 4509 7229
rect 4513 7225 4517 7229
rect 4477 7224 4517 7225
rect 4477 7220 4479 7224
rect 4483 7220 4489 7224
rect 4493 7220 4499 7224
rect 4503 7220 4509 7224
rect 4513 7220 4517 7224
rect 4477 7219 4517 7220
rect 4477 7215 4479 7219
rect 4483 7215 4489 7219
rect 4493 7215 4499 7219
rect 4503 7215 4509 7219
rect 4513 7215 4517 7219
rect 4477 7206 4517 7215
rect 4477 7202 4479 7206
rect 4483 7202 4489 7206
rect 4493 7202 4499 7206
rect 4503 7202 4509 7206
rect 4513 7202 4517 7206
rect 4477 7201 4517 7202
rect 4477 7197 4479 7201
rect 4483 7197 4489 7201
rect 4493 7197 4499 7201
rect 4503 7197 4509 7201
rect 4513 7197 4517 7201
rect 4477 7196 4517 7197
rect 4477 7192 4479 7196
rect 4483 7192 4489 7196
rect 4493 7192 4499 7196
rect 4503 7192 4509 7196
rect 4513 7192 4517 7196
rect 4477 7191 4517 7192
rect 4477 7187 4479 7191
rect 4483 7187 4489 7191
rect 4493 7187 4499 7191
rect 4503 7187 4509 7191
rect 4513 7187 4517 7191
rect 4477 7156 4517 7187
rect 4477 7152 4479 7156
rect 4483 7152 4489 7156
rect 4493 7152 4499 7156
rect 4503 7152 4509 7156
rect 4513 7152 4517 7156
rect 4477 6862 4517 7152
rect 4477 6858 4479 6862
rect 4483 6858 4489 6862
rect 4493 6858 4499 6862
rect 4503 6858 4509 6862
rect 4513 6858 4517 6862
rect 4477 6857 4517 6858
rect 4477 6853 4479 6857
rect 4483 6853 4489 6857
rect 4493 6853 4499 6857
rect 4503 6853 4509 6857
rect 4513 6853 4517 6857
rect 4477 6852 4517 6853
rect 4477 6848 4479 6852
rect 4483 6848 4489 6852
rect 4493 6848 4499 6852
rect 4503 6848 4509 6852
rect 4513 6848 4517 6852
rect 4477 6847 4517 6848
rect 4477 6843 4479 6847
rect 4483 6843 4489 6847
rect 4493 6843 4499 6847
rect 4503 6843 4509 6847
rect 4513 6843 4517 6847
rect 655 6536 659 6540
rect 663 6536 669 6540
rect 673 6536 679 6540
rect 683 6536 689 6540
rect 693 6536 695 6540
rect 655 6535 695 6536
rect 655 6531 659 6535
rect 663 6531 669 6535
rect 673 6531 679 6535
rect 683 6531 689 6535
rect 693 6531 695 6535
rect 655 6530 695 6531
rect 655 6526 659 6530
rect 663 6526 669 6530
rect 673 6526 679 6530
rect 683 6526 689 6530
rect 693 6526 695 6530
rect 655 6525 695 6526
rect 655 6521 659 6525
rect 663 6521 669 6525
rect 673 6521 679 6525
rect 683 6521 689 6525
rect 693 6521 695 6525
rect 655 6231 695 6521
rect 4477 6553 4517 6843
rect 4477 6549 4479 6553
rect 4483 6549 4489 6553
rect 4493 6549 4499 6553
rect 4503 6549 4509 6553
rect 4513 6549 4517 6553
rect 4477 6548 4517 6549
rect 4477 6544 4479 6548
rect 4483 6544 4489 6548
rect 4493 6544 4499 6548
rect 4503 6544 4509 6548
rect 4513 6544 4517 6548
rect 4477 6543 4517 6544
rect 4477 6539 4479 6543
rect 4483 6539 4489 6543
rect 4493 6539 4499 6543
rect 4503 6539 4509 6543
rect 4513 6539 4517 6543
rect 4477 6538 4517 6539
rect 4477 6534 4479 6538
rect 4483 6534 4489 6538
rect 4493 6534 4499 6538
rect 4503 6534 4509 6538
rect 4513 6534 4517 6538
rect 4477 6244 4517 6534
rect 4477 6240 4479 6244
rect 4483 6240 4489 6244
rect 4493 6240 4499 6244
rect 4503 6240 4509 6244
rect 4513 6240 4517 6244
rect 4477 6239 4517 6240
rect 4477 6235 4479 6239
rect 4483 6235 4489 6239
rect 4493 6235 4499 6239
rect 4503 6235 4509 6239
rect 4513 6235 4517 6239
rect 4477 6234 4517 6235
rect 655 6227 659 6231
rect 663 6227 669 6231
rect 673 6227 679 6231
rect 683 6227 689 6231
rect 693 6227 695 6231
rect 4477 6230 4479 6234
rect 4483 6230 4489 6234
rect 4493 6230 4499 6234
rect 4503 6230 4509 6234
rect 4513 6230 4517 6234
rect 4477 6229 4517 6230
rect 655 6226 695 6227
rect 655 6222 659 6226
rect 663 6222 669 6226
rect 673 6222 679 6226
rect 683 6222 689 6226
rect 693 6222 695 6226
rect 655 6221 695 6222
rect 655 6217 659 6221
rect 663 6217 669 6221
rect 673 6217 679 6221
rect 683 6217 689 6221
rect 693 6217 695 6221
rect 4477 6225 4479 6229
rect 4483 6225 4489 6229
rect 4493 6225 4499 6229
rect 4503 6225 4509 6229
rect 4513 6225 4517 6229
rect 655 6216 695 6217
rect 655 6212 659 6216
rect 663 6212 669 6216
rect 673 6212 679 6216
rect 683 6212 689 6216
rect 693 6212 695 6216
rect 655 6200 695 6212
rect 655 6196 659 6200
rect 663 6196 669 6200
rect 673 6196 679 6200
rect 683 6196 689 6200
rect 693 6196 695 6200
rect 655 6195 695 6196
rect 655 6191 659 6195
rect 663 6191 669 6195
rect 673 6191 679 6195
rect 683 6191 689 6195
rect 693 6191 695 6195
rect 655 6190 695 6191
rect 655 6186 659 6190
rect 663 6186 669 6190
rect 673 6186 679 6190
rect 683 6186 689 6190
rect 693 6186 695 6190
rect 655 6185 695 6186
rect 655 6181 659 6185
rect 663 6181 669 6185
rect 673 6181 679 6185
rect 683 6181 689 6185
rect 693 6181 695 6185
rect 655 5891 695 6181
rect 4477 5935 4517 6225
rect 4477 5931 4479 5935
rect 4483 5931 4489 5935
rect 4493 5931 4499 5935
rect 4503 5931 4509 5935
rect 4513 5931 4517 5935
rect 4477 5930 4517 5931
rect 4477 5926 4479 5930
rect 4483 5926 4489 5930
rect 4493 5926 4499 5930
rect 4503 5926 4509 5930
rect 4513 5926 4517 5930
rect 4477 5925 4517 5926
rect 4477 5921 4479 5925
rect 4483 5921 4489 5925
rect 4493 5921 4499 5925
rect 4503 5921 4509 5925
rect 4513 5921 4517 5925
rect 4477 5920 4517 5921
rect 4477 5916 4479 5920
rect 4483 5916 4489 5920
rect 4493 5916 4499 5920
rect 4503 5916 4509 5920
rect 4513 5916 4517 5920
rect 655 5887 659 5891
rect 663 5887 669 5891
rect 673 5887 679 5891
rect 683 5887 689 5891
rect 693 5887 695 5891
rect 655 5886 695 5887
rect 655 5882 659 5886
rect 663 5882 669 5886
rect 673 5882 679 5886
rect 683 5882 689 5886
rect 693 5882 695 5886
rect 655 5881 695 5882
rect 655 5877 659 5881
rect 663 5877 669 5881
rect 673 5877 679 5881
rect 683 5877 689 5881
rect 693 5877 695 5881
rect 655 5876 695 5877
rect 655 5872 659 5876
rect 663 5872 669 5876
rect 673 5872 679 5876
rect 683 5872 689 5876
rect 693 5872 695 5876
rect 655 5582 695 5872
rect 4477 5626 4517 5916
rect 4477 5622 4479 5626
rect 4483 5622 4489 5626
rect 4493 5622 4499 5626
rect 4503 5622 4509 5626
rect 4513 5622 4517 5626
rect 4477 5621 4517 5622
rect 4477 5617 4479 5621
rect 4483 5617 4489 5621
rect 4493 5617 4499 5621
rect 4503 5617 4509 5621
rect 4513 5617 4517 5621
rect 4477 5616 4517 5617
rect 4477 5612 4479 5616
rect 4483 5612 4489 5616
rect 4493 5612 4499 5616
rect 4503 5612 4509 5616
rect 4513 5612 4517 5616
rect 4477 5611 4517 5612
rect 4477 5607 4479 5611
rect 4483 5607 4489 5611
rect 4493 5607 4499 5611
rect 4503 5607 4509 5611
rect 4513 5607 4517 5611
rect 655 5578 659 5582
rect 663 5578 669 5582
rect 673 5578 679 5582
rect 683 5578 689 5582
rect 693 5578 695 5582
rect 655 5577 695 5578
rect 655 5573 659 5577
rect 663 5573 669 5577
rect 673 5573 679 5577
rect 683 5573 689 5577
rect 693 5573 695 5577
rect 655 5572 695 5573
rect 655 5568 659 5572
rect 663 5568 669 5572
rect 673 5568 679 5572
rect 683 5568 689 5572
rect 693 5568 695 5572
rect 655 5567 695 5568
rect 655 5563 659 5567
rect 663 5563 669 5567
rect 673 5563 679 5567
rect 683 5563 689 5567
rect 693 5563 695 5567
rect 655 5273 695 5563
rect 4477 5317 4517 5607
rect 4477 5313 4479 5317
rect 4483 5313 4489 5317
rect 4493 5313 4499 5317
rect 4503 5313 4509 5317
rect 4513 5313 4517 5317
rect 4477 5312 4517 5313
rect 4477 5308 4479 5312
rect 4483 5308 4489 5312
rect 4493 5308 4499 5312
rect 4503 5308 4509 5312
rect 4513 5308 4517 5312
rect 4477 5307 4517 5308
rect 4477 5303 4479 5307
rect 4483 5303 4489 5307
rect 4493 5303 4499 5307
rect 4503 5303 4509 5307
rect 4513 5303 4517 5307
rect 4477 5302 4517 5303
rect 4477 5298 4479 5302
rect 4483 5298 4489 5302
rect 4493 5298 4499 5302
rect 4503 5298 4509 5302
rect 4513 5298 4517 5302
rect 655 5269 659 5273
rect 663 5269 669 5273
rect 673 5269 679 5273
rect 683 5269 689 5273
rect 693 5269 695 5273
rect 655 5268 695 5269
rect 655 5264 659 5268
rect 663 5264 669 5268
rect 673 5264 679 5268
rect 683 5264 689 5268
rect 693 5264 695 5268
rect 655 5263 695 5264
rect 655 5259 659 5263
rect 663 5259 669 5263
rect 673 5259 679 5263
rect 683 5259 689 5263
rect 693 5259 695 5263
rect 655 5258 695 5259
rect 655 5254 659 5258
rect 663 5254 669 5258
rect 673 5254 679 5258
rect 683 5254 689 5258
rect 693 5254 695 5258
rect 655 4872 695 5254
rect 4477 5008 4517 5298
rect 4477 5004 4479 5008
rect 4483 5004 4489 5008
rect 4493 5004 4499 5008
rect 4503 5004 4509 5008
rect 4513 5004 4517 5008
rect 4477 5003 4517 5004
rect 4477 4999 4479 5003
rect 4483 4999 4489 5003
rect 4493 4999 4499 5003
rect 4503 4999 4509 5003
rect 4513 4999 4517 5003
rect 4477 4998 4517 4999
rect 4477 4994 4479 4998
rect 4483 4994 4489 4998
rect 4493 4994 4499 4998
rect 4503 4994 4509 4998
rect 4513 4994 4517 4998
rect 4477 4993 4517 4994
rect 4477 4989 4479 4993
rect 4483 4989 4489 4993
rect 4493 4989 4499 4993
rect 4503 4989 4509 4993
rect 4513 4989 4517 4993
rect 655 4868 659 4872
rect 663 4868 669 4872
rect 673 4868 679 4872
rect 683 4868 689 4872
rect 693 4868 695 4872
rect 655 4867 695 4868
rect 655 4863 659 4867
rect 663 4863 669 4867
rect 673 4863 679 4867
rect 683 4863 689 4867
rect 693 4863 695 4867
rect 655 4862 695 4863
rect 655 4858 659 4862
rect 663 4858 669 4862
rect 673 4858 679 4862
rect 683 4858 689 4862
rect 693 4858 695 4862
rect 655 4857 695 4858
rect 655 4853 659 4857
rect 663 4853 669 4857
rect 673 4853 679 4857
rect 683 4853 689 4857
rect 693 4853 695 4857
rect 655 4843 695 4853
rect 655 4839 659 4843
rect 663 4839 669 4843
rect 673 4839 679 4843
rect 683 4839 689 4843
rect 693 4839 695 4843
rect 655 4838 695 4839
rect 655 4834 659 4838
rect 663 4834 669 4838
rect 673 4834 679 4838
rect 683 4834 689 4838
rect 693 4834 695 4838
rect 655 4833 695 4834
rect 655 4829 659 4833
rect 663 4829 669 4833
rect 673 4829 679 4833
rect 683 4829 689 4833
rect 693 4829 695 4833
rect 655 4828 695 4829
rect 655 4824 659 4828
rect 663 4824 669 4828
rect 673 4824 679 4828
rect 683 4824 689 4828
rect 693 4824 695 4828
rect 655 4814 695 4824
rect 655 4810 659 4814
rect 663 4810 669 4814
rect 673 4810 679 4814
rect 683 4810 689 4814
rect 693 4810 695 4814
rect 655 4809 695 4810
rect 655 4805 659 4809
rect 663 4805 669 4809
rect 673 4805 679 4809
rect 683 4805 689 4809
rect 693 4805 695 4809
rect 655 4804 695 4805
rect 655 4800 659 4804
rect 663 4800 669 4804
rect 673 4800 679 4804
rect 683 4800 689 4804
rect 693 4800 695 4804
rect 655 4799 695 4800
rect 655 4795 659 4799
rect 663 4795 669 4799
rect 673 4795 679 4799
rect 683 4795 689 4799
rect 693 4795 695 4799
rect 655 4785 695 4795
rect 655 4781 659 4785
rect 663 4781 669 4785
rect 673 4781 679 4785
rect 683 4781 689 4785
rect 693 4781 695 4785
rect 655 4780 695 4781
rect 655 4776 659 4780
rect 663 4776 669 4780
rect 673 4776 679 4780
rect 683 4776 689 4780
rect 693 4776 695 4780
rect 655 4775 695 4776
rect 655 4771 659 4775
rect 663 4771 669 4775
rect 673 4771 679 4775
rect 683 4771 689 4775
rect 693 4771 695 4775
rect 655 4770 695 4771
rect 655 4766 659 4770
rect 663 4766 669 4770
rect 673 4766 679 4770
rect 683 4766 689 4770
rect 693 4766 695 4770
rect 655 4756 695 4766
rect 655 4752 659 4756
rect 663 4752 669 4756
rect 673 4752 679 4756
rect 683 4752 689 4756
rect 693 4752 695 4756
rect 655 4751 695 4752
rect 655 4747 659 4751
rect 663 4747 669 4751
rect 673 4747 679 4751
rect 683 4747 689 4751
rect 693 4747 695 4751
rect 655 4746 695 4747
rect 655 4742 659 4746
rect 663 4742 669 4746
rect 673 4742 679 4746
rect 683 4742 689 4746
rect 693 4742 695 4746
rect 655 4741 695 4742
rect 655 4737 659 4741
rect 663 4737 669 4741
rect 673 4737 679 4741
rect 683 4737 689 4741
rect 693 4737 695 4741
rect 655 4630 695 4737
rect 4477 4815 4517 4989
rect 4477 4811 4479 4815
rect 4483 4811 4489 4815
rect 4493 4811 4499 4815
rect 4503 4811 4509 4815
rect 4513 4811 4517 4815
rect 4477 4810 4517 4811
rect 4477 4806 4479 4810
rect 4483 4806 4489 4810
rect 4493 4806 4499 4810
rect 4503 4806 4509 4810
rect 4513 4806 4517 4810
rect 4477 4805 4517 4806
rect 4477 4801 4479 4805
rect 4483 4801 4489 4805
rect 4493 4801 4499 4805
rect 4503 4801 4509 4805
rect 4513 4801 4517 4805
rect 4477 4800 4517 4801
rect 4477 4796 4479 4800
rect 4483 4796 4489 4800
rect 4493 4796 4499 4800
rect 4503 4796 4509 4800
rect 4513 4796 4517 4800
rect 4477 4789 4517 4796
rect 4477 4785 4479 4789
rect 4483 4785 4489 4789
rect 4493 4785 4499 4789
rect 4503 4785 4509 4789
rect 4513 4785 4517 4789
rect 4477 4784 4517 4785
rect 4477 4780 4479 4784
rect 4483 4780 4489 4784
rect 4493 4780 4499 4784
rect 4503 4780 4509 4784
rect 4513 4780 4517 4784
rect 4477 4779 4517 4780
rect 4477 4775 4479 4779
rect 4483 4775 4489 4779
rect 4493 4775 4499 4779
rect 4503 4775 4509 4779
rect 4513 4775 4517 4779
rect 4477 4774 4517 4775
rect 4477 4770 4479 4774
rect 4483 4770 4489 4774
rect 4493 4770 4499 4774
rect 4503 4770 4509 4774
rect 4513 4770 4517 4774
rect 4477 4763 4517 4770
rect 4477 4759 4479 4763
rect 4483 4759 4489 4763
rect 4493 4759 4499 4763
rect 4503 4759 4509 4763
rect 4513 4759 4517 4763
rect 4477 4758 4517 4759
rect 4477 4754 4479 4758
rect 4483 4754 4489 4758
rect 4493 4754 4499 4758
rect 4503 4754 4509 4758
rect 4513 4754 4517 4758
rect 4477 4753 4517 4754
rect 4477 4749 4479 4753
rect 4483 4749 4489 4753
rect 4493 4749 4499 4753
rect 4503 4749 4509 4753
rect 4513 4749 4517 4753
rect 4477 4748 4517 4749
rect 4477 4744 4479 4748
rect 4483 4744 4489 4748
rect 4493 4744 4499 4748
rect 4503 4744 4509 4748
rect 4513 4744 4517 4748
rect 4477 4737 4517 4744
rect 4477 4733 4479 4737
rect 4483 4733 4489 4737
rect 4493 4733 4499 4737
rect 4503 4733 4509 4737
rect 4513 4733 4517 4737
rect 4477 4732 4517 4733
rect 4477 4728 4479 4732
rect 4483 4728 4489 4732
rect 4493 4728 4499 4732
rect 4503 4728 4509 4732
rect 4513 4728 4517 4732
rect 4477 4727 4517 4728
rect 4477 4723 4479 4727
rect 4483 4723 4489 4727
rect 4493 4723 4499 4727
rect 4503 4723 4509 4727
rect 4513 4723 4517 4727
rect 4477 4722 4517 4723
rect 4477 4718 4479 4722
rect 4483 4718 4489 4722
rect 4493 4718 4499 4722
rect 4503 4718 4509 4722
rect 4513 4718 4517 4722
rect 4477 4711 4517 4718
rect 4477 4707 4479 4711
rect 4483 4707 4489 4711
rect 4493 4707 4499 4711
rect 4503 4707 4509 4711
rect 4513 4707 4517 4711
rect 4477 4706 4517 4707
rect 4477 4702 4479 4706
rect 4483 4702 4489 4706
rect 4493 4702 4499 4706
rect 4503 4702 4509 4706
rect 4513 4702 4517 4706
rect 4477 4701 4517 4702
rect 4477 4697 4479 4701
rect 4483 4697 4489 4701
rect 4493 4697 4499 4701
rect 4503 4697 4509 4701
rect 4513 4697 4517 4701
rect 4477 4696 4517 4697
rect 4477 4692 4479 4696
rect 4483 4692 4489 4696
rect 4493 4692 4499 4696
rect 4503 4692 4509 4696
rect 4513 4692 4517 4696
rect 4477 4630 4517 4692
rect 655 4628 4517 4630
rect 655 4624 757 4628
rect 761 4624 762 4628
rect 766 4624 767 4628
rect 771 4624 772 4628
rect 776 4624 783 4628
rect 787 4624 788 4628
rect 792 4624 793 4628
rect 797 4624 798 4628
rect 802 4624 809 4628
rect 813 4624 814 4628
rect 818 4624 819 4628
rect 823 4624 824 4628
rect 828 4624 835 4628
rect 839 4624 840 4628
rect 844 4624 845 4628
rect 849 4624 850 4628
rect 854 4624 861 4628
rect 865 4624 866 4628
rect 870 4624 871 4628
rect 875 4624 876 4628
rect 880 4624 1053 4628
rect 1057 4624 1058 4628
rect 1062 4624 1063 4628
rect 1067 4624 1068 4628
rect 1072 4624 1362 4628
rect 1366 4624 1367 4628
rect 1371 4624 1372 4628
rect 1376 4624 1377 4628
rect 1381 4624 1671 4628
rect 1675 4624 1676 4628
rect 1680 4624 1681 4628
rect 1685 4624 1686 4628
rect 1690 4624 1980 4628
rect 1984 4624 1985 4628
rect 1989 4624 1990 4628
rect 1994 4624 1995 4628
rect 1999 4624 2289 4628
rect 2293 4624 2294 4628
rect 2298 4624 2299 4628
rect 2303 4624 2304 4628
rect 2308 4624 2598 4628
rect 2602 4624 2603 4628
rect 2607 4624 2608 4628
rect 2612 4624 2613 4628
rect 2617 4624 2907 4628
rect 2911 4624 2912 4628
rect 2916 4624 2917 4628
rect 2921 4624 2922 4628
rect 2926 4624 3216 4628
rect 3220 4624 3221 4628
rect 3225 4624 3226 4628
rect 3230 4624 3231 4628
rect 3235 4624 3525 4628
rect 3529 4624 3530 4628
rect 3534 4624 3535 4628
rect 3539 4624 3540 4628
rect 3544 4624 3834 4628
rect 3838 4624 3839 4628
rect 3843 4624 3844 4628
rect 3848 4624 3849 4628
rect 3853 4624 4235 4628
rect 4239 4624 4240 4628
rect 4244 4624 4245 4628
rect 4249 4624 4250 4628
rect 4254 4624 4264 4628
rect 4268 4624 4269 4628
rect 4273 4624 4274 4628
rect 4278 4624 4279 4628
rect 4283 4624 4293 4628
rect 4297 4624 4298 4628
rect 4302 4624 4303 4628
rect 4307 4624 4308 4628
rect 4312 4624 4322 4628
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4336 4624 4337 4628
rect 4341 4624 4351 4628
rect 4355 4624 4356 4628
rect 4360 4624 4361 4628
rect 4365 4624 4366 4628
rect 4370 4624 4517 4628
rect 655 4618 4517 4624
rect 655 4614 757 4618
rect 761 4614 762 4618
rect 766 4614 767 4618
rect 771 4614 772 4618
rect 776 4614 783 4618
rect 787 4614 788 4618
rect 792 4614 793 4618
rect 797 4614 798 4618
rect 802 4614 809 4618
rect 813 4614 814 4618
rect 818 4614 819 4618
rect 823 4614 824 4618
rect 828 4614 835 4618
rect 839 4614 840 4618
rect 844 4614 845 4618
rect 849 4614 850 4618
rect 854 4614 861 4618
rect 865 4614 866 4618
rect 870 4614 871 4618
rect 875 4614 876 4618
rect 880 4614 1053 4618
rect 1057 4614 1058 4618
rect 1062 4614 1063 4618
rect 1067 4614 1068 4618
rect 1072 4614 1362 4618
rect 1366 4614 1367 4618
rect 1371 4614 1372 4618
rect 1376 4614 1377 4618
rect 1381 4614 1671 4618
rect 1675 4614 1676 4618
rect 1680 4614 1681 4618
rect 1685 4614 1686 4618
rect 1690 4614 1980 4618
rect 1984 4614 1985 4618
rect 1989 4614 1990 4618
rect 1994 4614 1995 4618
rect 1999 4614 2289 4618
rect 2293 4614 2294 4618
rect 2298 4614 2299 4618
rect 2303 4614 2304 4618
rect 2308 4614 2598 4618
rect 2602 4614 2603 4618
rect 2607 4614 2608 4618
rect 2612 4614 2613 4618
rect 2617 4614 2907 4618
rect 2911 4614 2912 4618
rect 2916 4614 2917 4618
rect 2921 4614 2922 4618
rect 2926 4614 3216 4618
rect 3220 4614 3221 4618
rect 3225 4614 3226 4618
rect 3230 4614 3231 4618
rect 3235 4614 3525 4618
rect 3529 4614 3530 4618
rect 3534 4614 3535 4618
rect 3539 4614 3540 4618
rect 3544 4614 3834 4618
rect 3838 4614 3839 4618
rect 3843 4614 3844 4618
rect 3848 4614 3849 4618
rect 3853 4614 4235 4618
rect 4239 4614 4240 4618
rect 4244 4614 4245 4618
rect 4249 4614 4250 4618
rect 4254 4614 4264 4618
rect 4268 4614 4269 4618
rect 4273 4614 4274 4618
rect 4278 4614 4279 4618
rect 4283 4614 4293 4618
rect 4297 4614 4298 4618
rect 4302 4614 4303 4618
rect 4307 4614 4308 4618
rect 4312 4614 4322 4618
rect 4326 4614 4327 4618
rect 4331 4614 4332 4618
rect 4336 4614 4337 4618
rect 4341 4614 4351 4618
rect 4355 4614 4356 4618
rect 4360 4614 4361 4618
rect 4365 4614 4366 4618
rect 4370 4614 4517 4618
rect 655 4608 4517 4614
rect 655 4604 757 4608
rect 761 4604 762 4608
rect 766 4604 767 4608
rect 771 4604 772 4608
rect 776 4604 783 4608
rect 787 4604 788 4608
rect 792 4604 793 4608
rect 797 4604 798 4608
rect 802 4604 809 4608
rect 813 4604 814 4608
rect 818 4604 819 4608
rect 823 4604 824 4608
rect 828 4604 835 4608
rect 839 4604 840 4608
rect 844 4604 845 4608
rect 849 4604 850 4608
rect 854 4604 861 4608
rect 865 4604 866 4608
rect 870 4604 871 4608
rect 875 4604 876 4608
rect 880 4604 1053 4608
rect 1057 4604 1058 4608
rect 1062 4604 1063 4608
rect 1067 4604 1068 4608
rect 1072 4604 1362 4608
rect 1366 4604 1367 4608
rect 1371 4604 1372 4608
rect 1376 4604 1377 4608
rect 1381 4604 1671 4608
rect 1675 4604 1676 4608
rect 1680 4604 1681 4608
rect 1685 4604 1686 4608
rect 1690 4604 1980 4608
rect 1984 4604 1985 4608
rect 1989 4604 1990 4608
rect 1994 4604 1995 4608
rect 1999 4604 2289 4608
rect 2293 4604 2294 4608
rect 2298 4604 2299 4608
rect 2303 4604 2304 4608
rect 2308 4604 2598 4608
rect 2602 4604 2603 4608
rect 2607 4604 2608 4608
rect 2612 4604 2613 4608
rect 2617 4604 2907 4608
rect 2911 4604 2912 4608
rect 2916 4604 2917 4608
rect 2921 4604 2922 4608
rect 2926 4604 3216 4608
rect 3220 4604 3221 4608
rect 3225 4604 3226 4608
rect 3230 4604 3231 4608
rect 3235 4604 3525 4608
rect 3529 4604 3530 4608
rect 3534 4604 3535 4608
rect 3539 4604 3540 4608
rect 3544 4604 3834 4608
rect 3838 4604 3839 4608
rect 3843 4604 3844 4608
rect 3848 4604 3849 4608
rect 3853 4604 4235 4608
rect 4239 4604 4240 4608
rect 4244 4604 4245 4608
rect 4249 4604 4250 4608
rect 4254 4604 4264 4608
rect 4268 4604 4269 4608
rect 4273 4604 4274 4608
rect 4278 4604 4279 4608
rect 4283 4604 4293 4608
rect 4297 4604 4298 4608
rect 4302 4604 4303 4608
rect 4307 4604 4308 4608
rect 4312 4604 4322 4608
rect 4326 4604 4327 4608
rect 4331 4604 4332 4608
rect 4336 4604 4337 4608
rect 4341 4604 4351 4608
rect 4355 4604 4356 4608
rect 4360 4604 4361 4608
rect 4365 4604 4366 4608
rect 4370 4604 4517 4608
rect 655 4598 4517 4604
rect 655 4594 757 4598
rect 761 4594 762 4598
rect 766 4594 767 4598
rect 771 4594 772 4598
rect 776 4594 783 4598
rect 787 4594 788 4598
rect 792 4594 793 4598
rect 797 4594 798 4598
rect 802 4594 809 4598
rect 813 4594 814 4598
rect 818 4594 819 4598
rect 823 4594 824 4598
rect 828 4594 835 4598
rect 839 4594 840 4598
rect 844 4594 845 4598
rect 849 4594 850 4598
rect 854 4594 861 4598
rect 865 4594 866 4598
rect 870 4594 871 4598
rect 875 4594 876 4598
rect 880 4594 1053 4598
rect 1057 4594 1058 4598
rect 1062 4594 1063 4598
rect 1067 4594 1068 4598
rect 1072 4594 1362 4598
rect 1366 4594 1367 4598
rect 1371 4594 1372 4598
rect 1376 4594 1377 4598
rect 1381 4594 1671 4598
rect 1675 4594 1676 4598
rect 1680 4594 1681 4598
rect 1685 4594 1686 4598
rect 1690 4594 1980 4598
rect 1984 4594 1985 4598
rect 1989 4594 1990 4598
rect 1994 4594 1995 4598
rect 1999 4594 2289 4598
rect 2293 4594 2294 4598
rect 2298 4594 2299 4598
rect 2303 4594 2304 4598
rect 2308 4594 2598 4598
rect 2602 4594 2603 4598
rect 2607 4594 2608 4598
rect 2612 4594 2613 4598
rect 2617 4594 2907 4598
rect 2911 4594 2912 4598
rect 2916 4594 2917 4598
rect 2921 4594 2922 4598
rect 2926 4594 3216 4598
rect 3220 4594 3221 4598
rect 3225 4594 3226 4598
rect 3230 4594 3231 4598
rect 3235 4594 3525 4598
rect 3529 4594 3530 4598
rect 3534 4594 3535 4598
rect 3539 4594 3540 4598
rect 3544 4594 3834 4598
rect 3838 4594 3839 4598
rect 3843 4594 3844 4598
rect 3848 4594 3849 4598
rect 3853 4594 4235 4598
rect 4239 4594 4240 4598
rect 4244 4594 4245 4598
rect 4249 4594 4250 4598
rect 4254 4594 4264 4598
rect 4268 4594 4269 4598
rect 4273 4594 4274 4598
rect 4278 4594 4279 4598
rect 4283 4594 4293 4598
rect 4297 4594 4298 4598
rect 4302 4594 4303 4598
rect 4307 4594 4308 4598
rect 4312 4594 4322 4598
rect 4326 4594 4327 4598
rect 4331 4594 4332 4598
rect 4336 4594 4337 4598
rect 4341 4594 4351 4598
rect 4355 4594 4356 4598
rect 4360 4594 4361 4598
rect 4365 4594 4366 4598
rect 4370 4594 4517 4598
rect 655 4590 4517 4594
rect 4643 7477 4760 7479
rect 4643 7473 4645 7477
rect 4649 7473 4652 7477
rect 4656 7473 4657 7477
rect 4661 7473 4662 7477
rect 4666 7473 4667 7477
rect 4671 7473 4672 7477
rect 4676 7473 4677 7477
rect 4681 7473 4682 7477
rect 4686 7473 4687 7477
rect 4691 7473 4692 7477
rect 4696 7473 4697 7477
rect 4701 7473 4702 7477
rect 4706 7473 4707 7477
rect 4711 7473 4712 7477
rect 4716 7473 4717 7477
rect 4721 7473 4722 7477
rect 4726 7473 4727 7477
rect 4731 7473 4732 7477
rect 4736 7473 4737 7477
rect 4741 7473 4742 7477
rect 4746 7473 4747 7477
rect 4751 7473 4754 7477
rect 4758 7473 4760 7477
rect 4643 7471 4760 7473
rect 4643 7470 4651 7471
rect 4643 7466 4645 7470
rect 4649 7466 4651 7470
rect 4643 7465 4651 7466
rect 4752 7470 4760 7471
rect 4752 7466 4754 7470
rect 4758 7466 4760 7470
rect 4752 7465 4760 7466
rect 4643 7461 4645 7465
rect 4649 7461 4651 7465
rect 4643 7460 4651 7461
rect 4643 7456 4645 7460
rect 4649 7456 4651 7460
rect 4643 7455 4651 7456
rect 4643 7451 4645 7455
rect 4649 7451 4651 7455
rect 4643 7450 4651 7451
rect 4643 7446 4645 7450
rect 4649 7446 4651 7450
rect 4643 7445 4651 7446
rect 4643 7441 4645 7445
rect 4649 7441 4651 7445
rect 4643 7440 4651 7441
rect 4643 7436 4645 7440
rect 4649 7436 4651 7440
rect 4643 7435 4651 7436
rect 4643 7431 4645 7435
rect 4649 7431 4651 7435
rect 4643 7430 4651 7431
rect 4643 7426 4645 7430
rect 4649 7426 4651 7430
rect 4643 7425 4651 7426
rect 4643 7421 4645 7425
rect 4649 7421 4651 7425
rect 4752 7461 4754 7465
rect 4758 7461 4760 7465
rect 4752 7460 4760 7461
rect 4752 7456 4754 7460
rect 4758 7456 4760 7460
rect 4752 7455 4760 7456
rect 4752 7451 4754 7455
rect 4758 7451 4760 7455
rect 4752 7450 4760 7451
rect 4752 7446 4754 7450
rect 4758 7446 4760 7450
rect 4752 7445 4760 7446
rect 4752 7441 4754 7445
rect 4758 7441 4760 7445
rect 4752 7440 4760 7441
rect 4752 7436 4754 7440
rect 4758 7436 4760 7440
rect 4752 7435 4760 7436
rect 4752 7431 4754 7435
rect 4758 7431 4760 7435
rect 4752 7430 4760 7431
rect 4752 7426 4754 7430
rect 4758 7426 4760 7430
rect 4752 7425 4760 7426
rect 4752 7421 4754 7425
rect 4758 7421 4760 7425
rect 4643 7420 4651 7421
rect 4643 7416 4645 7420
rect 4649 7416 4651 7420
rect 4643 7415 4651 7416
rect 4752 7420 4760 7421
rect 4752 7416 4754 7420
rect 4758 7416 4760 7420
rect 4752 7415 4760 7416
rect 4643 7413 4760 7415
rect 4643 7409 4645 7413
rect 4649 7409 4652 7413
rect 4656 7409 4657 7413
rect 4661 7409 4662 7413
rect 4666 7409 4667 7413
rect 4671 7409 4672 7413
rect 4676 7409 4677 7413
rect 4681 7409 4682 7413
rect 4686 7409 4687 7413
rect 4691 7409 4692 7413
rect 4696 7409 4697 7413
rect 4701 7409 4702 7413
rect 4706 7409 4707 7413
rect 4711 7409 4712 7413
rect 4716 7409 4717 7413
rect 4721 7409 4722 7413
rect 4726 7409 4727 7413
rect 4731 7409 4732 7413
rect 4736 7409 4737 7413
rect 4741 7409 4742 7413
rect 4746 7409 4747 7413
rect 4751 7409 4754 7413
rect 4758 7409 4760 7413
rect 4643 7407 4760 7409
rect 4631 7330 4772 7331
rect 4631 7326 4632 7330
rect 4636 7326 4637 7330
rect 4641 7326 4642 7330
rect 4646 7326 4647 7330
rect 4651 7326 4652 7330
rect 4656 7326 4657 7330
rect 4661 7326 4662 7330
rect 4666 7326 4667 7330
rect 4671 7326 4672 7330
rect 4676 7326 4677 7330
rect 4681 7326 4682 7330
rect 4686 7326 4687 7330
rect 4691 7326 4692 7330
rect 4696 7326 4697 7330
rect 4701 7326 4702 7330
rect 4706 7326 4707 7330
rect 4711 7326 4712 7330
rect 4716 7326 4717 7330
rect 4721 7326 4722 7330
rect 4726 7326 4727 7330
rect 4731 7326 4732 7330
rect 4736 7326 4737 7330
rect 4741 7326 4742 7330
rect 4746 7326 4747 7330
rect 4751 7326 4752 7330
rect 4756 7326 4757 7330
rect 4761 7326 4762 7330
rect 4766 7326 4767 7330
rect 4771 7326 4772 7330
rect 4631 7325 4772 7326
rect 4631 7321 4632 7325
rect 4636 7321 4637 7325
rect 4631 7320 4637 7321
rect 4631 7316 4632 7320
rect 4636 7316 4637 7320
rect 4766 7321 4767 7325
rect 4771 7321 4772 7325
rect 4766 7320 4772 7321
rect 4631 7315 4637 7316
rect 4631 7311 4632 7315
rect 4636 7311 4637 7315
rect 4631 7310 4637 7311
rect 4631 7306 4632 7310
rect 4636 7306 4637 7310
rect 4631 7305 4637 7306
rect 4631 7301 4632 7305
rect 4636 7301 4637 7305
rect 4631 7300 4637 7301
rect 4631 7296 4632 7300
rect 4636 7296 4637 7300
rect 4631 7295 4637 7296
rect 4631 7291 4632 7295
rect 4636 7291 4637 7295
rect 4631 7290 4637 7291
rect 4631 7286 4632 7290
rect 4636 7286 4637 7290
rect 4631 7285 4637 7286
rect 4631 7281 4632 7285
rect 4636 7281 4637 7285
rect 4631 7280 4637 7281
rect 4631 7276 4632 7280
rect 4636 7276 4637 7280
rect 4631 7275 4637 7276
rect 4631 7271 4632 7275
rect 4636 7271 4637 7275
rect 4631 7270 4637 7271
rect 4631 7266 4632 7270
rect 4636 7266 4637 7270
rect 4631 7265 4637 7266
rect 4631 7261 4632 7265
rect 4636 7261 4637 7265
rect 4631 7260 4637 7261
rect 4631 7256 4632 7260
rect 4636 7256 4637 7260
rect 4631 7255 4637 7256
rect 4631 7251 4632 7255
rect 4636 7251 4637 7255
rect 4631 7250 4637 7251
rect 4631 7246 4632 7250
rect 4636 7246 4637 7250
rect 4766 7316 4767 7320
rect 4771 7316 4772 7320
rect 4766 7315 4772 7316
rect 4766 7311 4767 7315
rect 4771 7311 4772 7315
rect 4766 7310 4772 7311
rect 4766 7306 4767 7310
rect 4771 7306 4772 7310
rect 4766 7305 4772 7306
rect 4766 7301 4767 7305
rect 4771 7301 4772 7305
rect 4766 7300 4772 7301
rect 4766 7296 4767 7300
rect 4771 7296 4772 7300
rect 4766 7295 4772 7296
rect 4766 7291 4767 7295
rect 4771 7291 4772 7295
rect 4766 7290 4772 7291
rect 4766 7286 4767 7290
rect 4771 7286 4772 7290
rect 4766 7285 4772 7286
rect 4766 7281 4767 7285
rect 4771 7281 4772 7285
rect 4766 7280 4772 7281
rect 4766 7276 4767 7280
rect 4771 7276 4772 7280
rect 4766 7275 4772 7276
rect 4766 7271 4767 7275
rect 4771 7271 4772 7275
rect 4766 7270 4772 7271
rect 4766 7266 4767 7270
rect 4771 7266 4772 7270
rect 4766 7265 4772 7266
rect 4766 7261 4767 7265
rect 4771 7261 4772 7265
rect 4766 7260 4772 7261
rect 4766 7256 4767 7260
rect 4771 7256 4772 7260
rect 4766 7255 4772 7256
rect 4766 7251 4767 7255
rect 4771 7251 4772 7255
rect 4766 7250 4772 7251
rect 4631 7245 4637 7246
rect 4631 7241 4632 7245
rect 4636 7241 4637 7245
rect 4766 7246 4767 7250
rect 4771 7246 4772 7250
rect 4766 7245 4772 7246
rect 4766 7241 4767 7245
rect 4771 7241 4772 7245
rect 4631 7240 4772 7241
rect 4631 7236 4632 7240
rect 4636 7236 4637 7240
rect 4641 7236 4642 7240
rect 4646 7236 4647 7240
rect 4651 7236 4652 7240
rect 4656 7236 4657 7240
rect 4661 7236 4662 7240
rect 4666 7236 4667 7240
rect 4671 7236 4672 7240
rect 4676 7236 4677 7240
rect 4681 7236 4682 7240
rect 4686 7236 4687 7240
rect 4691 7236 4692 7240
rect 4696 7236 4697 7240
rect 4701 7236 4702 7240
rect 4706 7236 4707 7240
rect 4711 7236 4712 7240
rect 4716 7236 4717 7240
rect 4721 7236 4722 7240
rect 4726 7236 4727 7240
rect 4731 7236 4732 7240
rect 4736 7236 4737 7240
rect 4741 7236 4742 7240
rect 4746 7236 4747 7240
rect 4751 7236 4752 7240
rect 4756 7236 4757 7240
rect 4761 7236 4762 7240
rect 4766 7236 4767 7240
rect 4771 7236 4772 7240
rect 4631 7235 4772 7236
rect 1073 4475 1169 4476
rect 1073 4471 1074 4475
rect 1078 4471 1079 4475
rect 1083 4471 1084 4475
rect 1088 4471 1089 4475
rect 1093 4471 1094 4475
rect 1098 4471 1099 4475
rect 1103 4471 1104 4475
rect 1108 4471 1109 4475
rect 1113 4471 1114 4475
rect 1118 4471 1119 4475
rect 1123 4471 1124 4475
rect 1128 4471 1129 4475
rect 1133 4471 1134 4475
rect 1138 4471 1139 4475
rect 1143 4471 1144 4475
rect 1148 4471 1149 4475
rect 1153 4471 1154 4475
rect 1158 4471 1159 4475
rect 1163 4471 1164 4475
rect 1168 4471 1169 4475
rect 1073 4470 1169 4471
rect 1073 4466 1074 4470
rect 1078 4466 1079 4470
rect 1073 4465 1079 4466
rect 1073 4461 1074 4465
rect 1078 4461 1079 4465
rect 1163 4466 1164 4470
rect 1168 4466 1169 4470
rect 1163 4465 1169 4466
rect 1073 4460 1079 4461
rect 1073 4456 1074 4460
rect 1078 4456 1079 4460
rect 1073 4455 1079 4456
rect 1073 4451 1074 4455
rect 1078 4451 1079 4455
rect 1073 4450 1079 4451
rect 1073 4446 1074 4450
rect 1078 4446 1079 4450
rect 1073 4445 1079 4446
rect 1073 4441 1074 4445
rect 1078 4441 1079 4445
rect 1073 4440 1079 4441
rect 1073 4436 1074 4440
rect 1078 4436 1079 4440
rect 1073 4435 1079 4436
rect 1073 4431 1074 4435
rect 1078 4431 1079 4435
rect 1073 4430 1079 4431
rect 1073 4426 1074 4430
rect 1078 4426 1079 4430
rect 1073 4425 1079 4426
rect 1073 4421 1074 4425
rect 1078 4421 1079 4425
rect 1073 4420 1079 4421
rect 1073 4416 1074 4420
rect 1078 4416 1079 4420
rect 1073 4415 1079 4416
rect 1073 4411 1074 4415
rect 1078 4411 1079 4415
rect 1073 4410 1079 4411
rect 1073 4406 1074 4410
rect 1078 4406 1079 4410
rect 1073 4405 1079 4406
rect 1073 4401 1074 4405
rect 1078 4401 1079 4405
rect 1073 4400 1079 4401
rect 1073 4396 1074 4400
rect 1078 4396 1079 4400
rect 1073 4395 1079 4396
rect 1073 4391 1074 4395
rect 1078 4391 1079 4395
rect 1073 4390 1079 4391
rect 1073 4386 1074 4390
rect 1078 4386 1079 4390
rect 1073 4385 1079 4386
rect 1073 4381 1074 4385
rect 1078 4381 1079 4385
rect 1073 4380 1079 4381
rect 1073 4376 1074 4380
rect 1078 4376 1079 4380
rect 1073 4375 1079 4376
rect 1073 4371 1074 4375
rect 1078 4371 1079 4375
rect 1073 4370 1079 4371
rect 1073 4366 1074 4370
rect 1078 4366 1079 4370
rect 1073 4365 1079 4366
rect 1073 4361 1074 4365
rect 1078 4361 1079 4365
rect 1073 4360 1079 4361
rect 1073 4356 1074 4360
rect 1078 4356 1079 4360
rect 1073 4355 1079 4356
rect 1073 4351 1074 4355
rect 1078 4351 1079 4355
rect 1073 4350 1079 4351
rect 1073 4346 1074 4350
rect 1078 4346 1079 4350
rect 1163 4461 1164 4465
rect 1168 4461 1169 4465
rect 1163 4460 1169 4461
rect 1163 4456 1164 4460
rect 1168 4456 1169 4460
rect 1163 4455 1169 4456
rect 1163 4451 1164 4455
rect 1168 4451 1169 4455
rect 1163 4450 1169 4451
rect 1163 4446 1164 4450
rect 1168 4446 1169 4450
rect 1163 4445 1169 4446
rect 1163 4441 1164 4445
rect 1168 4441 1169 4445
rect 1163 4440 1169 4441
rect 1163 4436 1164 4440
rect 1168 4436 1169 4440
rect 1163 4435 1169 4436
rect 1163 4431 1164 4435
rect 1168 4431 1169 4435
rect 1163 4430 1169 4431
rect 1163 4426 1164 4430
rect 1168 4426 1169 4430
rect 1163 4425 1169 4426
rect 1163 4421 1164 4425
rect 1168 4421 1169 4425
rect 1163 4420 1169 4421
rect 1163 4416 1164 4420
rect 1168 4416 1169 4420
rect 1163 4415 1169 4416
rect 1163 4411 1164 4415
rect 1168 4411 1169 4415
rect 1163 4410 1169 4411
rect 1163 4406 1164 4410
rect 1168 4406 1169 4410
rect 1163 4405 1169 4406
rect 1163 4401 1164 4405
rect 1168 4401 1169 4405
rect 1163 4400 1169 4401
rect 1163 4396 1164 4400
rect 1168 4396 1169 4400
rect 1163 4395 1169 4396
rect 1163 4391 1164 4395
rect 1168 4391 1169 4395
rect 1163 4390 1169 4391
rect 1163 4386 1164 4390
rect 1168 4386 1169 4390
rect 1163 4385 1169 4386
rect 1163 4381 1164 4385
rect 1168 4381 1169 4385
rect 1163 4380 1169 4381
rect 1163 4376 1164 4380
rect 1168 4376 1169 4380
rect 1163 4375 1169 4376
rect 1163 4371 1164 4375
rect 1168 4371 1169 4375
rect 1163 4370 1169 4371
rect 1163 4366 1164 4370
rect 1168 4366 1169 4370
rect 1163 4365 1169 4366
rect 1163 4361 1164 4365
rect 1168 4361 1169 4365
rect 1163 4360 1169 4361
rect 1163 4356 1164 4360
rect 1168 4356 1169 4360
rect 1163 4355 1169 4356
rect 1163 4351 1164 4355
rect 1168 4351 1169 4355
rect 1163 4350 1169 4351
rect 1073 4345 1079 4346
rect 1073 4341 1074 4345
rect 1078 4341 1079 4345
rect 1163 4346 1164 4350
rect 1168 4346 1169 4350
rect 1163 4345 1169 4346
rect 1163 4341 1164 4345
rect 1168 4341 1169 4345
rect 1073 4340 1169 4341
rect 1073 4336 1074 4340
rect 1078 4336 1079 4340
rect 1083 4336 1084 4340
rect 1088 4336 1089 4340
rect 1093 4336 1094 4340
rect 1098 4336 1099 4340
rect 1103 4336 1104 4340
rect 1108 4336 1109 4340
rect 1113 4336 1114 4340
rect 1118 4336 1119 4340
rect 1123 4336 1124 4340
rect 1128 4336 1129 4340
rect 1133 4336 1134 4340
rect 1138 4336 1139 4340
rect 1143 4336 1144 4340
rect 1148 4336 1149 4340
rect 1153 4336 1154 4340
rect 1158 4336 1159 4340
rect 1163 4336 1164 4340
rect 1168 4336 1169 4340
rect 1073 4335 1169 4336
rect 1245 4462 1317 4464
rect 1245 4458 1247 4462
rect 1251 4458 1254 4462
rect 1258 4458 1259 4462
rect 1263 4458 1264 4462
rect 1268 4458 1269 4462
rect 1273 4458 1274 4462
rect 1278 4458 1279 4462
rect 1283 4458 1284 4462
rect 1288 4458 1289 4462
rect 1293 4458 1294 4462
rect 1298 4458 1299 4462
rect 1303 4458 1304 4462
rect 1308 4458 1311 4462
rect 1315 4458 1317 4462
rect 1245 4456 1317 4458
rect 1245 4455 1253 4456
rect 1245 4451 1247 4455
rect 1251 4451 1253 4455
rect 1245 4450 1253 4451
rect 1309 4455 1317 4456
rect 1309 4451 1311 4455
rect 1315 4451 1317 4455
rect 1309 4450 1317 4451
rect 1245 4446 1247 4450
rect 1251 4446 1253 4450
rect 1245 4445 1253 4446
rect 1245 4441 1247 4445
rect 1251 4441 1253 4445
rect 1245 4440 1253 4441
rect 1245 4436 1247 4440
rect 1251 4436 1253 4440
rect 1245 4435 1253 4436
rect 1245 4431 1247 4435
rect 1251 4431 1253 4435
rect 1245 4430 1253 4431
rect 1245 4426 1247 4430
rect 1251 4426 1253 4430
rect 1245 4425 1253 4426
rect 1245 4421 1247 4425
rect 1251 4421 1253 4425
rect 1245 4420 1253 4421
rect 1245 4416 1247 4420
rect 1251 4416 1253 4420
rect 1245 4415 1253 4416
rect 1245 4411 1247 4415
rect 1251 4411 1253 4415
rect 1245 4410 1253 4411
rect 1245 4406 1247 4410
rect 1251 4406 1253 4410
rect 1245 4405 1253 4406
rect 1245 4401 1247 4405
rect 1251 4401 1253 4405
rect 1245 4400 1253 4401
rect 1245 4396 1247 4400
rect 1251 4396 1253 4400
rect 1245 4395 1253 4396
rect 1245 4391 1247 4395
rect 1251 4391 1253 4395
rect 1245 4390 1253 4391
rect 1245 4386 1247 4390
rect 1251 4386 1253 4390
rect 1245 4385 1253 4386
rect 1245 4381 1247 4385
rect 1251 4381 1253 4385
rect 1245 4380 1253 4381
rect 1245 4376 1247 4380
rect 1251 4376 1253 4380
rect 1245 4375 1253 4376
rect 1245 4371 1247 4375
rect 1251 4371 1253 4375
rect 1245 4370 1253 4371
rect 1245 4366 1247 4370
rect 1251 4366 1253 4370
rect 1245 4365 1253 4366
rect 1245 4361 1247 4365
rect 1251 4361 1253 4365
rect 1309 4446 1311 4450
rect 1315 4446 1317 4450
rect 1309 4445 1317 4446
rect 1309 4441 1311 4445
rect 1315 4441 1317 4445
rect 1309 4440 1317 4441
rect 1309 4436 1311 4440
rect 1315 4436 1317 4440
rect 1309 4435 1317 4436
rect 1309 4431 1311 4435
rect 1315 4431 1317 4435
rect 1309 4430 1317 4431
rect 1309 4426 1311 4430
rect 1315 4426 1317 4430
rect 1309 4425 1317 4426
rect 1309 4421 1311 4425
rect 1315 4421 1317 4425
rect 1309 4420 1317 4421
rect 1309 4416 1311 4420
rect 1315 4416 1317 4420
rect 1309 4415 1317 4416
rect 1309 4411 1311 4415
rect 1315 4411 1317 4415
rect 1309 4410 1317 4411
rect 1309 4406 1311 4410
rect 1315 4406 1317 4410
rect 1309 4405 1317 4406
rect 1309 4401 1311 4405
rect 1315 4401 1317 4405
rect 1309 4400 1317 4401
rect 1309 4396 1311 4400
rect 1315 4396 1317 4400
rect 1309 4395 1317 4396
rect 1309 4391 1311 4395
rect 1315 4391 1317 4395
rect 1309 4390 1317 4391
rect 1309 4386 1311 4390
rect 1315 4386 1317 4390
rect 1309 4385 1317 4386
rect 1309 4381 1311 4385
rect 1315 4381 1317 4385
rect 1309 4380 1317 4381
rect 1309 4376 1311 4380
rect 1315 4376 1317 4380
rect 1309 4375 1317 4376
rect 1309 4371 1311 4375
rect 1315 4371 1317 4375
rect 1309 4370 1317 4371
rect 1309 4366 1311 4370
rect 1315 4366 1317 4370
rect 1309 4365 1317 4366
rect 1309 4361 1311 4365
rect 1315 4361 1317 4365
rect 1245 4360 1253 4361
rect 1245 4356 1247 4360
rect 1251 4356 1253 4360
rect 1245 4355 1253 4356
rect 1309 4360 1317 4361
rect 1309 4356 1311 4360
rect 1315 4356 1317 4360
rect 1309 4355 1317 4356
rect 1245 4353 1317 4355
rect 1245 4349 1247 4353
rect 1251 4349 1254 4353
rect 1258 4349 1259 4353
rect 1263 4349 1264 4353
rect 1268 4349 1269 4353
rect 1273 4349 1274 4353
rect 1278 4349 1279 4353
rect 1283 4349 1284 4353
rect 1288 4349 1289 4353
rect 1293 4349 1294 4353
rect 1298 4349 1299 4353
rect 1303 4349 1304 4353
rect 1308 4349 1311 4353
rect 1315 4349 1317 4353
rect 1245 4347 1317 4349
rect 1382 4475 1478 4476
rect 1382 4471 1383 4475
rect 1387 4471 1388 4475
rect 1392 4471 1393 4475
rect 1397 4471 1398 4475
rect 1402 4471 1403 4475
rect 1407 4471 1408 4475
rect 1412 4471 1413 4475
rect 1417 4471 1418 4475
rect 1422 4471 1423 4475
rect 1427 4471 1428 4475
rect 1432 4471 1433 4475
rect 1437 4471 1438 4475
rect 1442 4471 1443 4475
rect 1447 4471 1448 4475
rect 1452 4471 1453 4475
rect 1457 4471 1458 4475
rect 1462 4471 1463 4475
rect 1467 4471 1468 4475
rect 1472 4471 1473 4475
rect 1477 4471 1478 4475
rect 1382 4470 1478 4471
rect 1382 4466 1383 4470
rect 1387 4466 1388 4470
rect 1382 4465 1388 4466
rect 1382 4461 1383 4465
rect 1387 4461 1388 4465
rect 1472 4466 1473 4470
rect 1477 4466 1478 4470
rect 1472 4465 1478 4466
rect 1382 4460 1388 4461
rect 1382 4456 1383 4460
rect 1387 4456 1388 4460
rect 1382 4455 1388 4456
rect 1382 4451 1383 4455
rect 1387 4451 1388 4455
rect 1382 4450 1388 4451
rect 1382 4446 1383 4450
rect 1387 4446 1388 4450
rect 1382 4445 1388 4446
rect 1382 4441 1383 4445
rect 1387 4441 1388 4445
rect 1382 4440 1388 4441
rect 1382 4436 1383 4440
rect 1387 4436 1388 4440
rect 1382 4435 1388 4436
rect 1382 4431 1383 4435
rect 1387 4431 1388 4435
rect 1382 4430 1388 4431
rect 1382 4426 1383 4430
rect 1387 4426 1388 4430
rect 1382 4425 1388 4426
rect 1382 4421 1383 4425
rect 1387 4421 1388 4425
rect 1382 4420 1388 4421
rect 1382 4416 1383 4420
rect 1387 4416 1388 4420
rect 1382 4415 1388 4416
rect 1382 4411 1383 4415
rect 1387 4411 1388 4415
rect 1382 4410 1388 4411
rect 1382 4406 1383 4410
rect 1387 4406 1388 4410
rect 1382 4405 1388 4406
rect 1382 4401 1383 4405
rect 1387 4401 1388 4405
rect 1382 4400 1388 4401
rect 1382 4396 1383 4400
rect 1387 4396 1388 4400
rect 1382 4395 1388 4396
rect 1382 4391 1383 4395
rect 1387 4391 1388 4395
rect 1382 4390 1388 4391
rect 1382 4386 1383 4390
rect 1387 4386 1388 4390
rect 1382 4385 1388 4386
rect 1382 4381 1383 4385
rect 1387 4381 1388 4385
rect 1382 4380 1388 4381
rect 1382 4376 1383 4380
rect 1387 4376 1388 4380
rect 1382 4375 1388 4376
rect 1382 4371 1383 4375
rect 1387 4371 1388 4375
rect 1382 4370 1388 4371
rect 1382 4366 1383 4370
rect 1387 4366 1388 4370
rect 1382 4365 1388 4366
rect 1382 4361 1383 4365
rect 1387 4361 1388 4365
rect 1382 4360 1388 4361
rect 1382 4356 1383 4360
rect 1387 4356 1388 4360
rect 1382 4355 1388 4356
rect 1382 4351 1383 4355
rect 1387 4351 1388 4355
rect 1382 4350 1388 4351
rect 1382 4346 1383 4350
rect 1387 4346 1388 4350
rect 1472 4461 1473 4465
rect 1477 4461 1478 4465
rect 1472 4460 1478 4461
rect 1472 4456 1473 4460
rect 1477 4456 1478 4460
rect 1472 4455 1478 4456
rect 1472 4451 1473 4455
rect 1477 4451 1478 4455
rect 1472 4450 1478 4451
rect 1472 4446 1473 4450
rect 1477 4446 1478 4450
rect 1472 4445 1478 4446
rect 1472 4441 1473 4445
rect 1477 4441 1478 4445
rect 1472 4440 1478 4441
rect 1472 4436 1473 4440
rect 1477 4436 1478 4440
rect 1472 4435 1478 4436
rect 1472 4431 1473 4435
rect 1477 4431 1478 4435
rect 1472 4430 1478 4431
rect 1472 4426 1473 4430
rect 1477 4426 1478 4430
rect 1472 4425 1478 4426
rect 1472 4421 1473 4425
rect 1477 4421 1478 4425
rect 1472 4420 1478 4421
rect 1472 4416 1473 4420
rect 1477 4416 1478 4420
rect 1472 4415 1478 4416
rect 1472 4411 1473 4415
rect 1477 4411 1478 4415
rect 1472 4410 1478 4411
rect 1472 4406 1473 4410
rect 1477 4406 1478 4410
rect 1472 4405 1478 4406
rect 1472 4401 1473 4405
rect 1477 4401 1478 4405
rect 1472 4400 1478 4401
rect 1472 4396 1473 4400
rect 1477 4396 1478 4400
rect 1472 4395 1478 4396
rect 1472 4391 1473 4395
rect 1477 4391 1478 4395
rect 1472 4390 1478 4391
rect 1472 4386 1473 4390
rect 1477 4386 1478 4390
rect 1472 4385 1478 4386
rect 1472 4381 1473 4385
rect 1477 4381 1478 4385
rect 1472 4380 1478 4381
rect 1472 4376 1473 4380
rect 1477 4376 1478 4380
rect 1472 4375 1478 4376
rect 1472 4371 1473 4375
rect 1477 4371 1478 4375
rect 1472 4370 1478 4371
rect 1472 4366 1473 4370
rect 1477 4366 1478 4370
rect 1472 4365 1478 4366
rect 1472 4361 1473 4365
rect 1477 4361 1478 4365
rect 1472 4360 1478 4361
rect 1472 4356 1473 4360
rect 1477 4356 1478 4360
rect 1472 4355 1478 4356
rect 1472 4351 1473 4355
rect 1477 4351 1478 4355
rect 1472 4350 1478 4351
rect 1382 4345 1388 4346
rect 1382 4341 1383 4345
rect 1387 4341 1388 4345
rect 1472 4346 1473 4350
rect 1477 4346 1478 4350
rect 1472 4345 1478 4346
rect 1472 4341 1473 4345
rect 1477 4341 1478 4345
rect 1382 4340 1478 4341
rect 1382 4336 1383 4340
rect 1387 4336 1388 4340
rect 1392 4336 1393 4340
rect 1397 4336 1398 4340
rect 1402 4336 1403 4340
rect 1407 4336 1408 4340
rect 1412 4336 1413 4340
rect 1417 4336 1418 4340
rect 1422 4336 1423 4340
rect 1427 4336 1428 4340
rect 1432 4336 1433 4340
rect 1437 4336 1438 4340
rect 1442 4336 1443 4340
rect 1447 4336 1448 4340
rect 1452 4336 1453 4340
rect 1457 4336 1458 4340
rect 1462 4336 1463 4340
rect 1467 4336 1468 4340
rect 1472 4336 1473 4340
rect 1477 4336 1478 4340
rect 1382 4335 1478 4336
rect 1554 4462 1626 4464
rect 1554 4458 1556 4462
rect 1560 4458 1563 4462
rect 1567 4458 1568 4462
rect 1572 4458 1573 4462
rect 1577 4458 1578 4462
rect 1582 4458 1583 4462
rect 1587 4458 1588 4462
rect 1592 4458 1593 4462
rect 1597 4458 1598 4462
rect 1602 4458 1603 4462
rect 1607 4458 1608 4462
rect 1612 4458 1613 4462
rect 1617 4458 1620 4462
rect 1624 4458 1626 4462
rect 1554 4456 1626 4458
rect 1554 4455 1562 4456
rect 1554 4451 1556 4455
rect 1560 4451 1562 4455
rect 1554 4450 1562 4451
rect 1618 4455 1626 4456
rect 1618 4451 1620 4455
rect 1624 4451 1626 4455
rect 1618 4450 1626 4451
rect 1554 4446 1556 4450
rect 1560 4446 1562 4450
rect 1554 4445 1562 4446
rect 1554 4441 1556 4445
rect 1560 4441 1562 4445
rect 1554 4440 1562 4441
rect 1554 4436 1556 4440
rect 1560 4436 1562 4440
rect 1554 4435 1562 4436
rect 1554 4431 1556 4435
rect 1560 4431 1562 4435
rect 1554 4430 1562 4431
rect 1554 4426 1556 4430
rect 1560 4426 1562 4430
rect 1554 4425 1562 4426
rect 1554 4421 1556 4425
rect 1560 4421 1562 4425
rect 1554 4420 1562 4421
rect 1554 4416 1556 4420
rect 1560 4416 1562 4420
rect 1554 4415 1562 4416
rect 1554 4411 1556 4415
rect 1560 4411 1562 4415
rect 1554 4410 1562 4411
rect 1554 4406 1556 4410
rect 1560 4406 1562 4410
rect 1554 4405 1562 4406
rect 1554 4401 1556 4405
rect 1560 4401 1562 4405
rect 1554 4400 1562 4401
rect 1554 4396 1556 4400
rect 1560 4396 1562 4400
rect 1554 4395 1562 4396
rect 1554 4391 1556 4395
rect 1560 4391 1562 4395
rect 1554 4390 1562 4391
rect 1554 4386 1556 4390
rect 1560 4386 1562 4390
rect 1554 4385 1562 4386
rect 1554 4381 1556 4385
rect 1560 4381 1562 4385
rect 1554 4380 1562 4381
rect 1554 4376 1556 4380
rect 1560 4376 1562 4380
rect 1554 4375 1562 4376
rect 1554 4371 1556 4375
rect 1560 4371 1562 4375
rect 1554 4370 1562 4371
rect 1554 4366 1556 4370
rect 1560 4366 1562 4370
rect 1554 4365 1562 4366
rect 1554 4361 1556 4365
rect 1560 4361 1562 4365
rect 1618 4446 1620 4450
rect 1624 4446 1626 4450
rect 1618 4445 1626 4446
rect 1618 4441 1620 4445
rect 1624 4441 1626 4445
rect 1618 4440 1626 4441
rect 1618 4436 1620 4440
rect 1624 4436 1626 4440
rect 1618 4435 1626 4436
rect 1618 4431 1620 4435
rect 1624 4431 1626 4435
rect 1618 4430 1626 4431
rect 1618 4426 1620 4430
rect 1624 4426 1626 4430
rect 1618 4425 1626 4426
rect 1618 4421 1620 4425
rect 1624 4421 1626 4425
rect 1618 4420 1626 4421
rect 1618 4416 1620 4420
rect 1624 4416 1626 4420
rect 1618 4415 1626 4416
rect 1618 4411 1620 4415
rect 1624 4411 1626 4415
rect 1618 4410 1626 4411
rect 1618 4406 1620 4410
rect 1624 4406 1626 4410
rect 1618 4405 1626 4406
rect 1618 4401 1620 4405
rect 1624 4401 1626 4405
rect 1618 4400 1626 4401
rect 1618 4396 1620 4400
rect 1624 4396 1626 4400
rect 1618 4395 1626 4396
rect 1618 4391 1620 4395
rect 1624 4391 1626 4395
rect 1618 4390 1626 4391
rect 1618 4386 1620 4390
rect 1624 4386 1626 4390
rect 1618 4385 1626 4386
rect 1618 4381 1620 4385
rect 1624 4381 1626 4385
rect 1618 4380 1626 4381
rect 1618 4376 1620 4380
rect 1624 4376 1626 4380
rect 1618 4375 1626 4376
rect 1618 4371 1620 4375
rect 1624 4371 1626 4375
rect 1618 4370 1626 4371
rect 1618 4366 1620 4370
rect 1624 4366 1626 4370
rect 1618 4365 1626 4366
rect 1618 4361 1620 4365
rect 1624 4361 1626 4365
rect 1554 4360 1562 4361
rect 1554 4356 1556 4360
rect 1560 4356 1562 4360
rect 1554 4355 1562 4356
rect 1618 4360 1626 4361
rect 1618 4356 1620 4360
rect 1624 4356 1626 4360
rect 1618 4355 1626 4356
rect 1554 4353 1626 4355
rect 1554 4349 1556 4353
rect 1560 4349 1563 4353
rect 1567 4349 1568 4353
rect 1572 4349 1573 4353
rect 1577 4349 1578 4353
rect 1582 4349 1583 4353
rect 1587 4349 1588 4353
rect 1592 4349 1593 4353
rect 1597 4349 1598 4353
rect 1602 4349 1603 4353
rect 1607 4349 1608 4353
rect 1612 4349 1613 4353
rect 1617 4349 1620 4353
rect 1624 4349 1626 4353
rect 1554 4347 1626 4349
rect 1691 4475 1787 4476
rect 1691 4471 1692 4475
rect 1696 4471 1697 4475
rect 1701 4471 1702 4475
rect 1706 4471 1707 4475
rect 1711 4471 1712 4475
rect 1716 4471 1717 4475
rect 1721 4471 1722 4475
rect 1726 4471 1727 4475
rect 1731 4471 1732 4475
rect 1736 4471 1737 4475
rect 1741 4471 1742 4475
rect 1746 4471 1747 4475
rect 1751 4471 1752 4475
rect 1756 4471 1757 4475
rect 1761 4471 1762 4475
rect 1766 4471 1767 4475
rect 1771 4471 1772 4475
rect 1776 4471 1777 4475
rect 1781 4471 1782 4475
rect 1786 4471 1787 4475
rect 1691 4470 1787 4471
rect 1691 4466 1692 4470
rect 1696 4466 1697 4470
rect 1691 4465 1697 4466
rect 1691 4461 1692 4465
rect 1696 4461 1697 4465
rect 1781 4466 1782 4470
rect 1786 4466 1787 4470
rect 1781 4465 1787 4466
rect 1691 4460 1697 4461
rect 1691 4456 1692 4460
rect 1696 4456 1697 4460
rect 1691 4455 1697 4456
rect 1691 4451 1692 4455
rect 1696 4451 1697 4455
rect 1691 4450 1697 4451
rect 1691 4446 1692 4450
rect 1696 4446 1697 4450
rect 1691 4445 1697 4446
rect 1691 4441 1692 4445
rect 1696 4441 1697 4445
rect 1691 4440 1697 4441
rect 1691 4436 1692 4440
rect 1696 4436 1697 4440
rect 1691 4435 1697 4436
rect 1691 4431 1692 4435
rect 1696 4431 1697 4435
rect 1691 4430 1697 4431
rect 1691 4426 1692 4430
rect 1696 4426 1697 4430
rect 1691 4425 1697 4426
rect 1691 4421 1692 4425
rect 1696 4421 1697 4425
rect 1691 4420 1697 4421
rect 1691 4416 1692 4420
rect 1696 4416 1697 4420
rect 1691 4415 1697 4416
rect 1691 4411 1692 4415
rect 1696 4411 1697 4415
rect 1691 4410 1697 4411
rect 1691 4406 1692 4410
rect 1696 4406 1697 4410
rect 1691 4405 1697 4406
rect 1691 4401 1692 4405
rect 1696 4401 1697 4405
rect 1691 4400 1697 4401
rect 1691 4396 1692 4400
rect 1696 4396 1697 4400
rect 1691 4395 1697 4396
rect 1691 4391 1692 4395
rect 1696 4391 1697 4395
rect 1691 4390 1697 4391
rect 1691 4386 1692 4390
rect 1696 4386 1697 4390
rect 1691 4385 1697 4386
rect 1691 4381 1692 4385
rect 1696 4381 1697 4385
rect 1691 4380 1697 4381
rect 1691 4376 1692 4380
rect 1696 4376 1697 4380
rect 1691 4375 1697 4376
rect 1691 4371 1692 4375
rect 1696 4371 1697 4375
rect 1691 4370 1697 4371
rect 1691 4366 1692 4370
rect 1696 4366 1697 4370
rect 1691 4365 1697 4366
rect 1691 4361 1692 4365
rect 1696 4361 1697 4365
rect 1691 4360 1697 4361
rect 1691 4356 1692 4360
rect 1696 4356 1697 4360
rect 1691 4355 1697 4356
rect 1691 4351 1692 4355
rect 1696 4351 1697 4355
rect 1691 4350 1697 4351
rect 1691 4346 1692 4350
rect 1696 4346 1697 4350
rect 1781 4461 1782 4465
rect 1786 4461 1787 4465
rect 1781 4460 1787 4461
rect 1781 4456 1782 4460
rect 1786 4456 1787 4460
rect 1781 4455 1787 4456
rect 1781 4451 1782 4455
rect 1786 4451 1787 4455
rect 1781 4450 1787 4451
rect 1781 4446 1782 4450
rect 1786 4446 1787 4450
rect 1781 4445 1787 4446
rect 1781 4441 1782 4445
rect 1786 4441 1787 4445
rect 1781 4440 1787 4441
rect 1781 4436 1782 4440
rect 1786 4436 1787 4440
rect 1781 4435 1787 4436
rect 1781 4431 1782 4435
rect 1786 4431 1787 4435
rect 1781 4430 1787 4431
rect 1781 4426 1782 4430
rect 1786 4426 1787 4430
rect 1781 4425 1787 4426
rect 1781 4421 1782 4425
rect 1786 4421 1787 4425
rect 1781 4420 1787 4421
rect 1781 4416 1782 4420
rect 1786 4416 1787 4420
rect 1781 4415 1787 4416
rect 1781 4411 1782 4415
rect 1786 4411 1787 4415
rect 1781 4410 1787 4411
rect 1781 4406 1782 4410
rect 1786 4406 1787 4410
rect 1781 4405 1787 4406
rect 1781 4401 1782 4405
rect 1786 4401 1787 4405
rect 1781 4400 1787 4401
rect 1781 4396 1782 4400
rect 1786 4396 1787 4400
rect 1781 4395 1787 4396
rect 1781 4391 1782 4395
rect 1786 4391 1787 4395
rect 1781 4390 1787 4391
rect 1781 4386 1782 4390
rect 1786 4386 1787 4390
rect 1781 4385 1787 4386
rect 1781 4381 1782 4385
rect 1786 4381 1787 4385
rect 1781 4380 1787 4381
rect 1781 4376 1782 4380
rect 1786 4376 1787 4380
rect 1781 4375 1787 4376
rect 1781 4371 1782 4375
rect 1786 4371 1787 4375
rect 1781 4370 1787 4371
rect 1781 4366 1782 4370
rect 1786 4366 1787 4370
rect 1781 4365 1787 4366
rect 1781 4361 1782 4365
rect 1786 4361 1787 4365
rect 1781 4360 1787 4361
rect 1781 4356 1782 4360
rect 1786 4356 1787 4360
rect 1781 4355 1787 4356
rect 1781 4351 1782 4355
rect 1786 4351 1787 4355
rect 1781 4350 1787 4351
rect 1691 4345 1697 4346
rect 1691 4341 1692 4345
rect 1696 4341 1697 4345
rect 1781 4346 1782 4350
rect 1786 4346 1787 4350
rect 1781 4345 1787 4346
rect 1781 4341 1782 4345
rect 1786 4341 1787 4345
rect 1691 4340 1787 4341
rect 1691 4336 1692 4340
rect 1696 4336 1697 4340
rect 1701 4336 1702 4340
rect 1706 4336 1707 4340
rect 1711 4336 1712 4340
rect 1716 4336 1717 4340
rect 1721 4336 1722 4340
rect 1726 4336 1727 4340
rect 1731 4336 1732 4340
rect 1736 4336 1737 4340
rect 1741 4336 1742 4340
rect 1746 4336 1747 4340
rect 1751 4336 1752 4340
rect 1756 4336 1757 4340
rect 1761 4336 1762 4340
rect 1766 4336 1767 4340
rect 1771 4336 1772 4340
rect 1776 4336 1777 4340
rect 1781 4336 1782 4340
rect 1786 4336 1787 4340
rect 1691 4335 1787 4336
rect 1863 4462 1935 4464
rect 1863 4458 1865 4462
rect 1869 4458 1872 4462
rect 1876 4458 1877 4462
rect 1881 4458 1882 4462
rect 1886 4458 1887 4462
rect 1891 4458 1892 4462
rect 1896 4458 1897 4462
rect 1901 4458 1902 4462
rect 1906 4458 1907 4462
rect 1911 4458 1912 4462
rect 1916 4458 1917 4462
rect 1921 4458 1922 4462
rect 1926 4458 1929 4462
rect 1933 4458 1935 4462
rect 1863 4456 1935 4458
rect 1863 4455 1871 4456
rect 1863 4451 1865 4455
rect 1869 4451 1871 4455
rect 1863 4450 1871 4451
rect 1927 4455 1935 4456
rect 1927 4451 1929 4455
rect 1933 4451 1935 4455
rect 1927 4450 1935 4451
rect 1863 4446 1865 4450
rect 1869 4446 1871 4450
rect 1863 4445 1871 4446
rect 1863 4441 1865 4445
rect 1869 4441 1871 4445
rect 1863 4440 1871 4441
rect 1863 4436 1865 4440
rect 1869 4436 1871 4440
rect 1863 4435 1871 4436
rect 1863 4431 1865 4435
rect 1869 4431 1871 4435
rect 1863 4430 1871 4431
rect 1863 4426 1865 4430
rect 1869 4426 1871 4430
rect 1863 4425 1871 4426
rect 1863 4421 1865 4425
rect 1869 4421 1871 4425
rect 1863 4420 1871 4421
rect 1863 4416 1865 4420
rect 1869 4416 1871 4420
rect 1863 4415 1871 4416
rect 1863 4411 1865 4415
rect 1869 4411 1871 4415
rect 1863 4410 1871 4411
rect 1863 4406 1865 4410
rect 1869 4406 1871 4410
rect 1863 4405 1871 4406
rect 1863 4401 1865 4405
rect 1869 4401 1871 4405
rect 1863 4400 1871 4401
rect 1863 4396 1865 4400
rect 1869 4396 1871 4400
rect 1863 4395 1871 4396
rect 1863 4391 1865 4395
rect 1869 4391 1871 4395
rect 1863 4390 1871 4391
rect 1863 4386 1865 4390
rect 1869 4386 1871 4390
rect 1863 4385 1871 4386
rect 1863 4381 1865 4385
rect 1869 4381 1871 4385
rect 1863 4380 1871 4381
rect 1863 4376 1865 4380
rect 1869 4376 1871 4380
rect 1863 4375 1871 4376
rect 1863 4371 1865 4375
rect 1869 4371 1871 4375
rect 1863 4370 1871 4371
rect 1863 4366 1865 4370
rect 1869 4366 1871 4370
rect 1863 4365 1871 4366
rect 1863 4361 1865 4365
rect 1869 4361 1871 4365
rect 1927 4446 1929 4450
rect 1933 4446 1935 4450
rect 1927 4445 1935 4446
rect 1927 4441 1929 4445
rect 1933 4441 1935 4445
rect 1927 4440 1935 4441
rect 1927 4436 1929 4440
rect 1933 4436 1935 4440
rect 1927 4435 1935 4436
rect 1927 4431 1929 4435
rect 1933 4431 1935 4435
rect 1927 4430 1935 4431
rect 1927 4426 1929 4430
rect 1933 4426 1935 4430
rect 1927 4425 1935 4426
rect 1927 4421 1929 4425
rect 1933 4421 1935 4425
rect 1927 4420 1935 4421
rect 1927 4416 1929 4420
rect 1933 4416 1935 4420
rect 1927 4415 1935 4416
rect 1927 4411 1929 4415
rect 1933 4411 1935 4415
rect 1927 4410 1935 4411
rect 1927 4406 1929 4410
rect 1933 4406 1935 4410
rect 1927 4405 1935 4406
rect 1927 4401 1929 4405
rect 1933 4401 1935 4405
rect 1927 4400 1935 4401
rect 1927 4396 1929 4400
rect 1933 4396 1935 4400
rect 1927 4395 1935 4396
rect 1927 4391 1929 4395
rect 1933 4391 1935 4395
rect 1927 4390 1935 4391
rect 1927 4386 1929 4390
rect 1933 4386 1935 4390
rect 1927 4385 1935 4386
rect 1927 4381 1929 4385
rect 1933 4381 1935 4385
rect 1927 4380 1935 4381
rect 1927 4376 1929 4380
rect 1933 4376 1935 4380
rect 1927 4375 1935 4376
rect 1927 4371 1929 4375
rect 1933 4371 1935 4375
rect 1927 4370 1935 4371
rect 1927 4366 1929 4370
rect 1933 4366 1935 4370
rect 1927 4365 1935 4366
rect 1927 4361 1929 4365
rect 1933 4361 1935 4365
rect 1863 4360 1871 4361
rect 1863 4356 1865 4360
rect 1869 4356 1871 4360
rect 1863 4355 1871 4356
rect 1927 4360 1935 4361
rect 1927 4356 1929 4360
rect 1933 4356 1935 4360
rect 1927 4355 1935 4356
rect 1863 4353 1935 4355
rect 1863 4349 1865 4353
rect 1869 4349 1872 4353
rect 1876 4349 1877 4353
rect 1881 4349 1882 4353
rect 1886 4349 1887 4353
rect 1891 4349 1892 4353
rect 1896 4349 1897 4353
rect 1901 4349 1902 4353
rect 1906 4349 1907 4353
rect 1911 4349 1912 4353
rect 1916 4349 1917 4353
rect 1921 4349 1922 4353
rect 1926 4349 1929 4353
rect 1933 4349 1935 4353
rect 1863 4347 1935 4349
rect 2000 4475 2096 4476
rect 2000 4471 2001 4475
rect 2005 4471 2006 4475
rect 2010 4471 2011 4475
rect 2015 4471 2016 4475
rect 2020 4471 2021 4475
rect 2025 4471 2026 4475
rect 2030 4471 2031 4475
rect 2035 4471 2036 4475
rect 2040 4471 2041 4475
rect 2045 4471 2046 4475
rect 2050 4471 2051 4475
rect 2055 4471 2056 4475
rect 2060 4471 2061 4475
rect 2065 4471 2066 4475
rect 2070 4471 2071 4475
rect 2075 4471 2076 4475
rect 2080 4471 2081 4475
rect 2085 4471 2086 4475
rect 2090 4471 2091 4475
rect 2095 4471 2096 4475
rect 2000 4470 2096 4471
rect 2000 4466 2001 4470
rect 2005 4466 2006 4470
rect 2000 4465 2006 4466
rect 2000 4461 2001 4465
rect 2005 4461 2006 4465
rect 2090 4466 2091 4470
rect 2095 4466 2096 4470
rect 2090 4465 2096 4466
rect 2000 4460 2006 4461
rect 2000 4456 2001 4460
rect 2005 4456 2006 4460
rect 2000 4455 2006 4456
rect 2000 4451 2001 4455
rect 2005 4451 2006 4455
rect 2000 4450 2006 4451
rect 2000 4446 2001 4450
rect 2005 4446 2006 4450
rect 2000 4445 2006 4446
rect 2000 4441 2001 4445
rect 2005 4441 2006 4445
rect 2000 4440 2006 4441
rect 2000 4436 2001 4440
rect 2005 4436 2006 4440
rect 2000 4435 2006 4436
rect 2000 4431 2001 4435
rect 2005 4431 2006 4435
rect 2000 4430 2006 4431
rect 2000 4426 2001 4430
rect 2005 4426 2006 4430
rect 2000 4425 2006 4426
rect 2000 4421 2001 4425
rect 2005 4421 2006 4425
rect 2000 4420 2006 4421
rect 2000 4416 2001 4420
rect 2005 4416 2006 4420
rect 2000 4415 2006 4416
rect 2000 4411 2001 4415
rect 2005 4411 2006 4415
rect 2000 4410 2006 4411
rect 2000 4406 2001 4410
rect 2005 4406 2006 4410
rect 2000 4405 2006 4406
rect 2000 4401 2001 4405
rect 2005 4401 2006 4405
rect 2000 4400 2006 4401
rect 2000 4396 2001 4400
rect 2005 4396 2006 4400
rect 2000 4395 2006 4396
rect 2000 4391 2001 4395
rect 2005 4391 2006 4395
rect 2000 4390 2006 4391
rect 2000 4386 2001 4390
rect 2005 4386 2006 4390
rect 2000 4385 2006 4386
rect 2000 4381 2001 4385
rect 2005 4381 2006 4385
rect 2000 4380 2006 4381
rect 2000 4376 2001 4380
rect 2005 4376 2006 4380
rect 2000 4375 2006 4376
rect 2000 4371 2001 4375
rect 2005 4371 2006 4375
rect 2000 4370 2006 4371
rect 2000 4366 2001 4370
rect 2005 4366 2006 4370
rect 2000 4365 2006 4366
rect 2000 4361 2001 4365
rect 2005 4361 2006 4365
rect 2000 4360 2006 4361
rect 2000 4356 2001 4360
rect 2005 4356 2006 4360
rect 2000 4355 2006 4356
rect 2000 4351 2001 4355
rect 2005 4351 2006 4355
rect 2000 4350 2006 4351
rect 2000 4346 2001 4350
rect 2005 4346 2006 4350
rect 2090 4461 2091 4465
rect 2095 4461 2096 4465
rect 2090 4460 2096 4461
rect 2090 4456 2091 4460
rect 2095 4456 2096 4460
rect 2090 4455 2096 4456
rect 2090 4451 2091 4455
rect 2095 4451 2096 4455
rect 2090 4450 2096 4451
rect 2090 4446 2091 4450
rect 2095 4446 2096 4450
rect 2090 4445 2096 4446
rect 2090 4441 2091 4445
rect 2095 4441 2096 4445
rect 2090 4440 2096 4441
rect 2090 4436 2091 4440
rect 2095 4436 2096 4440
rect 2090 4435 2096 4436
rect 2090 4431 2091 4435
rect 2095 4431 2096 4435
rect 2090 4430 2096 4431
rect 2090 4426 2091 4430
rect 2095 4426 2096 4430
rect 2090 4425 2096 4426
rect 2090 4421 2091 4425
rect 2095 4421 2096 4425
rect 2090 4420 2096 4421
rect 2090 4416 2091 4420
rect 2095 4416 2096 4420
rect 2090 4415 2096 4416
rect 2090 4411 2091 4415
rect 2095 4411 2096 4415
rect 2090 4410 2096 4411
rect 2090 4406 2091 4410
rect 2095 4406 2096 4410
rect 2090 4405 2096 4406
rect 2090 4401 2091 4405
rect 2095 4401 2096 4405
rect 2090 4400 2096 4401
rect 2090 4396 2091 4400
rect 2095 4396 2096 4400
rect 2090 4395 2096 4396
rect 2090 4391 2091 4395
rect 2095 4391 2096 4395
rect 2090 4390 2096 4391
rect 2090 4386 2091 4390
rect 2095 4386 2096 4390
rect 2090 4385 2096 4386
rect 2090 4381 2091 4385
rect 2095 4381 2096 4385
rect 2090 4380 2096 4381
rect 2090 4376 2091 4380
rect 2095 4376 2096 4380
rect 2090 4375 2096 4376
rect 2090 4371 2091 4375
rect 2095 4371 2096 4375
rect 2090 4370 2096 4371
rect 2090 4366 2091 4370
rect 2095 4366 2096 4370
rect 2090 4365 2096 4366
rect 2090 4361 2091 4365
rect 2095 4361 2096 4365
rect 2090 4360 2096 4361
rect 2090 4356 2091 4360
rect 2095 4356 2096 4360
rect 2090 4355 2096 4356
rect 2090 4351 2091 4355
rect 2095 4351 2096 4355
rect 2090 4350 2096 4351
rect 2000 4345 2006 4346
rect 2000 4341 2001 4345
rect 2005 4341 2006 4345
rect 2090 4346 2091 4350
rect 2095 4346 2096 4350
rect 2090 4345 2096 4346
rect 2090 4341 2091 4345
rect 2095 4341 2096 4345
rect 2000 4340 2096 4341
rect 2000 4336 2001 4340
rect 2005 4336 2006 4340
rect 2010 4336 2011 4340
rect 2015 4336 2016 4340
rect 2020 4336 2021 4340
rect 2025 4336 2026 4340
rect 2030 4336 2031 4340
rect 2035 4336 2036 4340
rect 2040 4336 2041 4340
rect 2045 4336 2046 4340
rect 2050 4336 2051 4340
rect 2055 4336 2056 4340
rect 2060 4336 2061 4340
rect 2065 4336 2066 4340
rect 2070 4336 2071 4340
rect 2075 4336 2076 4340
rect 2080 4336 2081 4340
rect 2085 4336 2086 4340
rect 2090 4336 2091 4340
rect 2095 4336 2096 4340
rect 2000 4335 2096 4336
rect 2172 4462 2244 4464
rect 2172 4458 2174 4462
rect 2178 4458 2181 4462
rect 2185 4458 2186 4462
rect 2190 4458 2191 4462
rect 2195 4458 2196 4462
rect 2200 4458 2201 4462
rect 2205 4458 2206 4462
rect 2210 4458 2211 4462
rect 2215 4458 2216 4462
rect 2220 4458 2221 4462
rect 2225 4458 2226 4462
rect 2230 4458 2231 4462
rect 2235 4458 2238 4462
rect 2242 4458 2244 4462
rect 2172 4456 2244 4458
rect 2172 4455 2180 4456
rect 2172 4451 2174 4455
rect 2178 4451 2180 4455
rect 2172 4450 2180 4451
rect 2236 4455 2244 4456
rect 2236 4451 2238 4455
rect 2242 4451 2244 4455
rect 2236 4450 2244 4451
rect 2172 4446 2174 4450
rect 2178 4446 2180 4450
rect 2172 4445 2180 4446
rect 2172 4441 2174 4445
rect 2178 4441 2180 4445
rect 2172 4440 2180 4441
rect 2172 4436 2174 4440
rect 2178 4436 2180 4440
rect 2172 4435 2180 4436
rect 2172 4431 2174 4435
rect 2178 4431 2180 4435
rect 2172 4430 2180 4431
rect 2172 4426 2174 4430
rect 2178 4426 2180 4430
rect 2172 4425 2180 4426
rect 2172 4421 2174 4425
rect 2178 4421 2180 4425
rect 2172 4420 2180 4421
rect 2172 4416 2174 4420
rect 2178 4416 2180 4420
rect 2172 4415 2180 4416
rect 2172 4411 2174 4415
rect 2178 4411 2180 4415
rect 2172 4410 2180 4411
rect 2172 4406 2174 4410
rect 2178 4406 2180 4410
rect 2172 4405 2180 4406
rect 2172 4401 2174 4405
rect 2178 4401 2180 4405
rect 2172 4400 2180 4401
rect 2172 4396 2174 4400
rect 2178 4396 2180 4400
rect 2172 4395 2180 4396
rect 2172 4391 2174 4395
rect 2178 4391 2180 4395
rect 2172 4390 2180 4391
rect 2172 4386 2174 4390
rect 2178 4386 2180 4390
rect 2172 4385 2180 4386
rect 2172 4381 2174 4385
rect 2178 4381 2180 4385
rect 2172 4380 2180 4381
rect 2172 4376 2174 4380
rect 2178 4376 2180 4380
rect 2172 4375 2180 4376
rect 2172 4371 2174 4375
rect 2178 4371 2180 4375
rect 2172 4370 2180 4371
rect 2172 4366 2174 4370
rect 2178 4366 2180 4370
rect 2172 4365 2180 4366
rect 2172 4361 2174 4365
rect 2178 4361 2180 4365
rect 2236 4446 2238 4450
rect 2242 4446 2244 4450
rect 2236 4445 2244 4446
rect 2236 4441 2238 4445
rect 2242 4441 2244 4445
rect 2236 4440 2244 4441
rect 2236 4436 2238 4440
rect 2242 4436 2244 4440
rect 2236 4435 2244 4436
rect 2236 4431 2238 4435
rect 2242 4431 2244 4435
rect 2236 4430 2244 4431
rect 2236 4426 2238 4430
rect 2242 4426 2244 4430
rect 2236 4425 2244 4426
rect 2236 4421 2238 4425
rect 2242 4421 2244 4425
rect 2236 4420 2244 4421
rect 2236 4416 2238 4420
rect 2242 4416 2244 4420
rect 2236 4415 2244 4416
rect 2236 4411 2238 4415
rect 2242 4411 2244 4415
rect 2236 4410 2244 4411
rect 2236 4406 2238 4410
rect 2242 4406 2244 4410
rect 2236 4405 2244 4406
rect 2236 4401 2238 4405
rect 2242 4401 2244 4405
rect 2236 4400 2244 4401
rect 2236 4396 2238 4400
rect 2242 4396 2244 4400
rect 2236 4395 2244 4396
rect 2236 4391 2238 4395
rect 2242 4391 2244 4395
rect 2236 4390 2244 4391
rect 2236 4386 2238 4390
rect 2242 4386 2244 4390
rect 2236 4385 2244 4386
rect 2236 4381 2238 4385
rect 2242 4381 2244 4385
rect 2236 4380 2244 4381
rect 2236 4376 2238 4380
rect 2242 4376 2244 4380
rect 2236 4375 2244 4376
rect 2236 4371 2238 4375
rect 2242 4371 2244 4375
rect 2236 4370 2244 4371
rect 2236 4366 2238 4370
rect 2242 4366 2244 4370
rect 2236 4365 2244 4366
rect 2236 4361 2238 4365
rect 2242 4361 2244 4365
rect 2172 4360 2180 4361
rect 2172 4356 2174 4360
rect 2178 4356 2180 4360
rect 2172 4355 2180 4356
rect 2236 4360 2244 4361
rect 2236 4356 2238 4360
rect 2242 4356 2244 4360
rect 2236 4355 2244 4356
rect 2172 4353 2244 4355
rect 2172 4349 2174 4353
rect 2178 4349 2181 4353
rect 2185 4349 2186 4353
rect 2190 4349 2191 4353
rect 2195 4349 2196 4353
rect 2200 4349 2201 4353
rect 2205 4349 2206 4353
rect 2210 4349 2211 4353
rect 2215 4349 2216 4353
rect 2220 4349 2221 4353
rect 2225 4349 2226 4353
rect 2230 4349 2231 4353
rect 2235 4349 2238 4353
rect 2242 4349 2244 4353
rect 2172 4347 2244 4349
rect 2309 4475 2405 4476
rect 2309 4471 2310 4475
rect 2314 4471 2315 4475
rect 2319 4471 2320 4475
rect 2324 4471 2325 4475
rect 2329 4471 2330 4475
rect 2334 4471 2335 4475
rect 2339 4471 2340 4475
rect 2344 4471 2345 4475
rect 2349 4471 2350 4475
rect 2354 4471 2355 4475
rect 2359 4471 2360 4475
rect 2364 4471 2365 4475
rect 2369 4471 2370 4475
rect 2374 4471 2375 4475
rect 2379 4471 2380 4475
rect 2384 4471 2385 4475
rect 2389 4471 2390 4475
rect 2394 4471 2395 4475
rect 2399 4471 2400 4475
rect 2404 4471 2405 4475
rect 2309 4470 2405 4471
rect 2309 4466 2310 4470
rect 2314 4466 2315 4470
rect 2309 4465 2315 4466
rect 2309 4461 2310 4465
rect 2314 4461 2315 4465
rect 2399 4466 2400 4470
rect 2404 4466 2405 4470
rect 2399 4465 2405 4466
rect 2309 4460 2315 4461
rect 2309 4456 2310 4460
rect 2314 4456 2315 4460
rect 2309 4455 2315 4456
rect 2309 4451 2310 4455
rect 2314 4451 2315 4455
rect 2309 4450 2315 4451
rect 2309 4446 2310 4450
rect 2314 4446 2315 4450
rect 2309 4445 2315 4446
rect 2309 4441 2310 4445
rect 2314 4441 2315 4445
rect 2309 4440 2315 4441
rect 2309 4436 2310 4440
rect 2314 4436 2315 4440
rect 2309 4435 2315 4436
rect 2309 4431 2310 4435
rect 2314 4431 2315 4435
rect 2309 4430 2315 4431
rect 2309 4426 2310 4430
rect 2314 4426 2315 4430
rect 2309 4425 2315 4426
rect 2309 4421 2310 4425
rect 2314 4421 2315 4425
rect 2309 4420 2315 4421
rect 2309 4416 2310 4420
rect 2314 4416 2315 4420
rect 2309 4415 2315 4416
rect 2309 4411 2310 4415
rect 2314 4411 2315 4415
rect 2309 4410 2315 4411
rect 2309 4406 2310 4410
rect 2314 4406 2315 4410
rect 2309 4405 2315 4406
rect 2309 4401 2310 4405
rect 2314 4401 2315 4405
rect 2309 4400 2315 4401
rect 2309 4396 2310 4400
rect 2314 4396 2315 4400
rect 2309 4395 2315 4396
rect 2309 4391 2310 4395
rect 2314 4391 2315 4395
rect 2309 4390 2315 4391
rect 2309 4386 2310 4390
rect 2314 4386 2315 4390
rect 2309 4385 2315 4386
rect 2309 4381 2310 4385
rect 2314 4381 2315 4385
rect 2309 4380 2315 4381
rect 2309 4376 2310 4380
rect 2314 4376 2315 4380
rect 2309 4375 2315 4376
rect 2309 4371 2310 4375
rect 2314 4371 2315 4375
rect 2309 4370 2315 4371
rect 2309 4366 2310 4370
rect 2314 4366 2315 4370
rect 2309 4365 2315 4366
rect 2309 4361 2310 4365
rect 2314 4361 2315 4365
rect 2309 4360 2315 4361
rect 2309 4356 2310 4360
rect 2314 4356 2315 4360
rect 2309 4355 2315 4356
rect 2309 4351 2310 4355
rect 2314 4351 2315 4355
rect 2309 4350 2315 4351
rect 2309 4346 2310 4350
rect 2314 4346 2315 4350
rect 2399 4461 2400 4465
rect 2404 4461 2405 4465
rect 2399 4460 2405 4461
rect 2399 4456 2400 4460
rect 2404 4456 2405 4460
rect 2399 4455 2405 4456
rect 2399 4451 2400 4455
rect 2404 4451 2405 4455
rect 2399 4450 2405 4451
rect 2399 4446 2400 4450
rect 2404 4446 2405 4450
rect 2399 4445 2405 4446
rect 2399 4441 2400 4445
rect 2404 4441 2405 4445
rect 2399 4440 2405 4441
rect 2399 4436 2400 4440
rect 2404 4436 2405 4440
rect 2399 4435 2405 4436
rect 2399 4431 2400 4435
rect 2404 4431 2405 4435
rect 2399 4430 2405 4431
rect 2399 4426 2400 4430
rect 2404 4426 2405 4430
rect 2399 4425 2405 4426
rect 2399 4421 2400 4425
rect 2404 4421 2405 4425
rect 2399 4420 2405 4421
rect 2399 4416 2400 4420
rect 2404 4416 2405 4420
rect 2399 4415 2405 4416
rect 2399 4411 2400 4415
rect 2404 4411 2405 4415
rect 2399 4410 2405 4411
rect 2399 4406 2400 4410
rect 2404 4406 2405 4410
rect 2399 4405 2405 4406
rect 2399 4401 2400 4405
rect 2404 4401 2405 4405
rect 2399 4400 2405 4401
rect 2399 4396 2400 4400
rect 2404 4396 2405 4400
rect 2399 4395 2405 4396
rect 2399 4391 2400 4395
rect 2404 4391 2405 4395
rect 2399 4390 2405 4391
rect 2399 4386 2400 4390
rect 2404 4386 2405 4390
rect 2399 4385 2405 4386
rect 2399 4381 2400 4385
rect 2404 4381 2405 4385
rect 2399 4380 2405 4381
rect 2399 4376 2400 4380
rect 2404 4376 2405 4380
rect 2399 4375 2405 4376
rect 2399 4371 2400 4375
rect 2404 4371 2405 4375
rect 2399 4370 2405 4371
rect 2399 4366 2400 4370
rect 2404 4366 2405 4370
rect 2399 4365 2405 4366
rect 2399 4361 2400 4365
rect 2404 4361 2405 4365
rect 2399 4360 2405 4361
rect 2399 4356 2400 4360
rect 2404 4356 2405 4360
rect 2399 4355 2405 4356
rect 2399 4351 2400 4355
rect 2404 4351 2405 4355
rect 2399 4350 2405 4351
rect 2309 4345 2315 4346
rect 2309 4341 2310 4345
rect 2314 4341 2315 4345
rect 2399 4346 2400 4350
rect 2404 4346 2405 4350
rect 2399 4345 2405 4346
rect 2399 4341 2400 4345
rect 2404 4341 2405 4345
rect 2309 4340 2405 4341
rect 2309 4336 2310 4340
rect 2314 4336 2315 4340
rect 2319 4336 2320 4340
rect 2324 4336 2325 4340
rect 2329 4336 2330 4340
rect 2334 4336 2335 4340
rect 2339 4336 2340 4340
rect 2344 4336 2345 4340
rect 2349 4336 2350 4340
rect 2354 4336 2355 4340
rect 2359 4336 2360 4340
rect 2364 4336 2365 4340
rect 2369 4336 2370 4340
rect 2374 4336 2375 4340
rect 2379 4336 2380 4340
rect 2384 4336 2385 4340
rect 2389 4336 2390 4340
rect 2394 4336 2395 4340
rect 2399 4336 2400 4340
rect 2404 4336 2405 4340
rect 2309 4335 2405 4336
rect 2481 4462 2553 4464
rect 2481 4458 2483 4462
rect 2487 4458 2490 4462
rect 2494 4458 2495 4462
rect 2499 4458 2500 4462
rect 2504 4458 2505 4462
rect 2509 4458 2510 4462
rect 2514 4458 2515 4462
rect 2519 4458 2520 4462
rect 2524 4458 2525 4462
rect 2529 4458 2530 4462
rect 2534 4458 2535 4462
rect 2539 4458 2540 4462
rect 2544 4458 2547 4462
rect 2551 4458 2553 4462
rect 2481 4456 2553 4458
rect 2481 4455 2489 4456
rect 2481 4451 2483 4455
rect 2487 4451 2489 4455
rect 2481 4450 2489 4451
rect 2545 4455 2553 4456
rect 2545 4451 2547 4455
rect 2551 4451 2553 4455
rect 2545 4450 2553 4451
rect 2481 4446 2483 4450
rect 2487 4446 2489 4450
rect 2481 4445 2489 4446
rect 2481 4441 2483 4445
rect 2487 4441 2489 4445
rect 2481 4440 2489 4441
rect 2481 4436 2483 4440
rect 2487 4436 2489 4440
rect 2481 4435 2489 4436
rect 2481 4431 2483 4435
rect 2487 4431 2489 4435
rect 2481 4430 2489 4431
rect 2481 4426 2483 4430
rect 2487 4426 2489 4430
rect 2481 4425 2489 4426
rect 2481 4421 2483 4425
rect 2487 4421 2489 4425
rect 2481 4420 2489 4421
rect 2481 4416 2483 4420
rect 2487 4416 2489 4420
rect 2481 4415 2489 4416
rect 2481 4411 2483 4415
rect 2487 4411 2489 4415
rect 2481 4410 2489 4411
rect 2481 4406 2483 4410
rect 2487 4406 2489 4410
rect 2481 4405 2489 4406
rect 2481 4401 2483 4405
rect 2487 4401 2489 4405
rect 2481 4400 2489 4401
rect 2481 4396 2483 4400
rect 2487 4396 2489 4400
rect 2481 4395 2489 4396
rect 2481 4391 2483 4395
rect 2487 4391 2489 4395
rect 2481 4390 2489 4391
rect 2481 4386 2483 4390
rect 2487 4386 2489 4390
rect 2481 4385 2489 4386
rect 2481 4381 2483 4385
rect 2487 4381 2489 4385
rect 2481 4380 2489 4381
rect 2481 4376 2483 4380
rect 2487 4376 2489 4380
rect 2481 4375 2489 4376
rect 2481 4371 2483 4375
rect 2487 4371 2489 4375
rect 2481 4370 2489 4371
rect 2481 4366 2483 4370
rect 2487 4366 2489 4370
rect 2481 4365 2489 4366
rect 2481 4361 2483 4365
rect 2487 4361 2489 4365
rect 2545 4446 2547 4450
rect 2551 4446 2553 4450
rect 2545 4445 2553 4446
rect 2545 4441 2547 4445
rect 2551 4441 2553 4445
rect 2545 4440 2553 4441
rect 2545 4436 2547 4440
rect 2551 4436 2553 4440
rect 2545 4435 2553 4436
rect 2545 4431 2547 4435
rect 2551 4431 2553 4435
rect 2545 4430 2553 4431
rect 2545 4426 2547 4430
rect 2551 4426 2553 4430
rect 2545 4425 2553 4426
rect 2545 4421 2547 4425
rect 2551 4421 2553 4425
rect 2545 4420 2553 4421
rect 2545 4416 2547 4420
rect 2551 4416 2553 4420
rect 2545 4415 2553 4416
rect 2545 4411 2547 4415
rect 2551 4411 2553 4415
rect 2545 4410 2553 4411
rect 2545 4406 2547 4410
rect 2551 4406 2553 4410
rect 2545 4405 2553 4406
rect 2545 4401 2547 4405
rect 2551 4401 2553 4405
rect 2545 4400 2553 4401
rect 2545 4396 2547 4400
rect 2551 4396 2553 4400
rect 2545 4395 2553 4396
rect 2545 4391 2547 4395
rect 2551 4391 2553 4395
rect 2545 4390 2553 4391
rect 2545 4386 2547 4390
rect 2551 4386 2553 4390
rect 2545 4385 2553 4386
rect 2545 4381 2547 4385
rect 2551 4381 2553 4385
rect 2545 4380 2553 4381
rect 2545 4376 2547 4380
rect 2551 4376 2553 4380
rect 2545 4375 2553 4376
rect 2545 4371 2547 4375
rect 2551 4371 2553 4375
rect 2545 4370 2553 4371
rect 2545 4366 2547 4370
rect 2551 4366 2553 4370
rect 2545 4365 2553 4366
rect 2545 4361 2547 4365
rect 2551 4361 2553 4365
rect 2481 4360 2489 4361
rect 2481 4356 2483 4360
rect 2487 4356 2489 4360
rect 2481 4355 2489 4356
rect 2545 4360 2553 4361
rect 2545 4356 2547 4360
rect 2551 4356 2553 4360
rect 2545 4355 2553 4356
rect 2481 4353 2553 4355
rect 2481 4349 2483 4353
rect 2487 4349 2490 4353
rect 2494 4349 2495 4353
rect 2499 4349 2500 4353
rect 2504 4349 2505 4353
rect 2509 4349 2510 4353
rect 2514 4349 2515 4353
rect 2519 4349 2520 4353
rect 2524 4349 2525 4353
rect 2529 4349 2530 4353
rect 2534 4349 2535 4353
rect 2539 4349 2540 4353
rect 2544 4349 2547 4353
rect 2551 4349 2553 4353
rect 2481 4347 2553 4349
rect 2618 4475 2714 4476
rect 2618 4471 2619 4475
rect 2623 4471 2624 4475
rect 2628 4471 2629 4475
rect 2633 4471 2634 4475
rect 2638 4471 2639 4475
rect 2643 4471 2644 4475
rect 2648 4471 2649 4475
rect 2653 4471 2654 4475
rect 2658 4471 2659 4475
rect 2663 4471 2664 4475
rect 2668 4471 2669 4475
rect 2673 4471 2674 4475
rect 2678 4471 2679 4475
rect 2683 4471 2684 4475
rect 2688 4471 2689 4475
rect 2693 4471 2694 4475
rect 2698 4471 2699 4475
rect 2703 4471 2704 4475
rect 2708 4471 2709 4475
rect 2713 4471 2714 4475
rect 2618 4470 2714 4471
rect 2618 4466 2619 4470
rect 2623 4466 2624 4470
rect 2618 4465 2624 4466
rect 2618 4461 2619 4465
rect 2623 4461 2624 4465
rect 2708 4466 2709 4470
rect 2713 4466 2714 4470
rect 2708 4465 2714 4466
rect 2618 4460 2624 4461
rect 2618 4456 2619 4460
rect 2623 4456 2624 4460
rect 2618 4455 2624 4456
rect 2618 4451 2619 4455
rect 2623 4451 2624 4455
rect 2618 4450 2624 4451
rect 2618 4446 2619 4450
rect 2623 4446 2624 4450
rect 2618 4445 2624 4446
rect 2618 4441 2619 4445
rect 2623 4441 2624 4445
rect 2618 4440 2624 4441
rect 2618 4436 2619 4440
rect 2623 4436 2624 4440
rect 2618 4435 2624 4436
rect 2618 4431 2619 4435
rect 2623 4431 2624 4435
rect 2618 4430 2624 4431
rect 2618 4426 2619 4430
rect 2623 4426 2624 4430
rect 2618 4425 2624 4426
rect 2618 4421 2619 4425
rect 2623 4421 2624 4425
rect 2618 4420 2624 4421
rect 2618 4416 2619 4420
rect 2623 4416 2624 4420
rect 2618 4415 2624 4416
rect 2618 4411 2619 4415
rect 2623 4411 2624 4415
rect 2618 4410 2624 4411
rect 2618 4406 2619 4410
rect 2623 4406 2624 4410
rect 2618 4405 2624 4406
rect 2618 4401 2619 4405
rect 2623 4401 2624 4405
rect 2618 4400 2624 4401
rect 2618 4396 2619 4400
rect 2623 4396 2624 4400
rect 2618 4395 2624 4396
rect 2618 4391 2619 4395
rect 2623 4391 2624 4395
rect 2618 4390 2624 4391
rect 2618 4386 2619 4390
rect 2623 4386 2624 4390
rect 2618 4385 2624 4386
rect 2618 4381 2619 4385
rect 2623 4381 2624 4385
rect 2618 4380 2624 4381
rect 2618 4376 2619 4380
rect 2623 4376 2624 4380
rect 2618 4375 2624 4376
rect 2618 4371 2619 4375
rect 2623 4371 2624 4375
rect 2618 4370 2624 4371
rect 2618 4366 2619 4370
rect 2623 4366 2624 4370
rect 2618 4365 2624 4366
rect 2618 4361 2619 4365
rect 2623 4361 2624 4365
rect 2618 4360 2624 4361
rect 2618 4356 2619 4360
rect 2623 4356 2624 4360
rect 2618 4355 2624 4356
rect 2618 4351 2619 4355
rect 2623 4351 2624 4355
rect 2618 4350 2624 4351
rect 2618 4346 2619 4350
rect 2623 4346 2624 4350
rect 2708 4461 2709 4465
rect 2713 4461 2714 4465
rect 2708 4460 2714 4461
rect 2708 4456 2709 4460
rect 2713 4456 2714 4460
rect 2708 4455 2714 4456
rect 2708 4451 2709 4455
rect 2713 4451 2714 4455
rect 2708 4450 2714 4451
rect 2708 4446 2709 4450
rect 2713 4446 2714 4450
rect 2708 4445 2714 4446
rect 2708 4441 2709 4445
rect 2713 4441 2714 4445
rect 2708 4440 2714 4441
rect 2708 4436 2709 4440
rect 2713 4436 2714 4440
rect 2708 4435 2714 4436
rect 2708 4431 2709 4435
rect 2713 4431 2714 4435
rect 2708 4430 2714 4431
rect 2708 4426 2709 4430
rect 2713 4426 2714 4430
rect 2708 4425 2714 4426
rect 2708 4421 2709 4425
rect 2713 4421 2714 4425
rect 2708 4420 2714 4421
rect 2708 4416 2709 4420
rect 2713 4416 2714 4420
rect 2708 4415 2714 4416
rect 2708 4411 2709 4415
rect 2713 4411 2714 4415
rect 2708 4410 2714 4411
rect 2708 4406 2709 4410
rect 2713 4406 2714 4410
rect 2708 4405 2714 4406
rect 2708 4401 2709 4405
rect 2713 4401 2714 4405
rect 2708 4400 2714 4401
rect 2708 4396 2709 4400
rect 2713 4396 2714 4400
rect 2708 4395 2714 4396
rect 2708 4391 2709 4395
rect 2713 4391 2714 4395
rect 2708 4390 2714 4391
rect 2708 4386 2709 4390
rect 2713 4386 2714 4390
rect 2708 4385 2714 4386
rect 2708 4381 2709 4385
rect 2713 4381 2714 4385
rect 2708 4380 2714 4381
rect 2708 4376 2709 4380
rect 2713 4376 2714 4380
rect 2708 4375 2714 4376
rect 2708 4371 2709 4375
rect 2713 4371 2714 4375
rect 2708 4370 2714 4371
rect 2708 4366 2709 4370
rect 2713 4366 2714 4370
rect 2708 4365 2714 4366
rect 2708 4361 2709 4365
rect 2713 4361 2714 4365
rect 2708 4360 2714 4361
rect 2708 4356 2709 4360
rect 2713 4356 2714 4360
rect 2708 4355 2714 4356
rect 2708 4351 2709 4355
rect 2713 4351 2714 4355
rect 2708 4350 2714 4351
rect 2618 4345 2624 4346
rect 2618 4341 2619 4345
rect 2623 4341 2624 4345
rect 2708 4346 2709 4350
rect 2713 4346 2714 4350
rect 2708 4345 2714 4346
rect 2708 4341 2709 4345
rect 2713 4341 2714 4345
rect 2618 4340 2714 4341
rect 2618 4336 2619 4340
rect 2623 4336 2624 4340
rect 2628 4336 2629 4340
rect 2633 4336 2634 4340
rect 2638 4336 2639 4340
rect 2643 4336 2644 4340
rect 2648 4336 2649 4340
rect 2653 4336 2654 4340
rect 2658 4336 2659 4340
rect 2663 4336 2664 4340
rect 2668 4336 2669 4340
rect 2673 4336 2674 4340
rect 2678 4336 2679 4340
rect 2683 4336 2684 4340
rect 2688 4336 2689 4340
rect 2693 4336 2694 4340
rect 2698 4336 2699 4340
rect 2703 4336 2704 4340
rect 2708 4336 2709 4340
rect 2713 4336 2714 4340
rect 2618 4335 2714 4336
rect 2790 4462 2862 4464
rect 2790 4458 2792 4462
rect 2796 4458 2799 4462
rect 2803 4458 2804 4462
rect 2808 4458 2809 4462
rect 2813 4458 2814 4462
rect 2818 4458 2819 4462
rect 2823 4458 2824 4462
rect 2828 4458 2829 4462
rect 2833 4458 2834 4462
rect 2838 4458 2839 4462
rect 2843 4458 2844 4462
rect 2848 4458 2849 4462
rect 2853 4458 2856 4462
rect 2860 4458 2862 4462
rect 2790 4456 2862 4458
rect 2790 4455 2798 4456
rect 2790 4451 2792 4455
rect 2796 4451 2798 4455
rect 2790 4450 2798 4451
rect 2854 4455 2862 4456
rect 2854 4451 2856 4455
rect 2860 4451 2862 4455
rect 2854 4450 2862 4451
rect 2790 4446 2792 4450
rect 2796 4446 2798 4450
rect 2790 4445 2798 4446
rect 2790 4441 2792 4445
rect 2796 4441 2798 4445
rect 2790 4440 2798 4441
rect 2790 4436 2792 4440
rect 2796 4436 2798 4440
rect 2790 4435 2798 4436
rect 2790 4431 2792 4435
rect 2796 4431 2798 4435
rect 2790 4430 2798 4431
rect 2790 4426 2792 4430
rect 2796 4426 2798 4430
rect 2790 4425 2798 4426
rect 2790 4421 2792 4425
rect 2796 4421 2798 4425
rect 2790 4420 2798 4421
rect 2790 4416 2792 4420
rect 2796 4416 2798 4420
rect 2790 4415 2798 4416
rect 2790 4411 2792 4415
rect 2796 4411 2798 4415
rect 2790 4410 2798 4411
rect 2790 4406 2792 4410
rect 2796 4406 2798 4410
rect 2790 4405 2798 4406
rect 2790 4401 2792 4405
rect 2796 4401 2798 4405
rect 2790 4400 2798 4401
rect 2790 4396 2792 4400
rect 2796 4396 2798 4400
rect 2790 4395 2798 4396
rect 2790 4391 2792 4395
rect 2796 4391 2798 4395
rect 2790 4390 2798 4391
rect 2790 4386 2792 4390
rect 2796 4386 2798 4390
rect 2790 4385 2798 4386
rect 2790 4381 2792 4385
rect 2796 4381 2798 4385
rect 2790 4380 2798 4381
rect 2790 4376 2792 4380
rect 2796 4376 2798 4380
rect 2790 4375 2798 4376
rect 2790 4371 2792 4375
rect 2796 4371 2798 4375
rect 2790 4370 2798 4371
rect 2790 4366 2792 4370
rect 2796 4366 2798 4370
rect 2790 4365 2798 4366
rect 2790 4361 2792 4365
rect 2796 4361 2798 4365
rect 2854 4446 2856 4450
rect 2860 4446 2862 4450
rect 2854 4445 2862 4446
rect 2854 4441 2856 4445
rect 2860 4441 2862 4445
rect 2854 4440 2862 4441
rect 2854 4436 2856 4440
rect 2860 4436 2862 4440
rect 2854 4435 2862 4436
rect 2854 4431 2856 4435
rect 2860 4431 2862 4435
rect 2854 4430 2862 4431
rect 2854 4426 2856 4430
rect 2860 4426 2862 4430
rect 2854 4425 2862 4426
rect 2854 4421 2856 4425
rect 2860 4421 2862 4425
rect 2854 4420 2862 4421
rect 2854 4416 2856 4420
rect 2860 4416 2862 4420
rect 2854 4415 2862 4416
rect 2854 4411 2856 4415
rect 2860 4411 2862 4415
rect 2854 4410 2862 4411
rect 2854 4406 2856 4410
rect 2860 4406 2862 4410
rect 2854 4405 2862 4406
rect 2854 4401 2856 4405
rect 2860 4401 2862 4405
rect 2854 4400 2862 4401
rect 2854 4396 2856 4400
rect 2860 4396 2862 4400
rect 2854 4395 2862 4396
rect 2854 4391 2856 4395
rect 2860 4391 2862 4395
rect 2854 4390 2862 4391
rect 2854 4386 2856 4390
rect 2860 4386 2862 4390
rect 2854 4385 2862 4386
rect 2854 4381 2856 4385
rect 2860 4381 2862 4385
rect 2854 4380 2862 4381
rect 2854 4376 2856 4380
rect 2860 4376 2862 4380
rect 2854 4375 2862 4376
rect 2854 4371 2856 4375
rect 2860 4371 2862 4375
rect 2854 4370 2862 4371
rect 2854 4366 2856 4370
rect 2860 4366 2862 4370
rect 2854 4365 2862 4366
rect 2854 4361 2856 4365
rect 2860 4361 2862 4365
rect 2790 4360 2798 4361
rect 2790 4356 2792 4360
rect 2796 4356 2798 4360
rect 2790 4355 2798 4356
rect 2854 4360 2862 4361
rect 2854 4356 2856 4360
rect 2860 4356 2862 4360
rect 2854 4355 2862 4356
rect 2790 4353 2862 4355
rect 2790 4349 2792 4353
rect 2796 4349 2799 4353
rect 2803 4349 2804 4353
rect 2808 4349 2809 4353
rect 2813 4349 2814 4353
rect 2818 4349 2819 4353
rect 2823 4349 2824 4353
rect 2828 4349 2829 4353
rect 2833 4349 2834 4353
rect 2838 4349 2839 4353
rect 2843 4349 2844 4353
rect 2848 4349 2849 4353
rect 2853 4349 2856 4353
rect 2860 4349 2862 4353
rect 2790 4347 2862 4349
rect 2927 4475 3023 4476
rect 2927 4471 2928 4475
rect 2932 4471 2933 4475
rect 2937 4471 2938 4475
rect 2942 4471 2943 4475
rect 2947 4471 2948 4475
rect 2952 4471 2953 4475
rect 2957 4471 2958 4475
rect 2962 4471 2963 4475
rect 2967 4471 2968 4475
rect 2972 4471 2973 4475
rect 2977 4471 2978 4475
rect 2982 4471 2983 4475
rect 2987 4471 2988 4475
rect 2992 4471 2993 4475
rect 2997 4471 2998 4475
rect 3002 4471 3003 4475
rect 3007 4471 3008 4475
rect 3012 4471 3013 4475
rect 3017 4471 3018 4475
rect 3022 4471 3023 4475
rect 2927 4470 3023 4471
rect 2927 4466 2928 4470
rect 2932 4466 2933 4470
rect 2927 4465 2933 4466
rect 2927 4461 2928 4465
rect 2932 4461 2933 4465
rect 3017 4466 3018 4470
rect 3022 4466 3023 4470
rect 3017 4465 3023 4466
rect 2927 4460 2933 4461
rect 2927 4456 2928 4460
rect 2932 4456 2933 4460
rect 2927 4455 2933 4456
rect 2927 4451 2928 4455
rect 2932 4451 2933 4455
rect 2927 4450 2933 4451
rect 2927 4446 2928 4450
rect 2932 4446 2933 4450
rect 2927 4445 2933 4446
rect 2927 4441 2928 4445
rect 2932 4441 2933 4445
rect 2927 4440 2933 4441
rect 2927 4436 2928 4440
rect 2932 4436 2933 4440
rect 2927 4435 2933 4436
rect 2927 4431 2928 4435
rect 2932 4431 2933 4435
rect 2927 4430 2933 4431
rect 2927 4426 2928 4430
rect 2932 4426 2933 4430
rect 2927 4425 2933 4426
rect 2927 4421 2928 4425
rect 2932 4421 2933 4425
rect 2927 4420 2933 4421
rect 2927 4416 2928 4420
rect 2932 4416 2933 4420
rect 2927 4415 2933 4416
rect 2927 4411 2928 4415
rect 2932 4411 2933 4415
rect 2927 4410 2933 4411
rect 2927 4406 2928 4410
rect 2932 4406 2933 4410
rect 2927 4405 2933 4406
rect 2927 4401 2928 4405
rect 2932 4401 2933 4405
rect 2927 4400 2933 4401
rect 2927 4396 2928 4400
rect 2932 4396 2933 4400
rect 2927 4395 2933 4396
rect 2927 4391 2928 4395
rect 2932 4391 2933 4395
rect 2927 4390 2933 4391
rect 2927 4386 2928 4390
rect 2932 4386 2933 4390
rect 2927 4385 2933 4386
rect 2927 4381 2928 4385
rect 2932 4381 2933 4385
rect 2927 4380 2933 4381
rect 2927 4376 2928 4380
rect 2932 4376 2933 4380
rect 2927 4375 2933 4376
rect 2927 4371 2928 4375
rect 2932 4371 2933 4375
rect 2927 4370 2933 4371
rect 2927 4366 2928 4370
rect 2932 4366 2933 4370
rect 2927 4365 2933 4366
rect 2927 4361 2928 4365
rect 2932 4361 2933 4365
rect 2927 4360 2933 4361
rect 2927 4356 2928 4360
rect 2932 4356 2933 4360
rect 2927 4355 2933 4356
rect 2927 4351 2928 4355
rect 2932 4351 2933 4355
rect 2927 4350 2933 4351
rect 2927 4346 2928 4350
rect 2932 4346 2933 4350
rect 3017 4461 3018 4465
rect 3022 4461 3023 4465
rect 3017 4460 3023 4461
rect 3017 4456 3018 4460
rect 3022 4456 3023 4460
rect 3017 4455 3023 4456
rect 3017 4451 3018 4455
rect 3022 4451 3023 4455
rect 3017 4450 3023 4451
rect 3017 4446 3018 4450
rect 3022 4446 3023 4450
rect 3017 4445 3023 4446
rect 3017 4441 3018 4445
rect 3022 4441 3023 4445
rect 3017 4440 3023 4441
rect 3017 4436 3018 4440
rect 3022 4436 3023 4440
rect 3017 4435 3023 4436
rect 3017 4431 3018 4435
rect 3022 4431 3023 4435
rect 3017 4430 3023 4431
rect 3017 4426 3018 4430
rect 3022 4426 3023 4430
rect 3017 4425 3023 4426
rect 3017 4421 3018 4425
rect 3022 4421 3023 4425
rect 3017 4420 3023 4421
rect 3017 4416 3018 4420
rect 3022 4416 3023 4420
rect 3017 4415 3023 4416
rect 3017 4411 3018 4415
rect 3022 4411 3023 4415
rect 3017 4410 3023 4411
rect 3017 4406 3018 4410
rect 3022 4406 3023 4410
rect 3017 4405 3023 4406
rect 3017 4401 3018 4405
rect 3022 4401 3023 4405
rect 3017 4400 3023 4401
rect 3017 4396 3018 4400
rect 3022 4396 3023 4400
rect 3017 4395 3023 4396
rect 3017 4391 3018 4395
rect 3022 4391 3023 4395
rect 3017 4390 3023 4391
rect 3017 4386 3018 4390
rect 3022 4386 3023 4390
rect 3017 4385 3023 4386
rect 3017 4381 3018 4385
rect 3022 4381 3023 4385
rect 3017 4380 3023 4381
rect 3017 4376 3018 4380
rect 3022 4376 3023 4380
rect 3017 4375 3023 4376
rect 3017 4371 3018 4375
rect 3022 4371 3023 4375
rect 3017 4370 3023 4371
rect 3017 4366 3018 4370
rect 3022 4366 3023 4370
rect 3017 4365 3023 4366
rect 3017 4361 3018 4365
rect 3022 4361 3023 4365
rect 3017 4360 3023 4361
rect 3017 4356 3018 4360
rect 3022 4356 3023 4360
rect 3017 4355 3023 4356
rect 3017 4351 3018 4355
rect 3022 4351 3023 4355
rect 3017 4350 3023 4351
rect 2927 4345 2933 4346
rect 2927 4341 2928 4345
rect 2932 4341 2933 4345
rect 3017 4346 3018 4350
rect 3022 4346 3023 4350
rect 3017 4345 3023 4346
rect 3017 4341 3018 4345
rect 3022 4341 3023 4345
rect 2927 4340 3023 4341
rect 2927 4336 2928 4340
rect 2932 4336 2933 4340
rect 2937 4336 2938 4340
rect 2942 4336 2943 4340
rect 2947 4336 2948 4340
rect 2952 4336 2953 4340
rect 2957 4336 2958 4340
rect 2962 4336 2963 4340
rect 2967 4336 2968 4340
rect 2972 4336 2973 4340
rect 2977 4336 2978 4340
rect 2982 4336 2983 4340
rect 2987 4336 2988 4340
rect 2992 4336 2993 4340
rect 2997 4336 2998 4340
rect 3002 4336 3003 4340
rect 3007 4336 3008 4340
rect 3012 4336 3013 4340
rect 3017 4336 3018 4340
rect 3022 4336 3023 4340
rect 2927 4335 3023 4336
rect 3099 4462 3171 4464
rect 3099 4458 3101 4462
rect 3105 4458 3108 4462
rect 3112 4458 3113 4462
rect 3117 4458 3118 4462
rect 3122 4458 3123 4462
rect 3127 4458 3128 4462
rect 3132 4458 3133 4462
rect 3137 4458 3138 4462
rect 3142 4458 3143 4462
rect 3147 4458 3148 4462
rect 3152 4458 3153 4462
rect 3157 4458 3158 4462
rect 3162 4458 3165 4462
rect 3169 4458 3171 4462
rect 3099 4456 3171 4458
rect 3099 4455 3107 4456
rect 3099 4451 3101 4455
rect 3105 4451 3107 4455
rect 3099 4450 3107 4451
rect 3163 4455 3171 4456
rect 3163 4451 3165 4455
rect 3169 4451 3171 4455
rect 3163 4450 3171 4451
rect 3099 4446 3101 4450
rect 3105 4446 3107 4450
rect 3099 4445 3107 4446
rect 3099 4441 3101 4445
rect 3105 4441 3107 4445
rect 3099 4440 3107 4441
rect 3099 4436 3101 4440
rect 3105 4436 3107 4440
rect 3099 4435 3107 4436
rect 3099 4431 3101 4435
rect 3105 4431 3107 4435
rect 3099 4430 3107 4431
rect 3099 4426 3101 4430
rect 3105 4426 3107 4430
rect 3099 4425 3107 4426
rect 3099 4421 3101 4425
rect 3105 4421 3107 4425
rect 3099 4420 3107 4421
rect 3099 4416 3101 4420
rect 3105 4416 3107 4420
rect 3099 4415 3107 4416
rect 3099 4411 3101 4415
rect 3105 4411 3107 4415
rect 3099 4410 3107 4411
rect 3099 4406 3101 4410
rect 3105 4406 3107 4410
rect 3099 4405 3107 4406
rect 3099 4401 3101 4405
rect 3105 4401 3107 4405
rect 3099 4400 3107 4401
rect 3099 4396 3101 4400
rect 3105 4396 3107 4400
rect 3099 4395 3107 4396
rect 3099 4391 3101 4395
rect 3105 4391 3107 4395
rect 3099 4390 3107 4391
rect 3099 4386 3101 4390
rect 3105 4386 3107 4390
rect 3099 4385 3107 4386
rect 3099 4381 3101 4385
rect 3105 4381 3107 4385
rect 3099 4380 3107 4381
rect 3099 4376 3101 4380
rect 3105 4376 3107 4380
rect 3099 4375 3107 4376
rect 3099 4371 3101 4375
rect 3105 4371 3107 4375
rect 3099 4370 3107 4371
rect 3099 4366 3101 4370
rect 3105 4366 3107 4370
rect 3099 4365 3107 4366
rect 3099 4361 3101 4365
rect 3105 4361 3107 4365
rect 3163 4446 3165 4450
rect 3169 4446 3171 4450
rect 3163 4445 3171 4446
rect 3163 4441 3165 4445
rect 3169 4441 3171 4445
rect 3163 4440 3171 4441
rect 3163 4436 3165 4440
rect 3169 4436 3171 4440
rect 3163 4435 3171 4436
rect 3163 4431 3165 4435
rect 3169 4431 3171 4435
rect 3163 4430 3171 4431
rect 3163 4426 3165 4430
rect 3169 4426 3171 4430
rect 3163 4425 3171 4426
rect 3163 4421 3165 4425
rect 3169 4421 3171 4425
rect 3163 4420 3171 4421
rect 3163 4416 3165 4420
rect 3169 4416 3171 4420
rect 3163 4415 3171 4416
rect 3163 4411 3165 4415
rect 3169 4411 3171 4415
rect 3163 4410 3171 4411
rect 3163 4406 3165 4410
rect 3169 4406 3171 4410
rect 3163 4405 3171 4406
rect 3163 4401 3165 4405
rect 3169 4401 3171 4405
rect 3163 4400 3171 4401
rect 3163 4396 3165 4400
rect 3169 4396 3171 4400
rect 3163 4395 3171 4396
rect 3163 4391 3165 4395
rect 3169 4391 3171 4395
rect 3163 4390 3171 4391
rect 3163 4386 3165 4390
rect 3169 4386 3171 4390
rect 3163 4385 3171 4386
rect 3163 4381 3165 4385
rect 3169 4381 3171 4385
rect 3163 4380 3171 4381
rect 3163 4376 3165 4380
rect 3169 4376 3171 4380
rect 3163 4375 3171 4376
rect 3163 4371 3165 4375
rect 3169 4371 3171 4375
rect 3163 4370 3171 4371
rect 3163 4366 3165 4370
rect 3169 4366 3171 4370
rect 3163 4365 3171 4366
rect 3163 4361 3165 4365
rect 3169 4361 3171 4365
rect 3099 4360 3107 4361
rect 3099 4356 3101 4360
rect 3105 4356 3107 4360
rect 3099 4355 3107 4356
rect 3163 4360 3171 4361
rect 3163 4356 3165 4360
rect 3169 4356 3171 4360
rect 3163 4355 3171 4356
rect 3099 4353 3171 4355
rect 3099 4349 3101 4353
rect 3105 4349 3108 4353
rect 3112 4349 3113 4353
rect 3117 4349 3118 4353
rect 3122 4349 3123 4353
rect 3127 4349 3128 4353
rect 3132 4349 3133 4353
rect 3137 4349 3138 4353
rect 3142 4349 3143 4353
rect 3147 4349 3148 4353
rect 3152 4349 3153 4353
rect 3157 4349 3158 4353
rect 3162 4349 3165 4353
rect 3169 4349 3171 4353
rect 3099 4347 3171 4349
rect 3236 4475 3332 4476
rect 3236 4471 3237 4475
rect 3241 4471 3242 4475
rect 3246 4471 3247 4475
rect 3251 4471 3252 4475
rect 3256 4471 3257 4475
rect 3261 4471 3262 4475
rect 3266 4471 3267 4475
rect 3271 4471 3272 4475
rect 3276 4471 3277 4475
rect 3281 4471 3282 4475
rect 3286 4471 3287 4475
rect 3291 4471 3292 4475
rect 3296 4471 3297 4475
rect 3301 4471 3302 4475
rect 3306 4471 3307 4475
rect 3311 4471 3312 4475
rect 3316 4471 3317 4475
rect 3321 4471 3322 4475
rect 3326 4471 3327 4475
rect 3331 4471 3332 4475
rect 3236 4470 3332 4471
rect 3236 4466 3237 4470
rect 3241 4466 3242 4470
rect 3236 4465 3242 4466
rect 3236 4461 3237 4465
rect 3241 4461 3242 4465
rect 3326 4466 3327 4470
rect 3331 4466 3332 4470
rect 3326 4465 3332 4466
rect 3236 4460 3242 4461
rect 3236 4456 3237 4460
rect 3241 4456 3242 4460
rect 3236 4455 3242 4456
rect 3236 4451 3237 4455
rect 3241 4451 3242 4455
rect 3236 4450 3242 4451
rect 3236 4446 3237 4450
rect 3241 4446 3242 4450
rect 3236 4445 3242 4446
rect 3236 4441 3237 4445
rect 3241 4441 3242 4445
rect 3236 4440 3242 4441
rect 3236 4436 3237 4440
rect 3241 4436 3242 4440
rect 3236 4435 3242 4436
rect 3236 4431 3237 4435
rect 3241 4431 3242 4435
rect 3236 4430 3242 4431
rect 3236 4426 3237 4430
rect 3241 4426 3242 4430
rect 3236 4425 3242 4426
rect 3236 4421 3237 4425
rect 3241 4421 3242 4425
rect 3236 4420 3242 4421
rect 3236 4416 3237 4420
rect 3241 4416 3242 4420
rect 3236 4415 3242 4416
rect 3236 4411 3237 4415
rect 3241 4411 3242 4415
rect 3236 4410 3242 4411
rect 3236 4406 3237 4410
rect 3241 4406 3242 4410
rect 3236 4405 3242 4406
rect 3236 4401 3237 4405
rect 3241 4401 3242 4405
rect 3236 4400 3242 4401
rect 3236 4396 3237 4400
rect 3241 4396 3242 4400
rect 3236 4395 3242 4396
rect 3236 4391 3237 4395
rect 3241 4391 3242 4395
rect 3236 4390 3242 4391
rect 3236 4386 3237 4390
rect 3241 4386 3242 4390
rect 3236 4385 3242 4386
rect 3236 4381 3237 4385
rect 3241 4381 3242 4385
rect 3236 4380 3242 4381
rect 3236 4376 3237 4380
rect 3241 4376 3242 4380
rect 3236 4375 3242 4376
rect 3236 4371 3237 4375
rect 3241 4371 3242 4375
rect 3236 4370 3242 4371
rect 3236 4366 3237 4370
rect 3241 4366 3242 4370
rect 3236 4365 3242 4366
rect 3236 4361 3237 4365
rect 3241 4361 3242 4365
rect 3236 4360 3242 4361
rect 3236 4356 3237 4360
rect 3241 4356 3242 4360
rect 3236 4355 3242 4356
rect 3236 4351 3237 4355
rect 3241 4351 3242 4355
rect 3236 4350 3242 4351
rect 3236 4346 3237 4350
rect 3241 4346 3242 4350
rect 3326 4461 3327 4465
rect 3331 4461 3332 4465
rect 3326 4460 3332 4461
rect 3326 4456 3327 4460
rect 3331 4456 3332 4460
rect 3326 4455 3332 4456
rect 3326 4451 3327 4455
rect 3331 4451 3332 4455
rect 3326 4450 3332 4451
rect 3326 4446 3327 4450
rect 3331 4446 3332 4450
rect 3326 4445 3332 4446
rect 3326 4441 3327 4445
rect 3331 4441 3332 4445
rect 3326 4440 3332 4441
rect 3326 4436 3327 4440
rect 3331 4436 3332 4440
rect 3326 4435 3332 4436
rect 3326 4431 3327 4435
rect 3331 4431 3332 4435
rect 3326 4430 3332 4431
rect 3326 4426 3327 4430
rect 3331 4426 3332 4430
rect 3326 4425 3332 4426
rect 3326 4421 3327 4425
rect 3331 4421 3332 4425
rect 3326 4420 3332 4421
rect 3326 4416 3327 4420
rect 3331 4416 3332 4420
rect 3326 4415 3332 4416
rect 3326 4411 3327 4415
rect 3331 4411 3332 4415
rect 3326 4410 3332 4411
rect 3326 4406 3327 4410
rect 3331 4406 3332 4410
rect 3326 4405 3332 4406
rect 3326 4401 3327 4405
rect 3331 4401 3332 4405
rect 3326 4400 3332 4401
rect 3326 4396 3327 4400
rect 3331 4396 3332 4400
rect 3326 4395 3332 4396
rect 3326 4391 3327 4395
rect 3331 4391 3332 4395
rect 3326 4390 3332 4391
rect 3326 4386 3327 4390
rect 3331 4386 3332 4390
rect 3326 4385 3332 4386
rect 3326 4381 3327 4385
rect 3331 4381 3332 4385
rect 3326 4380 3332 4381
rect 3326 4376 3327 4380
rect 3331 4376 3332 4380
rect 3326 4375 3332 4376
rect 3326 4371 3327 4375
rect 3331 4371 3332 4375
rect 3326 4370 3332 4371
rect 3326 4366 3327 4370
rect 3331 4366 3332 4370
rect 3326 4365 3332 4366
rect 3326 4361 3327 4365
rect 3331 4361 3332 4365
rect 3326 4360 3332 4361
rect 3326 4356 3327 4360
rect 3331 4356 3332 4360
rect 3326 4355 3332 4356
rect 3326 4351 3327 4355
rect 3331 4351 3332 4355
rect 3326 4350 3332 4351
rect 3236 4345 3242 4346
rect 3236 4341 3237 4345
rect 3241 4341 3242 4345
rect 3326 4346 3327 4350
rect 3331 4346 3332 4350
rect 3326 4345 3332 4346
rect 3326 4341 3327 4345
rect 3331 4341 3332 4345
rect 3236 4340 3332 4341
rect 3236 4336 3237 4340
rect 3241 4336 3242 4340
rect 3246 4336 3247 4340
rect 3251 4336 3252 4340
rect 3256 4336 3257 4340
rect 3261 4336 3262 4340
rect 3266 4336 3267 4340
rect 3271 4336 3272 4340
rect 3276 4336 3277 4340
rect 3281 4336 3282 4340
rect 3286 4336 3287 4340
rect 3291 4336 3292 4340
rect 3296 4336 3297 4340
rect 3301 4336 3302 4340
rect 3306 4336 3307 4340
rect 3311 4336 3312 4340
rect 3316 4336 3317 4340
rect 3321 4336 3322 4340
rect 3326 4336 3327 4340
rect 3331 4336 3332 4340
rect 3236 4335 3332 4336
rect 3408 4462 3480 4464
rect 3408 4458 3410 4462
rect 3414 4458 3417 4462
rect 3421 4458 3422 4462
rect 3426 4458 3427 4462
rect 3431 4458 3432 4462
rect 3436 4458 3437 4462
rect 3441 4458 3442 4462
rect 3446 4458 3447 4462
rect 3451 4458 3452 4462
rect 3456 4458 3457 4462
rect 3461 4458 3462 4462
rect 3466 4458 3467 4462
rect 3471 4458 3474 4462
rect 3478 4458 3480 4462
rect 3408 4456 3480 4458
rect 3408 4455 3416 4456
rect 3408 4451 3410 4455
rect 3414 4451 3416 4455
rect 3408 4450 3416 4451
rect 3472 4455 3480 4456
rect 3472 4451 3474 4455
rect 3478 4451 3480 4455
rect 3472 4450 3480 4451
rect 3408 4446 3410 4450
rect 3414 4446 3416 4450
rect 3408 4445 3416 4446
rect 3408 4441 3410 4445
rect 3414 4441 3416 4445
rect 3408 4440 3416 4441
rect 3408 4436 3410 4440
rect 3414 4436 3416 4440
rect 3408 4435 3416 4436
rect 3408 4431 3410 4435
rect 3414 4431 3416 4435
rect 3408 4430 3416 4431
rect 3408 4426 3410 4430
rect 3414 4426 3416 4430
rect 3408 4425 3416 4426
rect 3408 4421 3410 4425
rect 3414 4421 3416 4425
rect 3408 4420 3416 4421
rect 3408 4416 3410 4420
rect 3414 4416 3416 4420
rect 3408 4415 3416 4416
rect 3408 4411 3410 4415
rect 3414 4411 3416 4415
rect 3408 4410 3416 4411
rect 3408 4406 3410 4410
rect 3414 4406 3416 4410
rect 3408 4405 3416 4406
rect 3408 4401 3410 4405
rect 3414 4401 3416 4405
rect 3408 4400 3416 4401
rect 3408 4396 3410 4400
rect 3414 4396 3416 4400
rect 3408 4395 3416 4396
rect 3408 4391 3410 4395
rect 3414 4391 3416 4395
rect 3408 4390 3416 4391
rect 3408 4386 3410 4390
rect 3414 4386 3416 4390
rect 3408 4385 3416 4386
rect 3408 4381 3410 4385
rect 3414 4381 3416 4385
rect 3408 4380 3416 4381
rect 3408 4376 3410 4380
rect 3414 4376 3416 4380
rect 3408 4375 3416 4376
rect 3408 4371 3410 4375
rect 3414 4371 3416 4375
rect 3408 4370 3416 4371
rect 3408 4366 3410 4370
rect 3414 4366 3416 4370
rect 3408 4365 3416 4366
rect 3408 4361 3410 4365
rect 3414 4361 3416 4365
rect 3472 4446 3474 4450
rect 3478 4446 3480 4450
rect 3472 4445 3480 4446
rect 3472 4441 3474 4445
rect 3478 4441 3480 4445
rect 3472 4440 3480 4441
rect 3472 4436 3474 4440
rect 3478 4436 3480 4440
rect 3472 4435 3480 4436
rect 3472 4431 3474 4435
rect 3478 4431 3480 4435
rect 3472 4430 3480 4431
rect 3472 4426 3474 4430
rect 3478 4426 3480 4430
rect 3472 4425 3480 4426
rect 3472 4421 3474 4425
rect 3478 4421 3480 4425
rect 3472 4420 3480 4421
rect 3472 4416 3474 4420
rect 3478 4416 3480 4420
rect 3472 4415 3480 4416
rect 3472 4411 3474 4415
rect 3478 4411 3480 4415
rect 3472 4410 3480 4411
rect 3472 4406 3474 4410
rect 3478 4406 3480 4410
rect 3472 4405 3480 4406
rect 3472 4401 3474 4405
rect 3478 4401 3480 4405
rect 3472 4400 3480 4401
rect 3472 4396 3474 4400
rect 3478 4396 3480 4400
rect 3472 4395 3480 4396
rect 3472 4391 3474 4395
rect 3478 4391 3480 4395
rect 3472 4390 3480 4391
rect 3472 4386 3474 4390
rect 3478 4386 3480 4390
rect 3472 4385 3480 4386
rect 3472 4381 3474 4385
rect 3478 4381 3480 4385
rect 3472 4380 3480 4381
rect 3472 4376 3474 4380
rect 3478 4376 3480 4380
rect 3472 4375 3480 4376
rect 3472 4371 3474 4375
rect 3478 4371 3480 4375
rect 3472 4370 3480 4371
rect 3472 4366 3474 4370
rect 3478 4366 3480 4370
rect 3472 4365 3480 4366
rect 3472 4361 3474 4365
rect 3478 4361 3480 4365
rect 3408 4360 3416 4361
rect 3408 4356 3410 4360
rect 3414 4356 3416 4360
rect 3408 4355 3416 4356
rect 3472 4360 3480 4361
rect 3472 4356 3474 4360
rect 3478 4356 3480 4360
rect 3472 4355 3480 4356
rect 3408 4353 3480 4355
rect 3408 4349 3410 4353
rect 3414 4349 3417 4353
rect 3421 4349 3422 4353
rect 3426 4349 3427 4353
rect 3431 4349 3432 4353
rect 3436 4349 3437 4353
rect 3441 4349 3442 4353
rect 3446 4349 3447 4353
rect 3451 4349 3452 4353
rect 3456 4349 3457 4353
rect 3461 4349 3462 4353
rect 3466 4349 3467 4353
rect 3471 4349 3474 4353
rect 3478 4349 3480 4353
rect 3408 4347 3480 4349
rect 3545 4475 3641 4476
rect 3545 4471 3546 4475
rect 3550 4471 3551 4475
rect 3555 4471 3556 4475
rect 3560 4471 3561 4475
rect 3565 4471 3566 4475
rect 3570 4471 3571 4475
rect 3575 4471 3576 4475
rect 3580 4471 3581 4475
rect 3585 4471 3586 4475
rect 3590 4471 3591 4475
rect 3595 4471 3596 4475
rect 3600 4471 3601 4475
rect 3605 4471 3606 4475
rect 3610 4471 3611 4475
rect 3615 4471 3616 4475
rect 3620 4471 3621 4475
rect 3625 4471 3626 4475
rect 3630 4471 3631 4475
rect 3635 4471 3636 4475
rect 3640 4471 3641 4475
rect 3545 4470 3641 4471
rect 3545 4466 3546 4470
rect 3550 4466 3551 4470
rect 3545 4465 3551 4466
rect 3545 4461 3546 4465
rect 3550 4461 3551 4465
rect 3635 4466 3636 4470
rect 3640 4466 3641 4470
rect 3635 4465 3641 4466
rect 3545 4460 3551 4461
rect 3545 4456 3546 4460
rect 3550 4456 3551 4460
rect 3545 4455 3551 4456
rect 3545 4451 3546 4455
rect 3550 4451 3551 4455
rect 3545 4450 3551 4451
rect 3545 4446 3546 4450
rect 3550 4446 3551 4450
rect 3545 4445 3551 4446
rect 3545 4441 3546 4445
rect 3550 4441 3551 4445
rect 3545 4440 3551 4441
rect 3545 4436 3546 4440
rect 3550 4436 3551 4440
rect 3545 4435 3551 4436
rect 3545 4431 3546 4435
rect 3550 4431 3551 4435
rect 3545 4430 3551 4431
rect 3545 4426 3546 4430
rect 3550 4426 3551 4430
rect 3545 4425 3551 4426
rect 3545 4421 3546 4425
rect 3550 4421 3551 4425
rect 3545 4420 3551 4421
rect 3545 4416 3546 4420
rect 3550 4416 3551 4420
rect 3545 4415 3551 4416
rect 3545 4411 3546 4415
rect 3550 4411 3551 4415
rect 3545 4410 3551 4411
rect 3545 4406 3546 4410
rect 3550 4406 3551 4410
rect 3545 4405 3551 4406
rect 3545 4401 3546 4405
rect 3550 4401 3551 4405
rect 3545 4400 3551 4401
rect 3545 4396 3546 4400
rect 3550 4396 3551 4400
rect 3545 4395 3551 4396
rect 3545 4391 3546 4395
rect 3550 4391 3551 4395
rect 3545 4390 3551 4391
rect 3545 4386 3546 4390
rect 3550 4386 3551 4390
rect 3545 4385 3551 4386
rect 3545 4381 3546 4385
rect 3550 4381 3551 4385
rect 3545 4380 3551 4381
rect 3545 4376 3546 4380
rect 3550 4376 3551 4380
rect 3545 4375 3551 4376
rect 3545 4371 3546 4375
rect 3550 4371 3551 4375
rect 3545 4370 3551 4371
rect 3545 4366 3546 4370
rect 3550 4366 3551 4370
rect 3545 4365 3551 4366
rect 3545 4361 3546 4365
rect 3550 4361 3551 4365
rect 3545 4360 3551 4361
rect 3545 4356 3546 4360
rect 3550 4356 3551 4360
rect 3545 4355 3551 4356
rect 3545 4351 3546 4355
rect 3550 4351 3551 4355
rect 3545 4350 3551 4351
rect 3545 4346 3546 4350
rect 3550 4346 3551 4350
rect 3635 4461 3636 4465
rect 3640 4461 3641 4465
rect 3635 4460 3641 4461
rect 3635 4456 3636 4460
rect 3640 4456 3641 4460
rect 3635 4455 3641 4456
rect 3635 4451 3636 4455
rect 3640 4451 3641 4455
rect 3635 4450 3641 4451
rect 3635 4446 3636 4450
rect 3640 4446 3641 4450
rect 3635 4445 3641 4446
rect 3635 4441 3636 4445
rect 3640 4441 3641 4445
rect 3635 4440 3641 4441
rect 3635 4436 3636 4440
rect 3640 4436 3641 4440
rect 3635 4435 3641 4436
rect 3635 4431 3636 4435
rect 3640 4431 3641 4435
rect 3635 4430 3641 4431
rect 3635 4426 3636 4430
rect 3640 4426 3641 4430
rect 3635 4425 3641 4426
rect 3635 4421 3636 4425
rect 3640 4421 3641 4425
rect 3635 4420 3641 4421
rect 3635 4416 3636 4420
rect 3640 4416 3641 4420
rect 3635 4415 3641 4416
rect 3635 4411 3636 4415
rect 3640 4411 3641 4415
rect 3635 4410 3641 4411
rect 3635 4406 3636 4410
rect 3640 4406 3641 4410
rect 3635 4405 3641 4406
rect 3635 4401 3636 4405
rect 3640 4401 3641 4405
rect 3635 4400 3641 4401
rect 3635 4396 3636 4400
rect 3640 4396 3641 4400
rect 3635 4395 3641 4396
rect 3635 4391 3636 4395
rect 3640 4391 3641 4395
rect 3635 4390 3641 4391
rect 3635 4386 3636 4390
rect 3640 4386 3641 4390
rect 3635 4385 3641 4386
rect 3635 4381 3636 4385
rect 3640 4381 3641 4385
rect 3635 4380 3641 4381
rect 3635 4376 3636 4380
rect 3640 4376 3641 4380
rect 3635 4375 3641 4376
rect 3635 4371 3636 4375
rect 3640 4371 3641 4375
rect 3635 4370 3641 4371
rect 3635 4366 3636 4370
rect 3640 4366 3641 4370
rect 3635 4365 3641 4366
rect 3635 4361 3636 4365
rect 3640 4361 3641 4365
rect 3635 4360 3641 4361
rect 3635 4356 3636 4360
rect 3640 4356 3641 4360
rect 3635 4355 3641 4356
rect 3635 4351 3636 4355
rect 3640 4351 3641 4355
rect 3635 4350 3641 4351
rect 3545 4345 3551 4346
rect 3545 4341 3546 4345
rect 3550 4341 3551 4345
rect 3635 4346 3636 4350
rect 3640 4346 3641 4350
rect 3635 4345 3641 4346
rect 3635 4341 3636 4345
rect 3640 4341 3641 4345
rect 3545 4340 3641 4341
rect 3545 4336 3546 4340
rect 3550 4336 3551 4340
rect 3555 4336 3556 4340
rect 3560 4336 3561 4340
rect 3565 4336 3566 4340
rect 3570 4336 3571 4340
rect 3575 4336 3576 4340
rect 3580 4336 3581 4340
rect 3585 4336 3586 4340
rect 3590 4336 3591 4340
rect 3595 4336 3596 4340
rect 3600 4336 3601 4340
rect 3605 4336 3606 4340
rect 3610 4336 3611 4340
rect 3615 4336 3616 4340
rect 3620 4336 3621 4340
rect 3625 4336 3626 4340
rect 3630 4336 3631 4340
rect 3635 4336 3636 4340
rect 3640 4336 3641 4340
rect 3545 4335 3641 4336
rect 3717 4462 3789 4464
rect 3717 4458 3719 4462
rect 3723 4458 3726 4462
rect 3730 4458 3731 4462
rect 3735 4458 3736 4462
rect 3740 4458 3741 4462
rect 3745 4458 3746 4462
rect 3750 4458 3751 4462
rect 3755 4458 3756 4462
rect 3760 4458 3761 4462
rect 3765 4458 3766 4462
rect 3770 4458 3771 4462
rect 3775 4458 3776 4462
rect 3780 4458 3783 4462
rect 3787 4458 3789 4462
rect 3717 4456 3789 4458
rect 3717 4455 3725 4456
rect 3717 4451 3719 4455
rect 3723 4451 3725 4455
rect 3717 4450 3725 4451
rect 3781 4455 3789 4456
rect 3781 4451 3783 4455
rect 3787 4451 3789 4455
rect 3781 4450 3789 4451
rect 3717 4446 3719 4450
rect 3723 4446 3725 4450
rect 3717 4445 3725 4446
rect 3717 4441 3719 4445
rect 3723 4441 3725 4445
rect 3717 4440 3725 4441
rect 3717 4436 3719 4440
rect 3723 4436 3725 4440
rect 3717 4435 3725 4436
rect 3717 4431 3719 4435
rect 3723 4431 3725 4435
rect 3717 4430 3725 4431
rect 3717 4426 3719 4430
rect 3723 4426 3725 4430
rect 3717 4425 3725 4426
rect 3717 4421 3719 4425
rect 3723 4421 3725 4425
rect 3717 4420 3725 4421
rect 3717 4416 3719 4420
rect 3723 4416 3725 4420
rect 3717 4415 3725 4416
rect 3717 4411 3719 4415
rect 3723 4411 3725 4415
rect 3717 4410 3725 4411
rect 3717 4406 3719 4410
rect 3723 4406 3725 4410
rect 3717 4405 3725 4406
rect 3717 4401 3719 4405
rect 3723 4401 3725 4405
rect 3717 4400 3725 4401
rect 3717 4396 3719 4400
rect 3723 4396 3725 4400
rect 3717 4395 3725 4396
rect 3717 4391 3719 4395
rect 3723 4391 3725 4395
rect 3717 4390 3725 4391
rect 3717 4386 3719 4390
rect 3723 4386 3725 4390
rect 3717 4385 3725 4386
rect 3717 4381 3719 4385
rect 3723 4381 3725 4385
rect 3717 4380 3725 4381
rect 3717 4376 3719 4380
rect 3723 4376 3725 4380
rect 3717 4375 3725 4376
rect 3717 4371 3719 4375
rect 3723 4371 3725 4375
rect 3717 4370 3725 4371
rect 3717 4366 3719 4370
rect 3723 4366 3725 4370
rect 3717 4365 3725 4366
rect 3717 4361 3719 4365
rect 3723 4361 3725 4365
rect 3781 4446 3783 4450
rect 3787 4446 3789 4450
rect 3781 4445 3789 4446
rect 3781 4441 3783 4445
rect 3787 4441 3789 4445
rect 3781 4440 3789 4441
rect 3781 4436 3783 4440
rect 3787 4436 3789 4440
rect 3781 4435 3789 4436
rect 3781 4431 3783 4435
rect 3787 4431 3789 4435
rect 3781 4430 3789 4431
rect 3781 4426 3783 4430
rect 3787 4426 3789 4430
rect 3781 4425 3789 4426
rect 3781 4421 3783 4425
rect 3787 4421 3789 4425
rect 3781 4420 3789 4421
rect 3781 4416 3783 4420
rect 3787 4416 3789 4420
rect 3781 4415 3789 4416
rect 3781 4411 3783 4415
rect 3787 4411 3789 4415
rect 3781 4410 3789 4411
rect 3781 4406 3783 4410
rect 3787 4406 3789 4410
rect 3781 4405 3789 4406
rect 3781 4401 3783 4405
rect 3787 4401 3789 4405
rect 3781 4400 3789 4401
rect 3781 4396 3783 4400
rect 3787 4396 3789 4400
rect 3781 4395 3789 4396
rect 3781 4391 3783 4395
rect 3787 4391 3789 4395
rect 3781 4390 3789 4391
rect 3781 4386 3783 4390
rect 3787 4386 3789 4390
rect 3781 4385 3789 4386
rect 3781 4381 3783 4385
rect 3787 4381 3789 4385
rect 3781 4380 3789 4381
rect 3781 4376 3783 4380
rect 3787 4376 3789 4380
rect 3781 4375 3789 4376
rect 3781 4371 3783 4375
rect 3787 4371 3789 4375
rect 3781 4370 3789 4371
rect 3781 4366 3783 4370
rect 3787 4366 3789 4370
rect 3781 4365 3789 4366
rect 3781 4361 3783 4365
rect 3787 4361 3789 4365
rect 3717 4360 3725 4361
rect 3717 4356 3719 4360
rect 3723 4356 3725 4360
rect 3717 4355 3725 4356
rect 3781 4360 3789 4361
rect 3781 4356 3783 4360
rect 3787 4356 3789 4360
rect 3781 4355 3789 4356
rect 3717 4353 3789 4355
rect 3717 4349 3719 4353
rect 3723 4349 3726 4353
rect 3730 4349 3731 4353
rect 3735 4349 3736 4353
rect 3740 4349 3741 4353
rect 3745 4349 3746 4353
rect 3750 4349 3751 4353
rect 3755 4349 3756 4353
rect 3760 4349 3761 4353
rect 3765 4349 3766 4353
rect 3770 4349 3771 4353
rect 3775 4349 3776 4353
rect 3780 4349 3783 4353
rect 3787 4349 3789 4353
rect 3717 4347 3789 4349
<< nsubstratendiff >>
rect 1371 9978 1467 9979
rect 1371 9974 1372 9978
rect 1376 9974 1377 9978
rect 1381 9974 1382 9978
rect 1386 9974 1387 9978
rect 1391 9974 1392 9978
rect 1396 9974 1397 9978
rect 1401 9974 1402 9978
rect 1406 9974 1407 9978
rect 1411 9974 1412 9978
rect 1416 9974 1417 9978
rect 1421 9974 1422 9978
rect 1426 9974 1427 9978
rect 1431 9974 1432 9978
rect 1436 9974 1437 9978
rect 1441 9974 1442 9978
rect 1446 9974 1447 9978
rect 1451 9974 1452 9978
rect 1456 9974 1457 9978
rect 1461 9974 1462 9978
rect 1466 9974 1467 9978
rect 1371 9973 1467 9974
rect 1371 9969 1372 9973
rect 1376 9969 1377 9973
rect 1371 9968 1377 9969
rect 1371 9964 1372 9968
rect 1376 9964 1377 9968
rect 1461 9969 1462 9973
rect 1466 9969 1467 9973
rect 1461 9968 1467 9969
rect 1371 9963 1377 9964
rect 1371 9959 1372 9963
rect 1376 9959 1377 9963
rect 1371 9958 1377 9959
rect 1371 9954 1372 9958
rect 1376 9954 1377 9958
rect 1371 9953 1377 9954
rect 1371 9949 1372 9953
rect 1376 9949 1377 9953
rect 1371 9948 1377 9949
rect 1371 9944 1372 9948
rect 1376 9944 1377 9948
rect 1371 9943 1377 9944
rect 1371 9939 1372 9943
rect 1376 9939 1377 9943
rect 1371 9938 1377 9939
rect 1371 9934 1372 9938
rect 1376 9934 1377 9938
rect 1371 9933 1377 9934
rect 1371 9929 1372 9933
rect 1376 9929 1377 9933
rect 1371 9928 1377 9929
rect 1371 9924 1372 9928
rect 1376 9924 1377 9928
rect 1371 9923 1377 9924
rect 1371 9919 1372 9923
rect 1376 9919 1377 9923
rect 1371 9918 1377 9919
rect 1371 9914 1372 9918
rect 1376 9914 1377 9918
rect 1371 9913 1377 9914
rect 1371 9909 1372 9913
rect 1376 9909 1377 9913
rect 1371 9908 1377 9909
rect 1371 9904 1372 9908
rect 1376 9904 1377 9908
rect 1371 9903 1377 9904
rect 1371 9899 1372 9903
rect 1376 9899 1377 9903
rect 1371 9898 1377 9899
rect 1371 9894 1372 9898
rect 1376 9894 1377 9898
rect 1371 9893 1377 9894
rect 1371 9889 1372 9893
rect 1376 9889 1377 9893
rect 1371 9888 1377 9889
rect 1371 9884 1372 9888
rect 1376 9884 1377 9888
rect 1371 9883 1377 9884
rect 1371 9879 1372 9883
rect 1376 9879 1377 9883
rect 1371 9878 1377 9879
rect 1371 9874 1372 9878
rect 1376 9874 1377 9878
rect 1371 9873 1377 9874
rect 1371 9869 1372 9873
rect 1376 9869 1377 9873
rect 1371 9868 1377 9869
rect 1371 9864 1372 9868
rect 1376 9864 1377 9868
rect 1371 9863 1377 9864
rect 1371 9859 1372 9863
rect 1376 9859 1377 9863
rect 1371 9858 1377 9859
rect 1371 9854 1372 9858
rect 1376 9854 1377 9858
rect 1371 9853 1377 9854
rect 1371 9849 1372 9853
rect 1376 9849 1377 9853
rect 1461 9964 1462 9968
rect 1466 9964 1467 9968
rect 1461 9963 1467 9964
rect 1461 9959 1462 9963
rect 1466 9959 1467 9963
rect 1461 9958 1467 9959
rect 1461 9954 1462 9958
rect 1466 9954 1467 9958
rect 1461 9953 1467 9954
rect 1461 9949 1462 9953
rect 1466 9949 1467 9953
rect 1461 9948 1467 9949
rect 1461 9944 1462 9948
rect 1466 9944 1467 9948
rect 1461 9943 1467 9944
rect 1461 9939 1462 9943
rect 1466 9939 1467 9943
rect 1461 9938 1467 9939
rect 1461 9934 1462 9938
rect 1466 9934 1467 9938
rect 1461 9933 1467 9934
rect 1461 9929 1462 9933
rect 1466 9929 1467 9933
rect 1461 9928 1467 9929
rect 1461 9924 1462 9928
rect 1466 9924 1467 9928
rect 1461 9923 1467 9924
rect 1461 9919 1462 9923
rect 1466 9919 1467 9923
rect 1461 9918 1467 9919
rect 1461 9914 1462 9918
rect 1466 9914 1467 9918
rect 1461 9913 1467 9914
rect 1461 9909 1462 9913
rect 1466 9909 1467 9913
rect 1461 9908 1467 9909
rect 1461 9904 1462 9908
rect 1466 9904 1467 9908
rect 1461 9903 1467 9904
rect 1461 9899 1462 9903
rect 1466 9899 1467 9903
rect 1461 9898 1467 9899
rect 1461 9894 1462 9898
rect 1466 9894 1467 9898
rect 1461 9893 1467 9894
rect 1461 9889 1462 9893
rect 1466 9889 1467 9893
rect 1461 9888 1467 9889
rect 1461 9884 1462 9888
rect 1466 9884 1467 9888
rect 1461 9883 1467 9884
rect 1461 9879 1462 9883
rect 1466 9879 1467 9883
rect 1461 9878 1467 9879
rect 1461 9874 1462 9878
rect 1466 9874 1467 9878
rect 1461 9873 1467 9874
rect 1461 9869 1462 9873
rect 1466 9869 1467 9873
rect 1461 9868 1467 9869
rect 1461 9864 1462 9868
rect 1466 9864 1467 9868
rect 1461 9863 1467 9864
rect 1461 9859 1462 9863
rect 1466 9859 1467 9863
rect 1461 9858 1467 9859
rect 1461 9854 1462 9858
rect 1466 9854 1467 9858
rect 1461 9853 1467 9854
rect 1371 9848 1377 9849
rect 1371 9844 1372 9848
rect 1376 9844 1377 9848
rect 1461 9849 1462 9853
rect 1466 9849 1467 9853
rect 1461 9848 1467 9849
rect 1461 9844 1462 9848
rect 1466 9844 1467 9848
rect 1371 9843 1467 9844
rect 1371 9839 1372 9843
rect 1376 9839 1377 9843
rect 1381 9839 1382 9843
rect 1386 9839 1387 9843
rect 1391 9839 1392 9843
rect 1396 9839 1397 9843
rect 1401 9839 1402 9843
rect 1406 9839 1407 9843
rect 1411 9839 1412 9843
rect 1416 9839 1417 9843
rect 1421 9839 1422 9843
rect 1426 9839 1427 9843
rect 1431 9839 1432 9843
rect 1436 9839 1437 9843
rect 1441 9839 1442 9843
rect 1446 9839 1447 9843
rect 1451 9839 1452 9843
rect 1456 9839 1457 9843
rect 1461 9839 1462 9843
rect 1466 9839 1467 9843
rect 1371 9838 1467 9839
rect 1543 9965 1615 9967
rect 1543 9961 1545 9965
rect 1549 9961 1552 9965
rect 1556 9961 1557 9965
rect 1561 9961 1562 9965
rect 1566 9961 1567 9965
rect 1571 9961 1572 9965
rect 1576 9961 1577 9965
rect 1581 9961 1582 9965
rect 1586 9961 1587 9965
rect 1591 9961 1592 9965
rect 1596 9961 1597 9965
rect 1601 9961 1602 9965
rect 1606 9961 1609 9965
rect 1613 9961 1615 9965
rect 1543 9959 1615 9961
rect 1543 9958 1551 9959
rect 1543 9954 1545 9958
rect 1549 9954 1551 9958
rect 1543 9953 1551 9954
rect 1607 9958 1615 9959
rect 1607 9954 1609 9958
rect 1613 9954 1615 9958
rect 1607 9953 1615 9954
rect 1543 9949 1545 9953
rect 1549 9949 1551 9953
rect 1543 9948 1551 9949
rect 1543 9944 1545 9948
rect 1549 9944 1551 9948
rect 1543 9943 1551 9944
rect 1543 9939 1545 9943
rect 1549 9939 1551 9943
rect 1543 9938 1551 9939
rect 1543 9934 1545 9938
rect 1549 9934 1551 9938
rect 1543 9933 1551 9934
rect 1543 9929 1545 9933
rect 1549 9929 1551 9933
rect 1543 9928 1551 9929
rect 1543 9924 1545 9928
rect 1549 9924 1551 9928
rect 1543 9923 1551 9924
rect 1543 9919 1545 9923
rect 1549 9919 1551 9923
rect 1543 9918 1551 9919
rect 1543 9914 1545 9918
rect 1549 9914 1551 9918
rect 1543 9913 1551 9914
rect 1543 9909 1545 9913
rect 1549 9909 1551 9913
rect 1543 9908 1551 9909
rect 1543 9904 1545 9908
rect 1549 9904 1551 9908
rect 1543 9903 1551 9904
rect 1543 9899 1545 9903
rect 1549 9899 1551 9903
rect 1543 9898 1551 9899
rect 1543 9894 1545 9898
rect 1549 9894 1551 9898
rect 1543 9893 1551 9894
rect 1543 9889 1545 9893
rect 1549 9889 1551 9893
rect 1543 9888 1551 9889
rect 1543 9884 1545 9888
rect 1549 9884 1551 9888
rect 1543 9883 1551 9884
rect 1543 9879 1545 9883
rect 1549 9879 1551 9883
rect 1543 9878 1551 9879
rect 1543 9874 1545 9878
rect 1549 9874 1551 9878
rect 1543 9873 1551 9874
rect 1543 9869 1545 9873
rect 1549 9869 1551 9873
rect 1543 9868 1551 9869
rect 1543 9864 1545 9868
rect 1549 9864 1551 9868
rect 1607 9949 1609 9953
rect 1613 9949 1615 9953
rect 1607 9948 1615 9949
rect 1607 9944 1609 9948
rect 1613 9944 1615 9948
rect 1607 9943 1615 9944
rect 1607 9939 1609 9943
rect 1613 9939 1615 9943
rect 1607 9938 1615 9939
rect 1607 9934 1609 9938
rect 1613 9934 1615 9938
rect 1607 9933 1615 9934
rect 1607 9929 1609 9933
rect 1613 9929 1615 9933
rect 1607 9928 1615 9929
rect 1607 9924 1609 9928
rect 1613 9924 1615 9928
rect 1607 9923 1615 9924
rect 1607 9919 1609 9923
rect 1613 9919 1615 9923
rect 1607 9918 1615 9919
rect 1607 9914 1609 9918
rect 1613 9914 1615 9918
rect 1607 9913 1615 9914
rect 1607 9909 1609 9913
rect 1613 9909 1615 9913
rect 1607 9908 1615 9909
rect 1607 9904 1609 9908
rect 1613 9904 1615 9908
rect 1607 9903 1615 9904
rect 1607 9899 1609 9903
rect 1613 9899 1615 9903
rect 1607 9898 1615 9899
rect 1607 9894 1609 9898
rect 1613 9894 1615 9898
rect 1607 9893 1615 9894
rect 1607 9889 1609 9893
rect 1613 9889 1615 9893
rect 1607 9888 1615 9889
rect 1607 9884 1609 9888
rect 1613 9884 1615 9888
rect 1607 9883 1615 9884
rect 1607 9879 1609 9883
rect 1613 9879 1615 9883
rect 1607 9878 1615 9879
rect 1607 9874 1609 9878
rect 1613 9874 1615 9878
rect 1607 9873 1615 9874
rect 1607 9869 1609 9873
rect 1613 9869 1615 9873
rect 1607 9868 1615 9869
rect 1607 9864 1609 9868
rect 1613 9864 1615 9868
rect 1543 9863 1551 9864
rect 1543 9859 1545 9863
rect 1549 9859 1551 9863
rect 1543 9858 1551 9859
rect 1607 9863 1615 9864
rect 1607 9859 1609 9863
rect 1613 9859 1615 9863
rect 1607 9858 1615 9859
rect 1543 9856 1615 9858
rect 1543 9852 1545 9856
rect 1549 9852 1552 9856
rect 1556 9852 1557 9856
rect 1561 9852 1562 9856
rect 1566 9852 1567 9856
rect 1571 9852 1572 9856
rect 1576 9852 1577 9856
rect 1581 9852 1582 9856
rect 1586 9852 1587 9856
rect 1591 9852 1592 9856
rect 1596 9852 1597 9856
rect 1601 9852 1602 9856
rect 1606 9852 1609 9856
rect 1613 9852 1615 9856
rect 1543 9850 1615 9852
rect 1680 9978 1776 9979
rect 1680 9974 1681 9978
rect 1685 9974 1686 9978
rect 1690 9974 1691 9978
rect 1695 9974 1696 9978
rect 1700 9974 1701 9978
rect 1705 9974 1706 9978
rect 1710 9974 1711 9978
rect 1715 9974 1716 9978
rect 1720 9974 1721 9978
rect 1725 9974 1726 9978
rect 1730 9974 1731 9978
rect 1735 9974 1736 9978
rect 1740 9974 1741 9978
rect 1745 9974 1746 9978
rect 1750 9974 1751 9978
rect 1755 9974 1756 9978
rect 1760 9974 1761 9978
rect 1765 9974 1766 9978
rect 1770 9974 1771 9978
rect 1775 9974 1776 9978
rect 1680 9973 1776 9974
rect 1680 9969 1681 9973
rect 1685 9969 1686 9973
rect 1680 9968 1686 9969
rect 1680 9964 1681 9968
rect 1685 9964 1686 9968
rect 1770 9969 1771 9973
rect 1775 9969 1776 9973
rect 1770 9968 1776 9969
rect 1680 9963 1686 9964
rect 1680 9959 1681 9963
rect 1685 9959 1686 9963
rect 1680 9958 1686 9959
rect 1680 9954 1681 9958
rect 1685 9954 1686 9958
rect 1680 9953 1686 9954
rect 1680 9949 1681 9953
rect 1685 9949 1686 9953
rect 1680 9948 1686 9949
rect 1680 9944 1681 9948
rect 1685 9944 1686 9948
rect 1680 9943 1686 9944
rect 1680 9939 1681 9943
rect 1685 9939 1686 9943
rect 1680 9938 1686 9939
rect 1680 9934 1681 9938
rect 1685 9934 1686 9938
rect 1680 9933 1686 9934
rect 1680 9929 1681 9933
rect 1685 9929 1686 9933
rect 1680 9928 1686 9929
rect 1680 9924 1681 9928
rect 1685 9924 1686 9928
rect 1680 9923 1686 9924
rect 1680 9919 1681 9923
rect 1685 9919 1686 9923
rect 1680 9918 1686 9919
rect 1680 9914 1681 9918
rect 1685 9914 1686 9918
rect 1680 9913 1686 9914
rect 1680 9909 1681 9913
rect 1685 9909 1686 9913
rect 1680 9908 1686 9909
rect 1680 9904 1681 9908
rect 1685 9904 1686 9908
rect 1680 9903 1686 9904
rect 1680 9899 1681 9903
rect 1685 9899 1686 9903
rect 1680 9898 1686 9899
rect 1680 9894 1681 9898
rect 1685 9894 1686 9898
rect 1680 9893 1686 9894
rect 1680 9889 1681 9893
rect 1685 9889 1686 9893
rect 1680 9888 1686 9889
rect 1680 9884 1681 9888
rect 1685 9884 1686 9888
rect 1680 9883 1686 9884
rect 1680 9879 1681 9883
rect 1685 9879 1686 9883
rect 1680 9878 1686 9879
rect 1680 9874 1681 9878
rect 1685 9874 1686 9878
rect 1680 9873 1686 9874
rect 1680 9869 1681 9873
rect 1685 9869 1686 9873
rect 1680 9868 1686 9869
rect 1680 9864 1681 9868
rect 1685 9864 1686 9868
rect 1680 9863 1686 9864
rect 1680 9859 1681 9863
rect 1685 9859 1686 9863
rect 1680 9858 1686 9859
rect 1680 9854 1681 9858
rect 1685 9854 1686 9858
rect 1680 9853 1686 9854
rect 1680 9849 1681 9853
rect 1685 9849 1686 9853
rect 1770 9964 1771 9968
rect 1775 9964 1776 9968
rect 1770 9963 1776 9964
rect 1770 9959 1771 9963
rect 1775 9959 1776 9963
rect 1770 9958 1776 9959
rect 1770 9954 1771 9958
rect 1775 9954 1776 9958
rect 1770 9953 1776 9954
rect 1770 9949 1771 9953
rect 1775 9949 1776 9953
rect 1770 9948 1776 9949
rect 1770 9944 1771 9948
rect 1775 9944 1776 9948
rect 1770 9943 1776 9944
rect 1770 9939 1771 9943
rect 1775 9939 1776 9943
rect 1770 9938 1776 9939
rect 1770 9934 1771 9938
rect 1775 9934 1776 9938
rect 1770 9933 1776 9934
rect 1770 9929 1771 9933
rect 1775 9929 1776 9933
rect 1770 9928 1776 9929
rect 1770 9924 1771 9928
rect 1775 9924 1776 9928
rect 1770 9923 1776 9924
rect 1770 9919 1771 9923
rect 1775 9919 1776 9923
rect 1770 9918 1776 9919
rect 1770 9914 1771 9918
rect 1775 9914 1776 9918
rect 1770 9913 1776 9914
rect 1770 9909 1771 9913
rect 1775 9909 1776 9913
rect 1770 9908 1776 9909
rect 1770 9904 1771 9908
rect 1775 9904 1776 9908
rect 1770 9903 1776 9904
rect 1770 9899 1771 9903
rect 1775 9899 1776 9903
rect 1770 9898 1776 9899
rect 1770 9894 1771 9898
rect 1775 9894 1776 9898
rect 1770 9893 1776 9894
rect 1770 9889 1771 9893
rect 1775 9889 1776 9893
rect 1770 9888 1776 9889
rect 1770 9884 1771 9888
rect 1775 9884 1776 9888
rect 1770 9883 1776 9884
rect 1770 9879 1771 9883
rect 1775 9879 1776 9883
rect 1770 9878 1776 9879
rect 1770 9874 1771 9878
rect 1775 9874 1776 9878
rect 1770 9873 1776 9874
rect 1770 9869 1771 9873
rect 1775 9869 1776 9873
rect 1770 9868 1776 9869
rect 1770 9864 1771 9868
rect 1775 9864 1776 9868
rect 1770 9863 1776 9864
rect 1770 9859 1771 9863
rect 1775 9859 1776 9863
rect 1770 9858 1776 9859
rect 1770 9854 1771 9858
rect 1775 9854 1776 9858
rect 1770 9853 1776 9854
rect 1680 9848 1686 9849
rect 1680 9844 1681 9848
rect 1685 9844 1686 9848
rect 1770 9849 1771 9853
rect 1775 9849 1776 9853
rect 1770 9848 1776 9849
rect 1770 9844 1771 9848
rect 1775 9844 1776 9848
rect 1680 9843 1776 9844
rect 1680 9839 1681 9843
rect 1685 9839 1686 9843
rect 1690 9839 1691 9843
rect 1695 9839 1696 9843
rect 1700 9839 1701 9843
rect 1705 9839 1706 9843
rect 1710 9839 1711 9843
rect 1715 9839 1716 9843
rect 1720 9839 1721 9843
rect 1725 9839 1726 9843
rect 1730 9839 1731 9843
rect 1735 9839 1736 9843
rect 1740 9839 1741 9843
rect 1745 9839 1746 9843
rect 1750 9839 1751 9843
rect 1755 9839 1756 9843
rect 1760 9839 1761 9843
rect 1765 9839 1766 9843
rect 1770 9839 1771 9843
rect 1775 9839 1776 9843
rect 1680 9838 1776 9839
rect 1852 9965 1924 9967
rect 1852 9961 1854 9965
rect 1858 9961 1861 9965
rect 1865 9961 1866 9965
rect 1870 9961 1871 9965
rect 1875 9961 1876 9965
rect 1880 9961 1881 9965
rect 1885 9961 1886 9965
rect 1890 9961 1891 9965
rect 1895 9961 1896 9965
rect 1900 9961 1901 9965
rect 1905 9961 1906 9965
rect 1910 9961 1911 9965
rect 1915 9961 1918 9965
rect 1922 9961 1924 9965
rect 1852 9959 1924 9961
rect 1852 9958 1860 9959
rect 1852 9954 1854 9958
rect 1858 9954 1860 9958
rect 1852 9953 1860 9954
rect 1916 9958 1924 9959
rect 1916 9954 1918 9958
rect 1922 9954 1924 9958
rect 1916 9953 1924 9954
rect 1852 9949 1854 9953
rect 1858 9949 1860 9953
rect 1852 9948 1860 9949
rect 1852 9944 1854 9948
rect 1858 9944 1860 9948
rect 1852 9943 1860 9944
rect 1852 9939 1854 9943
rect 1858 9939 1860 9943
rect 1852 9938 1860 9939
rect 1852 9934 1854 9938
rect 1858 9934 1860 9938
rect 1852 9933 1860 9934
rect 1852 9929 1854 9933
rect 1858 9929 1860 9933
rect 1852 9928 1860 9929
rect 1852 9924 1854 9928
rect 1858 9924 1860 9928
rect 1852 9923 1860 9924
rect 1852 9919 1854 9923
rect 1858 9919 1860 9923
rect 1852 9918 1860 9919
rect 1852 9914 1854 9918
rect 1858 9914 1860 9918
rect 1852 9913 1860 9914
rect 1852 9909 1854 9913
rect 1858 9909 1860 9913
rect 1852 9908 1860 9909
rect 1852 9904 1854 9908
rect 1858 9904 1860 9908
rect 1852 9903 1860 9904
rect 1852 9899 1854 9903
rect 1858 9899 1860 9903
rect 1852 9898 1860 9899
rect 1852 9894 1854 9898
rect 1858 9894 1860 9898
rect 1852 9893 1860 9894
rect 1852 9889 1854 9893
rect 1858 9889 1860 9893
rect 1852 9888 1860 9889
rect 1852 9884 1854 9888
rect 1858 9884 1860 9888
rect 1852 9883 1860 9884
rect 1852 9879 1854 9883
rect 1858 9879 1860 9883
rect 1852 9878 1860 9879
rect 1852 9874 1854 9878
rect 1858 9874 1860 9878
rect 1852 9873 1860 9874
rect 1852 9869 1854 9873
rect 1858 9869 1860 9873
rect 1852 9868 1860 9869
rect 1852 9864 1854 9868
rect 1858 9864 1860 9868
rect 1916 9949 1918 9953
rect 1922 9949 1924 9953
rect 1916 9948 1924 9949
rect 1916 9944 1918 9948
rect 1922 9944 1924 9948
rect 1916 9943 1924 9944
rect 1916 9939 1918 9943
rect 1922 9939 1924 9943
rect 1916 9938 1924 9939
rect 1916 9934 1918 9938
rect 1922 9934 1924 9938
rect 1916 9933 1924 9934
rect 1916 9929 1918 9933
rect 1922 9929 1924 9933
rect 1916 9928 1924 9929
rect 1916 9924 1918 9928
rect 1922 9924 1924 9928
rect 1916 9923 1924 9924
rect 1916 9919 1918 9923
rect 1922 9919 1924 9923
rect 1916 9918 1924 9919
rect 1916 9914 1918 9918
rect 1922 9914 1924 9918
rect 1916 9913 1924 9914
rect 1916 9909 1918 9913
rect 1922 9909 1924 9913
rect 1916 9908 1924 9909
rect 1916 9904 1918 9908
rect 1922 9904 1924 9908
rect 1916 9903 1924 9904
rect 1916 9899 1918 9903
rect 1922 9899 1924 9903
rect 1916 9898 1924 9899
rect 1916 9894 1918 9898
rect 1922 9894 1924 9898
rect 1916 9893 1924 9894
rect 1916 9889 1918 9893
rect 1922 9889 1924 9893
rect 1916 9888 1924 9889
rect 1916 9884 1918 9888
rect 1922 9884 1924 9888
rect 1916 9883 1924 9884
rect 1916 9879 1918 9883
rect 1922 9879 1924 9883
rect 1916 9878 1924 9879
rect 1916 9874 1918 9878
rect 1922 9874 1924 9878
rect 1916 9873 1924 9874
rect 1916 9869 1918 9873
rect 1922 9869 1924 9873
rect 1916 9868 1924 9869
rect 1916 9864 1918 9868
rect 1922 9864 1924 9868
rect 1852 9863 1860 9864
rect 1852 9859 1854 9863
rect 1858 9859 1860 9863
rect 1852 9858 1860 9859
rect 1916 9863 1924 9864
rect 1916 9859 1918 9863
rect 1922 9859 1924 9863
rect 1916 9858 1924 9859
rect 1852 9856 1924 9858
rect 1852 9852 1854 9856
rect 1858 9852 1861 9856
rect 1865 9852 1866 9856
rect 1870 9852 1871 9856
rect 1875 9852 1876 9856
rect 1880 9852 1881 9856
rect 1885 9852 1886 9856
rect 1890 9852 1891 9856
rect 1895 9852 1896 9856
rect 1900 9852 1901 9856
rect 1905 9852 1906 9856
rect 1910 9852 1911 9856
rect 1915 9852 1918 9856
rect 1922 9852 1924 9856
rect 1852 9850 1924 9852
rect 1989 9978 2085 9979
rect 1989 9974 1990 9978
rect 1994 9974 1995 9978
rect 1999 9974 2000 9978
rect 2004 9974 2005 9978
rect 2009 9974 2010 9978
rect 2014 9974 2015 9978
rect 2019 9974 2020 9978
rect 2024 9974 2025 9978
rect 2029 9974 2030 9978
rect 2034 9974 2035 9978
rect 2039 9974 2040 9978
rect 2044 9974 2045 9978
rect 2049 9974 2050 9978
rect 2054 9974 2055 9978
rect 2059 9974 2060 9978
rect 2064 9974 2065 9978
rect 2069 9974 2070 9978
rect 2074 9974 2075 9978
rect 2079 9974 2080 9978
rect 2084 9974 2085 9978
rect 1989 9973 2085 9974
rect 1989 9969 1990 9973
rect 1994 9969 1995 9973
rect 1989 9968 1995 9969
rect 1989 9964 1990 9968
rect 1994 9964 1995 9968
rect 2079 9969 2080 9973
rect 2084 9969 2085 9973
rect 2079 9968 2085 9969
rect 1989 9963 1995 9964
rect 1989 9959 1990 9963
rect 1994 9959 1995 9963
rect 1989 9958 1995 9959
rect 1989 9954 1990 9958
rect 1994 9954 1995 9958
rect 1989 9953 1995 9954
rect 1989 9949 1990 9953
rect 1994 9949 1995 9953
rect 1989 9948 1995 9949
rect 1989 9944 1990 9948
rect 1994 9944 1995 9948
rect 1989 9943 1995 9944
rect 1989 9939 1990 9943
rect 1994 9939 1995 9943
rect 1989 9938 1995 9939
rect 1989 9934 1990 9938
rect 1994 9934 1995 9938
rect 1989 9933 1995 9934
rect 1989 9929 1990 9933
rect 1994 9929 1995 9933
rect 1989 9928 1995 9929
rect 1989 9924 1990 9928
rect 1994 9924 1995 9928
rect 1989 9923 1995 9924
rect 1989 9919 1990 9923
rect 1994 9919 1995 9923
rect 1989 9918 1995 9919
rect 1989 9914 1990 9918
rect 1994 9914 1995 9918
rect 1989 9913 1995 9914
rect 1989 9909 1990 9913
rect 1994 9909 1995 9913
rect 1989 9908 1995 9909
rect 1989 9904 1990 9908
rect 1994 9904 1995 9908
rect 1989 9903 1995 9904
rect 1989 9899 1990 9903
rect 1994 9899 1995 9903
rect 1989 9898 1995 9899
rect 1989 9894 1990 9898
rect 1994 9894 1995 9898
rect 1989 9893 1995 9894
rect 1989 9889 1990 9893
rect 1994 9889 1995 9893
rect 1989 9888 1995 9889
rect 1989 9884 1990 9888
rect 1994 9884 1995 9888
rect 1989 9883 1995 9884
rect 1989 9879 1990 9883
rect 1994 9879 1995 9883
rect 1989 9878 1995 9879
rect 1989 9874 1990 9878
rect 1994 9874 1995 9878
rect 1989 9873 1995 9874
rect 1989 9869 1990 9873
rect 1994 9869 1995 9873
rect 1989 9868 1995 9869
rect 1989 9864 1990 9868
rect 1994 9864 1995 9868
rect 1989 9863 1995 9864
rect 1989 9859 1990 9863
rect 1994 9859 1995 9863
rect 1989 9858 1995 9859
rect 1989 9854 1990 9858
rect 1994 9854 1995 9858
rect 1989 9853 1995 9854
rect 1989 9849 1990 9853
rect 1994 9849 1995 9853
rect 2079 9964 2080 9968
rect 2084 9964 2085 9968
rect 2079 9963 2085 9964
rect 2079 9959 2080 9963
rect 2084 9959 2085 9963
rect 2079 9958 2085 9959
rect 2079 9954 2080 9958
rect 2084 9954 2085 9958
rect 2079 9953 2085 9954
rect 2079 9949 2080 9953
rect 2084 9949 2085 9953
rect 2079 9948 2085 9949
rect 2079 9944 2080 9948
rect 2084 9944 2085 9948
rect 2079 9943 2085 9944
rect 2079 9939 2080 9943
rect 2084 9939 2085 9943
rect 2079 9938 2085 9939
rect 2079 9934 2080 9938
rect 2084 9934 2085 9938
rect 2079 9933 2085 9934
rect 2079 9929 2080 9933
rect 2084 9929 2085 9933
rect 2079 9928 2085 9929
rect 2079 9924 2080 9928
rect 2084 9924 2085 9928
rect 2079 9923 2085 9924
rect 2079 9919 2080 9923
rect 2084 9919 2085 9923
rect 2079 9918 2085 9919
rect 2079 9914 2080 9918
rect 2084 9914 2085 9918
rect 2079 9913 2085 9914
rect 2079 9909 2080 9913
rect 2084 9909 2085 9913
rect 2079 9908 2085 9909
rect 2079 9904 2080 9908
rect 2084 9904 2085 9908
rect 2079 9903 2085 9904
rect 2079 9899 2080 9903
rect 2084 9899 2085 9903
rect 2079 9898 2085 9899
rect 2079 9894 2080 9898
rect 2084 9894 2085 9898
rect 2079 9893 2085 9894
rect 2079 9889 2080 9893
rect 2084 9889 2085 9893
rect 2079 9888 2085 9889
rect 2079 9884 2080 9888
rect 2084 9884 2085 9888
rect 2079 9883 2085 9884
rect 2079 9879 2080 9883
rect 2084 9879 2085 9883
rect 2079 9878 2085 9879
rect 2079 9874 2080 9878
rect 2084 9874 2085 9878
rect 2079 9873 2085 9874
rect 2079 9869 2080 9873
rect 2084 9869 2085 9873
rect 2079 9868 2085 9869
rect 2079 9864 2080 9868
rect 2084 9864 2085 9868
rect 2079 9863 2085 9864
rect 2079 9859 2080 9863
rect 2084 9859 2085 9863
rect 2079 9858 2085 9859
rect 2079 9854 2080 9858
rect 2084 9854 2085 9858
rect 2079 9853 2085 9854
rect 1989 9848 1995 9849
rect 1989 9844 1990 9848
rect 1994 9844 1995 9848
rect 2079 9849 2080 9853
rect 2084 9849 2085 9853
rect 2079 9848 2085 9849
rect 2079 9844 2080 9848
rect 2084 9844 2085 9848
rect 1989 9843 2085 9844
rect 1989 9839 1990 9843
rect 1994 9839 1995 9843
rect 1999 9839 2000 9843
rect 2004 9839 2005 9843
rect 2009 9839 2010 9843
rect 2014 9839 2015 9843
rect 2019 9839 2020 9843
rect 2024 9839 2025 9843
rect 2029 9839 2030 9843
rect 2034 9839 2035 9843
rect 2039 9839 2040 9843
rect 2044 9839 2045 9843
rect 2049 9839 2050 9843
rect 2054 9839 2055 9843
rect 2059 9839 2060 9843
rect 2064 9839 2065 9843
rect 2069 9839 2070 9843
rect 2074 9839 2075 9843
rect 2079 9839 2080 9843
rect 2084 9839 2085 9843
rect 1989 9838 2085 9839
rect 2161 9965 2233 9967
rect 2161 9961 2163 9965
rect 2167 9961 2170 9965
rect 2174 9961 2175 9965
rect 2179 9961 2180 9965
rect 2184 9961 2185 9965
rect 2189 9961 2190 9965
rect 2194 9961 2195 9965
rect 2199 9961 2200 9965
rect 2204 9961 2205 9965
rect 2209 9961 2210 9965
rect 2214 9961 2215 9965
rect 2219 9961 2220 9965
rect 2224 9961 2227 9965
rect 2231 9961 2233 9965
rect 2161 9959 2233 9961
rect 2161 9958 2169 9959
rect 2161 9954 2163 9958
rect 2167 9954 2169 9958
rect 2161 9953 2169 9954
rect 2225 9958 2233 9959
rect 2225 9954 2227 9958
rect 2231 9954 2233 9958
rect 2225 9953 2233 9954
rect 2161 9949 2163 9953
rect 2167 9949 2169 9953
rect 2161 9948 2169 9949
rect 2161 9944 2163 9948
rect 2167 9944 2169 9948
rect 2161 9943 2169 9944
rect 2161 9939 2163 9943
rect 2167 9939 2169 9943
rect 2161 9938 2169 9939
rect 2161 9934 2163 9938
rect 2167 9934 2169 9938
rect 2161 9933 2169 9934
rect 2161 9929 2163 9933
rect 2167 9929 2169 9933
rect 2161 9928 2169 9929
rect 2161 9924 2163 9928
rect 2167 9924 2169 9928
rect 2161 9923 2169 9924
rect 2161 9919 2163 9923
rect 2167 9919 2169 9923
rect 2161 9918 2169 9919
rect 2161 9914 2163 9918
rect 2167 9914 2169 9918
rect 2161 9913 2169 9914
rect 2161 9909 2163 9913
rect 2167 9909 2169 9913
rect 2161 9908 2169 9909
rect 2161 9904 2163 9908
rect 2167 9904 2169 9908
rect 2161 9903 2169 9904
rect 2161 9899 2163 9903
rect 2167 9899 2169 9903
rect 2161 9898 2169 9899
rect 2161 9894 2163 9898
rect 2167 9894 2169 9898
rect 2161 9893 2169 9894
rect 2161 9889 2163 9893
rect 2167 9889 2169 9893
rect 2161 9888 2169 9889
rect 2161 9884 2163 9888
rect 2167 9884 2169 9888
rect 2161 9883 2169 9884
rect 2161 9879 2163 9883
rect 2167 9879 2169 9883
rect 2161 9878 2169 9879
rect 2161 9874 2163 9878
rect 2167 9874 2169 9878
rect 2161 9873 2169 9874
rect 2161 9869 2163 9873
rect 2167 9869 2169 9873
rect 2161 9868 2169 9869
rect 2161 9864 2163 9868
rect 2167 9864 2169 9868
rect 2225 9949 2227 9953
rect 2231 9949 2233 9953
rect 2225 9948 2233 9949
rect 2225 9944 2227 9948
rect 2231 9944 2233 9948
rect 2225 9943 2233 9944
rect 2225 9939 2227 9943
rect 2231 9939 2233 9943
rect 2225 9938 2233 9939
rect 2225 9934 2227 9938
rect 2231 9934 2233 9938
rect 2225 9933 2233 9934
rect 2225 9929 2227 9933
rect 2231 9929 2233 9933
rect 2225 9928 2233 9929
rect 2225 9924 2227 9928
rect 2231 9924 2233 9928
rect 2225 9923 2233 9924
rect 2225 9919 2227 9923
rect 2231 9919 2233 9923
rect 2225 9918 2233 9919
rect 2225 9914 2227 9918
rect 2231 9914 2233 9918
rect 2225 9913 2233 9914
rect 2225 9909 2227 9913
rect 2231 9909 2233 9913
rect 2225 9908 2233 9909
rect 2225 9904 2227 9908
rect 2231 9904 2233 9908
rect 2225 9903 2233 9904
rect 2225 9899 2227 9903
rect 2231 9899 2233 9903
rect 2225 9898 2233 9899
rect 2225 9894 2227 9898
rect 2231 9894 2233 9898
rect 2225 9893 2233 9894
rect 2225 9889 2227 9893
rect 2231 9889 2233 9893
rect 2225 9888 2233 9889
rect 2225 9884 2227 9888
rect 2231 9884 2233 9888
rect 2225 9883 2233 9884
rect 2225 9879 2227 9883
rect 2231 9879 2233 9883
rect 2225 9878 2233 9879
rect 2225 9874 2227 9878
rect 2231 9874 2233 9878
rect 2225 9873 2233 9874
rect 2225 9869 2227 9873
rect 2231 9869 2233 9873
rect 2225 9868 2233 9869
rect 2225 9864 2227 9868
rect 2231 9864 2233 9868
rect 2161 9863 2169 9864
rect 2161 9859 2163 9863
rect 2167 9859 2169 9863
rect 2161 9858 2169 9859
rect 2225 9863 2233 9864
rect 2225 9859 2227 9863
rect 2231 9859 2233 9863
rect 2225 9858 2233 9859
rect 2161 9856 2233 9858
rect 2161 9852 2163 9856
rect 2167 9852 2170 9856
rect 2174 9852 2175 9856
rect 2179 9852 2180 9856
rect 2184 9852 2185 9856
rect 2189 9852 2190 9856
rect 2194 9852 2195 9856
rect 2199 9852 2200 9856
rect 2204 9852 2205 9856
rect 2209 9852 2210 9856
rect 2214 9852 2215 9856
rect 2219 9852 2220 9856
rect 2224 9852 2227 9856
rect 2231 9852 2233 9856
rect 2161 9850 2233 9852
rect 2298 9978 2394 9979
rect 2298 9974 2299 9978
rect 2303 9974 2304 9978
rect 2308 9974 2309 9978
rect 2313 9974 2314 9978
rect 2318 9974 2319 9978
rect 2323 9974 2324 9978
rect 2328 9974 2329 9978
rect 2333 9974 2334 9978
rect 2338 9974 2339 9978
rect 2343 9974 2344 9978
rect 2348 9974 2349 9978
rect 2353 9974 2354 9978
rect 2358 9974 2359 9978
rect 2363 9974 2364 9978
rect 2368 9974 2369 9978
rect 2373 9974 2374 9978
rect 2378 9974 2379 9978
rect 2383 9974 2384 9978
rect 2388 9974 2389 9978
rect 2393 9974 2394 9978
rect 2298 9973 2394 9974
rect 2298 9969 2299 9973
rect 2303 9969 2304 9973
rect 2298 9968 2304 9969
rect 2298 9964 2299 9968
rect 2303 9964 2304 9968
rect 2388 9969 2389 9973
rect 2393 9969 2394 9973
rect 2388 9968 2394 9969
rect 2298 9963 2304 9964
rect 2298 9959 2299 9963
rect 2303 9959 2304 9963
rect 2298 9958 2304 9959
rect 2298 9954 2299 9958
rect 2303 9954 2304 9958
rect 2298 9953 2304 9954
rect 2298 9949 2299 9953
rect 2303 9949 2304 9953
rect 2298 9948 2304 9949
rect 2298 9944 2299 9948
rect 2303 9944 2304 9948
rect 2298 9943 2304 9944
rect 2298 9939 2299 9943
rect 2303 9939 2304 9943
rect 2298 9938 2304 9939
rect 2298 9934 2299 9938
rect 2303 9934 2304 9938
rect 2298 9933 2304 9934
rect 2298 9929 2299 9933
rect 2303 9929 2304 9933
rect 2298 9928 2304 9929
rect 2298 9924 2299 9928
rect 2303 9924 2304 9928
rect 2298 9923 2304 9924
rect 2298 9919 2299 9923
rect 2303 9919 2304 9923
rect 2298 9918 2304 9919
rect 2298 9914 2299 9918
rect 2303 9914 2304 9918
rect 2298 9913 2304 9914
rect 2298 9909 2299 9913
rect 2303 9909 2304 9913
rect 2298 9908 2304 9909
rect 2298 9904 2299 9908
rect 2303 9904 2304 9908
rect 2298 9903 2304 9904
rect 2298 9899 2299 9903
rect 2303 9899 2304 9903
rect 2298 9898 2304 9899
rect 2298 9894 2299 9898
rect 2303 9894 2304 9898
rect 2298 9893 2304 9894
rect 2298 9889 2299 9893
rect 2303 9889 2304 9893
rect 2298 9888 2304 9889
rect 2298 9884 2299 9888
rect 2303 9884 2304 9888
rect 2298 9883 2304 9884
rect 2298 9879 2299 9883
rect 2303 9879 2304 9883
rect 2298 9878 2304 9879
rect 2298 9874 2299 9878
rect 2303 9874 2304 9878
rect 2298 9873 2304 9874
rect 2298 9869 2299 9873
rect 2303 9869 2304 9873
rect 2298 9868 2304 9869
rect 2298 9864 2299 9868
rect 2303 9864 2304 9868
rect 2298 9863 2304 9864
rect 2298 9859 2299 9863
rect 2303 9859 2304 9863
rect 2298 9858 2304 9859
rect 2298 9854 2299 9858
rect 2303 9854 2304 9858
rect 2298 9853 2304 9854
rect 2298 9849 2299 9853
rect 2303 9849 2304 9853
rect 2388 9964 2389 9968
rect 2393 9964 2394 9968
rect 2388 9963 2394 9964
rect 2388 9959 2389 9963
rect 2393 9959 2394 9963
rect 2388 9958 2394 9959
rect 2388 9954 2389 9958
rect 2393 9954 2394 9958
rect 2388 9953 2394 9954
rect 2388 9949 2389 9953
rect 2393 9949 2394 9953
rect 2388 9948 2394 9949
rect 2388 9944 2389 9948
rect 2393 9944 2394 9948
rect 2388 9943 2394 9944
rect 2388 9939 2389 9943
rect 2393 9939 2394 9943
rect 2388 9938 2394 9939
rect 2388 9934 2389 9938
rect 2393 9934 2394 9938
rect 2388 9933 2394 9934
rect 2388 9929 2389 9933
rect 2393 9929 2394 9933
rect 2388 9928 2394 9929
rect 2388 9924 2389 9928
rect 2393 9924 2394 9928
rect 2388 9923 2394 9924
rect 2388 9919 2389 9923
rect 2393 9919 2394 9923
rect 2388 9918 2394 9919
rect 2388 9914 2389 9918
rect 2393 9914 2394 9918
rect 2388 9913 2394 9914
rect 2388 9909 2389 9913
rect 2393 9909 2394 9913
rect 2388 9908 2394 9909
rect 2388 9904 2389 9908
rect 2393 9904 2394 9908
rect 2388 9903 2394 9904
rect 2388 9899 2389 9903
rect 2393 9899 2394 9903
rect 2388 9898 2394 9899
rect 2388 9894 2389 9898
rect 2393 9894 2394 9898
rect 2388 9893 2394 9894
rect 2388 9889 2389 9893
rect 2393 9889 2394 9893
rect 2388 9888 2394 9889
rect 2388 9884 2389 9888
rect 2393 9884 2394 9888
rect 2388 9883 2394 9884
rect 2388 9879 2389 9883
rect 2393 9879 2394 9883
rect 2388 9878 2394 9879
rect 2388 9874 2389 9878
rect 2393 9874 2394 9878
rect 2388 9873 2394 9874
rect 2388 9869 2389 9873
rect 2393 9869 2394 9873
rect 2388 9868 2394 9869
rect 2388 9864 2389 9868
rect 2393 9864 2394 9868
rect 2388 9863 2394 9864
rect 2388 9859 2389 9863
rect 2393 9859 2394 9863
rect 2388 9858 2394 9859
rect 2388 9854 2389 9858
rect 2393 9854 2394 9858
rect 2388 9853 2394 9854
rect 2298 9848 2304 9849
rect 2298 9844 2299 9848
rect 2303 9844 2304 9848
rect 2388 9849 2389 9853
rect 2393 9849 2394 9853
rect 2388 9848 2394 9849
rect 2388 9844 2389 9848
rect 2393 9844 2394 9848
rect 2298 9843 2394 9844
rect 2298 9839 2299 9843
rect 2303 9839 2304 9843
rect 2308 9839 2309 9843
rect 2313 9839 2314 9843
rect 2318 9839 2319 9843
rect 2323 9839 2324 9843
rect 2328 9839 2329 9843
rect 2333 9839 2334 9843
rect 2338 9839 2339 9843
rect 2343 9839 2344 9843
rect 2348 9839 2349 9843
rect 2353 9839 2354 9843
rect 2358 9839 2359 9843
rect 2363 9839 2364 9843
rect 2368 9839 2369 9843
rect 2373 9839 2374 9843
rect 2378 9839 2379 9843
rect 2383 9839 2384 9843
rect 2388 9839 2389 9843
rect 2393 9839 2394 9843
rect 2298 9838 2394 9839
rect 2470 9965 2542 9967
rect 2470 9961 2472 9965
rect 2476 9961 2479 9965
rect 2483 9961 2484 9965
rect 2488 9961 2489 9965
rect 2493 9961 2494 9965
rect 2498 9961 2499 9965
rect 2503 9961 2504 9965
rect 2508 9961 2509 9965
rect 2513 9961 2514 9965
rect 2518 9961 2519 9965
rect 2523 9961 2524 9965
rect 2528 9961 2529 9965
rect 2533 9961 2536 9965
rect 2540 9961 2542 9965
rect 2470 9959 2542 9961
rect 2470 9958 2478 9959
rect 2470 9954 2472 9958
rect 2476 9954 2478 9958
rect 2470 9953 2478 9954
rect 2534 9958 2542 9959
rect 2534 9954 2536 9958
rect 2540 9954 2542 9958
rect 2534 9953 2542 9954
rect 2470 9949 2472 9953
rect 2476 9949 2478 9953
rect 2470 9948 2478 9949
rect 2470 9944 2472 9948
rect 2476 9944 2478 9948
rect 2470 9943 2478 9944
rect 2470 9939 2472 9943
rect 2476 9939 2478 9943
rect 2470 9938 2478 9939
rect 2470 9934 2472 9938
rect 2476 9934 2478 9938
rect 2470 9933 2478 9934
rect 2470 9929 2472 9933
rect 2476 9929 2478 9933
rect 2470 9928 2478 9929
rect 2470 9924 2472 9928
rect 2476 9924 2478 9928
rect 2470 9923 2478 9924
rect 2470 9919 2472 9923
rect 2476 9919 2478 9923
rect 2470 9918 2478 9919
rect 2470 9914 2472 9918
rect 2476 9914 2478 9918
rect 2470 9913 2478 9914
rect 2470 9909 2472 9913
rect 2476 9909 2478 9913
rect 2470 9908 2478 9909
rect 2470 9904 2472 9908
rect 2476 9904 2478 9908
rect 2470 9903 2478 9904
rect 2470 9899 2472 9903
rect 2476 9899 2478 9903
rect 2470 9898 2478 9899
rect 2470 9894 2472 9898
rect 2476 9894 2478 9898
rect 2470 9893 2478 9894
rect 2470 9889 2472 9893
rect 2476 9889 2478 9893
rect 2470 9888 2478 9889
rect 2470 9884 2472 9888
rect 2476 9884 2478 9888
rect 2470 9883 2478 9884
rect 2470 9879 2472 9883
rect 2476 9879 2478 9883
rect 2470 9878 2478 9879
rect 2470 9874 2472 9878
rect 2476 9874 2478 9878
rect 2470 9873 2478 9874
rect 2470 9869 2472 9873
rect 2476 9869 2478 9873
rect 2470 9868 2478 9869
rect 2470 9864 2472 9868
rect 2476 9864 2478 9868
rect 2534 9949 2536 9953
rect 2540 9949 2542 9953
rect 2534 9948 2542 9949
rect 2534 9944 2536 9948
rect 2540 9944 2542 9948
rect 2534 9943 2542 9944
rect 2534 9939 2536 9943
rect 2540 9939 2542 9943
rect 2534 9938 2542 9939
rect 2534 9934 2536 9938
rect 2540 9934 2542 9938
rect 2534 9933 2542 9934
rect 2534 9929 2536 9933
rect 2540 9929 2542 9933
rect 2534 9928 2542 9929
rect 2534 9924 2536 9928
rect 2540 9924 2542 9928
rect 2534 9923 2542 9924
rect 2534 9919 2536 9923
rect 2540 9919 2542 9923
rect 2534 9918 2542 9919
rect 2534 9914 2536 9918
rect 2540 9914 2542 9918
rect 2534 9913 2542 9914
rect 2534 9909 2536 9913
rect 2540 9909 2542 9913
rect 2534 9908 2542 9909
rect 2534 9904 2536 9908
rect 2540 9904 2542 9908
rect 2534 9903 2542 9904
rect 2534 9899 2536 9903
rect 2540 9899 2542 9903
rect 2534 9898 2542 9899
rect 2534 9894 2536 9898
rect 2540 9894 2542 9898
rect 2534 9893 2542 9894
rect 2534 9889 2536 9893
rect 2540 9889 2542 9893
rect 2534 9888 2542 9889
rect 2534 9884 2536 9888
rect 2540 9884 2542 9888
rect 2534 9883 2542 9884
rect 2534 9879 2536 9883
rect 2540 9879 2542 9883
rect 2534 9878 2542 9879
rect 2534 9874 2536 9878
rect 2540 9874 2542 9878
rect 2534 9873 2542 9874
rect 2534 9869 2536 9873
rect 2540 9869 2542 9873
rect 2534 9868 2542 9869
rect 2534 9864 2536 9868
rect 2540 9864 2542 9868
rect 2470 9863 2478 9864
rect 2470 9859 2472 9863
rect 2476 9859 2478 9863
rect 2470 9858 2478 9859
rect 2534 9863 2542 9864
rect 2534 9859 2536 9863
rect 2540 9859 2542 9863
rect 2534 9858 2542 9859
rect 2470 9856 2542 9858
rect 2470 9852 2472 9856
rect 2476 9852 2479 9856
rect 2483 9852 2484 9856
rect 2488 9852 2489 9856
rect 2493 9852 2494 9856
rect 2498 9852 2499 9856
rect 2503 9852 2504 9856
rect 2508 9852 2509 9856
rect 2513 9852 2514 9856
rect 2518 9852 2519 9856
rect 2523 9852 2524 9856
rect 2528 9852 2529 9856
rect 2533 9852 2536 9856
rect 2540 9852 2542 9856
rect 2470 9850 2542 9852
rect 2607 9978 2703 9979
rect 2607 9974 2608 9978
rect 2612 9974 2613 9978
rect 2617 9974 2618 9978
rect 2622 9974 2623 9978
rect 2627 9974 2628 9978
rect 2632 9974 2633 9978
rect 2637 9974 2638 9978
rect 2642 9974 2643 9978
rect 2647 9974 2648 9978
rect 2652 9974 2653 9978
rect 2657 9974 2658 9978
rect 2662 9974 2663 9978
rect 2667 9974 2668 9978
rect 2672 9974 2673 9978
rect 2677 9974 2678 9978
rect 2682 9974 2683 9978
rect 2687 9974 2688 9978
rect 2692 9974 2693 9978
rect 2697 9974 2698 9978
rect 2702 9974 2703 9978
rect 2607 9973 2703 9974
rect 2607 9969 2608 9973
rect 2612 9969 2613 9973
rect 2607 9968 2613 9969
rect 2607 9964 2608 9968
rect 2612 9964 2613 9968
rect 2697 9969 2698 9973
rect 2702 9969 2703 9973
rect 2697 9968 2703 9969
rect 2607 9963 2613 9964
rect 2607 9959 2608 9963
rect 2612 9959 2613 9963
rect 2607 9958 2613 9959
rect 2607 9954 2608 9958
rect 2612 9954 2613 9958
rect 2607 9953 2613 9954
rect 2607 9949 2608 9953
rect 2612 9949 2613 9953
rect 2607 9948 2613 9949
rect 2607 9944 2608 9948
rect 2612 9944 2613 9948
rect 2607 9943 2613 9944
rect 2607 9939 2608 9943
rect 2612 9939 2613 9943
rect 2607 9938 2613 9939
rect 2607 9934 2608 9938
rect 2612 9934 2613 9938
rect 2607 9933 2613 9934
rect 2607 9929 2608 9933
rect 2612 9929 2613 9933
rect 2607 9928 2613 9929
rect 2607 9924 2608 9928
rect 2612 9924 2613 9928
rect 2607 9923 2613 9924
rect 2607 9919 2608 9923
rect 2612 9919 2613 9923
rect 2607 9918 2613 9919
rect 2607 9914 2608 9918
rect 2612 9914 2613 9918
rect 2607 9913 2613 9914
rect 2607 9909 2608 9913
rect 2612 9909 2613 9913
rect 2607 9908 2613 9909
rect 2607 9904 2608 9908
rect 2612 9904 2613 9908
rect 2607 9903 2613 9904
rect 2607 9899 2608 9903
rect 2612 9899 2613 9903
rect 2607 9898 2613 9899
rect 2607 9894 2608 9898
rect 2612 9894 2613 9898
rect 2607 9893 2613 9894
rect 2607 9889 2608 9893
rect 2612 9889 2613 9893
rect 2607 9888 2613 9889
rect 2607 9884 2608 9888
rect 2612 9884 2613 9888
rect 2607 9883 2613 9884
rect 2607 9879 2608 9883
rect 2612 9879 2613 9883
rect 2607 9878 2613 9879
rect 2607 9874 2608 9878
rect 2612 9874 2613 9878
rect 2607 9873 2613 9874
rect 2607 9869 2608 9873
rect 2612 9869 2613 9873
rect 2607 9868 2613 9869
rect 2607 9864 2608 9868
rect 2612 9864 2613 9868
rect 2607 9863 2613 9864
rect 2607 9859 2608 9863
rect 2612 9859 2613 9863
rect 2607 9858 2613 9859
rect 2607 9854 2608 9858
rect 2612 9854 2613 9858
rect 2607 9853 2613 9854
rect 2607 9849 2608 9853
rect 2612 9849 2613 9853
rect 2697 9964 2698 9968
rect 2702 9964 2703 9968
rect 2697 9963 2703 9964
rect 2697 9959 2698 9963
rect 2702 9959 2703 9963
rect 2697 9958 2703 9959
rect 2697 9954 2698 9958
rect 2702 9954 2703 9958
rect 2697 9953 2703 9954
rect 2697 9949 2698 9953
rect 2702 9949 2703 9953
rect 2697 9948 2703 9949
rect 2697 9944 2698 9948
rect 2702 9944 2703 9948
rect 2697 9943 2703 9944
rect 2697 9939 2698 9943
rect 2702 9939 2703 9943
rect 2697 9938 2703 9939
rect 2697 9934 2698 9938
rect 2702 9934 2703 9938
rect 2697 9933 2703 9934
rect 2697 9929 2698 9933
rect 2702 9929 2703 9933
rect 2697 9928 2703 9929
rect 2697 9924 2698 9928
rect 2702 9924 2703 9928
rect 2697 9923 2703 9924
rect 2697 9919 2698 9923
rect 2702 9919 2703 9923
rect 2697 9918 2703 9919
rect 2697 9914 2698 9918
rect 2702 9914 2703 9918
rect 2697 9913 2703 9914
rect 2697 9909 2698 9913
rect 2702 9909 2703 9913
rect 2697 9908 2703 9909
rect 2697 9904 2698 9908
rect 2702 9904 2703 9908
rect 2697 9903 2703 9904
rect 2697 9899 2698 9903
rect 2702 9899 2703 9903
rect 2697 9898 2703 9899
rect 2697 9894 2698 9898
rect 2702 9894 2703 9898
rect 2697 9893 2703 9894
rect 2697 9889 2698 9893
rect 2702 9889 2703 9893
rect 2697 9888 2703 9889
rect 2697 9884 2698 9888
rect 2702 9884 2703 9888
rect 2697 9883 2703 9884
rect 2697 9879 2698 9883
rect 2702 9879 2703 9883
rect 2697 9878 2703 9879
rect 2697 9874 2698 9878
rect 2702 9874 2703 9878
rect 2697 9873 2703 9874
rect 2697 9869 2698 9873
rect 2702 9869 2703 9873
rect 2697 9868 2703 9869
rect 2697 9864 2698 9868
rect 2702 9864 2703 9868
rect 2697 9863 2703 9864
rect 2697 9859 2698 9863
rect 2702 9859 2703 9863
rect 2697 9858 2703 9859
rect 2697 9854 2698 9858
rect 2702 9854 2703 9858
rect 2697 9853 2703 9854
rect 2607 9848 2613 9849
rect 2607 9844 2608 9848
rect 2612 9844 2613 9848
rect 2697 9849 2698 9853
rect 2702 9849 2703 9853
rect 2697 9848 2703 9849
rect 2697 9844 2698 9848
rect 2702 9844 2703 9848
rect 2607 9843 2703 9844
rect 2607 9839 2608 9843
rect 2612 9839 2613 9843
rect 2617 9839 2618 9843
rect 2622 9839 2623 9843
rect 2627 9839 2628 9843
rect 2632 9839 2633 9843
rect 2637 9839 2638 9843
rect 2642 9839 2643 9843
rect 2647 9839 2648 9843
rect 2652 9839 2653 9843
rect 2657 9839 2658 9843
rect 2662 9839 2663 9843
rect 2667 9839 2668 9843
rect 2672 9839 2673 9843
rect 2677 9839 2678 9843
rect 2682 9839 2683 9843
rect 2687 9839 2688 9843
rect 2692 9839 2693 9843
rect 2697 9839 2698 9843
rect 2702 9839 2703 9843
rect 2607 9838 2703 9839
rect 2779 9965 2851 9967
rect 2779 9961 2781 9965
rect 2785 9961 2788 9965
rect 2792 9961 2793 9965
rect 2797 9961 2798 9965
rect 2802 9961 2803 9965
rect 2807 9961 2808 9965
rect 2812 9961 2813 9965
rect 2817 9961 2818 9965
rect 2822 9961 2823 9965
rect 2827 9961 2828 9965
rect 2832 9961 2833 9965
rect 2837 9961 2838 9965
rect 2842 9961 2845 9965
rect 2849 9961 2851 9965
rect 2779 9959 2851 9961
rect 2779 9958 2787 9959
rect 2779 9954 2781 9958
rect 2785 9954 2787 9958
rect 2779 9953 2787 9954
rect 2843 9958 2851 9959
rect 2843 9954 2845 9958
rect 2849 9954 2851 9958
rect 2843 9953 2851 9954
rect 2779 9949 2781 9953
rect 2785 9949 2787 9953
rect 2779 9948 2787 9949
rect 2779 9944 2781 9948
rect 2785 9944 2787 9948
rect 2779 9943 2787 9944
rect 2779 9939 2781 9943
rect 2785 9939 2787 9943
rect 2779 9938 2787 9939
rect 2779 9934 2781 9938
rect 2785 9934 2787 9938
rect 2779 9933 2787 9934
rect 2779 9929 2781 9933
rect 2785 9929 2787 9933
rect 2779 9928 2787 9929
rect 2779 9924 2781 9928
rect 2785 9924 2787 9928
rect 2779 9923 2787 9924
rect 2779 9919 2781 9923
rect 2785 9919 2787 9923
rect 2779 9918 2787 9919
rect 2779 9914 2781 9918
rect 2785 9914 2787 9918
rect 2779 9913 2787 9914
rect 2779 9909 2781 9913
rect 2785 9909 2787 9913
rect 2779 9908 2787 9909
rect 2779 9904 2781 9908
rect 2785 9904 2787 9908
rect 2779 9903 2787 9904
rect 2779 9899 2781 9903
rect 2785 9899 2787 9903
rect 2779 9898 2787 9899
rect 2779 9894 2781 9898
rect 2785 9894 2787 9898
rect 2779 9893 2787 9894
rect 2779 9889 2781 9893
rect 2785 9889 2787 9893
rect 2779 9888 2787 9889
rect 2779 9884 2781 9888
rect 2785 9884 2787 9888
rect 2779 9883 2787 9884
rect 2779 9879 2781 9883
rect 2785 9879 2787 9883
rect 2779 9878 2787 9879
rect 2779 9874 2781 9878
rect 2785 9874 2787 9878
rect 2779 9873 2787 9874
rect 2779 9869 2781 9873
rect 2785 9869 2787 9873
rect 2779 9868 2787 9869
rect 2779 9864 2781 9868
rect 2785 9864 2787 9868
rect 2843 9949 2845 9953
rect 2849 9949 2851 9953
rect 2843 9948 2851 9949
rect 2843 9944 2845 9948
rect 2849 9944 2851 9948
rect 2843 9943 2851 9944
rect 2843 9939 2845 9943
rect 2849 9939 2851 9943
rect 2843 9938 2851 9939
rect 2843 9934 2845 9938
rect 2849 9934 2851 9938
rect 2843 9933 2851 9934
rect 2843 9929 2845 9933
rect 2849 9929 2851 9933
rect 2843 9928 2851 9929
rect 2843 9924 2845 9928
rect 2849 9924 2851 9928
rect 2843 9923 2851 9924
rect 2843 9919 2845 9923
rect 2849 9919 2851 9923
rect 2843 9918 2851 9919
rect 2843 9914 2845 9918
rect 2849 9914 2851 9918
rect 2843 9913 2851 9914
rect 2843 9909 2845 9913
rect 2849 9909 2851 9913
rect 2843 9908 2851 9909
rect 2843 9904 2845 9908
rect 2849 9904 2851 9908
rect 2843 9903 2851 9904
rect 2843 9899 2845 9903
rect 2849 9899 2851 9903
rect 2843 9898 2851 9899
rect 2843 9894 2845 9898
rect 2849 9894 2851 9898
rect 2843 9893 2851 9894
rect 2843 9889 2845 9893
rect 2849 9889 2851 9893
rect 2843 9888 2851 9889
rect 2843 9884 2845 9888
rect 2849 9884 2851 9888
rect 2843 9883 2851 9884
rect 2843 9879 2845 9883
rect 2849 9879 2851 9883
rect 2843 9878 2851 9879
rect 2843 9874 2845 9878
rect 2849 9874 2851 9878
rect 2843 9873 2851 9874
rect 2843 9869 2845 9873
rect 2849 9869 2851 9873
rect 2843 9868 2851 9869
rect 2843 9864 2845 9868
rect 2849 9864 2851 9868
rect 2779 9863 2787 9864
rect 2779 9859 2781 9863
rect 2785 9859 2787 9863
rect 2779 9858 2787 9859
rect 2843 9863 2851 9864
rect 2843 9859 2845 9863
rect 2849 9859 2851 9863
rect 2843 9858 2851 9859
rect 2779 9856 2851 9858
rect 2779 9852 2781 9856
rect 2785 9852 2788 9856
rect 2792 9852 2793 9856
rect 2797 9852 2798 9856
rect 2802 9852 2803 9856
rect 2807 9852 2808 9856
rect 2812 9852 2813 9856
rect 2817 9852 2818 9856
rect 2822 9852 2823 9856
rect 2827 9852 2828 9856
rect 2832 9852 2833 9856
rect 2837 9852 2838 9856
rect 2842 9852 2845 9856
rect 2849 9852 2851 9856
rect 2779 9850 2851 9852
rect 2916 9978 3012 9979
rect 2916 9974 2917 9978
rect 2921 9974 2922 9978
rect 2926 9974 2927 9978
rect 2931 9974 2932 9978
rect 2936 9974 2937 9978
rect 2941 9974 2942 9978
rect 2946 9974 2947 9978
rect 2951 9974 2952 9978
rect 2956 9974 2957 9978
rect 2961 9974 2962 9978
rect 2966 9974 2967 9978
rect 2971 9974 2972 9978
rect 2976 9974 2977 9978
rect 2981 9974 2982 9978
rect 2986 9974 2987 9978
rect 2991 9974 2992 9978
rect 2996 9974 2997 9978
rect 3001 9974 3002 9978
rect 3006 9974 3007 9978
rect 3011 9974 3012 9978
rect 2916 9973 3012 9974
rect 2916 9969 2917 9973
rect 2921 9969 2922 9973
rect 2916 9968 2922 9969
rect 2916 9964 2917 9968
rect 2921 9964 2922 9968
rect 3006 9969 3007 9973
rect 3011 9969 3012 9973
rect 3006 9968 3012 9969
rect 2916 9963 2922 9964
rect 2916 9959 2917 9963
rect 2921 9959 2922 9963
rect 2916 9958 2922 9959
rect 2916 9954 2917 9958
rect 2921 9954 2922 9958
rect 2916 9953 2922 9954
rect 2916 9949 2917 9953
rect 2921 9949 2922 9953
rect 2916 9948 2922 9949
rect 2916 9944 2917 9948
rect 2921 9944 2922 9948
rect 2916 9943 2922 9944
rect 2916 9939 2917 9943
rect 2921 9939 2922 9943
rect 2916 9938 2922 9939
rect 2916 9934 2917 9938
rect 2921 9934 2922 9938
rect 2916 9933 2922 9934
rect 2916 9929 2917 9933
rect 2921 9929 2922 9933
rect 2916 9928 2922 9929
rect 2916 9924 2917 9928
rect 2921 9924 2922 9928
rect 2916 9923 2922 9924
rect 2916 9919 2917 9923
rect 2921 9919 2922 9923
rect 2916 9918 2922 9919
rect 2916 9914 2917 9918
rect 2921 9914 2922 9918
rect 2916 9913 2922 9914
rect 2916 9909 2917 9913
rect 2921 9909 2922 9913
rect 2916 9908 2922 9909
rect 2916 9904 2917 9908
rect 2921 9904 2922 9908
rect 2916 9903 2922 9904
rect 2916 9899 2917 9903
rect 2921 9899 2922 9903
rect 2916 9898 2922 9899
rect 2916 9894 2917 9898
rect 2921 9894 2922 9898
rect 2916 9893 2922 9894
rect 2916 9889 2917 9893
rect 2921 9889 2922 9893
rect 2916 9888 2922 9889
rect 2916 9884 2917 9888
rect 2921 9884 2922 9888
rect 2916 9883 2922 9884
rect 2916 9879 2917 9883
rect 2921 9879 2922 9883
rect 2916 9878 2922 9879
rect 2916 9874 2917 9878
rect 2921 9874 2922 9878
rect 2916 9873 2922 9874
rect 2916 9869 2917 9873
rect 2921 9869 2922 9873
rect 2916 9868 2922 9869
rect 2916 9864 2917 9868
rect 2921 9864 2922 9868
rect 2916 9863 2922 9864
rect 2916 9859 2917 9863
rect 2921 9859 2922 9863
rect 2916 9858 2922 9859
rect 2916 9854 2917 9858
rect 2921 9854 2922 9858
rect 2916 9853 2922 9854
rect 2916 9849 2917 9853
rect 2921 9849 2922 9853
rect 3006 9964 3007 9968
rect 3011 9964 3012 9968
rect 3006 9963 3012 9964
rect 3006 9959 3007 9963
rect 3011 9959 3012 9963
rect 3006 9958 3012 9959
rect 3006 9954 3007 9958
rect 3011 9954 3012 9958
rect 3006 9953 3012 9954
rect 3006 9949 3007 9953
rect 3011 9949 3012 9953
rect 3006 9948 3012 9949
rect 3006 9944 3007 9948
rect 3011 9944 3012 9948
rect 3006 9943 3012 9944
rect 3006 9939 3007 9943
rect 3011 9939 3012 9943
rect 3006 9938 3012 9939
rect 3006 9934 3007 9938
rect 3011 9934 3012 9938
rect 3006 9933 3012 9934
rect 3006 9929 3007 9933
rect 3011 9929 3012 9933
rect 3006 9928 3012 9929
rect 3006 9924 3007 9928
rect 3011 9924 3012 9928
rect 3006 9923 3012 9924
rect 3006 9919 3007 9923
rect 3011 9919 3012 9923
rect 3006 9918 3012 9919
rect 3006 9914 3007 9918
rect 3011 9914 3012 9918
rect 3006 9913 3012 9914
rect 3006 9909 3007 9913
rect 3011 9909 3012 9913
rect 3006 9908 3012 9909
rect 3006 9904 3007 9908
rect 3011 9904 3012 9908
rect 3006 9903 3012 9904
rect 3006 9899 3007 9903
rect 3011 9899 3012 9903
rect 3006 9898 3012 9899
rect 3006 9894 3007 9898
rect 3011 9894 3012 9898
rect 3006 9893 3012 9894
rect 3006 9889 3007 9893
rect 3011 9889 3012 9893
rect 3006 9888 3012 9889
rect 3006 9884 3007 9888
rect 3011 9884 3012 9888
rect 3006 9883 3012 9884
rect 3006 9879 3007 9883
rect 3011 9879 3012 9883
rect 3006 9878 3012 9879
rect 3006 9874 3007 9878
rect 3011 9874 3012 9878
rect 3006 9873 3012 9874
rect 3006 9869 3007 9873
rect 3011 9869 3012 9873
rect 3006 9868 3012 9869
rect 3006 9864 3007 9868
rect 3011 9864 3012 9868
rect 3006 9863 3012 9864
rect 3006 9859 3007 9863
rect 3011 9859 3012 9863
rect 3006 9858 3012 9859
rect 3006 9854 3007 9858
rect 3011 9854 3012 9858
rect 3006 9853 3012 9854
rect 2916 9848 2922 9849
rect 2916 9844 2917 9848
rect 2921 9844 2922 9848
rect 3006 9849 3007 9853
rect 3011 9849 3012 9853
rect 3006 9848 3012 9849
rect 3006 9844 3007 9848
rect 3011 9844 3012 9848
rect 2916 9843 3012 9844
rect 2916 9839 2917 9843
rect 2921 9839 2922 9843
rect 2926 9839 2927 9843
rect 2931 9839 2932 9843
rect 2936 9839 2937 9843
rect 2941 9839 2942 9843
rect 2946 9839 2947 9843
rect 2951 9839 2952 9843
rect 2956 9839 2957 9843
rect 2961 9839 2962 9843
rect 2966 9839 2967 9843
rect 2971 9839 2972 9843
rect 2976 9839 2977 9843
rect 2981 9839 2982 9843
rect 2986 9839 2987 9843
rect 2991 9839 2992 9843
rect 2996 9839 2997 9843
rect 3001 9839 3002 9843
rect 3006 9839 3007 9843
rect 3011 9839 3012 9843
rect 2916 9838 3012 9839
rect 3088 9965 3160 9967
rect 3088 9961 3090 9965
rect 3094 9961 3097 9965
rect 3101 9961 3102 9965
rect 3106 9961 3107 9965
rect 3111 9961 3112 9965
rect 3116 9961 3117 9965
rect 3121 9961 3122 9965
rect 3126 9961 3127 9965
rect 3131 9961 3132 9965
rect 3136 9961 3137 9965
rect 3141 9961 3142 9965
rect 3146 9961 3147 9965
rect 3151 9961 3154 9965
rect 3158 9961 3160 9965
rect 3088 9959 3160 9961
rect 3088 9958 3096 9959
rect 3088 9954 3090 9958
rect 3094 9954 3096 9958
rect 3088 9953 3096 9954
rect 3152 9958 3160 9959
rect 3152 9954 3154 9958
rect 3158 9954 3160 9958
rect 3152 9953 3160 9954
rect 3088 9949 3090 9953
rect 3094 9949 3096 9953
rect 3088 9948 3096 9949
rect 3088 9944 3090 9948
rect 3094 9944 3096 9948
rect 3088 9943 3096 9944
rect 3088 9939 3090 9943
rect 3094 9939 3096 9943
rect 3088 9938 3096 9939
rect 3088 9934 3090 9938
rect 3094 9934 3096 9938
rect 3088 9933 3096 9934
rect 3088 9929 3090 9933
rect 3094 9929 3096 9933
rect 3088 9928 3096 9929
rect 3088 9924 3090 9928
rect 3094 9924 3096 9928
rect 3088 9923 3096 9924
rect 3088 9919 3090 9923
rect 3094 9919 3096 9923
rect 3088 9918 3096 9919
rect 3088 9914 3090 9918
rect 3094 9914 3096 9918
rect 3088 9913 3096 9914
rect 3088 9909 3090 9913
rect 3094 9909 3096 9913
rect 3088 9908 3096 9909
rect 3088 9904 3090 9908
rect 3094 9904 3096 9908
rect 3088 9903 3096 9904
rect 3088 9899 3090 9903
rect 3094 9899 3096 9903
rect 3088 9898 3096 9899
rect 3088 9894 3090 9898
rect 3094 9894 3096 9898
rect 3088 9893 3096 9894
rect 3088 9889 3090 9893
rect 3094 9889 3096 9893
rect 3088 9888 3096 9889
rect 3088 9884 3090 9888
rect 3094 9884 3096 9888
rect 3088 9883 3096 9884
rect 3088 9879 3090 9883
rect 3094 9879 3096 9883
rect 3088 9878 3096 9879
rect 3088 9874 3090 9878
rect 3094 9874 3096 9878
rect 3088 9873 3096 9874
rect 3088 9869 3090 9873
rect 3094 9869 3096 9873
rect 3088 9868 3096 9869
rect 3088 9864 3090 9868
rect 3094 9864 3096 9868
rect 3152 9949 3154 9953
rect 3158 9949 3160 9953
rect 3152 9948 3160 9949
rect 3152 9944 3154 9948
rect 3158 9944 3160 9948
rect 3152 9943 3160 9944
rect 3152 9939 3154 9943
rect 3158 9939 3160 9943
rect 3152 9938 3160 9939
rect 3152 9934 3154 9938
rect 3158 9934 3160 9938
rect 3152 9933 3160 9934
rect 3152 9929 3154 9933
rect 3158 9929 3160 9933
rect 3152 9928 3160 9929
rect 3152 9924 3154 9928
rect 3158 9924 3160 9928
rect 3152 9923 3160 9924
rect 3152 9919 3154 9923
rect 3158 9919 3160 9923
rect 3152 9918 3160 9919
rect 3152 9914 3154 9918
rect 3158 9914 3160 9918
rect 3152 9913 3160 9914
rect 3152 9909 3154 9913
rect 3158 9909 3160 9913
rect 3152 9908 3160 9909
rect 3152 9904 3154 9908
rect 3158 9904 3160 9908
rect 3152 9903 3160 9904
rect 3152 9899 3154 9903
rect 3158 9899 3160 9903
rect 3152 9898 3160 9899
rect 3152 9894 3154 9898
rect 3158 9894 3160 9898
rect 3152 9893 3160 9894
rect 3152 9889 3154 9893
rect 3158 9889 3160 9893
rect 3152 9888 3160 9889
rect 3152 9884 3154 9888
rect 3158 9884 3160 9888
rect 3152 9883 3160 9884
rect 3152 9879 3154 9883
rect 3158 9879 3160 9883
rect 3152 9878 3160 9879
rect 3152 9874 3154 9878
rect 3158 9874 3160 9878
rect 3152 9873 3160 9874
rect 3152 9869 3154 9873
rect 3158 9869 3160 9873
rect 3152 9868 3160 9869
rect 3152 9864 3154 9868
rect 3158 9864 3160 9868
rect 3088 9863 3096 9864
rect 3088 9859 3090 9863
rect 3094 9859 3096 9863
rect 3088 9858 3096 9859
rect 3152 9863 3160 9864
rect 3152 9859 3154 9863
rect 3158 9859 3160 9863
rect 3152 9858 3160 9859
rect 3088 9856 3160 9858
rect 3088 9852 3090 9856
rect 3094 9852 3097 9856
rect 3101 9852 3102 9856
rect 3106 9852 3107 9856
rect 3111 9852 3112 9856
rect 3116 9852 3117 9856
rect 3121 9852 3122 9856
rect 3126 9852 3127 9856
rect 3131 9852 3132 9856
rect 3136 9852 3137 9856
rect 3141 9852 3142 9856
rect 3146 9852 3147 9856
rect 3151 9852 3154 9856
rect 3158 9852 3160 9856
rect 3088 9850 3160 9852
rect 3225 9978 3321 9979
rect 3225 9974 3226 9978
rect 3230 9974 3231 9978
rect 3235 9974 3236 9978
rect 3240 9974 3241 9978
rect 3245 9974 3246 9978
rect 3250 9974 3251 9978
rect 3255 9974 3256 9978
rect 3260 9974 3261 9978
rect 3265 9974 3266 9978
rect 3270 9974 3271 9978
rect 3275 9974 3276 9978
rect 3280 9974 3281 9978
rect 3285 9974 3286 9978
rect 3290 9974 3291 9978
rect 3295 9974 3296 9978
rect 3300 9974 3301 9978
rect 3305 9974 3306 9978
rect 3310 9974 3311 9978
rect 3315 9974 3316 9978
rect 3320 9974 3321 9978
rect 3225 9973 3321 9974
rect 3225 9969 3226 9973
rect 3230 9969 3231 9973
rect 3225 9968 3231 9969
rect 3225 9964 3226 9968
rect 3230 9964 3231 9968
rect 3315 9969 3316 9973
rect 3320 9969 3321 9973
rect 3315 9968 3321 9969
rect 3225 9963 3231 9964
rect 3225 9959 3226 9963
rect 3230 9959 3231 9963
rect 3225 9958 3231 9959
rect 3225 9954 3226 9958
rect 3230 9954 3231 9958
rect 3225 9953 3231 9954
rect 3225 9949 3226 9953
rect 3230 9949 3231 9953
rect 3225 9948 3231 9949
rect 3225 9944 3226 9948
rect 3230 9944 3231 9948
rect 3225 9943 3231 9944
rect 3225 9939 3226 9943
rect 3230 9939 3231 9943
rect 3225 9938 3231 9939
rect 3225 9934 3226 9938
rect 3230 9934 3231 9938
rect 3225 9933 3231 9934
rect 3225 9929 3226 9933
rect 3230 9929 3231 9933
rect 3225 9928 3231 9929
rect 3225 9924 3226 9928
rect 3230 9924 3231 9928
rect 3225 9923 3231 9924
rect 3225 9919 3226 9923
rect 3230 9919 3231 9923
rect 3225 9918 3231 9919
rect 3225 9914 3226 9918
rect 3230 9914 3231 9918
rect 3225 9913 3231 9914
rect 3225 9909 3226 9913
rect 3230 9909 3231 9913
rect 3225 9908 3231 9909
rect 3225 9904 3226 9908
rect 3230 9904 3231 9908
rect 3225 9903 3231 9904
rect 3225 9899 3226 9903
rect 3230 9899 3231 9903
rect 3225 9898 3231 9899
rect 3225 9894 3226 9898
rect 3230 9894 3231 9898
rect 3225 9893 3231 9894
rect 3225 9889 3226 9893
rect 3230 9889 3231 9893
rect 3225 9888 3231 9889
rect 3225 9884 3226 9888
rect 3230 9884 3231 9888
rect 3225 9883 3231 9884
rect 3225 9879 3226 9883
rect 3230 9879 3231 9883
rect 3225 9878 3231 9879
rect 3225 9874 3226 9878
rect 3230 9874 3231 9878
rect 3225 9873 3231 9874
rect 3225 9869 3226 9873
rect 3230 9869 3231 9873
rect 3225 9868 3231 9869
rect 3225 9864 3226 9868
rect 3230 9864 3231 9868
rect 3225 9863 3231 9864
rect 3225 9859 3226 9863
rect 3230 9859 3231 9863
rect 3225 9858 3231 9859
rect 3225 9854 3226 9858
rect 3230 9854 3231 9858
rect 3225 9853 3231 9854
rect 3225 9849 3226 9853
rect 3230 9849 3231 9853
rect 3315 9964 3316 9968
rect 3320 9964 3321 9968
rect 3315 9963 3321 9964
rect 3315 9959 3316 9963
rect 3320 9959 3321 9963
rect 3315 9958 3321 9959
rect 3315 9954 3316 9958
rect 3320 9954 3321 9958
rect 3315 9953 3321 9954
rect 3315 9949 3316 9953
rect 3320 9949 3321 9953
rect 3315 9948 3321 9949
rect 3315 9944 3316 9948
rect 3320 9944 3321 9948
rect 3315 9943 3321 9944
rect 3315 9939 3316 9943
rect 3320 9939 3321 9943
rect 3315 9938 3321 9939
rect 3315 9934 3316 9938
rect 3320 9934 3321 9938
rect 3315 9933 3321 9934
rect 3315 9929 3316 9933
rect 3320 9929 3321 9933
rect 3315 9928 3321 9929
rect 3315 9924 3316 9928
rect 3320 9924 3321 9928
rect 3315 9923 3321 9924
rect 3315 9919 3316 9923
rect 3320 9919 3321 9923
rect 3315 9918 3321 9919
rect 3315 9914 3316 9918
rect 3320 9914 3321 9918
rect 3315 9913 3321 9914
rect 3315 9909 3316 9913
rect 3320 9909 3321 9913
rect 3315 9908 3321 9909
rect 3315 9904 3316 9908
rect 3320 9904 3321 9908
rect 3315 9903 3321 9904
rect 3315 9899 3316 9903
rect 3320 9899 3321 9903
rect 3315 9898 3321 9899
rect 3315 9894 3316 9898
rect 3320 9894 3321 9898
rect 3315 9893 3321 9894
rect 3315 9889 3316 9893
rect 3320 9889 3321 9893
rect 3315 9888 3321 9889
rect 3315 9884 3316 9888
rect 3320 9884 3321 9888
rect 3315 9883 3321 9884
rect 3315 9879 3316 9883
rect 3320 9879 3321 9883
rect 3315 9878 3321 9879
rect 3315 9874 3316 9878
rect 3320 9874 3321 9878
rect 3315 9873 3321 9874
rect 3315 9869 3316 9873
rect 3320 9869 3321 9873
rect 3315 9868 3321 9869
rect 3315 9864 3316 9868
rect 3320 9864 3321 9868
rect 3315 9863 3321 9864
rect 3315 9859 3316 9863
rect 3320 9859 3321 9863
rect 3315 9858 3321 9859
rect 3315 9854 3316 9858
rect 3320 9854 3321 9858
rect 3315 9853 3321 9854
rect 3225 9848 3231 9849
rect 3225 9844 3226 9848
rect 3230 9844 3231 9848
rect 3315 9849 3316 9853
rect 3320 9849 3321 9853
rect 3315 9848 3321 9849
rect 3315 9844 3316 9848
rect 3320 9844 3321 9848
rect 3225 9843 3321 9844
rect 3225 9839 3226 9843
rect 3230 9839 3231 9843
rect 3235 9839 3236 9843
rect 3240 9839 3241 9843
rect 3245 9839 3246 9843
rect 3250 9839 3251 9843
rect 3255 9839 3256 9843
rect 3260 9839 3261 9843
rect 3265 9839 3266 9843
rect 3270 9839 3271 9843
rect 3275 9839 3276 9843
rect 3280 9839 3281 9843
rect 3285 9839 3286 9843
rect 3290 9839 3291 9843
rect 3295 9839 3296 9843
rect 3300 9839 3301 9843
rect 3305 9839 3306 9843
rect 3310 9839 3311 9843
rect 3315 9839 3316 9843
rect 3320 9839 3321 9843
rect 3225 9838 3321 9839
rect 3397 9965 3469 9967
rect 3397 9961 3399 9965
rect 3403 9961 3406 9965
rect 3410 9961 3411 9965
rect 3415 9961 3416 9965
rect 3420 9961 3421 9965
rect 3425 9961 3426 9965
rect 3430 9961 3431 9965
rect 3435 9961 3436 9965
rect 3440 9961 3441 9965
rect 3445 9961 3446 9965
rect 3450 9961 3451 9965
rect 3455 9961 3456 9965
rect 3460 9961 3463 9965
rect 3467 9961 3469 9965
rect 3397 9959 3469 9961
rect 3397 9958 3405 9959
rect 3397 9954 3399 9958
rect 3403 9954 3405 9958
rect 3397 9953 3405 9954
rect 3461 9958 3469 9959
rect 3461 9954 3463 9958
rect 3467 9954 3469 9958
rect 3461 9953 3469 9954
rect 3397 9949 3399 9953
rect 3403 9949 3405 9953
rect 3397 9948 3405 9949
rect 3397 9944 3399 9948
rect 3403 9944 3405 9948
rect 3397 9943 3405 9944
rect 3397 9939 3399 9943
rect 3403 9939 3405 9943
rect 3397 9938 3405 9939
rect 3397 9934 3399 9938
rect 3403 9934 3405 9938
rect 3397 9933 3405 9934
rect 3397 9929 3399 9933
rect 3403 9929 3405 9933
rect 3397 9928 3405 9929
rect 3397 9924 3399 9928
rect 3403 9924 3405 9928
rect 3397 9923 3405 9924
rect 3397 9919 3399 9923
rect 3403 9919 3405 9923
rect 3397 9918 3405 9919
rect 3397 9914 3399 9918
rect 3403 9914 3405 9918
rect 3397 9913 3405 9914
rect 3397 9909 3399 9913
rect 3403 9909 3405 9913
rect 3397 9908 3405 9909
rect 3397 9904 3399 9908
rect 3403 9904 3405 9908
rect 3397 9903 3405 9904
rect 3397 9899 3399 9903
rect 3403 9899 3405 9903
rect 3397 9898 3405 9899
rect 3397 9894 3399 9898
rect 3403 9894 3405 9898
rect 3397 9893 3405 9894
rect 3397 9889 3399 9893
rect 3403 9889 3405 9893
rect 3397 9888 3405 9889
rect 3397 9884 3399 9888
rect 3403 9884 3405 9888
rect 3397 9883 3405 9884
rect 3397 9879 3399 9883
rect 3403 9879 3405 9883
rect 3397 9878 3405 9879
rect 3397 9874 3399 9878
rect 3403 9874 3405 9878
rect 3397 9873 3405 9874
rect 3397 9869 3399 9873
rect 3403 9869 3405 9873
rect 3397 9868 3405 9869
rect 3397 9864 3399 9868
rect 3403 9864 3405 9868
rect 3461 9949 3463 9953
rect 3467 9949 3469 9953
rect 3461 9948 3469 9949
rect 3461 9944 3463 9948
rect 3467 9944 3469 9948
rect 3461 9943 3469 9944
rect 3461 9939 3463 9943
rect 3467 9939 3469 9943
rect 3461 9938 3469 9939
rect 3461 9934 3463 9938
rect 3467 9934 3469 9938
rect 3461 9933 3469 9934
rect 3461 9929 3463 9933
rect 3467 9929 3469 9933
rect 3461 9928 3469 9929
rect 3461 9924 3463 9928
rect 3467 9924 3469 9928
rect 3461 9923 3469 9924
rect 3461 9919 3463 9923
rect 3467 9919 3469 9923
rect 3461 9918 3469 9919
rect 3461 9914 3463 9918
rect 3467 9914 3469 9918
rect 3461 9913 3469 9914
rect 3461 9909 3463 9913
rect 3467 9909 3469 9913
rect 3461 9908 3469 9909
rect 3461 9904 3463 9908
rect 3467 9904 3469 9908
rect 3461 9903 3469 9904
rect 3461 9899 3463 9903
rect 3467 9899 3469 9903
rect 3461 9898 3469 9899
rect 3461 9894 3463 9898
rect 3467 9894 3469 9898
rect 3461 9893 3469 9894
rect 3461 9889 3463 9893
rect 3467 9889 3469 9893
rect 3461 9888 3469 9889
rect 3461 9884 3463 9888
rect 3467 9884 3469 9888
rect 3461 9883 3469 9884
rect 3461 9879 3463 9883
rect 3467 9879 3469 9883
rect 3461 9878 3469 9879
rect 3461 9874 3463 9878
rect 3467 9874 3469 9878
rect 3461 9873 3469 9874
rect 3461 9869 3463 9873
rect 3467 9869 3469 9873
rect 3461 9868 3469 9869
rect 3461 9864 3463 9868
rect 3467 9864 3469 9868
rect 3397 9863 3405 9864
rect 3397 9859 3399 9863
rect 3403 9859 3405 9863
rect 3397 9858 3405 9859
rect 3461 9863 3469 9864
rect 3461 9859 3463 9863
rect 3467 9859 3469 9863
rect 3461 9858 3469 9859
rect 3397 9856 3469 9858
rect 3397 9852 3399 9856
rect 3403 9852 3406 9856
rect 3410 9852 3411 9856
rect 3415 9852 3416 9856
rect 3420 9852 3421 9856
rect 3425 9852 3426 9856
rect 3430 9852 3431 9856
rect 3435 9852 3436 9856
rect 3440 9852 3441 9856
rect 3445 9852 3446 9856
rect 3450 9852 3451 9856
rect 3455 9852 3456 9856
rect 3460 9852 3463 9856
rect 3467 9852 3469 9856
rect 3397 9850 3469 9852
rect 3534 9978 3630 9979
rect 3534 9974 3535 9978
rect 3539 9974 3540 9978
rect 3544 9974 3545 9978
rect 3549 9974 3550 9978
rect 3554 9974 3555 9978
rect 3559 9974 3560 9978
rect 3564 9974 3565 9978
rect 3569 9974 3570 9978
rect 3574 9974 3575 9978
rect 3579 9974 3580 9978
rect 3584 9974 3585 9978
rect 3589 9974 3590 9978
rect 3594 9974 3595 9978
rect 3599 9974 3600 9978
rect 3604 9974 3605 9978
rect 3609 9974 3610 9978
rect 3614 9974 3615 9978
rect 3619 9974 3620 9978
rect 3624 9974 3625 9978
rect 3629 9974 3630 9978
rect 3534 9973 3630 9974
rect 3534 9969 3535 9973
rect 3539 9969 3540 9973
rect 3534 9968 3540 9969
rect 3534 9964 3535 9968
rect 3539 9964 3540 9968
rect 3624 9969 3625 9973
rect 3629 9969 3630 9973
rect 3624 9968 3630 9969
rect 3534 9963 3540 9964
rect 3534 9959 3535 9963
rect 3539 9959 3540 9963
rect 3534 9958 3540 9959
rect 3534 9954 3535 9958
rect 3539 9954 3540 9958
rect 3534 9953 3540 9954
rect 3534 9949 3535 9953
rect 3539 9949 3540 9953
rect 3534 9948 3540 9949
rect 3534 9944 3535 9948
rect 3539 9944 3540 9948
rect 3534 9943 3540 9944
rect 3534 9939 3535 9943
rect 3539 9939 3540 9943
rect 3534 9938 3540 9939
rect 3534 9934 3535 9938
rect 3539 9934 3540 9938
rect 3534 9933 3540 9934
rect 3534 9929 3535 9933
rect 3539 9929 3540 9933
rect 3534 9928 3540 9929
rect 3534 9924 3535 9928
rect 3539 9924 3540 9928
rect 3534 9923 3540 9924
rect 3534 9919 3535 9923
rect 3539 9919 3540 9923
rect 3534 9918 3540 9919
rect 3534 9914 3535 9918
rect 3539 9914 3540 9918
rect 3534 9913 3540 9914
rect 3534 9909 3535 9913
rect 3539 9909 3540 9913
rect 3534 9908 3540 9909
rect 3534 9904 3535 9908
rect 3539 9904 3540 9908
rect 3534 9903 3540 9904
rect 3534 9899 3535 9903
rect 3539 9899 3540 9903
rect 3534 9898 3540 9899
rect 3534 9894 3535 9898
rect 3539 9894 3540 9898
rect 3534 9893 3540 9894
rect 3534 9889 3535 9893
rect 3539 9889 3540 9893
rect 3534 9888 3540 9889
rect 3534 9884 3535 9888
rect 3539 9884 3540 9888
rect 3534 9883 3540 9884
rect 3534 9879 3535 9883
rect 3539 9879 3540 9883
rect 3534 9878 3540 9879
rect 3534 9874 3535 9878
rect 3539 9874 3540 9878
rect 3534 9873 3540 9874
rect 3534 9869 3535 9873
rect 3539 9869 3540 9873
rect 3534 9868 3540 9869
rect 3534 9864 3535 9868
rect 3539 9864 3540 9868
rect 3534 9863 3540 9864
rect 3534 9859 3535 9863
rect 3539 9859 3540 9863
rect 3534 9858 3540 9859
rect 3534 9854 3535 9858
rect 3539 9854 3540 9858
rect 3534 9853 3540 9854
rect 3534 9849 3535 9853
rect 3539 9849 3540 9853
rect 3624 9964 3625 9968
rect 3629 9964 3630 9968
rect 3624 9963 3630 9964
rect 3624 9959 3625 9963
rect 3629 9959 3630 9963
rect 3624 9958 3630 9959
rect 3624 9954 3625 9958
rect 3629 9954 3630 9958
rect 3624 9953 3630 9954
rect 3624 9949 3625 9953
rect 3629 9949 3630 9953
rect 3624 9948 3630 9949
rect 3624 9944 3625 9948
rect 3629 9944 3630 9948
rect 3624 9943 3630 9944
rect 3624 9939 3625 9943
rect 3629 9939 3630 9943
rect 3624 9938 3630 9939
rect 3624 9934 3625 9938
rect 3629 9934 3630 9938
rect 3624 9933 3630 9934
rect 3624 9929 3625 9933
rect 3629 9929 3630 9933
rect 3624 9928 3630 9929
rect 3624 9924 3625 9928
rect 3629 9924 3630 9928
rect 3624 9923 3630 9924
rect 3624 9919 3625 9923
rect 3629 9919 3630 9923
rect 3624 9918 3630 9919
rect 3624 9914 3625 9918
rect 3629 9914 3630 9918
rect 3624 9913 3630 9914
rect 3624 9909 3625 9913
rect 3629 9909 3630 9913
rect 3624 9908 3630 9909
rect 3624 9904 3625 9908
rect 3629 9904 3630 9908
rect 3624 9903 3630 9904
rect 3624 9899 3625 9903
rect 3629 9899 3630 9903
rect 3624 9898 3630 9899
rect 3624 9894 3625 9898
rect 3629 9894 3630 9898
rect 3624 9893 3630 9894
rect 3624 9889 3625 9893
rect 3629 9889 3630 9893
rect 3624 9888 3630 9889
rect 3624 9884 3625 9888
rect 3629 9884 3630 9888
rect 3624 9883 3630 9884
rect 3624 9879 3625 9883
rect 3629 9879 3630 9883
rect 3624 9878 3630 9879
rect 3624 9874 3625 9878
rect 3629 9874 3630 9878
rect 3624 9873 3630 9874
rect 3624 9869 3625 9873
rect 3629 9869 3630 9873
rect 3624 9868 3630 9869
rect 3624 9864 3625 9868
rect 3629 9864 3630 9868
rect 3624 9863 3630 9864
rect 3624 9859 3625 9863
rect 3629 9859 3630 9863
rect 3624 9858 3630 9859
rect 3624 9854 3625 9858
rect 3629 9854 3630 9858
rect 3624 9853 3630 9854
rect 3534 9848 3540 9849
rect 3534 9844 3535 9848
rect 3539 9844 3540 9848
rect 3624 9849 3625 9853
rect 3629 9849 3630 9853
rect 3624 9848 3630 9849
rect 3624 9844 3625 9848
rect 3629 9844 3630 9848
rect 3534 9843 3630 9844
rect 3534 9839 3535 9843
rect 3539 9839 3540 9843
rect 3544 9839 3545 9843
rect 3549 9839 3550 9843
rect 3554 9839 3555 9843
rect 3559 9839 3560 9843
rect 3564 9839 3565 9843
rect 3569 9839 3570 9843
rect 3574 9839 3575 9843
rect 3579 9839 3580 9843
rect 3584 9839 3585 9843
rect 3589 9839 3590 9843
rect 3594 9839 3595 9843
rect 3599 9839 3600 9843
rect 3604 9839 3605 9843
rect 3609 9839 3610 9843
rect 3614 9839 3615 9843
rect 3619 9839 3620 9843
rect 3624 9839 3625 9843
rect 3629 9839 3630 9843
rect 3534 9838 3630 9839
rect 3706 9965 3778 9967
rect 3706 9961 3708 9965
rect 3712 9961 3715 9965
rect 3719 9961 3720 9965
rect 3724 9961 3725 9965
rect 3729 9961 3730 9965
rect 3734 9961 3735 9965
rect 3739 9961 3740 9965
rect 3744 9961 3745 9965
rect 3749 9961 3750 9965
rect 3754 9961 3755 9965
rect 3759 9961 3760 9965
rect 3764 9961 3765 9965
rect 3769 9961 3772 9965
rect 3776 9961 3778 9965
rect 3706 9959 3778 9961
rect 3706 9958 3714 9959
rect 3706 9954 3708 9958
rect 3712 9954 3714 9958
rect 3706 9953 3714 9954
rect 3770 9958 3778 9959
rect 3770 9954 3772 9958
rect 3776 9954 3778 9958
rect 3770 9953 3778 9954
rect 3706 9949 3708 9953
rect 3712 9949 3714 9953
rect 3706 9948 3714 9949
rect 3706 9944 3708 9948
rect 3712 9944 3714 9948
rect 3706 9943 3714 9944
rect 3706 9939 3708 9943
rect 3712 9939 3714 9943
rect 3706 9938 3714 9939
rect 3706 9934 3708 9938
rect 3712 9934 3714 9938
rect 3706 9933 3714 9934
rect 3706 9929 3708 9933
rect 3712 9929 3714 9933
rect 3706 9928 3714 9929
rect 3706 9924 3708 9928
rect 3712 9924 3714 9928
rect 3706 9923 3714 9924
rect 3706 9919 3708 9923
rect 3712 9919 3714 9923
rect 3706 9918 3714 9919
rect 3706 9914 3708 9918
rect 3712 9914 3714 9918
rect 3706 9913 3714 9914
rect 3706 9909 3708 9913
rect 3712 9909 3714 9913
rect 3706 9908 3714 9909
rect 3706 9904 3708 9908
rect 3712 9904 3714 9908
rect 3706 9903 3714 9904
rect 3706 9899 3708 9903
rect 3712 9899 3714 9903
rect 3706 9898 3714 9899
rect 3706 9894 3708 9898
rect 3712 9894 3714 9898
rect 3706 9893 3714 9894
rect 3706 9889 3708 9893
rect 3712 9889 3714 9893
rect 3706 9888 3714 9889
rect 3706 9884 3708 9888
rect 3712 9884 3714 9888
rect 3706 9883 3714 9884
rect 3706 9879 3708 9883
rect 3712 9879 3714 9883
rect 3706 9878 3714 9879
rect 3706 9874 3708 9878
rect 3712 9874 3714 9878
rect 3706 9873 3714 9874
rect 3706 9869 3708 9873
rect 3712 9869 3714 9873
rect 3706 9868 3714 9869
rect 3706 9864 3708 9868
rect 3712 9864 3714 9868
rect 3770 9949 3772 9953
rect 3776 9949 3778 9953
rect 3770 9948 3778 9949
rect 3770 9944 3772 9948
rect 3776 9944 3778 9948
rect 3770 9943 3778 9944
rect 3770 9939 3772 9943
rect 3776 9939 3778 9943
rect 3770 9938 3778 9939
rect 3770 9934 3772 9938
rect 3776 9934 3778 9938
rect 3770 9933 3778 9934
rect 3770 9929 3772 9933
rect 3776 9929 3778 9933
rect 3770 9928 3778 9929
rect 3770 9924 3772 9928
rect 3776 9924 3778 9928
rect 3770 9923 3778 9924
rect 3770 9919 3772 9923
rect 3776 9919 3778 9923
rect 3770 9918 3778 9919
rect 3770 9914 3772 9918
rect 3776 9914 3778 9918
rect 3770 9913 3778 9914
rect 3770 9909 3772 9913
rect 3776 9909 3778 9913
rect 3770 9908 3778 9909
rect 3770 9904 3772 9908
rect 3776 9904 3778 9908
rect 3770 9903 3778 9904
rect 3770 9899 3772 9903
rect 3776 9899 3778 9903
rect 3770 9898 3778 9899
rect 3770 9894 3772 9898
rect 3776 9894 3778 9898
rect 3770 9893 3778 9894
rect 3770 9889 3772 9893
rect 3776 9889 3778 9893
rect 3770 9888 3778 9889
rect 3770 9884 3772 9888
rect 3776 9884 3778 9888
rect 3770 9883 3778 9884
rect 3770 9879 3772 9883
rect 3776 9879 3778 9883
rect 3770 9878 3778 9879
rect 3770 9874 3772 9878
rect 3776 9874 3778 9878
rect 3770 9873 3778 9874
rect 3770 9869 3772 9873
rect 3776 9869 3778 9873
rect 3770 9868 3778 9869
rect 3770 9864 3772 9868
rect 3776 9864 3778 9868
rect 3706 9863 3714 9864
rect 3706 9859 3708 9863
rect 3712 9859 3714 9863
rect 3706 9858 3714 9859
rect 3770 9863 3778 9864
rect 3770 9859 3772 9863
rect 3776 9859 3778 9863
rect 3770 9858 3778 9859
rect 3706 9856 3778 9858
rect 3706 9852 3708 9856
rect 3712 9852 3715 9856
rect 3719 9852 3720 9856
rect 3724 9852 3725 9856
rect 3729 9852 3730 9856
rect 3734 9852 3735 9856
rect 3739 9852 3740 9856
rect 3744 9852 3745 9856
rect 3749 9852 3750 9856
rect 3754 9852 3755 9856
rect 3759 9852 3760 9856
rect 3764 9852 3765 9856
rect 3769 9852 3772 9856
rect 3776 9852 3778 9856
rect 3706 9850 3778 9852
rect 3843 9978 3939 9979
rect 3843 9974 3844 9978
rect 3848 9974 3849 9978
rect 3853 9974 3854 9978
rect 3858 9974 3859 9978
rect 3863 9974 3864 9978
rect 3868 9974 3869 9978
rect 3873 9974 3874 9978
rect 3878 9974 3879 9978
rect 3883 9974 3884 9978
rect 3888 9974 3889 9978
rect 3893 9974 3894 9978
rect 3898 9974 3899 9978
rect 3903 9974 3904 9978
rect 3908 9974 3909 9978
rect 3913 9974 3914 9978
rect 3918 9974 3919 9978
rect 3923 9974 3924 9978
rect 3928 9974 3929 9978
rect 3933 9974 3934 9978
rect 3938 9974 3939 9978
rect 3843 9973 3939 9974
rect 3843 9969 3844 9973
rect 3848 9969 3849 9973
rect 3843 9968 3849 9969
rect 3843 9964 3844 9968
rect 3848 9964 3849 9968
rect 3933 9969 3934 9973
rect 3938 9969 3939 9973
rect 3933 9968 3939 9969
rect 3843 9963 3849 9964
rect 3843 9959 3844 9963
rect 3848 9959 3849 9963
rect 3843 9958 3849 9959
rect 3843 9954 3844 9958
rect 3848 9954 3849 9958
rect 3843 9953 3849 9954
rect 3843 9949 3844 9953
rect 3848 9949 3849 9953
rect 3843 9948 3849 9949
rect 3843 9944 3844 9948
rect 3848 9944 3849 9948
rect 3843 9943 3849 9944
rect 3843 9939 3844 9943
rect 3848 9939 3849 9943
rect 3843 9938 3849 9939
rect 3843 9934 3844 9938
rect 3848 9934 3849 9938
rect 3843 9933 3849 9934
rect 3843 9929 3844 9933
rect 3848 9929 3849 9933
rect 3843 9928 3849 9929
rect 3843 9924 3844 9928
rect 3848 9924 3849 9928
rect 3843 9923 3849 9924
rect 3843 9919 3844 9923
rect 3848 9919 3849 9923
rect 3843 9918 3849 9919
rect 3843 9914 3844 9918
rect 3848 9914 3849 9918
rect 3843 9913 3849 9914
rect 3843 9909 3844 9913
rect 3848 9909 3849 9913
rect 3843 9908 3849 9909
rect 3843 9904 3844 9908
rect 3848 9904 3849 9908
rect 3843 9903 3849 9904
rect 3843 9899 3844 9903
rect 3848 9899 3849 9903
rect 3843 9898 3849 9899
rect 3843 9894 3844 9898
rect 3848 9894 3849 9898
rect 3843 9893 3849 9894
rect 3843 9889 3844 9893
rect 3848 9889 3849 9893
rect 3843 9888 3849 9889
rect 3843 9884 3844 9888
rect 3848 9884 3849 9888
rect 3843 9883 3849 9884
rect 3843 9879 3844 9883
rect 3848 9879 3849 9883
rect 3843 9878 3849 9879
rect 3843 9874 3844 9878
rect 3848 9874 3849 9878
rect 3843 9873 3849 9874
rect 3843 9869 3844 9873
rect 3848 9869 3849 9873
rect 3843 9868 3849 9869
rect 3843 9864 3844 9868
rect 3848 9864 3849 9868
rect 3843 9863 3849 9864
rect 3843 9859 3844 9863
rect 3848 9859 3849 9863
rect 3843 9858 3849 9859
rect 3843 9854 3844 9858
rect 3848 9854 3849 9858
rect 3843 9853 3849 9854
rect 3843 9849 3844 9853
rect 3848 9849 3849 9853
rect 3933 9964 3934 9968
rect 3938 9964 3939 9968
rect 3933 9963 3939 9964
rect 3933 9959 3934 9963
rect 3938 9959 3939 9963
rect 3933 9958 3939 9959
rect 3933 9954 3934 9958
rect 3938 9954 3939 9958
rect 3933 9953 3939 9954
rect 3933 9949 3934 9953
rect 3938 9949 3939 9953
rect 3933 9948 3939 9949
rect 3933 9944 3934 9948
rect 3938 9944 3939 9948
rect 3933 9943 3939 9944
rect 3933 9939 3934 9943
rect 3938 9939 3939 9943
rect 3933 9938 3939 9939
rect 3933 9934 3934 9938
rect 3938 9934 3939 9938
rect 3933 9933 3939 9934
rect 3933 9929 3934 9933
rect 3938 9929 3939 9933
rect 3933 9928 3939 9929
rect 3933 9924 3934 9928
rect 3938 9924 3939 9928
rect 3933 9923 3939 9924
rect 3933 9919 3934 9923
rect 3938 9919 3939 9923
rect 3933 9918 3939 9919
rect 3933 9914 3934 9918
rect 3938 9914 3939 9918
rect 3933 9913 3939 9914
rect 3933 9909 3934 9913
rect 3938 9909 3939 9913
rect 3933 9908 3939 9909
rect 3933 9904 3934 9908
rect 3938 9904 3939 9908
rect 3933 9903 3939 9904
rect 3933 9899 3934 9903
rect 3938 9899 3939 9903
rect 3933 9898 3939 9899
rect 3933 9894 3934 9898
rect 3938 9894 3939 9898
rect 3933 9893 3939 9894
rect 3933 9889 3934 9893
rect 3938 9889 3939 9893
rect 3933 9888 3939 9889
rect 3933 9884 3934 9888
rect 3938 9884 3939 9888
rect 3933 9883 3939 9884
rect 3933 9879 3934 9883
rect 3938 9879 3939 9883
rect 3933 9878 3939 9879
rect 3933 9874 3934 9878
rect 3938 9874 3939 9878
rect 3933 9873 3939 9874
rect 3933 9869 3934 9873
rect 3938 9869 3939 9873
rect 3933 9868 3939 9869
rect 3933 9864 3934 9868
rect 3938 9864 3939 9868
rect 3933 9863 3939 9864
rect 3933 9859 3934 9863
rect 3938 9859 3939 9863
rect 3933 9858 3939 9859
rect 3933 9854 3934 9858
rect 3938 9854 3939 9858
rect 3933 9853 3939 9854
rect 3843 9848 3849 9849
rect 3843 9844 3844 9848
rect 3848 9844 3849 9848
rect 3933 9849 3934 9853
rect 3938 9849 3939 9853
rect 3933 9848 3939 9849
rect 3933 9844 3934 9848
rect 3938 9844 3939 9848
rect 3843 9843 3939 9844
rect 3843 9839 3844 9843
rect 3848 9839 3849 9843
rect 3853 9839 3854 9843
rect 3858 9839 3859 9843
rect 3863 9839 3864 9843
rect 3868 9839 3869 9843
rect 3873 9839 3874 9843
rect 3878 9839 3879 9843
rect 3883 9839 3884 9843
rect 3888 9839 3889 9843
rect 3893 9839 3894 9843
rect 3898 9839 3899 9843
rect 3903 9839 3904 9843
rect 3908 9839 3909 9843
rect 3913 9839 3914 9843
rect 3918 9839 3919 9843
rect 3923 9839 3924 9843
rect 3928 9839 3929 9843
rect 3933 9839 3934 9843
rect 3938 9839 3939 9843
rect 3843 9838 3939 9839
rect 4015 9965 4087 9967
rect 4015 9961 4017 9965
rect 4021 9961 4024 9965
rect 4028 9961 4029 9965
rect 4033 9961 4034 9965
rect 4038 9961 4039 9965
rect 4043 9961 4044 9965
rect 4048 9961 4049 9965
rect 4053 9961 4054 9965
rect 4058 9961 4059 9965
rect 4063 9961 4064 9965
rect 4068 9961 4069 9965
rect 4073 9961 4074 9965
rect 4078 9961 4081 9965
rect 4085 9961 4087 9965
rect 4015 9959 4087 9961
rect 4015 9958 4023 9959
rect 4015 9954 4017 9958
rect 4021 9954 4023 9958
rect 4015 9953 4023 9954
rect 4079 9958 4087 9959
rect 4079 9954 4081 9958
rect 4085 9954 4087 9958
rect 4079 9953 4087 9954
rect 4015 9949 4017 9953
rect 4021 9949 4023 9953
rect 4015 9948 4023 9949
rect 4015 9944 4017 9948
rect 4021 9944 4023 9948
rect 4015 9943 4023 9944
rect 4015 9939 4017 9943
rect 4021 9939 4023 9943
rect 4015 9938 4023 9939
rect 4015 9934 4017 9938
rect 4021 9934 4023 9938
rect 4015 9933 4023 9934
rect 4015 9929 4017 9933
rect 4021 9929 4023 9933
rect 4015 9928 4023 9929
rect 4015 9924 4017 9928
rect 4021 9924 4023 9928
rect 4015 9923 4023 9924
rect 4015 9919 4017 9923
rect 4021 9919 4023 9923
rect 4015 9918 4023 9919
rect 4015 9914 4017 9918
rect 4021 9914 4023 9918
rect 4015 9913 4023 9914
rect 4015 9909 4017 9913
rect 4021 9909 4023 9913
rect 4015 9908 4023 9909
rect 4015 9904 4017 9908
rect 4021 9904 4023 9908
rect 4015 9903 4023 9904
rect 4015 9899 4017 9903
rect 4021 9899 4023 9903
rect 4015 9898 4023 9899
rect 4015 9894 4017 9898
rect 4021 9894 4023 9898
rect 4015 9893 4023 9894
rect 4015 9889 4017 9893
rect 4021 9889 4023 9893
rect 4015 9888 4023 9889
rect 4015 9884 4017 9888
rect 4021 9884 4023 9888
rect 4015 9883 4023 9884
rect 4015 9879 4017 9883
rect 4021 9879 4023 9883
rect 4015 9878 4023 9879
rect 4015 9874 4017 9878
rect 4021 9874 4023 9878
rect 4015 9873 4023 9874
rect 4015 9869 4017 9873
rect 4021 9869 4023 9873
rect 4015 9868 4023 9869
rect 4015 9864 4017 9868
rect 4021 9864 4023 9868
rect 4079 9949 4081 9953
rect 4085 9949 4087 9953
rect 4079 9948 4087 9949
rect 4079 9944 4081 9948
rect 4085 9944 4087 9948
rect 4079 9943 4087 9944
rect 4079 9939 4081 9943
rect 4085 9939 4087 9943
rect 4079 9938 4087 9939
rect 4079 9934 4081 9938
rect 4085 9934 4087 9938
rect 4079 9933 4087 9934
rect 4079 9929 4081 9933
rect 4085 9929 4087 9933
rect 4079 9928 4087 9929
rect 4079 9924 4081 9928
rect 4085 9924 4087 9928
rect 4079 9923 4087 9924
rect 4079 9919 4081 9923
rect 4085 9919 4087 9923
rect 4079 9918 4087 9919
rect 4079 9914 4081 9918
rect 4085 9914 4087 9918
rect 4079 9913 4087 9914
rect 4079 9909 4081 9913
rect 4085 9909 4087 9913
rect 4079 9908 4087 9909
rect 4079 9904 4081 9908
rect 4085 9904 4087 9908
rect 4079 9903 4087 9904
rect 4079 9899 4081 9903
rect 4085 9899 4087 9903
rect 4079 9898 4087 9899
rect 4079 9894 4081 9898
rect 4085 9894 4087 9898
rect 4079 9893 4087 9894
rect 4079 9889 4081 9893
rect 4085 9889 4087 9893
rect 4079 9888 4087 9889
rect 4079 9884 4081 9888
rect 4085 9884 4087 9888
rect 4079 9883 4087 9884
rect 4079 9879 4081 9883
rect 4085 9879 4087 9883
rect 4079 9878 4087 9879
rect 4079 9874 4081 9878
rect 4085 9874 4087 9878
rect 4079 9873 4087 9874
rect 4079 9869 4081 9873
rect 4085 9869 4087 9873
rect 4079 9868 4087 9869
rect 4079 9864 4081 9868
rect 4085 9864 4087 9868
rect 4015 9863 4023 9864
rect 4015 9859 4017 9863
rect 4021 9859 4023 9863
rect 4015 9858 4023 9859
rect 4079 9863 4087 9864
rect 4079 9859 4081 9863
rect 4085 9859 4087 9863
rect 4079 9858 4087 9859
rect 4015 9856 4087 9858
rect 4015 9852 4017 9856
rect 4021 9852 4024 9856
rect 4028 9852 4029 9856
rect 4033 9852 4034 9856
rect 4038 9852 4039 9856
rect 4043 9852 4044 9856
rect 4048 9852 4049 9856
rect 4053 9852 4054 9856
rect 4058 9852 4059 9856
rect 4063 9852 4064 9856
rect 4068 9852 4069 9856
rect 4073 9852 4074 9856
rect 4078 9852 4081 9856
rect 4085 9852 4087 9856
rect 4015 9850 4087 9852
rect 609 9766 4563 9770
rect 609 9762 802 9766
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 821 9762 831 9766
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 850 9762 860 9766
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 879 9762 889 9766
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 908 9762 918 9766
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 937 9762 1319 9766
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1338 9762 1628 9766
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1647 9762 1937 9766
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1956 9762 2246 9766
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2265 9762 2555 9766
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2574 9762 2864 9766
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2883 9762 3173 9766
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3192 9762 3482 9766
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3501 9762 3791 9766
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3810 9762 4100 9766
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4119 9762 4292 9766
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4311 9762 4318 9766
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4337 9762 4344 9766
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4363 9762 4370 9766
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4389 9762 4396 9766
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4415 9762 4563 9766
rect 609 9756 4563 9762
rect 609 9752 802 9756
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 821 9752 831 9756
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 850 9752 860 9756
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 879 9752 889 9756
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 908 9752 918 9756
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 937 9752 1319 9756
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1338 9752 1628 9756
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1647 9752 1937 9756
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1956 9752 2246 9756
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2265 9752 2555 9756
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2574 9752 2864 9756
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2883 9752 3173 9756
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3192 9752 3482 9756
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3501 9752 3791 9756
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3810 9752 4100 9756
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4119 9752 4292 9756
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4311 9752 4318 9756
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4337 9752 4344 9756
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4363 9752 4370 9756
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4389 9752 4396 9756
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4415 9752 4563 9756
rect 609 9746 4563 9752
rect 609 9742 802 9746
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 821 9742 831 9746
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 850 9742 860 9746
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 879 9742 889 9746
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 908 9742 918 9746
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 937 9742 1319 9746
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1338 9742 1628 9746
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1647 9742 1937 9746
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1956 9742 2246 9746
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2265 9742 2555 9746
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2574 9742 2864 9746
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2883 9742 3173 9746
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3192 9742 3482 9746
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3501 9742 3791 9746
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3810 9742 4100 9746
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4119 9742 4292 9746
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4311 9742 4318 9746
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4337 9742 4344 9746
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4363 9742 4370 9746
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4389 9742 4396 9746
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4415 9742 4563 9746
rect 609 9736 4563 9742
rect 609 9732 802 9736
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 821 9732 831 9736
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 850 9732 860 9736
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 879 9732 889 9736
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 908 9732 918 9736
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 937 9732 1319 9736
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1338 9732 1628 9736
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1647 9732 1937 9736
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1956 9732 2246 9736
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2265 9732 2555 9736
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2574 9732 2864 9736
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2883 9732 3173 9736
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3192 9732 3482 9736
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3501 9732 3791 9736
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3810 9732 4100 9736
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4119 9732 4292 9736
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4311 9732 4318 9736
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4337 9732 4344 9736
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4363 9732 4370 9736
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4389 9732 4396 9736
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 4415 9732 4563 9736
rect 609 9730 4563 9732
rect 609 9622 649 9730
rect 609 9618 613 9622
rect 617 9618 623 9622
rect 627 9618 633 9622
rect 637 9618 643 9622
rect 647 9618 649 9622
rect 609 9617 649 9618
rect 609 9613 613 9617
rect 617 9613 623 9617
rect 627 9613 633 9617
rect 637 9613 643 9617
rect 647 9613 649 9617
rect 609 9612 649 9613
rect 609 9608 613 9612
rect 617 9608 623 9612
rect 627 9608 633 9612
rect 637 9608 643 9612
rect 647 9608 649 9612
rect 609 9607 649 9608
rect 609 9603 613 9607
rect 617 9603 623 9607
rect 627 9603 633 9607
rect 637 9603 643 9607
rect 647 9603 649 9607
rect 609 9596 649 9603
rect 609 9592 613 9596
rect 617 9592 623 9596
rect 627 9592 633 9596
rect 637 9592 643 9596
rect 647 9592 649 9596
rect 609 9591 649 9592
rect 609 9587 613 9591
rect 617 9587 623 9591
rect 627 9587 633 9591
rect 637 9587 643 9591
rect 647 9587 649 9591
rect 609 9586 649 9587
rect 609 9582 613 9586
rect 617 9582 623 9586
rect 627 9582 633 9586
rect 637 9582 643 9586
rect 647 9582 649 9586
rect 609 9581 649 9582
rect 609 9577 613 9581
rect 617 9577 623 9581
rect 627 9577 633 9581
rect 637 9577 643 9581
rect 647 9577 649 9581
rect 609 9570 649 9577
rect 609 9566 613 9570
rect 617 9566 623 9570
rect 627 9566 633 9570
rect 637 9566 643 9570
rect 647 9566 649 9570
rect 609 9565 649 9566
rect 609 9561 613 9565
rect 617 9561 623 9565
rect 627 9561 633 9565
rect 637 9561 643 9565
rect 647 9561 649 9565
rect 609 9560 649 9561
rect 609 9556 613 9560
rect 617 9556 623 9560
rect 627 9556 633 9560
rect 637 9556 643 9560
rect 647 9556 649 9560
rect 609 9555 649 9556
rect 609 9551 613 9555
rect 617 9551 623 9555
rect 627 9551 633 9555
rect 637 9551 643 9555
rect 647 9551 649 9555
rect 609 9544 649 9551
rect 609 9540 613 9544
rect 617 9540 623 9544
rect 627 9540 633 9544
rect 637 9540 643 9544
rect 647 9540 649 9544
rect 609 9539 649 9540
rect 609 9535 613 9539
rect 617 9535 623 9539
rect 627 9535 633 9539
rect 637 9535 643 9539
rect 647 9535 649 9539
rect 609 9534 649 9535
rect 609 9530 613 9534
rect 617 9530 623 9534
rect 627 9530 633 9534
rect 637 9530 643 9534
rect 647 9530 649 9534
rect 609 9529 649 9530
rect 609 9525 613 9529
rect 617 9525 623 9529
rect 627 9525 633 9529
rect 637 9525 643 9529
rect 647 9525 649 9529
rect 609 9518 649 9525
rect 609 9514 613 9518
rect 617 9514 623 9518
rect 627 9514 633 9518
rect 637 9514 643 9518
rect 647 9514 649 9518
rect 609 9513 649 9514
rect 609 9509 613 9513
rect 617 9509 623 9513
rect 627 9509 633 9513
rect 637 9509 643 9513
rect 647 9509 649 9513
rect 609 9508 649 9509
rect 609 9504 613 9508
rect 617 9504 623 9508
rect 627 9504 633 9508
rect 637 9504 643 9508
rect 647 9504 649 9508
rect 609 9503 649 9504
rect 609 9499 613 9503
rect 617 9499 623 9503
rect 627 9499 633 9503
rect 637 9499 643 9503
rect 647 9499 649 9503
rect 609 9325 649 9499
rect 609 9321 613 9325
rect 617 9321 623 9325
rect 627 9321 633 9325
rect 637 9321 643 9325
rect 647 9321 649 9325
rect 609 9320 649 9321
rect 609 9316 613 9320
rect 617 9316 623 9320
rect 627 9316 633 9320
rect 637 9316 643 9320
rect 647 9316 649 9320
rect 609 9315 649 9316
rect 609 9311 613 9315
rect 617 9311 623 9315
rect 627 9311 633 9315
rect 637 9311 643 9315
rect 647 9311 649 9315
rect 609 9310 649 9311
rect 609 9306 613 9310
rect 617 9306 623 9310
rect 627 9306 633 9310
rect 637 9306 643 9310
rect 647 9306 649 9310
rect 609 9016 649 9306
rect 609 9012 613 9016
rect 617 9012 623 9016
rect 627 9012 633 9016
rect 637 9012 643 9016
rect 647 9012 649 9016
rect 609 9011 649 9012
rect 609 9007 613 9011
rect 617 9007 623 9011
rect 627 9007 633 9011
rect 637 9007 643 9011
rect 647 9007 649 9011
rect 609 9006 649 9007
rect 609 9002 613 9006
rect 617 9002 623 9006
rect 627 9002 633 9006
rect 637 9002 643 9006
rect 647 9002 649 9006
rect 609 9001 649 9002
rect 609 8997 613 9001
rect 617 8997 623 9001
rect 627 8997 633 9001
rect 637 8997 643 9001
rect 647 8997 649 9001
rect 609 8707 649 8997
rect 609 8703 613 8707
rect 617 8703 623 8707
rect 627 8703 633 8707
rect 637 8703 643 8707
rect 647 8703 649 8707
rect 609 8702 649 8703
rect 609 8698 613 8702
rect 617 8698 623 8702
rect 627 8698 633 8702
rect 637 8698 643 8702
rect 647 8698 649 8702
rect 609 8697 649 8698
rect 609 8693 613 8697
rect 617 8693 623 8697
rect 627 8693 633 8697
rect 637 8693 643 8697
rect 647 8693 649 8697
rect 609 8692 649 8693
rect 609 8688 613 8692
rect 617 8688 623 8692
rect 627 8688 633 8692
rect 637 8688 643 8692
rect 647 8688 649 8692
rect 609 8398 649 8688
rect 609 8394 613 8398
rect 617 8394 623 8398
rect 627 8394 633 8398
rect 637 8394 643 8398
rect 647 8394 649 8398
rect 609 8393 649 8394
rect 609 8389 613 8393
rect 617 8389 623 8393
rect 627 8389 633 8393
rect 637 8389 643 8393
rect 647 8389 649 8393
rect 609 8388 649 8389
rect 609 8384 613 8388
rect 617 8384 623 8388
rect 627 8384 633 8388
rect 637 8384 643 8388
rect 647 8384 649 8388
rect 609 8383 649 8384
rect 609 8379 613 8383
rect 617 8379 623 8383
rect 627 8379 633 8383
rect 637 8379 643 8383
rect 647 8379 649 8383
rect 609 8089 649 8379
rect 609 8085 613 8089
rect 617 8085 623 8089
rect 627 8085 633 8089
rect 637 8085 643 8089
rect 647 8085 649 8089
rect 609 8084 649 8085
rect 609 8080 613 8084
rect 617 8080 623 8084
rect 627 8080 633 8084
rect 637 8080 643 8084
rect 647 8080 649 8084
rect 609 8079 649 8080
rect 609 8075 613 8079
rect 617 8075 623 8079
rect 627 8075 633 8079
rect 637 8075 643 8079
rect 647 8075 649 8079
rect 609 8074 649 8075
rect 609 8070 613 8074
rect 617 8070 623 8074
rect 627 8070 633 8074
rect 637 8070 643 8074
rect 647 8070 649 8074
rect 609 7780 649 8070
rect 609 7776 613 7780
rect 617 7776 623 7780
rect 627 7776 633 7780
rect 637 7776 643 7780
rect 647 7776 649 7780
rect 609 7775 649 7776
rect 609 7771 613 7775
rect 617 7771 623 7775
rect 627 7771 633 7775
rect 637 7771 643 7775
rect 647 7771 649 7775
rect 609 7770 649 7771
rect 609 7766 613 7770
rect 617 7766 623 7770
rect 627 7766 633 7770
rect 637 7766 643 7770
rect 647 7766 649 7770
rect 609 7765 649 7766
rect 609 7761 613 7765
rect 617 7761 623 7765
rect 627 7761 633 7765
rect 637 7761 643 7765
rect 647 7761 649 7765
rect 609 7471 649 7761
rect 609 7467 613 7471
rect 617 7467 623 7471
rect 627 7467 633 7471
rect 637 7467 643 7471
rect 647 7467 649 7471
rect 609 7466 649 7467
rect 609 7462 613 7466
rect 617 7462 623 7466
rect 627 7462 633 7466
rect 637 7462 643 7466
rect 647 7462 649 7466
rect 609 7461 649 7462
rect 609 7457 613 7461
rect 617 7457 623 7461
rect 627 7457 633 7461
rect 637 7457 643 7461
rect 647 7457 649 7461
rect 609 7456 649 7457
rect 609 7452 613 7456
rect 617 7452 623 7456
rect 627 7452 633 7456
rect 637 7452 643 7456
rect 647 7452 649 7456
rect 609 7162 649 7452
rect 609 7158 613 7162
rect 617 7158 623 7162
rect 627 7158 633 7162
rect 637 7158 643 7162
rect 647 7158 649 7162
rect 609 7127 649 7158
rect 609 7123 613 7127
rect 617 7123 623 7127
rect 627 7123 633 7127
rect 637 7123 643 7127
rect 647 7123 649 7127
rect 609 7122 649 7123
rect 609 7118 613 7122
rect 617 7118 623 7122
rect 627 7118 633 7122
rect 637 7118 643 7122
rect 647 7118 649 7122
rect 609 7117 649 7118
rect 609 7113 613 7117
rect 617 7113 623 7117
rect 627 7113 633 7117
rect 637 7113 643 7117
rect 647 7113 649 7117
rect 609 7112 649 7113
rect 609 7108 613 7112
rect 617 7108 623 7112
rect 627 7108 633 7112
rect 637 7108 643 7112
rect 647 7108 649 7112
rect 609 6540 649 7108
rect 609 6536 613 6540
rect 617 6536 623 6540
rect 627 6536 633 6540
rect 637 6536 643 6540
rect 647 6536 649 6540
rect 609 6535 649 6536
rect 609 6531 613 6535
rect 617 6531 623 6535
rect 627 6531 633 6535
rect 637 6531 643 6535
rect 647 6531 649 6535
rect 609 6530 649 6531
rect 609 6526 613 6530
rect 617 6526 623 6530
rect 627 6526 633 6530
rect 637 6526 643 6530
rect 647 6526 649 6530
rect 609 6525 649 6526
rect 609 6521 613 6525
rect 617 6521 623 6525
rect 627 6521 633 6525
rect 637 6521 643 6525
rect 647 6521 649 6525
rect 609 6231 649 6521
rect 609 6227 613 6231
rect 617 6227 623 6231
rect 627 6227 633 6231
rect 637 6227 643 6231
rect 647 6227 649 6231
rect 609 6226 649 6227
rect 609 6222 613 6226
rect 617 6222 623 6226
rect 627 6222 633 6226
rect 637 6222 643 6226
rect 647 6222 649 6226
rect 609 6221 649 6222
rect 609 6217 613 6221
rect 617 6217 623 6221
rect 627 6217 633 6221
rect 637 6217 643 6221
rect 647 6217 649 6221
rect 609 6216 649 6217
rect 609 6212 613 6216
rect 617 6212 623 6216
rect 627 6212 633 6216
rect 637 6212 643 6216
rect 647 6212 649 6216
rect 609 6200 649 6212
rect 609 6196 613 6200
rect 617 6196 623 6200
rect 627 6196 633 6200
rect 637 6196 643 6200
rect 647 6196 649 6200
rect 609 6195 649 6196
rect 609 6191 613 6195
rect 617 6191 623 6195
rect 627 6191 633 6195
rect 637 6191 643 6195
rect 647 6191 649 6195
rect 609 6190 649 6191
rect 609 6186 613 6190
rect 617 6186 623 6190
rect 627 6186 633 6190
rect 637 6186 643 6190
rect 647 6186 649 6190
rect 609 6185 649 6186
rect 609 6181 613 6185
rect 617 6181 623 6185
rect 627 6181 633 6185
rect 637 6181 643 6185
rect 647 6181 649 6185
rect 609 5891 649 6181
rect 609 5887 613 5891
rect 617 5887 623 5891
rect 627 5887 633 5891
rect 637 5887 643 5891
rect 647 5887 649 5891
rect 609 5886 649 5887
rect 609 5882 613 5886
rect 617 5882 623 5886
rect 627 5882 633 5886
rect 637 5882 643 5886
rect 647 5882 649 5886
rect 609 5881 649 5882
rect 609 5877 613 5881
rect 617 5877 623 5881
rect 627 5877 633 5881
rect 637 5877 643 5881
rect 647 5877 649 5881
rect 609 5876 649 5877
rect 609 5872 613 5876
rect 617 5872 623 5876
rect 627 5872 633 5876
rect 637 5872 643 5876
rect 647 5872 649 5876
rect 609 5582 649 5872
rect 609 5578 613 5582
rect 617 5578 623 5582
rect 627 5578 633 5582
rect 637 5578 643 5582
rect 647 5578 649 5582
rect 609 5577 649 5578
rect 609 5573 613 5577
rect 617 5573 623 5577
rect 627 5573 633 5577
rect 637 5573 643 5577
rect 647 5573 649 5577
rect 609 5572 649 5573
rect 609 5568 613 5572
rect 617 5568 623 5572
rect 627 5568 633 5572
rect 637 5568 643 5572
rect 647 5568 649 5572
rect 609 5567 649 5568
rect 609 5563 613 5567
rect 617 5563 623 5567
rect 627 5563 633 5567
rect 637 5563 643 5567
rect 647 5563 649 5567
rect 609 5273 649 5563
rect 609 5269 613 5273
rect 617 5269 623 5273
rect 627 5269 633 5273
rect 637 5269 643 5273
rect 647 5269 649 5273
rect 609 5268 649 5269
rect 609 5264 613 5268
rect 617 5264 623 5268
rect 627 5264 633 5268
rect 637 5264 643 5268
rect 647 5264 649 5268
rect 609 5263 649 5264
rect 609 5259 613 5263
rect 617 5259 623 5263
rect 627 5259 633 5263
rect 637 5259 643 5263
rect 647 5259 649 5263
rect 609 5258 649 5259
rect 609 5254 613 5258
rect 617 5254 623 5258
rect 627 5254 633 5258
rect 637 5254 643 5258
rect 647 5254 649 5258
rect 609 4872 649 5254
rect 609 4868 613 4872
rect 617 4868 623 4872
rect 627 4868 633 4872
rect 637 4868 643 4872
rect 647 4868 649 4872
rect 609 4867 649 4868
rect 609 4863 613 4867
rect 617 4863 623 4867
rect 627 4863 633 4867
rect 637 4863 643 4867
rect 647 4863 649 4867
rect 609 4862 649 4863
rect 609 4858 613 4862
rect 617 4858 623 4862
rect 627 4858 633 4862
rect 637 4858 643 4862
rect 647 4858 649 4862
rect 609 4857 649 4858
rect 609 4853 613 4857
rect 617 4853 623 4857
rect 627 4853 633 4857
rect 637 4853 643 4857
rect 647 4853 649 4857
rect 609 4843 649 4853
rect 609 4839 613 4843
rect 617 4839 623 4843
rect 627 4839 633 4843
rect 637 4839 643 4843
rect 647 4839 649 4843
rect 609 4838 649 4839
rect 609 4834 613 4838
rect 617 4834 623 4838
rect 627 4834 633 4838
rect 637 4834 643 4838
rect 647 4834 649 4838
rect 609 4833 649 4834
rect 609 4829 613 4833
rect 617 4829 623 4833
rect 627 4829 633 4833
rect 637 4829 643 4833
rect 647 4829 649 4833
rect 609 4828 649 4829
rect 609 4824 613 4828
rect 617 4824 623 4828
rect 627 4824 633 4828
rect 637 4824 643 4828
rect 647 4824 649 4828
rect 609 4814 649 4824
rect 609 4810 613 4814
rect 617 4810 623 4814
rect 627 4810 633 4814
rect 637 4810 643 4814
rect 647 4810 649 4814
rect 609 4809 649 4810
rect 609 4805 613 4809
rect 617 4805 623 4809
rect 627 4805 633 4809
rect 637 4805 643 4809
rect 647 4805 649 4809
rect 609 4804 649 4805
rect 609 4800 613 4804
rect 617 4800 623 4804
rect 627 4800 633 4804
rect 637 4800 643 4804
rect 647 4800 649 4804
rect 609 4799 649 4800
rect 609 4795 613 4799
rect 617 4795 623 4799
rect 627 4795 633 4799
rect 637 4795 643 4799
rect 647 4795 649 4799
rect 609 4785 649 4795
rect 609 4781 613 4785
rect 617 4781 623 4785
rect 627 4781 633 4785
rect 637 4781 643 4785
rect 647 4781 649 4785
rect 609 4780 649 4781
rect 609 4776 613 4780
rect 617 4776 623 4780
rect 627 4776 633 4780
rect 637 4776 643 4780
rect 647 4776 649 4780
rect 609 4775 649 4776
rect 609 4771 613 4775
rect 617 4771 623 4775
rect 627 4771 633 4775
rect 637 4771 643 4775
rect 647 4771 649 4775
rect 609 4770 649 4771
rect 609 4766 613 4770
rect 617 4766 623 4770
rect 627 4766 633 4770
rect 637 4766 643 4770
rect 647 4766 649 4770
rect 609 4756 649 4766
rect 609 4752 613 4756
rect 617 4752 623 4756
rect 627 4752 633 4756
rect 637 4752 643 4756
rect 647 4752 649 4756
rect 609 4751 649 4752
rect 609 4747 613 4751
rect 617 4747 623 4751
rect 627 4747 633 4751
rect 637 4747 643 4751
rect 647 4747 649 4751
rect 609 4746 649 4747
rect 609 4742 613 4746
rect 617 4742 623 4746
rect 627 4742 633 4746
rect 637 4742 643 4746
rect 647 4742 649 4746
rect 609 4741 649 4742
rect 609 4737 613 4741
rect 617 4737 623 4741
rect 627 4737 633 4741
rect 637 4737 643 4741
rect 647 4737 649 4741
rect 609 4584 649 4737
rect 4523 9577 4563 9730
rect 4523 9573 4525 9577
rect 4529 9573 4535 9577
rect 4539 9573 4545 9577
rect 4549 9573 4555 9577
rect 4559 9573 4563 9577
rect 4523 9572 4563 9573
rect 4523 9568 4525 9572
rect 4529 9568 4535 9572
rect 4539 9568 4545 9572
rect 4549 9568 4555 9572
rect 4559 9568 4563 9572
rect 4523 9567 4563 9568
rect 4523 9563 4525 9567
rect 4529 9563 4535 9567
rect 4539 9563 4545 9567
rect 4549 9563 4555 9567
rect 4559 9563 4563 9567
rect 4523 9562 4563 9563
rect 4523 9558 4525 9562
rect 4529 9558 4535 9562
rect 4539 9558 4545 9562
rect 4549 9558 4555 9562
rect 4559 9558 4563 9562
rect 4523 9548 4563 9558
rect 4523 9544 4525 9548
rect 4529 9544 4535 9548
rect 4539 9544 4545 9548
rect 4549 9544 4555 9548
rect 4559 9544 4563 9548
rect 4523 9543 4563 9544
rect 4523 9539 4525 9543
rect 4529 9539 4535 9543
rect 4539 9539 4545 9543
rect 4549 9539 4555 9543
rect 4559 9539 4563 9543
rect 4523 9538 4563 9539
rect 4523 9534 4525 9538
rect 4529 9534 4535 9538
rect 4539 9534 4545 9538
rect 4549 9534 4555 9538
rect 4559 9534 4563 9538
rect 4523 9533 4563 9534
rect 4523 9529 4525 9533
rect 4529 9529 4535 9533
rect 4539 9529 4545 9533
rect 4549 9529 4555 9533
rect 4559 9529 4563 9533
rect 4523 9519 4563 9529
rect 4523 9515 4525 9519
rect 4529 9515 4535 9519
rect 4539 9515 4545 9519
rect 4549 9515 4555 9519
rect 4559 9515 4563 9519
rect 4523 9514 4563 9515
rect 4523 9510 4525 9514
rect 4529 9510 4535 9514
rect 4539 9510 4545 9514
rect 4549 9510 4555 9514
rect 4559 9510 4563 9514
rect 4523 9509 4563 9510
rect 4523 9505 4525 9509
rect 4529 9505 4535 9509
rect 4539 9505 4545 9509
rect 4549 9505 4555 9509
rect 4559 9505 4563 9509
rect 4523 9504 4563 9505
rect 4523 9500 4525 9504
rect 4529 9500 4535 9504
rect 4539 9500 4545 9504
rect 4549 9500 4555 9504
rect 4559 9500 4563 9504
rect 4523 9490 4563 9500
rect 4523 9486 4525 9490
rect 4529 9486 4535 9490
rect 4539 9486 4545 9490
rect 4549 9486 4555 9490
rect 4559 9486 4563 9490
rect 4523 9485 4563 9486
rect 4523 9481 4525 9485
rect 4529 9481 4535 9485
rect 4539 9481 4545 9485
rect 4549 9481 4555 9485
rect 4559 9481 4563 9485
rect 4523 9480 4563 9481
rect 4523 9476 4525 9480
rect 4529 9476 4535 9480
rect 4539 9476 4545 9480
rect 4549 9476 4555 9480
rect 4559 9476 4563 9480
rect 4523 9475 4563 9476
rect 4523 9471 4525 9475
rect 4529 9471 4535 9475
rect 4539 9471 4545 9475
rect 4549 9471 4555 9475
rect 4559 9471 4563 9475
rect 4523 9461 4563 9471
rect 4523 9457 4525 9461
rect 4529 9457 4535 9461
rect 4539 9457 4545 9461
rect 4549 9457 4555 9461
rect 4559 9457 4563 9461
rect 4523 9456 4563 9457
rect 4523 9452 4525 9456
rect 4529 9452 4535 9456
rect 4539 9452 4545 9456
rect 4549 9452 4555 9456
rect 4559 9452 4563 9456
rect 4523 9451 4563 9452
rect 4523 9447 4525 9451
rect 4529 9447 4535 9451
rect 4539 9447 4545 9451
rect 4549 9447 4555 9451
rect 4559 9447 4563 9451
rect 4523 9446 4563 9447
rect 4523 9442 4525 9446
rect 4529 9442 4535 9446
rect 4539 9442 4545 9446
rect 4549 9442 4555 9446
rect 4559 9442 4563 9446
rect 4523 9060 4563 9442
rect 4523 9056 4525 9060
rect 4529 9056 4535 9060
rect 4539 9056 4545 9060
rect 4549 9056 4555 9060
rect 4559 9056 4563 9060
rect 4523 9055 4563 9056
rect 4523 9051 4525 9055
rect 4529 9051 4535 9055
rect 4539 9051 4545 9055
rect 4549 9051 4555 9055
rect 4559 9051 4563 9055
rect 4523 9050 4563 9051
rect 4523 9046 4525 9050
rect 4529 9046 4535 9050
rect 4539 9046 4545 9050
rect 4549 9046 4555 9050
rect 4559 9046 4563 9050
rect 4523 9045 4563 9046
rect 4523 9041 4525 9045
rect 4529 9041 4535 9045
rect 4539 9041 4545 9045
rect 4549 9041 4555 9045
rect 4559 9041 4563 9045
rect 4523 8751 4563 9041
rect 4523 8747 4525 8751
rect 4529 8747 4535 8751
rect 4539 8747 4545 8751
rect 4549 8747 4555 8751
rect 4559 8747 4563 8751
rect 4523 8746 4563 8747
rect 4523 8742 4525 8746
rect 4529 8742 4535 8746
rect 4539 8742 4545 8746
rect 4549 8742 4555 8746
rect 4559 8742 4563 8746
rect 4523 8741 4563 8742
rect 4523 8737 4525 8741
rect 4529 8737 4535 8741
rect 4539 8737 4545 8741
rect 4549 8737 4555 8741
rect 4559 8737 4563 8741
rect 4523 8736 4563 8737
rect 4523 8732 4525 8736
rect 4529 8732 4535 8736
rect 4539 8732 4545 8736
rect 4549 8732 4555 8736
rect 4559 8732 4563 8736
rect 4523 8442 4563 8732
rect 4523 8438 4525 8442
rect 4529 8438 4535 8442
rect 4539 8438 4545 8442
rect 4549 8438 4555 8442
rect 4559 8438 4563 8442
rect 4523 8437 4563 8438
rect 4523 8433 4525 8437
rect 4529 8433 4535 8437
rect 4539 8433 4545 8437
rect 4549 8433 4555 8437
rect 4559 8433 4563 8437
rect 4523 8432 4563 8433
rect 4523 8428 4525 8432
rect 4529 8428 4535 8432
rect 4539 8428 4545 8432
rect 4549 8428 4555 8432
rect 4559 8428 4563 8432
rect 4523 8427 4563 8428
rect 4523 8423 4525 8427
rect 4529 8423 4535 8427
rect 4539 8423 4545 8427
rect 4549 8423 4555 8427
rect 4559 8423 4563 8427
rect 4523 8133 4563 8423
rect 4523 8129 4525 8133
rect 4529 8129 4535 8133
rect 4539 8129 4545 8133
rect 4549 8129 4555 8133
rect 4559 8129 4563 8133
rect 4523 8128 4563 8129
rect 4523 8124 4525 8128
rect 4529 8124 4535 8128
rect 4539 8124 4545 8128
rect 4549 8124 4555 8128
rect 4559 8124 4563 8128
rect 4523 8123 4563 8124
rect 4523 8119 4525 8123
rect 4529 8119 4535 8123
rect 4539 8119 4545 8123
rect 4549 8119 4555 8123
rect 4559 8119 4563 8123
rect 4523 8118 4563 8119
rect 4523 8114 4525 8118
rect 4529 8114 4535 8118
rect 4539 8114 4545 8118
rect 4549 8114 4555 8118
rect 4559 8114 4563 8118
rect 4523 8102 4563 8114
rect 4523 8098 4525 8102
rect 4529 8098 4535 8102
rect 4539 8098 4545 8102
rect 4549 8098 4555 8102
rect 4559 8098 4563 8102
rect 4523 8097 4563 8098
rect 4523 8093 4525 8097
rect 4529 8093 4535 8097
rect 4539 8093 4545 8097
rect 4549 8093 4555 8097
rect 4559 8093 4563 8097
rect 4523 8092 4563 8093
rect 4523 8088 4525 8092
rect 4529 8088 4535 8092
rect 4539 8088 4545 8092
rect 4549 8088 4555 8092
rect 4559 8088 4563 8092
rect 4523 8087 4563 8088
rect 4523 8083 4525 8087
rect 4529 8083 4535 8087
rect 4539 8083 4545 8087
rect 4549 8083 4555 8087
rect 4559 8083 4563 8087
rect 4523 7793 4563 8083
rect 4523 7789 4525 7793
rect 4529 7789 4535 7793
rect 4539 7789 4545 7793
rect 4549 7789 4555 7793
rect 4559 7789 4563 7793
rect 4523 7788 4563 7789
rect 4523 7784 4525 7788
rect 4529 7784 4535 7788
rect 4539 7784 4545 7788
rect 4549 7784 4555 7788
rect 4559 7784 4563 7788
rect 4523 7783 4563 7784
rect 4523 7779 4525 7783
rect 4529 7779 4535 7783
rect 4539 7779 4545 7783
rect 4549 7779 4555 7783
rect 4559 7779 4563 7783
rect 4523 7778 4563 7779
rect 4523 7774 4525 7778
rect 4529 7774 4535 7778
rect 4539 7774 4545 7778
rect 4549 7774 4555 7778
rect 4559 7774 4563 7778
rect 4523 7234 4563 7774
rect 4631 7490 4772 7491
rect 4631 7486 4632 7490
rect 4636 7486 4637 7490
rect 4641 7486 4642 7490
rect 4646 7486 4647 7490
rect 4651 7486 4652 7490
rect 4656 7486 4657 7490
rect 4661 7486 4662 7490
rect 4666 7486 4667 7490
rect 4671 7486 4672 7490
rect 4676 7486 4677 7490
rect 4681 7486 4682 7490
rect 4686 7486 4687 7490
rect 4691 7486 4692 7490
rect 4696 7486 4697 7490
rect 4701 7486 4702 7490
rect 4706 7486 4707 7490
rect 4711 7486 4712 7490
rect 4716 7486 4717 7490
rect 4721 7486 4722 7490
rect 4726 7486 4727 7490
rect 4731 7486 4732 7490
rect 4736 7486 4737 7490
rect 4741 7486 4742 7490
rect 4746 7486 4747 7490
rect 4751 7486 4752 7490
rect 4756 7486 4757 7490
rect 4761 7486 4762 7490
rect 4766 7486 4767 7490
rect 4771 7486 4772 7490
rect 4631 7485 4772 7486
rect 4631 7481 4632 7485
rect 4636 7481 4637 7485
rect 4631 7480 4637 7481
rect 4631 7476 4632 7480
rect 4636 7476 4637 7480
rect 4766 7481 4767 7485
rect 4771 7481 4772 7485
rect 4766 7480 4772 7481
rect 4631 7475 4637 7476
rect 4631 7471 4632 7475
rect 4636 7471 4637 7475
rect 4631 7470 4637 7471
rect 4631 7466 4632 7470
rect 4636 7466 4637 7470
rect 4631 7465 4637 7466
rect 4631 7461 4632 7465
rect 4636 7461 4637 7465
rect 4631 7460 4637 7461
rect 4631 7456 4632 7460
rect 4636 7456 4637 7460
rect 4631 7455 4637 7456
rect 4631 7451 4632 7455
rect 4636 7451 4637 7455
rect 4631 7450 4637 7451
rect 4631 7446 4632 7450
rect 4636 7446 4637 7450
rect 4631 7445 4637 7446
rect 4631 7441 4632 7445
rect 4636 7441 4637 7445
rect 4631 7440 4637 7441
rect 4631 7436 4632 7440
rect 4636 7436 4637 7440
rect 4631 7435 4637 7436
rect 4631 7431 4632 7435
rect 4636 7431 4637 7435
rect 4631 7430 4637 7431
rect 4631 7426 4632 7430
rect 4636 7426 4637 7430
rect 4631 7425 4637 7426
rect 4631 7421 4632 7425
rect 4636 7421 4637 7425
rect 4631 7420 4637 7421
rect 4631 7416 4632 7420
rect 4636 7416 4637 7420
rect 4631 7415 4637 7416
rect 4631 7411 4632 7415
rect 4636 7411 4637 7415
rect 4631 7410 4637 7411
rect 4631 7406 4632 7410
rect 4636 7406 4637 7410
rect 4766 7476 4767 7480
rect 4771 7476 4772 7480
rect 4766 7475 4772 7476
rect 4766 7471 4767 7475
rect 4771 7471 4772 7475
rect 4766 7470 4772 7471
rect 4766 7466 4767 7470
rect 4771 7466 4772 7470
rect 4766 7465 4772 7466
rect 4766 7461 4767 7465
rect 4771 7461 4772 7465
rect 4766 7460 4772 7461
rect 4766 7456 4767 7460
rect 4771 7456 4772 7460
rect 4766 7455 4772 7456
rect 4766 7451 4767 7455
rect 4771 7451 4772 7455
rect 4766 7450 4772 7451
rect 4766 7446 4767 7450
rect 4771 7446 4772 7450
rect 4766 7445 4772 7446
rect 4766 7441 4767 7445
rect 4771 7441 4772 7445
rect 4766 7440 4772 7441
rect 4766 7436 4767 7440
rect 4771 7436 4772 7440
rect 4766 7435 4772 7436
rect 4766 7431 4767 7435
rect 4771 7431 4772 7435
rect 4766 7430 4772 7431
rect 4766 7426 4767 7430
rect 4771 7426 4772 7430
rect 4766 7425 4772 7426
rect 4766 7421 4767 7425
rect 4771 7421 4772 7425
rect 4766 7420 4772 7421
rect 4766 7416 4767 7420
rect 4771 7416 4772 7420
rect 4766 7415 4772 7416
rect 4766 7411 4767 7415
rect 4771 7411 4772 7415
rect 4766 7410 4772 7411
rect 4631 7405 4637 7406
rect 4631 7401 4632 7405
rect 4636 7401 4637 7405
rect 4766 7406 4767 7410
rect 4771 7406 4772 7410
rect 4766 7405 4772 7406
rect 4766 7401 4767 7405
rect 4771 7401 4772 7405
rect 4631 7400 4772 7401
rect 4631 7396 4632 7400
rect 4636 7396 4637 7400
rect 4641 7396 4642 7400
rect 4646 7396 4647 7400
rect 4651 7396 4652 7400
rect 4656 7396 4657 7400
rect 4661 7396 4662 7400
rect 4666 7396 4667 7400
rect 4671 7396 4672 7400
rect 4676 7396 4677 7400
rect 4681 7396 4682 7400
rect 4686 7396 4687 7400
rect 4691 7396 4692 7400
rect 4696 7396 4697 7400
rect 4701 7396 4702 7400
rect 4706 7396 4707 7400
rect 4711 7396 4712 7400
rect 4716 7396 4717 7400
rect 4721 7396 4722 7400
rect 4726 7396 4727 7400
rect 4731 7396 4732 7400
rect 4736 7396 4737 7400
rect 4741 7396 4742 7400
rect 4746 7396 4747 7400
rect 4751 7396 4752 7400
rect 4756 7396 4757 7400
rect 4761 7396 4762 7400
rect 4766 7396 4767 7400
rect 4771 7396 4772 7400
rect 4631 7395 4772 7396
rect 4643 7317 4760 7319
rect 4643 7313 4645 7317
rect 4649 7313 4652 7317
rect 4656 7313 4657 7317
rect 4661 7313 4662 7317
rect 4666 7313 4667 7317
rect 4671 7313 4672 7317
rect 4676 7313 4677 7317
rect 4681 7313 4682 7317
rect 4686 7313 4687 7317
rect 4691 7313 4692 7317
rect 4696 7313 4697 7317
rect 4701 7313 4702 7317
rect 4706 7313 4707 7317
rect 4711 7313 4712 7317
rect 4716 7313 4717 7317
rect 4721 7313 4722 7317
rect 4726 7313 4727 7317
rect 4731 7313 4732 7317
rect 4736 7313 4737 7317
rect 4741 7313 4742 7317
rect 4746 7313 4747 7317
rect 4751 7313 4754 7317
rect 4758 7313 4760 7317
rect 4643 7311 4760 7313
rect 4643 7310 4651 7311
rect 4643 7306 4645 7310
rect 4649 7306 4651 7310
rect 4752 7310 4760 7311
rect 4752 7306 4754 7310
rect 4758 7306 4760 7310
rect 4643 7305 4651 7306
rect 4643 7301 4645 7305
rect 4649 7301 4651 7305
rect 4643 7300 4651 7301
rect 4643 7296 4645 7300
rect 4649 7296 4651 7300
rect 4643 7295 4651 7296
rect 4643 7291 4645 7295
rect 4649 7291 4651 7295
rect 4643 7290 4651 7291
rect 4643 7286 4645 7290
rect 4649 7286 4651 7290
rect 4643 7285 4651 7286
rect 4643 7281 4645 7285
rect 4649 7281 4651 7285
rect 4643 7280 4651 7281
rect 4643 7276 4645 7280
rect 4649 7276 4651 7280
rect 4643 7275 4651 7276
rect 4643 7271 4645 7275
rect 4649 7271 4651 7275
rect 4643 7270 4651 7271
rect 4643 7266 4645 7270
rect 4649 7266 4651 7270
rect 4643 7265 4651 7266
rect 4643 7261 4645 7265
rect 4649 7261 4651 7265
rect 4752 7305 4760 7306
rect 4752 7301 4754 7305
rect 4758 7301 4760 7305
rect 4752 7300 4760 7301
rect 4752 7296 4754 7300
rect 4758 7296 4760 7300
rect 4752 7295 4760 7296
rect 4752 7291 4754 7295
rect 4758 7291 4760 7295
rect 4752 7290 4760 7291
rect 4752 7286 4754 7290
rect 4758 7286 4760 7290
rect 4752 7285 4760 7286
rect 4752 7281 4754 7285
rect 4758 7281 4760 7285
rect 4752 7280 4760 7281
rect 4752 7276 4754 7280
rect 4758 7276 4760 7280
rect 4752 7275 4760 7276
rect 4752 7271 4754 7275
rect 4758 7271 4760 7275
rect 4752 7270 4760 7271
rect 4752 7266 4754 7270
rect 4758 7266 4760 7270
rect 4752 7265 4760 7266
rect 4752 7261 4754 7265
rect 4758 7261 4760 7265
rect 4643 7260 4651 7261
rect 4643 7256 4645 7260
rect 4649 7256 4651 7260
rect 4643 7255 4651 7256
rect 4752 7260 4760 7261
rect 4752 7256 4754 7260
rect 4758 7256 4760 7260
rect 4752 7255 4760 7256
rect 4643 7253 4760 7255
rect 4643 7249 4645 7253
rect 4649 7249 4652 7253
rect 4656 7249 4657 7253
rect 4661 7249 4662 7253
rect 4666 7249 4667 7253
rect 4671 7249 4672 7253
rect 4676 7249 4677 7253
rect 4681 7249 4682 7253
rect 4686 7249 4687 7253
rect 4691 7249 4692 7253
rect 4696 7249 4697 7253
rect 4701 7249 4702 7253
rect 4706 7249 4707 7253
rect 4711 7249 4712 7253
rect 4716 7249 4717 7253
rect 4721 7249 4722 7253
rect 4726 7249 4727 7253
rect 4731 7249 4732 7253
rect 4736 7249 4737 7253
rect 4741 7249 4742 7253
rect 4746 7249 4747 7253
rect 4751 7249 4754 7253
rect 4758 7249 4760 7253
rect 4643 7247 4760 7249
rect 4523 7230 4525 7234
rect 4529 7230 4535 7234
rect 4539 7230 4545 7234
rect 4549 7230 4555 7234
rect 4559 7230 4563 7234
rect 4523 7229 4563 7230
rect 4523 7225 4525 7229
rect 4529 7225 4535 7229
rect 4539 7225 4545 7229
rect 4549 7225 4555 7229
rect 4559 7225 4563 7229
rect 4523 7224 4563 7225
rect 4523 7220 4525 7224
rect 4529 7220 4535 7224
rect 4539 7220 4545 7224
rect 4549 7220 4555 7224
rect 4559 7220 4563 7224
rect 4523 7219 4563 7220
rect 4523 7215 4525 7219
rect 4529 7215 4535 7219
rect 4539 7215 4545 7219
rect 4549 7215 4555 7219
rect 4559 7215 4563 7219
rect 4523 7206 4563 7215
rect 4523 7202 4525 7206
rect 4529 7202 4535 7206
rect 4539 7202 4545 7206
rect 4549 7202 4555 7206
rect 4559 7202 4563 7206
rect 4523 7201 4563 7202
rect 4523 7197 4525 7201
rect 4529 7197 4535 7201
rect 4539 7197 4545 7201
rect 4549 7197 4555 7201
rect 4559 7197 4563 7201
rect 4523 7196 4563 7197
rect 4523 7192 4525 7196
rect 4529 7192 4535 7196
rect 4539 7192 4545 7196
rect 4549 7192 4555 7196
rect 4559 7192 4563 7196
rect 4523 7191 4563 7192
rect 4523 7187 4525 7191
rect 4529 7187 4535 7191
rect 4539 7187 4545 7191
rect 4549 7187 4555 7191
rect 4559 7187 4563 7191
rect 4523 7156 4563 7187
rect 4523 7152 4525 7156
rect 4529 7152 4535 7156
rect 4539 7152 4545 7156
rect 4549 7152 4555 7156
rect 4559 7152 4563 7156
rect 4523 6862 4563 7152
rect 4523 6858 4525 6862
rect 4529 6858 4535 6862
rect 4539 6858 4545 6862
rect 4549 6858 4555 6862
rect 4559 6858 4563 6862
rect 4523 6857 4563 6858
rect 4523 6853 4525 6857
rect 4529 6853 4535 6857
rect 4539 6853 4545 6857
rect 4549 6853 4555 6857
rect 4559 6853 4563 6857
rect 4523 6852 4563 6853
rect 4523 6848 4525 6852
rect 4529 6848 4535 6852
rect 4539 6848 4545 6852
rect 4549 6848 4555 6852
rect 4559 6848 4563 6852
rect 4523 6847 4563 6848
rect 4523 6843 4525 6847
rect 4529 6843 4535 6847
rect 4539 6843 4545 6847
rect 4549 6843 4555 6847
rect 4559 6843 4563 6847
rect 4523 6553 4563 6843
rect 4523 6549 4525 6553
rect 4529 6549 4535 6553
rect 4539 6549 4545 6553
rect 4549 6549 4555 6553
rect 4559 6549 4563 6553
rect 4523 6548 4563 6549
rect 4523 6544 4525 6548
rect 4529 6544 4535 6548
rect 4539 6544 4545 6548
rect 4549 6544 4555 6548
rect 4559 6544 4563 6548
rect 4523 6543 4563 6544
rect 4523 6539 4525 6543
rect 4529 6539 4535 6543
rect 4539 6539 4545 6543
rect 4549 6539 4555 6543
rect 4559 6539 4563 6543
rect 4523 6538 4563 6539
rect 4523 6534 4525 6538
rect 4529 6534 4535 6538
rect 4539 6534 4545 6538
rect 4549 6534 4555 6538
rect 4559 6534 4563 6538
rect 4523 6244 4563 6534
rect 4523 6240 4525 6244
rect 4529 6240 4535 6244
rect 4539 6240 4545 6244
rect 4549 6240 4555 6244
rect 4559 6240 4563 6244
rect 4523 6239 4563 6240
rect 4523 6235 4525 6239
rect 4529 6235 4535 6239
rect 4539 6235 4545 6239
rect 4549 6235 4555 6239
rect 4559 6235 4563 6239
rect 4523 6234 4563 6235
rect 4523 6230 4525 6234
rect 4529 6230 4535 6234
rect 4539 6230 4545 6234
rect 4549 6230 4555 6234
rect 4559 6230 4563 6234
rect 4523 6229 4563 6230
rect 4523 6225 4525 6229
rect 4529 6225 4535 6229
rect 4539 6225 4545 6229
rect 4549 6225 4555 6229
rect 4559 6225 4563 6229
rect 4523 5935 4563 6225
rect 4523 5931 4525 5935
rect 4529 5931 4535 5935
rect 4539 5931 4545 5935
rect 4549 5931 4555 5935
rect 4559 5931 4563 5935
rect 4523 5930 4563 5931
rect 4523 5926 4525 5930
rect 4529 5926 4535 5930
rect 4539 5926 4545 5930
rect 4549 5926 4555 5930
rect 4559 5926 4563 5930
rect 4523 5925 4563 5926
rect 4523 5921 4525 5925
rect 4529 5921 4535 5925
rect 4539 5921 4545 5925
rect 4549 5921 4555 5925
rect 4559 5921 4563 5925
rect 4523 5920 4563 5921
rect 4523 5916 4525 5920
rect 4529 5916 4535 5920
rect 4539 5916 4545 5920
rect 4549 5916 4555 5920
rect 4559 5916 4563 5920
rect 4523 5626 4563 5916
rect 4523 5622 4525 5626
rect 4529 5622 4535 5626
rect 4539 5622 4545 5626
rect 4549 5622 4555 5626
rect 4559 5622 4563 5626
rect 4523 5621 4563 5622
rect 4523 5617 4525 5621
rect 4529 5617 4535 5621
rect 4539 5617 4545 5621
rect 4549 5617 4555 5621
rect 4559 5617 4563 5621
rect 4523 5616 4563 5617
rect 4523 5612 4525 5616
rect 4529 5612 4535 5616
rect 4539 5612 4545 5616
rect 4549 5612 4555 5616
rect 4559 5612 4563 5616
rect 4523 5611 4563 5612
rect 4523 5607 4525 5611
rect 4529 5607 4535 5611
rect 4539 5607 4545 5611
rect 4549 5607 4555 5611
rect 4559 5607 4563 5611
rect 4523 5317 4563 5607
rect 4523 5313 4525 5317
rect 4529 5313 4535 5317
rect 4539 5313 4545 5317
rect 4549 5313 4555 5317
rect 4559 5313 4563 5317
rect 4523 5312 4563 5313
rect 4523 5308 4525 5312
rect 4529 5308 4535 5312
rect 4539 5308 4545 5312
rect 4549 5308 4555 5312
rect 4559 5308 4563 5312
rect 4523 5307 4563 5308
rect 4523 5303 4525 5307
rect 4529 5303 4535 5307
rect 4539 5303 4545 5307
rect 4549 5303 4555 5307
rect 4559 5303 4563 5307
rect 4523 5302 4563 5303
rect 4523 5298 4525 5302
rect 4529 5298 4535 5302
rect 4539 5298 4545 5302
rect 4549 5298 4555 5302
rect 4559 5298 4563 5302
rect 4523 5008 4563 5298
rect 4523 5004 4525 5008
rect 4529 5004 4535 5008
rect 4539 5004 4545 5008
rect 4549 5004 4555 5008
rect 4559 5004 4563 5008
rect 4523 5003 4563 5004
rect 4523 4999 4525 5003
rect 4529 4999 4535 5003
rect 4539 4999 4545 5003
rect 4549 4999 4555 5003
rect 4559 4999 4563 5003
rect 4523 4998 4563 4999
rect 4523 4994 4525 4998
rect 4529 4994 4535 4998
rect 4539 4994 4545 4998
rect 4549 4994 4555 4998
rect 4559 4994 4563 4998
rect 4523 4993 4563 4994
rect 4523 4989 4525 4993
rect 4529 4989 4535 4993
rect 4539 4989 4545 4993
rect 4549 4989 4555 4993
rect 4559 4989 4563 4993
rect 4523 4815 4563 4989
rect 4523 4811 4525 4815
rect 4529 4811 4535 4815
rect 4539 4811 4545 4815
rect 4549 4811 4555 4815
rect 4559 4811 4563 4815
rect 4523 4810 4563 4811
rect 4523 4806 4525 4810
rect 4529 4806 4535 4810
rect 4539 4806 4545 4810
rect 4549 4806 4555 4810
rect 4559 4806 4563 4810
rect 4523 4805 4563 4806
rect 4523 4801 4525 4805
rect 4529 4801 4535 4805
rect 4539 4801 4545 4805
rect 4549 4801 4555 4805
rect 4559 4801 4563 4805
rect 4523 4800 4563 4801
rect 4523 4796 4525 4800
rect 4529 4796 4535 4800
rect 4539 4796 4545 4800
rect 4549 4796 4555 4800
rect 4559 4796 4563 4800
rect 4523 4789 4563 4796
rect 4523 4785 4525 4789
rect 4529 4785 4535 4789
rect 4539 4785 4545 4789
rect 4549 4785 4555 4789
rect 4559 4785 4563 4789
rect 4523 4784 4563 4785
rect 4523 4780 4525 4784
rect 4529 4780 4535 4784
rect 4539 4780 4545 4784
rect 4549 4780 4555 4784
rect 4559 4780 4563 4784
rect 4523 4779 4563 4780
rect 4523 4775 4525 4779
rect 4529 4775 4535 4779
rect 4539 4775 4545 4779
rect 4549 4775 4555 4779
rect 4559 4775 4563 4779
rect 4523 4774 4563 4775
rect 4523 4770 4525 4774
rect 4529 4770 4535 4774
rect 4539 4770 4545 4774
rect 4549 4770 4555 4774
rect 4559 4770 4563 4774
rect 4523 4763 4563 4770
rect 4523 4759 4525 4763
rect 4529 4759 4535 4763
rect 4539 4759 4545 4763
rect 4549 4759 4555 4763
rect 4559 4759 4563 4763
rect 4523 4758 4563 4759
rect 4523 4754 4525 4758
rect 4529 4754 4535 4758
rect 4539 4754 4545 4758
rect 4549 4754 4555 4758
rect 4559 4754 4563 4758
rect 4523 4753 4563 4754
rect 4523 4749 4525 4753
rect 4529 4749 4535 4753
rect 4539 4749 4545 4753
rect 4549 4749 4555 4753
rect 4559 4749 4563 4753
rect 4523 4748 4563 4749
rect 4523 4744 4525 4748
rect 4529 4744 4535 4748
rect 4539 4744 4545 4748
rect 4549 4744 4555 4748
rect 4559 4744 4563 4748
rect 4523 4737 4563 4744
rect 4523 4733 4525 4737
rect 4529 4733 4535 4737
rect 4539 4733 4545 4737
rect 4549 4733 4555 4737
rect 4559 4733 4563 4737
rect 4523 4732 4563 4733
rect 4523 4728 4525 4732
rect 4529 4728 4535 4732
rect 4539 4728 4545 4732
rect 4549 4728 4555 4732
rect 4559 4728 4563 4732
rect 4523 4727 4563 4728
rect 4523 4723 4525 4727
rect 4529 4723 4535 4727
rect 4539 4723 4545 4727
rect 4549 4723 4555 4727
rect 4559 4723 4563 4727
rect 4523 4722 4563 4723
rect 4523 4718 4525 4722
rect 4529 4718 4535 4722
rect 4539 4718 4545 4722
rect 4549 4718 4555 4722
rect 4559 4718 4563 4722
rect 4523 4711 4563 4718
rect 4523 4707 4525 4711
rect 4529 4707 4535 4711
rect 4539 4707 4545 4711
rect 4549 4707 4555 4711
rect 4559 4707 4563 4711
rect 4523 4706 4563 4707
rect 4523 4702 4525 4706
rect 4529 4702 4535 4706
rect 4539 4702 4545 4706
rect 4549 4702 4555 4706
rect 4559 4702 4563 4706
rect 4523 4701 4563 4702
rect 4523 4697 4525 4701
rect 4529 4697 4535 4701
rect 4539 4697 4545 4701
rect 4549 4697 4555 4701
rect 4559 4697 4563 4701
rect 4523 4696 4563 4697
rect 4523 4692 4525 4696
rect 4529 4692 4535 4696
rect 4539 4692 4545 4696
rect 4549 4692 4555 4696
rect 4559 4692 4563 4696
rect 4523 4584 4563 4692
rect 609 4582 4563 4584
rect 609 4578 757 4582
rect 761 4578 762 4582
rect 766 4578 767 4582
rect 771 4578 772 4582
rect 776 4578 783 4582
rect 787 4578 788 4582
rect 792 4578 793 4582
rect 797 4578 798 4582
rect 802 4578 809 4582
rect 813 4578 814 4582
rect 818 4578 819 4582
rect 823 4578 824 4582
rect 828 4578 835 4582
rect 839 4578 840 4582
rect 844 4578 845 4582
rect 849 4578 850 4582
rect 854 4578 861 4582
rect 865 4578 866 4582
rect 870 4578 871 4582
rect 875 4578 876 4582
rect 880 4578 1053 4582
rect 1057 4578 1058 4582
rect 1062 4578 1063 4582
rect 1067 4578 1068 4582
rect 1072 4578 1362 4582
rect 1366 4578 1367 4582
rect 1371 4578 1372 4582
rect 1376 4578 1377 4582
rect 1381 4578 1671 4582
rect 1675 4578 1676 4582
rect 1680 4578 1681 4582
rect 1685 4578 1686 4582
rect 1690 4578 1980 4582
rect 1984 4578 1985 4582
rect 1989 4578 1990 4582
rect 1994 4578 1995 4582
rect 1999 4578 2289 4582
rect 2293 4578 2294 4582
rect 2298 4578 2299 4582
rect 2303 4578 2304 4582
rect 2308 4578 2598 4582
rect 2602 4578 2603 4582
rect 2607 4578 2608 4582
rect 2612 4578 2613 4582
rect 2617 4578 2907 4582
rect 2911 4578 2912 4582
rect 2916 4578 2917 4582
rect 2921 4578 2922 4582
rect 2926 4578 3216 4582
rect 3220 4578 3221 4582
rect 3225 4578 3226 4582
rect 3230 4578 3231 4582
rect 3235 4578 3525 4582
rect 3529 4578 3530 4582
rect 3534 4578 3535 4582
rect 3539 4578 3540 4582
rect 3544 4578 3834 4582
rect 3838 4578 3839 4582
rect 3843 4578 3844 4582
rect 3848 4578 3849 4582
rect 3853 4578 4235 4582
rect 4239 4578 4240 4582
rect 4244 4578 4245 4582
rect 4249 4578 4250 4582
rect 4254 4578 4264 4582
rect 4268 4578 4269 4582
rect 4273 4578 4274 4582
rect 4278 4578 4279 4582
rect 4283 4578 4293 4582
rect 4297 4578 4298 4582
rect 4302 4578 4303 4582
rect 4307 4578 4308 4582
rect 4312 4578 4322 4582
rect 4326 4578 4327 4582
rect 4331 4578 4332 4582
rect 4336 4578 4337 4582
rect 4341 4578 4351 4582
rect 4355 4578 4356 4582
rect 4360 4578 4361 4582
rect 4365 4578 4366 4582
rect 4370 4578 4563 4582
rect 609 4572 4563 4578
rect 609 4568 757 4572
rect 761 4568 762 4572
rect 766 4568 767 4572
rect 771 4568 772 4572
rect 776 4568 783 4572
rect 787 4568 788 4572
rect 792 4568 793 4572
rect 797 4568 798 4572
rect 802 4568 809 4572
rect 813 4568 814 4572
rect 818 4568 819 4572
rect 823 4568 824 4572
rect 828 4568 835 4572
rect 839 4568 840 4572
rect 844 4568 845 4572
rect 849 4568 850 4572
rect 854 4568 861 4572
rect 865 4568 866 4572
rect 870 4568 871 4572
rect 875 4568 876 4572
rect 880 4568 1053 4572
rect 1057 4568 1058 4572
rect 1062 4568 1063 4572
rect 1067 4568 1068 4572
rect 1072 4568 1362 4572
rect 1366 4568 1367 4572
rect 1371 4568 1372 4572
rect 1376 4568 1377 4572
rect 1381 4568 1671 4572
rect 1675 4568 1676 4572
rect 1680 4568 1681 4572
rect 1685 4568 1686 4572
rect 1690 4568 1980 4572
rect 1984 4568 1985 4572
rect 1989 4568 1990 4572
rect 1994 4568 1995 4572
rect 1999 4568 2289 4572
rect 2293 4568 2294 4572
rect 2298 4568 2299 4572
rect 2303 4568 2304 4572
rect 2308 4568 2598 4572
rect 2602 4568 2603 4572
rect 2607 4568 2608 4572
rect 2612 4568 2613 4572
rect 2617 4568 2907 4572
rect 2911 4568 2912 4572
rect 2916 4568 2917 4572
rect 2921 4568 2922 4572
rect 2926 4568 3216 4572
rect 3220 4568 3221 4572
rect 3225 4568 3226 4572
rect 3230 4568 3231 4572
rect 3235 4568 3525 4572
rect 3529 4568 3530 4572
rect 3534 4568 3535 4572
rect 3539 4568 3540 4572
rect 3544 4568 3834 4572
rect 3838 4568 3839 4572
rect 3843 4568 3844 4572
rect 3848 4568 3849 4572
rect 3853 4568 4235 4572
rect 4239 4568 4240 4572
rect 4244 4568 4245 4572
rect 4249 4568 4250 4572
rect 4254 4568 4264 4572
rect 4268 4568 4269 4572
rect 4273 4568 4274 4572
rect 4278 4568 4279 4572
rect 4283 4568 4293 4572
rect 4297 4568 4298 4572
rect 4302 4568 4303 4572
rect 4307 4568 4308 4572
rect 4312 4568 4322 4572
rect 4326 4568 4327 4572
rect 4331 4568 4332 4572
rect 4336 4568 4337 4572
rect 4341 4568 4351 4572
rect 4355 4568 4356 4572
rect 4360 4568 4361 4572
rect 4365 4568 4366 4572
rect 4370 4568 4563 4572
rect 609 4562 4563 4568
rect 609 4558 757 4562
rect 761 4558 762 4562
rect 766 4558 767 4562
rect 771 4558 772 4562
rect 776 4558 783 4562
rect 787 4558 788 4562
rect 792 4558 793 4562
rect 797 4558 798 4562
rect 802 4558 809 4562
rect 813 4558 814 4562
rect 818 4558 819 4562
rect 823 4558 824 4562
rect 828 4558 835 4562
rect 839 4558 840 4562
rect 844 4558 845 4562
rect 849 4558 850 4562
rect 854 4558 861 4562
rect 865 4558 866 4562
rect 870 4558 871 4562
rect 875 4558 876 4562
rect 880 4558 1053 4562
rect 1057 4558 1058 4562
rect 1062 4558 1063 4562
rect 1067 4558 1068 4562
rect 1072 4558 1362 4562
rect 1366 4558 1367 4562
rect 1371 4558 1372 4562
rect 1376 4558 1377 4562
rect 1381 4558 1671 4562
rect 1675 4558 1676 4562
rect 1680 4558 1681 4562
rect 1685 4558 1686 4562
rect 1690 4558 1980 4562
rect 1984 4558 1985 4562
rect 1989 4558 1990 4562
rect 1994 4558 1995 4562
rect 1999 4558 2289 4562
rect 2293 4558 2294 4562
rect 2298 4558 2299 4562
rect 2303 4558 2304 4562
rect 2308 4558 2598 4562
rect 2602 4558 2603 4562
rect 2607 4558 2608 4562
rect 2612 4558 2613 4562
rect 2617 4558 2907 4562
rect 2911 4558 2912 4562
rect 2916 4558 2917 4562
rect 2921 4558 2922 4562
rect 2926 4558 3216 4562
rect 3220 4558 3221 4562
rect 3225 4558 3226 4562
rect 3230 4558 3231 4562
rect 3235 4558 3525 4562
rect 3529 4558 3530 4562
rect 3534 4558 3535 4562
rect 3539 4558 3540 4562
rect 3544 4558 3834 4562
rect 3838 4558 3839 4562
rect 3843 4558 3844 4562
rect 3848 4558 3849 4562
rect 3853 4558 4235 4562
rect 4239 4558 4240 4562
rect 4244 4558 4245 4562
rect 4249 4558 4250 4562
rect 4254 4558 4264 4562
rect 4268 4558 4269 4562
rect 4273 4558 4274 4562
rect 4278 4558 4279 4562
rect 4283 4558 4293 4562
rect 4297 4558 4298 4562
rect 4302 4558 4303 4562
rect 4307 4558 4308 4562
rect 4312 4558 4322 4562
rect 4326 4558 4327 4562
rect 4331 4558 4332 4562
rect 4336 4558 4337 4562
rect 4341 4558 4351 4562
rect 4355 4558 4356 4562
rect 4360 4558 4361 4562
rect 4365 4558 4366 4562
rect 4370 4558 4563 4562
rect 609 4552 4563 4558
rect 609 4548 757 4552
rect 761 4548 762 4552
rect 766 4548 767 4552
rect 771 4548 772 4552
rect 776 4548 783 4552
rect 787 4548 788 4552
rect 792 4548 793 4552
rect 797 4548 798 4552
rect 802 4548 809 4552
rect 813 4548 814 4552
rect 818 4548 819 4552
rect 823 4548 824 4552
rect 828 4548 835 4552
rect 839 4548 840 4552
rect 844 4548 845 4552
rect 849 4548 850 4552
rect 854 4548 861 4552
rect 865 4548 866 4552
rect 870 4548 871 4552
rect 875 4548 876 4552
rect 880 4548 1053 4552
rect 1057 4548 1058 4552
rect 1062 4548 1063 4552
rect 1067 4548 1068 4552
rect 1072 4548 1362 4552
rect 1366 4548 1367 4552
rect 1371 4548 1372 4552
rect 1376 4548 1377 4552
rect 1381 4548 1671 4552
rect 1675 4548 1676 4552
rect 1680 4548 1681 4552
rect 1685 4548 1686 4552
rect 1690 4548 1980 4552
rect 1984 4548 1985 4552
rect 1989 4548 1990 4552
rect 1994 4548 1995 4552
rect 1999 4548 2289 4552
rect 2293 4548 2294 4552
rect 2298 4548 2299 4552
rect 2303 4548 2304 4552
rect 2308 4548 2598 4552
rect 2602 4548 2603 4552
rect 2607 4548 2608 4552
rect 2612 4548 2613 4552
rect 2617 4548 2907 4552
rect 2911 4548 2912 4552
rect 2916 4548 2917 4552
rect 2921 4548 2922 4552
rect 2926 4548 3216 4552
rect 3220 4548 3221 4552
rect 3225 4548 3226 4552
rect 3230 4548 3231 4552
rect 3235 4548 3525 4552
rect 3529 4548 3530 4552
rect 3534 4548 3535 4552
rect 3539 4548 3540 4552
rect 3544 4548 3834 4552
rect 3838 4548 3839 4552
rect 3843 4548 3844 4552
rect 3848 4548 3849 4552
rect 3853 4548 4235 4552
rect 4239 4548 4240 4552
rect 4244 4548 4245 4552
rect 4249 4548 4250 4552
rect 4254 4548 4264 4552
rect 4268 4548 4269 4552
rect 4273 4548 4274 4552
rect 4278 4548 4279 4552
rect 4283 4548 4293 4552
rect 4297 4548 4298 4552
rect 4302 4548 4303 4552
rect 4307 4548 4308 4552
rect 4312 4548 4322 4552
rect 4326 4548 4327 4552
rect 4331 4548 4332 4552
rect 4336 4548 4337 4552
rect 4341 4548 4351 4552
rect 4355 4548 4356 4552
rect 4360 4548 4361 4552
rect 4365 4548 4366 4552
rect 4370 4548 4563 4552
rect 609 4544 4563 4548
rect 1085 4462 1157 4464
rect 1085 4458 1087 4462
rect 1091 4458 1094 4462
rect 1098 4458 1099 4462
rect 1103 4458 1104 4462
rect 1108 4458 1109 4462
rect 1113 4458 1114 4462
rect 1118 4458 1119 4462
rect 1123 4458 1124 4462
rect 1128 4458 1129 4462
rect 1133 4458 1134 4462
rect 1138 4458 1139 4462
rect 1143 4458 1144 4462
rect 1148 4458 1151 4462
rect 1155 4458 1157 4462
rect 1085 4456 1157 4458
rect 1085 4455 1093 4456
rect 1085 4451 1087 4455
rect 1091 4451 1093 4455
rect 1085 4450 1093 4451
rect 1149 4455 1157 4456
rect 1149 4451 1151 4455
rect 1155 4451 1157 4455
rect 1149 4450 1157 4451
rect 1085 4446 1087 4450
rect 1091 4446 1093 4450
rect 1085 4445 1093 4446
rect 1085 4441 1087 4445
rect 1091 4441 1093 4445
rect 1085 4440 1093 4441
rect 1085 4436 1087 4440
rect 1091 4436 1093 4440
rect 1085 4435 1093 4436
rect 1085 4431 1087 4435
rect 1091 4431 1093 4435
rect 1085 4430 1093 4431
rect 1085 4426 1087 4430
rect 1091 4426 1093 4430
rect 1085 4425 1093 4426
rect 1085 4421 1087 4425
rect 1091 4421 1093 4425
rect 1085 4420 1093 4421
rect 1085 4416 1087 4420
rect 1091 4416 1093 4420
rect 1085 4415 1093 4416
rect 1085 4411 1087 4415
rect 1091 4411 1093 4415
rect 1085 4410 1093 4411
rect 1085 4406 1087 4410
rect 1091 4406 1093 4410
rect 1085 4405 1093 4406
rect 1085 4401 1087 4405
rect 1091 4401 1093 4405
rect 1085 4400 1093 4401
rect 1085 4396 1087 4400
rect 1091 4396 1093 4400
rect 1085 4395 1093 4396
rect 1085 4391 1087 4395
rect 1091 4391 1093 4395
rect 1085 4390 1093 4391
rect 1085 4386 1087 4390
rect 1091 4386 1093 4390
rect 1085 4385 1093 4386
rect 1085 4381 1087 4385
rect 1091 4381 1093 4385
rect 1085 4380 1093 4381
rect 1085 4376 1087 4380
rect 1091 4376 1093 4380
rect 1085 4375 1093 4376
rect 1085 4371 1087 4375
rect 1091 4371 1093 4375
rect 1085 4370 1093 4371
rect 1085 4366 1087 4370
rect 1091 4366 1093 4370
rect 1085 4365 1093 4366
rect 1085 4361 1087 4365
rect 1091 4361 1093 4365
rect 1149 4446 1151 4450
rect 1155 4446 1157 4450
rect 1149 4445 1157 4446
rect 1149 4441 1151 4445
rect 1155 4441 1157 4445
rect 1149 4440 1157 4441
rect 1149 4436 1151 4440
rect 1155 4436 1157 4440
rect 1149 4435 1157 4436
rect 1149 4431 1151 4435
rect 1155 4431 1157 4435
rect 1149 4430 1157 4431
rect 1149 4426 1151 4430
rect 1155 4426 1157 4430
rect 1149 4425 1157 4426
rect 1149 4421 1151 4425
rect 1155 4421 1157 4425
rect 1149 4420 1157 4421
rect 1149 4416 1151 4420
rect 1155 4416 1157 4420
rect 1149 4415 1157 4416
rect 1149 4411 1151 4415
rect 1155 4411 1157 4415
rect 1149 4410 1157 4411
rect 1149 4406 1151 4410
rect 1155 4406 1157 4410
rect 1149 4405 1157 4406
rect 1149 4401 1151 4405
rect 1155 4401 1157 4405
rect 1149 4400 1157 4401
rect 1149 4396 1151 4400
rect 1155 4396 1157 4400
rect 1149 4395 1157 4396
rect 1149 4391 1151 4395
rect 1155 4391 1157 4395
rect 1149 4390 1157 4391
rect 1149 4386 1151 4390
rect 1155 4386 1157 4390
rect 1149 4385 1157 4386
rect 1149 4381 1151 4385
rect 1155 4381 1157 4385
rect 1149 4380 1157 4381
rect 1149 4376 1151 4380
rect 1155 4376 1157 4380
rect 1149 4375 1157 4376
rect 1149 4371 1151 4375
rect 1155 4371 1157 4375
rect 1149 4370 1157 4371
rect 1149 4366 1151 4370
rect 1155 4366 1157 4370
rect 1149 4365 1157 4366
rect 1149 4361 1151 4365
rect 1155 4361 1157 4365
rect 1085 4360 1093 4361
rect 1085 4356 1087 4360
rect 1091 4356 1093 4360
rect 1085 4355 1093 4356
rect 1149 4360 1157 4361
rect 1149 4356 1151 4360
rect 1155 4356 1157 4360
rect 1149 4355 1157 4356
rect 1085 4353 1157 4355
rect 1085 4349 1087 4353
rect 1091 4349 1094 4353
rect 1098 4349 1099 4353
rect 1103 4349 1104 4353
rect 1108 4349 1109 4353
rect 1113 4349 1114 4353
rect 1118 4349 1119 4353
rect 1123 4349 1124 4353
rect 1128 4349 1129 4353
rect 1133 4349 1134 4353
rect 1138 4349 1139 4353
rect 1143 4349 1144 4353
rect 1148 4349 1151 4353
rect 1155 4349 1157 4353
rect 1085 4347 1157 4349
rect 1233 4475 1329 4476
rect 1233 4471 1234 4475
rect 1238 4471 1239 4475
rect 1243 4471 1244 4475
rect 1248 4471 1249 4475
rect 1253 4471 1254 4475
rect 1258 4471 1259 4475
rect 1263 4471 1264 4475
rect 1268 4471 1269 4475
rect 1273 4471 1274 4475
rect 1278 4471 1279 4475
rect 1283 4471 1284 4475
rect 1288 4471 1289 4475
rect 1293 4471 1294 4475
rect 1298 4471 1299 4475
rect 1303 4471 1304 4475
rect 1308 4471 1309 4475
rect 1313 4471 1314 4475
rect 1318 4471 1319 4475
rect 1323 4471 1324 4475
rect 1328 4471 1329 4475
rect 1233 4470 1329 4471
rect 1233 4466 1234 4470
rect 1238 4466 1239 4470
rect 1233 4465 1239 4466
rect 1233 4461 1234 4465
rect 1238 4461 1239 4465
rect 1323 4466 1324 4470
rect 1328 4466 1329 4470
rect 1323 4465 1329 4466
rect 1233 4460 1239 4461
rect 1233 4456 1234 4460
rect 1238 4456 1239 4460
rect 1233 4455 1239 4456
rect 1233 4451 1234 4455
rect 1238 4451 1239 4455
rect 1233 4450 1239 4451
rect 1233 4446 1234 4450
rect 1238 4446 1239 4450
rect 1233 4445 1239 4446
rect 1233 4441 1234 4445
rect 1238 4441 1239 4445
rect 1233 4440 1239 4441
rect 1233 4436 1234 4440
rect 1238 4436 1239 4440
rect 1233 4435 1239 4436
rect 1233 4431 1234 4435
rect 1238 4431 1239 4435
rect 1233 4430 1239 4431
rect 1233 4426 1234 4430
rect 1238 4426 1239 4430
rect 1233 4425 1239 4426
rect 1233 4421 1234 4425
rect 1238 4421 1239 4425
rect 1233 4420 1239 4421
rect 1233 4416 1234 4420
rect 1238 4416 1239 4420
rect 1233 4415 1239 4416
rect 1233 4411 1234 4415
rect 1238 4411 1239 4415
rect 1233 4410 1239 4411
rect 1233 4406 1234 4410
rect 1238 4406 1239 4410
rect 1233 4405 1239 4406
rect 1233 4401 1234 4405
rect 1238 4401 1239 4405
rect 1233 4400 1239 4401
rect 1233 4396 1234 4400
rect 1238 4396 1239 4400
rect 1233 4395 1239 4396
rect 1233 4391 1234 4395
rect 1238 4391 1239 4395
rect 1233 4390 1239 4391
rect 1233 4386 1234 4390
rect 1238 4386 1239 4390
rect 1233 4385 1239 4386
rect 1233 4381 1234 4385
rect 1238 4381 1239 4385
rect 1233 4380 1239 4381
rect 1233 4376 1234 4380
rect 1238 4376 1239 4380
rect 1233 4375 1239 4376
rect 1233 4371 1234 4375
rect 1238 4371 1239 4375
rect 1233 4370 1239 4371
rect 1233 4366 1234 4370
rect 1238 4366 1239 4370
rect 1233 4365 1239 4366
rect 1233 4361 1234 4365
rect 1238 4361 1239 4365
rect 1233 4360 1239 4361
rect 1233 4356 1234 4360
rect 1238 4356 1239 4360
rect 1233 4355 1239 4356
rect 1233 4351 1234 4355
rect 1238 4351 1239 4355
rect 1233 4350 1239 4351
rect 1233 4346 1234 4350
rect 1238 4346 1239 4350
rect 1323 4461 1324 4465
rect 1328 4461 1329 4465
rect 1323 4460 1329 4461
rect 1323 4456 1324 4460
rect 1328 4456 1329 4460
rect 1323 4455 1329 4456
rect 1323 4451 1324 4455
rect 1328 4451 1329 4455
rect 1323 4450 1329 4451
rect 1323 4446 1324 4450
rect 1328 4446 1329 4450
rect 1323 4445 1329 4446
rect 1323 4441 1324 4445
rect 1328 4441 1329 4445
rect 1323 4440 1329 4441
rect 1323 4436 1324 4440
rect 1328 4436 1329 4440
rect 1323 4435 1329 4436
rect 1323 4431 1324 4435
rect 1328 4431 1329 4435
rect 1323 4430 1329 4431
rect 1323 4426 1324 4430
rect 1328 4426 1329 4430
rect 1323 4425 1329 4426
rect 1323 4421 1324 4425
rect 1328 4421 1329 4425
rect 1323 4420 1329 4421
rect 1323 4416 1324 4420
rect 1328 4416 1329 4420
rect 1323 4415 1329 4416
rect 1323 4411 1324 4415
rect 1328 4411 1329 4415
rect 1323 4410 1329 4411
rect 1323 4406 1324 4410
rect 1328 4406 1329 4410
rect 1323 4405 1329 4406
rect 1323 4401 1324 4405
rect 1328 4401 1329 4405
rect 1323 4400 1329 4401
rect 1323 4396 1324 4400
rect 1328 4396 1329 4400
rect 1323 4395 1329 4396
rect 1323 4391 1324 4395
rect 1328 4391 1329 4395
rect 1323 4390 1329 4391
rect 1323 4386 1324 4390
rect 1328 4386 1329 4390
rect 1323 4385 1329 4386
rect 1323 4381 1324 4385
rect 1328 4381 1329 4385
rect 1323 4380 1329 4381
rect 1323 4376 1324 4380
rect 1328 4376 1329 4380
rect 1323 4375 1329 4376
rect 1323 4371 1324 4375
rect 1328 4371 1329 4375
rect 1323 4370 1329 4371
rect 1323 4366 1324 4370
rect 1328 4366 1329 4370
rect 1323 4365 1329 4366
rect 1323 4361 1324 4365
rect 1328 4361 1329 4365
rect 1323 4360 1329 4361
rect 1323 4356 1324 4360
rect 1328 4356 1329 4360
rect 1323 4355 1329 4356
rect 1323 4351 1324 4355
rect 1328 4351 1329 4355
rect 1323 4350 1329 4351
rect 1233 4345 1239 4346
rect 1233 4341 1234 4345
rect 1238 4341 1239 4345
rect 1323 4346 1324 4350
rect 1328 4346 1329 4350
rect 1323 4345 1329 4346
rect 1323 4341 1324 4345
rect 1328 4341 1329 4345
rect 1233 4340 1329 4341
rect 1233 4336 1234 4340
rect 1238 4336 1239 4340
rect 1243 4336 1244 4340
rect 1248 4336 1249 4340
rect 1253 4336 1254 4340
rect 1258 4336 1259 4340
rect 1263 4336 1264 4340
rect 1268 4336 1269 4340
rect 1273 4336 1274 4340
rect 1278 4336 1279 4340
rect 1283 4336 1284 4340
rect 1288 4336 1289 4340
rect 1293 4336 1294 4340
rect 1298 4336 1299 4340
rect 1303 4336 1304 4340
rect 1308 4336 1309 4340
rect 1313 4336 1314 4340
rect 1318 4336 1319 4340
rect 1323 4336 1324 4340
rect 1328 4336 1329 4340
rect 1233 4335 1329 4336
rect 1394 4462 1466 4464
rect 1394 4458 1396 4462
rect 1400 4458 1403 4462
rect 1407 4458 1408 4462
rect 1412 4458 1413 4462
rect 1417 4458 1418 4462
rect 1422 4458 1423 4462
rect 1427 4458 1428 4462
rect 1432 4458 1433 4462
rect 1437 4458 1438 4462
rect 1442 4458 1443 4462
rect 1447 4458 1448 4462
rect 1452 4458 1453 4462
rect 1457 4458 1460 4462
rect 1464 4458 1466 4462
rect 1394 4456 1466 4458
rect 1394 4455 1402 4456
rect 1394 4451 1396 4455
rect 1400 4451 1402 4455
rect 1394 4450 1402 4451
rect 1458 4455 1466 4456
rect 1458 4451 1460 4455
rect 1464 4451 1466 4455
rect 1458 4450 1466 4451
rect 1394 4446 1396 4450
rect 1400 4446 1402 4450
rect 1394 4445 1402 4446
rect 1394 4441 1396 4445
rect 1400 4441 1402 4445
rect 1394 4440 1402 4441
rect 1394 4436 1396 4440
rect 1400 4436 1402 4440
rect 1394 4435 1402 4436
rect 1394 4431 1396 4435
rect 1400 4431 1402 4435
rect 1394 4430 1402 4431
rect 1394 4426 1396 4430
rect 1400 4426 1402 4430
rect 1394 4425 1402 4426
rect 1394 4421 1396 4425
rect 1400 4421 1402 4425
rect 1394 4420 1402 4421
rect 1394 4416 1396 4420
rect 1400 4416 1402 4420
rect 1394 4415 1402 4416
rect 1394 4411 1396 4415
rect 1400 4411 1402 4415
rect 1394 4410 1402 4411
rect 1394 4406 1396 4410
rect 1400 4406 1402 4410
rect 1394 4405 1402 4406
rect 1394 4401 1396 4405
rect 1400 4401 1402 4405
rect 1394 4400 1402 4401
rect 1394 4396 1396 4400
rect 1400 4396 1402 4400
rect 1394 4395 1402 4396
rect 1394 4391 1396 4395
rect 1400 4391 1402 4395
rect 1394 4390 1402 4391
rect 1394 4386 1396 4390
rect 1400 4386 1402 4390
rect 1394 4385 1402 4386
rect 1394 4381 1396 4385
rect 1400 4381 1402 4385
rect 1394 4380 1402 4381
rect 1394 4376 1396 4380
rect 1400 4376 1402 4380
rect 1394 4375 1402 4376
rect 1394 4371 1396 4375
rect 1400 4371 1402 4375
rect 1394 4370 1402 4371
rect 1394 4366 1396 4370
rect 1400 4366 1402 4370
rect 1394 4365 1402 4366
rect 1394 4361 1396 4365
rect 1400 4361 1402 4365
rect 1458 4446 1460 4450
rect 1464 4446 1466 4450
rect 1458 4445 1466 4446
rect 1458 4441 1460 4445
rect 1464 4441 1466 4445
rect 1458 4440 1466 4441
rect 1458 4436 1460 4440
rect 1464 4436 1466 4440
rect 1458 4435 1466 4436
rect 1458 4431 1460 4435
rect 1464 4431 1466 4435
rect 1458 4430 1466 4431
rect 1458 4426 1460 4430
rect 1464 4426 1466 4430
rect 1458 4425 1466 4426
rect 1458 4421 1460 4425
rect 1464 4421 1466 4425
rect 1458 4420 1466 4421
rect 1458 4416 1460 4420
rect 1464 4416 1466 4420
rect 1458 4415 1466 4416
rect 1458 4411 1460 4415
rect 1464 4411 1466 4415
rect 1458 4410 1466 4411
rect 1458 4406 1460 4410
rect 1464 4406 1466 4410
rect 1458 4405 1466 4406
rect 1458 4401 1460 4405
rect 1464 4401 1466 4405
rect 1458 4400 1466 4401
rect 1458 4396 1460 4400
rect 1464 4396 1466 4400
rect 1458 4395 1466 4396
rect 1458 4391 1460 4395
rect 1464 4391 1466 4395
rect 1458 4390 1466 4391
rect 1458 4386 1460 4390
rect 1464 4386 1466 4390
rect 1458 4385 1466 4386
rect 1458 4381 1460 4385
rect 1464 4381 1466 4385
rect 1458 4380 1466 4381
rect 1458 4376 1460 4380
rect 1464 4376 1466 4380
rect 1458 4375 1466 4376
rect 1458 4371 1460 4375
rect 1464 4371 1466 4375
rect 1458 4370 1466 4371
rect 1458 4366 1460 4370
rect 1464 4366 1466 4370
rect 1458 4365 1466 4366
rect 1458 4361 1460 4365
rect 1464 4361 1466 4365
rect 1394 4360 1402 4361
rect 1394 4356 1396 4360
rect 1400 4356 1402 4360
rect 1394 4355 1402 4356
rect 1458 4360 1466 4361
rect 1458 4356 1460 4360
rect 1464 4356 1466 4360
rect 1458 4355 1466 4356
rect 1394 4353 1466 4355
rect 1394 4349 1396 4353
rect 1400 4349 1403 4353
rect 1407 4349 1408 4353
rect 1412 4349 1413 4353
rect 1417 4349 1418 4353
rect 1422 4349 1423 4353
rect 1427 4349 1428 4353
rect 1432 4349 1433 4353
rect 1437 4349 1438 4353
rect 1442 4349 1443 4353
rect 1447 4349 1448 4353
rect 1452 4349 1453 4353
rect 1457 4349 1460 4353
rect 1464 4349 1466 4353
rect 1394 4347 1466 4349
rect 1542 4475 1638 4476
rect 1542 4471 1543 4475
rect 1547 4471 1548 4475
rect 1552 4471 1553 4475
rect 1557 4471 1558 4475
rect 1562 4471 1563 4475
rect 1567 4471 1568 4475
rect 1572 4471 1573 4475
rect 1577 4471 1578 4475
rect 1582 4471 1583 4475
rect 1587 4471 1588 4475
rect 1592 4471 1593 4475
rect 1597 4471 1598 4475
rect 1602 4471 1603 4475
rect 1607 4471 1608 4475
rect 1612 4471 1613 4475
rect 1617 4471 1618 4475
rect 1622 4471 1623 4475
rect 1627 4471 1628 4475
rect 1632 4471 1633 4475
rect 1637 4471 1638 4475
rect 1542 4470 1638 4471
rect 1542 4466 1543 4470
rect 1547 4466 1548 4470
rect 1542 4465 1548 4466
rect 1542 4461 1543 4465
rect 1547 4461 1548 4465
rect 1632 4466 1633 4470
rect 1637 4466 1638 4470
rect 1632 4465 1638 4466
rect 1542 4460 1548 4461
rect 1542 4456 1543 4460
rect 1547 4456 1548 4460
rect 1542 4455 1548 4456
rect 1542 4451 1543 4455
rect 1547 4451 1548 4455
rect 1542 4450 1548 4451
rect 1542 4446 1543 4450
rect 1547 4446 1548 4450
rect 1542 4445 1548 4446
rect 1542 4441 1543 4445
rect 1547 4441 1548 4445
rect 1542 4440 1548 4441
rect 1542 4436 1543 4440
rect 1547 4436 1548 4440
rect 1542 4435 1548 4436
rect 1542 4431 1543 4435
rect 1547 4431 1548 4435
rect 1542 4430 1548 4431
rect 1542 4426 1543 4430
rect 1547 4426 1548 4430
rect 1542 4425 1548 4426
rect 1542 4421 1543 4425
rect 1547 4421 1548 4425
rect 1542 4420 1548 4421
rect 1542 4416 1543 4420
rect 1547 4416 1548 4420
rect 1542 4415 1548 4416
rect 1542 4411 1543 4415
rect 1547 4411 1548 4415
rect 1542 4410 1548 4411
rect 1542 4406 1543 4410
rect 1547 4406 1548 4410
rect 1542 4405 1548 4406
rect 1542 4401 1543 4405
rect 1547 4401 1548 4405
rect 1542 4400 1548 4401
rect 1542 4396 1543 4400
rect 1547 4396 1548 4400
rect 1542 4395 1548 4396
rect 1542 4391 1543 4395
rect 1547 4391 1548 4395
rect 1542 4390 1548 4391
rect 1542 4386 1543 4390
rect 1547 4386 1548 4390
rect 1542 4385 1548 4386
rect 1542 4381 1543 4385
rect 1547 4381 1548 4385
rect 1542 4380 1548 4381
rect 1542 4376 1543 4380
rect 1547 4376 1548 4380
rect 1542 4375 1548 4376
rect 1542 4371 1543 4375
rect 1547 4371 1548 4375
rect 1542 4370 1548 4371
rect 1542 4366 1543 4370
rect 1547 4366 1548 4370
rect 1542 4365 1548 4366
rect 1542 4361 1543 4365
rect 1547 4361 1548 4365
rect 1542 4360 1548 4361
rect 1542 4356 1543 4360
rect 1547 4356 1548 4360
rect 1542 4355 1548 4356
rect 1542 4351 1543 4355
rect 1547 4351 1548 4355
rect 1542 4350 1548 4351
rect 1542 4346 1543 4350
rect 1547 4346 1548 4350
rect 1632 4461 1633 4465
rect 1637 4461 1638 4465
rect 1632 4460 1638 4461
rect 1632 4456 1633 4460
rect 1637 4456 1638 4460
rect 1632 4455 1638 4456
rect 1632 4451 1633 4455
rect 1637 4451 1638 4455
rect 1632 4450 1638 4451
rect 1632 4446 1633 4450
rect 1637 4446 1638 4450
rect 1632 4445 1638 4446
rect 1632 4441 1633 4445
rect 1637 4441 1638 4445
rect 1632 4440 1638 4441
rect 1632 4436 1633 4440
rect 1637 4436 1638 4440
rect 1632 4435 1638 4436
rect 1632 4431 1633 4435
rect 1637 4431 1638 4435
rect 1632 4430 1638 4431
rect 1632 4426 1633 4430
rect 1637 4426 1638 4430
rect 1632 4425 1638 4426
rect 1632 4421 1633 4425
rect 1637 4421 1638 4425
rect 1632 4420 1638 4421
rect 1632 4416 1633 4420
rect 1637 4416 1638 4420
rect 1632 4415 1638 4416
rect 1632 4411 1633 4415
rect 1637 4411 1638 4415
rect 1632 4410 1638 4411
rect 1632 4406 1633 4410
rect 1637 4406 1638 4410
rect 1632 4405 1638 4406
rect 1632 4401 1633 4405
rect 1637 4401 1638 4405
rect 1632 4400 1638 4401
rect 1632 4396 1633 4400
rect 1637 4396 1638 4400
rect 1632 4395 1638 4396
rect 1632 4391 1633 4395
rect 1637 4391 1638 4395
rect 1632 4390 1638 4391
rect 1632 4386 1633 4390
rect 1637 4386 1638 4390
rect 1632 4385 1638 4386
rect 1632 4381 1633 4385
rect 1637 4381 1638 4385
rect 1632 4380 1638 4381
rect 1632 4376 1633 4380
rect 1637 4376 1638 4380
rect 1632 4375 1638 4376
rect 1632 4371 1633 4375
rect 1637 4371 1638 4375
rect 1632 4370 1638 4371
rect 1632 4366 1633 4370
rect 1637 4366 1638 4370
rect 1632 4365 1638 4366
rect 1632 4361 1633 4365
rect 1637 4361 1638 4365
rect 1632 4360 1638 4361
rect 1632 4356 1633 4360
rect 1637 4356 1638 4360
rect 1632 4355 1638 4356
rect 1632 4351 1633 4355
rect 1637 4351 1638 4355
rect 1632 4350 1638 4351
rect 1542 4345 1548 4346
rect 1542 4341 1543 4345
rect 1547 4341 1548 4345
rect 1632 4346 1633 4350
rect 1637 4346 1638 4350
rect 1632 4345 1638 4346
rect 1632 4341 1633 4345
rect 1637 4341 1638 4345
rect 1542 4340 1638 4341
rect 1542 4336 1543 4340
rect 1547 4336 1548 4340
rect 1552 4336 1553 4340
rect 1557 4336 1558 4340
rect 1562 4336 1563 4340
rect 1567 4336 1568 4340
rect 1572 4336 1573 4340
rect 1577 4336 1578 4340
rect 1582 4336 1583 4340
rect 1587 4336 1588 4340
rect 1592 4336 1593 4340
rect 1597 4336 1598 4340
rect 1602 4336 1603 4340
rect 1607 4336 1608 4340
rect 1612 4336 1613 4340
rect 1617 4336 1618 4340
rect 1622 4336 1623 4340
rect 1627 4336 1628 4340
rect 1632 4336 1633 4340
rect 1637 4336 1638 4340
rect 1542 4335 1638 4336
rect 1703 4462 1775 4464
rect 1703 4458 1705 4462
rect 1709 4458 1712 4462
rect 1716 4458 1717 4462
rect 1721 4458 1722 4462
rect 1726 4458 1727 4462
rect 1731 4458 1732 4462
rect 1736 4458 1737 4462
rect 1741 4458 1742 4462
rect 1746 4458 1747 4462
rect 1751 4458 1752 4462
rect 1756 4458 1757 4462
rect 1761 4458 1762 4462
rect 1766 4458 1769 4462
rect 1773 4458 1775 4462
rect 1703 4456 1775 4458
rect 1703 4455 1711 4456
rect 1703 4451 1705 4455
rect 1709 4451 1711 4455
rect 1703 4450 1711 4451
rect 1767 4455 1775 4456
rect 1767 4451 1769 4455
rect 1773 4451 1775 4455
rect 1767 4450 1775 4451
rect 1703 4446 1705 4450
rect 1709 4446 1711 4450
rect 1703 4445 1711 4446
rect 1703 4441 1705 4445
rect 1709 4441 1711 4445
rect 1703 4440 1711 4441
rect 1703 4436 1705 4440
rect 1709 4436 1711 4440
rect 1703 4435 1711 4436
rect 1703 4431 1705 4435
rect 1709 4431 1711 4435
rect 1703 4430 1711 4431
rect 1703 4426 1705 4430
rect 1709 4426 1711 4430
rect 1703 4425 1711 4426
rect 1703 4421 1705 4425
rect 1709 4421 1711 4425
rect 1703 4420 1711 4421
rect 1703 4416 1705 4420
rect 1709 4416 1711 4420
rect 1703 4415 1711 4416
rect 1703 4411 1705 4415
rect 1709 4411 1711 4415
rect 1703 4410 1711 4411
rect 1703 4406 1705 4410
rect 1709 4406 1711 4410
rect 1703 4405 1711 4406
rect 1703 4401 1705 4405
rect 1709 4401 1711 4405
rect 1703 4400 1711 4401
rect 1703 4396 1705 4400
rect 1709 4396 1711 4400
rect 1703 4395 1711 4396
rect 1703 4391 1705 4395
rect 1709 4391 1711 4395
rect 1703 4390 1711 4391
rect 1703 4386 1705 4390
rect 1709 4386 1711 4390
rect 1703 4385 1711 4386
rect 1703 4381 1705 4385
rect 1709 4381 1711 4385
rect 1703 4380 1711 4381
rect 1703 4376 1705 4380
rect 1709 4376 1711 4380
rect 1703 4375 1711 4376
rect 1703 4371 1705 4375
rect 1709 4371 1711 4375
rect 1703 4370 1711 4371
rect 1703 4366 1705 4370
rect 1709 4366 1711 4370
rect 1703 4365 1711 4366
rect 1703 4361 1705 4365
rect 1709 4361 1711 4365
rect 1767 4446 1769 4450
rect 1773 4446 1775 4450
rect 1767 4445 1775 4446
rect 1767 4441 1769 4445
rect 1773 4441 1775 4445
rect 1767 4440 1775 4441
rect 1767 4436 1769 4440
rect 1773 4436 1775 4440
rect 1767 4435 1775 4436
rect 1767 4431 1769 4435
rect 1773 4431 1775 4435
rect 1767 4430 1775 4431
rect 1767 4426 1769 4430
rect 1773 4426 1775 4430
rect 1767 4425 1775 4426
rect 1767 4421 1769 4425
rect 1773 4421 1775 4425
rect 1767 4420 1775 4421
rect 1767 4416 1769 4420
rect 1773 4416 1775 4420
rect 1767 4415 1775 4416
rect 1767 4411 1769 4415
rect 1773 4411 1775 4415
rect 1767 4410 1775 4411
rect 1767 4406 1769 4410
rect 1773 4406 1775 4410
rect 1767 4405 1775 4406
rect 1767 4401 1769 4405
rect 1773 4401 1775 4405
rect 1767 4400 1775 4401
rect 1767 4396 1769 4400
rect 1773 4396 1775 4400
rect 1767 4395 1775 4396
rect 1767 4391 1769 4395
rect 1773 4391 1775 4395
rect 1767 4390 1775 4391
rect 1767 4386 1769 4390
rect 1773 4386 1775 4390
rect 1767 4385 1775 4386
rect 1767 4381 1769 4385
rect 1773 4381 1775 4385
rect 1767 4380 1775 4381
rect 1767 4376 1769 4380
rect 1773 4376 1775 4380
rect 1767 4375 1775 4376
rect 1767 4371 1769 4375
rect 1773 4371 1775 4375
rect 1767 4370 1775 4371
rect 1767 4366 1769 4370
rect 1773 4366 1775 4370
rect 1767 4365 1775 4366
rect 1767 4361 1769 4365
rect 1773 4361 1775 4365
rect 1703 4360 1711 4361
rect 1703 4356 1705 4360
rect 1709 4356 1711 4360
rect 1703 4355 1711 4356
rect 1767 4360 1775 4361
rect 1767 4356 1769 4360
rect 1773 4356 1775 4360
rect 1767 4355 1775 4356
rect 1703 4353 1775 4355
rect 1703 4349 1705 4353
rect 1709 4349 1712 4353
rect 1716 4349 1717 4353
rect 1721 4349 1722 4353
rect 1726 4349 1727 4353
rect 1731 4349 1732 4353
rect 1736 4349 1737 4353
rect 1741 4349 1742 4353
rect 1746 4349 1747 4353
rect 1751 4349 1752 4353
rect 1756 4349 1757 4353
rect 1761 4349 1762 4353
rect 1766 4349 1769 4353
rect 1773 4349 1775 4353
rect 1703 4347 1775 4349
rect 1851 4475 1947 4476
rect 1851 4471 1852 4475
rect 1856 4471 1857 4475
rect 1861 4471 1862 4475
rect 1866 4471 1867 4475
rect 1871 4471 1872 4475
rect 1876 4471 1877 4475
rect 1881 4471 1882 4475
rect 1886 4471 1887 4475
rect 1891 4471 1892 4475
rect 1896 4471 1897 4475
rect 1901 4471 1902 4475
rect 1906 4471 1907 4475
rect 1911 4471 1912 4475
rect 1916 4471 1917 4475
rect 1921 4471 1922 4475
rect 1926 4471 1927 4475
rect 1931 4471 1932 4475
rect 1936 4471 1937 4475
rect 1941 4471 1942 4475
rect 1946 4471 1947 4475
rect 1851 4470 1947 4471
rect 1851 4466 1852 4470
rect 1856 4466 1857 4470
rect 1851 4465 1857 4466
rect 1851 4461 1852 4465
rect 1856 4461 1857 4465
rect 1941 4466 1942 4470
rect 1946 4466 1947 4470
rect 1941 4465 1947 4466
rect 1851 4460 1857 4461
rect 1851 4456 1852 4460
rect 1856 4456 1857 4460
rect 1851 4455 1857 4456
rect 1851 4451 1852 4455
rect 1856 4451 1857 4455
rect 1851 4450 1857 4451
rect 1851 4446 1852 4450
rect 1856 4446 1857 4450
rect 1851 4445 1857 4446
rect 1851 4441 1852 4445
rect 1856 4441 1857 4445
rect 1851 4440 1857 4441
rect 1851 4436 1852 4440
rect 1856 4436 1857 4440
rect 1851 4435 1857 4436
rect 1851 4431 1852 4435
rect 1856 4431 1857 4435
rect 1851 4430 1857 4431
rect 1851 4426 1852 4430
rect 1856 4426 1857 4430
rect 1851 4425 1857 4426
rect 1851 4421 1852 4425
rect 1856 4421 1857 4425
rect 1851 4420 1857 4421
rect 1851 4416 1852 4420
rect 1856 4416 1857 4420
rect 1851 4415 1857 4416
rect 1851 4411 1852 4415
rect 1856 4411 1857 4415
rect 1851 4410 1857 4411
rect 1851 4406 1852 4410
rect 1856 4406 1857 4410
rect 1851 4405 1857 4406
rect 1851 4401 1852 4405
rect 1856 4401 1857 4405
rect 1851 4400 1857 4401
rect 1851 4396 1852 4400
rect 1856 4396 1857 4400
rect 1851 4395 1857 4396
rect 1851 4391 1852 4395
rect 1856 4391 1857 4395
rect 1851 4390 1857 4391
rect 1851 4386 1852 4390
rect 1856 4386 1857 4390
rect 1851 4385 1857 4386
rect 1851 4381 1852 4385
rect 1856 4381 1857 4385
rect 1851 4380 1857 4381
rect 1851 4376 1852 4380
rect 1856 4376 1857 4380
rect 1851 4375 1857 4376
rect 1851 4371 1852 4375
rect 1856 4371 1857 4375
rect 1851 4370 1857 4371
rect 1851 4366 1852 4370
rect 1856 4366 1857 4370
rect 1851 4365 1857 4366
rect 1851 4361 1852 4365
rect 1856 4361 1857 4365
rect 1851 4360 1857 4361
rect 1851 4356 1852 4360
rect 1856 4356 1857 4360
rect 1851 4355 1857 4356
rect 1851 4351 1852 4355
rect 1856 4351 1857 4355
rect 1851 4350 1857 4351
rect 1851 4346 1852 4350
rect 1856 4346 1857 4350
rect 1941 4461 1942 4465
rect 1946 4461 1947 4465
rect 1941 4460 1947 4461
rect 1941 4456 1942 4460
rect 1946 4456 1947 4460
rect 1941 4455 1947 4456
rect 1941 4451 1942 4455
rect 1946 4451 1947 4455
rect 1941 4450 1947 4451
rect 1941 4446 1942 4450
rect 1946 4446 1947 4450
rect 1941 4445 1947 4446
rect 1941 4441 1942 4445
rect 1946 4441 1947 4445
rect 1941 4440 1947 4441
rect 1941 4436 1942 4440
rect 1946 4436 1947 4440
rect 1941 4435 1947 4436
rect 1941 4431 1942 4435
rect 1946 4431 1947 4435
rect 1941 4430 1947 4431
rect 1941 4426 1942 4430
rect 1946 4426 1947 4430
rect 1941 4425 1947 4426
rect 1941 4421 1942 4425
rect 1946 4421 1947 4425
rect 1941 4420 1947 4421
rect 1941 4416 1942 4420
rect 1946 4416 1947 4420
rect 1941 4415 1947 4416
rect 1941 4411 1942 4415
rect 1946 4411 1947 4415
rect 1941 4410 1947 4411
rect 1941 4406 1942 4410
rect 1946 4406 1947 4410
rect 1941 4405 1947 4406
rect 1941 4401 1942 4405
rect 1946 4401 1947 4405
rect 1941 4400 1947 4401
rect 1941 4396 1942 4400
rect 1946 4396 1947 4400
rect 1941 4395 1947 4396
rect 1941 4391 1942 4395
rect 1946 4391 1947 4395
rect 1941 4390 1947 4391
rect 1941 4386 1942 4390
rect 1946 4386 1947 4390
rect 1941 4385 1947 4386
rect 1941 4381 1942 4385
rect 1946 4381 1947 4385
rect 1941 4380 1947 4381
rect 1941 4376 1942 4380
rect 1946 4376 1947 4380
rect 1941 4375 1947 4376
rect 1941 4371 1942 4375
rect 1946 4371 1947 4375
rect 1941 4370 1947 4371
rect 1941 4366 1942 4370
rect 1946 4366 1947 4370
rect 1941 4365 1947 4366
rect 1941 4361 1942 4365
rect 1946 4361 1947 4365
rect 1941 4360 1947 4361
rect 1941 4356 1942 4360
rect 1946 4356 1947 4360
rect 1941 4355 1947 4356
rect 1941 4351 1942 4355
rect 1946 4351 1947 4355
rect 1941 4350 1947 4351
rect 1851 4345 1857 4346
rect 1851 4341 1852 4345
rect 1856 4341 1857 4345
rect 1941 4346 1942 4350
rect 1946 4346 1947 4350
rect 1941 4345 1947 4346
rect 1941 4341 1942 4345
rect 1946 4341 1947 4345
rect 1851 4340 1947 4341
rect 1851 4336 1852 4340
rect 1856 4336 1857 4340
rect 1861 4336 1862 4340
rect 1866 4336 1867 4340
rect 1871 4336 1872 4340
rect 1876 4336 1877 4340
rect 1881 4336 1882 4340
rect 1886 4336 1887 4340
rect 1891 4336 1892 4340
rect 1896 4336 1897 4340
rect 1901 4336 1902 4340
rect 1906 4336 1907 4340
rect 1911 4336 1912 4340
rect 1916 4336 1917 4340
rect 1921 4336 1922 4340
rect 1926 4336 1927 4340
rect 1931 4336 1932 4340
rect 1936 4336 1937 4340
rect 1941 4336 1942 4340
rect 1946 4336 1947 4340
rect 1851 4335 1947 4336
rect 2012 4462 2084 4464
rect 2012 4458 2014 4462
rect 2018 4458 2021 4462
rect 2025 4458 2026 4462
rect 2030 4458 2031 4462
rect 2035 4458 2036 4462
rect 2040 4458 2041 4462
rect 2045 4458 2046 4462
rect 2050 4458 2051 4462
rect 2055 4458 2056 4462
rect 2060 4458 2061 4462
rect 2065 4458 2066 4462
rect 2070 4458 2071 4462
rect 2075 4458 2078 4462
rect 2082 4458 2084 4462
rect 2012 4456 2084 4458
rect 2012 4455 2020 4456
rect 2012 4451 2014 4455
rect 2018 4451 2020 4455
rect 2012 4450 2020 4451
rect 2076 4455 2084 4456
rect 2076 4451 2078 4455
rect 2082 4451 2084 4455
rect 2076 4450 2084 4451
rect 2012 4446 2014 4450
rect 2018 4446 2020 4450
rect 2012 4445 2020 4446
rect 2012 4441 2014 4445
rect 2018 4441 2020 4445
rect 2012 4440 2020 4441
rect 2012 4436 2014 4440
rect 2018 4436 2020 4440
rect 2012 4435 2020 4436
rect 2012 4431 2014 4435
rect 2018 4431 2020 4435
rect 2012 4430 2020 4431
rect 2012 4426 2014 4430
rect 2018 4426 2020 4430
rect 2012 4425 2020 4426
rect 2012 4421 2014 4425
rect 2018 4421 2020 4425
rect 2012 4420 2020 4421
rect 2012 4416 2014 4420
rect 2018 4416 2020 4420
rect 2012 4415 2020 4416
rect 2012 4411 2014 4415
rect 2018 4411 2020 4415
rect 2012 4410 2020 4411
rect 2012 4406 2014 4410
rect 2018 4406 2020 4410
rect 2012 4405 2020 4406
rect 2012 4401 2014 4405
rect 2018 4401 2020 4405
rect 2012 4400 2020 4401
rect 2012 4396 2014 4400
rect 2018 4396 2020 4400
rect 2012 4395 2020 4396
rect 2012 4391 2014 4395
rect 2018 4391 2020 4395
rect 2012 4390 2020 4391
rect 2012 4386 2014 4390
rect 2018 4386 2020 4390
rect 2012 4385 2020 4386
rect 2012 4381 2014 4385
rect 2018 4381 2020 4385
rect 2012 4380 2020 4381
rect 2012 4376 2014 4380
rect 2018 4376 2020 4380
rect 2012 4375 2020 4376
rect 2012 4371 2014 4375
rect 2018 4371 2020 4375
rect 2012 4370 2020 4371
rect 2012 4366 2014 4370
rect 2018 4366 2020 4370
rect 2012 4365 2020 4366
rect 2012 4361 2014 4365
rect 2018 4361 2020 4365
rect 2076 4446 2078 4450
rect 2082 4446 2084 4450
rect 2076 4445 2084 4446
rect 2076 4441 2078 4445
rect 2082 4441 2084 4445
rect 2076 4440 2084 4441
rect 2076 4436 2078 4440
rect 2082 4436 2084 4440
rect 2076 4435 2084 4436
rect 2076 4431 2078 4435
rect 2082 4431 2084 4435
rect 2076 4430 2084 4431
rect 2076 4426 2078 4430
rect 2082 4426 2084 4430
rect 2076 4425 2084 4426
rect 2076 4421 2078 4425
rect 2082 4421 2084 4425
rect 2076 4420 2084 4421
rect 2076 4416 2078 4420
rect 2082 4416 2084 4420
rect 2076 4415 2084 4416
rect 2076 4411 2078 4415
rect 2082 4411 2084 4415
rect 2076 4410 2084 4411
rect 2076 4406 2078 4410
rect 2082 4406 2084 4410
rect 2076 4405 2084 4406
rect 2076 4401 2078 4405
rect 2082 4401 2084 4405
rect 2076 4400 2084 4401
rect 2076 4396 2078 4400
rect 2082 4396 2084 4400
rect 2076 4395 2084 4396
rect 2076 4391 2078 4395
rect 2082 4391 2084 4395
rect 2076 4390 2084 4391
rect 2076 4386 2078 4390
rect 2082 4386 2084 4390
rect 2076 4385 2084 4386
rect 2076 4381 2078 4385
rect 2082 4381 2084 4385
rect 2076 4380 2084 4381
rect 2076 4376 2078 4380
rect 2082 4376 2084 4380
rect 2076 4375 2084 4376
rect 2076 4371 2078 4375
rect 2082 4371 2084 4375
rect 2076 4370 2084 4371
rect 2076 4366 2078 4370
rect 2082 4366 2084 4370
rect 2076 4365 2084 4366
rect 2076 4361 2078 4365
rect 2082 4361 2084 4365
rect 2012 4360 2020 4361
rect 2012 4356 2014 4360
rect 2018 4356 2020 4360
rect 2012 4355 2020 4356
rect 2076 4360 2084 4361
rect 2076 4356 2078 4360
rect 2082 4356 2084 4360
rect 2076 4355 2084 4356
rect 2012 4353 2084 4355
rect 2012 4349 2014 4353
rect 2018 4349 2021 4353
rect 2025 4349 2026 4353
rect 2030 4349 2031 4353
rect 2035 4349 2036 4353
rect 2040 4349 2041 4353
rect 2045 4349 2046 4353
rect 2050 4349 2051 4353
rect 2055 4349 2056 4353
rect 2060 4349 2061 4353
rect 2065 4349 2066 4353
rect 2070 4349 2071 4353
rect 2075 4349 2078 4353
rect 2082 4349 2084 4353
rect 2012 4347 2084 4349
rect 2160 4475 2256 4476
rect 2160 4471 2161 4475
rect 2165 4471 2166 4475
rect 2170 4471 2171 4475
rect 2175 4471 2176 4475
rect 2180 4471 2181 4475
rect 2185 4471 2186 4475
rect 2190 4471 2191 4475
rect 2195 4471 2196 4475
rect 2200 4471 2201 4475
rect 2205 4471 2206 4475
rect 2210 4471 2211 4475
rect 2215 4471 2216 4475
rect 2220 4471 2221 4475
rect 2225 4471 2226 4475
rect 2230 4471 2231 4475
rect 2235 4471 2236 4475
rect 2240 4471 2241 4475
rect 2245 4471 2246 4475
rect 2250 4471 2251 4475
rect 2255 4471 2256 4475
rect 2160 4470 2256 4471
rect 2160 4466 2161 4470
rect 2165 4466 2166 4470
rect 2160 4465 2166 4466
rect 2160 4461 2161 4465
rect 2165 4461 2166 4465
rect 2250 4466 2251 4470
rect 2255 4466 2256 4470
rect 2250 4465 2256 4466
rect 2160 4460 2166 4461
rect 2160 4456 2161 4460
rect 2165 4456 2166 4460
rect 2160 4455 2166 4456
rect 2160 4451 2161 4455
rect 2165 4451 2166 4455
rect 2160 4450 2166 4451
rect 2160 4446 2161 4450
rect 2165 4446 2166 4450
rect 2160 4445 2166 4446
rect 2160 4441 2161 4445
rect 2165 4441 2166 4445
rect 2160 4440 2166 4441
rect 2160 4436 2161 4440
rect 2165 4436 2166 4440
rect 2160 4435 2166 4436
rect 2160 4431 2161 4435
rect 2165 4431 2166 4435
rect 2160 4430 2166 4431
rect 2160 4426 2161 4430
rect 2165 4426 2166 4430
rect 2160 4425 2166 4426
rect 2160 4421 2161 4425
rect 2165 4421 2166 4425
rect 2160 4420 2166 4421
rect 2160 4416 2161 4420
rect 2165 4416 2166 4420
rect 2160 4415 2166 4416
rect 2160 4411 2161 4415
rect 2165 4411 2166 4415
rect 2160 4410 2166 4411
rect 2160 4406 2161 4410
rect 2165 4406 2166 4410
rect 2160 4405 2166 4406
rect 2160 4401 2161 4405
rect 2165 4401 2166 4405
rect 2160 4400 2166 4401
rect 2160 4396 2161 4400
rect 2165 4396 2166 4400
rect 2160 4395 2166 4396
rect 2160 4391 2161 4395
rect 2165 4391 2166 4395
rect 2160 4390 2166 4391
rect 2160 4386 2161 4390
rect 2165 4386 2166 4390
rect 2160 4385 2166 4386
rect 2160 4381 2161 4385
rect 2165 4381 2166 4385
rect 2160 4380 2166 4381
rect 2160 4376 2161 4380
rect 2165 4376 2166 4380
rect 2160 4375 2166 4376
rect 2160 4371 2161 4375
rect 2165 4371 2166 4375
rect 2160 4370 2166 4371
rect 2160 4366 2161 4370
rect 2165 4366 2166 4370
rect 2160 4365 2166 4366
rect 2160 4361 2161 4365
rect 2165 4361 2166 4365
rect 2160 4360 2166 4361
rect 2160 4356 2161 4360
rect 2165 4356 2166 4360
rect 2160 4355 2166 4356
rect 2160 4351 2161 4355
rect 2165 4351 2166 4355
rect 2160 4350 2166 4351
rect 2160 4346 2161 4350
rect 2165 4346 2166 4350
rect 2250 4461 2251 4465
rect 2255 4461 2256 4465
rect 2250 4460 2256 4461
rect 2250 4456 2251 4460
rect 2255 4456 2256 4460
rect 2250 4455 2256 4456
rect 2250 4451 2251 4455
rect 2255 4451 2256 4455
rect 2250 4450 2256 4451
rect 2250 4446 2251 4450
rect 2255 4446 2256 4450
rect 2250 4445 2256 4446
rect 2250 4441 2251 4445
rect 2255 4441 2256 4445
rect 2250 4440 2256 4441
rect 2250 4436 2251 4440
rect 2255 4436 2256 4440
rect 2250 4435 2256 4436
rect 2250 4431 2251 4435
rect 2255 4431 2256 4435
rect 2250 4430 2256 4431
rect 2250 4426 2251 4430
rect 2255 4426 2256 4430
rect 2250 4425 2256 4426
rect 2250 4421 2251 4425
rect 2255 4421 2256 4425
rect 2250 4420 2256 4421
rect 2250 4416 2251 4420
rect 2255 4416 2256 4420
rect 2250 4415 2256 4416
rect 2250 4411 2251 4415
rect 2255 4411 2256 4415
rect 2250 4410 2256 4411
rect 2250 4406 2251 4410
rect 2255 4406 2256 4410
rect 2250 4405 2256 4406
rect 2250 4401 2251 4405
rect 2255 4401 2256 4405
rect 2250 4400 2256 4401
rect 2250 4396 2251 4400
rect 2255 4396 2256 4400
rect 2250 4395 2256 4396
rect 2250 4391 2251 4395
rect 2255 4391 2256 4395
rect 2250 4390 2256 4391
rect 2250 4386 2251 4390
rect 2255 4386 2256 4390
rect 2250 4385 2256 4386
rect 2250 4381 2251 4385
rect 2255 4381 2256 4385
rect 2250 4380 2256 4381
rect 2250 4376 2251 4380
rect 2255 4376 2256 4380
rect 2250 4375 2256 4376
rect 2250 4371 2251 4375
rect 2255 4371 2256 4375
rect 2250 4370 2256 4371
rect 2250 4366 2251 4370
rect 2255 4366 2256 4370
rect 2250 4365 2256 4366
rect 2250 4361 2251 4365
rect 2255 4361 2256 4365
rect 2250 4360 2256 4361
rect 2250 4356 2251 4360
rect 2255 4356 2256 4360
rect 2250 4355 2256 4356
rect 2250 4351 2251 4355
rect 2255 4351 2256 4355
rect 2250 4350 2256 4351
rect 2160 4345 2166 4346
rect 2160 4341 2161 4345
rect 2165 4341 2166 4345
rect 2250 4346 2251 4350
rect 2255 4346 2256 4350
rect 2250 4345 2256 4346
rect 2250 4341 2251 4345
rect 2255 4341 2256 4345
rect 2160 4340 2256 4341
rect 2160 4336 2161 4340
rect 2165 4336 2166 4340
rect 2170 4336 2171 4340
rect 2175 4336 2176 4340
rect 2180 4336 2181 4340
rect 2185 4336 2186 4340
rect 2190 4336 2191 4340
rect 2195 4336 2196 4340
rect 2200 4336 2201 4340
rect 2205 4336 2206 4340
rect 2210 4336 2211 4340
rect 2215 4336 2216 4340
rect 2220 4336 2221 4340
rect 2225 4336 2226 4340
rect 2230 4336 2231 4340
rect 2235 4336 2236 4340
rect 2240 4336 2241 4340
rect 2245 4336 2246 4340
rect 2250 4336 2251 4340
rect 2255 4336 2256 4340
rect 2160 4335 2256 4336
rect 2321 4462 2393 4464
rect 2321 4458 2323 4462
rect 2327 4458 2330 4462
rect 2334 4458 2335 4462
rect 2339 4458 2340 4462
rect 2344 4458 2345 4462
rect 2349 4458 2350 4462
rect 2354 4458 2355 4462
rect 2359 4458 2360 4462
rect 2364 4458 2365 4462
rect 2369 4458 2370 4462
rect 2374 4458 2375 4462
rect 2379 4458 2380 4462
rect 2384 4458 2387 4462
rect 2391 4458 2393 4462
rect 2321 4456 2393 4458
rect 2321 4455 2329 4456
rect 2321 4451 2323 4455
rect 2327 4451 2329 4455
rect 2321 4450 2329 4451
rect 2385 4455 2393 4456
rect 2385 4451 2387 4455
rect 2391 4451 2393 4455
rect 2385 4450 2393 4451
rect 2321 4446 2323 4450
rect 2327 4446 2329 4450
rect 2321 4445 2329 4446
rect 2321 4441 2323 4445
rect 2327 4441 2329 4445
rect 2321 4440 2329 4441
rect 2321 4436 2323 4440
rect 2327 4436 2329 4440
rect 2321 4435 2329 4436
rect 2321 4431 2323 4435
rect 2327 4431 2329 4435
rect 2321 4430 2329 4431
rect 2321 4426 2323 4430
rect 2327 4426 2329 4430
rect 2321 4425 2329 4426
rect 2321 4421 2323 4425
rect 2327 4421 2329 4425
rect 2321 4420 2329 4421
rect 2321 4416 2323 4420
rect 2327 4416 2329 4420
rect 2321 4415 2329 4416
rect 2321 4411 2323 4415
rect 2327 4411 2329 4415
rect 2321 4410 2329 4411
rect 2321 4406 2323 4410
rect 2327 4406 2329 4410
rect 2321 4405 2329 4406
rect 2321 4401 2323 4405
rect 2327 4401 2329 4405
rect 2321 4400 2329 4401
rect 2321 4396 2323 4400
rect 2327 4396 2329 4400
rect 2321 4395 2329 4396
rect 2321 4391 2323 4395
rect 2327 4391 2329 4395
rect 2321 4390 2329 4391
rect 2321 4386 2323 4390
rect 2327 4386 2329 4390
rect 2321 4385 2329 4386
rect 2321 4381 2323 4385
rect 2327 4381 2329 4385
rect 2321 4380 2329 4381
rect 2321 4376 2323 4380
rect 2327 4376 2329 4380
rect 2321 4375 2329 4376
rect 2321 4371 2323 4375
rect 2327 4371 2329 4375
rect 2321 4370 2329 4371
rect 2321 4366 2323 4370
rect 2327 4366 2329 4370
rect 2321 4365 2329 4366
rect 2321 4361 2323 4365
rect 2327 4361 2329 4365
rect 2385 4446 2387 4450
rect 2391 4446 2393 4450
rect 2385 4445 2393 4446
rect 2385 4441 2387 4445
rect 2391 4441 2393 4445
rect 2385 4440 2393 4441
rect 2385 4436 2387 4440
rect 2391 4436 2393 4440
rect 2385 4435 2393 4436
rect 2385 4431 2387 4435
rect 2391 4431 2393 4435
rect 2385 4430 2393 4431
rect 2385 4426 2387 4430
rect 2391 4426 2393 4430
rect 2385 4425 2393 4426
rect 2385 4421 2387 4425
rect 2391 4421 2393 4425
rect 2385 4420 2393 4421
rect 2385 4416 2387 4420
rect 2391 4416 2393 4420
rect 2385 4415 2393 4416
rect 2385 4411 2387 4415
rect 2391 4411 2393 4415
rect 2385 4410 2393 4411
rect 2385 4406 2387 4410
rect 2391 4406 2393 4410
rect 2385 4405 2393 4406
rect 2385 4401 2387 4405
rect 2391 4401 2393 4405
rect 2385 4400 2393 4401
rect 2385 4396 2387 4400
rect 2391 4396 2393 4400
rect 2385 4395 2393 4396
rect 2385 4391 2387 4395
rect 2391 4391 2393 4395
rect 2385 4390 2393 4391
rect 2385 4386 2387 4390
rect 2391 4386 2393 4390
rect 2385 4385 2393 4386
rect 2385 4381 2387 4385
rect 2391 4381 2393 4385
rect 2385 4380 2393 4381
rect 2385 4376 2387 4380
rect 2391 4376 2393 4380
rect 2385 4375 2393 4376
rect 2385 4371 2387 4375
rect 2391 4371 2393 4375
rect 2385 4370 2393 4371
rect 2385 4366 2387 4370
rect 2391 4366 2393 4370
rect 2385 4365 2393 4366
rect 2385 4361 2387 4365
rect 2391 4361 2393 4365
rect 2321 4360 2329 4361
rect 2321 4356 2323 4360
rect 2327 4356 2329 4360
rect 2321 4355 2329 4356
rect 2385 4360 2393 4361
rect 2385 4356 2387 4360
rect 2391 4356 2393 4360
rect 2385 4355 2393 4356
rect 2321 4353 2393 4355
rect 2321 4349 2323 4353
rect 2327 4349 2330 4353
rect 2334 4349 2335 4353
rect 2339 4349 2340 4353
rect 2344 4349 2345 4353
rect 2349 4349 2350 4353
rect 2354 4349 2355 4353
rect 2359 4349 2360 4353
rect 2364 4349 2365 4353
rect 2369 4349 2370 4353
rect 2374 4349 2375 4353
rect 2379 4349 2380 4353
rect 2384 4349 2387 4353
rect 2391 4349 2393 4353
rect 2321 4347 2393 4349
rect 2469 4475 2565 4476
rect 2469 4471 2470 4475
rect 2474 4471 2475 4475
rect 2479 4471 2480 4475
rect 2484 4471 2485 4475
rect 2489 4471 2490 4475
rect 2494 4471 2495 4475
rect 2499 4471 2500 4475
rect 2504 4471 2505 4475
rect 2509 4471 2510 4475
rect 2514 4471 2515 4475
rect 2519 4471 2520 4475
rect 2524 4471 2525 4475
rect 2529 4471 2530 4475
rect 2534 4471 2535 4475
rect 2539 4471 2540 4475
rect 2544 4471 2545 4475
rect 2549 4471 2550 4475
rect 2554 4471 2555 4475
rect 2559 4471 2560 4475
rect 2564 4471 2565 4475
rect 2469 4470 2565 4471
rect 2469 4466 2470 4470
rect 2474 4466 2475 4470
rect 2469 4465 2475 4466
rect 2469 4461 2470 4465
rect 2474 4461 2475 4465
rect 2559 4466 2560 4470
rect 2564 4466 2565 4470
rect 2559 4465 2565 4466
rect 2469 4460 2475 4461
rect 2469 4456 2470 4460
rect 2474 4456 2475 4460
rect 2469 4455 2475 4456
rect 2469 4451 2470 4455
rect 2474 4451 2475 4455
rect 2469 4450 2475 4451
rect 2469 4446 2470 4450
rect 2474 4446 2475 4450
rect 2469 4445 2475 4446
rect 2469 4441 2470 4445
rect 2474 4441 2475 4445
rect 2469 4440 2475 4441
rect 2469 4436 2470 4440
rect 2474 4436 2475 4440
rect 2469 4435 2475 4436
rect 2469 4431 2470 4435
rect 2474 4431 2475 4435
rect 2469 4430 2475 4431
rect 2469 4426 2470 4430
rect 2474 4426 2475 4430
rect 2469 4425 2475 4426
rect 2469 4421 2470 4425
rect 2474 4421 2475 4425
rect 2469 4420 2475 4421
rect 2469 4416 2470 4420
rect 2474 4416 2475 4420
rect 2469 4415 2475 4416
rect 2469 4411 2470 4415
rect 2474 4411 2475 4415
rect 2469 4410 2475 4411
rect 2469 4406 2470 4410
rect 2474 4406 2475 4410
rect 2469 4405 2475 4406
rect 2469 4401 2470 4405
rect 2474 4401 2475 4405
rect 2469 4400 2475 4401
rect 2469 4396 2470 4400
rect 2474 4396 2475 4400
rect 2469 4395 2475 4396
rect 2469 4391 2470 4395
rect 2474 4391 2475 4395
rect 2469 4390 2475 4391
rect 2469 4386 2470 4390
rect 2474 4386 2475 4390
rect 2469 4385 2475 4386
rect 2469 4381 2470 4385
rect 2474 4381 2475 4385
rect 2469 4380 2475 4381
rect 2469 4376 2470 4380
rect 2474 4376 2475 4380
rect 2469 4375 2475 4376
rect 2469 4371 2470 4375
rect 2474 4371 2475 4375
rect 2469 4370 2475 4371
rect 2469 4366 2470 4370
rect 2474 4366 2475 4370
rect 2469 4365 2475 4366
rect 2469 4361 2470 4365
rect 2474 4361 2475 4365
rect 2469 4360 2475 4361
rect 2469 4356 2470 4360
rect 2474 4356 2475 4360
rect 2469 4355 2475 4356
rect 2469 4351 2470 4355
rect 2474 4351 2475 4355
rect 2469 4350 2475 4351
rect 2469 4346 2470 4350
rect 2474 4346 2475 4350
rect 2559 4461 2560 4465
rect 2564 4461 2565 4465
rect 2559 4460 2565 4461
rect 2559 4456 2560 4460
rect 2564 4456 2565 4460
rect 2559 4455 2565 4456
rect 2559 4451 2560 4455
rect 2564 4451 2565 4455
rect 2559 4450 2565 4451
rect 2559 4446 2560 4450
rect 2564 4446 2565 4450
rect 2559 4445 2565 4446
rect 2559 4441 2560 4445
rect 2564 4441 2565 4445
rect 2559 4440 2565 4441
rect 2559 4436 2560 4440
rect 2564 4436 2565 4440
rect 2559 4435 2565 4436
rect 2559 4431 2560 4435
rect 2564 4431 2565 4435
rect 2559 4430 2565 4431
rect 2559 4426 2560 4430
rect 2564 4426 2565 4430
rect 2559 4425 2565 4426
rect 2559 4421 2560 4425
rect 2564 4421 2565 4425
rect 2559 4420 2565 4421
rect 2559 4416 2560 4420
rect 2564 4416 2565 4420
rect 2559 4415 2565 4416
rect 2559 4411 2560 4415
rect 2564 4411 2565 4415
rect 2559 4410 2565 4411
rect 2559 4406 2560 4410
rect 2564 4406 2565 4410
rect 2559 4405 2565 4406
rect 2559 4401 2560 4405
rect 2564 4401 2565 4405
rect 2559 4400 2565 4401
rect 2559 4396 2560 4400
rect 2564 4396 2565 4400
rect 2559 4395 2565 4396
rect 2559 4391 2560 4395
rect 2564 4391 2565 4395
rect 2559 4390 2565 4391
rect 2559 4386 2560 4390
rect 2564 4386 2565 4390
rect 2559 4385 2565 4386
rect 2559 4381 2560 4385
rect 2564 4381 2565 4385
rect 2559 4380 2565 4381
rect 2559 4376 2560 4380
rect 2564 4376 2565 4380
rect 2559 4375 2565 4376
rect 2559 4371 2560 4375
rect 2564 4371 2565 4375
rect 2559 4370 2565 4371
rect 2559 4366 2560 4370
rect 2564 4366 2565 4370
rect 2559 4365 2565 4366
rect 2559 4361 2560 4365
rect 2564 4361 2565 4365
rect 2559 4360 2565 4361
rect 2559 4356 2560 4360
rect 2564 4356 2565 4360
rect 2559 4355 2565 4356
rect 2559 4351 2560 4355
rect 2564 4351 2565 4355
rect 2559 4350 2565 4351
rect 2469 4345 2475 4346
rect 2469 4341 2470 4345
rect 2474 4341 2475 4345
rect 2559 4346 2560 4350
rect 2564 4346 2565 4350
rect 2559 4345 2565 4346
rect 2559 4341 2560 4345
rect 2564 4341 2565 4345
rect 2469 4340 2565 4341
rect 2469 4336 2470 4340
rect 2474 4336 2475 4340
rect 2479 4336 2480 4340
rect 2484 4336 2485 4340
rect 2489 4336 2490 4340
rect 2494 4336 2495 4340
rect 2499 4336 2500 4340
rect 2504 4336 2505 4340
rect 2509 4336 2510 4340
rect 2514 4336 2515 4340
rect 2519 4336 2520 4340
rect 2524 4336 2525 4340
rect 2529 4336 2530 4340
rect 2534 4336 2535 4340
rect 2539 4336 2540 4340
rect 2544 4336 2545 4340
rect 2549 4336 2550 4340
rect 2554 4336 2555 4340
rect 2559 4336 2560 4340
rect 2564 4336 2565 4340
rect 2469 4335 2565 4336
rect 2630 4462 2702 4464
rect 2630 4458 2632 4462
rect 2636 4458 2639 4462
rect 2643 4458 2644 4462
rect 2648 4458 2649 4462
rect 2653 4458 2654 4462
rect 2658 4458 2659 4462
rect 2663 4458 2664 4462
rect 2668 4458 2669 4462
rect 2673 4458 2674 4462
rect 2678 4458 2679 4462
rect 2683 4458 2684 4462
rect 2688 4458 2689 4462
rect 2693 4458 2696 4462
rect 2700 4458 2702 4462
rect 2630 4456 2702 4458
rect 2630 4455 2638 4456
rect 2630 4451 2632 4455
rect 2636 4451 2638 4455
rect 2630 4450 2638 4451
rect 2694 4455 2702 4456
rect 2694 4451 2696 4455
rect 2700 4451 2702 4455
rect 2694 4450 2702 4451
rect 2630 4446 2632 4450
rect 2636 4446 2638 4450
rect 2630 4445 2638 4446
rect 2630 4441 2632 4445
rect 2636 4441 2638 4445
rect 2630 4440 2638 4441
rect 2630 4436 2632 4440
rect 2636 4436 2638 4440
rect 2630 4435 2638 4436
rect 2630 4431 2632 4435
rect 2636 4431 2638 4435
rect 2630 4430 2638 4431
rect 2630 4426 2632 4430
rect 2636 4426 2638 4430
rect 2630 4425 2638 4426
rect 2630 4421 2632 4425
rect 2636 4421 2638 4425
rect 2630 4420 2638 4421
rect 2630 4416 2632 4420
rect 2636 4416 2638 4420
rect 2630 4415 2638 4416
rect 2630 4411 2632 4415
rect 2636 4411 2638 4415
rect 2630 4410 2638 4411
rect 2630 4406 2632 4410
rect 2636 4406 2638 4410
rect 2630 4405 2638 4406
rect 2630 4401 2632 4405
rect 2636 4401 2638 4405
rect 2630 4400 2638 4401
rect 2630 4396 2632 4400
rect 2636 4396 2638 4400
rect 2630 4395 2638 4396
rect 2630 4391 2632 4395
rect 2636 4391 2638 4395
rect 2630 4390 2638 4391
rect 2630 4386 2632 4390
rect 2636 4386 2638 4390
rect 2630 4385 2638 4386
rect 2630 4381 2632 4385
rect 2636 4381 2638 4385
rect 2630 4380 2638 4381
rect 2630 4376 2632 4380
rect 2636 4376 2638 4380
rect 2630 4375 2638 4376
rect 2630 4371 2632 4375
rect 2636 4371 2638 4375
rect 2630 4370 2638 4371
rect 2630 4366 2632 4370
rect 2636 4366 2638 4370
rect 2630 4365 2638 4366
rect 2630 4361 2632 4365
rect 2636 4361 2638 4365
rect 2694 4446 2696 4450
rect 2700 4446 2702 4450
rect 2694 4445 2702 4446
rect 2694 4441 2696 4445
rect 2700 4441 2702 4445
rect 2694 4440 2702 4441
rect 2694 4436 2696 4440
rect 2700 4436 2702 4440
rect 2694 4435 2702 4436
rect 2694 4431 2696 4435
rect 2700 4431 2702 4435
rect 2694 4430 2702 4431
rect 2694 4426 2696 4430
rect 2700 4426 2702 4430
rect 2694 4425 2702 4426
rect 2694 4421 2696 4425
rect 2700 4421 2702 4425
rect 2694 4420 2702 4421
rect 2694 4416 2696 4420
rect 2700 4416 2702 4420
rect 2694 4415 2702 4416
rect 2694 4411 2696 4415
rect 2700 4411 2702 4415
rect 2694 4410 2702 4411
rect 2694 4406 2696 4410
rect 2700 4406 2702 4410
rect 2694 4405 2702 4406
rect 2694 4401 2696 4405
rect 2700 4401 2702 4405
rect 2694 4400 2702 4401
rect 2694 4396 2696 4400
rect 2700 4396 2702 4400
rect 2694 4395 2702 4396
rect 2694 4391 2696 4395
rect 2700 4391 2702 4395
rect 2694 4390 2702 4391
rect 2694 4386 2696 4390
rect 2700 4386 2702 4390
rect 2694 4385 2702 4386
rect 2694 4381 2696 4385
rect 2700 4381 2702 4385
rect 2694 4380 2702 4381
rect 2694 4376 2696 4380
rect 2700 4376 2702 4380
rect 2694 4375 2702 4376
rect 2694 4371 2696 4375
rect 2700 4371 2702 4375
rect 2694 4370 2702 4371
rect 2694 4366 2696 4370
rect 2700 4366 2702 4370
rect 2694 4365 2702 4366
rect 2694 4361 2696 4365
rect 2700 4361 2702 4365
rect 2630 4360 2638 4361
rect 2630 4356 2632 4360
rect 2636 4356 2638 4360
rect 2630 4355 2638 4356
rect 2694 4360 2702 4361
rect 2694 4356 2696 4360
rect 2700 4356 2702 4360
rect 2694 4355 2702 4356
rect 2630 4353 2702 4355
rect 2630 4349 2632 4353
rect 2636 4349 2639 4353
rect 2643 4349 2644 4353
rect 2648 4349 2649 4353
rect 2653 4349 2654 4353
rect 2658 4349 2659 4353
rect 2663 4349 2664 4353
rect 2668 4349 2669 4353
rect 2673 4349 2674 4353
rect 2678 4349 2679 4353
rect 2683 4349 2684 4353
rect 2688 4349 2689 4353
rect 2693 4349 2696 4353
rect 2700 4349 2702 4353
rect 2630 4347 2702 4349
rect 2778 4475 2874 4476
rect 2778 4471 2779 4475
rect 2783 4471 2784 4475
rect 2788 4471 2789 4475
rect 2793 4471 2794 4475
rect 2798 4471 2799 4475
rect 2803 4471 2804 4475
rect 2808 4471 2809 4475
rect 2813 4471 2814 4475
rect 2818 4471 2819 4475
rect 2823 4471 2824 4475
rect 2828 4471 2829 4475
rect 2833 4471 2834 4475
rect 2838 4471 2839 4475
rect 2843 4471 2844 4475
rect 2848 4471 2849 4475
rect 2853 4471 2854 4475
rect 2858 4471 2859 4475
rect 2863 4471 2864 4475
rect 2868 4471 2869 4475
rect 2873 4471 2874 4475
rect 2778 4470 2874 4471
rect 2778 4466 2779 4470
rect 2783 4466 2784 4470
rect 2778 4465 2784 4466
rect 2778 4461 2779 4465
rect 2783 4461 2784 4465
rect 2868 4466 2869 4470
rect 2873 4466 2874 4470
rect 2868 4465 2874 4466
rect 2778 4460 2784 4461
rect 2778 4456 2779 4460
rect 2783 4456 2784 4460
rect 2778 4455 2784 4456
rect 2778 4451 2779 4455
rect 2783 4451 2784 4455
rect 2778 4450 2784 4451
rect 2778 4446 2779 4450
rect 2783 4446 2784 4450
rect 2778 4445 2784 4446
rect 2778 4441 2779 4445
rect 2783 4441 2784 4445
rect 2778 4440 2784 4441
rect 2778 4436 2779 4440
rect 2783 4436 2784 4440
rect 2778 4435 2784 4436
rect 2778 4431 2779 4435
rect 2783 4431 2784 4435
rect 2778 4430 2784 4431
rect 2778 4426 2779 4430
rect 2783 4426 2784 4430
rect 2778 4425 2784 4426
rect 2778 4421 2779 4425
rect 2783 4421 2784 4425
rect 2778 4420 2784 4421
rect 2778 4416 2779 4420
rect 2783 4416 2784 4420
rect 2778 4415 2784 4416
rect 2778 4411 2779 4415
rect 2783 4411 2784 4415
rect 2778 4410 2784 4411
rect 2778 4406 2779 4410
rect 2783 4406 2784 4410
rect 2778 4405 2784 4406
rect 2778 4401 2779 4405
rect 2783 4401 2784 4405
rect 2778 4400 2784 4401
rect 2778 4396 2779 4400
rect 2783 4396 2784 4400
rect 2778 4395 2784 4396
rect 2778 4391 2779 4395
rect 2783 4391 2784 4395
rect 2778 4390 2784 4391
rect 2778 4386 2779 4390
rect 2783 4386 2784 4390
rect 2778 4385 2784 4386
rect 2778 4381 2779 4385
rect 2783 4381 2784 4385
rect 2778 4380 2784 4381
rect 2778 4376 2779 4380
rect 2783 4376 2784 4380
rect 2778 4375 2784 4376
rect 2778 4371 2779 4375
rect 2783 4371 2784 4375
rect 2778 4370 2784 4371
rect 2778 4366 2779 4370
rect 2783 4366 2784 4370
rect 2778 4365 2784 4366
rect 2778 4361 2779 4365
rect 2783 4361 2784 4365
rect 2778 4360 2784 4361
rect 2778 4356 2779 4360
rect 2783 4356 2784 4360
rect 2778 4355 2784 4356
rect 2778 4351 2779 4355
rect 2783 4351 2784 4355
rect 2778 4350 2784 4351
rect 2778 4346 2779 4350
rect 2783 4346 2784 4350
rect 2868 4461 2869 4465
rect 2873 4461 2874 4465
rect 2868 4460 2874 4461
rect 2868 4456 2869 4460
rect 2873 4456 2874 4460
rect 2868 4455 2874 4456
rect 2868 4451 2869 4455
rect 2873 4451 2874 4455
rect 2868 4450 2874 4451
rect 2868 4446 2869 4450
rect 2873 4446 2874 4450
rect 2868 4445 2874 4446
rect 2868 4441 2869 4445
rect 2873 4441 2874 4445
rect 2868 4440 2874 4441
rect 2868 4436 2869 4440
rect 2873 4436 2874 4440
rect 2868 4435 2874 4436
rect 2868 4431 2869 4435
rect 2873 4431 2874 4435
rect 2868 4430 2874 4431
rect 2868 4426 2869 4430
rect 2873 4426 2874 4430
rect 2868 4425 2874 4426
rect 2868 4421 2869 4425
rect 2873 4421 2874 4425
rect 2868 4420 2874 4421
rect 2868 4416 2869 4420
rect 2873 4416 2874 4420
rect 2868 4415 2874 4416
rect 2868 4411 2869 4415
rect 2873 4411 2874 4415
rect 2868 4410 2874 4411
rect 2868 4406 2869 4410
rect 2873 4406 2874 4410
rect 2868 4405 2874 4406
rect 2868 4401 2869 4405
rect 2873 4401 2874 4405
rect 2868 4400 2874 4401
rect 2868 4396 2869 4400
rect 2873 4396 2874 4400
rect 2868 4395 2874 4396
rect 2868 4391 2869 4395
rect 2873 4391 2874 4395
rect 2868 4390 2874 4391
rect 2868 4386 2869 4390
rect 2873 4386 2874 4390
rect 2868 4385 2874 4386
rect 2868 4381 2869 4385
rect 2873 4381 2874 4385
rect 2868 4380 2874 4381
rect 2868 4376 2869 4380
rect 2873 4376 2874 4380
rect 2868 4375 2874 4376
rect 2868 4371 2869 4375
rect 2873 4371 2874 4375
rect 2868 4370 2874 4371
rect 2868 4366 2869 4370
rect 2873 4366 2874 4370
rect 2868 4365 2874 4366
rect 2868 4361 2869 4365
rect 2873 4361 2874 4365
rect 2868 4360 2874 4361
rect 2868 4356 2869 4360
rect 2873 4356 2874 4360
rect 2868 4355 2874 4356
rect 2868 4351 2869 4355
rect 2873 4351 2874 4355
rect 2868 4350 2874 4351
rect 2778 4345 2784 4346
rect 2778 4341 2779 4345
rect 2783 4341 2784 4345
rect 2868 4346 2869 4350
rect 2873 4346 2874 4350
rect 2868 4345 2874 4346
rect 2868 4341 2869 4345
rect 2873 4341 2874 4345
rect 2778 4340 2874 4341
rect 2778 4336 2779 4340
rect 2783 4336 2784 4340
rect 2788 4336 2789 4340
rect 2793 4336 2794 4340
rect 2798 4336 2799 4340
rect 2803 4336 2804 4340
rect 2808 4336 2809 4340
rect 2813 4336 2814 4340
rect 2818 4336 2819 4340
rect 2823 4336 2824 4340
rect 2828 4336 2829 4340
rect 2833 4336 2834 4340
rect 2838 4336 2839 4340
rect 2843 4336 2844 4340
rect 2848 4336 2849 4340
rect 2853 4336 2854 4340
rect 2858 4336 2859 4340
rect 2863 4336 2864 4340
rect 2868 4336 2869 4340
rect 2873 4336 2874 4340
rect 2778 4335 2874 4336
rect 2939 4462 3011 4464
rect 2939 4458 2941 4462
rect 2945 4458 2948 4462
rect 2952 4458 2953 4462
rect 2957 4458 2958 4462
rect 2962 4458 2963 4462
rect 2967 4458 2968 4462
rect 2972 4458 2973 4462
rect 2977 4458 2978 4462
rect 2982 4458 2983 4462
rect 2987 4458 2988 4462
rect 2992 4458 2993 4462
rect 2997 4458 2998 4462
rect 3002 4458 3005 4462
rect 3009 4458 3011 4462
rect 2939 4456 3011 4458
rect 2939 4455 2947 4456
rect 2939 4451 2941 4455
rect 2945 4451 2947 4455
rect 2939 4450 2947 4451
rect 3003 4455 3011 4456
rect 3003 4451 3005 4455
rect 3009 4451 3011 4455
rect 3003 4450 3011 4451
rect 2939 4446 2941 4450
rect 2945 4446 2947 4450
rect 2939 4445 2947 4446
rect 2939 4441 2941 4445
rect 2945 4441 2947 4445
rect 2939 4440 2947 4441
rect 2939 4436 2941 4440
rect 2945 4436 2947 4440
rect 2939 4435 2947 4436
rect 2939 4431 2941 4435
rect 2945 4431 2947 4435
rect 2939 4430 2947 4431
rect 2939 4426 2941 4430
rect 2945 4426 2947 4430
rect 2939 4425 2947 4426
rect 2939 4421 2941 4425
rect 2945 4421 2947 4425
rect 2939 4420 2947 4421
rect 2939 4416 2941 4420
rect 2945 4416 2947 4420
rect 2939 4415 2947 4416
rect 2939 4411 2941 4415
rect 2945 4411 2947 4415
rect 2939 4410 2947 4411
rect 2939 4406 2941 4410
rect 2945 4406 2947 4410
rect 2939 4405 2947 4406
rect 2939 4401 2941 4405
rect 2945 4401 2947 4405
rect 2939 4400 2947 4401
rect 2939 4396 2941 4400
rect 2945 4396 2947 4400
rect 2939 4395 2947 4396
rect 2939 4391 2941 4395
rect 2945 4391 2947 4395
rect 2939 4390 2947 4391
rect 2939 4386 2941 4390
rect 2945 4386 2947 4390
rect 2939 4385 2947 4386
rect 2939 4381 2941 4385
rect 2945 4381 2947 4385
rect 2939 4380 2947 4381
rect 2939 4376 2941 4380
rect 2945 4376 2947 4380
rect 2939 4375 2947 4376
rect 2939 4371 2941 4375
rect 2945 4371 2947 4375
rect 2939 4370 2947 4371
rect 2939 4366 2941 4370
rect 2945 4366 2947 4370
rect 2939 4365 2947 4366
rect 2939 4361 2941 4365
rect 2945 4361 2947 4365
rect 3003 4446 3005 4450
rect 3009 4446 3011 4450
rect 3003 4445 3011 4446
rect 3003 4441 3005 4445
rect 3009 4441 3011 4445
rect 3003 4440 3011 4441
rect 3003 4436 3005 4440
rect 3009 4436 3011 4440
rect 3003 4435 3011 4436
rect 3003 4431 3005 4435
rect 3009 4431 3011 4435
rect 3003 4430 3011 4431
rect 3003 4426 3005 4430
rect 3009 4426 3011 4430
rect 3003 4425 3011 4426
rect 3003 4421 3005 4425
rect 3009 4421 3011 4425
rect 3003 4420 3011 4421
rect 3003 4416 3005 4420
rect 3009 4416 3011 4420
rect 3003 4415 3011 4416
rect 3003 4411 3005 4415
rect 3009 4411 3011 4415
rect 3003 4410 3011 4411
rect 3003 4406 3005 4410
rect 3009 4406 3011 4410
rect 3003 4405 3011 4406
rect 3003 4401 3005 4405
rect 3009 4401 3011 4405
rect 3003 4400 3011 4401
rect 3003 4396 3005 4400
rect 3009 4396 3011 4400
rect 3003 4395 3011 4396
rect 3003 4391 3005 4395
rect 3009 4391 3011 4395
rect 3003 4390 3011 4391
rect 3003 4386 3005 4390
rect 3009 4386 3011 4390
rect 3003 4385 3011 4386
rect 3003 4381 3005 4385
rect 3009 4381 3011 4385
rect 3003 4380 3011 4381
rect 3003 4376 3005 4380
rect 3009 4376 3011 4380
rect 3003 4375 3011 4376
rect 3003 4371 3005 4375
rect 3009 4371 3011 4375
rect 3003 4370 3011 4371
rect 3003 4366 3005 4370
rect 3009 4366 3011 4370
rect 3003 4365 3011 4366
rect 3003 4361 3005 4365
rect 3009 4361 3011 4365
rect 2939 4360 2947 4361
rect 2939 4356 2941 4360
rect 2945 4356 2947 4360
rect 2939 4355 2947 4356
rect 3003 4360 3011 4361
rect 3003 4356 3005 4360
rect 3009 4356 3011 4360
rect 3003 4355 3011 4356
rect 2939 4353 3011 4355
rect 2939 4349 2941 4353
rect 2945 4349 2948 4353
rect 2952 4349 2953 4353
rect 2957 4349 2958 4353
rect 2962 4349 2963 4353
rect 2967 4349 2968 4353
rect 2972 4349 2973 4353
rect 2977 4349 2978 4353
rect 2982 4349 2983 4353
rect 2987 4349 2988 4353
rect 2992 4349 2993 4353
rect 2997 4349 2998 4353
rect 3002 4349 3005 4353
rect 3009 4349 3011 4353
rect 2939 4347 3011 4349
rect 3087 4475 3183 4476
rect 3087 4471 3088 4475
rect 3092 4471 3093 4475
rect 3097 4471 3098 4475
rect 3102 4471 3103 4475
rect 3107 4471 3108 4475
rect 3112 4471 3113 4475
rect 3117 4471 3118 4475
rect 3122 4471 3123 4475
rect 3127 4471 3128 4475
rect 3132 4471 3133 4475
rect 3137 4471 3138 4475
rect 3142 4471 3143 4475
rect 3147 4471 3148 4475
rect 3152 4471 3153 4475
rect 3157 4471 3158 4475
rect 3162 4471 3163 4475
rect 3167 4471 3168 4475
rect 3172 4471 3173 4475
rect 3177 4471 3178 4475
rect 3182 4471 3183 4475
rect 3087 4470 3183 4471
rect 3087 4466 3088 4470
rect 3092 4466 3093 4470
rect 3087 4465 3093 4466
rect 3087 4461 3088 4465
rect 3092 4461 3093 4465
rect 3177 4466 3178 4470
rect 3182 4466 3183 4470
rect 3177 4465 3183 4466
rect 3087 4460 3093 4461
rect 3087 4456 3088 4460
rect 3092 4456 3093 4460
rect 3087 4455 3093 4456
rect 3087 4451 3088 4455
rect 3092 4451 3093 4455
rect 3087 4450 3093 4451
rect 3087 4446 3088 4450
rect 3092 4446 3093 4450
rect 3087 4445 3093 4446
rect 3087 4441 3088 4445
rect 3092 4441 3093 4445
rect 3087 4440 3093 4441
rect 3087 4436 3088 4440
rect 3092 4436 3093 4440
rect 3087 4435 3093 4436
rect 3087 4431 3088 4435
rect 3092 4431 3093 4435
rect 3087 4430 3093 4431
rect 3087 4426 3088 4430
rect 3092 4426 3093 4430
rect 3087 4425 3093 4426
rect 3087 4421 3088 4425
rect 3092 4421 3093 4425
rect 3087 4420 3093 4421
rect 3087 4416 3088 4420
rect 3092 4416 3093 4420
rect 3087 4415 3093 4416
rect 3087 4411 3088 4415
rect 3092 4411 3093 4415
rect 3087 4410 3093 4411
rect 3087 4406 3088 4410
rect 3092 4406 3093 4410
rect 3087 4405 3093 4406
rect 3087 4401 3088 4405
rect 3092 4401 3093 4405
rect 3087 4400 3093 4401
rect 3087 4396 3088 4400
rect 3092 4396 3093 4400
rect 3087 4395 3093 4396
rect 3087 4391 3088 4395
rect 3092 4391 3093 4395
rect 3087 4390 3093 4391
rect 3087 4386 3088 4390
rect 3092 4386 3093 4390
rect 3087 4385 3093 4386
rect 3087 4381 3088 4385
rect 3092 4381 3093 4385
rect 3087 4380 3093 4381
rect 3087 4376 3088 4380
rect 3092 4376 3093 4380
rect 3087 4375 3093 4376
rect 3087 4371 3088 4375
rect 3092 4371 3093 4375
rect 3087 4370 3093 4371
rect 3087 4366 3088 4370
rect 3092 4366 3093 4370
rect 3087 4365 3093 4366
rect 3087 4361 3088 4365
rect 3092 4361 3093 4365
rect 3087 4360 3093 4361
rect 3087 4356 3088 4360
rect 3092 4356 3093 4360
rect 3087 4355 3093 4356
rect 3087 4351 3088 4355
rect 3092 4351 3093 4355
rect 3087 4350 3093 4351
rect 3087 4346 3088 4350
rect 3092 4346 3093 4350
rect 3177 4461 3178 4465
rect 3182 4461 3183 4465
rect 3177 4460 3183 4461
rect 3177 4456 3178 4460
rect 3182 4456 3183 4460
rect 3177 4455 3183 4456
rect 3177 4451 3178 4455
rect 3182 4451 3183 4455
rect 3177 4450 3183 4451
rect 3177 4446 3178 4450
rect 3182 4446 3183 4450
rect 3177 4445 3183 4446
rect 3177 4441 3178 4445
rect 3182 4441 3183 4445
rect 3177 4440 3183 4441
rect 3177 4436 3178 4440
rect 3182 4436 3183 4440
rect 3177 4435 3183 4436
rect 3177 4431 3178 4435
rect 3182 4431 3183 4435
rect 3177 4430 3183 4431
rect 3177 4426 3178 4430
rect 3182 4426 3183 4430
rect 3177 4425 3183 4426
rect 3177 4421 3178 4425
rect 3182 4421 3183 4425
rect 3177 4420 3183 4421
rect 3177 4416 3178 4420
rect 3182 4416 3183 4420
rect 3177 4415 3183 4416
rect 3177 4411 3178 4415
rect 3182 4411 3183 4415
rect 3177 4410 3183 4411
rect 3177 4406 3178 4410
rect 3182 4406 3183 4410
rect 3177 4405 3183 4406
rect 3177 4401 3178 4405
rect 3182 4401 3183 4405
rect 3177 4400 3183 4401
rect 3177 4396 3178 4400
rect 3182 4396 3183 4400
rect 3177 4395 3183 4396
rect 3177 4391 3178 4395
rect 3182 4391 3183 4395
rect 3177 4390 3183 4391
rect 3177 4386 3178 4390
rect 3182 4386 3183 4390
rect 3177 4385 3183 4386
rect 3177 4381 3178 4385
rect 3182 4381 3183 4385
rect 3177 4380 3183 4381
rect 3177 4376 3178 4380
rect 3182 4376 3183 4380
rect 3177 4375 3183 4376
rect 3177 4371 3178 4375
rect 3182 4371 3183 4375
rect 3177 4370 3183 4371
rect 3177 4366 3178 4370
rect 3182 4366 3183 4370
rect 3177 4365 3183 4366
rect 3177 4361 3178 4365
rect 3182 4361 3183 4365
rect 3177 4360 3183 4361
rect 3177 4356 3178 4360
rect 3182 4356 3183 4360
rect 3177 4355 3183 4356
rect 3177 4351 3178 4355
rect 3182 4351 3183 4355
rect 3177 4350 3183 4351
rect 3087 4345 3093 4346
rect 3087 4341 3088 4345
rect 3092 4341 3093 4345
rect 3177 4346 3178 4350
rect 3182 4346 3183 4350
rect 3177 4345 3183 4346
rect 3177 4341 3178 4345
rect 3182 4341 3183 4345
rect 3087 4340 3183 4341
rect 3087 4336 3088 4340
rect 3092 4336 3093 4340
rect 3097 4336 3098 4340
rect 3102 4336 3103 4340
rect 3107 4336 3108 4340
rect 3112 4336 3113 4340
rect 3117 4336 3118 4340
rect 3122 4336 3123 4340
rect 3127 4336 3128 4340
rect 3132 4336 3133 4340
rect 3137 4336 3138 4340
rect 3142 4336 3143 4340
rect 3147 4336 3148 4340
rect 3152 4336 3153 4340
rect 3157 4336 3158 4340
rect 3162 4336 3163 4340
rect 3167 4336 3168 4340
rect 3172 4336 3173 4340
rect 3177 4336 3178 4340
rect 3182 4336 3183 4340
rect 3087 4335 3183 4336
rect 3248 4462 3320 4464
rect 3248 4458 3250 4462
rect 3254 4458 3257 4462
rect 3261 4458 3262 4462
rect 3266 4458 3267 4462
rect 3271 4458 3272 4462
rect 3276 4458 3277 4462
rect 3281 4458 3282 4462
rect 3286 4458 3287 4462
rect 3291 4458 3292 4462
rect 3296 4458 3297 4462
rect 3301 4458 3302 4462
rect 3306 4458 3307 4462
rect 3311 4458 3314 4462
rect 3318 4458 3320 4462
rect 3248 4456 3320 4458
rect 3248 4455 3256 4456
rect 3248 4451 3250 4455
rect 3254 4451 3256 4455
rect 3248 4450 3256 4451
rect 3312 4455 3320 4456
rect 3312 4451 3314 4455
rect 3318 4451 3320 4455
rect 3312 4450 3320 4451
rect 3248 4446 3250 4450
rect 3254 4446 3256 4450
rect 3248 4445 3256 4446
rect 3248 4441 3250 4445
rect 3254 4441 3256 4445
rect 3248 4440 3256 4441
rect 3248 4436 3250 4440
rect 3254 4436 3256 4440
rect 3248 4435 3256 4436
rect 3248 4431 3250 4435
rect 3254 4431 3256 4435
rect 3248 4430 3256 4431
rect 3248 4426 3250 4430
rect 3254 4426 3256 4430
rect 3248 4425 3256 4426
rect 3248 4421 3250 4425
rect 3254 4421 3256 4425
rect 3248 4420 3256 4421
rect 3248 4416 3250 4420
rect 3254 4416 3256 4420
rect 3248 4415 3256 4416
rect 3248 4411 3250 4415
rect 3254 4411 3256 4415
rect 3248 4410 3256 4411
rect 3248 4406 3250 4410
rect 3254 4406 3256 4410
rect 3248 4405 3256 4406
rect 3248 4401 3250 4405
rect 3254 4401 3256 4405
rect 3248 4400 3256 4401
rect 3248 4396 3250 4400
rect 3254 4396 3256 4400
rect 3248 4395 3256 4396
rect 3248 4391 3250 4395
rect 3254 4391 3256 4395
rect 3248 4390 3256 4391
rect 3248 4386 3250 4390
rect 3254 4386 3256 4390
rect 3248 4385 3256 4386
rect 3248 4381 3250 4385
rect 3254 4381 3256 4385
rect 3248 4380 3256 4381
rect 3248 4376 3250 4380
rect 3254 4376 3256 4380
rect 3248 4375 3256 4376
rect 3248 4371 3250 4375
rect 3254 4371 3256 4375
rect 3248 4370 3256 4371
rect 3248 4366 3250 4370
rect 3254 4366 3256 4370
rect 3248 4365 3256 4366
rect 3248 4361 3250 4365
rect 3254 4361 3256 4365
rect 3312 4446 3314 4450
rect 3318 4446 3320 4450
rect 3312 4445 3320 4446
rect 3312 4441 3314 4445
rect 3318 4441 3320 4445
rect 3312 4440 3320 4441
rect 3312 4436 3314 4440
rect 3318 4436 3320 4440
rect 3312 4435 3320 4436
rect 3312 4431 3314 4435
rect 3318 4431 3320 4435
rect 3312 4430 3320 4431
rect 3312 4426 3314 4430
rect 3318 4426 3320 4430
rect 3312 4425 3320 4426
rect 3312 4421 3314 4425
rect 3318 4421 3320 4425
rect 3312 4420 3320 4421
rect 3312 4416 3314 4420
rect 3318 4416 3320 4420
rect 3312 4415 3320 4416
rect 3312 4411 3314 4415
rect 3318 4411 3320 4415
rect 3312 4410 3320 4411
rect 3312 4406 3314 4410
rect 3318 4406 3320 4410
rect 3312 4405 3320 4406
rect 3312 4401 3314 4405
rect 3318 4401 3320 4405
rect 3312 4400 3320 4401
rect 3312 4396 3314 4400
rect 3318 4396 3320 4400
rect 3312 4395 3320 4396
rect 3312 4391 3314 4395
rect 3318 4391 3320 4395
rect 3312 4390 3320 4391
rect 3312 4386 3314 4390
rect 3318 4386 3320 4390
rect 3312 4385 3320 4386
rect 3312 4381 3314 4385
rect 3318 4381 3320 4385
rect 3312 4380 3320 4381
rect 3312 4376 3314 4380
rect 3318 4376 3320 4380
rect 3312 4375 3320 4376
rect 3312 4371 3314 4375
rect 3318 4371 3320 4375
rect 3312 4370 3320 4371
rect 3312 4366 3314 4370
rect 3318 4366 3320 4370
rect 3312 4365 3320 4366
rect 3312 4361 3314 4365
rect 3318 4361 3320 4365
rect 3248 4360 3256 4361
rect 3248 4356 3250 4360
rect 3254 4356 3256 4360
rect 3248 4355 3256 4356
rect 3312 4360 3320 4361
rect 3312 4356 3314 4360
rect 3318 4356 3320 4360
rect 3312 4355 3320 4356
rect 3248 4353 3320 4355
rect 3248 4349 3250 4353
rect 3254 4349 3257 4353
rect 3261 4349 3262 4353
rect 3266 4349 3267 4353
rect 3271 4349 3272 4353
rect 3276 4349 3277 4353
rect 3281 4349 3282 4353
rect 3286 4349 3287 4353
rect 3291 4349 3292 4353
rect 3296 4349 3297 4353
rect 3301 4349 3302 4353
rect 3306 4349 3307 4353
rect 3311 4349 3314 4353
rect 3318 4349 3320 4353
rect 3248 4347 3320 4349
rect 3396 4475 3492 4476
rect 3396 4471 3397 4475
rect 3401 4471 3402 4475
rect 3406 4471 3407 4475
rect 3411 4471 3412 4475
rect 3416 4471 3417 4475
rect 3421 4471 3422 4475
rect 3426 4471 3427 4475
rect 3431 4471 3432 4475
rect 3436 4471 3437 4475
rect 3441 4471 3442 4475
rect 3446 4471 3447 4475
rect 3451 4471 3452 4475
rect 3456 4471 3457 4475
rect 3461 4471 3462 4475
rect 3466 4471 3467 4475
rect 3471 4471 3472 4475
rect 3476 4471 3477 4475
rect 3481 4471 3482 4475
rect 3486 4471 3487 4475
rect 3491 4471 3492 4475
rect 3396 4470 3492 4471
rect 3396 4466 3397 4470
rect 3401 4466 3402 4470
rect 3396 4465 3402 4466
rect 3396 4461 3397 4465
rect 3401 4461 3402 4465
rect 3486 4466 3487 4470
rect 3491 4466 3492 4470
rect 3486 4465 3492 4466
rect 3396 4460 3402 4461
rect 3396 4456 3397 4460
rect 3401 4456 3402 4460
rect 3396 4455 3402 4456
rect 3396 4451 3397 4455
rect 3401 4451 3402 4455
rect 3396 4450 3402 4451
rect 3396 4446 3397 4450
rect 3401 4446 3402 4450
rect 3396 4445 3402 4446
rect 3396 4441 3397 4445
rect 3401 4441 3402 4445
rect 3396 4440 3402 4441
rect 3396 4436 3397 4440
rect 3401 4436 3402 4440
rect 3396 4435 3402 4436
rect 3396 4431 3397 4435
rect 3401 4431 3402 4435
rect 3396 4430 3402 4431
rect 3396 4426 3397 4430
rect 3401 4426 3402 4430
rect 3396 4425 3402 4426
rect 3396 4421 3397 4425
rect 3401 4421 3402 4425
rect 3396 4420 3402 4421
rect 3396 4416 3397 4420
rect 3401 4416 3402 4420
rect 3396 4415 3402 4416
rect 3396 4411 3397 4415
rect 3401 4411 3402 4415
rect 3396 4410 3402 4411
rect 3396 4406 3397 4410
rect 3401 4406 3402 4410
rect 3396 4405 3402 4406
rect 3396 4401 3397 4405
rect 3401 4401 3402 4405
rect 3396 4400 3402 4401
rect 3396 4396 3397 4400
rect 3401 4396 3402 4400
rect 3396 4395 3402 4396
rect 3396 4391 3397 4395
rect 3401 4391 3402 4395
rect 3396 4390 3402 4391
rect 3396 4386 3397 4390
rect 3401 4386 3402 4390
rect 3396 4385 3402 4386
rect 3396 4381 3397 4385
rect 3401 4381 3402 4385
rect 3396 4380 3402 4381
rect 3396 4376 3397 4380
rect 3401 4376 3402 4380
rect 3396 4375 3402 4376
rect 3396 4371 3397 4375
rect 3401 4371 3402 4375
rect 3396 4370 3402 4371
rect 3396 4366 3397 4370
rect 3401 4366 3402 4370
rect 3396 4365 3402 4366
rect 3396 4361 3397 4365
rect 3401 4361 3402 4365
rect 3396 4360 3402 4361
rect 3396 4356 3397 4360
rect 3401 4356 3402 4360
rect 3396 4355 3402 4356
rect 3396 4351 3397 4355
rect 3401 4351 3402 4355
rect 3396 4350 3402 4351
rect 3396 4346 3397 4350
rect 3401 4346 3402 4350
rect 3486 4461 3487 4465
rect 3491 4461 3492 4465
rect 3486 4460 3492 4461
rect 3486 4456 3487 4460
rect 3491 4456 3492 4460
rect 3486 4455 3492 4456
rect 3486 4451 3487 4455
rect 3491 4451 3492 4455
rect 3486 4450 3492 4451
rect 3486 4446 3487 4450
rect 3491 4446 3492 4450
rect 3486 4445 3492 4446
rect 3486 4441 3487 4445
rect 3491 4441 3492 4445
rect 3486 4440 3492 4441
rect 3486 4436 3487 4440
rect 3491 4436 3492 4440
rect 3486 4435 3492 4436
rect 3486 4431 3487 4435
rect 3491 4431 3492 4435
rect 3486 4430 3492 4431
rect 3486 4426 3487 4430
rect 3491 4426 3492 4430
rect 3486 4425 3492 4426
rect 3486 4421 3487 4425
rect 3491 4421 3492 4425
rect 3486 4420 3492 4421
rect 3486 4416 3487 4420
rect 3491 4416 3492 4420
rect 3486 4415 3492 4416
rect 3486 4411 3487 4415
rect 3491 4411 3492 4415
rect 3486 4410 3492 4411
rect 3486 4406 3487 4410
rect 3491 4406 3492 4410
rect 3486 4405 3492 4406
rect 3486 4401 3487 4405
rect 3491 4401 3492 4405
rect 3486 4400 3492 4401
rect 3486 4396 3487 4400
rect 3491 4396 3492 4400
rect 3486 4395 3492 4396
rect 3486 4391 3487 4395
rect 3491 4391 3492 4395
rect 3486 4390 3492 4391
rect 3486 4386 3487 4390
rect 3491 4386 3492 4390
rect 3486 4385 3492 4386
rect 3486 4381 3487 4385
rect 3491 4381 3492 4385
rect 3486 4380 3492 4381
rect 3486 4376 3487 4380
rect 3491 4376 3492 4380
rect 3486 4375 3492 4376
rect 3486 4371 3487 4375
rect 3491 4371 3492 4375
rect 3486 4370 3492 4371
rect 3486 4366 3487 4370
rect 3491 4366 3492 4370
rect 3486 4365 3492 4366
rect 3486 4361 3487 4365
rect 3491 4361 3492 4365
rect 3486 4360 3492 4361
rect 3486 4356 3487 4360
rect 3491 4356 3492 4360
rect 3486 4355 3492 4356
rect 3486 4351 3487 4355
rect 3491 4351 3492 4355
rect 3486 4350 3492 4351
rect 3396 4345 3402 4346
rect 3396 4341 3397 4345
rect 3401 4341 3402 4345
rect 3486 4346 3487 4350
rect 3491 4346 3492 4350
rect 3486 4345 3492 4346
rect 3486 4341 3487 4345
rect 3491 4341 3492 4345
rect 3396 4340 3492 4341
rect 3396 4336 3397 4340
rect 3401 4336 3402 4340
rect 3406 4336 3407 4340
rect 3411 4336 3412 4340
rect 3416 4336 3417 4340
rect 3421 4336 3422 4340
rect 3426 4336 3427 4340
rect 3431 4336 3432 4340
rect 3436 4336 3437 4340
rect 3441 4336 3442 4340
rect 3446 4336 3447 4340
rect 3451 4336 3452 4340
rect 3456 4336 3457 4340
rect 3461 4336 3462 4340
rect 3466 4336 3467 4340
rect 3471 4336 3472 4340
rect 3476 4336 3477 4340
rect 3481 4336 3482 4340
rect 3486 4336 3487 4340
rect 3491 4336 3492 4340
rect 3396 4335 3492 4336
rect 3557 4462 3629 4464
rect 3557 4458 3559 4462
rect 3563 4458 3566 4462
rect 3570 4458 3571 4462
rect 3575 4458 3576 4462
rect 3580 4458 3581 4462
rect 3585 4458 3586 4462
rect 3590 4458 3591 4462
rect 3595 4458 3596 4462
rect 3600 4458 3601 4462
rect 3605 4458 3606 4462
rect 3610 4458 3611 4462
rect 3615 4458 3616 4462
rect 3620 4458 3623 4462
rect 3627 4458 3629 4462
rect 3557 4456 3629 4458
rect 3557 4455 3565 4456
rect 3557 4451 3559 4455
rect 3563 4451 3565 4455
rect 3557 4450 3565 4451
rect 3621 4455 3629 4456
rect 3621 4451 3623 4455
rect 3627 4451 3629 4455
rect 3621 4450 3629 4451
rect 3557 4446 3559 4450
rect 3563 4446 3565 4450
rect 3557 4445 3565 4446
rect 3557 4441 3559 4445
rect 3563 4441 3565 4445
rect 3557 4440 3565 4441
rect 3557 4436 3559 4440
rect 3563 4436 3565 4440
rect 3557 4435 3565 4436
rect 3557 4431 3559 4435
rect 3563 4431 3565 4435
rect 3557 4430 3565 4431
rect 3557 4426 3559 4430
rect 3563 4426 3565 4430
rect 3557 4425 3565 4426
rect 3557 4421 3559 4425
rect 3563 4421 3565 4425
rect 3557 4420 3565 4421
rect 3557 4416 3559 4420
rect 3563 4416 3565 4420
rect 3557 4415 3565 4416
rect 3557 4411 3559 4415
rect 3563 4411 3565 4415
rect 3557 4410 3565 4411
rect 3557 4406 3559 4410
rect 3563 4406 3565 4410
rect 3557 4405 3565 4406
rect 3557 4401 3559 4405
rect 3563 4401 3565 4405
rect 3557 4400 3565 4401
rect 3557 4396 3559 4400
rect 3563 4396 3565 4400
rect 3557 4395 3565 4396
rect 3557 4391 3559 4395
rect 3563 4391 3565 4395
rect 3557 4390 3565 4391
rect 3557 4386 3559 4390
rect 3563 4386 3565 4390
rect 3557 4385 3565 4386
rect 3557 4381 3559 4385
rect 3563 4381 3565 4385
rect 3557 4380 3565 4381
rect 3557 4376 3559 4380
rect 3563 4376 3565 4380
rect 3557 4375 3565 4376
rect 3557 4371 3559 4375
rect 3563 4371 3565 4375
rect 3557 4370 3565 4371
rect 3557 4366 3559 4370
rect 3563 4366 3565 4370
rect 3557 4365 3565 4366
rect 3557 4361 3559 4365
rect 3563 4361 3565 4365
rect 3621 4446 3623 4450
rect 3627 4446 3629 4450
rect 3621 4445 3629 4446
rect 3621 4441 3623 4445
rect 3627 4441 3629 4445
rect 3621 4440 3629 4441
rect 3621 4436 3623 4440
rect 3627 4436 3629 4440
rect 3621 4435 3629 4436
rect 3621 4431 3623 4435
rect 3627 4431 3629 4435
rect 3621 4430 3629 4431
rect 3621 4426 3623 4430
rect 3627 4426 3629 4430
rect 3621 4425 3629 4426
rect 3621 4421 3623 4425
rect 3627 4421 3629 4425
rect 3621 4420 3629 4421
rect 3621 4416 3623 4420
rect 3627 4416 3629 4420
rect 3621 4415 3629 4416
rect 3621 4411 3623 4415
rect 3627 4411 3629 4415
rect 3621 4410 3629 4411
rect 3621 4406 3623 4410
rect 3627 4406 3629 4410
rect 3621 4405 3629 4406
rect 3621 4401 3623 4405
rect 3627 4401 3629 4405
rect 3621 4400 3629 4401
rect 3621 4396 3623 4400
rect 3627 4396 3629 4400
rect 3621 4395 3629 4396
rect 3621 4391 3623 4395
rect 3627 4391 3629 4395
rect 3621 4390 3629 4391
rect 3621 4386 3623 4390
rect 3627 4386 3629 4390
rect 3621 4385 3629 4386
rect 3621 4381 3623 4385
rect 3627 4381 3629 4385
rect 3621 4380 3629 4381
rect 3621 4376 3623 4380
rect 3627 4376 3629 4380
rect 3621 4375 3629 4376
rect 3621 4371 3623 4375
rect 3627 4371 3629 4375
rect 3621 4370 3629 4371
rect 3621 4366 3623 4370
rect 3627 4366 3629 4370
rect 3621 4365 3629 4366
rect 3621 4361 3623 4365
rect 3627 4361 3629 4365
rect 3557 4360 3565 4361
rect 3557 4356 3559 4360
rect 3563 4356 3565 4360
rect 3557 4355 3565 4356
rect 3621 4360 3629 4361
rect 3621 4356 3623 4360
rect 3627 4356 3629 4360
rect 3621 4355 3629 4356
rect 3557 4353 3629 4355
rect 3557 4349 3559 4353
rect 3563 4349 3566 4353
rect 3570 4349 3571 4353
rect 3575 4349 3576 4353
rect 3580 4349 3581 4353
rect 3585 4349 3586 4353
rect 3590 4349 3591 4353
rect 3595 4349 3596 4353
rect 3600 4349 3601 4353
rect 3605 4349 3606 4353
rect 3610 4349 3611 4353
rect 3615 4349 3616 4353
rect 3620 4349 3623 4353
rect 3627 4349 3629 4353
rect 3557 4347 3629 4349
rect 3705 4475 3801 4476
rect 3705 4471 3706 4475
rect 3710 4471 3711 4475
rect 3715 4471 3716 4475
rect 3720 4471 3721 4475
rect 3725 4471 3726 4475
rect 3730 4471 3731 4475
rect 3735 4471 3736 4475
rect 3740 4471 3741 4475
rect 3745 4471 3746 4475
rect 3750 4471 3751 4475
rect 3755 4471 3756 4475
rect 3760 4471 3761 4475
rect 3765 4471 3766 4475
rect 3770 4471 3771 4475
rect 3775 4471 3776 4475
rect 3780 4471 3781 4475
rect 3785 4471 3786 4475
rect 3790 4471 3791 4475
rect 3795 4471 3796 4475
rect 3800 4471 3801 4475
rect 3705 4470 3801 4471
rect 3705 4466 3706 4470
rect 3710 4466 3711 4470
rect 3705 4465 3711 4466
rect 3705 4461 3706 4465
rect 3710 4461 3711 4465
rect 3795 4466 3796 4470
rect 3800 4466 3801 4470
rect 3795 4465 3801 4466
rect 3705 4460 3711 4461
rect 3705 4456 3706 4460
rect 3710 4456 3711 4460
rect 3705 4455 3711 4456
rect 3705 4451 3706 4455
rect 3710 4451 3711 4455
rect 3705 4450 3711 4451
rect 3705 4446 3706 4450
rect 3710 4446 3711 4450
rect 3705 4445 3711 4446
rect 3705 4441 3706 4445
rect 3710 4441 3711 4445
rect 3705 4440 3711 4441
rect 3705 4436 3706 4440
rect 3710 4436 3711 4440
rect 3705 4435 3711 4436
rect 3705 4431 3706 4435
rect 3710 4431 3711 4435
rect 3705 4430 3711 4431
rect 3705 4426 3706 4430
rect 3710 4426 3711 4430
rect 3705 4425 3711 4426
rect 3705 4421 3706 4425
rect 3710 4421 3711 4425
rect 3705 4420 3711 4421
rect 3705 4416 3706 4420
rect 3710 4416 3711 4420
rect 3705 4415 3711 4416
rect 3705 4411 3706 4415
rect 3710 4411 3711 4415
rect 3705 4410 3711 4411
rect 3705 4406 3706 4410
rect 3710 4406 3711 4410
rect 3705 4405 3711 4406
rect 3705 4401 3706 4405
rect 3710 4401 3711 4405
rect 3705 4400 3711 4401
rect 3705 4396 3706 4400
rect 3710 4396 3711 4400
rect 3705 4395 3711 4396
rect 3705 4391 3706 4395
rect 3710 4391 3711 4395
rect 3705 4390 3711 4391
rect 3705 4386 3706 4390
rect 3710 4386 3711 4390
rect 3705 4385 3711 4386
rect 3705 4381 3706 4385
rect 3710 4381 3711 4385
rect 3705 4380 3711 4381
rect 3705 4376 3706 4380
rect 3710 4376 3711 4380
rect 3705 4375 3711 4376
rect 3705 4371 3706 4375
rect 3710 4371 3711 4375
rect 3705 4370 3711 4371
rect 3705 4366 3706 4370
rect 3710 4366 3711 4370
rect 3705 4365 3711 4366
rect 3705 4361 3706 4365
rect 3710 4361 3711 4365
rect 3705 4360 3711 4361
rect 3705 4356 3706 4360
rect 3710 4356 3711 4360
rect 3705 4355 3711 4356
rect 3705 4351 3706 4355
rect 3710 4351 3711 4355
rect 3705 4350 3711 4351
rect 3705 4346 3706 4350
rect 3710 4346 3711 4350
rect 3795 4461 3796 4465
rect 3800 4461 3801 4465
rect 3795 4460 3801 4461
rect 3795 4456 3796 4460
rect 3800 4456 3801 4460
rect 3795 4455 3801 4456
rect 3795 4451 3796 4455
rect 3800 4451 3801 4455
rect 3795 4450 3801 4451
rect 3795 4446 3796 4450
rect 3800 4446 3801 4450
rect 3795 4445 3801 4446
rect 3795 4441 3796 4445
rect 3800 4441 3801 4445
rect 3795 4440 3801 4441
rect 3795 4436 3796 4440
rect 3800 4436 3801 4440
rect 3795 4435 3801 4436
rect 3795 4431 3796 4435
rect 3800 4431 3801 4435
rect 3795 4430 3801 4431
rect 3795 4426 3796 4430
rect 3800 4426 3801 4430
rect 3795 4425 3801 4426
rect 3795 4421 3796 4425
rect 3800 4421 3801 4425
rect 3795 4420 3801 4421
rect 3795 4416 3796 4420
rect 3800 4416 3801 4420
rect 3795 4415 3801 4416
rect 3795 4411 3796 4415
rect 3800 4411 3801 4415
rect 3795 4410 3801 4411
rect 3795 4406 3796 4410
rect 3800 4406 3801 4410
rect 3795 4405 3801 4406
rect 3795 4401 3796 4405
rect 3800 4401 3801 4405
rect 3795 4400 3801 4401
rect 3795 4396 3796 4400
rect 3800 4396 3801 4400
rect 3795 4395 3801 4396
rect 3795 4391 3796 4395
rect 3800 4391 3801 4395
rect 3795 4390 3801 4391
rect 3795 4386 3796 4390
rect 3800 4386 3801 4390
rect 3795 4385 3801 4386
rect 3795 4381 3796 4385
rect 3800 4381 3801 4385
rect 3795 4380 3801 4381
rect 3795 4376 3796 4380
rect 3800 4376 3801 4380
rect 3795 4375 3801 4376
rect 3795 4371 3796 4375
rect 3800 4371 3801 4375
rect 3795 4370 3801 4371
rect 3795 4366 3796 4370
rect 3800 4366 3801 4370
rect 3795 4365 3801 4366
rect 3795 4361 3796 4365
rect 3800 4361 3801 4365
rect 3795 4360 3801 4361
rect 3795 4356 3796 4360
rect 3800 4356 3801 4360
rect 3795 4355 3801 4356
rect 3795 4351 3796 4355
rect 3800 4351 3801 4355
rect 3795 4350 3801 4351
rect 3705 4345 3711 4346
rect 3705 4341 3706 4345
rect 3710 4341 3711 4345
rect 3795 4346 3796 4350
rect 3800 4346 3801 4350
rect 3795 4345 3801 4346
rect 3795 4341 3796 4345
rect 3800 4341 3801 4345
rect 3705 4340 3801 4341
rect 3705 4336 3706 4340
rect 3710 4336 3711 4340
rect 3715 4336 3716 4340
rect 3720 4336 3721 4340
rect 3725 4336 3726 4340
rect 3730 4336 3731 4340
rect 3735 4336 3736 4340
rect 3740 4336 3741 4340
rect 3745 4336 3746 4340
rect 3750 4336 3751 4340
rect 3755 4336 3756 4340
rect 3760 4336 3761 4340
rect 3765 4336 3766 4340
rect 3770 4336 3771 4340
rect 3775 4336 3776 4340
rect 3780 4336 3781 4340
rect 3785 4336 3786 4340
rect 3790 4336 3791 4340
rect 3795 4336 3796 4340
rect 3800 4336 3801 4340
rect 3705 4335 3801 4336
<< psubstratepcontact >>
rect 1385 9961 1389 9965
rect 1392 9961 1396 9965
rect 1397 9961 1401 9965
rect 1402 9961 1406 9965
rect 1407 9961 1411 9965
rect 1412 9961 1416 9965
rect 1417 9961 1421 9965
rect 1422 9961 1426 9965
rect 1427 9961 1431 9965
rect 1432 9961 1436 9965
rect 1437 9961 1441 9965
rect 1442 9961 1446 9965
rect 1449 9961 1453 9965
rect 1385 9954 1389 9958
rect 1449 9954 1453 9958
rect 1385 9949 1389 9953
rect 1385 9944 1389 9948
rect 1385 9939 1389 9943
rect 1385 9934 1389 9938
rect 1385 9929 1389 9933
rect 1385 9924 1389 9928
rect 1385 9919 1389 9923
rect 1385 9914 1389 9918
rect 1385 9909 1389 9913
rect 1385 9904 1389 9908
rect 1385 9899 1389 9903
rect 1385 9894 1389 9898
rect 1385 9889 1389 9893
rect 1385 9884 1389 9888
rect 1385 9879 1389 9883
rect 1385 9874 1389 9878
rect 1385 9869 1389 9873
rect 1385 9864 1389 9868
rect 1449 9949 1453 9953
rect 1449 9944 1453 9948
rect 1449 9939 1453 9943
rect 1449 9934 1453 9938
rect 1449 9929 1453 9933
rect 1449 9924 1453 9928
rect 1449 9919 1453 9923
rect 1449 9914 1453 9918
rect 1449 9909 1453 9913
rect 1449 9904 1453 9908
rect 1449 9899 1453 9903
rect 1449 9894 1453 9898
rect 1449 9889 1453 9893
rect 1449 9884 1453 9888
rect 1449 9879 1453 9883
rect 1449 9874 1453 9878
rect 1449 9869 1453 9873
rect 1449 9864 1453 9868
rect 1385 9859 1389 9863
rect 1449 9859 1453 9863
rect 1385 9852 1389 9856
rect 1392 9852 1396 9856
rect 1397 9852 1401 9856
rect 1402 9852 1406 9856
rect 1407 9852 1411 9856
rect 1412 9852 1416 9856
rect 1417 9852 1421 9856
rect 1422 9852 1426 9856
rect 1427 9852 1431 9856
rect 1432 9852 1436 9856
rect 1437 9852 1441 9856
rect 1442 9852 1446 9856
rect 1449 9852 1453 9856
rect 1532 9974 1536 9978
rect 1537 9974 1541 9978
rect 1542 9974 1546 9978
rect 1547 9974 1551 9978
rect 1552 9974 1556 9978
rect 1557 9974 1561 9978
rect 1562 9974 1566 9978
rect 1567 9974 1571 9978
rect 1572 9974 1576 9978
rect 1577 9974 1581 9978
rect 1582 9974 1586 9978
rect 1587 9974 1591 9978
rect 1592 9974 1596 9978
rect 1597 9974 1601 9978
rect 1602 9974 1606 9978
rect 1607 9974 1611 9978
rect 1612 9974 1616 9978
rect 1617 9974 1621 9978
rect 1622 9974 1626 9978
rect 1532 9969 1536 9973
rect 1532 9964 1536 9968
rect 1622 9969 1626 9973
rect 1532 9959 1536 9963
rect 1532 9954 1536 9958
rect 1532 9949 1536 9953
rect 1532 9944 1536 9948
rect 1532 9939 1536 9943
rect 1532 9934 1536 9938
rect 1532 9929 1536 9933
rect 1532 9924 1536 9928
rect 1532 9919 1536 9923
rect 1532 9914 1536 9918
rect 1532 9909 1536 9913
rect 1532 9904 1536 9908
rect 1532 9899 1536 9903
rect 1532 9894 1536 9898
rect 1532 9889 1536 9893
rect 1532 9884 1536 9888
rect 1532 9879 1536 9883
rect 1532 9874 1536 9878
rect 1532 9869 1536 9873
rect 1532 9864 1536 9868
rect 1532 9859 1536 9863
rect 1532 9854 1536 9858
rect 1532 9849 1536 9853
rect 1622 9964 1626 9968
rect 1622 9959 1626 9963
rect 1622 9954 1626 9958
rect 1622 9949 1626 9953
rect 1622 9944 1626 9948
rect 1622 9939 1626 9943
rect 1622 9934 1626 9938
rect 1622 9929 1626 9933
rect 1622 9924 1626 9928
rect 1622 9919 1626 9923
rect 1622 9914 1626 9918
rect 1622 9909 1626 9913
rect 1622 9904 1626 9908
rect 1622 9899 1626 9903
rect 1622 9894 1626 9898
rect 1622 9889 1626 9893
rect 1622 9884 1626 9888
rect 1622 9879 1626 9883
rect 1622 9874 1626 9878
rect 1622 9869 1626 9873
rect 1622 9864 1626 9868
rect 1622 9859 1626 9863
rect 1622 9854 1626 9858
rect 1532 9844 1536 9848
rect 1622 9849 1626 9853
rect 1622 9844 1626 9848
rect 1532 9839 1536 9843
rect 1537 9839 1541 9843
rect 1542 9839 1546 9843
rect 1547 9839 1551 9843
rect 1552 9839 1556 9843
rect 1557 9839 1561 9843
rect 1562 9839 1566 9843
rect 1567 9839 1571 9843
rect 1572 9839 1576 9843
rect 1577 9839 1581 9843
rect 1582 9839 1586 9843
rect 1587 9839 1591 9843
rect 1592 9839 1596 9843
rect 1597 9839 1601 9843
rect 1602 9839 1606 9843
rect 1607 9839 1611 9843
rect 1612 9839 1616 9843
rect 1617 9839 1621 9843
rect 1622 9839 1626 9843
rect 1694 9961 1698 9965
rect 1701 9961 1705 9965
rect 1706 9961 1710 9965
rect 1711 9961 1715 9965
rect 1716 9961 1720 9965
rect 1721 9961 1725 9965
rect 1726 9961 1730 9965
rect 1731 9961 1735 9965
rect 1736 9961 1740 9965
rect 1741 9961 1745 9965
rect 1746 9961 1750 9965
rect 1751 9961 1755 9965
rect 1758 9961 1762 9965
rect 1694 9954 1698 9958
rect 1758 9954 1762 9958
rect 1694 9949 1698 9953
rect 1694 9944 1698 9948
rect 1694 9939 1698 9943
rect 1694 9934 1698 9938
rect 1694 9929 1698 9933
rect 1694 9924 1698 9928
rect 1694 9919 1698 9923
rect 1694 9914 1698 9918
rect 1694 9909 1698 9913
rect 1694 9904 1698 9908
rect 1694 9899 1698 9903
rect 1694 9894 1698 9898
rect 1694 9889 1698 9893
rect 1694 9884 1698 9888
rect 1694 9879 1698 9883
rect 1694 9874 1698 9878
rect 1694 9869 1698 9873
rect 1694 9864 1698 9868
rect 1758 9949 1762 9953
rect 1758 9944 1762 9948
rect 1758 9939 1762 9943
rect 1758 9934 1762 9938
rect 1758 9929 1762 9933
rect 1758 9924 1762 9928
rect 1758 9919 1762 9923
rect 1758 9914 1762 9918
rect 1758 9909 1762 9913
rect 1758 9904 1762 9908
rect 1758 9899 1762 9903
rect 1758 9894 1762 9898
rect 1758 9889 1762 9893
rect 1758 9884 1762 9888
rect 1758 9879 1762 9883
rect 1758 9874 1762 9878
rect 1758 9869 1762 9873
rect 1758 9864 1762 9868
rect 1694 9859 1698 9863
rect 1758 9859 1762 9863
rect 1694 9852 1698 9856
rect 1701 9852 1705 9856
rect 1706 9852 1710 9856
rect 1711 9852 1715 9856
rect 1716 9852 1720 9856
rect 1721 9852 1725 9856
rect 1726 9852 1730 9856
rect 1731 9852 1735 9856
rect 1736 9852 1740 9856
rect 1741 9852 1745 9856
rect 1746 9852 1750 9856
rect 1751 9852 1755 9856
rect 1758 9852 1762 9856
rect 1841 9974 1845 9978
rect 1846 9974 1850 9978
rect 1851 9974 1855 9978
rect 1856 9974 1860 9978
rect 1861 9974 1865 9978
rect 1866 9974 1870 9978
rect 1871 9974 1875 9978
rect 1876 9974 1880 9978
rect 1881 9974 1885 9978
rect 1886 9974 1890 9978
rect 1891 9974 1895 9978
rect 1896 9974 1900 9978
rect 1901 9974 1905 9978
rect 1906 9974 1910 9978
rect 1911 9974 1915 9978
rect 1916 9974 1920 9978
rect 1921 9974 1925 9978
rect 1926 9974 1930 9978
rect 1931 9974 1935 9978
rect 1841 9969 1845 9973
rect 1841 9964 1845 9968
rect 1931 9969 1935 9973
rect 1841 9959 1845 9963
rect 1841 9954 1845 9958
rect 1841 9949 1845 9953
rect 1841 9944 1845 9948
rect 1841 9939 1845 9943
rect 1841 9934 1845 9938
rect 1841 9929 1845 9933
rect 1841 9924 1845 9928
rect 1841 9919 1845 9923
rect 1841 9914 1845 9918
rect 1841 9909 1845 9913
rect 1841 9904 1845 9908
rect 1841 9899 1845 9903
rect 1841 9894 1845 9898
rect 1841 9889 1845 9893
rect 1841 9884 1845 9888
rect 1841 9879 1845 9883
rect 1841 9874 1845 9878
rect 1841 9869 1845 9873
rect 1841 9864 1845 9868
rect 1841 9859 1845 9863
rect 1841 9854 1845 9858
rect 1841 9849 1845 9853
rect 1931 9964 1935 9968
rect 1931 9959 1935 9963
rect 1931 9954 1935 9958
rect 1931 9949 1935 9953
rect 1931 9944 1935 9948
rect 1931 9939 1935 9943
rect 1931 9934 1935 9938
rect 1931 9929 1935 9933
rect 1931 9924 1935 9928
rect 1931 9919 1935 9923
rect 1931 9914 1935 9918
rect 1931 9909 1935 9913
rect 1931 9904 1935 9908
rect 1931 9899 1935 9903
rect 1931 9894 1935 9898
rect 1931 9889 1935 9893
rect 1931 9884 1935 9888
rect 1931 9879 1935 9883
rect 1931 9874 1935 9878
rect 1931 9869 1935 9873
rect 1931 9864 1935 9868
rect 1931 9859 1935 9863
rect 1931 9854 1935 9858
rect 1841 9844 1845 9848
rect 1931 9849 1935 9853
rect 1931 9844 1935 9848
rect 1841 9839 1845 9843
rect 1846 9839 1850 9843
rect 1851 9839 1855 9843
rect 1856 9839 1860 9843
rect 1861 9839 1865 9843
rect 1866 9839 1870 9843
rect 1871 9839 1875 9843
rect 1876 9839 1880 9843
rect 1881 9839 1885 9843
rect 1886 9839 1890 9843
rect 1891 9839 1895 9843
rect 1896 9839 1900 9843
rect 1901 9839 1905 9843
rect 1906 9839 1910 9843
rect 1911 9839 1915 9843
rect 1916 9839 1920 9843
rect 1921 9839 1925 9843
rect 1926 9839 1930 9843
rect 1931 9839 1935 9843
rect 2003 9961 2007 9965
rect 2010 9961 2014 9965
rect 2015 9961 2019 9965
rect 2020 9961 2024 9965
rect 2025 9961 2029 9965
rect 2030 9961 2034 9965
rect 2035 9961 2039 9965
rect 2040 9961 2044 9965
rect 2045 9961 2049 9965
rect 2050 9961 2054 9965
rect 2055 9961 2059 9965
rect 2060 9961 2064 9965
rect 2067 9961 2071 9965
rect 2003 9954 2007 9958
rect 2067 9954 2071 9958
rect 2003 9949 2007 9953
rect 2003 9944 2007 9948
rect 2003 9939 2007 9943
rect 2003 9934 2007 9938
rect 2003 9929 2007 9933
rect 2003 9924 2007 9928
rect 2003 9919 2007 9923
rect 2003 9914 2007 9918
rect 2003 9909 2007 9913
rect 2003 9904 2007 9908
rect 2003 9899 2007 9903
rect 2003 9894 2007 9898
rect 2003 9889 2007 9893
rect 2003 9884 2007 9888
rect 2003 9879 2007 9883
rect 2003 9874 2007 9878
rect 2003 9869 2007 9873
rect 2003 9864 2007 9868
rect 2067 9949 2071 9953
rect 2067 9944 2071 9948
rect 2067 9939 2071 9943
rect 2067 9934 2071 9938
rect 2067 9929 2071 9933
rect 2067 9924 2071 9928
rect 2067 9919 2071 9923
rect 2067 9914 2071 9918
rect 2067 9909 2071 9913
rect 2067 9904 2071 9908
rect 2067 9899 2071 9903
rect 2067 9894 2071 9898
rect 2067 9889 2071 9893
rect 2067 9884 2071 9888
rect 2067 9879 2071 9883
rect 2067 9874 2071 9878
rect 2067 9869 2071 9873
rect 2067 9864 2071 9868
rect 2003 9859 2007 9863
rect 2067 9859 2071 9863
rect 2003 9852 2007 9856
rect 2010 9852 2014 9856
rect 2015 9852 2019 9856
rect 2020 9852 2024 9856
rect 2025 9852 2029 9856
rect 2030 9852 2034 9856
rect 2035 9852 2039 9856
rect 2040 9852 2044 9856
rect 2045 9852 2049 9856
rect 2050 9852 2054 9856
rect 2055 9852 2059 9856
rect 2060 9852 2064 9856
rect 2067 9852 2071 9856
rect 2150 9974 2154 9978
rect 2155 9974 2159 9978
rect 2160 9974 2164 9978
rect 2165 9974 2169 9978
rect 2170 9974 2174 9978
rect 2175 9974 2179 9978
rect 2180 9974 2184 9978
rect 2185 9974 2189 9978
rect 2190 9974 2194 9978
rect 2195 9974 2199 9978
rect 2200 9974 2204 9978
rect 2205 9974 2209 9978
rect 2210 9974 2214 9978
rect 2215 9974 2219 9978
rect 2220 9974 2224 9978
rect 2225 9974 2229 9978
rect 2230 9974 2234 9978
rect 2235 9974 2239 9978
rect 2240 9974 2244 9978
rect 2150 9969 2154 9973
rect 2150 9964 2154 9968
rect 2240 9969 2244 9973
rect 2150 9959 2154 9963
rect 2150 9954 2154 9958
rect 2150 9949 2154 9953
rect 2150 9944 2154 9948
rect 2150 9939 2154 9943
rect 2150 9934 2154 9938
rect 2150 9929 2154 9933
rect 2150 9924 2154 9928
rect 2150 9919 2154 9923
rect 2150 9914 2154 9918
rect 2150 9909 2154 9913
rect 2150 9904 2154 9908
rect 2150 9899 2154 9903
rect 2150 9894 2154 9898
rect 2150 9889 2154 9893
rect 2150 9884 2154 9888
rect 2150 9879 2154 9883
rect 2150 9874 2154 9878
rect 2150 9869 2154 9873
rect 2150 9864 2154 9868
rect 2150 9859 2154 9863
rect 2150 9854 2154 9858
rect 2150 9849 2154 9853
rect 2240 9964 2244 9968
rect 2240 9959 2244 9963
rect 2240 9954 2244 9958
rect 2240 9949 2244 9953
rect 2240 9944 2244 9948
rect 2240 9939 2244 9943
rect 2240 9934 2244 9938
rect 2240 9929 2244 9933
rect 2240 9924 2244 9928
rect 2240 9919 2244 9923
rect 2240 9914 2244 9918
rect 2240 9909 2244 9913
rect 2240 9904 2244 9908
rect 2240 9899 2244 9903
rect 2240 9894 2244 9898
rect 2240 9889 2244 9893
rect 2240 9884 2244 9888
rect 2240 9879 2244 9883
rect 2240 9874 2244 9878
rect 2240 9869 2244 9873
rect 2240 9864 2244 9868
rect 2240 9859 2244 9863
rect 2240 9854 2244 9858
rect 2150 9844 2154 9848
rect 2240 9849 2244 9853
rect 2240 9844 2244 9848
rect 2150 9839 2154 9843
rect 2155 9839 2159 9843
rect 2160 9839 2164 9843
rect 2165 9839 2169 9843
rect 2170 9839 2174 9843
rect 2175 9839 2179 9843
rect 2180 9839 2184 9843
rect 2185 9839 2189 9843
rect 2190 9839 2194 9843
rect 2195 9839 2199 9843
rect 2200 9839 2204 9843
rect 2205 9839 2209 9843
rect 2210 9839 2214 9843
rect 2215 9839 2219 9843
rect 2220 9839 2224 9843
rect 2225 9839 2229 9843
rect 2230 9839 2234 9843
rect 2235 9839 2239 9843
rect 2240 9839 2244 9843
rect 2312 9961 2316 9965
rect 2319 9961 2323 9965
rect 2324 9961 2328 9965
rect 2329 9961 2333 9965
rect 2334 9961 2338 9965
rect 2339 9961 2343 9965
rect 2344 9961 2348 9965
rect 2349 9961 2353 9965
rect 2354 9961 2358 9965
rect 2359 9961 2363 9965
rect 2364 9961 2368 9965
rect 2369 9961 2373 9965
rect 2376 9961 2380 9965
rect 2312 9954 2316 9958
rect 2376 9954 2380 9958
rect 2312 9949 2316 9953
rect 2312 9944 2316 9948
rect 2312 9939 2316 9943
rect 2312 9934 2316 9938
rect 2312 9929 2316 9933
rect 2312 9924 2316 9928
rect 2312 9919 2316 9923
rect 2312 9914 2316 9918
rect 2312 9909 2316 9913
rect 2312 9904 2316 9908
rect 2312 9899 2316 9903
rect 2312 9894 2316 9898
rect 2312 9889 2316 9893
rect 2312 9884 2316 9888
rect 2312 9879 2316 9883
rect 2312 9874 2316 9878
rect 2312 9869 2316 9873
rect 2312 9864 2316 9868
rect 2376 9949 2380 9953
rect 2376 9944 2380 9948
rect 2376 9939 2380 9943
rect 2376 9934 2380 9938
rect 2376 9929 2380 9933
rect 2376 9924 2380 9928
rect 2376 9919 2380 9923
rect 2376 9914 2380 9918
rect 2376 9909 2380 9913
rect 2376 9904 2380 9908
rect 2376 9899 2380 9903
rect 2376 9894 2380 9898
rect 2376 9889 2380 9893
rect 2376 9884 2380 9888
rect 2376 9879 2380 9883
rect 2376 9874 2380 9878
rect 2376 9869 2380 9873
rect 2376 9864 2380 9868
rect 2312 9859 2316 9863
rect 2376 9859 2380 9863
rect 2312 9852 2316 9856
rect 2319 9852 2323 9856
rect 2324 9852 2328 9856
rect 2329 9852 2333 9856
rect 2334 9852 2338 9856
rect 2339 9852 2343 9856
rect 2344 9852 2348 9856
rect 2349 9852 2353 9856
rect 2354 9852 2358 9856
rect 2359 9852 2363 9856
rect 2364 9852 2368 9856
rect 2369 9852 2373 9856
rect 2376 9852 2380 9856
rect 2459 9974 2463 9978
rect 2464 9974 2468 9978
rect 2469 9974 2473 9978
rect 2474 9974 2478 9978
rect 2479 9974 2483 9978
rect 2484 9974 2488 9978
rect 2489 9974 2493 9978
rect 2494 9974 2498 9978
rect 2499 9974 2503 9978
rect 2504 9974 2508 9978
rect 2509 9974 2513 9978
rect 2514 9974 2518 9978
rect 2519 9974 2523 9978
rect 2524 9974 2528 9978
rect 2529 9974 2533 9978
rect 2534 9974 2538 9978
rect 2539 9974 2543 9978
rect 2544 9974 2548 9978
rect 2549 9974 2553 9978
rect 2459 9969 2463 9973
rect 2459 9964 2463 9968
rect 2549 9969 2553 9973
rect 2459 9959 2463 9963
rect 2459 9954 2463 9958
rect 2459 9949 2463 9953
rect 2459 9944 2463 9948
rect 2459 9939 2463 9943
rect 2459 9934 2463 9938
rect 2459 9929 2463 9933
rect 2459 9924 2463 9928
rect 2459 9919 2463 9923
rect 2459 9914 2463 9918
rect 2459 9909 2463 9913
rect 2459 9904 2463 9908
rect 2459 9899 2463 9903
rect 2459 9894 2463 9898
rect 2459 9889 2463 9893
rect 2459 9884 2463 9888
rect 2459 9879 2463 9883
rect 2459 9874 2463 9878
rect 2459 9869 2463 9873
rect 2459 9864 2463 9868
rect 2459 9859 2463 9863
rect 2459 9854 2463 9858
rect 2459 9849 2463 9853
rect 2549 9964 2553 9968
rect 2549 9959 2553 9963
rect 2549 9954 2553 9958
rect 2549 9949 2553 9953
rect 2549 9944 2553 9948
rect 2549 9939 2553 9943
rect 2549 9934 2553 9938
rect 2549 9929 2553 9933
rect 2549 9924 2553 9928
rect 2549 9919 2553 9923
rect 2549 9914 2553 9918
rect 2549 9909 2553 9913
rect 2549 9904 2553 9908
rect 2549 9899 2553 9903
rect 2549 9894 2553 9898
rect 2549 9889 2553 9893
rect 2549 9884 2553 9888
rect 2549 9879 2553 9883
rect 2549 9874 2553 9878
rect 2549 9869 2553 9873
rect 2549 9864 2553 9868
rect 2549 9859 2553 9863
rect 2549 9854 2553 9858
rect 2459 9844 2463 9848
rect 2549 9849 2553 9853
rect 2549 9844 2553 9848
rect 2459 9839 2463 9843
rect 2464 9839 2468 9843
rect 2469 9839 2473 9843
rect 2474 9839 2478 9843
rect 2479 9839 2483 9843
rect 2484 9839 2488 9843
rect 2489 9839 2493 9843
rect 2494 9839 2498 9843
rect 2499 9839 2503 9843
rect 2504 9839 2508 9843
rect 2509 9839 2513 9843
rect 2514 9839 2518 9843
rect 2519 9839 2523 9843
rect 2524 9839 2528 9843
rect 2529 9839 2533 9843
rect 2534 9839 2538 9843
rect 2539 9839 2543 9843
rect 2544 9839 2548 9843
rect 2549 9839 2553 9843
rect 2621 9961 2625 9965
rect 2628 9961 2632 9965
rect 2633 9961 2637 9965
rect 2638 9961 2642 9965
rect 2643 9961 2647 9965
rect 2648 9961 2652 9965
rect 2653 9961 2657 9965
rect 2658 9961 2662 9965
rect 2663 9961 2667 9965
rect 2668 9961 2672 9965
rect 2673 9961 2677 9965
rect 2678 9961 2682 9965
rect 2685 9961 2689 9965
rect 2621 9954 2625 9958
rect 2685 9954 2689 9958
rect 2621 9949 2625 9953
rect 2621 9944 2625 9948
rect 2621 9939 2625 9943
rect 2621 9934 2625 9938
rect 2621 9929 2625 9933
rect 2621 9924 2625 9928
rect 2621 9919 2625 9923
rect 2621 9914 2625 9918
rect 2621 9909 2625 9913
rect 2621 9904 2625 9908
rect 2621 9899 2625 9903
rect 2621 9894 2625 9898
rect 2621 9889 2625 9893
rect 2621 9884 2625 9888
rect 2621 9879 2625 9883
rect 2621 9874 2625 9878
rect 2621 9869 2625 9873
rect 2621 9864 2625 9868
rect 2685 9949 2689 9953
rect 2685 9944 2689 9948
rect 2685 9939 2689 9943
rect 2685 9934 2689 9938
rect 2685 9929 2689 9933
rect 2685 9924 2689 9928
rect 2685 9919 2689 9923
rect 2685 9914 2689 9918
rect 2685 9909 2689 9913
rect 2685 9904 2689 9908
rect 2685 9899 2689 9903
rect 2685 9894 2689 9898
rect 2685 9889 2689 9893
rect 2685 9884 2689 9888
rect 2685 9879 2689 9883
rect 2685 9874 2689 9878
rect 2685 9869 2689 9873
rect 2685 9864 2689 9868
rect 2621 9859 2625 9863
rect 2685 9859 2689 9863
rect 2621 9852 2625 9856
rect 2628 9852 2632 9856
rect 2633 9852 2637 9856
rect 2638 9852 2642 9856
rect 2643 9852 2647 9856
rect 2648 9852 2652 9856
rect 2653 9852 2657 9856
rect 2658 9852 2662 9856
rect 2663 9852 2667 9856
rect 2668 9852 2672 9856
rect 2673 9852 2677 9856
rect 2678 9852 2682 9856
rect 2685 9852 2689 9856
rect 2768 9974 2772 9978
rect 2773 9974 2777 9978
rect 2778 9974 2782 9978
rect 2783 9974 2787 9978
rect 2788 9974 2792 9978
rect 2793 9974 2797 9978
rect 2798 9974 2802 9978
rect 2803 9974 2807 9978
rect 2808 9974 2812 9978
rect 2813 9974 2817 9978
rect 2818 9974 2822 9978
rect 2823 9974 2827 9978
rect 2828 9974 2832 9978
rect 2833 9974 2837 9978
rect 2838 9974 2842 9978
rect 2843 9974 2847 9978
rect 2848 9974 2852 9978
rect 2853 9974 2857 9978
rect 2858 9974 2862 9978
rect 2768 9969 2772 9973
rect 2768 9964 2772 9968
rect 2858 9969 2862 9973
rect 2768 9959 2772 9963
rect 2768 9954 2772 9958
rect 2768 9949 2772 9953
rect 2768 9944 2772 9948
rect 2768 9939 2772 9943
rect 2768 9934 2772 9938
rect 2768 9929 2772 9933
rect 2768 9924 2772 9928
rect 2768 9919 2772 9923
rect 2768 9914 2772 9918
rect 2768 9909 2772 9913
rect 2768 9904 2772 9908
rect 2768 9899 2772 9903
rect 2768 9894 2772 9898
rect 2768 9889 2772 9893
rect 2768 9884 2772 9888
rect 2768 9879 2772 9883
rect 2768 9874 2772 9878
rect 2768 9869 2772 9873
rect 2768 9864 2772 9868
rect 2768 9859 2772 9863
rect 2768 9854 2772 9858
rect 2768 9849 2772 9853
rect 2858 9964 2862 9968
rect 2858 9959 2862 9963
rect 2858 9954 2862 9958
rect 2858 9949 2862 9953
rect 2858 9944 2862 9948
rect 2858 9939 2862 9943
rect 2858 9934 2862 9938
rect 2858 9929 2862 9933
rect 2858 9924 2862 9928
rect 2858 9919 2862 9923
rect 2858 9914 2862 9918
rect 2858 9909 2862 9913
rect 2858 9904 2862 9908
rect 2858 9899 2862 9903
rect 2858 9894 2862 9898
rect 2858 9889 2862 9893
rect 2858 9884 2862 9888
rect 2858 9879 2862 9883
rect 2858 9874 2862 9878
rect 2858 9869 2862 9873
rect 2858 9864 2862 9868
rect 2858 9859 2862 9863
rect 2858 9854 2862 9858
rect 2768 9844 2772 9848
rect 2858 9849 2862 9853
rect 2858 9844 2862 9848
rect 2768 9839 2772 9843
rect 2773 9839 2777 9843
rect 2778 9839 2782 9843
rect 2783 9839 2787 9843
rect 2788 9839 2792 9843
rect 2793 9839 2797 9843
rect 2798 9839 2802 9843
rect 2803 9839 2807 9843
rect 2808 9839 2812 9843
rect 2813 9839 2817 9843
rect 2818 9839 2822 9843
rect 2823 9839 2827 9843
rect 2828 9839 2832 9843
rect 2833 9839 2837 9843
rect 2838 9839 2842 9843
rect 2843 9839 2847 9843
rect 2848 9839 2852 9843
rect 2853 9839 2857 9843
rect 2858 9839 2862 9843
rect 2930 9961 2934 9965
rect 2937 9961 2941 9965
rect 2942 9961 2946 9965
rect 2947 9961 2951 9965
rect 2952 9961 2956 9965
rect 2957 9961 2961 9965
rect 2962 9961 2966 9965
rect 2967 9961 2971 9965
rect 2972 9961 2976 9965
rect 2977 9961 2981 9965
rect 2982 9961 2986 9965
rect 2987 9961 2991 9965
rect 2994 9961 2998 9965
rect 2930 9954 2934 9958
rect 2994 9954 2998 9958
rect 2930 9949 2934 9953
rect 2930 9944 2934 9948
rect 2930 9939 2934 9943
rect 2930 9934 2934 9938
rect 2930 9929 2934 9933
rect 2930 9924 2934 9928
rect 2930 9919 2934 9923
rect 2930 9914 2934 9918
rect 2930 9909 2934 9913
rect 2930 9904 2934 9908
rect 2930 9899 2934 9903
rect 2930 9894 2934 9898
rect 2930 9889 2934 9893
rect 2930 9884 2934 9888
rect 2930 9879 2934 9883
rect 2930 9874 2934 9878
rect 2930 9869 2934 9873
rect 2930 9864 2934 9868
rect 2994 9949 2998 9953
rect 2994 9944 2998 9948
rect 2994 9939 2998 9943
rect 2994 9934 2998 9938
rect 2994 9929 2998 9933
rect 2994 9924 2998 9928
rect 2994 9919 2998 9923
rect 2994 9914 2998 9918
rect 2994 9909 2998 9913
rect 2994 9904 2998 9908
rect 2994 9899 2998 9903
rect 2994 9894 2998 9898
rect 2994 9889 2998 9893
rect 2994 9884 2998 9888
rect 2994 9879 2998 9883
rect 2994 9874 2998 9878
rect 2994 9869 2998 9873
rect 2994 9864 2998 9868
rect 2930 9859 2934 9863
rect 2994 9859 2998 9863
rect 2930 9852 2934 9856
rect 2937 9852 2941 9856
rect 2942 9852 2946 9856
rect 2947 9852 2951 9856
rect 2952 9852 2956 9856
rect 2957 9852 2961 9856
rect 2962 9852 2966 9856
rect 2967 9852 2971 9856
rect 2972 9852 2976 9856
rect 2977 9852 2981 9856
rect 2982 9852 2986 9856
rect 2987 9852 2991 9856
rect 2994 9852 2998 9856
rect 3077 9974 3081 9978
rect 3082 9974 3086 9978
rect 3087 9974 3091 9978
rect 3092 9974 3096 9978
rect 3097 9974 3101 9978
rect 3102 9974 3106 9978
rect 3107 9974 3111 9978
rect 3112 9974 3116 9978
rect 3117 9974 3121 9978
rect 3122 9974 3126 9978
rect 3127 9974 3131 9978
rect 3132 9974 3136 9978
rect 3137 9974 3141 9978
rect 3142 9974 3146 9978
rect 3147 9974 3151 9978
rect 3152 9974 3156 9978
rect 3157 9974 3161 9978
rect 3162 9974 3166 9978
rect 3167 9974 3171 9978
rect 3077 9969 3081 9973
rect 3077 9964 3081 9968
rect 3167 9969 3171 9973
rect 3077 9959 3081 9963
rect 3077 9954 3081 9958
rect 3077 9949 3081 9953
rect 3077 9944 3081 9948
rect 3077 9939 3081 9943
rect 3077 9934 3081 9938
rect 3077 9929 3081 9933
rect 3077 9924 3081 9928
rect 3077 9919 3081 9923
rect 3077 9914 3081 9918
rect 3077 9909 3081 9913
rect 3077 9904 3081 9908
rect 3077 9899 3081 9903
rect 3077 9894 3081 9898
rect 3077 9889 3081 9893
rect 3077 9884 3081 9888
rect 3077 9879 3081 9883
rect 3077 9874 3081 9878
rect 3077 9869 3081 9873
rect 3077 9864 3081 9868
rect 3077 9859 3081 9863
rect 3077 9854 3081 9858
rect 3077 9849 3081 9853
rect 3167 9964 3171 9968
rect 3167 9959 3171 9963
rect 3167 9954 3171 9958
rect 3167 9949 3171 9953
rect 3167 9944 3171 9948
rect 3167 9939 3171 9943
rect 3167 9934 3171 9938
rect 3167 9929 3171 9933
rect 3167 9924 3171 9928
rect 3167 9919 3171 9923
rect 3167 9914 3171 9918
rect 3167 9909 3171 9913
rect 3167 9904 3171 9908
rect 3167 9899 3171 9903
rect 3167 9894 3171 9898
rect 3167 9889 3171 9893
rect 3167 9884 3171 9888
rect 3167 9879 3171 9883
rect 3167 9874 3171 9878
rect 3167 9869 3171 9873
rect 3167 9864 3171 9868
rect 3167 9859 3171 9863
rect 3167 9854 3171 9858
rect 3077 9844 3081 9848
rect 3167 9849 3171 9853
rect 3167 9844 3171 9848
rect 3077 9839 3081 9843
rect 3082 9839 3086 9843
rect 3087 9839 3091 9843
rect 3092 9839 3096 9843
rect 3097 9839 3101 9843
rect 3102 9839 3106 9843
rect 3107 9839 3111 9843
rect 3112 9839 3116 9843
rect 3117 9839 3121 9843
rect 3122 9839 3126 9843
rect 3127 9839 3131 9843
rect 3132 9839 3136 9843
rect 3137 9839 3141 9843
rect 3142 9839 3146 9843
rect 3147 9839 3151 9843
rect 3152 9839 3156 9843
rect 3157 9839 3161 9843
rect 3162 9839 3166 9843
rect 3167 9839 3171 9843
rect 3239 9961 3243 9965
rect 3246 9961 3250 9965
rect 3251 9961 3255 9965
rect 3256 9961 3260 9965
rect 3261 9961 3265 9965
rect 3266 9961 3270 9965
rect 3271 9961 3275 9965
rect 3276 9961 3280 9965
rect 3281 9961 3285 9965
rect 3286 9961 3290 9965
rect 3291 9961 3295 9965
rect 3296 9961 3300 9965
rect 3303 9961 3307 9965
rect 3239 9954 3243 9958
rect 3303 9954 3307 9958
rect 3239 9949 3243 9953
rect 3239 9944 3243 9948
rect 3239 9939 3243 9943
rect 3239 9934 3243 9938
rect 3239 9929 3243 9933
rect 3239 9924 3243 9928
rect 3239 9919 3243 9923
rect 3239 9914 3243 9918
rect 3239 9909 3243 9913
rect 3239 9904 3243 9908
rect 3239 9899 3243 9903
rect 3239 9894 3243 9898
rect 3239 9889 3243 9893
rect 3239 9884 3243 9888
rect 3239 9879 3243 9883
rect 3239 9874 3243 9878
rect 3239 9869 3243 9873
rect 3239 9864 3243 9868
rect 3303 9949 3307 9953
rect 3303 9944 3307 9948
rect 3303 9939 3307 9943
rect 3303 9934 3307 9938
rect 3303 9929 3307 9933
rect 3303 9924 3307 9928
rect 3303 9919 3307 9923
rect 3303 9914 3307 9918
rect 3303 9909 3307 9913
rect 3303 9904 3307 9908
rect 3303 9899 3307 9903
rect 3303 9894 3307 9898
rect 3303 9889 3307 9893
rect 3303 9884 3307 9888
rect 3303 9879 3307 9883
rect 3303 9874 3307 9878
rect 3303 9869 3307 9873
rect 3303 9864 3307 9868
rect 3239 9859 3243 9863
rect 3303 9859 3307 9863
rect 3239 9852 3243 9856
rect 3246 9852 3250 9856
rect 3251 9852 3255 9856
rect 3256 9852 3260 9856
rect 3261 9852 3265 9856
rect 3266 9852 3270 9856
rect 3271 9852 3275 9856
rect 3276 9852 3280 9856
rect 3281 9852 3285 9856
rect 3286 9852 3290 9856
rect 3291 9852 3295 9856
rect 3296 9852 3300 9856
rect 3303 9852 3307 9856
rect 3386 9974 3390 9978
rect 3391 9974 3395 9978
rect 3396 9974 3400 9978
rect 3401 9974 3405 9978
rect 3406 9974 3410 9978
rect 3411 9974 3415 9978
rect 3416 9974 3420 9978
rect 3421 9974 3425 9978
rect 3426 9974 3430 9978
rect 3431 9974 3435 9978
rect 3436 9974 3440 9978
rect 3441 9974 3445 9978
rect 3446 9974 3450 9978
rect 3451 9974 3455 9978
rect 3456 9974 3460 9978
rect 3461 9974 3465 9978
rect 3466 9974 3470 9978
rect 3471 9974 3475 9978
rect 3476 9974 3480 9978
rect 3386 9969 3390 9973
rect 3386 9964 3390 9968
rect 3476 9969 3480 9973
rect 3386 9959 3390 9963
rect 3386 9954 3390 9958
rect 3386 9949 3390 9953
rect 3386 9944 3390 9948
rect 3386 9939 3390 9943
rect 3386 9934 3390 9938
rect 3386 9929 3390 9933
rect 3386 9924 3390 9928
rect 3386 9919 3390 9923
rect 3386 9914 3390 9918
rect 3386 9909 3390 9913
rect 3386 9904 3390 9908
rect 3386 9899 3390 9903
rect 3386 9894 3390 9898
rect 3386 9889 3390 9893
rect 3386 9884 3390 9888
rect 3386 9879 3390 9883
rect 3386 9874 3390 9878
rect 3386 9869 3390 9873
rect 3386 9864 3390 9868
rect 3386 9859 3390 9863
rect 3386 9854 3390 9858
rect 3386 9849 3390 9853
rect 3476 9964 3480 9968
rect 3476 9959 3480 9963
rect 3476 9954 3480 9958
rect 3476 9949 3480 9953
rect 3476 9944 3480 9948
rect 3476 9939 3480 9943
rect 3476 9934 3480 9938
rect 3476 9929 3480 9933
rect 3476 9924 3480 9928
rect 3476 9919 3480 9923
rect 3476 9914 3480 9918
rect 3476 9909 3480 9913
rect 3476 9904 3480 9908
rect 3476 9899 3480 9903
rect 3476 9894 3480 9898
rect 3476 9889 3480 9893
rect 3476 9884 3480 9888
rect 3476 9879 3480 9883
rect 3476 9874 3480 9878
rect 3476 9869 3480 9873
rect 3476 9864 3480 9868
rect 3476 9859 3480 9863
rect 3476 9854 3480 9858
rect 3386 9844 3390 9848
rect 3476 9849 3480 9853
rect 3476 9844 3480 9848
rect 3386 9839 3390 9843
rect 3391 9839 3395 9843
rect 3396 9839 3400 9843
rect 3401 9839 3405 9843
rect 3406 9839 3410 9843
rect 3411 9839 3415 9843
rect 3416 9839 3420 9843
rect 3421 9839 3425 9843
rect 3426 9839 3430 9843
rect 3431 9839 3435 9843
rect 3436 9839 3440 9843
rect 3441 9839 3445 9843
rect 3446 9839 3450 9843
rect 3451 9839 3455 9843
rect 3456 9839 3460 9843
rect 3461 9839 3465 9843
rect 3466 9839 3470 9843
rect 3471 9839 3475 9843
rect 3476 9839 3480 9843
rect 3548 9961 3552 9965
rect 3555 9961 3559 9965
rect 3560 9961 3564 9965
rect 3565 9961 3569 9965
rect 3570 9961 3574 9965
rect 3575 9961 3579 9965
rect 3580 9961 3584 9965
rect 3585 9961 3589 9965
rect 3590 9961 3594 9965
rect 3595 9961 3599 9965
rect 3600 9961 3604 9965
rect 3605 9961 3609 9965
rect 3612 9961 3616 9965
rect 3548 9954 3552 9958
rect 3612 9954 3616 9958
rect 3548 9949 3552 9953
rect 3548 9944 3552 9948
rect 3548 9939 3552 9943
rect 3548 9934 3552 9938
rect 3548 9929 3552 9933
rect 3548 9924 3552 9928
rect 3548 9919 3552 9923
rect 3548 9914 3552 9918
rect 3548 9909 3552 9913
rect 3548 9904 3552 9908
rect 3548 9899 3552 9903
rect 3548 9894 3552 9898
rect 3548 9889 3552 9893
rect 3548 9884 3552 9888
rect 3548 9879 3552 9883
rect 3548 9874 3552 9878
rect 3548 9869 3552 9873
rect 3548 9864 3552 9868
rect 3612 9949 3616 9953
rect 3612 9944 3616 9948
rect 3612 9939 3616 9943
rect 3612 9934 3616 9938
rect 3612 9929 3616 9933
rect 3612 9924 3616 9928
rect 3612 9919 3616 9923
rect 3612 9914 3616 9918
rect 3612 9909 3616 9913
rect 3612 9904 3616 9908
rect 3612 9899 3616 9903
rect 3612 9894 3616 9898
rect 3612 9889 3616 9893
rect 3612 9884 3616 9888
rect 3612 9879 3616 9883
rect 3612 9874 3616 9878
rect 3612 9869 3616 9873
rect 3612 9864 3616 9868
rect 3548 9859 3552 9863
rect 3612 9859 3616 9863
rect 3548 9852 3552 9856
rect 3555 9852 3559 9856
rect 3560 9852 3564 9856
rect 3565 9852 3569 9856
rect 3570 9852 3574 9856
rect 3575 9852 3579 9856
rect 3580 9852 3584 9856
rect 3585 9852 3589 9856
rect 3590 9852 3594 9856
rect 3595 9852 3599 9856
rect 3600 9852 3604 9856
rect 3605 9852 3609 9856
rect 3612 9852 3616 9856
rect 3695 9974 3699 9978
rect 3700 9974 3704 9978
rect 3705 9974 3709 9978
rect 3710 9974 3714 9978
rect 3715 9974 3719 9978
rect 3720 9974 3724 9978
rect 3725 9974 3729 9978
rect 3730 9974 3734 9978
rect 3735 9974 3739 9978
rect 3740 9974 3744 9978
rect 3745 9974 3749 9978
rect 3750 9974 3754 9978
rect 3755 9974 3759 9978
rect 3760 9974 3764 9978
rect 3765 9974 3769 9978
rect 3770 9974 3774 9978
rect 3775 9974 3779 9978
rect 3780 9974 3784 9978
rect 3785 9974 3789 9978
rect 3695 9969 3699 9973
rect 3695 9964 3699 9968
rect 3785 9969 3789 9973
rect 3695 9959 3699 9963
rect 3695 9954 3699 9958
rect 3695 9949 3699 9953
rect 3695 9944 3699 9948
rect 3695 9939 3699 9943
rect 3695 9934 3699 9938
rect 3695 9929 3699 9933
rect 3695 9924 3699 9928
rect 3695 9919 3699 9923
rect 3695 9914 3699 9918
rect 3695 9909 3699 9913
rect 3695 9904 3699 9908
rect 3695 9899 3699 9903
rect 3695 9894 3699 9898
rect 3695 9889 3699 9893
rect 3695 9884 3699 9888
rect 3695 9879 3699 9883
rect 3695 9874 3699 9878
rect 3695 9869 3699 9873
rect 3695 9864 3699 9868
rect 3695 9859 3699 9863
rect 3695 9854 3699 9858
rect 3695 9849 3699 9853
rect 3785 9964 3789 9968
rect 3785 9959 3789 9963
rect 3785 9954 3789 9958
rect 3785 9949 3789 9953
rect 3785 9944 3789 9948
rect 3785 9939 3789 9943
rect 3785 9934 3789 9938
rect 3785 9929 3789 9933
rect 3785 9924 3789 9928
rect 3785 9919 3789 9923
rect 3785 9914 3789 9918
rect 3785 9909 3789 9913
rect 3785 9904 3789 9908
rect 3785 9899 3789 9903
rect 3785 9894 3789 9898
rect 3785 9889 3789 9893
rect 3785 9884 3789 9888
rect 3785 9879 3789 9883
rect 3785 9874 3789 9878
rect 3785 9869 3789 9873
rect 3785 9864 3789 9868
rect 3785 9859 3789 9863
rect 3785 9854 3789 9858
rect 3695 9844 3699 9848
rect 3785 9849 3789 9853
rect 3785 9844 3789 9848
rect 3695 9839 3699 9843
rect 3700 9839 3704 9843
rect 3705 9839 3709 9843
rect 3710 9839 3714 9843
rect 3715 9839 3719 9843
rect 3720 9839 3724 9843
rect 3725 9839 3729 9843
rect 3730 9839 3734 9843
rect 3735 9839 3739 9843
rect 3740 9839 3744 9843
rect 3745 9839 3749 9843
rect 3750 9839 3754 9843
rect 3755 9839 3759 9843
rect 3760 9839 3764 9843
rect 3765 9839 3769 9843
rect 3770 9839 3774 9843
rect 3775 9839 3779 9843
rect 3780 9839 3784 9843
rect 3785 9839 3789 9843
rect 3857 9961 3861 9965
rect 3864 9961 3868 9965
rect 3869 9961 3873 9965
rect 3874 9961 3878 9965
rect 3879 9961 3883 9965
rect 3884 9961 3888 9965
rect 3889 9961 3893 9965
rect 3894 9961 3898 9965
rect 3899 9961 3903 9965
rect 3904 9961 3908 9965
rect 3909 9961 3913 9965
rect 3914 9961 3918 9965
rect 3921 9961 3925 9965
rect 3857 9954 3861 9958
rect 3921 9954 3925 9958
rect 3857 9949 3861 9953
rect 3857 9944 3861 9948
rect 3857 9939 3861 9943
rect 3857 9934 3861 9938
rect 3857 9929 3861 9933
rect 3857 9924 3861 9928
rect 3857 9919 3861 9923
rect 3857 9914 3861 9918
rect 3857 9909 3861 9913
rect 3857 9904 3861 9908
rect 3857 9899 3861 9903
rect 3857 9894 3861 9898
rect 3857 9889 3861 9893
rect 3857 9884 3861 9888
rect 3857 9879 3861 9883
rect 3857 9874 3861 9878
rect 3857 9869 3861 9873
rect 3857 9864 3861 9868
rect 3921 9949 3925 9953
rect 3921 9944 3925 9948
rect 3921 9939 3925 9943
rect 3921 9934 3925 9938
rect 3921 9929 3925 9933
rect 3921 9924 3925 9928
rect 3921 9919 3925 9923
rect 3921 9914 3925 9918
rect 3921 9909 3925 9913
rect 3921 9904 3925 9908
rect 3921 9899 3925 9903
rect 3921 9894 3925 9898
rect 3921 9889 3925 9893
rect 3921 9884 3925 9888
rect 3921 9879 3925 9883
rect 3921 9874 3925 9878
rect 3921 9869 3925 9873
rect 3921 9864 3925 9868
rect 3857 9859 3861 9863
rect 3921 9859 3925 9863
rect 3857 9852 3861 9856
rect 3864 9852 3868 9856
rect 3869 9852 3873 9856
rect 3874 9852 3878 9856
rect 3879 9852 3883 9856
rect 3884 9852 3888 9856
rect 3889 9852 3893 9856
rect 3894 9852 3898 9856
rect 3899 9852 3903 9856
rect 3904 9852 3908 9856
rect 3909 9852 3913 9856
rect 3914 9852 3918 9856
rect 3921 9852 3925 9856
rect 4004 9974 4008 9978
rect 4009 9974 4013 9978
rect 4014 9974 4018 9978
rect 4019 9974 4023 9978
rect 4024 9974 4028 9978
rect 4029 9974 4033 9978
rect 4034 9974 4038 9978
rect 4039 9974 4043 9978
rect 4044 9974 4048 9978
rect 4049 9974 4053 9978
rect 4054 9974 4058 9978
rect 4059 9974 4063 9978
rect 4064 9974 4068 9978
rect 4069 9974 4073 9978
rect 4074 9974 4078 9978
rect 4079 9974 4083 9978
rect 4084 9974 4088 9978
rect 4089 9974 4093 9978
rect 4094 9974 4098 9978
rect 4004 9969 4008 9973
rect 4004 9964 4008 9968
rect 4094 9969 4098 9973
rect 4004 9959 4008 9963
rect 4004 9954 4008 9958
rect 4004 9949 4008 9953
rect 4004 9944 4008 9948
rect 4004 9939 4008 9943
rect 4004 9934 4008 9938
rect 4004 9929 4008 9933
rect 4004 9924 4008 9928
rect 4004 9919 4008 9923
rect 4004 9914 4008 9918
rect 4004 9909 4008 9913
rect 4004 9904 4008 9908
rect 4004 9899 4008 9903
rect 4004 9894 4008 9898
rect 4004 9889 4008 9893
rect 4004 9884 4008 9888
rect 4004 9879 4008 9883
rect 4004 9874 4008 9878
rect 4004 9869 4008 9873
rect 4004 9864 4008 9868
rect 4004 9859 4008 9863
rect 4004 9854 4008 9858
rect 4004 9849 4008 9853
rect 4094 9964 4098 9968
rect 4094 9959 4098 9963
rect 4094 9954 4098 9958
rect 4094 9949 4098 9953
rect 4094 9944 4098 9948
rect 4094 9939 4098 9943
rect 4094 9934 4098 9938
rect 4094 9929 4098 9933
rect 4094 9924 4098 9928
rect 4094 9919 4098 9923
rect 4094 9914 4098 9918
rect 4094 9909 4098 9913
rect 4094 9904 4098 9908
rect 4094 9899 4098 9903
rect 4094 9894 4098 9898
rect 4094 9889 4098 9893
rect 4094 9884 4098 9888
rect 4094 9879 4098 9883
rect 4094 9874 4098 9878
rect 4094 9869 4098 9873
rect 4094 9864 4098 9868
rect 4094 9859 4098 9863
rect 4094 9854 4098 9858
rect 4004 9844 4008 9848
rect 4094 9849 4098 9853
rect 4094 9844 4098 9848
rect 4004 9839 4008 9843
rect 4009 9839 4013 9843
rect 4014 9839 4018 9843
rect 4019 9839 4023 9843
rect 4024 9839 4028 9843
rect 4029 9839 4033 9843
rect 4034 9839 4038 9843
rect 4039 9839 4043 9843
rect 4044 9839 4048 9843
rect 4049 9839 4053 9843
rect 4054 9839 4058 9843
rect 4059 9839 4063 9843
rect 4064 9839 4068 9843
rect 4069 9839 4073 9843
rect 4074 9839 4078 9843
rect 4079 9839 4083 9843
rect 4084 9839 4088 9843
rect 4089 9839 4093 9843
rect 4094 9839 4098 9843
rect 418 6280 422 6339
rect 459 6280 463 6339
rect 502 6280 506 6339
rect 541 6299 545 6339
rect 802 9716 806 9720
rect 807 9716 811 9720
rect 812 9716 816 9720
rect 817 9716 821 9720
rect 831 9716 835 9720
rect 836 9716 840 9720
rect 841 9716 845 9720
rect 846 9716 850 9720
rect 860 9716 864 9720
rect 865 9716 869 9720
rect 870 9716 874 9720
rect 875 9716 879 9720
rect 889 9716 893 9720
rect 894 9716 898 9720
rect 899 9716 903 9720
rect 904 9716 908 9720
rect 918 9716 922 9720
rect 923 9716 927 9720
rect 928 9716 932 9720
rect 933 9716 937 9720
rect 1319 9716 1323 9720
rect 1324 9716 1328 9720
rect 1329 9716 1333 9720
rect 1334 9716 1338 9720
rect 1628 9716 1632 9720
rect 1633 9716 1637 9720
rect 1638 9716 1642 9720
rect 1643 9716 1647 9720
rect 1937 9716 1941 9720
rect 1942 9716 1946 9720
rect 1947 9716 1951 9720
rect 1952 9716 1956 9720
rect 2246 9716 2250 9720
rect 2251 9716 2255 9720
rect 2256 9716 2260 9720
rect 2261 9716 2265 9720
rect 2555 9716 2559 9720
rect 2560 9716 2564 9720
rect 2565 9716 2569 9720
rect 2570 9716 2574 9720
rect 2864 9716 2868 9720
rect 2869 9716 2873 9720
rect 2874 9716 2878 9720
rect 2879 9716 2883 9720
rect 3173 9716 3177 9720
rect 3178 9716 3182 9720
rect 3183 9716 3187 9720
rect 3188 9716 3192 9720
rect 3482 9716 3486 9720
rect 3487 9716 3491 9720
rect 3492 9716 3496 9720
rect 3497 9716 3501 9720
rect 3791 9716 3795 9720
rect 3796 9716 3800 9720
rect 3801 9716 3805 9720
rect 3806 9716 3810 9720
rect 4100 9716 4104 9720
rect 4105 9716 4109 9720
rect 4110 9716 4114 9720
rect 4115 9716 4119 9720
rect 4292 9716 4296 9720
rect 4297 9716 4301 9720
rect 4302 9716 4306 9720
rect 4307 9716 4311 9720
rect 4318 9716 4322 9720
rect 4323 9716 4327 9720
rect 4328 9716 4332 9720
rect 4333 9716 4337 9720
rect 4344 9716 4348 9720
rect 4349 9716 4353 9720
rect 4354 9716 4358 9720
rect 4359 9716 4363 9720
rect 4370 9716 4374 9720
rect 4375 9716 4379 9720
rect 4380 9716 4384 9720
rect 4385 9716 4389 9720
rect 4396 9716 4400 9720
rect 4401 9716 4405 9720
rect 4406 9716 4410 9720
rect 4411 9716 4415 9720
rect 802 9706 806 9710
rect 807 9706 811 9710
rect 812 9706 816 9710
rect 817 9706 821 9710
rect 831 9706 835 9710
rect 836 9706 840 9710
rect 841 9706 845 9710
rect 846 9706 850 9710
rect 860 9706 864 9710
rect 865 9706 869 9710
rect 870 9706 874 9710
rect 875 9706 879 9710
rect 889 9706 893 9710
rect 894 9706 898 9710
rect 899 9706 903 9710
rect 904 9706 908 9710
rect 918 9706 922 9710
rect 923 9706 927 9710
rect 928 9706 932 9710
rect 933 9706 937 9710
rect 1319 9706 1323 9710
rect 1324 9706 1328 9710
rect 1329 9706 1333 9710
rect 1334 9706 1338 9710
rect 1628 9706 1632 9710
rect 1633 9706 1637 9710
rect 1638 9706 1642 9710
rect 1643 9706 1647 9710
rect 1937 9706 1941 9710
rect 1942 9706 1946 9710
rect 1947 9706 1951 9710
rect 1952 9706 1956 9710
rect 2246 9706 2250 9710
rect 2251 9706 2255 9710
rect 2256 9706 2260 9710
rect 2261 9706 2265 9710
rect 2555 9706 2559 9710
rect 2560 9706 2564 9710
rect 2565 9706 2569 9710
rect 2570 9706 2574 9710
rect 2864 9706 2868 9710
rect 2869 9706 2873 9710
rect 2874 9706 2878 9710
rect 2879 9706 2883 9710
rect 3173 9706 3177 9710
rect 3178 9706 3182 9710
rect 3183 9706 3187 9710
rect 3188 9706 3192 9710
rect 3482 9706 3486 9710
rect 3487 9706 3491 9710
rect 3492 9706 3496 9710
rect 3497 9706 3501 9710
rect 3791 9706 3795 9710
rect 3796 9706 3800 9710
rect 3801 9706 3805 9710
rect 3806 9706 3810 9710
rect 4100 9706 4104 9710
rect 4105 9706 4109 9710
rect 4110 9706 4114 9710
rect 4115 9706 4119 9710
rect 4292 9706 4296 9710
rect 4297 9706 4301 9710
rect 4302 9706 4306 9710
rect 4307 9706 4311 9710
rect 4318 9706 4322 9710
rect 4323 9706 4327 9710
rect 4328 9706 4332 9710
rect 4333 9706 4337 9710
rect 4344 9706 4348 9710
rect 4349 9706 4353 9710
rect 4354 9706 4358 9710
rect 4359 9706 4363 9710
rect 4370 9706 4374 9710
rect 4375 9706 4379 9710
rect 4380 9706 4384 9710
rect 4385 9706 4389 9710
rect 4396 9706 4400 9710
rect 4401 9706 4405 9710
rect 4406 9706 4410 9710
rect 4411 9706 4415 9710
rect 802 9696 806 9700
rect 807 9696 811 9700
rect 812 9696 816 9700
rect 817 9696 821 9700
rect 831 9696 835 9700
rect 836 9696 840 9700
rect 841 9696 845 9700
rect 846 9696 850 9700
rect 860 9696 864 9700
rect 865 9696 869 9700
rect 870 9696 874 9700
rect 875 9696 879 9700
rect 889 9696 893 9700
rect 894 9696 898 9700
rect 899 9696 903 9700
rect 904 9696 908 9700
rect 918 9696 922 9700
rect 923 9696 927 9700
rect 928 9696 932 9700
rect 933 9696 937 9700
rect 1319 9696 1323 9700
rect 1324 9696 1328 9700
rect 1329 9696 1333 9700
rect 1334 9696 1338 9700
rect 1628 9696 1632 9700
rect 1633 9696 1637 9700
rect 1638 9696 1642 9700
rect 1643 9696 1647 9700
rect 1937 9696 1941 9700
rect 1942 9696 1946 9700
rect 1947 9696 1951 9700
rect 1952 9696 1956 9700
rect 2246 9696 2250 9700
rect 2251 9696 2255 9700
rect 2256 9696 2260 9700
rect 2261 9696 2265 9700
rect 2555 9696 2559 9700
rect 2560 9696 2564 9700
rect 2565 9696 2569 9700
rect 2570 9696 2574 9700
rect 2864 9696 2868 9700
rect 2869 9696 2873 9700
rect 2874 9696 2878 9700
rect 2879 9696 2883 9700
rect 3173 9696 3177 9700
rect 3178 9696 3182 9700
rect 3183 9696 3187 9700
rect 3188 9696 3192 9700
rect 3482 9696 3486 9700
rect 3487 9696 3491 9700
rect 3492 9696 3496 9700
rect 3497 9696 3501 9700
rect 3791 9696 3795 9700
rect 3796 9696 3800 9700
rect 3801 9696 3805 9700
rect 3806 9696 3810 9700
rect 4100 9696 4104 9700
rect 4105 9696 4109 9700
rect 4110 9696 4114 9700
rect 4115 9696 4119 9700
rect 4292 9696 4296 9700
rect 4297 9696 4301 9700
rect 4302 9696 4306 9700
rect 4307 9696 4311 9700
rect 4318 9696 4322 9700
rect 4323 9696 4327 9700
rect 4328 9696 4332 9700
rect 4333 9696 4337 9700
rect 4344 9696 4348 9700
rect 4349 9696 4353 9700
rect 4354 9696 4358 9700
rect 4359 9696 4363 9700
rect 4370 9696 4374 9700
rect 4375 9696 4379 9700
rect 4380 9696 4384 9700
rect 4385 9696 4389 9700
rect 4396 9696 4400 9700
rect 4401 9696 4405 9700
rect 4406 9696 4410 9700
rect 4411 9696 4415 9700
rect 802 9686 806 9690
rect 807 9686 811 9690
rect 812 9686 816 9690
rect 817 9686 821 9690
rect 831 9686 835 9690
rect 836 9686 840 9690
rect 841 9686 845 9690
rect 846 9686 850 9690
rect 860 9686 864 9690
rect 865 9686 869 9690
rect 870 9686 874 9690
rect 875 9686 879 9690
rect 889 9686 893 9690
rect 894 9686 898 9690
rect 899 9686 903 9690
rect 904 9686 908 9690
rect 918 9686 922 9690
rect 923 9686 927 9690
rect 928 9686 932 9690
rect 933 9686 937 9690
rect 1319 9686 1323 9690
rect 1324 9686 1328 9690
rect 1329 9686 1333 9690
rect 1334 9686 1338 9690
rect 1628 9686 1632 9690
rect 1633 9686 1637 9690
rect 1638 9686 1642 9690
rect 1643 9686 1647 9690
rect 1937 9686 1941 9690
rect 1942 9686 1946 9690
rect 1947 9686 1951 9690
rect 1952 9686 1956 9690
rect 2246 9686 2250 9690
rect 2251 9686 2255 9690
rect 2256 9686 2260 9690
rect 2261 9686 2265 9690
rect 2555 9686 2559 9690
rect 2560 9686 2564 9690
rect 2565 9686 2569 9690
rect 2570 9686 2574 9690
rect 2864 9686 2868 9690
rect 2869 9686 2873 9690
rect 2874 9686 2878 9690
rect 2879 9686 2883 9690
rect 3173 9686 3177 9690
rect 3178 9686 3182 9690
rect 3183 9686 3187 9690
rect 3188 9686 3192 9690
rect 3482 9686 3486 9690
rect 3487 9686 3491 9690
rect 3492 9686 3496 9690
rect 3497 9686 3501 9690
rect 3791 9686 3795 9690
rect 3796 9686 3800 9690
rect 3801 9686 3805 9690
rect 3806 9686 3810 9690
rect 4100 9686 4104 9690
rect 4105 9686 4109 9690
rect 4110 9686 4114 9690
rect 4115 9686 4119 9690
rect 4292 9686 4296 9690
rect 4297 9686 4301 9690
rect 4302 9686 4306 9690
rect 4307 9686 4311 9690
rect 4318 9686 4322 9690
rect 4323 9686 4327 9690
rect 4328 9686 4332 9690
rect 4333 9686 4337 9690
rect 4344 9686 4348 9690
rect 4349 9686 4353 9690
rect 4354 9686 4358 9690
rect 4359 9686 4363 9690
rect 4370 9686 4374 9690
rect 4375 9686 4379 9690
rect 4380 9686 4384 9690
rect 4385 9686 4389 9690
rect 4396 9686 4400 9690
rect 4401 9686 4405 9690
rect 4406 9686 4410 9690
rect 4411 9686 4415 9690
rect 659 9618 663 9622
rect 669 9618 673 9622
rect 679 9618 683 9622
rect 689 9618 693 9622
rect 659 9613 663 9617
rect 669 9613 673 9617
rect 679 9613 683 9617
rect 689 9613 693 9617
rect 659 9608 663 9612
rect 669 9608 673 9612
rect 679 9608 683 9612
rect 689 9608 693 9612
rect 659 9603 663 9607
rect 669 9603 673 9607
rect 679 9603 683 9607
rect 689 9603 693 9607
rect 659 9592 663 9596
rect 669 9592 673 9596
rect 679 9592 683 9596
rect 689 9592 693 9596
rect 659 9587 663 9591
rect 669 9587 673 9591
rect 679 9587 683 9591
rect 689 9587 693 9591
rect 659 9582 663 9586
rect 669 9582 673 9586
rect 679 9582 683 9586
rect 689 9582 693 9586
rect 659 9577 663 9581
rect 669 9577 673 9581
rect 679 9577 683 9581
rect 689 9577 693 9581
rect 659 9566 663 9570
rect 669 9566 673 9570
rect 679 9566 683 9570
rect 689 9566 693 9570
rect 659 9561 663 9565
rect 669 9561 673 9565
rect 679 9561 683 9565
rect 689 9561 693 9565
rect 659 9556 663 9560
rect 669 9556 673 9560
rect 679 9556 683 9560
rect 689 9556 693 9560
rect 659 9551 663 9555
rect 669 9551 673 9555
rect 679 9551 683 9555
rect 689 9551 693 9555
rect 659 9540 663 9544
rect 669 9540 673 9544
rect 679 9540 683 9544
rect 689 9540 693 9544
rect 659 9535 663 9539
rect 669 9535 673 9539
rect 679 9535 683 9539
rect 689 9535 693 9539
rect 659 9530 663 9534
rect 669 9530 673 9534
rect 679 9530 683 9534
rect 689 9530 693 9534
rect 659 9525 663 9529
rect 669 9525 673 9529
rect 679 9525 683 9529
rect 689 9525 693 9529
rect 659 9514 663 9518
rect 669 9514 673 9518
rect 679 9514 683 9518
rect 689 9514 693 9518
rect 659 9509 663 9513
rect 669 9509 673 9513
rect 679 9509 683 9513
rect 689 9509 693 9513
rect 659 9504 663 9508
rect 669 9504 673 9508
rect 679 9504 683 9508
rect 689 9504 693 9508
rect 659 9499 663 9503
rect 669 9499 673 9503
rect 679 9499 683 9503
rect 689 9499 693 9503
rect 4479 9573 4483 9577
rect 4489 9573 4493 9577
rect 4499 9573 4503 9577
rect 4509 9573 4513 9577
rect 4479 9568 4483 9572
rect 4489 9568 4493 9572
rect 4499 9568 4503 9572
rect 4509 9568 4513 9572
rect 4479 9563 4483 9567
rect 4489 9563 4493 9567
rect 4499 9563 4503 9567
rect 4509 9563 4513 9567
rect 4479 9558 4483 9562
rect 4489 9558 4493 9562
rect 4499 9558 4503 9562
rect 4509 9558 4513 9562
rect 4479 9544 4483 9548
rect 4489 9544 4493 9548
rect 4499 9544 4503 9548
rect 4509 9544 4513 9548
rect 4479 9539 4483 9543
rect 4489 9539 4493 9543
rect 4499 9539 4503 9543
rect 4509 9539 4513 9543
rect 4479 9534 4483 9538
rect 4489 9534 4493 9538
rect 4499 9534 4503 9538
rect 4509 9534 4513 9538
rect 4479 9529 4483 9533
rect 4489 9529 4493 9533
rect 4499 9529 4503 9533
rect 4509 9529 4513 9533
rect 4479 9515 4483 9519
rect 4489 9515 4493 9519
rect 4499 9515 4503 9519
rect 4509 9515 4513 9519
rect 4479 9510 4483 9514
rect 4489 9510 4493 9514
rect 4499 9510 4503 9514
rect 4509 9510 4513 9514
rect 4479 9505 4483 9509
rect 4489 9505 4493 9509
rect 4499 9505 4503 9509
rect 4509 9505 4513 9509
rect 4479 9500 4483 9504
rect 4489 9500 4493 9504
rect 4499 9500 4503 9504
rect 4509 9500 4513 9504
rect 4479 9486 4483 9490
rect 4489 9486 4493 9490
rect 4499 9486 4503 9490
rect 4509 9486 4513 9490
rect 4479 9481 4483 9485
rect 4489 9481 4493 9485
rect 4499 9481 4503 9485
rect 4509 9481 4513 9485
rect 4479 9476 4483 9480
rect 4489 9476 4493 9480
rect 4499 9476 4503 9480
rect 4509 9476 4513 9480
rect 4479 9471 4483 9475
rect 4489 9471 4493 9475
rect 4499 9471 4503 9475
rect 4509 9471 4513 9475
rect 4479 9457 4483 9461
rect 4489 9457 4493 9461
rect 4499 9457 4503 9461
rect 4509 9457 4513 9461
rect 4479 9452 4483 9456
rect 4489 9452 4493 9456
rect 4499 9452 4503 9456
rect 4509 9452 4513 9456
rect 4479 9447 4483 9451
rect 4489 9447 4493 9451
rect 4499 9447 4503 9451
rect 4509 9447 4513 9451
rect 4479 9442 4483 9446
rect 4489 9442 4493 9446
rect 4499 9442 4503 9446
rect 4509 9442 4513 9446
rect 659 9321 663 9325
rect 669 9321 673 9325
rect 679 9321 683 9325
rect 689 9321 693 9325
rect 659 9316 663 9320
rect 669 9316 673 9320
rect 679 9316 683 9320
rect 689 9316 693 9320
rect 659 9311 663 9315
rect 669 9311 673 9315
rect 679 9311 683 9315
rect 689 9311 693 9315
rect 659 9306 663 9310
rect 669 9306 673 9310
rect 679 9306 683 9310
rect 689 9306 693 9310
rect 2881 9283 2885 9287
rect 2909 9283 2913 9287
rect 2939 9283 2943 9287
rect 3013 9283 3017 9287
rect 3041 9283 3045 9287
rect 3071 9283 3075 9287
rect 3145 9283 3149 9287
rect 3173 9283 3177 9287
rect 3203 9283 3207 9287
rect 3277 9283 3281 9287
rect 3305 9283 3309 9287
rect 3335 9283 3339 9287
rect 3826 9283 3830 9287
rect 3854 9283 3858 9287
rect 3884 9283 3888 9287
rect 3958 9283 3962 9287
rect 3986 9283 3990 9287
rect 4016 9283 4020 9287
rect 4090 9283 4094 9287
rect 4118 9283 4122 9287
rect 4148 9283 4152 9287
rect 4222 9283 4226 9287
rect 4250 9283 4254 9287
rect 4280 9283 4284 9287
rect 2529 9250 2533 9254
rect 2557 9250 2561 9254
rect 2587 9250 2591 9254
rect 3474 9250 3478 9254
rect 3502 9250 3506 9254
rect 3532 9250 3536 9254
rect 2862 9197 2866 9201
rect 2897 9197 2901 9201
rect 3023 9197 3027 9201
rect 3047 9197 3051 9201
rect 3101 9197 3108 9201
rect 3128 9197 3132 9201
rect 3182 9197 3186 9201
rect 3807 9197 3811 9201
rect 3842 9197 3846 9201
rect 3968 9197 3972 9201
rect 3992 9197 3996 9201
rect 4046 9197 4053 9201
rect 4073 9197 4077 9201
rect 4127 9197 4131 9201
rect 2526 9148 2530 9152
rect 2556 9148 2560 9152
rect 2584 9148 2588 9152
rect 3471 9148 3475 9152
rect 3501 9148 3505 9152
rect 3529 9148 3533 9152
rect 2862 9065 2866 9069
rect 2897 9065 2901 9069
rect 3023 9065 3027 9069
rect 3047 9065 3051 9069
rect 3101 9065 3105 9069
rect 3128 9065 3132 9069
rect 3152 9065 3156 9069
rect 3807 9065 3811 9069
rect 3842 9065 3846 9069
rect 3968 9065 3972 9069
rect 3992 9065 3996 9069
rect 4046 9065 4050 9069
rect 4073 9065 4077 9069
rect 4097 9065 4101 9069
rect 4479 9056 4483 9060
rect 4489 9056 4493 9060
rect 4499 9056 4503 9060
rect 4509 9056 4513 9060
rect 4479 9051 4483 9055
rect 4489 9051 4493 9055
rect 4499 9051 4503 9055
rect 4509 9051 4513 9055
rect 4479 9046 4483 9050
rect 4489 9046 4493 9050
rect 4499 9046 4503 9050
rect 4509 9046 4513 9050
rect 4479 9041 4483 9045
rect 4489 9041 4493 9045
rect 4499 9041 4503 9045
rect 4509 9041 4513 9045
rect 3359 9022 3363 9026
rect 3383 9022 3387 9026
rect 3437 9022 3441 9026
rect 3580 9022 3584 9026
rect 659 9012 663 9016
rect 669 9012 673 9016
rect 679 9012 683 9016
rect 689 9012 693 9016
rect 659 9007 663 9011
rect 669 9007 673 9011
rect 679 9007 683 9011
rect 689 9007 693 9011
rect 659 9002 663 9006
rect 669 9002 673 9006
rect 679 9002 683 9006
rect 689 9002 693 9006
rect 659 8997 663 9001
rect 669 8997 673 9001
rect 679 8997 683 9001
rect 689 8997 693 9001
rect 2862 8933 2866 8937
rect 2897 8933 2901 8937
rect 3023 8933 3027 8937
rect 3047 8933 3051 8937
rect 3101 8933 3108 8937
rect 3128 8933 3132 8937
rect 3182 8933 3186 8937
rect 3218 8933 3222 8937
rect 3272 8933 3276 8937
rect 3807 8933 3811 8937
rect 3842 8933 3846 8937
rect 3968 8933 3972 8937
rect 3992 8933 3996 8937
rect 4046 8933 4053 8937
rect 4073 8933 4077 8937
rect 4127 8933 4131 8937
rect 4163 8933 4167 8937
rect 4217 8933 4221 8937
rect 3337 8892 3341 8896
rect 3359 8892 3363 8896
rect 3383 8892 3387 8896
rect 3437 8892 3441 8896
rect 3486 8892 3490 8896
rect 2862 8801 2866 8805
rect 2897 8801 2901 8805
rect 3023 8801 3027 8805
rect 3047 8801 3051 8805
rect 3158 8801 3162 8805
rect 3807 8801 3811 8805
rect 3842 8801 3846 8805
rect 3968 8801 3972 8805
rect 3992 8801 3996 8805
rect 4103 8801 4107 8805
rect 2397 8748 2401 8752
rect 2425 8748 2429 8752
rect 2455 8748 2459 8752
rect 2529 8748 2533 8752
rect 2557 8748 2561 8752
rect 2587 8748 2591 8752
rect 2661 8748 2665 8752
rect 2689 8748 2693 8752
rect 2719 8748 2723 8752
rect 3342 8748 3346 8752
rect 3370 8748 3374 8752
rect 3400 8748 3404 8752
rect 3474 8748 3478 8752
rect 3502 8748 3506 8752
rect 3532 8748 3536 8752
rect 3606 8748 3610 8752
rect 3634 8748 3638 8752
rect 3664 8748 3668 8752
rect 4479 8747 4483 8751
rect 4489 8747 4493 8751
rect 4499 8747 4503 8751
rect 4509 8747 4513 8751
rect 4479 8742 4483 8746
rect 4489 8742 4493 8746
rect 4499 8742 4503 8746
rect 4509 8742 4513 8746
rect 4479 8737 4483 8741
rect 4489 8737 4493 8741
rect 4499 8737 4503 8741
rect 4509 8737 4513 8741
rect 4479 8732 4483 8736
rect 4489 8732 4493 8736
rect 4499 8732 4503 8736
rect 4509 8732 4513 8736
rect 659 8703 663 8707
rect 669 8703 673 8707
rect 679 8703 683 8707
rect 689 8703 693 8707
rect 659 8698 663 8702
rect 669 8698 673 8702
rect 679 8698 683 8702
rect 689 8698 693 8702
rect 659 8693 663 8697
rect 669 8693 673 8697
rect 679 8693 683 8697
rect 689 8693 693 8697
rect 659 8688 663 8692
rect 669 8688 673 8692
rect 679 8688 683 8692
rect 689 8688 693 8692
rect 3180 8636 3184 8640
rect 3208 8636 3212 8640
rect 3238 8636 3242 8640
rect 4125 8636 4129 8640
rect 4153 8636 4157 8640
rect 4183 8636 4187 8640
rect 2397 8606 2401 8610
rect 2425 8606 2429 8610
rect 2455 8606 2459 8610
rect 2529 8606 2533 8610
rect 2557 8606 2561 8610
rect 2587 8606 2591 8610
rect 2661 8606 2665 8610
rect 2689 8606 2693 8610
rect 2719 8606 2723 8610
rect 3342 8606 3346 8610
rect 3370 8606 3374 8610
rect 3400 8606 3404 8610
rect 3474 8606 3478 8610
rect 3502 8606 3506 8610
rect 3532 8606 3536 8610
rect 3606 8606 3610 8610
rect 3634 8606 3638 8610
rect 3664 8606 3668 8610
rect 3180 8550 3184 8554
rect 3208 8550 3212 8554
rect 3238 8550 3242 8554
rect 4125 8550 4129 8554
rect 4153 8550 4157 8554
rect 4183 8550 4187 8554
rect 2397 8520 2401 8524
rect 2425 8520 2429 8524
rect 2455 8520 2459 8524
rect 2529 8520 2533 8524
rect 2557 8520 2561 8524
rect 2587 8520 2591 8524
rect 2661 8520 2665 8524
rect 2689 8520 2693 8524
rect 2719 8520 2723 8524
rect 3342 8520 3346 8524
rect 3370 8520 3374 8524
rect 3400 8520 3404 8524
rect 3474 8520 3478 8524
rect 3502 8520 3506 8524
rect 3532 8520 3536 8524
rect 3606 8520 3610 8524
rect 3634 8520 3638 8524
rect 3664 8520 3668 8524
rect 4479 8438 4483 8442
rect 4489 8438 4493 8442
rect 4499 8438 4503 8442
rect 4509 8438 4513 8442
rect 4479 8433 4483 8437
rect 4489 8433 4493 8437
rect 4499 8433 4503 8437
rect 4509 8433 4513 8437
rect 4479 8428 4483 8432
rect 4489 8428 4493 8432
rect 4499 8428 4503 8432
rect 4509 8428 4513 8432
rect 4479 8423 4483 8427
rect 4489 8423 4493 8427
rect 4499 8423 4503 8427
rect 4509 8423 4513 8427
rect 659 8394 663 8398
rect 669 8394 673 8398
rect 679 8394 683 8398
rect 689 8394 693 8398
rect 659 8389 663 8393
rect 669 8389 673 8393
rect 679 8389 683 8393
rect 689 8389 693 8393
rect 659 8384 663 8388
rect 669 8384 673 8388
rect 679 8384 683 8388
rect 689 8384 693 8388
rect 659 8379 663 8383
rect 669 8379 673 8383
rect 679 8379 683 8383
rect 689 8379 693 8383
rect 2397 8380 2401 8384
rect 2425 8380 2429 8384
rect 2455 8380 2459 8384
rect 2529 8380 2533 8384
rect 2557 8380 2561 8384
rect 2587 8380 2591 8384
rect 2661 8380 2665 8384
rect 2689 8380 2693 8384
rect 2719 8380 2723 8384
rect 3342 8380 3346 8384
rect 3370 8380 3374 8384
rect 3400 8380 3404 8384
rect 3474 8380 3478 8384
rect 3502 8380 3506 8384
rect 3532 8380 3536 8384
rect 3606 8380 3610 8384
rect 3634 8380 3638 8384
rect 3664 8380 3668 8384
rect 2881 8301 2885 8305
rect 2909 8301 2913 8305
rect 2939 8301 2943 8305
rect 3013 8301 3017 8305
rect 3041 8301 3045 8305
rect 3071 8301 3075 8305
rect 3145 8301 3149 8305
rect 3173 8301 3177 8305
rect 3203 8301 3207 8305
rect 3277 8301 3281 8305
rect 3305 8301 3309 8305
rect 3335 8301 3339 8305
rect 3826 8301 3830 8305
rect 3854 8301 3858 8305
rect 3884 8301 3888 8305
rect 3958 8301 3962 8305
rect 3986 8301 3990 8305
rect 4016 8301 4020 8305
rect 4090 8301 4094 8305
rect 4118 8301 4122 8305
rect 4148 8301 4152 8305
rect 4222 8301 4226 8305
rect 4250 8301 4254 8305
rect 4280 8301 4284 8305
rect 2529 8268 2533 8272
rect 2557 8268 2561 8272
rect 2587 8268 2591 8272
rect 3474 8268 3478 8272
rect 3502 8268 3506 8272
rect 3532 8268 3536 8272
rect 2862 8215 2866 8219
rect 2897 8215 2901 8219
rect 3023 8215 3027 8219
rect 3047 8215 3051 8219
rect 3101 8215 3108 8219
rect 3128 8215 3132 8219
rect 3182 8215 3186 8219
rect 3807 8215 3811 8219
rect 3842 8215 3846 8219
rect 3968 8215 3972 8219
rect 3992 8215 3996 8219
rect 4046 8215 4053 8219
rect 4073 8215 4077 8219
rect 4127 8215 4131 8219
rect 2526 8166 2530 8170
rect 2556 8166 2560 8170
rect 2584 8166 2588 8170
rect 3471 8166 3475 8170
rect 3501 8166 3505 8170
rect 3529 8166 3533 8170
rect 4479 8129 4483 8133
rect 4489 8129 4493 8133
rect 4499 8129 4503 8133
rect 4509 8129 4513 8133
rect 4479 8124 4483 8128
rect 4489 8124 4493 8128
rect 4499 8124 4503 8128
rect 4509 8124 4513 8128
rect 4479 8119 4483 8123
rect 4489 8119 4493 8123
rect 4499 8119 4503 8123
rect 4509 8119 4513 8123
rect 4479 8114 4483 8118
rect 4489 8114 4493 8118
rect 4499 8114 4503 8118
rect 4509 8114 4513 8118
rect 4479 8098 4483 8102
rect 4489 8098 4493 8102
rect 4499 8098 4503 8102
rect 4509 8098 4513 8102
rect 659 8085 663 8089
rect 669 8085 673 8089
rect 679 8085 683 8089
rect 689 8085 693 8089
rect 4479 8093 4483 8097
rect 4489 8093 4493 8097
rect 4499 8093 4503 8097
rect 4509 8093 4513 8097
rect 4479 8088 4483 8092
rect 4489 8088 4493 8092
rect 4499 8088 4503 8092
rect 4509 8088 4513 8092
rect 659 8080 663 8084
rect 669 8080 673 8084
rect 679 8080 683 8084
rect 689 8080 693 8084
rect 2862 8083 2866 8087
rect 2897 8083 2901 8087
rect 3023 8083 3027 8087
rect 3047 8083 3051 8087
rect 3101 8083 3105 8087
rect 3128 8083 3132 8087
rect 3152 8083 3156 8087
rect 3807 8083 3811 8087
rect 3842 8083 3846 8087
rect 3968 8083 3972 8087
rect 3992 8083 3996 8087
rect 4046 8083 4050 8087
rect 4073 8083 4077 8087
rect 4097 8083 4101 8087
rect 4479 8083 4483 8087
rect 4489 8083 4493 8087
rect 4499 8083 4503 8087
rect 4509 8083 4513 8087
rect 659 8075 663 8079
rect 669 8075 673 8079
rect 679 8075 683 8079
rect 689 8075 693 8079
rect 659 8070 663 8074
rect 669 8070 673 8074
rect 679 8070 683 8074
rect 689 8070 693 8074
rect 2862 7951 2866 7955
rect 2897 7951 2901 7955
rect 3023 7951 3027 7955
rect 3047 7951 3051 7955
rect 3101 7951 3108 7955
rect 3128 7951 3132 7955
rect 3182 7951 3186 7955
rect 3218 7951 3222 7955
rect 3272 7951 3276 7955
rect 3807 7951 3811 7955
rect 3842 7951 3846 7955
rect 3968 7951 3972 7955
rect 3992 7951 3996 7955
rect 4046 7951 4053 7955
rect 4073 7951 4077 7955
rect 4127 7951 4131 7955
rect 4163 7951 4167 7955
rect 4217 7951 4221 7955
rect 2862 7819 2866 7823
rect 2897 7819 2901 7823
rect 3023 7819 3027 7823
rect 3047 7819 3051 7823
rect 3158 7819 3162 7823
rect 3807 7819 3811 7823
rect 3842 7819 3846 7823
rect 3968 7819 3972 7823
rect 3992 7819 3996 7823
rect 4103 7819 4107 7823
rect 659 7776 663 7780
rect 669 7776 673 7780
rect 679 7776 683 7780
rect 689 7776 693 7780
rect 659 7771 663 7775
rect 669 7771 673 7775
rect 679 7771 683 7775
rect 689 7771 693 7775
rect 659 7766 663 7770
rect 669 7766 673 7770
rect 679 7766 683 7770
rect 689 7766 693 7770
rect 2397 7766 2401 7770
rect 2425 7766 2429 7770
rect 2455 7766 2459 7770
rect 2529 7766 2533 7770
rect 2557 7766 2561 7770
rect 2587 7766 2591 7770
rect 2661 7766 2665 7770
rect 2689 7766 2693 7770
rect 2719 7766 2723 7770
rect 659 7761 663 7765
rect 669 7761 673 7765
rect 679 7761 683 7765
rect 689 7761 693 7765
rect 4479 7789 4483 7793
rect 4489 7789 4493 7793
rect 4499 7789 4503 7793
rect 4509 7789 4513 7793
rect 4479 7784 4483 7788
rect 4489 7784 4493 7788
rect 4499 7784 4503 7788
rect 4509 7784 4513 7788
rect 3342 7766 3346 7770
rect 3370 7766 3374 7770
rect 3400 7766 3404 7770
rect 3474 7766 3478 7770
rect 3502 7766 3506 7770
rect 3532 7766 3536 7770
rect 3606 7766 3610 7770
rect 3634 7766 3638 7770
rect 3664 7766 3668 7770
rect 4479 7779 4483 7783
rect 4489 7779 4493 7783
rect 4499 7779 4503 7783
rect 4509 7779 4513 7783
rect 4479 7774 4483 7778
rect 4489 7774 4493 7778
rect 4499 7774 4503 7778
rect 4509 7774 4513 7778
rect 3180 7654 3184 7658
rect 3208 7654 3212 7658
rect 3238 7654 3242 7658
rect 4125 7654 4129 7658
rect 4153 7654 4157 7658
rect 4183 7654 4187 7658
rect 2397 7624 2401 7628
rect 2425 7624 2429 7628
rect 2455 7624 2459 7628
rect 2529 7624 2533 7628
rect 2557 7624 2561 7628
rect 2587 7624 2591 7628
rect 2661 7624 2665 7628
rect 2689 7624 2693 7628
rect 2719 7624 2723 7628
rect 3342 7624 3346 7628
rect 3370 7624 3374 7628
rect 3400 7624 3404 7628
rect 3474 7624 3478 7628
rect 3502 7624 3506 7628
rect 3532 7624 3536 7628
rect 3606 7624 3610 7628
rect 3634 7624 3638 7628
rect 3664 7624 3668 7628
rect 3180 7568 3184 7572
rect 3208 7568 3212 7572
rect 3238 7568 3242 7572
rect 4125 7568 4129 7572
rect 4153 7568 4157 7572
rect 4183 7568 4187 7572
rect 2397 7538 2401 7542
rect 2425 7538 2429 7542
rect 2455 7538 2459 7542
rect 2529 7538 2533 7542
rect 2557 7538 2561 7542
rect 2587 7538 2591 7542
rect 2661 7538 2665 7542
rect 2689 7538 2693 7542
rect 2719 7538 2723 7542
rect 3342 7538 3346 7542
rect 3370 7538 3374 7542
rect 3400 7538 3404 7542
rect 3474 7538 3478 7542
rect 3502 7538 3506 7542
rect 3532 7538 3536 7542
rect 3606 7538 3610 7542
rect 3634 7538 3638 7542
rect 3664 7538 3668 7542
rect 659 7467 663 7471
rect 669 7467 673 7471
rect 679 7467 683 7471
rect 689 7467 693 7471
rect 659 7462 663 7466
rect 669 7462 673 7466
rect 679 7462 683 7466
rect 689 7462 693 7466
rect 659 7457 663 7461
rect 669 7457 673 7461
rect 679 7457 683 7461
rect 689 7457 693 7461
rect 659 7452 663 7456
rect 669 7452 673 7456
rect 679 7452 683 7456
rect 689 7452 693 7456
rect 2397 7398 2401 7402
rect 2425 7398 2429 7402
rect 2455 7398 2459 7402
rect 2529 7398 2533 7402
rect 2557 7398 2561 7402
rect 2587 7398 2591 7402
rect 2661 7398 2665 7402
rect 2689 7398 2693 7402
rect 2719 7398 2723 7402
rect 3342 7398 3346 7402
rect 3370 7398 3374 7402
rect 3400 7398 3404 7402
rect 3474 7398 3478 7402
rect 3502 7398 3506 7402
rect 3532 7398 3536 7402
rect 3606 7398 3610 7402
rect 3634 7398 3638 7402
rect 3664 7398 3668 7402
rect 659 7158 663 7162
rect 669 7158 673 7162
rect 679 7158 683 7162
rect 689 7158 693 7162
rect 659 7123 663 7127
rect 669 7123 673 7127
rect 679 7123 683 7127
rect 689 7123 693 7127
rect 659 7118 663 7122
rect 669 7118 673 7122
rect 679 7118 683 7122
rect 689 7118 693 7122
rect 659 7113 663 7117
rect 669 7113 673 7117
rect 679 7113 683 7117
rect 689 7113 693 7117
rect 659 7108 663 7112
rect 669 7108 673 7112
rect 679 7108 683 7112
rect 689 7108 693 7112
rect 4479 7230 4483 7234
rect 4489 7230 4493 7234
rect 4499 7230 4503 7234
rect 4509 7230 4513 7234
rect 4479 7225 4483 7229
rect 4489 7225 4493 7229
rect 4499 7225 4503 7229
rect 4509 7225 4513 7229
rect 4479 7220 4483 7224
rect 4489 7220 4493 7224
rect 4499 7220 4503 7224
rect 4509 7220 4513 7224
rect 4479 7215 4483 7219
rect 4489 7215 4493 7219
rect 4499 7215 4503 7219
rect 4509 7215 4513 7219
rect 4479 7202 4483 7206
rect 4489 7202 4493 7206
rect 4499 7202 4503 7206
rect 4509 7202 4513 7206
rect 4479 7197 4483 7201
rect 4489 7197 4493 7201
rect 4499 7197 4503 7201
rect 4509 7197 4513 7201
rect 4479 7192 4483 7196
rect 4489 7192 4493 7196
rect 4499 7192 4503 7196
rect 4509 7192 4513 7196
rect 4479 7187 4483 7191
rect 4489 7187 4493 7191
rect 4499 7187 4503 7191
rect 4509 7187 4513 7191
rect 4479 7152 4483 7156
rect 4489 7152 4493 7156
rect 4499 7152 4503 7156
rect 4509 7152 4513 7156
rect 1504 6912 1508 6916
rect 1534 6912 1538 6916
rect 1562 6912 1566 6916
rect 1636 6912 1640 6916
rect 1666 6912 1670 6916
rect 1694 6912 1698 6916
rect 1768 6912 1772 6916
rect 1798 6912 1802 6916
rect 1826 6912 1830 6916
rect 2449 6912 2453 6916
rect 2479 6912 2483 6916
rect 2507 6912 2511 6916
rect 2581 6912 2585 6916
rect 2611 6912 2615 6916
rect 2639 6912 2643 6916
rect 2713 6912 2717 6916
rect 2743 6912 2747 6916
rect 2771 6912 2775 6916
rect 4479 6858 4483 6862
rect 4489 6858 4493 6862
rect 4499 6858 4503 6862
rect 4509 6858 4513 6862
rect 4479 6853 4483 6857
rect 4489 6853 4493 6857
rect 4499 6853 4503 6857
rect 4509 6853 4513 6857
rect 4479 6848 4483 6852
rect 4489 6848 4493 6852
rect 4499 6848 4503 6852
rect 4509 6848 4513 6852
rect 4479 6843 4483 6847
rect 4489 6843 4493 6847
rect 4499 6843 4503 6847
rect 4509 6843 4513 6847
rect 1504 6772 1508 6776
rect 1534 6772 1538 6776
rect 1562 6772 1566 6776
rect 1636 6772 1640 6776
rect 1666 6772 1670 6776
rect 1694 6772 1698 6776
rect 1768 6772 1772 6776
rect 1798 6772 1802 6776
rect 1826 6772 1830 6776
rect 2449 6772 2453 6776
rect 2479 6772 2483 6776
rect 2507 6772 2511 6776
rect 2581 6772 2585 6776
rect 2611 6772 2615 6776
rect 2639 6772 2643 6776
rect 2713 6772 2717 6776
rect 2743 6772 2747 6776
rect 2771 6772 2775 6776
rect 985 6742 989 6746
rect 1015 6742 1019 6746
rect 1043 6742 1047 6746
rect 1930 6742 1934 6746
rect 1960 6742 1964 6746
rect 1988 6742 1992 6746
rect 1504 6686 1508 6690
rect 1534 6686 1538 6690
rect 1562 6686 1566 6690
rect 1636 6686 1640 6690
rect 1666 6686 1670 6690
rect 1694 6686 1698 6690
rect 1768 6686 1772 6690
rect 1798 6686 1802 6690
rect 1826 6686 1830 6690
rect 2449 6686 2453 6690
rect 2479 6686 2483 6690
rect 2507 6686 2511 6690
rect 2581 6686 2585 6690
rect 2611 6686 2615 6690
rect 2639 6686 2643 6690
rect 2713 6686 2717 6690
rect 2743 6686 2747 6690
rect 2771 6686 2775 6690
rect 985 6656 989 6660
rect 1015 6656 1019 6660
rect 1043 6656 1047 6660
rect 1930 6656 1934 6660
rect 1960 6656 1964 6660
rect 1988 6656 1992 6660
rect 659 6536 663 6540
rect 669 6536 673 6540
rect 679 6536 683 6540
rect 689 6536 693 6540
rect 659 6531 663 6535
rect 669 6531 673 6535
rect 679 6531 683 6535
rect 689 6531 693 6535
rect 1504 6544 1508 6548
rect 1534 6544 1538 6548
rect 1562 6544 1566 6548
rect 1636 6544 1640 6548
rect 1666 6544 1670 6548
rect 1694 6544 1698 6548
rect 1768 6544 1772 6548
rect 1798 6544 1802 6548
rect 1826 6544 1830 6548
rect 659 6526 663 6530
rect 669 6526 673 6530
rect 679 6526 683 6530
rect 689 6526 693 6530
rect 659 6521 663 6525
rect 669 6521 673 6525
rect 679 6521 683 6525
rect 689 6521 693 6525
rect 4479 6549 4483 6553
rect 4489 6549 4493 6553
rect 4499 6549 4503 6553
rect 4509 6549 4513 6553
rect 2449 6544 2453 6548
rect 2479 6544 2483 6548
rect 2507 6544 2511 6548
rect 2581 6544 2585 6548
rect 2611 6544 2615 6548
rect 2639 6544 2643 6548
rect 2713 6544 2717 6548
rect 2743 6544 2747 6548
rect 2771 6544 2775 6548
rect 4479 6544 4483 6548
rect 4489 6544 4493 6548
rect 4499 6544 4503 6548
rect 4509 6544 4513 6548
rect 4479 6539 4483 6543
rect 4489 6539 4493 6543
rect 4499 6539 4503 6543
rect 4509 6539 4513 6543
rect 4479 6534 4483 6538
rect 4489 6534 4493 6538
rect 4499 6534 4503 6538
rect 4509 6534 4513 6538
rect 1065 6491 1069 6495
rect 1176 6491 1180 6495
rect 1200 6491 1204 6495
rect 1326 6491 1330 6495
rect 1361 6491 1365 6495
rect 2010 6491 2014 6495
rect 2121 6491 2125 6495
rect 2145 6491 2149 6495
rect 2271 6491 2275 6495
rect 2306 6491 2310 6495
rect 951 6359 955 6363
rect 1005 6359 1009 6363
rect 1041 6359 1045 6363
rect 1095 6359 1099 6363
rect 1119 6359 1126 6363
rect 1176 6359 1180 6363
rect 1200 6359 1204 6363
rect 1326 6359 1330 6363
rect 1361 6359 1365 6363
rect 1896 6359 1900 6363
rect 1950 6359 1954 6363
rect 1986 6359 1990 6363
rect 2040 6359 2044 6363
rect 2064 6359 2071 6363
rect 2121 6359 2125 6363
rect 2145 6359 2149 6363
rect 2271 6359 2275 6363
rect 2306 6359 2310 6363
rect 4479 6240 4483 6244
rect 4489 6240 4493 6244
rect 4499 6240 4503 6244
rect 4509 6240 4513 6244
rect 4479 6235 4483 6239
rect 4489 6235 4493 6239
rect 4499 6235 4503 6239
rect 4509 6235 4513 6239
rect 659 6227 663 6231
rect 669 6227 673 6231
rect 679 6227 683 6231
rect 689 6227 693 6231
rect 1071 6227 1075 6231
rect 1095 6227 1099 6231
rect 1122 6227 1126 6231
rect 1176 6227 1180 6231
rect 1200 6227 1204 6231
rect 1326 6227 1330 6231
rect 1361 6227 1365 6231
rect 2016 6227 2020 6231
rect 2040 6227 2044 6231
rect 2067 6227 2071 6231
rect 2121 6227 2125 6231
rect 2145 6227 2149 6231
rect 2271 6227 2275 6231
rect 2306 6227 2310 6231
rect 4479 6230 4483 6234
rect 4489 6230 4493 6234
rect 4499 6230 4503 6234
rect 4509 6230 4513 6234
rect 659 6222 663 6226
rect 669 6222 673 6226
rect 679 6222 683 6226
rect 689 6222 693 6226
rect 659 6217 663 6221
rect 669 6217 673 6221
rect 679 6217 683 6221
rect 689 6217 693 6221
rect 4479 6225 4483 6229
rect 4489 6225 4493 6229
rect 4499 6225 4503 6229
rect 4509 6225 4513 6229
rect 659 6212 663 6216
rect 669 6212 673 6216
rect 679 6212 683 6216
rect 689 6212 693 6216
rect 659 6196 663 6200
rect 669 6196 673 6200
rect 679 6196 683 6200
rect 689 6196 693 6200
rect 659 6191 663 6195
rect 669 6191 673 6195
rect 679 6191 683 6195
rect 689 6191 693 6195
rect 659 6186 663 6190
rect 669 6186 673 6190
rect 679 6186 683 6190
rect 689 6186 693 6190
rect 659 6181 663 6185
rect 669 6181 673 6185
rect 679 6181 683 6185
rect 689 6181 693 6185
rect 1639 6144 1643 6148
rect 1667 6144 1671 6148
rect 1697 6144 1701 6148
rect 2584 6144 2588 6148
rect 2612 6144 2616 6148
rect 2642 6144 2646 6148
rect 1041 6095 1045 6099
rect 1095 6095 1099 6099
rect 1119 6095 1126 6099
rect 1176 6095 1180 6099
rect 1200 6095 1204 6099
rect 1326 6095 1330 6099
rect 1361 6095 1365 6099
rect 1986 6095 1990 6099
rect 2040 6095 2044 6099
rect 2064 6095 2071 6099
rect 2121 6095 2125 6099
rect 2145 6095 2149 6099
rect 2271 6095 2275 6099
rect 2306 6095 2310 6099
rect 1636 6042 1640 6046
rect 1666 6042 1670 6046
rect 1694 6042 1698 6046
rect 2581 6042 2585 6046
rect 2611 6042 2615 6046
rect 2639 6042 2643 6046
rect 888 6009 892 6013
rect 918 6009 922 6013
rect 946 6009 950 6013
rect 1020 6009 1024 6013
rect 1050 6009 1054 6013
rect 1078 6009 1082 6013
rect 1152 6009 1156 6013
rect 1182 6009 1186 6013
rect 1210 6009 1214 6013
rect 1284 6009 1288 6013
rect 1314 6009 1318 6013
rect 1342 6009 1346 6013
rect 1833 6009 1837 6013
rect 1863 6009 1867 6013
rect 1891 6009 1895 6013
rect 1965 6009 1969 6013
rect 1995 6009 1999 6013
rect 2023 6009 2027 6013
rect 2097 6009 2101 6013
rect 2127 6009 2131 6013
rect 2155 6009 2159 6013
rect 2229 6009 2233 6013
rect 2259 6009 2263 6013
rect 2287 6009 2291 6013
rect 1504 5930 1508 5934
rect 1534 5930 1538 5934
rect 1562 5930 1566 5934
rect 1636 5930 1640 5934
rect 1666 5930 1670 5934
rect 1694 5930 1698 5934
rect 1768 5930 1772 5934
rect 1798 5930 1802 5934
rect 1826 5930 1830 5934
rect 2449 5930 2453 5934
rect 2479 5930 2483 5934
rect 2507 5930 2511 5934
rect 2581 5930 2585 5934
rect 2611 5930 2615 5934
rect 2639 5930 2643 5934
rect 2713 5930 2717 5934
rect 2743 5930 2747 5934
rect 2771 5930 2775 5934
rect 4479 5931 4483 5935
rect 4489 5931 4493 5935
rect 4499 5931 4503 5935
rect 4509 5931 4513 5935
rect 4479 5926 4483 5930
rect 4489 5926 4493 5930
rect 4499 5926 4503 5930
rect 4509 5926 4513 5930
rect 4479 5921 4483 5925
rect 4489 5921 4493 5925
rect 4499 5921 4503 5925
rect 4509 5921 4513 5925
rect 4479 5916 4483 5920
rect 4489 5916 4493 5920
rect 4499 5916 4503 5920
rect 4509 5916 4513 5920
rect 659 5887 663 5891
rect 669 5887 673 5891
rect 679 5887 683 5891
rect 689 5887 693 5891
rect 659 5882 663 5886
rect 669 5882 673 5886
rect 679 5882 683 5886
rect 689 5882 693 5886
rect 659 5877 663 5881
rect 669 5877 673 5881
rect 679 5877 683 5881
rect 689 5877 693 5881
rect 659 5872 663 5876
rect 669 5872 673 5876
rect 679 5872 683 5876
rect 689 5872 693 5876
rect 1504 5790 1508 5794
rect 1534 5790 1538 5794
rect 1562 5790 1566 5794
rect 1636 5790 1640 5794
rect 1666 5790 1670 5794
rect 1694 5790 1698 5794
rect 1768 5790 1772 5794
rect 1798 5790 1802 5794
rect 1826 5790 1830 5794
rect 2449 5790 2453 5794
rect 2479 5790 2483 5794
rect 2507 5790 2511 5794
rect 2581 5790 2585 5794
rect 2611 5790 2615 5794
rect 2639 5790 2643 5794
rect 2713 5790 2717 5794
rect 2743 5790 2747 5794
rect 2771 5790 2775 5794
rect 985 5760 989 5764
rect 1015 5760 1019 5764
rect 1043 5760 1047 5764
rect 1930 5760 1934 5764
rect 1960 5760 1964 5764
rect 1988 5760 1992 5764
rect 1504 5704 1508 5708
rect 1534 5704 1538 5708
rect 1562 5704 1566 5708
rect 1636 5704 1640 5708
rect 1666 5704 1670 5708
rect 1694 5704 1698 5708
rect 1768 5704 1772 5708
rect 1798 5704 1802 5708
rect 1826 5704 1830 5708
rect 2449 5704 2453 5708
rect 2479 5704 2483 5708
rect 2507 5704 2511 5708
rect 2581 5704 2585 5708
rect 2611 5704 2615 5708
rect 2639 5704 2643 5708
rect 2713 5704 2717 5708
rect 2743 5704 2747 5708
rect 2771 5704 2775 5708
rect 985 5674 989 5678
rect 1015 5674 1019 5678
rect 1043 5674 1047 5678
rect 1930 5674 1934 5678
rect 1960 5674 1964 5678
rect 1988 5674 1992 5678
rect 4479 5622 4483 5626
rect 4489 5622 4493 5626
rect 4499 5622 4503 5626
rect 4509 5622 4513 5626
rect 4479 5617 4483 5621
rect 4489 5617 4493 5621
rect 4499 5617 4503 5621
rect 4509 5617 4513 5621
rect 4479 5612 4483 5616
rect 4489 5612 4493 5616
rect 4499 5612 4503 5616
rect 4509 5612 4513 5616
rect 4479 5607 4483 5611
rect 4489 5607 4493 5611
rect 4499 5607 4503 5611
rect 4509 5607 4513 5611
rect 659 5578 663 5582
rect 669 5578 673 5582
rect 679 5578 683 5582
rect 689 5578 693 5582
rect 659 5573 663 5577
rect 669 5573 673 5577
rect 679 5573 683 5577
rect 689 5573 693 5577
rect 659 5568 663 5572
rect 669 5568 673 5572
rect 679 5568 683 5572
rect 689 5568 693 5572
rect 659 5563 663 5567
rect 669 5563 673 5567
rect 679 5563 683 5567
rect 689 5563 693 5567
rect 1504 5562 1508 5566
rect 1534 5562 1538 5566
rect 1562 5562 1566 5566
rect 1636 5562 1640 5566
rect 1666 5562 1670 5566
rect 1694 5562 1698 5566
rect 1768 5562 1772 5566
rect 1798 5562 1802 5566
rect 1826 5562 1830 5566
rect 2449 5562 2453 5566
rect 2479 5562 2483 5566
rect 2507 5562 2511 5566
rect 2581 5562 2585 5566
rect 2611 5562 2615 5566
rect 2639 5562 2643 5566
rect 2713 5562 2717 5566
rect 2743 5562 2747 5566
rect 2771 5562 2775 5566
rect 1065 5509 1069 5513
rect 1176 5509 1180 5513
rect 1200 5509 1204 5513
rect 1326 5509 1330 5513
rect 1361 5509 1365 5513
rect 2010 5509 2014 5513
rect 2121 5509 2125 5513
rect 2145 5509 2149 5513
rect 2271 5509 2275 5513
rect 2306 5509 2310 5513
rect 1682 5418 1686 5422
rect 1731 5418 1735 5422
rect 1785 5418 1789 5422
rect 1809 5418 1813 5422
rect 1831 5418 1835 5422
rect 951 5377 955 5381
rect 1005 5377 1009 5381
rect 1041 5377 1045 5381
rect 1095 5377 1099 5381
rect 1119 5377 1126 5381
rect 1176 5377 1180 5381
rect 1200 5377 1204 5381
rect 1326 5377 1330 5381
rect 1361 5377 1365 5381
rect 1896 5377 1900 5381
rect 1950 5377 1954 5381
rect 1986 5377 1990 5381
rect 2040 5377 2044 5381
rect 2064 5377 2071 5381
rect 2121 5377 2125 5381
rect 2145 5377 2149 5381
rect 2271 5377 2275 5381
rect 2306 5377 2310 5381
rect 4479 5313 4483 5317
rect 4489 5313 4493 5317
rect 4499 5313 4503 5317
rect 4509 5313 4513 5317
rect 4479 5308 4483 5312
rect 4489 5308 4493 5312
rect 4499 5308 4503 5312
rect 4509 5308 4513 5312
rect 4479 5303 4483 5307
rect 4489 5303 4493 5307
rect 4499 5303 4503 5307
rect 4509 5303 4513 5307
rect 4479 5298 4483 5302
rect 4489 5298 4493 5302
rect 4499 5298 4503 5302
rect 4509 5298 4513 5302
rect 1588 5288 1592 5292
rect 1731 5288 1735 5292
rect 1785 5288 1789 5292
rect 1809 5288 1813 5292
rect 659 5269 663 5273
rect 669 5269 673 5273
rect 679 5269 683 5273
rect 689 5269 693 5273
rect 659 5264 663 5268
rect 669 5264 673 5268
rect 679 5264 683 5268
rect 689 5264 693 5268
rect 659 5259 663 5263
rect 669 5259 673 5263
rect 679 5259 683 5263
rect 689 5259 693 5263
rect 659 5254 663 5258
rect 669 5254 673 5258
rect 679 5254 683 5258
rect 689 5254 693 5258
rect 1071 5245 1075 5249
rect 1095 5245 1099 5249
rect 1122 5245 1126 5249
rect 1176 5245 1180 5249
rect 1200 5245 1204 5249
rect 1326 5245 1330 5249
rect 1361 5245 1365 5249
rect 2016 5245 2020 5249
rect 2040 5245 2044 5249
rect 2067 5245 2071 5249
rect 2121 5245 2125 5249
rect 2145 5245 2149 5249
rect 2271 5245 2275 5249
rect 2306 5245 2310 5249
rect 1639 5162 1643 5166
rect 1667 5162 1671 5166
rect 1697 5162 1701 5166
rect 2584 5162 2588 5166
rect 2612 5162 2616 5166
rect 2642 5162 2646 5166
rect 1041 5113 1045 5117
rect 1095 5113 1099 5117
rect 1119 5113 1126 5117
rect 1176 5113 1180 5117
rect 1200 5113 1204 5117
rect 1326 5113 1330 5117
rect 1361 5113 1365 5117
rect 1986 5113 1990 5117
rect 2040 5113 2044 5117
rect 2064 5113 2071 5117
rect 2121 5113 2125 5117
rect 2145 5113 2149 5117
rect 2271 5113 2275 5117
rect 2306 5113 2310 5117
rect 1636 5060 1640 5064
rect 1666 5060 1670 5064
rect 1694 5060 1698 5064
rect 2581 5060 2585 5064
rect 2611 5060 2615 5064
rect 2639 5060 2643 5064
rect 888 5027 892 5031
rect 918 5027 922 5031
rect 946 5027 950 5031
rect 1020 5027 1024 5031
rect 1050 5027 1054 5031
rect 1078 5027 1082 5031
rect 1152 5027 1156 5031
rect 1182 5027 1186 5031
rect 1210 5027 1214 5031
rect 1284 5027 1288 5031
rect 1314 5027 1318 5031
rect 1342 5027 1346 5031
rect 1833 5027 1837 5031
rect 1863 5027 1867 5031
rect 1891 5027 1895 5031
rect 1965 5027 1969 5031
rect 1995 5027 1999 5031
rect 2023 5027 2027 5031
rect 2097 5027 2101 5031
rect 2127 5027 2131 5031
rect 2155 5027 2159 5031
rect 2229 5027 2233 5031
rect 2259 5027 2263 5031
rect 2287 5027 2291 5031
rect 4479 5004 4483 5008
rect 4489 5004 4493 5008
rect 4499 5004 4503 5008
rect 4509 5004 4513 5008
rect 4479 4999 4483 5003
rect 4489 4999 4493 5003
rect 4499 4999 4503 5003
rect 4509 4999 4513 5003
rect 4479 4994 4483 4998
rect 4489 4994 4493 4998
rect 4499 4994 4503 4998
rect 4509 4994 4513 4998
rect 4479 4989 4483 4993
rect 4489 4989 4493 4993
rect 4499 4989 4503 4993
rect 4509 4989 4513 4993
rect 659 4868 663 4872
rect 669 4868 673 4872
rect 679 4868 683 4872
rect 689 4868 693 4872
rect 659 4863 663 4867
rect 669 4863 673 4867
rect 679 4863 683 4867
rect 689 4863 693 4867
rect 659 4858 663 4862
rect 669 4858 673 4862
rect 679 4858 683 4862
rect 689 4858 693 4862
rect 659 4853 663 4857
rect 669 4853 673 4857
rect 679 4853 683 4857
rect 689 4853 693 4857
rect 659 4839 663 4843
rect 669 4839 673 4843
rect 679 4839 683 4843
rect 689 4839 693 4843
rect 659 4834 663 4838
rect 669 4834 673 4838
rect 679 4834 683 4838
rect 689 4834 693 4838
rect 659 4829 663 4833
rect 669 4829 673 4833
rect 679 4829 683 4833
rect 689 4829 693 4833
rect 659 4824 663 4828
rect 669 4824 673 4828
rect 679 4824 683 4828
rect 689 4824 693 4828
rect 659 4810 663 4814
rect 669 4810 673 4814
rect 679 4810 683 4814
rect 689 4810 693 4814
rect 659 4805 663 4809
rect 669 4805 673 4809
rect 679 4805 683 4809
rect 689 4805 693 4809
rect 659 4800 663 4804
rect 669 4800 673 4804
rect 679 4800 683 4804
rect 689 4800 693 4804
rect 659 4795 663 4799
rect 669 4795 673 4799
rect 679 4795 683 4799
rect 689 4795 693 4799
rect 659 4781 663 4785
rect 669 4781 673 4785
rect 679 4781 683 4785
rect 689 4781 693 4785
rect 659 4776 663 4780
rect 669 4776 673 4780
rect 679 4776 683 4780
rect 689 4776 693 4780
rect 659 4771 663 4775
rect 669 4771 673 4775
rect 679 4771 683 4775
rect 689 4771 693 4775
rect 659 4766 663 4770
rect 669 4766 673 4770
rect 679 4766 683 4770
rect 689 4766 693 4770
rect 659 4752 663 4756
rect 669 4752 673 4756
rect 679 4752 683 4756
rect 689 4752 693 4756
rect 659 4747 663 4751
rect 669 4747 673 4751
rect 679 4747 683 4751
rect 689 4747 693 4751
rect 659 4742 663 4746
rect 669 4742 673 4746
rect 679 4742 683 4746
rect 689 4742 693 4746
rect 659 4737 663 4741
rect 669 4737 673 4741
rect 679 4737 683 4741
rect 689 4737 693 4741
rect 4479 4811 4483 4815
rect 4489 4811 4493 4815
rect 4499 4811 4503 4815
rect 4509 4811 4513 4815
rect 4479 4806 4483 4810
rect 4489 4806 4493 4810
rect 4499 4806 4503 4810
rect 4509 4806 4513 4810
rect 4479 4801 4483 4805
rect 4489 4801 4493 4805
rect 4499 4801 4503 4805
rect 4509 4801 4513 4805
rect 4479 4796 4483 4800
rect 4489 4796 4493 4800
rect 4499 4796 4503 4800
rect 4509 4796 4513 4800
rect 4479 4785 4483 4789
rect 4489 4785 4493 4789
rect 4499 4785 4503 4789
rect 4509 4785 4513 4789
rect 4479 4780 4483 4784
rect 4489 4780 4493 4784
rect 4499 4780 4503 4784
rect 4509 4780 4513 4784
rect 4479 4775 4483 4779
rect 4489 4775 4493 4779
rect 4499 4775 4503 4779
rect 4509 4775 4513 4779
rect 4479 4770 4483 4774
rect 4489 4770 4493 4774
rect 4499 4770 4503 4774
rect 4509 4770 4513 4774
rect 4479 4759 4483 4763
rect 4489 4759 4493 4763
rect 4499 4759 4503 4763
rect 4509 4759 4513 4763
rect 4479 4754 4483 4758
rect 4489 4754 4493 4758
rect 4499 4754 4503 4758
rect 4509 4754 4513 4758
rect 4479 4749 4483 4753
rect 4489 4749 4493 4753
rect 4499 4749 4503 4753
rect 4509 4749 4513 4753
rect 4479 4744 4483 4748
rect 4489 4744 4493 4748
rect 4499 4744 4503 4748
rect 4509 4744 4513 4748
rect 4479 4733 4483 4737
rect 4489 4733 4493 4737
rect 4499 4733 4503 4737
rect 4509 4733 4513 4737
rect 4479 4728 4483 4732
rect 4489 4728 4493 4732
rect 4499 4728 4503 4732
rect 4509 4728 4513 4732
rect 4479 4723 4483 4727
rect 4489 4723 4493 4727
rect 4499 4723 4503 4727
rect 4509 4723 4513 4727
rect 4479 4718 4483 4722
rect 4489 4718 4493 4722
rect 4499 4718 4503 4722
rect 4509 4718 4513 4722
rect 4479 4707 4483 4711
rect 4489 4707 4493 4711
rect 4499 4707 4503 4711
rect 4509 4707 4513 4711
rect 4479 4702 4483 4706
rect 4489 4702 4493 4706
rect 4499 4702 4503 4706
rect 4509 4702 4513 4706
rect 4479 4697 4483 4701
rect 4489 4697 4493 4701
rect 4499 4697 4503 4701
rect 4509 4697 4513 4701
rect 4479 4692 4483 4696
rect 4489 4692 4493 4696
rect 4499 4692 4503 4696
rect 4509 4692 4513 4696
rect 757 4624 761 4628
rect 762 4624 766 4628
rect 767 4624 771 4628
rect 772 4624 776 4628
rect 783 4624 787 4628
rect 788 4624 792 4628
rect 793 4624 797 4628
rect 798 4624 802 4628
rect 809 4624 813 4628
rect 814 4624 818 4628
rect 819 4624 823 4628
rect 824 4624 828 4628
rect 835 4624 839 4628
rect 840 4624 844 4628
rect 845 4624 849 4628
rect 850 4624 854 4628
rect 861 4624 865 4628
rect 866 4624 870 4628
rect 871 4624 875 4628
rect 876 4624 880 4628
rect 1053 4624 1057 4628
rect 1058 4624 1062 4628
rect 1063 4624 1067 4628
rect 1068 4624 1072 4628
rect 1362 4624 1366 4628
rect 1367 4624 1371 4628
rect 1372 4624 1376 4628
rect 1377 4624 1381 4628
rect 1671 4624 1675 4628
rect 1676 4624 1680 4628
rect 1681 4624 1685 4628
rect 1686 4624 1690 4628
rect 1980 4624 1984 4628
rect 1985 4624 1989 4628
rect 1990 4624 1994 4628
rect 1995 4624 1999 4628
rect 2289 4624 2293 4628
rect 2294 4624 2298 4628
rect 2299 4624 2303 4628
rect 2304 4624 2308 4628
rect 2598 4624 2602 4628
rect 2603 4624 2607 4628
rect 2608 4624 2612 4628
rect 2613 4624 2617 4628
rect 2907 4624 2911 4628
rect 2912 4624 2916 4628
rect 2917 4624 2921 4628
rect 2922 4624 2926 4628
rect 3216 4624 3220 4628
rect 3221 4624 3225 4628
rect 3226 4624 3230 4628
rect 3231 4624 3235 4628
rect 3525 4624 3529 4628
rect 3530 4624 3534 4628
rect 3535 4624 3539 4628
rect 3540 4624 3544 4628
rect 3834 4624 3838 4628
rect 3839 4624 3843 4628
rect 3844 4624 3848 4628
rect 3849 4624 3853 4628
rect 4235 4624 4239 4628
rect 4240 4624 4244 4628
rect 4245 4624 4249 4628
rect 4250 4624 4254 4628
rect 4264 4624 4268 4628
rect 4269 4624 4273 4628
rect 4274 4624 4278 4628
rect 4279 4624 4283 4628
rect 4293 4624 4297 4628
rect 4298 4624 4302 4628
rect 4303 4624 4307 4628
rect 4308 4624 4312 4628
rect 4322 4624 4326 4628
rect 4327 4624 4331 4628
rect 4332 4624 4336 4628
rect 4337 4624 4341 4628
rect 4351 4624 4355 4628
rect 4356 4624 4360 4628
rect 4361 4624 4365 4628
rect 4366 4624 4370 4628
rect 757 4614 761 4618
rect 762 4614 766 4618
rect 767 4614 771 4618
rect 772 4614 776 4618
rect 783 4614 787 4618
rect 788 4614 792 4618
rect 793 4614 797 4618
rect 798 4614 802 4618
rect 809 4614 813 4618
rect 814 4614 818 4618
rect 819 4614 823 4618
rect 824 4614 828 4618
rect 835 4614 839 4618
rect 840 4614 844 4618
rect 845 4614 849 4618
rect 850 4614 854 4618
rect 861 4614 865 4618
rect 866 4614 870 4618
rect 871 4614 875 4618
rect 876 4614 880 4618
rect 1053 4614 1057 4618
rect 1058 4614 1062 4618
rect 1063 4614 1067 4618
rect 1068 4614 1072 4618
rect 1362 4614 1366 4618
rect 1367 4614 1371 4618
rect 1372 4614 1376 4618
rect 1377 4614 1381 4618
rect 1671 4614 1675 4618
rect 1676 4614 1680 4618
rect 1681 4614 1685 4618
rect 1686 4614 1690 4618
rect 1980 4614 1984 4618
rect 1985 4614 1989 4618
rect 1990 4614 1994 4618
rect 1995 4614 1999 4618
rect 2289 4614 2293 4618
rect 2294 4614 2298 4618
rect 2299 4614 2303 4618
rect 2304 4614 2308 4618
rect 2598 4614 2602 4618
rect 2603 4614 2607 4618
rect 2608 4614 2612 4618
rect 2613 4614 2617 4618
rect 2907 4614 2911 4618
rect 2912 4614 2916 4618
rect 2917 4614 2921 4618
rect 2922 4614 2926 4618
rect 3216 4614 3220 4618
rect 3221 4614 3225 4618
rect 3226 4614 3230 4618
rect 3231 4614 3235 4618
rect 3525 4614 3529 4618
rect 3530 4614 3534 4618
rect 3535 4614 3539 4618
rect 3540 4614 3544 4618
rect 3834 4614 3838 4618
rect 3839 4614 3843 4618
rect 3844 4614 3848 4618
rect 3849 4614 3853 4618
rect 4235 4614 4239 4618
rect 4240 4614 4244 4618
rect 4245 4614 4249 4618
rect 4250 4614 4254 4618
rect 4264 4614 4268 4618
rect 4269 4614 4273 4618
rect 4274 4614 4278 4618
rect 4279 4614 4283 4618
rect 4293 4614 4297 4618
rect 4298 4614 4302 4618
rect 4303 4614 4307 4618
rect 4308 4614 4312 4618
rect 4322 4614 4326 4618
rect 4327 4614 4331 4618
rect 4332 4614 4336 4618
rect 4337 4614 4341 4618
rect 4351 4614 4355 4618
rect 4356 4614 4360 4618
rect 4361 4614 4365 4618
rect 4366 4614 4370 4618
rect 757 4604 761 4608
rect 762 4604 766 4608
rect 767 4604 771 4608
rect 772 4604 776 4608
rect 783 4604 787 4608
rect 788 4604 792 4608
rect 793 4604 797 4608
rect 798 4604 802 4608
rect 809 4604 813 4608
rect 814 4604 818 4608
rect 819 4604 823 4608
rect 824 4604 828 4608
rect 835 4604 839 4608
rect 840 4604 844 4608
rect 845 4604 849 4608
rect 850 4604 854 4608
rect 861 4604 865 4608
rect 866 4604 870 4608
rect 871 4604 875 4608
rect 876 4604 880 4608
rect 1053 4604 1057 4608
rect 1058 4604 1062 4608
rect 1063 4604 1067 4608
rect 1068 4604 1072 4608
rect 1362 4604 1366 4608
rect 1367 4604 1371 4608
rect 1372 4604 1376 4608
rect 1377 4604 1381 4608
rect 1671 4604 1675 4608
rect 1676 4604 1680 4608
rect 1681 4604 1685 4608
rect 1686 4604 1690 4608
rect 1980 4604 1984 4608
rect 1985 4604 1989 4608
rect 1990 4604 1994 4608
rect 1995 4604 1999 4608
rect 2289 4604 2293 4608
rect 2294 4604 2298 4608
rect 2299 4604 2303 4608
rect 2304 4604 2308 4608
rect 2598 4604 2602 4608
rect 2603 4604 2607 4608
rect 2608 4604 2612 4608
rect 2613 4604 2617 4608
rect 2907 4604 2911 4608
rect 2912 4604 2916 4608
rect 2917 4604 2921 4608
rect 2922 4604 2926 4608
rect 3216 4604 3220 4608
rect 3221 4604 3225 4608
rect 3226 4604 3230 4608
rect 3231 4604 3235 4608
rect 3525 4604 3529 4608
rect 3530 4604 3534 4608
rect 3535 4604 3539 4608
rect 3540 4604 3544 4608
rect 3834 4604 3838 4608
rect 3839 4604 3843 4608
rect 3844 4604 3848 4608
rect 3849 4604 3853 4608
rect 4235 4604 4239 4608
rect 4240 4604 4244 4608
rect 4245 4604 4249 4608
rect 4250 4604 4254 4608
rect 4264 4604 4268 4608
rect 4269 4604 4273 4608
rect 4274 4604 4278 4608
rect 4279 4604 4283 4608
rect 4293 4604 4297 4608
rect 4298 4604 4302 4608
rect 4303 4604 4307 4608
rect 4308 4604 4312 4608
rect 4322 4604 4326 4608
rect 4327 4604 4331 4608
rect 4332 4604 4336 4608
rect 4337 4604 4341 4608
rect 4351 4604 4355 4608
rect 4356 4604 4360 4608
rect 4361 4604 4365 4608
rect 4366 4604 4370 4608
rect 757 4594 761 4598
rect 762 4594 766 4598
rect 767 4594 771 4598
rect 772 4594 776 4598
rect 783 4594 787 4598
rect 788 4594 792 4598
rect 793 4594 797 4598
rect 798 4594 802 4598
rect 809 4594 813 4598
rect 814 4594 818 4598
rect 819 4594 823 4598
rect 824 4594 828 4598
rect 835 4594 839 4598
rect 840 4594 844 4598
rect 845 4594 849 4598
rect 850 4594 854 4598
rect 861 4594 865 4598
rect 866 4594 870 4598
rect 871 4594 875 4598
rect 876 4594 880 4598
rect 1053 4594 1057 4598
rect 1058 4594 1062 4598
rect 1063 4594 1067 4598
rect 1068 4594 1072 4598
rect 1362 4594 1366 4598
rect 1367 4594 1371 4598
rect 1372 4594 1376 4598
rect 1377 4594 1381 4598
rect 1671 4594 1675 4598
rect 1676 4594 1680 4598
rect 1681 4594 1685 4598
rect 1686 4594 1690 4598
rect 1980 4594 1984 4598
rect 1985 4594 1989 4598
rect 1990 4594 1994 4598
rect 1995 4594 1999 4598
rect 2289 4594 2293 4598
rect 2294 4594 2298 4598
rect 2299 4594 2303 4598
rect 2304 4594 2308 4598
rect 2598 4594 2602 4598
rect 2603 4594 2607 4598
rect 2608 4594 2612 4598
rect 2613 4594 2617 4598
rect 2907 4594 2911 4598
rect 2912 4594 2916 4598
rect 2917 4594 2921 4598
rect 2922 4594 2926 4598
rect 3216 4594 3220 4598
rect 3221 4594 3225 4598
rect 3226 4594 3230 4598
rect 3231 4594 3235 4598
rect 3525 4594 3529 4598
rect 3530 4594 3534 4598
rect 3535 4594 3539 4598
rect 3540 4594 3544 4598
rect 3834 4594 3838 4598
rect 3839 4594 3843 4598
rect 3844 4594 3848 4598
rect 3849 4594 3853 4598
rect 4235 4594 4239 4598
rect 4240 4594 4244 4598
rect 4245 4594 4249 4598
rect 4250 4594 4254 4598
rect 4264 4594 4268 4598
rect 4269 4594 4273 4598
rect 4274 4594 4278 4598
rect 4279 4594 4283 4598
rect 4293 4594 4297 4598
rect 4298 4594 4302 4598
rect 4303 4594 4307 4598
rect 4308 4594 4312 4598
rect 4322 4594 4326 4598
rect 4327 4594 4331 4598
rect 4332 4594 4336 4598
rect 4337 4594 4341 4598
rect 4351 4594 4355 4598
rect 4356 4594 4360 4598
rect 4361 4594 4365 4598
rect 4366 4594 4370 4598
rect 4627 7975 4631 8015
rect 4666 7975 4670 8034
rect 4709 7975 4713 8034
rect 4750 7975 4754 8034
rect 4645 7473 4649 7477
rect 4652 7473 4656 7477
rect 4657 7473 4661 7477
rect 4662 7473 4666 7477
rect 4667 7473 4671 7477
rect 4672 7473 4676 7477
rect 4677 7473 4681 7477
rect 4682 7473 4686 7477
rect 4687 7473 4691 7477
rect 4692 7473 4696 7477
rect 4697 7473 4701 7477
rect 4702 7473 4706 7477
rect 4707 7473 4711 7477
rect 4712 7473 4716 7477
rect 4717 7473 4721 7477
rect 4722 7473 4726 7477
rect 4727 7473 4731 7477
rect 4732 7473 4736 7477
rect 4737 7473 4741 7477
rect 4742 7473 4746 7477
rect 4747 7473 4751 7477
rect 4754 7473 4758 7477
rect 4645 7466 4649 7470
rect 4754 7466 4758 7470
rect 4645 7461 4649 7465
rect 4645 7456 4649 7460
rect 4645 7451 4649 7455
rect 4645 7446 4649 7450
rect 4645 7441 4649 7445
rect 4645 7436 4649 7440
rect 4645 7431 4649 7435
rect 4645 7426 4649 7430
rect 4645 7421 4649 7425
rect 4754 7461 4758 7465
rect 4754 7456 4758 7460
rect 4754 7451 4758 7455
rect 4754 7446 4758 7450
rect 4754 7441 4758 7445
rect 4754 7436 4758 7440
rect 4754 7431 4758 7435
rect 4754 7426 4758 7430
rect 4754 7421 4758 7425
rect 4645 7416 4649 7420
rect 4754 7416 4758 7420
rect 4645 7409 4649 7413
rect 4652 7409 4656 7413
rect 4657 7409 4661 7413
rect 4662 7409 4666 7413
rect 4667 7409 4671 7413
rect 4672 7409 4676 7413
rect 4677 7409 4681 7413
rect 4682 7409 4686 7413
rect 4687 7409 4691 7413
rect 4692 7409 4696 7413
rect 4697 7409 4701 7413
rect 4702 7409 4706 7413
rect 4707 7409 4711 7413
rect 4712 7409 4716 7413
rect 4717 7409 4721 7413
rect 4722 7409 4726 7413
rect 4727 7409 4731 7413
rect 4732 7409 4736 7413
rect 4737 7409 4741 7413
rect 4742 7409 4746 7413
rect 4747 7409 4751 7413
rect 4754 7409 4758 7413
rect 4632 7326 4636 7330
rect 4637 7326 4641 7330
rect 4642 7326 4646 7330
rect 4647 7326 4651 7330
rect 4652 7326 4656 7330
rect 4657 7326 4661 7330
rect 4662 7326 4666 7330
rect 4667 7326 4671 7330
rect 4672 7326 4676 7330
rect 4677 7326 4681 7330
rect 4682 7326 4686 7330
rect 4687 7326 4691 7330
rect 4692 7326 4696 7330
rect 4697 7326 4701 7330
rect 4702 7326 4706 7330
rect 4707 7326 4711 7330
rect 4712 7326 4716 7330
rect 4717 7326 4721 7330
rect 4722 7326 4726 7330
rect 4727 7326 4731 7330
rect 4732 7326 4736 7330
rect 4737 7326 4741 7330
rect 4742 7326 4746 7330
rect 4747 7326 4751 7330
rect 4752 7326 4756 7330
rect 4757 7326 4761 7330
rect 4762 7326 4766 7330
rect 4767 7326 4771 7330
rect 4632 7321 4636 7325
rect 4632 7316 4636 7320
rect 4767 7321 4771 7325
rect 4632 7311 4636 7315
rect 4632 7306 4636 7310
rect 4632 7301 4636 7305
rect 4632 7296 4636 7300
rect 4632 7291 4636 7295
rect 4632 7286 4636 7290
rect 4632 7281 4636 7285
rect 4632 7276 4636 7280
rect 4632 7271 4636 7275
rect 4632 7266 4636 7270
rect 4632 7261 4636 7265
rect 4632 7256 4636 7260
rect 4632 7251 4636 7255
rect 4632 7246 4636 7250
rect 4767 7316 4771 7320
rect 4767 7311 4771 7315
rect 4767 7306 4771 7310
rect 4767 7301 4771 7305
rect 4767 7296 4771 7300
rect 4767 7291 4771 7295
rect 4767 7286 4771 7290
rect 4767 7281 4771 7285
rect 4767 7276 4771 7280
rect 4767 7271 4771 7275
rect 4767 7266 4771 7270
rect 4767 7261 4771 7265
rect 4767 7256 4771 7260
rect 4767 7251 4771 7255
rect 4632 7241 4636 7245
rect 4767 7246 4771 7250
rect 4767 7241 4771 7245
rect 4632 7236 4636 7240
rect 4637 7236 4641 7240
rect 4642 7236 4646 7240
rect 4647 7236 4651 7240
rect 4652 7236 4656 7240
rect 4657 7236 4661 7240
rect 4662 7236 4666 7240
rect 4667 7236 4671 7240
rect 4672 7236 4676 7240
rect 4677 7236 4681 7240
rect 4682 7236 4686 7240
rect 4687 7236 4691 7240
rect 4692 7236 4696 7240
rect 4697 7236 4701 7240
rect 4702 7236 4706 7240
rect 4707 7236 4711 7240
rect 4712 7236 4716 7240
rect 4717 7236 4721 7240
rect 4722 7236 4726 7240
rect 4727 7236 4731 7240
rect 4732 7236 4736 7240
rect 4737 7236 4741 7240
rect 4742 7236 4746 7240
rect 4747 7236 4751 7240
rect 4752 7236 4756 7240
rect 4757 7236 4761 7240
rect 4762 7236 4766 7240
rect 4767 7236 4771 7240
rect 1074 4471 1078 4475
rect 1079 4471 1083 4475
rect 1084 4471 1088 4475
rect 1089 4471 1093 4475
rect 1094 4471 1098 4475
rect 1099 4471 1103 4475
rect 1104 4471 1108 4475
rect 1109 4471 1113 4475
rect 1114 4471 1118 4475
rect 1119 4471 1123 4475
rect 1124 4471 1128 4475
rect 1129 4471 1133 4475
rect 1134 4471 1138 4475
rect 1139 4471 1143 4475
rect 1144 4471 1148 4475
rect 1149 4471 1153 4475
rect 1154 4471 1158 4475
rect 1159 4471 1163 4475
rect 1164 4471 1168 4475
rect 1074 4466 1078 4470
rect 1074 4461 1078 4465
rect 1164 4466 1168 4470
rect 1074 4456 1078 4460
rect 1074 4451 1078 4455
rect 1074 4446 1078 4450
rect 1074 4441 1078 4445
rect 1074 4436 1078 4440
rect 1074 4431 1078 4435
rect 1074 4426 1078 4430
rect 1074 4421 1078 4425
rect 1074 4416 1078 4420
rect 1074 4411 1078 4415
rect 1074 4406 1078 4410
rect 1074 4401 1078 4405
rect 1074 4396 1078 4400
rect 1074 4391 1078 4395
rect 1074 4386 1078 4390
rect 1074 4381 1078 4385
rect 1074 4376 1078 4380
rect 1074 4371 1078 4375
rect 1074 4366 1078 4370
rect 1074 4361 1078 4365
rect 1074 4356 1078 4360
rect 1074 4351 1078 4355
rect 1074 4346 1078 4350
rect 1164 4461 1168 4465
rect 1164 4456 1168 4460
rect 1164 4451 1168 4455
rect 1164 4446 1168 4450
rect 1164 4441 1168 4445
rect 1164 4436 1168 4440
rect 1164 4431 1168 4435
rect 1164 4426 1168 4430
rect 1164 4421 1168 4425
rect 1164 4416 1168 4420
rect 1164 4411 1168 4415
rect 1164 4406 1168 4410
rect 1164 4401 1168 4405
rect 1164 4396 1168 4400
rect 1164 4391 1168 4395
rect 1164 4386 1168 4390
rect 1164 4381 1168 4385
rect 1164 4376 1168 4380
rect 1164 4371 1168 4375
rect 1164 4366 1168 4370
rect 1164 4361 1168 4365
rect 1164 4356 1168 4360
rect 1164 4351 1168 4355
rect 1074 4341 1078 4345
rect 1164 4346 1168 4350
rect 1164 4341 1168 4345
rect 1074 4336 1078 4340
rect 1079 4336 1083 4340
rect 1084 4336 1088 4340
rect 1089 4336 1093 4340
rect 1094 4336 1098 4340
rect 1099 4336 1103 4340
rect 1104 4336 1108 4340
rect 1109 4336 1113 4340
rect 1114 4336 1118 4340
rect 1119 4336 1123 4340
rect 1124 4336 1128 4340
rect 1129 4336 1133 4340
rect 1134 4336 1138 4340
rect 1139 4336 1143 4340
rect 1144 4336 1148 4340
rect 1149 4336 1153 4340
rect 1154 4336 1158 4340
rect 1159 4336 1163 4340
rect 1164 4336 1168 4340
rect 1247 4458 1251 4462
rect 1254 4458 1258 4462
rect 1259 4458 1263 4462
rect 1264 4458 1268 4462
rect 1269 4458 1273 4462
rect 1274 4458 1278 4462
rect 1279 4458 1283 4462
rect 1284 4458 1288 4462
rect 1289 4458 1293 4462
rect 1294 4458 1298 4462
rect 1299 4458 1303 4462
rect 1304 4458 1308 4462
rect 1311 4458 1315 4462
rect 1247 4451 1251 4455
rect 1311 4451 1315 4455
rect 1247 4446 1251 4450
rect 1247 4441 1251 4445
rect 1247 4436 1251 4440
rect 1247 4431 1251 4435
rect 1247 4426 1251 4430
rect 1247 4421 1251 4425
rect 1247 4416 1251 4420
rect 1247 4411 1251 4415
rect 1247 4406 1251 4410
rect 1247 4401 1251 4405
rect 1247 4396 1251 4400
rect 1247 4391 1251 4395
rect 1247 4386 1251 4390
rect 1247 4381 1251 4385
rect 1247 4376 1251 4380
rect 1247 4371 1251 4375
rect 1247 4366 1251 4370
rect 1247 4361 1251 4365
rect 1311 4446 1315 4450
rect 1311 4441 1315 4445
rect 1311 4436 1315 4440
rect 1311 4431 1315 4435
rect 1311 4426 1315 4430
rect 1311 4421 1315 4425
rect 1311 4416 1315 4420
rect 1311 4411 1315 4415
rect 1311 4406 1315 4410
rect 1311 4401 1315 4405
rect 1311 4396 1315 4400
rect 1311 4391 1315 4395
rect 1311 4386 1315 4390
rect 1311 4381 1315 4385
rect 1311 4376 1315 4380
rect 1311 4371 1315 4375
rect 1311 4366 1315 4370
rect 1311 4361 1315 4365
rect 1247 4356 1251 4360
rect 1311 4356 1315 4360
rect 1247 4349 1251 4353
rect 1254 4349 1258 4353
rect 1259 4349 1263 4353
rect 1264 4349 1268 4353
rect 1269 4349 1273 4353
rect 1274 4349 1278 4353
rect 1279 4349 1283 4353
rect 1284 4349 1288 4353
rect 1289 4349 1293 4353
rect 1294 4349 1298 4353
rect 1299 4349 1303 4353
rect 1304 4349 1308 4353
rect 1311 4349 1315 4353
rect 1383 4471 1387 4475
rect 1388 4471 1392 4475
rect 1393 4471 1397 4475
rect 1398 4471 1402 4475
rect 1403 4471 1407 4475
rect 1408 4471 1412 4475
rect 1413 4471 1417 4475
rect 1418 4471 1422 4475
rect 1423 4471 1427 4475
rect 1428 4471 1432 4475
rect 1433 4471 1437 4475
rect 1438 4471 1442 4475
rect 1443 4471 1447 4475
rect 1448 4471 1452 4475
rect 1453 4471 1457 4475
rect 1458 4471 1462 4475
rect 1463 4471 1467 4475
rect 1468 4471 1472 4475
rect 1473 4471 1477 4475
rect 1383 4466 1387 4470
rect 1383 4461 1387 4465
rect 1473 4466 1477 4470
rect 1383 4456 1387 4460
rect 1383 4451 1387 4455
rect 1383 4446 1387 4450
rect 1383 4441 1387 4445
rect 1383 4436 1387 4440
rect 1383 4431 1387 4435
rect 1383 4426 1387 4430
rect 1383 4421 1387 4425
rect 1383 4416 1387 4420
rect 1383 4411 1387 4415
rect 1383 4406 1387 4410
rect 1383 4401 1387 4405
rect 1383 4396 1387 4400
rect 1383 4391 1387 4395
rect 1383 4386 1387 4390
rect 1383 4381 1387 4385
rect 1383 4376 1387 4380
rect 1383 4371 1387 4375
rect 1383 4366 1387 4370
rect 1383 4361 1387 4365
rect 1383 4356 1387 4360
rect 1383 4351 1387 4355
rect 1383 4346 1387 4350
rect 1473 4461 1477 4465
rect 1473 4456 1477 4460
rect 1473 4451 1477 4455
rect 1473 4446 1477 4450
rect 1473 4441 1477 4445
rect 1473 4436 1477 4440
rect 1473 4431 1477 4435
rect 1473 4426 1477 4430
rect 1473 4421 1477 4425
rect 1473 4416 1477 4420
rect 1473 4411 1477 4415
rect 1473 4406 1477 4410
rect 1473 4401 1477 4405
rect 1473 4396 1477 4400
rect 1473 4391 1477 4395
rect 1473 4386 1477 4390
rect 1473 4381 1477 4385
rect 1473 4376 1477 4380
rect 1473 4371 1477 4375
rect 1473 4366 1477 4370
rect 1473 4361 1477 4365
rect 1473 4356 1477 4360
rect 1473 4351 1477 4355
rect 1383 4341 1387 4345
rect 1473 4346 1477 4350
rect 1473 4341 1477 4345
rect 1383 4336 1387 4340
rect 1388 4336 1392 4340
rect 1393 4336 1397 4340
rect 1398 4336 1402 4340
rect 1403 4336 1407 4340
rect 1408 4336 1412 4340
rect 1413 4336 1417 4340
rect 1418 4336 1422 4340
rect 1423 4336 1427 4340
rect 1428 4336 1432 4340
rect 1433 4336 1437 4340
rect 1438 4336 1442 4340
rect 1443 4336 1447 4340
rect 1448 4336 1452 4340
rect 1453 4336 1457 4340
rect 1458 4336 1462 4340
rect 1463 4336 1467 4340
rect 1468 4336 1472 4340
rect 1473 4336 1477 4340
rect 1556 4458 1560 4462
rect 1563 4458 1567 4462
rect 1568 4458 1572 4462
rect 1573 4458 1577 4462
rect 1578 4458 1582 4462
rect 1583 4458 1587 4462
rect 1588 4458 1592 4462
rect 1593 4458 1597 4462
rect 1598 4458 1602 4462
rect 1603 4458 1607 4462
rect 1608 4458 1612 4462
rect 1613 4458 1617 4462
rect 1620 4458 1624 4462
rect 1556 4451 1560 4455
rect 1620 4451 1624 4455
rect 1556 4446 1560 4450
rect 1556 4441 1560 4445
rect 1556 4436 1560 4440
rect 1556 4431 1560 4435
rect 1556 4426 1560 4430
rect 1556 4421 1560 4425
rect 1556 4416 1560 4420
rect 1556 4411 1560 4415
rect 1556 4406 1560 4410
rect 1556 4401 1560 4405
rect 1556 4396 1560 4400
rect 1556 4391 1560 4395
rect 1556 4386 1560 4390
rect 1556 4381 1560 4385
rect 1556 4376 1560 4380
rect 1556 4371 1560 4375
rect 1556 4366 1560 4370
rect 1556 4361 1560 4365
rect 1620 4446 1624 4450
rect 1620 4441 1624 4445
rect 1620 4436 1624 4440
rect 1620 4431 1624 4435
rect 1620 4426 1624 4430
rect 1620 4421 1624 4425
rect 1620 4416 1624 4420
rect 1620 4411 1624 4415
rect 1620 4406 1624 4410
rect 1620 4401 1624 4405
rect 1620 4396 1624 4400
rect 1620 4391 1624 4395
rect 1620 4386 1624 4390
rect 1620 4381 1624 4385
rect 1620 4376 1624 4380
rect 1620 4371 1624 4375
rect 1620 4366 1624 4370
rect 1620 4361 1624 4365
rect 1556 4356 1560 4360
rect 1620 4356 1624 4360
rect 1556 4349 1560 4353
rect 1563 4349 1567 4353
rect 1568 4349 1572 4353
rect 1573 4349 1577 4353
rect 1578 4349 1582 4353
rect 1583 4349 1587 4353
rect 1588 4349 1592 4353
rect 1593 4349 1597 4353
rect 1598 4349 1602 4353
rect 1603 4349 1607 4353
rect 1608 4349 1612 4353
rect 1613 4349 1617 4353
rect 1620 4349 1624 4353
rect 1692 4471 1696 4475
rect 1697 4471 1701 4475
rect 1702 4471 1706 4475
rect 1707 4471 1711 4475
rect 1712 4471 1716 4475
rect 1717 4471 1721 4475
rect 1722 4471 1726 4475
rect 1727 4471 1731 4475
rect 1732 4471 1736 4475
rect 1737 4471 1741 4475
rect 1742 4471 1746 4475
rect 1747 4471 1751 4475
rect 1752 4471 1756 4475
rect 1757 4471 1761 4475
rect 1762 4471 1766 4475
rect 1767 4471 1771 4475
rect 1772 4471 1776 4475
rect 1777 4471 1781 4475
rect 1782 4471 1786 4475
rect 1692 4466 1696 4470
rect 1692 4461 1696 4465
rect 1782 4466 1786 4470
rect 1692 4456 1696 4460
rect 1692 4451 1696 4455
rect 1692 4446 1696 4450
rect 1692 4441 1696 4445
rect 1692 4436 1696 4440
rect 1692 4431 1696 4435
rect 1692 4426 1696 4430
rect 1692 4421 1696 4425
rect 1692 4416 1696 4420
rect 1692 4411 1696 4415
rect 1692 4406 1696 4410
rect 1692 4401 1696 4405
rect 1692 4396 1696 4400
rect 1692 4391 1696 4395
rect 1692 4386 1696 4390
rect 1692 4381 1696 4385
rect 1692 4376 1696 4380
rect 1692 4371 1696 4375
rect 1692 4366 1696 4370
rect 1692 4361 1696 4365
rect 1692 4356 1696 4360
rect 1692 4351 1696 4355
rect 1692 4346 1696 4350
rect 1782 4461 1786 4465
rect 1782 4456 1786 4460
rect 1782 4451 1786 4455
rect 1782 4446 1786 4450
rect 1782 4441 1786 4445
rect 1782 4436 1786 4440
rect 1782 4431 1786 4435
rect 1782 4426 1786 4430
rect 1782 4421 1786 4425
rect 1782 4416 1786 4420
rect 1782 4411 1786 4415
rect 1782 4406 1786 4410
rect 1782 4401 1786 4405
rect 1782 4396 1786 4400
rect 1782 4391 1786 4395
rect 1782 4386 1786 4390
rect 1782 4381 1786 4385
rect 1782 4376 1786 4380
rect 1782 4371 1786 4375
rect 1782 4366 1786 4370
rect 1782 4361 1786 4365
rect 1782 4356 1786 4360
rect 1782 4351 1786 4355
rect 1692 4341 1696 4345
rect 1782 4346 1786 4350
rect 1782 4341 1786 4345
rect 1692 4336 1696 4340
rect 1697 4336 1701 4340
rect 1702 4336 1706 4340
rect 1707 4336 1711 4340
rect 1712 4336 1716 4340
rect 1717 4336 1721 4340
rect 1722 4336 1726 4340
rect 1727 4336 1731 4340
rect 1732 4336 1736 4340
rect 1737 4336 1741 4340
rect 1742 4336 1746 4340
rect 1747 4336 1751 4340
rect 1752 4336 1756 4340
rect 1757 4336 1761 4340
rect 1762 4336 1766 4340
rect 1767 4336 1771 4340
rect 1772 4336 1776 4340
rect 1777 4336 1781 4340
rect 1782 4336 1786 4340
rect 1865 4458 1869 4462
rect 1872 4458 1876 4462
rect 1877 4458 1881 4462
rect 1882 4458 1886 4462
rect 1887 4458 1891 4462
rect 1892 4458 1896 4462
rect 1897 4458 1901 4462
rect 1902 4458 1906 4462
rect 1907 4458 1911 4462
rect 1912 4458 1916 4462
rect 1917 4458 1921 4462
rect 1922 4458 1926 4462
rect 1929 4458 1933 4462
rect 1865 4451 1869 4455
rect 1929 4451 1933 4455
rect 1865 4446 1869 4450
rect 1865 4441 1869 4445
rect 1865 4436 1869 4440
rect 1865 4431 1869 4435
rect 1865 4426 1869 4430
rect 1865 4421 1869 4425
rect 1865 4416 1869 4420
rect 1865 4411 1869 4415
rect 1865 4406 1869 4410
rect 1865 4401 1869 4405
rect 1865 4396 1869 4400
rect 1865 4391 1869 4395
rect 1865 4386 1869 4390
rect 1865 4381 1869 4385
rect 1865 4376 1869 4380
rect 1865 4371 1869 4375
rect 1865 4366 1869 4370
rect 1865 4361 1869 4365
rect 1929 4446 1933 4450
rect 1929 4441 1933 4445
rect 1929 4436 1933 4440
rect 1929 4431 1933 4435
rect 1929 4426 1933 4430
rect 1929 4421 1933 4425
rect 1929 4416 1933 4420
rect 1929 4411 1933 4415
rect 1929 4406 1933 4410
rect 1929 4401 1933 4405
rect 1929 4396 1933 4400
rect 1929 4391 1933 4395
rect 1929 4386 1933 4390
rect 1929 4381 1933 4385
rect 1929 4376 1933 4380
rect 1929 4371 1933 4375
rect 1929 4366 1933 4370
rect 1929 4361 1933 4365
rect 1865 4356 1869 4360
rect 1929 4356 1933 4360
rect 1865 4349 1869 4353
rect 1872 4349 1876 4353
rect 1877 4349 1881 4353
rect 1882 4349 1886 4353
rect 1887 4349 1891 4353
rect 1892 4349 1896 4353
rect 1897 4349 1901 4353
rect 1902 4349 1906 4353
rect 1907 4349 1911 4353
rect 1912 4349 1916 4353
rect 1917 4349 1921 4353
rect 1922 4349 1926 4353
rect 1929 4349 1933 4353
rect 2001 4471 2005 4475
rect 2006 4471 2010 4475
rect 2011 4471 2015 4475
rect 2016 4471 2020 4475
rect 2021 4471 2025 4475
rect 2026 4471 2030 4475
rect 2031 4471 2035 4475
rect 2036 4471 2040 4475
rect 2041 4471 2045 4475
rect 2046 4471 2050 4475
rect 2051 4471 2055 4475
rect 2056 4471 2060 4475
rect 2061 4471 2065 4475
rect 2066 4471 2070 4475
rect 2071 4471 2075 4475
rect 2076 4471 2080 4475
rect 2081 4471 2085 4475
rect 2086 4471 2090 4475
rect 2091 4471 2095 4475
rect 2001 4466 2005 4470
rect 2001 4461 2005 4465
rect 2091 4466 2095 4470
rect 2001 4456 2005 4460
rect 2001 4451 2005 4455
rect 2001 4446 2005 4450
rect 2001 4441 2005 4445
rect 2001 4436 2005 4440
rect 2001 4431 2005 4435
rect 2001 4426 2005 4430
rect 2001 4421 2005 4425
rect 2001 4416 2005 4420
rect 2001 4411 2005 4415
rect 2001 4406 2005 4410
rect 2001 4401 2005 4405
rect 2001 4396 2005 4400
rect 2001 4391 2005 4395
rect 2001 4386 2005 4390
rect 2001 4381 2005 4385
rect 2001 4376 2005 4380
rect 2001 4371 2005 4375
rect 2001 4366 2005 4370
rect 2001 4361 2005 4365
rect 2001 4356 2005 4360
rect 2001 4351 2005 4355
rect 2001 4346 2005 4350
rect 2091 4461 2095 4465
rect 2091 4456 2095 4460
rect 2091 4451 2095 4455
rect 2091 4446 2095 4450
rect 2091 4441 2095 4445
rect 2091 4436 2095 4440
rect 2091 4431 2095 4435
rect 2091 4426 2095 4430
rect 2091 4421 2095 4425
rect 2091 4416 2095 4420
rect 2091 4411 2095 4415
rect 2091 4406 2095 4410
rect 2091 4401 2095 4405
rect 2091 4396 2095 4400
rect 2091 4391 2095 4395
rect 2091 4386 2095 4390
rect 2091 4381 2095 4385
rect 2091 4376 2095 4380
rect 2091 4371 2095 4375
rect 2091 4366 2095 4370
rect 2091 4361 2095 4365
rect 2091 4356 2095 4360
rect 2091 4351 2095 4355
rect 2001 4341 2005 4345
rect 2091 4346 2095 4350
rect 2091 4341 2095 4345
rect 2001 4336 2005 4340
rect 2006 4336 2010 4340
rect 2011 4336 2015 4340
rect 2016 4336 2020 4340
rect 2021 4336 2025 4340
rect 2026 4336 2030 4340
rect 2031 4336 2035 4340
rect 2036 4336 2040 4340
rect 2041 4336 2045 4340
rect 2046 4336 2050 4340
rect 2051 4336 2055 4340
rect 2056 4336 2060 4340
rect 2061 4336 2065 4340
rect 2066 4336 2070 4340
rect 2071 4336 2075 4340
rect 2076 4336 2080 4340
rect 2081 4336 2085 4340
rect 2086 4336 2090 4340
rect 2091 4336 2095 4340
rect 2174 4458 2178 4462
rect 2181 4458 2185 4462
rect 2186 4458 2190 4462
rect 2191 4458 2195 4462
rect 2196 4458 2200 4462
rect 2201 4458 2205 4462
rect 2206 4458 2210 4462
rect 2211 4458 2215 4462
rect 2216 4458 2220 4462
rect 2221 4458 2225 4462
rect 2226 4458 2230 4462
rect 2231 4458 2235 4462
rect 2238 4458 2242 4462
rect 2174 4451 2178 4455
rect 2238 4451 2242 4455
rect 2174 4446 2178 4450
rect 2174 4441 2178 4445
rect 2174 4436 2178 4440
rect 2174 4431 2178 4435
rect 2174 4426 2178 4430
rect 2174 4421 2178 4425
rect 2174 4416 2178 4420
rect 2174 4411 2178 4415
rect 2174 4406 2178 4410
rect 2174 4401 2178 4405
rect 2174 4396 2178 4400
rect 2174 4391 2178 4395
rect 2174 4386 2178 4390
rect 2174 4381 2178 4385
rect 2174 4376 2178 4380
rect 2174 4371 2178 4375
rect 2174 4366 2178 4370
rect 2174 4361 2178 4365
rect 2238 4446 2242 4450
rect 2238 4441 2242 4445
rect 2238 4436 2242 4440
rect 2238 4431 2242 4435
rect 2238 4426 2242 4430
rect 2238 4421 2242 4425
rect 2238 4416 2242 4420
rect 2238 4411 2242 4415
rect 2238 4406 2242 4410
rect 2238 4401 2242 4405
rect 2238 4396 2242 4400
rect 2238 4391 2242 4395
rect 2238 4386 2242 4390
rect 2238 4381 2242 4385
rect 2238 4376 2242 4380
rect 2238 4371 2242 4375
rect 2238 4366 2242 4370
rect 2238 4361 2242 4365
rect 2174 4356 2178 4360
rect 2238 4356 2242 4360
rect 2174 4349 2178 4353
rect 2181 4349 2185 4353
rect 2186 4349 2190 4353
rect 2191 4349 2195 4353
rect 2196 4349 2200 4353
rect 2201 4349 2205 4353
rect 2206 4349 2210 4353
rect 2211 4349 2215 4353
rect 2216 4349 2220 4353
rect 2221 4349 2225 4353
rect 2226 4349 2230 4353
rect 2231 4349 2235 4353
rect 2238 4349 2242 4353
rect 2310 4471 2314 4475
rect 2315 4471 2319 4475
rect 2320 4471 2324 4475
rect 2325 4471 2329 4475
rect 2330 4471 2334 4475
rect 2335 4471 2339 4475
rect 2340 4471 2344 4475
rect 2345 4471 2349 4475
rect 2350 4471 2354 4475
rect 2355 4471 2359 4475
rect 2360 4471 2364 4475
rect 2365 4471 2369 4475
rect 2370 4471 2374 4475
rect 2375 4471 2379 4475
rect 2380 4471 2384 4475
rect 2385 4471 2389 4475
rect 2390 4471 2394 4475
rect 2395 4471 2399 4475
rect 2400 4471 2404 4475
rect 2310 4466 2314 4470
rect 2310 4461 2314 4465
rect 2400 4466 2404 4470
rect 2310 4456 2314 4460
rect 2310 4451 2314 4455
rect 2310 4446 2314 4450
rect 2310 4441 2314 4445
rect 2310 4436 2314 4440
rect 2310 4431 2314 4435
rect 2310 4426 2314 4430
rect 2310 4421 2314 4425
rect 2310 4416 2314 4420
rect 2310 4411 2314 4415
rect 2310 4406 2314 4410
rect 2310 4401 2314 4405
rect 2310 4396 2314 4400
rect 2310 4391 2314 4395
rect 2310 4386 2314 4390
rect 2310 4381 2314 4385
rect 2310 4376 2314 4380
rect 2310 4371 2314 4375
rect 2310 4366 2314 4370
rect 2310 4361 2314 4365
rect 2310 4356 2314 4360
rect 2310 4351 2314 4355
rect 2310 4346 2314 4350
rect 2400 4461 2404 4465
rect 2400 4456 2404 4460
rect 2400 4451 2404 4455
rect 2400 4446 2404 4450
rect 2400 4441 2404 4445
rect 2400 4436 2404 4440
rect 2400 4431 2404 4435
rect 2400 4426 2404 4430
rect 2400 4421 2404 4425
rect 2400 4416 2404 4420
rect 2400 4411 2404 4415
rect 2400 4406 2404 4410
rect 2400 4401 2404 4405
rect 2400 4396 2404 4400
rect 2400 4391 2404 4395
rect 2400 4386 2404 4390
rect 2400 4381 2404 4385
rect 2400 4376 2404 4380
rect 2400 4371 2404 4375
rect 2400 4366 2404 4370
rect 2400 4361 2404 4365
rect 2400 4356 2404 4360
rect 2400 4351 2404 4355
rect 2310 4341 2314 4345
rect 2400 4346 2404 4350
rect 2400 4341 2404 4345
rect 2310 4336 2314 4340
rect 2315 4336 2319 4340
rect 2320 4336 2324 4340
rect 2325 4336 2329 4340
rect 2330 4336 2334 4340
rect 2335 4336 2339 4340
rect 2340 4336 2344 4340
rect 2345 4336 2349 4340
rect 2350 4336 2354 4340
rect 2355 4336 2359 4340
rect 2360 4336 2364 4340
rect 2365 4336 2369 4340
rect 2370 4336 2374 4340
rect 2375 4336 2379 4340
rect 2380 4336 2384 4340
rect 2385 4336 2389 4340
rect 2390 4336 2394 4340
rect 2395 4336 2399 4340
rect 2400 4336 2404 4340
rect 2483 4458 2487 4462
rect 2490 4458 2494 4462
rect 2495 4458 2499 4462
rect 2500 4458 2504 4462
rect 2505 4458 2509 4462
rect 2510 4458 2514 4462
rect 2515 4458 2519 4462
rect 2520 4458 2524 4462
rect 2525 4458 2529 4462
rect 2530 4458 2534 4462
rect 2535 4458 2539 4462
rect 2540 4458 2544 4462
rect 2547 4458 2551 4462
rect 2483 4451 2487 4455
rect 2547 4451 2551 4455
rect 2483 4446 2487 4450
rect 2483 4441 2487 4445
rect 2483 4436 2487 4440
rect 2483 4431 2487 4435
rect 2483 4426 2487 4430
rect 2483 4421 2487 4425
rect 2483 4416 2487 4420
rect 2483 4411 2487 4415
rect 2483 4406 2487 4410
rect 2483 4401 2487 4405
rect 2483 4396 2487 4400
rect 2483 4391 2487 4395
rect 2483 4386 2487 4390
rect 2483 4381 2487 4385
rect 2483 4376 2487 4380
rect 2483 4371 2487 4375
rect 2483 4366 2487 4370
rect 2483 4361 2487 4365
rect 2547 4446 2551 4450
rect 2547 4441 2551 4445
rect 2547 4436 2551 4440
rect 2547 4431 2551 4435
rect 2547 4426 2551 4430
rect 2547 4421 2551 4425
rect 2547 4416 2551 4420
rect 2547 4411 2551 4415
rect 2547 4406 2551 4410
rect 2547 4401 2551 4405
rect 2547 4396 2551 4400
rect 2547 4391 2551 4395
rect 2547 4386 2551 4390
rect 2547 4381 2551 4385
rect 2547 4376 2551 4380
rect 2547 4371 2551 4375
rect 2547 4366 2551 4370
rect 2547 4361 2551 4365
rect 2483 4356 2487 4360
rect 2547 4356 2551 4360
rect 2483 4349 2487 4353
rect 2490 4349 2494 4353
rect 2495 4349 2499 4353
rect 2500 4349 2504 4353
rect 2505 4349 2509 4353
rect 2510 4349 2514 4353
rect 2515 4349 2519 4353
rect 2520 4349 2524 4353
rect 2525 4349 2529 4353
rect 2530 4349 2534 4353
rect 2535 4349 2539 4353
rect 2540 4349 2544 4353
rect 2547 4349 2551 4353
rect 2619 4471 2623 4475
rect 2624 4471 2628 4475
rect 2629 4471 2633 4475
rect 2634 4471 2638 4475
rect 2639 4471 2643 4475
rect 2644 4471 2648 4475
rect 2649 4471 2653 4475
rect 2654 4471 2658 4475
rect 2659 4471 2663 4475
rect 2664 4471 2668 4475
rect 2669 4471 2673 4475
rect 2674 4471 2678 4475
rect 2679 4471 2683 4475
rect 2684 4471 2688 4475
rect 2689 4471 2693 4475
rect 2694 4471 2698 4475
rect 2699 4471 2703 4475
rect 2704 4471 2708 4475
rect 2709 4471 2713 4475
rect 2619 4466 2623 4470
rect 2619 4461 2623 4465
rect 2709 4466 2713 4470
rect 2619 4456 2623 4460
rect 2619 4451 2623 4455
rect 2619 4446 2623 4450
rect 2619 4441 2623 4445
rect 2619 4436 2623 4440
rect 2619 4431 2623 4435
rect 2619 4426 2623 4430
rect 2619 4421 2623 4425
rect 2619 4416 2623 4420
rect 2619 4411 2623 4415
rect 2619 4406 2623 4410
rect 2619 4401 2623 4405
rect 2619 4396 2623 4400
rect 2619 4391 2623 4395
rect 2619 4386 2623 4390
rect 2619 4381 2623 4385
rect 2619 4376 2623 4380
rect 2619 4371 2623 4375
rect 2619 4366 2623 4370
rect 2619 4361 2623 4365
rect 2619 4356 2623 4360
rect 2619 4351 2623 4355
rect 2619 4346 2623 4350
rect 2709 4461 2713 4465
rect 2709 4456 2713 4460
rect 2709 4451 2713 4455
rect 2709 4446 2713 4450
rect 2709 4441 2713 4445
rect 2709 4436 2713 4440
rect 2709 4431 2713 4435
rect 2709 4426 2713 4430
rect 2709 4421 2713 4425
rect 2709 4416 2713 4420
rect 2709 4411 2713 4415
rect 2709 4406 2713 4410
rect 2709 4401 2713 4405
rect 2709 4396 2713 4400
rect 2709 4391 2713 4395
rect 2709 4386 2713 4390
rect 2709 4381 2713 4385
rect 2709 4376 2713 4380
rect 2709 4371 2713 4375
rect 2709 4366 2713 4370
rect 2709 4361 2713 4365
rect 2709 4356 2713 4360
rect 2709 4351 2713 4355
rect 2619 4341 2623 4345
rect 2709 4346 2713 4350
rect 2709 4341 2713 4345
rect 2619 4336 2623 4340
rect 2624 4336 2628 4340
rect 2629 4336 2633 4340
rect 2634 4336 2638 4340
rect 2639 4336 2643 4340
rect 2644 4336 2648 4340
rect 2649 4336 2653 4340
rect 2654 4336 2658 4340
rect 2659 4336 2663 4340
rect 2664 4336 2668 4340
rect 2669 4336 2673 4340
rect 2674 4336 2678 4340
rect 2679 4336 2683 4340
rect 2684 4336 2688 4340
rect 2689 4336 2693 4340
rect 2694 4336 2698 4340
rect 2699 4336 2703 4340
rect 2704 4336 2708 4340
rect 2709 4336 2713 4340
rect 2792 4458 2796 4462
rect 2799 4458 2803 4462
rect 2804 4458 2808 4462
rect 2809 4458 2813 4462
rect 2814 4458 2818 4462
rect 2819 4458 2823 4462
rect 2824 4458 2828 4462
rect 2829 4458 2833 4462
rect 2834 4458 2838 4462
rect 2839 4458 2843 4462
rect 2844 4458 2848 4462
rect 2849 4458 2853 4462
rect 2856 4458 2860 4462
rect 2792 4451 2796 4455
rect 2856 4451 2860 4455
rect 2792 4446 2796 4450
rect 2792 4441 2796 4445
rect 2792 4436 2796 4440
rect 2792 4431 2796 4435
rect 2792 4426 2796 4430
rect 2792 4421 2796 4425
rect 2792 4416 2796 4420
rect 2792 4411 2796 4415
rect 2792 4406 2796 4410
rect 2792 4401 2796 4405
rect 2792 4396 2796 4400
rect 2792 4391 2796 4395
rect 2792 4386 2796 4390
rect 2792 4381 2796 4385
rect 2792 4376 2796 4380
rect 2792 4371 2796 4375
rect 2792 4366 2796 4370
rect 2792 4361 2796 4365
rect 2856 4446 2860 4450
rect 2856 4441 2860 4445
rect 2856 4436 2860 4440
rect 2856 4431 2860 4435
rect 2856 4426 2860 4430
rect 2856 4421 2860 4425
rect 2856 4416 2860 4420
rect 2856 4411 2860 4415
rect 2856 4406 2860 4410
rect 2856 4401 2860 4405
rect 2856 4396 2860 4400
rect 2856 4391 2860 4395
rect 2856 4386 2860 4390
rect 2856 4381 2860 4385
rect 2856 4376 2860 4380
rect 2856 4371 2860 4375
rect 2856 4366 2860 4370
rect 2856 4361 2860 4365
rect 2792 4356 2796 4360
rect 2856 4356 2860 4360
rect 2792 4349 2796 4353
rect 2799 4349 2803 4353
rect 2804 4349 2808 4353
rect 2809 4349 2813 4353
rect 2814 4349 2818 4353
rect 2819 4349 2823 4353
rect 2824 4349 2828 4353
rect 2829 4349 2833 4353
rect 2834 4349 2838 4353
rect 2839 4349 2843 4353
rect 2844 4349 2848 4353
rect 2849 4349 2853 4353
rect 2856 4349 2860 4353
rect 2928 4471 2932 4475
rect 2933 4471 2937 4475
rect 2938 4471 2942 4475
rect 2943 4471 2947 4475
rect 2948 4471 2952 4475
rect 2953 4471 2957 4475
rect 2958 4471 2962 4475
rect 2963 4471 2967 4475
rect 2968 4471 2972 4475
rect 2973 4471 2977 4475
rect 2978 4471 2982 4475
rect 2983 4471 2987 4475
rect 2988 4471 2992 4475
rect 2993 4471 2997 4475
rect 2998 4471 3002 4475
rect 3003 4471 3007 4475
rect 3008 4471 3012 4475
rect 3013 4471 3017 4475
rect 3018 4471 3022 4475
rect 2928 4466 2932 4470
rect 2928 4461 2932 4465
rect 3018 4466 3022 4470
rect 2928 4456 2932 4460
rect 2928 4451 2932 4455
rect 2928 4446 2932 4450
rect 2928 4441 2932 4445
rect 2928 4436 2932 4440
rect 2928 4431 2932 4435
rect 2928 4426 2932 4430
rect 2928 4421 2932 4425
rect 2928 4416 2932 4420
rect 2928 4411 2932 4415
rect 2928 4406 2932 4410
rect 2928 4401 2932 4405
rect 2928 4396 2932 4400
rect 2928 4391 2932 4395
rect 2928 4386 2932 4390
rect 2928 4381 2932 4385
rect 2928 4376 2932 4380
rect 2928 4371 2932 4375
rect 2928 4366 2932 4370
rect 2928 4361 2932 4365
rect 2928 4356 2932 4360
rect 2928 4351 2932 4355
rect 2928 4346 2932 4350
rect 3018 4461 3022 4465
rect 3018 4456 3022 4460
rect 3018 4451 3022 4455
rect 3018 4446 3022 4450
rect 3018 4441 3022 4445
rect 3018 4436 3022 4440
rect 3018 4431 3022 4435
rect 3018 4426 3022 4430
rect 3018 4421 3022 4425
rect 3018 4416 3022 4420
rect 3018 4411 3022 4415
rect 3018 4406 3022 4410
rect 3018 4401 3022 4405
rect 3018 4396 3022 4400
rect 3018 4391 3022 4395
rect 3018 4386 3022 4390
rect 3018 4381 3022 4385
rect 3018 4376 3022 4380
rect 3018 4371 3022 4375
rect 3018 4366 3022 4370
rect 3018 4361 3022 4365
rect 3018 4356 3022 4360
rect 3018 4351 3022 4355
rect 2928 4341 2932 4345
rect 3018 4346 3022 4350
rect 3018 4341 3022 4345
rect 2928 4336 2932 4340
rect 2933 4336 2937 4340
rect 2938 4336 2942 4340
rect 2943 4336 2947 4340
rect 2948 4336 2952 4340
rect 2953 4336 2957 4340
rect 2958 4336 2962 4340
rect 2963 4336 2967 4340
rect 2968 4336 2972 4340
rect 2973 4336 2977 4340
rect 2978 4336 2982 4340
rect 2983 4336 2987 4340
rect 2988 4336 2992 4340
rect 2993 4336 2997 4340
rect 2998 4336 3002 4340
rect 3003 4336 3007 4340
rect 3008 4336 3012 4340
rect 3013 4336 3017 4340
rect 3018 4336 3022 4340
rect 3101 4458 3105 4462
rect 3108 4458 3112 4462
rect 3113 4458 3117 4462
rect 3118 4458 3122 4462
rect 3123 4458 3127 4462
rect 3128 4458 3132 4462
rect 3133 4458 3137 4462
rect 3138 4458 3142 4462
rect 3143 4458 3147 4462
rect 3148 4458 3152 4462
rect 3153 4458 3157 4462
rect 3158 4458 3162 4462
rect 3165 4458 3169 4462
rect 3101 4451 3105 4455
rect 3165 4451 3169 4455
rect 3101 4446 3105 4450
rect 3101 4441 3105 4445
rect 3101 4436 3105 4440
rect 3101 4431 3105 4435
rect 3101 4426 3105 4430
rect 3101 4421 3105 4425
rect 3101 4416 3105 4420
rect 3101 4411 3105 4415
rect 3101 4406 3105 4410
rect 3101 4401 3105 4405
rect 3101 4396 3105 4400
rect 3101 4391 3105 4395
rect 3101 4386 3105 4390
rect 3101 4381 3105 4385
rect 3101 4376 3105 4380
rect 3101 4371 3105 4375
rect 3101 4366 3105 4370
rect 3101 4361 3105 4365
rect 3165 4446 3169 4450
rect 3165 4441 3169 4445
rect 3165 4436 3169 4440
rect 3165 4431 3169 4435
rect 3165 4426 3169 4430
rect 3165 4421 3169 4425
rect 3165 4416 3169 4420
rect 3165 4411 3169 4415
rect 3165 4406 3169 4410
rect 3165 4401 3169 4405
rect 3165 4396 3169 4400
rect 3165 4391 3169 4395
rect 3165 4386 3169 4390
rect 3165 4381 3169 4385
rect 3165 4376 3169 4380
rect 3165 4371 3169 4375
rect 3165 4366 3169 4370
rect 3165 4361 3169 4365
rect 3101 4356 3105 4360
rect 3165 4356 3169 4360
rect 3101 4349 3105 4353
rect 3108 4349 3112 4353
rect 3113 4349 3117 4353
rect 3118 4349 3122 4353
rect 3123 4349 3127 4353
rect 3128 4349 3132 4353
rect 3133 4349 3137 4353
rect 3138 4349 3142 4353
rect 3143 4349 3147 4353
rect 3148 4349 3152 4353
rect 3153 4349 3157 4353
rect 3158 4349 3162 4353
rect 3165 4349 3169 4353
rect 3237 4471 3241 4475
rect 3242 4471 3246 4475
rect 3247 4471 3251 4475
rect 3252 4471 3256 4475
rect 3257 4471 3261 4475
rect 3262 4471 3266 4475
rect 3267 4471 3271 4475
rect 3272 4471 3276 4475
rect 3277 4471 3281 4475
rect 3282 4471 3286 4475
rect 3287 4471 3291 4475
rect 3292 4471 3296 4475
rect 3297 4471 3301 4475
rect 3302 4471 3306 4475
rect 3307 4471 3311 4475
rect 3312 4471 3316 4475
rect 3317 4471 3321 4475
rect 3322 4471 3326 4475
rect 3327 4471 3331 4475
rect 3237 4466 3241 4470
rect 3237 4461 3241 4465
rect 3327 4466 3331 4470
rect 3237 4456 3241 4460
rect 3237 4451 3241 4455
rect 3237 4446 3241 4450
rect 3237 4441 3241 4445
rect 3237 4436 3241 4440
rect 3237 4431 3241 4435
rect 3237 4426 3241 4430
rect 3237 4421 3241 4425
rect 3237 4416 3241 4420
rect 3237 4411 3241 4415
rect 3237 4406 3241 4410
rect 3237 4401 3241 4405
rect 3237 4396 3241 4400
rect 3237 4391 3241 4395
rect 3237 4386 3241 4390
rect 3237 4381 3241 4385
rect 3237 4376 3241 4380
rect 3237 4371 3241 4375
rect 3237 4366 3241 4370
rect 3237 4361 3241 4365
rect 3237 4356 3241 4360
rect 3237 4351 3241 4355
rect 3237 4346 3241 4350
rect 3327 4461 3331 4465
rect 3327 4456 3331 4460
rect 3327 4451 3331 4455
rect 3327 4446 3331 4450
rect 3327 4441 3331 4445
rect 3327 4436 3331 4440
rect 3327 4431 3331 4435
rect 3327 4426 3331 4430
rect 3327 4421 3331 4425
rect 3327 4416 3331 4420
rect 3327 4411 3331 4415
rect 3327 4406 3331 4410
rect 3327 4401 3331 4405
rect 3327 4396 3331 4400
rect 3327 4391 3331 4395
rect 3327 4386 3331 4390
rect 3327 4381 3331 4385
rect 3327 4376 3331 4380
rect 3327 4371 3331 4375
rect 3327 4366 3331 4370
rect 3327 4361 3331 4365
rect 3327 4356 3331 4360
rect 3327 4351 3331 4355
rect 3237 4341 3241 4345
rect 3327 4346 3331 4350
rect 3327 4341 3331 4345
rect 3237 4336 3241 4340
rect 3242 4336 3246 4340
rect 3247 4336 3251 4340
rect 3252 4336 3256 4340
rect 3257 4336 3261 4340
rect 3262 4336 3266 4340
rect 3267 4336 3271 4340
rect 3272 4336 3276 4340
rect 3277 4336 3281 4340
rect 3282 4336 3286 4340
rect 3287 4336 3291 4340
rect 3292 4336 3296 4340
rect 3297 4336 3301 4340
rect 3302 4336 3306 4340
rect 3307 4336 3311 4340
rect 3312 4336 3316 4340
rect 3317 4336 3321 4340
rect 3322 4336 3326 4340
rect 3327 4336 3331 4340
rect 3410 4458 3414 4462
rect 3417 4458 3421 4462
rect 3422 4458 3426 4462
rect 3427 4458 3431 4462
rect 3432 4458 3436 4462
rect 3437 4458 3441 4462
rect 3442 4458 3446 4462
rect 3447 4458 3451 4462
rect 3452 4458 3456 4462
rect 3457 4458 3461 4462
rect 3462 4458 3466 4462
rect 3467 4458 3471 4462
rect 3474 4458 3478 4462
rect 3410 4451 3414 4455
rect 3474 4451 3478 4455
rect 3410 4446 3414 4450
rect 3410 4441 3414 4445
rect 3410 4436 3414 4440
rect 3410 4431 3414 4435
rect 3410 4426 3414 4430
rect 3410 4421 3414 4425
rect 3410 4416 3414 4420
rect 3410 4411 3414 4415
rect 3410 4406 3414 4410
rect 3410 4401 3414 4405
rect 3410 4396 3414 4400
rect 3410 4391 3414 4395
rect 3410 4386 3414 4390
rect 3410 4381 3414 4385
rect 3410 4376 3414 4380
rect 3410 4371 3414 4375
rect 3410 4366 3414 4370
rect 3410 4361 3414 4365
rect 3474 4446 3478 4450
rect 3474 4441 3478 4445
rect 3474 4436 3478 4440
rect 3474 4431 3478 4435
rect 3474 4426 3478 4430
rect 3474 4421 3478 4425
rect 3474 4416 3478 4420
rect 3474 4411 3478 4415
rect 3474 4406 3478 4410
rect 3474 4401 3478 4405
rect 3474 4396 3478 4400
rect 3474 4391 3478 4395
rect 3474 4386 3478 4390
rect 3474 4381 3478 4385
rect 3474 4376 3478 4380
rect 3474 4371 3478 4375
rect 3474 4366 3478 4370
rect 3474 4361 3478 4365
rect 3410 4356 3414 4360
rect 3474 4356 3478 4360
rect 3410 4349 3414 4353
rect 3417 4349 3421 4353
rect 3422 4349 3426 4353
rect 3427 4349 3431 4353
rect 3432 4349 3436 4353
rect 3437 4349 3441 4353
rect 3442 4349 3446 4353
rect 3447 4349 3451 4353
rect 3452 4349 3456 4353
rect 3457 4349 3461 4353
rect 3462 4349 3466 4353
rect 3467 4349 3471 4353
rect 3474 4349 3478 4353
rect 3546 4471 3550 4475
rect 3551 4471 3555 4475
rect 3556 4471 3560 4475
rect 3561 4471 3565 4475
rect 3566 4471 3570 4475
rect 3571 4471 3575 4475
rect 3576 4471 3580 4475
rect 3581 4471 3585 4475
rect 3586 4471 3590 4475
rect 3591 4471 3595 4475
rect 3596 4471 3600 4475
rect 3601 4471 3605 4475
rect 3606 4471 3610 4475
rect 3611 4471 3615 4475
rect 3616 4471 3620 4475
rect 3621 4471 3625 4475
rect 3626 4471 3630 4475
rect 3631 4471 3635 4475
rect 3636 4471 3640 4475
rect 3546 4466 3550 4470
rect 3546 4461 3550 4465
rect 3636 4466 3640 4470
rect 3546 4456 3550 4460
rect 3546 4451 3550 4455
rect 3546 4446 3550 4450
rect 3546 4441 3550 4445
rect 3546 4436 3550 4440
rect 3546 4431 3550 4435
rect 3546 4426 3550 4430
rect 3546 4421 3550 4425
rect 3546 4416 3550 4420
rect 3546 4411 3550 4415
rect 3546 4406 3550 4410
rect 3546 4401 3550 4405
rect 3546 4396 3550 4400
rect 3546 4391 3550 4395
rect 3546 4386 3550 4390
rect 3546 4381 3550 4385
rect 3546 4376 3550 4380
rect 3546 4371 3550 4375
rect 3546 4366 3550 4370
rect 3546 4361 3550 4365
rect 3546 4356 3550 4360
rect 3546 4351 3550 4355
rect 3546 4346 3550 4350
rect 3636 4461 3640 4465
rect 3636 4456 3640 4460
rect 3636 4451 3640 4455
rect 3636 4446 3640 4450
rect 3636 4441 3640 4445
rect 3636 4436 3640 4440
rect 3636 4431 3640 4435
rect 3636 4426 3640 4430
rect 3636 4421 3640 4425
rect 3636 4416 3640 4420
rect 3636 4411 3640 4415
rect 3636 4406 3640 4410
rect 3636 4401 3640 4405
rect 3636 4396 3640 4400
rect 3636 4391 3640 4395
rect 3636 4386 3640 4390
rect 3636 4381 3640 4385
rect 3636 4376 3640 4380
rect 3636 4371 3640 4375
rect 3636 4366 3640 4370
rect 3636 4361 3640 4365
rect 3636 4356 3640 4360
rect 3636 4351 3640 4355
rect 3546 4341 3550 4345
rect 3636 4346 3640 4350
rect 3636 4341 3640 4345
rect 3546 4336 3550 4340
rect 3551 4336 3555 4340
rect 3556 4336 3560 4340
rect 3561 4336 3565 4340
rect 3566 4336 3570 4340
rect 3571 4336 3575 4340
rect 3576 4336 3580 4340
rect 3581 4336 3585 4340
rect 3586 4336 3590 4340
rect 3591 4336 3595 4340
rect 3596 4336 3600 4340
rect 3601 4336 3605 4340
rect 3606 4336 3610 4340
rect 3611 4336 3615 4340
rect 3616 4336 3620 4340
rect 3621 4336 3625 4340
rect 3626 4336 3630 4340
rect 3631 4336 3635 4340
rect 3636 4336 3640 4340
rect 3719 4458 3723 4462
rect 3726 4458 3730 4462
rect 3731 4458 3735 4462
rect 3736 4458 3740 4462
rect 3741 4458 3745 4462
rect 3746 4458 3750 4462
rect 3751 4458 3755 4462
rect 3756 4458 3760 4462
rect 3761 4458 3765 4462
rect 3766 4458 3770 4462
rect 3771 4458 3775 4462
rect 3776 4458 3780 4462
rect 3783 4458 3787 4462
rect 3719 4451 3723 4455
rect 3783 4451 3787 4455
rect 3719 4446 3723 4450
rect 3719 4441 3723 4445
rect 3719 4436 3723 4440
rect 3719 4431 3723 4435
rect 3719 4426 3723 4430
rect 3719 4421 3723 4425
rect 3719 4416 3723 4420
rect 3719 4411 3723 4415
rect 3719 4406 3723 4410
rect 3719 4401 3723 4405
rect 3719 4396 3723 4400
rect 3719 4391 3723 4395
rect 3719 4386 3723 4390
rect 3719 4381 3723 4385
rect 3719 4376 3723 4380
rect 3719 4371 3723 4375
rect 3719 4366 3723 4370
rect 3719 4361 3723 4365
rect 3783 4446 3787 4450
rect 3783 4441 3787 4445
rect 3783 4436 3787 4440
rect 3783 4431 3787 4435
rect 3783 4426 3787 4430
rect 3783 4421 3787 4425
rect 3783 4416 3787 4420
rect 3783 4411 3787 4415
rect 3783 4406 3787 4410
rect 3783 4401 3787 4405
rect 3783 4396 3787 4400
rect 3783 4391 3787 4395
rect 3783 4386 3787 4390
rect 3783 4381 3787 4385
rect 3783 4376 3787 4380
rect 3783 4371 3787 4375
rect 3783 4366 3787 4370
rect 3783 4361 3787 4365
rect 3719 4356 3723 4360
rect 3783 4356 3787 4360
rect 3719 4349 3723 4353
rect 3726 4349 3730 4353
rect 3731 4349 3735 4353
rect 3736 4349 3740 4353
rect 3741 4349 3745 4353
rect 3746 4349 3750 4353
rect 3751 4349 3755 4353
rect 3756 4349 3760 4353
rect 3761 4349 3765 4353
rect 3766 4349 3770 4353
rect 3771 4349 3775 4353
rect 3776 4349 3780 4353
rect 3783 4349 3787 4353
<< nsubstratencontact >>
rect 1372 9974 1376 9978
rect 1377 9974 1381 9978
rect 1382 9974 1386 9978
rect 1387 9974 1391 9978
rect 1392 9974 1396 9978
rect 1397 9974 1401 9978
rect 1402 9974 1406 9978
rect 1407 9974 1411 9978
rect 1412 9974 1416 9978
rect 1417 9974 1421 9978
rect 1422 9974 1426 9978
rect 1427 9974 1431 9978
rect 1432 9974 1436 9978
rect 1437 9974 1441 9978
rect 1442 9974 1446 9978
rect 1447 9974 1451 9978
rect 1452 9974 1456 9978
rect 1457 9974 1461 9978
rect 1462 9974 1466 9978
rect 1372 9969 1376 9973
rect 1372 9964 1376 9968
rect 1462 9969 1466 9973
rect 1372 9959 1376 9963
rect 1372 9954 1376 9958
rect 1372 9949 1376 9953
rect 1372 9944 1376 9948
rect 1372 9939 1376 9943
rect 1372 9934 1376 9938
rect 1372 9929 1376 9933
rect 1372 9924 1376 9928
rect 1372 9919 1376 9923
rect 1372 9914 1376 9918
rect 1372 9909 1376 9913
rect 1372 9904 1376 9908
rect 1372 9899 1376 9903
rect 1372 9894 1376 9898
rect 1372 9889 1376 9893
rect 1372 9884 1376 9888
rect 1372 9879 1376 9883
rect 1372 9874 1376 9878
rect 1372 9869 1376 9873
rect 1372 9864 1376 9868
rect 1372 9859 1376 9863
rect 1372 9854 1376 9858
rect 1372 9849 1376 9853
rect 1462 9964 1466 9968
rect 1462 9959 1466 9963
rect 1462 9954 1466 9958
rect 1462 9949 1466 9953
rect 1462 9944 1466 9948
rect 1462 9939 1466 9943
rect 1462 9934 1466 9938
rect 1462 9929 1466 9933
rect 1462 9924 1466 9928
rect 1462 9919 1466 9923
rect 1462 9914 1466 9918
rect 1462 9909 1466 9913
rect 1462 9904 1466 9908
rect 1462 9899 1466 9903
rect 1462 9894 1466 9898
rect 1462 9889 1466 9893
rect 1462 9884 1466 9888
rect 1462 9879 1466 9883
rect 1462 9874 1466 9878
rect 1462 9869 1466 9873
rect 1462 9864 1466 9868
rect 1462 9859 1466 9863
rect 1462 9854 1466 9858
rect 1372 9844 1376 9848
rect 1462 9849 1466 9853
rect 1462 9844 1466 9848
rect 1372 9839 1376 9843
rect 1377 9839 1381 9843
rect 1382 9839 1386 9843
rect 1387 9839 1391 9843
rect 1392 9839 1396 9843
rect 1397 9839 1401 9843
rect 1402 9839 1406 9843
rect 1407 9839 1411 9843
rect 1412 9839 1416 9843
rect 1417 9839 1421 9843
rect 1422 9839 1426 9843
rect 1427 9839 1431 9843
rect 1432 9839 1436 9843
rect 1437 9839 1441 9843
rect 1442 9839 1446 9843
rect 1447 9839 1451 9843
rect 1452 9839 1456 9843
rect 1457 9839 1461 9843
rect 1462 9839 1466 9843
rect 1545 9961 1549 9965
rect 1552 9961 1556 9965
rect 1557 9961 1561 9965
rect 1562 9961 1566 9965
rect 1567 9961 1571 9965
rect 1572 9961 1576 9965
rect 1577 9961 1581 9965
rect 1582 9961 1586 9965
rect 1587 9961 1591 9965
rect 1592 9961 1596 9965
rect 1597 9961 1601 9965
rect 1602 9961 1606 9965
rect 1609 9961 1613 9965
rect 1545 9954 1549 9958
rect 1609 9954 1613 9958
rect 1545 9949 1549 9953
rect 1545 9944 1549 9948
rect 1545 9939 1549 9943
rect 1545 9934 1549 9938
rect 1545 9929 1549 9933
rect 1545 9924 1549 9928
rect 1545 9919 1549 9923
rect 1545 9914 1549 9918
rect 1545 9909 1549 9913
rect 1545 9904 1549 9908
rect 1545 9899 1549 9903
rect 1545 9894 1549 9898
rect 1545 9889 1549 9893
rect 1545 9884 1549 9888
rect 1545 9879 1549 9883
rect 1545 9874 1549 9878
rect 1545 9869 1549 9873
rect 1545 9864 1549 9868
rect 1609 9949 1613 9953
rect 1609 9944 1613 9948
rect 1609 9939 1613 9943
rect 1609 9934 1613 9938
rect 1609 9929 1613 9933
rect 1609 9924 1613 9928
rect 1609 9919 1613 9923
rect 1609 9914 1613 9918
rect 1609 9909 1613 9913
rect 1609 9904 1613 9908
rect 1609 9899 1613 9903
rect 1609 9894 1613 9898
rect 1609 9889 1613 9893
rect 1609 9884 1613 9888
rect 1609 9879 1613 9883
rect 1609 9874 1613 9878
rect 1609 9869 1613 9873
rect 1609 9864 1613 9868
rect 1545 9859 1549 9863
rect 1609 9859 1613 9863
rect 1545 9852 1549 9856
rect 1552 9852 1556 9856
rect 1557 9852 1561 9856
rect 1562 9852 1566 9856
rect 1567 9852 1571 9856
rect 1572 9852 1576 9856
rect 1577 9852 1581 9856
rect 1582 9852 1586 9856
rect 1587 9852 1591 9856
rect 1592 9852 1596 9856
rect 1597 9852 1601 9856
rect 1602 9852 1606 9856
rect 1609 9852 1613 9856
rect 1681 9974 1685 9978
rect 1686 9974 1690 9978
rect 1691 9974 1695 9978
rect 1696 9974 1700 9978
rect 1701 9974 1705 9978
rect 1706 9974 1710 9978
rect 1711 9974 1715 9978
rect 1716 9974 1720 9978
rect 1721 9974 1725 9978
rect 1726 9974 1730 9978
rect 1731 9974 1735 9978
rect 1736 9974 1740 9978
rect 1741 9974 1745 9978
rect 1746 9974 1750 9978
rect 1751 9974 1755 9978
rect 1756 9974 1760 9978
rect 1761 9974 1765 9978
rect 1766 9974 1770 9978
rect 1771 9974 1775 9978
rect 1681 9969 1685 9973
rect 1681 9964 1685 9968
rect 1771 9969 1775 9973
rect 1681 9959 1685 9963
rect 1681 9954 1685 9958
rect 1681 9949 1685 9953
rect 1681 9944 1685 9948
rect 1681 9939 1685 9943
rect 1681 9934 1685 9938
rect 1681 9929 1685 9933
rect 1681 9924 1685 9928
rect 1681 9919 1685 9923
rect 1681 9914 1685 9918
rect 1681 9909 1685 9913
rect 1681 9904 1685 9908
rect 1681 9899 1685 9903
rect 1681 9894 1685 9898
rect 1681 9889 1685 9893
rect 1681 9884 1685 9888
rect 1681 9879 1685 9883
rect 1681 9874 1685 9878
rect 1681 9869 1685 9873
rect 1681 9864 1685 9868
rect 1681 9859 1685 9863
rect 1681 9854 1685 9858
rect 1681 9849 1685 9853
rect 1771 9964 1775 9968
rect 1771 9959 1775 9963
rect 1771 9954 1775 9958
rect 1771 9949 1775 9953
rect 1771 9944 1775 9948
rect 1771 9939 1775 9943
rect 1771 9934 1775 9938
rect 1771 9929 1775 9933
rect 1771 9924 1775 9928
rect 1771 9919 1775 9923
rect 1771 9914 1775 9918
rect 1771 9909 1775 9913
rect 1771 9904 1775 9908
rect 1771 9899 1775 9903
rect 1771 9894 1775 9898
rect 1771 9889 1775 9893
rect 1771 9884 1775 9888
rect 1771 9879 1775 9883
rect 1771 9874 1775 9878
rect 1771 9869 1775 9873
rect 1771 9864 1775 9868
rect 1771 9859 1775 9863
rect 1771 9854 1775 9858
rect 1681 9844 1685 9848
rect 1771 9849 1775 9853
rect 1771 9844 1775 9848
rect 1681 9839 1685 9843
rect 1686 9839 1690 9843
rect 1691 9839 1695 9843
rect 1696 9839 1700 9843
rect 1701 9839 1705 9843
rect 1706 9839 1710 9843
rect 1711 9839 1715 9843
rect 1716 9839 1720 9843
rect 1721 9839 1725 9843
rect 1726 9839 1730 9843
rect 1731 9839 1735 9843
rect 1736 9839 1740 9843
rect 1741 9839 1745 9843
rect 1746 9839 1750 9843
rect 1751 9839 1755 9843
rect 1756 9839 1760 9843
rect 1761 9839 1765 9843
rect 1766 9839 1770 9843
rect 1771 9839 1775 9843
rect 1854 9961 1858 9965
rect 1861 9961 1865 9965
rect 1866 9961 1870 9965
rect 1871 9961 1875 9965
rect 1876 9961 1880 9965
rect 1881 9961 1885 9965
rect 1886 9961 1890 9965
rect 1891 9961 1895 9965
rect 1896 9961 1900 9965
rect 1901 9961 1905 9965
rect 1906 9961 1910 9965
rect 1911 9961 1915 9965
rect 1918 9961 1922 9965
rect 1854 9954 1858 9958
rect 1918 9954 1922 9958
rect 1854 9949 1858 9953
rect 1854 9944 1858 9948
rect 1854 9939 1858 9943
rect 1854 9934 1858 9938
rect 1854 9929 1858 9933
rect 1854 9924 1858 9928
rect 1854 9919 1858 9923
rect 1854 9914 1858 9918
rect 1854 9909 1858 9913
rect 1854 9904 1858 9908
rect 1854 9899 1858 9903
rect 1854 9894 1858 9898
rect 1854 9889 1858 9893
rect 1854 9884 1858 9888
rect 1854 9879 1858 9883
rect 1854 9874 1858 9878
rect 1854 9869 1858 9873
rect 1854 9864 1858 9868
rect 1918 9949 1922 9953
rect 1918 9944 1922 9948
rect 1918 9939 1922 9943
rect 1918 9934 1922 9938
rect 1918 9929 1922 9933
rect 1918 9924 1922 9928
rect 1918 9919 1922 9923
rect 1918 9914 1922 9918
rect 1918 9909 1922 9913
rect 1918 9904 1922 9908
rect 1918 9899 1922 9903
rect 1918 9894 1922 9898
rect 1918 9889 1922 9893
rect 1918 9884 1922 9888
rect 1918 9879 1922 9883
rect 1918 9874 1922 9878
rect 1918 9869 1922 9873
rect 1918 9864 1922 9868
rect 1854 9859 1858 9863
rect 1918 9859 1922 9863
rect 1854 9852 1858 9856
rect 1861 9852 1865 9856
rect 1866 9852 1870 9856
rect 1871 9852 1875 9856
rect 1876 9852 1880 9856
rect 1881 9852 1885 9856
rect 1886 9852 1890 9856
rect 1891 9852 1895 9856
rect 1896 9852 1900 9856
rect 1901 9852 1905 9856
rect 1906 9852 1910 9856
rect 1911 9852 1915 9856
rect 1918 9852 1922 9856
rect 1990 9974 1994 9978
rect 1995 9974 1999 9978
rect 2000 9974 2004 9978
rect 2005 9974 2009 9978
rect 2010 9974 2014 9978
rect 2015 9974 2019 9978
rect 2020 9974 2024 9978
rect 2025 9974 2029 9978
rect 2030 9974 2034 9978
rect 2035 9974 2039 9978
rect 2040 9974 2044 9978
rect 2045 9974 2049 9978
rect 2050 9974 2054 9978
rect 2055 9974 2059 9978
rect 2060 9974 2064 9978
rect 2065 9974 2069 9978
rect 2070 9974 2074 9978
rect 2075 9974 2079 9978
rect 2080 9974 2084 9978
rect 1990 9969 1994 9973
rect 1990 9964 1994 9968
rect 2080 9969 2084 9973
rect 1990 9959 1994 9963
rect 1990 9954 1994 9958
rect 1990 9949 1994 9953
rect 1990 9944 1994 9948
rect 1990 9939 1994 9943
rect 1990 9934 1994 9938
rect 1990 9929 1994 9933
rect 1990 9924 1994 9928
rect 1990 9919 1994 9923
rect 1990 9914 1994 9918
rect 1990 9909 1994 9913
rect 1990 9904 1994 9908
rect 1990 9899 1994 9903
rect 1990 9894 1994 9898
rect 1990 9889 1994 9893
rect 1990 9884 1994 9888
rect 1990 9879 1994 9883
rect 1990 9874 1994 9878
rect 1990 9869 1994 9873
rect 1990 9864 1994 9868
rect 1990 9859 1994 9863
rect 1990 9854 1994 9858
rect 1990 9849 1994 9853
rect 2080 9964 2084 9968
rect 2080 9959 2084 9963
rect 2080 9954 2084 9958
rect 2080 9949 2084 9953
rect 2080 9944 2084 9948
rect 2080 9939 2084 9943
rect 2080 9934 2084 9938
rect 2080 9929 2084 9933
rect 2080 9924 2084 9928
rect 2080 9919 2084 9923
rect 2080 9914 2084 9918
rect 2080 9909 2084 9913
rect 2080 9904 2084 9908
rect 2080 9899 2084 9903
rect 2080 9894 2084 9898
rect 2080 9889 2084 9893
rect 2080 9884 2084 9888
rect 2080 9879 2084 9883
rect 2080 9874 2084 9878
rect 2080 9869 2084 9873
rect 2080 9864 2084 9868
rect 2080 9859 2084 9863
rect 2080 9854 2084 9858
rect 1990 9844 1994 9848
rect 2080 9849 2084 9853
rect 2080 9844 2084 9848
rect 1990 9839 1994 9843
rect 1995 9839 1999 9843
rect 2000 9839 2004 9843
rect 2005 9839 2009 9843
rect 2010 9839 2014 9843
rect 2015 9839 2019 9843
rect 2020 9839 2024 9843
rect 2025 9839 2029 9843
rect 2030 9839 2034 9843
rect 2035 9839 2039 9843
rect 2040 9839 2044 9843
rect 2045 9839 2049 9843
rect 2050 9839 2054 9843
rect 2055 9839 2059 9843
rect 2060 9839 2064 9843
rect 2065 9839 2069 9843
rect 2070 9839 2074 9843
rect 2075 9839 2079 9843
rect 2080 9839 2084 9843
rect 2163 9961 2167 9965
rect 2170 9961 2174 9965
rect 2175 9961 2179 9965
rect 2180 9961 2184 9965
rect 2185 9961 2189 9965
rect 2190 9961 2194 9965
rect 2195 9961 2199 9965
rect 2200 9961 2204 9965
rect 2205 9961 2209 9965
rect 2210 9961 2214 9965
rect 2215 9961 2219 9965
rect 2220 9961 2224 9965
rect 2227 9961 2231 9965
rect 2163 9954 2167 9958
rect 2227 9954 2231 9958
rect 2163 9949 2167 9953
rect 2163 9944 2167 9948
rect 2163 9939 2167 9943
rect 2163 9934 2167 9938
rect 2163 9929 2167 9933
rect 2163 9924 2167 9928
rect 2163 9919 2167 9923
rect 2163 9914 2167 9918
rect 2163 9909 2167 9913
rect 2163 9904 2167 9908
rect 2163 9899 2167 9903
rect 2163 9894 2167 9898
rect 2163 9889 2167 9893
rect 2163 9884 2167 9888
rect 2163 9879 2167 9883
rect 2163 9874 2167 9878
rect 2163 9869 2167 9873
rect 2163 9864 2167 9868
rect 2227 9949 2231 9953
rect 2227 9944 2231 9948
rect 2227 9939 2231 9943
rect 2227 9934 2231 9938
rect 2227 9929 2231 9933
rect 2227 9924 2231 9928
rect 2227 9919 2231 9923
rect 2227 9914 2231 9918
rect 2227 9909 2231 9913
rect 2227 9904 2231 9908
rect 2227 9899 2231 9903
rect 2227 9894 2231 9898
rect 2227 9889 2231 9893
rect 2227 9884 2231 9888
rect 2227 9879 2231 9883
rect 2227 9874 2231 9878
rect 2227 9869 2231 9873
rect 2227 9864 2231 9868
rect 2163 9859 2167 9863
rect 2227 9859 2231 9863
rect 2163 9852 2167 9856
rect 2170 9852 2174 9856
rect 2175 9852 2179 9856
rect 2180 9852 2184 9856
rect 2185 9852 2189 9856
rect 2190 9852 2194 9856
rect 2195 9852 2199 9856
rect 2200 9852 2204 9856
rect 2205 9852 2209 9856
rect 2210 9852 2214 9856
rect 2215 9852 2219 9856
rect 2220 9852 2224 9856
rect 2227 9852 2231 9856
rect 2299 9974 2303 9978
rect 2304 9974 2308 9978
rect 2309 9974 2313 9978
rect 2314 9974 2318 9978
rect 2319 9974 2323 9978
rect 2324 9974 2328 9978
rect 2329 9974 2333 9978
rect 2334 9974 2338 9978
rect 2339 9974 2343 9978
rect 2344 9974 2348 9978
rect 2349 9974 2353 9978
rect 2354 9974 2358 9978
rect 2359 9974 2363 9978
rect 2364 9974 2368 9978
rect 2369 9974 2373 9978
rect 2374 9974 2378 9978
rect 2379 9974 2383 9978
rect 2384 9974 2388 9978
rect 2389 9974 2393 9978
rect 2299 9969 2303 9973
rect 2299 9964 2303 9968
rect 2389 9969 2393 9973
rect 2299 9959 2303 9963
rect 2299 9954 2303 9958
rect 2299 9949 2303 9953
rect 2299 9944 2303 9948
rect 2299 9939 2303 9943
rect 2299 9934 2303 9938
rect 2299 9929 2303 9933
rect 2299 9924 2303 9928
rect 2299 9919 2303 9923
rect 2299 9914 2303 9918
rect 2299 9909 2303 9913
rect 2299 9904 2303 9908
rect 2299 9899 2303 9903
rect 2299 9894 2303 9898
rect 2299 9889 2303 9893
rect 2299 9884 2303 9888
rect 2299 9879 2303 9883
rect 2299 9874 2303 9878
rect 2299 9869 2303 9873
rect 2299 9864 2303 9868
rect 2299 9859 2303 9863
rect 2299 9854 2303 9858
rect 2299 9849 2303 9853
rect 2389 9964 2393 9968
rect 2389 9959 2393 9963
rect 2389 9954 2393 9958
rect 2389 9949 2393 9953
rect 2389 9944 2393 9948
rect 2389 9939 2393 9943
rect 2389 9934 2393 9938
rect 2389 9929 2393 9933
rect 2389 9924 2393 9928
rect 2389 9919 2393 9923
rect 2389 9914 2393 9918
rect 2389 9909 2393 9913
rect 2389 9904 2393 9908
rect 2389 9899 2393 9903
rect 2389 9894 2393 9898
rect 2389 9889 2393 9893
rect 2389 9884 2393 9888
rect 2389 9879 2393 9883
rect 2389 9874 2393 9878
rect 2389 9869 2393 9873
rect 2389 9864 2393 9868
rect 2389 9859 2393 9863
rect 2389 9854 2393 9858
rect 2299 9844 2303 9848
rect 2389 9849 2393 9853
rect 2389 9844 2393 9848
rect 2299 9839 2303 9843
rect 2304 9839 2308 9843
rect 2309 9839 2313 9843
rect 2314 9839 2318 9843
rect 2319 9839 2323 9843
rect 2324 9839 2328 9843
rect 2329 9839 2333 9843
rect 2334 9839 2338 9843
rect 2339 9839 2343 9843
rect 2344 9839 2348 9843
rect 2349 9839 2353 9843
rect 2354 9839 2358 9843
rect 2359 9839 2363 9843
rect 2364 9839 2368 9843
rect 2369 9839 2373 9843
rect 2374 9839 2378 9843
rect 2379 9839 2383 9843
rect 2384 9839 2388 9843
rect 2389 9839 2393 9843
rect 2472 9961 2476 9965
rect 2479 9961 2483 9965
rect 2484 9961 2488 9965
rect 2489 9961 2493 9965
rect 2494 9961 2498 9965
rect 2499 9961 2503 9965
rect 2504 9961 2508 9965
rect 2509 9961 2513 9965
rect 2514 9961 2518 9965
rect 2519 9961 2523 9965
rect 2524 9961 2528 9965
rect 2529 9961 2533 9965
rect 2536 9961 2540 9965
rect 2472 9954 2476 9958
rect 2536 9954 2540 9958
rect 2472 9949 2476 9953
rect 2472 9944 2476 9948
rect 2472 9939 2476 9943
rect 2472 9934 2476 9938
rect 2472 9929 2476 9933
rect 2472 9924 2476 9928
rect 2472 9919 2476 9923
rect 2472 9914 2476 9918
rect 2472 9909 2476 9913
rect 2472 9904 2476 9908
rect 2472 9899 2476 9903
rect 2472 9894 2476 9898
rect 2472 9889 2476 9893
rect 2472 9884 2476 9888
rect 2472 9879 2476 9883
rect 2472 9874 2476 9878
rect 2472 9869 2476 9873
rect 2472 9864 2476 9868
rect 2536 9949 2540 9953
rect 2536 9944 2540 9948
rect 2536 9939 2540 9943
rect 2536 9934 2540 9938
rect 2536 9929 2540 9933
rect 2536 9924 2540 9928
rect 2536 9919 2540 9923
rect 2536 9914 2540 9918
rect 2536 9909 2540 9913
rect 2536 9904 2540 9908
rect 2536 9899 2540 9903
rect 2536 9894 2540 9898
rect 2536 9889 2540 9893
rect 2536 9884 2540 9888
rect 2536 9879 2540 9883
rect 2536 9874 2540 9878
rect 2536 9869 2540 9873
rect 2536 9864 2540 9868
rect 2472 9859 2476 9863
rect 2536 9859 2540 9863
rect 2472 9852 2476 9856
rect 2479 9852 2483 9856
rect 2484 9852 2488 9856
rect 2489 9852 2493 9856
rect 2494 9852 2498 9856
rect 2499 9852 2503 9856
rect 2504 9852 2508 9856
rect 2509 9852 2513 9856
rect 2514 9852 2518 9856
rect 2519 9852 2523 9856
rect 2524 9852 2528 9856
rect 2529 9852 2533 9856
rect 2536 9852 2540 9856
rect 2608 9974 2612 9978
rect 2613 9974 2617 9978
rect 2618 9974 2622 9978
rect 2623 9974 2627 9978
rect 2628 9974 2632 9978
rect 2633 9974 2637 9978
rect 2638 9974 2642 9978
rect 2643 9974 2647 9978
rect 2648 9974 2652 9978
rect 2653 9974 2657 9978
rect 2658 9974 2662 9978
rect 2663 9974 2667 9978
rect 2668 9974 2672 9978
rect 2673 9974 2677 9978
rect 2678 9974 2682 9978
rect 2683 9974 2687 9978
rect 2688 9974 2692 9978
rect 2693 9974 2697 9978
rect 2698 9974 2702 9978
rect 2608 9969 2612 9973
rect 2608 9964 2612 9968
rect 2698 9969 2702 9973
rect 2608 9959 2612 9963
rect 2608 9954 2612 9958
rect 2608 9949 2612 9953
rect 2608 9944 2612 9948
rect 2608 9939 2612 9943
rect 2608 9934 2612 9938
rect 2608 9929 2612 9933
rect 2608 9924 2612 9928
rect 2608 9919 2612 9923
rect 2608 9914 2612 9918
rect 2608 9909 2612 9913
rect 2608 9904 2612 9908
rect 2608 9899 2612 9903
rect 2608 9894 2612 9898
rect 2608 9889 2612 9893
rect 2608 9884 2612 9888
rect 2608 9879 2612 9883
rect 2608 9874 2612 9878
rect 2608 9869 2612 9873
rect 2608 9864 2612 9868
rect 2608 9859 2612 9863
rect 2608 9854 2612 9858
rect 2608 9849 2612 9853
rect 2698 9964 2702 9968
rect 2698 9959 2702 9963
rect 2698 9954 2702 9958
rect 2698 9949 2702 9953
rect 2698 9944 2702 9948
rect 2698 9939 2702 9943
rect 2698 9934 2702 9938
rect 2698 9929 2702 9933
rect 2698 9924 2702 9928
rect 2698 9919 2702 9923
rect 2698 9914 2702 9918
rect 2698 9909 2702 9913
rect 2698 9904 2702 9908
rect 2698 9899 2702 9903
rect 2698 9894 2702 9898
rect 2698 9889 2702 9893
rect 2698 9884 2702 9888
rect 2698 9879 2702 9883
rect 2698 9874 2702 9878
rect 2698 9869 2702 9873
rect 2698 9864 2702 9868
rect 2698 9859 2702 9863
rect 2698 9854 2702 9858
rect 2608 9844 2612 9848
rect 2698 9849 2702 9853
rect 2698 9844 2702 9848
rect 2608 9839 2612 9843
rect 2613 9839 2617 9843
rect 2618 9839 2622 9843
rect 2623 9839 2627 9843
rect 2628 9839 2632 9843
rect 2633 9839 2637 9843
rect 2638 9839 2642 9843
rect 2643 9839 2647 9843
rect 2648 9839 2652 9843
rect 2653 9839 2657 9843
rect 2658 9839 2662 9843
rect 2663 9839 2667 9843
rect 2668 9839 2672 9843
rect 2673 9839 2677 9843
rect 2678 9839 2682 9843
rect 2683 9839 2687 9843
rect 2688 9839 2692 9843
rect 2693 9839 2697 9843
rect 2698 9839 2702 9843
rect 2781 9961 2785 9965
rect 2788 9961 2792 9965
rect 2793 9961 2797 9965
rect 2798 9961 2802 9965
rect 2803 9961 2807 9965
rect 2808 9961 2812 9965
rect 2813 9961 2817 9965
rect 2818 9961 2822 9965
rect 2823 9961 2827 9965
rect 2828 9961 2832 9965
rect 2833 9961 2837 9965
rect 2838 9961 2842 9965
rect 2845 9961 2849 9965
rect 2781 9954 2785 9958
rect 2845 9954 2849 9958
rect 2781 9949 2785 9953
rect 2781 9944 2785 9948
rect 2781 9939 2785 9943
rect 2781 9934 2785 9938
rect 2781 9929 2785 9933
rect 2781 9924 2785 9928
rect 2781 9919 2785 9923
rect 2781 9914 2785 9918
rect 2781 9909 2785 9913
rect 2781 9904 2785 9908
rect 2781 9899 2785 9903
rect 2781 9894 2785 9898
rect 2781 9889 2785 9893
rect 2781 9884 2785 9888
rect 2781 9879 2785 9883
rect 2781 9874 2785 9878
rect 2781 9869 2785 9873
rect 2781 9864 2785 9868
rect 2845 9949 2849 9953
rect 2845 9944 2849 9948
rect 2845 9939 2849 9943
rect 2845 9934 2849 9938
rect 2845 9929 2849 9933
rect 2845 9924 2849 9928
rect 2845 9919 2849 9923
rect 2845 9914 2849 9918
rect 2845 9909 2849 9913
rect 2845 9904 2849 9908
rect 2845 9899 2849 9903
rect 2845 9894 2849 9898
rect 2845 9889 2849 9893
rect 2845 9884 2849 9888
rect 2845 9879 2849 9883
rect 2845 9874 2849 9878
rect 2845 9869 2849 9873
rect 2845 9864 2849 9868
rect 2781 9859 2785 9863
rect 2845 9859 2849 9863
rect 2781 9852 2785 9856
rect 2788 9852 2792 9856
rect 2793 9852 2797 9856
rect 2798 9852 2802 9856
rect 2803 9852 2807 9856
rect 2808 9852 2812 9856
rect 2813 9852 2817 9856
rect 2818 9852 2822 9856
rect 2823 9852 2827 9856
rect 2828 9852 2832 9856
rect 2833 9852 2837 9856
rect 2838 9852 2842 9856
rect 2845 9852 2849 9856
rect 2917 9974 2921 9978
rect 2922 9974 2926 9978
rect 2927 9974 2931 9978
rect 2932 9974 2936 9978
rect 2937 9974 2941 9978
rect 2942 9974 2946 9978
rect 2947 9974 2951 9978
rect 2952 9974 2956 9978
rect 2957 9974 2961 9978
rect 2962 9974 2966 9978
rect 2967 9974 2971 9978
rect 2972 9974 2976 9978
rect 2977 9974 2981 9978
rect 2982 9974 2986 9978
rect 2987 9974 2991 9978
rect 2992 9974 2996 9978
rect 2997 9974 3001 9978
rect 3002 9974 3006 9978
rect 3007 9974 3011 9978
rect 2917 9969 2921 9973
rect 2917 9964 2921 9968
rect 3007 9969 3011 9973
rect 2917 9959 2921 9963
rect 2917 9954 2921 9958
rect 2917 9949 2921 9953
rect 2917 9944 2921 9948
rect 2917 9939 2921 9943
rect 2917 9934 2921 9938
rect 2917 9929 2921 9933
rect 2917 9924 2921 9928
rect 2917 9919 2921 9923
rect 2917 9914 2921 9918
rect 2917 9909 2921 9913
rect 2917 9904 2921 9908
rect 2917 9899 2921 9903
rect 2917 9894 2921 9898
rect 2917 9889 2921 9893
rect 2917 9884 2921 9888
rect 2917 9879 2921 9883
rect 2917 9874 2921 9878
rect 2917 9869 2921 9873
rect 2917 9864 2921 9868
rect 2917 9859 2921 9863
rect 2917 9854 2921 9858
rect 2917 9849 2921 9853
rect 3007 9964 3011 9968
rect 3007 9959 3011 9963
rect 3007 9954 3011 9958
rect 3007 9949 3011 9953
rect 3007 9944 3011 9948
rect 3007 9939 3011 9943
rect 3007 9934 3011 9938
rect 3007 9929 3011 9933
rect 3007 9924 3011 9928
rect 3007 9919 3011 9923
rect 3007 9914 3011 9918
rect 3007 9909 3011 9913
rect 3007 9904 3011 9908
rect 3007 9899 3011 9903
rect 3007 9894 3011 9898
rect 3007 9889 3011 9893
rect 3007 9884 3011 9888
rect 3007 9879 3011 9883
rect 3007 9874 3011 9878
rect 3007 9869 3011 9873
rect 3007 9864 3011 9868
rect 3007 9859 3011 9863
rect 3007 9854 3011 9858
rect 2917 9844 2921 9848
rect 3007 9849 3011 9853
rect 3007 9844 3011 9848
rect 2917 9839 2921 9843
rect 2922 9839 2926 9843
rect 2927 9839 2931 9843
rect 2932 9839 2936 9843
rect 2937 9839 2941 9843
rect 2942 9839 2946 9843
rect 2947 9839 2951 9843
rect 2952 9839 2956 9843
rect 2957 9839 2961 9843
rect 2962 9839 2966 9843
rect 2967 9839 2971 9843
rect 2972 9839 2976 9843
rect 2977 9839 2981 9843
rect 2982 9839 2986 9843
rect 2987 9839 2991 9843
rect 2992 9839 2996 9843
rect 2997 9839 3001 9843
rect 3002 9839 3006 9843
rect 3007 9839 3011 9843
rect 3090 9961 3094 9965
rect 3097 9961 3101 9965
rect 3102 9961 3106 9965
rect 3107 9961 3111 9965
rect 3112 9961 3116 9965
rect 3117 9961 3121 9965
rect 3122 9961 3126 9965
rect 3127 9961 3131 9965
rect 3132 9961 3136 9965
rect 3137 9961 3141 9965
rect 3142 9961 3146 9965
rect 3147 9961 3151 9965
rect 3154 9961 3158 9965
rect 3090 9954 3094 9958
rect 3154 9954 3158 9958
rect 3090 9949 3094 9953
rect 3090 9944 3094 9948
rect 3090 9939 3094 9943
rect 3090 9934 3094 9938
rect 3090 9929 3094 9933
rect 3090 9924 3094 9928
rect 3090 9919 3094 9923
rect 3090 9914 3094 9918
rect 3090 9909 3094 9913
rect 3090 9904 3094 9908
rect 3090 9899 3094 9903
rect 3090 9894 3094 9898
rect 3090 9889 3094 9893
rect 3090 9884 3094 9888
rect 3090 9879 3094 9883
rect 3090 9874 3094 9878
rect 3090 9869 3094 9873
rect 3090 9864 3094 9868
rect 3154 9949 3158 9953
rect 3154 9944 3158 9948
rect 3154 9939 3158 9943
rect 3154 9934 3158 9938
rect 3154 9929 3158 9933
rect 3154 9924 3158 9928
rect 3154 9919 3158 9923
rect 3154 9914 3158 9918
rect 3154 9909 3158 9913
rect 3154 9904 3158 9908
rect 3154 9899 3158 9903
rect 3154 9894 3158 9898
rect 3154 9889 3158 9893
rect 3154 9884 3158 9888
rect 3154 9879 3158 9883
rect 3154 9874 3158 9878
rect 3154 9869 3158 9873
rect 3154 9864 3158 9868
rect 3090 9859 3094 9863
rect 3154 9859 3158 9863
rect 3090 9852 3094 9856
rect 3097 9852 3101 9856
rect 3102 9852 3106 9856
rect 3107 9852 3111 9856
rect 3112 9852 3116 9856
rect 3117 9852 3121 9856
rect 3122 9852 3126 9856
rect 3127 9852 3131 9856
rect 3132 9852 3136 9856
rect 3137 9852 3141 9856
rect 3142 9852 3146 9856
rect 3147 9852 3151 9856
rect 3154 9852 3158 9856
rect 3226 9974 3230 9978
rect 3231 9974 3235 9978
rect 3236 9974 3240 9978
rect 3241 9974 3245 9978
rect 3246 9974 3250 9978
rect 3251 9974 3255 9978
rect 3256 9974 3260 9978
rect 3261 9974 3265 9978
rect 3266 9974 3270 9978
rect 3271 9974 3275 9978
rect 3276 9974 3280 9978
rect 3281 9974 3285 9978
rect 3286 9974 3290 9978
rect 3291 9974 3295 9978
rect 3296 9974 3300 9978
rect 3301 9974 3305 9978
rect 3306 9974 3310 9978
rect 3311 9974 3315 9978
rect 3316 9974 3320 9978
rect 3226 9969 3230 9973
rect 3226 9964 3230 9968
rect 3316 9969 3320 9973
rect 3226 9959 3230 9963
rect 3226 9954 3230 9958
rect 3226 9949 3230 9953
rect 3226 9944 3230 9948
rect 3226 9939 3230 9943
rect 3226 9934 3230 9938
rect 3226 9929 3230 9933
rect 3226 9924 3230 9928
rect 3226 9919 3230 9923
rect 3226 9914 3230 9918
rect 3226 9909 3230 9913
rect 3226 9904 3230 9908
rect 3226 9899 3230 9903
rect 3226 9894 3230 9898
rect 3226 9889 3230 9893
rect 3226 9884 3230 9888
rect 3226 9879 3230 9883
rect 3226 9874 3230 9878
rect 3226 9869 3230 9873
rect 3226 9864 3230 9868
rect 3226 9859 3230 9863
rect 3226 9854 3230 9858
rect 3226 9849 3230 9853
rect 3316 9964 3320 9968
rect 3316 9959 3320 9963
rect 3316 9954 3320 9958
rect 3316 9949 3320 9953
rect 3316 9944 3320 9948
rect 3316 9939 3320 9943
rect 3316 9934 3320 9938
rect 3316 9929 3320 9933
rect 3316 9924 3320 9928
rect 3316 9919 3320 9923
rect 3316 9914 3320 9918
rect 3316 9909 3320 9913
rect 3316 9904 3320 9908
rect 3316 9899 3320 9903
rect 3316 9894 3320 9898
rect 3316 9889 3320 9893
rect 3316 9884 3320 9888
rect 3316 9879 3320 9883
rect 3316 9874 3320 9878
rect 3316 9869 3320 9873
rect 3316 9864 3320 9868
rect 3316 9859 3320 9863
rect 3316 9854 3320 9858
rect 3226 9844 3230 9848
rect 3316 9849 3320 9853
rect 3316 9844 3320 9848
rect 3226 9839 3230 9843
rect 3231 9839 3235 9843
rect 3236 9839 3240 9843
rect 3241 9839 3245 9843
rect 3246 9839 3250 9843
rect 3251 9839 3255 9843
rect 3256 9839 3260 9843
rect 3261 9839 3265 9843
rect 3266 9839 3270 9843
rect 3271 9839 3275 9843
rect 3276 9839 3280 9843
rect 3281 9839 3285 9843
rect 3286 9839 3290 9843
rect 3291 9839 3295 9843
rect 3296 9839 3300 9843
rect 3301 9839 3305 9843
rect 3306 9839 3310 9843
rect 3311 9839 3315 9843
rect 3316 9839 3320 9843
rect 3399 9961 3403 9965
rect 3406 9961 3410 9965
rect 3411 9961 3415 9965
rect 3416 9961 3420 9965
rect 3421 9961 3425 9965
rect 3426 9961 3430 9965
rect 3431 9961 3435 9965
rect 3436 9961 3440 9965
rect 3441 9961 3445 9965
rect 3446 9961 3450 9965
rect 3451 9961 3455 9965
rect 3456 9961 3460 9965
rect 3463 9961 3467 9965
rect 3399 9954 3403 9958
rect 3463 9954 3467 9958
rect 3399 9949 3403 9953
rect 3399 9944 3403 9948
rect 3399 9939 3403 9943
rect 3399 9934 3403 9938
rect 3399 9929 3403 9933
rect 3399 9924 3403 9928
rect 3399 9919 3403 9923
rect 3399 9914 3403 9918
rect 3399 9909 3403 9913
rect 3399 9904 3403 9908
rect 3399 9899 3403 9903
rect 3399 9894 3403 9898
rect 3399 9889 3403 9893
rect 3399 9884 3403 9888
rect 3399 9879 3403 9883
rect 3399 9874 3403 9878
rect 3399 9869 3403 9873
rect 3399 9864 3403 9868
rect 3463 9949 3467 9953
rect 3463 9944 3467 9948
rect 3463 9939 3467 9943
rect 3463 9934 3467 9938
rect 3463 9929 3467 9933
rect 3463 9924 3467 9928
rect 3463 9919 3467 9923
rect 3463 9914 3467 9918
rect 3463 9909 3467 9913
rect 3463 9904 3467 9908
rect 3463 9899 3467 9903
rect 3463 9894 3467 9898
rect 3463 9889 3467 9893
rect 3463 9884 3467 9888
rect 3463 9879 3467 9883
rect 3463 9874 3467 9878
rect 3463 9869 3467 9873
rect 3463 9864 3467 9868
rect 3399 9859 3403 9863
rect 3463 9859 3467 9863
rect 3399 9852 3403 9856
rect 3406 9852 3410 9856
rect 3411 9852 3415 9856
rect 3416 9852 3420 9856
rect 3421 9852 3425 9856
rect 3426 9852 3430 9856
rect 3431 9852 3435 9856
rect 3436 9852 3440 9856
rect 3441 9852 3445 9856
rect 3446 9852 3450 9856
rect 3451 9852 3455 9856
rect 3456 9852 3460 9856
rect 3463 9852 3467 9856
rect 3535 9974 3539 9978
rect 3540 9974 3544 9978
rect 3545 9974 3549 9978
rect 3550 9974 3554 9978
rect 3555 9974 3559 9978
rect 3560 9974 3564 9978
rect 3565 9974 3569 9978
rect 3570 9974 3574 9978
rect 3575 9974 3579 9978
rect 3580 9974 3584 9978
rect 3585 9974 3589 9978
rect 3590 9974 3594 9978
rect 3595 9974 3599 9978
rect 3600 9974 3604 9978
rect 3605 9974 3609 9978
rect 3610 9974 3614 9978
rect 3615 9974 3619 9978
rect 3620 9974 3624 9978
rect 3625 9974 3629 9978
rect 3535 9969 3539 9973
rect 3535 9964 3539 9968
rect 3625 9969 3629 9973
rect 3535 9959 3539 9963
rect 3535 9954 3539 9958
rect 3535 9949 3539 9953
rect 3535 9944 3539 9948
rect 3535 9939 3539 9943
rect 3535 9934 3539 9938
rect 3535 9929 3539 9933
rect 3535 9924 3539 9928
rect 3535 9919 3539 9923
rect 3535 9914 3539 9918
rect 3535 9909 3539 9913
rect 3535 9904 3539 9908
rect 3535 9899 3539 9903
rect 3535 9894 3539 9898
rect 3535 9889 3539 9893
rect 3535 9884 3539 9888
rect 3535 9879 3539 9883
rect 3535 9874 3539 9878
rect 3535 9869 3539 9873
rect 3535 9864 3539 9868
rect 3535 9859 3539 9863
rect 3535 9854 3539 9858
rect 3535 9849 3539 9853
rect 3625 9964 3629 9968
rect 3625 9959 3629 9963
rect 3625 9954 3629 9958
rect 3625 9949 3629 9953
rect 3625 9944 3629 9948
rect 3625 9939 3629 9943
rect 3625 9934 3629 9938
rect 3625 9929 3629 9933
rect 3625 9924 3629 9928
rect 3625 9919 3629 9923
rect 3625 9914 3629 9918
rect 3625 9909 3629 9913
rect 3625 9904 3629 9908
rect 3625 9899 3629 9903
rect 3625 9894 3629 9898
rect 3625 9889 3629 9893
rect 3625 9884 3629 9888
rect 3625 9879 3629 9883
rect 3625 9874 3629 9878
rect 3625 9869 3629 9873
rect 3625 9864 3629 9868
rect 3625 9859 3629 9863
rect 3625 9854 3629 9858
rect 3535 9844 3539 9848
rect 3625 9849 3629 9853
rect 3625 9844 3629 9848
rect 3535 9839 3539 9843
rect 3540 9839 3544 9843
rect 3545 9839 3549 9843
rect 3550 9839 3554 9843
rect 3555 9839 3559 9843
rect 3560 9839 3564 9843
rect 3565 9839 3569 9843
rect 3570 9839 3574 9843
rect 3575 9839 3579 9843
rect 3580 9839 3584 9843
rect 3585 9839 3589 9843
rect 3590 9839 3594 9843
rect 3595 9839 3599 9843
rect 3600 9839 3604 9843
rect 3605 9839 3609 9843
rect 3610 9839 3614 9843
rect 3615 9839 3619 9843
rect 3620 9839 3624 9843
rect 3625 9839 3629 9843
rect 3708 9961 3712 9965
rect 3715 9961 3719 9965
rect 3720 9961 3724 9965
rect 3725 9961 3729 9965
rect 3730 9961 3734 9965
rect 3735 9961 3739 9965
rect 3740 9961 3744 9965
rect 3745 9961 3749 9965
rect 3750 9961 3754 9965
rect 3755 9961 3759 9965
rect 3760 9961 3764 9965
rect 3765 9961 3769 9965
rect 3772 9961 3776 9965
rect 3708 9954 3712 9958
rect 3772 9954 3776 9958
rect 3708 9949 3712 9953
rect 3708 9944 3712 9948
rect 3708 9939 3712 9943
rect 3708 9934 3712 9938
rect 3708 9929 3712 9933
rect 3708 9924 3712 9928
rect 3708 9919 3712 9923
rect 3708 9914 3712 9918
rect 3708 9909 3712 9913
rect 3708 9904 3712 9908
rect 3708 9899 3712 9903
rect 3708 9894 3712 9898
rect 3708 9889 3712 9893
rect 3708 9884 3712 9888
rect 3708 9879 3712 9883
rect 3708 9874 3712 9878
rect 3708 9869 3712 9873
rect 3708 9864 3712 9868
rect 3772 9949 3776 9953
rect 3772 9944 3776 9948
rect 3772 9939 3776 9943
rect 3772 9934 3776 9938
rect 3772 9929 3776 9933
rect 3772 9924 3776 9928
rect 3772 9919 3776 9923
rect 3772 9914 3776 9918
rect 3772 9909 3776 9913
rect 3772 9904 3776 9908
rect 3772 9899 3776 9903
rect 3772 9894 3776 9898
rect 3772 9889 3776 9893
rect 3772 9884 3776 9888
rect 3772 9879 3776 9883
rect 3772 9874 3776 9878
rect 3772 9869 3776 9873
rect 3772 9864 3776 9868
rect 3708 9859 3712 9863
rect 3772 9859 3776 9863
rect 3708 9852 3712 9856
rect 3715 9852 3719 9856
rect 3720 9852 3724 9856
rect 3725 9852 3729 9856
rect 3730 9852 3734 9856
rect 3735 9852 3739 9856
rect 3740 9852 3744 9856
rect 3745 9852 3749 9856
rect 3750 9852 3754 9856
rect 3755 9852 3759 9856
rect 3760 9852 3764 9856
rect 3765 9852 3769 9856
rect 3772 9852 3776 9856
rect 3844 9974 3848 9978
rect 3849 9974 3853 9978
rect 3854 9974 3858 9978
rect 3859 9974 3863 9978
rect 3864 9974 3868 9978
rect 3869 9974 3873 9978
rect 3874 9974 3878 9978
rect 3879 9974 3883 9978
rect 3884 9974 3888 9978
rect 3889 9974 3893 9978
rect 3894 9974 3898 9978
rect 3899 9974 3903 9978
rect 3904 9974 3908 9978
rect 3909 9974 3913 9978
rect 3914 9974 3918 9978
rect 3919 9974 3923 9978
rect 3924 9974 3928 9978
rect 3929 9974 3933 9978
rect 3934 9974 3938 9978
rect 3844 9969 3848 9973
rect 3844 9964 3848 9968
rect 3934 9969 3938 9973
rect 3844 9959 3848 9963
rect 3844 9954 3848 9958
rect 3844 9949 3848 9953
rect 3844 9944 3848 9948
rect 3844 9939 3848 9943
rect 3844 9934 3848 9938
rect 3844 9929 3848 9933
rect 3844 9924 3848 9928
rect 3844 9919 3848 9923
rect 3844 9914 3848 9918
rect 3844 9909 3848 9913
rect 3844 9904 3848 9908
rect 3844 9899 3848 9903
rect 3844 9894 3848 9898
rect 3844 9889 3848 9893
rect 3844 9884 3848 9888
rect 3844 9879 3848 9883
rect 3844 9874 3848 9878
rect 3844 9869 3848 9873
rect 3844 9864 3848 9868
rect 3844 9859 3848 9863
rect 3844 9854 3848 9858
rect 3844 9849 3848 9853
rect 3934 9964 3938 9968
rect 3934 9959 3938 9963
rect 3934 9954 3938 9958
rect 3934 9949 3938 9953
rect 3934 9944 3938 9948
rect 3934 9939 3938 9943
rect 3934 9934 3938 9938
rect 3934 9929 3938 9933
rect 3934 9924 3938 9928
rect 3934 9919 3938 9923
rect 3934 9914 3938 9918
rect 3934 9909 3938 9913
rect 3934 9904 3938 9908
rect 3934 9899 3938 9903
rect 3934 9894 3938 9898
rect 3934 9889 3938 9893
rect 3934 9884 3938 9888
rect 3934 9879 3938 9883
rect 3934 9874 3938 9878
rect 3934 9869 3938 9873
rect 3934 9864 3938 9868
rect 3934 9859 3938 9863
rect 3934 9854 3938 9858
rect 3844 9844 3848 9848
rect 3934 9849 3938 9853
rect 3934 9844 3938 9848
rect 3844 9839 3848 9843
rect 3849 9839 3853 9843
rect 3854 9839 3858 9843
rect 3859 9839 3863 9843
rect 3864 9839 3868 9843
rect 3869 9839 3873 9843
rect 3874 9839 3878 9843
rect 3879 9839 3883 9843
rect 3884 9839 3888 9843
rect 3889 9839 3893 9843
rect 3894 9839 3898 9843
rect 3899 9839 3903 9843
rect 3904 9839 3908 9843
rect 3909 9839 3913 9843
rect 3914 9839 3918 9843
rect 3919 9839 3923 9843
rect 3924 9839 3928 9843
rect 3929 9839 3933 9843
rect 3934 9839 3938 9843
rect 4017 9961 4021 9965
rect 4024 9961 4028 9965
rect 4029 9961 4033 9965
rect 4034 9961 4038 9965
rect 4039 9961 4043 9965
rect 4044 9961 4048 9965
rect 4049 9961 4053 9965
rect 4054 9961 4058 9965
rect 4059 9961 4063 9965
rect 4064 9961 4068 9965
rect 4069 9961 4073 9965
rect 4074 9961 4078 9965
rect 4081 9961 4085 9965
rect 4017 9954 4021 9958
rect 4081 9954 4085 9958
rect 4017 9949 4021 9953
rect 4017 9944 4021 9948
rect 4017 9939 4021 9943
rect 4017 9934 4021 9938
rect 4017 9929 4021 9933
rect 4017 9924 4021 9928
rect 4017 9919 4021 9923
rect 4017 9914 4021 9918
rect 4017 9909 4021 9913
rect 4017 9904 4021 9908
rect 4017 9899 4021 9903
rect 4017 9894 4021 9898
rect 4017 9889 4021 9893
rect 4017 9884 4021 9888
rect 4017 9879 4021 9883
rect 4017 9874 4021 9878
rect 4017 9869 4021 9873
rect 4017 9864 4021 9868
rect 4081 9949 4085 9953
rect 4081 9944 4085 9948
rect 4081 9939 4085 9943
rect 4081 9934 4085 9938
rect 4081 9929 4085 9933
rect 4081 9924 4085 9928
rect 4081 9919 4085 9923
rect 4081 9914 4085 9918
rect 4081 9909 4085 9913
rect 4081 9904 4085 9908
rect 4081 9899 4085 9903
rect 4081 9894 4085 9898
rect 4081 9889 4085 9893
rect 4081 9884 4085 9888
rect 4081 9879 4085 9883
rect 4081 9874 4085 9878
rect 4081 9869 4085 9873
rect 4081 9864 4085 9868
rect 4017 9859 4021 9863
rect 4081 9859 4085 9863
rect 4017 9852 4021 9856
rect 4024 9852 4028 9856
rect 4029 9852 4033 9856
rect 4034 9852 4038 9856
rect 4039 9852 4043 9856
rect 4044 9852 4048 9856
rect 4049 9852 4053 9856
rect 4054 9852 4058 9856
rect 4059 9852 4063 9856
rect 4064 9852 4068 9856
rect 4069 9852 4073 9856
rect 4074 9852 4078 9856
rect 4081 9852 4085 9856
rect 802 9762 806 9766
rect 807 9762 811 9766
rect 812 9762 816 9766
rect 817 9762 821 9766
rect 831 9762 835 9766
rect 836 9762 840 9766
rect 841 9762 845 9766
rect 846 9762 850 9766
rect 860 9762 864 9766
rect 865 9762 869 9766
rect 870 9762 874 9766
rect 875 9762 879 9766
rect 889 9762 893 9766
rect 894 9762 898 9766
rect 899 9762 903 9766
rect 904 9762 908 9766
rect 918 9762 922 9766
rect 923 9762 927 9766
rect 928 9762 932 9766
rect 933 9762 937 9766
rect 1319 9762 1323 9766
rect 1324 9762 1328 9766
rect 1329 9762 1333 9766
rect 1334 9762 1338 9766
rect 1628 9762 1632 9766
rect 1633 9762 1637 9766
rect 1638 9762 1642 9766
rect 1643 9762 1647 9766
rect 1937 9762 1941 9766
rect 1942 9762 1946 9766
rect 1947 9762 1951 9766
rect 1952 9762 1956 9766
rect 2246 9762 2250 9766
rect 2251 9762 2255 9766
rect 2256 9762 2260 9766
rect 2261 9762 2265 9766
rect 2555 9762 2559 9766
rect 2560 9762 2564 9766
rect 2565 9762 2569 9766
rect 2570 9762 2574 9766
rect 2864 9762 2868 9766
rect 2869 9762 2873 9766
rect 2874 9762 2878 9766
rect 2879 9762 2883 9766
rect 3173 9762 3177 9766
rect 3178 9762 3182 9766
rect 3183 9762 3187 9766
rect 3188 9762 3192 9766
rect 3482 9762 3486 9766
rect 3487 9762 3491 9766
rect 3492 9762 3496 9766
rect 3497 9762 3501 9766
rect 3791 9762 3795 9766
rect 3796 9762 3800 9766
rect 3801 9762 3805 9766
rect 3806 9762 3810 9766
rect 4100 9762 4104 9766
rect 4105 9762 4109 9766
rect 4110 9762 4114 9766
rect 4115 9762 4119 9766
rect 4292 9762 4296 9766
rect 4297 9762 4301 9766
rect 4302 9762 4306 9766
rect 4307 9762 4311 9766
rect 4318 9762 4322 9766
rect 4323 9762 4327 9766
rect 4328 9762 4332 9766
rect 4333 9762 4337 9766
rect 4344 9762 4348 9766
rect 4349 9762 4353 9766
rect 4354 9762 4358 9766
rect 4359 9762 4363 9766
rect 4370 9762 4374 9766
rect 4375 9762 4379 9766
rect 4380 9762 4384 9766
rect 4385 9762 4389 9766
rect 4396 9762 4400 9766
rect 4401 9762 4405 9766
rect 4406 9762 4410 9766
rect 4411 9762 4415 9766
rect 802 9752 806 9756
rect 807 9752 811 9756
rect 812 9752 816 9756
rect 817 9752 821 9756
rect 831 9752 835 9756
rect 836 9752 840 9756
rect 841 9752 845 9756
rect 846 9752 850 9756
rect 860 9752 864 9756
rect 865 9752 869 9756
rect 870 9752 874 9756
rect 875 9752 879 9756
rect 889 9752 893 9756
rect 894 9752 898 9756
rect 899 9752 903 9756
rect 904 9752 908 9756
rect 918 9752 922 9756
rect 923 9752 927 9756
rect 928 9752 932 9756
rect 933 9752 937 9756
rect 1319 9752 1323 9756
rect 1324 9752 1328 9756
rect 1329 9752 1333 9756
rect 1334 9752 1338 9756
rect 1628 9752 1632 9756
rect 1633 9752 1637 9756
rect 1638 9752 1642 9756
rect 1643 9752 1647 9756
rect 1937 9752 1941 9756
rect 1942 9752 1946 9756
rect 1947 9752 1951 9756
rect 1952 9752 1956 9756
rect 2246 9752 2250 9756
rect 2251 9752 2255 9756
rect 2256 9752 2260 9756
rect 2261 9752 2265 9756
rect 2555 9752 2559 9756
rect 2560 9752 2564 9756
rect 2565 9752 2569 9756
rect 2570 9752 2574 9756
rect 2864 9752 2868 9756
rect 2869 9752 2873 9756
rect 2874 9752 2878 9756
rect 2879 9752 2883 9756
rect 3173 9752 3177 9756
rect 3178 9752 3182 9756
rect 3183 9752 3187 9756
rect 3188 9752 3192 9756
rect 3482 9752 3486 9756
rect 3487 9752 3491 9756
rect 3492 9752 3496 9756
rect 3497 9752 3501 9756
rect 3791 9752 3795 9756
rect 3796 9752 3800 9756
rect 3801 9752 3805 9756
rect 3806 9752 3810 9756
rect 4100 9752 4104 9756
rect 4105 9752 4109 9756
rect 4110 9752 4114 9756
rect 4115 9752 4119 9756
rect 4292 9752 4296 9756
rect 4297 9752 4301 9756
rect 4302 9752 4306 9756
rect 4307 9752 4311 9756
rect 4318 9752 4322 9756
rect 4323 9752 4327 9756
rect 4328 9752 4332 9756
rect 4333 9752 4337 9756
rect 4344 9752 4348 9756
rect 4349 9752 4353 9756
rect 4354 9752 4358 9756
rect 4359 9752 4363 9756
rect 4370 9752 4374 9756
rect 4375 9752 4379 9756
rect 4380 9752 4384 9756
rect 4385 9752 4389 9756
rect 4396 9752 4400 9756
rect 4401 9752 4405 9756
rect 4406 9752 4410 9756
rect 4411 9752 4415 9756
rect 802 9742 806 9746
rect 807 9742 811 9746
rect 812 9742 816 9746
rect 817 9742 821 9746
rect 831 9742 835 9746
rect 836 9742 840 9746
rect 841 9742 845 9746
rect 846 9742 850 9746
rect 860 9742 864 9746
rect 865 9742 869 9746
rect 870 9742 874 9746
rect 875 9742 879 9746
rect 889 9742 893 9746
rect 894 9742 898 9746
rect 899 9742 903 9746
rect 904 9742 908 9746
rect 918 9742 922 9746
rect 923 9742 927 9746
rect 928 9742 932 9746
rect 933 9742 937 9746
rect 1319 9742 1323 9746
rect 1324 9742 1328 9746
rect 1329 9742 1333 9746
rect 1334 9742 1338 9746
rect 1628 9742 1632 9746
rect 1633 9742 1637 9746
rect 1638 9742 1642 9746
rect 1643 9742 1647 9746
rect 1937 9742 1941 9746
rect 1942 9742 1946 9746
rect 1947 9742 1951 9746
rect 1952 9742 1956 9746
rect 2246 9742 2250 9746
rect 2251 9742 2255 9746
rect 2256 9742 2260 9746
rect 2261 9742 2265 9746
rect 2555 9742 2559 9746
rect 2560 9742 2564 9746
rect 2565 9742 2569 9746
rect 2570 9742 2574 9746
rect 2864 9742 2868 9746
rect 2869 9742 2873 9746
rect 2874 9742 2878 9746
rect 2879 9742 2883 9746
rect 3173 9742 3177 9746
rect 3178 9742 3182 9746
rect 3183 9742 3187 9746
rect 3188 9742 3192 9746
rect 3482 9742 3486 9746
rect 3487 9742 3491 9746
rect 3492 9742 3496 9746
rect 3497 9742 3501 9746
rect 3791 9742 3795 9746
rect 3796 9742 3800 9746
rect 3801 9742 3805 9746
rect 3806 9742 3810 9746
rect 4100 9742 4104 9746
rect 4105 9742 4109 9746
rect 4110 9742 4114 9746
rect 4115 9742 4119 9746
rect 4292 9742 4296 9746
rect 4297 9742 4301 9746
rect 4302 9742 4306 9746
rect 4307 9742 4311 9746
rect 4318 9742 4322 9746
rect 4323 9742 4327 9746
rect 4328 9742 4332 9746
rect 4333 9742 4337 9746
rect 4344 9742 4348 9746
rect 4349 9742 4353 9746
rect 4354 9742 4358 9746
rect 4359 9742 4363 9746
rect 4370 9742 4374 9746
rect 4375 9742 4379 9746
rect 4380 9742 4384 9746
rect 4385 9742 4389 9746
rect 4396 9742 4400 9746
rect 4401 9742 4405 9746
rect 4406 9742 4410 9746
rect 4411 9742 4415 9746
rect 802 9732 806 9736
rect 807 9732 811 9736
rect 812 9732 816 9736
rect 817 9732 821 9736
rect 831 9732 835 9736
rect 836 9732 840 9736
rect 841 9732 845 9736
rect 846 9732 850 9736
rect 860 9732 864 9736
rect 865 9732 869 9736
rect 870 9732 874 9736
rect 875 9732 879 9736
rect 889 9732 893 9736
rect 894 9732 898 9736
rect 899 9732 903 9736
rect 904 9732 908 9736
rect 918 9732 922 9736
rect 923 9732 927 9736
rect 928 9732 932 9736
rect 933 9732 937 9736
rect 1319 9732 1323 9736
rect 1324 9732 1328 9736
rect 1329 9732 1333 9736
rect 1334 9732 1338 9736
rect 1628 9732 1632 9736
rect 1633 9732 1637 9736
rect 1638 9732 1642 9736
rect 1643 9732 1647 9736
rect 1937 9732 1941 9736
rect 1942 9732 1946 9736
rect 1947 9732 1951 9736
rect 1952 9732 1956 9736
rect 2246 9732 2250 9736
rect 2251 9732 2255 9736
rect 2256 9732 2260 9736
rect 2261 9732 2265 9736
rect 2555 9732 2559 9736
rect 2560 9732 2564 9736
rect 2565 9732 2569 9736
rect 2570 9732 2574 9736
rect 2864 9732 2868 9736
rect 2869 9732 2873 9736
rect 2874 9732 2878 9736
rect 2879 9732 2883 9736
rect 3173 9732 3177 9736
rect 3178 9732 3182 9736
rect 3183 9732 3187 9736
rect 3188 9732 3192 9736
rect 3482 9732 3486 9736
rect 3487 9732 3491 9736
rect 3492 9732 3496 9736
rect 3497 9732 3501 9736
rect 3791 9732 3795 9736
rect 3796 9732 3800 9736
rect 3801 9732 3805 9736
rect 3806 9732 3810 9736
rect 4100 9732 4104 9736
rect 4105 9732 4109 9736
rect 4110 9732 4114 9736
rect 4115 9732 4119 9736
rect 4292 9732 4296 9736
rect 4297 9732 4301 9736
rect 4302 9732 4306 9736
rect 4307 9732 4311 9736
rect 4318 9732 4322 9736
rect 4323 9732 4327 9736
rect 4328 9732 4332 9736
rect 4333 9732 4337 9736
rect 4344 9732 4348 9736
rect 4349 9732 4353 9736
rect 4354 9732 4358 9736
rect 4359 9732 4363 9736
rect 4370 9732 4374 9736
rect 4375 9732 4379 9736
rect 4380 9732 4384 9736
rect 4385 9732 4389 9736
rect 4396 9732 4400 9736
rect 4401 9732 4405 9736
rect 4406 9732 4410 9736
rect 4411 9732 4415 9736
rect 613 9618 617 9622
rect 623 9618 627 9622
rect 633 9618 637 9622
rect 643 9618 647 9622
rect 613 9613 617 9617
rect 623 9613 627 9617
rect 633 9613 637 9617
rect 643 9613 647 9617
rect 613 9608 617 9612
rect 623 9608 627 9612
rect 633 9608 637 9612
rect 643 9608 647 9612
rect 613 9603 617 9607
rect 623 9603 627 9607
rect 633 9603 637 9607
rect 643 9603 647 9607
rect 613 9592 617 9596
rect 623 9592 627 9596
rect 633 9592 637 9596
rect 643 9592 647 9596
rect 613 9587 617 9591
rect 623 9587 627 9591
rect 633 9587 637 9591
rect 643 9587 647 9591
rect 613 9582 617 9586
rect 623 9582 627 9586
rect 633 9582 637 9586
rect 643 9582 647 9586
rect 613 9577 617 9581
rect 623 9577 627 9581
rect 633 9577 637 9581
rect 643 9577 647 9581
rect 613 9566 617 9570
rect 623 9566 627 9570
rect 633 9566 637 9570
rect 643 9566 647 9570
rect 613 9561 617 9565
rect 623 9561 627 9565
rect 633 9561 637 9565
rect 643 9561 647 9565
rect 613 9556 617 9560
rect 623 9556 627 9560
rect 633 9556 637 9560
rect 643 9556 647 9560
rect 613 9551 617 9555
rect 623 9551 627 9555
rect 633 9551 637 9555
rect 643 9551 647 9555
rect 613 9540 617 9544
rect 623 9540 627 9544
rect 633 9540 637 9544
rect 643 9540 647 9544
rect 613 9535 617 9539
rect 623 9535 627 9539
rect 633 9535 637 9539
rect 643 9535 647 9539
rect 613 9530 617 9534
rect 623 9530 627 9534
rect 633 9530 637 9534
rect 643 9530 647 9534
rect 613 9525 617 9529
rect 623 9525 627 9529
rect 633 9525 637 9529
rect 643 9525 647 9529
rect 613 9514 617 9518
rect 623 9514 627 9518
rect 633 9514 637 9518
rect 643 9514 647 9518
rect 613 9509 617 9513
rect 623 9509 627 9513
rect 633 9509 637 9513
rect 643 9509 647 9513
rect 613 9504 617 9508
rect 623 9504 627 9508
rect 633 9504 637 9508
rect 643 9504 647 9508
rect 613 9499 617 9503
rect 623 9499 627 9503
rect 633 9499 637 9503
rect 643 9499 647 9503
rect 613 9321 617 9325
rect 623 9321 627 9325
rect 633 9321 637 9325
rect 643 9321 647 9325
rect 613 9316 617 9320
rect 623 9316 627 9320
rect 633 9316 637 9320
rect 643 9316 647 9320
rect 613 9311 617 9315
rect 623 9311 627 9315
rect 633 9311 637 9315
rect 643 9311 647 9315
rect 613 9306 617 9310
rect 623 9306 627 9310
rect 633 9306 637 9310
rect 643 9306 647 9310
rect 613 9012 617 9016
rect 623 9012 627 9016
rect 633 9012 637 9016
rect 643 9012 647 9016
rect 613 9007 617 9011
rect 623 9007 627 9011
rect 633 9007 637 9011
rect 643 9007 647 9011
rect 613 9002 617 9006
rect 623 9002 627 9006
rect 633 9002 637 9006
rect 643 9002 647 9006
rect 613 8997 617 9001
rect 623 8997 627 9001
rect 633 8997 637 9001
rect 643 8997 647 9001
rect 613 8703 617 8707
rect 623 8703 627 8707
rect 633 8703 637 8707
rect 643 8703 647 8707
rect 613 8698 617 8702
rect 623 8698 627 8702
rect 633 8698 637 8702
rect 643 8698 647 8702
rect 613 8693 617 8697
rect 623 8693 627 8697
rect 633 8693 637 8697
rect 643 8693 647 8697
rect 613 8688 617 8692
rect 623 8688 627 8692
rect 633 8688 637 8692
rect 643 8688 647 8692
rect 613 8394 617 8398
rect 623 8394 627 8398
rect 633 8394 637 8398
rect 643 8394 647 8398
rect 613 8389 617 8393
rect 623 8389 627 8393
rect 633 8389 637 8393
rect 643 8389 647 8393
rect 613 8384 617 8388
rect 623 8384 627 8388
rect 633 8384 637 8388
rect 643 8384 647 8388
rect 613 8379 617 8383
rect 623 8379 627 8383
rect 633 8379 637 8383
rect 643 8379 647 8383
rect 613 8085 617 8089
rect 623 8085 627 8089
rect 633 8085 637 8089
rect 643 8085 647 8089
rect 613 8080 617 8084
rect 623 8080 627 8084
rect 633 8080 637 8084
rect 643 8080 647 8084
rect 613 8075 617 8079
rect 623 8075 627 8079
rect 633 8075 637 8079
rect 643 8075 647 8079
rect 613 8070 617 8074
rect 623 8070 627 8074
rect 633 8070 637 8074
rect 643 8070 647 8074
rect 613 7776 617 7780
rect 623 7776 627 7780
rect 633 7776 637 7780
rect 643 7776 647 7780
rect 613 7771 617 7775
rect 623 7771 627 7775
rect 633 7771 637 7775
rect 643 7771 647 7775
rect 613 7766 617 7770
rect 623 7766 627 7770
rect 633 7766 637 7770
rect 643 7766 647 7770
rect 613 7761 617 7765
rect 623 7761 627 7765
rect 633 7761 637 7765
rect 643 7761 647 7765
rect 613 7467 617 7471
rect 623 7467 627 7471
rect 633 7467 637 7471
rect 643 7467 647 7471
rect 613 7462 617 7466
rect 623 7462 627 7466
rect 633 7462 637 7466
rect 643 7462 647 7466
rect 613 7457 617 7461
rect 623 7457 627 7461
rect 633 7457 637 7461
rect 643 7457 647 7461
rect 613 7452 617 7456
rect 623 7452 627 7456
rect 633 7452 637 7456
rect 643 7452 647 7456
rect 613 7158 617 7162
rect 623 7158 627 7162
rect 633 7158 637 7162
rect 643 7158 647 7162
rect 613 7123 617 7127
rect 623 7123 627 7127
rect 633 7123 637 7127
rect 643 7123 647 7127
rect 613 7118 617 7122
rect 623 7118 627 7122
rect 633 7118 637 7122
rect 643 7118 647 7122
rect 613 7113 617 7117
rect 623 7113 627 7117
rect 633 7113 637 7117
rect 643 7113 647 7117
rect 613 7108 617 7112
rect 623 7108 627 7112
rect 633 7108 637 7112
rect 643 7108 647 7112
rect 613 6536 617 6540
rect 623 6536 627 6540
rect 633 6536 637 6540
rect 643 6536 647 6540
rect 613 6531 617 6535
rect 623 6531 627 6535
rect 633 6531 637 6535
rect 643 6531 647 6535
rect 613 6526 617 6530
rect 623 6526 627 6530
rect 633 6526 637 6530
rect 643 6526 647 6530
rect 613 6521 617 6525
rect 623 6521 627 6525
rect 633 6521 637 6525
rect 643 6521 647 6525
rect 418 6369 422 6457
rect 459 6369 463 6457
rect 502 6369 506 6457
rect 541 6369 545 6425
rect 613 6227 617 6231
rect 623 6227 627 6231
rect 633 6227 637 6231
rect 643 6227 647 6231
rect 613 6222 617 6226
rect 623 6222 627 6226
rect 633 6222 637 6226
rect 643 6222 647 6226
rect 613 6217 617 6221
rect 623 6217 627 6221
rect 633 6217 637 6221
rect 643 6217 647 6221
rect 613 6212 617 6216
rect 623 6212 627 6216
rect 633 6212 637 6216
rect 643 6212 647 6216
rect 613 6196 617 6200
rect 623 6196 627 6200
rect 633 6196 637 6200
rect 643 6196 647 6200
rect 613 6191 617 6195
rect 623 6191 627 6195
rect 633 6191 637 6195
rect 643 6191 647 6195
rect 613 6186 617 6190
rect 623 6186 627 6190
rect 633 6186 637 6190
rect 643 6186 647 6190
rect 613 6181 617 6185
rect 623 6181 627 6185
rect 633 6181 637 6185
rect 643 6181 647 6185
rect 613 5887 617 5891
rect 623 5887 627 5891
rect 633 5887 637 5891
rect 643 5887 647 5891
rect 613 5882 617 5886
rect 623 5882 627 5886
rect 633 5882 637 5886
rect 643 5882 647 5886
rect 613 5877 617 5881
rect 623 5877 627 5881
rect 633 5877 637 5881
rect 643 5877 647 5881
rect 613 5872 617 5876
rect 623 5872 627 5876
rect 633 5872 637 5876
rect 643 5872 647 5876
rect 613 5578 617 5582
rect 623 5578 627 5582
rect 633 5578 637 5582
rect 643 5578 647 5582
rect 613 5573 617 5577
rect 623 5573 627 5577
rect 633 5573 637 5577
rect 643 5573 647 5577
rect 613 5568 617 5572
rect 623 5568 627 5572
rect 633 5568 637 5572
rect 643 5568 647 5572
rect 613 5563 617 5567
rect 623 5563 627 5567
rect 633 5563 637 5567
rect 643 5563 647 5567
rect 613 5269 617 5273
rect 623 5269 627 5273
rect 633 5269 637 5273
rect 643 5269 647 5273
rect 613 5264 617 5268
rect 623 5264 627 5268
rect 633 5264 637 5268
rect 643 5264 647 5268
rect 613 5259 617 5263
rect 623 5259 627 5263
rect 633 5259 637 5263
rect 643 5259 647 5263
rect 613 5254 617 5258
rect 623 5254 627 5258
rect 633 5254 637 5258
rect 643 5254 647 5258
rect 613 4868 617 4872
rect 623 4868 627 4872
rect 633 4868 637 4872
rect 643 4868 647 4872
rect 613 4863 617 4867
rect 623 4863 627 4867
rect 633 4863 637 4867
rect 643 4863 647 4867
rect 613 4858 617 4862
rect 623 4858 627 4862
rect 633 4858 637 4862
rect 643 4858 647 4862
rect 613 4853 617 4857
rect 623 4853 627 4857
rect 633 4853 637 4857
rect 643 4853 647 4857
rect 613 4839 617 4843
rect 623 4839 627 4843
rect 633 4839 637 4843
rect 643 4839 647 4843
rect 613 4834 617 4838
rect 623 4834 627 4838
rect 633 4834 637 4838
rect 643 4834 647 4838
rect 613 4829 617 4833
rect 623 4829 627 4833
rect 633 4829 637 4833
rect 643 4829 647 4833
rect 613 4824 617 4828
rect 623 4824 627 4828
rect 633 4824 637 4828
rect 643 4824 647 4828
rect 613 4810 617 4814
rect 623 4810 627 4814
rect 633 4810 637 4814
rect 643 4810 647 4814
rect 613 4805 617 4809
rect 623 4805 627 4809
rect 633 4805 637 4809
rect 643 4805 647 4809
rect 613 4800 617 4804
rect 623 4800 627 4804
rect 633 4800 637 4804
rect 643 4800 647 4804
rect 613 4795 617 4799
rect 623 4795 627 4799
rect 633 4795 637 4799
rect 643 4795 647 4799
rect 613 4781 617 4785
rect 623 4781 627 4785
rect 633 4781 637 4785
rect 643 4781 647 4785
rect 613 4776 617 4780
rect 623 4776 627 4780
rect 633 4776 637 4780
rect 643 4776 647 4780
rect 613 4771 617 4775
rect 623 4771 627 4775
rect 633 4771 637 4775
rect 643 4771 647 4775
rect 613 4766 617 4770
rect 623 4766 627 4770
rect 633 4766 637 4770
rect 643 4766 647 4770
rect 613 4752 617 4756
rect 623 4752 627 4756
rect 633 4752 637 4756
rect 643 4752 647 4756
rect 613 4747 617 4751
rect 623 4747 627 4751
rect 633 4747 637 4751
rect 643 4747 647 4751
rect 613 4742 617 4746
rect 623 4742 627 4746
rect 633 4742 637 4746
rect 643 4742 647 4746
rect 613 4737 617 4741
rect 623 4737 627 4741
rect 633 4737 637 4741
rect 643 4737 647 4741
rect 2881 9340 2885 9344
rect 2909 9340 2913 9344
rect 2939 9340 2943 9344
rect 2976 9340 2980 9344
rect 3013 9340 3017 9344
rect 3041 9340 3045 9344
rect 3071 9340 3075 9344
rect 3108 9340 3112 9344
rect 3145 9340 3149 9344
rect 3173 9340 3177 9344
rect 3203 9340 3207 9344
rect 3240 9340 3244 9344
rect 3277 9340 3281 9344
rect 3305 9340 3309 9344
rect 3335 9340 3339 9344
rect 3372 9340 3376 9344
rect 3826 9340 3830 9344
rect 3854 9340 3858 9344
rect 3884 9340 3888 9344
rect 3921 9340 3925 9344
rect 3958 9340 3962 9344
rect 3986 9340 3990 9344
rect 4016 9340 4020 9344
rect 4053 9340 4057 9344
rect 4090 9340 4094 9344
rect 4118 9340 4122 9344
rect 4148 9340 4152 9344
rect 4185 9340 4189 9344
rect 4222 9340 4226 9344
rect 4250 9340 4254 9344
rect 4280 9340 4284 9344
rect 4317 9340 4321 9344
rect 2529 9307 2533 9311
rect 2557 9307 2561 9311
rect 2587 9307 2591 9311
rect 2624 9307 2628 9311
rect 3474 9307 3478 9311
rect 3502 9307 3506 9311
rect 3532 9307 3536 9311
rect 3569 9307 3573 9311
rect 2871 9263 2875 9267
rect 2900 9263 2904 9267
rect 2925 9263 2929 9267
rect 2967 9263 2971 9267
rect 3023 9263 3027 9267
rect 3047 9263 3051 9267
rect 3101 9263 3105 9267
rect 3128 9263 3132 9267
rect 3182 9263 3186 9267
rect 3816 9263 3820 9267
rect 3845 9263 3849 9267
rect 3870 9263 3874 9267
rect 3912 9263 3916 9267
rect 3968 9263 3972 9267
rect 3992 9263 3996 9267
rect 4046 9263 4050 9267
rect 4073 9263 4077 9267
rect 4127 9263 4131 9267
rect 2489 9205 2493 9209
rect 2526 9205 2530 9209
rect 2556 9205 2560 9209
rect 2584 9205 2588 9209
rect 3434 9205 3438 9209
rect 3471 9205 3475 9209
rect 3501 9205 3505 9209
rect 3529 9205 3533 9209
rect 2871 9131 2875 9135
rect 2900 9131 2904 9135
rect 2925 9131 2929 9135
rect 2967 9131 2971 9135
rect 3023 9131 3027 9135
rect 3047 9131 3051 9135
rect 3101 9131 3105 9135
rect 3128 9131 3132 9135
rect 3190 9131 3194 9135
rect 3816 9131 3820 9135
rect 3845 9131 3849 9135
rect 3870 9131 3874 9135
rect 3912 9131 3916 9135
rect 3968 9131 3972 9135
rect 3992 9131 3996 9135
rect 4046 9131 4050 9135
rect 4073 9131 4077 9135
rect 4135 9131 4139 9135
rect 3359 9102 3363 9106
rect 3383 9102 3387 9106
rect 3437 9102 3441 9106
rect 3580 9102 3584 9106
rect 2871 8999 2875 9003
rect 2900 8999 2904 9003
rect 2925 8999 2929 9003
rect 2967 8999 2971 9003
rect 3023 8999 3027 9003
rect 3047 8999 3051 9003
rect 3101 8999 3105 9003
rect 3128 8999 3132 9003
rect 3182 8999 3186 9003
rect 3190 8999 3194 9003
rect 3218 8999 3222 9003
rect 3272 8999 3276 9003
rect 3816 8999 3820 9003
rect 3845 8999 3849 9003
rect 3870 8999 3874 9003
rect 3912 8999 3916 9003
rect 3968 8999 3972 9003
rect 3992 8999 3996 9003
rect 4046 8999 4050 9003
rect 4073 8999 4077 9003
rect 4127 8999 4131 9003
rect 4135 8999 4139 9003
rect 4163 8999 4167 9003
rect 4217 8999 4221 9003
rect 3337 8972 3341 8976
rect 3359 8972 3363 8976
rect 3383 8972 3387 8976
rect 3437 8972 3441 8976
rect 3486 8972 3490 8976
rect 2871 8867 2875 8871
rect 2900 8867 2904 8871
rect 2925 8867 2929 8871
rect 2967 8867 2971 8871
rect 3023 8867 3027 8871
rect 3047 8867 3051 8871
rect 3101 8867 3105 8871
rect 3128 8867 3132 8871
rect 3218 8867 3222 8871
rect 3816 8867 3820 8871
rect 3845 8867 3849 8871
rect 3870 8867 3874 8871
rect 3912 8867 3916 8871
rect 3968 8867 3972 8871
rect 3992 8867 3996 8871
rect 4046 8867 4050 8871
rect 4073 8867 4077 8871
rect 4163 8867 4167 8871
rect 3383 8842 3387 8846
rect 2397 8805 2401 8809
rect 2425 8805 2429 8809
rect 2455 8805 2459 8809
rect 2492 8805 2496 8809
rect 2529 8805 2533 8809
rect 2557 8805 2561 8809
rect 2587 8805 2591 8809
rect 2624 8805 2628 8809
rect 2661 8805 2665 8809
rect 2689 8805 2693 8809
rect 2719 8805 2723 8809
rect 2756 8805 2760 8809
rect 3342 8805 3346 8809
rect 3370 8805 3374 8809
rect 3400 8805 3404 8809
rect 3437 8805 3441 8809
rect 3474 8805 3478 8809
rect 3502 8805 3506 8809
rect 3532 8805 3536 8809
rect 3569 8805 3573 8809
rect 3606 8805 3610 8809
rect 3634 8805 3638 8809
rect 3664 8805 3668 8809
rect 3701 8805 3705 8809
rect 2871 8735 2875 8739
rect 2900 8735 2904 8739
rect 2925 8735 2929 8739
rect 2967 8735 2971 8739
rect 3047 8735 3051 8739
rect 3101 8735 3105 8739
rect 3132 8735 3136 8739
rect 3161 8735 3165 8739
rect 3186 8735 3190 8739
rect 3228 8735 3232 8739
rect 3816 8735 3820 8739
rect 3845 8735 3849 8739
rect 3870 8735 3874 8739
rect 3912 8735 3916 8739
rect 3992 8735 3996 8739
rect 4046 8735 4050 8739
rect 4077 8735 4081 8739
rect 4106 8735 4110 8739
rect 4131 8735 4135 8739
rect 4173 8735 4177 8739
rect 3180 8693 3184 8697
rect 3208 8693 3212 8697
rect 3238 8693 3242 8697
rect 3275 8693 3279 8697
rect 4125 8693 4129 8697
rect 4153 8693 4157 8697
rect 4183 8693 4187 8697
rect 4220 8693 4224 8697
rect 2397 8663 2401 8667
rect 2425 8663 2429 8667
rect 2455 8663 2459 8667
rect 2492 8663 2496 8667
rect 2529 8663 2533 8667
rect 2557 8663 2561 8667
rect 2587 8663 2591 8667
rect 2624 8663 2628 8667
rect 2661 8663 2665 8667
rect 2689 8663 2693 8667
rect 2719 8663 2723 8667
rect 2756 8663 2760 8667
rect 3342 8663 3346 8667
rect 3370 8663 3374 8667
rect 3400 8663 3404 8667
rect 3437 8663 3441 8667
rect 3474 8663 3478 8667
rect 3502 8663 3506 8667
rect 3532 8663 3536 8667
rect 3569 8663 3573 8667
rect 3606 8663 3610 8667
rect 3634 8663 3638 8667
rect 3664 8663 3668 8667
rect 3701 8663 3705 8667
rect 3180 8607 3184 8611
rect 3208 8607 3212 8611
rect 3238 8607 3242 8611
rect 3275 8607 3279 8611
rect 4125 8607 4129 8611
rect 4153 8607 4157 8611
rect 4183 8607 4187 8611
rect 4220 8607 4224 8611
rect 2397 8577 2401 8581
rect 2425 8577 2429 8581
rect 2455 8577 2459 8581
rect 2492 8577 2496 8581
rect 2529 8577 2533 8581
rect 2557 8577 2561 8581
rect 2587 8577 2591 8581
rect 2624 8577 2628 8581
rect 2661 8577 2665 8581
rect 2689 8577 2693 8581
rect 2719 8577 2723 8581
rect 2756 8577 2760 8581
rect 3342 8577 3346 8581
rect 3370 8577 3374 8581
rect 3400 8577 3404 8581
rect 3437 8577 3441 8581
rect 3474 8577 3478 8581
rect 3502 8577 3506 8581
rect 3532 8577 3536 8581
rect 3569 8577 3573 8581
rect 3606 8577 3610 8581
rect 3634 8577 3638 8581
rect 3664 8577 3668 8581
rect 3701 8577 3705 8581
rect 2397 8437 2401 8441
rect 2425 8437 2429 8441
rect 2455 8437 2459 8441
rect 2492 8437 2496 8441
rect 2529 8437 2533 8441
rect 2557 8437 2561 8441
rect 2587 8437 2591 8441
rect 2624 8437 2628 8441
rect 2661 8437 2665 8441
rect 2689 8437 2693 8441
rect 2719 8437 2723 8441
rect 2756 8437 2760 8441
rect 3342 8437 3346 8441
rect 3370 8437 3374 8441
rect 3400 8437 3404 8441
rect 3437 8437 3441 8441
rect 3474 8437 3478 8441
rect 3502 8437 3506 8441
rect 3532 8437 3536 8441
rect 3569 8437 3573 8441
rect 3606 8437 3610 8441
rect 3634 8437 3638 8441
rect 3664 8437 3668 8441
rect 3701 8437 3705 8441
rect 2881 8358 2885 8362
rect 2909 8358 2913 8362
rect 2939 8358 2943 8362
rect 2976 8358 2980 8362
rect 3013 8358 3017 8362
rect 3041 8358 3045 8362
rect 3071 8358 3075 8362
rect 3108 8358 3112 8362
rect 3145 8358 3149 8362
rect 3173 8358 3177 8362
rect 3203 8358 3207 8362
rect 3240 8358 3244 8362
rect 3277 8358 3281 8362
rect 3305 8358 3309 8362
rect 3335 8358 3339 8362
rect 3372 8358 3376 8362
rect 3826 8358 3830 8362
rect 3854 8358 3858 8362
rect 3884 8358 3888 8362
rect 3921 8358 3925 8362
rect 3958 8358 3962 8362
rect 3986 8358 3990 8362
rect 4016 8358 4020 8362
rect 4053 8358 4057 8362
rect 4090 8358 4094 8362
rect 4118 8358 4122 8362
rect 4148 8358 4152 8362
rect 4185 8358 4189 8362
rect 4222 8358 4226 8362
rect 4250 8358 4254 8362
rect 4280 8358 4284 8362
rect 4317 8358 4321 8362
rect 2529 8325 2533 8329
rect 2557 8325 2561 8329
rect 2587 8325 2591 8329
rect 2624 8325 2628 8329
rect 3474 8325 3478 8329
rect 3502 8325 3506 8329
rect 3532 8325 3536 8329
rect 3569 8325 3573 8329
rect 2871 8281 2875 8285
rect 2900 8281 2904 8285
rect 2925 8281 2929 8285
rect 2967 8281 2971 8285
rect 3023 8281 3027 8285
rect 3047 8281 3051 8285
rect 3101 8281 3105 8285
rect 3128 8281 3132 8285
rect 3182 8281 3186 8285
rect 3816 8281 3820 8285
rect 3845 8281 3849 8285
rect 3870 8281 3874 8285
rect 3912 8281 3916 8285
rect 3968 8281 3972 8285
rect 3992 8281 3996 8285
rect 4046 8281 4050 8285
rect 4073 8281 4077 8285
rect 4127 8281 4131 8285
rect 2489 8223 2493 8227
rect 2526 8223 2530 8227
rect 2556 8223 2560 8227
rect 2584 8223 2588 8227
rect 3434 8223 3438 8227
rect 3471 8223 3475 8227
rect 3501 8223 3505 8227
rect 3529 8223 3533 8227
rect 2871 8149 2875 8153
rect 2900 8149 2904 8153
rect 2925 8149 2929 8153
rect 2967 8149 2971 8153
rect 3023 8149 3027 8153
rect 3047 8149 3051 8153
rect 3101 8149 3105 8153
rect 3128 8149 3132 8153
rect 3190 8149 3194 8153
rect 3816 8149 3820 8153
rect 3845 8149 3849 8153
rect 3870 8149 3874 8153
rect 3912 8149 3916 8153
rect 3968 8149 3972 8153
rect 3992 8149 3996 8153
rect 4046 8149 4050 8153
rect 4073 8149 4077 8153
rect 4135 8149 4139 8153
rect 2871 8017 2875 8021
rect 2900 8017 2904 8021
rect 2925 8017 2929 8021
rect 2967 8017 2971 8021
rect 3023 8017 3027 8021
rect 3047 8017 3051 8021
rect 3101 8017 3105 8021
rect 3128 8017 3132 8021
rect 3182 8017 3186 8021
rect 3190 8017 3194 8021
rect 3218 8017 3222 8021
rect 3272 8017 3276 8021
rect 3816 8017 3820 8021
rect 3845 8017 3849 8021
rect 3870 8017 3874 8021
rect 3912 8017 3916 8021
rect 3968 8017 3972 8021
rect 3992 8017 3996 8021
rect 4046 8017 4050 8021
rect 4073 8017 4077 8021
rect 4127 8017 4131 8021
rect 4135 8017 4139 8021
rect 4163 8017 4167 8021
rect 4217 8017 4221 8021
rect 2871 7885 2875 7889
rect 2900 7885 2904 7889
rect 2925 7885 2929 7889
rect 2967 7885 2971 7889
rect 3023 7885 3027 7889
rect 3047 7885 3051 7889
rect 3101 7885 3105 7889
rect 3128 7885 3132 7889
rect 3218 7885 3222 7889
rect 3816 7885 3820 7889
rect 3845 7885 3849 7889
rect 3870 7885 3874 7889
rect 3912 7885 3916 7889
rect 3968 7885 3972 7889
rect 3992 7885 3996 7889
rect 4046 7885 4050 7889
rect 4073 7885 4077 7889
rect 4163 7885 4167 7889
rect 2397 7823 2401 7827
rect 2425 7823 2429 7827
rect 2455 7823 2459 7827
rect 2492 7823 2496 7827
rect 2529 7823 2533 7827
rect 2557 7823 2561 7827
rect 2587 7823 2591 7827
rect 2624 7823 2628 7827
rect 2661 7823 2665 7827
rect 2689 7823 2693 7827
rect 2719 7823 2723 7827
rect 2756 7823 2760 7827
rect 3342 7823 3346 7827
rect 3370 7823 3374 7827
rect 3400 7823 3404 7827
rect 3437 7823 3441 7827
rect 3474 7823 3478 7827
rect 3502 7823 3506 7827
rect 3532 7823 3536 7827
rect 3569 7823 3573 7827
rect 3606 7823 3610 7827
rect 3634 7823 3638 7827
rect 3664 7823 3668 7827
rect 3701 7823 3705 7827
rect 2871 7753 2875 7757
rect 2900 7753 2904 7757
rect 2925 7753 2929 7757
rect 2967 7753 2971 7757
rect 3047 7753 3051 7757
rect 3101 7753 3105 7757
rect 3132 7753 3136 7757
rect 3161 7753 3165 7757
rect 3186 7753 3190 7757
rect 3228 7753 3232 7757
rect 3816 7753 3820 7757
rect 3845 7753 3849 7757
rect 3870 7753 3874 7757
rect 3912 7753 3916 7757
rect 3992 7753 3996 7757
rect 4046 7753 4050 7757
rect 4077 7753 4081 7757
rect 4106 7753 4110 7757
rect 4131 7753 4135 7757
rect 4173 7753 4177 7757
rect 3180 7711 3184 7715
rect 3208 7711 3212 7715
rect 3238 7711 3242 7715
rect 3275 7711 3279 7715
rect 4125 7711 4129 7715
rect 4153 7711 4157 7715
rect 4183 7711 4187 7715
rect 4220 7711 4224 7715
rect 2397 7681 2401 7685
rect 2425 7681 2429 7685
rect 2455 7681 2459 7685
rect 2492 7681 2496 7685
rect 2529 7681 2533 7685
rect 2557 7681 2561 7685
rect 2587 7681 2591 7685
rect 2624 7681 2628 7685
rect 2661 7681 2665 7685
rect 2689 7681 2693 7685
rect 2719 7681 2723 7685
rect 2756 7681 2760 7685
rect 3342 7681 3346 7685
rect 3370 7681 3374 7685
rect 3400 7681 3404 7685
rect 3437 7681 3441 7685
rect 3474 7681 3478 7685
rect 3502 7681 3506 7685
rect 3532 7681 3536 7685
rect 3569 7681 3573 7685
rect 3606 7681 3610 7685
rect 3634 7681 3638 7685
rect 3664 7681 3668 7685
rect 3701 7681 3705 7685
rect 3180 7625 3184 7629
rect 3208 7625 3212 7629
rect 3238 7625 3242 7629
rect 3275 7625 3279 7629
rect 4125 7625 4129 7629
rect 4153 7625 4157 7629
rect 4183 7625 4187 7629
rect 4220 7625 4224 7629
rect 2397 7595 2401 7599
rect 2425 7595 2429 7599
rect 2455 7595 2459 7599
rect 2492 7595 2496 7599
rect 2529 7595 2533 7599
rect 2557 7595 2561 7599
rect 2587 7595 2591 7599
rect 2624 7595 2628 7599
rect 2661 7595 2665 7599
rect 2689 7595 2693 7599
rect 2719 7595 2723 7599
rect 2756 7595 2760 7599
rect 3342 7595 3346 7599
rect 3370 7595 3374 7599
rect 3400 7595 3404 7599
rect 3437 7595 3441 7599
rect 3474 7595 3478 7599
rect 3502 7595 3506 7599
rect 3532 7595 3536 7599
rect 3569 7595 3573 7599
rect 3606 7595 3610 7599
rect 3634 7595 3638 7599
rect 3664 7595 3668 7599
rect 3701 7595 3705 7599
rect 2397 7455 2401 7459
rect 2425 7455 2429 7459
rect 2455 7455 2459 7459
rect 2492 7455 2496 7459
rect 2529 7455 2533 7459
rect 2557 7455 2561 7459
rect 2587 7455 2591 7459
rect 2624 7455 2628 7459
rect 2661 7455 2665 7459
rect 2689 7455 2693 7459
rect 2719 7455 2723 7459
rect 2756 7455 2760 7459
rect 3342 7455 3346 7459
rect 3370 7455 3374 7459
rect 3400 7455 3404 7459
rect 3437 7455 3441 7459
rect 3474 7455 3478 7459
rect 3502 7455 3506 7459
rect 3532 7455 3536 7459
rect 3569 7455 3573 7459
rect 3606 7455 3610 7459
rect 3634 7455 3638 7459
rect 3664 7455 3668 7459
rect 3701 7455 3705 7459
rect 1467 6855 1471 6859
rect 1504 6855 1508 6859
rect 1534 6855 1538 6859
rect 1562 6855 1566 6859
rect 1599 6855 1603 6859
rect 1636 6855 1640 6859
rect 1666 6855 1670 6859
rect 1694 6855 1698 6859
rect 1731 6855 1735 6859
rect 1768 6855 1772 6859
rect 1798 6855 1802 6859
rect 1826 6855 1830 6859
rect 2412 6855 2416 6859
rect 2449 6855 2453 6859
rect 2479 6855 2483 6859
rect 2507 6855 2511 6859
rect 2544 6855 2548 6859
rect 2581 6855 2585 6859
rect 2611 6855 2615 6859
rect 2639 6855 2643 6859
rect 2676 6855 2680 6859
rect 2713 6855 2717 6859
rect 2743 6855 2747 6859
rect 2771 6855 2775 6859
rect 1467 6715 1471 6719
rect 1504 6715 1508 6719
rect 1534 6715 1538 6719
rect 1562 6715 1566 6719
rect 1599 6715 1603 6719
rect 1636 6715 1640 6719
rect 1666 6715 1670 6719
rect 1694 6715 1698 6719
rect 1731 6715 1735 6719
rect 1768 6715 1772 6719
rect 1798 6715 1802 6719
rect 1826 6715 1830 6719
rect 2412 6715 2416 6719
rect 2449 6715 2453 6719
rect 2479 6715 2483 6719
rect 2507 6715 2511 6719
rect 2544 6715 2548 6719
rect 2581 6715 2585 6719
rect 2611 6715 2615 6719
rect 2639 6715 2643 6719
rect 2676 6715 2680 6719
rect 2713 6715 2717 6719
rect 2743 6715 2747 6719
rect 2771 6715 2775 6719
rect 948 6685 952 6689
rect 985 6685 989 6689
rect 1015 6685 1019 6689
rect 1043 6685 1047 6689
rect 1893 6685 1897 6689
rect 1930 6685 1934 6689
rect 1960 6685 1964 6689
rect 1988 6685 1992 6689
rect 1467 6629 1471 6633
rect 1504 6629 1508 6633
rect 1534 6629 1538 6633
rect 1562 6629 1566 6633
rect 1599 6629 1603 6633
rect 1636 6629 1640 6633
rect 1666 6629 1670 6633
rect 1694 6629 1698 6633
rect 1731 6629 1735 6633
rect 1768 6629 1772 6633
rect 1798 6629 1802 6633
rect 1826 6629 1830 6633
rect 2412 6629 2416 6633
rect 2449 6629 2453 6633
rect 2479 6629 2483 6633
rect 2507 6629 2511 6633
rect 2544 6629 2548 6633
rect 2581 6629 2585 6633
rect 2611 6629 2615 6633
rect 2639 6629 2643 6633
rect 2676 6629 2680 6633
rect 2713 6629 2717 6633
rect 2743 6629 2747 6633
rect 2771 6629 2775 6633
rect 948 6599 952 6603
rect 985 6599 989 6603
rect 1015 6599 1019 6603
rect 1043 6599 1047 6603
rect 1893 6599 1897 6603
rect 1930 6599 1934 6603
rect 1960 6599 1964 6603
rect 1988 6599 1992 6603
rect 995 6557 999 6561
rect 1037 6557 1041 6561
rect 1062 6557 1066 6561
rect 1091 6557 1095 6561
rect 1122 6557 1126 6561
rect 1176 6557 1180 6561
rect 1256 6557 1260 6561
rect 1298 6557 1302 6561
rect 1323 6557 1327 6561
rect 1352 6557 1356 6561
rect 1940 6557 1944 6561
rect 1982 6557 1986 6561
rect 2007 6557 2011 6561
rect 2036 6557 2040 6561
rect 2067 6557 2071 6561
rect 2121 6557 2125 6561
rect 2201 6557 2205 6561
rect 2243 6557 2247 6561
rect 2268 6557 2272 6561
rect 2297 6557 2301 6561
rect 1467 6487 1471 6491
rect 1504 6487 1508 6491
rect 1534 6487 1538 6491
rect 1562 6487 1566 6491
rect 1599 6487 1603 6491
rect 1636 6487 1640 6491
rect 1666 6487 1670 6491
rect 1694 6487 1698 6491
rect 1731 6487 1735 6491
rect 1768 6487 1772 6491
rect 1798 6487 1802 6491
rect 1826 6487 1830 6491
rect 2412 6487 2416 6491
rect 2449 6487 2453 6491
rect 2479 6487 2483 6491
rect 2507 6487 2511 6491
rect 2544 6487 2548 6491
rect 2581 6487 2585 6491
rect 2611 6487 2615 6491
rect 2639 6487 2643 6491
rect 2676 6487 2680 6491
rect 2713 6487 2717 6491
rect 2743 6487 2747 6491
rect 2771 6487 2775 6491
rect 1005 6425 1009 6429
rect 1095 6425 1099 6429
rect 1122 6425 1126 6429
rect 1176 6425 1180 6429
rect 1200 6425 1204 6429
rect 1256 6425 1260 6429
rect 1298 6425 1302 6429
rect 1323 6425 1327 6429
rect 1352 6425 1356 6429
rect 1950 6425 1954 6429
rect 2040 6425 2044 6429
rect 2067 6425 2071 6429
rect 2121 6425 2125 6429
rect 2145 6425 2149 6429
rect 2201 6425 2205 6429
rect 2243 6425 2247 6429
rect 2268 6425 2272 6429
rect 2297 6425 2301 6429
rect 951 6293 955 6297
rect 1005 6293 1009 6297
rect 1033 6293 1037 6297
rect 1041 6293 1045 6297
rect 1095 6293 1099 6297
rect 1122 6293 1126 6297
rect 1176 6293 1180 6297
rect 1200 6293 1204 6297
rect 1256 6293 1260 6297
rect 1298 6293 1302 6297
rect 1323 6293 1327 6297
rect 1352 6293 1356 6297
rect 1896 6293 1900 6297
rect 1950 6293 1954 6297
rect 1978 6293 1982 6297
rect 1986 6293 1990 6297
rect 2040 6293 2044 6297
rect 2067 6293 2071 6297
rect 2121 6293 2125 6297
rect 2145 6293 2149 6297
rect 2201 6293 2205 6297
rect 2243 6293 2247 6297
rect 2268 6293 2272 6297
rect 2297 6293 2301 6297
rect 1033 6161 1037 6165
rect 1095 6161 1099 6165
rect 1122 6161 1126 6165
rect 1176 6161 1180 6165
rect 1200 6161 1204 6165
rect 1256 6161 1260 6165
rect 1298 6161 1302 6165
rect 1323 6161 1327 6165
rect 1352 6161 1356 6165
rect 1978 6161 1982 6165
rect 2040 6161 2044 6165
rect 2067 6161 2071 6165
rect 2121 6161 2125 6165
rect 2145 6161 2149 6165
rect 2201 6161 2205 6165
rect 2243 6161 2247 6165
rect 2268 6161 2272 6165
rect 2297 6161 2301 6165
rect 1639 6087 1643 6091
rect 1667 6087 1671 6091
rect 1697 6087 1701 6091
rect 1734 6087 1738 6091
rect 2584 6087 2588 6091
rect 2612 6087 2616 6091
rect 2642 6087 2646 6091
rect 2679 6087 2683 6091
rect 1041 6029 1045 6033
rect 1095 6029 1099 6033
rect 1122 6029 1126 6033
rect 1176 6029 1180 6033
rect 1200 6029 1204 6033
rect 1256 6029 1260 6033
rect 1298 6029 1302 6033
rect 1323 6029 1327 6033
rect 1352 6029 1356 6033
rect 1986 6029 1990 6033
rect 2040 6029 2044 6033
rect 2067 6029 2071 6033
rect 2121 6029 2125 6033
rect 2145 6029 2149 6033
rect 2201 6029 2205 6033
rect 2243 6029 2247 6033
rect 2268 6029 2272 6033
rect 2297 6029 2301 6033
rect 1599 5985 1603 5989
rect 1636 5985 1640 5989
rect 1666 5985 1670 5989
rect 1694 5985 1698 5989
rect 2544 5985 2548 5989
rect 2581 5985 2585 5989
rect 2611 5985 2615 5989
rect 2639 5985 2643 5989
rect 851 5952 855 5956
rect 888 5952 892 5956
rect 918 5952 922 5956
rect 946 5952 950 5956
rect 983 5952 987 5956
rect 1020 5952 1024 5956
rect 1050 5952 1054 5956
rect 1078 5952 1082 5956
rect 1115 5952 1119 5956
rect 1152 5952 1156 5956
rect 1182 5952 1186 5956
rect 1210 5952 1214 5956
rect 1247 5952 1251 5956
rect 1284 5952 1288 5956
rect 1314 5952 1318 5956
rect 1342 5952 1346 5956
rect 1796 5952 1800 5956
rect 1833 5952 1837 5956
rect 1863 5952 1867 5956
rect 1891 5952 1895 5956
rect 1928 5952 1932 5956
rect 1965 5952 1969 5956
rect 1995 5952 1999 5956
rect 2023 5952 2027 5956
rect 2060 5952 2064 5956
rect 2097 5952 2101 5956
rect 2127 5952 2131 5956
rect 2155 5952 2159 5956
rect 2192 5952 2196 5956
rect 2229 5952 2233 5956
rect 2259 5952 2263 5956
rect 2287 5952 2291 5956
rect 1467 5873 1471 5877
rect 1504 5873 1508 5877
rect 1534 5873 1538 5877
rect 1562 5873 1566 5877
rect 1599 5873 1603 5877
rect 1636 5873 1640 5877
rect 1666 5873 1670 5877
rect 1694 5873 1698 5877
rect 1731 5873 1735 5877
rect 1768 5873 1772 5877
rect 1798 5873 1802 5877
rect 1826 5873 1830 5877
rect 2412 5873 2416 5877
rect 2449 5873 2453 5877
rect 2479 5873 2483 5877
rect 2507 5873 2511 5877
rect 2544 5873 2548 5877
rect 2581 5873 2585 5877
rect 2611 5873 2615 5877
rect 2639 5873 2643 5877
rect 2676 5873 2680 5877
rect 2713 5873 2717 5877
rect 2743 5873 2747 5877
rect 2771 5873 2775 5877
rect 1467 5733 1471 5737
rect 1504 5733 1508 5737
rect 1534 5733 1538 5737
rect 1562 5733 1566 5737
rect 1599 5733 1603 5737
rect 1636 5733 1640 5737
rect 1666 5733 1670 5737
rect 1694 5733 1698 5737
rect 1731 5733 1735 5737
rect 1768 5733 1772 5737
rect 1798 5733 1802 5737
rect 1826 5733 1830 5737
rect 2412 5733 2416 5737
rect 2449 5733 2453 5737
rect 2479 5733 2483 5737
rect 2507 5733 2511 5737
rect 2544 5733 2548 5737
rect 2581 5733 2585 5737
rect 2611 5733 2615 5737
rect 2639 5733 2643 5737
rect 2676 5733 2680 5737
rect 2713 5733 2717 5737
rect 2743 5733 2747 5737
rect 2771 5733 2775 5737
rect 948 5703 952 5707
rect 985 5703 989 5707
rect 1015 5703 1019 5707
rect 1043 5703 1047 5707
rect 1893 5703 1897 5707
rect 1930 5703 1934 5707
rect 1960 5703 1964 5707
rect 1988 5703 1992 5707
rect 1467 5647 1471 5651
rect 1504 5647 1508 5651
rect 1534 5647 1538 5651
rect 1562 5647 1566 5651
rect 1599 5647 1603 5651
rect 1636 5647 1640 5651
rect 1666 5647 1670 5651
rect 1694 5647 1698 5651
rect 1731 5647 1735 5651
rect 1768 5647 1772 5651
rect 1798 5647 1802 5651
rect 1826 5647 1830 5651
rect 2412 5647 2416 5651
rect 2449 5647 2453 5651
rect 2479 5647 2483 5651
rect 2507 5647 2511 5651
rect 2544 5647 2548 5651
rect 2581 5647 2585 5651
rect 2611 5647 2615 5651
rect 2639 5647 2643 5651
rect 2676 5647 2680 5651
rect 2713 5647 2717 5651
rect 2743 5647 2747 5651
rect 2771 5647 2775 5651
rect 948 5617 952 5621
rect 985 5617 989 5621
rect 1015 5617 1019 5621
rect 1043 5617 1047 5621
rect 1893 5617 1897 5621
rect 1930 5617 1934 5621
rect 1960 5617 1964 5621
rect 1988 5617 1992 5621
rect 995 5575 999 5579
rect 1037 5575 1041 5579
rect 1062 5575 1066 5579
rect 1091 5575 1095 5579
rect 1122 5575 1126 5579
rect 1176 5575 1180 5579
rect 1256 5575 1260 5579
rect 1298 5575 1302 5579
rect 1323 5575 1327 5579
rect 1352 5575 1356 5579
rect 1940 5575 1944 5579
rect 1982 5575 1986 5579
rect 2007 5575 2011 5579
rect 2036 5575 2040 5579
rect 2067 5575 2071 5579
rect 2121 5575 2125 5579
rect 2201 5575 2205 5579
rect 2243 5575 2247 5579
rect 2268 5575 2272 5579
rect 2297 5575 2301 5579
rect 1467 5505 1471 5509
rect 1504 5505 1508 5509
rect 1534 5505 1538 5509
rect 1562 5505 1566 5509
rect 1599 5505 1603 5509
rect 1636 5505 1640 5509
rect 1666 5505 1670 5509
rect 1694 5505 1698 5509
rect 1731 5505 1735 5509
rect 1768 5505 1772 5509
rect 1798 5505 1802 5509
rect 1826 5505 1830 5509
rect 2412 5505 2416 5509
rect 2449 5505 2453 5509
rect 2479 5505 2483 5509
rect 2507 5505 2511 5509
rect 2544 5505 2548 5509
rect 2581 5505 2585 5509
rect 2611 5505 2615 5509
rect 2639 5505 2643 5509
rect 2676 5505 2680 5509
rect 2713 5505 2717 5509
rect 2743 5505 2747 5509
rect 2771 5505 2775 5509
rect 1785 5468 1789 5472
rect 1005 5443 1009 5447
rect 1095 5443 1099 5447
rect 1122 5443 1126 5447
rect 1176 5443 1180 5447
rect 1200 5443 1204 5447
rect 1256 5443 1260 5447
rect 1298 5443 1302 5447
rect 1323 5443 1327 5447
rect 1352 5443 1356 5447
rect 1950 5443 1954 5447
rect 2040 5443 2044 5447
rect 2067 5443 2071 5447
rect 2121 5443 2125 5447
rect 2145 5443 2149 5447
rect 2201 5443 2205 5447
rect 2243 5443 2247 5447
rect 2268 5443 2272 5447
rect 2297 5443 2301 5447
rect 1682 5338 1686 5342
rect 1731 5338 1735 5342
rect 1785 5338 1789 5342
rect 1809 5338 1813 5342
rect 1831 5338 1835 5342
rect 951 5311 955 5315
rect 1005 5311 1009 5315
rect 1033 5311 1037 5315
rect 1041 5311 1045 5315
rect 1095 5311 1099 5315
rect 1122 5311 1126 5315
rect 1176 5311 1180 5315
rect 1200 5311 1204 5315
rect 1256 5311 1260 5315
rect 1298 5311 1302 5315
rect 1323 5311 1327 5315
rect 1352 5311 1356 5315
rect 1896 5311 1900 5315
rect 1950 5311 1954 5315
rect 1978 5311 1982 5315
rect 1986 5311 1990 5315
rect 2040 5311 2044 5315
rect 2067 5311 2071 5315
rect 2121 5311 2125 5315
rect 2145 5311 2149 5315
rect 2201 5311 2205 5315
rect 2243 5311 2247 5315
rect 2268 5311 2272 5315
rect 2297 5311 2301 5315
rect 1588 5208 1592 5212
rect 1731 5208 1735 5212
rect 1785 5208 1789 5212
rect 1809 5208 1813 5212
rect 1033 5179 1037 5183
rect 1095 5179 1099 5183
rect 1122 5179 1126 5183
rect 1176 5179 1180 5183
rect 1200 5179 1204 5183
rect 1256 5179 1260 5183
rect 1298 5179 1302 5183
rect 1323 5179 1327 5183
rect 1352 5179 1356 5183
rect 1978 5179 1982 5183
rect 2040 5179 2044 5183
rect 2067 5179 2071 5183
rect 2121 5179 2125 5183
rect 2145 5179 2149 5183
rect 2201 5179 2205 5183
rect 2243 5179 2247 5183
rect 2268 5179 2272 5183
rect 2297 5179 2301 5183
rect 1639 5105 1643 5109
rect 1667 5105 1671 5109
rect 1697 5105 1701 5109
rect 1734 5105 1738 5109
rect 2584 5105 2588 5109
rect 2612 5105 2616 5109
rect 2642 5105 2646 5109
rect 2679 5105 2683 5109
rect 1041 5047 1045 5051
rect 1095 5047 1099 5051
rect 1122 5047 1126 5051
rect 1176 5047 1180 5051
rect 1200 5047 1204 5051
rect 1256 5047 1260 5051
rect 1298 5047 1302 5051
rect 1323 5047 1327 5051
rect 1352 5047 1356 5051
rect 1986 5047 1990 5051
rect 2040 5047 2044 5051
rect 2067 5047 2071 5051
rect 2121 5047 2125 5051
rect 2145 5047 2149 5051
rect 2201 5047 2205 5051
rect 2243 5047 2247 5051
rect 2268 5047 2272 5051
rect 2297 5047 2301 5051
rect 1599 5003 1603 5007
rect 1636 5003 1640 5007
rect 1666 5003 1670 5007
rect 1694 5003 1698 5007
rect 2544 5003 2548 5007
rect 2581 5003 2585 5007
rect 2611 5003 2615 5007
rect 2639 5003 2643 5007
rect 851 4970 855 4974
rect 888 4970 892 4974
rect 918 4970 922 4974
rect 946 4970 950 4974
rect 983 4970 987 4974
rect 1020 4970 1024 4974
rect 1050 4970 1054 4974
rect 1078 4970 1082 4974
rect 1115 4970 1119 4974
rect 1152 4970 1156 4974
rect 1182 4970 1186 4974
rect 1210 4970 1214 4974
rect 1247 4970 1251 4974
rect 1284 4970 1288 4974
rect 1314 4970 1318 4974
rect 1342 4970 1346 4974
rect 1796 4970 1800 4974
rect 1833 4970 1837 4974
rect 1863 4970 1867 4974
rect 1891 4970 1895 4974
rect 1928 4970 1932 4974
rect 1965 4970 1969 4974
rect 1995 4970 1999 4974
rect 2023 4970 2027 4974
rect 2060 4970 2064 4974
rect 2097 4970 2101 4974
rect 2127 4970 2131 4974
rect 2155 4970 2159 4974
rect 2192 4970 2196 4974
rect 2229 4970 2233 4974
rect 2259 4970 2263 4974
rect 2287 4970 2291 4974
rect 4525 9573 4529 9577
rect 4535 9573 4539 9577
rect 4545 9573 4549 9577
rect 4555 9573 4559 9577
rect 4525 9568 4529 9572
rect 4535 9568 4539 9572
rect 4545 9568 4549 9572
rect 4555 9568 4559 9572
rect 4525 9563 4529 9567
rect 4535 9563 4539 9567
rect 4545 9563 4549 9567
rect 4555 9563 4559 9567
rect 4525 9558 4529 9562
rect 4535 9558 4539 9562
rect 4545 9558 4549 9562
rect 4555 9558 4559 9562
rect 4525 9544 4529 9548
rect 4535 9544 4539 9548
rect 4545 9544 4549 9548
rect 4555 9544 4559 9548
rect 4525 9539 4529 9543
rect 4535 9539 4539 9543
rect 4545 9539 4549 9543
rect 4555 9539 4559 9543
rect 4525 9534 4529 9538
rect 4535 9534 4539 9538
rect 4545 9534 4549 9538
rect 4555 9534 4559 9538
rect 4525 9529 4529 9533
rect 4535 9529 4539 9533
rect 4545 9529 4549 9533
rect 4555 9529 4559 9533
rect 4525 9515 4529 9519
rect 4535 9515 4539 9519
rect 4545 9515 4549 9519
rect 4555 9515 4559 9519
rect 4525 9510 4529 9514
rect 4535 9510 4539 9514
rect 4545 9510 4549 9514
rect 4555 9510 4559 9514
rect 4525 9505 4529 9509
rect 4535 9505 4539 9509
rect 4545 9505 4549 9509
rect 4555 9505 4559 9509
rect 4525 9500 4529 9504
rect 4535 9500 4539 9504
rect 4545 9500 4549 9504
rect 4555 9500 4559 9504
rect 4525 9486 4529 9490
rect 4535 9486 4539 9490
rect 4545 9486 4549 9490
rect 4555 9486 4559 9490
rect 4525 9481 4529 9485
rect 4535 9481 4539 9485
rect 4545 9481 4549 9485
rect 4555 9481 4559 9485
rect 4525 9476 4529 9480
rect 4535 9476 4539 9480
rect 4545 9476 4549 9480
rect 4555 9476 4559 9480
rect 4525 9471 4529 9475
rect 4535 9471 4539 9475
rect 4545 9471 4549 9475
rect 4555 9471 4559 9475
rect 4525 9457 4529 9461
rect 4535 9457 4539 9461
rect 4545 9457 4549 9461
rect 4555 9457 4559 9461
rect 4525 9452 4529 9456
rect 4535 9452 4539 9456
rect 4545 9452 4549 9456
rect 4555 9452 4559 9456
rect 4525 9447 4529 9451
rect 4535 9447 4539 9451
rect 4545 9447 4549 9451
rect 4555 9447 4559 9451
rect 4525 9442 4529 9446
rect 4535 9442 4539 9446
rect 4545 9442 4549 9446
rect 4555 9442 4559 9446
rect 4525 9056 4529 9060
rect 4535 9056 4539 9060
rect 4545 9056 4549 9060
rect 4555 9056 4559 9060
rect 4525 9051 4529 9055
rect 4535 9051 4539 9055
rect 4545 9051 4549 9055
rect 4555 9051 4559 9055
rect 4525 9046 4529 9050
rect 4535 9046 4539 9050
rect 4545 9046 4549 9050
rect 4555 9046 4559 9050
rect 4525 9041 4529 9045
rect 4535 9041 4539 9045
rect 4545 9041 4549 9045
rect 4555 9041 4559 9045
rect 4525 8747 4529 8751
rect 4535 8747 4539 8751
rect 4545 8747 4549 8751
rect 4555 8747 4559 8751
rect 4525 8742 4529 8746
rect 4535 8742 4539 8746
rect 4545 8742 4549 8746
rect 4555 8742 4559 8746
rect 4525 8737 4529 8741
rect 4535 8737 4539 8741
rect 4545 8737 4549 8741
rect 4555 8737 4559 8741
rect 4525 8732 4529 8736
rect 4535 8732 4539 8736
rect 4545 8732 4549 8736
rect 4555 8732 4559 8736
rect 4525 8438 4529 8442
rect 4535 8438 4539 8442
rect 4545 8438 4549 8442
rect 4555 8438 4559 8442
rect 4525 8433 4529 8437
rect 4535 8433 4539 8437
rect 4545 8433 4549 8437
rect 4555 8433 4559 8437
rect 4525 8428 4529 8432
rect 4535 8428 4539 8432
rect 4545 8428 4549 8432
rect 4555 8428 4559 8432
rect 4525 8423 4529 8427
rect 4535 8423 4539 8427
rect 4545 8423 4549 8427
rect 4555 8423 4559 8427
rect 4525 8129 4529 8133
rect 4535 8129 4539 8133
rect 4545 8129 4549 8133
rect 4555 8129 4559 8133
rect 4525 8124 4529 8128
rect 4535 8124 4539 8128
rect 4545 8124 4549 8128
rect 4555 8124 4559 8128
rect 4525 8119 4529 8123
rect 4535 8119 4539 8123
rect 4545 8119 4549 8123
rect 4555 8119 4559 8123
rect 4525 8114 4529 8118
rect 4535 8114 4539 8118
rect 4545 8114 4549 8118
rect 4555 8114 4559 8118
rect 4525 8098 4529 8102
rect 4535 8098 4539 8102
rect 4545 8098 4549 8102
rect 4555 8098 4559 8102
rect 4525 8093 4529 8097
rect 4535 8093 4539 8097
rect 4545 8093 4549 8097
rect 4555 8093 4559 8097
rect 4525 8088 4529 8092
rect 4535 8088 4539 8092
rect 4545 8088 4549 8092
rect 4555 8088 4559 8092
rect 4525 8083 4529 8087
rect 4535 8083 4539 8087
rect 4545 8083 4549 8087
rect 4555 8083 4559 8087
rect 4627 7889 4631 7945
rect 4666 7857 4670 7945
rect 4709 7857 4713 7945
rect 4750 7857 4754 7945
rect 4525 7789 4529 7793
rect 4535 7789 4539 7793
rect 4545 7789 4549 7793
rect 4555 7789 4559 7793
rect 4525 7784 4529 7788
rect 4535 7784 4539 7788
rect 4545 7784 4549 7788
rect 4555 7784 4559 7788
rect 4525 7779 4529 7783
rect 4535 7779 4539 7783
rect 4545 7779 4549 7783
rect 4555 7779 4559 7783
rect 4525 7774 4529 7778
rect 4535 7774 4539 7778
rect 4545 7774 4549 7778
rect 4555 7774 4559 7778
rect 4632 7486 4636 7490
rect 4637 7486 4641 7490
rect 4642 7486 4646 7490
rect 4647 7486 4651 7490
rect 4652 7486 4656 7490
rect 4657 7486 4661 7490
rect 4662 7486 4666 7490
rect 4667 7486 4671 7490
rect 4672 7486 4676 7490
rect 4677 7486 4681 7490
rect 4682 7486 4686 7490
rect 4687 7486 4691 7490
rect 4692 7486 4696 7490
rect 4697 7486 4701 7490
rect 4702 7486 4706 7490
rect 4707 7486 4711 7490
rect 4712 7486 4716 7490
rect 4717 7486 4721 7490
rect 4722 7486 4726 7490
rect 4727 7486 4731 7490
rect 4732 7486 4736 7490
rect 4737 7486 4741 7490
rect 4742 7486 4746 7490
rect 4747 7486 4751 7490
rect 4752 7486 4756 7490
rect 4757 7486 4761 7490
rect 4762 7486 4766 7490
rect 4767 7486 4771 7490
rect 4632 7481 4636 7485
rect 4632 7476 4636 7480
rect 4767 7481 4771 7485
rect 4632 7471 4636 7475
rect 4632 7466 4636 7470
rect 4632 7461 4636 7465
rect 4632 7456 4636 7460
rect 4632 7451 4636 7455
rect 4632 7446 4636 7450
rect 4632 7441 4636 7445
rect 4632 7436 4636 7440
rect 4632 7431 4636 7435
rect 4632 7426 4636 7430
rect 4632 7421 4636 7425
rect 4632 7416 4636 7420
rect 4632 7411 4636 7415
rect 4632 7406 4636 7410
rect 4767 7476 4771 7480
rect 4767 7471 4771 7475
rect 4767 7466 4771 7470
rect 4767 7461 4771 7465
rect 4767 7456 4771 7460
rect 4767 7451 4771 7455
rect 4767 7446 4771 7450
rect 4767 7441 4771 7445
rect 4767 7436 4771 7440
rect 4767 7431 4771 7435
rect 4767 7426 4771 7430
rect 4767 7421 4771 7425
rect 4767 7416 4771 7420
rect 4767 7411 4771 7415
rect 4632 7401 4636 7405
rect 4767 7406 4771 7410
rect 4767 7401 4771 7405
rect 4632 7396 4636 7400
rect 4637 7396 4641 7400
rect 4642 7396 4646 7400
rect 4647 7396 4651 7400
rect 4652 7396 4656 7400
rect 4657 7396 4661 7400
rect 4662 7396 4666 7400
rect 4667 7396 4671 7400
rect 4672 7396 4676 7400
rect 4677 7396 4681 7400
rect 4682 7396 4686 7400
rect 4687 7396 4691 7400
rect 4692 7396 4696 7400
rect 4697 7396 4701 7400
rect 4702 7396 4706 7400
rect 4707 7396 4711 7400
rect 4712 7396 4716 7400
rect 4717 7396 4721 7400
rect 4722 7396 4726 7400
rect 4727 7396 4731 7400
rect 4732 7396 4736 7400
rect 4737 7396 4741 7400
rect 4742 7396 4746 7400
rect 4747 7396 4751 7400
rect 4752 7396 4756 7400
rect 4757 7396 4761 7400
rect 4762 7396 4766 7400
rect 4767 7396 4771 7400
rect 4645 7313 4649 7317
rect 4652 7313 4656 7317
rect 4657 7313 4661 7317
rect 4662 7313 4666 7317
rect 4667 7313 4671 7317
rect 4672 7313 4676 7317
rect 4677 7313 4681 7317
rect 4682 7313 4686 7317
rect 4687 7313 4691 7317
rect 4692 7313 4696 7317
rect 4697 7313 4701 7317
rect 4702 7313 4706 7317
rect 4707 7313 4711 7317
rect 4712 7313 4716 7317
rect 4717 7313 4721 7317
rect 4722 7313 4726 7317
rect 4727 7313 4731 7317
rect 4732 7313 4736 7317
rect 4737 7313 4741 7317
rect 4742 7313 4746 7317
rect 4747 7313 4751 7317
rect 4754 7313 4758 7317
rect 4645 7306 4649 7310
rect 4754 7306 4758 7310
rect 4645 7301 4649 7305
rect 4645 7296 4649 7300
rect 4645 7291 4649 7295
rect 4645 7286 4649 7290
rect 4645 7281 4649 7285
rect 4645 7276 4649 7280
rect 4645 7271 4649 7275
rect 4645 7266 4649 7270
rect 4645 7261 4649 7265
rect 4754 7301 4758 7305
rect 4754 7296 4758 7300
rect 4754 7291 4758 7295
rect 4754 7286 4758 7290
rect 4754 7281 4758 7285
rect 4754 7276 4758 7280
rect 4754 7271 4758 7275
rect 4754 7266 4758 7270
rect 4754 7261 4758 7265
rect 4645 7256 4649 7260
rect 4754 7256 4758 7260
rect 4645 7249 4649 7253
rect 4652 7249 4656 7253
rect 4657 7249 4661 7253
rect 4662 7249 4666 7253
rect 4667 7249 4671 7253
rect 4672 7249 4676 7253
rect 4677 7249 4681 7253
rect 4682 7249 4686 7253
rect 4687 7249 4691 7253
rect 4692 7249 4696 7253
rect 4697 7249 4701 7253
rect 4702 7249 4706 7253
rect 4707 7249 4711 7253
rect 4712 7249 4716 7253
rect 4717 7249 4721 7253
rect 4722 7249 4726 7253
rect 4727 7249 4731 7253
rect 4732 7249 4736 7253
rect 4737 7249 4741 7253
rect 4742 7249 4746 7253
rect 4747 7249 4751 7253
rect 4754 7249 4758 7253
rect 4525 7230 4529 7234
rect 4535 7230 4539 7234
rect 4545 7230 4549 7234
rect 4555 7230 4559 7234
rect 4525 7225 4529 7229
rect 4535 7225 4539 7229
rect 4545 7225 4549 7229
rect 4555 7225 4559 7229
rect 4525 7220 4529 7224
rect 4535 7220 4539 7224
rect 4545 7220 4549 7224
rect 4555 7220 4559 7224
rect 4525 7215 4529 7219
rect 4535 7215 4539 7219
rect 4545 7215 4549 7219
rect 4555 7215 4559 7219
rect 4525 7202 4529 7206
rect 4535 7202 4539 7206
rect 4545 7202 4549 7206
rect 4555 7202 4559 7206
rect 4525 7197 4529 7201
rect 4535 7197 4539 7201
rect 4545 7197 4549 7201
rect 4555 7197 4559 7201
rect 4525 7192 4529 7196
rect 4535 7192 4539 7196
rect 4545 7192 4549 7196
rect 4555 7192 4559 7196
rect 4525 7187 4529 7191
rect 4535 7187 4539 7191
rect 4545 7187 4549 7191
rect 4555 7187 4559 7191
rect 4525 7152 4529 7156
rect 4535 7152 4539 7156
rect 4545 7152 4549 7156
rect 4555 7152 4559 7156
rect 4525 6858 4529 6862
rect 4535 6858 4539 6862
rect 4545 6858 4549 6862
rect 4555 6858 4559 6862
rect 4525 6853 4529 6857
rect 4535 6853 4539 6857
rect 4545 6853 4549 6857
rect 4555 6853 4559 6857
rect 4525 6848 4529 6852
rect 4535 6848 4539 6852
rect 4545 6848 4549 6852
rect 4555 6848 4559 6852
rect 4525 6843 4529 6847
rect 4535 6843 4539 6847
rect 4545 6843 4549 6847
rect 4555 6843 4559 6847
rect 4525 6549 4529 6553
rect 4535 6549 4539 6553
rect 4545 6549 4549 6553
rect 4555 6549 4559 6553
rect 4525 6544 4529 6548
rect 4535 6544 4539 6548
rect 4545 6544 4549 6548
rect 4555 6544 4559 6548
rect 4525 6539 4529 6543
rect 4535 6539 4539 6543
rect 4545 6539 4549 6543
rect 4555 6539 4559 6543
rect 4525 6534 4529 6538
rect 4535 6534 4539 6538
rect 4545 6534 4549 6538
rect 4555 6534 4559 6538
rect 4525 6240 4529 6244
rect 4535 6240 4539 6244
rect 4545 6240 4549 6244
rect 4555 6240 4559 6244
rect 4525 6235 4529 6239
rect 4535 6235 4539 6239
rect 4545 6235 4549 6239
rect 4555 6235 4559 6239
rect 4525 6230 4529 6234
rect 4535 6230 4539 6234
rect 4545 6230 4549 6234
rect 4555 6230 4559 6234
rect 4525 6225 4529 6229
rect 4535 6225 4539 6229
rect 4545 6225 4549 6229
rect 4555 6225 4559 6229
rect 4525 5931 4529 5935
rect 4535 5931 4539 5935
rect 4545 5931 4549 5935
rect 4555 5931 4559 5935
rect 4525 5926 4529 5930
rect 4535 5926 4539 5930
rect 4545 5926 4549 5930
rect 4555 5926 4559 5930
rect 4525 5921 4529 5925
rect 4535 5921 4539 5925
rect 4545 5921 4549 5925
rect 4555 5921 4559 5925
rect 4525 5916 4529 5920
rect 4535 5916 4539 5920
rect 4545 5916 4549 5920
rect 4555 5916 4559 5920
rect 4525 5622 4529 5626
rect 4535 5622 4539 5626
rect 4545 5622 4549 5626
rect 4555 5622 4559 5626
rect 4525 5617 4529 5621
rect 4535 5617 4539 5621
rect 4545 5617 4549 5621
rect 4555 5617 4559 5621
rect 4525 5612 4529 5616
rect 4535 5612 4539 5616
rect 4545 5612 4549 5616
rect 4555 5612 4559 5616
rect 4525 5607 4529 5611
rect 4535 5607 4539 5611
rect 4545 5607 4549 5611
rect 4555 5607 4559 5611
rect 4525 5313 4529 5317
rect 4535 5313 4539 5317
rect 4545 5313 4549 5317
rect 4555 5313 4559 5317
rect 4525 5308 4529 5312
rect 4535 5308 4539 5312
rect 4545 5308 4549 5312
rect 4555 5308 4559 5312
rect 4525 5303 4529 5307
rect 4535 5303 4539 5307
rect 4545 5303 4549 5307
rect 4555 5303 4559 5307
rect 4525 5298 4529 5302
rect 4535 5298 4539 5302
rect 4545 5298 4549 5302
rect 4555 5298 4559 5302
rect 4525 5004 4529 5008
rect 4535 5004 4539 5008
rect 4545 5004 4549 5008
rect 4555 5004 4559 5008
rect 4525 4999 4529 5003
rect 4535 4999 4539 5003
rect 4545 4999 4549 5003
rect 4555 4999 4559 5003
rect 4525 4994 4529 4998
rect 4535 4994 4539 4998
rect 4545 4994 4549 4998
rect 4555 4994 4559 4998
rect 4525 4989 4529 4993
rect 4535 4989 4539 4993
rect 4545 4989 4549 4993
rect 4555 4989 4559 4993
rect 4525 4811 4529 4815
rect 4535 4811 4539 4815
rect 4545 4811 4549 4815
rect 4555 4811 4559 4815
rect 4525 4806 4529 4810
rect 4535 4806 4539 4810
rect 4545 4806 4549 4810
rect 4555 4806 4559 4810
rect 4525 4801 4529 4805
rect 4535 4801 4539 4805
rect 4545 4801 4549 4805
rect 4555 4801 4559 4805
rect 4525 4796 4529 4800
rect 4535 4796 4539 4800
rect 4545 4796 4549 4800
rect 4555 4796 4559 4800
rect 4525 4785 4529 4789
rect 4535 4785 4539 4789
rect 4545 4785 4549 4789
rect 4555 4785 4559 4789
rect 4525 4780 4529 4784
rect 4535 4780 4539 4784
rect 4545 4780 4549 4784
rect 4555 4780 4559 4784
rect 4525 4775 4529 4779
rect 4535 4775 4539 4779
rect 4545 4775 4549 4779
rect 4555 4775 4559 4779
rect 4525 4770 4529 4774
rect 4535 4770 4539 4774
rect 4545 4770 4549 4774
rect 4555 4770 4559 4774
rect 4525 4759 4529 4763
rect 4535 4759 4539 4763
rect 4545 4759 4549 4763
rect 4555 4759 4559 4763
rect 4525 4754 4529 4758
rect 4535 4754 4539 4758
rect 4545 4754 4549 4758
rect 4555 4754 4559 4758
rect 4525 4749 4529 4753
rect 4535 4749 4539 4753
rect 4545 4749 4549 4753
rect 4555 4749 4559 4753
rect 4525 4744 4529 4748
rect 4535 4744 4539 4748
rect 4545 4744 4549 4748
rect 4555 4744 4559 4748
rect 4525 4733 4529 4737
rect 4535 4733 4539 4737
rect 4545 4733 4549 4737
rect 4555 4733 4559 4737
rect 4525 4728 4529 4732
rect 4535 4728 4539 4732
rect 4545 4728 4549 4732
rect 4555 4728 4559 4732
rect 4525 4723 4529 4727
rect 4535 4723 4539 4727
rect 4545 4723 4549 4727
rect 4555 4723 4559 4727
rect 4525 4718 4529 4722
rect 4535 4718 4539 4722
rect 4545 4718 4549 4722
rect 4555 4718 4559 4722
rect 4525 4707 4529 4711
rect 4535 4707 4539 4711
rect 4545 4707 4549 4711
rect 4555 4707 4559 4711
rect 4525 4702 4529 4706
rect 4535 4702 4539 4706
rect 4545 4702 4549 4706
rect 4555 4702 4559 4706
rect 4525 4697 4529 4701
rect 4535 4697 4539 4701
rect 4545 4697 4549 4701
rect 4555 4697 4559 4701
rect 4525 4692 4529 4696
rect 4535 4692 4539 4696
rect 4545 4692 4549 4696
rect 4555 4692 4559 4696
rect 757 4578 761 4582
rect 762 4578 766 4582
rect 767 4578 771 4582
rect 772 4578 776 4582
rect 783 4578 787 4582
rect 788 4578 792 4582
rect 793 4578 797 4582
rect 798 4578 802 4582
rect 809 4578 813 4582
rect 814 4578 818 4582
rect 819 4578 823 4582
rect 824 4578 828 4582
rect 835 4578 839 4582
rect 840 4578 844 4582
rect 845 4578 849 4582
rect 850 4578 854 4582
rect 861 4578 865 4582
rect 866 4578 870 4582
rect 871 4578 875 4582
rect 876 4578 880 4582
rect 1053 4578 1057 4582
rect 1058 4578 1062 4582
rect 1063 4578 1067 4582
rect 1068 4578 1072 4582
rect 1362 4578 1366 4582
rect 1367 4578 1371 4582
rect 1372 4578 1376 4582
rect 1377 4578 1381 4582
rect 1671 4578 1675 4582
rect 1676 4578 1680 4582
rect 1681 4578 1685 4582
rect 1686 4578 1690 4582
rect 1980 4578 1984 4582
rect 1985 4578 1989 4582
rect 1990 4578 1994 4582
rect 1995 4578 1999 4582
rect 2289 4578 2293 4582
rect 2294 4578 2298 4582
rect 2299 4578 2303 4582
rect 2304 4578 2308 4582
rect 2598 4578 2602 4582
rect 2603 4578 2607 4582
rect 2608 4578 2612 4582
rect 2613 4578 2617 4582
rect 2907 4578 2911 4582
rect 2912 4578 2916 4582
rect 2917 4578 2921 4582
rect 2922 4578 2926 4582
rect 3216 4578 3220 4582
rect 3221 4578 3225 4582
rect 3226 4578 3230 4582
rect 3231 4578 3235 4582
rect 3525 4578 3529 4582
rect 3530 4578 3534 4582
rect 3535 4578 3539 4582
rect 3540 4578 3544 4582
rect 3834 4578 3838 4582
rect 3839 4578 3843 4582
rect 3844 4578 3848 4582
rect 3849 4578 3853 4582
rect 4235 4578 4239 4582
rect 4240 4578 4244 4582
rect 4245 4578 4249 4582
rect 4250 4578 4254 4582
rect 4264 4578 4268 4582
rect 4269 4578 4273 4582
rect 4274 4578 4278 4582
rect 4279 4578 4283 4582
rect 4293 4578 4297 4582
rect 4298 4578 4302 4582
rect 4303 4578 4307 4582
rect 4308 4578 4312 4582
rect 4322 4578 4326 4582
rect 4327 4578 4331 4582
rect 4332 4578 4336 4582
rect 4337 4578 4341 4582
rect 4351 4578 4355 4582
rect 4356 4578 4360 4582
rect 4361 4578 4365 4582
rect 4366 4578 4370 4582
rect 757 4568 761 4572
rect 762 4568 766 4572
rect 767 4568 771 4572
rect 772 4568 776 4572
rect 783 4568 787 4572
rect 788 4568 792 4572
rect 793 4568 797 4572
rect 798 4568 802 4572
rect 809 4568 813 4572
rect 814 4568 818 4572
rect 819 4568 823 4572
rect 824 4568 828 4572
rect 835 4568 839 4572
rect 840 4568 844 4572
rect 845 4568 849 4572
rect 850 4568 854 4572
rect 861 4568 865 4572
rect 866 4568 870 4572
rect 871 4568 875 4572
rect 876 4568 880 4572
rect 1053 4568 1057 4572
rect 1058 4568 1062 4572
rect 1063 4568 1067 4572
rect 1068 4568 1072 4572
rect 1362 4568 1366 4572
rect 1367 4568 1371 4572
rect 1372 4568 1376 4572
rect 1377 4568 1381 4572
rect 1671 4568 1675 4572
rect 1676 4568 1680 4572
rect 1681 4568 1685 4572
rect 1686 4568 1690 4572
rect 1980 4568 1984 4572
rect 1985 4568 1989 4572
rect 1990 4568 1994 4572
rect 1995 4568 1999 4572
rect 2289 4568 2293 4572
rect 2294 4568 2298 4572
rect 2299 4568 2303 4572
rect 2304 4568 2308 4572
rect 2598 4568 2602 4572
rect 2603 4568 2607 4572
rect 2608 4568 2612 4572
rect 2613 4568 2617 4572
rect 2907 4568 2911 4572
rect 2912 4568 2916 4572
rect 2917 4568 2921 4572
rect 2922 4568 2926 4572
rect 3216 4568 3220 4572
rect 3221 4568 3225 4572
rect 3226 4568 3230 4572
rect 3231 4568 3235 4572
rect 3525 4568 3529 4572
rect 3530 4568 3534 4572
rect 3535 4568 3539 4572
rect 3540 4568 3544 4572
rect 3834 4568 3838 4572
rect 3839 4568 3843 4572
rect 3844 4568 3848 4572
rect 3849 4568 3853 4572
rect 4235 4568 4239 4572
rect 4240 4568 4244 4572
rect 4245 4568 4249 4572
rect 4250 4568 4254 4572
rect 4264 4568 4268 4572
rect 4269 4568 4273 4572
rect 4274 4568 4278 4572
rect 4279 4568 4283 4572
rect 4293 4568 4297 4572
rect 4298 4568 4302 4572
rect 4303 4568 4307 4572
rect 4308 4568 4312 4572
rect 4322 4568 4326 4572
rect 4327 4568 4331 4572
rect 4332 4568 4336 4572
rect 4337 4568 4341 4572
rect 4351 4568 4355 4572
rect 4356 4568 4360 4572
rect 4361 4568 4365 4572
rect 4366 4568 4370 4572
rect 757 4558 761 4562
rect 762 4558 766 4562
rect 767 4558 771 4562
rect 772 4558 776 4562
rect 783 4558 787 4562
rect 788 4558 792 4562
rect 793 4558 797 4562
rect 798 4558 802 4562
rect 809 4558 813 4562
rect 814 4558 818 4562
rect 819 4558 823 4562
rect 824 4558 828 4562
rect 835 4558 839 4562
rect 840 4558 844 4562
rect 845 4558 849 4562
rect 850 4558 854 4562
rect 861 4558 865 4562
rect 866 4558 870 4562
rect 871 4558 875 4562
rect 876 4558 880 4562
rect 1053 4558 1057 4562
rect 1058 4558 1062 4562
rect 1063 4558 1067 4562
rect 1068 4558 1072 4562
rect 1362 4558 1366 4562
rect 1367 4558 1371 4562
rect 1372 4558 1376 4562
rect 1377 4558 1381 4562
rect 1671 4558 1675 4562
rect 1676 4558 1680 4562
rect 1681 4558 1685 4562
rect 1686 4558 1690 4562
rect 1980 4558 1984 4562
rect 1985 4558 1989 4562
rect 1990 4558 1994 4562
rect 1995 4558 1999 4562
rect 2289 4558 2293 4562
rect 2294 4558 2298 4562
rect 2299 4558 2303 4562
rect 2304 4558 2308 4562
rect 2598 4558 2602 4562
rect 2603 4558 2607 4562
rect 2608 4558 2612 4562
rect 2613 4558 2617 4562
rect 2907 4558 2911 4562
rect 2912 4558 2916 4562
rect 2917 4558 2921 4562
rect 2922 4558 2926 4562
rect 3216 4558 3220 4562
rect 3221 4558 3225 4562
rect 3226 4558 3230 4562
rect 3231 4558 3235 4562
rect 3525 4558 3529 4562
rect 3530 4558 3534 4562
rect 3535 4558 3539 4562
rect 3540 4558 3544 4562
rect 3834 4558 3838 4562
rect 3839 4558 3843 4562
rect 3844 4558 3848 4562
rect 3849 4558 3853 4562
rect 4235 4558 4239 4562
rect 4240 4558 4244 4562
rect 4245 4558 4249 4562
rect 4250 4558 4254 4562
rect 4264 4558 4268 4562
rect 4269 4558 4273 4562
rect 4274 4558 4278 4562
rect 4279 4558 4283 4562
rect 4293 4558 4297 4562
rect 4298 4558 4302 4562
rect 4303 4558 4307 4562
rect 4308 4558 4312 4562
rect 4322 4558 4326 4562
rect 4327 4558 4331 4562
rect 4332 4558 4336 4562
rect 4337 4558 4341 4562
rect 4351 4558 4355 4562
rect 4356 4558 4360 4562
rect 4361 4558 4365 4562
rect 4366 4558 4370 4562
rect 757 4548 761 4552
rect 762 4548 766 4552
rect 767 4548 771 4552
rect 772 4548 776 4552
rect 783 4548 787 4552
rect 788 4548 792 4552
rect 793 4548 797 4552
rect 798 4548 802 4552
rect 809 4548 813 4552
rect 814 4548 818 4552
rect 819 4548 823 4552
rect 824 4548 828 4552
rect 835 4548 839 4552
rect 840 4548 844 4552
rect 845 4548 849 4552
rect 850 4548 854 4552
rect 861 4548 865 4552
rect 866 4548 870 4552
rect 871 4548 875 4552
rect 876 4548 880 4552
rect 1053 4548 1057 4552
rect 1058 4548 1062 4552
rect 1063 4548 1067 4552
rect 1068 4548 1072 4552
rect 1362 4548 1366 4552
rect 1367 4548 1371 4552
rect 1372 4548 1376 4552
rect 1377 4548 1381 4552
rect 1671 4548 1675 4552
rect 1676 4548 1680 4552
rect 1681 4548 1685 4552
rect 1686 4548 1690 4552
rect 1980 4548 1984 4552
rect 1985 4548 1989 4552
rect 1990 4548 1994 4552
rect 1995 4548 1999 4552
rect 2289 4548 2293 4552
rect 2294 4548 2298 4552
rect 2299 4548 2303 4552
rect 2304 4548 2308 4552
rect 2598 4548 2602 4552
rect 2603 4548 2607 4552
rect 2608 4548 2612 4552
rect 2613 4548 2617 4552
rect 2907 4548 2911 4552
rect 2912 4548 2916 4552
rect 2917 4548 2921 4552
rect 2922 4548 2926 4552
rect 3216 4548 3220 4552
rect 3221 4548 3225 4552
rect 3226 4548 3230 4552
rect 3231 4548 3235 4552
rect 3525 4548 3529 4552
rect 3530 4548 3534 4552
rect 3535 4548 3539 4552
rect 3540 4548 3544 4552
rect 3834 4548 3838 4552
rect 3839 4548 3843 4552
rect 3844 4548 3848 4552
rect 3849 4548 3853 4552
rect 4235 4548 4239 4552
rect 4240 4548 4244 4552
rect 4245 4548 4249 4552
rect 4250 4548 4254 4552
rect 4264 4548 4268 4552
rect 4269 4548 4273 4552
rect 4274 4548 4278 4552
rect 4279 4548 4283 4552
rect 4293 4548 4297 4552
rect 4298 4548 4302 4552
rect 4303 4548 4307 4552
rect 4308 4548 4312 4552
rect 4322 4548 4326 4552
rect 4327 4548 4331 4552
rect 4332 4548 4336 4552
rect 4337 4548 4341 4552
rect 4351 4548 4355 4552
rect 4356 4548 4360 4552
rect 4361 4548 4365 4552
rect 4366 4548 4370 4552
rect 1087 4458 1091 4462
rect 1094 4458 1098 4462
rect 1099 4458 1103 4462
rect 1104 4458 1108 4462
rect 1109 4458 1113 4462
rect 1114 4458 1118 4462
rect 1119 4458 1123 4462
rect 1124 4458 1128 4462
rect 1129 4458 1133 4462
rect 1134 4458 1138 4462
rect 1139 4458 1143 4462
rect 1144 4458 1148 4462
rect 1151 4458 1155 4462
rect 1087 4451 1091 4455
rect 1151 4451 1155 4455
rect 1087 4446 1091 4450
rect 1087 4441 1091 4445
rect 1087 4436 1091 4440
rect 1087 4431 1091 4435
rect 1087 4426 1091 4430
rect 1087 4421 1091 4425
rect 1087 4416 1091 4420
rect 1087 4411 1091 4415
rect 1087 4406 1091 4410
rect 1087 4401 1091 4405
rect 1087 4396 1091 4400
rect 1087 4391 1091 4395
rect 1087 4386 1091 4390
rect 1087 4381 1091 4385
rect 1087 4376 1091 4380
rect 1087 4371 1091 4375
rect 1087 4366 1091 4370
rect 1087 4361 1091 4365
rect 1151 4446 1155 4450
rect 1151 4441 1155 4445
rect 1151 4436 1155 4440
rect 1151 4431 1155 4435
rect 1151 4426 1155 4430
rect 1151 4421 1155 4425
rect 1151 4416 1155 4420
rect 1151 4411 1155 4415
rect 1151 4406 1155 4410
rect 1151 4401 1155 4405
rect 1151 4396 1155 4400
rect 1151 4391 1155 4395
rect 1151 4386 1155 4390
rect 1151 4381 1155 4385
rect 1151 4376 1155 4380
rect 1151 4371 1155 4375
rect 1151 4366 1155 4370
rect 1151 4361 1155 4365
rect 1087 4356 1091 4360
rect 1151 4356 1155 4360
rect 1087 4349 1091 4353
rect 1094 4349 1098 4353
rect 1099 4349 1103 4353
rect 1104 4349 1108 4353
rect 1109 4349 1113 4353
rect 1114 4349 1118 4353
rect 1119 4349 1123 4353
rect 1124 4349 1128 4353
rect 1129 4349 1133 4353
rect 1134 4349 1138 4353
rect 1139 4349 1143 4353
rect 1144 4349 1148 4353
rect 1151 4349 1155 4353
rect 1234 4471 1238 4475
rect 1239 4471 1243 4475
rect 1244 4471 1248 4475
rect 1249 4471 1253 4475
rect 1254 4471 1258 4475
rect 1259 4471 1263 4475
rect 1264 4471 1268 4475
rect 1269 4471 1273 4475
rect 1274 4471 1278 4475
rect 1279 4471 1283 4475
rect 1284 4471 1288 4475
rect 1289 4471 1293 4475
rect 1294 4471 1298 4475
rect 1299 4471 1303 4475
rect 1304 4471 1308 4475
rect 1309 4471 1313 4475
rect 1314 4471 1318 4475
rect 1319 4471 1323 4475
rect 1324 4471 1328 4475
rect 1234 4466 1238 4470
rect 1234 4461 1238 4465
rect 1324 4466 1328 4470
rect 1234 4456 1238 4460
rect 1234 4451 1238 4455
rect 1234 4446 1238 4450
rect 1234 4441 1238 4445
rect 1234 4436 1238 4440
rect 1234 4431 1238 4435
rect 1234 4426 1238 4430
rect 1234 4421 1238 4425
rect 1234 4416 1238 4420
rect 1234 4411 1238 4415
rect 1234 4406 1238 4410
rect 1234 4401 1238 4405
rect 1234 4396 1238 4400
rect 1234 4391 1238 4395
rect 1234 4386 1238 4390
rect 1234 4381 1238 4385
rect 1234 4376 1238 4380
rect 1234 4371 1238 4375
rect 1234 4366 1238 4370
rect 1234 4361 1238 4365
rect 1234 4356 1238 4360
rect 1234 4351 1238 4355
rect 1234 4346 1238 4350
rect 1324 4461 1328 4465
rect 1324 4456 1328 4460
rect 1324 4451 1328 4455
rect 1324 4446 1328 4450
rect 1324 4441 1328 4445
rect 1324 4436 1328 4440
rect 1324 4431 1328 4435
rect 1324 4426 1328 4430
rect 1324 4421 1328 4425
rect 1324 4416 1328 4420
rect 1324 4411 1328 4415
rect 1324 4406 1328 4410
rect 1324 4401 1328 4405
rect 1324 4396 1328 4400
rect 1324 4391 1328 4395
rect 1324 4386 1328 4390
rect 1324 4381 1328 4385
rect 1324 4376 1328 4380
rect 1324 4371 1328 4375
rect 1324 4366 1328 4370
rect 1324 4361 1328 4365
rect 1324 4356 1328 4360
rect 1324 4351 1328 4355
rect 1234 4341 1238 4345
rect 1324 4346 1328 4350
rect 1324 4341 1328 4345
rect 1234 4336 1238 4340
rect 1239 4336 1243 4340
rect 1244 4336 1248 4340
rect 1249 4336 1253 4340
rect 1254 4336 1258 4340
rect 1259 4336 1263 4340
rect 1264 4336 1268 4340
rect 1269 4336 1273 4340
rect 1274 4336 1278 4340
rect 1279 4336 1283 4340
rect 1284 4336 1288 4340
rect 1289 4336 1293 4340
rect 1294 4336 1298 4340
rect 1299 4336 1303 4340
rect 1304 4336 1308 4340
rect 1309 4336 1313 4340
rect 1314 4336 1318 4340
rect 1319 4336 1323 4340
rect 1324 4336 1328 4340
rect 1396 4458 1400 4462
rect 1403 4458 1407 4462
rect 1408 4458 1412 4462
rect 1413 4458 1417 4462
rect 1418 4458 1422 4462
rect 1423 4458 1427 4462
rect 1428 4458 1432 4462
rect 1433 4458 1437 4462
rect 1438 4458 1442 4462
rect 1443 4458 1447 4462
rect 1448 4458 1452 4462
rect 1453 4458 1457 4462
rect 1460 4458 1464 4462
rect 1396 4451 1400 4455
rect 1460 4451 1464 4455
rect 1396 4446 1400 4450
rect 1396 4441 1400 4445
rect 1396 4436 1400 4440
rect 1396 4431 1400 4435
rect 1396 4426 1400 4430
rect 1396 4421 1400 4425
rect 1396 4416 1400 4420
rect 1396 4411 1400 4415
rect 1396 4406 1400 4410
rect 1396 4401 1400 4405
rect 1396 4396 1400 4400
rect 1396 4391 1400 4395
rect 1396 4386 1400 4390
rect 1396 4381 1400 4385
rect 1396 4376 1400 4380
rect 1396 4371 1400 4375
rect 1396 4366 1400 4370
rect 1396 4361 1400 4365
rect 1460 4446 1464 4450
rect 1460 4441 1464 4445
rect 1460 4436 1464 4440
rect 1460 4431 1464 4435
rect 1460 4426 1464 4430
rect 1460 4421 1464 4425
rect 1460 4416 1464 4420
rect 1460 4411 1464 4415
rect 1460 4406 1464 4410
rect 1460 4401 1464 4405
rect 1460 4396 1464 4400
rect 1460 4391 1464 4395
rect 1460 4386 1464 4390
rect 1460 4381 1464 4385
rect 1460 4376 1464 4380
rect 1460 4371 1464 4375
rect 1460 4366 1464 4370
rect 1460 4361 1464 4365
rect 1396 4356 1400 4360
rect 1460 4356 1464 4360
rect 1396 4349 1400 4353
rect 1403 4349 1407 4353
rect 1408 4349 1412 4353
rect 1413 4349 1417 4353
rect 1418 4349 1422 4353
rect 1423 4349 1427 4353
rect 1428 4349 1432 4353
rect 1433 4349 1437 4353
rect 1438 4349 1442 4353
rect 1443 4349 1447 4353
rect 1448 4349 1452 4353
rect 1453 4349 1457 4353
rect 1460 4349 1464 4353
rect 1543 4471 1547 4475
rect 1548 4471 1552 4475
rect 1553 4471 1557 4475
rect 1558 4471 1562 4475
rect 1563 4471 1567 4475
rect 1568 4471 1572 4475
rect 1573 4471 1577 4475
rect 1578 4471 1582 4475
rect 1583 4471 1587 4475
rect 1588 4471 1592 4475
rect 1593 4471 1597 4475
rect 1598 4471 1602 4475
rect 1603 4471 1607 4475
rect 1608 4471 1612 4475
rect 1613 4471 1617 4475
rect 1618 4471 1622 4475
rect 1623 4471 1627 4475
rect 1628 4471 1632 4475
rect 1633 4471 1637 4475
rect 1543 4466 1547 4470
rect 1543 4461 1547 4465
rect 1633 4466 1637 4470
rect 1543 4456 1547 4460
rect 1543 4451 1547 4455
rect 1543 4446 1547 4450
rect 1543 4441 1547 4445
rect 1543 4436 1547 4440
rect 1543 4431 1547 4435
rect 1543 4426 1547 4430
rect 1543 4421 1547 4425
rect 1543 4416 1547 4420
rect 1543 4411 1547 4415
rect 1543 4406 1547 4410
rect 1543 4401 1547 4405
rect 1543 4396 1547 4400
rect 1543 4391 1547 4395
rect 1543 4386 1547 4390
rect 1543 4381 1547 4385
rect 1543 4376 1547 4380
rect 1543 4371 1547 4375
rect 1543 4366 1547 4370
rect 1543 4361 1547 4365
rect 1543 4356 1547 4360
rect 1543 4351 1547 4355
rect 1543 4346 1547 4350
rect 1633 4461 1637 4465
rect 1633 4456 1637 4460
rect 1633 4451 1637 4455
rect 1633 4446 1637 4450
rect 1633 4441 1637 4445
rect 1633 4436 1637 4440
rect 1633 4431 1637 4435
rect 1633 4426 1637 4430
rect 1633 4421 1637 4425
rect 1633 4416 1637 4420
rect 1633 4411 1637 4415
rect 1633 4406 1637 4410
rect 1633 4401 1637 4405
rect 1633 4396 1637 4400
rect 1633 4391 1637 4395
rect 1633 4386 1637 4390
rect 1633 4381 1637 4385
rect 1633 4376 1637 4380
rect 1633 4371 1637 4375
rect 1633 4366 1637 4370
rect 1633 4361 1637 4365
rect 1633 4356 1637 4360
rect 1633 4351 1637 4355
rect 1543 4341 1547 4345
rect 1633 4346 1637 4350
rect 1633 4341 1637 4345
rect 1543 4336 1547 4340
rect 1548 4336 1552 4340
rect 1553 4336 1557 4340
rect 1558 4336 1562 4340
rect 1563 4336 1567 4340
rect 1568 4336 1572 4340
rect 1573 4336 1577 4340
rect 1578 4336 1582 4340
rect 1583 4336 1587 4340
rect 1588 4336 1592 4340
rect 1593 4336 1597 4340
rect 1598 4336 1602 4340
rect 1603 4336 1607 4340
rect 1608 4336 1612 4340
rect 1613 4336 1617 4340
rect 1618 4336 1622 4340
rect 1623 4336 1627 4340
rect 1628 4336 1632 4340
rect 1633 4336 1637 4340
rect 1705 4458 1709 4462
rect 1712 4458 1716 4462
rect 1717 4458 1721 4462
rect 1722 4458 1726 4462
rect 1727 4458 1731 4462
rect 1732 4458 1736 4462
rect 1737 4458 1741 4462
rect 1742 4458 1746 4462
rect 1747 4458 1751 4462
rect 1752 4458 1756 4462
rect 1757 4458 1761 4462
rect 1762 4458 1766 4462
rect 1769 4458 1773 4462
rect 1705 4451 1709 4455
rect 1769 4451 1773 4455
rect 1705 4446 1709 4450
rect 1705 4441 1709 4445
rect 1705 4436 1709 4440
rect 1705 4431 1709 4435
rect 1705 4426 1709 4430
rect 1705 4421 1709 4425
rect 1705 4416 1709 4420
rect 1705 4411 1709 4415
rect 1705 4406 1709 4410
rect 1705 4401 1709 4405
rect 1705 4396 1709 4400
rect 1705 4391 1709 4395
rect 1705 4386 1709 4390
rect 1705 4381 1709 4385
rect 1705 4376 1709 4380
rect 1705 4371 1709 4375
rect 1705 4366 1709 4370
rect 1705 4361 1709 4365
rect 1769 4446 1773 4450
rect 1769 4441 1773 4445
rect 1769 4436 1773 4440
rect 1769 4431 1773 4435
rect 1769 4426 1773 4430
rect 1769 4421 1773 4425
rect 1769 4416 1773 4420
rect 1769 4411 1773 4415
rect 1769 4406 1773 4410
rect 1769 4401 1773 4405
rect 1769 4396 1773 4400
rect 1769 4391 1773 4395
rect 1769 4386 1773 4390
rect 1769 4381 1773 4385
rect 1769 4376 1773 4380
rect 1769 4371 1773 4375
rect 1769 4366 1773 4370
rect 1769 4361 1773 4365
rect 1705 4356 1709 4360
rect 1769 4356 1773 4360
rect 1705 4349 1709 4353
rect 1712 4349 1716 4353
rect 1717 4349 1721 4353
rect 1722 4349 1726 4353
rect 1727 4349 1731 4353
rect 1732 4349 1736 4353
rect 1737 4349 1741 4353
rect 1742 4349 1746 4353
rect 1747 4349 1751 4353
rect 1752 4349 1756 4353
rect 1757 4349 1761 4353
rect 1762 4349 1766 4353
rect 1769 4349 1773 4353
rect 1852 4471 1856 4475
rect 1857 4471 1861 4475
rect 1862 4471 1866 4475
rect 1867 4471 1871 4475
rect 1872 4471 1876 4475
rect 1877 4471 1881 4475
rect 1882 4471 1886 4475
rect 1887 4471 1891 4475
rect 1892 4471 1896 4475
rect 1897 4471 1901 4475
rect 1902 4471 1906 4475
rect 1907 4471 1911 4475
rect 1912 4471 1916 4475
rect 1917 4471 1921 4475
rect 1922 4471 1926 4475
rect 1927 4471 1931 4475
rect 1932 4471 1936 4475
rect 1937 4471 1941 4475
rect 1942 4471 1946 4475
rect 1852 4466 1856 4470
rect 1852 4461 1856 4465
rect 1942 4466 1946 4470
rect 1852 4456 1856 4460
rect 1852 4451 1856 4455
rect 1852 4446 1856 4450
rect 1852 4441 1856 4445
rect 1852 4436 1856 4440
rect 1852 4431 1856 4435
rect 1852 4426 1856 4430
rect 1852 4421 1856 4425
rect 1852 4416 1856 4420
rect 1852 4411 1856 4415
rect 1852 4406 1856 4410
rect 1852 4401 1856 4405
rect 1852 4396 1856 4400
rect 1852 4391 1856 4395
rect 1852 4386 1856 4390
rect 1852 4381 1856 4385
rect 1852 4376 1856 4380
rect 1852 4371 1856 4375
rect 1852 4366 1856 4370
rect 1852 4361 1856 4365
rect 1852 4356 1856 4360
rect 1852 4351 1856 4355
rect 1852 4346 1856 4350
rect 1942 4461 1946 4465
rect 1942 4456 1946 4460
rect 1942 4451 1946 4455
rect 1942 4446 1946 4450
rect 1942 4441 1946 4445
rect 1942 4436 1946 4440
rect 1942 4431 1946 4435
rect 1942 4426 1946 4430
rect 1942 4421 1946 4425
rect 1942 4416 1946 4420
rect 1942 4411 1946 4415
rect 1942 4406 1946 4410
rect 1942 4401 1946 4405
rect 1942 4396 1946 4400
rect 1942 4391 1946 4395
rect 1942 4386 1946 4390
rect 1942 4381 1946 4385
rect 1942 4376 1946 4380
rect 1942 4371 1946 4375
rect 1942 4366 1946 4370
rect 1942 4361 1946 4365
rect 1942 4356 1946 4360
rect 1942 4351 1946 4355
rect 1852 4341 1856 4345
rect 1942 4346 1946 4350
rect 1942 4341 1946 4345
rect 1852 4336 1856 4340
rect 1857 4336 1861 4340
rect 1862 4336 1866 4340
rect 1867 4336 1871 4340
rect 1872 4336 1876 4340
rect 1877 4336 1881 4340
rect 1882 4336 1886 4340
rect 1887 4336 1891 4340
rect 1892 4336 1896 4340
rect 1897 4336 1901 4340
rect 1902 4336 1906 4340
rect 1907 4336 1911 4340
rect 1912 4336 1916 4340
rect 1917 4336 1921 4340
rect 1922 4336 1926 4340
rect 1927 4336 1931 4340
rect 1932 4336 1936 4340
rect 1937 4336 1941 4340
rect 1942 4336 1946 4340
rect 2014 4458 2018 4462
rect 2021 4458 2025 4462
rect 2026 4458 2030 4462
rect 2031 4458 2035 4462
rect 2036 4458 2040 4462
rect 2041 4458 2045 4462
rect 2046 4458 2050 4462
rect 2051 4458 2055 4462
rect 2056 4458 2060 4462
rect 2061 4458 2065 4462
rect 2066 4458 2070 4462
rect 2071 4458 2075 4462
rect 2078 4458 2082 4462
rect 2014 4451 2018 4455
rect 2078 4451 2082 4455
rect 2014 4446 2018 4450
rect 2014 4441 2018 4445
rect 2014 4436 2018 4440
rect 2014 4431 2018 4435
rect 2014 4426 2018 4430
rect 2014 4421 2018 4425
rect 2014 4416 2018 4420
rect 2014 4411 2018 4415
rect 2014 4406 2018 4410
rect 2014 4401 2018 4405
rect 2014 4396 2018 4400
rect 2014 4391 2018 4395
rect 2014 4386 2018 4390
rect 2014 4381 2018 4385
rect 2014 4376 2018 4380
rect 2014 4371 2018 4375
rect 2014 4366 2018 4370
rect 2014 4361 2018 4365
rect 2078 4446 2082 4450
rect 2078 4441 2082 4445
rect 2078 4436 2082 4440
rect 2078 4431 2082 4435
rect 2078 4426 2082 4430
rect 2078 4421 2082 4425
rect 2078 4416 2082 4420
rect 2078 4411 2082 4415
rect 2078 4406 2082 4410
rect 2078 4401 2082 4405
rect 2078 4396 2082 4400
rect 2078 4391 2082 4395
rect 2078 4386 2082 4390
rect 2078 4381 2082 4385
rect 2078 4376 2082 4380
rect 2078 4371 2082 4375
rect 2078 4366 2082 4370
rect 2078 4361 2082 4365
rect 2014 4356 2018 4360
rect 2078 4356 2082 4360
rect 2014 4349 2018 4353
rect 2021 4349 2025 4353
rect 2026 4349 2030 4353
rect 2031 4349 2035 4353
rect 2036 4349 2040 4353
rect 2041 4349 2045 4353
rect 2046 4349 2050 4353
rect 2051 4349 2055 4353
rect 2056 4349 2060 4353
rect 2061 4349 2065 4353
rect 2066 4349 2070 4353
rect 2071 4349 2075 4353
rect 2078 4349 2082 4353
rect 2161 4471 2165 4475
rect 2166 4471 2170 4475
rect 2171 4471 2175 4475
rect 2176 4471 2180 4475
rect 2181 4471 2185 4475
rect 2186 4471 2190 4475
rect 2191 4471 2195 4475
rect 2196 4471 2200 4475
rect 2201 4471 2205 4475
rect 2206 4471 2210 4475
rect 2211 4471 2215 4475
rect 2216 4471 2220 4475
rect 2221 4471 2225 4475
rect 2226 4471 2230 4475
rect 2231 4471 2235 4475
rect 2236 4471 2240 4475
rect 2241 4471 2245 4475
rect 2246 4471 2250 4475
rect 2251 4471 2255 4475
rect 2161 4466 2165 4470
rect 2161 4461 2165 4465
rect 2251 4466 2255 4470
rect 2161 4456 2165 4460
rect 2161 4451 2165 4455
rect 2161 4446 2165 4450
rect 2161 4441 2165 4445
rect 2161 4436 2165 4440
rect 2161 4431 2165 4435
rect 2161 4426 2165 4430
rect 2161 4421 2165 4425
rect 2161 4416 2165 4420
rect 2161 4411 2165 4415
rect 2161 4406 2165 4410
rect 2161 4401 2165 4405
rect 2161 4396 2165 4400
rect 2161 4391 2165 4395
rect 2161 4386 2165 4390
rect 2161 4381 2165 4385
rect 2161 4376 2165 4380
rect 2161 4371 2165 4375
rect 2161 4366 2165 4370
rect 2161 4361 2165 4365
rect 2161 4356 2165 4360
rect 2161 4351 2165 4355
rect 2161 4346 2165 4350
rect 2251 4461 2255 4465
rect 2251 4456 2255 4460
rect 2251 4451 2255 4455
rect 2251 4446 2255 4450
rect 2251 4441 2255 4445
rect 2251 4436 2255 4440
rect 2251 4431 2255 4435
rect 2251 4426 2255 4430
rect 2251 4421 2255 4425
rect 2251 4416 2255 4420
rect 2251 4411 2255 4415
rect 2251 4406 2255 4410
rect 2251 4401 2255 4405
rect 2251 4396 2255 4400
rect 2251 4391 2255 4395
rect 2251 4386 2255 4390
rect 2251 4381 2255 4385
rect 2251 4376 2255 4380
rect 2251 4371 2255 4375
rect 2251 4366 2255 4370
rect 2251 4361 2255 4365
rect 2251 4356 2255 4360
rect 2251 4351 2255 4355
rect 2161 4341 2165 4345
rect 2251 4346 2255 4350
rect 2251 4341 2255 4345
rect 2161 4336 2165 4340
rect 2166 4336 2170 4340
rect 2171 4336 2175 4340
rect 2176 4336 2180 4340
rect 2181 4336 2185 4340
rect 2186 4336 2190 4340
rect 2191 4336 2195 4340
rect 2196 4336 2200 4340
rect 2201 4336 2205 4340
rect 2206 4336 2210 4340
rect 2211 4336 2215 4340
rect 2216 4336 2220 4340
rect 2221 4336 2225 4340
rect 2226 4336 2230 4340
rect 2231 4336 2235 4340
rect 2236 4336 2240 4340
rect 2241 4336 2245 4340
rect 2246 4336 2250 4340
rect 2251 4336 2255 4340
rect 2323 4458 2327 4462
rect 2330 4458 2334 4462
rect 2335 4458 2339 4462
rect 2340 4458 2344 4462
rect 2345 4458 2349 4462
rect 2350 4458 2354 4462
rect 2355 4458 2359 4462
rect 2360 4458 2364 4462
rect 2365 4458 2369 4462
rect 2370 4458 2374 4462
rect 2375 4458 2379 4462
rect 2380 4458 2384 4462
rect 2387 4458 2391 4462
rect 2323 4451 2327 4455
rect 2387 4451 2391 4455
rect 2323 4446 2327 4450
rect 2323 4441 2327 4445
rect 2323 4436 2327 4440
rect 2323 4431 2327 4435
rect 2323 4426 2327 4430
rect 2323 4421 2327 4425
rect 2323 4416 2327 4420
rect 2323 4411 2327 4415
rect 2323 4406 2327 4410
rect 2323 4401 2327 4405
rect 2323 4396 2327 4400
rect 2323 4391 2327 4395
rect 2323 4386 2327 4390
rect 2323 4381 2327 4385
rect 2323 4376 2327 4380
rect 2323 4371 2327 4375
rect 2323 4366 2327 4370
rect 2323 4361 2327 4365
rect 2387 4446 2391 4450
rect 2387 4441 2391 4445
rect 2387 4436 2391 4440
rect 2387 4431 2391 4435
rect 2387 4426 2391 4430
rect 2387 4421 2391 4425
rect 2387 4416 2391 4420
rect 2387 4411 2391 4415
rect 2387 4406 2391 4410
rect 2387 4401 2391 4405
rect 2387 4396 2391 4400
rect 2387 4391 2391 4395
rect 2387 4386 2391 4390
rect 2387 4381 2391 4385
rect 2387 4376 2391 4380
rect 2387 4371 2391 4375
rect 2387 4366 2391 4370
rect 2387 4361 2391 4365
rect 2323 4356 2327 4360
rect 2387 4356 2391 4360
rect 2323 4349 2327 4353
rect 2330 4349 2334 4353
rect 2335 4349 2339 4353
rect 2340 4349 2344 4353
rect 2345 4349 2349 4353
rect 2350 4349 2354 4353
rect 2355 4349 2359 4353
rect 2360 4349 2364 4353
rect 2365 4349 2369 4353
rect 2370 4349 2374 4353
rect 2375 4349 2379 4353
rect 2380 4349 2384 4353
rect 2387 4349 2391 4353
rect 2470 4471 2474 4475
rect 2475 4471 2479 4475
rect 2480 4471 2484 4475
rect 2485 4471 2489 4475
rect 2490 4471 2494 4475
rect 2495 4471 2499 4475
rect 2500 4471 2504 4475
rect 2505 4471 2509 4475
rect 2510 4471 2514 4475
rect 2515 4471 2519 4475
rect 2520 4471 2524 4475
rect 2525 4471 2529 4475
rect 2530 4471 2534 4475
rect 2535 4471 2539 4475
rect 2540 4471 2544 4475
rect 2545 4471 2549 4475
rect 2550 4471 2554 4475
rect 2555 4471 2559 4475
rect 2560 4471 2564 4475
rect 2470 4466 2474 4470
rect 2470 4461 2474 4465
rect 2560 4466 2564 4470
rect 2470 4456 2474 4460
rect 2470 4451 2474 4455
rect 2470 4446 2474 4450
rect 2470 4441 2474 4445
rect 2470 4436 2474 4440
rect 2470 4431 2474 4435
rect 2470 4426 2474 4430
rect 2470 4421 2474 4425
rect 2470 4416 2474 4420
rect 2470 4411 2474 4415
rect 2470 4406 2474 4410
rect 2470 4401 2474 4405
rect 2470 4396 2474 4400
rect 2470 4391 2474 4395
rect 2470 4386 2474 4390
rect 2470 4381 2474 4385
rect 2470 4376 2474 4380
rect 2470 4371 2474 4375
rect 2470 4366 2474 4370
rect 2470 4361 2474 4365
rect 2470 4356 2474 4360
rect 2470 4351 2474 4355
rect 2470 4346 2474 4350
rect 2560 4461 2564 4465
rect 2560 4456 2564 4460
rect 2560 4451 2564 4455
rect 2560 4446 2564 4450
rect 2560 4441 2564 4445
rect 2560 4436 2564 4440
rect 2560 4431 2564 4435
rect 2560 4426 2564 4430
rect 2560 4421 2564 4425
rect 2560 4416 2564 4420
rect 2560 4411 2564 4415
rect 2560 4406 2564 4410
rect 2560 4401 2564 4405
rect 2560 4396 2564 4400
rect 2560 4391 2564 4395
rect 2560 4386 2564 4390
rect 2560 4381 2564 4385
rect 2560 4376 2564 4380
rect 2560 4371 2564 4375
rect 2560 4366 2564 4370
rect 2560 4361 2564 4365
rect 2560 4356 2564 4360
rect 2560 4351 2564 4355
rect 2470 4341 2474 4345
rect 2560 4346 2564 4350
rect 2560 4341 2564 4345
rect 2470 4336 2474 4340
rect 2475 4336 2479 4340
rect 2480 4336 2484 4340
rect 2485 4336 2489 4340
rect 2490 4336 2494 4340
rect 2495 4336 2499 4340
rect 2500 4336 2504 4340
rect 2505 4336 2509 4340
rect 2510 4336 2514 4340
rect 2515 4336 2519 4340
rect 2520 4336 2524 4340
rect 2525 4336 2529 4340
rect 2530 4336 2534 4340
rect 2535 4336 2539 4340
rect 2540 4336 2544 4340
rect 2545 4336 2549 4340
rect 2550 4336 2554 4340
rect 2555 4336 2559 4340
rect 2560 4336 2564 4340
rect 2632 4458 2636 4462
rect 2639 4458 2643 4462
rect 2644 4458 2648 4462
rect 2649 4458 2653 4462
rect 2654 4458 2658 4462
rect 2659 4458 2663 4462
rect 2664 4458 2668 4462
rect 2669 4458 2673 4462
rect 2674 4458 2678 4462
rect 2679 4458 2683 4462
rect 2684 4458 2688 4462
rect 2689 4458 2693 4462
rect 2696 4458 2700 4462
rect 2632 4451 2636 4455
rect 2696 4451 2700 4455
rect 2632 4446 2636 4450
rect 2632 4441 2636 4445
rect 2632 4436 2636 4440
rect 2632 4431 2636 4435
rect 2632 4426 2636 4430
rect 2632 4421 2636 4425
rect 2632 4416 2636 4420
rect 2632 4411 2636 4415
rect 2632 4406 2636 4410
rect 2632 4401 2636 4405
rect 2632 4396 2636 4400
rect 2632 4391 2636 4395
rect 2632 4386 2636 4390
rect 2632 4381 2636 4385
rect 2632 4376 2636 4380
rect 2632 4371 2636 4375
rect 2632 4366 2636 4370
rect 2632 4361 2636 4365
rect 2696 4446 2700 4450
rect 2696 4441 2700 4445
rect 2696 4436 2700 4440
rect 2696 4431 2700 4435
rect 2696 4426 2700 4430
rect 2696 4421 2700 4425
rect 2696 4416 2700 4420
rect 2696 4411 2700 4415
rect 2696 4406 2700 4410
rect 2696 4401 2700 4405
rect 2696 4396 2700 4400
rect 2696 4391 2700 4395
rect 2696 4386 2700 4390
rect 2696 4381 2700 4385
rect 2696 4376 2700 4380
rect 2696 4371 2700 4375
rect 2696 4366 2700 4370
rect 2696 4361 2700 4365
rect 2632 4356 2636 4360
rect 2696 4356 2700 4360
rect 2632 4349 2636 4353
rect 2639 4349 2643 4353
rect 2644 4349 2648 4353
rect 2649 4349 2653 4353
rect 2654 4349 2658 4353
rect 2659 4349 2663 4353
rect 2664 4349 2668 4353
rect 2669 4349 2673 4353
rect 2674 4349 2678 4353
rect 2679 4349 2683 4353
rect 2684 4349 2688 4353
rect 2689 4349 2693 4353
rect 2696 4349 2700 4353
rect 2779 4471 2783 4475
rect 2784 4471 2788 4475
rect 2789 4471 2793 4475
rect 2794 4471 2798 4475
rect 2799 4471 2803 4475
rect 2804 4471 2808 4475
rect 2809 4471 2813 4475
rect 2814 4471 2818 4475
rect 2819 4471 2823 4475
rect 2824 4471 2828 4475
rect 2829 4471 2833 4475
rect 2834 4471 2838 4475
rect 2839 4471 2843 4475
rect 2844 4471 2848 4475
rect 2849 4471 2853 4475
rect 2854 4471 2858 4475
rect 2859 4471 2863 4475
rect 2864 4471 2868 4475
rect 2869 4471 2873 4475
rect 2779 4466 2783 4470
rect 2779 4461 2783 4465
rect 2869 4466 2873 4470
rect 2779 4456 2783 4460
rect 2779 4451 2783 4455
rect 2779 4446 2783 4450
rect 2779 4441 2783 4445
rect 2779 4436 2783 4440
rect 2779 4431 2783 4435
rect 2779 4426 2783 4430
rect 2779 4421 2783 4425
rect 2779 4416 2783 4420
rect 2779 4411 2783 4415
rect 2779 4406 2783 4410
rect 2779 4401 2783 4405
rect 2779 4396 2783 4400
rect 2779 4391 2783 4395
rect 2779 4386 2783 4390
rect 2779 4381 2783 4385
rect 2779 4376 2783 4380
rect 2779 4371 2783 4375
rect 2779 4366 2783 4370
rect 2779 4361 2783 4365
rect 2779 4356 2783 4360
rect 2779 4351 2783 4355
rect 2779 4346 2783 4350
rect 2869 4461 2873 4465
rect 2869 4456 2873 4460
rect 2869 4451 2873 4455
rect 2869 4446 2873 4450
rect 2869 4441 2873 4445
rect 2869 4436 2873 4440
rect 2869 4431 2873 4435
rect 2869 4426 2873 4430
rect 2869 4421 2873 4425
rect 2869 4416 2873 4420
rect 2869 4411 2873 4415
rect 2869 4406 2873 4410
rect 2869 4401 2873 4405
rect 2869 4396 2873 4400
rect 2869 4391 2873 4395
rect 2869 4386 2873 4390
rect 2869 4381 2873 4385
rect 2869 4376 2873 4380
rect 2869 4371 2873 4375
rect 2869 4366 2873 4370
rect 2869 4361 2873 4365
rect 2869 4356 2873 4360
rect 2869 4351 2873 4355
rect 2779 4341 2783 4345
rect 2869 4346 2873 4350
rect 2869 4341 2873 4345
rect 2779 4336 2783 4340
rect 2784 4336 2788 4340
rect 2789 4336 2793 4340
rect 2794 4336 2798 4340
rect 2799 4336 2803 4340
rect 2804 4336 2808 4340
rect 2809 4336 2813 4340
rect 2814 4336 2818 4340
rect 2819 4336 2823 4340
rect 2824 4336 2828 4340
rect 2829 4336 2833 4340
rect 2834 4336 2838 4340
rect 2839 4336 2843 4340
rect 2844 4336 2848 4340
rect 2849 4336 2853 4340
rect 2854 4336 2858 4340
rect 2859 4336 2863 4340
rect 2864 4336 2868 4340
rect 2869 4336 2873 4340
rect 2941 4458 2945 4462
rect 2948 4458 2952 4462
rect 2953 4458 2957 4462
rect 2958 4458 2962 4462
rect 2963 4458 2967 4462
rect 2968 4458 2972 4462
rect 2973 4458 2977 4462
rect 2978 4458 2982 4462
rect 2983 4458 2987 4462
rect 2988 4458 2992 4462
rect 2993 4458 2997 4462
rect 2998 4458 3002 4462
rect 3005 4458 3009 4462
rect 2941 4451 2945 4455
rect 3005 4451 3009 4455
rect 2941 4446 2945 4450
rect 2941 4441 2945 4445
rect 2941 4436 2945 4440
rect 2941 4431 2945 4435
rect 2941 4426 2945 4430
rect 2941 4421 2945 4425
rect 2941 4416 2945 4420
rect 2941 4411 2945 4415
rect 2941 4406 2945 4410
rect 2941 4401 2945 4405
rect 2941 4396 2945 4400
rect 2941 4391 2945 4395
rect 2941 4386 2945 4390
rect 2941 4381 2945 4385
rect 2941 4376 2945 4380
rect 2941 4371 2945 4375
rect 2941 4366 2945 4370
rect 2941 4361 2945 4365
rect 3005 4446 3009 4450
rect 3005 4441 3009 4445
rect 3005 4436 3009 4440
rect 3005 4431 3009 4435
rect 3005 4426 3009 4430
rect 3005 4421 3009 4425
rect 3005 4416 3009 4420
rect 3005 4411 3009 4415
rect 3005 4406 3009 4410
rect 3005 4401 3009 4405
rect 3005 4396 3009 4400
rect 3005 4391 3009 4395
rect 3005 4386 3009 4390
rect 3005 4381 3009 4385
rect 3005 4376 3009 4380
rect 3005 4371 3009 4375
rect 3005 4366 3009 4370
rect 3005 4361 3009 4365
rect 2941 4356 2945 4360
rect 3005 4356 3009 4360
rect 2941 4349 2945 4353
rect 2948 4349 2952 4353
rect 2953 4349 2957 4353
rect 2958 4349 2962 4353
rect 2963 4349 2967 4353
rect 2968 4349 2972 4353
rect 2973 4349 2977 4353
rect 2978 4349 2982 4353
rect 2983 4349 2987 4353
rect 2988 4349 2992 4353
rect 2993 4349 2997 4353
rect 2998 4349 3002 4353
rect 3005 4349 3009 4353
rect 3088 4471 3092 4475
rect 3093 4471 3097 4475
rect 3098 4471 3102 4475
rect 3103 4471 3107 4475
rect 3108 4471 3112 4475
rect 3113 4471 3117 4475
rect 3118 4471 3122 4475
rect 3123 4471 3127 4475
rect 3128 4471 3132 4475
rect 3133 4471 3137 4475
rect 3138 4471 3142 4475
rect 3143 4471 3147 4475
rect 3148 4471 3152 4475
rect 3153 4471 3157 4475
rect 3158 4471 3162 4475
rect 3163 4471 3167 4475
rect 3168 4471 3172 4475
rect 3173 4471 3177 4475
rect 3178 4471 3182 4475
rect 3088 4466 3092 4470
rect 3088 4461 3092 4465
rect 3178 4466 3182 4470
rect 3088 4456 3092 4460
rect 3088 4451 3092 4455
rect 3088 4446 3092 4450
rect 3088 4441 3092 4445
rect 3088 4436 3092 4440
rect 3088 4431 3092 4435
rect 3088 4426 3092 4430
rect 3088 4421 3092 4425
rect 3088 4416 3092 4420
rect 3088 4411 3092 4415
rect 3088 4406 3092 4410
rect 3088 4401 3092 4405
rect 3088 4396 3092 4400
rect 3088 4391 3092 4395
rect 3088 4386 3092 4390
rect 3088 4381 3092 4385
rect 3088 4376 3092 4380
rect 3088 4371 3092 4375
rect 3088 4366 3092 4370
rect 3088 4361 3092 4365
rect 3088 4356 3092 4360
rect 3088 4351 3092 4355
rect 3088 4346 3092 4350
rect 3178 4461 3182 4465
rect 3178 4456 3182 4460
rect 3178 4451 3182 4455
rect 3178 4446 3182 4450
rect 3178 4441 3182 4445
rect 3178 4436 3182 4440
rect 3178 4431 3182 4435
rect 3178 4426 3182 4430
rect 3178 4421 3182 4425
rect 3178 4416 3182 4420
rect 3178 4411 3182 4415
rect 3178 4406 3182 4410
rect 3178 4401 3182 4405
rect 3178 4396 3182 4400
rect 3178 4391 3182 4395
rect 3178 4386 3182 4390
rect 3178 4381 3182 4385
rect 3178 4376 3182 4380
rect 3178 4371 3182 4375
rect 3178 4366 3182 4370
rect 3178 4361 3182 4365
rect 3178 4356 3182 4360
rect 3178 4351 3182 4355
rect 3088 4341 3092 4345
rect 3178 4346 3182 4350
rect 3178 4341 3182 4345
rect 3088 4336 3092 4340
rect 3093 4336 3097 4340
rect 3098 4336 3102 4340
rect 3103 4336 3107 4340
rect 3108 4336 3112 4340
rect 3113 4336 3117 4340
rect 3118 4336 3122 4340
rect 3123 4336 3127 4340
rect 3128 4336 3132 4340
rect 3133 4336 3137 4340
rect 3138 4336 3142 4340
rect 3143 4336 3147 4340
rect 3148 4336 3152 4340
rect 3153 4336 3157 4340
rect 3158 4336 3162 4340
rect 3163 4336 3167 4340
rect 3168 4336 3172 4340
rect 3173 4336 3177 4340
rect 3178 4336 3182 4340
rect 3250 4458 3254 4462
rect 3257 4458 3261 4462
rect 3262 4458 3266 4462
rect 3267 4458 3271 4462
rect 3272 4458 3276 4462
rect 3277 4458 3281 4462
rect 3282 4458 3286 4462
rect 3287 4458 3291 4462
rect 3292 4458 3296 4462
rect 3297 4458 3301 4462
rect 3302 4458 3306 4462
rect 3307 4458 3311 4462
rect 3314 4458 3318 4462
rect 3250 4451 3254 4455
rect 3314 4451 3318 4455
rect 3250 4446 3254 4450
rect 3250 4441 3254 4445
rect 3250 4436 3254 4440
rect 3250 4431 3254 4435
rect 3250 4426 3254 4430
rect 3250 4421 3254 4425
rect 3250 4416 3254 4420
rect 3250 4411 3254 4415
rect 3250 4406 3254 4410
rect 3250 4401 3254 4405
rect 3250 4396 3254 4400
rect 3250 4391 3254 4395
rect 3250 4386 3254 4390
rect 3250 4381 3254 4385
rect 3250 4376 3254 4380
rect 3250 4371 3254 4375
rect 3250 4366 3254 4370
rect 3250 4361 3254 4365
rect 3314 4446 3318 4450
rect 3314 4441 3318 4445
rect 3314 4436 3318 4440
rect 3314 4431 3318 4435
rect 3314 4426 3318 4430
rect 3314 4421 3318 4425
rect 3314 4416 3318 4420
rect 3314 4411 3318 4415
rect 3314 4406 3318 4410
rect 3314 4401 3318 4405
rect 3314 4396 3318 4400
rect 3314 4391 3318 4395
rect 3314 4386 3318 4390
rect 3314 4381 3318 4385
rect 3314 4376 3318 4380
rect 3314 4371 3318 4375
rect 3314 4366 3318 4370
rect 3314 4361 3318 4365
rect 3250 4356 3254 4360
rect 3314 4356 3318 4360
rect 3250 4349 3254 4353
rect 3257 4349 3261 4353
rect 3262 4349 3266 4353
rect 3267 4349 3271 4353
rect 3272 4349 3276 4353
rect 3277 4349 3281 4353
rect 3282 4349 3286 4353
rect 3287 4349 3291 4353
rect 3292 4349 3296 4353
rect 3297 4349 3301 4353
rect 3302 4349 3306 4353
rect 3307 4349 3311 4353
rect 3314 4349 3318 4353
rect 3397 4471 3401 4475
rect 3402 4471 3406 4475
rect 3407 4471 3411 4475
rect 3412 4471 3416 4475
rect 3417 4471 3421 4475
rect 3422 4471 3426 4475
rect 3427 4471 3431 4475
rect 3432 4471 3436 4475
rect 3437 4471 3441 4475
rect 3442 4471 3446 4475
rect 3447 4471 3451 4475
rect 3452 4471 3456 4475
rect 3457 4471 3461 4475
rect 3462 4471 3466 4475
rect 3467 4471 3471 4475
rect 3472 4471 3476 4475
rect 3477 4471 3481 4475
rect 3482 4471 3486 4475
rect 3487 4471 3491 4475
rect 3397 4466 3401 4470
rect 3397 4461 3401 4465
rect 3487 4466 3491 4470
rect 3397 4456 3401 4460
rect 3397 4451 3401 4455
rect 3397 4446 3401 4450
rect 3397 4441 3401 4445
rect 3397 4436 3401 4440
rect 3397 4431 3401 4435
rect 3397 4426 3401 4430
rect 3397 4421 3401 4425
rect 3397 4416 3401 4420
rect 3397 4411 3401 4415
rect 3397 4406 3401 4410
rect 3397 4401 3401 4405
rect 3397 4396 3401 4400
rect 3397 4391 3401 4395
rect 3397 4386 3401 4390
rect 3397 4381 3401 4385
rect 3397 4376 3401 4380
rect 3397 4371 3401 4375
rect 3397 4366 3401 4370
rect 3397 4361 3401 4365
rect 3397 4356 3401 4360
rect 3397 4351 3401 4355
rect 3397 4346 3401 4350
rect 3487 4461 3491 4465
rect 3487 4456 3491 4460
rect 3487 4451 3491 4455
rect 3487 4446 3491 4450
rect 3487 4441 3491 4445
rect 3487 4436 3491 4440
rect 3487 4431 3491 4435
rect 3487 4426 3491 4430
rect 3487 4421 3491 4425
rect 3487 4416 3491 4420
rect 3487 4411 3491 4415
rect 3487 4406 3491 4410
rect 3487 4401 3491 4405
rect 3487 4396 3491 4400
rect 3487 4391 3491 4395
rect 3487 4386 3491 4390
rect 3487 4381 3491 4385
rect 3487 4376 3491 4380
rect 3487 4371 3491 4375
rect 3487 4366 3491 4370
rect 3487 4361 3491 4365
rect 3487 4356 3491 4360
rect 3487 4351 3491 4355
rect 3397 4341 3401 4345
rect 3487 4346 3491 4350
rect 3487 4341 3491 4345
rect 3397 4336 3401 4340
rect 3402 4336 3406 4340
rect 3407 4336 3411 4340
rect 3412 4336 3416 4340
rect 3417 4336 3421 4340
rect 3422 4336 3426 4340
rect 3427 4336 3431 4340
rect 3432 4336 3436 4340
rect 3437 4336 3441 4340
rect 3442 4336 3446 4340
rect 3447 4336 3451 4340
rect 3452 4336 3456 4340
rect 3457 4336 3461 4340
rect 3462 4336 3466 4340
rect 3467 4336 3471 4340
rect 3472 4336 3476 4340
rect 3477 4336 3481 4340
rect 3482 4336 3486 4340
rect 3487 4336 3491 4340
rect 3559 4458 3563 4462
rect 3566 4458 3570 4462
rect 3571 4458 3575 4462
rect 3576 4458 3580 4462
rect 3581 4458 3585 4462
rect 3586 4458 3590 4462
rect 3591 4458 3595 4462
rect 3596 4458 3600 4462
rect 3601 4458 3605 4462
rect 3606 4458 3610 4462
rect 3611 4458 3615 4462
rect 3616 4458 3620 4462
rect 3623 4458 3627 4462
rect 3559 4451 3563 4455
rect 3623 4451 3627 4455
rect 3559 4446 3563 4450
rect 3559 4441 3563 4445
rect 3559 4436 3563 4440
rect 3559 4431 3563 4435
rect 3559 4426 3563 4430
rect 3559 4421 3563 4425
rect 3559 4416 3563 4420
rect 3559 4411 3563 4415
rect 3559 4406 3563 4410
rect 3559 4401 3563 4405
rect 3559 4396 3563 4400
rect 3559 4391 3563 4395
rect 3559 4386 3563 4390
rect 3559 4381 3563 4385
rect 3559 4376 3563 4380
rect 3559 4371 3563 4375
rect 3559 4366 3563 4370
rect 3559 4361 3563 4365
rect 3623 4446 3627 4450
rect 3623 4441 3627 4445
rect 3623 4436 3627 4440
rect 3623 4431 3627 4435
rect 3623 4426 3627 4430
rect 3623 4421 3627 4425
rect 3623 4416 3627 4420
rect 3623 4411 3627 4415
rect 3623 4406 3627 4410
rect 3623 4401 3627 4405
rect 3623 4396 3627 4400
rect 3623 4391 3627 4395
rect 3623 4386 3627 4390
rect 3623 4381 3627 4385
rect 3623 4376 3627 4380
rect 3623 4371 3627 4375
rect 3623 4366 3627 4370
rect 3623 4361 3627 4365
rect 3559 4356 3563 4360
rect 3623 4356 3627 4360
rect 3559 4349 3563 4353
rect 3566 4349 3570 4353
rect 3571 4349 3575 4353
rect 3576 4349 3580 4353
rect 3581 4349 3585 4353
rect 3586 4349 3590 4353
rect 3591 4349 3595 4353
rect 3596 4349 3600 4353
rect 3601 4349 3605 4353
rect 3606 4349 3610 4353
rect 3611 4349 3615 4353
rect 3616 4349 3620 4353
rect 3623 4349 3627 4353
rect 3706 4471 3710 4475
rect 3711 4471 3715 4475
rect 3716 4471 3720 4475
rect 3721 4471 3725 4475
rect 3726 4471 3730 4475
rect 3731 4471 3735 4475
rect 3736 4471 3740 4475
rect 3741 4471 3745 4475
rect 3746 4471 3750 4475
rect 3751 4471 3755 4475
rect 3756 4471 3760 4475
rect 3761 4471 3765 4475
rect 3766 4471 3770 4475
rect 3771 4471 3775 4475
rect 3776 4471 3780 4475
rect 3781 4471 3785 4475
rect 3786 4471 3790 4475
rect 3791 4471 3795 4475
rect 3796 4471 3800 4475
rect 3706 4466 3710 4470
rect 3706 4461 3710 4465
rect 3796 4466 3800 4470
rect 3706 4456 3710 4460
rect 3706 4451 3710 4455
rect 3706 4446 3710 4450
rect 3706 4441 3710 4445
rect 3706 4436 3710 4440
rect 3706 4431 3710 4435
rect 3706 4426 3710 4430
rect 3706 4421 3710 4425
rect 3706 4416 3710 4420
rect 3706 4411 3710 4415
rect 3706 4406 3710 4410
rect 3706 4401 3710 4405
rect 3706 4396 3710 4400
rect 3706 4391 3710 4395
rect 3706 4386 3710 4390
rect 3706 4381 3710 4385
rect 3706 4376 3710 4380
rect 3706 4371 3710 4375
rect 3706 4366 3710 4370
rect 3706 4361 3710 4365
rect 3706 4356 3710 4360
rect 3706 4351 3710 4355
rect 3706 4346 3710 4350
rect 3796 4461 3800 4465
rect 3796 4456 3800 4460
rect 3796 4451 3800 4455
rect 3796 4446 3800 4450
rect 3796 4441 3800 4445
rect 3796 4436 3800 4440
rect 3796 4431 3800 4435
rect 3796 4426 3800 4430
rect 3796 4421 3800 4425
rect 3796 4416 3800 4420
rect 3796 4411 3800 4415
rect 3796 4406 3800 4410
rect 3796 4401 3800 4405
rect 3796 4396 3800 4400
rect 3796 4391 3800 4395
rect 3796 4386 3800 4390
rect 3796 4381 3800 4385
rect 3796 4376 3800 4380
rect 3796 4371 3800 4375
rect 3796 4366 3800 4370
rect 3796 4361 3800 4365
rect 3796 4356 3800 4360
rect 3796 4351 3800 4355
rect 3706 4341 3710 4345
rect 3796 4346 3800 4350
rect 3796 4341 3800 4345
rect 3706 4336 3710 4340
rect 3711 4336 3715 4340
rect 3716 4336 3720 4340
rect 3721 4336 3725 4340
rect 3726 4336 3730 4340
rect 3731 4336 3735 4340
rect 3736 4336 3740 4340
rect 3741 4336 3745 4340
rect 3746 4336 3750 4340
rect 3751 4336 3755 4340
rect 3756 4336 3760 4340
rect 3761 4336 3765 4340
rect 3766 4336 3770 4340
rect 3771 4336 3775 4340
rect 3776 4336 3780 4340
rect 3781 4336 3785 4340
rect 3786 4336 3790 4340
rect 3791 4336 3795 4340
rect 3796 4336 3800 4340
<< polysilicon >>
rect 118 9786 1024 10280
rect 1797 9883 1818 9952
rect 2106 9883 2127 9952
rect 2415 9883 2436 9952
rect 2724 9883 2745 9952
rect 3033 9883 3054 9952
rect 3960 9883 3981 9952
rect 1803 9826 1812 9827
rect 2112 9826 2121 9827
rect 2421 9826 2430 9827
rect 2730 9826 2739 9827
rect 3039 9826 3048 9827
rect 3966 9826 3975 9827
rect 1741 9824 1743 9826
rect 1799 9824 1829 9826
rect 1869 9824 1871 9826
rect 2050 9824 2052 9826
rect 2108 9824 2138 9826
rect 2178 9824 2180 9826
rect 2359 9824 2361 9826
rect 2417 9824 2447 9826
rect 2487 9824 2489 9826
rect 2668 9824 2670 9826
rect 2726 9824 2756 9826
rect 2796 9824 2798 9826
rect 2977 9824 2979 9826
rect 3035 9824 3065 9826
rect 3105 9824 3107 9826
rect 3904 9824 3906 9826
rect 3962 9824 3992 9826
rect 4032 9824 4034 9826
rect 1806 9818 1808 9824
rect 2115 9818 2117 9824
rect 2424 9818 2426 9824
rect 2733 9818 2735 9824
rect 3042 9818 3044 9824
rect 3969 9818 3971 9824
rect 1741 9816 1743 9818
rect 1799 9816 1829 9818
rect 1869 9816 1871 9818
rect 2050 9816 2052 9818
rect 2108 9816 2138 9818
rect 2178 9816 2180 9818
rect 2359 9816 2361 9818
rect 2417 9816 2447 9818
rect 2487 9816 2489 9818
rect 2668 9816 2670 9818
rect 2726 9816 2756 9818
rect 2796 9816 2798 9818
rect 2977 9816 2979 9818
rect 3035 9816 3065 9818
rect 3105 9816 3107 9818
rect 3904 9816 3906 9818
rect 3962 9816 3992 9818
rect 4032 9816 4034 9818
rect 1740 9808 1743 9810
rect 1799 9808 1813 9810
rect 1819 9808 1829 9810
rect 1869 9808 1872 9810
rect 1740 9802 1742 9808
rect 1800 9806 1828 9808
rect 1800 9802 1802 9806
rect 1740 9800 1743 9802
rect 1799 9800 1802 9802
rect 1740 9794 1742 9800
rect 1800 9794 1802 9800
rect 1740 9792 1743 9794
rect 1799 9792 1802 9794
rect 1740 9786 1742 9792
rect 1800 9786 1802 9792
rect 118 9348 593 9786
rect 1740 9784 1743 9786
rect 1799 9784 1802 9786
rect 1826 9802 1828 9806
rect 1870 9802 1872 9808
rect 1826 9800 1829 9802
rect 1869 9800 1872 9802
rect 1826 9794 1828 9800
rect 1870 9794 1872 9800
rect 1826 9792 1829 9794
rect 1869 9792 1872 9794
rect 1826 9786 1828 9792
rect 1870 9786 1872 9792
rect 1826 9784 1829 9786
rect 1869 9784 1872 9786
rect 2049 9808 2052 9810
rect 2108 9808 2122 9810
rect 2128 9808 2138 9810
rect 2178 9808 2181 9810
rect 2049 9802 2051 9808
rect 2109 9806 2137 9808
rect 2109 9802 2111 9806
rect 2049 9800 2052 9802
rect 2108 9800 2111 9802
rect 2049 9794 2051 9800
rect 2109 9794 2111 9800
rect 2049 9792 2052 9794
rect 2108 9792 2111 9794
rect 2049 9786 2051 9792
rect 2109 9786 2111 9792
rect 2049 9784 2052 9786
rect 2108 9784 2111 9786
rect 2135 9802 2137 9806
rect 2179 9802 2181 9808
rect 2135 9800 2138 9802
rect 2178 9800 2181 9802
rect 2135 9794 2137 9800
rect 2179 9794 2181 9800
rect 2135 9792 2138 9794
rect 2178 9792 2181 9794
rect 2135 9786 2137 9792
rect 2179 9786 2181 9792
rect 2135 9784 2138 9786
rect 2178 9784 2181 9786
rect 2358 9808 2361 9810
rect 2417 9808 2431 9810
rect 2437 9808 2447 9810
rect 2487 9808 2490 9810
rect 2358 9802 2360 9808
rect 2418 9806 2446 9808
rect 2418 9802 2420 9806
rect 2358 9800 2361 9802
rect 2417 9800 2420 9802
rect 2358 9794 2360 9800
rect 2418 9794 2420 9800
rect 2358 9792 2361 9794
rect 2417 9792 2420 9794
rect 2358 9786 2360 9792
rect 2418 9786 2420 9792
rect 2358 9784 2361 9786
rect 2417 9784 2420 9786
rect 2444 9802 2446 9806
rect 2488 9802 2490 9808
rect 2444 9800 2447 9802
rect 2487 9800 2490 9802
rect 2444 9794 2446 9800
rect 2488 9794 2490 9800
rect 2444 9792 2447 9794
rect 2487 9792 2490 9794
rect 2444 9786 2446 9792
rect 2488 9786 2490 9792
rect 2444 9784 2447 9786
rect 2487 9784 2490 9786
rect 2667 9808 2670 9810
rect 2726 9808 2740 9810
rect 2746 9808 2756 9810
rect 2796 9808 2799 9810
rect 2667 9802 2669 9808
rect 2727 9806 2755 9808
rect 2727 9802 2729 9806
rect 2667 9800 2670 9802
rect 2726 9800 2729 9802
rect 2667 9794 2669 9800
rect 2727 9794 2729 9800
rect 2667 9792 2670 9794
rect 2726 9792 2729 9794
rect 2667 9786 2669 9792
rect 2727 9786 2729 9792
rect 2667 9784 2670 9786
rect 2726 9784 2729 9786
rect 2753 9802 2755 9806
rect 2797 9802 2799 9808
rect 2753 9800 2756 9802
rect 2796 9800 2799 9802
rect 2753 9794 2755 9800
rect 2797 9794 2799 9800
rect 2753 9792 2756 9794
rect 2796 9792 2799 9794
rect 2753 9786 2755 9792
rect 2797 9786 2799 9792
rect 2753 9784 2756 9786
rect 2796 9784 2799 9786
rect 2976 9808 2979 9810
rect 3035 9808 3049 9810
rect 3055 9808 3065 9810
rect 3105 9808 3108 9810
rect 2976 9802 2978 9808
rect 3036 9806 3064 9808
rect 3036 9802 3038 9806
rect 2976 9800 2979 9802
rect 3035 9800 3038 9802
rect 2976 9794 2978 9800
rect 3036 9794 3038 9800
rect 2976 9792 2979 9794
rect 3035 9792 3038 9794
rect 2976 9786 2978 9792
rect 3036 9786 3038 9792
rect 2976 9784 2979 9786
rect 3035 9784 3038 9786
rect 3062 9802 3064 9806
rect 3106 9802 3108 9808
rect 3062 9800 3065 9802
rect 3105 9800 3108 9802
rect 3062 9794 3064 9800
rect 3106 9794 3108 9800
rect 3062 9792 3065 9794
rect 3105 9792 3108 9794
rect 3062 9786 3064 9792
rect 3106 9786 3108 9792
rect 3062 9784 3065 9786
rect 3105 9784 3108 9786
rect 3903 9808 3906 9810
rect 3962 9808 3976 9810
rect 3982 9808 3992 9810
rect 4032 9808 4035 9810
rect 3903 9802 3905 9808
rect 3963 9806 3991 9808
rect 3963 9802 3965 9806
rect 3903 9800 3906 9802
rect 3962 9800 3965 9802
rect 3903 9794 3905 9800
rect 3963 9794 3965 9800
rect 3903 9792 3906 9794
rect 3962 9792 3965 9794
rect 3903 9786 3905 9792
rect 3963 9786 3965 9792
rect 3903 9784 3906 9786
rect 3962 9784 3965 9786
rect 3989 9802 3991 9806
rect 4033 9802 4035 9808
rect 3989 9800 3992 9802
rect 4032 9800 4035 9802
rect 3989 9794 3991 9800
rect 4033 9794 4035 9800
rect 3989 9792 3992 9794
rect 4032 9792 4035 9794
rect 3989 9786 3991 9792
rect 4033 9786 4035 9792
rect 4141 9786 5073 10261
rect 3989 9784 3992 9786
rect 4032 9784 4035 9786
rect 428 6458 454 6460
rect 428 6457 430 6458
rect 436 6457 438 6458
rect 444 6457 446 6458
rect 452 6457 454 6458
rect 469 6458 495 6460
rect 469 6457 471 6458
rect 477 6457 479 6458
rect 485 6457 487 6458
rect 493 6457 495 6458
rect 512 6458 538 6460
rect 512 6457 514 6458
rect 520 6457 522 6458
rect 528 6457 530 6458
rect 536 6457 538 6458
rect 551 6426 577 6428
rect 551 6425 553 6426
rect 559 6425 561 6426
rect 567 6425 569 6426
rect 575 6425 577 6426
rect 583 6425 585 6427
rect 591 6425 593 6427
rect 428 6366 430 6369
rect 436 6366 438 6369
rect 444 6366 446 6369
rect 452 6366 454 6369
rect 428 6364 454 6366
rect 469 6366 471 6369
rect 477 6366 479 6369
rect 485 6366 487 6369
rect 493 6366 495 6369
rect 512 6368 514 6369
rect 520 6368 522 6369
rect 528 6368 530 6369
rect 536 6368 538 6369
rect 512 6366 538 6368
rect 551 6368 553 6369
rect 559 6368 561 6369
rect 567 6368 569 6369
rect 575 6368 577 6369
rect 551 6366 577 6368
rect 469 6364 495 6366
rect 428 6362 495 6364
rect 428 6360 490 6362
rect 428 6351 455 6360
rect 461 6351 490 6360
rect 428 6349 490 6351
rect 494 6349 495 6362
rect 428 6340 495 6349
rect 531 6364 538 6366
rect 531 6351 533 6364
rect 537 6351 538 6364
rect 531 6342 538 6351
rect 573 6355 577 6366
rect 583 6362 585 6369
rect 591 6362 593 6369
rect 583 6360 593 6362
rect 573 6349 575 6355
rect 573 6342 577 6349
rect 428 6339 430 6340
rect 436 6339 438 6340
rect 444 6339 446 6340
rect 452 6339 454 6340
rect 469 6339 471 6340
rect 477 6339 479 6340
rect 485 6339 487 6340
rect 493 6339 495 6340
rect 512 6340 538 6342
rect 512 6339 514 6340
rect 520 6339 522 6340
rect 528 6339 530 6340
rect 536 6339 538 6340
rect 551 6340 577 6342
rect 551 6339 553 6340
rect 559 6339 561 6340
rect 567 6339 569 6340
rect 575 6339 577 6340
rect 583 6339 585 6360
rect 591 6354 596 6360
rect 591 6339 593 6354
rect 551 6298 553 6299
rect 559 6298 561 6299
rect 567 6298 569 6299
rect 575 6298 577 6299
rect 551 6296 577 6298
rect 583 6297 585 6299
rect 591 6297 593 6299
rect 428 6279 430 6280
rect 436 6279 438 6280
rect 428 6277 438 6279
rect 444 6279 446 6280
rect 452 6279 454 6280
rect 444 6277 454 6279
rect 469 6279 471 6280
rect 477 6279 479 6280
rect 469 6277 479 6279
rect 485 6279 487 6280
rect 493 6279 495 6280
rect 485 6277 495 6279
rect 512 6279 514 6280
rect 520 6279 522 6280
rect 512 6277 522 6279
rect 528 6279 530 6280
rect 536 6279 538 6280
rect 528 6277 538 6279
rect 99 4528 593 4959
rect 2856 9330 2858 9332
rect 2861 9330 2863 9333
rect 2877 9330 2879 9332
rect 2893 9330 2895 9332
rect 2898 9330 2900 9333
rect 2919 9330 2921 9333
rect 2935 9330 2937 9333
rect 2951 9330 2953 9332
rect 2956 9330 2958 9333
rect 2972 9330 2974 9332
rect 2988 9330 2990 9332
rect 2993 9330 2995 9333
rect 3009 9330 3011 9332
rect 3025 9330 3027 9332
rect 3030 9330 3032 9333
rect 3051 9330 3053 9333
rect 3067 9330 3069 9333
rect 3083 9330 3085 9332
rect 3088 9330 3090 9333
rect 3104 9330 3106 9332
rect 3120 9330 3122 9332
rect 3125 9330 3127 9333
rect 3141 9330 3143 9332
rect 3157 9330 3159 9332
rect 3162 9330 3164 9333
rect 3183 9330 3185 9333
rect 3199 9330 3201 9333
rect 3215 9330 3217 9332
rect 3220 9330 3222 9333
rect 3236 9330 3238 9332
rect 3252 9330 3254 9332
rect 3257 9330 3259 9333
rect 3273 9330 3275 9332
rect 3289 9330 3291 9332
rect 3294 9330 3296 9333
rect 3315 9330 3317 9333
rect 3331 9330 3333 9333
rect 3347 9330 3349 9332
rect 3352 9330 3354 9333
rect 3368 9330 3370 9332
rect 3801 9330 3803 9332
rect 3806 9330 3808 9333
rect 3822 9330 3824 9332
rect 3838 9330 3840 9332
rect 3843 9330 3845 9333
rect 3864 9330 3866 9333
rect 3880 9330 3882 9333
rect 3896 9330 3898 9332
rect 3901 9330 3903 9333
rect 3917 9330 3919 9332
rect 3933 9330 3935 9332
rect 3938 9330 3940 9333
rect 3954 9330 3956 9332
rect 3970 9330 3972 9332
rect 3975 9330 3977 9333
rect 3996 9330 3998 9333
rect 4012 9330 4014 9333
rect 4028 9330 4030 9332
rect 4033 9330 4035 9333
rect 4049 9330 4051 9332
rect 4065 9330 4067 9332
rect 4070 9330 4072 9333
rect 4086 9330 4088 9332
rect 4102 9330 4104 9332
rect 4107 9330 4109 9333
rect 4128 9330 4130 9333
rect 4144 9330 4146 9333
rect 4160 9330 4162 9332
rect 4165 9330 4167 9333
rect 4181 9330 4183 9332
rect 4197 9330 4199 9332
rect 4202 9330 4204 9333
rect 4218 9330 4220 9332
rect 4234 9330 4236 9332
rect 4239 9330 4241 9333
rect 4260 9330 4262 9333
rect 4276 9330 4278 9333
rect 4292 9330 4294 9332
rect 4297 9330 4299 9333
rect 4313 9330 4315 9332
rect 2856 9317 2858 9322
rect 2861 9320 2863 9322
rect 2856 9303 2858 9313
rect 2861 9303 2863 9310
rect 2877 9303 2879 9322
rect 2893 9313 2895 9322
rect 2898 9320 2900 9322
rect 2919 9320 2921 9322
rect 2935 9319 2937 9322
rect 2893 9303 2895 9306
rect 2898 9303 2900 9305
rect 2919 9303 2921 9305
rect 2935 9303 2937 9315
rect 2951 9313 2953 9322
rect 2956 9320 2958 9322
rect 2972 9314 2974 9322
rect 2988 9317 2990 9322
rect 2993 9320 2995 9322
rect 2951 9303 2953 9306
rect 2956 9303 2958 9305
rect 2972 9303 2974 9310
rect 2988 9303 2990 9313
rect 2993 9303 2995 9310
rect 3009 9303 3011 9322
rect 3025 9313 3027 9322
rect 3030 9320 3032 9322
rect 3051 9320 3053 9322
rect 3067 9319 3069 9322
rect 3025 9303 3027 9306
rect 3030 9303 3032 9305
rect 3051 9303 3053 9305
rect 3067 9303 3069 9315
rect 3083 9313 3085 9322
rect 3088 9320 3090 9322
rect 3104 9314 3106 9322
rect 3120 9317 3122 9322
rect 3125 9320 3127 9322
rect 3083 9303 3085 9306
rect 3088 9303 3090 9305
rect 3104 9303 3106 9310
rect 3120 9303 3122 9313
rect 3125 9303 3127 9310
rect 3141 9303 3143 9322
rect 3157 9313 3159 9322
rect 3162 9320 3164 9322
rect 3183 9320 3185 9322
rect 3199 9319 3201 9322
rect 3157 9303 3159 9306
rect 3162 9303 3164 9305
rect 3183 9303 3185 9305
rect 3199 9303 3201 9315
rect 3215 9313 3217 9322
rect 3220 9320 3222 9322
rect 3236 9314 3238 9322
rect 3252 9317 3254 9322
rect 3257 9320 3259 9322
rect 3215 9303 3217 9306
rect 3220 9303 3222 9305
rect 3236 9303 3238 9310
rect 3252 9303 3254 9313
rect 3257 9303 3259 9310
rect 3273 9303 3275 9322
rect 3289 9313 3291 9322
rect 3294 9320 3296 9322
rect 3315 9320 3317 9322
rect 3331 9319 3333 9322
rect 3289 9303 3291 9306
rect 3294 9303 3296 9305
rect 3315 9303 3317 9305
rect 3331 9303 3333 9315
rect 3347 9313 3349 9322
rect 3352 9320 3354 9322
rect 3368 9314 3370 9322
rect 3801 9317 3803 9322
rect 3806 9320 3808 9322
rect 3347 9303 3349 9306
rect 3352 9303 3354 9305
rect 3368 9303 3370 9310
rect 2504 9297 2506 9299
rect 2509 9297 2511 9300
rect 2525 9297 2527 9299
rect 2541 9297 2543 9299
rect 2546 9297 2548 9300
rect 2567 9297 2569 9300
rect 2583 9297 2585 9300
rect 2599 9297 2601 9299
rect 2604 9297 2606 9300
rect 3801 9303 3803 9313
rect 3806 9303 3808 9310
rect 3822 9303 3824 9322
rect 3838 9313 3840 9322
rect 3843 9320 3845 9322
rect 3864 9320 3866 9322
rect 3880 9319 3882 9322
rect 3838 9303 3840 9306
rect 3843 9303 3845 9305
rect 3864 9303 3866 9305
rect 3880 9303 3882 9315
rect 3896 9313 3898 9322
rect 3901 9320 3903 9322
rect 3917 9314 3919 9322
rect 3933 9317 3935 9322
rect 3938 9320 3940 9322
rect 3896 9303 3898 9306
rect 3901 9303 3903 9305
rect 3917 9303 3919 9310
rect 3933 9303 3935 9313
rect 3938 9303 3940 9310
rect 3954 9303 3956 9322
rect 3970 9313 3972 9322
rect 3975 9320 3977 9322
rect 3996 9320 3998 9322
rect 4012 9319 4014 9322
rect 3970 9303 3972 9306
rect 3975 9303 3977 9305
rect 3996 9303 3998 9305
rect 4012 9303 4014 9315
rect 4028 9313 4030 9322
rect 4033 9320 4035 9322
rect 4049 9314 4051 9322
rect 4065 9317 4067 9322
rect 4070 9320 4072 9322
rect 4028 9303 4030 9306
rect 4033 9303 4035 9305
rect 4049 9303 4051 9310
rect 4065 9303 4067 9313
rect 4070 9303 4072 9310
rect 4086 9303 4088 9322
rect 4102 9313 4104 9322
rect 4107 9320 4109 9322
rect 4128 9320 4130 9322
rect 4144 9319 4146 9322
rect 4102 9303 4104 9306
rect 4107 9303 4109 9305
rect 4128 9303 4130 9305
rect 4144 9303 4146 9315
rect 4160 9313 4162 9322
rect 4165 9320 4167 9322
rect 4181 9314 4183 9322
rect 4197 9317 4199 9322
rect 4202 9320 4204 9322
rect 4160 9303 4162 9306
rect 4165 9303 4167 9305
rect 4181 9303 4183 9310
rect 4197 9303 4199 9313
rect 4202 9303 4204 9310
rect 4218 9303 4220 9322
rect 4234 9313 4236 9322
rect 4239 9320 4241 9322
rect 4260 9320 4262 9322
rect 4276 9319 4278 9322
rect 4234 9303 4236 9306
rect 4239 9303 4241 9305
rect 4260 9303 4262 9305
rect 4276 9303 4278 9315
rect 4292 9313 4294 9322
rect 4297 9320 4299 9322
rect 4313 9314 4315 9322
rect 4292 9303 4294 9306
rect 4297 9303 4299 9305
rect 4313 9303 4315 9310
rect 2620 9297 2622 9299
rect 2856 9297 2858 9299
rect 2861 9296 2863 9299
rect 2877 9297 2879 9299
rect 2893 9297 2895 9299
rect 2898 9294 2900 9299
rect 2919 9294 2921 9299
rect 2935 9297 2937 9299
rect 2951 9297 2953 9299
rect 2956 9294 2958 9299
rect 2972 9297 2974 9299
rect 2988 9297 2990 9299
rect 2993 9296 2995 9299
rect 3009 9297 3011 9299
rect 3025 9297 3027 9299
rect 3030 9294 3032 9299
rect 3051 9294 3053 9299
rect 3067 9297 3069 9299
rect 3083 9297 3085 9299
rect 3088 9294 3090 9299
rect 3104 9297 3106 9299
rect 3120 9297 3122 9299
rect 3125 9296 3127 9299
rect 3141 9297 3143 9299
rect 3157 9297 3159 9299
rect 3162 9294 3164 9299
rect 3183 9294 3185 9299
rect 3199 9297 3201 9299
rect 3215 9297 3217 9299
rect 3220 9294 3222 9299
rect 3236 9297 3238 9299
rect 3252 9297 3254 9299
rect 3257 9296 3259 9299
rect 3273 9297 3275 9299
rect 3289 9297 3291 9299
rect 3294 9294 3296 9299
rect 3315 9294 3317 9299
rect 3331 9297 3333 9299
rect 3347 9297 3349 9299
rect 3352 9294 3354 9299
rect 3368 9297 3370 9299
rect 3449 9297 3451 9299
rect 3454 9297 3456 9300
rect 3470 9297 3472 9299
rect 3486 9297 3488 9299
rect 3491 9297 3493 9300
rect 3512 9297 3514 9300
rect 3528 9297 3530 9300
rect 3544 9297 3546 9299
rect 3549 9297 3551 9300
rect 3565 9297 3567 9299
rect 3801 9297 3803 9299
rect 3806 9296 3808 9299
rect 3822 9297 3824 9299
rect 3838 9297 3840 9299
rect 3843 9294 3845 9299
rect 3864 9294 3866 9299
rect 3880 9297 3882 9299
rect 3896 9297 3898 9299
rect 3901 9294 3903 9299
rect 3917 9297 3919 9299
rect 3933 9297 3935 9299
rect 3938 9296 3940 9299
rect 3954 9297 3956 9299
rect 3970 9297 3972 9299
rect 3975 9294 3977 9299
rect 3996 9294 3998 9299
rect 4012 9297 4014 9299
rect 4028 9297 4030 9299
rect 4033 9294 4035 9299
rect 4049 9297 4051 9299
rect 4065 9297 4067 9299
rect 4070 9296 4072 9299
rect 4086 9297 4088 9299
rect 4102 9297 4104 9299
rect 4107 9294 4109 9299
rect 4128 9294 4130 9299
rect 4144 9297 4146 9299
rect 4160 9297 4162 9299
rect 4165 9294 4167 9299
rect 4181 9297 4183 9299
rect 4197 9297 4199 9299
rect 4202 9296 4204 9299
rect 4218 9297 4220 9299
rect 4234 9297 4236 9299
rect 4239 9294 4241 9299
rect 4260 9294 4262 9299
rect 4276 9297 4278 9299
rect 4292 9297 4294 9299
rect 4297 9294 4299 9299
rect 4313 9297 4315 9299
rect 2504 9284 2506 9289
rect 2509 9287 2511 9289
rect 2504 9270 2506 9280
rect 2509 9270 2511 9277
rect 2525 9270 2527 9289
rect 2541 9280 2543 9289
rect 2546 9287 2548 9289
rect 2567 9287 2569 9289
rect 2583 9286 2585 9289
rect 2541 9270 2543 9273
rect 2546 9270 2548 9272
rect 2567 9270 2569 9272
rect 2583 9270 2585 9282
rect 2599 9280 2601 9289
rect 2604 9287 2606 9289
rect 2599 9270 2601 9273
rect 2604 9270 2606 9272
rect 2620 9270 2622 9289
rect 3449 9284 3451 9289
rect 3454 9287 3456 9289
rect 3449 9270 3451 9280
rect 3454 9270 3456 9277
rect 3470 9270 3472 9289
rect 3486 9280 3488 9289
rect 3491 9287 3493 9289
rect 3512 9287 3514 9289
rect 3528 9286 3530 9289
rect 3486 9270 3488 9273
rect 3491 9270 3493 9272
rect 3512 9270 3514 9272
rect 3528 9270 3530 9282
rect 3544 9280 3546 9289
rect 3549 9287 3551 9289
rect 3544 9270 3546 9273
rect 3549 9270 3551 9272
rect 3565 9270 3567 9289
rect 2504 9264 2506 9266
rect 2509 9263 2511 9266
rect 2525 9264 2527 9266
rect 2541 9264 2543 9266
rect 2546 9261 2548 9266
rect 2567 9261 2569 9266
rect 2583 9264 2585 9266
rect 2599 9264 2601 9266
rect 2604 9261 2606 9266
rect 2620 9264 2622 9266
rect 3449 9264 3451 9266
rect 3454 9263 3456 9266
rect 3470 9264 3472 9266
rect 3486 9264 3488 9266
rect 3035 9259 3037 9261
rect 2877 9253 2879 9256
rect 2921 9253 2923 9256
rect 2947 9253 2949 9256
rect 2993 9253 2995 9256
rect 2947 9249 2948 9253
rect 3061 9253 3063 9257
rect 3089 9259 3091 9261
rect 3116 9259 3118 9261
rect 3066 9253 3068 9256
rect 2861 9246 2863 9248
rect 2877 9246 2879 9249
rect 2893 9246 2895 9248
rect 2916 9246 2918 9248
rect 2921 9246 2923 9249
rect 2947 9246 2949 9249
rect 2968 9246 2970 9249
rect 2988 9246 2990 9248
rect 2993 9246 2995 9249
rect 3011 9246 3013 9248
rect 2628 9233 2630 9236
rect 2628 9227 2630 9229
rect 2511 9224 2513 9227
rect 2861 9224 2863 9238
rect 2877 9236 2879 9238
rect 2877 9224 2879 9226
rect 2893 9224 2895 9238
rect 2916 9233 2918 9238
rect 2921 9236 2923 9238
rect 2947 9236 2949 9238
rect 2912 9229 2918 9233
rect 2916 9224 2918 9229
rect 2921 9224 2923 9226
rect 2947 9224 2949 9226
rect 2968 9224 2970 9238
rect 2988 9233 2990 9238
rect 2993 9236 2995 9238
rect 2984 9229 2990 9233
rect 2988 9224 2990 9229
rect 2993 9224 2995 9226
rect 3011 9224 3013 9238
rect 3035 9237 3037 9251
rect 3142 9253 3144 9257
rect 3170 9259 3172 9261
rect 3491 9261 3493 9266
rect 3512 9261 3514 9266
rect 3528 9264 3530 9266
rect 3544 9264 3546 9266
rect 3549 9261 3551 9266
rect 3565 9264 3567 9266
rect 3147 9253 3149 9256
rect 3061 9242 3063 9245
rect 3066 9243 3068 9245
rect 3062 9238 3063 9242
rect 3061 9233 3063 9238
rect 3066 9233 3068 9235
rect 3035 9231 3037 9233
rect 3089 9229 3091 9251
rect 3116 9237 3118 9251
rect 3980 9259 3982 9261
rect 3142 9242 3144 9245
rect 3147 9243 3149 9245
rect 3143 9238 3144 9242
rect 3142 9233 3144 9238
rect 3147 9233 3149 9235
rect 3116 9231 3118 9233
rect 3170 9229 3172 9251
rect 3822 9253 3824 9256
rect 3866 9253 3868 9256
rect 3892 9253 3894 9256
rect 3938 9253 3940 9256
rect 3892 9249 3893 9253
rect 4006 9253 4008 9257
rect 4034 9259 4036 9261
rect 4061 9259 4063 9261
rect 4011 9253 4013 9256
rect 3806 9246 3808 9248
rect 3822 9246 3824 9249
rect 3838 9246 3840 9248
rect 3861 9246 3863 9248
rect 3866 9246 3868 9249
rect 3892 9246 3894 9249
rect 3913 9246 3915 9249
rect 3933 9246 3935 9248
rect 3938 9246 3940 9249
rect 3956 9246 3958 9248
rect 3573 9233 3575 9236
rect 3061 9227 3063 9229
rect 3066 9224 3068 9229
rect 3142 9227 3144 9229
rect 3089 9223 3091 9225
rect 3147 9224 3149 9229
rect 3573 9227 3575 9229
rect 3170 9223 3172 9225
rect 3456 9224 3458 9227
rect 3806 9224 3808 9238
rect 3822 9236 3824 9238
rect 3822 9224 3824 9226
rect 3838 9224 3840 9238
rect 3861 9233 3863 9238
rect 3866 9236 3868 9238
rect 3892 9236 3894 9238
rect 3857 9229 3863 9233
rect 3861 9224 3863 9229
rect 3866 9224 3868 9226
rect 3892 9224 3894 9226
rect 3913 9224 3915 9238
rect 3933 9233 3935 9238
rect 3938 9236 3940 9238
rect 3929 9229 3935 9233
rect 3933 9224 3935 9229
rect 3938 9224 3940 9226
rect 3956 9224 3958 9238
rect 3980 9237 3982 9251
rect 4087 9253 4089 9257
rect 4115 9259 4117 9261
rect 4092 9253 4094 9256
rect 4006 9242 4008 9245
rect 4011 9243 4013 9245
rect 4007 9238 4008 9242
rect 4006 9233 4008 9238
rect 4011 9233 4013 9235
rect 3980 9231 3982 9233
rect 4034 9229 4036 9251
rect 4061 9237 4063 9251
rect 4087 9242 4089 9245
rect 4092 9243 4094 9245
rect 4088 9238 4089 9242
rect 4087 9233 4089 9238
rect 4092 9233 4094 9235
rect 4061 9231 4063 9233
rect 4115 9229 4117 9251
rect 4006 9227 4008 9229
rect 4011 9224 4013 9229
rect 4087 9227 4089 9229
rect 4034 9223 4036 9225
rect 4092 9224 4094 9229
rect 4115 9223 4117 9225
rect 2511 9218 2513 9220
rect 2861 9218 2863 9220
rect 2877 9216 2879 9220
rect 2893 9218 2895 9220
rect 2916 9218 2918 9220
rect 2878 9212 2879 9216
rect 2921 9215 2923 9220
rect 2947 9216 2949 9220
rect 2968 9218 2970 9220
rect 2988 9218 2990 9220
rect 2877 9209 2879 9212
rect 2922 9211 2923 9215
rect 2948 9212 2949 9216
rect 2993 9215 2995 9220
rect 3011 9218 3013 9220
rect 3456 9218 3458 9220
rect 3806 9218 3808 9220
rect 3822 9216 3824 9220
rect 3838 9218 3840 9220
rect 3861 9218 3863 9220
rect 2921 9209 2923 9211
rect 2947 9208 2949 9212
rect 2994 9211 2995 9215
rect 3823 9212 3824 9216
rect 3866 9215 3868 9220
rect 3892 9216 3894 9220
rect 3913 9218 3915 9220
rect 3933 9218 3935 9220
rect 2993 9209 2995 9211
rect 3822 9209 3824 9212
rect 3867 9211 3868 9215
rect 3893 9212 3894 9216
rect 3938 9215 3940 9220
rect 3956 9218 3958 9220
rect 3866 9209 3868 9211
rect 3892 9208 3894 9212
rect 3939 9211 3940 9215
rect 3938 9209 3940 9211
rect 2495 9195 2497 9197
rect 2511 9195 2513 9198
rect 2516 9195 2518 9197
rect 2532 9195 2534 9198
rect 2548 9195 2550 9198
rect 2569 9195 2571 9198
rect 2574 9195 2576 9197
rect 2590 9195 2592 9197
rect 2606 9195 2608 9198
rect 2611 9195 2613 9197
rect 3440 9195 3442 9197
rect 3456 9195 3458 9198
rect 3461 9195 3463 9197
rect 3477 9195 3479 9198
rect 3493 9195 3495 9198
rect 3514 9195 3516 9198
rect 3519 9195 3521 9197
rect 3535 9195 3537 9197
rect 3551 9195 3553 9198
rect 3556 9195 3558 9197
rect 2495 9168 2497 9187
rect 2511 9185 2513 9187
rect 2516 9178 2518 9187
rect 2532 9184 2534 9187
rect 2548 9185 2550 9187
rect 2569 9185 2571 9187
rect 2511 9168 2513 9170
rect 2516 9168 2518 9171
rect 2532 9168 2534 9180
rect 2574 9178 2576 9187
rect 2548 9168 2550 9170
rect 2569 9168 2571 9170
rect 2574 9168 2576 9171
rect 2590 9168 2592 9187
rect 2606 9185 2608 9187
rect 2611 9182 2613 9187
rect 2877 9186 2879 9189
rect 2921 9187 2923 9189
rect 2878 9182 2879 9186
rect 2922 9183 2923 9187
rect 2947 9186 2949 9190
rect 2993 9187 2995 9189
rect 2861 9178 2863 9180
rect 2877 9178 2879 9182
rect 2893 9178 2895 9180
rect 2916 9178 2918 9180
rect 2921 9178 2923 9183
rect 2948 9182 2949 9186
rect 2994 9183 2995 9187
rect 2947 9178 2949 9182
rect 2968 9178 2970 9180
rect 2988 9178 2990 9180
rect 2993 9178 2995 9183
rect 3011 9178 3013 9180
rect 2606 9168 2608 9175
rect 2611 9168 2613 9178
rect 3061 9177 3063 9180
rect 3066 9177 3068 9180
rect 3142 9177 3144 9180
rect 3147 9177 3149 9180
rect 2495 9162 2497 9164
rect 2511 9159 2513 9164
rect 2516 9162 2518 9164
rect 2532 9162 2534 9164
rect 2548 9159 2550 9164
rect 2569 9159 2571 9164
rect 2574 9162 2576 9164
rect 2590 9162 2592 9164
rect 2606 9161 2608 9164
rect 2611 9162 2613 9164
rect 2861 9160 2863 9174
rect 2877 9172 2879 9174
rect 2877 9160 2879 9162
rect 2893 9160 2895 9174
rect 2916 9169 2918 9174
rect 2921 9172 2923 9174
rect 2947 9172 2949 9174
rect 2912 9165 2918 9169
rect 2916 9160 2918 9165
rect 2921 9160 2923 9162
rect 2947 9160 2949 9162
rect 2968 9160 2970 9174
rect 2988 9169 2990 9174
rect 2993 9172 2995 9174
rect 2984 9165 2990 9169
rect 2988 9160 2990 9165
rect 2993 9160 2995 9162
rect 3011 9160 3013 9174
rect 3061 9161 3063 9173
rect 3066 9171 3068 9173
rect 3066 9161 3068 9163
rect 3142 9161 3144 9173
rect 3147 9171 3149 9173
rect 3440 9168 3442 9187
rect 3456 9185 3458 9187
rect 3461 9178 3463 9187
rect 3477 9184 3479 9187
rect 3493 9185 3495 9187
rect 3514 9185 3516 9187
rect 3456 9168 3458 9170
rect 3461 9168 3463 9171
rect 3477 9168 3479 9180
rect 3519 9178 3521 9187
rect 3493 9168 3495 9170
rect 3514 9168 3516 9170
rect 3519 9168 3521 9171
rect 3535 9168 3537 9187
rect 3551 9185 3553 9187
rect 3556 9182 3558 9187
rect 3822 9186 3824 9189
rect 3866 9187 3868 9189
rect 3823 9182 3824 9186
rect 3867 9183 3868 9187
rect 3892 9186 3894 9190
rect 3938 9187 3940 9189
rect 3806 9178 3808 9180
rect 3822 9178 3824 9182
rect 3838 9178 3840 9180
rect 3861 9178 3863 9180
rect 3866 9178 3868 9183
rect 3893 9182 3894 9186
rect 3939 9183 3940 9187
rect 3892 9178 3894 9182
rect 3913 9178 3915 9180
rect 3933 9178 3935 9180
rect 3938 9178 3940 9183
rect 3956 9178 3958 9180
rect 3551 9168 3553 9175
rect 3556 9168 3558 9178
rect 4006 9177 4008 9180
rect 4011 9177 4013 9180
rect 4087 9177 4089 9180
rect 4092 9177 4094 9180
rect 3147 9161 3149 9163
rect 3440 9162 3442 9164
rect 3456 9159 3458 9164
rect 3461 9162 3463 9164
rect 3477 9162 3479 9164
rect 3493 9159 3495 9164
rect 3514 9159 3516 9164
rect 3519 9162 3521 9164
rect 3535 9162 3537 9164
rect 3551 9161 3553 9164
rect 3556 9162 3558 9164
rect 3806 9160 3808 9174
rect 3822 9172 3824 9174
rect 3822 9160 3824 9162
rect 3838 9160 3840 9174
rect 3861 9169 3863 9174
rect 3866 9172 3868 9174
rect 3892 9172 3894 9174
rect 3857 9165 3863 9169
rect 3861 9160 3863 9165
rect 3866 9160 3868 9162
rect 3892 9160 3894 9162
rect 3913 9160 3915 9174
rect 3933 9169 3935 9174
rect 3938 9172 3940 9174
rect 3929 9165 3935 9169
rect 3933 9160 3935 9165
rect 3938 9160 3940 9162
rect 3956 9160 3958 9174
rect 4006 9161 4008 9173
rect 4011 9171 4013 9173
rect 4011 9161 4013 9163
rect 4087 9161 4089 9173
rect 4092 9171 4094 9173
rect 4092 9161 4094 9163
rect 2861 9150 2863 9152
rect 2877 9149 2879 9152
rect 2893 9150 2895 9152
rect 2916 9150 2918 9152
rect 2921 9149 2923 9152
rect 2947 9149 2949 9152
rect 2968 9149 2970 9152
rect 2988 9150 2990 9152
rect 2993 9149 2995 9152
rect 3011 9150 3013 9152
rect 3061 9151 3063 9153
rect 2947 9145 2948 9149
rect 3066 9148 3068 9153
rect 3142 9151 3144 9153
rect 3147 9148 3149 9153
rect 3806 9150 3808 9152
rect 3822 9149 3824 9152
rect 3838 9150 3840 9152
rect 3861 9150 3863 9152
rect 3866 9149 3868 9152
rect 3892 9149 3894 9152
rect 3913 9149 3915 9152
rect 3933 9150 3935 9152
rect 3938 9149 3940 9152
rect 3956 9150 3958 9152
rect 4006 9151 4008 9153
rect 2877 9142 2879 9145
rect 2921 9142 2923 9145
rect 2947 9142 2949 9145
rect 2993 9142 2995 9145
rect 3892 9145 3893 9149
rect 4011 9148 4013 9153
rect 4087 9151 4089 9153
rect 4092 9148 4094 9153
rect 3822 9142 3824 9145
rect 3866 9142 3868 9145
rect 3892 9142 3894 9145
rect 3938 9142 3940 9145
rect 2877 9121 2879 9124
rect 2921 9121 2923 9124
rect 2947 9121 2949 9124
rect 2993 9121 2995 9124
rect 3061 9121 3063 9125
rect 3089 9127 3091 9129
rect 3140 9127 3142 9129
rect 3066 9121 3068 9124
rect 2947 9117 2948 9121
rect 2861 9114 2863 9116
rect 2877 9114 2879 9117
rect 2893 9114 2895 9116
rect 2916 9114 2918 9116
rect 2921 9114 2923 9117
rect 2947 9114 2949 9117
rect 2968 9114 2970 9117
rect 2988 9114 2990 9116
rect 2993 9114 2995 9117
rect 3011 9114 3013 9116
rect 3166 9121 3168 9125
rect 3194 9127 3196 9129
rect 3171 9121 3173 9124
rect 3061 9110 3063 9113
rect 3066 9111 3068 9113
rect 3062 9106 3063 9110
rect 2861 9092 2863 9106
rect 2877 9104 2879 9106
rect 2877 9092 2879 9094
rect 2893 9092 2895 9106
rect 2916 9101 2918 9106
rect 2921 9104 2923 9106
rect 2947 9104 2949 9106
rect 2912 9097 2918 9101
rect 2916 9092 2918 9097
rect 2921 9092 2923 9094
rect 2947 9092 2949 9094
rect 2968 9092 2970 9106
rect 2988 9101 2990 9106
rect 2993 9104 2995 9106
rect 2984 9097 2990 9101
rect 2988 9092 2990 9097
rect 2993 9092 2995 9094
rect 3011 9092 3013 9106
rect 3061 9101 3063 9106
rect 3066 9101 3068 9103
rect 3089 9097 3091 9119
rect 3140 9105 3142 9119
rect 3822 9121 3824 9124
rect 3866 9121 3868 9124
rect 3892 9121 3894 9124
rect 3938 9121 3940 9124
rect 4006 9121 4008 9125
rect 4034 9127 4036 9129
rect 4085 9127 4087 9129
rect 4011 9121 4013 9124
rect 3166 9110 3168 9113
rect 3171 9111 3173 9113
rect 3167 9106 3168 9110
rect 3166 9101 3168 9106
rect 3171 9101 3173 9103
rect 3140 9099 3142 9101
rect 3194 9097 3196 9119
rect 3892 9117 3893 9121
rect 3806 9114 3808 9116
rect 3822 9114 3824 9117
rect 3838 9114 3840 9116
rect 3861 9114 3863 9116
rect 3866 9114 3868 9117
rect 3892 9114 3894 9117
rect 3913 9114 3915 9117
rect 3933 9114 3935 9116
rect 3938 9114 3940 9117
rect 3956 9114 3958 9116
rect 4111 9121 4113 9125
rect 4139 9127 4141 9129
rect 4116 9121 4118 9124
rect 4006 9110 4008 9113
rect 4011 9111 4013 9113
rect 4007 9106 4008 9110
rect 3371 9098 3373 9100
rect 3061 9095 3063 9097
rect 3066 9092 3068 9097
rect 3166 9095 3168 9097
rect 3089 9091 3091 9093
rect 3171 9092 3173 9097
rect 3194 9091 3196 9093
rect 3397 9092 3399 9096
rect 3425 9098 3427 9100
rect 3402 9092 3404 9095
rect 2861 9086 2863 9088
rect 2877 9084 2879 9088
rect 2893 9086 2895 9088
rect 2916 9086 2918 9088
rect 2878 9080 2879 9084
rect 2921 9083 2923 9088
rect 2947 9084 2949 9088
rect 2968 9086 2970 9088
rect 2988 9086 2990 9088
rect 2877 9077 2879 9080
rect 2922 9079 2923 9083
rect 2948 9080 2949 9084
rect 2993 9083 2995 9088
rect 3011 9086 3013 9088
rect 2921 9077 2923 9079
rect 2947 9076 2949 9080
rect 2994 9079 2995 9083
rect 2993 9077 2995 9079
rect 3371 9076 3373 9090
rect 3557 9095 3559 9098
rect 3610 9095 3612 9098
rect 3397 9081 3399 9084
rect 3402 9082 3404 9084
rect 3398 9077 3399 9081
rect 3397 9072 3399 9077
rect 3402 9072 3404 9074
rect 3371 9070 3373 9072
rect 3425 9068 3427 9090
rect 3397 9066 3399 9068
rect 3402 9063 3404 9068
rect 3806 9092 3808 9106
rect 3822 9104 3824 9106
rect 3822 9092 3824 9094
rect 3838 9092 3840 9106
rect 3861 9101 3863 9106
rect 3866 9104 3868 9106
rect 3892 9104 3894 9106
rect 3857 9097 3863 9101
rect 3861 9092 3863 9097
rect 3866 9092 3868 9094
rect 3892 9092 3894 9094
rect 3913 9092 3915 9106
rect 3933 9101 3935 9106
rect 3938 9104 3940 9106
rect 3929 9097 3935 9101
rect 3933 9092 3935 9097
rect 3938 9092 3940 9094
rect 3956 9092 3958 9106
rect 4006 9101 4008 9106
rect 4011 9101 4013 9103
rect 4034 9097 4036 9119
rect 4085 9105 4087 9119
rect 4111 9110 4113 9113
rect 4116 9111 4118 9113
rect 4112 9106 4113 9110
rect 4111 9101 4113 9106
rect 4116 9101 4118 9103
rect 4085 9099 4087 9101
rect 4139 9097 4141 9119
rect 4006 9095 4008 9097
rect 4011 9092 4013 9097
rect 4111 9095 4113 9097
rect 4034 9091 4036 9093
rect 4116 9092 4118 9097
rect 4139 9091 4141 9093
rect 3806 9086 3808 9088
rect 3822 9084 3824 9088
rect 3838 9086 3840 9088
rect 3861 9086 3863 9088
rect 3823 9080 3824 9084
rect 3866 9083 3868 9088
rect 3892 9084 3894 9088
rect 3913 9086 3915 9088
rect 3933 9086 3935 9088
rect 3822 9077 3824 9080
rect 3867 9079 3868 9083
rect 3893 9080 3894 9084
rect 3938 9083 3940 9088
rect 3956 9086 3958 9088
rect 3866 9077 3868 9079
rect 3892 9076 3894 9080
rect 3939 9079 3940 9083
rect 3938 9077 3940 9079
rect 3425 9062 3427 9064
rect 2877 9054 2879 9057
rect 2921 9055 2923 9057
rect 2878 9050 2879 9054
rect 2922 9051 2923 9055
rect 2947 9054 2949 9058
rect 3557 9057 3559 9065
rect 3610 9057 3612 9065
rect 2993 9055 2995 9057
rect 2861 9046 2863 9048
rect 2877 9046 2879 9050
rect 2893 9046 2895 9048
rect 2916 9046 2918 9048
rect 2921 9046 2923 9051
rect 2948 9050 2949 9054
rect 2994 9051 2995 9055
rect 3822 9054 3824 9057
rect 3866 9055 3868 9057
rect 2947 9046 2949 9050
rect 2968 9046 2970 9048
rect 2988 9046 2990 9048
rect 2993 9046 2995 9051
rect 3011 9046 3013 9048
rect 3061 9046 3063 9049
rect 3066 9046 3068 9049
rect 3166 9046 3168 9049
rect 3171 9046 3173 9049
rect 3557 9045 3559 9053
rect 3610 9045 3612 9053
rect 3823 9050 3824 9054
rect 3867 9051 3868 9055
rect 3892 9054 3894 9058
rect 3938 9055 3940 9057
rect 3806 9046 3808 9048
rect 3822 9046 3824 9050
rect 3838 9046 3840 9048
rect 3861 9046 3863 9048
rect 3866 9046 3868 9051
rect 3893 9050 3894 9054
rect 3939 9051 3940 9055
rect 3892 9046 3894 9050
rect 3913 9046 3915 9048
rect 3933 9046 3935 9048
rect 3938 9046 3940 9051
rect 3956 9046 3958 9048
rect 4006 9046 4008 9049
rect 4011 9046 4013 9049
rect 4111 9046 4113 9049
rect 4116 9046 4118 9049
rect 2861 9028 2863 9042
rect 2877 9040 2879 9042
rect 2877 9028 2879 9030
rect 2893 9028 2895 9042
rect 2916 9037 2918 9042
rect 2921 9040 2923 9042
rect 2947 9040 2949 9042
rect 2912 9033 2918 9037
rect 2916 9028 2918 9033
rect 2921 9028 2923 9030
rect 2947 9028 2949 9030
rect 2968 9028 2970 9042
rect 2988 9037 2990 9042
rect 2993 9040 2995 9042
rect 2984 9033 2990 9037
rect 2988 9028 2990 9033
rect 2993 9028 2995 9030
rect 3011 9028 3013 9042
rect 3061 9030 3063 9042
rect 3066 9040 3068 9042
rect 3066 9030 3068 9032
rect 3166 9030 3168 9042
rect 3171 9040 3173 9042
rect 3171 9030 3173 9032
rect 3557 9031 3559 9033
rect 3610 9031 3612 9033
rect 3806 9028 3808 9042
rect 3822 9040 3824 9042
rect 3822 9028 3824 9030
rect 3838 9028 3840 9042
rect 3861 9037 3863 9042
rect 3866 9040 3868 9042
rect 3892 9040 3894 9042
rect 3857 9033 3863 9037
rect 3861 9028 3863 9033
rect 3866 9028 3868 9030
rect 3892 9028 3894 9030
rect 3913 9028 3915 9042
rect 3933 9037 3935 9042
rect 3938 9040 3940 9042
rect 3929 9033 3935 9037
rect 3933 9028 3935 9033
rect 3938 9028 3940 9030
rect 3956 9028 3958 9042
rect 4006 9030 4008 9042
rect 4011 9040 4013 9042
rect 4011 9030 4013 9032
rect 4111 9030 4113 9042
rect 4116 9040 4118 9042
rect 4116 9030 4118 9032
rect 3061 9020 3063 9022
rect 2861 9018 2863 9020
rect 2877 9017 2879 9020
rect 2893 9018 2895 9020
rect 2916 9018 2918 9020
rect 2921 9017 2923 9020
rect 2947 9017 2949 9020
rect 2968 9017 2970 9020
rect 2988 9018 2990 9020
rect 2993 9017 2995 9020
rect 3011 9018 3013 9020
rect 3066 9017 3068 9022
rect 3166 9020 3168 9022
rect 3171 9017 3173 9022
rect 4006 9020 4008 9022
rect 2947 9013 2948 9017
rect 3806 9018 3808 9020
rect 3822 9017 3824 9020
rect 3838 9018 3840 9020
rect 3861 9018 3863 9020
rect 3866 9017 3868 9020
rect 3892 9017 3894 9020
rect 3913 9017 3915 9020
rect 3933 9018 3935 9020
rect 3938 9017 3940 9020
rect 3956 9018 3958 9020
rect 4011 9017 4013 9022
rect 4111 9020 4113 9022
rect 4116 9017 4118 9022
rect 2877 9010 2879 9013
rect 2921 9010 2923 9013
rect 2947 9010 2949 9013
rect 2993 9010 2995 9013
rect 3397 9012 3399 9015
rect 3402 9012 3404 9015
rect 3892 9013 3893 9017
rect 3822 9010 3824 9013
rect 3866 9010 3868 9013
rect 3892 9010 3894 9013
rect 3938 9010 3940 9013
rect 2877 8989 2879 8992
rect 2921 8989 2923 8992
rect 2947 8989 2949 8992
rect 2993 8989 2995 8992
rect 3061 8989 3063 8993
rect 3089 8995 3091 8997
rect 3116 8995 3118 8997
rect 3066 8989 3068 8992
rect 2947 8985 2948 8989
rect 2861 8982 2863 8984
rect 2877 8982 2879 8985
rect 2893 8982 2895 8984
rect 2916 8982 2918 8984
rect 2921 8982 2923 8985
rect 2947 8982 2949 8985
rect 2968 8982 2970 8985
rect 2988 8982 2990 8984
rect 2993 8982 2995 8985
rect 3011 8982 3013 8984
rect 3142 8989 3144 8993
rect 3170 8995 3172 8997
rect 3206 8995 3208 8997
rect 3147 8989 3149 8992
rect 3061 8978 3063 8981
rect 3066 8979 3068 8981
rect 3062 8974 3063 8978
rect 2861 8960 2863 8974
rect 2877 8972 2879 8974
rect 2877 8960 2879 8962
rect 2893 8960 2895 8974
rect 2916 8969 2918 8974
rect 2921 8972 2923 8974
rect 2947 8972 2949 8974
rect 2912 8965 2918 8969
rect 2916 8960 2918 8965
rect 2921 8960 2923 8962
rect 2947 8960 2949 8962
rect 2968 8960 2970 8974
rect 2988 8969 2990 8974
rect 2993 8972 2995 8974
rect 2984 8965 2990 8969
rect 2988 8960 2990 8965
rect 2993 8960 2995 8962
rect 3011 8960 3013 8974
rect 3061 8969 3063 8974
rect 3066 8969 3068 8971
rect 3089 8965 3091 8987
rect 3116 8973 3118 8987
rect 3232 8989 3234 8993
rect 3260 8995 3262 8997
rect 3397 8996 3399 9008
rect 3402 9006 3404 9008
rect 3402 8996 3404 8998
rect 3237 8989 3239 8992
rect 3142 8978 3144 8981
rect 3147 8979 3149 8981
rect 3143 8974 3144 8978
rect 3142 8969 3144 8974
rect 3147 8969 3149 8971
rect 3116 8967 3118 8969
rect 3170 8965 3172 8987
rect 3206 8973 3208 8987
rect 3822 8989 3824 8992
rect 3866 8989 3868 8992
rect 3892 8989 3894 8992
rect 3938 8989 3940 8992
rect 4006 8989 4008 8993
rect 4034 8995 4036 8997
rect 4061 8995 4063 8997
rect 4011 8989 4013 8992
rect 3232 8978 3234 8981
rect 3237 8979 3239 8981
rect 3233 8974 3234 8978
rect 3232 8969 3234 8974
rect 3237 8969 3239 8971
rect 3206 8967 3208 8969
rect 3260 8965 3262 8987
rect 3397 8986 3399 8988
rect 3402 8983 3404 8988
rect 3892 8985 3893 8989
rect 3806 8982 3808 8984
rect 3822 8982 3824 8985
rect 3838 8982 3840 8984
rect 3861 8982 3863 8984
rect 3866 8982 3868 8985
rect 3892 8982 3894 8985
rect 3913 8982 3915 8985
rect 3933 8982 3935 8984
rect 3938 8982 3940 8985
rect 3956 8982 3958 8984
rect 4087 8989 4089 8993
rect 4115 8995 4117 8997
rect 4151 8995 4153 8997
rect 4092 8989 4094 8992
rect 4006 8978 4008 8981
rect 4011 8979 4013 8981
rect 4007 8974 4008 8978
rect 3349 8968 3351 8970
rect 3371 8968 3373 8970
rect 3061 8963 3063 8965
rect 3066 8960 3068 8965
rect 3142 8963 3144 8965
rect 3089 8959 3091 8961
rect 3147 8960 3149 8965
rect 3232 8963 3234 8965
rect 3170 8959 3172 8961
rect 3237 8960 3239 8965
rect 3260 8959 3262 8961
rect 3397 8962 3399 8966
rect 3425 8968 3427 8970
rect 3402 8962 3404 8965
rect 2861 8954 2863 8956
rect 2877 8952 2879 8956
rect 2893 8954 2895 8956
rect 2916 8954 2918 8956
rect 2878 8948 2879 8952
rect 2921 8951 2923 8956
rect 2947 8952 2949 8956
rect 2968 8954 2970 8956
rect 2988 8954 2990 8956
rect 2877 8945 2879 8948
rect 2922 8947 2923 8951
rect 2948 8948 2949 8952
rect 2993 8951 2995 8956
rect 3011 8954 3013 8956
rect 2921 8945 2923 8947
rect 2947 8944 2949 8948
rect 2994 8947 2995 8951
rect 2993 8945 2995 8947
rect 3349 8946 3351 8960
rect 3371 8946 3373 8960
rect 3463 8965 3465 8968
rect 3516 8965 3518 8968
rect 3397 8951 3399 8954
rect 3402 8952 3404 8954
rect 3398 8947 3399 8951
rect 3397 8942 3399 8947
rect 3402 8942 3404 8944
rect 3349 8940 3351 8942
rect 3371 8940 3373 8942
rect 3425 8938 3427 8960
rect 3397 8936 3399 8938
rect 3402 8933 3404 8938
rect 3806 8960 3808 8974
rect 3822 8972 3824 8974
rect 3822 8960 3824 8962
rect 3838 8960 3840 8974
rect 3861 8969 3863 8974
rect 3866 8972 3868 8974
rect 3892 8972 3894 8974
rect 3857 8965 3863 8969
rect 3861 8960 3863 8965
rect 3866 8960 3868 8962
rect 3892 8960 3894 8962
rect 3913 8960 3915 8974
rect 3933 8969 3935 8974
rect 3938 8972 3940 8974
rect 3929 8965 3935 8969
rect 3933 8960 3935 8965
rect 3938 8960 3940 8962
rect 3956 8960 3958 8974
rect 4006 8969 4008 8974
rect 4011 8969 4013 8971
rect 4034 8965 4036 8987
rect 4061 8973 4063 8987
rect 4177 8989 4179 8993
rect 4205 8995 4207 8997
rect 4182 8989 4184 8992
rect 4087 8978 4089 8981
rect 4092 8979 4094 8981
rect 4088 8974 4089 8978
rect 4087 8969 4089 8974
rect 4092 8969 4094 8971
rect 4061 8967 4063 8969
rect 4115 8965 4117 8987
rect 4151 8973 4153 8987
rect 4177 8978 4179 8981
rect 4182 8979 4184 8981
rect 4178 8974 4179 8978
rect 4177 8969 4179 8974
rect 4182 8969 4184 8971
rect 4151 8967 4153 8969
rect 4205 8965 4207 8987
rect 4006 8963 4008 8965
rect 4011 8960 4013 8965
rect 4087 8963 4089 8965
rect 4034 8959 4036 8961
rect 4092 8960 4094 8965
rect 4177 8963 4179 8965
rect 4115 8959 4117 8961
rect 4182 8960 4184 8965
rect 4205 8959 4207 8961
rect 3806 8954 3808 8956
rect 3822 8952 3824 8956
rect 3838 8954 3840 8956
rect 3861 8954 3863 8956
rect 3823 8948 3824 8952
rect 3866 8951 3868 8956
rect 3892 8952 3894 8956
rect 3913 8954 3915 8956
rect 3933 8954 3935 8956
rect 3822 8945 3824 8948
rect 3867 8947 3868 8951
rect 3893 8948 3894 8952
rect 3938 8951 3940 8956
rect 3956 8954 3958 8956
rect 3866 8945 3868 8947
rect 3892 8944 3894 8948
rect 3939 8947 3940 8951
rect 3938 8945 3940 8947
rect 3425 8932 3427 8934
rect 3463 8927 3465 8935
rect 3516 8927 3518 8935
rect 2877 8922 2879 8925
rect 2921 8923 2923 8925
rect 2878 8918 2879 8922
rect 2922 8919 2923 8923
rect 2947 8922 2949 8926
rect 2993 8923 2995 8925
rect 2861 8914 2863 8916
rect 2877 8914 2879 8918
rect 2893 8914 2895 8916
rect 2916 8914 2918 8916
rect 2921 8914 2923 8919
rect 2948 8918 2949 8922
rect 2994 8919 2995 8923
rect 2947 8914 2949 8918
rect 2968 8914 2970 8916
rect 2988 8914 2990 8916
rect 2993 8914 2995 8919
rect 3011 8914 3013 8916
rect 3463 8915 3465 8923
rect 3516 8915 3518 8923
rect 3822 8922 3824 8925
rect 3866 8923 3868 8925
rect 3823 8918 3824 8922
rect 3867 8919 3868 8923
rect 3892 8922 3894 8926
rect 3938 8923 3940 8925
rect 3061 8911 3063 8914
rect 3066 8911 3068 8914
rect 3142 8911 3144 8914
rect 3147 8911 3149 8914
rect 3232 8911 3234 8914
rect 3237 8911 3239 8914
rect 2861 8896 2863 8910
rect 2877 8908 2879 8910
rect 2877 8896 2879 8898
rect 2893 8896 2895 8910
rect 2916 8905 2918 8910
rect 2921 8908 2923 8910
rect 2947 8908 2949 8910
rect 2912 8901 2918 8905
rect 2916 8896 2918 8901
rect 2921 8896 2923 8898
rect 2947 8896 2949 8898
rect 2968 8896 2970 8910
rect 2988 8905 2990 8910
rect 2993 8908 2995 8910
rect 2984 8901 2990 8905
rect 2988 8896 2990 8901
rect 2993 8896 2995 8898
rect 3011 8896 3013 8910
rect 3061 8895 3063 8907
rect 3066 8905 3068 8907
rect 3066 8895 3068 8897
rect 3142 8895 3144 8907
rect 3147 8905 3149 8907
rect 3147 8895 3149 8897
rect 3232 8895 3234 8907
rect 3237 8905 3239 8907
rect 3806 8914 3808 8916
rect 3822 8914 3824 8918
rect 3838 8914 3840 8916
rect 3861 8914 3863 8916
rect 3866 8914 3868 8919
rect 3893 8918 3894 8922
rect 3939 8919 3940 8923
rect 3892 8914 3894 8918
rect 3913 8914 3915 8916
rect 3933 8914 3935 8916
rect 3938 8914 3940 8919
rect 3956 8914 3958 8916
rect 4006 8911 4008 8914
rect 4011 8911 4013 8914
rect 4087 8911 4089 8914
rect 4092 8911 4094 8914
rect 4177 8911 4179 8914
rect 4182 8911 4184 8914
rect 3463 8901 3465 8903
rect 3516 8901 3518 8903
rect 3237 8895 3239 8897
rect 3806 8896 3808 8910
rect 3822 8908 3824 8910
rect 3822 8896 3824 8898
rect 3838 8896 3840 8910
rect 3861 8905 3863 8910
rect 3866 8908 3868 8910
rect 3892 8908 3894 8910
rect 3857 8901 3863 8905
rect 3861 8896 3863 8901
rect 3866 8896 3868 8898
rect 3892 8896 3894 8898
rect 3913 8896 3915 8910
rect 3933 8905 3935 8910
rect 3938 8908 3940 8910
rect 3929 8901 3935 8905
rect 3933 8896 3935 8901
rect 3938 8896 3940 8898
rect 3956 8896 3958 8910
rect 2861 8886 2863 8888
rect 2877 8885 2879 8888
rect 2893 8886 2895 8888
rect 2916 8886 2918 8888
rect 2921 8885 2923 8888
rect 2947 8885 2949 8888
rect 2968 8885 2970 8888
rect 2988 8886 2990 8888
rect 2993 8885 2995 8888
rect 3011 8886 3013 8888
rect 3061 8885 3063 8887
rect 2947 8881 2948 8885
rect 3066 8882 3068 8887
rect 3142 8885 3144 8887
rect 3147 8882 3149 8887
rect 3232 8885 3234 8887
rect 3237 8882 3239 8887
rect 4006 8895 4008 8907
rect 4011 8905 4013 8907
rect 4011 8895 4013 8897
rect 4087 8895 4089 8907
rect 4092 8905 4094 8907
rect 4092 8895 4094 8897
rect 4177 8895 4179 8907
rect 4182 8905 4184 8907
rect 4182 8895 4184 8897
rect 3806 8886 3808 8888
rect 3822 8885 3824 8888
rect 3838 8886 3840 8888
rect 3861 8886 3863 8888
rect 3866 8885 3868 8888
rect 3892 8885 3894 8888
rect 3913 8885 3915 8888
rect 3933 8886 3935 8888
rect 3938 8885 3940 8888
rect 3956 8886 3958 8888
rect 4006 8885 4008 8887
rect 3397 8882 3399 8885
rect 3402 8882 3404 8885
rect 2877 8878 2879 8881
rect 2921 8878 2923 8881
rect 2947 8878 2949 8881
rect 2993 8878 2995 8881
rect 3892 8881 3893 8885
rect 4011 8882 4013 8887
rect 4087 8885 4089 8887
rect 4092 8882 4094 8887
rect 4177 8885 4179 8887
rect 4182 8882 4184 8887
rect 3822 8878 3824 8881
rect 3866 8878 3868 8881
rect 3892 8878 3894 8881
rect 3938 8878 3940 8881
rect 3397 8866 3399 8878
rect 3402 8876 3404 8878
rect 3402 8866 3404 8868
rect 2877 8857 2879 8860
rect 2921 8857 2923 8860
rect 2947 8857 2949 8860
rect 2993 8857 2995 8860
rect 3061 8857 3063 8861
rect 3089 8863 3091 8865
rect 3066 8857 3068 8860
rect 2947 8853 2948 8857
rect 2861 8850 2863 8852
rect 2877 8850 2879 8853
rect 2893 8850 2895 8852
rect 2916 8850 2918 8852
rect 2921 8850 2923 8853
rect 2947 8850 2949 8853
rect 2968 8850 2970 8853
rect 2988 8850 2990 8852
rect 2993 8850 2995 8853
rect 3011 8850 3013 8852
rect 3397 8856 3399 8858
rect 3061 8846 3063 8849
rect 3066 8847 3068 8849
rect 3062 8842 3063 8846
rect 2861 8828 2863 8842
rect 2877 8840 2879 8842
rect 2877 8828 2879 8830
rect 2893 8828 2895 8842
rect 2916 8837 2918 8842
rect 2921 8840 2923 8842
rect 2947 8840 2949 8842
rect 2912 8833 2918 8837
rect 2916 8828 2918 8833
rect 2921 8828 2923 8830
rect 2947 8828 2949 8830
rect 2968 8828 2970 8842
rect 2988 8837 2990 8842
rect 2993 8840 2995 8842
rect 2984 8833 2990 8837
rect 2988 8828 2990 8833
rect 2993 8828 2995 8830
rect 3011 8828 3013 8842
rect 3061 8837 3063 8842
rect 3066 8837 3068 8839
rect 3089 8833 3091 8855
rect 3402 8853 3404 8858
rect 3822 8857 3824 8860
rect 3866 8857 3868 8860
rect 3892 8857 3894 8860
rect 3938 8857 3940 8860
rect 4006 8857 4008 8861
rect 4034 8863 4036 8865
rect 4011 8857 4013 8860
rect 3892 8853 3893 8857
rect 3806 8850 3808 8852
rect 3822 8850 3824 8853
rect 3838 8850 3840 8852
rect 3861 8850 3863 8852
rect 3866 8850 3868 8853
rect 3892 8850 3894 8853
rect 3913 8850 3915 8853
rect 3933 8850 3935 8852
rect 3938 8850 3940 8853
rect 3956 8850 3958 8852
rect 4006 8846 4008 8849
rect 4011 8847 4013 8849
rect 4007 8842 4008 8846
rect 3061 8831 3063 8833
rect 3066 8828 3068 8833
rect 3089 8827 3091 8829
rect 3806 8828 3808 8842
rect 3822 8840 3824 8842
rect 3822 8828 3824 8830
rect 3838 8828 3840 8842
rect 3861 8837 3863 8842
rect 3866 8840 3868 8842
rect 3892 8840 3894 8842
rect 3857 8833 3863 8837
rect 3861 8828 3863 8833
rect 3866 8828 3868 8830
rect 3892 8828 3894 8830
rect 3913 8828 3915 8842
rect 3933 8837 3935 8842
rect 3938 8840 3940 8842
rect 3929 8833 3935 8837
rect 3933 8828 3935 8833
rect 3938 8828 3940 8830
rect 3956 8828 3958 8842
rect 4006 8837 4008 8842
rect 4011 8837 4013 8839
rect 4034 8833 4036 8855
rect 4006 8831 4008 8833
rect 4011 8828 4013 8833
rect 4034 8827 4036 8829
rect 2861 8822 2863 8824
rect 2877 8820 2879 8824
rect 2893 8822 2895 8824
rect 2916 8822 2918 8824
rect 2878 8816 2879 8820
rect 2921 8819 2923 8824
rect 2947 8820 2949 8824
rect 2968 8822 2970 8824
rect 2988 8822 2990 8824
rect 2877 8813 2879 8816
rect 2922 8815 2923 8819
rect 2948 8816 2949 8820
rect 2993 8819 2995 8824
rect 3011 8822 3013 8824
rect 3806 8822 3808 8824
rect 3822 8820 3824 8824
rect 3838 8822 3840 8824
rect 3861 8822 3863 8824
rect 2921 8813 2923 8815
rect 2947 8812 2949 8816
rect 2994 8815 2995 8819
rect 3823 8816 3824 8820
rect 3866 8819 3868 8824
rect 3892 8820 3894 8824
rect 3913 8822 3915 8824
rect 3933 8822 3935 8824
rect 2993 8813 2995 8815
rect 3822 8813 3824 8816
rect 3867 8815 3868 8819
rect 3893 8816 3894 8820
rect 3938 8819 3940 8824
rect 3956 8822 3958 8824
rect 3866 8813 3868 8815
rect 3892 8812 3894 8816
rect 3939 8815 3940 8819
rect 3938 8813 3940 8815
rect 2372 8795 2374 8797
rect 2377 8795 2379 8798
rect 2393 8795 2395 8797
rect 2409 8795 2411 8797
rect 2414 8795 2416 8798
rect 2435 8795 2437 8798
rect 2451 8795 2453 8798
rect 2467 8795 2469 8797
rect 2472 8795 2474 8798
rect 2488 8795 2490 8797
rect 2504 8795 2506 8797
rect 2509 8795 2511 8798
rect 2525 8795 2527 8797
rect 2541 8795 2543 8797
rect 2546 8795 2548 8798
rect 2567 8795 2569 8798
rect 2583 8795 2585 8798
rect 2599 8795 2601 8797
rect 2604 8795 2606 8798
rect 2620 8795 2622 8797
rect 2636 8795 2638 8797
rect 2641 8795 2643 8798
rect 2657 8795 2659 8797
rect 2673 8795 2675 8797
rect 2678 8795 2680 8798
rect 2699 8795 2701 8798
rect 2715 8795 2717 8798
rect 2731 8795 2733 8797
rect 2736 8795 2738 8798
rect 2752 8795 2754 8797
rect 3317 8795 3319 8797
rect 3322 8795 3324 8798
rect 3338 8795 3340 8797
rect 3354 8795 3356 8797
rect 3359 8795 3361 8798
rect 3380 8795 3382 8798
rect 3396 8795 3398 8798
rect 3412 8795 3414 8797
rect 3417 8795 3419 8798
rect 3433 8795 3435 8797
rect 3449 8795 3451 8797
rect 3454 8795 3456 8798
rect 3470 8795 3472 8797
rect 3486 8795 3488 8797
rect 3491 8795 3493 8798
rect 3512 8795 3514 8798
rect 3528 8795 3530 8798
rect 3544 8795 3546 8797
rect 3549 8795 3551 8798
rect 3565 8795 3567 8797
rect 3581 8795 3583 8797
rect 3586 8795 3588 8798
rect 3602 8795 3604 8797
rect 3618 8795 3620 8797
rect 3623 8795 3625 8798
rect 3644 8795 3646 8798
rect 3660 8795 3662 8798
rect 3676 8795 3678 8797
rect 3681 8795 3683 8798
rect 3697 8795 3699 8797
rect 2877 8790 2879 8793
rect 2921 8791 2923 8793
rect 2372 8782 2374 8787
rect 2377 8785 2379 8787
rect 2372 8768 2374 8778
rect 2377 8768 2379 8775
rect 2393 8768 2395 8787
rect 2409 8778 2411 8787
rect 2414 8785 2416 8787
rect 2435 8785 2437 8787
rect 2451 8784 2453 8787
rect 2409 8768 2411 8771
rect 2414 8768 2416 8770
rect 2435 8768 2437 8770
rect 2451 8768 2453 8780
rect 2467 8778 2469 8787
rect 2472 8785 2474 8787
rect 2467 8768 2469 8771
rect 2472 8768 2474 8770
rect 2488 8768 2490 8787
rect 2504 8784 2506 8787
rect 2509 8785 2511 8787
rect 2504 8768 2506 8780
rect 2509 8768 2511 8775
rect 2525 8768 2527 8787
rect 2541 8778 2543 8787
rect 2546 8785 2548 8787
rect 2567 8785 2569 8787
rect 2583 8784 2585 8787
rect 2541 8768 2543 8771
rect 2546 8768 2548 8770
rect 2567 8768 2569 8770
rect 2583 8768 2585 8780
rect 2599 8778 2601 8787
rect 2604 8785 2606 8787
rect 2599 8768 2601 8771
rect 2604 8768 2606 8770
rect 2620 8768 2622 8787
rect 2636 8784 2638 8787
rect 2641 8785 2643 8787
rect 2636 8768 2638 8780
rect 2641 8768 2643 8775
rect 2657 8768 2659 8787
rect 2673 8778 2675 8787
rect 2678 8785 2680 8787
rect 2699 8785 2701 8787
rect 2715 8784 2717 8787
rect 2673 8768 2675 8771
rect 2678 8768 2680 8770
rect 2699 8768 2701 8770
rect 2715 8768 2717 8780
rect 2731 8778 2733 8787
rect 2736 8785 2738 8787
rect 2752 8779 2754 8787
rect 2878 8786 2879 8790
rect 2922 8787 2923 8791
rect 2947 8790 2949 8794
rect 2993 8791 2995 8793
rect 2861 8782 2863 8784
rect 2877 8782 2879 8786
rect 2893 8782 2895 8784
rect 2916 8782 2918 8784
rect 2921 8782 2923 8787
rect 2948 8786 2949 8790
rect 2994 8787 2995 8791
rect 3138 8790 3140 8793
rect 3182 8791 3184 8793
rect 2947 8782 2949 8786
rect 2968 8782 2970 8784
rect 2988 8782 2990 8784
rect 2993 8782 2995 8787
rect 3139 8786 3140 8790
rect 3183 8787 3184 8791
rect 3208 8790 3210 8794
rect 3254 8791 3256 8793
rect 3011 8782 3013 8784
rect 3095 8782 3097 8785
rect 3113 8782 3115 8785
rect 3138 8782 3140 8786
rect 3154 8782 3156 8784
rect 3177 8782 3179 8784
rect 3182 8782 3184 8787
rect 3209 8786 3210 8790
rect 3255 8787 3256 8791
rect 3822 8790 3824 8793
rect 3866 8791 3868 8793
rect 3208 8782 3210 8786
rect 3229 8782 3231 8784
rect 3249 8782 3251 8784
rect 3254 8782 3256 8787
rect 3272 8782 3274 8784
rect 3317 8782 3319 8787
rect 3322 8785 3324 8787
rect 2731 8768 2733 8771
rect 2736 8768 2738 8770
rect 2752 8768 2754 8775
rect 2861 8764 2863 8778
rect 2877 8776 2879 8778
rect 2877 8764 2879 8766
rect 2893 8764 2895 8778
rect 2916 8773 2918 8778
rect 2921 8776 2923 8778
rect 2947 8776 2949 8778
rect 2912 8769 2918 8773
rect 2916 8764 2918 8769
rect 2921 8764 2923 8766
rect 2947 8764 2949 8766
rect 2968 8764 2970 8778
rect 2988 8773 2990 8778
rect 2993 8776 2995 8778
rect 2984 8769 2990 8773
rect 2988 8764 2990 8769
rect 2993 8764 2995 8766
rect 3011 8764 3013 8778
rect 3061 8775 3063 8778
rect 3066 8775 3068 8778
rect 3095 8773 3097 8778
rect 2372 8762 2374 8764
rect 2377 8761 2379 8764
rect 2393 8762 2395 8764
rect 2409 8762 2411 8764
rect 2414 8759 2416 8764
rect 2435 8759 2437 8764
rect 2451 8762 2453 8764
rect 2467 8762 2469 8764
rect 2472 8759 2474 8764
rect 2488 8762 2490 8764
rect 2504 8762 2506 8764
rect 2509 8761 2511 8764
rect 2525 8762 2527 8764
rect 2541 8762 2543 8764
rect 2546 8759 2548 8764
rect 2567 8759 2569 8764
rect 2583 8762 2585 8764
rect 2599 8762 2601 8764
rect 2604 8759 2606 8764
rect 2620 8762 2622 8764
rect 2636 8762 2638 8764
rect 2641 8761 2643 8764
rect 2657 8762 2659 8764
rect 2673 8762 2675 8764
rect 2678 8759 2680 8764
rect 2699 8759 2701 8764
rect 2715 8762 2717 8764
rect 2731 8762 2733 8764
rect 2736 8759 2738 8764
rect 2752 8762 2754 8764
rect 3061 8759 3063 8771
rect 3066 8769 3068 8771
rect 3095 8764 3097 8769
rect 3113 8764 3115 8778
rect 3138 8776 3140 8778
rect 3138 8764 3140 8766
rect 3154 8764 3156 8778
rect 3177 8773 3179 8778
rect 3182 8776 3184 8778
rect 3208 8776 3210 8778
rect 3173 8769 3179 8773
rect 3177 8764 3179 8769
rect 3182 8764 3184 8766
rect 3208 8764 3210 8766
rect 3229 8764 3231 8778
rect 3249 8773 3251 8778
rect 3254 8776 3256 8778
rect 3245 8769 3251 8773
rect 3249 8764 3251 8769
rect 3254 8764 3256 8766
rect 3272 8764 3274 8778
rect 3317 8768 3319 8778
rect 3322 8768 3324 8775
rect 3338 8768 3340 8787
rect 3354 8778 3356 8787
rect 3359 8785 3361 8787
rect 3380 8785 3382 8787
rect 3396 8784 3398 8787
rect 3354 8768 3356 8771
rect 3359 8768 3361 8770
rect 3380 8768 3382 8770
rect 3396 8768 3398 8780
rect 3412 8778 3414 8787
rect 3417 8785 3419 8787
rect 3412 8768 3414 8771
rect 3417 8768 3419 8770
rect 3433 8768 3435 8787
rect 3449 8784 3451 8787
rect 3454 8785 3456 8787
rect 3449 8768 3451 8780
rect 3454 8768 3456 8775
rect 3470 8768 3472 8787
rect 3486 8778 3488 8787
rect 3491 8785 3493 8787
rect 3512 8785 3514 8787
rect 3528 8784 3530 8787
rect 3486 8768 3488 8771
rect 3491 8768 3493 8770
rect 3512 8768 3514 8770
rect 3528 8768 3530 8780
rect 3544 8778 3546 8787
rect 3549 8785 3551 8787
rect 3544 8768 3546 8771
rect 3549 8768 3551 8770
rect 3565 8768 3567 8787
rect 3581 8784 3583 8787
rect 3586 8785 3588 8787
rect 3581 8768 3583 8780
rect 3586 8768 3588 8775
rect 3602 8768 3604 8787
rect 3618 8778 3620 8787
rect 3623 8785 3625 8787
rect 3644 8785 3646 8787
rect 3660 8784 3662 8787
rect 3618 8768 3620 8771
rect 3623 8768 3625 8770
rect 3644 8768 3646 8770
rect 3660 8768 3662 8780
rect 3676 8778 3678 8787
rect 3681 8785 3683 8787
rect 3697 8779 3699 8787
rect 3823 8786 3824 8790
rect 3867 8787 3868 8791
rect 3892 8790 3894 8794
rect 3938 8791 3940 8793
rect 3806 8782 3808 8784
rect 3822 8782 3824 8786
rect 3838 8782 3840 8784
rect 3861 8782 3863 8784
rect 3866 8782 3868 8787
rect 3893 8786 3894 8790
rect 3939 8787 3940 8791
rect 4083 8790 4085 8793
rect 4127 8791 4129 8793
rect 3892 8782 3894 8786
rect 3913 8782 3915 8784
rect 3933 8782 3935 8784
rect 3938 8782 3940 8787
rect 4084 8786 4085 8790
rect 4128 8787 4129 8791
rect 4153 8790 4155 8794
rect 4199 8791 4201 8793
rect 3956 8782 3958 8784
rect 4040 8782 4042 8785
rect 4058 8782 4060 8785
rect 4083 8782 4085 8786
rect 4099 8782 4101 8784
rect 4122 8782 4124 8784
rect 4127 8782 4129 8787
rect 4154 8786 4155 8790
rect 4200 8787 4201 8791
rect 4153 8782 4155 8786
rect 4174 8782 4176 8784
rect 4194 8782 4196 8784
rect 4199 8782 4201 8787
rect 4217 8782 4219 8784
rect 3676 8768 3678 8771
rect 3681 8768 3683 8770
rect 3697 8768 3699 8775
rect 3806 8764 3808 8778
rect 3822 8776 3824 8778
rect 3822 8764 3824 8766
rect 3838 8764 3840 8778
rect 3861 8773 3863 8778
rect 3866 8776 3868 8778
rect 3892 8776 3894 8778
rect 3857 8769 3863 8773
rect 3861 8764 3863 8769
rect 3866 8764 3868 8766
rect 3892 8764 3894 8766
rect 3913 8764 3915 8778
rect 3933 8773 3935 8778
rect 3938 8776 3940 8778
rect 3929 8769 3935 8773
rect 3933 8764 3935 8769
rect 3938 8764 3940 8766
rect 3956 8764 3958 8778
rect 4006 8775 4008 8778
rect 4011 8775 4013 8778
rect 4040 8773 4042 8778
rect 3066 8759 3068 8761
rect 2861 8754 2863 8756
rect 2877 8753 2879 8756
rect 2893 8754 2895 8756
rect 2916 8754 2918 8756
rect 2921 8753 2923 8756
rect 2947 8753 2949 8756
rect 2968 8753 2970 8756
rect 2988 8754 2990 8756
rect 2993 8753 2995 8756
rect 3011 8754 3013 8756
rect 2947 8749 2948 8753
rect 3317 8762 3319 8764
rect 3322 8761 3324 8764
rect 3338 8762 3340 8764
rect 3354 8762 3356 8764
rect 3359 8759 3361 8764
rect 3380 8759 3382 8764
rect 3396 8762 3398 8764
rect 3412 8762 3414 8764
rect 3417 8759 3419 8764
rect 3433 8762 3435 8764
rect 3449 8762 3451 8764
rect 3095 8753 3097 8756
rect 3061 8749 3063 8751
rect 2877 8746 2879 8749
rect 2921 8746 2923 8749
rect 2947 8746 2949 8749
rect 2993 8746 2995 8749
rect 3066 8746 3068 8751
rect 2487 8724 2489 8727
rect 2511 8724 2513 8727
rect 2487 8717 2489 8720
rect 2511 8717 2513 8720
rect 3113 8714 3115 8756
rect 3138 8753 3140 8756
rect 3154 8754 3156 8756
rect 3177 8754 3179 8756
rect 3182 8753 3184 8756
rect 3208 8753 3210 8756
rect 3229 8753 3231 8756
rect 3249 8754 3251 8756
rect 3254 8753 3256 8756
rect 3272 8754 3274 8756
rect 3454 8761 3456 8764
rect 3470 8762 3472 8764
rect 3486 8762 3488 8764
rect 3491 8759 3493 8764
rect 3512 8759 3514 8764
rect 3528 8762 3530 8764
rect 3544 8762 3546 8764
rect 3549 8759 3551 8764
rect 3565 8762 3567 8764
rect 3581 8762 3583 8764
rect 3586 8761 3588 8764
rect 3602 8762 3604 8764
rect 3618 8762 3620 8764
rect 3623 8759 3625 8764
rect 3644 8759 3646 8764
rect 3660 8762 3662 8764
rect 3676 8762 3678 8764
rect 3681 8759 3683 8764
rect 3697 8762 3699 8764
rect 4006 8759 4008 8771
rect 4011 8769 4013 8771
rect 4040 8764 4042 8769
rect 4058 8764 4060 8778
rect 4083 8776 4085 8778
rect 4083 8764 4085 8766
rect 4099 8764 4101 8778
rect 4122 8773 4124 8778
rect 4127 8776 4129 8778
rect 4153 8776 4155 8778
rect 4118 8769 4124 8773
rect 4122 8764 4124 8769
rect 4127 8764 4129 8766
rect 4153 8764 4155 8766
rect 4174 8764 4176 8778
rect 4194 8773 4196 8778
rect 4199 8776 4201 8778
rect 4190 8769 4196 8773
rect 4194 8764 4196 8769
rect 4199 8764 4201 8766
rect 4217 8764 4219 8778
rect 4011 8759 4013 8761
rect 3806 8754 3808 8756
rect 3822 8753 3824 8756
rect 3838 8754 3840 8756
rect 3861 8754 3863 8756
rect 3866 8753 3868 8756
rect 3892 8753 3894 8756
rect 3913 8753 3915 8756
rect 3933 8754 3935 8756
rect 3938 8753 3940 8756
rect 3956 8754 3958 8756
rect 3208 8749 3209 8753
rect 3138 8746 3140 8749
rect 3182 8746 3184 8749
rect 3208 8746 3210 8749
rect 3254 8746 3256 8749
rect 3892 8749 3893 8753
rect 4040 8753 4042 8756
rect 4006 8749 4008 8751
rect 3822 8746 3824 8749
rect 3866 8746 3868 8749
rect 3892 8746 3894 8749
rect 3938 8746 3940 8749
rect 4011 8746 4013 8751
rect 3432 8724 3434 8727
rect 3456 8724 3458 8727
rect 3281 8722 3284 8724
rect 3288 8722 3291 8724
rect 3432 8717 3434 8720
rect 3456 8717 3458 8720
rect 4058 8718 4060 8756
rect 4083 8753 4085 8756
rect 4099 8754 4101 8756
rect 4122 8754 4124 8756
rect 4127 8753 4129 8756
rect 4153 8753 4155 8756
rect 4174 8753 4176 8756
rect 4194 8754 4196 8756
rect 4199 8753 4201 8756
rect 4217 8754 4219 8756
rect 4153 8749 4154 8753
rect 4083 8746 4085 8749
rect 4127 8746 4129 8749
rect 4153 8746 4155 8749
rect 4199 8746 4201 8749
rect 4226 8722 4229 8724
rect 4233 8722 4236 8724
rect 2507 8711 2509 8713
rect 3452 8711 3454 8713
rect 2507 8704 2509 8707
rect 3452 8704 3454 8707
rect 2496 8693 2498 8695
rect 2502 8693 2521 8695
rect 3441 8693 3443 8695
rect 3447 8693 3466 8695
rect 2487 8688 2489 8690
rect 2511 8688 2513 8690
rect 3432 8688 3434 8690
rect 3456 8688 3458 8690
rect 2487 8681 2489 8684
rect 2511 8681 2513 8684
rect 3155 8683 3157 8685
rect 3160 8683 3162 8686
rect 3176 8683 3178 8685
rect 3192 8683 3194 8685
rect 3197 8683 3199 8686
rect 3218 8683 3220 8686
rect 3234 8683 3236 8686
rect 3250 8683 3252 8685
rect 3255 8683 3257 8686
rect 3271 8683 3273 8685
rect 3432 8681 3434 8684
rect 3456 8681 3458 8684
rect 4100 8683 4102 8685
rect 4105 8683 4107 8686
rect 4121 8683 4123 8685
rect 4137 8683 4139 8685
rect 4142 8683 4144 8686
rect 4163 8683 4165 8686
rect 4179 8683 4181 8686
rect 4195 8683 4197 8685
rect 4200 8683 4202 8686
rect 4216 8683 4218 8685
rect 3155 8670 3157 8675
rect 3160 8673 3162 8675
rect 3155 8656 3157 8666
rect 3160 8656 3162 8663
rect 3176 8656 3178 8675
rect 3192 8666 3194 8675
rect 3197 8673 3199 8675
rect 3218 8673 3220 8675
rect 3234 8672 3236 8675
rect 3192 8656 3194 8659
rect 3197 8656 3199 8658
rect 3218 8656 3220 8658
rect 3234 8656 3236 8668
rect 3250 8666 3252 8675
rect 3255 8673 3257 8675
rect 3250 8656 3252 8659
rect 3255 8656 3257 8658
rect 3271 8656 3273 8675
rect 4100 8670 4102 8675
rect 4105 8673 4107 8675
rect 4100 8656 4102 8666
rect 4105 8656 4107 8663
rect 4121 8656 4123 8675
rect 4137 8666 4139 8675
rect 4142 8673 4144 8675
rect 4163 8673 4165 8675
rect 4179 8672 4181 8675
rect 4137 8656 4139 8659
rect 4142 8656 4144 8658
rect 4163 8656 4165 8658
rect 4179 8656 4181 8668
rect 4195 8666 4197 8675
rect 4200 8673 4202 8675
rect 4195 8656 4197 8659
rect 4200 8656 4202 8658
rect 4216 8656 4218 8675
rect 2372 8653 2374 8655
rect 2377 8653 2379 8656
rect 2393 8653 2395 8655
rect 2409 8653 2411 8655
rect 2414 8653 2416 8656
rect 2435 8653 2437 8656
rect 2451 8653 2453 8656
rect 2467 8653 2469 8655
rect 2472 8653 2474 8656
rect 2488 8653 2490 8655
rect 2504 8653 2506 8655
rect 2509 8653 2511 8656
rect 2525 8653 2527 8655
rect 2541 8653 2543 8655
rect 2546 8653 2548 8656
rect 2567 8653 2569 8656
rect 2583 8653 2585 8656
rect 2599 8653 2601 8655
rect 2604 8653 2606 8656
rect 2620 8653 2622 8655
rect 2636 8653 2638 8655
rect 2641 8653 2643 8656
rect 2657 8653 2659 8655
rect 2673 8653 2675 8655
rect 2678 8653 2680 8656
rect 2699 8653 2701 8656
rect 2715 8653 2717 8656
rect 2731 8653 2733 8655
rect 2736 8653 2738 8656
rect 2752 8653 2754 8655
rect 3317 8653 3319 8655
rect 3322 8653 3324 8656
rect 3338 8653 3340 8655
rect 3354 8653 3356 8655
rect 3359 8653 3361 8656
rect 3380 8653 3382 8656
rect 3396 8653 3398 8656
rect 3412 8653 3414 8655
rect 3417 8653 3419 8656
rect 3433 8653 3435 8655
rect 3449 8653 3451 8655
rect 3454 8653 3456 8656
rect 3470 8653 3472 8655
rect 3486 8653 3488 8655
rect 3491 8653 3493 8656
rect 3512 8653 3514 8656
rect 3528 8653 3530 8656
rect 3544 8653 3546 8655
rect 3549 8653 3551 8656
rect 3565 8653 3567 8655
rect 3581 8653 3583 8655
rect 3586 8653 3588 8656
rect 3602 8653 3604 8655
rect 3618 8653 3620 8655
rect 3623 8653 3625 8656
rect 3644 8653 3646 8656
rect 3660 8653 3662 8656
rect 3676 8653 3678 8655
rect 3681 8653 3683 8656
rect 3697 8653 3699 8655
rect 3155 8650 3157 8652
rect 3160 8649 3162 8652
rect 3176 8650 3178 8652
rect 3192 8650 3194 8652
rect 3197 8647 3199 8652
rect 3218 8647 3220 8652
rect 3234 8650 3236 8652
rect 3250 8650 3252 8652
rect 3255 8647 3257 8652
rect 3271 8650 3273 8652
rect 2372 8640 2374 8645
rect 2377 8643 2379 8645
rect 2372 8626 2374 8636
rect 2377 8626 2379 8633
rect 2393 8626 2395 8645
rect 2409 8636 2411 8645
rect 2414 8643 2416 8645
rect 2435 8643 2437 8645
rect 2451 8642 2453 8645
rect 2409 8626 2411 8629
rect 2414 8626 2416 8628
rect 2435 8626 2437 8628
rect 2451 8626 2453 8638
rect 2467 8636 2469 8645
rect 2472 8643 2474 8645
rect 2467 8626 2469 8629
rect 2472 8626 2474 8628
rect 2488 8626 2490 8645
rect 2504 8642 2506 8645
rect 2509 8643 2511 8645
rect 2504 8626 2506 8638
rect 2509 8626 2511 8633
rect 2525 8626 2527 8645
rect 2541 8636 2543 8645
rect 2546 8643 2548 8645
rect 2567 8643 2569 8645
rect 2583 8642 2585 8645
rect 2541 8626 2543 8629
rect 2546 8626 2548 8628
rect 2567 8626 2569 8628
rect 2583 8626 2585 8638
rect 2599 8636 2601 8645
rect 2604 8643 2606 8645
rect 2599 8626 2601 8629
rect 2604 8626 2606 8628
rect 2620 8626 2622 8645
rect 2636 8642 2638 8645
rect 2641 8643 2643 8645
rect 2636 8626 2638 8638
rect 2641 8626 2643 8633
rect 2657 8626 2659 8645
rect 2673 8636 2675 8645
rect 2678 8643 2680 8645
rect 2699 8643 2701 8645
rect 2715 8642 2717 8645
rect 2673 8626 2675 8629
rect 2678 8626 2680 8628
rect 2699 8626 2701 8628
rect 2715 8626 2717 8638
rect 2731 8636 2733 8645
rect 2736 8643 2738 8645
rect 2752 8637 2754 8645
rect 4100 8650 4102 8652
rect 4105 8649 4107 8652
rect 4121 8650 4123 8652
rect 4137 8650 4139 8652
rect 4142 8647 4144 8652
rect 4163 8647 4165 8652
rect 4179 8650 4181 8652
rect 4195 8650 4197 8652
rect 4200 8647 4202 8652
rect 4216 8650 4218 8652
rect 3317 8640 3319 8645
rect 3322 8643 3324 8645
rect 2731 8626 2733 8629
rect 2736 8626 2738 8628
rect 2752 8626 2754 8633
rect 3317 8626 3319 8636
rect 3322 8626 3324 8633
rect 3338 8626 3340 8645
rect 3354 8636 3356 8645
rect 3359 8643 3361 8645
rect 3380 8643 3382 8645
rect 3396 8642 3398 8645
rect 3354 8626 3356 8629
rect 3359 8626 3361 8628
rect 3380 8626 3382 8628
rect 3396 8626 3398 8638
rect 3412 8636 3414 8645
rect 3417 8643 3419 8645
rect 3412 8626 3414 8629
rect 3417 8626 3419 8628
rect 3433 8626 3435 8645
rect 3449 8642 3451 8645
rect 3454 8643 3456 8645
rect 3449 8626 3451 8638
rect 3454 8626 3456 8633
rect 3470 8626 3472 8645
rect 3486 8636 3488 8645
rect 3491 8643 3493 8645
rect 3512 8643 3514 8645
rect 3528 8642 3530 8645
rect 3486 8626 3488 8629
rect 3491 8626 3493 8628
rect 3512 8626 3514 8628
rect 3528 8626 3530 8638
rect 3544 8636 3546 8645
rect 3549 8643 3551 8645
rect 3544 8626 3546 8629
rect 3549 8626 3551 8628
rect 3565 8626 3567 8645
rect 3581 8642 3583 8645
rect 3586 8643 3588 8645
rect 3581 8626 3583 8638
rect 3586 8626 3588 8633
rect 3602 8626 3604 8645
rect 3618 8636 3620 8645
rect 3623 8643 3625 8645
rect 3644 8643 3646 8645
rect 3660 8642 3662 8645
rect 3618 8626 3620 8629
rect 3623 8626 3625 8628
rect 3644 8626 3646 8628
rect 3660 8626 3662 8638
rect 3676 8636 3678 8645
rect 3681 8643 3683 8645
rect 3697 8637 3699 8645
rect 3676 8626 3678 8629
rect 3681 8626 3683 8628
rect 3697 8626 3699 8633
rect 2372 8620 2374 8622
rect 2377 8619 2379 8622
rect 2393 8620 2395 8622
rect 2409 8620 2411 8622
rect 2414 8617 2416 8622
rect 2435 8617 2437 8622
rect 2451 8620 2453 8622
rect 2467 8620 2469 8622
rect 2472 8617 2474 8622
rect 2488 8620 2490 8622
rect 2504 8620 2506 8622
rect 2509 8619 2511 8622
rect 2525 8620 2527 8622
rect 2541 8620 2543 8622
rect 2546 8617 2548 8622
rect 2567 8617 2569 8622
rect 2583 8620 2585 8622
rect 2599 8620 2601 8622
rect 2604 8617 2606 8622
rect 2620 8620 2622 8622
rect 2636 8620 2638 8622
rect 2641 8619 2643 8622
rect 2657 8620 2659 8622
rect 2673 8620 2675 8622
rect 2678 8617 2680 8622
rect 2699 8617 2701 8622
rect 2715 8620 2717 8622
rect 2731 8620 2733 8622
rect 2736 8617 2738 8622
rect 2752 8620 2754 8622
rect 3317 8620 3319 8622
rect 3322 8619 3324 8622
rect 3338 8620 3340 8622
rect 3354 8620 3356 8622
rect 3359 8617 3361 8622
rect 3380 8617 3382 8622
rect 3396 8620 3398 8622
rect 3412 8620 3414 8622
rect 3417 8617 3419 8622
rect 3433 8620 3435 8622
rect 3449 8620 3451 8622
rect 3454 8619 3456 8622
rect 3470 8620 3472 8622
rect 3486 8620 3488 8622
rect 3491 8617 3493 8622
rect 3512 8617 3514 8622
rect 3528 8620 3530 8622
rect 3544 8620 3546 8622
rect 3549 8617 3551 8622
rect 3565 8620 3567 8622
rect 3581 8620 3583 8622
rect 3586 8619 3588 8622
rect 3602 8620 3604 8622
rect 3618 8620 3620 8622
rect 3623 8617 3625 8622
rect 3644 8617 3646 8622
rect 3660 8620 3662 8622
rect 3676 8620 3678 8622
rect 3681 8617 3683 8622
rect 3697 8620 3699 8622
rect 3155 8597 3157 8599
rect 3160 8597 3162 8600
rect 3176 8597 3178 8599
rect 3192 8597 3194 8599
rect 3197 8597 3199 8600
rect 3218 8597 3220 8600
rect 3234 8597 3236 8600
rect 3250 8597 3252 8599
rect 3255 8597 3257 8600
rect 3271 8597 3273 8599
rect 4100 8597 4102 8599
rect 4105 8597 4107 8600
rect 4121 8597 4123 8599
rect 4137 8597 4139 8599
rect 4142 8597 4144 8600
rect 4163 8597 4165 8600
rect 4179 8597 4181 8600
rect 4195 8597 4197 8599
rect 4200 8597 4202 8600
rect 4216 8597 4218 8599
rect 3155 8584 3157 8589
rect 3160 8587 3162 8589
rect 3155 8570 3157 8580
rect 3160 8570 3162 8577
rect 3176 8570 3178 8589
rect 3192 8580 3194 8589
rect 3197 8587 3199 8589
rect 3218 8587 3220 8589
rect 3234 8586 3236 8589
rect 3192 8570 3194 8573
rect 3197 8570 3199 8572
rect 3218 8570 3220 8572
rect 3234 8570 3236 8582
rect 3250 8580 3252 8589
rect 3255 8587 3257 8589
rect 3250 8570 3252 8573
rect 3255 8570 3257 8572
rect 3271 8570 3273 8589
rect 4100 8584 4102 8589
rect 4105 8587 4107 8589
rect 3293 8576 3296 8578
rect 3300 8576 3303 8578
rect 4100 8570 4102 8580
rect 4105 8570 4107 8577
rect 4121 8570 4123 8589
rect 4137 8580 4139 8589
rect 4142 8587 4144 8589
rect 4163 8587 4165 8589
rect 4179 8586 4181 8589
rect 4137 8570 4139 8573
rect 4142 8570 4144 8572
rect 4163 8570 4165 8572
rect 4179 8570 4181 8582
rect 4195 8580 4197 8589
rect 4200 8587 4202 8589
rect 4195 8570 4197 8573
rect 4200 8570 4202 8572
rect 4216 8570 4218 8589
rect 4238 8576 4241 8578
rect 4245 8576 4248 8578
rect 2372 8567 2374 8569
rect 2377 8567 2379 8570
rect 2393 8567 2395 8569
rect 2409 8567 2411 8569
rect 2414 8567 2416 8570
rect 2435 8567 2437 8570
rect 2451 8567 2453 8570
rect 2467 8567 2469 8569
rect 2472 8567 2474 8570
rect 2488 8567 2490 8569
rect 2504 8567 2506 8569
rect 2509 8567 2511 8570
rect 2525 8567 2527 8569
rect 2541 8567 2543 8569
rect 2546 8567 2548 8570
rect 2567 8567 2569 8570
rect 2583 8567 2585 8570
rect 2599 8567 2601 8569
rect 2604 8567 2606 8570
rect 2620 8567 2622 8569
rect 2636 8567 2638 8569
rect 2641 8567 2643 8570
rect 2657 8567 2659 8569
rect 2673 8567 2675 8569
rect 2678 8567 2680 8570
rect 2699 8567 2701 8570
rect 2715 8567 2717 8570
rect 2731 8567 2733 8569
rect 2736 8567 2738 8570
rect 2752 8567 2754 8569
rect 3317 8567 3319 8569
rect 3322 8567 3324 8570
rect 3338 8567 3340 8569
rect 3354 8567 3356 8569
rect 3359 8567 3361 8570
rect 3380 8567 3382 8570
rect 3396 8567 3398 8570
rect 3412 8567 3414 8569
rect 3417 8567 3419 8570
rect 3433 8567 3435 8569
rect 3449 8567 3451 8569
rect 3454 8567 3456 8570
rect 3470 8567 3472 8569
rect 3486 8567 3488 8569
rect 3491 8567 3493 8570
rect 3512 8567 3514 8570
rect 3528 8567 3530 8570
rect 3544 8567 3546 8569
rect 3549 8567 3551 8570
rect 3565 8567 3567 8569
rect 3581 8567 3583 8569
rect 3586 8567 3588 8570
rect 3602 8567 3604 8569
rect 3618 8567 3620 8569
rect 3623 8567 3625 8570
rect 3644 8567 3646 8570
rect 3660 8567 3662 8570
rect 3676 8567 3678 8569
rect 3681 8567 3683 8570
rect 3697 8567 3699 8569
rect 3155 8564 3157 8566
rect 3160 8563 3162 8566
rect 3176 8564 3178 8566
rect 3192 8564 3194 8566
rect 3197 8561 3199 8566
rect 3218 8561 3220 8566
rect 3234 8564 3236 8566
rect 3250 8564 3252 8566
rect 3255 8561 3257 8566
rect 3271 8564 3273 8566
rect 2372 8554 2374 8559
rect 2377 8557 2379 8559
rect 2372 8540 2374 8550
rect 2377 8540 2379 8547
rect 2393 8540 2395 8559
rect 2409 8550 2411 8559
rect 2414 8557 2416 8559
rect 2435 8557 2437 8559
rect 2451 8556 2453 8559
rect 2409 8540 2411 8543
rect 2414 8540 2416 8542
rect 2435 8540 2437 8542
rect 2451 8540 2453 8552
rect 2467 8550 2469 8559
rect 2472 8557 2474 8559
rect 2467 8540 2469 8543
rect 2472 8540 2474 8542
rect 2488 8540 2490 8559
rect 2504 8556 2506 8559
rect 2509 8557 2511 8559
rect 2504 8540 2506 8552
rect 2509 8540 2511 8547
rect 2525 8540 2527 8559
rect 2541 8550 2543 8559
rect 2546 8557 2548 8559
rect 2567 8557 2569 8559
rect 2583 8556 2585 8559
rect 2541 8540 2543 8543
rect 2546 8540 2548 8542
rect 2567 8540 2569 8542
rect 2583 8540 2585 8552
rect 2599 8550 2601 8559
rect 2604 8557 2606 8559
rect 2599 8540 2601 8543
rect 2604 8540 2606 8542
rect 2620 8540 2622 8559
rect 2636 8556 2638 8559
rect 2641 8557 2643 8559
rect 2636 8540 2638 8552
rect 2641 8540 2643 8547
rect 2657 8540 2659 8559
rect 2673 8550 2675 8559
rect 2678 8557 2680 8559
rect 2699 8557 2701 8559
rect 2715 8556 2717 8559
rect 2673 8540 2675 8543
rect 2678 8540 2680 8542
rect 2699 8540 2701 8542
rect 2715 8540 2717 8552
rect 2731 8550 2733 8559
rect 2736 8557 2738 8559
rect 2752 8551 2754 8559
rect 4100 8564 4102 8566
rect 4105 8563 4107 8566
rect 4121 8564 4123 8566
rect 4137 8564 4139 8566
rect 4142 8561 4144 8566
rect 4163 8561 4165 8566
rect 4179 8564 4181 8566
rect 4195 8564 4197 8566
rect 4200 8561 4202 8566
rect 4216 8564 4218 8566
rect 3317 8554 3319 8559
rect 3322 8557 3324 8559
rect 2731 8540 2733 8543
rect 2736 8540 2738 8542
rect 2752 8540 2754 8547
rect 3317 8540 3319 8550
rect 3322 8540 3324 8547
rect 3338 8540 3340 8559
rect 3354 8550 3356 8559
rect 3359 8557 3361 8559
rect 3380 8557 3382 8559
rect 3396 8556 3398 8559
rect 3354 8540 3356 8543
rect 3359 8540 3361 8542
rect 3380 8540 3382 8542
rect 3396 8540 3398 8552
rect 3412 8550 3414 8559
rect 3417 8557 3419 8559
rect 3412 8540 3414 8543
rect 3417 8540 3419 8542
rect 3433 8540 3435 8559
rect 3449 8556 3451 8559
rect 3454 8557 3456 8559
rect 3449 8540 3451 8552
rect 3454 8540 3456 8547
rect 3470 8540 3472 8559
rect 3486 8550 3488 8559
rect 3491 8557 3493 8559
rect 3512 8557 3514 8559
rect 3528 8556 3530 8559
rect 3486 8540 3488 8543
rect 3491 8540 3493 8542
rect 3512 8540 3514 8542
rect 3528 8540 3530 8552
rect 3544 8550 3546 8559
rect 3549 8557 3551 8559
rect 3544 8540 3546 8543
rect 3549 8540 3551 8542
rect 3565 8540 3567 8559
rect 3581 8556 3583 8559
rect 3586 8557 3588 8559
rect 3581 8540 3583 8552
rect 3586 8540 3588 8547
rect 3602 8540 3604 8559
rect 3618 8550 3620 8559
rect 3623 8557 3625 8559
rect 3644 8557 3646 8559
rect 3660 8556 3662 8559
rect 3618 8540 3620 8543
rect 3623 8540 3625 8542
rect 3644 8540 3646 8542
rect 3660 8540 3662 8552
rect 3676 8550 3678 8559
rect 3681 8557 3683 8559
rect 3697 8551 3699 8559
rect 3676 8540 3678 8543
rect 3681 8540 3683 8542
rect 3697 8540 3699 8547
rect 2372 8534 2374 8536
rect 2377 8533 2379 8536
rect 2393 8534 2395 8536
rect 2409 8534 2411 8536
rect 2414 8531 2416 8536
rect 2435 8531 2437 8536
rect 2451 8534 2453 8536
rect 2467 8534 2469 8536
rect 2472 8531 2474 8536
rect 2488 8534 2490 8536
rect 2504 8534 2506 8536
rect 2509 8533 2511 8536
rect 2525 8534 2527 8536
rect 2541 8534 2543 8536
rect 2546 8531 2548 8536
rect 2567 8531 2569 8536
rect 2583 8534 2585 8536
rect 2599 8534 2601 8536
rect 2604 8531 2606 8536
rect 2620 8534 2622 8536
rect 2636 8534 2638 8536
rect 2641 8533 2643 8536
rect 2657 8534 2659 8536
rect 2673 8534 2675 8536
rect 2678 8531 2680 8536
rect 2699 8531 2701 8536
rect 2715 8534 2717 8536
rect 2731 8534 2733 8536
rect 2736 8531 2738 8536
rect 2752 8534 2754 8536
rect 3317 8534 3319 8536
rect 3322 8533 3324 8536
rect 3338 8534 3340 8536
rect 3354 8534 3356 8536
rect 3359 8531 3361 8536
rect 3380 8531 3382 8536
rect 3396 8534 3398 8536
rect 3412 8534 3414 8536
rect 3417 8531 3419 8536
rect 3433 8534 3435 8536
rect 3449 8534 3451 8536
rect 3454 8533 3456 8536
rect 3470 8534 3472 8536
rect 3486 8534 3488 8536
rect 3491 8531 3493 8536
rect 3512 8531 3514 8536
rect 3528 8534 3530 8536
rect 3544 8534 3546 8536
rect 3549 8531 3551 8536
rect 3565 8534 3567 8536
rect 3581 8534 3583 8536
rect 3586 8533 3588 8536
rect 3602 8534 3604 8536
rect 3618 8534 3620 8536
rect 3623 8531 3625 8536
rect 3644 8531 3646 8536
rect 3660 8534 3662 8536
rect 3676 8534 3678 8536
rect 3681 8531 3683 8536
rect 3697 8534 3699 8536
rect 2604 8496 2606 8499
rect 2628 8496 2630 8499
rect 3549 8496 3551 8499
rect 3573 8496 3575 8499
rect 2604 8490 2606 8492
rect 2628 8490 2630 8492
rect 3549 8490 3551 8492
rect 3573 8490 3575 8492
rect 2624 8485 2626 8487
rect 3569 8485 3571 8487
rect 2624 8478 2626 8481
rect 3569 8478 3571 8481
rect 2613 8467 2615 8469
rect 2619 8467 2638 8469
rect 3558 8467 3560 8469
rect 3564 8467 3583 8469
rect 2604 8462 2606 8464
rect 2628 8462 2630 8464
rect 3549 8462 3551 8464
rect 3573 8462 3575 8464
rect 2604 8455 2606 8458
rect 2628 8455 2630 8458
rect 3549 8455 3551 8458
rect 3573 8455 3575 8458
rect 2372 8427 2374 8429
rect 2377 8427 2379 8430
rect 2393 8427 2395 8429
rect 2409 8427 2411 8429
rect 2414 8427 2416 8430
rect 2435 8427 2437 8430
rect 2451 8427 2453 8430
rect 2467 8427 2469 8429
rect 2472 8427 2474 8430
rect 2488 8427 2490 8429
rect 2504 8427 2506 8429
rect 2509 8427 2511 8430
rect 2525 8427 2527 8429
rect 2541 8427 2543 8429
rect 2546 8427 2548 8430
rect 2567 8427 2569 8430
rect 2583 8427 2585 8430
rect 2599 8427 2601 8429
rect 2604 8427 2606 8430
rect 2620 8427 2622 8429
rect 2636 8427 2638 8429
rect 2641 8427 2643 8430
rect 2657 8427 2659 8429
rect 2673 8427 2675 8429
rect 2678 8427 2680 8430
rect 2699 8427 2701 8430
rect 2715 8427 2717 8430
rect 2731 8427 2733 8429
rect 2736 8427 2738 8430
rect 2752 8427 2754 8429
rect 3317 8427 3319 8429
rect 3322 8427 3324 8430
rect 3338 8427 3340 8429
rect 3354 8427 3356 8429
rect 3359 8427 3361 8430
rect 3380 8427 3382 8430
rect 3396 8427 3398 8430
rect 3412 8427 3414 8429
rect 3417 8427 3419 8430
rect 3433 8427 3435 8429
rect 3449 8427 3451 8429
rect 3454 8427 3456 8430
rect 3470 8427 3472 8429
rect 3486 8427 3488 8429
rect 3491 8427 3493 8430
rect 3512 8427 3514 8430
rect 3528 8427 3530 8430
rect 3544 8427 3546 8429
rect 3549 8427 3551 8430
rect 3565 8427 3567 8429
rect 3581 8427 3583 8429
rect 3586 8427 3588 8430
rect 3602 8427 3604 8429
rect 3618 8427 3620 8429
rect 3623 8427 3625 8430
rect 3644 8427 3646 8430
rect 3660 8427 3662 8430
rect 3676 8427 3678 8429
rect 3681 8427 3683 8430
rect 3697 8427 3699 8429
rect 2372 8414 2374 8419
rect 2377 8417 2379 8419
rect 2372 8400 2374 8410
rect 2377 8400 2379 8407
rect 2393 8400 2395 8419
rect 2409 8410 2411 8419
rect 2414 8417 2416 8419
rect 2435 8417 2437 8419
rect 2451 8416 2453 8419
rect 2409 8400 2411 8403
rect 2414 8400 2416 8402
rect 2435 8400 2437 8402
rect 2451 8400 2453 8412
rect 2467 8410 2469 8419
rect 2472 8417 2474 8419
rect 2467 8400 2469 8403
rect 2472 8400 2474 8402
rect 2488 8400 2490 8419
rect 2504 8416 2506 8419
rect 2509 8417 2511 8419
rect 2504 8400 2506 8412
rect 2509 8400 2511 8407
rect 2525 8400 2527 8419
rect 2541 8410 2543 8419
rect 2546 8417 2548 8419
rect 2567 8417 2569 8419
rect 2583 8416 2585 8419
rect 2541 8400 2543 8403
rect 2546 8400 2548 8402
rect 2567 8400 2569 8402
rect 2583 8400 2585 8412
rect 2599 8410 2601 8419
rect 2604 8417 2606 8419
rect 2599 8400 2601 8403
rect 2604 8400 2606 8402
rect 2620 8400 2622 8419
rect 2636 8416 2638 8419
rect 2641 8417 2643 8419
rect 2636 8400 2638 8412
rect 2641 8400 2643 8407
rect 2657 8400 2659 8419
rect 2673 8410 2675 8419
rect 2678 8417 2680 8419
rect 2699 8417 2701 8419
rect 2715 8416 2717 8419
rect 2673 8400 2675 8403
rect 2678 8400 2680 8402
rect 2699 8400 2701 8402
rect 2715 8400 2717 8412
rect 2731 8410 2733 8419
rect 2736 8417 2738 8419
rect 2752 8411 2754 8419
rect 3317 8414 3319 8419
rect 3322 8417 3324 8419
rect 2731 8400 2733 8403
rect 2736 8400 2738 8402
rect 2752 8400 2754 8407
rect 3317 8400 3319 8410
rect 3322 8400 3324 8407
rect 3338 8400 3340 8419
rect 3354 8410 3356 8419
rect 3359 8417 3361 8419
rect 3380 8417 3382 8419
rect 3396 8416 3398 8419
rect 3354 8400 3356 8403
rect 3359 8400 3361 8402
rect 3380 8400 3382 8402
rect 3396 8400 3398 8412
rect 3412 8410 3414 8419
rect 3417 8417 3419 8419
rect 3412 8400 3414 8403
rect 3417 8400 3419 8402
rect 3433 8400 3435 8419
rect 3449 8416 3451 8419
rect 3454 8417 3456 8419
rect 3449 8400 3451 8412
rect 3454 8400 3456 8407
rect 3470 8400 3472 8419
rect 3486 8410 3488 8419
rect 3491 8417 3493 8419
rect 3512 8417 3514 8419
rect 3528 8416 3530 8419
rect 3486 8400 3488 8403
rect 3491 8400 3493 8402
rect 3512 8400 3514 8402
rect 3528 8400 3530 8412
rect 3544 8410 3546 8419
rect 3549 8417 3551 8419
rect 3544 8400 3546 8403
rect 3549 8400 3551 8402
rect 3565 8400 3567 8419
rect 3581 8416 3583 8419
rect 3586 8417 3588 8419
rect 3581 8400 3583 8412
rect 3586 8400 3588 8407
rect 3602 8400 3604 8419
rect 3618 8410 3620 8419
rect 3623 8417 3625 8419
rect 3644 8417 3646 8419
rect 3660 8416 3662 8419
rect 3618 8400 3620 8403
rect 3623 8400 3625 8402
rect 3644 8400 3646 8402
rect 3660 8400 3662 8412
rect 3676 8410 3678 8419
rect 3681 8417 3683 8419
rect 3697 8411 3699 8419
rect 3676 8400 3678 8403
rect 3681 8400 3683 8402
rect 3697 8400 3699 8407
rect 2372 8394 2374 8396
rect 2377 8393 2379 8396
rect 2393 8394 2395 8396
rect 2409 8394 2411 8396
rect 2414 8391 2416 8396
rect 2435 8391 2437 8396
rect 2451 8394 2453 8396
rect 2467 8394 2469 8396
rect 2472 8391 2474 8396
rect 2488 8394 2490 8396
rect 2504 8394 2506 8396
rect 2509 8393 2511 8396
rect 2525 8394 2527 8396
rect 2541 8394 2543 8396
rect 2546 8391 2548 8396
rect 2567 8391 2569 8396
rect 2583 8394 2585 8396
rect 2599 8394 2601 8396
rect 2604 8391 2606 8396
rect 2620 8394 2622 8396
rect 2636 8394 2638 8396
rect 2641 8393 2643 8396
rect 2657 8394 2659 8396
rect 2673 8394 2675 8396
rect 2678 8391 2680 8396
rect 2699 8391 2701 8396
rect 2715 8394 2717 8396
rect 2731 8394 2733 8396
rect 2736 8391 2738 8396
rect 2752 8394 2754 8396
rect 3317 8394 3319 8396
rect 3322 8393 3324 8396
rect 3338 8394 3340 8396
rect 3354 8394 3356 8396
rect 3359 8391 3361 8396
rect 3380 8391 3382 8396
rect 3396 8394 3398 8396
rect 3412 8394 3414 8396
rect 3417 8391 3419 8396
rect 3433 8394 3435 8396
rect 3449 8394 3451 8396
rect 3454 8393 3456 8396
rect 3470 8394 3472 8396
rect 3486 8394 3488 8396
rect 3491 8391 3493 8396
rect 3512 8391 3514 8396
rect 3528 8394 3530 8396
rect 3544 8394 3546 8396
rect 3549 8391 3551 8396
rect 3565 8394 3567 8396
rect 3581 8394 3583 8396
rect 3586 8393 3588 8396
rect 3602 8394 3604 8396
rect 3618 8394 3620 8396
rect 3623 8391 3625 8396
rect 3644 8391 3646 8396
rect 3660 8394 3662 8396
rect 3676 8394 3678 8396
rect 3681 8391 3683 8396
rect 3697 8394 3699 8396
rect 2856 8348 2858 8350
rect 2861 8348 2863 8351
rect 2877 8348 2879 8350
rect 2893 8348 2895 8350
rect 2898 8348 2900 8351
rect 2919 8348 2921 8351
rect 2935 8348 2937 8351
rect 2951 8348 2953 8350
rect 2956 8348 2958 8351
rect 2972 8348 2974 8350
rect 2988 8348 2990 8350
rect 2993 8348 2995 8351
rect 3009 8348 3011 8350
rect 3025 8348 3027 8350
rect 3030 8348 3032 8351
rect 3051 8348 3053 8351
rect 3067 8348 3069 8351
rect 3083 8348 3085 8350
rect 3088 8348 3090 8351
rect 3104 8348 3106 8350
rect 3120 8348 3122 8350
rect 3125 8348 3127 8351
rect 3141 8348 3143 8350
rect 3157 8348 3159 8350
rect 3162 8348 3164 8351
rect 3183 8348 3185 8351
rect 3199 8348 3201 8351
rect 3215 8348 3217 8350
rect 3220 8348 3222 8351
rect 3236 8348 3238 8350
rect 3252 8348 3254 8350
rect 3257 8348 3259 8351
rect 3273 8348 3275 8350
rect 3289 8348 3291 8350
rect 3294 8348 3296 8351
rect 3315 8348 3317 8351
rect 3331 8348 3333 8351
rect 3347 8348 3349 8350
rect 3352 8348 3354 8351
rect 3368 8348 3370 8350
rect 3801 8348 3803 8350
rect 3806 8348 3808 8351
rect 3822 8348 3824 8350
rect 3838 8348 3840 8350
rect 3843 8348 3845 8351
rect 3864 8348 3866 8351
rect 3880 8348 3882 8351
rect 3896 8348 3898 8350
rect 3901 8348 3903 8351
rect 3917 8348 3919 8350
rect 3933 8348 3935 8350
rect 3938 8348 3940 8351
rect 3954 8348 3956 8350
rect 3970 8348 3972 8350
rect 3975 8348 3977 8351
rect 3996 8348 3998 8351
rect 4012 8348 4014 8351
rect 4028 8348 4030 8350
rect 4033 8348 4035 8351
rect 4049 8348 4051 8350
rect 4065 8348 4067 8350
rect 4070 8348 4072 8351
rect 4086 8348 4088 8350
rect 4102 8348 4104 8350
rect 4107 8348 4109 8351
rect 4128 8348 4130 8351
rect 4144 8348 4146 8351
rect 4160 8348 4162 8350
rect 4165 8348 4167 8351
rect 4181 8348 4183 8350
rect 4197 8348 4199 8350
rect 4202 8348 4204 8351
rect 4218 8348 4220 8350
rect 4234 8348 4236 8350
rect 4239 8348 4241 8351
rect 4260 8348 4262 8351
rect 4276 8348 4278 8351
rect 4292 8348 4294 8350
rect 4297 8348 4299 8351
rect 4313 8348 4315 8350
rect 2856 8335 2858 8340
rect 2861 8338 2863 8340
rect 2856 8321 2858 8331
rect 2861 8321 2863 8328
rect 2877 8321 2879 8340
rect 2893 8331 2895 8340
rect 2898 8338 2900 8340
rect 2919 8338 2921 8340
rect 2935 8337 2937 8340
rect 2893 8321 2895 8324
rect 2898 8321 2900 8323
rect 2919 8321 2921 8323
rect 2935 8321 2937 8333
rect 2951 8331 2953 8340
rect 2956 8338 2958 8340
rect 2972 8332 2974 8340
rect 2988 8335 2990 8340
rect 2993 8338 2995 8340
rect 2951 8321 2953 8324
rect 2956 8321 2958 8323
rect 2972 8321 2974 8328
rect 2988 8321 2990 8331
rect 2993 8321 2995 8328
rect 3009 8321 3011 8340
rect 3025 8331 3027 8340
rect 3030 8338 3032 8340
rect 3051 8338 3053 8340
rect 3067 8337 3069 8340
rect 3025 8321 3027 8324
rect 3030 8321 3032 8323
rect 3051 8321 3053 8323
rect 3067 8321 3069 8333
rect 3083 8331 3085 8340
rect 3088 8338 3090 8340
rect 3104 8332 3106 8340
rect 3120 8335 3122 8340
rect 3125 8338 3127 8340
rect 3083 8321 3085 8324
rect 3088 8321 3090 8323
rect 3104 8321 3106 8328
rect 3120 8321 3122 8331
rect 3125 8321 3127 8328
rect 3141 8321 3143 8340
rect 3157 8331 3159 8340
rect 3162 8338 3164 8340
rect 3183 8338 3185 8340
rect 3199 8337 3201 8340
rect 3157 8321 3159 8324
rect 3162 8321 3164 8323
rect 3183 8321 3185 8323
rect 3199 8321 3201 8333
rect 3215 8331 3217 8340
rect 3220 8338 3222 8340
rect 3236 8332 3238 8340
rect 3252 8335 3254 8340
rect 3257 8338 3259 8340
rect 3215 8321 3217 8324
rect 3220 8321 3222 8323
rect 3236 8321 3238 8328
rect 3252 8321 3254 8331
rect 3257 8321 3259 8328
rect 3273 8321 3275 8340
rect 3289 8331 3291 8340
rect 3294 8338 3296 8340
rect 3315 8338 3317 8340
rect 3331 8337 3333 8340
rect 3289 8321 3291 8324
rect 3294 8321 3296 8323
rect 3315 8321 3317 8323
rect 3331 8321 3333 8333
rect 3347 8331 3349 8340
rect 3352 8338 3354 8340
rect 3368 8332 3370 8340
rect 3801 8335 3803 8340
rect 3806 8338 3808 8340
rect 3347 8321 3349 8324
rect 3352 8321 3354 8323
rect 3368 8321 3370 8328
rect 2504 8315 2506 8317
rect 2509 8315 2511 8318
rect 2525 8315 2527 8317
rect 2541 8315 2543 8317
rect 2546 8315 2548 8318
rect 2567 8315 2569 8318
rect 2583 8315 2585 8318
rect 2599 8315 2601 8317
rect 2604 8315 2606 8318
rect 3801 8321 3803 8331
rect 3806 8321 3808 8328
rect 3822 8321 3824 8340
rect 3838 8331 3840 8340
rect 3843 8338 3845 8340
rect 3864 8338 3866 8340
rect 3880 8337 3882 8340
rect 3838 8321 3840 8324
rect 3843 8321 3845 8323
rect 3864 8321 3866 8323
rect 3880 8321 3882 8333
rect 3896 8331 3898 8340
rect 3901 8338 3903 8340
rect 3917 8332 3919 8340
rect 3933 8335 3935 8340
rect 3938 8338 3940 8340
rect 3896 8321 3898 8324
rect 3901 8321 3903 8323
rect 3917 8321 3919 8328
rect 3933 8321 3935 8331
rect 3938 8321 3940 8328
rect 3954 8321 3956 8340
rect 3970 8331 3972 8340
rect 3975 8338 3977 8340
rect 3996 8338 3998 8340
rect 4012 8337 4014 8340
rect 3970 8321 3972 8324
rect 3975 8321 3977 8323
rect 3996 8321 3998 8323
rect 4012 8321 4014 8333
rect 4028 8331 4030 8340
rect 4033 8338 4035 8340
rect 4049 8332 4051 8340
rect 4065 8335 4067 8340
rect 4070 8338 4072 8340
rect 4028 8321 4030 8324
rect 4033 8321 4035 8323
rect 4049 8321 4051 8328
rect 4065 8321 4067 8331
rect 4070 8321 4072 8328
rect 4086 8321 4088 8340
rect 4102 8331 4104 8340
rect 4107 8338 4109 8340
rect 4128 8338 4130 8340
rect 4144 8337 4146 8340
rect 4102 8321 4104 8324
rect 4107 8321 4109 8323
rect 4128 8321 4130 8323
rect 4144 8321 4146 8333
rect 4160 8331 4162 8340
rect 4165 8338 4167 8340
rect 4181 8332 4183 8340
rect 4197 8335 4199 8340
rect 4202 8338 4204 8340
rect 4160 8321 4162 8324
rect 4165 8321 4167 8323
rect 4181 8321 4183 8328
rect 4197 8321 4199 8331
rect 4202 8321 4204 8328
rect 4218 8321 4220 8340
rect 4234 8331 4236 8340
rect 4239 8338 4241 8340
rect 4260 8338 4262 8340
rect 4276 8337 4278 8340
rect 4234 8321 4236 8324
rect 4239 8321 4241 8323
rect 4260 8321 4262 8323
rect 4276 8321 4278 8333
rect 4292 8331 4294 8340
rect 4297 8338 4299 8340
rect 4313 8332 4315 8340
rect 4292 8321 4294 8324
rect 4297 8321 4299 8323
rect 4313 8321 4315 8328
rect 2620 8315 2622 8317
rect 2856 8315 2858 8317
rect 2861 8314 2863 8317
rect 2877 8315 2879 8317
rect 2893 8315 2895 8317
rect 2898 8312 2900 8317
rect 2919 8312 2921 8317
rect 2935 8315 2937 8317
rect 2951 8315 2953 8317
rect 2956 8312 2958 8317
rect 2972 8315 2974 8317
rect 2988 8315 2990 8317
rect 2993 8314 2995 8317
rect 3009 8315 3011 8317
rect 3025 8315 3027 8317
rect 3030 8312 3032 8317
rect 3051 8312 3053 8317
rect 3067 8315 3069 8317
rect 3083 8315 3085 8317
rect 3088 8312 3090 8317
rect 3104 8315 3106 8317
rect 3120 8315 3122 8317
rect 3125 8314 3127 8317
rect 3141 8315 3143 8317
rect 3157 8315 3159 8317
rect 3162 8312 3164 8317
rect 3183 8312 3185 8317
rect 3199 8315 3201 8317
rect 3215 8315 3217 8317
rect 3220 8312 3222 8317
rect 3236 8315 3238 8317
rect 3252 8315 3254 8317
rect 3257 8314 3259 8317
rect 3273 8315 3275 8317
rect 3289 8315 3291 8317
rect 3294 8312 3296 8317
rect 3315 8312 3317 8317
rect 3331 8315 3333 8317
rect 3347 8315 3349 8317
rect 3352 8312 3354 8317
rect 3368 8315 3370 8317
rect 3449 8315 3451 8317
rect 3454 8315 3456 8318
rect 3470 8315 3472 8317
rect 3486 8315 3488 8317
rect 3491 8315 3493 8318
rect 3512 8315 3514 8318
rect 3528 8315 3530 8318
rect 3544 8315 3546 8317
rect 3549 8315 3551 8318
rect 3565 8315 3567 8317
rect 3801 8315 3803 8317
rect 3806 8314 3808 8317
rect 3822 8315 3824 8317
rect 3838 8315 3840 8317
rect 3843 8312 3845 8317
rect 3864 8312 3866 8317
rect 3880 8315 3882 8317
rect 3896 8315 3898 8317
rect 3901 8312 3903 8317
rect 3917 8315 3919 8317
rect 3933 8315 3935 8317
rect 3938 8314 3940 8317
rect 3954 8315 3956 8317
rect 3970 8315 3972 8317
rect 3975 8312 3977 8317
rect 3996 8312 3998 8317
rect 4012 8315 4014 8317
rect 4028 8315 4030 8317
rect 4033 8312 4035 8317
rect 4049 8315 4051 8317
rect 4065 8315 4067 8317
rect 4070 8314 4072 8317
rect 4086 8315 4088 8317
rect 4102 8315 4104 8317
rect 4107 8312 4109 8317
rect 4128 8312 4130 8317
rect 4144 8315 4146 8317
rect 4160 8315 4162 8317
rect 4165 8312 4167 8317
rect 4181 8315 4183 8317
rect 4197 8315 4199 8317
rect 4202 8314 4204 8317
rect 4218 8315 4220 8317
rect 4234 8315 4236 8317
rect 4239 8312 4241 8317
rect 4260 8312 4262 8317
rect 4276 8315 4278 8317
rect 4292 8315 4294 8317
rect 4297 8312 4299 8317
rect 4313 8315 4315 8317
rect 2504 8302 2506 8307
rect 2509 8305 2511 8307
rect 2504 8288 2506 8298
rect 2509 8288 2511 8295
rect 2525 8288 2527 8307
rect 2541 8298 2543 8307
rect 2546 8305 2548 8307
rect 2567 8305 2569 8307
rect 2583 8304 2585 8307
rect 2541 8288 2543 8291
rect 2546 8288 2548 8290
rect 2567 8288 2569 8290
rect 2583 8288 2585 8300
rect 2599 8298 2601 8307
rect 2604 8305 2606 8307
rect 2599 8288 2601 8291
rect 2604 8288 2606 8290
rect 2620 8288 2622 8307
rect 3449 8302 3451 8307
rect 3454 8305 3456 8307
rect 3449 8288 3451 8298
rect 3454 8288 3456 8295
rect 3470 8288 3472 8307
rect 3486 8298 3488 8307
rect 3491 8305 3493 8307
rect 3512 8305 3514 8307
rect 3528 8304 3530 8307
rect 3486 8288 3488 8291
rect 3491 8288 3493 8290
rect 3512 8288 3514 8290
rect 3528 8288 3530 8300
rect 3544 8298 3546 8307
rect 3549 8305 3551 8307
rect 3544 8288 3546 8291
rect 3549 8288 3551 8290
rect 3565 8288 3567 8307
rect 2504 8282 2506 8284
rect 2509 8281 2511 8284
rect 2525 8282 2527 8284
rect 2541 8282 2543 8284
rect 2546 8279 2548 8284
rect 2567 8279 2569 8284
rect 2583 8282 2585 8284
rect 2599 8282 2601 8284
rect 2604 8279 2606 8284
rect 2620 8282 2622 8284
rect 3449 8282 3451 8284
rect 3454 8281 3456 8284
rect 3470 8282 3472 8284
rect 3486 8282 3488 8284
rect 3035 8277 3037 8279
rect 2877 8271 2879 8274
rect 2921 8271 2923 8274
rect 2947 8271 2949 8274
rect 2993 8271 2995 8274
rect 2947 8267 2948 8271
rect 3061 8271 3063 8275
rect 3089 8277 3091 8279
rect 3116 8277 3118 8279
rect 3066 8271 3068 8274
rect 2861 8264 2863 8266
rect 2877 8264 2879 8267
rect 2893 8264 2895 8266
rect 2916 8264 2918 8266
rect 2921 8264 2923 8267
rect 2947 8264 2949 8267
rect 2968 8264 2970 8267
rect 2988 8264 2990 8266
rect 2993 8264 2995 8267
rect 3011 8264 3013 8266
rect 2628 8251 2630 8254
rect 2628 8245 2630 8247
rect 2511 8242 2513 8245
rect 2861 8242 2863 8256
rect 2877 8254 2879 8256
rect 2877 8242 2879 8244
rect 2893 8242 2895 8256
rect 2916 8251 2918 8256
rect 2921 8254 2923 8256
rect 2947 8254 2949 8256
rect 2912 8247 2918 8251
rect 2916 8242 2918 8247
rect 2921 8242 2923 8244
rect 2947 8242 2949 8244
rect 2968 8242 2970 8256
rect 2988 8251 2990 8256
rect 2993 8254 2995 8256
rect 2984 8247 2990 8251
rect 2988 8242 2990 8247
rect 2993 8242 2995 8244
rect 3011 8242 3013 8256
rect 3035 8255 3037 8269
rect 3142 8271 3144 8275
rect 3170 8277 3172 8279
rect 3491 8279 3493 8284
rect 3512 8279 3514 8284
rect 3528 8282 3530 8284
rect 3544 8282 3546 8284
rect 3549 8279 3551 8284
rect 3565 8282 3567 8284
rect 3147 8271 3149 8274
rect 3061 8260 3063 8263
rect 3066 8261 3068 8263
rect 3062 8256 3063 8260
rect 3061 8251 3063 8256
rect 3066 8251 3068 8253
rect 3035 8249 3037 8251
rect 3089 8247 3091 8269
rect 3116 8255 3118 8269
rect 3980 8277 3982 8279
rect 3142 8260 3144 8263
rect 3147 8261 3149 8263
rect 3143 8256 3144 8260
rect 3142 8251 3144 8256
rect 3147 8251 3149 8253
rect 3116 8249 3118 8251
rect 3170 8247 3172 8269
rect 3822 8271 3824 8274
rect 3866 8271 3868 8274
rect 3892 8271 3894 8274
rect 3938 8271 3940 8274
rect 3892 8267 3893 8271
rect 4006 8271 4008 8275
rect 4034 8277 4036 8279
rect 4061 8277 4063 8279
rect 4011 8271 4013 8274
rect 3806 8264 3808 8266
rect 3822 8264 3824 8267
rect 3838 8264 3840 8266
rect 3861 8264 3863 8266
rect 3866 8264 3868 8267
rect 3892 8264 3894 8267
rect 3913 8264 3915 8267
rect 3933 8264 3935 8266
rect 3938 8264 3940 8267
rect 3956 8264 3958 8266
rect 3573 8251 3575 8254
rect 3061 8245 3063 8247
rect 3066 8242 3068 8247
rect 3142 8245 3144 8247
rect 3089 8241 3091 8243
rect 3147 8242 3149 8247
rect 3573 8245 3575 8247
rect 3170 8241 3172 8243
rect 3456 8242 3458 8245
rect 3806 8242 3808 8256
rect 3822 8254 3824 8256
rect 3822 8242 3824 8244
rect 3838 8242 3840 8256
rect 3861 8251 3863 8256
rect 3866 8254 3868 8256
rect 3892 8254 3894 8256
rect 3857 8247 3863 8251
rect 3861 8242 3863 8247
rect 3866 8242 3868 8244
rect 3892 8242 3894 8244
rect 3913 8242 3915 8256
rect 3933 8251 3935 8256
rect 3938 8254 3940 8256
rect 3929 8247 3935 8251
rect 3933 8242 3935 8247
rect 3938 8242 3940 8244
rect 3956 8242 3958 8256
rect 3980 8255 3982 8269
rect 4087 8271 4089 8275
rect 4115 8277 4117 8279
rect 4092 8271 4094 8274
rect 4006 8260 4008 8263
rect 4011 8261 4013 8263
rect 4007 8256 4008 8260
rect 4006 8251 4008 8256
rect 4011 8251 4013 8253
rect 3980 8249 3982 8251
rect 4034 8247 4036 8269
rect 4061 8255 4063 8269
rect 4087 8260 4089 8263
rect 4092 8261 4094 8263
rect 4088 8256 4089 8260
rect 4087 8251 4089 8256
rect 4092 8251 4094 8253
rect 4061 8249 4063 8251
rect 4115 8247 4117 8269
rect 4006 8245 4008 8247
rect 4011 8242 4013 8247
rect 4087 8245 4089 8247
rect 4034 8241 4036 8243
rect 4092 8242 4094 8247
rect 4115 8241 4117 8243
rect 2511 8236 2513 8238
rect 2861 8236 2863 8238
rect 2877 8234 2879 8238
rect 2893 8236 2895 8238
rect 2916 8236 2918 8238
rect 2878 8230 2879 8234
rect 2921 8233 2923 8238
rect 2947 8234 2949 8238
rect 2968 8236 2970 8238
rect 2988 8236 2990 8238
rect 2877 8227 2879 8230
rect 2922 8229 2923 8233
rect 2948 8230 2949 8234
rect 2993 8233 2995 8238
rect 3011 8236 3013 8238
rect 3456 8236 3458 8238
rect 3806 8236 3808 8238
rect 3822 8234 3824 8238
rect 3838 8236 3840 8238
rect 3861 8236 3863 8238
rect 2921 8227 2923 8229
rect 2947 8226 2949 8230
rect 2994 8229 2995 8233
rect 3823 8230 3824 8234
rect 3866 8233 3868 8238
rect 3892 8234 3894 8238
rect 3913 8236 3915 8238
rect 3933 8236 3935 8238
rect 2993 8227 2995 8229
rect 3822 8227 3824 8230
rect 3867 8229 3868 8233
rect 3893 8230 3894 8234
rect 3938 8233 3940 8238
rect 3956 8236 3958 8238
rect 3866 8227 3868 8229
rect 3892 8226 3894 8230
rect 3939 8229 3940 8233
rect 3938 8227 3940 8229
rect 2495 8213 2497 8215
rect 2511 8213 2513 8216
rect 2516 8213 2518 8215
rect 2532 8213 2534 8216
rect 2548 8213 2550 8216
rect 2569 8213 2571 8216
rect 2574 8213 2576 8215
rect 2590 8213 2592 8215
rect 2606 8213 2608 8216
rect 2611 8213 2613 8215
rect 3440 8213 3442 8215
rect 3456 8213 3458 8216
rect 3461 8213 3463 8215
rect 3477 8213 3479 8216
rect 3493 8213 3495 8216
rect 3514 8213 3516 8216
rect 3519 8213 3521 8215
rect 3535 8213 3537 8215
rect 3551 8213 3553 8216
rect 3556 8213 3558 8215
rect 2495 8186 2497 8205
rect 2511 8203 2513 8205
rect 2516 8196 2518 8205
rect 2532 8202 2534 8205
rect 2548 8203 2550 8205
rect 2569 8203 2571 8205
rect 2511 8186 2513 8188
rect 2516 8186 2518 8189
rect 2532 8186 2534 8198
rect 2574 8196 2576 8205
rect 2548 8186 2550 8188
rect 2569 8186 2571 8188
rect 2574 8186 2576 8189
rect 2590 8186 2592 8205
rect 2606 8203 2608 8205
rect 2611 8200 2613 8205
rect 2877 8204 2879 8207
rect 2921 8205 2923 8207
rect 2878 8200 2879 8204
rect 2922 8201 2923 8205
rect 2947 8204 2949 8208
rect 2993 8205 2995 8207
rect 2861 8196 2863 8198
rect 2877 8196 2879 8200
rect 2893 8196 2895 8198
rect 2916 8196 2918 8198
rect 2921 8196 2923 8201
rect 2948 8200 2949 8204
rect 2994 8201 2995 8205
rect 2947 8196 2949 8200
rect 2968 8196 2970 8198
rect 2988 8196 2990 8198
rect 2993 8196 2995 8201
rect 3011 8196 3013 8198
rect 2606 8186 2608 8193
rect 2611 8186 2613 8196
rect 3061 8195 3063 8198
rect 3066 8195 3068 8198
rect 3142 8195 3144 8198
rect 3147 8195 3149 8198
rect 2495 8180 2497 8182
rect 2511 8177 2513 8182
rect 2516 8180 2518 8182
rect 2532 8180 2534 8182
rect 2548 8177 2550 8182
rect 2569 8177 2571 8182
rect 2574 8180 2576 8182
rect 2590 8180 2592 8182
rect 2606 8179 2608 8182
rect 2611 8180 2613 8182
rect 2861 8178 2863 8192
rect 2877 8190 2879 8192
rect 2877 8178 2879 8180
rect 2893 8178 2895 8192
rect 2916 8187 2918 8192
rect 2921 8190 2923 8192
rect 2947 8190 2949 8192
rect 2912 8183 2918 8187
rect 2916 8178 2918 8183
rect 2921 8178 2923 8180
rect 2947 8178 2949 8180
rect 2968 8178 2970 8192
rect 2988 8187 2990 8192
rect 2993 8190 2995 8192
rect 2984 8183 2990 8187
rect 2988 8178 2990 8183
rect 2993 8178 2995 8180
rect 3011 8178 3013 8192
rect 3061 8179 3063 8191
rect 3066 8189 3068 8191
rect 3066 8179 3068 8181
rect 3142 8179 3144 8191
rect 3147 8189 3149 8191
rect 3440 8186 3442 8205
rect 3456 8203 3458 8205
rect 3461 8196 3463 8205
rect 3477 8202 3479 8205
rect 3493 8203 3495 8205
rect 3514 8203 3516 8205
rect 3456 8186 3458 8188
rect 3461 8186 3463 8189
rect 3477 8186 3479 8198
rect 3519 8196 3521 8205
rect 3493 8186 3495 8188
rect 3514 8186 3516 8188
rect 3519 8186 3521 8189
rect 3535 8186 3537 8205
rect 3551 8203 3553 8205
rect 3556 8200 3558 8205
rect 3822 8204 3824 8207
rect 3866 8205 3868 8207
rect 3823 8200 3824 8204
rect 3867 8201 3868 8205
rect 3892 8204 3894 8208
rect 3938 8205 3940 8207
rect 3806 8196 3808 8198
rect 3822 8196 3824 8200
rect 3838 8196 3840 8198
rect 3861 8196 3863 8198
rect 3866 8196 3868 8201
rect 3893 8200 3894 8204
rect 3939 8201 3940 8205
rect 3892 8196 3894 8200
rect 3913 8196 3915 8198
rect 3933 8196 3935 8198
rect 3938 8196 3940 8201
rect 3956 8196 3958 8198
rect 3551 8186 3553 8193
rect 3556 8186 3558 8196
rect 4006 8195 4008 8198
rect 4011 8195 4013 8198
rect 4087 8195 4089 8198
rect 4092 8195 4094 8198
rect 3147 8179 3149 8181
rect 3440 8180 3442 8182
rect 3456 8177 3458 8182
rect 3461 8180 3463 8182
rect 3477 8180 3479 8182
rect 3493 8177 3495 8182
rect 3514 8177 3516 8182
rect 3519 8180 3521 8182
rect 3535 8180 3537 8182
rect 3551 8179 3553 8182
rect 3556 8180 3558 8182
rect 3806 8178 3808 8192
rect 3822 8190 3824 8192
rect 3822 8178 3824 8180
rect 3838 8178 3840 8192
rect 3861 8187 3863 8192
rect 3866 8190 3868 8192
rect 3892 8190 3894 8192
rect 3857 8183 3863 8187
rect 3861 8178 3863 8183
rect 3866 8178 3868 8180
rect 3892 8178 3894 8180
rect 3913 8178 3915 8192
rect 3933 8187 3935 8192
rect 3938 8190 3940 8192
rect 3929 8183 3935 8187
rect 3933 8178 3935 8183
rect 3938 8178 3940 8180
rect 3956 8178 3958 8192
rect 4006 8179 4008 8191
rect 4011 8189 4013 8191
rect 4011 8179 4013 8181
rect 4087 8179 4089 8191
rect 4092 8189 4094 8191
rect 4092 8179 4094 8181
rect 2861 8168 2863 8170
rect 2877 8167 2879 8170
rect 2893 8168 2895 8170
rect 2916 8168 2918 8170
rect 2921 8167 2923 8170
rect 2947 8167 2949 8170
rect 2968 8167 2970 8170
rect 2988 8168 2990 8170
rect 2993 8167 2995 8170
rect 3011 8168 3013 8170
rect 3061 8169 3063 8171
rect 2947 8163 2948 8167
rect 3066 8166 3068 8171
rect 3142 8169 3144 8171
rect 3147 8166 3149 8171
rect 3806 8168 3808 8170
rect 3822 8167 3824 8170
rect 3838 8168 3840 8170
rect 3861 8168 3863 8170
rect 3866 8167 3868 8170
rect 3892 8167 3894 8170
rect 3913 8167 3915 8170
rect 3933 8168 3935 8170
rect 3938 8167 3940 8170
rect 3956 8168 3958 8170
rect 4006 8169 4008 8171
rect 2877 8160 2879 8163
rect 2921 8160 2923 8163
rect 2947 8160 2949 8163
rect 2993 8160 2995 8163
rect 3892 8163 3893 8167
rect 4011 8166 4013 8171
rect 4087 8169 4089 8171
rect 4092 8166 4094 8171
rect 3822 8160 3824 8163
rect 3866 8160 3868 8163
rect 3892 8160 3894 8163
rect 3938 8160 3940 8163
rect 2877 8139 2879 8142
rect 2921 8139 2923 8142
rect 2947 8139 2949 8142
rect 2993 8139 2995 8142
rect 3061 8139 3063 8143
rect 3089 8145 3091 8147
rect 3140 8145 3142 8147
rect 3066 8139 3068 8142
rect 2947 8135 2948 8139
rect 2861 8132 2863 8134
rect 2877 8132 2879 8135
rect 2893 8132 2895 8134
rect 2916 8132 2918 8134
rect 2921 8132 2923 8135
rect 2947 8132 2949 8135
rect 2968 8132 2970 8135
rect 2988 8132 2990 8134
rect 2993 8132 2995 8135
rect 3011 8132 3013 8134
rect 3166 8139 3168 8143
rect 3194 8145 3196 8147
rect 3171 8139 3173 8142
rect 3061 8128 3063 8131
rect 3066 8129 3068 8131
rect 3062 8124 3063 8128
rect 2861 8110 2863 8124
rect 2877 8122 2879 8124
rect 2877 8110 2879 8112
rect 2893 8110 2895 8124
rect 2916 8119 2918 8124
rect 2921 8122 2923 8124
rect 2947 8122 2949 8124
rect 2912 8115 2918 8119
rect 2916 8110 2918 8115
rect 2921 8110 2923 8112
rect 2947 8110 2949 8112
rect 2968 8110 2970 8124
rect 2988 8119 2990 8124
rect 2993 8122 2995 8124
rect 2984 8115 2990 8119
rect 2988 8110 2990 8115
rect 2993 8110 2995 8112
rect 3011 8110 3013 8124
rect 3061 8119 3063 8124
rect 3066 8119 3068 8121
rect 3089 8115 3091 8137
rect 3140 8123 3142 8137
rect 3822 8139 3824 8142
rect 3866 8139 3868 8142
rect 3892 8139 3894 8142
rect 3938 8139 3940 8142
rect 4006 8139 4008 8143
rect 4034 8145 4036 8147
rect 4085 8145 4087 8147
rect 4011 8139 4013 8142
rect 3166 8128 3168 8131
rect 3171 8129 3173 8131
rect 3167 8124 3168 8128
rect 3166 8119 3168 8124
rect 3171 8119 3173 8121
rect 3140 8117 3142 8119
rect 3194 8115 3196 8137
rect 3892 8135 3893 8139
rect 3806 8132 3808 8134
rect 3822 8132 3824 8135
rect 3838 8132 3840 8134
rect 3861 8132 3863 8134
rect 3866 8132 3868 8135
rect 3892 8132 3894 8135
rect 3913 8132 3915 8135
rect 3933 8132 3935 8134
rect 3938 8132 3940 8135
rect 3956 8132 3958 8134
rect 4111 8139 4113 8143
rect 4139 8145 4141 8147
rect 4116 8139 4118 8142
rect 4006 8128 4008 8131
rect 4011 8129 4013 8131
rect 4007 8124 4008 8128
rect 3061 8113 3063 8115
rect 3066 8110 3068 8115
rect 3166 8113 3168 8115
rect 3089 8109 3091 8111
rect 3171 8110 3173 8115
rect 3194 8109 3196 8111
rect 3806 8110 3808 8124
rect 3822 8122 3824 8124
rect 3822 8110 3824 8112
rect 3838 8110 3840 8124
rect 3861 8119 3863 8124
rect 3866 8122 3868 8124
rect 3892 8122 3894 8124
rect 3857 8115 3863 8119
rect 3861 8110 3863 8115
rect 3866 8110 3868 8112
rect 3892 8110 3894 8112
rect 3913 8110 3915 8124
rect 3933 8119 3935 8124
rect 3938 8122 3940 8124
rect 3929 8115 3935 8119
rect 3933 8110 3935 8115
rect 3938 8110 3940 8112
rect 3956 8110 3958 8124
rect 4006 8119 4008 8124
rect 4011 8119 4013 8121
rect 4034 8115 4036 8137
rect 4085 8123 4087 8137
rect 4111 8128 4113 8131
rect 4116 8129 4118 8131
rect 4112 8124 4113 8128
rect 4111 8119 4113 8124
rect 4116 8119 4118 8121
rect 4085 8117 4087 8119
rect 4139 8115 4141 8137
rect 4006 8113 4008 8115
rect 4011 8110 4013 8115
rect 4111 8113 4113 8115
rect 4034 8109 4036 8111
rect 4116 8110 4118 8115
rect 4139 8109 4141 8111
rect 2861 8104 2863 8106
rect 2877 8102 2879 8106
rect 2893 8104 2895 8106
rect 2916 8104 2918 8106
rect 2878 8098 2879 8102
rect 2921 8101 2923 8106
rect 2947 8102 2949 8106
rect 2968 8104 2970 8106
rect 2988 8104 2990 8106
rect 2877 8095 2879 8098
rect 2922 8097 2923 8101
rect 2948 8098 2949 8102
rect 2993 8101 2995 8106
rect 3011 8104 3013 8106
rect 3806 8104 3808 8106
rect 3822 8102 3824 8106
rect 3838 8104 3840 8106
rect 3861 8104 3863 8106
rect 2921 8095 2923 8097
rect 2947 8094 2949 8098
rect 2994 8097 2995 8101
rect 3823 8098 3824 8102
rect 3866 8101 3868 8106
rect 3892 8102 3894 8106
rect 3913 8104 3915 8106
rect 3933 8104 3935 8106
rect 2993 8095 2995 8097
rect 3822 8095 3824 8098
rect 3867 8097 3868 8101
rect 3893 8098 3894 8102
rect 3938 8101 3940 8106
rect 3956 8104 3958 8106
rect 3866 8095 3868 8097
rect 3892 8094 3894 8098
rect 3939 8097 3940 8101
rect 3938 8095 3940 8097
rect 2877 8072 2879 8075
rect 2921 8073 2923 8075
rect 2878 8068 2879 8072
rect 2922 8069 2923 8073
rect 2947 8072 2949 8076
rect 2993 8073 2995 8075
rect 2861 8064 2863 8066
rect 2877 8064 2879 8068
rect 2893 8064 2895 8066
rect 2916 8064 2918 8066
rect 2921 8064 2923 8069
rect 2948 8068 2949 8072
rect 2994 8069 2995 8073
rect 3822 8072 3824 8075
rect 3866 8073 3868 8075
rect 2947 8064 2949 8068
rect 2968 8064 2970 8066
rect 2988 8064 2990 8066
rect 2993 8064 2995 8069
rect 3823 8068 3824 8072
rect 3867 8069 3868 8073
rect 3892 8072 3894 8076
rect 3938 8073 3940 8075
rect 3011 8064 3013 8066
rect 3061 8064 3063 8067
rect 3066 8064 3068 8067
rect 3166 8064 3168 8067
rect 3171 8064 3173 8067
rect 3806 8064 3808 8066
rect 3822 8064 3824 8068
rect 3838 8064 3840 8066
rect 3861 8064 3863 8066
rect 3866 8064 3868 8069
rect 3893 8068 3894 8072
rect 3939 8069 3940 8073
rect 3892 8064 3894 8068
rect 3913 8064 3915 8066
rect 3933 8064 3935 8066
rect 3938 8064 3940 8069
rect 3956 8064 3958 8066
rect 4006 8064 4008 8067
rect 4011 8064 4013 8067
rect 4111 8064 4113 8067
rect 4116 8064 4118 8067
rect 2861 8046 2863 8060
rect 2877 8058 2879 8060
rect 2877 8046 2879 8048
rect 2893 8046 2895 8060
rect 2916 8055 2918 8060
rect 2921 8058 2923 8060
rect 2947 8058 2949 8060
rect 2912 8051 2918 8055
rect 2916 8046 2918 8051
rect 2921 8046 2923 8048
rect 2947 8046 2949 8048
rect 2968 8046 2970 8060
rect 2988 8055 2990 8060
rect 2993 8058 2995 8060
rect 2984 8051 2990 8055
rect 2988 8046 2990 8051
rect 2993 8046 2995 8048
rect 3011 8046 3013 8060
rect 3061 8048 3063 8060
rect 3066 8058 3068 8060
rect 3066 8048 3068 8050
rect 3166 8048 3168 8060
rect 3171 8058 3173 8060
rect 3171 8048 3173 8050
rect 3806 8046 3808 8060
rect 3822 8058 3824 8060
rect 3822 8046 3824 8048
rect 3838 8046 3840 8060
rect 3861 8055 3863 8060
rect 3866 8058 3868 8060
rect 3892 8058 3894 8060
rect 3857 8051 3863 8055
rect 3861 8046 3863 8051
rect 3866 8046 3868 8048
rect 3892 8046 3894 8048
rect 3913 8046 3915 8060
rect 3933 8055 3935 8060
rect 3938 8058 3940 8060
rect 3929 8051 3935 8055
rect 3933 8046 3935 8051
rect 3938 8046 3940 8048
rect 3956 8046 3958 8060
rect 4006 8048 4008 8060
rect 4011 8058 4013 8060
rect 4011 8048 4013 8050
rect 4111 8048 4113 8060
rect 4116 8058 4118 8060
rect 4116 8048 4118 8050
rect 3061 8038 3063 8040
rect 2861 8036 2863 8038
rect 2877 8035 2879 8038
rect 2893 8036 2895 8038
rect 2916 8036 2918 8038
rect 2921 8035 2923 8038
rect 2947 8035 2949 8038
rect 2968 8035 2970 8038
rect 2988 8036 2990 8038
rect 2993 8035 2995 8038
rect 3011 8036 3013 8038
rect 3066 8035 3068 8040
rect 3166 8038 3168 8040
rect 3171 8035 3173 8040
rect 4006 8038 4008 8040
rect 3806 8036 3808 8038
rect 2947 8031 2948 8035
rect 3822 8035 3824 8038
rect 3838 8036 3840 8038
rect 3861 8036 3863 8038
rect 3866 8035 3868 8038
rect 3892 8035 3894 8038
rect 3913 8035 3915 8038
rect 3933 8036 3935 8038
rect 3938 8035 3940 8038
rect 3956 8036 3958 8038
rect 4011 8035 4013 8040
rect 4111 8038 4113 8040
rect 4116 8035 4118 8040
rect 3892 8031 3893 8035
rect 2877 8028 2879 8031
rect 2921 8028 2923 8031
rect 2947 8028 2949 8031
rect 2993 8028 2995 8031
rect 3822 8028 3824 8031
rect 3866 8028 3868 8031
rect 3892 8028 3894 8031
rect 3938 8028 3940 8031
rect 2877 8007 2879 8010
rect 2921 8007 2923 8010
rect 2947 8007 2949 8010
rect 2993 8007 2995 8010
rect 3061 8007 3063 8011
rect 3089 8013 3091 8015
rect 3116 8013 3118 8015
rect 3066 8007 3068 8010
rect 2947 8003 2948 8007
rect 2861 8000 2863 8002
rect 2877 8000 2879 8003
rect 2893 8000 2895 8002
rect 2916 8000 2918 8002
rect 2921 8000 2923 8003
rect 2947 8000 2949 8003
rect 2968 8000 2970 8003
rect 2988 8000 2990 8002
rect 2993 8000 2995 8003
rect 3011 8000 3013 8002
rect 3142 8007 3144 8011
rect 3170 8013 3172 8015
rect 3206 8013 3208 8015
rect 3147 8007 3149 8010
rect 3061 7996 3063 7999
rect 3066 7997 3068 7999
rect 3062 7992 3063 7996
rect 2861 7978 2863 7992
rect 2877 7990 2879 7992
rect 2877 7978 2879 7980
rect 2893 7978 2895 7992
rect 2916 7987 2918 7992
rect 2921 7990 2923 7992
rect 2947 7990 2949 7992
rect 2912 7983 2918 7987
rect 2916 7978 2918 7983
rect 2921 7978 2923 7980
rect 2947 7978 2949 7980
rect 2968 7978 2970 7992
rect 2988 7987 2990 7992
rect 2993 7990 2995 7992
rect 2984 7983 2990 7987
rect 2988 7978 2990 7983
rect 2993 7978 2995 7980
rect 3011 7978 3013 7992
rect 3061 7987 3063 7992
rect 3066 7987 3068 7989
rect 3089 7983 3091 8005
rect 3116 7991 3118 8005
rect 3232 8007 3234 8011
rect 3260 8013 3262 8015
rect 3237 8007 3239 8010
rect 3142 7996 3144 7999
rect 3147 7997 3149 7999
rect 3143 7992 3144 7996
rect 3142 7987 3144 7992
rect 3147 7987 3149 7989
rect 3116 7985 3118 7987
rect 3170 7983 3172 8005
rect 3206 7991 3208 8005
rect 3822 8007 3824 8010
rect 3866 8007 3868 8010
rect 3892 8007 3894 8010
rect 3938 8007 3940 8010
rect 4006 8007 4008 8011
rect 4034 8013 4036 8015
rect 4061 8013 4063 8015
rect 4011 8007 4013 8010
rect 3232 7996 3234 7999
rect 3237 7997 3239 7999
rect 3233 7992 3234 7996
rect 3232 7987 3234 7992
rect 3237 7987 3239 7989
rect 3206 7985 3208 7987
rect 3260 7983 3262 8005
rect 3892 8003 3893 8007
rect 3806 8000 3808 8002
rect 3822 8000 3824 8003
rect 3838 8000 3840 8002
rect 3861 8000 3863 8002
rect 3866 8000 3868 8003
rect 3892 8000 3894 8003
rect 3913 8000 3915 8003
rect 3933 8000 3935 8002
rect 3938 8000 3940 8003
rect 3956 8000 3958 8002
rect 4087 8007 4089 8011
rect 4115 8013 4117 8015
rect 4151 8013 4153 8015
rect 4092 8007 4094 8010
rect 4006 7996 4008 7999
rect 4011 7997 4013 7999
rect 4007 7992 4008 7996
rect 3061 7981 3063 7983
rect 3066 7978 3068 7983
rect 3142 7981 3144 7983
rect 3089 7977 3091 7979
rect 3147 7978 3149 7983
rect 3232 7981 3234 7983
rect 3170 7977 3172 7979
rect 3237 7978 3239 7983
rect 3260 7977 3262 7979
rect 3806 7978 3808 7992
rect 3822 7990 3824 7992
rect 3822 7978 3824 7980
rect 3838 7978 3840 7992
rect 3861 7987 3863 7992
rect 3866 7990 3868 7992
rect 3892 7990 3894 7992
rect 3857 7983 3863 7987
rect 3861 7978 3863 7983
rect 3866 7978 3868 7980
rect 3892 7978 3894 7980
rect 3913 7978 3915 7992
rect 3933 7987 3935 7992
rect 3938 7990 3940 7992
rect 3929 7983 3935 7987
rect 3933 7978 3935 7983
rect 3938 7978 3940 7980
rect 3956 7978 3958 7992
rect 4006 7987 4008 7992
rect 4011 7987 4013 7989
rect 4034 7983 4036 8005
rect 4061 7991 4063 8005
rect 4177 8007 4179 8011
rect 4205 8013 4207 8015
rect 4182 8007 4184 8010
rect 4087 7996 4089 7999
rect 4092 7997 4094 7999
rect 4088 7992 4089 7996
rect 4087 7987 4089 7992
rect 4092 7987 4094 7989
rect 4061 7985 4063 7987
rect 4115 7983 4117 8005
rect 4151 7991 4153 8005
rect 4177 7996 4179 7999
rect 4182 7997 4184 7999
rect 4178 7992 4179 7996
rect 4177 7987 4179 7992
rect 4182 7987 4184 7989
rect 4151 7985 4153 7987
rect 4205 7983 4207 8005
rect 4006 7981 4008 7983
rect 4011 7978 4013 7983
rect 4087 7981 4089 7983
rect 4034 7977 4036 7979
rect 4092 7978 4094 7983
rect 4177 7981 4179 7983
rect 4115 7977 4117 7979
rect 4182 7978 4184 7983
rect 4205 7977 4207 7979
rect 2861 7972 2863 7974
rect 2877 7970 2879 7974
rect 2893 7972 2895 7974
rect 2916 7972 2918 7974
rect 2878 7966 2879 7970
rect 2921 7969 2923 7974
rect 2947 7970 2949 7974
rect 2968 7972 2970 7974
rect 2988 7972 2990 7974
rect 2877 7963 2879 7966
rect 2922 7965 2923 7969
rect 2948 7966 2949 7970
rect 2993 7969 2995 7974
rect 3011 7972 3013 7974
rect 3806 7972 3808 7974
rect 3822 7970 3824 7974
rect 3838 7972 3840 7974
rect 3861 7972 3863 7974
rect 2921 7963 2923 7965
rect 2947 7962 2949 7966
rect 2994 7965 2995 7969
rect 3823 7966 3824 7970
rect 3866 7969 3868 7974
rect 3892 7970 3894 7974
rect 3913 7972 3915 7974
rect 3933 7972 3935 7974
rect 2993 7963 2995 7965
rect 3822 7963 3824 7966
rect 3867 7965 3868 7969
rect 3893 7966 3894 7970
rect 3938 7969 3940 7974
rect 3956 7972 3958 7974
rect 3866 7963 3868 7965
rect 3892 7962 3894 7966
rect 3939 7965 3940 7969
rect 3938 7963 3940 7965
rect 2877 7940 2879 7943
rect 2921 7941 2923 7943
rect 2878 7936 2879 7940
rect 2922 7937 2923 7941
rect 2947 7940 2949 7944
rect 2993 7941 2995 7943
rect 2861 7932 2863 7934
rect 2877 7932 2879 7936
rect 2893 7932 2895 7934
rect 2916 7932 2918 7934
rect 2921 7932 2923 7937
rect 2948 7936 2949 7940
rect 2994 7937 2995 7941
rect 3822 7940 3824 7943
rect 3866 7941 3868 7943
rect 2947 7932 2949 7936
rect 2968 7932 2970 7934
rect 2988 7932 2990 7934
rect 2993 7932 2995 7937
rect 3823 7936 3824 7940
rect 3867 7937 3868 7941
rect 3892 7940 3894 7944
rect 3938 7941 3940 7943
rect 3011 7932 3013 7934
rect 3806 7932 3808 7934
rect 3822 7932 3824 7936
rect 3838 7932 3840 7934
rect 3861 7932 3863 7934
rect 3866 7932 3868 7937
rect 3893 7936 3894 7940
rect 3939 7937 3940 7941
rect 3892 7932 3894 7936
rect 3913 7932 3915 7934
rect 3933 7932 3935 7934
rect 3938 7932 3940 7937
rect 3956 7932 3958 7934
rect 3061 7929 3063 7932
rect 3066 7929 3068 7932
rect 3142 7929 3144 7932
rect 3147 7929 3149 7932
rect 3232 7929 3234 7932
rect 3237 7929 3239 7932
rect 2861 7914 2863 7928
rect 2877 7926 2879 7928
rect 2877 7914 2879 7916
rect 2893 7914 2895 7928
rect 2916 7923 2918 7928
rect 2921 7926 2923 7928
rect 2947 7926 2949 7928
rect 2912 7919 2918 7923
rect 2916 7914 2918 7919
rect 2921 7914 2923 7916
rect 2947 7914 2949 7916
rect 2968 7914 2970 7928
rect 2988 7923 2990 7928
rect 2993 7926 2995 7928
rect 2984 7919 2990 7923
rect 2988 7914 2990 7919
rect 2993 7914 2995 7916
rect 3011 7914 3013 7928
rect 4006 7929 4008 7932
rect 4011 7929 4013 7932
rect 4087 7929 4089 7932
rect 4092 7929 4094 7932
rect 4177 7929 4179 7932
rect 4182 7929 4184 7932
rect 3061 7913 3063 7925
rect 3066 7923 3068 7925
rect 3066 7913 3068 7915
rect 3142 7913 3144 7925
rect 3147 7923 3149 7925
rect 3147 7913 3149 7915
rect 3232 7913 3234 7925
rect 3237 7923 3239 7925
rect 3237 7913 3239 7915
rect 3806 7914 3808 7928
rect 3822 7926 3824 7928
rect 3822 7914 3824 7916
rect 3838 7914 3840 7928
rect 3861 7923 3863 7928
rect 3866 7926 3868 7928
rect 3892 7926 3894 7928
rect 3857 7919 3863 7923
rect 3861 7914 3863 7919
rect 3866 7914 3868 7916
rect 3892 7914 3894 7916
rect 3913 7914 3915 7928
rect 3933 7923 3935 7928
rect 3938 7926 3940 7928
rect 3929 7919 3935 7923
rect 3933 7914 3935 7919
rect 3938 7914 3940 7916
rect 3956 7914 3958 7928
rect 2861 7904 2863 7906
rect 2877 7903 2879 7906
rect 2893 7904 2895 7906
rect 2916 7904 2918 7906
rect 2921 7903 2923 7906
rect 2947 7903 2949 7906
rect 2968 7903 2970 7906
rect 2988 7904 2990 7906
rect 2993 7903 2995 7906
rect 3011 7904 3013 7906
rect 4006 7913 4008 7925
rect 4011 7923 4013 7925
rect 4011 7913 4013 7915
rect 4087 7913 4089 7925
rect 4092 7923 4094 7925
rect 4092 7913 4094 7915
rect 4177 7913 4179 7925
rect 4182 7923 4184 7925
rect 4182 7913 4184 7915
rect 3061 7903 3063 7905
rect 2947 7899 2948 7903
rect 3066 7900 3068 7905
rect 3142 7903 3144 7905
rect 3147 7900 3149 7905
rect 3232 7903 3234 7905
rect 3237 7900 3239 7905
rect 3806 7904 3808 7906
rect 2877 7896 2879 7899
rect 2921 7896 2923 7899
rect 2947 7896 2949 7899
rect 2993 7896 2995 7899
rect 3822 7903 3824 7906
rect 3838 7904 3840 7906
rect 3861 7904 3863 7906
rect 3866 7903 3868 7906
rect 3892 7903 3894 7906
rect 3913 7903 3915 7906
rect 3933 7904 3935 7906
rect 3938 7903 3940 7906
rect 3956 7904 3958 7906
rect 4006 7903 4008 7905
rect 3892 7899 3893 7903
rect 4011 7900 4013 7905
rect 4087 7903 4089 7905
rect 4092 7900 4094 7905
rect 4177 7903 4179 7905
rect 4182 7900 4184 7905
rect 3822 7896 3824 7899
rect 3866 7896 3868 7899
rect 3892 7896 3894 7899
rect 3938 7896 3940 7899
rect 2877 7875 2879 7878
rect 2921 7875 2923 7878
rect 2947 7875 2949 7878
rect 2993 7875 2995 7878
rect 3061 7875 3063 7879
rect 3089 7881 3091 7883
rect 3066 7875 3068 7878
rect 2947 7871 2948 7875
rect 2861 7868 2863 7870
rect 2877 7868 2879 7871
rect 2893 7868 2895 7870
rect 2916 7868 2918 7870
rect 2921 7868 2923 7871
rect 2947 7868 2949 7871
rect 2968 7868 2970 7871
rect 2988 7868 2990 7870
rect 2993 7868 2995 7871
rect 3011 7868 3013 7870
rect 3822 7875 3824 7878
rect 3866 7875 3868 7878
rect 3892 7875 3894 7878
rect 3938 7875 3940 7878
rect 4006 7875 4008 7879
rect 4034 7881 4036 7883
rect 4011 7875 4013 7878
rect 3061 7864 3063 7867
rect 3066 7865 3068 7867
rect 3062 7860 3063 7864
rect 2861 7846 2863 7860
rect 2877 7858 2879 7860
rect 2877 7846 2879 7848
rect 2893 7846 2895 7860
rect 2916 7855 2918 7860
rect 2921 7858 2923 7860
rect 2947 7858 2949 7860
rect 2912 7851 2918 7855
rect 2916 7846 2918 7851
rect 2921 7846 2923 7848
rect 2947 7846 2949 7848
rect 2968 7846 2970 7860
rect 2988 7855 2990 7860
rect 2993 7858 2995 7860
rect 2984 7851 2990 7855
rect 2988 7846 2990 7851
rect 2993 7846 2995 7848
rect 3011 7846 3013 7860
rect 3061 7855 3063 7860
rect 3066 7855 3068 7857
rect 3089 7851 3091 7873
rect 3892 7871 3893 7875
rect 3806 7868 3808 7870
rect 3822 7868 3824 7871
rect 3838 7868 3840 7870
rect 3861 7868 3863 7870
rect 3866 7868 3868 7871
rect 3892 7868 3894 7871
rect 3913 7868 3915 7871
rect 3933 7868 3935 7870
rect 3938 7868 3940 7871
rect 3956 7868 3958 7870
rect 4006 7864 4008 7867
rect 4011 7865 4013 7867
rect 4007 7860 4008 7864
rect 3061 7849 3063 7851
rect 3066 7846 3068 7851
rect 3089 7845 3091 7847
rect 3806 7846 3808 7860
rect 3822 7858 3824 7860
rect 3822 7846 3824 7848
rect 3838 7846 3840 7860
rect 3861 7855 3863 7860
rect 3866 7858 3868 7860
rect 3892 7858 3894 7860
rect 3857 7851 3863 7855
rect 3861 7846 3863 7851
rect 3866 7846 3868 7848
rect 3892 7846 3894 7848
rect 3913 7846 3915 7860
rect 3933 7855 3935 7860
rect 3938 7858 3940 7860
rect 3929 7851 3935 7855
rect 3933 7846 3935 7851
rect 3938 7846 3940 7848
rect 3956 7846 3958 7860
rect 4006 7855 4008 7860
rect 4011 7855 4013 7857
rect 4034 7851 4036 7873
rect 4006 7849 4008 7851
rect 4011 7846 4013 7851
rect 4034 7845 4036 7847
rect 2861 7840 2863 7842
rect 2877 7838 2879 7842
rect 2893 7840 2895 7842
rect 2916 7840 2918 7842
rect 2878 7834 2879 7838
rect 2921 7837 2923 7842
rect 2947 7838 2949 7842
rect 2968 7840 2970 7842
rect 2988 7840 2990 7842
rect 2877 7831 2879 7834
rect 2922 7833 2923 7837
rect 2948 7834 2949 7838
rect 2993 7837 2995 7842
rect 3011 7840 3013 7842
rect 3806 7840 3808 7842
rect 3822 7838 3824 7842
rect 3838 7840 3840 7842
rect 3861 7840 3863 7842
rect 2921 7831 2923 7833
rect 2947 7830 2949 7834
rect 2994 7833 2995 7837
rect 3823 7834 3824 7838
rect 3866 7837 3868 7842
rect 3892 7838 3894 7842
rect 3913 7840 3915 7842
rect 3933 7840 3935 7842
rect 2993 7831 2995 7833
rect 3822 7831 3824 7834
rect 3867 7833 3868 7837
rect 3893 7834 3894 7838
rect 3938 7837 3940 7842
rect 3956 7840 3958 7842
rect 3866 7831 3868 7833
rect 3892 7830 3894 7834
rect 3939 7833 3940 7837
rect 3938 7831 3940 7833
rect 2372 7813 2374 7815
rect 2377 7813 2379 7816
rect 2393 7813 2395 7815
rect 2409 7813 2411 7815
rect 2414 7813 2416 7816
rect 2435 7813 2437 7816
rect 2451 7813 2453 7816
rect 2467 7813 2469 7815
rect 2472 7813 2474 7816
rect 2488 7813 2490 7815
rect 2504 7813 2506 7815
rect 2509 7813 2511 7816
rect 2525 7813 2527 7815
rect 2541 7813 2543 7815
rect 2546 7813 2548 7816
rect 2567 7813 2569 7816
rect 2583 7813 2585 7816
rect 2599 7813 2601 7815
rect 2604 7813 2606 7816
rect 2620 7813 2622 7815
rect 2636 7813 2638 7815
rect 2641 7813 2643 7816
rect 2657 7813 2659 7815
rect 2673 7813 2675 7815
rect 2678 7813 2680 7816
rect 2699 7813 2701 7816
rect 2715 7813 2717 7816
rect 2731 7813 2733 7815
rect 2736 7813 2738 7816
rect 2752 7813 2754 7815
rect 3317 7813 3319 7815
rect 3322 7813 3324 7816
rect 3338 7813 3340 7815
rect 3354 7813 3356 7815
rect 3359 7813 3361 7816
rect 3380 7813 3382 7816
rect 3396 7813 3398 7816
rect 3412 7813 3414 7815
rect 3417 7813 3419 7816
rect 3433 7813 3435 7815
rect 3449 7813 3451 7815
rect 3454 7813 3456 7816
rect 3470 7813 3472 7815
rect 3486 7813 3488 7815
rect 3491 7813 3493 7816
rect 3512 7813 3514 7816
rect 3528 7813 3530 7816
rect 3544 7813 3546 7815
rect 3549 7813 3551 7816
rect 3565 7813 3567 7815
rect 3581 7813 3583 7815
rect 3586 7813 3588 7816
rect 3602 7813 3604 7815
rect 3618 7813 3620 7815
rect 3623 7813 3625 7816
rect 3644 7813 3646 7816
rect 3660 7813 3662 7816
rect 3676 7813 3678 7815
rect 3681 7813 3683 7816
rect 3697 7813 3699 7815
rect 2877 7808 2879 7811
rect 2921 7809 2923 7811
rect 2372 7800 2374 7805
rect 2377 7803 2379 7805
rect 2372 7786 2374 7796
rect 2377 7786 2379 7793
rect 2393 7786 2395 7805
rect 2409 7796 2411 7805
rect 2414 7803 2416 7805
rect 2435 7803 2437 7805
rect 2451 7802 2453 7805
rect 2409 7786 2411 7789
rect 2414 7786 2416 7788
rect 2435 7786 2437 7788
rect 2451 7786 2453 7798
rect 2467 7796 2469 7805
rect 2472 7803 2474 7805
rect 2467 7786 2469 7789
rect 2472 7786 2474 7788
rect 2488 7786 2490 7805
rect 2504 7802 2506 7805
rect 2509 7803 2511 7805
rect 2504 7786 2506 7798
rect 2509 7786 2511 7793
rect 2525 7786 2527 7805
rect 2541 7796 2543 7805
rect 2546 7803 2548 7805
rect 2567 7803 2569 7805
rect 2583 7802 2585 7805
rect 2541 7786 2543 7789
rect 2546 7786 2548 7788
rect 2567 7786 2569 7788
rect 2583 7786 2585 7798
rect 2599 7796 2601 7805
rect 2604 7803 2606 7805
rect 2599 7786 2601 7789
rect 2604 7786 2606 7788
rect 2620 7786 2622 7805
rect 2636 7802 2638 7805
rect 2641 7803 2643 7805
rect 2636 7786 2638 7798
rect 2641 7786 2643 7793
rect 2657 7786 2659 7805
rect 2673 7796 2675 7805
rect 2678 7803 2680 7805
rect 2699 7803 2701 7805
rect 2715 7802 2717 7805
rect 2673 7786 2675 7789
rect 2678 7786 2680 7788
rect 2699 7786 2701 7788
rect 2715 7786 2717 7798
rect 2731 7796 2733 7805
rect 2736 7803 2738 7805
rect 2752 7797 2754 7805
rect 2878 7804 2879 7808
rect 2922 7805 2923 7809
rect 2947 7808 2949 7812
rect 2993 7809 2995 7811
rect 2861 7800 2863 7802
rect 2877 7800 2879 7804
rect 2893 7800 2895 7802
rect 2916 7800 2918 7802
rect 2921 7800 2923 7805
rect 2948 7804 2949 7808
rect 2994 7805 2995 7809
rect 3138 7808 3140 7811
rect 3182 7809 3184 7811
rect 2947 7800 2949 7804
rect 2968 7800 2970 7802
rect 2988 7800 2990 7802
rect 2993 7800 2995 7805
rect 3139 7804 3140 7808
rect 3183 7805 3184 7809
rect 3208 7808 3210 7812
rect 3254 7809 3256 7811
rect 3011 7800 3013 7802
rect 3095 7800 3097 7803
rect 3113 7800 3115 7803
rect 3138 7800 3140 7804
rect 3154 7800 3156 7802
rect 3177 7800 3179 7802
rect 3182 7800 3184 7805
rect 3209 7804 3210 7808
rect 3255 7805 3256 7809
rect 3822 7808 3824 7811
rect 3866 7809 3868 7811
rect 3208 7800 3210 7804
rect 3229 7800 3231 7802
rect 3249 7800 3251 7802
rect 3254 7800 3256 7805
rect 3272 7800 3274 7802
rect 3317 7800 3319 7805
rect 3322 7803 3324 7805
rect 2731 7786 2733 7789
rect 2736 7786 2738 7788
rect 2752 7786 2754 7793
rect 2861 7782 2863 7796
rect 2877 7794 2879 7796
rect 2877 7782 2879 7784
rect 2893 7782 2895 7796
rect 2916 7791 2918 7796
rect 2921 7794 2923 7796
rect 2947 7794 2949 7796
rect 2912 7787 2918 7791
rect 2916 7782 2918 7787
rect 2921 7782 2923 7784
rect 2947 7782 2949 7784
rect 2968 7782 2970 7796
rect 2988 7791 2990 7796
rect 2993 7794 2995 7796
rect 2984 7787 2990 7791
rect 2988 7782 2990 7787
rect 2993 7782 2995 7784
rect 3011 7782 3013 7796
rect 3061 7793 3063 7796
rect 3066 7793 3068 7796
rect 3095 7791 3097 7796
rect 2372 7780 2374 7782
rect 2377 7779 2379 7782
rect 2393 7780 2395 7782
rect 2409 7780 2411 7782
rect 2414 7777 2416 7782
rect 2435 7777 2437 7782
rect 2451 7780 2453 7782
rect 2467 7780 2469 7782
rect 2472 7777 2474 7782
rect 2488 7780 2490 7782
rect 2504 7780 2506 7782
rect 2509 7779 2511 7782
rect 2525 7780 2527 7782
rect 2541 7780 2543 7782
rect 2546 7777 2548 7782
rect 2567 7777 2569 7782
rect 2583 7780 2585 7782
rect 2599 7780 2601 7782
rect 2604 7777 2606 7782
rect 2620 7780 2622 7782
rect 2636 7780 2638 7782
rect 2641 7779 2643 7782
rect 2657 7780 2659 7782
rect 2673 7780 2675 7782
rect 2678 7777 2680 7782
rect 2699 7777 2701 7782
rect 2715 7780 2717 7782
rect 2731 7780 2733 7782
rect 2736 7777 2738 7782
rect 2752 7780 2754 7782
rect 3061 7777 3063 7789
rect 3066 7787 3068 7789
rect 3095 7782 3097 7787
rect 3113 7782 3115 7796
rect 3138 7794 3140 7796
rect 3138 7782 3140 7784
rect 3154 7782 3156 7796
rect 3177 7791 3179 7796
rect 3182 7794 3184 7796
rect 3208 7794 3210 7796
rect 3173 7787 3179 7791
rect 3177 7782 3179 7787
rect 3182 7782 3184 7784
rect 3208 7782 3210 7784
rect 3229 7782 3231 7796
rect 3249 7791 3251 7796
rect 3254 7794 3256 7796
rect 3245 7787 3251 7791
rect 3249 7782 3251 7787
rect 3254 7782 3256 7784
rect 3272 7782 3274 7796
rect 3317 7786 3319 7796
rect 3322 7786 3324 7793
rect 3338 7786 3340 7805
rect 3354 7796 3356 7805
rect 3359 7803 3361 7805
rect 3380 7803 3382 7805
rect 3396 7802 3398 7805
rect 3354 7786 3356 7789
rect 3359 7786 3361 7788
rect 3380 7786 3382 7788
rect 3396 7786 3398 7798
rect 3412 7796 3414 7805
rect 3417 7803 3419 7805
rect 3412 7786 3414 7789
rect 3417 7786 3419 7788
rect 3433 7786 3435 7805
rect 3449 7802 3451 7805
rect 3454 7803 3456 7805
rect 3449 7786 3451 7798
rect 3454 7786 3456 7793
rect 3470 7786 3472 7805
rect 3486 7796 3488 7805
rect 3491 7803 3493 7805
rect 3512 7803 3514 7805
rect 3528 7802 3530 7805
rect 3486 7786 3488 7789
rect 3491 7786 3493 7788
rect 3512 7786 3514 7788
rect 3528 7786 3530 7798
rect 3544 7796 3546 7805
rect 3549 7803 3551 7805
rect 3544 7786 3546 7789
rect 3549 7786 3551 7788
rect 3565 7786 3567 7805
rect 3581 7802 3583 7805
rect 3586 7803 3588 7805
rect 3581 7786 3583 7798
rect 3586 7786 3588 7793
rect 3602 7786 3604 7805
rect 3618 7796 3620 7805
rect 3623 7803 3625 7805
rect 3644 7803 3646 7805
rect 3660 7802 3662 7805
rect 3618 7786 3620 7789
rect 3623 7786 3625 7788
rect 3644 7786 3646 7788
rect 3660 7786 3662 7798
rect 3676 7796 3678 7805
rect 3681 7803 3683 7805
rect 3697 7797 3699 7805
rect 3823 7804 3824 7808
rect 3867 7805 3868 7809
rect 3892 7808 3894 7812
rect 3938 7809 3940 7811
rect 3806 7800 3808 7802
rect 3822 7800 3824 7804
rect 3838 7800 3840 7802
rect 3861 7800 3863 7802
rect 3866 7800 3868 7805
rect 3893 7804 3894 7808
rect 3939 7805 3940 7809
rect 4083 7808 4085 7811
rect 4127 7809 4129 7811
rect 3892 7800 3894 7804
rect 3913 7800 3915 7802
rect 3933 7800 3935 7802
rect 3938 7800 3940 7805
rect 4084 7804 4085 7808
rect 4128 7805 4129 7809
rect 4153 7808 4155 7812
rect 4199 7809 4201 7811
rect 3956 7800 3958 7802
rect 4040 7800 4042 7803
rect 4058 7800 4060 7803
rect 4083 7800 4085 7804
rect 4099 7800 4101 7802
rect 4122 7800 4124 7802
rect 4127 7800 4129 7805
rect 4154 7804 4155 7808
rect 4200 7805 4201 7809
rect 4153 7800 4155 7804
rect 4174 7800 4176 7802
rect 4194 7800 4196 7802
rect 4199 7800 4201 7805
rect 4217 7800 4219 7802
rect 3676 7786 3678 7789
rect 3681 7786 3683 7788
rect 3697 7786 3699 7793
rect 3806 7782 3808 7796
rect 3822 7794 3824 7796
rect 3822 7782 3824 7784
rect 3838 7782 3840 7796
rect 3861 7791 3863 7796
rect 3866 7794 3868 7796
rect 3892 7794 3894 7796
rect 3857 7787 3863 7791
rect 3861 7782 3863 7787
rect 3866 7782 3868 7784
rect 3892 7782 3894 7784
rect 3913 7782 3915 7796
rect 3933 7791 3935 7796
rect 3938 7794 3940 7796
rect 3929 7787 3935 7791
rect 3933 7782 3935 7787
rect 3938 7782 3940 7784
rect 3956 7782 3958 7796
rect 4006 7793 4008 7796
rect 4011 7793 4013 7796
rect 4040 7791 4042 7796
rect 3066 7777 3068 7779
rect 2861 7772 2863 7774
rect 2877 7771 2879 7774
rect 2893 7772 2895 7774
rect 2916 7772 2918 7774
rect 2921 7771 2923 7774
rect 2947 7771 2949 7774
rect 2968 7771 2970 7774
rect 2988 7772 2990 7774
rect 2993 7771 2995 7774
rect 3011 7772 3013 7774
rect 2947 7767 2948 7771
rect 3317 7780 3319 7782
rect 3322 7779 3324 7782
rect 3338 7780 3340 7782
rect 3354 7780 3356 7782
rect 3359 7777 3361 7782
rect 3380 7777 3382 7782
rect 3396 7780 3398 7782
rect 3412 7780 3414 7782
rect 3417 7777 3419 7782
rect 3433 7780 3435 7782
rect 3449 7780 3451 7782
rect 3095 7771 3097 7774
rect 3061 7767 3063 7769
rect 2877 7764 2879 7767
rect 2921 7764 2923 7767
rect 2947 7764 2949 7767
rect 2993 7764 2995 7767
rect 3066 7764 3068 7769
rect 2487 7742 2489 7745
rect 2511 7742 2513 7745
rect 2487 7736 2489 7738
rect 2511 7736 2513 7738
rect 3113 7732 3115 7774
rect 3138 7771 3140 7774
rect 3154 7772 3156 7774
rect 3177 7772 3179 7774
rect 3182 7771 3184 7774
rect 3208 7771 3210 7774
rect 3229 7771 3231 7774
rect 3249 7772 3251 7774
rect 3254 7771 3256 7774
rect 3272 7772 3274 7774
rect 3454 7779 3456 7782
rect 3470 7780 3472 7782
rect 3486 7780 3488 7782
rect 3491 7777 3493 7782
rect 3512 7777 3514 7782
rect 3528 7780 3530 7782
rect 3544 7780 3546 7782
rect 3549 7777 3551 7782
rect 3565 7780 3567 7782
rect 3581 7780 3583 7782
rect 3586 7779 3588 7782
rect 3602 7780 3604 7782
rect 3618 7780 3620 7782
rect 3623 7777 3625 7782
rect 3644 7777 3646 7782
rect 3660 7780 3662 7782
rect 3676 7780 3678 7782
rect 3681 7777 3683 7782
rect 3697 7780 3699 7782
rect 4006 7777 4008 7789
rect 4011 7787 4013 7789
rect 4040 7782 4042 7787
rect 4058 7782 4060 7796
rect 4083 7794 4085 7796
rect 4083 7782 4085 7784
rect 4099 7782 4101 7796
rect 4122 7791 4124 7796
rect 4127 7794 4129 7796
rect 4153 7794 4155 7796
rect 4118 7787 4124 7791
rect 4122 7782 4124 7787
rect 4127 7782 4129 7784
rect 4153 7782 4155 7784
rect 4174 7782 4176 7796
rect 4194 7791 4196 7796
rect 4199 7794 4201 7796
rect 4190 7787 4196 7791
rect 4194 7782 4196 7787
rect 4199 7782 4201 7784
rect 4217 7782 4219 7796
rect 4011 7777 4013 7779
rect 3806 7772 3808 7774
rect 3822 7771 3824 7774
rect 3838 7772 3840 7774
rect 3861 7772 3863 7774
rect 3866 7771 3868 7774
rect 3892 7771 3894 7774
rect 3913 7771 3915 7774
rect 3933 7772 3935 7774
rect 3938 7771 3940 7774
rect 3956 7772 3958 7774
rect 3208 7767 3209 7771
rect 3138 7764 3140 7767
rect 3182 7764 3184 7767
rect 3208 7764 3210 7767
rect 3254 7764 3256 7767
rect 3892 7767 3893 7771
rect 4040 7771 4042 7774
rect 4006 7767 4008 7769
rect 3822 7764 3824 7767
rect 3866 7764 3868 7767
rect 3892 7764 3894 7767
rect 3938 7764 3940 7767
rect 4011 7764 4013 7769
rect 3432 7742 3434 7745
rect 3456 7742 3458 7745
rect 3281 7740 3284 7742
rect 3288 7740 3291 7742
rect 3432 7736 3434 7738
rect 3456 7736 3458 7738
rect 4058 7736 4060 7774
rect 4083 7771 4085 7774
rect 4099 7772 4101 7774
rect 4122 7772 4124 7774
rect 4127 7771 4129 7774
rect 4153 7771 4155 7774
rect 4174 7771 4176 7774
rect 4194 7772 4196 7774
rect 4199 7771 4201 7774
rect 4217 7772 4219 7774
rect 4153 7767 4154 7771
rect 4083 7764 4085 7767
rect 4127 7764 4129 7767
rect 4153 7764 4155 7767
rect 4199 7764 4201 7767
rect 4226 7740 4229 7742
rect 4233 7740 4236 7742
rect 2507 7729 2509 7731
rect 3452 7729 3454 7731
rect 2507 7722 2509 7725
rect 3452 7722 3454 7725
rect 2496 7711 2498 7713
rect 2502 7711 2521 7713
rect 3441 7711 3443 7713
rect 3447 7711 3466 7713
rect 2487 7706 2489 7708
rect 2511 7706 2513 7708
rect 3432 7706 3434 7708
rect 3456 7706 3458 7708
rect 2487 7699 2489 7702
rect 2511 7699 2513 7702
rect 3155 7701 3157 7703
rect 3160 7701 3162 7704
rect 3176 7701 3178 7703
rect 3192 7701 3194 7703
rect 3197 7701 3199 7704
rect 3218 7701 3220 7704
rect 3234 7701 3236 7704
rect 3250 7701 3252 7703
rect 3255 7701 3257 7704
rect 3271 7701 3273 7703
rect 3432 7699 3434 7702
rect 3456 7699 3458 7702
rect 4100 7701 4102 7703
rect 4105 7701 4107 7704
rect 4121 7701 4123 7703
rect 4137 7701 4139 7703
rect 4142 7701 4144 7704
rect 4163 7701 4165 7704
rect 4179 7701 4181 7704
rect 4195 7701 4197 7703
rect 4200 7701 4202 7704
rect 4216 7701 4218 7703
rect 3155 7688 3157 7693
rect 3160 7691 3162 7693
rect 3155 7674 3157 7684
rect 3160 7674 3162 7681
rect 3176 7674 3178 7693
rect 3192 7684 3194 7693
rect 3197 7691 3199 7693
rect 3218 7691 3220 7693
rect 3234 7690 3236 7693
rect 3192 7674 3194 7677
rect 3197 7674 3199 7676
rect 3218 7674 3220 7676
rect 3234 7674 3236 7686
rect 3250 7684 3252 7693
rect 3255 7691 3257 7693
rect 3250 7674 3252 7677
rect 3255 7674 3257 7676
rect 3271 7674 3273 7693
rect 4100 7688 4102 7693
rect 4105 7691 4107 7693
rect 4100 7674 4102 7684
rect 4105 7674 4107 7681
rect 4121 7674 4123 7693
rect 4137 7684 4139 7693
rect 4142 7691 4144 7693
rect 4163 7691 4165 7693
rect 4179 7690 4181 7693
rect 4137 7674 4139 7677
rect 4142 7674 4144 7676
rect 4163 7674 4165 7676
rect 4179 7674 4181 7686
rect 4195 7684 4197 7693
rect 4200 7691 4202 7693
rect 4195 7674 4197 7677
rect 4200 7674 4202 7676
rect 4216 7674 4218 7693
rect 2372 7671 2374 7673
rect 2377 7671 2379 7674
rect 2393 7671 2395 7673
rect 2409 7671 2411 7673
rect 2414 7671 2416 7674
rect 2435 7671 2437 7674
rect 2451 7671 2453 7674
rect 2467 7671 2469 7673
rect 2472 7671 2474 7674
rect 2488 7671 2490 7673
rect 2504 7671 2506 7673
rect 2509 7671 2511 7674
rect 2525 7671 2527 7673
rect 2541 7671 2543 7673
rect 2546 7671 2548 7674
rect 2567 7671 2569 7674
rect 2583 7671 2585 7674
rect 2599 7671 2601 7673
rect 2604 7671 2606 7674
rect 2620 7671 2622 7673
rect 2636 7671 2638 7673
rect 2641 7671 2643 7674
rect 2657 7671 2659 7673
rect 2673 7671 2675 7673
rect 2678 7671 2680 7674
rect 2699 7671 2701 7674
rect 2715 7671 2717 7674
rect 2731 7671 2733 7673
rect 2736 7671 2738 7674
rect 2752 7671 2754 7673
rect 3317 7671 3319 7673
rect 3322 7671 3324 7674
rect 3338 7671 3340 7673
rect 3354 7671 3356 7673
rect 3359 7671 3361 7674
rect 3380 7671 3382 7674
rect 3396 7671 3398 7674
rect 3412 7671 3414 7673
rect 3417 7671 3419 7674
rect 3433 7671 3435 7673
rect 3449 7671 3451 7673
rect 3454 7671 3456 7674
rect 3470 7671 3472 7673
rect 3486 7671 3488 7673
rect 3491 7671 3493 7674
rect 3512 7671 3514 7674
rect 3528 7671 3530 7674
rect 3544 7671 3546 7673
rect 3549 7671 3551 7674
rect 3565 7671 3567 7673
rect 3581 7671 3583 7673
rect 3586 7671 3588 7674
rect 3602 7671 3604 7673
rect 3618 7671 3620 7673
rect 3623 7671 3625 7674
rect 3644 7671 3646 7674
rect 3660 7671 3662 7674
rect 3676 7671 3678 7673
rect 3681 7671 3683 7674
rect 3697 7671 3699 7673
rect 3155 7668 3157 7670
rect 3160 7667 3162 7670
rect 3176 7668 3178 7670
rect 3192 7668 3194 7670
rect 3197 7665 3199 7670
rect 3218 7665 3220 7670
rect 3234 7668 3236 7670
rect 3250 7668 3252 7670
rect 3255 7665 3257 7670
rect 3271 7668 3273 7670
rect 2372 7658 2374 7663
rect 2377 7661 2379 7663
rect 2372 7644 2374 7654
rect 2377 7644 2379 7651
rect 2393 7644 2395 7663
rect 2409 7654 2411 7663
rect 2414 7661 2416 7663
rect 2435 7661 2437 7663
rect 2451 7660 2453 7663
rect 2409 7644 2411 7647
rect 2414 7644 2416 7646
rect 2435 7644 2437 7646
rect 2451 7644 2453 7656
rect 2467 7654 2469 7663
rect 2472 7661 2474 7663
rect 2467 7644 2469 7647
rect 2472 7644 2474 7646
rect 2488 7644 2490 7663
rect 2504 7660 2506 7663
rect 2509 7661 2511 7663
rect 2504 7644 2506 7656
rect 2509 7644 2511 7651
rect 2525 7644 2527 7663
rect 2541 7654 2543 7663
rect 2546 7661 2548 7663
rect 2567 7661 2569 7663
rect 2583 7660 2585 7663
rect 2541 7644 2543 7647
rect 2546 7644 2548 7646
rect 2567 7644 2569 7646
rect 2583 7644 2585 7656
rect 2599 7654 2601 7663
rect 2604 7661 2606 7663
rect 2599 7644 2601 7647
rect 2604 7644 2606 7646
rect 2620 7644 2622 7663
rect 2636 7660 2638 7663
rect 2641 7661 2643 7663
rect 2636 7644 2638 7656
rect 2641 7644 2643 7651
rect 2657 7644 2659 7663
rect 2673 7654 2675 7663
rect 2678 7661 2680 7663
rect 2699 7661 2701 7663
rect 2715 7660 2717 7663
rect 2673 7644 2675 7647
rect 2678 7644 2680 7646
rect 2699 7644 2701 7646
rect 2715 7644 2717 7656
rect 2731 7654 2733 7663
rect 2736 7661 2738 7663
rect 2752 7655 2754 7663
rect 4100 7668 4102 7670
rect 4105 7667 4107 7670
rect 4121 7668 4123 7670
rect 4137 7668 4139 7670
rect 4142 7665 4144 7670
rect 4163 7665 4165 7670
rect 4179 7668 4181 7670
rect 4195 7668 4197 7670
rect 4200 7665 4202 7670
rect 4216 7668 4218 7670
rect 3317 7658 3319 7663
rect 3322 7661 3324 7663
rect 2731 7644 2733 7647
rect 2736 7644 2738 7646
rect 2752 7644 2754 7651
rect 3317 7644 3319 7654
rect 3322 7644 3324 7651
rect 3338 7644 3340 7663
rect 3354 7654 3356 7663
rect 3359 7661 3361 7663
rect 3380 7661 3382 7663
rect 3396 7660 3398 7663
rect 3354 7644 3356 7647
rect 3359 7644 3361 7646
rect 3380 7644 3382 7646
rect 3396 7644 3398 7656
rect 3412 7654 3414 7663
rect 3417 7661 3419 7663
rect 3412 7644 3414 7647
rect 3417 7644 3419 7646
rect 3433 7644 3435 7663
rect 3449 7660 3451 7663
rect 3454 7661 3456 7663
rect 3449 7644 3451 7656
rect 3454 7644 3456 7651
rect 3470 7644 3472 7663
rect 3486 7654 3488 7663
rect 3491 7661 3493 7663
rect 3512 7661 3514 7663
rect 3528 7660 3530 7663
rect 3486 7644 3488 7647
rect 3491 7644 3493 7646
rect 3512 7644 3514 7646
rect 3528 7644 3530 7656
rect 3544 7654 3546 7663
rect 3549 7661 3551 7663
rect 3544 7644 3546 7647
rect 3549 7644 3551 7646
rect 3565 7644 3567 7663
rect 3581 7660 3583 7663
rect 3586 7661 3588 7663
rect 3581 7644 3583 7656
rect 3586 7644 3588 7651
rect 3602 7644 3604 7663
rect 3618 7654 3620 7663
rect 3623 7661 3625 7663
rect 3644 7661 3646 7663
rect 3660 7660 3662 7663
rect 3618 7644 3620 7647
rect 3623 7644 3625 7646
rect 3644 7644 3646 7646
rect 3660 7644 3662 7656
rect 3676 7654 3678 7663
rect 3681 7661 3683 7663
rect 3697 7655 3699 7663
rect 3676 7644 3678 7647
rect 3681 7644 3683 7646
rect 3697 7644 3699 7651
rect 2372 7638 2374 7640
rect 2377 7637 2379 7640
rect 2393 7638 2395 7640
rect 2409 7638 2411 7640
rect 2414 7635 2416 7640
rect 2435 7635 2437 7640
rect 2451 7638 2453 7640
rect 2467 7638 2469 7640
rect 2472 7635 2474 7640
rect 2488 7638 2490 7640
rect 2504 7638 2506 7640
rect 2509 7637 2511 7640
rect 2525 7638 2527 7640
rect 2541 7638 2543 7640
rect 2546 7635 2548 7640
rect 2567 7635 2569 7640
rect 2583 7638 2585 7640
rect 2599 7638 2601 7640
rect 2604 7635 2606 7640
rect 2620 7638 2622 7640
rect 2636 7638 2638 7640
rect 2641 7637 2643 7640
rect 2657 7638 2659 7640
rect 2673 7638 2675 7640
rect 2678 7635 2680 7640
rect 2699 7635 2701 7640
rect 2715 7638 2717 7640
rect 2731 7638 2733 7640
rect 2736 7635 2738 7640
rect 2752 7638 2754 7640
rect 3317 7638 3319 7640
rect 3322 7637 3324 7640
rect 3338 7638 3340 7640
rect 3354 7638 3356 7640
rect 3359 7635 3361 7640
rect 3380 7635 3382 7640
rect 3396 7638 3398 7640
rect 3412 7638 3414 7640
rect 3417 7635 3419 7640
rect 3433 7638 3435 7640
rect 3449 7638 3451 7640
rect 3454 7637 3456 7640
rect 3470 7638 3472 7640
rect 3486 7638 3488 7640
rect 3491 7635 3493 7640
rect 3512 7635 3514 7640
rect 3528 7638 3530 7640
rect 3544 7638 3546 7640
rect 3549 7635 3551 7640
rect 3565 7638 3567 7640
rect 3581 7638 3583 7640
rect 3586 7637 3588 7640
rect 3602 7638 3604 7640
rect 3618 7638 3620 7640
rect 3623 7635 3625 7640
rect 3644 7635 3646 7640
rect 3660 7638 3662 7640
rect 3676 7638 3678 7640
rect 3681 7635 3683 7640
rect 3697 7638 3699 7640
rect 3155 7615 3157 7617
rect 3160 7615 3162 7618
rect 3176 7615 3178 7617
rect 3192 7615 3194 7617
rect 3197 7615 3199 7618
rect 3218 7615 3220 7618
rect 3234 7615 3236 7618
rect 3250 7615 3252 7617
rect 3255 7615 3257 7618
rect 3271 7615 3273 7617
rect 4100 7615 4102 7617
rect 4105 7615 4107 7618
rect 4121 7615 4123 7617
rect 4137 7615 4139 7617
rect 4142 7615 4144 7618
rect 4163 7615 4165 7618
rect 4179 7615 4181 7618
rect 4195 7615 4197 7617
rect 4200 7615 4202 7618
rect 4216 7615 4218 7617
rect 3155 7602 3157 7607
rect 3160 7605 3162 7607
rect 3155 7588 3157 7598
rect 3160 7588 3162 7595
rect 3176 7588 3178 7607
rect 3192 7598 3194 7607
rect 3197 7605 3199 7607
rect 3218 7605 3220 7607
rect 3234 7604 3236 7607
rect 3192 7588 3194 7591
rect 3197 7588 3199 7590
rect 3218 7588 3220 7590
rect 3234 7588 3236 7600
rect 3250 7598 3252 7607
rect 3255 7605 3257 7607
rect 3250 7588 3252 7591
rect 3255 7588 3257 7590
rect 3271 7588 3273 7607
rect 4100 7602 4102 7607
rect 4105 7605 4107 7607
rect 3293 7594 3296 7596
rect 3300 7594 3303 7596
rect 4100 7588 4102 7598
rect 4105 7588 4107 7595
rect 4121 7588 4123 7607
rect 4137 7598 4139 7607
rect 4142 7605 4144 7607
rect 4163 7605 4165 7607
rect 4179 7604 4181 7607
rect 4137 7588 4139 7591
rect 4142 7588 4144 7590
rect 4163 7588 4165 7590
rect 4179 7588 4181 7600
rect 4195 7598 4197 7607
rect 4200 7605 4202 7607
rect 4195 7588 4197 7591
rect 4200 7588 4202 7590
rect 4216 7588 4218 7607
rect 4238 7594 4241 7596
rect 4245 7594 4248 7596
rect 2372 7585 2374 7587
rect 2377 7585 2379 7588
rect 2393 7585 2395 7587
rect 2409 7585 2411 7587
rect 2414 7585 2416 7588
rect 2435 7585 2437 7588
rect 2451 7585 2453 7588
rect 2467 7585 2469 7587
rect 2472 7585 2474 7588
rect 2488 7585 2490 7587
rect 2504 7585 2506 7587
rect 2509 7585 2511 7588
rect 2525 7585 2527 7587
rect 2541 7585 2543 7587
rect 2546 7585 2548 7588
rect 2567 7585 2569 7588
rect 2583 7585 2585 7588
rect 2599 7585 2601 7587
rect 2604 7585 2606 7588
rect 2620 7585 2622 7587
rect 2636 7585 2638 7587
rect 2641 7585 2643 7588
rect 2657 7585 2659 7587
rect 2673 7585 2675 7587
rect 2678 7585 2680 7588
rect 2699 7585 2701 7588
rect 2715 7585 2717 7588
rect 2731 7585 2733 7587
rect 2736 7585 2738 7588
rect 2752 7585 2754 7587
rect 3317 7585 3319 7587
rect 3322 7585 3324 7588
rect 3338 7585 3340 7587
rect 3354 7585 3356 7587
rect 3359 7585 3361 7588
rect 3380 7585 3382 7588
rect 3396 7585 3398 7588
rect 3412 7585 3414 7587
rect 3417 7585 3419 7588
rect 3433 7585 3435 7587
rect 3449 7585 3451 7587
rect 3454 7585 3456 7588
rect 3470 7585 3472 7587
rect 3486 7585 3488 7587
rect 3491 7585 3493 7588
rect 3512 7585 3514 7588
rect 3528 7585 3530 7588
rect 3544 7585 3546 7587
rect 3549 7585 3551 7588
rect 3565 7585 3567 7587
rect 3581 7585 3583 7587
rect 3586 7585 3588 7588
rect 3602 7585 3604 7587
rect 3618 7585 3620 7587
rect 3623 7585 3625 7588
rect 3644 7585 3646 7588
rect 3660 7585 3662 7588
rect 3676 7585 3678 7587
rect 3681 7585 3683 7588
rect 3697 7585 3699 7587
rect 3155 7582 3157 7584
rect 3160 7581 3162 7584
rect 3176 7582 3178 7584
rect 3192 7582 3194 7584
rect 3197 7579 3199 7584
rect 3218 7579 3220 7584
rect 3234 7582 3236 7584
rect 3250 7582 3252 7584
rect 3255 7579 3257 7584
rect 3271 7582 3273 7584
rect 2372 7572 2374 7577
rect 2377 7575 2379 7577
rect 2372 7558 2374 7568
rect 2377 7558 2379 7565
rect 2393 7558 2395 7577
rect 2409 7568 2411 7577
rect 2414 7575 2416 7577
rect 2435 7575 2437 7577
rect 2451 7574 2453 7577
rect 2409 7558 2411 7561
rect 2414 7558 2416 7560
rect 2435 7558 2437 7560
rect 2451 7558 2453 7570
rect 2467 7568 2469 7577
rect 2472 7575 2474 7577
rect 2467 7558 2469 7561
rect 2472 7558 2474 7560
rect 2488 7558 2490 7577
rect 2504 7574 2506 7577
rect 2509 7575 2511 7577
rect 2504 7558 2506 7570
rect 2509 7558 2511 7565
rect 2525 7558 2527 7577
rect 2541 7568 2543 7577
rect 2546 7575 2548 7577
rect 2567 7575 2569 7577
rect 2583 7574 2585 7577
rect 2541 7558 2543 7561
rect 2546 7558 2548 7560
rect 2567 7558 2569 7560
rect 2583 7558 2585 7570
rect 2599 7568 2601 7577
rect 2604 7575 2606 7577
rect 2599 7558 2601 7561
rect 2604 7558 2606 7560
rect 2620 7558 2622 7577
rect 2636 7574 2638 7577
rect 2641 7575 2643 7577
rect 2636 7558 2638 7570
rect 2641 7558 2643 7565
rect 2657 7558 2659 7577
rect 2673 7568 2675 7577
rect 2678 7575 2680 7577
rect 2699 7575 2701 7577
rect 2715 7574 2717 7577
rect 2673 7558 2675 7561
rect 2678 7558 2680 7560
rect 2699 7558 2701 7560
rect 2715 7558 2717 7570
rect 2731 7568 2733 7577
rect 2736 7575 2738 7577
rect 2752 7569 2754 7577
rect 4100 7582 4102 7584
rect 4105 7581 4107 7584
rect 4121 7582 4123 7584
rect 4137 7582 4139 7584
rect 4142 7579 4144 7584
rect 4163 7579 4165 7584
rect 4179 7582 4181 7584
rect 4195 7582 4197 7584
rect 4200 7579 4202 7584
rect 4216 7582 4218 7584
rect 3317 7572 3319 7577
rect 3322 7575 3324 7577
rect 2731 7558 2733 7561
rect 2736 7558 2738 7560
rect 2752 7558 2754 7565
rect 3317 7558 3319 7568
rect 3322 7558 3324 7565
rect 3338 7558 3340 7577
rect 3354 7568 3356 7577
rect 3359 7575 3361 7577
rect 3380 7575 3382 7577
rect 3396 7574 3398 7577
rect 3354 7558 3356 7561
rect 3359 7558 3361 7560
rect 3380 7558 3382 7560
rect 3396 7558 3398 7570
rect 3412 7568 3414 7577
rect 3417 7575 3419 7577
rect 3412 7558 3414 7561
rect 3417 7558 3419 7560
rect 3433 7558 3435 7577
rect 3449 7574 3451 7577
rect 3454 7575 3456 7577
rect 3449 7558 3451 7570
rect 3454 7558 3456 7565
rect 3470 7558 3472 7577
rect 3486 7568 3488 7577
rect 3491 7575 3493 7577
rect 3512 7575 3514 7577
rect 3528 7574 3530 7577
rect 3486 7558 3488 7561
rect 3491 7558 3493 7560
rect 3512 7558 3514 7560
rect 3528 7558 3530 7570
rect 3544 7568 3546 7577
rect 3549 7575 3551 7577
rect 3544 7558 3546 7561
rect 3549 7558 3551 7560
rect 3565 7558 3567 7577
rect 3581 7574 3583 7577
rect 3586 7575 3588 7577
rect 3581 7558 3583 7570
rect 3586 7558 3588 7565
rect 3602 7558 3604 7577
rect 3618 7568 3620 7577
rect 3623 7575 3625 7577
rect 3644 7575 3646 7577
rect 3660 7574 3662 7577
rect 3618 7558 3620 7561
rect 3623 7558 3625 7560
rect 3644 7558 3646 7560
rect 3660 7558 3662 7570
rect 3676 7568 3678 7577
rect 3681 7575 3683 7577
rect 3697 7569 3699 7577
rect 3676 7558 3678 7561
rect 3681 7558 3683 7560
rect 3697 7558 3699 7565
rect 2372 7552 2374 7554
rect 2377 7551 2379 7554
rect 2393 7552 2395 7554
rect 2409 7552 2411 7554
rect 2414 7549 2416 7554
rect 2435 7549 2437 7554
rect 2451 7552 2453 7554
rect 2467 7552 2469 7554
rect 2472 7549 2474 7554
rect 2488 7552 2490 7554
rect 2504 7552 2506 7554
rect 2509 7551 2511 7554
rect 2525 7552 2527 7554
rect 2541 7552 2543 7554
rect 2546 7549 2548 7554
rect 2567 7549 2569 7554
rect 2583 7552 2585 7554
rect 2599 7552 2601 7554
rect 2604 7549 2606 7554
rect 2620 7552 2622 7554
rect 2636 7552 2638 7554
rect 2641 7551 2643 7554
rect 2657 7552 2659 7554
rect 2673 7552 2675 7554
rect 2678 7549 2680 7554
rect 2699 7549 2701 7554
rect 2715 7552 2717 7554
rect 2731 7552 2733 7554
rect 2736 7549 2738 7554
rect 2752 7552 2754 7554
rect 3317 7552 3319 7554
rect 3322 7551 3324 7554
rect 3338 7552 3340 7554
rect 3354 7552 3356 7554
rect 3359 7549 3361 7554
rect 3380 7549 3382 7554
rect 3396 7552 3398 7554
rect 3412 7552 3414 7554
rect 3417 7549 3419 7554
rect 3433 7552 3435 7554
rect 3449 7552 3451 7554
rect 3454 7551 3456 7554
rect 3470 7552 3472 7554
rect 3486 7552 3488 7554
rect 3491 7549 3493 7554
rect 3512 7549 3514 7554
rect 3528 7552 3530 7554
rect 3544 7552 3546 7554
rect 3549 7549 3551 7554
rect 3565 7552 3567 7554
rect 3581 7552 3583 7554
rect 3586 7551 3588 7554
rect 3602 7552 3604 7554
rect 3618 7552 3620 7554
rect 3623 7549 3625 7554
rect 3644 7549 3646 7554
rect 3660 7552 3662 7554
rect 3676 7552 3678 7554
rect 3681 7549 3683 7554
rect 3697 7552 3699 7554
rect 2604 7514 2606 7517
rect 2628 7514 2630 7517
rect 3549 7514 3551 7517
rect 3573 7514 3575 7517
rect 2604 7508 2606 7510
rect 2628 7508 2630 7510
rect 3549 7508 3551 7510
rect 3573 7508 3575 7510
rect 2624 7503 2626 7505
rect 3569 7503 3571 7505
rect 2624 7496 2626 7499
rect 3569 7496 3571 7499
rect 2613 7485 2615 7487
rect 2619 7485 2638 7487
rect 3558 7485 3560 7487
rect 3564 7485 3583 7487
rect 2604 7480 2606 7482
rect 2628 7480 2630 7482
rect 3549 7480 3551 7482
rect 3573 7480 3575 7482
rect 2604 7473 2606 7476
rect 2628 7473 2630 7476
rect 3549 7473 3551 7476
rect 3573 7473 3575 7476
rect 3832 7473 3836 7475
rect 3844 7473 3847 7475
rect 2372 7445 2374 7447
rect 2377 7445 2379 7448
rect 2393 7445 2395 7447
rect 2409 7445 2411 7447
rect 2414 7445 2416 7448
rect 2435 7445 2437 7448
rect 2451 7445 2453 7448
rect 2467 7445 2469 7447
rect 2472 7445 2474 7448
rect 2488 7445 2490 7447
rect 2504 7445 2506 7447
rect 2509 7445 2511 7448
rect 2525 7445 2527 7447
rect 2541 7445 2543 7447
rect 2546 7445 2548 7448
rect 2567 7445 2569 7448
rect 2583 7445 2585 7448
rect 2599 7445 2601 7447
rect 2604 7445 2606 7448
rect 2620 7445 2622 7447
rect 2636 7445 2638 7447
rect 2641 7445 2643 7448
rect 2657 7445 2659 7447
rect 2673 7445 2675 7447
rect 2678 7445 2680 7448
rect 2699 7445 2701 7448
rect 2715 7445 2717 7448
rect 2731 7445 2733 7447
rect 2736 7445 2738 7448
rect 2752 7445 2754 7447
rect 3317 7445 3319 7447
rect 3322 7445 3324 7448
rect 3338 7445 3340 7447
rect 3354 7445 3356 7447
rect 3359 7445 3361 7448
rect 3380 7445 3382 7448
rect 3396 7445 3398 7448
rect 3412 7445 3414 7447
rect 3417 7445 3419 7448
rect 3433 7445 3435 7447
rect 3449 7445 3451 7447
rect 3454 7445 3456 7448
rect 3470 7445 3472 7447
rect 3486 7445 3488 7447
rect 3491 7445 3493 7448
rect 3512 7445 3514 7448
rect 3528 7445 3530 7448
rect 3544 7445 3546 7447
rect 3549 7445 3551 7448
rect 3565 7445 3567 7447
rect 3581 7445 3583 7447
rect 3586 7445 3588 7448
rect 3602 7445 3604 7447
rect 3618 7445 3620 7447
rect 3623 7445 3625 7448
rect 3644 7445 3646 7448
rect 3660 7445 3662 7448
rect 3676 7445 3678 7447
rect 3681 7445 3683 7448
rect 3697 7445 3699 7447
rect 2372 7432 2374 7437
rect 2377 7435 2379 7437
rect 2372 7418 2374 7428
rect 2377 7418 2379 7425
rect 2393 7418 2395 7437
rect 2409 7428 2411 7437
rect 2414 7435 2416 7437
rect 2435 7435 2437 7437
rect 2451 7434 2453 7437
rect 2409 7418 2411 7421
rect 2414 7418 2416 7420
rect 2435 7418 2437 7420
rect 2451 7418 2453 7430
rect 2467 7428 2469 7437
rect 2472 7435 2474 7437
rect 2467 7418 2469 7421
rect 2472 7418 2474 7420
rect 2488 7418 2490 7437
rect 2504 7434 2506 7437
rect 2509 7435 2511 7437
rect 2504 7418 2506 7430
rect 2509 7418 2511 7425
rect 2525 7418 2527 7437
rect 2541 7428 2543 7437
rect 2546 7435 2548 7437
rect 2567 7435 2569 7437
rect 2583 7434 2585 7437
rect 2541 7418 2543 7421
rect 2546 7418 2548 7420
rect 2567 7418 2569 7420
rect 2583 7418 2585 7430
rect 2599 7428 2601 7437
rect 2604 7435 2606 7437
rect 2599 7418 2601 7421
rect 2604 7418 2606 7420
rect 2620 7418 2622 7437
rect 2636 7434 2638 7437
rect 2641 7435 2643 7437
rect 2636 7418 2638 7430
rect 2641 7418 2643 7425
rect 2657 7418 2659 7437
rect 2673 7428 2675 7437
rect 2678 7435 2680 7437
rect 2699 7435 2701 7437
rect 2715 7434 2717 7437
rect 2673 7418 2675 7421
rect 2678 7418 2680 7420
rect 2699 7418 2701 7420
rect 2715 7418 2717 7430
rect 2731 7428 2733 7437
rect 2736 7435 2738 7437
rect 2752 7429 2754 7437
rect 3317 7432 3319 7437
rect 3322 7435 3324 7437
rect 2731 7418 2733 7421
rect 2736 7418 2738 7420
rect 2752 7418 2754 7425
rect 3317 7418 3319 7428
rect 3322 7418 3324 7425
rect 3338 7418 3340 7437
rect 3354 7428 3356 7437
rect 3359 7435 3361 7437
rect 3380 7435 3382 7437
rect 3396 7434 3398 7437
rect 3354 7418 3356 7421
rect 3359 7418 3361 7420
rect 3380 7418 3382 7420
rect 3396 7418 3398 7430
rect 3412 7428 3414 7437
rect 3417 7435 3419 7437
rect 3412 7418 3414 7421
rect 3417 7418 3419 7420
rect 3433 7418 3435 7437
rect 3449 7434 3451 7437
rect 3454 7435 3456 7437
rect 3449 7418 3451 7430
rect 3454 7418 3456 7425
rect 3470 7418 3472 7437
rect 3486 7428 3488 7437
rect 3491 7435 3493 7437
rect 3512 7435 3514 7437
rect 3528 7434 3530 7437
rect 3486 7418 3488 7421
rect 3491 7418 3493 7420
rect 3512 7418 3514 7420
rect 3528 7418 3530 7430
rect 3544 7428 3546 7437
rect 3549 7435 3551 7437
rect 3544 7418 3546 7421
rect 3549 7418 3551 7420
rect 3565 7418 3567 7437
rect 3581 7434 3583 7437
rect 3586 7435 3588 7437
rect 3581 7418 3583 7430
rect 3586 7418 3588 7425
rect 3602 7418 3604 7437
rect 3618 7428 3620 7437
rect 3623 7435 3625 7437
rect 3644 7435 3646 7437
rect 3660 7434 3662 7437
rect 3618 7418 3620 7421
rect 3623 7418 3625 7420
rect 3644 7418 3646 7420
rect 3660 7418 3662 7430
rect 3676 7428 3678 7437
rect 3681 7435 3683 7437
rect 3697 7429 3699 7437
rect 3676 7418 3678 7421
rect 3681 7418 3683 7420
rect 3697 7418 3699 7425
rect 2372 7412 2374 7414
rect 2377 7411 2379 7414
rect 2393 7412 2395 7414
rect 2409 7412 2411 7414
rect 2414 7409 2416 7414
rect 2435 7409 2437 7414
rect 2451 7412 2453 7414
rect 2467 7412 2469 7414
rect 2472 7409 2474 7414
rect 2488 7412 2490 7414
rect 2504 7412 2506 7414
rect 2509 7411 2511 7414
rect 2525 7412 2527 7414
rect 2541 7412 2543 7414
rect 2546 7409 2548 7414
rect 2567 7409 2569 7414
rect 2583 7412 2585 7414
rect 2599 7412 2601 7414
rect 2604 7409 2606 7414
rect 2620 7412 2622 7414
rect 2636 7412 2638 7414
rect 2641 7411 2643 7414
rect 2657 7412 2659 7414
rect 2673 7412 2675 7414
rect 2678 7409 2680 7414
rect 2699 7409 2701 7414
rect 2715 7412 2717 7414
rect 2731 7412 2733 7414
rect 2736 7409 2738 7414
rect 2752 7412 2754 7414
rect 3317 7412 3319 7414
rect 3322 7411 3324 7414
rect 3338 7412 3340 7414
rect 3354 7412 3356 7414
rect 3359 7409 3361 7414
rect 3380 7409 3382 7414
rect 3396 7412 3398 7414
rect 3412 7412 3414 7414
rect 3417 7409 3419 7414
rect 3433 7412 3435 7414
rect 3449 7412 3451 7414
rect 3454 7411 3456 7414
rect 3470 7412 3472 7414
rect 3486 7412 3488 7414
rect 3491 7409 3493 7414
rect 3512 7409 3514 7414
rect 3528 7412 3530 7414
rect 3544 7412 3546 7414
rect 3549 7409 3551 7414
rect 3565 7412 3567 7414
rect 3581 7412 3583 7414
rect 3586 7411 3588 7414
rect 3602 7412 3604 7414
rect 3618 7412 3620 7414
rect 3623 7409 3625 7414
rect 3644 7409 3646 7414
rect 3660 7412 3662 7414
rect 3676 7412 3678 7414
rect 3681 7409 3683 7414
rect 3697 7412 3699 7414
rect 1473 6900 1475 6902
rect 1489 6900 1491 6905
rect 1494 6900 1496 6902
rect 1510 6900 1512 6902
rect 1526 6900 1528 6905
rect 1547 6900 1549 6905
rect 1552 6900 1554 6902
rect 1568 6900 1570 6902
rect 1584 6900 1586 6903
rect 1589 6900 1591 6902
rect 1605 6900 1607 6902
rect 1621 6900 1623 6905
rect 1626 6900 1628 6902
rect 1642 6900 1644 6902
rect 1658 6900 1660 6905
rect 1679 6900 1681 6905
rect 1684 6900 1686 6902
rect 1700 6900 1702 6902
rect 1716 6900 1718 6903
rect 1721 6900 1723 6902
rect 1737 6900 1739 6902
rect 1753 6900 1755 6905
rect 1758 6900 1760 6902
rect 1774 6900 1776 6902
rect 1790 6900 1792 6905
rect 1811 6900 1813 6905
rect 1816 6900 1818 6902
rect 1832 6900 1834 6902
rect 1848 6900 1850 6903
rect 1853 6900 1855 6902
rect 2418 6900 2420 6902
rect 2434 6900 2436 6905
rect 2439 6900 2441 6902
rect 2455 6900 2457 6902
rect 2471 6900 2473 6905
rect 2492 6900 2494 6905
rect 2497 6900 2499 6902
rect 2513 6900 2515 6902
rect 2529 6900 2531 6903
rect 2534 6900 2536 6902
rect 2550 6900 2552 6902
rect 2566 6900 2568 6905
rect 2571 6900 2573 6902
rect 2587 6900 2589 6902
rect 2603 6900 2605 6905
rect 2624 6900 2626 6905
rect 2629 6900 2631 6902
rect 2645 6900 2647 6902
rect 2661 6900 2663 6903
rect 2666 6900 2668 6902
rect 2682 6900 2684 6902
rect 2698 6900 2700 6905
rect 2703 6900 2705 6902
rect 2719 6900 2721 6902
rect 2735 6900 2737 6905
rect 2756 6900 2758 6905
rect 2761 6900 2763 6902
rect 2777 6900 2779 6902
rect 2793 6900 2795 6903
rect 2798 6900 2800 6902
rect 1473 6889 1475 6896
rect 1489 6894 1491 6896
rect 1494 6893 1496 6896
rect 1473 6877 1475 6885
rect 1489 6877 1491 6879
rect 1494 6877 1496 6886
rect 1510 6884 1512 6896
rect 1526 6894 1528 6896
rect 1547 6894 1549 6896
rect 1552 6893 1554 6896
rect 1510 6877 1512 6880
rect 1526 6877 1528 6879
rect 1547 6877 1549 6879
rect 1552 6877 1554 6886
rect 1568 6877 1570 6896
rect 1584 6889 1586 6896
rect 1589 6884 1591 6896
rect 1584 6877 1586 6879
rect 1589 6877 1591 6880
rect 1605 6877 1607 6896
rect 1621 6894 1623 6896
rect 1626 6893 1628 6896
rect 1621 6877 1623 6879
rect 1626 6877 1628 6886
rect 1642 6884 1644 6896
rect 1658 6894 1660 6896
rect 1679 6894 1681 6896
rect 1684 6893 1686 6896
rect 1642 6877 1644 6880
rect 1658 6877 1660 6879
rect 1679 6877 1681 6879
rect 1684 6877 1686 6886
rect 1700 6877 1702 6896
rect 1716 6889 1718 6896
rect 1721 6884 1723 6896
rect 1716 6877 1718 6879
rect 1721 6877 1723 6880
rect 1737 6877 1739 6896
rect 1753 6894 1755 6896
rect 1758 6893 1760 6896
rect 1753 6877 1755 6879
rect 1758 6877 1760 6886
rect 1774 6884 1776 6896
rect 1790 6894 1792 6896
rect 1811 6894 1813 6896
rect 1816 6893 1818 6896
rect 1774 6877 1776 6880
rect 1790 6877 1792 6879
rect 1811 6877 1813 6879
rect 1816 6877 1818 6886
rect 1832 6877 1834 6896
rect 1848 6889 1850 6896
rect 1853 6886 1855 6896
rect 2418 6889 2420 6896
rect 2434 6894 2436 6896
rect 2439 6893 2441 6896
rect 1848 6877 1850 6879
rect 1853 6877 1855 6882
rect 2418 6877 2420 6885
rect 2434 6877 2436 6879
rect 2439 6877 2441 6886
rect 2455 6884 2457 6896
rect 2471 6894 2473 6896
rect 2492 6894 2494 6896
rect 2497 6893 2499 6896
rect 2455 6877 2457 6880
rect 2471 6877 2473 6879
rect 2492 6877 2494 6879
rect 2497 6877 2499 6886
rect 2513 6877 2515 6896
rect 2529 6889 2531 6896
rect 2534 6884 2536 6896
rect 2529 6877 2531 6879
rect 2534 6877 2536 6880
rect 2550 6877 2552 6896
rect 2566 6894 2568 6896
rect 2571 6893 2573 6896
rect 2566 6877 2568 6879
rect 2571 6877 2573 6886
rect 2587 6884 2589 6896
rect 2603 6894 2605 6896
rect 2624 6894 2626 6896
rect 2629 6893 2631 6896
rect 2587 6877 2589 6880
rect 2603 6877 2605 6879
rect 2624 6877 2626 6879
rect 2629 6877 2631 6886
rect 2645 6877 2647 6896
rect 2661 6889 2663 6896
rect 2666 6884 2668 6896
rect 2661 6877 2663 6879
rect 2666 6877 2668 6880
rect 2682 6877 2684 6896
rect 2698 6894 2700 6896
rect 2703 6893 2705 6896
rect 2698 6877 2700 6879
rect 2703 6877 2705 6886
rect 2719 6884 2721 6896
rect 2735 6894 2737 6896
rect 2756 6894 2758 6896
rect 2761 6893 2763 6896
rect 2719 6877 2721 6880
rect 2735 6877 2737 6879
rect 2756 6877 2758 6879
rect 2761 6877 2763 6886
rect 2777 6877 2779 6896
rect 2793 6889 2795 6896
rect 2798 6886 2800 6896
rect 2793 6877 2795 6879
rect 2798 6877 2800 6882
rect 1473 6867 1475 6869
rect 1489 6866 1491 6869
rect 1494 6867 1496 6869
rect 1510 6866 1512 6869
rect 1526 6866 1528 6869
rect 1547 6866 1549 6869
rect 1552 6867 1554 6869
rect 1568 6867 1570 6869
rect 1584 6866 1586 6869
rect 1589 6867 1591 6869
rect 1605 6867 1607 6869
rect 1621 6866 1623 6869
rect 1626 6867 1628 6869
rect 1642 6866 1644 6869
rect 1658 6866 1660 6869
rect 1679 6866 1681 6869
rect 1684 6867 1686 6869
rect 1700 6867 1702 6869
rect 1716 6866 1718 6869
rect 1721 6867 1723 6869
rect 1737 6867 1739 6869
rect 1753 6866 1755 6869
rect 1758 6867 1760 6869
rect 1774 6866 1776 6869
rect 1790 6866 1792 6869
rect 1811 6866 1813 6869
rect 1816 6867 1818 6869
rect 1832 6867 1834 6869
rect 1848 6866 1850 6869
rect 1853 6867 1855 6869
rect 2418 6867 2420 6869
rect 2434 6866 2436 6869
rect 2439 6867 2441 6869
rect 2455 6866 2457 6869
rect 2471 6866 2473 6869
rect 2492 6866 2494 6869
rect 2497 6867 2499 6869
rect 2513 6867 2515 6869
rect 2529 6866 2531 6869
rect 2534 6867 2536 6869
rect 2550 6867 2552 6869
rect 2566 6866 2568 6869
rect 2571 6867 2573 6869
rect 2587 6866 2589 6869
rect 2603 6866 2605 6869
rect 2624 6866 2626 6869
rect 2629 6867 2631 6869
rect 2645 6867 2647 6869
rect 2661 6866 2663 6869
rect 2666 6867 2668 6869
rect 2682 6867 2684 6869
rect 2698 6866 2700 6869
rect 2703 6867 2705 6869
rect 2719 6866 2721 6869
rect 2735 6866 2737 6869
rect 2756 6866 2758 6869
rect 2761 6867 2763 6869
rect 2777 6867 2779 6869
rect 2793 6866 2795 6869
rect 2798 6867 2800 6869
rect 1597 6838 1599 6841
rect 1621 6838 1623 6841
rect 2542 6838 2544 6841
rect 2566 6838 2568 6841
rect 1597 6832 1599 6834
rect 1621 6832 1623 6834
rect 2542 6832 2544 6834
rect 2566 6832 2568 6834
rect 1589 6827 1608 6829
rect 1612 6827 1614 6829
rect 2534 6827 2553 6829
rect 2557 6827 2559 6829
rect 1601 6815 1603 6818
rect 2546 6815 2548 6818
rect 1601 6809 1603 6811
rect 2546 6809 2548 6811
rect 1597 6804 1599 6806
rect 1621 6804 1623 6806
rect 2542 6804 2544 6806
rect 2566 6804 2568 6806
rect 1597 6797 1599 6800
rect 1621 6797 1623 6800
rect 2542 6797 2544 6800
rect 2566 6797 2568 6800
rect 1473 6760 1475 6762
rect 1489 6760 1491 6765
rect 1494 6760 1496 6762
rect 1510 6760 1512 6762
rect 1526 6760 1528 6765
rect 1547 6760 1549 6765
rect 1552 6760 1554 6762
rect 1568 6760 1570 6762
rect 1584 6760 1586 6763
rect 1589 6760 1591 6762
rect 1605 6760 1607 6762
rect 1621 6760 1623 6765
rect 1626 6760 1628 6762
rect 1642 6760 1644 6762
rect 1658 6760 1660 6765
rect 1679 6760 1681 6765
rect 1684 6760 1686 6762
rect 1700 6760 1702 6762
rect 1716 6760 1718 6763
rect 1721 6760 1723 6762
rect 1737 6760 1739 6762
rect 1753 6760 1755 6765
rect 1758 6760 1760 6762
rect 1774 6760 1776 6762
rect 1790 6760 1792 6765
rect 1811 6760 1813 6765
rect 1816 6760 1818 6762
rect 1832 6760 1834 6762
rect 1848 6760 1850 6763
rect 1853 6760 1855 6762
rect 2418 6760 2420 6762
rect 2434 6760 2436 6765
rect 2439 6760 2441 6762
rect 2455 6760 2457 6762
rect 2471 6760 2473 6765
rect 2492 6760 2494 6765
rect 2497 6760 2499 6762
rect 2513 6760 2515 6762
rect 2529 6760 2531 6763
rect 2534 6760 2536 6762
rect 2550 6760 2552 6762
rect 2566 6760 2568 6765
rect 2571 6760 2573 6762
rect 2587 6760 2589 6762
rect 2603 6760 2605 6765
rect 2624 6760 2626 6765
rect 2629 6760 2631 6762
rect 2645 6760 2647 6762
rect 2661 6760 2663 6763
rect 2666 6760 2668 6762
rect 2682 6760 2684 6762
rect 2698 6760 2700 6765
rect 2703 6760 2705 6762
rect 2719 6760 2721 6762
rect 2735 6760 2737 6765
rect 2756 6760 2758 6765
rect 2761 6760 2763 6762
rect 2777 6760 2779 6762
rect 2793 6760 2795 6763
rect 2798 6760 2800 6762
rect 1473 6749 1475 6756
rect 1489 6754 1491 6756
rect 1494 6753 1496 6756
rect 1473 6737 1475 6745
rect 1489 6737 1491 6739
rect 1494 6737 1496 6746
rect 1510 6744 1512 6756
rect 1526 6754 1528 6756
rect 1547 6754 1549 6756
rect 1552 6753 1554 6756
rect 1510 6737 1512 6740
rect 1526 6737 1528 6739
rect 1547 6737 1549 6739
rect 1552 6737 1554 6746
rect 1568 6737 1570 6756
rect 1584 6749 1586 6756
rect 1589 6744 1591 6756
rect 1584 6737 1586 6739
rect 1589 6737 1591 6740
rect 1605 6737 1607 6756
rect 1621 6754 1623 6756
rect 1626 6753 1628 6756
rect 1621 6737 1623 6739
rect 1626 6737 1628 6746
rect 1642 6744 1644 6756
rect 1658 6754 1660 6756
rect 1679 6754 1681 6756
rect 1684 6753 1686 6756
rect 1642 6737 1644 6740
rect 1658 6737 1660 6739
rect 1679 6737 1681 6739
rect 1684 6737 1686 6746
rect 1700 6737 1702 6756
rect 1716 6749 1718 6756
rect 1721 6744 1723 6756
rect 1716 6737 1718 6739
rect 1721 6737 1723 6740
rect 1737 6737 1739 6756
rect 1753 6754 1755 6756
rect 1758 6753 1760 6756
rect 1753 6737 1755 6739
rect 1758 6737 1760 6746
rect 1774 6744 1776 6756
rect 1790 6754 1792 6756
rect 1811 6754 1813 6756
rect 1816 6753 1818 6756
rect 1774 6737 1776 6740
rect 1790 6737 1792 6739
rect 1811 6737 1813 6739
rect 1816 6737 1818 6746
rect 1832 6737 1834 6756
rect 1848 6749 1850 6756
rect 1853 6746 1855 6756
rect 2418 6749 2420 6756
rect 2434 6754 2436 6756
rect 2439 6753 2441 6756
rect 1848 6737 1850 6739
rect 1853 6737 1855 6742
rect 954 6730 956 6732
rect 970 6730 972 6735
rect 975 6730 977 6732
rect 991 6730 993 6732
rect 1007 6730 1009 6735
rect 1028 6730 1030 6735
rect 1033 6730 1035 6732
rect 1049 6730 1051 6732
rect 1065 6730 1067 6733
rect 1070 6730 1072 6732
rect 2418 6737 2420 6745
rect 2434 6737 2436 6739
rect 2439 6737 2441 6746
rect 2455 6744 2457 6756
rect 2471 6754 2473 6756
rect 2492 6754 2494 6756
rect 2497 6753 2499 6756
rect 2455 6737 2457 6740
rect 2471 6737 2473 6739
rect 2492 6737 2494 6739
rect 2497 6737 2499 6746
rect 2513 6737 2515 6756
rect 2529 6749 2531 6756
rect 2534 6744 2536 6756
rect 2529 6737 2531 6739
rect 2534 6737 2536 6740
rect 2550 6737 2552 6756
rect 2566 6754 2568 6756
rect 2571 6753 2573 6756
rect 2566 6737 2568 6739
rect 2571 6737 2573 6746
rect 2587 6744 2589 6756
rect 2603 6754 2605 6756
rect 2624 6754 2626 6756
rect 2629 6753 2631 6756
rect 2587 6737 2589 6740
rect 2603 6737 2605 6739
rect 2624 6737 2626 6739
rect 2629 6737 2631 6746
rect 2645 6737 2647 6756
rect 2661 6749 2663 6756
rect 2666 6744 2668 6756
rect 2661 6737 2663 6739
rect 2666 6737 2668 6740
rect 2682 6737 2684 6756
rect 2698 6754 2700 6756
rect 2703 6753 2705 6756
rect 2698 6737 2700 6739
rect 2703 6737 2705 6746
rect 2719 6744 2721 6756
rect 2735 6754 2737 6756
rect 2756 6754 2758 6756
rect 2761 6753 2763 6756
rect 2719 6737 2721 6740
rect 2735 6737 2737 6739
rect 2756 6737 2758 6739
rect 2761 6737 2763 6746
rect 2777 6737 2779 6756
rect 2793 6749 2795 6756
rect 2798 6746 2800 6756
rect 2793 6737 2795 6739
rect 2798 6737 2800 6742
rect 1899 6730 1901 6732
rect 1915 6730 1917 6735
rect 1920 6730 1922 6732
rect 1936 6730 1938 6732
rect 1952 6730 1954 6735
rect 1973 6730 1975 6735
rect 1978 6730 1980 6732
rect 1994 6730 1996 6732
rect 2010 6730 2012 6733
rect 2015 6730 2017 6732
rect 1473 6727 1475 6729
rect 1489 6726 1491 6729
rect 1494 6727 1496 6729
rect 1510 6726 1512 6729
rect 1526 6726 1528 6729
rect 1547 6726 1549 6729
rect 1552 6727 1554 6729
rect 1568 6727 1570 6729
rect 1584 6726 1586 6729
rect 1589 6727 1591 6729
rect 1605 6727 1607 6729
rect 1621 6726 1623 6729
rect 1626 6727 1628 6729
rect 1642 6726 1644 6729
rect 1658 6726 1660 6729
rect 1679 6726 1681 6729
rect 1684 6727 1686 6729
rect 1700 6727 1702 6729
rect 1716 6726 1718 6729
rect 1721 6727 1723 6729
rect 1737 6727 1739 6729
rect 1753 6726 1755 6729
rect 1758 6727 1760 6729
rect 1774 6726 1776 6729
rect 1790 6726 1792 6729
rect 1811 6726 1813 6729
rect 1816 6727 1818 6729
rect 1832 6727 1834 6729
rect 1848 6726 1850 6729
rect 1853 6727 1855 6729
rect 2418 6727 2420 6729
rect 2434 6726 2436 6729
rect 2439 6727 2441 6729
rect 2455 6726 2457 6729
rect 2471 6726 2473 6729
rect 2492 6726 2494 6729
rect 2497 6727 2499 6729
rect 2513 6727 2515 6729
rect 2529 6726 2531 6729
rect 2534 6727 2536 6729
rect 2550 6727 2552 6729
rect 2566 6726 2568 6729
rect 2571 6727 2573 6729
rect 2587 6726 2589 6729
rect 2603 6726 2605 6729
rect 2624 6726 2626 6729
rect 2629 6727 2631 6729
rect 2645 6727 2647 6729
rect 2661 6726 2663 6729
rect 2666 6727 2668 6729
rect 2682 6727 2684 6729
rect 2698 6726 2700 6729
rect 2703 6727 2705 6729
rect 2719 6726 2721 6729
rect 2735 6726 2737 6729
rect 2756 6726 2758 6729
rect 2761 6727 2763 6729
rect 2777 6727 2779 6729
rect 2793 6726 2795 6729
rect 2798 6727 2800 6729
rect 924 6718 927 6720
rect 931 6718 934 6720
rect 954 6707 956 6726
rect 970 6724 972 6726
rect 975 6723 977 6726
rect 970 6707 972 6709
rect 975 6707 977 6716
rect 991 6714 993 6726
rect 1007 6724 1009 6726
rect 1028 6724 1030 6726
rect 1033 6723 1035 6726
rect 991 6707 993 6710
rect 1007 6707 1009 6709
rect 1028 6707 1030 6709
rect 1033 6707 1035 6716
rect 1049 6707 1051 6726
rect 1065 6719 1067 6726
rect 1070 6716 1072 6726
rect 1869 6718 1872 6720
rect 1876 6718 1879 6720
rect 1065 6707 1067 6709
rect 1070 6707 1072 6712
rect 1899 6707 1901 6726
rect 1915 6724 1917 6726
rect 1920 6723 1922 6726
rect 1915 6707 1917 6709
rect 1920 6707 1922 6716
rect 1936 6714 1938 6726
rect 1952 6724 1954 6726
rect 1973 6724 1975 6726
rect 1978 6723 1980 6726
rect 1936 6707 1938 6710
rect 1952 6707 1954 6709
rect 1973 6707 1975 6709
rect 1978 6707 1980 6716
rect 1994 6707 1996 6726
rect 2010 6719 2012 6726
rect 2015 6716 2017 6726
rect 2010 6707 2012 6709
rect 2015 6707 2017 6712
rect 954 6697 956 6699
rect 970 6696 972 6699
rect 975 6697 977 6699
rect 991 6696 993 6699
rect 1007 6696 1009 6699
rect 1028 6696 1030 6699
rect 1033 6697 1035 6699
rect 1049 6697 1051 6699
rect 1065 6696 1067 6699
rect 1070 6697 1072 6699
rect 1899 6697 1901 6699
rect 1915 6696 1917 6699
rect 1920 6697 1922 6699
rect 1936 6696 1938 6699
rect 1952 6696 1954 6699
rect 1973 6696 1975 6699
rect 1978 6697 1980 6699
rect 1994 6697 1996 6699
rect 2010 6696 2012 6699
rect 2015 6697 2017 6699
rect 1473 6674 1475 6676
rect 1489 6674 1491 6679
rect 1494 6674 1496 6676
rect 1510 6674 1512 6676
rect 1526 6674 1528 6679
rect 1547 6674 1549 6679
rect 1552 6674 1554 6676
rect 1568 6674 1570 6676
rect 1584 6674 1586 6677
rect 1589 6674 1591 6676
rect 1605 6674 1607 6676
rect 1621 6674 1623 6679
rect 1626 6674 1628 6676
rect 1642 6674 1644 6676
rect 1658 6674 1660 6679
rect 1679 6674 1681 6679
rect 1684 6674 1686 6676
rect 1700 6674 1702 6676
rect 1716 6674 1718 6677
rect 1721 6674 1723 6676
rect 1737 6674 1739 6676
rect 1753 6674 1755 6679
rect 1758 6674 1760 6676
rect 1774 6674 1776 6676
rect 1790 6674 1792 6679
rect 1811 6674 1813 6679
rect 1816 6674 1818 6676
rect 1832 6674 1834 6676
rect 1848 6674 1850 6677
rect 1853 6674 1855 6676
rect 2418 6674 2420 6676
rect 2434 6674 2436 6679
rect 2439 6674 2441 6676
rect 2455 6674 2457 6676
rect 2471 6674 2473 6679
rect 2492 6674 2494 6679
rect 2497 6674 2499 6676
rect 2513 6674 2515 6676
rect 2529 6674 2531 6677
rect 2534 6674 2536 6676
rect 2550 6674 2552 6676
rect 2566 6674 2568 6679
rect 2571 6674 2573 6676
rect 2587 6674 2589 6676
rect 2603 6674 2605 6679
rect 2624 6674 2626 6679
rect 2629 6674 2631 6676
rect 2645 6674 2647 6676
rect 2661 6674 2663 6677
rect 2666 6674 2668 6676
rect 2682 6674 2684 6676
rect 2698 6674 2700 6679
rect 2703 6674 2705 6676
rect 2719 6674 2721 6676
rect 2735 6674 2737 6679
rect 2756 6674 2758 6679
rect 2761 6674 2763 6676
rect 2777 6674 2779 6676
rect 2793 6674 2795 6677
rect 2798 6674 2800 6676
rect 1473 6663 1475 6670
rect 1489 6668 1491 6670
rect 1494 6667 1496 6670
rect 1473 6651 1475 6659
rect 1489 6651 1491 6653
rect 1494 6651 1496 6660
rect 1510 6658 1512 6670
rect 1526 6668 1528 6670
rect 1547 6668 1549 6670
rect 1552 6667 1554 6670
rect 1510 6651 1512 6654
rect 1526 6651 1528 6653
rect 1547 6651 1549 6653
rect 1552 6651 1554 6660
rect 1568 6651 1570 6670
rect 1584 6663 1586 6670
rect 1589 6658 1591 6670
rect 1584 6651 1586 6653
rect 1589 6651 1591 6654
rect 1605 6651 1607 6670
rect 1621 6668 1623 6670
rect 1626 6667 1628 6670
rect 1621 6651 1623 6653
rect 1626 6651 1628 6660
rect 1642 6658 1644 6670
rect 1658 6668 1660 6670
rect 1679 6668 1681 6670
rect 1684 6667 1686 6670
rect 1642 6651 1644 6654
rect 1658 6651 1660 6653
rect 1679 6651 1681 6653
rect 1684 6651 1686 6660
rect 1700 6651 1702 6670
rect 1716 6663 1718 6670
rect 1721 6658 1723 6670
rect 1716 6651 1718 6653
rect 1721 6651 1723 6654
rect 1737 6651 1739 6670
rect 1753 6668 1755 6670
rect 1758 6667 1760 6670
rect 1753 6651 1755 6653
rect 1758 6651 1760 6660
rect 1774 6658 1776 6670
rect 1790 6668 1792 6670
rect 1811 6668 1813 6670
rect 1816 6667 1818 6670
rect 1774 6651 1776 6654
rect 1790 6651 1792 6653
rect 1811 6651 1813 6653
rect 1816 6651 1818 6660
rect 1832 6651 1834 6670
rect 1848 6663 1850 6670
rect 1853 6660 1855 6670
rect 2418 6663 2420 6670
rect 2434 6668 2436 6670
rect 2439 6667 2441 6670
rect 1848 6651 1850 6653
rect 1853 6651 1855 6656
rect 954 6644 956 6646
rect 970 6644 972 6649
rect 975 6644 977 6646
rect 991 6644 993 6646
rect 1007 6644 1009 6649
rect 1028 6644 1030 6649
rect 1033 6644 1035 6646
rect 1049 6644 1051 6646
rect 1065 6644 1067 6647
rect 1070 6644 1072 6646
rect 2418 6651 2420 6659
rect 2434 6651 2436 6653
rect 2439 6651 2441 6660
rect 2455 6658 2457 6670
rect 2471 6668 2473 6670
rect 2492 6668 2494 6670
rect 2497 6667 2499 6670
rect 2455 6651 2457 6654
rect 2471 6651 2473 6653
rect 2492 6651 2494 6653
rect 2497 6651 2499 6660
rect 2513 6651 2515 6670
rect 2529 6663 2531 6670
rect 2534 6658 2536 6670
rect 2529 6651 2531 6653
rect 2534 6651 2536 6654
rect 2550 6651 2552 6670
rect 2566 6668 2568 6670
rect 2571 6667 2573 6670
rect 2566 6651 2568 6653
rect 2571 6651 2573 6660
rect 2587 6658 2589 6670
rect 2603 6668 2605 6670
rect 2624 6668 2626 6670
rect 2629 6667 2631 6670
rect 2587 6651 2589 6654
rect 2603 6651 2605 6653
rect 2624 6651 2626 6653
rect 2629 6651 2631 6660
rect 2645 6651 2647 6670
rect 2661 6663 2663 6670
rect 2666 6658 2668 6670
rect 2661 6651 2663 6653
rect 2666 6651 2668 6654
rect 2682 6651 2684 6670
rect 2698 6668 2700 6670
rect 2703 6667 2705 6670
rect 2698 6651 2700 6653
rect 2703 6651 2705 6660
rect 2719 6658 2721 6670
rect 2735 6668 2737 6670
rect 2756 6668 2758 6670
rect 2761 6667 2763 6670
rect 2719 6651 2721 6654
rect 2735 6651 2737 6653
rect 2756 6651 2758 6653
rect 2761 6651 2763 6660
rect 2777 6651 2779 6670
rect 2793 6663 2795 6670
rect 2798 6660 2800 6670
rect 2793 6651 2795 6653
rect 2798 6651 2800 6656
rect 1899 6644 1901 6646
rect 1915 6644 1917 6649
rect 1920 6644 1922 6646
rect 1936 6644 1938 6646
rect 1952 6644 1954 6649
rect 1973 6644 1975 6649
rect 1978 6644 1980 6646
rect 1994 6644 1996 6646
rect 2010 6644 2012 6647
rect 2015 6644 2017 6646
rect 1473 6641 1475 6643
rect 1489 6640 1491 6643
rect 1494 6641 1496 6643
rect 1510 6640 1512 6643
rect 1526 6640 1528 6643
rect 1547 6640 1549 6643
rect 1552 6641 1554 6643
rect 1568 6641 1570 6643
rect 1584 6640 1586 6643
rect 1589 6641 1591 6643
rect 1605 6641 1607 6643
rect 1621 6640 1623 6643
rect 1626 6641 1628 6643
rect 1642 6640 1644 6643
rect 1658 6640 1660 6643
rect 1679 6640 1681 6643
rect 1684 6641 1686 6643
rect 1700 6641 1702 6643
rect 1716 6640 1718 6643
rect 1721 6641 1723 6643
rect 1737 6641 1739 6643
rect 1753 6640 1755 6643
rect 1758 6641 1760 6643
rect 1774 6640 1776 6643
rect 1790 6640 1792 6643
rect 1811 6640 1813 6643
rect 1816 6641 1818 6643
rect 1832 6641 1834 6643
rect 1848 6640 1850 6643
rect 1853 6641 1855 6643
rect 2418 6641 2420 6643
rect 2434 6640 2436 6643
rect 2439 6641 2441 6643
rect 2455 6640 2457 6643
rect 2471 6640 2473 6643
rect 2492 6640 2494 6643
rect 2497 6641 2499 6643
rect 2513 6641 2515 6643
rect 2529 6640 2531 6643
rect 2534 6641 2536 6643
rect 2550 6641 2552 6643
rect 2566 6640 2568 6643
rect 2571 6641 2573 6643
rect 2587 6640 2589 6643
rect 2603 6640 2605 6643
rect 2624 6640 2626 6643
rect 2629 6641 2631 6643
rect 2645 6641 2647 6643
rect 2661 6640 2663 6643
rect 2666 6641 2668 6643
rect 2682 6641 2684 6643
rect 2698 6640 2700 6643
rect 2703 6641 2705 6643
rect 2719 6640 2721 6643
rect 2735 6640 2737 6643
rect 2756 6640 2758 6643
rect 2761 6641 2763 6643
rect 2777 6641 2779 6643
rect 2793 6640 2795 6643
rect 2798 6641 2800 6643
rect 954 6621 956 6640
rect 970 6638 972 6640
rect 975 6637 977 6640
rect 970 6621 972 6623
rect 975 6621 977 6630
rect 991 6628 993 6640
rect 1007 6638 1009 6640
rect 1028 6638 1030 6640
rect 1033 6637 1035 6640
rect 991 6621 993 6624
rect 1007 6621 1009 6623
rect 1028 6621 1030 6623
rect 1033 6621 1035 6630
rect 1049 6621 1051 6640
rect 1065 6633 1067 6640
rect 1070 6630 1072 6640
rect 1065 6621 1067 6623
rect 1070 6621 1072 6626
rect 1899 6621 1901 6640
rect 1915 6638 1917 6640
rect 1920 6637 1922 6640
rect 1915 6621 1917 6623
rect 1920 6621 1922 6630
rect 1936 6628 1938 6640
rect 1952 6638 1954 6640
rect 1973 6638 1975 6640
rect 1978 6637 1980 6640
rect 1936 6621 1938 6624
rect 1952 6621 1954 6623
rect 1973 6621 1975 6623
rect 1978 6621 1980 6630
rect 1994 6621 1996 6640
rect 2010 6633 2012 6640
rect 2015 6630 2017 6640
rect 2010 6621 2012 6623
rect 2015 6621 2017 6626
rect 954 6611 956 6613
rect 970 6610 972 6613
rect 975 6611 977 6613
rect 991 6610 993 6613
rect 1007 6610 1009 6613
rect 1028 6610 1030 6613
rect 1033 6611 1035 6613
rect 1049 6611 1051 6613
rect 1065 6610 1067 6613
rect 1070 6611 1072 6613
rect 1714 6612 1716 6615
rect 1738 6612 1740 6615
rect 1899 6611 1901 6613
rect 1915 6610 1917 6613
rect 1920 6611 1922 6613
rect 1936 6610 1938 6613
rect 1952 6610 1954 6613
rect 1973 6610 1975 6613
rect 1978 6611 1980 6613
rect 1994 6611 1996 6613
rect 2010 6610 2012 6613
rect 2015 6611 2017 6613
rect 2659 6612 2661 6615
rect 2683 6612 2685 6615
rect 1714 6606 1716 6608
rect 1738 6606 1740 6608
rect 2659 6606 2661 6608
rect 2683 6606 2685 6608
rect 1706 6601 1725 6603
rect 1729 6601 1731 6603
rect 2651 6601 2670 6603
rect 2674 6601 2676 6603
rect 1718 6589 1720 6592
rect 2663 6589 2665 6592
rect 1718 6583 1720 6585
rect 2663 6583 2665 6585
rect 936 6572 939 6574
rect 943 6572 946 6574
rect 971 6547 973 6550
rect 1017 6547 1019 6550
rect 1043 6547 1045 6550
rect 1087 6547 1089 6550
rect 1018 6543 1019 6547
rect 953 6540 955 6542
rect 971 6540 973 6543
rect 976 6540 978 6542
rect 996 6540 998 6543
rect 1017 6540 1019 6543
rect 1043 6540 1045 6543
rect 1048 6540 1050 6542
rect 1071 6540 1073 6542
rect 1087 6540 1089 6543
rect 1112 6540 1114 6578
rect 1714 6576 1716 6578
rect 1738 6576 1740 6578
rect 1881 6572 1884 6574
rect 1888 6572 1891 6574
rect 1714 6569 1716 6572
rect 1738 6569 1740 6572
rect 1159 6545 1161 6550
rect 1232 6547 1234 6550
rect 1278 6547 1280 6550
rect 1304 6547 1306 6550
rect 1348 6547 1350 6550
rect 1164 6545 1166 6547
rect 1130 6540 1132 6543
rect 1279 6543 1280 6547
rect 1916 6547 1918 6550
rect 1962 6547 1964 6550
rect 1988 6547 1990 6550
rect 2032 6547 2034 6550
rect 1963 6543 1964 6547
rect 1214 6540 1216 6542
rect 1232 6540 1234 6543
rect 1237 6540 1239 6542
rect 1257 6540 1259 6543
rect 1278 6540 1280 6543
rect 1304 6540 1306 6543
rect 1309 6540 1311 6542
rect 1332 6540 1334 6542
rect 1348 6540 1350 6543
rect 1364 6540 1366 6542
rect 1159 6535 1161 6537
rect 953 6518 955 6532
rect 971 6530 973 6532
rect 976 6527 978 6532
rect 976 6523 982 6527
rect 971 6518 973 6520
rect 976 6518 978 6523
rect 996 6518 998 6532
rect 1017 6530 1019 6532
rect 1043 6530 1045 6532
rect 1048 6527 1050 6532
rect 1048 6523 1054 6527
rect 1017 6518 1019 6520
rect 1043 6518 1045 6520
rect 1048 6518 1050 6523
rect 1071 6518 1073 6532
rect 1087 6530 1089 6532
rect 1087 6518 1089 6520
rect 1112 6518 1114 6532
rect 1130 6527 1132 6532
rect 1159 6525 1161 6527
rect 1164 6525 1166 6537
rect 1473 6532 1475 6534
rect 1489 6532 1491 6537
rect 1494 6532 1496 6534
rect 1510 6532 1512 6534
rect 1526 6532 1528 6537
rect 1547 6532 1549 6537
rect 1552 6532 1554 6534
rect 1568 6532 1570 6534
rect 1584 6532 1586 6535
rect 1589 6532 1591 6534
rect 1605 6532 1607 6534
rect 1621 6532 1623 6537
rect 1626 6532 1628 6534
rect 1642 6532 1644 6534
rect 1658 6532 1660 6537
rect 1679 6532 1681 6537
rect 1684 6532 1686 6534
rect 1700 6532 1702 6534
rect 1716 6532 1718 6535
rect 1898 6540 1900 6542
rect 1916 6540 1918 6543
rect 1921 6540 1923 6542
rect 1941 6540 1943 6543
rect 1962 6540 1964 6543
rect 1988 6540 1990 6543
rect 1993 6540 1995 6542
rect 2016 6540 2018 6542
rect 2032 6540 2034 6543
rect 2057 6540 2059 6582
rect 2659 6576 2661 6578
rect 2683 6576 2685 6578
rect 2659 6569 2661 6572
rect 2683 6569 2685 6572
rect 2104 6545 2106 6550
rect 2177 6547 2179 6550
rect 2223 6547 2225 6550
rect 2249 6547 2251 6550
rect 2293 6547 2295 6550
rect 2109 6545 2111 6547
rect 2075 6540 2077 6543
rect 1721 6532 1723 6534
rect 1737 6532 1739 6534
rect 1753 6532 1755 6537
rect 1758 6532 1760 6534
rect 1774 6532 1776 6534
rect 1790 6532 1792 6537
rect 1811 6532 1813 6537
rect 1816 6532 1818 6534
rect 1832 6532 1834 6534
rect 1848 6532 1850 6535
rect 1853 6532 1855 6534
rect 2224 6543 2225 6547
rect 2159 6540 2161 6542
rect 2177 6540 2179 6543
rect 2182 6540 2184 6542
rect 2202 6540 2204 6543
rect 2223 6540 2225 6543
rect 2249 6540 2251 6543
rect 2254 6540 2256 6542
rect 2277 6540 2279 6542
rect 2293 6540 2295 6543
rect 2309 6540 2311 6542
rect 2104 6535 2106 6537
rect 1130 6518 1132 6523
rect 1159 6518 1161 6521
rect 1164 6518 1166 6521
rect 1214 6518 1216 6532
rect 1232 6530 1234 6532
rect 1237 6527 1239 6532
rect 1237 6523 1243 6527
rect 1232 6518 1234 6520
rect 1237 6518 1239 6523
rect 1257 6518 1259 6532
rect 1278 6530 1280 6532
rect 1304 6530 1306 6532
rect 1309 6527 1311 6532
rect 1309 6523 1315 6527
rect 1278 6518 1280 6520
rect 1304 6518 1306 6520
rect 1309 6518 1311 6523
rect 1332 6518 1334 6532
rect 1348 6530 1350 6532
rect 1348 6518 1350 6520
rect 1364 6518 1366 6532
rect 1473 6521 1475 6528
rect 1489 6526 1491 6528
rect 1494 6525 1496 6528
rect 953 6512 955 6514
rect 971 6509 973 6514
rect 976 6512 978 6514
rect 996 6512 998 6514
rect 1017 6510 1019 6514
rect 971 6505 972 6509
rect 1017 6506 1018 6510
rect 1043 6509 1045 6514
rect 1048 6512 1050 6514
rect 1071 6512 1073 6514
rect 1087 6510 1089 6514
rect 1112 6511 1114 6514
rect 1130 6511 1132 6514
rect 1214 6512 1216 6514
rect 971 6503 973 6505
rect 1017 6502 1019 6506
rect 1043 6505 1044 6509
rect 1087 6506 1088 6510
rect 1232 6509 1234 6514
rect 1237 6512 1239 6514
rect 1257 6512 1259 6514
rect 1278 6510 1280 6514
rect 1043 6503 1045 6505
rect 1087 6503 1089 6506
rect 1232 6505 1233 6509
rect 1278 6506 1279 6510
rect 1304 6509 1306 6514
rect 1309 6512 1311 6514
rect 1332 6512 1334 6514
rect 1348 6510 1350 6514
rect 1364 6512 1366 6514
rect 1232 6503 1234 6505
rect 1278 6502 1280 6506
rect 1304 6505 1305 6509
rect 1348 6506 1349 6510
rect 1473 6509 1475 6517
rect 1489 6509 1491 6511
rect 1494 6509 1496 6518
rect 1510 6516 1512 6528
rect 1526 6526 1528 6528
rect 1547 6526 1549 6528
rect 1552 6525 1554 6528
rect 1510 6509 1512 6512
rect 1526 6509 1528 6511
rect 1547 6509 1549 6511
rect 1552 6509 1554 6518
rect 1568 6509 1570 6528
rect 1584 6521 1586 6528
rect 1589 6516 1591 6528
rect 1584 6509 1586 6511
rect 1589 6509 1591 6512
rect 1605 6509 1607 6528
rect 1621 6526 1623 6528
rect 1626 6525 1628 6528
rect 1621 6509 1623 6511
rect 1626 6509 1628 6518
rect 1642 6516 1644 6528
rect 1658 6526 1660 6528
rect 1679 6526 1681 6528
rect 1684 6525 1686 6528
rect 1642 6509 1644 6512
rect 1658 6509 1660 6511
rect 1679 6509 1681 6511
rect 1684 6509 1686 6518
rect 1700 6509 1702 6528
rect 1716 6521 1718 6528
rect 1721 6516 1723 6528
rect 1716 6509 1718 6511
rect 1721 6509 1723 6512
rect 1737 6509 1739 6528
rect 1753 6526 1755 6528
rect 1758 6525 1760 6528
rect 1753 6509 1755 6511
rect 1758 6509 1760 6518
rect 1774 6516 1776 6528
rect 1790 6526 1792 6528
rect 1811 6526 1813 6528
rect 1816 6525 1818 6528
rect 1774 6509 1776 6512
rect 1790 6509 1792 6511
rect 1811 6509 1813 6511
rect 1816 6509 1818 6518
rect 1832 6509 1834 6528
rect 1848 6521 1850 6528
rect 1853 6518 1855 6528
rect 1898 6518 1900 6532
rect 1916 6530 1918 6532
rect 1921 6527 1923 6532
rect 1921 6523 1927 6527
rect 1916 6518 1918 6520
rect 1921 6518 1923 6523
rect 1941 6518 1943 6532
rect 1962 6530 1964 6532
rect 1988 6530 1990 6532
rect 1993 6527 1995 6532
rect 1993 6523 1999 6527
rect 1962 6518 1964 6520
rect 1988 6518 1990 6520
rect 1993 6518 1995 6523
rect 2016 6518 2018 6532
rect 2032 6530 2034 6532
rect 2032 6518 2034 6520
rect 2057 6518 2059 6532
rect 2075 6527 2077 6532
rect 2104 6525 2106 6527
rect 2109 6525 2111 6537
rect 2418 6532 2420 6534
rect 2434 6532 2436 6537
rect 2439 6532 2441 6534
rect 2455 6532 2457 6534
rect 2471 6532 2473 6537
rect 2492 6532 2494 6537
rect 2497 6532 2499 6534
rect 2513 6532 2515 6534
rect 2529 6532 2531 6535
rect 2534 6532 2536 6534
rect 2550 6532 2552 6534
rect 2566 6532 2568 6537
rect 2571 6532 2573 6534
rect 2587 6532 2589 6534
rect 2603 6532 2605 6537
rect 2624 6532 2626 6537
rect 2629 6532 2631 6534
rect 2645 6532 2647 6534
rect 2661 6532 2663 6535
rect 2666 6532 2668 6534
rect 2682 6532 2684 6534
rect 2698 6532 2700 6537
rect 2703 6532 2705 6534
rect 2719 6532 2721 6534
rect 2735 6532 2737 6537
rect 2756 6532 2758 6537
rect 2761 6532 2763 6534
rect 2777 6532 2779 6534
rect 2793 6532 2795 6535
rect 2798 6532 2800 6534
rect 2075 6518 2077 6523
rect 2104 6518 2106 6521
rect 2109 6518 2111 6521
rect 2159 6518 2161 6532
rect 2177 6530 2179 6532
rect 2182 6527 2184 6532
rect 2182 6523 2188 6527
rect 2177 6518 2179 6520
rect 2182 6518 2184 6523
rect 2202 6518 2204 6532
rect 2223 6530 2225 6532
rect 2249 6530 2251 6532
rect 2254 6527 2256 6532
rect 2254 6523 2260 6527
rect 2223 6518 2225 6520
rect 2249 6518 2251 6520
rect 2254 6518 2256 6523
rect 2277 6518 2279 6532
rect 2293 6530 2295 6532
rect 2293 6518 2295 6520
rect 2309 6518 2311 6532
rect 2418 6521 2420 6528
rect 2434 6526 2436 6528
rect 2439 6525 2441 6528
rect 1848 6509 1850 6511
rect 1853 6509 1855 6514
rect 1898 6512 1900 6514
rect 1916 6509 1918 6514
rect 1921 6512 1923 6514
rect 1941 6512 1943 6514
rect 1962 6510 1964 6514
rect 1304 6503 1306 6505
rect 1348 6503 1350 6506
rect 1916 6505 1917 6509
rect 1962 6506 1963 6510
rect 1988 6509 1990 6514
rect 1993 6512 1995 6514
rect 2016 6512 2018 6514
rect 2032 6510 2034 6514
rect 2057 6511 2059 6514
rect 2075 6511 2077 6514
rect 2159 6512 2161 6514
rect 1916 6503 1918 6505
rect 1962 6502 1964 6506
rect 1988 6505 1989 6509
rect 2032 6506 2033 6510
rect 2177 6509 2179 6514
rect 2182 6512 2184 6514
rect 2202 6512 2204 6514
rect 2223 6510 2225 6514
rect 1988 6503 1990 6505
rect 2032 6503 2034 6506
rect 2177 6505 2178 6509
rect 2223 6506 2224 6510
rect 2249 6509 2251 6514
rect 2254 6512 2256 6514
rect 2277 6512 2279 6514
rect 2293 6510 2295 6514
rect 2309 6512 2311 6514
rect 2177 6503 2179 6505
rect 2223 6502 2225 6506
rect 2249 6505 2250 6509
rect 2293 6506 2294 6510
rect 2418 6509 2420 6517
rect 2434 6509 2436 6511
rect 2439 6509 2441 6518
rect 2455 6516 2457 6528
rect 2471 6526 2473 6528
rect 2492 6526 2494 6528
rect 2497 6525 2499 6528
rect 2455 6509 2457 6512
rect 2471 6509 2473 6511
rect 2492 6509 2494 6511
rect 2497 6509 2499 6518
rect 2513 6509 2515 6528
rect 2529 6521 2531 6528
rect 2534 6516 2536 6528
rect 2529 6509 2531 6511
rect 2534 6509 2536 6512
rect 2550 6509 2552 6528
rect 2566 6526 2568 6528
rect 2571 6525 2573 6528
rect 2566 6509 2568 6511
rect 2571 6509 2573 6518
rect 2587 6516 2589 6528
rect 2603 6526 2605 6528
rect 2624 6526 2626 6528
rect 2629 6525 2631 6528
rect 2587 6509 2589 6512
rect 2603 6509 2605 6511
rect 2624 6509 2626 6511
rect 2629 6509 2631 6518
rect 2645 6509 2647 6528
rect 2661 6521 2663 6528
rect 2666 6516 2668 6528
rect 2661 6509 2663 6511
rect 2666 6509 2668 6512
rect 2682 6509 2684 6528
rect 2698 6526 2700 6528
rect 2703 6525 2705 6528
rect 2698 6509 2700 6511
rect 2703 6509 2705 6518
rect 2719 6516 2721 6528
rect 2735 6526 2737 6528
rect 2756 6526 2758 6528
rect 2761 6525 2763 6528
rect 2719 6509 2721 6512
rect 2735 6509 2737 6511
rect 2756 6509 2758 6511
rect 2761 6509 2763 6518
rect 2777 6509 2779 6528
rect 2793 6521 2795 6528
rect 2798 6518 2800 6528
rect 2793 6509 2795 6511
rect 2798 6509 2800 6514
rect 2249 6503 2251 6505
rect 2293 6503 2295 6506
rect 1473 6499 1475 6501
rect 1489 6498 1491 6501
rect 1494 6499 1496 6501
rect 1510 6498 1512 6501
rect 1526 6498 1528 6501
rect 1547 6498 1549 6501
rect 1552 6499 1554 6501
rect 1568 6499 1570 6501
rect 1584 6498 1586 6501
rect 1589 6499 1591 6501
rect 1605 6499 1607 6501
rect 1621 6498 1623 6501
rect 1626 6499 1628 6501
rect 1642 6498 1644 6501
rect 1658 6498 1660 6501
rect 1679 6498 1681 6501
rect 1684 6499 1686 6501
rect 1700 6499 1702 6501
rect 1716 6498 1718 6501
rect 1721 6499 1723 6501
rect 1737 6499 1739 6501
rect 1753 6498 1755 6501
rect 1758 6499 1760 6501
rect 1774 6498 1776 6501
rect 1790 6498 1792 6501
rect 1811 6498 1813 6501
rect 1816 6499 1818 6501
rect 1832 6499 1834 6501
rect 1848 6498 1850 6501
rect 1853 6499 1855 6501
rect 2418 6499 2420 6501
rect 2434 6498 2436 6501
rect 2439 6499 2441 6501
rect 2455 6498 2457 6501
rect 2471 6498 2473 6501
rect 2492 6498 2494 6501
rect 2497 6499 2499 6501
rect 2513 6499 2515 6501
rect 2529 6498 2531 6501
rect 2534 6499 2536 6501
rect 2550 6499 2552 6501
rect 2566 6498 2568 6501
rect 2571 6499 2573 6501
rect 2587 6498 2589 6501
rect 2603 6498 2605 6501
rect 2624 6498 2626 6501
rect 2629 6499 2631 6501
rect 2645 6499 2647 6501
rect 2661 6498 2663 6501
rect 2666 6499 2668 6501
rect 2682 6499 2684 6501
rect 2698 6498 2700 6501
rect 2703 6499 2705 6501
rect 2719 6498 2721 6501
rect 2735 6498 2737 6501
rect 2756 6498 2758 6501
rect 2761 6499 2763 6501
rect 2777 6499 2779 6501
rect 2793 6498 2795 6501
rect 2798 6499 2800 6501
rect 1232 6481 1234 6483
rect 1232 6477 1233 6481
rect 1278 6480 1280 6484
rect 1304 6481 1306 6483
rect 1214 6472 1216 6474
rect 1232 6472 1234 6477
rect 1278 6476 1279 6480
rect 1304 6477 1305 6481
rect 1348 6480 1350 6483
rect 2177 6481 2179 6483
rect 1237 6472 1239 6474
rect 1257 6472 1259 6474
rect 1278 6472 1280 6476
rect 1304 6472 1306 6477
rect 1348 6476 1349 6480
rect 2177 6477 2178 6481
rect 2223 6480 2225 6484
rect 2249 6481 2251 6483
rect 1309 6472 1311 6474
rect 1332 6472 1334 6474
rect 1348 6472 1350 6476
rect 1364 6472 1366 6474
rect 2159 6472 2161 6474
rect 2177 6472 2179 6477
rect 2223 6476 2224 6480
rect 2249 6477 2250 6481
rect 2293 6480 2295 6483
rect 2182 6472 2184 6474
rect 2202 6472 2204 6474
rect 2223 6472 2225 6476
rect 2249 6472 2251 6477
rect 2293 6476 2294 6480
rect 2254 6472 2256 6474
rect 2277 6472 2279 6474
rect 2293 6472 2295 6476
rect 2309 6472 2311 6474
rect 1136 6467 1138 6469
rect 1159 6463 1161 6468
rect 1164 6463 1166 6465
rect 1136 6441 1138 6463
rect 1159 6457 1161 6459
rect 1164 6454 1166 6459
rect 1214 6454 1216 6468
rect 1232 6466 1234 6468
rect 1237 6463 1239 6468
rect 1237 6459 1243 6463
rect 1232 6454 1234 6456
rect 1237 6454 1239 6459
rect 1257 6454 1259 6468
rect 1278 6466 1280 6468
rect 1304 6466 1306 6468
rect 1309 6463 1311 6468
rect 1309 6459 1315 6463
rect 1278 6454 1280 6456
rect 1304 6454 1306 6456
rect 1309 6454 1311 6459
rect 1332 6454 1334 6468
rect 1348 6466 1350 6468
rect 1348 6454 1350 6456
rect 1364 6454 1366 6468
rect 2081 6467 2083 6469
rect 2104 6463 2106 6468
rect 2109 6463 2111 6465
rect 1164 6450 1165 6454
rect 1159 6447 1161 6449
rect 1164 6447 1166 6450
rect 1214 6444 1216 6446
rect 1232 6443 1234 6446
rect 1237 6444 1239 6446
rect 1257 6443 1259 6446
rect 1278 6443 1280 6446
rect 1304 6443 1306 6446
rect 1309 6444 1311 6446
rect 1332 6444 1334 6446
rect 1348 6443 1350 6446
rect 1364 6444 1366 6446
rect 1279 6439 1280 6443
rect 2081 6441 2083 6463
rect 2104 6457 2106 6459
rect 2109 6454 2111 6459
rect 2159 6454 2161 6468
rect 2177 6466 2179 6468
rect 2182 6463 2184 6468
rect 2182 6459 2188 6463
rect 2177 6454 2179 6456
rect 2182 6454 2184 6459
rect 2202 6454 2204 6468
rect 2223 6466 2225 6468
rect 2249 6466 2251 6468
rect 2254 6463 2256 6468
rect 2254 6459 2260 6463
rect 2223 6454 2225 6456
rect 2249 6454 2251 6456
rect 2254 6454 2256 6459
rect 2277 6454 2279 6468
rect 2293 6466 2295 6468
rect 2293 6454 2295 6456
rect 2309 6454 2311 6468
rect 2109 6450 2110 6454
rect 2104 6447 2106 6449
rect 2109 6447 2111 6450
rect 1159 6436 1161 6439
rect 1136 6431 1138 6433
rect 1164 6435 1166 6439
rect 1232 6436 1234 6439
rect 1278 6436 1280 6439
rect 1304 6436 1306 6439
rect 1348 6436 1350 6439
rect 2159 6444 2161 6446
rect 2177 6443 2179 6446
rect 2182 6444 2184 6446
rect 2202 6443 2204 6446
rect 2223 6443 2225 6446
rect 2249 6443 2251 6446
rect 2254 6444 2256 6446
rect 2277 6444 2279 6446
rect 2293 6443 2295 6446
rect 2309 6444 2311 6446
rect 2224 6439 2225 6443
rect 2104 6436 2106 6439
rect 2081 6431 2083 6433
rect 2109 6435 2111 6439
rect 2177 6436 2179 6439
rect 2223 6436 2225 6439
rect 2249 6436 2251 6439
rect 2293 6436 2295 6439
rect 1232 6415 1234 6418
rect 1278 6415 1280 6418
rect 1304 6415 1306 6418
rect 1348 6415 1350 6418
rect 988 6409 990 6414
rect 993 6409 995 6411
rect 1078 6409 1080 6414
rect 1083 6409 1085 6411
rect 1159 6409 1161 6414
rect 1279 6411 1280 6415
rect 1164 6409 1166 6411
rect 1214 6408 1216 6410
rect 1232 6408 1234 6411
rect 1237 6408 1239 6410
rect 1257 6408 1259 6411
rect 1278 6408 1280 6411
rect 1304 6408 1306 6411
rect 1309 6408 1311 6410
rect 1332 6408 1334 6410
rect 1348 6408 1350 6411
rect 2177 6415 2179 6418
rect 2223 6415 2225 6418
rect 2249 6415 2251 6418
rect 2293 6415 2295 6418
rect 1364 6408 1366 6410
rect 1933 6409 1935 6414
rect 1938 6409 1940 6411
rect 2023 6409 2025 6414
rect 2028 6409 2030 6411
rect 2104 6409 2106 6414
rect 2224 6411 2225 6415
rect 2109 6409 2111 6411
rect 988 6399 990 6401
rect 988 6389 990 6391
rect 993 6389 995 6401
rect 1078 6399 1080 6401
rect 1078 6389 1080 6391
rect 1083 6389 1085 6401
rect 1159 6399 1161 6401
rect 1159 6389 1161 6391
rect 1164 6389 1166 6401
rect 2159 6408 2161 6410
rect 2177 6408 2179 6411
rect 2182 6408 2184 6410
rect 2202 6408 2204 6411
rect 2223 6408 2225 6411
rect 2249 6408 2251 6411
rect 2254 6408 2256 6410
rect 2277 6408 2279 6410
rect 2293 6408 2295 6411
rect 2309 6408 2311 6410
rect 1214 6386 1216 6400
rect 1232 6398 1234 6400
rect 1237 6395 1239 6400
rect 1237 6391 1243 6395
rect 1232 6386 1234 6388
rect 1237 6386 1239 6391
rect 1257 6386 1259 6400
rect 1278 6398 1280 6400
rect 1304 6398 1306 6400
rect 1309 6395 1311 6400
rect 1309 6391 1315 6395
rect 1278 6386 1280 6388
rect 1304 6386 1306 6388
rect 1309 6386 1311 6391
rect 1332 6386 1334 6400
rect 1348 6398 1350 6400
rect 1348 6386 1350 6388
rect 1364 6386 1366 6400
rect 1933 6399 1935 6401
rect 1933 6389 1935 6391
rect 1938 6389 1940 6401
rect 2023 6399 2025 6401
rect 2023 6389 2025 6391
rect 2028 6389 2030 6401
rect 2104 6399 2106 6401
rect 2104 6389 2106 6391
rect 2109 6389 2111 6401
rect 988 6382 990 6385
rect 993 6382 995 6385
rect 1078 6382 1080 6385
rect 1083 6382 1085 6385
rect 1159 6382 1161 6385
rect 1164 6382 1166 6385
rect 2159 6386 2161 6400
rect 2177 6398 2179 6400
rect 2182 6395 2184 6400
rect 2182 6391 2188 6395
rect 2177 6386 2179 6388
rect 2182 6386 2184 6391
rect 2202 6386 2204 6400
rect 2223 6398 2225 6400
rect 2249 6398 2251 6400
rect 2254 6395 2256 6400
rect 2254 6391 2260 6395
rect 2223 6386 2225 6388
rect 2249 6386 2251 6388
rect 2254 6386 2256 6391
rect 2277 6386 2279 6400
rect 2293 6398 2295 6400
rect 2293 6386 2295 6388
rect 2309 6386 2311 6400
rect 1933 6382 1935 6385
rect 1938 6382 1940 6385
rect 2023 6382 2025 6385
rect 2028 6382 2030 6385
rect 2104 6382 2106 6385
rect 2109 6382 2111 6385
rect 1214 6380 1216 6382
rect 1232 6377 1234 6382
rect 1237 6380 1239 6382
rect 1257 6380 1259 6382
rect 1278 6378 1280 6382
rect 1232 6373 1233 6377
rect 1278 6374 1279 6378
rect 1304 6377 1306 6382
rect 1309 6380 1311 6382
rect 1332 6380 1334 6382
rect 1348 6378 1350 6382
rect 1364 6380 1366 6382
rect 2159 6380 2161 6382
rect 1232 6371 1234 6373
rect 1278 6370 1280 6374
rect 1304 6373 1305 6377
rect 1348 6374 1349 6378
rect 2177 6377 2179 6382
rect 2182 6380 2184 6382
rect 2202 6380 2204 6382
rect 2223 6378 2225 6382
rect 1304 6371 1306 6373
rect 1348 6371 1350 6374
rect 2177 6373 2178 6377
rect 2223 6374 2224 6378
rect 2249 6377 2251 6382
rect 2254 6380 2256 6382
rect 2277 6380 2279 6382
rect 2293 6378 2295 6382
rect 2309 6380 2311 6382
rect 2177 6371 2179 6373
rect 2223 6370 2225 6374
rect 2249 6373 2250 6377
rect 2293 6374 2294 6378
rect 2249 6371 2251 6373
rect 2293 6371 2295 6374
rect 1232 6349 1234 6351
rect 1232 6345 1233 6349
rect 1278 6348 1280 6352
rect 1304 6349 1306 6351
rect 1214 6340 1216 6342
rect 1232 6340 1234 6345
rect 1278 6344 1279 6348
rect 1304 6345 1305 6349
rect 1348 6348 1350 6351
rect 2177 6349 2179 6351
rect 1237 6340 1239 6342
rect 1257 6340 1259 6342
rect 1278 6340 1280 6344
rect 1304 6340 1306 6345
rect 1348 6344 1349 6348
rect 2177 6345 2178 6349
rect 2223 6348 2225 6352
rect 2249 6349 2251 6351
rect 1309 6340 1311 6342
rect 1332 6340 1334 6342
rect 1348 6340 1350 6344
rect 1364 6340 1366 6342
rect 2159 6340 2161 6342
rect 2177 6340 2179 6345
rect 2223 6344 2224 6348
rect 2249 6345 2250 6349
rect 2293 6348 2295 6351
rect 2182 6340 2184 6342
rect 2202 6340 2204 6342
rect 2223 6340 2225 6344
rect 2249 6340 2251 6345
rect 2293 6344 2294 6348
rect 2254 6340 2256 6342
rect 2277 6340 2279 6342
rect 2293 6340 2295 6344
rect 2309 6340 2311 6342
rect 965 6335 967 6337
rect 988 6331 990 6336
rect 1055 6335 1057 6337
rect 993 6331 995 6333
rect 1078 6331 1080 6336
rect 1136 6335 1138 6337
rect 1083 6331 1085 6333
rect 1159 6331 1161 6336
rect 1164 6331 1166 6333
rect 965 6309 967 6331
rect 1019 6327 1021 6329
rect 988 6325 990 6327
rect 993 6322 995 6327
rect 993 6318 994 6322
rect 988 6315 990 6317
rect 993 6315 995 6318
rect 1019 6309 1021 6323
rect 1055 6309 1057 6331
rect 1109 6327 1111 6329
rect 1078 6325 1080 6327
rect 1083 6322 1085 6327
rect 1083 6318 1084 6322
rect 1078 6315 1080 6317
rect 1083 6315 1085 6318
rect 988 6304 990 6307
rect 965 6299 967 6301
rect 993 6303 995 6307
rect 1109 6309 1111 6323
rect 1136 6309 1138 6331
rect 1159 6325 1161 6327
rect 1164 6322 1166 6327
rect 1214 6322 1216 6336
rect 1232 6334 1234 6336
rect 1237 6331 1239 6336
rect 1237 6327 1243 6331
rect 1232 6322 1234 6324
rect 1237 6322 1239 6327
rect 1257 6322 1259 6336
rect 1278 6334 1280 6336
rect 1304 6334 1306 6336
rect 1309 6331 1311 6336
rect 1309 6327 1315 6331
rect 1278 6322 1280 6324
rect 1304 6322 1306 6324
rect 1309 6322 1311 6327
rect 1332 6322 1334 6336
rect 1348 6334 1350 6336
rect 1348 6322 1350 6324
rect 1364 6322 1366 6336
rect 1910 6335 1912 6337
rect 1933 6331 1935 6336
rect 2000 6335 2002 6337
rect 1938 6331 1940 6333
rect 2023 6331 2025 6336
rect 2081 6335 2083 6337
rect 2028 6331 2030 6333
rect 2104 6331 2106 6336
rect 2109 6331 2111 6333
rect 1164 6318 1165 6322
rect 1159 6315 1161 6317
rect 1164 6315 1166 6318
rect 1078 6304 1080 6307
rect 1019 6299 1021 6301
rect 1055 6299 1057 6301
rect 1083 6303 1085 6307
rect 1214 6312 1216 6314
rect 1232 6311 1234 6314
rect 1237 6312 1239 6314
rect 1257 6311 1259 6314
rect 1278 6311 1280 6314
rect 1304 6311 1306 6314
rect 1309 6312 1311 6314
rect 1332 6312 1334 6314
rect 1348 6311 1350 6314
rect 1364 6312 1366 6314
rect 1279 6307 1280 6311
rect 1910 6309 1912 6331
rect 1964 6327 1966 6329
rect 1933 6325 1935 6327
rect 1938 6322 1940 6327
rect 1938 6318 1939 6322
rect 1933 6315 1935 6317
rect 1938 6315 1940 6318
rect 1159 6304 1161 6307
rect 1109 6299 1111 6301
rect 1136 6299 1138 6301
rect 1164 6303 1166 6307
rect 1232 6304 1234 6307
rect 1278 6304 1280 6307
rect 1304 6304 1306 6307
rect 1348 6304 1350 6307
rect 1964 6309 1966 6323
rect 2000 6309 2002 6331
rect 2054 6327 2056 6329
rect 2023 6325 2025 6327
rect 2028 6322 2030 6327
rect 2028 6318 2029 6322
rect 2023 6315 2025 6317
rect 2028 6315 2030 6318
rect 1933 6304 1935 6307
rect 1910 6299 1912 6301
rect 1938 6303 1940 6307
rect 2054 6309 2056 6323
rect 2081 6309 2083 6331
rect 2104 6325 2106 6327
rect 2109 6322 2111 6327
rect 2159 6322 2161 6336
rect 2177 6334 2179 6336
rect 2182 6331 2184 6336
rect 2182 6327 2188 6331
rect 2177 6322 2179 6324
rect 2182 6322 2184 6327
rect 2202 6322 2204 6336
rect 2223 6334 2225 6336
rect 2249 6334 2251 6336
rect 2254 6331 2256 6336
rect 2254 6327 2260 6331
rect 2223 6322 2225 6324
rect 2249 6322 2251 6324
rect 2254 6322 2256 6327
rect 2277 6322 2279 6336
rect 2293 6334 2295 6336
rect 2293 6322 2295 6324
rect 2309 6322 2311 6336
rect 2109 6318 2110 6322
rect 2104 6315 2106 6317
rect 2109 6315 2111 6318
rect 2023 6304 2025 6307
rect 1964 6299 1966 6301
rect 2000 6299 2002 6301
rect 2028 6303 2030 6307
rect 2159 6312 2161 6314
rect 2177 6311 2179 6314
rect 2182 6312 2184 6314
rect 2202 6311 2204 6314
rect 2223 6311 2225 6314
rect 2249 6311 2251 6314
rect 2254 6312 2256 6314
rect 2277 6312 2279 6314
rect 2293 6311 2295 6314
rect 2309 6312 2311 6314
rect 2224 6307 2225 6311
rect 2104 6304 2106 6307
rect 2054 6299 2056 6301
rect 2081 6299 2083 6301
rect 2109 6303 2111 6307
rect 2177 6304 2179 6307
rect 2223 6304 2225 6307
rect 2249 6304 2251 6307
rect 2293 6304 2295 6307
rect 1232 6283 1234 6286
rect 1278 6283 1280 6286
rect 1304 6283 1306 6286
rect 1348 6283 1350 6286
rect 2177 6283 2179 6286
rect 2223 6283 2225 6286
rect 2249 6283 2251 6286
rect 2293 6283 2295 6286
rect 1279 6279 1280 6283
rect 1054 6274 1056 6279
rect 1059 6274 1061 6276
rect 1159 6274 1161 6279
rect 1214 6276 1216 6278
rect 1232 6276 1234 6279
rect 1237 6276 1239 6278
rect 1257 6276 1259 6279
rect 1278 6276 1280 6279
rect 1304 6276 1306 6279
rect 1309 6276 1311 6278
rect 1332 6276 1334 6278
rect 1348 6276 1350 6279
rect 2224 6279 2225 6283
rect 1364 6276 1366 6278
rect 1164 6274 1166 6276
rect 1999 6274 2001 6279
rect 2004 6274 2006 6276
rect 2104 6274 2106 6279
rect 2159 6276 2161 6278
rect 2177 6276 2179 6279
rect 2182 6276 2184 6278
rect 2202 6276 2204 6279
rect 2223 6276 2225 6279
rect 2249 6276 2251 6279
rect 2254 6276 2256 6278
rect 2277 6276 2279 6278
rect 2293 6276 2295 6279
rect 2309 6276 2311 6278
rect 2109 6274 2111 6276
rect 1054 6264 1056 6266
rect 1054 6254 1056 6256
rect 1059 6254 1061 6266
rect 1159 6264 1161 6266
rect 1159 6254 1161 6256
rect 1164 6254 1166 6266
rect 1214 6254 1216 6268
rect 1232 6266 1234 6268
rect 1237 6263 1239 6268
rect 1237 6259 1243 6263
rect 1232 6254 1234 6256
rect 1237 6254 1239 6259
rect 1257 6254 1259 6268
rect 1278 6266 1280 6268
rect 1304 6266 1306 6268
rect 1309 6263 1311 6268
rect 1309 6259 1315 6263
rect 1278 6254 1280 6256
rect 1304 6254 1306 6256
rect 1309 6254 1311 6259
rect 1332 6254 1334 6268
rect 1348 6266 1350 6268
rect 1348 6254 1350 6256
rect 1364 6254 1366 6268
rect 1999 6264 2001 6266
rect 1999 6254 2001 6256
rect 2004 6254 2006 6266
rect 2104 6264 2106 6266
rect 2104 6254 2106 6256
rect 2109 6254 2111 6266
rect 2159 6254 2161 6268
rect 2177 6266 2179 6268
rect 2182 6263 2184 6268
rect 2182 6259 2188 6263
rect 2177 6254 2179 6256
rect 2182 6254 2184 6259
rect 2202 6254 2204 6268
rect 2223 6266 2225 6268
rect 2249 6266 2251 6268
rect 2254 6263 2256 6268
rect 2254 6259 2260 6263
rect 2223 6254 2225 6256
rect 2249 6254 2251 6256
rect 2254 6254 2256 6259
rect 2277 6254 2279 6268
rect 2293 6266 2295 6268
rect 2293 6254 2295 6256
rect 2309 6254 2311 6268
rect 1054 6247 1056 6250
rect 1059 6247 1061 6250
rect 1159 6247 1161 6250
rect 1164 6247 1166 6250
rect 1214 6248 1216 6250
rect 1232 6245 1234 6250
rect 1237 6248 1239 6250
rect 1257 6248 1259 6250
rect 1278 6246 1280 6250
rect 1232 6241 1233 6245
rect 1278 6242 1279 6246
rect 1304 6245 1306 6250
rect 1309 6248 1311 6250
rect 1332 6248 1334 6250
rect 1348 6246 1350 6250
rect 1364 6248 1366 6250
rect 1999 6247 2001 6250
rect 2004 6247 2006 6250
rect 2104 6247 2106 6250
rect 2109 6247 2111 6250
rect 2159 6248 2161 6250
rect 1232 6239 1234 6241
rect 1278 6238 1280 6242
rect 1304 6241 1305 6245
rect 1348 6242 1349 6246
rect 2177 6245 2179 6250
rect 2182 6248 2184 6250
rect 2202 6248 2204 6250
rect 2223 6246 2225 6250
rect 1304 6239 1306 6241
rect 1348 6239 1350 6242
rect 2177 6241 2178 6245
rect 2223 6242 2224 6246
rect 2249 6245 2251 6250
rect 2254 6248 2256 6250
rect 2277 6248 2279 6250
rect 2293 6246 2295 6250
rect 2309 6248 2311 6250
rect 2177 6239 2179 6241
rect 2223 6238 2225 6242
rect 2249 6241 2250 6245
rect 2293 6242 2294 6246
rect 2249 6239 2251 6241
rect 2293 6239 2295 6242
rect 1232 6217 1234 6219
rect 1232 6213 1233 6217
rect 1278 6216 1280 6220
rect 1304 6217 1306 6219
rect 1214 6208 1216 6210
rect 1232 6208 1234 6213
rect 1278 6212 1279 6216
rect 1304 6213 1305 6217
rect 1348 6216 1350 6219
rect 2177 6217 2179 6219
rect 1237 6208 1239 6210
rect 1257 6208 1259 6210
rect 1278 6208 1280 6212
rect 1304 6208 1306 6213
rect 1348 6212 1349 6216
rect 2177 6213 2178 6217
rect 2223 6216 2225 6220
rect 2249 6217 2251 6219
rect 1309 6208 1311 6210
rect 1332 6208 1334 6210
rect 1348 6208 1350 6212
rect 1364 6208 1366 6210
rect 2159 6208 2161 6210
rect 2177 6208 2179 6213
rect 2223 6212 2224 6216
rect 2249 6213 2250 6217
rect 2293 6216 2295 6219
rect 2182 6208 2184 6210
rect 2202 6208 2204 6210
rect 2223 6208 2225 6212
rect 2249 6208 2251 6213
rect 2293 6212 2294 6216
rect 2254 6208 2256 6210
rect 2277 6208 2279 6210
rect 2293 6208 2295 6212
rect 2309 6208 2311 6210
rect 1031 6203 1033 6205
rect 1054 6199 1056 6204
rect 1136 6203 1138 6205
rect 1059 6199 1061 6201
rect 1159 6199 1161 6204
rect 1164 6199 1166 6201
rect 1031 6177 1033 6199
rect 1085 6195 1087 6197
rect 1054 6193 1056 6195
rect 1059 6190 1061 6195
rect 1059 6186 1060 6190
rect 1054 6183 1056 6185
rect 1059 6183 1061 6186
rect 1085 6177 1087 6191
rect 1136 6177 1138 6199
rect 1159 6193 1161 6195
rect 1164 6190 1166 6195
rect 1214 6190 1216 6204
rect 1232 6202 1234 6204
rect 1237 6199 1239 6204
rect 1237 6195 1243 6199
rect 1232 6190 1234 6192
rect 1237 6190 1239 6195
rect 1257 6190 1259 6204
rect 1278 6202 1280 6204
rect 1304 6202 1306 6204
rect 1309 6199 1311 6204
rect 1309 6195 1315 6199
rect 1278 6190 1280 6192
rect 1304 6190 1306 6192
rect 1309 6190 1311 6195
rect 1332 6190 1334 6204
rect 1348 6202 1350 6204
rect 1348 6190 1350 6192
rect 1364 6190 1366 6204
rect 1976 6203 1978 6205
rect 1999 6199 2001 6204
rect 2081 6203 2083 6205
rect 2004 6199 2006 6201
rect 2104 6199 2106 6204
rect 2109 6199 2111 6201
rect 1164 6186 1165 6190
rect 1159 6183 1161 6185
rect 1164 6183 1166 6186
rect 1054 6172 1056 6175
rect 1031 6167 1033 6169
rect 1059 6171 1061 6175
rect 1214 6180 1216 6182
rect 1232 6179 1234 6182
rect 1237 6180 1239 6182
rect 1257 6179 1259 6182
rect 1278 6179 1280 6182
rect 1304 6179 1306 6182
rect 1309 6180 1311 6182
rect 1332 6180 1334 6182
rect 1348 6179 1350 6182
rect 1364 6180 1366 6182
rect 1279 6175 1280 6179
rect 1976 6177 1978 6199
rect 2030 6195 2032 6197
rect 1999 6193 2001 6195
rect 2004 6190 2006 6195
rect 2004 6186 2005 6190
rect 1999 6183 2001 6185
rect 2004 6183 2006 6186
rect 1159 6172 1161 6175
rect 1085 6167 1087 6169
rect 1136 6167 1138 6169
rect 1164 6171 1166 6175
rect 1232 6172 1234 6175
rect 1278 6172 1280 6175
rect 1304 6172 1306 6175
rect 1348 6172 1350 6175
rect 2030 6177 2032 6191
rect 2081 6177 2083 6199
rect 2104 6193 2106 6195
rect 2109 6190 2111 6195
rect 2159 6190 2161 6204
rect 2177 6202 2179 6204
rect 2182 6199 2184 6204
rect 2182 6195 2188 6199
rect 2177 6190 2179 6192
rect 2182 6190 2184 6195
rect 2202 6190 2204 6204
rect 2223 6202 2225 6204
rect 2249 6202 2251 6204
rect 2254 6199 2256 6204
rect 2254 6195 2260 6199
rect 2223 6190 2225 6192
rect 2249 6190 2251 6192
rect 2254 6190 2256 6195
rect 2277 6190 2279 6204
rect 2293 6202 2295 6204
rect 2293 6190 2295 6192
rect 2309 6190 2311 6204
rect 2109 6186 2110 6190
rect 2104 6183 2106 6185
rect 2109 6183 2111 6186
rect 1999 6172 2001 6175
rect 1976 6167 1978 6169
rect 2004 6171 2006 6175
rect 2159 6180 2161 6182
rect 2177 6179 2179 6182
rect 2182 6180 2184 6182
rect 2202 6179 2204 6182
rect 2223 6179 2225 6182
rect 2249 6179 2251 6182
rect 2254 6180 2256 6182
rect 2277 6180 2279 6182
rect 2293 6179 2295 6182
rect 2309 6180 2311 6182
rect 2224 6175 2225 6179
rect 2104 6172 2106 6175
rect 2030 6167 2032 6169
rect 2081 6167 2083 6169
rect 2109 6171 2111 6175
rect 2177 6172 2179 6175
rect 2223 6172 2225 6175
rect 2249 6172 2251 6175
rect 2293 6172 2295 6175
rect 1232 6151 1234 6154
rect 1278 6151 1280 6154
rect 1304 6151 1306 6154
rect 1348 6151 1350 6154
rect 1078 6143 1080 6148
rect 1083 6143 1085 6145
rect 1159 6143 1161 6148
rect 1279 6147 1280 6151
rect 2177 6151 2179 6154
rect 2223 6151 2225 6154
rect 2249 6151 2251 6154
rect 2293 6151 2295 6154
rect 1164 6143 1166 6145
rect 1214 6144 1216 6146
rect 1232 6144 1234 6147
rect 1237 6144 1239 6146
rect 1257 6144 1259 6147
rect 1278 6144 1280 6147
rect 1304 6144 1306 6147
rect 1309 6144 1311 6146
rect 1332 6144 1334 6146
rect 1348 6144 1350 6147
rect 1364 6144 1366 6146
rect 2023 6143 2025 6148
rect 2028 6143 2030 6145
rect 2104 6143 2106 6148
rect 2224 6147 2225 6151
rect 2109 6143 2111 6145
rect 2159 6144 2161 6146
rect 2177 6144 2179 6147
rect 2182 6144 2184 6146
rect 2202 6144 2204 6147
rect 2223 6144 2225 6147
rect 2249 6144 2251 6147
rect 2254 6144 2256 6146
rect 2277 6144 2279 6146
rect 2293 6144 2295 6147
rect 2309 6144 2311 6146
rect 1078 6133 1080 6135
rect 1078 6123 1080 6125
rect 1083 6123 1085 6135
rect 1159 6133 1161 6135
rect 1159 6123 1161 6125
rect 1164 6123 1166 6135
rect 1214 6122 1216 6136
rect 1232 6134 1234 6136
rect 1237 6131 1239 6136
rect 1237 6127 1243 6131
rect 1232 6122 1234 6124
rect 1237 6122 1239 6127
rect 1257 6122 1259 6136
rect 1278 6134 1280 6136
rect 1304 6134 1306 6136
rect 1309 6131 1311 6136
rect 1309 6127 1315 6131
rect 1278 6122 1280 6124
rect 1304 6122 1306 6124
rect 1309 6122 1311 6127
rect 1332 6122 1334 6136
rect 1348 6134 1350 6136
rect 1348 6122 1350 6124
rect 1364 6122 1366 6136
rect 1614 6132 1616 6134
rect 1619 6132 1621 6135
rect 1635 6132 1637 6134
rect 1651 6132 1653 6134
rect 1656 6132 1658 6137
rect 1677 6132 1679 6137
rect 1693 6132 1695 6134
rect 1709 6132 1711 6134
rect 1714 6132 1716 6137
rect 1730 6132 1732 6134
rect 2023 6133 2025 6135
rect 1078 6116 1080 6119
rect 1083 6116 1085 6119
rect 1159 6116 1161 6119
rect 1164 6116 1166 6119
rect 1614 6118 1616 6128
rect 1619 6121 1621 6128
rect 1214 6116 1216 6118
rect 1232 6113 1234 6118
rect 1237 6116 1239 6118
rect 1257 6116 1259 6118
rect 1278 6114 1280 6118
rect 1232 6109 1233 6113
rect 1278 6110 1279 6114
rect 1304 6113 1306 6118
rect 1309 6116 1311 6118
rect 1332 6116 1334 6118
rect 1348 6114 1350 6118
rect 1364 6116 1366 6118
rect 1232 6107 1234 6109
rect 1278 6106 1280 6110
rect 1304 6109 1305 6113
rect 1348 6110 1349 6114
rect 1304 6107 1306 6109
rect 1348 6107 1350 6110
rect 1614 6109 1616 6114
rect 1619 6109 1621 6111
rect 1635 6109 1637 6128
rect 1651 6125 1653 6128
rect 1656 6126 1658 6128
rect 1677 6126 1679 6128
rect 1651 6109 1653 6118
rect 1693 6116 1695 6128
rect 1709 6125 1711 6128
rect 1714 6126 1716 6128
rect 1656 6109 1658 6111
rect 1677 6109 1679 6111
rect 1693 6109 1695 6112
rect 1709 6109 1711 6118
rect 1714 6109 1716 6111
rect 1730 6109 1732 6128
rect 2023 6123 2025 6125
rect 2028 6123 2030 6135
rect 2104 6133 2106 6135
rect 2104 6123 2106 6125
rect 2109 6123 2111 6135
rect 2159 6122 2161 6136
rect 2177 6134 2179 6136
rect 2182 6131 2184 6136
rect 2182 6127 2188 6131
rect 2177 6122 2179 6124
rect 2182 6122 2184 6127
rect 2202 6122 2204 6136
rect 2223 6134 2225 6136
rect 2249 6134 2251 6136
rect 2254 6131 2256 6136
rect 2254 6127 2260 6131
rect 2223 6122 2225 6124
rect 2249 6122 2251 6124
rect 2254 6122 2256 6127
rect 2277 6122 2279 6136
rect 2293 6134 2295 6136
rect 2293 6122 2295 6124
rect 2309 6122 2311 6136
rect 2559 6132 2561 6134
rect 2564 6132 2566 6135
rect 2580 6132 2582 6134
rect 2596 6132 2598 6134
rect 2601 6132 2603 6137
rect 2622 6132 2624 6137
rect 2638 6132 2640 6134
rect 2654 6132 2656 6134
rect 2659 6132 2661 6137
rect 2675 6132 2677 6134
rect 2023 6116 2025 6119
rect 2028 6116 2030 6119
rect 2104 6116 2106 6119
rect 2109 6116 2111 6119
rect 2559 6118 2561 6128
rect 2564 6121 2566 6128
rect 2159 6116 2161 6118
rect 2177 6113 2179 6118
rect 2182 6116 2184 6118
rect 2202 6116 2204 6118
rect 2223 6114 2225 6118
rect 2177 6109 2178 6113
rect 2223 6110 2224 6114
rect 2249 6113 2251 6118
rect 2254 6116 2256 6118
rect 2277 6116 2279 6118
rect 2293 6114 2295 6118
rect 2309 6116 2311 6118
rect 2177 6107 2179 6109
rect 2223 6106 2225 6110
rect 2249 6109 2250 6113
rect 2293 6110 2294 6114
rect 2249 6107 2251 6109
rect 2293 6107 2295 6110
rect 2559 6109 2561 6114
rect 2564 6109 2566 6111
rect 2580 6109 2582 6128
rect 2596 6125 2598 6128
rect 2601 6126 2603 6128
rect 2622 6126 2624 6128
rect 2596 6109 2598 6118
rect 2638 6116 2640 6128
rect 2654 6125 2656 6128
rect 2659 6126 2661 6128
rect 2601 6109 2603 6111
rect 2622 6109 2624 6111
rect 2638 6109 2640 6112
rect 2654 6109 2656 6118
rect 2659 6109 2661 6111
rect 2675 6109 2677 6128
rect 1614 6099 1616 6101
rect 1619 6098 1621 6101
rect 1635 6099 1637 6101
rect 1651 6099 1653 6101
rect 1656 6098 1658 6101
rect 1677 6098 1679 6101
rect 1693 6098 1695 6101
rect 1709 6099 1711 6101
rect 1714 6098 1716 6101
rect 1730 6099 1732 6101
rect 2559 6099 2561 6101
rect 2564 6098 2566 6101
rect 2580 6099 2582 6101
rect 2596 6099 2598 6101
rect 2601 6098 2603 6101
rect 2622 6098 2624 6101
rect 2638 6098 2640 6101
rect 2654 6099 2656 6101
rect 2659 6098 2661 6101
rect 2675 6099 2677 6101
rect 1232 6085 1234 6087
rect 1232 6081 1233 6085
rect 1278 6084 1280 6088
rect 1304 6085 1306 6087
rect 1214 6076 1216 6078
rect 1232 6076 1234 6081
rect 1278 6080 1279 6084
rect 1304 6081 1305 6085
rect 1348 6084 1350 6087
rect 2177 6085 2179 6087
rect 1237 6076 1239 6078
rect 1257 6076 1259 6078
rect 1278 6076 1280 6080
rect 1304 6076 1306 6081
rect 1348 6080 1349 6084
rect 2177 6081 2178 6085
rect 2223 6084 2225 6088
rect 2249 6085 2251 6087
rect 1309 6076 1311 6078
rect 1332 6076 1334 6078
rect 1348 6076 1350 6080
rect 1364 6076 1366 6078
rect 1714 6076 1716 6078
rect 2159 6076 2161 6078
rect 2177 6076 2179 6081
rect 2223 6080 2224 6084
rect 2249 6081 2250 6085
rect 2293 6084 2295 6087
rect 2182 6076 2184 6078
rect 2202 6076 2204 6078
rect 2223 6076 2225 6080
rect 2249 6076 2251 6081
rect 2293 6080 2294 6084
rect 2254 6076 2256 6078
rect 2277 6076 2279 6078
rect 2293 6076 2295 6080
rect 2309 6076 2311 6078
rect 2659 6076 2661 6078
rect 1055 6071 1057 6073
rect 1078 6067 1080 6072
rect 1136 6071 1138 6073
rect 1083 6067 1085 6069
rect 1159 6067 1161 6072
rect 1164 6067 1166 6069
rect 1055 6045 1057 6067
rect 1109 6063 1111 6065
rect 1078 6061 1080 6063
rect 1083 6058 1085 6063
rect 1083 6054 1084 6058
rect 1078 6051 1080 6053
rect 1083 6051 1085 6054
rect 1109 6045 1111 6059
rect 1136 6045 1138 6067
rect 1190 6063 1192 6065
rect 1159 6061 1161 6063
rect 1164 6058 1166 6063
rect 1164 6054 1165 6058
rect 1159 6051 1161 6053
rect 1164 6051 1166 6054
rect 1078 6040 1080 6043
rect 1055 6035 1057 6037
rect 1083 6039 1085 6043
rect 1190 6045 1192 6059
rect 1214 6058 1216 6072
rect 1232 6070 1234 6072
rect 1237 6067 1239 6072
rect 1237 6063 1243 6067
rect 1232 6058 1234 6060
rect 1237 6058 1239 6063
rect 1257 6058 1259 6072
rect 1278 6070 1280 6072
rect 1304 6070 1306 6072
rect 1309 6067 1311 6072
rect 1309 6063 1315 6067
rect 1278 6058 1280 6060
rect 1304 6058 1306 6060
rect 1309 6058 1311 6063
rect 1332 6058 1334 6072
rect 1348 6070 1350 6072
rect 1348 6058 1350 6060
rect 1364 6058 1366 6072
rect 1714 6069 1716 6072
rect 2000 6071 2002 6073
rect 1597 6067 1599 6069
rect 2023 6067 2025 6072
rect 2081 6071 2083 6073
rect 2028 6067 2030 6069
rect 2104 6067 2106 6072
rect 2109 6067 2111 6069
rect 1597 6060 1599 6063
rect 1214 6048 1216 6050
rect 1232 6047 1234 6050
rect 1237 6048 1239 6050
rect 1257 6047 1259 6050
rect 1278 6047 1280 6050
rect 1304 6047 1306 6050
rect 1309 6048 1311 6050
rect 1332 6048 1334 6050
rect 1348 6047 1350 6050
rect 1364 6048 1366 6050
rect 1159 6040 1161 6043
rect 1109 6035 1111 6037
rect 1136 6035 1138 6037
rect 1164 6039 1166 6043
rect 1279 6043 1280 6047
rect 1232 6040 1234 6043
rect 1278 6040 1280 6043
rect 1304 6040 1306 6043
rect 1348 6040 1350 6043
rect 2000 6045 2002 6067
rect 2054 6063 2056 6065
rect 2023 6061 2025 6063
rect 2028 6058 2030 6063
rect 2028 6054 2029 6058
rect 2023 6051 2025 6053
rect 2028 6051 2030 6054
rect 1190 6035 1192 6037
rect 2054 6045 2056 6059
rect 2081 6045 2083 6067
rect 2135 6063 2137 6065
rect 2104 6061 2106 6063
rect 2109 6058 2111 6063
rect 2109 6054 2110 6058
rect 2104 6051 2106 6053
rect 2109 6051 2111 6054
rect 2023 6040 2025 6043
rect 1605 6030 1607 6032
rect 1621 6030 1623 6035
rect 1626 6030 1628 6032
rect 1642 6030 1644 6032
rect 1658 6030 1660 6035
rect 1679 6030 1681 6035
rect 2000 6035 2002 6037
rect 2028 6039 2030 6043
rect 2135 6045 2137 6059
rect 2159 6058 2161 6072
rect 2177 6070 2179 6072
rect 2182 6067 2184 6072
rect 2182 6063 2188 6067
rect 2177 6058 2179 6060
rect 2182 6058 2184 6063
rect 2202 6058 2204 6072
rect 2223 6070 2225 6072
rect 2249 6070 2251 6072
rect 2254 6067 2256 6072
rect 2254 6063 2260 6067
rect 2223 6058 2225 6060
rect 2249 6058 2251 6060
rect 2254 6058 2256 6063
rect 2277 6058 2279 6072
rect 2293 6070 2295 6072
rect 2293 6058 2295 6060
rect 2309 6058 2311 6072
rect 2659 6069 2661 6072
rect 2542 6067 2544 6069
rect 2542 6060 2544 6063
rect 2159 6048 2161 6050
rect 2177 6047 2179 6050
rect 2182 6048 2184 6050
rect 2202 6047 2204 6050
rect 2223 6047 2225 6050
rect 2249 6047 2251 6050
rect 2254 6048 2256 6050
rect 2277 6048 2279 6050
rect 2293 6047 2295 6050
rect 2309 6048 2311 6050
rect 2104 6040 2106 6043
rect 2054 6035 2056 6037
rect 2081 6035 2083 6037
rect 2109 6039 2111 6043
rect 2224 6043 2225 6047
rect 2177 6040 2179 6043
rect 2223 6040 2225 6043
rect 2249 6040 2251 6043
rect 2293 6040 2295 6043
rect 2135 6035 2137 6037
rect 1684 6030 1686 6032
rect 1700 6030 1702 6032
rect 1716 6030 1718 6033
rect 1721 6030 1723 6032
rect 2550 6030 2552 6032
rect 2566 6030 2568 6035
rect 2571 6030 2573 6032
rect 2587 6030 2589 6032
rect 2603 6030 2605 6035
rect 2624 6030 2626 6035
rect 2629 6030 2631 6032
rect 2645 6030 2647 6032
rect 2661 6030 2663 6033
rect 2666 6030 2668 6032
rect 1605 6007 1607 6026
rect 1621 6024 1623 6026
rect 1626 6023 1628 6026
rect 1621 6007 1623 6009
rect 1626 6007 1628 6016
rect 1642 6014 1644 6026
rect 1658 6024 1660 6026
rect 1679 6024 1681 6026
rect 1684 6023 1686 6026
rect 1642 6007 1644 6010
rect 1658 6007 1660 6009
rect 1679 6007 1681 6009
rect 1684 6007 1686 6016
rect 1700 6007 1702 6026
rect 1716 6019 1718 6026
rect 1721 6016 1723 6026
rect 1716 6007 1718 6009
rect 1721 6007 1723 6012
rect 2550 6007 2552 6026
rect 2566 6024 2568 6026
rect 2571 6023 2573 6026
rect 2566 6007 2568 6009
rect 2571 6007 2573 6016
rect 2587 6014 2589 6026
rect 2603 6024 2605 6026
rect 2624 6024 2626 6026
rect 2629 6023 2631 6026
rect 2587 6007 2589 6010
rect 2603 6007 2605 6009
rect 2624 6007 2626 6009
rect 2629 6007 2631 6016
rect 2645 6007 2647 6026
rect 2661 6019 2663 6026
rect 2666 6016 2668 6026
rect 2661 6007 2663 6009
rect 2666 6007 2668 6012
rect 857 5997 859 5999
rect 873 5997 875 6002
rect 878 5997 880 5999
rect 894 5997 896 5999
rect 910 5997 912 6002
rect 931 5997 933 6002
rect 936 5997 938 5999
rect 952 5997 954 5999
rect 968 5997 970 6000
rect 973 5997 975 5999
rect 989 5997 991 5999
rect 1005 5997 1007 6002
rect 1010 5997 1012 5999
rect 1026 5997 1028 5999
rect 1042 5997 1044 6002
rect 1063 5997 1065 6002
rect 1068 5997 1070 5999
rect 1084 5997 1086 5999
rect 1100 5997 1102 6000
rect 1105 5997 1107 5999
rect 1121 5997 1123 5999
rect 1137 5997 1139 6002
rect 1142 5997 1144 5999
rect 1158 5997 1160 5999
rect 1174 5997 1176 6002
rect 1195 5997 1197 6002
rect 1200 5997 1202 5999
rect 1216 5997 1218 5999
rect 1232 5997 1234 6000
rect 1237 5997 1239 5999
rect 1253 5997 1255 5999
rect 1269 5997 1271 6002
rect 1274 5997 1276 5999
rect 1290 5997 1292 5999
rect 1306 5997 1308 6002
rect 1327 5997 1329 6002
rect 1332 5997 1334 5999
rect 1348 5997 1350 5999
rect 1364 5997 1366 6000
rect 1369 5997 1371 5999
rect 1605 5997 1607 5999
rect 1621 5996 1623 5999
rect 1626 5997 1628 5999
rect 1642 5996 1644 5999
rect 1658 5996 1660 5999
rect 1679 5996 1681 5999
rect 1684 5997 1686 5999
rect 1700 5997 1702 5999
rect 1716 5996 1718 5999
rect 1721 5997 1723 5999
rect 1802 5997 1804 5999
rect 1818 5997 1820 6002
rect 1823 5997 1825 5999
rect 1839 5997 1841 5999
rect 1855 5997 1857 6002
rect 1876 5997 1878 6002
rect 1881 5997 1883 5999
rect 1897 5997 1899 5999
rect 1913 5997 1915 6000
rect 1918 5997 1920 5999
rect 1934 5997 1936 5999
rect 1950 5997 1952 6002
rect 1955 5997 1957 5999
rect 1971 5997 1973 5999
rect 1987 5997 1989 6002
rect 2008 5997 2010 6002
rect 2013 5997 2015 5999
rect 2029 5997 2031 5999
rect 2045 5997 2047 6000
rect 2050 5997 2052 5999
rect 2066 5997 2068 5999
rect 2082 5997 2084 6002
rect 2087 5997 2089 5999
rect 2103 5997 2105 5999
rect 2119 5997 2121 6002
rect 2140 5997 2142 6002
rect 2145 5997 2147 5999
rect 2161 5997 2163 5999
rect 2177 5997 2179 6000
rect 2182 5997 2184 5999
rect 2198 5997 2200 5999
rect 2214 5997 2216 6002
rect 2219 5997 2221 5999
rect 2235 5997 2237 5999
rect 2251 5997 2253 6002
rect 2272 5997 2274 6002
rect 2277 5997 2279 5999
rect 2293 5997 2295 5999
rect 2309 5997 2311 6000
rect 2314 5997 2316 5999
rect 2550 5997 2552 5999
rect 857 5986 859 5993
rect 873 5991 875 5993
rect 878 5990 880 5993
rect 857 5974 859 5982
rect 873 5974 875 5976
rect 878 5974 880 5983
rect 894 5981 896 5993
rect 910 5991 912 5993
rect 931 5991 933 5993
rect 936 5990 938 5993
rect 894 5974 896 5977
rect 910 5974 912 5976
rect 931 5974 933 5976
rect 936 5974 938 5983
rect 952 5974 954 5993
rect 968 5986 970 5993
rect 973 5983 975 5993
rect 989 5986 991 5993
rect 1005 5991 1007 5993
rect 1010 5990 1012 5993
rect 968 5974 970 5976
rect 973 5974 975 5979
rect 989 5974 991 5982
rect 1005 5974 1007 5976
rect 1010 5974 1012 5983
rect 1026 5981 1028 5993
rect 1042 5991 1044 5993
rect 1063 5991 1065 5993
rect 1068 5990 1070 5993
rect 1026 5974 1028 5977
rect 1042 5974 1044 5976
rect 1063 5974 1065 5976
rect 1068 5974 1070 5983
rect 1084 5974 1086 5993
rect 1100 5986 1102 5993
rect 1105 5983 1107 5993
rect 1121 5986 1123 5993
rect 1137 5991 1139 5993
rect 1142 5990 1144 5993
rect 1100 5974 1102 5976
rect 1105 5974 1107 5979
rect 1121 5974 1123 5982
rect 1137 5974 1139 5976
rect 1142 5974 1144 5983
rect 1158 5981 1160 5993
rect 1174 5991 1176 5993
rect 1195 5991 1197 5993
rect 1200 5990 1202 5993
rect 1158 5974 1160 5977
rect 1174 5974 1176 5976
rect 1195 5974 1197 5976
rect 1200 5974 1202 5983
rect 1216 5974 1218 5993
rect 1232 5986 1234 5993
rect 1237 5983 1239 5993
rect 1253 5986 1255 5993
rect 1269 5991 1271 5993
rect 1274 5990 1276 5993
rect 1232 5974 1234 5976
rect 1237 5974 1239 5979
rect 1253 5974 1255 5982
rect 1269 5974 1271 5976
rect 1274 5974 1276 5983
rect 1290 5981 1292 5993
rect 1306 5991 1308 5993
rect 1327 5991 1329 5993
rect 1332 5990 1334 5993
rect 1290 5974 1292 5977
rect 1306 5974 1308 5976
rect 1327 5974 1329 5976
rect 1332 5974 1334 5983
rect 1348 5974 1350 5993
rect 1364 5986 1366 5993
rect 1369 5983 1371 5993
rect 2566 5996 2568 5999
rect 2571 5997 2573 5999
rect 2587 5996 2589 5999
rect 2603 5996 2605 5999
rect 2624 5996 2626 5999
rect 2629 5997 2631 5999
rect 2645 5997 2647 5999
rect 2661 5996 2663 5999
rect 2666 5997 2668 5999
rect 1802 5986 1804 5993
rect 1818 5991 1820 5993
rect 1823 5990 1825 5993
rect 1364 5974 1366 5976
rect 1369 5974 1371 5979
rect 1802 5974 1804 5982
rect 1818 5974 1820 5976
rect 1823 5974 1825 5983
rect 1839 5981 1841 5993
rect 1855 5991 1857 5993
rect 1876 5991 1878 5993
rect 1881 5990 1883 5993
rect 1839 5974 1841 5977
rect 1855 5974 1857 5976
rect 1876 5974 1878 5976
rect 1881 5974 1883 5983
rect 1897 5974 1899 5993
rect 1913 5986 1915 5993
rect 1918 5983 1920 5993
rect 1934 5986 1936 5993
rect 1950 5991 1952 5993
rect 1955 5990 1957 5993
rect 1913 5974 1915 5976
rect 1918 5974 1920 5979
rect 1934 5974 1936 5982
rect 1950 5974 1952 5976
rect 1955 5974 1957 5983
rect 1971 5981 1973 5993
rect 1987 5991 1989 5993
rect 2008 5991 2010 5993
rect 2013 5990 2015 5993
rect 1971 5974 1973 5977
rect 1987 5974 1989 5976
rect 2008 5974 2010 5976
rect 2013 5974 2015 5983
rect 2029 5974 2031 5993
rect 2045 5986 2047 5993
rect 2050 5983 2052 5993
rect 2066 5986 2068 5993
rect 2082 5991 2084 5993
rect 2087 5990 2089 5993
rect 2045 5974 2047 5976
rect 2050 5974 2052 5979
rect 2066 5974 2068 5982
rect 2082 5974 2084 5976
rect 2087 5974 2089 5983
rect 2103 5981 2105 5993
rect 2119 5991 2121 5993
rect 2140 5991 2142 5993
rect 2145 5990 2147 5993
rect 2103 5974 2105 5977
rect 2119 5974 2121 5976
rect 2140 5974 2142 5976
rect 2145 5974 2147 5983
rect 2161 5974 2163 5993
rect 2177 5986 2179 5993
rect 2182 5983 2184 5993
rect 2198 5986 2200 5993
rect 2214 5991 2216 5993
rect 2219 5990 2221 5993
rect 2177 5974 2179 5976
rect 2182 5974 2184 5979
rect 2198 5974 2200 5982
rect 2214 5974 2216 5976
rect 2219 5974 2221 5983
rect 2235 5981 2237 5993
rect 2251 5991 2253 5993
rect 2272 5991 2274 5993
rect 2277 5990 2279 5993
rect 2235 5974 2237 5977
rect 2251 5974 2253 5976
rect 2272 5974 2274 5976
rect 2277 5974 2279 5983
rect 2293 5974 2295 5993
rect 2309 5986 2311 5993
rect 2314 5983 2316 5993
rect 2309 5974 2311 5976
rect 2314 5974 2316 5979
rect 857 5964 859 5966
rect 873 5963 875 5966
rect 878 5964 880 5966
rect 894 5963 896 5966
rect 910 5963 912 5966
rect 931 5963 933 5966
rect 936 5964 938 5966
rect 952 5964 954 5966
rect 968 5963 970 5966
rect 973 5964 975 5966
rect 989 5964 991 5966
rect 1005 5963 1007 5966
rect 1010 5964 1012 5966
rect 1026 5963 1028 5966
rect 1042 5963 1044 5966
rect 1063 5963 1065 5966
rect 1068 5964 1070 5966
rect 1084 5964 1086 5966
rect 1100 5963 1102 5966
rect 1105 5964 1107 5966
rect 1121 5964 1123 5966
rect 1137 5963 1139 5966
rect 1142 5964 1144 5966
rect 1158 5963 1160 5966
rect 1174 5963 1176 5966
rect 1195 5963 1197 5966
rect 1200 5964 1202 5966
rect 1216 5964 1218 5966
rect 1232 5963 1234 5966
rect 1237 5964 1239 5966
rect 1253 5964 1255 5966
rect 1269 5963 1271 5966
rect 1274 5964 1276 5966
rect 1290 5963 1292 5966
rect 1306 5963 1308 5966
rect 1327 5963 1329 5966
rect 1332 5964 1334 5966
rect 1348 5964 1350 5966
rect 1364 5963 1366 5966
rect 1369 5964 1371 5966
rect 1802 5964 1804 5966
rect 1818 5963 1820 5966
rect 1823 5964 1825 5966
rect 1839 5963 1841 5966
rect 1855 5963 1857 5966
rect 1876 5963 1878 5966
rect 1881 5964 1883 5966
rect 1897 5964 1899 5966
rect 1913 5963 1915 5966
rect 1918 5964 1920 5966
rect 1934 5964 1936 5966
rect 1950 5963 1952 5966
rect 1955 5964 1957 5966
rect 1971 5963 1973 5966
rect 1987 5963 1989 5966
rect 2008 5963 2010 5966
rect 2013 5964 2015 5966
rect 2029 5964 2031 5966
rect 2045 5963 2047 5966
rect 2050 5964 2052 5966
rect 2066 5964 2068 5966
rect 2082 5963 2084 5966
rect 2087 5964 2089 5966
rect 2103 5963 2105 5966
rect 2119 5963 2121 5966
rect 2140 5963 2142 5966
rect 2145 5964 2147 5966
rect 2161 5964 2163 5966
rect 2177 5963 2179 5966
rect 2182 5964 2184 5966
rect 2198 5964 2200 5966
rect 2214 5963 2216 5966
rect 2219 5964 2221 5966
rect 2235 5963 2237 5966
rect 2251 5963 2253 5966
rect 2272 5963 2274 5966
rect 2277 5964 2279 5966
rect 2293 5964 2295 5966
rect 2309 5963 2311 5966
rect 2314 5964 2316 5966
rect 1473 5918 1475 5920
rect 1489 5918 1491 5923
rect 1494 5918 1496 5920
rect 1510 5918 1512 5920
rect 1526 5918 1528 5923
rect 1547 5918 1549 5923
rect 1552 5918 1554 5920
rect 1568 5918 1570 5920
rect 1584 5918 1586 5921
rect 1589 5918 1591 5920
rect 1605 5918 1607 5920
rect 1621 5918 1623 5923
rect 1626 5918 1628 5920
rect 1642 5918 1644 5920
rect 1658 5918 1660 5923
rect 1679 5918 1681 5923
rect 1684 5918 1686 5920
rect 1700 5918 1702 5920
rect 1716 5918 1718 5921
rect 1721 5918 1723 5920
rect 1737 5918 1739 5920
rect 1753 5918 1755 5923
rect 1758 5918 1760 5920
rect 1774 5918 1776 5920
rect 1790 5918 1792 5923
rect 1811 5918 1813 5923
rect 1816 5918 1818 5920
rect 1832 5918 1834 5920
rect 1848 5918 1850 5921
rect 1853 5918 1855 5920
rect 2418 5918 2420 5920
rect 2434 5918 2436 5923
rect 2439 5918 2441 5920
rect 2455 5918 2457 5920
rect 2471 5918 2473 5923
rect 2492 5918 2494 5923
rect 2497 5918 2499 5920
rect 2513 5918 2515 5920
rect 2529 5918 2531 5921
rect 2534 5918 2536 5920
rect 2550 5918 2552 5920
rect 2566 5918 2568 5923
rect 2571 5918 2573 5920
rect 2587 5918 2589 5920
rect 2603 5918 2605 5923
rect 2624 5918 2626 5923
rect 2629 5918 2631 5920
rect 2645 5918 2647 5920
rect 2661 5918 2663 5921
rect 2666 5918 2668 5920
rect 2682 5918 2684 5920
rect 2698 5918 2700 5923
rect 2703 5918 2705 5920
rect 2719 5918 2721 5920
rect 2735 5918 2737 5923
rect 2756 5918 2758 5923
rect 2761 5918 2763 5920
rect 2777 5918 2779 5920
rect 2793 5918 2795 5921
rect 2798 5918 2800 5920
rect 1473 5907 1475 5914
rect 1489 5912 1491 5914
rect 1494 5911 1496 5914
rect 1473 5895 1475 5903
rect 1489 5895 1491 5897
rect 1494 5895 1496 5904
rect 1510 5902 1512 5914
rect 1526 5912 1528 5914
rect 1547 5912 1549 5914
rect 1552 5911 1554 5914
rect 1510 5895 1512 5898
rect 1526 5895 1528 5897
rect 1547 5895 1549 5897
rect 1552 5895 1554 5904
rect 1568 5895 1570 5914
rect 1584 5907 1586 5914
rect 1589 5902 1591 5914
rect 1584 5895 1586 5897
rect 1589 5895 1591 5898
rect 1605 5895 1607 5914
rect 1621 5912 1623 5914
rect 1626 5911 1628 5914
rect 1621 5895 1623 5897
rect 1626 5895 1628 5904
rect 1642 5902 1644 5914
rect 1658 5912 1660 5914
rect 1679 5912 1681 5914
rect 1684 5911 1686 5914
rect 1642 5895 1644 5898
rect 1658 5895 1660 5897
rect 1679 5895 1681 5897
rect 1684 5895 1686 5904
rect 1700 5895 1702 5914
rect 1716 5907 1718 5914
rect 1721 5902 1723 5914
rect 1716 5895 1718 5897
rect 1721 5895 1723 5898
rect 1737 5895 1739 5914
rect 1753 5912 1755 5914
rect 1758 5911 1760 5914
rect 1753 5895 1755 5897
rect 1758 5895 1760 5904
rect 1774 5902 1776 5914
rect 1790 5912 1792 5914
rect 1811 5912 1813 5914
rect 1816 5911 1818 5914
rect 1774 5895 1776 5898
rect 1790 5895 1792 5897
rect 1811 5895 1813 5897
rect 1816 5895 1818 5904
rect 1832 5895 1834 5914
rect 1848 5907 1850 5914
rect 1853 5904 1855 5914
rect 2418 5907 2420 5914
rect 2434 5912 2436 5914
rect 2439 5911 2441 5914
rect 1848 5895 1850 5897
rect 1853 5895 1855 5900
rect 2418 5895 2420 5903
rect 2434 5895 2436 5897
rect 2439 5895 2441 5904
rect 2455 5902 2457 5914
rect 2471 5912 2473 5914
rect 2492 5912 2494 5914
rect 2497 5911 2499 5914
rect 2455 5895 2457 5898
rect 2471 5895 2473 5897
rect 2492 5895 2494 5897
rect 2497 5895 2499 5904
rect 2513 5895 2515 5914
rect 2529 5907 2531 5914
rect 2534 5902 2536 5914
rect 2529 5895 2531 5897
rect 2534 5895 2536 5898
rect 2550 5895 2552 5914
rect 2566 5912 2568 5914
rect 2571 5911 2573 5914
rect 2566 5895 2568 5897
rect 2571 5895 2573 5904
rect 2587 5902 2589 5914
rect 2603 5912 2605 5914
rect 2624 5912 2626 5914
rect 2629 5911 2631 5914
rect 2587 5895 2589 5898
rect 2603 5895 2605 5897
rect 2624 5895 2626 5897
rect 2629 5895 2631 5904
rect 2645 5895 2647 5914
rect 2661 5907 2663 5914
rect 2666 5902 2668 5914
rect 2661 5895 2663 5897
rect 2666 5895 2668 5898
rect 2682 5895 2684 5914
rect 2698 5912 2700 5914
rect 2703 5911 2705 5914
rect 2698 5895 2700 5897
rect 2703 5895 2705 5904
rect 2719 5902 2721 5914
rect 2735 5912 2737 5914
rect 2756 5912 2758 5914
rect 2761 5911 2763 5914
rect 2719 5895 2721 5898
rect 2735 5895 2737 5897
rect 2756 5895 2758 5897
rect 2761 5895 2763 5904
rect 2777 5895 2779 5914
rect 2793 5907 2795 5914
rect 2798 5904 2800 5914
rect 2793 5895 2795 5897
rect 2798 5895 2800 5900
rect 1473 5885 1475 5887
rect 1489 5884 1491 5887
rect 1494 5885 1496 5887
rect 1510 5884 1512 5887
rect 1526 5884 1528 5887
rect 1547 5884 1549 5887
rect 1552 5885 1554 5887
rect 1568 5885 1570 5887
rect 1584 5884 1586 5887
rect 1589 5885 1591 5887
rect 1605 5885 1607 5887
rect 1621 5884 1623 5887
rect 1626 5885 1628 5887
rect 1642 5884 1644 5887
rect 1658 5884 1660 5887
rect 1679 5884 1681 5887
rect 1684 5885 1686 5887
rect 1700 5885 1702 5887
rect 1716 5884 1718 5887
rect 1721 5885 1723 5887
rect 1737 5885 1739 5887
rect 1753 5884 1755 5887
rect 1758 5885 1760 5887
rect 1774 5884 1776 5887
rect 1790 5884 1792 5887
rect 1811 5884 1813 5887
rect 1816 5885 1818 5887
rect 1832 5885 1834 5887
rect 1848 5884 1850 5887
rect 1853 5885 1855 5887
rect 2418 5885 2420 5887
rect 2434 5884 2436 5887
rect 2439 5885 2441 5887
rect 2455 5884 2457 5887
rect 2471 5884 2473 5887
rect 2492 5884 2494 5887
rect 2497 5885 2499 5887
rect 2513 5885 2515 5887
rect 2529 5884 2531 5887
rect 2534 5885 2536 5887
rect 2550 5885 2552 5887
rect 2566 5884 2568 5887
rect 2571 5885 2573 5887
rect 2587 5884 2589 5887
rect 2603 5884 2605 5887
rect 2624 5884 2626 5887
rect 2629 5885 2631 5887
rect 2645 5885 2647 5887
rect 2661 5884 2663 5887
rect 2666 5885 2668 5887
rect 2682 5885 2684 5887
rect 2698 5884 2700 5887
rect 2703 5885 2705 5887
rect 2719 5884 2721 5887
rect 2735 5884 2737 5887
rect 2756 5884 2758 5887
rect 2761 5885 2763 5887
rect 2777 5885 2779 5887
rect 2793 5884 2795 5887
rect 2798 5885 2800 5887
rect 1597 5856 1599 5859
rect 1621 5856 1623 5859
rect 2542 5856 2544 5859
rect 2566 5856 2568 5859
rect 1597 5850 1599 5852
rect 1621 5850 1623 5852
rect 2542 5850 2544 5852
rect 2566 5850 2568 5852
rect 1589 5845 1608 5847
rect 1612 5845 1614 5847
rect 2534 5845 2553 5847
rect 2557 5845 2559 5847
rect 1601 5833 1603 5836
rect 2546 5833 2548 5836
rect 1601 5827 1603 5829
rect 2546 5827 2548 5829
rect 1597 5822 1599 5824
rect 1621 5822 1623 5824
rect 2542 5822 2544 5824
rect 2566 5822 2568 5824
rect 1597 5815 1599 5818
rect 1621 5815 1623 5818
rect 2542 5815 2544 5818
rect 2566 5815 2568 5818
rect 1473 5778 1475 5780
rect 1489 5778 1491 5783
rect 1494 5778 1496 5780
rect 1510 5778 1512 5780
rect 1526 5778 1528 5783
rect 1547 5778 1549 5783
rect 1552 5778 1554 5780
rect 1568 5778 1570 5780
rect 1584 5778 1586 5781
rect 1589 5778 1591 5780
rect 1605 5778 1607 5780
rect 1621 5778 1623 5783
rect 1626 5778 1628 5780
rect 1642 5778 1644 5780
rect 1658 5778 1660 5783
rect 1679 5778 1681 5783
rect 1684 5778 1686 5780
rect 1700 5778 1702 5780
rect 1716 5778 1718 5781
rect 1721 5778 1723 5780
rect 1737 5778 1739 5780
rect 1753 5778 1755 5783
rect 1758 5778 1760 5780
rect 1774 5778 1776 5780
rect 1790 5778 1792 5783
rect 1811 5778 1813 5783
rect 1816 5778 1818 5780
rect 1832 5778 1834 5780
rect 1848 5778 1850 5781
rect 1853 5778 1855 5780
rect 2418 5778 2420 5780
rect 2434 5778 2436 5783
rect 2439 5778 2441 5780
rect 2455 5778 2457 5780
rect 2471 5778 2473 5783
rect 2492 5778 2494 5783
rect 2497 5778 2499 5780
rect 2513 5778 2515 5780
rect 2529 5778 2531 5781
rect 2534 5778 2536 5780
rect 2550 5778 2552 5780
rect 2566 5778 2568 5783
rect 2571 5778 2573 5780
rect 2587 5778 2589 5780
rect 2603 5778 2605 5783
rect 2624 5778 2626 5783
rect 2629 5778 2631 5780
rect 2645 5778 2647 5780
rect 2661 5778 2663 5781
rect 2666 5778 2668 5780
rect 2682 5778 2684 5780
rect 2698 5778 2700 5783
rect 2703 5778 2705 5780
rect 2719 5778 2721 5780
rect 2735 5778 2737 5783
rect 2756 5778 2758 5783
rect 2761 5778 2763 5780
rect 2777 5778 2779 5780
rect 2793 5778 2795 5781
rect 2798 5778 2800 5780
rect 1473 5767 1475 5774
rect 1489 5772 1491 5774
rect 1494 5771 1496 5774
rect 1473 5755 1475 5763
rect 1489 5755 1491 5757
rect 1494 5755 1496 5764
rect 1510 5762 1512 5774
rect 1526 5772 1528 5774
rect 1547 5772 1549 5774
rect 1552 5771 1554 5774
rect 1510 5755 1512 5758
rect 1526 5755 1528 5757
rect 1547 5755 1549 5757
rect 1552 5755 1554 5764
rect 1568 5755 1570 5774
rect 1584 5767 1586 5774
rect 1589 5762 1591 5774
rect 1584 5755 1586 5757
rect 1589 5755 1591 5758
rect 1605 5755 1607 5774
rect 1621 5772 1623 5774
rect 1626 5771 1628 5774
rect 1621 5755 1623 5757
rect 1626 5755 1628 5764
rect 1642 5762 1644 5774
rect 1658 5772 1660 5774
rect 1679 5772 1681 5774
rect 1684 5771 1686 5774
rect 1642 5755 1644 5758
rect 1658 5755 1660 5757
rect 1679 5755 1681 5757
rect 1684 5755 1686 5764
rect 1700 5755 1702 5774
rect 1716 5767 1718 5774
rect 1721 5762 1723 5774
rect 1716 5755 1718 5757
rect 1721 5755 1723 5758
rect 1737 5755 1739 5774
rect 1753 5772 1755 5774
rect 1758 5771 1760 5774
rect 1753 5755 1755 5757
rect 1758 5755 1760 5764
rect 1774 5762 1776 5774
rect 1790 5772 1792 5774
rect 1811 5772 1813 5774
rect 1816 5771 1818 5774
rect 1774 5755 1776 5758
rect 1790 5755 1792 5757
rect 1811 5755 1813 5757
rect 1816 5755 1818 5764
rect 1832 5755 1834 5774
rect 1848 5767 1850 5774
rect 1853 5764 1855 5774
rect 2418 5767 2420 5774
rect 2434 5772 2436 5774
rect 2439 5771 2441 5774
rect 1848 5755 1850 5757
rect 1853 5755 1855 5760
rect 954 5748 956 5750
rect 970 5748 972 5753
rect 975 5748 977 5750
rect 991 5748 993 5750
rect 1007 5748 1009 5753
rect 1028 5748 1030 5753
rect 1033 5748 1035 5750
rect 1049 5748 1051 5750
rect 1065 5748 1067 5751
rect 1070 5748 1072 5750
rect 2418 5755 2420 5763
rect 2434 5755 2436 5757
rect 2439 5755 2441 5764
rect 2455 5762 2457 5774
rect 2471 5772 2473 5774
rect 2492 5772 2494 5774
rect 2497 5771 2499 5774
rect 2455 5755 2457 5758
rect 2471 5755 2473 5757
rect 2492 5755 2494 5757
rect 2497 5755 2499 5764
rect 2513 5755 2515 5774
rect 2529 5767 2531 5774
rect 2534 5762 2536 5774
rect 2529 5755 2531 5757
rect 2534 5755 2536 5758
rect 2550 5755 2552 5774
rect 2566 5772 2568 5774
rect 2571 5771 2573 5774
rect 2566 5755 2568 5757
rect 2571 5755 2573 5764
rect 2587 5762 2589 5774
rect 2603 5772 2605 5774
rect 2624 5772 2626 5774
rect 2629 5771 2631 5774
rect 2587 5755 2589 5758
rect 2603 5755 2605 5757
rect 2624 5755 2626 5757
rect 2629 5755 2631 5764
rect 2645 5755 2647 5774
rect 2661 5767 2663 5774
rect 2666 5762 2668 5774
rect 2661 5755 2663 5757
rect 2666 5755 2668 5758
rect 2682 5755 2684 5774
rect 2698 5772 2700 5774
rect 2703 5771 2705 5774
rect 2698 5755 2700 5757
rect 2703 5755 2705 5764
rect 2719 5762 2721 5774
rect 2735 5772 2737 5774
rect 2756 5772 2758 5774
rect 2761 5771 2763 5774
rect 2719 5755 2721 5758
rect 2735 5755 2737 5757
rect 2756 5755 2758 5757
rect 2761 5755 2763 5764
rect 2777 5755 2779 5774
rect 2793 5767 2795 5774
rect 2798 5764 2800 5774
rect 2793 5755 2795 5757
rect 2798 5755 2800 5760
rect 1899 5748 1901 5750
rect 1915 5748 1917 5753
rect 1920 5748 1922 5750
rect 1936 5748 1938 5750
rect 1952 5748 1954 5753
rect 1973 5748 1975 5753
rect 1978 5748 1980 5750
rect 1994 5748 1996 5750
rect 2010 5748 2012 5751
rect 2015 5748 2017 5750
rect 1473 5745 1475 5747
rect 1489 5744 1491 5747
rect 1494 5745 1496 5747
rect 1510 5744 1512 5747
rect 1526 5744 1528 5747
rect 1547 5744 1549 5747
rect 1552 5745 1554 5747
rect 1568 5745 1570 5747
rect 1584 5744 1586 5747
rect 1589 5745 1591 5747
rect 1605 5745 1607 5747
rect 1621 5744 1623 5747
rect 1626 5745 1628 5747
rect 1642 5744 1644 5747
rect 1658 5744 1660 5747
rect 1679 5744 1681 5747
rect 1684 5745 1686 5747
rect 1700 5745 1702 5747
rect 1716 5744 1718 5747
rect 1721 5745 1723 5747
rect 1737 5745 1739 5747
rect 1753 5744 1755 5747
rect 1758 5745 1760 5747
rect 1774 5744 1776 5747
rect 1790 5744 1792 5747
rect 1811 5744 1813 5747
rect 1816 5745 1818 5747
rect 1832 5745 1834 5747
rect 1848 5744 1850 5747
rect 1853 5745 1855 5747
rect 2418 5745 2420 5747
rect 2434 5744 2436 5747
rect 2439 5745 2441 5747
rect 2455 5744 2457 5747
rect 2471 5744 2473 5747
rect 2492 5744 2494 5747
rect 2497 5745 2499 5747
rect 2513 5745 2515 5747
rect 2529 5744 2531 5747
rect 2534 5745 2536 5747
rect 2550 5745 2552 5747
rect 2566 5744 2568 5747
rect 2571 5745 2573 5747
rect 2587 5744 2589 5747
rect 2603 5744 2605 5747
rect 2624 5744 2626 5747
rect 2629 5745 2631 5747
rect 2645 5745 2647 5747
rect 2661 5744 2663 5747
rect 2666 5745 2668 5747
rect 2682 5745 2684 5747
rect 2698 5744 2700 5747
rect 2703 5745 2705 5747
rect 2719 5744 2721 5747
rect 2735 5744 2737 5747
rect 2756 5744 2758 5747
rect 2761 5745 2763 5747
rect 2777 5745 2779 5747
rect 2793 5744 2795 5747
rect 2798 5745 2800 5747
rect 924 5736 927 5738
rect 931 5736 934 5738
rect 954 5725 956 5744
rect 970 5742 972 5744
rect 975 5741 977 5744
rect 970 5725 972 5727
rect 975 5725 977 5734
rect 991 5732 993 5744
rect 1007 5742 1009 5744
rect 1028 5742 1030 5744
rect 1033 5741 1035 5744
rect 991 5725 993 5728
rect 1007 5725 1009 5727
rect 1028 5725 1030 5727
rect 1033 5725 1035 5734
rect 1049 5725 1051 5744
rect 1065 5737 1067 5744
rect 1070 5734 1072 5744
rect 1869 5736 1872 5738
rect 1876 5736 1879 5738
rect 1065 5725 1067 5727
rect 1070 5725 1072 5730
rect 1899 5725 1901 5744
rect 1915 5742 1917 5744
rect 1920 5741 1922 5744
rect 1915 5725 1917 5727
rect 1920 5725 1922 5734
rect 1936 5732 1938 5744
rect 1952 5742 1954 5744
rect 1973 5742 1975 5744
rect 1978 5741 1980 5744
rect 1936 5725 1938 5728
rect 1952 5725 1954 5727
rect 1973 5725 1975 5727
rect 1978 5725 1980 5734
rect 1994 5725 1996 5744
rect 2010 5737 2012 5744
rect 2015 5734 2017 5744
rect 2010 5725 2012 5727
rect 2015 5725 2017 5730
rect 954 5715 956 5717
rect 970 5714 972 5717
rect 975 5715 977 5717
rect 991 5714 993 5717
rect 1007 5714 1009 5717
rect 1028 5714 1030 5717
rect 1033 5715 1035 5717
rect 1049 5715 1051 5717
rect 1065 5714 1067 5717
rect 1070 5715 1072 5717
rect 1899 5715 1901 5717
rect 1915 5714 1917 5717
rect 1920 5715 1922 5717
rect 1936 5714 1938 5717
rect 1952 5714 1954 5717
rect 1973 5714 1975 5717
rect 1978 5715 1980 5717
rect 1994 5715 1996 5717
rect 2010 5714 2012 5717
rect 2015 5715 2017 5717
rect 1473 5692 1475 5694
rect 1489 5692 1491 5697
rect 1494 5692 1496 5694
rect 1510 5692 1512 5694
rect 1526 5692 1528 5697
rect 1547 5692 1549 5697
rect 1552 5692 1554 5694
rect 1568 5692 1570 5694
rect 1584 5692 1586 5695
rect 1589 5692 1591 5694
rect 1605 5692 1607 5694
rect 1621 5692 1623 5697
rect 1626 5692 1628 5694
rect 1642 5692 1644 5694
rect 1658 5692 1660 5697
rect 1679 5692 1681 5697
rect 1684 5692 1686 5694
rect 1700 5692 1702 5694
rect 1716 5692 1718 5695
rect 1721 5692 1723 5694
rect 1737 5692 1739 5694
rect 1753 5692 1755 5697
rect 1758 5692 1760 5694
rect 1774 5692 1776 5694
rect 1790 5692 1792 5697
rect 1811 5692 1813 5697
rect 1816 5692 1818 5694
rect 1832 5692 1834 5694
rect 1848 5692 1850 5695
rect 1853 5692 1855 5694
rect 2418 5692 2420 5694
rect 2434 5692 2436 5697
rect 2439 5692 2441 5694
rect 2455 5692 2457 5694
rect 2471 5692 2473 5697
rect 2492 5692 2494 5697
rect 2497 5692 2499 5694
rect 2513 5692 2515 5694
rect 2529 5692 2531 5695
rect 2534 5692 2536 5694
rect 2550 5692 2552 5694
rect 2566 5692 2568 5697
rect 2571 5692 2573 5694
rect 2587 5692 2589 5694
rect 2603 5692 2605 5697
rect 2624 5692 2626 5697
rect 2629 5692 2631 5694
rect 2645 5692 2647 5694
rect 2661 5692 2663 5695
rect 2666 5692 2668 5694
rect 2682 5692 2684 5694
rect 2698 5692 2700 5697
rect 2703 5692 2705 5694
rect 2719 5692 2721 5694
rect 2735 5692 2737 5697
rect 2756 5692 2758 5697
rect 2761 5692 2763 5694
rect 2777 5692 2779 5694
rect 2793 5692 2795 5695
rect 2798 5692 2800 5694
rect 1473 5681 1475 5688
rect 1489 5686 1491 5688
rect 1494 5685 1496 5688
rect 1473 5669 1475 5677
rect 1489 5669 1491 5671
rect 1494 5669 1496 5678
rect 1510 5676 1512 5688
rect 1526 5686 1528 5688
rect 1547 5686 1549 5688
rect 1552 5685 1554 5688
rect 1510 5669 1512 5672
rect 1526 5669 1528 5671
rect 1547 5669 1549 5671
rect 1552 5669 1554 5678
rect 1568 5669 1570 5688
rect 1584 5681 1586 5688
rect 1589 5676 1591 5688
rect 1584 5669 1586 5671
rect 1589 5669 1591 5672
rect 1605 5669 1607 5688
rect 1621 5686 1623 5688
rect 1626 5685 1628 5688
rect 1621 5669 1623 5671
rect 1626 5669 1628 5678
rect 1642 5676 1644 5688
rect 1658 5686 1660 5688
rect 1679 5686 1681 5688
rect 1684 5685 1686 5688
rect 1642 5669 1644 5672
rect 1658 5669 1660 5671
rect 1679 5669 1681 5671
rect 1684 5669 1686 5678
rect 1700 5669 1702 5688
rect 1716 5681 1718 5688
rect 1721 5676 1723 5688
rect 1716 5669 1718 5671
rect 1721 5669 1723 5672
rect 1737 5669 1739 5688
rect 1753 5686 1755 5688
rect 1758 5685 1760 5688
rect 1753 5669 1755 5671
rect 1758 5669 1760 5678
rect 1774 5676 1776 5688
rect 1790 5686 1792 5688
rect 1811 5686 1813 5688
rect 1816 5685 1818 5688
rect 1774 5669 1776 5672
rect 1790 5669 1792 5671
rect 1811 5669 1813 5671
rect 1816 5669 1818 5678
rect 1832 5669 1834 5688
rect 1848 5681 1850 5688
rect 1853 5678 1855 5688
rect 2418 5681 2420 5688
rect 2434 5686 2436 5688
rect 2439 5685 2441 5688
rect 1848 5669 1850 5671
rect 1853 5669 1855 5674
rect 954 5662 956 5664
rect 970 5662 972 5667
rect 975 5662 977 5664
rect 991 5662 993 5664
rect 1007 5662 1009 5667
rect 1028 5662 1030 5667
rect 1033 5662 1035 5664
rect 1049 5662 1051 5664
rect 1065 5662 1067 5665
rect 1070 5662 1072 5664
rect 2418 5669 2420 5677
rect 2434 5669 2436 5671
rect 2439 5669 2441 5678
rect 2455 5676 2457 5688
rect 2471 5686 2473 5688
rect 2492 5686 2494 5688
rect 2497 5685 2499 5688
rect 2455 5669 2457 5672
rect 2471 5669 2473 5671
rect 2492 5669 2494 5671
rect 2497 5669 2499 5678
rect 2513 5669 2515 5688
rect 2529 5681 2531 5688
rect 2534 5676 2536 5688
rect 2529 5669 2531 5671
rect 2534 5669 2536 5672
rect 2550 5669 2552 5688
rect 2566 5686 2568 5688
rect 2571 5685 2573 5688
rect 2566 5669 2568 5671
rect 2571 5669 2573 5678
rect 2587 5676 2589 5688
rect 2603 5686 2605 5688
rect 2624 5686 2626 5688
rect 2629 5685 2631 5688
rect 2587 5669 2589 5672
rect 2603 5669 2605 5671
rect 2624 5669 2626 5671
rect 2629 5669 2631 5678
rect 2645 5669 2647 5688
rect 2661 5681 2663 5688
rect 2666 5676 2668 5688
rect 2661 5669 2663 5671
rect 2666 5669 2668 5672
rect 2682 5669 2684 5688
rect 2698 5686 2700 5688
rect 2703 5685 2705 5688
rect 2698 5669 2700 5671
rect 2703 5669 2705 5678
rect 2719 5676 2721 5688
rect 2735 5686 2737 5688
rect 2756 5686 2758 5688
rect 2761 5685 2763 5688
rect 2719 5669 2721 5672
rect 2735 5669 2737 5671
rect 2756 5669 2758 5671
rect 2761 5669 2763 5678
rect 2777 5669 2779 5688
rect 2793 5681 2795 5688
rect 2798 5678 2800 5688
rect 2793 5669 2795 5671
rect 2798 5669 2800 5674
rect 1899 5662 1901 5664
rect 1915 5662 1917 5667
rect 1920 5662 1922 5664
rect 1936 5662 1938 5664
rect 1952 5662 1954 5667
rect 1973 5662 1975 5667
rect 1978 5662 1980 5664
rect 1994 5662 1996 5664
rect 2010 5662 2012 5665
rect 2015 5662 2017 5664
rect 1473 5659 1475 5661
rect 1489 5658 1491 5661
rect 1494 5659 1496 5661
rect 1510 5658 1512 5661
rect 1526 5658 1528 5661
rect 1547 5658 1549 5661
rect 1552 5659 1554 5661
rect 1568 5659 1570 5661
rect 1584 5658 1586 5661
rect 1589 5659 1591 5661
rect 1605 5659 1607 5661
rect 1621 5658 1623 5661
rect 1626 5659 1628 5661
rect 1642 5658 1644 5661
rect 1658 5658 1660 5661
rect 1679 5658 1681 5661
rect 1684 5659 1686 5661
rect 1700 5659 1702 5661
rect 1716 5658 1718 5661
rect 1721 5659 1723 5661
rect 1737 5659 1739 5661
rect 1753 5658 1755 5661
rect 1758 5659 1760 5661
rect 1774 5658 1776 5661
rect 1790 5658 1792 5661
rect 1811 5658 1813 5661
rect 1816 5659 1818 5661
rect 1832 5659 1834 5661
rect 1848 5658 1850 5661
rect 1853 5659 1855 5661
rect 2418 5659 2420 5661
rect 2434 5658 2436 5661
rect 2439 5659 2441 5661
rect 2455 5658 2457 5661
rect 2471 5658 2473 5661
rect 2492 5658 2494 5661
rect 2497 5659 2499 5661
rect 2513 5659 2515 5661
rect 2529 5658 2531 5661
rect 2534 5659 2536 5661
rect 2550 5659 2552 5661
rect 2566 5658 2568 5661
rect 2571 5659 2573 5661
rect 2587 5658 2589 5661
rect 2603 5658 2605 5661
rect 2624 5658 2626 5661
rect 2629 5659 2631 5661
rect 2645 5659 2647 5661
rect 2661 5658 2663 5661
rect 2666 5659 2668 5661
rect 2682 5659 2684 5661
rect 2698 5658 2700 5661
rect 2703 5659 2705 5661
rect 2719 5658 2721 5661
rect 2735 5658 2737 5661
rect 2756 5658 2758 5661
rect 2761 5659 2763 5661
rect 2777 5659 2779 5661
rect 2793 5658 2795 5661
rect 2798 5659 2800 5661
rect 954 5639 956 5658
rect 970 5656 972 5658
rect 975 5655 977 5658
rect 970 5639 972 5641
rect 975 5639 977 5648
rect 991 5646 993 5658
rect 1007 5656 1009 5658
rect 1028 5656 1030 5658
rect 1033 5655 1035 5658
rect 991 5639 993 5642
rect 1007 5639 1009 5641
rect 1028 5639 1030 5641
rect 1033 5639 1035 5648
rect 1049 5639 1051 5658
rect 1065 5651 1067 5658
rect 1070 5648 1072 5658
rect 1065 5639 1067 5641
rect 1070 5639 1072 5644
rect 1899 5639 1901 5658
rect 1915 5656 1917 5658
rect 1920 5655 1922 5658
rect 1915 5639 1917 5641
rect 1920 5639 1922 5648
rect 1936 5646 1938 5658
rect 1952 5656 1954 5658
rect 1973 5656 1975 5658
rect 1978 5655 1980 5658
rect 1936 5639 1938 5642
rect 1952 5639 1954 5641
rect 1973 5639 1975 5641
rect 1978 5639 1980 5648
rect 1994 5639 1996 5658
rect 2010 5651 2012 5658
rect 2015 5648 2017 5658
rect 2010 5639 2012 5641
rect 2015 5639 2017 5644
rect 954 5629 956 5631
rect 970 5628 972 5631
rect 975 5629 977 5631
rect 991 5628 993 5631
rect 1007 5628 1009 5631
rect 1028 5628 1030 5631
rect 1033 5629 1035 5631
rect 1049 5629 1051 5631
rect 1065 5628 1067 5631
rect 1070 5629 1072 5631
rect 1714 5630 1716 5633
rect 1738 5630 1740 5633
rect 1899 5629 1901 5631
rect 1915 5628 1917 5631
rect 1920 5629 1922 5631
rect 1936 5628 1938 5631
rect 1952 5628 1954 5631
rect 1973 5628 1975 5631
rect 1978 5629 1980 5631
rect 1994 5629 1996 5631
rect 2010 5628 2012 5631
rect 2015 5629 2017 5631
rect 2659 5630 2661 5633
rect 2683 5630 2685 5633
rect 1714 5624 1716 5626
rect 1738 5624 1740 5626
rect 2659 5624 2661 5626
rect 2683 5624 2685 5626
rect 1706 5619 1725 5621
rect 1729 5619 1731 5621
rect 2651 5619 2670 5621
rect 2674 5619 2676 5621
rect 1718 5607 1720 5610
rect 2663 5607 2665 5610
rect 1718 5601 1720 5603
rect 2663 5601 2665 5603
rect 936 5590 939 5592
rect 943 5590 946 5592
rect 971 5565 973 5568
rect 1017 5565 1019 5568
rect 1043 5565 1045 5568
rect 1087 5565 1089 5568
rect 1018 5561 1019 5565
rect 953 5558 955 5560
rect 971 5558 973 5561
rect 976 5558 978 5560
rect 996 5558 998 5561
rect 1017 5558 1019 5561
rect 1043 5558 1045 5561
rect 1048 5558 1050 5560
rect 1071 5558 1073 5560
rect 1087 5558 1089 5561
rect 1112 5558 1114 5596
rect 1714 5594 1716 5597
rect 1738 5594 1740 5597
rect 1881 5590 1884 5592
rect 1888 5590 1891 5592
rect 1714 5587 1716 5590
rect 1738 5587 1740 5590
rect 1159 5563 1161 5568
rect 1232 5565 1234 5568
rect 1278 5565 1280 5568
rect 1304 5565 1306 5568
rect 1348 5565 1350 5568
rect 1164 5563 1166 5565
rect 1130 5558 1132 5561
rect 1279 5561 1280 5565
rect 1916 5565 1918 5568
rect 1962 5565 1964 5568
rect 1988 5565 1990 5568
rect 2032 5565 2034 5568
rect 1963 5561 1964 5565
rect 1214 5558 1216 5560
rect 1232 5558 1234 5561
rect 1237 5558 1239 5560
rect 1257 5558 1259 5561
rect 1278 5558 1280 5561
rect 1304 5558 1306 5561
rect 1309 5558 1311 5560
rect 1332 5558 1334 5560
rect 1348 5558 1350 5561
rect 1364 5558 1366 5560
rect 1159 5553 1161 5555
rect 953 5536 955 5550
rect 971 5548 973 5550
rect 976 5545 978 5550
rect 976 5541 982 5545
rect 971 5536 973 5538
rect 976 5536 978 5541
rect 996 5536 998 5550
rect 1017 5548 1019 5550
rect 1043 5548 1045 5550
rect 1048 5545 1050 5550
rect 1048 5541 1054 5545
rect 1017 5536 1019 5538
rect 1043 5536 1045 5538
rect 1048 5536 1050 5541
rect 1071 5536 1073 5550
rect 1087 5548 1089 5550
rect 1087 5536 1089 5538
rect 1112 5536 1114 5550
rect 1130 5545 1132 5550
rect 1159 5543 1161 5545
rect 1164 5543 1166 5555
rect 1473 5550 1475 5552
rect 1489 5550 1491 5555
rect 1494 5550 1496 5552
rect 1510 5550 1512 5552
rect 1526 5550 1528 5555
rect 1547 5550 1549 5555
rect 1552 5550 1554 5552
rect 1568 5550 1570 5552
rect 1584 5550 1586 5553
rect 1589 5550 1591 5552
rect 1605 5550 1607 5552
rect 1621 5550 1623 5555
rect 1626 5550 1628 5552
rect 1642 5550 1644 5552
rect 1658 5550 1660 5555
rect 1679 5550 1681 5555
rect 1684 5550 1686 5552
rect 1700 5550 1702 5552
rect 1716 5550 1718 5553
rect 1898 5558 1900 5560
rect 1916 5558 1918 5561
rect 1921 5558 1923 5560
rect 1941 5558 1943 5561
rect 1962 5558 1964 5561
rect 1988 5558 1990 5561
rect 1993 5558 1995 5560
rect 2016 5558 2018 5560
rect 2032 5558 2034 5561
rect 2057 5558 2059 5600
rect 2659 5594 2661 5597
rect 2683 5594 2685 5597
rect 2659 5587 2661 5590
rect 2683 5587 2685 5590
rect 2104 5563 2106 5568
rect 2177 5565 2179 5568
rect 2223 5565 2225 5568
rect 2249 5565 2251 5568
rect 2293 5565 2295 5568
rect 2109 5563 2111 5565
rect 2075 5558 2077 5561
rect 1721 5550 1723 5552
rect 1737 5550 1739 5552
rect 1753 5550 1755 5555
rect 1758 5550 1760 5552
rect 1774 5550 1776 5552
rect 1790 5550 1792 5555
rect 1811 5550 1813 5555
rect 1816 5550 1818 5552
rect 1832 5550 1834 5552
rect 1848 5550 1850 5553
rect 1853 5550 1855 5552
rect 2224 5561 2225 5565
rect 2159 5558 2161 5560
rect 2177 5558 2179 5561
rect 2182 5558 2184 5560
rect 2202 5558 2204 5561
rect 2223 5558 2225 5561
rect 2249 5558 2251 5561
rect 2254 5558 2256 5560
rect 2277 5558 2279 5560
rect 2293 5558 2295 5561
rect 2309 5558 2311 5560
rect 2104 5553 2106 5555
rect 1130 5536 1132 5541
rect 1159 5536 1161 5539
rect 1164 5536 1166 5539
rect 1214 5536 1216 5550
rect 1232 5548 1234 5550
rect 1237 5545 1239 5550
rect 1237 5541 1243 5545
rect 1232 5536 1234 5538
rect 1237 5536 1239 5541
rect 1257 5536 1259 5550
rect 1278 5548 1280 5550
rect 1304 5548 1306 5550
rect 1309 5545 1311 5550
rect 1309 5541 1315 5545
rect 1278 5536 1280 5538
rect 1304 5536 1306 5538
rect 1309 5536 1311 5541
rect 1332 5536 1334 5550
rect 1348 5548 1350 5550
rect 1348 5536 1350 5538
rect 1364 5536 1366 5550
rect 1473 5539 1475 5546
rect 1489 5544 1491 5546
rect 1494 5543 1496 5546
rect 953 5530 955 5532
rect 971 5527 973 5532
rect 976 5530 978 5532
rect 996 5530 998 5532
rect 1017 5528 1019 5532
rect 971 5523 972 5527
rect 1017 5524 1018 5528
rect 1043 5527 1045 5532
rect 1048 5530 1050 5532
rect 1071 5530 1073 5532
rect 1087 5528 1089 5532
rect 1112 5529 1114 5532
rect 1130 5529 1132 5532
rect 1214 5530 1216 5532
rect 971 5521 973 5523
rect 1017 5520 1019 5524
rect 1043 5523 1044 5527
rect 1087 5524 1088 5528
rect 1232 5527 1234 5532
rect 1237 5530 1239 5532
rect 1257 5530 1259 5532
rect 1278 5528 1280 5532
rect 1043 5521 1045 5523
rect 1087 5521 1089 5524
rect 1232 5523 1233 5527
rect 1278 5524 1279 5528
rect 1304 5527 1306 5532
rect 1309 5530 1311 5532
rect 1332 5530 1334 5532
rect 1348 5528 1350 5532
rect 1364 5530 1366 5532
rect 1232 5521 1234 5523
rect 1278 5520 1280 5524
rect 1304 5523 1305 5527
rect 1348 5524 1349 5528
rect 1473 5527 1475 5535
rect 1489 5527 1491 5529
rect 1494 5527 1496 5536
rect 1510 5534 1512 5546
rect 1526 5544 1528 5546
rect 1547 5544 1549 5546
rect 1552 5543 1554 5546
rect 1510 5527 1512 5530
rect 1526 5527 1528 5529
rect 1547 5527 1549 5529
rect 1552 5527 1554 5536
rect 1568 5527 1570 5546
rect 1584 5539 1586 5546
rect 1589 5534 1591 5546
rect 1584 5527 1586 5529
rect 1589 5527 1591 5530
rect 1605 5527 1607 5546
rect 1621 5544 1623 5546
rect 1626 5543 1628 5546
rect 1621 5527 1623 5529
rect 1626 5527 1628 5536
rect 1642 5534 1644 5546
rect 1658 5544 1660 5546
rect 1679 5544 1681 5546
rect 1684 5543 1686 5546
rect 1642 5527 1644 5530
rect 1658 5527 1660 5529
rect 1679 5527 1681 5529
rect 1684 5527 1686 5536
rect 1700 5527 1702 5546
rect 1716 5539 1718 5546
rect 1721 5534 1723 5546
rect 1716 5527 1718 5529
rect 1721 5527 1723 5530
rect 1737 5527 1739 5546
rect 1753 5544 1755 5546
rect 1758 5543 1760 5546
rect 1753 5527 1755 5529
rect 1758 5527 1760 5536
rect 1774 5534 1776 5546
rect 1790 5544 1792 5546
rect 1811 5544 1813 5546
rect 1816 5543 1818 5546
rect 1774 5527 1776 5530
rect 1790 5527 1792 5529
rect 1811 5527 1813 5529
rect 1816 5527 1818 5536
rect 1832 5527 1834 5546
rect 1848 5539 1850 5546
rect 1853 5536 1855 5546
rect 1898 5536 1900 5550
rect 1916 5548 1918 5550
rect 1921 5545 1923 5550
rect 1921 5541 1927 5545
rect 1916 5536 1918 5538
rect 1921 5536 1923 5541
rect 1941 5536 1943 5550
rect 1962 5548 1964 5550
rect 1988 5548 1990 5550
rect 1993 5545 1995 5550
rect 1993 5541 1999 5545
rect 1962 5536 1964 5538
rect 1988 5536 1990 5538
rect 1993 5536 1995 5541
rect 2016 5536 2018 5550
rect 2032 5548 2034 5550
rect 2032 5536 2034 5538
rect 2057 5536 2059 5550
rect 2075 5545 2077 5550
rect 2104 5543 2106 5545
rect 2109 5543 2111 5555
rect 2418 5550 2420 5552
rect 2434 5550 2436 5555
rect 2439 5550 2441 5552
rect 2455 5550 2457 5552
rect 2471 5550 2473 5555
rect 2492 5550 2494 5555
rect 2497 5550 2499 5552
rect 2513 5550 2515 5552
rect 2529 5550 2531 5553
rect 2534 5550 2536 5552
rect 2550 5550 2552 5552
rect 2566 5550 2568 5555
rect 2571 5550 2573 5552
rect 2587 5550 2589 5552
rect 2603 5550 2605 5555
rect 2624 5550 2626 5555
rect 2629 5550 2631 5552
rect 2645 5550 2647 5552
rect 2661 5550 2663 5553
rect 2666 5550 2668 5552
rect 2682 5550 2684 5552
rect 2698 5550 2700 5555
rect 2703 5550 2705 5552
rect 2719 5550 2721 5552
rect 2735 5550 2737 5555
rect 2756 5550 2758 5555
rect 2761 5550 2763 5552
rect 2777 5550 2779 5552
rect 2793 5550 2795 5553
rect 2798 5550 2800 5552
rect 2075 5536 2077 5541
rect 2104 5536 2106 5539
rect 2109 5536 2111 5539
rect 2159 5536 2161 5550
rect 2177 5548 2179 5550
rect 2182 5545 2184 5550
rect 2182 5541 2188 5545
rect 2177 5536 2179 5538
rect 2182 5536 2184 5541
rect 2202 5536 2204 5550
rect 2223 5548 2225 5550
rect 2249 5548 2251 5550
rect 2254 5545 2256 5550
rect 2254 5541 2260 5545
rect 2223 5536 2225 5538
rect 2249 5536 2251 5538
rect 2254 5536 2256 5541
rect 2277 5536 2279 5550
rect 2293 5548 2295 5550
rect 2293 5536 2295 5538
rect 2309 5536 2311 5550
rect 2418 5539 2420 5546
rect 2434 5544 2436 5546
rect 2439 5543 2441 5546
rect 1848 5527 1850 5529
rect 1853 5527 1855 5532
rect 1898 5530 1900 5532
rect 1916 5527 1918 5532
rect 1921 5530 1923 5532
rect 1941 5530 1943 5532
rect 1962 5528 1964 5532
rect 1304 5521 1306 5523
rect 1348 5521 1350 5524
rect 1916 5523 1917 5527
rect 1962 5524 1963 5528
rect 1988 5527 1990 5532
rect 1993 5530 1995 5532
rect 2016 5530 2018 5532
rect 2032 5528 2034 5532
rect 2057 5529 2059 5532
rect 2075 5529 2077 5532
rect 2159 5530 2161 5532
rect 1916 5521 1918 5523
rect 1962 5520 1964 5524
rect 1988 5523 1989 5527
rect 2032 5524 2033 5528
rect 2177 5527 2179 5532
rect 2182 5530 2184 5532
rect 2202 5530 2204 5532
rect 2223 5528 2225 5532
rect 1988 5521 1990 5523
rect 2032 5521 2034 5524
rect 2177 5523 2178 5527
rect 2223 5524 2224 5528
rect 2249 5527 2251 5532
rect 2254 5530 2256 5532
rect 2277 5530 2279 5532
rect 2293 5528 2295 5532
rect 2309 5530 2311 5532
rect 2177 5521 2179 5523
rect 2223 5520 2225 5524
rect 2249 5523 2250 5527
rect 2293 5524 2294 5528
rect 2418 5527 2420 5535
rect 2434 5527 2436 5529
rect 2439 5527 2441 5536
rect 2455 5534 2457 5546
rect 2471 5544 2473 5546
rect 2492 5544 2494 5546
rect 2497 5543 2499 5546
rect 2455 5527 2457 5530
rect 2471 5527 2473 5529
rect 2492 5527 2494 5529
rect 2497 5527 2499 5536
rect 2513 5527 2515 5546
rect 2529 5539 2531 5546
rect 2534 5534 2536 5546
rect 2529 5527 2531 5529
rect 2534 5527 2536 5530
rect 2550 5527 2552 5546
rect 2566 5544 2568 5546
rect 2571 5543 2573 5546
rect 2566 5527 2568 5529
rect 2571 5527 2573 5536
rect 2587 5534 2589 5546
rect 2603 5544 2605 5546
rect 2624 5544 2626 5546
rect 2629 5543 2631 5546
rect 2587 5527 2589 5530
rect 2603 5527 2605 5529
rect 2624 5527 2626 5529
rect 2629 5527 2631 5536
rect 2645 5527 2647 5546
rect 2661 5539 2663 5546
rect 2666 5534 2668 5546
rect 2661 5527 2663 5529
rect 2666 5527 2668 5530
rect 2682 5527 2684 5546
rect 2698 5544 2700 5546
rect 2703 5543 2705 5546
rect 2698 5527 2700 5529
rect 2703 5527 2705 5536
rect 2719 5534 2721 5546
rect 2735 5544 2737 5546
rect 2756 5544 2758 5546
rect 2761 5543 2763 5546
rect 2719 5527 2721 5530
rect 2735 5527 2737 5529
rect 2756 5527 2758 5529
rect 2761 5527 2763 5536
rect 2777 5527 2779 5546
rect 2793 5539 2795 5546
rect 2798 5536 2800 5546
rect 2793 5527 2795 5529
rect 2798 5527 2800 5532
rect 2249 5521 2251 5523
rect 2293 5521 2295 5524
rect 1473 5517 1475 5519
rect 1489 5516 1491 5519
rect 1494 5517 1496 5519
rect 1510 5516 1512 5519
rect 1526 5516 1528 5519
rect 1547 5516 1549 5519
rect 1552 5517 1554 5519
rect 1568 5517 1570 5519
rect 1584 5516 1586 5519
rect 1589 5517 1591 5519
rect 1605 5517 1607 5519
rect 1621 5516 1623 5519
rect 1626 5517 1628 5519
rect 1642 5516 1644 5519
rect 1658 5516 1660 5519
rect 1679 5516 1681 5519
rect 1684 5517 1686 5519
rect 1700 5517 1702 5519
rect 1716 5516 1718 5519
rect 1721 5517 1723 5519
rect 1737 5517 1739 5519
rect 1753 5516 1755 5519
rect 1758 5517 1760 5519
rect 1774 5516 1776 5519
rect 1790 5516 1792 5519
rect 1811 5516 1813 5519
rect 1816 5517 1818 5519
rect 1832 5517 1834 5519
rect 1848 5516 1850 5519
rect 1853 5517 1855 5519
rect 2418 5517 2420 5519
rect 2434 5516 2436 5519
rect 2439 5517 2441 5519
rect 2455 5516 2457 5519
rect 2471 5516 2473 5519
rect 2492 5516 2494 5519
rect 2497 5517 2499 5519
rect 2513 5517 2515 5519
rect 2529 5516 2531 5519
rect 2534 5517 2536 5519
rect 2550 5517 2552 5519
rect 2566 5516 2568 5519
rect 2571 5517 2573 5519
rect 2587 5516 2589 5519
rect 2603 5516 2605 5519
rect 2624 5516 2626 5519
rect 2629 5517 2631 5519
rect 2645 5517 2647 5519
rect 2661 5516 2663 5519
rect 2666 5517 2668 5519
rect 2682 5517 2684 5519
rect 2698 5516 2700 5519
rect 2703 5517 2705 5519
rect 2719 5516 2721 5519
rect 2735 5516 2737 5519
rect 2756 5516 2758 5519
rect 2761 5517 2763 5519
rect 2777 5517 2779 5519
rect 2793 5516 2795 5519
rect 2798 5517 2800 5519
rect 1232 5499 1234 5501
rect 1232 5495 1233 5499
rect 1278 5498 1280 5502
rect 1304 5499 1306 5501
rect 1214 5490 1216 5492
rect 1232 5490 1234 5495
rect 1278 5494 1279 5498
rect 1304 5495 1305 5499
rect 1348 5498 1350 5501
rect 2177 5499 2179 5501
rect 1237 5490 1239 5492
rect 1257 5490 1259 5492
rect 1278 5490 1280 5494
rect 1304 5490 1306 5495
rect 1348 5494 1349 5498
rect 2177 5495 2178 5499
rect 2223 5498 2225 5502
rect 2249 5499 2251 5501
rect 1309 5490 1311 5492
rect 1332 5490 1334 5492
rect 1348 5490 1350 5494
rect 1364 5490 1366 5492
rect 2159 5490 2161 5492
rect 2177 5490 2179 5495
rect 2223 5494 2224 5498
rect 2249 5495 2250 5499
rect 2293 5498 2295 5501
rect 2182 5490 2184 5492
rect 2202 5490 2204 5492
rect 2223 5490 2225 5494
rect 2249 5490 2251 5495
rect 2293 5494 2294 5498
rect 2254 5490 2256 5492
rect 2277 5490 2279 5492
rect 2293 5490 2295 5494
rect 2309 5490 2311 5492
rect 1136 5485 1138 5487
rect 1159 5481 1161 5486
rect 1164 5481 1166 5483
rect 1136 5459 1138 5481
rect 1159 5475 1161 5477
rect 1164 5472 1166 5477
rect 1214 5472 1216 5486
rect 1232 5484 1234 5486
rect 1237 5481 1239 5486
rect 1237 5477 1243 5481
rect 1232 5472 1234 5474
rect 1237 5472 1239 5477
rect 1257 5472 1259 5486
rect 1278 5484 1280 5486
rect 1304 5484 1306 5486
rect 1309 5481 1311 5486
rect 1309 5477 1315 5481
rect 1278 5472 1280 5474
rect 1304 5472 1306 5474
rect 1309 5472 1311 5477
rect 1332 5472 1334 5486
rect 1348 5484 1350 5486
rect 1348 5472 1350 5474
rect 1364 5472 1366 5486
rect 2081 5485 2083 5487
rect 2104 5481 2106 5486
rect 2109 5481 2111 5483
rect 1164 5468 1165 5472
rect 1159 5465 1161 5467
rect 1164 5465 1166 5468
rect 1214 5462 1216 5464
rect 1232 5461 1234 5464
rect 1237 5462 1239 5464
rect 1257 5461 1259 5464
rect 1278 5461 1280 5464
rect 1304 5461 1306 5464
rect 1309 5462 1311 5464
rect 1332 5462 1334 5464
rect 1348 5461 1350 5464
rect 1364 5462 1366 5464
rect 1279 5457 1280 5461
rect 1159 5454 1161 5457
rect 1136 5449 1138 5451
rect 1164 5453 1166 5457
rect 1232 5454 1234 5457
rect 1278 5454 1280 5457
rect 1304 5454 1306 5457
rect 1348 5454 1350 5457
rect 1768 5456 1770 5461
rect 2081 5459 2083 5481
rect 2104 5475 2106 5477
rect 2109 5472 2111 5477
rect 2159 5472 2161 5486
rect 2177 5484 2179 5486
rect 2182 5481 2184 5486
rect 2182 5477 2188 5481
rect 2177 5472 2179 5474
rect 2182 5472 2184 5477
rect 2202 5472 2204 5486
rect 2223 5484 2225 5486
rect 2249 5484 2251 5486
rect 2254 5481 2256 5486
rect 2254 5477 2260 5481
rect 2223 5472 2225 5474
rect 2249 5472 2251 5474
rect 2254 5472 2256 5477
rect 2277 5472 2279 5486
rect 2293 5484 2295 5486
rect 2293 5472 2295 5474
rect 2309 5472 2311 5486
rect 2109 5468 2110 5472
rect 2104 5465 2106 5467
rect 2109 5465 2111 5468
rect 1773 5456 1775 5458
rect 2159 5462 2161 5464
rect 2177 5461 2179 5464
rect 2182 5462 2184 5464
rect 2202 5461 2204 5464
rect 2223 5461 2225 5464
rect 2249 5461 2251 5464
rect 2254 5462 2256 5464
rect 2277 5462 2279 5464
rect 2293 5461 2295 5464
rect 2309 5462 2311 5464
rect 2224 5457 2225 5461
rect 2104 5454 2106 5457
rect 2081 5449 2083 5451
rect 2109 5453 2111 5457
rect 2177 5454 2179 5457
rect 2223 5454 2225 5457
rect 2249 5454 2251 5457
rect 2293 5454 2295 5457
rect 1768 5446 1770 5448
rect 1768 5436 1770 5438
rect 1773 5436 1775 5448
rect 1232 5433 1234 5436
rect 1278 5433 1280 5436
rect 1304 5433 1306 5436
rect 1348 5433 1350 5436
rect 988 5427 990 5432
rect 993 5427 995 5429
rect 1078 5427 1080 5432
rect 1083 5427 1085 5429
rect 1159 5427 1161 5432
rect 1279 5429 1280 5433
rect 2177 5433 2179 5436
rect 2223 5433 2225 5436
rect 2249 5433 2251 5436
rect 2293 5433 2295 5436
rect 1768 5429 1770 5432
rect 1773 5429 1775 5432
rect 1164 5427 1166 5429
rect 1214 5426 1216 5428
rect 1232 5426 1234 5429
rect 1237 5426 1239 5428
rect 1257 5426 1259 5429
rect 1278 5426 1280 5429
rect 1304 5426 1306 5429
rect 1309 5426 1311 5428
rect 1332 5426 1334 5428
rect 1348 5426 1350 5429
rect 1364 5426 1366 5428
rect 988 5417 990 5419
rect 988 5407 990 5409
rect 993 5407 995 5419
rect 1078 5417 1080 5419
rect 1078 5407 1080 5409
rect 1083 5407 1085 5419
rect 1159 5417 1161 5419
rect 1159 5407 1161 5409
rect 1164 5407 1166 5419
rect 1933 5427 1935 5432
rect 1938 5427 1940 5429
rect 2023 5427 2025 5432
rect 2028 5427 2030 5429
rect 2104 5427 2106 5432
rect 2224 5429 2225 5433
rect 2109 5427 2111 5429
rect 2159 5426 2161 5428
rect 2177 5426 2179 5429
rect 2182 5426 2184 5428
rect 2202 5426 2204 5429
rect 2223 5426 2225 5429
rect 2249 5426 2251 5429
rect 2254 5426 2256 5428
rect 2277 5426 2279 5428
rect 2293 5426 2295 5429
rect 2309 5426 2311 5428
rect 1214 5404 1216 5418
rect 1232 5416 1234 5418
rect 1237 5413 1239 5418
rect 1237 5409 1243 5413
rect 1232 5404 1234 5406
rect 1237 5404 1239 5409
rect 1257 5404 1259 5418
rect 1278 5416 1280 5418
rect 1304 5416 1306 5418
rect 1309 5413 1311 5418
rect 1309 5409 1315 5413
rect 1278 5404 1280 5406
rect 1304 5404 1306 5406
rect 1309 5404 1311 5409
rect 1332 5404 1334 5418
rect 1348 5416 1350 5418
rect 1348 5404 1350 5406
rect 1364 5404 1366 5418
rect 1933 5417 1935 5419
rect 1654 5411 1656 5413
rect 1707 5411 1709 5413
rect 988 5400 990 5403
rect 993 5400 995 5403
rect 1078 5400 1080 5403
rect 1083 5400 1085 5403
rect 1159 5400 1161 5403
rect 1164 5400 1166 5403
rect 1214 5398 1216 5400
rect 1232 5395 1234 5400
rect 1237 5398 1239 5400
rect 1257 5398 1259 5400
rect 1278 5396 1280 5400
rect 1232 5391 1233 5395
rect 1278 5392 1279 5396
rect 1304 5395 1306 5400
rect 1309 5398 1311 5400
rect 1332 5398 1334 5400
rect 1348 5396 1350 5400
rect 1364 5398 1366 5400
rect 1933 5407 1935 5409
rect 1938 5407 1940 5419
rect 2023 5417 2025 5419
rect 2023 5407 2025 5409
rect 2028 5407 2030 5419
rect 2104 5417 2106 5419
rect 2104 5407 2106 5409
rect 2109 5407 2111 5419
rect 2159 5404 2161 5418
rect 2177 5416 2179 5418
rect 2182 5413 2184 5418
rect 2182 5409 2188 5413
rect 2177 5404 2179 5406
rect 2182 5404 2184 5409
rect 2202 5404 2204 5418
rect 2223 5416 2225 5418
rect 2249 5416 2251 5418
rect 2254 5413 2256 5418
rect 2254 5409 2260 5413
rect 2223 5404 2225 5406
rect 2249 5404 2251 5406
rect 2254 5404 2256 5409
rect 2277 5404 2279 5418
rect 2293 5416 2295 5418
rect 2293 5404 2295 5406
rect 2309 5404 2311 5418
rect 1933 5400 1935 5403
rect 1938 5400 1940 5403
rect 2023 5400 2025 5403
rect 2028 5400 2030 5403
rect 2104 5400 2106 5403
rect 2109 5400 2111 5403
rect 1232 5389 1234 5391
rect 1278 5388 1280 5392
rect 1304 5391 1305 5395
rect 1348 5392 1349 5396
rect 1304 5389 1306 5391
rect 1348 5389 1350 5392
rect 1654 5391 1656 5399
rect 1707 5391 1709 5399
rect 2159 5398 2161 5400
rect 2177 5395 2179 5400
rect 2182 5398 2184 5400
rect 2202 5398 2204 5400
rect 2223 5396 2225 5400
rect 2177 5391 2178 5395
rect 2223 5392 2224 5396
rect 2249 5395 2251 5400
rect 2254 5398 2256 5400
rect 2277 5398 2279 5400
rect 2293 5396 2295 5400
rect 2309 5398 2311 5400
rect 2177 5389 2179 5391
rect 2223 5388 2225 5392
rect 2249 5391 2250 5395
rect 2293 5392 2294 5396
rect 2249 5389 2251 5391
rect 2293 5389 2295 5392
rect 1654 5379 1656 5387
rect 1707 5379 1709 5387
rect 1745 5380 1747 5382
rect 1232 5367 1234 5369
rect 1232 5363 1233 5367
rect 1278 5366 1280 5370
rect 1304 5367 1306 5369
rect 1214 5358 1216 5360
rect 1232 5358 1234 5363
rect 1278 5362 1279 5366
rect 1304 5363 1305 5367
rect 1348 5366 1350 5369
rect 1237 5358 1239 5360
rect 1257 5358 1259 5360
rect 1278 5358 1280 5362
rect 1304 5358 1306 5363
rect 1348 5362 1349 5366
rect 1309 5358 1311 5360
rect 1332 5358 1334 5360
rect 1348 5358 1350 5362
rect 1364 5358 1366 5360
rect 965 5353 967 5355
rect 988 5349 990 5354
rect 1055 5353 1057 5355
rect 993 5349 995 5351
rect 1078 5349 1080 5354
rect 1136 5353 1138 5355
rect 1083 5349 1085 5351
rect 1159 5349 1161 5354
rect 1164 5349 1166 5351
rect 965 5327 967 5349
rect 1019 5345 1021 5347
rect 988 5343 990 5345
rect 993 5340 995 5345
rect 993 5336 994 5340
rect 988 5333 990 5335
rect 993 5333 995 5336
rect 1019 5327 1021 5341
rect 1055 5327 1057 5349
rect 1109 5345 1111 5347
rect 1078 5343 1080 5345
rect 1083 5340 1085 5345
rect 1083 5336 1084 5340
rect 1078 5333 1080 5335
rect 1083 5333 1085 5336
rect 988 5322 990 5325
rect 965 5317 967 5319
rect 993 5321 995 5325
rect 1109 5327 1111 5341
rect 1136 5327 1138 5349
rect 1159 5343 1161 5345
rect 1164 5340 1166 5345
rect 1214 5340 1216 5354
rect 1232 5352 1234 5354
rect 1237 5349 1239 5354
rect 1237 5345 1243 5349
rect 1232 5340 1234 5342
rect 1237 5340 1239 5345
rect 1257 5340 1259 5354
rect 1278 5352 1280 5354
rect 1304 5352 1306 5354
rect 1309 5349 1311 5354
rect 1309 5345 1315 5349
rect 1278 5340 1280 5342
rect 1304 5340 1306 5342
rect 1309 5340 1311 5345
rect 1332 5340 1334 5354
rect 1348 5352 1350 5354
rect 1348 5340 1350 5342
rect 1364 5340 1366 5354
rect 1768 5376 1770 5381
rect 1773 5376 1775 5378
rect 1745 5354 1747 5376
rect 1799 5372 1801 5374
rect 1821 5372 1823 5374
rect 1768 5370 1770 5372
rect 1773 5367 1775 5372
rect 1773 5363 1774 5367
rect 1768 5360 1770 5362
rect 1773 5360 1775 5363
rect 1654 5346 1656 5349
rect 1707 5346 1709 5349
rect 1799 5354 1801 5368
rect 1821 5354 1823 5368
rect 2177 5367 2179 5369
rect 2177 5363 2178 5367
rect 2223 5366 2225 5370
rect 2249 5367 2251 5369
rect 2159 5358 2161 5360
rect 2177 5358 2179 5363
rect 2223 5362 2224 5366
rect 2249 5363 2250 5367
rect 2293 5366 2295 5369
rect 2182 5358 2184 5360
rect 2202 5358 2204 5360
rect 2223 5358 2225 5362
rect 2249 5358 2251 5363
rect 2293 5362 2294 5366
rect 2254 5358 2256 5360
rect 2277 5358 2279 5360
rect 2293 5358 2295 5362
rect 2309 5358 2311 5360
rect 1768 5349 1770 5352
rect 1745 5344 1747 5346
rect 1773 5348 1775 5352
rect 1910 5353 1912 5355
rect 1933 5349 1935 5354
rect 2000 5353 2002 5355
rect 1938 5349 1940 5351
rect 2023 5349 2025 5354
rect 2081 5353 2083 5355
rect 2028 5349 2030 5351
rect 2104 5349 2106 5354
rect 2109 5349 2111 5351
rect 1799 5344 1801 5346
rect 1821 5344 1823 5346
rect 1164 5336 1165 5340
rect 1159 5333 1161 5335
rect 1164 5333 1166 5336
rect 1078 5322 1080 5325
rect 1019 5317 1021 5319
rect 1055 5317 1057 5319
rect 1083 5321 1085 5325
rect 1214 5330 1216 5332
rect 1232 5329 1234 5332
rect 1237 5330 1239 5332
rect 1257 5329 1259 5332
rect 1278 5329 1280 5332
rect 1304 5329 1306 5332
rect 1309 5330 1311 5332
rect 1332 5330 1334 5332
rect 1348 5329 1350 5332
rect 1364 5330 1366 5332
rect 1279 5325 1280 5329
rect 1768 5326 1770 5331
rect 1773 5326 1775 5328
rect 1910 5327 1912 5349
rect 1964 5345 1966 5347
rect 1933 5343 1935 5345
rect 1938 5340 1940 5345
rect 1938 5336 1939 5340
rect 1933 5333 1935 5335
rect 1938 5333 1940 5336
rect 1159 5322 1161 5325
rect 1109 5317 1111 5319
rect 1136 5317 1138 5319
rect 1164 5321 1166 5325
rect 1232 5322 1234 5325
rect 1278 5322 1280 5325
rect 1304 5322 1306 5325
rect 1348 5322 1350 5325
rect 1964 5327 1966 5341
rect 2000 5327 2002 5349
rect 2054 5345 2056 5347
rect 2023 5343 2025 5345
rect 2028 5340 2030 5345
rect 2028 5336 2029 5340
rect 2023 5333 2025 5335
rect 2028 5333 2030 5336
rect 1933 5322 1935 5325
rect 1768 5316 1770 5318
rect 1768 5306 1770 5308
rect 1773 5306 1775 5318
rect 1910 5317 1912 5319
rect 1938 5321 1940 5325
rect 2054 5327 2056 5341
rect 2081 5327 2083 5349
rect 2104 5343 2106 5345
rect 2109 5340 2111 5345
rect 2159 5340 2161 5354
rect 2177 5352 2179 5354
rect 2182 5349 2184 5354
rect 2182 5345 2188 5349
rect 2177 5340 2179 5342
rect 2182 5340 2184 5345
rect 2202 5340 2204 5354
rect 2223 5352 2225 5354
rect 2249 5352 2251 5354
rect 2254 5349 2256 5354
rect 2254 5345 2260 5349
rect 2223 5340 2225 5342
rect 2249 5340 2251 5342
rect 2254 5340 2256 5345
rect 2277 5340 2279 5354
rect 2293 5352 2295 5354
rect 2293 5340 2295 5342
rect 2309 5340 2311 5354
rect 2109 5336 2110 5340
rect 2104 5333 2106 5335
rect 2109 5333 2111 5336
rect 2023 5322 2025 5325
rect 1964 5317 1966 5319
rect 2000 5317 2002 5319
rect 2028 5321 2030 5325
rect 2159 5330 2161 5332
rect 2177 5329 2179 5332
rect 2182 5330 2184 5332
rect 2202 5329 2204 5332
rect 2223 5329 2225 5332
rect 2249 5329 2251 5332
rect 2254 5330 2256 5332
rect 2277 5330 2279 5332
rect 2293 5329 2295 5332
rect 2309 5330 2311 5332
rect 2224 5325 2225 5329
rect 2104 5322 2106 5325
rect 2054 5317 2056 5319
rect 2081 5317 2083 5319
rect 2109 5321 2111 5325
rect 2177 5322 2179 5325
rect 2223 5322 2225 5325
rect 2249 5322 2251 5325
rect 2293 5322 2295 5325
rect 1232 5301 1234 5304
rect 1278 5301 1280 5304
rect 1304 5301 1306 5304
rect 1348 5301 1350 5304
rect 1279 5297 1280 5301
rect 1768 5299 1770 5302
rect 1773 5299 1775 5302
rect 2177 5301 2179 5304
rect 2223 5301 2225 5304
rect 2249 5301 2251 5304
rect 2293 5301 2295 5304
rect 1054 5292 1056 5297
rect 1059 5292 1061 5294
rect 1159 5292 1161 5297
rect 1214 5294 1216 5296
rect 1232 5294 1234 5297
rect 1237 5294 1239 5296
rect 1257 5294 1259 5297
rect 1278 5294 1280 5297
rect 1304 5294 1306 5297
rect 1309 5294 1311 5296
rect 1332 5294 1334 5296
rect 1348 5294 1350 5297
rect 1364 5294 1366 5296
rect 2224 5297 2225 5301
rect 1164 5292 1166 5294
rect 1999 5292 2001 5297
rect 2004 5292 2006 5294
rect 2104 5292 2106 5297
rect 2159 5294 2161 5296
rect 2177 5294 2179 5297
rect 2182 5294 2184 5296
rect 2202 5294 2204 5297
rect 2223 5294 2225 5297
rect 2249 5294 2251 5297
rect 2254 5294 2256 5296
rect 2277 5294 2279 5296
rect 2293 5294 2295 5297
rect 2309 5294 2311 5296
rect 2109 5292 2111 5294
rect 1054 5282 1056 5284
rect 1054 5272 1056 5274
rect 1059 5272 1061 5284
rect 1159 5282 1161 5284
rect 1159 5272 1161 5274
rect 1164 5272 1166 5284
rect 1214 5272 1216 5286
rect 1232 5284 1234 5286
rect 1237 5281 1239 5286
rect 1237 5277 1243 5281
rect 1232 5272 1234 5274
rect 1237 5272 1239 5277
rect 1257 5272 1259 5286
rect 1278 5284 1280 5286
rect 1304 5284 1306 5286
rect 1309 5281 1311 5286
rect 1309 5277 1315 5281
rect 1278 5272 1280 5274
rect 1304 5272 1306 5274
rect 1309 5272 1311 5277
rect 1332 5272 1334 5286
rect 1348 5284 1350 5286
rect 1348 5272 1350 5274
rect 1364 5272 1366 5286
rect 1560 5281 1562 5283
rect 1613 5281 1615 5283
rect 1999 5282 2001 5284
rect 1999 5272 2001 5274
rect 2004 5272 2006 5284
rect 2104 5282 2106 5284
rect 2104 5272 2106 5274
rect 2109 5272 2111 5284
rect 2159 5272 2161 5286
rect 2177 5284 2179 5286
rect 2182 5281 2184 5286
rect 2182 5277 2188 5281
rect 2177 5272 2179 5274
rect 2182 5272 2184 5277
rect 2202 5272 2204 5286
rect 2223 5284 2225 5286
rect 2249 5284 2251 5286
rect 2254 5281 2256 5286
rect 2254 5277 2260 5281
rect 2223 5272 2225 5274
rect 2249 5272 2251 5274
rect 2254 5272 2256 5277
rect 2277 5272 2279 5286
rect 2293 5284 2295 5286
rect 2293 5272 2295 5274
rect 2309 5272 2311 5286
rect 1054 5265 1056 5268
rect 1059 5265 1061 5268
rect 1159 5265 1161 5268
rect 1164 5265 1166 5268
rect 1214 5266 1216 5268
rect 1232 5263 1234 5268
rect 1237 5266 1239 5268
rect 1257 5266 1259 5268
rect 1278 5264 1280 5268
rect 1232 5259 1233 5263
rect 1278 5260 1279 5264
rect 1304 5263 1306 5268
rect 1309 5266 1311 5268
rect 1332 5266 1334 5268
rect 1348 5264 1350 5268
rect 1364 5266 1366 5268
rect 1232 5257 1234 5259
rect 1278 5256 1280 5260
rect 1304 5259 1305 5263
rect 1348 5260 1349 5264
rect 1560 5261 1562 5269
rect 1613 5261 1615 5269
rect 1999 5265 2001 5268
rect 2004 5265 2006 5268
rect 2104 5265 2106 5268
rect 2109 5265 2111 5268
rect 2159 5266 2161 5268
rect 2177 5263 2179 5268
rect 2182 5266 2184 5268
rect 2202 5266 2204 5268
rect 2223 5264 2225 5268
rect 1304 5257 1306 5259
rect 1348 5257 1350 5260
rect 2177 5259 2178 5263
rect 2223 5260 2224 5264
rect 2249 5263 2251 5268
rect 2254 5266 2256 5268
rect 2277 5266 2279 5268
rect 2293 5264 2295 5268
rect 2309 5266 2311 5268
rect 2177 5257 2179 5259
rect 1560 5249 1562 5257
rect 1613 5249 1615 5257
rect 2223 5256 2225 5260
rect 2249 5259 2250 5263
rect 2293 5260 2294 5264
rect 2249 5257 2251 5259
rect 2293 5257 2295 5260
rect 1745 5250 1747 5252
rect 1232 5235 1234 5237
rect 1232 5231 1233 5235
rect 1278 5234 1280 5238
rect 1304 5235 1306 5237
rect 1214 5226 1216 5228
rect 1232 5226 1234 5231
rect 1278 5230 1279 5234
rect 1304 5231 1305 5235
rect 1348 5234 1350 5237
rect 1237 5226 1239 5228
rect 1257 5226 1259 5228
rect 1278 5226 1280 5230
rect 1304 5226 1306 5231
rect 1348 5230 1349 5234
rect 1309 5226 1311 5228
rect 1332 5226 1334 5228
rect 1348 5226 1350 5230
rect 1364 5226 1366 5228
rect 1031 5221 1033 5223
rect 1054 5217 1056 5222
rect 1136 5221 1138 5223
rect 1059 5217 1061 5219
rect 1159 5217 1161 5222
rect 1164 5217 1166 5219
rect 1031 5195 1033 5217
rect 1085 5213 1087 5215
rect 1054 5211 1056 5213
rect 1059 5208 1061 5213
rect 1059 5204 1060 5208
rect 1054 5201 1056 5203
rect 1059 5201 1061 5204
rect 1085 5195 1087 5209
rect 1136 5195 1138 5217
rect 1159 5211 1161 5213
rect 1164 5208 1166 5213
rect 1214 5208 1216 5222
rect 1232 5220 1234 5222
rect 1237 5217 1239 5222
rect 1237 5213 1243 5217
rect 1232 5208 1234 5210
rect 1237 5208 1239 5213
rect 1257 5208 1259 5222
rect 1278 5220 1280 5222
rect 1304 5220 1306 5222
rect 1309 5217 1311 5222
rect 1309 5213 1315 5217
rect 1278 5208 1280 5210
rect 1304 5208 1306 5210
rect 1309 5208 1311 5213
rect 1332 5208 1334 5222
rect 1348 5220 1350 5222
rect 1348 5208 1350 5210
rect 1364 5208 1366 5222
rect 1768 5246 1770 5251
rect 1773 5246 1775 5248
rect 1745 5224 1747 5246
rect 1799 5242 1801 5244
rect 1768 5240 1770 5242
rect 1773 5237 1775 5242
rect 1773 5233 1774 5237
rect 1768 5230 1770 5232
rect 1773 5230 1775 5233
rect 1560 5216 1562 5219
rect 1613 5216 1615 5219
rect 1799 5224 1801 5238
rect 2177 5235 2179 5237
rect 2177 5231 2178 5235
rect 2223 5234 2225 5238
rect 2249 5235 2251 5237
rect 2159 5226 2161 5228
rect 2177 5226 2179 5231
rect 2223 5230 2224 5234
rect 2249 5231 2250 5235
rect 2293 5234 2295 5237
rect 2182 5226 2184 5228
rect 2202 5226 2204 5228
rect 2223 5226 2225 5230
rect 2249 5226 2251 5231
rect 2293 5230 2294 5234
rect 2254 5226 2256 5228
rect 2277 5226 2279 5228
rect 2293 5226 2295 5230
rect 2309 5226 2311 5228
rect 1768 5219 1770 5222
rect 1745 5214 1747 5216
rect 1773 5218 1775 5222
rect 1976 5221 1978 5223
rect 1999 5217 2001 5222
rect 2081 5221 2083 5223
rect 2004 5217 2006 5219
rect 2104 5217 2106 5222
rect 2109 5217 2111 5219
rect 1799 5214 1801 5216
rect 1164 5204 1165 5208
rect 1159 5201 1161 5203
rect 1164 5201 1166 5204
rect 1054 5190 1056 5193
rect 1031 5185 1033 5187
rect 1059 5189 1061 5193
rect 1214 5198 1216 5200
rect 1232 5197 1234 5200
rect 1237 5198 1239 5200
rect 1257 5197 1259 5200
rect 1278 5197 1280 5200
rect 1304 5197 1306 5200
rect 1309 5198 1311 5200
rect 1332 5198 1334 5200
rect 1348 5197 1350 5200
rect 1364 5198 1366 5200
rect 1279 5193 1280 5197
rect 1976 5195 1978 5217
rect 2030 5213 2032 5215
rect 1999 5211 2001 5213
rect 2004 5208 2006 5213
rect 2004 5204 2005 5208
rect 1999 5201 2001 5203
rect 2004 5201 2006 5204
rect 1159 5190 1161 5193
rect 1085 5185 1087 5187
rect 1136 5185 1138 5187
rect 1164 5189 1166 5193
rect 1232 5190 1234 5193
rect 1278 5190 1280 5193
rect 1304 5190 1306 5193
rect 1348 5190 1350 5193
rect 2030 5195 2032 5209
rect 2081 5195 2083 5217
rect 2104 5211 2106 5213
rect 2109 5208 2111 5213
rect 2159 5208 2161 5222
rect 2177 5220 2179 5222
rect 2182 5217 2184 5222
rect 2182 5213 2188 5217
rect 2177 5208 2179 5210
rect 2182 5208 2184 5213
rect 2202 5208 2204 5222
rect 2223 5220 2225 5222
rect 2249 5220 2251 5222
rect 2254 5217 2256 5222
rect 2254 5213 2260 5217
rect 2223 5208 2225 5210
rect 2249 5208 2251 5210
rect 2254 5208 2256 5213
rect 2277 5208 2279 5222
rect 2293 5220 2295 5222
rect 2293 5208 2295 5210
rect 2309 5208 2311 5222
rect 2109 5204 2110 5208
rect 2104 5201 2106 5203
rect 2109 5201 2111 5204
rect 1999 5190 2001 5193
rect 1976 5185 1978 5187
rect 2004 5189 2006 5193
rect 2159 5198 2161 5200
rect 2177 5197 2179 5200
rect 2182 5198 2184 5200
rect 2202 5197 2204 5200
rect 2223 5197 2225 5200
rect 2249 5197 2251 5200
rect 2254 5198 2256 5200
rect 2277 5198 2279 5200
rect 2293 5197 2295 5200
rect 2309 5198 2311 5200
rect 2224 5193 2225 5197
rect 2104 5190 2106 5193
rect 2030 5185 2032 5187
rect 2081 5185 2083 5187
rect 2109 5189 2111 5193
rect 2177 5190 2179 5193
rect 2223 5190 2225 5193
rect 2249 5190 2251 5193
rect 2293 5190 2295 5193
rect 1232 5169 1234 5172
rect 1278 5169 1280 5172
rect 1304 5169 1306 5172
rect 1348 5169 1350 5172
rect 1078 5161 1080 5166
rect 1083 5161 1085 5163
rect 1159 5161 1161 5166
rect 1279 5165 1280 5169
rect 2177 5169 2179 5172
rect 2223 5169 2225 5172
rect 2249 5169 2251 5172
rect 2293 5169 2295 5172
rect 1164 5161 1166 5163
rect 1214 5162 1216 5164
rect 1232 5162 1234 5165
rect 1237 5162 1239 5164
rect 1257 5162 1259 5165
rect 1278 5162 1280 5165
rect 1304 5162 1306 5165
rect 1309 5162 1311 5164
rect 1332 5162 1334 5164
rect 1348 5162 1350 5165
rect 1364 5162 1366 5164
rect 2023 5161 2025 5166
rect 2028 5161 2030 5163
rect 2104 5161 2106 5166
rect 2224 5165 2225 5169
rect 2109 5161 2111 5163
rect 2159 5162 2161 5164
rect 2177 5162 2179 5165
rect 2182 5162 2184 5164
rect 2202 5162 2204 5165
rect 2223 5162 2225 5165
rect 2249 5162 2251 5165
rect 2254 5162 2256 5164
rect 2277 5162 2279 5164
rect 2293 5162 2295 5165
rect 2309 5162 2311 5164
rect 1078 5151 1080 5153
rect 1078 5141 1080 5143
rect 1083 5141 1085 5153
rect 1159 5151 1161 5153
rect 1159 5141 1161 5143
rect 1164 5141 1166 5153
rect 1214 5140 1216 5154
rect 1232 5152 1234 5154
rect 1237 5149 1239 5154
rect 1237 5145 1243 5149
rect 1232 5140 1234 5142
rect 1237 5140 1239 5145
rect 1257 5140 1259 5154
rect 1278 5152 1280 5154
rect 1304 5152 1306 5154
rect 1309 5149 1311 5154
rect 1309 5145 1315 5149
rect 1278 5140 1280 5142
rect 1304 5140 1306 5142
rect 1309 5140 1311 5145
rect 1332 5140 1334 5154
rect 1348 5152 1350 5154
rect 1348 5140 1350 5142
rect 1364 5140 1366 5154
rect 1614 5150 1616 5152
rect 1619 5150 1621 5153
rect 1635 5150 1637 5152
rect 1651 5150 1653 5152
rect 1656 5150 1658 5155
rect 1677 5150 1679 5155
rect 1693 5150 1695 5152
rect 1709 5150 1711 5152
rect 1714 5150 1716 5155
rect 1730 5150 1732 5152
rect 2023 5151 2025 5153
rect 1078 5134 1080 5137
rect 1083 5134 1085 5137
rect 1159 5134 1161 5137
rect 1164 5134 1166 5137
rect 1614 5136 1616 5146
rect 1619 5139 1621 5146
rect 1214 5134 1216 5136
rect 1232 5131 1234 5136
rect 1237 5134 1239 5136
rect 1257 5134 1259 5136
rect 1278 5132 1280 5136
rect 1232 5127 1233 5131
rect 1278 5128 1279 5132
rect 1304 5131 1306 5136
rect 1309 5134 1311 5136
rect 1332 5134 1334 5136
rect 1348 5132 1350 5136
rect 1364 5134 1366 5136
rect 1232 5125 1234 5127
rect 1278 5124 1280 5128
rect 1304 5127 1305 5131
rect 1348 5128 1349 5132
rect 1304 5125 1306 5127
rect 1348 5125 1350 5128
rect 1614 5127 1616 5132
rect 1619 5127 1621 5129
rect 1635 5127 1637 5146
rect 1651 5143 1653 5146
rect 1656 5144 1658 5146
rect 1677 5144 1679 5146
rect 1651 5127 1653 5136
rect 1693 5134 1695 5146
rect 1709 5143 1711 5146
rect 1714 5144 1716 5146
rect 1656 5127 1658 5129
rect 1677 5127 1679 5129
rect 1693 5127 1695 5130
rect 1709 5127 1711 5136
rect 1714 5127 1716 5129
rect 1730 5127 1732 5146
rect 2023 5141 2025 5143
rect 2028 5141 2030 5153
rect 2104 5151 2106 5153
rect 2104 5141 2106 5143
rect 2109 5141 2111 5153
rect 2159 5140 2161 5154
rect 2177 5152 2179 5154
rect 2182 5149 2184 5154
rect 2182 5145 2188 5149
rect 2177 5140 2179 5142
rect 2182 5140 2184 5145
rect 2202 5140 2204 5154
rect 2223 5152 2225 5154
rect 2249 5152 2251 5154
rect 2254 5149 2256 5154
rect 2254 5145 2260 5149
rect 2223 5140 2225 5142
rect 2249 5140 2251 5142
rect 2254 5140 2256 5145
rect 2277 5140 2279 5154
rect 2293 5152 2295 5154
rect 2293 5140 2295 5142
rect 2309 5140 2311 5154
rect 2559 5150 2561 5152
rect 2564 5150 2566 5153
rect 2580 5150 2582 5152
rect 2596 5150 2598 5152
rect 2601 5150 2603 5155
rect 2622 5150 2624 5155
rect 2638 5150 2640 5152
rect 2654 5150 2656 5152
rect 2659 5150 2661 5155
rect 2675 5150 2677 5152
rect 2023 5134 2025 5137
rect 2028 5134 2030 5137
rect 2104 5134 2106 5137
rect 2109 5134 2111 5137
rect 2559 5136 2561 5146
rect 2564 5139 2566 5146
rect 2159 5134 2161 5136
rect 2177 5131 2179 5136
rect 2182 5134 2184 5136
rect 2202 5134 2204 5136
rect 2223 5132 2225 5136
rect 2177 5127 2178 5131
rect 2223 5128 2224 5132
rect 2249 5131 2251 5136
rect 2254 5134 2256 5136
rect 2277 5134 2279 5136
rect 2293 5132 2295 5136
rect 2309 5134 2311 5136
rect 2177 5125 2179 5127
rect 2223 5124 2225 5128
rect 2249 5127 2250 5131
rect 2293 5128 2294 5132
rect 2249 5125 2251 5127
rect 2293 5125 2295 5128
rect 2559 5127 2561 5132
rect 2564 5127 2566 5129
rect 2580 5127 2582 5146
rect 2596 5143 2598 5146
rect 2601 5144 2603 5146
rect 2622 5144 2624 5146
rect 2596 5127 2598 5136
rect 2638 5134 2640 5146
rect 2654 5143 2656 5146
rect 2659 5144 2661 5146
rect 2601 5127 2603 5129
rect 2622 5127 2624 5129
rect 2638 5127 2640 5130
rect 2654 5127 2656 5136
rect 2659 5127 2661 5129
rect 2675 5127 2677 5146
rect 1614 5117 1616 5119
rect 1619 5116 1621 5119
rect 1635 5117 1637 5119
rect 1651 5117 1653 5119
rect 1656 5116 1658 5119
rect 1677 5116 1679 5119
rect 1693 5116 1695 5119
rect 1709 5117 1711 5119
rect 1714 5116 1716 5119
rect 1730 5117 1732 5119
rect 2559 5117 2561 5119
rect 2564 5116 2566 5119
rect 2580 5117 2582 5119
rect 2596 5117 2598 5119
rect 2601 5116 2603 5119
rect 2622 5116 2624 5119
rect 2638 5116 2640 5119
rect 2654 5117 2656 5119
rect 2659 5116 2661 5119
rect 2675 5117 2677 5119
rect 1232 5103 1234 5105
rect 1232 5099 1233 5103
rect 1278 5102 1280 5106
rect 1304 5103 1306 5105
rect 1214 5094 1216 5096
rect 1232 5094 1234 5099
rect 1278 5098 1279 5102
rect 1304 5099 1305 5103
rect 1348 5102 1350 5105
rect 2177 5103 2179 5105
rect 1237 5094 1239 5096
rect 1257 5094 1259 5096
rect 1278 5094 1280 5098
rect 1304 5094 1306 5099
rect 1348 5098 1349 5102
rect 2177 5099 2178 5103
rect 2223 5102 2225 5106
rect 2249 5103 2251 5105
rect 1309 5094 1311 5096
rect 1332 5094 1334 5096
rect 1348 5094 1350 5098
rect 1364 5094 1366 5096
rect 1714 5094 1716 5096
rect 2159 5094 2161 5096
rect 2177 5094 2179 5099
rect 2223 5098 2224 5102
rect 2249 5099 2250 5103
rect 2293 5102 2295 5105
rect 2182 5094 2184 5096
rect 2202 5094 2204 5096
rect 2223 5094 2225 5098
rect 2249 5094 2251 5099
rect 2293 5098 2294 5102
rect 2254 5094 2256 5096
rect 2277 5094 2279 5096
rect 2293 5094 2295 5098
rect 2309 5094 2311 5096
rect 2659 5094 2661 5096
rect 1055 5089 1057 5091
rect 1078 5085 1080 5090
rect 1136 5089 1138 5091
rect 1083 5085 1085 5087
rect 1159 5085 1161 5090
rect 1164 5085 1166 5087
rect 1055 5063 1057 5085
rect 1109 5081 1111 5083
rect 1078 5079 1080 5081
rect 1083 5076 1085 5081
rect 1083 5072 1084 5076
rect 1078 5069 1080 5071
rect 1083 5069 1085 5072
rect 1109 5063 1111 5077
rect 1136 5063 1138 5085
rect 1190 5081 1192 5083
rect 1159 5079 1161 5081
rect 1164 5076 1166 5081
rect 1164 5072 1165 5076
rect 1159 5069 1161 5071
rect 1164 5069 1166 5072
rect 1078 5058 1080 5061
rect 1055 5053 1057 5055
rect 1083 5057 1085 5061
rect 1190 5063 1192 5077
rect 1214 5076 1216 5090
rect 1232 5088 1234 5090
rect 1237 5085 1239 5090
rect 1237 5081 1243 5085
rect 1232 5076 1234 5078
rect 1237 5076 1239 5081
rect 1257 5076 1259 5090
rect 1278 5088 1280 5090
rect 1304 5088 1306 5090
rect 1309 5085 1311 5090
rect 1309 5081 1315 5085
rect 1278 5076 1280 5078
rect 1304 5076 1306 5078
rect 1309 5076 1311 5081
rect 1332 5076 1334 5090
rect 1348 5088 1350 5090
rect 1348 5076 1350 5078
rect 1364 5076 1366 5090
rect 1714 5087 1716 5090
rect 2000 5089 2002 5091
rect 1597 5085 1599 5087
rect 2023 5085 2025 5090
rect 2081 5089 2083 5091
rect 2028 5085 2030 5087
rect 2104 5085 2106 5090
rect 2109 5085 2111 5087
rect 1597 5078 1599 5081
rect 1214 5066 1216 5068
rect 1232 5065 1234 5068
rect 1237 5066 1239 5068
rect 1257 5065 1259 5068
rect 1278 5065 1280 5068
rect 1304 5065 1306 5068
rect 1309 5066 1311 5068
rect 1332 5066 1334 5068
rect 1348 5065 1350 5068
rect 1364 5066 1366 5068
rect 1159 5058 1161 5061
rect 1109 5053 1111 5055
rect 1136 5053 1138 5055
rect 1164 5057 1166 5061
rect 1279 5061 1280 5065
rect 1232 5058 1234 5061
rect 1278 5058 1280 5061
rect 1304 5058 1306 5061
rect 1348 5058 1350 5061
rect 2000 5063 2002 5085
rect 2054 5081 2056 5083
rect 2023 5079 2025 5081
rect 2028 5076 2030 5081
rect 2028 5072 2029 5076
rect 2023 5069 2025 5071
rect 2028 5069 2030 5072
rect 1190 5053 1192 5055
rect 2054 5063 2056 5077
rect 2081 5063 2083 5085
rect 2135 5081 2137 5083
rect 2104 5079 2106 5081
rect 2109 5076 2111 5081
rect 2109 5072 2110 5076
rect 2104 5069 2106 5071
rect 2109 5069 2111 5072
rect 2023 5058 2025 5061
rect 1605 5048 1607 5050
rect 1621 5048 1623 5053
rect 1626 5048 1628 5050
rect 1642 5048 1644 5050
rect 1658 5048 1660 5053
rect 1679 5048 1681 5053
rect 2000 5053 2002 5055
rect 2028 5057 2030 5061
rect 2135 5063 2137 5077
rect 2159 5076 2161 5090
rect 2177 5088 2179 5090
rect 2182 5085 2184 5090
rect 2182 5081 2188 5085
rect 2177 5076 2179 5078
rect 2182 5076 2184 5081
rect 2202 5076 2204 5090
rect 2223 5088 2225 5090
rect 2249 5088 2251 5090
rect 2254 5085 2256 5090
rect 2254 5081 2260 5085
rect 2223 5076 2225 5078
rect 2249 5076 2251 5078
rect 2254 5076 2256 5081
rect 2277 5076 2279 5090
rect 2293 5088 2295 5090
rect 2293 5076 2295 5078
rect 2309 5076 2311 5090
rect 2659 5087 2661 5090
rect 2542 5085 2544 5087
rect 2542 5078 2544 5081
rect 2159 5066 2161 5068
rect 2177 5065 2179 5068
rect 2182 5066 2184 5068
rect 2202 5065 2204 5068
rect 2223 5065 2225 5068
rect 2249 5065 2251 5068
rect 2254 5066 2256 5068
rect 2277 5066 2279 5068
rect 2293 5065 2295 5068
rect 2309 5066 2311 5068
rect 2104 5058 2106 5061
rect 2054 5053 2056 5055
rect 2081 5053 2083 5055
rect 2109 5057 2111 5061
rect 2224 5061 2225 5065
rect 2177 5058 2179 5061
rect 2223 5058 2225 5061
rect 2249 5058 2251 5061
rect 2293 5058 2295 5061
rect 2135 5053 2137 5055
rect 1684 5048 1686 5050
rect 1700 5048 1702 5050
rect 1716 5048 1718 5051
rect 1721 5048 1723 5050
rect 2550 5048 2552 5050
rect 2566 5048 2568 5053
rect 2571 5048 2573 5050
rect 2587 5048 2589 5050
rect 2603 5048 2605 5053
rect 2624 5048 2626 5053
rect 2629 5048 2631 5050
rect 2645 5048 2647 5050
rect 2661 5048 2663 5051
rect 2666 5048 2668 5050
rect 1605 5025 1607 5044
rect 1621 5042 1623 5044
rect 1626 5041 1628 5044
rect 1621 5025 1623 5027
rect 1626 5025 1628 5034
rect 1642 5032 1644 5044
rect 1658 5042 1660 5044
rect 1679 5042 1681 5044
rect 1684 5041 1686 5044
rect 1642 5025 1644 5028
rect 1658 5025 1660 5027
rect 1679 5025 1681 5027
rect 1684 5025 1686 5034
rect 1700 5025 1702 5044
rect 1716 5037 1718 5044
rect 1721 5034 1723 5044
rect 1716 5025 1718 5027
rect 1721 5025 1723 5030
rect 2550 5025 2552 5044
rect 2566 5042 2568 5044
rect 2571 5041 2573 5044
rect 2566 5025 2568 5027
rect 2571 5025 2573 5034
rect 2587 5032 2589 5044
rect 2603 5042 2605 5044
rect 2624 5042 2626 5044
rect 2629 5041 2631 5044
rect 2587 5025 2589 5028
rect 2603 5025 2605 5027
rect 2624 5025 2626 5027
rect 2629 5025 2631 5034
rect 2645 5025 2647 5044
rect 2661 5037 2663 5044
rect 2666 5034 2668 5044
rect 2661 5025 2663 5027
rect 2666 5025 2668 5030
rect 857 5015 859 5017
rect 873 5015 875 5020
rect 878 5015 880 5017
rect 894 5015 896 5017
rect 910 5015 912 5020
rect 931 5015 933 5020
rect 936 5015 938 5017
rect 952 5015 954 5017
rect 968 5015 970 5018
rect 973 5015 975 5017
rect 989 5015 991 5017
rect 1005 5015 1007 5020
rect 1010 5015 1012 5017
rect 1026 5015 1028 5017
rect 1042 5015 1044 5020
rect 1063 5015 1065 5020
rect 1068 5015 1070 5017
rect 1084 5015 1086 5017
rect 1100 5015 1102 5018
rect 1105 5015 1107 5017
rect 1121 5015 1123 5017
rect 1137 5015 1139 5020
rect 1142 5015 1144 5017
rect 1158 5015 1160 5017
rect 1174 5015 1176 5020
rect 1195 5015 1197 5020
rect 1200 5015 1202 5017
rect 1216 5015 1218 5017
rect 1232 5015 1234 5018
rect 1237 5015 1239 5017
rect 1253 5015 1255 5017
rect 1269 5015 1271 5020
rect 1274 5015 1276 5017
rect 1290 5015 1292 5017
rect 1306 5015 1308 5020
rect 1327 5015 1329 5020
rect 1332 5015 1334 5017
rect 1348 5015 1350 5017
rect 1364 5015 1366 5018
rect 1369 5015 1371 5017
rect 1605 5015 1607 5017
rect 1621 5014 1623 5017
rect 1626 5015 1628 5017
rect 1642 5014 1644 5017
rect 1658 5014 1660 5017
rect 1679 5014 1681 5017
rect 1684 5015 1686 5017
rect 1700 5015 1702 5017
rect 1716 5014 1718 5017
rect 1721 5015 1723 5017
rect 1802 5015 1804 5017
rect 1818 5015 1820 5020
rect 1823 5015 1825 5017
rect 1839 5015 1841 5017
rect 1855 5015 1857 5020
rect 1876 5015 1878 5020
rect 1881 5015 1883 5017
rect 1897 5015 1899 5017
rect 1913 5015 1915 5018
rect 1918 5015 1920 5017
rect 1934 5015 1936 5017
rect 1950 5015 1952 5020
rect 1955 5015 1957 5017
rect 1971 5015 1973 5017
rect 1987 5015 1989 5020
rect 2008 5015 2010 5020
rect 2013 5015 2015 5017
rect 2029 5015 2031 5017
rect 2045 5015 2047 5018
rect 2050 5015 2052 5017
rect 2066 5015 2068 5017
rect 2082 5015 2084 5020
rect 2087 5015 2089 5017
rect 2103 5015 2105 5017
rect 2119 5015 2121 5020
rect 2140 5015 2142 5020
rect 2145 5015 2147 5017
rect 2161 5015 2163 5017
rect 2177 5015 2179 5018
rect 2182 5015 2184 5017
rect 2198 5015 2200 5017
rect 2214 5015 2216 5020
rect 2219 5015 2221 5017
rect 2235 5015 2237 5017
rect 2251 5015 2253 5020
rect 2272 5015 2274 5020
rect 2277 5015 2279 5017
rect 2293 5015 2295 5017
rect 2309 5015 2311 5018
rect 2314 5015 2316 5017
rect 2550 5015 2552 5017
rect 857 5004 859 5011
rect 873 5009 875 5011
rect 878 5008 880 5011
rect 857 4992 859 5000
rect 873 4992 875 4994
rect 878 4992 880 5001
rect 894 4999 896 5011
rect 910 5009 912 5011
rect 931 5009 933 5011
rect 936 5008 938 5011
rect 894 4992 896 4995
rect 910 4992 912 4994
rect 931 4992 933 4994
rect 936 4992 938 5001
rect 952 4992 954 5011
rect 968 5004 970 5011
rect 973 5001 975 5011
rect 989 5004 991 5011
rect 1005 5009 1007 5011
rect 1010 5008 1012 5011
rect 968 4992 970 4994
rect 973 4992 975 4997
rect 989 4992 991 5000
rect 1005 4992 1007 4994
rect 1010 4992 1012 5001
rect 1026 4999 1028 5011
rect 1042 5009 1044 5011
rect 1063 5009 1065 5011
rect 1068 5008 1070 5011
rect 1026 4992 1028 4995
rect 1042 4992 1044 4994
rect 1063 4992 1065 4994
rect 1068 4992 1070 5001
rect 1084 4992 1086 5011
rect 1100 5004 1102 5011
rect 1105 5001 1107 5011
rect 1121 5004 1123 5011
rect 1137 5009 1139 5011
rect 1142 5008 1144 5011
rect 1100 4992 1102 4994
rect 1105 4992 1107 4997
rect 1121 4992 1123 5000
rect 1137 4992 1139 4994
rect 1142 4992 1144 5001
rect 1158 4999 1160 5011
rect 1174 5009 1176 5011
rect 1195 5009 1197 5011
rect 1200 5008 1202 5011
rect 1158 4992 1160 4995
rect 1174 4992 1176 4994
rect 1195 4992 1197 4994
rect 1200 4992 1202 5001
rect 1216 4992 1218 5011
rect 1232 5004 1234 5011
rect 1237 5001 1239 5011
rect 1253 5004 1255 5011
rect 1269 5009 1271 5011
rect 1274 5008 1276 5011
rect 1232 4992 1234 4994
rect 1237 4992 1239 4997
rect 1253 4992 1255 5000
rect 1269 4992 1271 4994
rect 1274 4992 1276 5001
rect 1290 4999 1292 5011
rect 1306 5009 1308 5011
rect 1327 5009 1329 5011
rect 1332 5008 1334 5011
rect 1290 4992 1292 4995
rect 1306 4992 1308 4994
rect 1327 4992 1329 4994
rect 1332 4992 1334 5001
rect 1348 4992 1350 5011
rect 1364 5004 1366 5011
rect 1369 5001 1371 5011
rect 2566 5014 2568 5017
rect 2571 5015 2573 5017
rect 2587 5014 2589 5017
rect 2603 5014 2605 5017
rect 2624 5014 2626 5017
rect 2629 5015 2631 5017
rect 2645 5015 2647 5017
rect 2661 5014 2663 5017
rect 2666 5015 2668 5017
rect 1802 5004 1804 5011
rect 1818 5009 1820 5011
rect 1823 5008 1825 5011
rect 1364 4992 1366 4994
rect 1369 4992 1371 4997
rect 1802 4992 1804 5000
rect 1818 4992 1820 4994
rect 1823 4992 1825 5001
rect 1839 4999 1841 5011
rect 1855 5009 1857 5011
rect 1876 5009 1878 5011
rect 1881 5008 1883 5011
rect 1839 4992 1841 4995
rect 1855 4992 1857 4994
rect 1876 4992 1878 4994
rect 1881 4992 1883 5001
rect 1897 4992 1899 5011
rect 1913 5004 1915 5011
rect 1918 5001 1920 5011
rect 1934 5004 1936 5011
rect 1950 5009 1952 5011
rect 1955 5008 1957 5011
rect 1913 4992 1915 4994
rect 1918 4992 1920 4997
rect 1934 4992 1936 5000
rect 1950 4992 1952 4994
rect 1955 4992 1957 5001
rect 1971 4999 1973 5011
rect 1987 5009 1989 5011
rect 2008 5009 2010 5011
rect 2013 5008 2015 5011
rect 1971 4992 1973 4995
rect 1987 4992 1989 4994
rect 2008 4992 2010 4994
rect 2013 4992 2015 5001
rect 2029 4992 2031 5011
rect 2045 5004 2047 5011
rect 2050 5001 2052 5011
rect 2066 5004 2068 5011
rect 2082 5009 2084 5011
rect 2087 5008 2089 5011
rect 2045 4992 2047 4994
rect 2050 4992 2052 4997
rect 2066 4992 2068 5000
rect 2082 4992 2084 4994
rect 2087 4992 2089 5001
rect 2103 4999 2105 5011
rect 2119 5009 2121 5011
rect 2140 5009 2142 5011
rect 2145 5008 2147 5011
rect 2103 4992 2105 4995
rect 2119 4992 2121 4994
rect 2140 4992 2142 4994
rect 2145 4992 2147 5001
rect 2161 4992 2163 5011
rect 2177 5004 2179 5011
rect 2182 5001 2184 5011
rect 2198 5004 2200 5011
rect 2214 5009 2216 5011
rect 2219 5008 2221 5011
rect 2177 4992 2179 4994
rect 2182 4992 2184 4997
rect 2198 4992 2200 5000
rect 2214 4992 2216 4994
rect 2219 4992 2221 5001
rect 2235 4999 2237 5011
rect 2251 5009 2253 5011
rect 2272 5009 2274 5011
rect 2277 5008 2279 5011
rect 2235 4992 2237 4995
rect 2251 4992 2253 4994
rect 2272 4992 2274 4994
rect 2277 4992 2279 5001
rect 2293 4992 2295 5011
rect 2309 5004 2311 5011
rect 2314 5001 2316 5011
rect 2309 4992 2311 4994
rect 2314 4992 2316 4997
rect 857 4982 859 4984
rect 873 4981 875 4984
rect 878 4982 880 4984
rect 894 4981 896 4984
rect 910 4981 912 4984
rect 931 4981 933 4984
rect 936 4982 938 4984
rect 952 4982 954 4984
rect 968 4981 970 4984
rect 973 4982 975 4984
rect 989 4982 991 4984
rect 1005 4981 1007 4984
rect 1010 4982 1012 4984
rect 1026 4981 1028 4984
rect 1042 4981 1044 4984
rect 1063 4981 1065 4984
rect 1068 4982 1070 4984
rect 1084 4982 1086 4984
rect 1100 4981 1102 4984
rect 1105 4982 1107 4984
rect 1121 4982 1123 4984
rect 1137 4981 1139 4984
rect 1142 4982 1144 4984
rect 1158 4981 1160 4984
rect 1174 4981 1176 4984
rect 1195 4981 1197 4984
rect 1200 4982 1202 4984
rect 1216 4982 1218 4984
rect 1232 4981 1234 4984
rect 1237 4982 1239 4984
rect 1253 4982 1255 4984
rect 1269 4981 1271 4984
rect 1274 4982 1276 4984
rect 1290 4981 1292 4984
rect 1306 4981 1308 4984
rect 1327 4981 1329 4984
rect 1332 4982 1334 4984
rect 1348 4982 1350 4984
rect 1364 4981 1366 4984
rect 1369 4982 1371 4984
rect 1802 4982 1804 4984
rect 1818 4981 1820 4984
rect 1823 4982 1825 4984
rect 1839 4981 1841 4984
rect 1855 4981 1857 4984
rect 1876 4981 1878 4984
rect 1881 4982 1883 4984
rect 1897 4982 1899 4984
rect 1913 4981 1915 4984
rect 1918 4982 1920 4984
rect 1934 4982 1936 4984
rect 1950 4981 1952 4984
rect 1955 4982 1957 4984
rect 1971 4981 1973 4984
rect 1987 4981 1989 4984
rect 2008 4981 2010 4984
rect 2013 4982 2015 4984
rect 2029 4982 2031 4984
rect 2045 4981 2047 4984
rect 2050 4982 2052 4984
rect 2066 4982 2068 4984
rect 2082 4981 2084 4984
rect 2087 4982 2089 4984
rect 2103 4981 2105 4984
rect 2119 4981 2121 4984
rect 2140 4981 2142 4984
rect 2145 4982 2147 4984
rect 2161 4982 2163 4984
rect 2177 4981 2179 4984
rect 2182 4982 2184 4984
rect 2198 4982 2200 4984
rect 2214 4981 2216 4984
rect 2219 4982 2221 4984
rect 2235 4981 2237 4984
rect 2251 4981 2253 4984
rect 2272 4981 2274 4984
rect 2277 4982 2279 4984
rect 2293 4982 2295 4984
rect 2309 4981 2311 4984
rect 2314 4982 2316 4984
rect 4579 9355 5073 9786
rect 4634 8035 4644 8037
rect 4634 8034 4636 8035
rect 4642 8034 4644 8035
rect 4650 8035 4660 8037
rect 4650 8034 4652 8035
rect 4658 8034 4660 8035
rect 4677 8035 4687 8037
rect 4677 8034 4679 8035
rect 4685 8034 4687 8035
rect 4693 8035 4703 8037
rect 4693 8034 4695 8035
rect 4701 8034 4703 8035
rect 4718 8035 4728 8037
rect 4718 8034 4720 8035
rect 4726 8034 4728 8035
rect 4734 8035 4744 8037
rect 4734 8034 4736 8035
rect 4742 8034 4744 8035
rect 4579 8015 4581 8017
rect 4587 8015 4589 8017
rect 4595 8016 4621 8018
rect 4595 8015 4597 8016
rect 4603 8015 4605 8016
rect 4611 8015 4613 8016
rect 4619 8015 4621 8016
rect 4579 7960 4581 7975
rect 4576 7954 4581 7960
rect 4587 7954 4589 7975
rect 4595 7974 4597 7975
rect 4603 7974 4605 7975
rect 4611 7974 4613 7975
rect 4619 7974 4621 7975
rect 4595 7972 4621 7974
rect 4634 7974 4636 7975
rect 4642 7974 4644 7975
rect 4650 7974 4652 7975
rect 4658 7974 4660 7975
rect 4634 7972 4660 7974
rect 4677 7974 4679 7975
rect 4685 7974 4687 7975
rect 4693 7974 4695 7975
rect 4701 7974 4703 7975
rect 4718 7974 4720 7975
rect 4726 7974 4728 7975
rect 4734 7974 4736 7975
rect 4742 7974 4744 7975
rect 4595 7965 4599 7972
rect 4597 7959 4599 7965
rect 4579 7952 4589 7954
rect 4579 7945 4581 7952
rect 4587 7945 4589 7952
rect 4595 7948 4599 7959
rect 4634 7963 4641 7972
rect 4634 7950 4635 7963
rect 4639 7950 4641 7963
rect 4634 7948 4641 7950
rect 4677 7965 4744 7974
rect 4677 7952 4678 7965
rect 4682 7963 4744 7965
rect 4682 7954 4711 7963
rect 4717 7954 4744 7963
rect 4682 7952 4744 7954
rect 4677 7950 4744 7952
rect 4677 7948 4703 7950
rect 4595 7946 4621 7948
rect 4595 7945 4597 7946
rect 4603 7945 4605 7946
rect 4611 7945 4613 7946
rect 4619 7945 4621 7946
rect 4634 7946 4660 7948
rect 4634 7945 4636 7946
rect 4642 7945 4644 7946
rect 4650 7945 4652 7946
rect 4658 7945 4660 7946
rect 4677 7945 4679 7948
rect 4685 7945 4687 7948
rect 4693 7945 4695 7948
rect 4701 7945 4703 7948
rect 4718 7948 4744 7950
rect 4718 7945 4720 7948
rect 4726 7945 4728 7948
rect 4734 7945 4736 7948
rect 4742 7945 4744 7948
rect 4579 7887 4581 7889
rect 4587 7887 4589 7889
rect 4595 7888 4597 7889
rect 4603 7888 4605 7889
rect 4611 7888 4613 7889
rect 4619 7888 4621 7889
rect 4595 7886 4621 7888
rect 4634 7856 4636 7857
rect 4642 7856 4644 7857
rect 4650 7856 4652 7857
rect 4658 7856 4660 7857
rect 4634 7854 4660 7856
rect 4677 7856 4679 7857
rect 4685 7856 4687 7857
rect 4693 7856 4695 7857
rect 4701 7856 4703 7857
rect 4677 7854 4703 7856
rect 4718 7856 4720 7857
rect 4726 7856 4728 7857
rect 4734 7856 4736 7857
rect 4742 7856 4744 7857
rect 4718 7854 4744 7856
rect 4577 7429 4603 7431
rect 4577 7428 4579 7429
rect 4585 7428 4587 7429
rect 4593 7428 4595 7429
rect 4601 7428 4603 7429
rect 4609 7428 4611 7430
rect 4617 7428 4619 7430
rect 4577 7371 4579 7372
rect 4585 7371 4587 7372
rect 4593 7371 4595 7372
rect 4601 7371 4603 7372
rect 4577 7369 4603 7371
rect 4599 7358 4603 7369
rect 4609 7365 4611 7372
rect 4617 7368 4619 7372
rect 4617 7365 4620 7368
rect 4609 7363 4620 7365
rect 4599 7352 4601 7358
rect 4599 7345 4603 7352
rect 4577 7343 4603 7345
rect 4577 7342 4579 7343
rect 4585 7342 4587 7343
rect 4593 7342 4595 7343
rect 4601 7342 4603 7343
rect 4609 7342 4611 7363
rect 4617 7359 4620 7363
rect 4617 7342 4619 7359
rect 4676 7353 4745 7374
rect 4577 7301 4579 7302
rect 4585 7301 4587 7302
rect 4593 7301 4595 7302
rect 4601 7301 4603 7302
rect 4577 7299 4603 7301
rect 4609 7300 4611 7302
rect 4617 7300 4619 7302
rect 1137 4528 1140 4530
rect 1180 4528 1183 4530
rect 99 4053 1031 4528
rect 1137 4522 1139 4528
rect 1181 4522 1183 4528
rect 1137 4520 1140 4522
rect 1180 4520 1183 4522
rect 1137 4514 1139 4520
rect 1181 4514 1183 4520
rect 1137 4512 1140 4514
rect 1180 4512 1183 4514
rect 1137 4506 1139 4512
rect 1181 4508 1183 4512
rect 1207 4528 1210 4530
rect 1266 4528 1269 4530
rect 1207 4522 1209 4528
rect 1267 4522 1269 4528
rect 1207 4520 1210 4522
rect 1266 4520 1269 4522
rect 1207 4514 1209 4520
rect 1267 4514 1269 4520
rect 1207 4512 1210 4514
rect 1266 4512 1269 4514
rect 1207 4508 1209 4512
rect 1181 4506 1209 4508
rect 1267 4506 1269 4512
rect 1137 4504 1140 4506
rect 1180 4504 1190 4506
rect 1196 4504 1210 4506
rect 1266 4504 1269 4506
rect 2064 4528 2067 4530
rect 2107 4528 2110 4530
rect 2064 4522 2066 4528
rect 2108 4522 2110 4528
rect 2064 4520 2067 4522
rect 2107 4520 2110 4522
rect 2064 4514 2066 4520
rect 2108 4514 2110 4520
rect 2064 4512 2067 4514
rect 2107 4512 2110 4514
rect 2064 4506 2066 4512
rect 2108 4508 2110 4512
rect 2134 4528 2137 4530
rect 2193 4528 2196 4530
rect 2134 4522 2136 4528
rect 2194 4522 2196 4528
rect 2134 4520 2137 4522
rect 2193 4520 2196 4522
rect 2134 4514 2136 4520
rect 2194 4514 2196 4520
rect 2134 4512 2137 4514
rect 2193 4512 2196 4514
rect 2134 4508 2136 4512
rect 2108 4506 2136 4508
rect 2194 4506 2196 4512
rect 2064 4504 2067 4506
rect 2107 4504 2117 4506
rect 2123 4504 2137 4506
rect 2193 4504 2196 4506
rect 2373 4528 2376 4530
rect 2416 4528 2419 4530
rect 2373 4522 2375 4528
rect 2417 4522 2419 4528
rect 2373 4520 2376 4522
rect 2416 4520 2419 4522
rect 2373 4514 2375 4520
rect 2417 4514 2419 4520
rect 2373 4512 2376 4514
rect 2416 4512 2419 4514
rect 2373 4506 2375 4512
rect 2417 4508 2419 4512
rect 2443 4528 2446 4530
rect 2502 4528 2505 4530
rect 2443 4522 2445 4528
rect 2503 4522 2505 4528
rect 2443 4520 2446 4522
rect 2502 4520 2505 4522
rect 2443 4514 2445 4520
rect 2503 4514 2505 4520
rect 2443 4512 2446 4514
rect 2502 4512 2505 4514
rect 2443 4508 2445 4512
rect 2417 4506 2445 4508
rect 2503 4506 2505 4512
rect 2373 4504 2376 4506
rect 2416 4504 2426 4506
rect 2432 4504 2446 4506
rect 2502 4504 2505 4506
rect 2682 4528 2685 4530
rect 2725 4528 2728 4530
rect 2682 4522 2684 4528
rect 2726 4522 2728 4528
rect 2682 4520 2685 4522
rect 2725 4520 2728 4522
rect 2682 4514 2684 4520
rect 2726 4514 2728 4520
rect 2682 4512 2685 4514
rect 2725 4512 2728 4514
rect 2682 4506 2684 4512
rect 2726 4508 2728 4512
rect 2752 4528 2755 4530
rect 2811 4528 2814 4530
rect 2752 4522 2754 4528
rect 2812 4522 2814 4528
rect 2752 4520 2755 4522
rect 2811 4520 2814 4522
rect 2752 4514 2754 4520
rect 2812 4514 2814 4520
rect 2752 4512 2755 4514
rect 2811 4512 2814 4514
rect 2752 4508 2754 4512
rect 2726 4506 2754 4508
rect 2812 4506 2814 4512
rect 2682 4504 2685 4506
rect 2725 4504 2735 4506
rect 2741 4504 2755 4506
rect 2811 4504 2814 4506
rect 2991 4528 2994 4530
rect 3034 4528 3037 4530
rect 2991 4522 2993 4528
rect 3035 4522 3037 4528
rect 2991 4520 2994 4522
rect 3034 4520 3037 4522
rect 2991 4514 2993 4520
rect 3035 4514 3037 4520
rect 2991 4512 2994 4514
rect 3034 4512 3037 4514
rect 2991 4506 2993 4512
rect 3035 4508 3037 4512
rect 3061 4528 3064 4530
rect 3120 4528 3123 4530
rect 3061 4522 3063 4528
rect 3121 4522 3123 4528
rect 3061 4520 3064 4522
rect 3120 4520 3123 4522
rect 3061 4514 3063 4520
rect 3121 4514 3123 4520
rect 3061 4512 3064 4514
rect 3120 4512 3123 4514
rect 3061 4508 3063 4512
rect 3035 4506 3063 4508
rect 3121 4506 3123 4512
rect 2991 4504 2994 4506
rect 3034 4504 3044 4506
rect 3050 4504 3064 4506
rect 3120 4504 3123 4506
rect 3300 4528 3303 4530
rect 3343 4528 3346 4530
rect 3300 4522 3302 4528
rect 3344 4522 3346 4528
rect 3300 4520 3303 4522
rect 3343 4520 3346 4522
rect 3300 4514 3302 4520
rect 3344 4514 3346 4520
rect 3300 4512 3303 4514
rect 3343 4512 3346 4514
rect 3300 4506 3302 4512
rect 3344 4508 3346 4512
rect 3370 4528 3373 4530
rect 3429 4528 3432 4530
rect 4579 4528 5054 4966
rect 3370 4522 3372 4528
rect 3430 4522 3432 4528
rect 3370 4520 3373 4522
rect 3429 4520 3432 4522
rect 3370 4514 3372 4520
rect 3430 4514 3432 4520
rect 3370 4512 3373 4514
rect 3429 4512 3432 4514
rect 3370 4508 3372 4512
rect 3344 4506 3372 4508
rect 3430 4506 3432 4512
rect 3300 4504 3303 4506
rect 3343 4504 3353 4506
rect 3359 4504 3373 4506
rect 3429 4504 3432 4506
rect 1138 4496 1140 4498
rect 1180 4496 1210 4498
rect 1266 4496 1268 4498
rect 2065 4496 2067 4498
rect 2107 4496 2137 4498
rect 2193 4496 2195 4498
rect 2374 4496 2376 4498
rect 2416 4496 2446 4498
rect 2502 4496 2504 4498
rect 2683 4496 2685 4498
rect 2725 4496 2755 4498
rect 2811 4496 2813 4498
rect 2992 4496 2994 4498
rect 3034 4496 3064 4498
rect 3120 4496 3122 4498
rect 3301 4496 3303 4498
rect 3343 4496 3373 4498
rect 3429 4496 3431 4498
rect 1201 4490 1203 4496
rect 2128 4490 2130 4496
rect 2437 4490 2439 4496
rect 2746 4490 2748 4496
rect 3055 4490 3057 4496
rect 3364 4490 3366 4496
rect 1138 4488 1140 4490
rect 1180 4488 1210 4490
rect 1266 4488 1268 4490
rect 2065 4488 2067 4490
rect 2107 4488 2137 4490
rect 2193 4488 2195 4490
rect 2374 4488 2376 4490
rect 2416 4488 2446 4490
rect 2502 4488 2504 4490
rect 2683 4488 2685 4490
rect 2725 4488 2755 4490
rect 2811 4488 2813 4490
rect 2992 4488 2994 4490
rect 3034 4488 3064 4490
rect 3120 4488 3122 4490
rect 3301 4488 3303 4490
rect 3343 4488 3373 4490
rect 3429 4488 3431 4490
rect 1197 4487 1206 4488
rect 2124 4487 2133 4488
rect 2433 4487 2442 4488
rect 2742 4487 2751 4488
rect 3051 4487 3060 4488
rect 3360 4487 3369 4488
rect 1191 4362 1212 4431
rect 2118 4362 2139 4431
rect 2427 4362 2448 4431
rect 2736 4362 2757 4431
rect 3045 4362 3066 4431
rect 3354 4362 3375 4431
rect 4148 4034 5054 4528
<< polycontact >>
rect 1797 9952 1818 9961
rect 1797 9874 1818 9883
rect 2106 9952 2127 9961
rect 2106 9874 2127 9883
rect 2415 9952 2436 9961
rect 2415 9874 2436 9883
rect 2724 9952 2745 9961
rect 2724 9874 2745 9883
rect 3033 9952 3054 9961
rect 3033 9874 3054 9883
rect 3960 9952 3981 9961
rect 3960 9874 3981 9883
rect 1803 9827 1812 9831
rect 2112 9827 2121 9831
rect 2421 9827 2430 9831
rect 2730 9827 2739 9831
rect 3039 9827 3048 9831
rect 3966 9827 3975 9831
rect 1813 9808 1819 9812
rect 2122 9808 2128 9812
rect 2431 9808 2437 9812
rect 2740 9808 2746 9812
rect 3049 9808 3055 9812
rect 3976 9808 3982 9812
rect 455 6351 461 6360
rect 490 6349 494 6362
rect 533 6351 537 6364
rect 575 6349 579 6355
rect 596 6354 600 6360
rect 2861 9333 2865 9337
rect 2898 9333 2902 9337
rect 2918 9333 2922 9337
rect 2956 9333 2960 9337
rect 2993 9333 2997 9337
rect 3030 9333 3034 9337
rect 3050 9333 3054 9337
rect 3088 9333 3092 9337
rect 3125 9333 3129 9337
rect 3162 9333 3166 9337
rect 3182 9333 3186 9337
rect 3220 9333 3224 9337
rect 3257 9333 3261 9337
rect 3294 9333 3298 9337
rect 3314 9333 3318 9337
rect 3352 9333 3356 9337
rect 3806 9333 3810 9337
rect 3843 9333 3847 9337
rect 3863 9333 3867 9337
rect 3901 9333 3905 9337
rect 3938 9333 3942 9337
rect 3975 9333 3979 9337
rect 3995 9333 3999 9337
rect 4033 9333 4037 9337
rect 4070 9333 4074 9337
rect 4107 9333 4111 9337
rect 4127 9333 4131 9337
rect 4165 9333 4169 9337
rect 4202 9333 4206 9337
rect 4239 9333 4243 9337
rect 4259 9333 4263 9337
rect 4297 9333 4301 9337
rect 2855 9313 2859 9317
rect 2873 9315 2877 9319
rect 2509 9300 2513 9304
rect 2546 9300 2550 9304
rect 2566 9300 2570 9304
rect 2604 9300 2608 9304
rect 2933 9315 2937 9319
rect 2891 9306 2895 9313
rect 2949 9306 2953 9313
rect 2970 9310 2974 9314
rect 2987 9313 2991 9317
rect 3005 9315 3009 9319
rect 3065 9315 3069 9319
rect 3023 9306 3027 9313
rect 3081 9306 3085 9313
rect 3102 9310 3106 9314
rect 3119 9313 3123 9317
rect 3137 9315 3141 9319
rect 3197 9315 3201 9319
rect 3155 9306 3159 9313
rect 3213 9306 3217 9313
rect 3234 9310 3238 9314
rect 3251 9313 3255 9317
rect 3269 9315 3273 9319
rect 3329 9315 3333 9319
rect 3287 9306 3291 9313
rect 3345 9306 3349 9313
rect 3366 9310 3370 9314
rect 3800 9313 3804 9317
rect 3818 9315 3822 9319
rect 3454 9300 3458 9304
rect 3491 9300 3495 9304
rect 3511 9300 3515 9304
rect 3549 9300 3553 9304
rect 3878 9315 3882 9319
rect 3836 9306 3840 9313
rect 3894 9306 3898 9313
rect 3915 9310 3919 9314
rect 3932 9313 3936 9317
rect 3950 9315 3954 9319
rect 4010 9315 4014 9319
rect 3968 9306 3972 9313
rect 4026 9306 4030 9313
rect 4047 9310 4051 9314
rect 4064 9313 4068 9317
rect 4082 9315 4086 9319
rect 4142 9315 4146 9319
rect 4100 9306 4104 9313
rect 4158 9306 4162 9313
rect 4179 9310 4183 9314
rect 4196 9313 4200 9317
rect 4214 9315 4218 9319
rect 4274 9315 4278 9319
rect 4232 9306 4236 9313
rect 4290 9306 4294 9313
rect 4311 9310 4315 9314
rect 2861 9292 2865 9296
rect 2898 9290 2902 9294
rect 2918 9290 2922 9294
rect 2954 9290 2958 9294
rect 2993 9292 2997 9296
rect 3030 9290 3034 9294
rect 3050 9290 3054 9294
rect 3086 9290 3090 9294
rect 3125 9292 3129 9296
rect 3162 9290 3166 9294
rect 3182 9290 3186 9294
rect 3218 9290 3222 9294
rect 3257 9292 3261 9296
rect 3294 9290 3298 9294
rect 3314 9290 3318 9294
rect 3350 9290 3354 9294
rect 3806 9292 3810 9296
rect 3843 9290 3847 9294
rect 3863 9290 3867 9294
rect 3899 9290 3903 9294
rect 3938 9292 3942 9296
rect 3975 9290 3979 9294
rect 3995 9290 3999 9294
rect 4031 9290 4035 9294
rect 4070 9292 4074 9296
rect 4107 9290 4111 9294
rect 4127 9290 4131 9294
rect 4163 9290 4167 9294
rect 4202 9292 4206 9296
rect 4239 9290 4243 9294
rect 4259 9290 4263 9294
rect 4295 9290 4299 9294
rect 2503 9280 2507 9284
rect 2521 9282 2525 9286
rect 2581 9282 2585 9286
rect 2539 9273 2543 9280
rect 2597 9273 2601 9280
rect 2616 9277 2620 9281
rect 3448 9280 3452 9284
rect 3466 9282 3470 9286
rect 3526 9282 3530 9286
rect 3484 9273 3488 9280
rect 3542 9273 3546 9280
rect 3561 9277 3565 9281
rect 2509 9259 2513 9263
rect 2546 9257 2550 9261
rect 2566 9257 2570 9261
rect 2602 9257 2606 9261
rect 2877 9249 2881 9253
rect 2921 9249 2925 9253
rect 2948 9249 2952 9253
rect 2993 9249 2997 9253
rect 3066 9256 3070 9260
rect 2627 9236 2631 9240
rect 3031 9242 3035 9246
rect 2510 9227 2514 9231
rect 2857 9229 2861 9233
rect 2889 9230 2893 9234
rect 2908 9229 2912 9233
rect 2964 9230 2968 9234
rect 2980 9229 2984 9233
rect 3007 9229 3011 9233
rect 3147 9256 3151 9260
rect 3454 9259 3458 9263
rect 3058 9238 3062 9242
rect 3085 9234 3089 9238
rect 3112 9242 3116 9246
rect 3491 9257 3495 9261
rect 3511 9257 3515 9261
rect 3547 9257 3551 9261
rect 3139 9238 3143 9242
rect 3166 9234 3170 9238
rect 3822 9249 3826 9253
rect 3866 9249 3870 9253
rect 3893 9249 3897 9253
rect 3938 9249 3942 9253
rect 4011 9256 4015 9260
rect 3572 9236 3576 9240
rect 3976 9242 3980 9246
rect 3064 9220 3068 9224
rect 3455 9227 3459 9231
rect 3802 9229 3806 9233
rect 3145 9220 3149 9224
rect 3834 9230 3838 9234
rect 3853 9229 3857 9233
rect 3909 9230 3913 9234
rect 3925 9229 3929 9233
rect 3952 9229 3956 9233
rect 4092 9256 4096 9260
rect 4003 9238 4007 9242
rect 4030 9234 4034 9238
rect 4057 9242 4061 9246
rect 4084 9238 4088 9242
rect 4111 9234 4115 9238
rect 4009 9220 4013 9224
rect 4090 9220 4094 9224
rect 2874 9212 2878 9216
rect 2918 9211 2922 9215
rect 2943 9212 2948 9216
rect 2990 9211 2994 9215
rect 3819 9212 3823 9216
rect 3863 9211 3867 9215
rect 3888 9212 3893 9216
rect 3935 9211 3939 9215
rect 2509 9198 2513 9202
rect 2547 9198 2551 9202
rect 2567 9198 2571 9202
rect 2604 9198 2608 9202
rect 3454 9198 3458 9202
rect 3492 9198 3496 9202
rect 3512 9198 3516 9202
rect 3549 9198 3553 9202
rect 2497 9175 2501 9179
rect 2532 9180 2536 9184
rect 2516 9171 2520 9178
rect 2574 9171 2578 9178
rect 2592 9180 2596 9184
rect 2874 9182 2878 9186
rect 2918 9183 2922 9187
rect 2610 9178 2614 9182
rect 2943 9182 2948 9186
rect 2990 9183 2994 9187
rect 3066 9180 3070 9184
rect 3147 9180 3151 9184
rect 2857 9165 2861 9169
rect 2511 9155 2515 9159
rect 2547 9155 2551 9159
rect 2567 9155 2571 9159
rect 2604 9157 2608 9161
rect 2889 9164 2893 9168
rect 2908 9165 2912 9169
rect 2964 9164 2968 9168
rect 2980 9165 2984 9169
rect 3007 9165 3011 9169
rect 3055 9164 3061 9168
rect 3136 9164 3142 9168
rect 3442 9175 3446 9179
rect 3477 9180 3481 9184
rect 3461 9171 3465 9178
rect 3519 9171 3523 9178
rect 3537 9180 3541 9184
rect 3819 9182 3823 9186
rect 3863 9183 3867 9187
rect 3555 9178 3559 9182
rect 3888 9182 3893 9186
rect 3935 9183 3939 9187
rect 4011 9180 4015 9184
rect 4092 9180 4096 9184
rect 3802 9165 3806 9169
rect 3456 9155 3460 9159
rect 3492 9155 3496 9159
rect 3512 9155 3516 9159
rect 3549 9157 3553 9161
rect 3834 9164 3838 9168
rect 3853 9165 3857 9169
rect 3909 9164 3913 9168
rect 3925 9165 3929 9169
rect 3952 9165 3956 9169
rect 4000 9164 4006 9168
rect 4081 9164 4087 9168
rect 2877 9145 2881 9149
rect 2921 9145 2925 9149
rect 2948 9145 2952 9149
rect 2993 9145 2997 9149
rect 3064 9144 3068 9148
rect 3145 9144 3149 9148
rect 3822 9145 3826 9149
rect 3866 9145 3870 9149
rect 3893 9145 3897 9149
rect 3938 9145 3942 9149
rect 4009 9144 4013 9148
rect 4090 9144 4094 9148
rect 3066 9124 3070 9128
rect 2877 9117 2881 9121
rect 2921 9117 2925 9121
rect 2948 9117 2952 9121
rect 2993 9117 2997 9121
rect 3171 9124 3175 9128
rect 3058 9106 3062 9110
rect 2857 9097 2861 9101
rect 2889 9098 2893 9102
rect 2908 9097 2912 9101
rect 2964 9098 2968 9102
rect 2980 9097 2984 9101
rect 3007 9097 3011 9101
rect 3085 9102 3089 9106
rect 3136 9110 3140 9114
rect 4011 9124 4015 9128
rect 3163 9106 3167 9110
rect 3190 9102 3194 9106
rect 3822 9117 3826 9121
rect 3866 9117 3870 9121
rect 3893 9117 3897 9121
rect 3938 9117 3942 9121
rect 4116 9124 4120 9128
rect 4003 9106 4007 9110
rect 3064 9088 3068 9092
rect 3169 9088 3173 9092
rect 3402 9095 3406 9099
rect 2874 9080 2878 9084
rect 2918 9079 2922 9083
rect 2943 9080 2948 9084
rect 2990 9079 2994 9083
rect 3367 9081 3371 9085
rect 3802 9097 3806 9101
rect 3394 9077 3398 9081
rect 3421 9073 3425 9077
rect 3834 9098 3838 9102
rect 3853 9097 3857 9101
rect 3909 9098 3913 9102
rect 3925 9097 3929 9101
rect 3952 9097 3956 9101
rect 4030 9102 4034 9106
rect 4081 9110 4085 9114
rect 4108 9106 4112 9110
rect 4135 9102 4139 9106
rect 4009 9088 4013 9092
rect 4114 9088 4118 9092
rect 3819 9080 3823 9084
rect 3863 9079 3867 9083
rect 3888 9080 3893 9084
rect 3935 9079 3939 9083
rect 3400 9059 3404 9063
rect 2874 9050 2878 9054
rect 2918 9051 2922 9055
rect 2943 9050 2948 9054
rect 2990 9051 2994 9055
rect 3555 9053 3559 9057
rect 3608 9053 3612 9057
rect 3066 9049 3070 9053
rect 3171 9049 3175 9053
rect 3819 9050 3823 9054
rect 3863 9051 3867 9055
rect 3888 9050 3893 9054
rect 3935 9051 3939 9055
rect 4011 9049 4015 9053
rect 4116 9049 4120 9053
rect 2857 9033 2861 9037
rect 2889 9032 2893 9036
rect 2908 9033 2912 9037
rect 2964 9032 2968 9036
rect 2980 9033 2984 9037
rect 3007 9033 3011 9037
rect 3055 9033 3061 9037
rect 3160 9033 3166 9037
rect 3802 9033 3806 9037
rect 3834 9032 3838 9036
rect 3853 9033 3857 9037
rect 3909 9032 3913 9036
rect 3925 9033 3929 9037
rect 3952 9033 3956 9037
rect 4000 9033 4006 9037
rect 4105 9033 4111 9037
rect 2877 9013 2881 9017
rect 2921 9013 2925 9017
rect 2948 9013 2952 9017
rect 2993 9013 2997 9017
rect 3064 9013 3068 9017
rect 3169 9013 3173 9017
rect 3402 9015 3406 9019
rect 3822 9013 3826 9017
rect 3866 9013 3870 9017
rect 3893 9013 3897 9017
rect 3938 9013 3942 9017
rect 4009 9013 4013 9017
rect 4114 9013 4118 9017
rect 3391 8999 3397 9003
rect 3066 8992 3070 8996
rect 2877 8985 2881 8989
rect 2921 8985 2925 8989
rect 2948 8985 2952 8989
rect 2993 8985 2997 8989
rect 3147 8992 3151 8996
rect 3058 8974 3062 8978
rect 2857 8965 2861 8969
rect 2889 8966 2893 8970
rect 2908 8965 2912 8969
rect 2964 8966 2968 8970
rect 2980 8965 2984 8969
rect 3007 8965 3011 8969
rect 3085 8970 3089 8974
rect 3112 8978 3116 8982
rect 3237 8992 3241 8996
rect 3139 8974 3143 8978
rect 3166 8970 3170 8974
rect 3202 8978 3206 8982
rect 4011 8992 4015 8996
rect 3229 8974 3233 8978
rect 3256 8970 3260 8974
rect 3822 8985 3826 8989
rect 3866 8985 3870 8989
rect 3893 8985 3897 8989
rect 3938 8985 3942 8989
rect 3400 8979 3404 8983
rect 4092 8992 4096 8996
rect 4003 8974 4007 8978
rect 3064 8956 3068 8960
rect 3145 8956 3149 8960
rect 3235 8956 3239 8960
rect 3402 8965 3406 8969
rect 2874 8948 2878 8952
rect 2918 8947 2922 8951
rect 2943 8948 2948 8952
rect 3345 8951 3349 8955
rect 2990 8947 2994 8951
rect 3367 8951 3371 8955
rect 3802 8965 3806 8969
rect 3394 8947 3398 8951
rect 3421 8943 3425 8947
rect 3834 8966 3838 8970
rect 3853 8965 3857 8969
rect 3909 8966 3913 8970
rect 3925 8965 3929 8969
rect 3952 8965 3956 8969
rect 4030 8970 4034 8974
rect 4057 8978 4061 8982
rect 4182 8992 4186 8996
rect 4084 8974 4088 8978
rect 4111 8970 4115 8974
rect 4147 8978 4151 8982
rect 4174 8974 4178 8978
rect 4201 8970 4205 8974
rect 4009 8956 4013 8960
rect 4090 8956 4094 8960
rect 4180 8956 4184 8960
rect 3819 8948 3823 8952
rect 3863 8947 3867 8951
rect 3888 8948 3893 8952
rect 3935 8947 3939 8951
rect 3400 8929 3404 8933
rect 2874 8918 2878 8922
rect 2918 8919 2922 8923
rect 3461 8923 3465 8927
rect 3514 8923 3518 8927
rect 2943 8918 2948 8922
rect 2990 8919 2994 8923
rect 3066 8914 3070 8918
rect 3147 8914 3151 8918
rect 3237 8914 3241 8918
rect 3819 8918 3823 8922
rect 3863 8919 3867 8923
rect 2857 8901 2861 8905
rect 2889 8900 2893 8904
rect 2908 8901 2912 8905
rect 2964 8900 2968 8904
rect 2980 8901 2984 8905
rect 3007 8901 3011 8905
rect 3055 8898 3061 8902
rect 3136 8898 3142 8902
rect 3226 8898 3232 8902
rect 3888 8918 3893 8922
rect 3935 8919 3939 8923
rect 4011 8914 4015 8918
rect 4092 8914 4096 8918
rect 4182 8914 4186 8918
rect 3802 8901 3806 8905
rect 3834 8900 3838 8904
rect 3853 8901 3857 8905
rect 3909 8900 3913 8904
rect 3925 8901 3929 8905
rect 3952 8901 3956 8905
rect 4000 8898 4006 8902
rect 2877 8881 2881 8885
rect 2921 8881 2925 8885
rect 2948 8881 2952 8885
rect 2993 8881 2997 8885
rect 3402 8885 3406 8889
rect 4081 8898 4087 8902
rect 4171 8898 4177 8902
rect 3064 8878 3068 8882
rect 3145 8878 3149 8882
rect 3235 8878 3239 8882
rect 3822 8881 3826 8885
rect 3866 8881 3870 8885
rect 3893 8881 3897 8885
rect 3938 8881 3942 8885
rect 4009 8878 4013 8882
rect 4090 8878 4094 8882
rect 4180 8878 4184 8882
rect 3391 8869 3397 8873
rect 3066 8860 3070 8864
rect 2877 8853 2881 8857
rect 2921 8853 2925 8857
rect 2948 8853 2952 8857
rect 2993 8853 2997 8857
rect 3058 8842 3062 8846
rect 2857 8833 2861 8837
rect 2889 8834 2893 8838
rect 2908 8833 2912 8837
rect 2964 8834 2968 8838
rect 2980 8833 2984 8837
rect 3007 8833 3011 8837
rect 3085 8838 3089 8842
rect 3400 8849 3404 8853
rect 4011 8860 4015 8864
rect 3822 8853 3826 8857
rect 3866 8853 3870 8857
rect 3893 8853 3897 8857
rect 3938 8853 3942 8857
rect 4003 8842 4007 8846
rect 3802 8833 3806 8837
rect 3064 8824 3068 8828
rect 3834 8834 3838 8838
rect 3853 8833 3857 8837
rect 3909 8834 3913 8838
rect 3925 8833 3929 8837
rect 3952 8833 3956 8837
rect 4030 8838 4034 8842
rect 4009 8824 4013 8828
rect 2874 8816 2878 8820
rect 2918 8815 2922 8819
rect 2943 8816 2948 8820
rect 2990 8815 2994 8819
rect 3819 8816 3823 8820
rect 3863 8815 3867 8819
rect 3888 8816 3893 8820
rect 3935 8815 3939 8819
rect 2377 8798 2381 8802
rect 2414 8798 2418 8802
rect 2434 8798 2438 8802
rect 2472 8798 2476 8802
rect 2509 8798 2513 8802
rect 2546 8798 2550 8802
rect 2566 8798 2570 8802
rect 2604 8798 2608 8802
rect 2641 8798 2645 8802
rect 2678 8798 2682 8802
rect 2698 8798 2702 8802
rect 2736 8798 2740 8802
rect 3322 8798 3326 8802
rect 3359 8798 3363 8802
rect 3379 8798 3383 8802
rect 3417 8798 3421 8802
rect 3454 8798 3458 8802
rect 3491 8798 3495 8802
rect 3511 8798 3515 8802
rect 3549 8798 3553 8802
rect 3586 8798 3590 8802
rect 3623 8798 3627 8802
rect 3643 8798 3647 8802
rect 3681 8798 3685 8802
rect 2371 8778 2375 8782
rect 2389 8780 2393 8784
rect 2449 8780 2453 8784
rect 2407 8771 2411 8778
rect 2465 8771 2469 8778
rect 2484 8775 2488 8779
rect 2502 8780 2506 8784
rect 2521 8780 2525 8784
rect 2581 8780 2585 8784
rect 2539 8771 2543 8778
rect 2597 8771 2601 8778
rect 2616 8775 2620 8779
rect 2634 8780 2638 8784
rect 2653 8780 2657 8784
rect 2713 8780 2717 8784
rect 2671 8771 2675 8778
rect 2874 8786 2878 8790
rect 2918 8787 2922 8791
rect 2943 8786 2948 8790
rect 2990 8787 2994 8791
rect 3135 8786 3139 8790
rect 3179 8787 3183 8791
rect 3204 8786 3209 8790
rect 3251 8787 3255 8791
rect 2729 8771 2733 8778
rect 2750 8775 2754 8779
rect 3066 8778 3070 8782
rect 3316 8778 3320 8782
rect 3334 8780 3338 8784
rect 2857 8769 2861 8773
rect 2889 8768 2893 8772
rect 2908 8769 2912 8773
rect 2964 8768 2968 8772
rect 2980 8769 2984 8773
rect 3007 8769 3011 8773
rect 2377 8757 2381 8761
rect 2414 8755 2418 8759
rect 2434 8755 2438 8759
rect 2470 8755 2474 8759
rect 2509 8757 2513 8761
rect 2546 8755 2550 8759
rect 2566 8755 2570 8759
rect 2602 8755 2606 8759
rect 2641 8757 2645 8761
rect 2678 8755 2682 8759
rect 2698 8755 2702 8759
rect 2734 8755 2738 8759
rect 3055 8762 3061 8766
rect 3093 8769 3097 8773
rect 3150 8768 3154 8772
rect 3169 8769 3173 8773
rect 3225 8768 3229 8772
rect 3241 8769 3245 8773
rect 3268 8769 3272 8773
rect 3394 8780 3398 8784
rect 3352 8771 3356 8778
rect 3410 8771 3414 8778
rect 3429 8775 3433 8779
rect 3447 8780 3451 8784
rect 3466 8780 3470 8784
rect 3526 8780 3530 8784
rect 3484 8771 3488 8778
rect 3542 8771 3546 8778
rect 3561 8775 3565 8779
rect 3579 8780 3583 8784
rect 3598 8780 3602 8784
rect 3658 8780 3662 8784
rect 3616 8771 3620 8778
rect 3819 8786 3823 8790
rect 3863 8787 3867 8791
rect 3888 8786 3893 8790
rect 3935 8787 3939 8791
rect 4080 8786 4084 8790
rect 4124 8787 4128 8791
rect 4149 8786 4154 8790
rect 4196 8787 4200 8791
rect 3674 8771 3678 8778
rect 3695 8775 3699 8779
rect 4011 8778 4015 8782
rect 3802 8769 3806 8773
rect 3834 8768 3838 8772
rect 3853 8769 3857 8773
rect 3909 8768 3913 8772
rect 3925 8769 3929 8773
rect 3952 8769 3956 8773
rect 2877 8749 2881 8753
rect 2921 8749 2925 8753
rect 2948 8749 2952 8753
rect 2993 8749 2997 8753
rect 3322 8757 3326 8761
rect 3064 8742 3068 8746
rect 2486 8727 2490 8731
rect 2510 8727 2514 8731
rect 3359 8755 3363 8759
rect 3379 8755 3383 8759
rect 3415 8755 3419 8759
rect 3454 8757 3458 8761
rect 3491 8755 3495 8759
rect 3511 8755 3515 8759
rect 3547 8755 3551 8759
rect 3586 8757 3590 8761
rect 3623 8755 3627 8759
rect 3643 8755 3647 8759
rect 3679 8755 3683 8759
rect 4000 8762 4006 8766
rect 4038 8769 4042 8773
rect 4095 8768 4099 8772
rect 4114 8769 4118 8773
rect 4170 8768 4174 8772
rect 4186 8769 4190 8773
rect 4213 8769 4217 8773
rect 3138 8749 3142 8753
rect 3182 8749 3186 8753
rect 3209 8749 3213 8753
rect 3254 8749 3258 8753
rect 3822 8749 3826 8753
rect 3866 8749 3870 8753
rect 3893 8749 3897 8753
rect 3938 8749 3942 8753
rect 4009 8742 4013 8746
rect 3431 8727 3435 8731
rect 3455 8727 3459 8731
rect 3277 8721 3281 8725
rect 3115 8714 3119 8718
rect 4083 8749 4087 8753
rect 4127 8749 4131 8753
rect 4154 8749 4158 8753
rect 4199 8749 4203 8753
rect 4222 8721 4226 8725
rect 4058 8714 4062 8718
rect 2506 8700 2510 8704
rect 3451 8700 3455 8704
rect 2521 8692 2525 8696
rect 3466 8692 3470 8696
rect 3160 8686 3164 8690
rect 3197 8686 3201 8690
rect 3217 8686 3221 8690
rect 3255 8686 3259 8690
rect 4105 8686 4109 8690
rect 4142 8686 4146 8690
rect 4162 8686 4166 8690
rect 4200 8686 4204 8690
rect 2486 8677 2490 8681
rect 2510 8677 2514 8681
rect 3431 8677 3435 8681
rect 3455 8677 3459 8681
rect 3154 8666 3158 8670
rect 3172 8668 3176 8672
rect 2377 8656 2381 8660
rect 2414 8656 2418 8660
rect 2434 8656 2438 8660
rect 2472 8656 2476 8660
rect 2509 8656 2513 8660
rect 2546 8656 2550 8660
rect 2566 8656 2570 8660
rect 2604 8656 2608 8660
rect 2641 8656 2645 8660
rect 2678 8656 2682 8660
rect 2698 8656 2702 8660
rect 2736 8656 2740 8660
rect 3232 8668 3236 8672
rect 3190 8659 3194 8666
rect 3248 8659 3252 8666
rect 3267 8663 3271 8667
rect 4099 8666 4103 8670
rect 4117 8668 4121 8672
rect 3322 8656 3326 8660
rect 3359 8656 3363 8660
rect 3379 8656 3383 8660
rect 3417 8656 3421 8660
rect 3454 8656 3458 8660
rect 3491 8656 3495 8660
rect 3511 8656 3515 8660
rect 3549 8656 3553 8660
rect 3586 8656 3590 8660
rect 3623 8656 3627 8660
rect 3643 8656 3647 8660
rect 3681 8656 3685 8660
rect 4177 8668 4181 8672
rect 4135 8659 4139 8666
rect 4193 8659 4197 8666
rect 4212 8663 4216 8667
rect 3160 8645 3164 8649
rect 2371 8636 2375 8640
rect 2389 8638 2393 8642
rect 2449 8638 2453 8642
rect 2407 8629 2411 8636
rect 2465 8629 2469 8636
rect 2484 8633 2488 8637
rect 2502 8638 2506 8642
rect 2521 8638 2525 8642
rect 2581 8638 2585 8642
rect 2539 8629 2543 8636
rect 2597 8629 2601 8636
rect 2616 8633 2620 8637
rect 2634 8638 2638 8642
rect 2653 8638 2657 8642
rect 2713 8638 2717 8642
rect 2671 8629 2675 8636
rect 3197 8643 3201 8647
rect 3217 8643 3221 8647
rect 3253 8643 3257 8647
rect 4105 8645 4109 8649
rect 2729 8629 2733 8636
rect 2750 8633 2754 8637
rect 3316 8636 3320 8640
rect 3334 8638 3338 8642
rect 3394 8638 3398 8642
rect 3352 8629 3356 8636
rect 3410 8629 3414 8636
rect 3429 8633 3433 8637
rect 3447 8638 3451 8642
rect 3466 8638 3470 8642
rect 3526 8638 3530 8642
rect 3484 8629 3488 8636
rect 3542 8629 3546 8636
rect 3561 8633 3565 8637
rect 3579 8638 3583 8642
rect 3598 8638 3602 8642
rect 3658 8638 3662 8642
rect 3616 8629 3620 8636
rect 4142 8643 4146 8647
rect 4162 8643 4166 8647
rect 4198 8643 4202 8647
rect 3674 8629 3678 8636
rect 3695 8633 3699 8637
rect 2377 8615 2381 8619
rect 2414 8613 2418 8617
rect 2434 8613 2438 8617
rect 2470 8613 2474 8617
rect 2509 8615 2513 8619
rect 2546 8613 2550 8617
rect 2566 8613 2570 8617
rect 2602 8613 2606 8617
rect 2641 8615 2645 8619
rect 2678 8613 2682 8617
rect 2698 8613 2702 8617
rect 2734 8613 2738 8617
rect 3322 8615 3326 8619
rect 3359 8613 3363 8617
rect 3379 8613 3383 8617
rect 3415 8613 3419 8617
rect 3454 8615 3458 8619
rect 3491 8613 3495 8617
rect 3511 8613 3515 8617
rect 3547 8613 3551 8617
rect 3586 8615 3590 8619
rect 3623 8613 3627 8617
rect 3643 8613 3647 8617
rect 3679 8613 3683 8617
rect 3160 8600 3164 8604
rect 3197 8600 3201 8604
rect 3217 8600 3221 8604
rect 3255 8600 3259 8604
rect 4105 8600 4109 8604
rect 4142 8600 4146 8604
rect 4162 8600 4166 8604
rect 4200 8600 4204 8604
rect 3154 8580 3158 8584
rect 3172 8582 3176 8586
rect 2377 8570 2381 8574
rect 2414 8570 2418 8574
rect 2434 8570 2438 8574
rect 2472 8570 2476 8574
rect 2509 8570 2513 8574
rect 2546 8570 2550 8574
rect 2566 8570 2570 8574
rect 2604 8570 2608 8574
rect 2641 8570 2645 8574
rect 2678 8570 2682 8574
rect 2698 8570 2702 8574
rect 2736 8570 2740 8574
rect 3232 8582 3236 8586
rect 3190 8573 3194 8580
rect 3248 8573 3252 8580
rect 3267 8577 3271 8581
rect 3289 8575 3293 8579
rect 4099 8580 4103 8584
rect 4117 8582 4121 8586
rect 3322 8570 3326 8574
rect 3359 8570 3363 8574
rect 3379 8570 3383 8574
rect 3417 8570 3421 8574
rect 3454 8570 3458 8574
rect 3491 8570 3495 8574
rect 3511 8570 3515 8574
rect 3549 8570 3553 8574
rect 3586 8570 3590 8574
rect 3623 8570 3627 8574
rect 3643 8570 3647 8574
rect 3681 8570 3685 8574
rect 4177 8582 4181 8586
rect 4135 8573 4139 8580
rect 4193 8573 4197 8580
rect 4212 8577 4216 8581
rect 4234 8575 4238 8579
rect 3160 8559 3164 8563
rect 2371 8550 2375 8554
rect 2389 8552 2393 8556
rect 2449 8552 2453 8556
rect 2407 8543 2411 8550
rect 2465 8543 2469 8550
rect 2484 8547 2488 8551
rect 2502 8552 2506 8556
rect 2521 8552 2525 8556
rect 2581 8552 2585 8556
rect 2539 8543 2543 8550
rect 2597 8543 2601 8550
rect 2616 8547 2620 8551
rect 2634 8552 2638 8556
rect 2653 8552 2657 8556
rect 2713 8552 2717 8556
rect 2671 8543 2675 8550
rect 3197 8557 3201 8561
rect 3217 8557 3221 8561
rect 3253 8557 3257 8561
rect 4105 8559 4109 8563
rect 2729 8543 2733 8550
rect 2750 8547 2754 8551
rect 3316 8550 3320 8554
rect 3334 8552 3338 8556
rect 3394 8552 3398 8556
rect 3352 8543 3356 8550
rect 3410 8543 3414 8550
rect 3429 8547 3433 8551
rect 3447 8552 3451 8556
rect 3466 8552 3470 8556
rect 3526 8552 3530 8556
rect 3484 8543 3488 8550
rect 3542 8543 3546 8550
rect 3561 8547 3565 8551
rect 3579 8552 3583 8556
rect 3598 8552 3602 8556
rect 3658 8552 3662 8556
rect 3616 8543 3620 8550
rect 4142 8557 4146 8561
rect 4162 8557 4166 8561
rect 4198 8557 4202 8561
rect 3674 8543 3678 8550
rect 3695 8547 3699 8551
rect 2377 8529 2381 8533
rect 2414 8527 2418 8531
rect 2434 8527 2438 8531
rect 2470 8527 2474 8531
rect 2509 8529 2513 8533
rect 2546 8527 2550 8531
rect 2566 8527 2570 8531
rect 2602 8527 2606 8531
rect 2641 8529 2645 8533
rect 2678 8527 2682 8531
rect 2698 8527 2702 8531
rect 2734 8527 2738 8531
rect 3322 8529 3326 8533
rect 3359 8527 3363 8531
rect 3379 8527 3383 8531
rect 3415 8527 3419 8531
rect 3454 8529 3458 8533
rect 3491 8527 3495 8531
rect 3511 8527 3515 8531
rect 3547 8527 3551 8531
rect 3586 8529 3590 8533
rect 3623 8527 3627 8531
rect 3643 8527 3647 8531
rect 3679 8527 3683 8531
rect 2603 8499 2607 8503
rect 2627 8499 2631 8503
rect 3548 8499 3552 8503
rect 3572 8499 3576 8503
rect 2623 8474 2627 8478
rect 3568 8474 3572 8478
rect 2638 8466 2642 8470
rect 3583 8466 3587 8470
rect 2603 8451 2607 8455
rect 2627 8451 2631 8455
rect 3548 8451 3552 8455
rect 3572 8451 3576 8455
rect 2377 8430 2381 8434
rect 2414 8430 2418 8434
rect 2434 8430 2438 8434
rect 2472 8430 2476 8434
rect 2509 8430 2513 8434
rect 2546 8430 2550 8434
rect 2566 8430 2570 8434
rect 2604 8430 2608 8434
rect 2641 8430 2645 8434
rect 2678 8430 2682 8434
rect 2698 8430 2702 8434
rect 2736 8430 2740 8434
rect 3322 8430 3326 8434
rect 3359 8430 3363 8434
rect 3379 8430 3383 8434
rect 3417 8430 3421 8434
rect 3454 8430 3458 8434
rect 3491 8430 3495 8434
rect 3511 8430 3515 8434
rect 3549 8430 3553 8434
rect 3586 8430 3590 8434
rect 3623 8430 3627 8434
rect 3643 8430 3647 8434
rect 3681 8430 3685 8434
rect 2371 8410 2375 8414
rect 2389 8412 2393 8416
rect 2449 8412 2453 8416
rect 2407 8403 2411 8410
rect 2465 8403 2469 8410
rect 2484 8407 2488 8411
rect 2502 8412 2506 8416
rect 2521 8412 2525 8416
rect 2581 8412 2585 8416
rect 2539 8403 2543 8410
rect 2597 8403 2601 8410
rect 2616 8407 2620 8411
rect 2634 8412 2638 8416
rect 2653 8412 2657 8416
rect 2713 8412 2717 8416
rect 2671 8403 2675 8410
rect 2729 8403 2733 8410
rect 2750 8407 2754 8411
rect 3316 8410 3320 8414
rect 3334 8412 3338 8416
rect 3394 8412 3398 8416
rect 3352 8403 3356 8410
rect 3410 8403 3414 8410
rect 3429 8407 3433 8411
rect 3447 8412 3451 8416
rect 3466 8412 3470 8416
rect 3526 8412 3530 8416
rect 3484 8403 3488 8410
rect 3542 8403 3546 8410
rect 3561 8407 3565 8411
rect 3579 8412 3583 8416
rect 3598 8412 3602 8416
rect 3658 8412 3662 8416
rect 3616 8403 3620 8410
rect 3674 8403 3678 8410
rect 3695 8407 3699 8411
rect 2377 8389 2381 8393
rect 2414 8387 2418 8391
rect 2434 8387 2438 8391
rect 2470 8387 2474 8391
rect 2509 8389 2513 8393
rect 2546 8387 2550 8391
rect 2566 8387 2570 8391
rect 2602 8387 2606 8391
rect 2641 8389 2645 8393
rect 2678 8387 2682 8391
rect 2698 8387 2702 8391
rect 2734 8387 2738 8391
rect 3322 8389 3326 8393
rect 3359 8387 3363 8391
rect 3379 8387 3383 8391
rect 3415 8387 3419 8391
rect 3454 8389 3458 8393
rect 3491 8387 3495 8391
rect 3511 8387 3515 8391
rect 3547 8387 3551 8391
rect 3586 8389 3590 8393
rect 3623 8387 3627 8391
rect 3643 8387 3647 8391
rect 3679 8387 3683 8391
rect 2861 8351 2865 8355
rect 2898 8351 2902 8355
rect 2918 8351 2922 8355
rect 2956 8351 2960 8355
rect 2993 8351 2997 8355
rect 3030 8351 3034 8355
rect 3050 8351 3054 8355
rect 3088 8351 3092 8355
rect 3125 8351 3129 8355
rect 3162 8351 3166 8355
rect 3182 8351 3186 8355
rect 3220 8351 3224 8355
rect 3257 8351 3261 8355
rect 3294 8351 3298 8355
rect 3314 8351 3318 8355
rect 3352 8351 3356 8355
rect 3806 8351 3810 8355
rect 3843 8351 3847 8355
rect 3863 8351 3867 8355
rect 3901 8351 3905 8355
rect 3938 8351 3942 8355
rect 3975 8351 3979 8355
rect 3995 8351 3999 8355
rect 4033 8351 4037 8355
rect 4070 8351 4074 8355
rect 4107 8351 4111 8355
rect 4127 8351 4131 8355
rect 4165 8351 4169 8355
rect 4202 8351 4206 8355
rect 4239 8351 4243 8355
rect 4259 8351 4263 8355
rect 4297 8351 4301 8355
rect 2855 8331 2859 8335
rect 2873 8333 2877 8337
rect 2509 8318 2513 8322
rect 2546 8318 2550 8322
rect 2566 8318 2570 8322
rect 2604 8318 2608 8322
rect 2933 8333 2937 8337
rect 2891 8324 2895 8331
rect 2949 8324 2953 8331
rect 2970 8328 2974 8332
rect 2987 8331 2991 8335
rect 3005 8333 3009 8337
rect 3065 8333 3069 8337
rect 3023 8324 3027 8331
rect 3081 8324 3085 8331
rect 3102 8328 3106 8332
rect 3119 8331 3123 8335
rect 3137 8333 3141 8337
rect 3197 8333 3201 8337
rect 3155 8324 3159 8331
rect 3213 8324 3217 8331
rect 3234 8328 3238 8332
rect 3251 8331 3255 8335
rect 3269 8333 3273 8337
rect 3329 8333 3333 8337
rect 3287 8324 3291 8331
rect 3345 8324 3349 8331
rect 3366 8328 3370 8332
rect 3800 8331 3804 8335
rect 3818 8333 3822 8337
rect 3454 8318 3458 8322
rect 3491 8318 3495 8322
rect 3511 8318 3515 8322
rect 3549 8318 3553 8322
rect 3878 8333 3882 8337
rect 3836 8324 3840 8331
rect 3894 8324 3898 8331
rect 3915 8328 3919 8332
rect 3932 8331 3936 8335
rect 3950 8333 3954 8337
rect 4010 8333 4014 8337
rect 3968 8324 3972 8331
rect 4026 8324 4030 8331
rect 4047 8328 4051 8332
rect 4064 8331 4068 8335
rect 4082 8333 4086 8337
rect 4142 8333 4146 8337
rect 4100 8324 4104 8331
rect 4158 8324 4162 8331
rect 4179 8328 4183 8332
rect 4196 8331 4200 8335
rect 4214 8333 4218 8337
rect 4274 8333 4278 8337
rect 4232 8324 4236 8331
rect 4290 8324 4294 8331
rect 4311 8328 4315 8332
rect 2861 8310 2865 8314
rect 2898 8308 2902 8312
rect 2918 8308 2922 8312
rect 2954 8308 2958 8312
rect 2993 8310 2997 8314
rect 3030 8308 3034 8312
rect 3050 8308 3054 8312
rect 3086 8308 3090 8312
rect 3125 8310 3129 8314
rect 3162 8308 3166 8312
rect 3182 8308 3186 8312
rect 3218 8308 3222 8312
rect 3257 8310 3261 8314
rect 3294 8308 3298 8312
rect 3314 8308 3318 8312
rect 3350 8308 3354 8312
rect 3806 8310 3810 8314
rect 3843 8308 3847 8312
rect 3863 8308 3867 8312
rect 3899 8308 3903 8312
rect 3938 8310 3942 8314
rect 3975 8308 3979 8312
rect 3995 8308 3999 8312
rect 4031 8308 4035 8312
rect 4070 8310 4074 8314
rect 4107 8308 4111 8312
rect 4127 8308 4131 8312
rect 4163 8308 4167 8312
rect 4202 8310 4206 8314
rect 4239 8308 4243 8312
rect 4259 8308 4263 8312
rect 4295 8308 4299 8312
rect 2503 8298 2507 8302
rect 2521 8300 2525 8304
rect 2581 8300 2585 8304
rect 2539 8291 2543 8298
rect 2597 8291 2601 8298
rect 2616 8295 2620 8299
rect 3448 8298 3452 8302
rect 3466 8300 3470 8304
rect 3526 8300 3530 8304
rect 3484 8291 3488 8298
rect 3542 8291 3546 8298
rect 3561 8295 3565 8299
rect 2509 8277 2513 8281
rect 2546 8275 2550 8279
rect 2566 8275 2570 8279
rect 2602 8275 2606 8279
rect 2877 8267 2881 8271
rect 2921 8267 2925 8271
rect 2948 8267 2952 8271
rect 2993 8267 2997 8271
rect 3066 8274 3070 8278
rect 2627 8254 2631 8258
rect 3031 8260 3035 8264
rect 2510 8245 2514 8249
rect 2857 8247 2861 8251
rect 2889 8248 2893 8252
rect 2908 8247 2912 8251
rect 2964 8248 2968 8252
rect 2980 8247 2984 8251
rect 3007 8247 3011 8251
rect 3147 8274 3151 8278
rect 3454 8277 3458 8281
rect 3058 8256 3062 8260
rect 3085 8252 3089 8256
rect 3112 8260 3116 8264
rect 3491 8275 3495 8279
rect 3511 8275 3515 8279
rect 3547 8275 3551 8279
rect 3139 8256 3143 8260
rect 3166 8252 3170 8256
rect 3822 8267 3826 8271
rect 3866 8267 3870 8271
rect 3893 8267 3897 8271
rect 3938 8267 3942 8271
rect 4011 8274 4015 8278
rect 3572 8254 3576 8258
rect 3976 8260 3980 8264
rect 3064 8238 3068 8242
rect 3455 8245 3459 8249
rect 3802 8247 3806 8251
rect 3145 8238 3149 8242
rect 3834 8248 3838 8252
rect 3853 8247 3857 8251
rect 3909 8248 3913 8252
rect 3925 8247 3929 8251
rect 3952 8247 3956 8251
rect 4092 8274 4096 8278
rect 4003 8256 4007 8260
rect 4030 8252 4034 8256
rect 4057 8260 4061 8264
rect 4084 8256 4088 8260
rect 4111 8252 4115 8256
rect 4009 8238 4013 8242
rect 4090 8238 4094 8242
rect 2874 8230 2878 8234
rect 2918 8229 2922 8233
rect 2943 8230 2948 8234
rect 2990 8229 2994 8233
rect 3819 8230 3823 8234
rect 3863 8229 3867 8233
rect 3888 8230 3893 8234
rect 3935 8229 3939 8233
rect 2509 8216 2513 8220
rect 2547 8216 2551 8220
rect 2567 8216 2571 8220
rect 2604 8216 2608 8220
rect 3454 8216 3458 8220
rect 3492 8216 3496 8220
rect 3512 8216 3516 8220
rect 3549 8216 3553 8220
rect 2497 8193 2501 8197
rect 2532 8198 2536 8202
rect 2516 8189 2520 8196
rect 2574 8189 2578 8196
rect 2592 8198 2596 8202
rect 2874 8200 2878 8204
rect 2918 8201 2922 8205
rect 2610 8196 2614 8200
rect 2943 8200 2948 8204
rect 2990 8201 2994 8205
rect 3066 8198 3070 8202
rect 3147 8198 3151 8202
rect 2857 8183 2861 8187
rect 2511 8173 2515 8177
rect 2547 8173 2551 8177
rect 2567 8173 2571 8177
rect 2604 8175 2608 8179
rect 2889 8182 2893 8186
rect 2908 8183 2912 8187
rect 2964 8182 2968 8186
rect 2980 8183 2984 8187
rect 3007 8183 3011 8187
rect 3055 8182 3061 8186
rect 3136 8182 3142 8186
rect 3442 8193 3446 8197
rect 3477 8198 3481 8202
rect 3461 8189 3465 8196
rect 3519 8189 3523 8196
rect 3537 8198 3541 8202
rect 3819 8200 3823 8204
rect 3863 8201 3867 8205
rect 3555 8196 3559 8200
rect 3888 8200 3893 8204
rect 3935 8201 3939 8205
rect 4011 8198 4015 8202
rect 4092 8198 4096 8202
rect 3802 8183 3806 8187
rect 3456 8173 3460 8177
rect 3492 8173 3496 8177
rect 3512 8173 3516 8177
rect 3549 8175 3553 8179
rect 3834 8182 3838 8186
rect 3853 8183 3857 8187
rect 3909 8182 3913 8186
rect 3925 8183 3929 8187
rect 3952 8183 3956 8187
rect 4000 8182 4006 8186
rect 4081 8182 4087 8186
rect 2877 8163 2881 8167
rect 2921 8163 2925 8167
rect 2948 8163 2952 8167
rect 2993 8163 2997 8167
rect 3064 8162 3068 8166
rect 3145 8162 3149 8166
rect 3822 8163 3826 8167
rect 3866 8163 3870 8167
rect 3893 8163 3897 8167
rect 3938 8163 3942 8167
rect 4009 8162 4013 8166
rect 4090 8162 4094 8166
rect 3066 8142 3070 8146
rect 2877 8135 2881 8139
rect 2921 8135 2925 8139
rect 2948 8135 2952 8139
rect 2993 8135 2997 8139
rect 3171 8142 3175 8146
rect 3058 8124 3062 8128
rect 2857 8115 2861 8119
rect 2889 8116 2893 8120
rect 2908 8115 2912 8119
rect 2964 8116 2968 8120
rect 2980 8115 2984 8119
rect 3007 8115 3011 8119
rect 3085 8120 3089 8124
rect 3136 8128 3140 8132
rect 4011 8142 4015 8146
rect 3163 8124 3167 8128
rect 3190 8120 3194 8124
rect 3822 8135 3826 8139
rect 3866 8135 3870 8139
rect 3893 8135 3897 8139
rect 3938 8135 3942 8139
rect 4116 8142 4120 8146
rect 4003 8124 4007 8128
rect 3802 8115 3806 8119
rect 3064 8106 3068 8110
rect 3169 8106 3173 8110
rect 3834 8116 3838 8120
rect 3853 8115 3857 8119
rect 3909 8116 3913 8120
rect 3925 8115 3929 8119
rect 3952 8115 3956 8119
rect 4030 8120 4034 8124
rect 4081 8128 4085 8132
rect 4108 8124 4112 8128
rect 4135 8120 4139 8124
rect 4009 8106 4013 8110
rect 4114 8106 4118 8110
rect 2874 8098 2878 8102
rect 2918 8097 2922 8101
rect 2943 8098 2948 8102
rect 2990 8097 2994 8101
rect 3819 8098 3823 8102
rect 3863 8097 3867 8101
rect 3888 8098 3893 8102
rect 3935 8097 3939 8101
rect 2874 8068 2878 8072
rect 2918 8069 2922 8073
rect 2943 8068 2948 8072
rect 2990 8069 2994 8073
rect 3066 8067 3070 8071
rect 3171 8067 3175 8071
rect 3819 8068 3823 8072
rect 3863 8069 3867 8073
rect 3888 8068 3893 8072
rect 3935 8069 3939 8073
rect 4011 8067 4015 8071
rect 4116 8067 4120 8071
rect 2857 8051 2861 8055
rect 2889 8050 2893 8054
rect 2908 8051 2912 8055
rect 2964 8050 2968 8054
rect 2980 8051 2984 8055
rect 3007 8051 3011 8055
rect 3055 8051 3061 8055
rect 3160 8051 3166 8055
rect 3802 8051 3806 8055
rect 3834 8050 3838 8054
rect 3853 8051 3857 8055
rect 3909 8050 3913 8054
rect 3925 8051 3929 8055
rect 3952 8051 3956 8055
rect 4000 8051 4006 8055
rect 4105 8051 4111 8055
rect 2877 8031 2881 8035
rect 2921 8031 2925 8035
rect 2948 8031 2952 8035
rect 2993 8031 2997 8035
rect 3064 8031 3068 8035
rect 3169 8031 3173 8035
rect 3822 8031 3826 8035
rect 3866 8031 3870 8035
rect 3893 8031 3897 8035
rect 3938 8031 3942 8035
rect 4009 8031 4013 8035
rect 4114 8031 4118 8035
rect 3066 8010 3070 8014
rect 2877 8003 2881 8007
rect 2921 8003 2925 8007
rect 2948 8003 2952 8007
rect 2993 8003 2997 8007
rect 3147 8010 3151 8014
rect 3058 7992 3062 7996
rect 2857 7983 2861 7987
rect 2889 7984 2893 7988
rect 2908 7983 2912 7987
rect 2964 7984 2968 7988
rect 2980 7983 2984 7987
rect 3007 7983 3011 7987
rect 3085 7988 3089 7992
rect 3112 7996 3116 8000
rect 3237 8010 3241 8014
rect 3139 7992 3143 7996
rect 3166 7988 3170 7992
rect 3202 7996 3206 8000
rect 4011 8010 4015 8014
rect 3229 7992 3233 7996
rect 3256 7988 3260 7992
rect 3822 8003 3826 8007
rect 3866 8003 3870 8007
rect 3893 8003 3897 8007
rect 3938 8003 3942 8007
rect 4092 8010 4096 8014
rect 4003 7992 4007 7996
rect 3802 7983 3806 7987
rect 3064 7974 3068 7978
rect 3145 7974 3149 7978
rect 3235 7974 3239 7978
rect 3834 7984 3838 7988
rect 3853 7983 3857 7987
rect 3909 7984 3913 7988
rect 3925 7983 3929 7987
rect 3952 7983 3956 7987
rect 4030 7988 4034 7992
rect 4057 7996 4061 8000
rect 4182 8010 4186 8014
rect 4084 7992 4088 7996
rect 4111 7988 4115 7992
rect 4147 7996 4151 8000
rect 4174 7992 4178 7996
rect 4201 7988 4205 7992
rect 4009 7974 4013 7978
rect 4090 7974 4094 7978
rect 4180 7974 4184 7978
rect 2874 7966 2878 7970
rect 2918 7965 2922 7969
rect 2943 7966 2948 7970
rect 2990 7965 2994 7969
rect 3819 7966 3823 7970
rect 3863 7965 3867 7969
rect 3888 7966 3893 7970
rect 3935 7965 3939 7969
rect 2874 7936 2878 7940
rect 2918 7937 2922 7941
rect 2943 7936 2948 7940
rect 2990 7937 2994 7941
rect 3819 7936 3823 7940
rect 3863 7937 3867 7941
rect 3066 7932 3070 7936
rect 3147 7932 3151 7936
rect 3237 7932 3241 7936
rect 3888 7936 3893 7940
rect 3935 7937 3939 7941
rect 4011 7932 4015 7936
rect 4092 7932 4096 7936
rect 4182 7932 4186 7936
rect 2857 7919 2861 7923
rect 2889 7918 2893 7922
rect 2908 7919 2912 7923
rect 2964 7918 2968 7922
rect 2980 7919 2984 7923
rect 3007 7919 3011 7923
rect 3055 7916 3061 7920
rect 3136 7916 3142 7920
rect 3226 7916 3232 7920
rect 3802 7919 3806 7923
rect 3834 7918 3838 7922
rect 3853 7919 3857 7923
rect 3909 7918 3913 7922
rect 3925 7919 3929 7923
rect 3952 7919 3956 7923
rect 4000 7916 4006 7920
rect 4081 7916 4087 7920
rect 4171 7916 4177 7920
rect 2877 7899 2881 7903
rect 2921 7899 2925 7903
rect 2948 7899 2952 7903
rect 2993 7899 2997 7903
rect 3064 7896 3068 7900
rect 3145 7896 3149 7900
rect 3235 7896 3239 7900
rect 3822 7899 3826 7903
rect 3866 7899 3870 7903
rect 3893 7899 3897 7903
rect 3938 7899 3942 7903
rect 4009 7896 4013 7900
rect 4090 7896 4094 7900
rect 4180 7896 4184 7900
rect 3066 7878 3070 7882
rect 2877 7871 2881 7875
rect 2921 7871 2925 7875
rect 2948 7871 2952 7875
rect 2993 7871 2997 7875
rect 4011 7878 4015 7882
rect 3058 7860 3062 7864
rect 2857 7851 2861 7855
rect 2889 7852 2893 7856
rect 2908 7851 2912 7855
rect 2964 7852 2968 7856
rect 2980 7851 2984 7855
rect 3007 7851 3011 7855
rect 3085 7856 3089 7860
rect 3822 7871 3826 7875
rect 3866 7871 3870 7875
rect 3893 7871 3897 7875
rect 3938 7871 3942 7875
rect 4003 7860 4007 7864
rect 3802 7851 3806 7855
rect 3064 7842 3068 7846
rect 3834 7852 3838 7856
rect 3853 7851 3857 7855
rect 3909 7852 3913 7856
rect 3925 7851 3929 7855
rect 3952 7851 3956 7855
rect 4030 7856 4034 7860
rect 4009 7842 4013 7846
rect 2874 7834 2878 7838
rect 2918 7833 2922 7837
rect 2943 7834 2948 7838
rect 2990 7833 2994 7837
rect 3819 7834 3823 7838
rect 3863 7833 3867 7837
rect 3888 7834 3893 7838
rect 3935 7833 3939 7837
rect 2377 7816 2381 7820
rect 2414 7816 2418 7820
rect 2434 7816 2438 7820
rect 2472 7816 2476 7820
rect 2509 7816 2513 7820
rect 2546 7816 2550 7820
rect 2566 7816 2570 7820
rect 2604 7816 2608 7820
rect 2641 7816 2645 7820
rect 2678 7816 2682 7820
rect 2698 7816 2702 7820
rect 2736 7816 2740 7820
rect 3322 7816 3326 7820
rect 3359 7816 3363 7820
rect 3379 7816 3383 7820
rect 3417 7816 3421 7820
rect 3454 7816 3458 7820
rect 3491 7816 3495 7820
rect 3511 7816 3515 7820
rect 3549 7816 3553 7820
rect 3586 7816 3590 7820
rect 3623 7816 3627 7820
rect 3643 7816 3647 7820
rect 3681 7816 3685 7820
rect 2371 7796 2375 7800
rect 2389 7798 2393 7802
rect 2449 7798 2453 7802
rect 2407 7789 2411 7796
rect 2465 7789 2469 7796
rect 2484 7793 2488 7797
rect 2502 7798 2506 7802
rect 2521 7798 2525 7802
rect 2581 7798 2585 7802
rect 2539 7789 2543 7796
rect 2597 7789 2601 7796
rect 2616 7793 2620 7797
rect 2634 7798 2638 7802
rect 2653 7798 2657 7802
rect 2713 7798 2717 7802
rect 2671 7789 2675 7796
rect 2874 7804 2878 7808
rect 2918 7805 2922 7809
rect 2943 7804 2948 7808
rect 2990 7805 2994 7809
rect 3135 7804 3139 7808
rect 3179 7805 3183 7809
rect 3204 7804 3209 7808
rect 3251 7805 3255 7809
rect 2729 7789 2733 7796
rect 2750 7793 2754 7797
rect 3066 7796 3070 7800
rect 3316 7796 3320 7800
rect 3334 7798 3338 7802
rect 2857 7787 2861 7791
rect 2889 7786 2893 7790
rect 2908 7787 2912 7791
rect 2964 7786 2968 7790
rect 2980 7787 2984 7791
rect 3007 7787 3011 7791
rect 2377 7775 2381 7779
rect 2414 7773 2418 7777
rect 2434 7773 2438 7777
rect 2470 7773 2474 7777
rect 2509 7775 2513 7779
rect 2546 7773 2550 7777
rect 2566 7773 2570 7777
rect 2602 7773 2606 7777
rect 2641 7775 2645 7779
rect 2678 7773 2682 7777
rect 2698 7773 2702 7777
rect 2734 7773 2738 7777
rect 3055 7780 3061 7784
rect 3093 7787 3097 7791
rect 3150 7786 3154 7790
rect 3169 7787 3173 7791
rect 3225 7786 3229 7790
rect 3241 7787 3245 7791
rect 3268 7787 3272 7791
rect 3394 7798 3398 7802
rect 3352 7789 3356 7796
rect 3410 7789 3414 7796
rect 3429 7793 3433 7797
rect 3447 7798 3451 7802
rect 3466 7798 3470 7802
rect 3526 7798 3530 7802
rect 3484 7789 3488 7796
rect 3542 7789 3546 7796
rect 3561 7793 3565 7797
rect 3579 7798 3583 7802
rect 3598 7798 3602 7802
rect 3658 7798 3662 7802
rect 3616 7789 3620 7796
rect 3819 7804 3823 7808
rect 3863 7805 3867 7809
rect 3888 7804 3893 7808
rect 3935 7805 3939 7809
rect 4080 7804 4084 7808
rect 4124 7805 4128 7809
rect 4149 7804 4154 7808
rect 4196 7805 4200 7809
rect 3674 7789 3678 7796
rect 3695 7793 3699 7797
rect 4011 7796 4015 7800
rect 3802 7787 3806 7791
rect 3834 7786 3838 7790
rect 3853 7787 3857 7791
rect 3909 7786 3913 7790
rect 3925 7787 3929 7791
rect 3952 7787 3956 7791
rect 2877 7767 2881 7771
rect 2921 7767 2925 7771
rect 2948 7767 2952 7771
rect 2993 7767 2997 7771
rect 3322 7775 3326 7779
rect 3064 7760 3068 7764
rect 2486 7745 2490 7749
rect 2510 7745 2514 7749
rect 3359 7773 3363 7777
rect 3379 7773 3383 7777
rect 3415 7773 3419 7777
rect 3454 7775 3458 7779
rect 3491 7773 3495 7777
rect 3511 7773 3515 7777
rect 3547 7773 3551 7777
rect 3586 7775 3590 7779
rect 3623 7773 3627 7777
rect 3643 7773 3647 7777
rect 3679 7773 3683 7777
rect 4000 7780 4006 7784
rect 4038 7787 4042 7791
rect 4095 7786 4099 7790
rect 4114 7787 4118 7791
rect 4170 7786 4174 7790
rect 4186 7787 4190 7791
rect 4213 7787 4217 7791
rect 3138 7767 3142 7771
rect 3182 7767 3186 7771
rect 3209 7767 3213 7771
rect 3254 7767 3258 7771
rect 3822 7767 3826 7771
rect 3866 7767 3870 7771
rect 3893 7767 3897 7771
rect 3938 7767 3942 7771
rect 4009 7760 4013 7764
rect 3431 7745 3435 7749
rect 3455 7745 3459 7749
rect 3277 7739 3281 7743
rect 3115 7732 3119 7736
rect 4083 7767 4087 7771
rect 4127 7767 4131 7771
rect 4154 7767 4158 7771
rect 4199 7767 4203 7771
rect 4222 7739 4226 7743
rect 4058 7732 4062 7736
rect 2506 7718 2510 7722
rect 3451 7718 3455 7722
rect 2521 7710 2525 7714
rect 3466 7710 3470 7714
rect 3160 7704 3164 7708
rect 3197 7704 3201 7708
rect 3217 7704 3221 7708
rect 3255 7704 3259 7708
rect 4105 7704 4109 7708
rect 4142 7704 4146 7708
rect 4162 7704 4166 7708
rect 4200 7704 4204 7708
rect 2486 7695 2490 7699
rect 2510 7695 2514 7699
rect 3431 7695 3435 7699
rect 3455 7695 3459 7699
rect 3154 7684 3158 7688
rect 3172 7686 3176 7690
rect 2377 7674 2381 7678
rect 2414 7674 2418 7678
rect 2434 7674 2438 7678
rect 2472 7674 2476 7678
rect 2509 7674 2513 7678
rect 2546 7674 2550 7678
rect 2566 7674 2570 7678
rect 2604 7674 2608 7678
rect 2641 7674 2645 7678
rect 2678 7674 2682 7678
rect 2698 7674 2702 7678
rect 2736 7674 2740 7678
rect 3232 7686 3236 7690
rect 3190 7677 3194 7684
rect 3248 7677 3252 7684
rect 3267 7681 3271 7685
rect 4099 7684 4103 7688
rect 4117 7686 4121 7690
rect 3322 7674 3326 7678
rect 3359 7674 3363 7678
rect 3379 7674 3383 7678
rect 3417 7674 3421 7678
rect 3454 7674 3458 7678
rect 3491 7674 3495 7678
rect 3511 7674 3515 7678
rect 3549 7674 3553 7678
rect 3586 7674 3590 7678
rect 3623 7674 3627 7678
rect 3643 7674 3647 7678
rect 3681 7674 3685 7678
rect 4177 7686 4181 7690
rect 4135 7677 4139 7684
rect 4193 7677 4197 7684
rect 4212 7681 4216 7685
rect 3160 7663 3164 7667
rect 2371 7654 2375 7658
rect 2389 7656 2393 7660
rect 2449 7656 2453 7660
rect 2407 7647 2411 7654
rect 2465 7647 2469 7654
rect 2484 7651 2488 7655
rect 2502 7656 2506 7660
rect 2521 7656 2525 7660
rect 2581 7656 2585 7660
rect 2539 7647 2543 7654
rect 2597 7647 2601 7654
rect 2616 7651 2620 7655
rect 2634 7656 2638 7660
rect 2653 7656 2657 7660
rect 2713 7656 2717 7660
rect 2671 7647 2675 7654
rect 3197 7661 3201 7665
rect 3217 7661 3221 7665
rect 3253 7661 3257 7665
rect 4105 7663 4109 7667
rect 2729 7647 2733 7654
rect 2750 7651 2754 7655
rect 3316 7654 3320 7658
rect 3334 7656 3338 7660
rect 3394 7656 3398 7660
rect 3352 7647 3356 7654
rect 3410 7647 3414 7654
rect 3429 7651 3433 7655
rect 3447 7656 3451 7660
rect 3466 7656 3470 7660
rect 3526 7656 3530 7660
rect 3484 7647 3488 7654
rect 3542 7647 3546 7654
rect 3561 7651 3565 7655
rect 3579 7656 3583 7660
rect 3598 7656 3602 7660
rect 3658 7656 3662 7660
rect 3616 7647 3620 7654
rect 4142 7661 4146 7665
rect 4162 7661 4166 7665
rect 4198 7661 4202 7665
rect 3674 7647 3678 7654
rect 3695 7651 3699 7655
rect 2377 7633 2381 7637
rect 2414 7631 2418 7635
rect 2434 7631 2438 7635
rect 2470 7631 2474 7635
rect 2509 7633 2513 7637
rect 2546 7631 2550 7635
rect 2566 7631 2570 7635
rect 2602 7631 2606 7635
rect 2641 7633 2645 7637
rect 2678 7631 2682 7635
rect 2698 7631 2702 7635
rect 2734 7631 2738 7635
rect 3322 7633 3326 7637
rect 3359 7631 3363 7635
rect 3379 7631 3383 7635
rect 3415 7631 3419 7635
rect 3454 7633 3458 7637
rect 3491 7631 3495 7635
rect 3511 7631 3515 7635
rect 3547 7631 3551 7635
rect 3586 7633 3590 7637
rect 3623 7631 3627 7635
rect 3643 7631 3647 7635
rect 3679 7631 3683 7635
rect 3160 7618 3164 7622
rect 3197 7618 3201 7622
rect 3217 7618 3221 7622
rect 3255 7618 3259 7622
rect 4105 7618 4109 7622
rect 4142 7618 4146 7622
rect 4162 7618 4166 7622
rect 4200 7618 4204 7622
rect 3154 7598 3158 7602
rect 3172 7600 3176 7604
rect 2377 7588 2381 7592
rect 2414 7588 2418 7592
rect 2434 7588 2438 7592
rect 2472 7588 2476 7592
rect 2509 7588 2513 7592
rect 2546 7588 2550 7592
rect 2566 7588 2570 7592
rect 2604 7588 2608 7592
rect 2641 7588 2645 7592
rect 2678 7588 2682 7592
rect 2698 7588 2702 7592
rect 2736 7588 2740 7592
rect 3232 7600 3236 7604
rect 3190 7591 3194 7598
rect 3248 7591 3252 7598
rect 3267 7595 3271 7599
rect 3289 7593 3293 7597
rect 4099 7598 4103 7602
rect 4117 7600 4121 7604
rect 3322 7588 3326 7592
rect 3359 7588 3363 7592
rect 3379 7588 3383 7592
rect 3417 7588 3421 7592
rect 3454 7588 3458 7592
rect 3491 7588 3495 7592
rect 3511 7588 3515 7592
rect 3549 7588 3553 7592
rect 3586 7588 3590 7592
rect 3623 7588 3627 7592
rect 3643 7588 3647 7592
rect 3681 7588 3685 7592
rect 4177 7600 4181 7604
rect 4135 7591 4139 7598
rect 4193 7591 4197 7598
rect 4212 7595 4216 7599
rect 4234 7593 4238 7597
rect 3160 7577 3164 7581
rect 2371 7568 2375 7572
rect 2389 7570 2393 7574
rect 2449 7570 2453 7574
rect 2407 7561 2411 7568
rect 2465 7561 2469 7568
rect 2484 7565 2488 7569
rect 2502 7570 2506 7574
rect 2521 7570 2525 7574
rect 2581 7570 2585 7574
rect 2539 7561 2543 7568
rect 2597 7561 2601 7568
rect 2616 7565 2620 7569
rect 2634 7570 2638 7574
rect 2653 7570 2657 7574
rect 2713 7570 2717 7574
rect 2671 7561 2675 7568
rect 3197 7575 3201 7579
rect 3217 7575 3221 7579
rect 3253 7575 3257 7579
rect 4105 7577 4109 7581
rect 2729 7561 2733 7568
rect 2750 7565 2754 7569
rect 3316 7568 3320 7572
rect 3334 7570 3338 7574
rect 3394 7570 3398 7574
rect 3352 7561 3356 7568
rect 3410 7561 3414 7568
rect 3429 7565 3433 7569
rect 3447 7570 3451 7574
rect 3466 7570 3470 7574
rect 3526 7570 3530 7574
rect 3484 7561 3488 7568
rect 3542 7561 3546 7568
rect 3561 7565 3565 7569
rect 3579 7570 3583 7574
rect 3598 7570 3602 7574
rect 3658 7570 3662 7574
rect 3616 7561 3620 7568
rect 4142 7575 4146 7579
rect 4162 7575 4166 7579
rect 4198 7575 4202 7579
rect 3674 7561 3678 7568
rect 3695 7565 3699 7569
rect 2377 7547 2381 7551
rect 2414 7545 2418 7549
rect 2434 7545 2438 7549
rect 2470 7545 2474 7549
rect 2509 7547 2513 7551
rect 2546 7545 2550 7549
rect 2566 7545 2570 7549
rect 2602 7545 2606 7549
rect 2641 7547 2645 7551
rect 2678 7545 2682 7549
rect 2698 7545 2702 7549
rect 2734 7545 2738 7549
rect 3322 7547 3326 7551
rect 3359 7545 3363 7549
rect 3379 7545 3383 7549
rect 3415 7545 3419 7549
rect 3454 7547 3458 7551
rect 3491 7545 3495 7549
rect 3511 7545 3515 7549
rect 3547 7545 3551 7549
rect 3586 7547 3590 7551
rect 3623 7545 3627 7549
rect 3643 7545 3647 7549
rect 3679 7545 3683 7549
rect 2603 7517 2607 7521
rect 2627 7517 2631 7521
rect 3548 7517 3552 7521
rect 3572 7517 3576 7521
rect 2623 7492 2627 7496
rect 3568 7492 3572 7496
rect 2638 7484 2642 7488
rect 3583 7484 3587 7488
rect 2603 7469 2607 7473
rect 2627 7469 2631 7473
rect 3548 7469 3552 7473
rect 3572 7469 3576 7473
rect 3847 7472 3851 7476
rect 2377 7448 2381 7452
rect 2414 7448 2418 7452
rect 2434 7448 2438 7452
rect 2472 7448 2476 7452
rect 2509 7448 2513 7452
rect 2546 7448 2550 7452
rect 2566 7448 2570 7452
rect 2604 7448 2608 7452
rect 2641 7448 2645 7452
rect 2678 7448 2682 7452
rect 2698 7448 2702 7452
rect 2736 7448 2740 7452
rect 3322 7448 3326 7452
rect 3359 7448 3363 7452
rect 3379 7448 3383 7452
rect 3417 7448 3421 7452
rect 3454 7448 3458 7452
rect 3491 7448 3495 7452
rect 3511 7448 3515 7452
rect 3549 7448 3553 7452
rect 3586 7448 3590 7452
rect 3623 7448 3627 7452
rect 3643 7448 3647 7452
rect 3681 7448 3685 7452
rect 2371 7428 2375 7432
rect 2389 7430 2393 7434
rect 2449 7430 2453 7434
rect 2407 7421 2411 7428
rect 2465 7421 2469 7428
rect 2484 7425 2488 7429
rect 2502 7430 2506 7434
rect 2521 7430 2525 7434
rect 2581 7430 2585 7434
rect 2539 7421 2543 7428
rect 2597 7421 2601 7428
rect 2616 7425 2620 7429
rect 2634 7430 2638 7434
rect 2653 7430 2657 7434
rect 2713 7430 2717 7434
rect 2671 7421 2675 7428
rect 2729 7421 2733 7428
rect 2750 7425 2754 7429
rect 3316 7428 3320 7432
rect 3334 7430 3338 7434
rect 3394 7430 3398 7434
rect 3352 7421 3356 7428
rect 3410 7421 3414 7428
rect 3429 7425 3433 7429
rect 3447 7430 3451 7434
rect 3466 7430 3470 7434
rect 3526 7430 3530 7434
rect 3484 7421 3488 7428
rect 3542 7421 3546 7428
rect 3561 7425 3565 7429
rect 3579 7430 3583 7434
rect 3598 7430 3602 7434
rect 3658 7430 3662 7434
rect 3616 7421 3620 7428
rect 3674 7421 3678 7428
rect 3695 7425 3699 7429
rect 2377 7407 2381 7411
rect 2414 7405 2418 7409
rect 2434 7405 2438 7409
rect 2470 7405 2474 7409
rect 2509 7407 2513 7411
rect 2546 7405 2550 7409
rect 2566 7405 2570 7409
rect 2602 7405 2606 7409
rect 2641 7407 2645 7411
rect 2678 7405 2682 7409
rect 2698 7405 2702 7409
rect 2734 7405 2738 7409
rect 3322 7407 3326 7411
rect 3359 7405 3363 7409
rect 3379 7405 3383 7409
rect 3415 7405 3419 7409
rect 3454 7407 3458 7411
rect 3491 7405 3495 7409
rect 3511 7405 3515 7409
rect 3547 7405 3551 7409
rect 3586 7407 3590 7411
rect 3623 7405 3627 7409
rect 3643 7405 3647 7409
rect 3679 7405 3683 7409
rect 1489 6905 1493 6909
rect 1525 6905 1529 6909
rect 1545 6905 1549 6909
rect 1582 6903 1586 6907
rect 1621 6905 1625 6909
rect 1657 6905 1661 6909
rect 1677 6905 1681 6909
rect 1714 6903 1718 6907
rect 1753 6905 1757 6909
rect 1789 6905 1793 6909
rect 1809 6905 1813 6909
rect 1846 6903 1850 6907
rect 2434 6905 2438 6909
rect 2470 6905 2474 6909
rect 2490 6905 2494 6909
rect 2527 6903 2531 6907
rect 2566 6905 2570 6909
rect 2602 6905 2606 6909
rect 2622 6905 2626 6909
rect 2659 6903 2663 6907
rect 2698 6905 2702 6909
rect 2734 6905 2738 6909
rect 2754 6905 2758 6909
rect 2791 6903 2795 6907
rect 1473 6885 1477 6889
rect 1494 6886 1498 6893
rect 1552 6886 1556 6893
rect 1510 6880 1514 6884
rect 1570 6880 1574 6884
rect 1589 6880 1593 6884
rect 1607 6885 1611 6889
rect 1626 6886 1630 6893
rect 1684 6886 1688 6893
rect 1642 6880 1646 6884
rect 1702 6880 1706 6884
rect 1721 6880 1725 6884
rect 1739 6885 1743 6889
rect 1758 6886 1762 6893
rect 1816 6886 1820 6893
rect 1774 6880 1778 6884
rect 1834 6880 1838 6884
rect 1852 6882 1856 6886
rect 2418 6885 2422 6889
rect 2439 6886 2443 6893
rect 2497 6886 2501 6893
rect 2455 6880 2459 6884
rect 2515 6880 2519 6884
rect 2534 6880 2538 6884
rect 2552 6885 2556 6889
rect 2571 6886 2575 6893
rect 2629 6886 2633 6893
rect 2587 6880 2591 6884
rect 2647 6880 2651 6884
rect 2666 6880 2670 6884
rect 2684 6885 2688 6889
rect 2703 6886 2707 6893
rect 2761 6886 2765 6893
rect 2719 6880 2723 6884
rect 2779 6880 2783 6884
rect 2797 6882 2801 6886
rect 1487 6862 1491 6866
rect 1525 6862 1529 6866
rect 1545 6862 1549 6866
rect 1582 6862 1586 6866
rect 1619 6862 1623 6866
rect 1657 6862 1661 6866
rect 1677 6862 1681 6866
rect 1714 6862 1718 6866
rect 1751 6862 1755 6866
rect 1789 6862 1793 6866
rect 1809 6862 1813 6866
rect 1846 6862 1850 6866
rect 2432 6862 2436 6866
rect 2470 6862 2474 6866
rect 2490 6862 2494 6866
rect 2527 6862 2531 6866
rect 2564 6862 2568 6866
rect 2602 6862 2606 6866
rect 2622 6862 2626 6866
rect 2659 6862 2663 6866
rect 2696 6862 2700 6866
rect 2734 6862 2738 6866
rect 2754 6862 2758 6866
rect 2791 6862 2795 6866
rect 1596 6841 1600 6845
rect 1620 6841 1624 6845
rect 2541 6841 2545 6845
rect 2565 6841 2569 6845
rect 1585 6826 1589 6830
rect 2530 6826 2534 6830
rect 1600 6818 1604 6822
rect 2545 6818 2549 6822
rect 1596 6793 1600 6797
rect 1620 6793 1624 6797
rect 2541 6793 2545 6797
rect 2565 6793 2569 6797
rect 1489 6765 1493 6769
rect 1525 6765 1529 6769
rect 1545 6765 1549 6769
rect 1582 6763 1586 6767
rect 1621 6765 1625 6769
rect 1657 6765 1661 6769
rect 1677 6765 1681 6769
rect 1714 6763 1718 6767
rect 1753 6765 1757 6769
rect 1789 6765 1793 6769
rect 1809 6765 1813 6769
rect 1846 6763 1850 6767
rect 2434 6765 2438 6769
rect 2470 6765 2474 6769
rect 2490 6765 2494 6769
rect 2527 6763 2531 6767
rect 2566 6765 2570 6769
rect 2602 6765 2606 6769
rect 2622 6765 2626 6769
rect 2659 6763 2663 6767
rect 2698 6765 2702 6769
rect 2734 6765 2738 6769
rect 2754 6765 2758 6769
rect 2791 6763 2795 6767
rect 1473 6745 1477 6749
rect 1494 6746 1498 6753
rect 970 6735 974 6739
rect 1006 6735 1010 6739
rect 1026 6735 1030 6739
rect 1552 6746 1556 6753
rect 1510 6740 1514 6744
rect 1570 6740 1574 6744
rect 1589 6740 1593 6744
rect 1607 6745 1611 6749
rect 1626 6746 1630 6753
rect 1684 6746 1688 6753
rect 1642 6740 1646 6744
rect 1702 6740 1706 6744
rect 1721 6740 1725 6744
rect 1739 6745 1743 6749
rect 1758 6746 1762 6753
rect 1816 6746 1820 6753
rect 1774 6740 1778 6744
rect 1834 6740 1838 6744
rect 1852 6742 1856 6746
rect 2418 6745 2422 6749
rect 2439 6746 2443 6753
rect 1063 6733 1067 6737
rect 1915 6735 1919 6739
rect 1951 6735 1955 6739
rect 1971 6735 1975 6739
rect 2497 6746 2501 6753
rect 2455 6740 2459 6744
rect 2515 6740 2519 6744
rect 2534 6740 2538 6744
rect 2552 6745 2556 6749
rect 2571 6746 2575 6753
rect 2629 6746 2633 6753
rect 2587 6740 2591 6744
rect 2647 6740 2651 6744
rect 2666 6740 2670 6744
rect 2684 6745 2688 6749
rect 2703 6746 2707 6753
rect 2761 6746 2765 6753
rect 2719 6740 2723 6744
rect 2779 6740 2783 6744
rect 2797 6742 2801 6746
rect 2008 6733 2012 6737
rect 934 6717 938 6721
rect 956 6715 960 6719
rect 975 6716 979 6723
rect 1033 6716 1037 6723
rect 991 6710 995 6714
rect 1487 6722 1491 6726
rect 1525 6722 1529 6726
rect 1545 6722 1549 6726
rect 1582 6722 1586 6726
rect 1619 6722 1623 6726
rect 1657 6722 1661 6726
rect 1677 6722 1681 6726
rect 1714 6722 1718 6726
rect 1751 6722 1755 6726
rect 1789 6722 1793 6726
rect 1809 6722 1813 6726
rect 1846 6722 1850 6726
rect 1051 6710 1055 6714
rect 1069 6712 1073 6716
rect 1879 6717 1883 6721
rect 1901 6715 1905 6719
rect 1920 6716 1924 6723
rect 1978 6716 1982 6723
rect 1936 6710 1940 6714
rect 2432 6722 2436 6726
rect 2470 6722 2474 6726
rect 2490 6722 2494 6726
rect 2527 6722 2531 6726
rect 2564 6722 2568 6726
rect 2602 6722 2606 6726
rect 2622 6722 2626 6726
rect 2659 6722 2663 6726
rect 2696 6722 2700 6726
rect 2734 6722 2738 6726
rect 2754 6722 2758 6726
rect 2791 6722 2795 6726
rect 1996 6710 2000 6714
rect 2014 6712 2018 6716
rect 968 6692 972 6696
rect 1006 6692 1010 6696
rect 1026 6692 1030 6696
rect 1063 6692 1067 6696
rect 1913 6692 1917 6696
rect 1951 6692 1955 6696
rect 1971 6692 1975 6696
rect 2008 6692 2012 6696
rect 1489 6679 1493 6683
rect 1525 6679 1529 6683
rect 1545 6679 1549 6683
rect 1582 6677 1586 6681
rect 1621 6679 1625 6683
rect 1657 6679 1661 6683
rect 1677 6679 1681 6683
rect 1714 6677 1718 6681
rect 1753 6679 1757 6683
rect 1789 6679 1793 6683
rect 1809 6679 1813 6683
rect 1846 6677 1850 6681
rect 2434 6679 2438 6683
rect 2470 6679 2474 6683
rect 2490 6679 2494 6683
rect 2527 6677 2531 6681
rect 2566 6679 2570 6683
rect 2602 6679 2606 6683
rect 2622 6679 2626 6683
rect 2659 6677 2663 6681
rect 2698 6679 2702 6683
rect 2734 6679 2738 6683
rect 2754 6679 2758 6683
rect 2791 6677 2795 6681
rect 1473 6659 1477 6663
rect 1494 6660 1498 6667
rect 970 6649 974 6653
rect 1006 6649 1010 6653
rect 1026 6649 1030 6653
rect 1552 6660 1556 6667
rect 1510 6654 1514 6658
rect 1570 6654 1574 6658
rect 1589 6654 1593 6658
rect 1607 6659 1611 6663
rect 1626 6660 1630 6667
rect 1684 6660 1688 6667
rect 1642 6654 1646 6658
rect 1702 6654 1706 6658
rect 1721 6654 1725 6658
rect 1739 6659 1743 6663
rect 1758 6660 1762 6667
rect 1816 6660 1820 6667
rect 1774 6654 1778 6658
rect 1834 6654 1838 6658
rect 1852 6656 1856 6660
rect 2418 6659 2422 6663
rect 2439 6660 2443 6667
rect 1063 6647 1067 6651
rect 1915 6649 1919 6653
rect 1951 6649 1955 6653
rect 1971 6649 1975 6653
rect 2497 6660 2501 6667
rect 2455 6654 2459 6658
rect 2515 6654 2519 6658
rect 2534 6654 2538 6658
rect 2552 6659 2556 6663
rect 2571 6660 2575 6667
rect 2629 6660 2633 6667
rect 2587 6654 2591 6658
rect 2647 6654 2651 6658
rect 2666 6654 2670 6658
rect 2684 6659 2688 6663
rect 2703 6660 2707 6667
rect 2761 6660 2765 6667
rect 2719 6654 2723 6658
rect 2779 6654 2783 6658
rect 2797 6656 2801 6660
rect 2008 6647 2012 6651
rect 956 6629 960 6633
rect 975 6630 979 6637
rect 1033 6630 1037 6637
rect 991 6624 995 6628
rect 1487 6636 1491 6640
rect 1525 6636 1529 6640
rect 1545 6636 1549 6640
rect 1582 6636 1586 6640
rect 1619 6636 1623 6640
rect 1657 6636 1661 6640
rect 1677 6636 1681 6640
rect 1714 6636 1718 6640
rect 1751 6636 1755 6640
rect 1789 6636 1793 6640
rect 1809 6636 1813 6640
rect 1846 6636 1850 6640
rect 1051 6624 1055 6628
rect 1069 6626 1073 6630
rect 1901 6629 1905 6633
rect 1920 6630 1924 6637
rect 1978 6630 1982 6637
rect 1936 6624 1940 6628
rect 2432 6636 2436 6640
rect 2470 6636 2474 6640
rect 2490 6636 2494 6640
rect 2527 6636 2531 6640
rect 2564 6636 2568 6640
rect 2602 6636 2606 6640
rect 2622 6636 2626 6640
rect 2659 6636 2663 6640
rect 2696 6636 2700 6640
rect 2734 6636 2738 6640
rect 2754 6636 2758 6640
rect 2791 6636 2795 6640
rect 1996 6624 2000 6628
rect 2014 6626 2018 6630
rect 1713 6615 1717 6619
rect 1737 6615 1741 6619
rect 2658 6615 2662 6619
rect 2682 6615 2686 6619
rect 968 6606 972 6610
rect 1006 6606 1010 6610
rect 1026 6606 1030 6610
rect 1063 6606 1067 6610
rect 1913 6606 1917 6610
rect 1951 6606 1955 6610
rect 1971 6606 1975 6610
rect 2008 6606 2012 6610
rect 1702 6600 1706 6604
rect 2647 6600 2651 6604
rect 1717 6592 1721 6596
rect 2662 6592 2666 6596
rect 1110 6578 1114 6582
rect 946 6571 950 6575
rect 969 6543 973 6547
rect 1014 6543 1018 6547
rect 1041 6543 1045 6547
rect 1085 6543 1089 6547
rect 2053 6578 2057 6582
rect 1891 6571 1895 6575
rect 1713 6565 1717 6569
rect 1737 6565 1741 6569
rect 1159 6550 1163 6554
rect 1230 6543 1234 6547
rect 1275 6543 1279 6547
rect 1302 6543 1306 6547
rect 1346 6543 1350 6547
rect 1914 6543 1918 6547
rect 1959 6543 1963 6547
rect 1986 6543 1990 6547
rect 2030 6543 2034 6547
rect 955 6523 959 6527
rect 982 6523 986 6527
rect 998 6524 1002 6528
rect 1054 6523 1058 6527
rect 1073 6524 1077 6528
rect 1130 6523 1134 6527
rect 1166 6530 1172 6534
rect 1489 6537 1493 6541
rect 1525 6537 1529 6541
rect 1545 6537 1549 6541
rect 1582 6535 1586 6539
rect 1621 6537 1625 6541
rect 1657 6537 1661 6541
rect 1677 6537 1681 6541
rect 1714 6535 1718 6539
rect 1753 6537 1757 6541
rect 1789 6537 1793 6541
rect 1809 6537 1813 6541
rect 2658 6565 2662 6569
rect 2682 6565 2686 6569
rect 2104 6550 2108 6554
rect 1846 6535 1850 6539
rect 2175 6543 2179 6547
rect 2220 6543 2224 6547
rect 2247 6543 2251 6547
rect 2291 6543 2295 6547
rect 1216 6523 1220 6527
rect 1243 6523 1247 6527
rect 1259 6524 1263 6528
rect 1315 6523 1319 6527
rect 1334 6524 1338 6528
rect 1366 6523 1370 6527
rect 1157 6514 1161 6518
rect 1473 6517 1477 6521
rect 1494 6518 1498 6525
rect 972 6505 976 6509
rect 1018 6506 1023 6510
rect 1044 6505 1048 6509
rect 1088 6506 1092 6510
rect 1233 6505 1237 6509
rect 1279 6506 1284 6510
rect 1305 6505 1309 6509
rect 1349 6506 1353 6510
rect 1552 6518 1556 6525
rect 1510 6512 1514 6516
rect 1570 6512 1574 6516
rect 1589 6512 1593 6516
rect 1607 6517 1611 6521
rect 1626 6518 1630 6525
rect 1684 6518 1688 6525
rect 1642 6512 1646 6516
rect 1702 6512 1706 6516
rect 1721 6512 1725 6516
rect 1739 6517 1743 6521
rect 1758 6518 1762 6525
rect 1816 6518 1820 6525
rect 1774 6512 1778 6516
rect 1900 6523 1904 6527
rect 1927 6523 1931 6527
rect 1943 6524 1947 6528
rect 1999 6523 2003 6527
rect 2018 6524 2022 6528
rect 2075 6523 2079 6527
rect 2111 6530 2117 6534
rect 2434 6537 2438 6541
rect 2470 6537 2474 6541
rect 2490 6537 2494 6541
rect 2527 6535 2531 6539
rect 2566 6537 2570 6541
rect 2602 6537 2606 6541
rect 2622 6537 2626 6541
rect 2659 6535 2663 6539
rect 2698 6537 2702 6541
rect 2734 6537 2738 6541
rect 2754 6537 2758 6541
rect 2791 6535 2795 6539
rect 2161 6523 2165 6527
rect 2188 6523 2192 6527
rect 2204 6524 2208 6528
rect 2260 6523 2264 6527
rect 2279 6524 2283 6528
rect 2311 6523 2315 6527
rect 1834 6512 1838 6516
rect 1852 6514 1856 6518
rect 2102 6514 2106 6518
rect 2418 6517 2422 6521
rect 2439 6518 2443 6525
rect 1917 6505 1921 6509
rect 1963 6506 1968 6510
rect 1989 6505 1993 6509
rect 2033 6506 2037 6510
rect 2178 6505 2182 6509
rect 2224 6506 2229 6510
rect 2250 6505 2254 6509
rect 2294 6506 2298 6510
rect 2497 6518 2501 6525
rect 2455 6512 2459 6516
rect 2515 6512 2519 6516
rect 2534 6512 2538 6516
rect 2552 6517 2556 6521
rect 2571 6518 2575 6525
rect 2629 6518 2633 6525
rect 2587 6512 2591 6516
rect 2647 6512 2651 6516
rect 2666 6512 2670 6516
rect 2684 6517 2688 6521
rect 2703 6518 2707 6525
rect 2761 6518 2765 6525
rect 2719 6512 2723 6516
rect 2779 6512 2783 6516
rect 2797 6514 2801 6518
rect 1487 6494 1491 6498
rect 1525 6494 1529 6498
rect 1545 6494 1549 6498
rect 1582 6494 1586 6498
rect 1619 6494 1623 6498
rect 1657 6494 1661 6498
rect 1677 6494 1681 6498
rect 1714 6494 1718 6498
rect 1751 6494 1755 6498
rect 1789 6494 1793 6498
rect 1809 6494 1813 6498
rect 1846 6494 1850 6498
rect 2432 6494 2436 6498
rect 2470 6494 2474 6498
rect 2490 6494 2494 6498
rect 2527 6494 2531 6498
rect 2564 6494 2568 6498
rect 2602 6494 2606 6498
rect 2622 6494 2626 6498
rect 2659 6494 2663 6498
rect 2696 6494 2700 6498
rect 2734 6494 2738 6498
rect 2754 6494 2758 6498
rect 2791 6494 2795 6498
rect 1233 6477 1237 6481
rect 1279 6476 1284 6480
rect 1305 6477 1309 6481
rect 1349 6476 1353 6480
rect 2178 6477 2182 6481
rect 2224 6476 2229 6480
rect 2250 6477 2254 6481
rect 2294 6476 2298 6480
rect 1159 6468 1163 6472
rect 1138 6454 1142 6458
rect 1216 6459 1220 6463
rect 1243 6459 1247 6463
rect 1259 6458 1263 6462
rect 1315 6459 1319 6463
rect 1334 6458 1338 6462
rect 2104 6468 2108 6472
rect 1366 6459 1370 6463
rect 1165 6450 1169 6454
rect 1230 6439 1234 6443
rect 1275 6439 1279 6443
rect 1302 6439 1306 6443
rect 1346 6439 1350 6443
rect 2083 6454 2087 6458
rect 2161 6459 2165 6463
rect 2188 6459 2192 6463
rect 2204 6458 2208 6462
rect 2260 6459 2264 6463
rect 2279 6458 2283 6462
rect 2311 6459 2315 6463
rect 2110 6450 2114 6454
rect 1157 6432 1161 6436
rect 2175 6439 2179 6443
rect 2220 6439 2224 6443
rect 2247 6439 2251 6443
rect 2291 6439 2295 6443
rect 2102 6432 2106 6436
rect 988 6414 992 6418
rect 1078 6414 1082 6418
rect 1159 6414 1163 6418
rect 1230 6411 1234 6415
rect 1275 6411 1279 6415
rect 1302 6411 1306 6415
rect 1346 6411 1350 6415
rect 1933 6414 1937 6418
rect 2023 6414 2027 6418
rect 2104 6414 2108 6418
rect 2175 6411 2179 6415
rect 2220 6411 2224 6415
rect 2247 6411 2251 6415
rect 2291 6411 2295 6415
rect 995 6394 1001 6398
rect 1085 6394 1091 6398
rect 1166 6394 1172 6398
rect 1216 6391 1220 6395
rect 1243 6391 1247 6395
rect 1259 6392 1263 6396
rect 1315 6391 1319 6395
rect 1334 6392 1338 6396
rect 1366 6391 1370 6395
rect 1940 6394 1946 6398
rect 2030 6394 2036 6398
rect 2111 6394 2117 6398
rect 2161 6391 2165 6395
rect 2188 6391 2192 6395
rect 2204 6392 2208 6396
rect 2260 6391 2264 6395
rect 2279 6392 2283 6396
rect 2311 6391 2315 6395
rect 986 6378 990 6382
rect 1076 6378 1080 6382
rect 1157 6378 1161 6382
rect 1233 6373 1237 6377
rect 1279 6374 1284 6378
rect 1931 6378 1935 6382
rect 2021 6378 2025 6382
rect 2102 6378 2106 6382
rect 1305 6373 1309 6377
rect 1349 6374 1353 6378
rect 2178 6373 2182 6377
rect 2224 6374 2229 6378
rect 2250 6373 2254 6377
rect 2294 6374 2298 6378
rect 1233 6345 1237 6349
rect 1279 6344 1284 6348
rect 1305 6345 1309 6349
rect 1349 6344 1353 6348
rect 2178 6345 2182 6349
rect 2224 6344 2229 6348
rect 2250 6345 2254 6349
rect 2294 6344 2298 6348
rect 988 6336 992 6340
rect 1078 6336 1082 6340
rect 1159 6336 1163 6340
rect 967 6322 971 6326
rect 994 6318 998 6322
rect 1021 6314 1025 6318
rect 1057 6322 1061 6326
rect 1084 6318 1088 6322
rect 986 6300 990 6304
rect 1111 6314 1115 6318
rect 1138 6322 1142 6326
rect 1216 6327 1220 6331
rect 1243 6327 1247 6331
rect 1259 6326 1263 6330
rect 1315 6327 1319 6331
rect 1334 6326 1338 6330
rect 1933 6336 1937 6340
rect 2023 6336 2027 6340
rect 2104 6336 2108 6340
rect 1366 6327 1370 6331
rect 1165 6318 1169 6322
rect 1076 6300 1080 6304
rect 1230 6307 1234 6311
rect 1275 6307 1279 6311
rect 1302 6307 1306 6311
rect 1346 6307 1350 6311
rect 1912 6322 1916 6326
rect 1939 6318 1943 6322
rect 1157 6300 1161 6304
rect 1966 6314 1970 6318
rect 2002 6322 2006 6326
rect 2029 6318 2033 6322
rect 1931 6300 1935 6304
rect 2056 6314 2060 6318
rect 2083 6322 2087 6326
rect 2161 6327 2165 6331
rect 2188 6327 2192 6331
rect 2204 6326 2208 6330
rect 2260 6327 2264 6331
rect 2279 6326 2283 6330
rect 2311 6327 2315 6331
rect 2110 6318 2114 6322
rect 2021 6300 2025 6304
rect 2175 6307 2179 6311
rect 2220 6307 2224 6311
rect 2247 6307 2251 6311
rect 2291 6307 2295 6311
rect 2102 6300 2106 6304
rect 1054 6279 1058 6283
rect 1159 6279 1163 6283
rect 1230 6279 1234 6283
rect 1275 6279 1279 6283
rect 1302 6279 1306 6283
rect 1346 6279 1350 6283
rect 1999 6279 2003 6283
rect 2104 6279 2108 6283
rect 2175 6279 2179 6283
rect 2220 6279 2224 6283
rect 2247 6279 2251 6283
rect 2291 6279 2295 6283
rect 1061 6259 1067 6263
rect 1166 6259 1172 6263
rect 1216 6259 1220 6263
rect 1243 6259 1247 6263
rect 1259 6260 1263 6264
rect 1315 6259 1319 6263
rect 1334 6260 1338 6264
rect 1366 6259 1370 6263
rect 2006 6259 2012 6263
rect 2111 6259 2117 6263
rect 2161 6259 2165 6263
rect 2188 6259 2192 6263
rect 2204 6260 2208 6264
rect 2260 6259 2264 6263
rect 2279 6260 2283 6264
rect 2311 6259 2315 6263
rect 1052 6243 1056 6247
rect 1157 6243 1161 6247
rect 1233 6241 1237 6245
rect 1279 6242 1284 6246
rect 1305 6241 1309 6245
rect 1349 6242 1353 6246
rect 1997 6243 2001 6247
rect 2102 6243 2106 6247
rect 2178 6241 2182 6245
rect 2224 6242 2229 6246
rect 2250 6241 2254 6245
rect 2294 6242 2298 6246
rect 1233 6213 1237 6217
rect 1279 6212 1284 6216
rect 1305 6213 1309 6217
rect 1349 6212 1353 6216
rect 2178 6213 2182 6217
rect 2224 6212 2229 6216
rect 2250 6213 2254 6217
rect 2294 6212 2298 6216
rect 1054 6204 1058 6208
rect 1159 6204 1163 6208
rect 1033 6190 1037 6194
rect 1060 6186 1064 6190
rect 1087 6182 1091 6186
rect 1138 6190 1142 6194
rect 1216 6195 1220 6199
rect 1243 6195 1247 6199
rect 1259 6194 1263 6198
rect 1315 6195 1319 6199
rect 1334 6194 1338 6198
rect 1999 6204 2003 6208
rect 2104 6204 2108 6208
rect 1366 6195 1370 6199
rect 1165 6186 1169 6190
rect 1052 6168 1056 6172
rect 1230 6175 1234 6179
rect 1275 6175 1279 6179
rect 1302 6175 1306 6179
rect 1346 6175 1350 6179
rect 1978 6190 1982 6194
rect 2005 6186 2009 6190
rect 1157 6168 1161 6172
rect 2032 6182 2036 6186
rect 2083 6190 2087 6194
rect 2161 6195 2165 6199
rect 2188 6195 2192 6199
rect 2204 6194 2208 6198
rect 2260 6195 2264 6199
rect 2279 6194 2283 6198
rect 2311 6195 2315 6199
rect 2110 6186 2114 6190
rect 1997 6168 2001 6172
rect 2175 6175 2179 6179
rect 2220 6175 2224 6179
rect 2247 6175 2251 6179
rect 2291 6175 2295 6179
rect 2102 6168 2106 6172
rect 1078 6148 1082 6152
rect 1159 6148 1163 6152
rect 1230 6147 1234 6151
rect 1275 6147 1279 6151
rect 1302 6147 1306 6151
rect 1346 6147 1350 6151
rect 2023 6148 2027 6152
rect 2104 6148 2108 6152
rect 2175 6147 2179 6151
rect 2220 6147 2224 6151
rect 2247 6147 2251 6151
rect 2291 6147 2295 6151
rect 1085 6128 1091 6132
rect 1166 6128 1172 6132
rect 1216 6127 1220 6131
rect 1243 6127 1247 6131
rect 1259 6128 1263 6132
rect 1315 6127 1319 6131
rect 1334 6128 1338 6132
rect 1619 6135 1623 6139
rect 1656 6137 1660 6141
rect 1676 6137 1680 6141
rect 1712 6137 1716 6141
rect 1366 6127 1370 6131
rect 1076 6112 1080 6116
rect 1157 6112 1161 6116
rect 1233 6109 1237 6113
rect 1279 6110 1284 6114
rect 1613 6114 1617 6118
rect 1305 6109 1309 6113
rect 1349 6110 1353 6114
rect 1631 6112 1635 6116
rect 1649 6118 1653 6125
rect 1707 6118 1711 6125
rect 1691 6112 1695 6116
rect 1726 6117 1730 6121
rect 2030 6128 2036 6132
rect 2111 6128 2117 6132
rect 2161 6127 2165 6131
rect 2188 6127 2192 6131
rect 2204 6128 2208 6132
rect 2260 6127 2264 6131
rect 2279 6128 2283 6132
rect 2564 6135 2568 6139
rect 2601 6137 2605 6141
rect 2621 6137 2625 6141
rect 2657 6137 2661 6141
rect 2311 6127 2315 6131
rect 2021 6112 2025 6116
rect 2102 6112 2106 6116
rect 2178 6109 2182 6113
rect 2224 6110 2229 6114
rect 2558 6114 2562 6118
rect 2250 6109 2254 6113
rect 2294 6110 2298 6114
rect 2576 6112 2580 6116
rect 2594 6118 2598 6125
rect 2652 6118 2656 6125
rect 2636 6112 2640 6116
rect 2671 6117 2675 6121
rect 1619 6094 1623 6098
rect 1656 6094 1660 6098
rect 1676 6094 1680 6098
rect 1714 6094 1718 6098
rect 2564 6094 2568 6098
rect 2601 6094 2605 6098
rect 2621 6094 2625 6098
rect 2659 6094 2663 6098
rect 1233 6081 1237 6085
rect 1279 6080 1284 6084
rect 1305 6081 1309 6085
rect 1349 6080 1353 6084
rect 2178 6081 2182 6085
rect 2224 6080 2229 6084
rect 2250 6081 2254 6085
rect 2294 6080 2298 6084
rect 1078 6072 1082 6076
rect 1159 6072 1163 6076
rect 1057 6058 1061 6062
rect 1084 6054 1088 6058
rect 1111 6050 1115 6054
rect 1138 6058 1142 6062
rect 1165 6054 1169 6058
rect 1076 6036 1080 6040
rect 1216 6063 1220 6067
rect 1243 6063 1247 6067
rect 1259 6062 1263 6066
rect 1315 6063 1319 6067
rect 1334 6062 1338 6066
rect 2023 6072 2027 6076
rect 1366 6063 1370 6067
rect 1713 6065 1717 6069
rect 2104 6072 2108 6076
rect 1192 6050 1196 6054
rect 1596 6056 1600 6060
rect 1157 6036 1161 6040
rect 1230 6043 1234 6047
rect 1275 6043 1279 6047
rect 1302 6043 1306 6047
rect 1346 6043 1350 6047
rect 2002 6058 2006 6062
rect 2029 6054 2033 6058
rect 1621 6035 1625 6039
rect 1657 6035 1661 6039
rect 1677 6035 1681 6039
rect 2056 6050 2060 6054
rect 2083 6058 2087 6062
rect 2110 6054 2114 6058
rect 1714 6033 1718 6037
rect 2021 6036 2025 6040
rect 2161 6063 2165 6067
rect 2188 6063 2192 6067
rect 2204 6062 2208 6066
rect 2260 6063 2264 6067
rect 2279 6062 2283 6066
rect 2311 6063 2315 6067
rect 2658 6065 2662 6069
rect 2137 6050 2141 6054
rect 2541 6056 2545 6060
rect 2102 6036 2106 6040
rect 2175 6043 2179 6047
rect 2220 6043 2224 6047
rect 2247 6043 2251 6047
rect 2291 6043 2295 6047
rect 2566 6035 2570 6039
rect 2602 6035 2606 6039
rect 2622 6035 2626 6039
rect 2659 6033 2663 6037
rect 1607 6015 1611 6019
rect 1626 6016 1630 6023
rect 1684 6016 1688 6023
rect 1642 6010 1646 6014
rect 1702 6010 1706 6014
rect 1720 6012 1724 6016
rect 2552 6015 2556 6019
rect 2571 6016 2575 6023
rect 2629 6016 2633 6023
rect 2587 6010 2591 6014
rect 2647 6010 2651 6014
rect 2665 6012 2669 6016
rect 873 6002 877 6006
rect 909 6002 913 6006
rect 929 6002 933 6006
rect 966 6000 970 6004
rect 1005 6002 1009 6006
rect 1041 6002 1045 6006
rect 1061 6002 1065 6006
rect 1098 6000 1102 6004
rect 1137 6002 1141 6006
rect 1173 6002 1177 6006
rect 1193 6002 1197 6006
rect 1230 6000 1234 6004
rect 1269 6002 1273 6006
rect 1305 6002 1309 6006
rect 1325 6002 1329 6006
rect 1362 6000 1366 6004
rect 1818 6002 1822 6006
rect 1854 6002 1858 6006
rect 1874 6002 1878 6006
rect 1911 6000 1915 6004
rect 1950 6002 1954 6006
rect 1986 6002 1990 6006
rect 2006 6002 2010 6006
rect 2043 6000 2047 6004
rect 2082 6002 2086 6006
rect 2118 6002 2122 6006
rect 2138 6002 2142 6006
rect 2175 6000 2179 6004
rect 2214 6002 2218 6006
rect 2250 6002 2254 6006
rect 2270 6002 2274 6006
rect 2307 6000 2311 6004
rect 857 5982 861 5986
rect 878 5983 882 5990
rect 936 5983 940 5990
rect 894 5977 898 5981
rect 954 5977 958 5981
rect 972 5979 976 5983
rect 989 5982 993 5986
rect 1010 5983 1014 5990
rect 1068 5983 1072 5990
rect 1026 5977 1030 5981
rect 1086 5977 1090 5981
rect 1104 5979 1108 5983
rect 1121 5982 1125 5986
rect 1142 5983 1146 5990
rect 1200 5983 1204 5990
rect 1158 5977 1162 5981
rect 1218 5977 1222 5981
rect 1236 5979 1240 5983
rect 1253 5982 1257 5986
rect 1274 5983 1278 5990
rect 1332 5983 1336 5990
rect 1290 5977 1294 5981
rect 1619 5992 1623 5996
rect 1657 5992 1661 5996
rect 1677 5992 1681 5996
rect 1714 5992 1718 5996
rect 1350 5977 1354 5981
rect 1368 5979 1372 5983
rect 1802 5982 1806 5986
rect 1823 5983 1827 5990
rect 1881 5983 1885 5990
rect 1839 5977 1843 5981
rect 1899 5977 1903 5981
rect 1917 5979 1921 5983
rect 1934 5982 1938 5986
rect 1955 5983 1959 5990
rect 2013 5983 2017 5990
rect 1971 5977 1975 5981
rect 2031 5977 2035 5981
rect 2049 5979 2053 5983
rect 2066 5982 2070 5986
rect 2087 5983 2091 5990
rect 2145 5983 2149 5990
rect 2103 5977 2107 5981
rect 2163 5977 2167 5981
rect 2181 5979 2185 5983
rect 2198 5982 2202 5986
rect 2219 5983 2223 5990
rect 2277 5983 2281 5990
rect 2235 5977 2239 5981
rect 2564 5992 2568 5996
rect 2602 5992 2606 5996
rect 2622 5992 2626 5996
rect 2659 5992 2663 5996
rect 2295 5977 2299 5981
rect 2313 5979 2317 5983
rect 871 5959 875 5963
rect 909 5959 913 5963
rect 929 5959 933 5963
rect 966 5959 970 5963
rect 1003 5959 1007 5963
rect 1041 5959 1045 5963
rect 1061 5959 1065 5963
rect 1098 5959 1102 5963
rect 1135 5959 1139 5963
rect 1173 5959 1177 5963
rect 1193 5959 1197 5963
rect 1230 5959 1234 5963
rect 1267 5959 1271 5963
rect 1305 5959 1309 5963
rect 1325 5959 1329 5963
rect 1362 5959 1366 5963
rect 1816 5959 1820 5963
rect 1854 5959 1858 5963
rect 1874 5959 1878 5963
rect 1911 5959 1915 5963
rect 1948 5959 1952 5963
rect 1986 5959 1990 5963
rect 2006 5959 2010 5963
rect 2043 5959 2047 5963
rect 2080 5959 2084 5963
rect 2118 5959 2122 5963
rect 2138 5959 2142 5963
rect 2175 5959 2179 5963
rect 2212 5959 2216 5963
rect 2250 5959 2254 5963
rect 2270 5959 2274 5963
rect 2307 5959 2311 5963
rect 1489 5923 1493 5927
rect 1525 5923 1529 5927
rect 1545 5923 1549 5927
rect 1582 5921 1586 5925
rect 1621 5923 1625 5927
rect 1657 5923 1661 5927
rect 1677 5923 1681 5927
rect 1714 5921 1718 5925
rect 1753 5923 1757 5927
rect 1789 5923 1793 5927
rect 1809 5923 1813 5927
rect 1846 5921 1850 5925
rect 2434 5923 2438 5927
rect 2470 5923 2474 5927
rect 2490 5923 2494 5927
rect 2527 5921 2531 5925
rect 2566 5923 2570 5927
rect 2602 5923 2606 5927
rect 2622 5923 2626 5927
rect 2659 5921 2663 5925
rect 2698 5923 2702 5927
rect 2734 5923 2738 5927
rect 2754 5923 2758 5927
rect 2791 5921 2795 5925
rect 1473 5903 1477 5907
rect 1494 5904 1498 5911
rect 1552 5904 1556 5911
rect 1510 5898 1514 5902
rect 1570 5898 1574 5902
rect 1589 5898 1593 5902
rect 1607 5903 1611 5907
rect 1626 5904 1630 5911
rect 1684 5904 1688 5911
rect 1642 5898 1646 5902
rect 1702 5898 1706 5902
rect 1721 5898 1725 5902
rect 1739 5903 1743 5907
rect 1758 5904 1762 5911
rect 1816 5904 1820 5911
rect 1774 5898 1778 5902
rect 1834 5898 1838 5902
rect 1852 5900 1856 5904
rect 2418 5903 2422 5907
rect 2439 5904 2443 5911
rect 2497 5904 2501 5911
rect 2455 5898 2459 5902
rect 2515 5898 2519 5902
rect 2534 5898 2538 5902
rect 2552 5903 2556 5907
rect 2571 5904 2575 5911
rect 2629 5904 2633 5911
rect 2587 5898 2591 5902
rect 2647 5898 2651 5902
rect 2666 5898 2670 5902
rect 2684 5903 2688 5907
rect 2703 5904 2707 5911
rect 2761 5904 2765 5911
rect 2719 5898 2723 5902
rect 2779 5898 2783 5902
rect 2797 5900 2801 5904
rect 1487 5880 1491 5884
rect 1525 5880 1529 5884
rect 1545 5880 1549 5884
rect 1582 5880 1586 5884
rect 1619 5880 1623 5884
rect 1657 5880 1661 5884
rect 1677 5880 1681 5884
rect 1714 5880 1718 5884
rect 1751 5880 1755 5884
rect 1789 5880 1793 5884
rect 1809 5880 1813 5884
rect 1846 5880 1850 5884
rect 2432 5880 2436 5884
rect 2470 5880 2474 5884
rect 2490 5880 2494 5884
rect 2527 5880 2531 5884
rect 2564 5880 2568 5884
rect 2602 5880 2606 5884
rect 2622 5880 2626 5884
rect 2659 5880 2663 5884
rect 2696 5880 2700 5884
rect 2734 5880 2738 5884
rect 2754 5880 2758 5884
rect 2791 5880 2795 5884
rect 1596 5859 1600 5863
rect 1620 5859 1624 5863
rect 2541 5859 2545 5863
rect 2565 5859 2569 5863
rect 1585 5844 1589 5848
rect 2530 5844 2534 5848
rect 1600 5836 1604 5840
rect 2545 5836 2549 5840
rect 1596 5811 1600 5815
rect 1620 5811 1624 5815
rect 2541 5811 2545 5815
rect 2565 5811 2569 5815
rect 1489 5783 1493 5787
rect 1525 5783 1529 5787
rect 1545 5783 1549 5787
rect 1582 5781 1586 5785
rect 1621 5783 1625 5787
rect 1657 5783 1661 5787
rect 1677 5783 1681 5787
rect 1714 5781 1718 5785
rect 1753 5783 1757 5787
rect 1789 5783 1793 5787
rect 1809 5783 1813 5787
rect 1846 5781 1850 5785
rect 2434 5783 2438 5787
rect 2470 5783 2474 5787
rect 2490 5783 2494 5787
rect 2527 5781 2531 5785
rect 2566 5783 2570 5787
rect 2602 5783 2606 5787
rect 2622 5783 2626 5787
rect 2659 5781 2663 5785
rect 2698 5783 2702 5787
rect 2734 5783 2738 5787
rect 2754 5783 2758 5787
rect 2791 5781 2795 5785
rect 1473 5763 1477 5767
rect 1494 5764 1498 5771
rect 970 5753 974 5757
rect 1006 5753 1010 5757
rect 1026 5753 1030 5757
rect 1552 5764 1556 5771
rect 1510 5758 1514 5762
rect 1570 5758 1574 5762
rect 1589 5758 1593 5762
rect 1607 5763 1611 5767
rect 1626 5764 1630 5771
rect 1684 5764 1688 5771
rect 1642 5758 1646 5762
rect 1702 5758 1706 5762
rect 1721 5758 1725 5762
rect 1739 5763 1743 5767
rect 1758 5764 1762 5771
rect 1816 5764 1820 5771
rect 1774 5758 1778 5762
rect 1834 5758 1838 5762
rect 1852 5760 1856 5764
rect 2418 5763 2422 5767
rect 2439 5764 2443 5771
rect 1063 5751 1067 5755
rect 1915 5753 1919 5757
rect 1951 5753 1955 5757
rect 1971 5753 1975 5757
rect 2497 5764 2501 5771
rect 2455 5758 2459 5762
rect 2515 5758 2519 5762
rect 2534 5758 2538 5762
rect 2552 5763 2556 5767
rect 2571 5764 2575 5771
rect 2629 5764 2633 5771
rect 2587 5758 2591 5762
rect 2647 5758 2651 5762
rect 2666 5758 2670 5762
rect 2684 5763 2688 5767
rect 2703 5764 2707 5771
rect 2761 5764 2765 5771
rect 2719 5758 2723 5762
rect 2779 5758 2783 5762
rect 2797 5760 2801 5764
rect 2008 5751 2012 5755
rect 934 5735 938 5739
rect 956 5733 960 5737
rect 975 5734 979 5741
rect 1033 5734 1037 5741
rect 991 5728 995 5732
rect 1487 5740 1491 5744
rect 1525 5740 1529 5744
rect 1545 5740 1549 5744
rect 1582 5740 1586 5744
rect 1619 5740 1623 5744
rect 1657 5740 1661 5744
rect 1677 5740 1681 5744
rect 1714 5740 1718 5744
rect 1751 5740 1755 5744
rect 1789 5740 1793 5744
rect 1809 5740 1813 5744
rect 1846 5740 1850 5744
rect 1051 5728 1055 5732
rect 1069 5730 1073 5734
rect 1879 5735 1883 5739
rect 1901 5733 1905 5737
rect 1920 5734 1924 5741
rect 1978 5734 1982 5741
rect 1936 5728 1940 5732
rect 2432 5740 2436 5744
rect 2470 5740 2474 5744
rect 2490 5740 2494 5744
rect 2527 5740 2531 5744
rect 2564 5740 2568 5744
rect 2602 5740 2606 5744
rect 2622 5740 2626 5744
rect 2659 5740 2663 5744
rect 2696 5740 2700 5744
rect 2734 5740 2738 5744
rect 2754 5740 2758 5744
rect 2791 5740 2795 5744
rect 1996 5728 2000 5732
rect 2014 5730 2018 5734
rect 968 5710 972 5714
rect 1006 5710 1010 5714
rect 1026 5710 1030 5714
rect 1063 5710 1067 5714
rect 1913 5710 1917 5714
rect 1951 5710 1955 5714
rect 1971 5710 1975 5714
rect 2008 5710 2012 5714
rect 1489 5697 1493 5701
rect 1525 5697 1529 5701
rect 1545 5697 1549 5701
rect 1582 5695 1586 5699
rect 1621 5697 1625 5701
rect 1657 5697 1661 5701
rect 1677 5697 1681 5701
rect 1714 5695 1718 5699
rect 1753 5697 1757 5701
rect 1789 5697 1793 5701
rect 1809 5697 1813 5701
rect 1846 5695 1850 5699
rect 2434 5697 2438 5701
rect 2470 5697 2474 5701
rect 2490 5697 2494 5701
rect 2527 5695 2531 5699
rect 2566 5697 2570 5701
rect 2602 5697 2606 5701
rect 2622 5697 2626 5701
rect 2659 5695 2663 5699
rect 2698 5697 2702 5701
rect 2734 5697 2738 5701
rect 2754 5697 2758 5701
rect 2791 5695 2795 5699
rect 1473 5677 1477 5681
rect 1494 5678 1498 5685
rect 970 5667 974 5671
rect 1006 5667 1010 5671
rect 1026 5667 1030 5671
rect 1552 5678 1556 5685
rect 1510 5672 1514 5676
rect 1570 5672 1574 5676
rect 1589 5672 1593 5676
rect 1607 5677 1611 5681
rect 1626 5678 1630 5685
rect 1684 5678 1688 5685
rect 1642 5672 1646 5676
rect 1702 5672 1706 5676
rect 1721 5672 1725 5676
rect 1739 5677 1743 5681
rect 1758 5678 1762 5685
rect 1816 5678 1820 5685
rect 1774 5672 1778 5676
rect 1834 5672 1838 5676
rect 1852 5674 1856 5678
rect 2418 5677 2422 5681
rect 2439 5678 2443 5685
rect 1063 5665 1067 5669
rect 1915 5667 1919 5671
rect 1951 5667 1955 5671
rect 1971 5667 1975 5671
rect 2497 5678 2501 5685
rect 2455 5672 2459 5676
rect 2515 5672 2519 5676
rect 2534 5672 2538 5676
rect 2552 5677 2556 5681
rect 2571 5678 2575 5685
rect 2629 5678 2633 5685
rect 2587 5672 2591 5676
rect 2647 5672 2651 5676
rect 2666 5672 2670 5676
rect 2684 5677 2688 5681
rect 2703 5678 2707 5685
rect 2761 5678 2765 5685
rect 2719 5672 2723 5676
rect 2779 5672 2783 5676
rect 2797 5674 2801 5678
rect 2008 5665 2012 5669
rect 956 5647 960 5651
rect 975 5648 979 5655
rect 1033 5648 1037 5655
rect 991 5642 995 5646
rect 1487 5654 1491 5658
rect 1525 5654 1529 5658
rect 1545 5654 1549 5658
rect 1582 5654 1586 5658
rect 1619 5654 1623 5658
rect 1657 5654 1661 5658
rect 1677 5654 1681 5658
rect 1714 5654 1718 5658
rect 1751 5654 1755 5658
rect 1789 5654 1793 5658
rect 1809 5654 1813 5658
rect 1846 5654 1850 5658
rect 1051 5642 1055 5646
rect 1069 5644 1073 5648
rect 1901 5647 1905 5651
rect 1920 5648 1924 5655
rect 1978 5648 1982 5655
rect 1936 5642 1940 5646
rect 2432 5654 2436 5658
rect 2470 5654 2474 5658
rect 2490 5654 2494 5658
rect 2527 5654 2531 5658
rect 2564 5654 2568 5658
rect 2602 5654 2606 5658
rect 2622 5654 2626 5658
rect 2659 5654 2663 5658
rect 2696 5654 2700 5658
rect 2734 5654 2738 5658
rect 2754 5654 2758 5658
rect 2791 5654 2795 5658
rect 1996 5642 2000 5646
rect 2014 5644 2018 5648
rect 1713 5633 1717 5637
rect 1737 5633 1741 5637
rect 2658 5633 2662 5637
rect 2682 5633 2686 5637
rect 968 5624 972 5628
rect 1006 5624 1010 5628
rect 1026 5624 1030 5628
rect 1063 5624 1067 5628
rect 1913 5624 1917 5628
rect 1951 5624 1955 5628
rect 1971 5624 1975 5628
rect 2008 5624 2012 5628
rect 1702 5618 1706 5622
rect 2647 5618 2651 5622
rect 1717 5610 1721 5614
rect 2662 5610 2666 5614
rect 1110 5596 1114 5600
rect 946 5589 950 5593
rect 969 5561 973 5565
rect 1014 5561 1018 5565
rect 1041 5561 1045 5565
rect 1085 5561 1089 5565
rect 2053 5596 2057 5600
rect 1891 5589 1895 5593
rect 1713 5583 1717 5587
rect 1737 5583 1741 5587
rect 1159 5568 1163 5572
rect 1230 5561 1234 5565
rect 1275 5561 1279 5565
rect 1302 5561 1306 5565
rect 1346 5561 1350 5565
rect 1914 5561 1918 5565
rect 1959 5561 1963 5565
rect 1986 5561 1990 5565
rect 2030 5561 2034 5565
rect 955 5541 959 5545
rect 982 5541 986 5545
rect 998 5542 1002 5546
rect 1054 5541 1058 5545
rect 1073 5542 1077 5546
rect 1130 5541 1134 5545
rect 1166 5548 1172 5552
rect 1489 5555 1493 5559
rect 1525 5555 1529 5559
rect 1545 5555 1549 5559
rect 1582 5553 1586 5557
rect 1621 5555 1625 5559
rect 1657 5555 1661 5559
rect 1677 5555 1681 5559
rect 1714 5553 1718 5557
rect 1753 5555 1757 5559
rect 1789 5555 1793 5559
rect 1809 5555 1813 5559
rect 2658 5583 2662 5587
rect 2682 5583 2686 5587
rect 2104 5568 2108 5572
rect 1846 5553 1850 5557
rect 2175 5561 2179 5565
rect 2220 5561 2224 5565
rect 2247 5561 2251 5565
rect 2291 5561 2295 5565
rect 1216 5541 1220 5545
rect 1243 5541 1247 5545
rect 1259 5542 1263 5546
rect 1315 5541 1319 5545
rect 1334 5542 1338 5546
rect 1366 5541 1370 5545
rect 1157 5532 1161 5536
rect 1473 5535 1477 5539
rect 1494 5536 1498 5543
rect 972 5523 976 5527
rect 1018 5524 1023 5528
rect 1044 5523 1048 5527
rect 1088 5524 1092 5528
rect 1233 5523 1237 5527
rect 1279 5524 1284 5528
rect 1305 5523 1309 5527
rect 1349 5524 1353 5528
rect 1552 5536 1556 5543
rect 1510 5530 1514 5534
rect 1570 5530 1574 5534
rect 1589 5530 1593 5534
rect 1607 5535 1611 5539
rect 1626 5536 1630 5543
rect 1684 5536 1688 5543
rect 1642 5530 1646 5534
rect 1702 5530 1706 5534
rect 1721 5530 1725 5534
rect 1739 5535 1743 5539
rect 1758 5536 1762 5543
rect 1816 5536 1820 5543
rect 1774 5530 1778 5534
rect 1900 5541 1904 5545
rect 1927 5541 1931 5545
rect 1943 5542 1947 5546
rect 1999 5541 2003 5545
rect 2018 5542 2022 5546
rect 2075 5541 2079 5545
rect 2111 5548 2117 5552
rect 2434 5555 2438 5559
rect 2470 5555 2474 5559
rect 2490 5555 2494 5559
rect 2527 5553 2531 5557
rect 2566 5555 2570 5559
rect 2602 5555 2606 5559
rect 2622 5555 2626 5559
rect 2659 5553 2663 5557
rect 2698 5555 2702 5559
rect 2734 5555 2738 5559
rect 2754 5555 2758 5559
rect 2791 5553 2795 5557
rect 2161 5541 2165 5545
rect 2188 5541 2192 5545
rect 2204 5542 2208 5546
rect 2260 5541 2264 5545
rect 2279 5542 2283 5546
rect 2311 5541 2315 5545
rect 1834 5530 1838 5534
rect 1852 5532 1856 5536
rect 2102 5532 2106 5536
rect 2418 5535 2422 5539
rect 2439 5536 2443 5543
rect 1917 5523 1921 5527
rect 1963 5524 1968 5528
rect 1989 5523 1993 5527
rect 2033 5524 2037 5528
rect 2178 5523 2182 5527
rect 2224 5524 2229 5528
rect 2250 5523 2254 5527
rect 2294 5524 2298 5528
rect 2497 5536 2501 5543
rect 2455 5530 2459 5534
rect 2515 5530 2519 5534
rect 2534 5530 2538 5534
rect 2552 5535 2556 5539
rect 2571 5536 2575 5543
rect 2629 5536 2633 5543
rect 2587 5530 2591 5534
rect 2647 5530 2651 5534
rect 2666 5530 2670 5534
rect 2684 5535 2688 5539
rect 2703 5536 2707 5543
rect 2761 5536 2765 5543
rect 2719 5530 2723 5534
rect 2779 5530 2783 5534
rect 2797 5532 2801 5536
rect 1487 5512 1491 5516
rect 1525 5512 1529 5516
rect 1545 5512 1549 5516
rect 1582 5512 1586 5516
rect 1619 5512 1623 5516
rect 1657 5512 1661 5516
rect 1677 5512 1681 5516
rect 1714 5512 1718 5516
rect 1751 5512 1755 5516
rect 1789 5512 1793 5516
rect 1809 5512 1813 5516
rect 1846 5512 1850 5516
rect 2432 5512 2436 5516
rect 2470 5512 2474 5516
rect 2490 5512 2494 5516
rect 2527 5512 2531 5516
rect 2564 5512 2568 5516
rect 2602 5512 2606 5516
rect 2622 5512 2626 5516
rect 2659 5512 2663 5516
rect 2696 5512 2700 5516
rect 2734 5512 2738 5516
rect 2754 5512 2758 5516
rect 2791 5512 2795 5516
rect 1233 5495 1237 5499
rect 1279 5494 1284 5498
rect 1305 5495 1309 5499
rect 1349 5494 1353 5498
rect 2178 5495 2182 5499
rect 2224 5494 2229 5498
rect 2250 5495 2254 5499
rect 2294 5494 2298 5498
rect 1159 5486 1163 5490
rect 1138 5472 1142 5476
rect 1216 5477 1220 5481
rect 1243 5477 1247 5481
rect 1259 5476 1263 5480
rect 1315 5477 1319 5481
rect 1334 5476 1338 5480
rect 2104 5486 2108 5490
rect 1366 5477 1370 5481
rect 1165 5468 1169 5472
rect 1230 5457 1234 5461
rect 1275 5457 1279 5461
rect 1302 5457 1306 5461
rect 1346 5457 1350 5461
rect 1157 5450 1161 5454
rect 1768 5461 1772 5465
rect 2083 5472 2087 5476
rect 2161 5477 2165 5481
rect 2188 5477 2192 5481
rect 2204 5476 2208 5480
rect 2260 5477 2264 5481
rect 2279 5476 2283 5480
rect 2311 5477 2315 5481
rect 2110 5468 2114 5472
rect 2175 5457 2179 5461
rect 2220 5457 2224 5461
rect 2247 5457 2251 5461
rect 2291 5457 2295 5461
rect 2102 5450 2106 5454
rect 1775 5441 1781 5445
rect 988 5432 992 5436
rect 1078 5432 1082 5436
rect 1159 5432 1163 5436
rect 1230 5429 1234 5433
rect 1275 5429 1279 5433
rect 1302 5429 1306 5433
rect 1346 5429 1350 5433
rect 1933 5432 1937 5436
rect 2023 5432 2027 5436
rect 2104 5432 2108 5436
rect 995 5412 1001 5416
rect 1085 5412 1091 5416
rect 1766 5425 1770 5429
rect 2175 5429 2179 5433
rect 2220 5429 2224 5433
rect 2247 5429 2251 5433
rect 2291 5429 2295 5433
rect 1166 5412 1172 5416
rect 1216 5409 1220 5413
rect 1243 5409 1247 5413
rect 1259 5410 1263 5414
rect 1315 5409 1319 5413
rect 1334 5410 1338 5414
rect 1366 5409 1370 5413
rect 986 5396 990 5400
rect 1076 5396 1080 5400
rect 1157 5396 1161 5400
rect 1233 5391 1237 5395
rect 1279 5392 1284 5396
rect 1940 5412 1946 5416
rect 2030 5412 2036 5416
rect 2111 5412 2117 5416
rect 2161 5409 2165 5413
rect 2188 5409 2192 5413
rect 2204 5410 2208 5414
rect 2260 5409 2264 5413
rect 2279 5410 2283 5414
rect 2311 5409 2315 5413
rect 1305 5391 1309 5395
rect 1349 5392 1353 5396
rect 1931 5396 1935 5400
rect 2021 5396 2025 5400
rect 2102 5396 2106 5400
rect 2178 5391 2182 5395
rect 2224 5392 2229 5396
rect 1654 5387 1658 5391
rect 1707 5387 1711 5391
rect 2250 5391 2254 5395
rect 2294 5392 2298 5396
rect 1768 5381 1772 5385
rect 1233 5363 1237 5367
rect 1279 5362 1284 5366
rect 1305 5363 1309 5367
rect 1349 5362 1353 5366
rect 988 5354 992 5358
rect 1078 5354 1082 5358
rect 1159 5354 1163 5358
rect 967 5340 971 5344
rect 994 5336 998 5340
rect 1021 5332 1025 5336
rect 1057 5340 1061 5344
rect 1084 5336 1088 5340
rect 986 5318 990 5322
rect 1111 5332 1115 5336
rect 1138 5340 1142 5344
rect 1216 5345 1220 5349
rect 1243 5345 1247 5349
rect 1259 5344 1263 5348
rect 1315 5345 1319 5349
rect 1334 5344 1338 5348
rect 1747 5367 1751 5371
rect 1774 5363 1778 5367
rect 1366 5345 1370 5349
rect 1801 5359 1805 5363
rect 2178 5363 2182 5367
rect 1823 5359 1827 5363
rect 2224 5362 2229 5366
rect 2250 5363 2254 5367
rect 2294 5362 2298 5366
rect 1766 5345 1770 5349
rect 1933 5354 1937 5358
rect 2023 5354 2027 5358
rect 2104 5354 2108 5358
rect 1165 5336 1169 5340
rect 1076 5318 1080 5322
rect 1768 5331 1772 5335
rect 1230 5325 1234 5329
rect 1275 5325 1279 5329
rect 1302 5325 1306 5329
rect 1346 5325 1350 5329
rect 1912 5340 1916 5344
rect 1939 5336 1943 5340
rect 1157 5318 1161 5322
rect 1966 5332 1970 5336
rect 2002 5340 2006 5344
rect 2029 5336 2033 5340
rect 1931 5318 1935 5322
rect 2056 5332 2060 5336
rect 2083 5340 2087 5344
rect 2161 5345 2165 5349
rect 2188 5345 2192 5349
rect 2204 5344 2208 5348
rect 2260 5345 2264 5349
rect 2279 5344 2283 5348
rect 2311 5345 2315 5349
rect 2110 5336 2114 5340
rect 2021 5318 2025 5322
rect 2175 5325 2179 5329
rect 2220 5325 2224 5329
rect 2247 5325 2251 5329
rect 2291 5325 2295 5329
rect 2102 5318 2106 5322
rect 1775 5311 1781 5315
rect 1054 5297 1058 5301
rect 1159 5297 1163 5301
rect 1230 5297 1234 5301
rect 1275 5297 1279 5301
rect 1302 5297 1306 5301
rect 1346 5297 1350 5301
rect 1766 5295 1770 5299
rect 1999 5297 2003 5301
rect 2104 5297 2108 5301
rect 2175 5297 2179 5301
rect 2220 5297 2224 5301
rect 2247 5297 2251 5301
rect 2291 5297 2295 5301
rect 1061 5277 1067 5281
rect 1166 5277 1172 5281
rect 1216 5277 1220 5281
rect 1243 5277 1247 5281
rect 1259 5278 1263 5282
rect 1315 5277 1319 5281
rect 1334 5278 1338 5282
rect 1366 5277 1370 5281
rect 2006 5277 2012 5281
rect 2111 5277 2117 5281
rect 2161 5277 2165 5281
rect 2188 5277 2192 5281
rect 2204 5278 2208 5282
rect 2260 5277 2264 5281
rect 2279 5278 2283 5282
rect 2311 5277 2315 5281
rect 1052 5261 1056 5265
rect 1157 5261 1161 5265
rect 1233 5259 1237 5263
rect 1279 5260 1284 5264
rect 1305 5259 1309 5263
rect 1349 5260 1353 5264
rect 1997 5261 2001 5265
rect 2102 5261 2106 5265
rect 1560 5257 1564 5261
rect 1613 5257 1617 5261
rect 2178 5259 2182 5263
rect 2224 5260 2229 5264
rect 2250 5259 2254 5263
rect 2294 5260 2298 5264
rect 1768 5251 1772 5255
rect 1233 5231 1237 5235
rect 1279 5230 1284 5234
rect 1305 5231 1309 5235
rect 1349 5230 1353 5234
rect 1054 5222 1058 5226
rect 1159 5222 1163 5226
rect 1033 5208 1037 5212
rect 1060 5204 1064 5208
rect 1087 5200 1091 5204
rect 1138 5208 1142 5212
rect 1216 5213 1220 5217
rect 1243 5213 1247 5217
rect 1259 5212 1263 5216
rect 1315 5213 1319 5217
rect 1334 5212 1338 5216
rect 1747 5237 1751 5241
rect 1774 5233 1778 5237
rect 1366 5213 1370 5217
rect 1801 5229 1805 5233
rect 2178 5231 2182 5235
rect 2224 5230 2229 5234
rect 2250 5231 2254 5235
rect 2294 5230 2298 5234
rect 1766 5215 1770 5219
rect 1999 5222 2003 5226
rect 2104 5222 2108 5226
rect 1165 5204 1169 5208
rect 1052 5186 1056 5190
rect 1230 5193 1234 5197
rect 1275 5193 1279 5197
rect 1302 5193 1306 5197
rect 1346 5193 1350 5197
rect 1978 5208 1982 5212
rect 2005 5204 2009 5208
rect 1157 5186 1161 5190
rect 2032 5200 2036 5204
rect 2083 5208 2087 5212
rect 2161 5213 2165 5217
rect 2188 5213 2192 5217
rect 2204 5212 2208 5216
rect 2260 5213 2264 5217
rect 2279 5212 2283 5216
rect 2311 5213 2315 5217
rect 2110 5204 2114 5208
rect 1997 5186 2001 5190
rect 2175 5193 2179 5197
rect 2220 5193 2224 5197
rect 2247 5193 2251 5197
rect 2291 5193 2295 5197
rect 2102 5186 2106 5190
rect 1078 5166 1082 5170
rect 1159 5166 1163 5170
rect 1230 5165 1234 5169
rect 1275 5165 1279 5169
rect 1302 5165 1306 5169
rect 1346 5165 1350 5169
rect 2023 5166 2027 5170
rect 2104 5166 2108 5170
rect 2175 5165 2179 5169
rect 2220 5165 2224 5169
rect 2247 5165 2251 5169
rect 2291 5165 2295 5169
rect 1085 5146 1091 5150
rect 1166 5146 1172 5150
rect 1216 5145 1220 5149
rect 1243 5145 1247 5149
rect 1259 5146 1263 5150
rect 1315 5145 1319 5149
rect 1334 5146 1338 5150
rect 1619 5153 1623 5157
rect 1656 5155 1660 5159
rect 1676 5155 1680 5159
rect 1712 5155 1716 5159
rect 1366 5145 1370 5149
rect 1076 5130 1080 5134
rect 1157 5130 1161 5134
rect 1233 5127 1237 5131
rect 1279 5128 1284 5132
rect 1613 5132 1617 5136
rect 1305 5127 1309 5131
rect 1349 5128 1353 5132
rect 1631 5130 1635 5134
rect 1649 5136 1653 5143
rect 1707 5136 1711 5143
rect 1691 5130 1695 5134
rect 1726 5135 1730 5139
rect 2030 5146 2036 5150
rect 2111 5146 2117 5150
rect 2161 5145 2165 5149
rect 2188 5145 2192 5149
rect 2204 5146 2208 5150
rect 2260 5145 2264 5149
rect 2279 5146 2283 5150
rect 2564 5153 2568 5157
rect 2601 5155 2605 5159
rect 2621 5155 2625 5159
rect 2657 5155 2661 5159
rect 2311 5145 2315 5149
rect 2021 5130 2025 5134
rect 2102 5130 2106 5134
rect 2178 5127 2182 5131
rect 2224 5128 2229 5132
rect 2558 5132 2562 5136
rect 2250 5127 2254 5131
rect 2294 5128 2298 5132
rect 2576 5130 2580 5134
rect 2594 5136 2598 5143
rect 2652 5136 2656 5143
rect 2636 5130 2640 5134
rect 2671 5135 2675 5139
rect 1619 5112 1623 5116
rect 1656 5112 1660 5116
rect 1676 5112 1680 5116
rect 1714 5112 1718 5116
rect 2564 5112 2568 5116
rect 2601 5112 2605 5116
rect 2621 5112 2625 5116
rect 2659 5112 2663 5116
rect 1233 5099 1237 5103
rect 1279 5098 1284 5102
rect 1305 5099 1309 5103
rect 1349 5098 1353 5102
rect 2178 5099 2182 5103
rect 2224 5098 2229 5102
rect 2250 5099 2254 5103
rect 2294 5098 2298 5102
rect 1078 5090 1082 5094
rect 1159 5090 1163 5094
rect 1057 5076 1061 5080
rect 1084 5072 1088 5076
rect 1111 5068 1115 5072
rect 1138 5076 1142 5080
rect 1165 5072 1169 5076
rect 1076 5054 1080 5058
rect 1216 5081 1220 5085
rect 1243 5081 1247 5085
rect 1259 5080 1263 5084
rect 1315 5081 1319 5085
rect 1334 5080 1338 5084
rect 2023 5090 2027 5094
rect 1366 5081 1370 5085
rect 1713 5083 1717 5087
rect 2104 5090 2108 5094
rect 1192 5068 1196 5072
rect 1596 5074 1600 5078
rect 1157 5054 1161 5058
rect 1230 5061 1234 5065
rect 1275 5061 1279 5065
rect 1302 5061 1306 5065
rect 1346 5061 1350 5065
rect 2002 5076 2006 5080
rect 2029 5072 2033 5076
rect 1621 5053 1625 5057
rect 1657 5053 1661 5057
rect 1677 5053 1681 5057
rect 2056 5068 2060 5072
rect 2083 5076 2087 5080
rect 2110 5072 2114 5076
rect 1714 5051 1718 5055
rect 2021 5054 2025 5058
rect 2161 5081 2165 5085
rect 2188 5081 2192 5085
rect 2204 5080 2208 5084
rect 2260 5081 2264 5085
rect 2279 5080 2283 5084
rect 2311 5081 2315 5085
rect 2658 5083 2662 5087
rect 2137 5068 2141 5072
rect 2541 5074 2545 5078
rect 2102 5054 2106 5058
rect 2175 5061 2179 5065
rect 2220 5061 2224 5065
rect 2247 5061 2251 5065
rect 2291 5061 2295 5065
rect 2566 5053 2570 5057
rect 2602 5053 2606 5057
rect 2622 5053 2626 5057
rect 2659 5051 2663 5055
rect 1607 5033 1611 5037
rect 1626 5034 1630 5041
rect 1684 5034 1688 5041
rect 1642 5028 1646 5032
rect 1702 5028 1706 5032
rect 1720 5030 1724 5034
rect 2552 5033 2556 5037
rect 2571 5034 2575 5041
rect 2629 5034 2633 5041
rect 2587 5028 2591 5032
rect 2647 5028 2651 5032
rect 2665 5030 2669 5034
rect 873 5020 877 5024
rect 909 5020 913 5024
rect 929 5020 933 5024
rect 966 5018 970 5022
rect 1005 5020 1009 5024
rect 1041 5020 1045 5024
rect 1061 5020 1065 5024
rect 1098 5018 1102 5022
rect 1137 5020 1141 5024
rect 1173 5020 1177 5024
rect 1193 5020 1197 5024
rect 1230 5018 1234 5022
rect 1269 5020 1273 5024
rect 1305 5020 1309 5024
rect 1325 5020 1329 5024
rect 1362 5018 1366 5022
rect 1818 5020 1822 5024
rect 1854 5020 1858 5024
rect 1874 5020 1878 5024
rect 1911 5018 1915 5022
rect 1950 5020 1954 5024
rect 1986 5020 1990 5024
rect 2006 5020 2010 5024
rect 2043 5018 2047 5022
rect 2082 5020 2086 5024
rect 2118 5020 2122 5024
rect 2138 5020 2142 5024
rect 2175 5018 2179 5022
rect 2214 5020 2218 5024
rect 2250 5020 2254 5024
rect 2270 5020 2274 5024
rect 2307 5018 2311 5022
rect 857 5000 861 5004
rect 878 5001 882 5008
rect 936 5001 940 5008
rect 894 4995 898 4999
rect 954 4995 958 4999
rect 972 4997 976 5001
rect 989 5000 993 5004
rect 1010 5001 1014 5008
rect 1068 5001 1072 5008
rect 1026 4995 1030 4999
rect 1086 4995 1090 4999
rect 1104 4997 1108 5001
rect 1121 5000 1125 5004
rect 1142 5001 1146 5008
rect 1200 5001 1204 5008
rect 1158 4995 1162 4999
rect 1218 4995 1222 4999
rect 1236 4997 1240 5001
rect 1253 5000 1257 5004
rect 1274 5001 1278 5008
rect 1332 5001 1336 5008
rect 1290 4995 1294 4999
rect 1619 5010 1623 5014
rect 1657 5010 1661 5014
rect 1677 5010 1681 5014
rect 1714 5010 1718 5014
rect 1350 4995 1354 4999
rect 1368 4997 1372 5001
rect 1802 5000 1806 5004
rect 1823 5001 1827 5008
rect 1881 5001 1885 5008
rect 1839 4995 1843 4999
rect 1899 4995 1903 4999
rect 1917 4997 1921 5001
rect 1934 5000 1938 5004
rect 1955 5001 1959 5008
rect 2013 5001 2017 5008
rect 1971 4995 1975 4999
rect 2031 4995 2035 4999
rect 2049 4997 2053 5001
rect 2066 5000 2070 5004
rect 2087 5001 2091 5008
rect 2145 5001 2149 5008
rect 2103 4995 2107 4999
rect 2163 4995 2167 4999
rect 2181 4997 2185 5001
rect 2198 5000 2202 5004
rect 2219 5001 2223 5008
rect 2277 5001 2281 5008
rect 2235 4995 2239 4999
rect 2564 5010 2568 5014
rect 2602 5010 2606 5014
rect 2622 5010 2626 5014
rect 2659 5010 2663 5014
rect 2295 4995 2299 4999
rect 2313 4997 2317 5001
rect 871 4977 875 4981
rect 909 4977 913 4981
rect 929 4977 933 4981
rect 966 4977 970 4981
rect 1003 4977 1007 4981
rect 1041 4977 1045 4981
rect 1061 4977 1065 4981
rect 1098 4977 1102 4981
rect 1135 4977 1139 4981
rect 1173 4977 1177 4981
rect 1193 4977 1197 4981
rect 1230 4977 1234 4981
rect 1267 4977 1271 4981
rect 1305 4977 1309 4981
rect 1325 4977 1329 4981
rect 1362 4977 1366 4981
rect 1816 4977 1820 4981
rect 1854 4977 1858 4981
rect 1874 4977 1878 4981
rect 1911 4977 1915 4981
rect 1948 4977 1952 4981
rect 1986 4977 1990 4981
rect 2006 4977 2010 4981
rect 2043 4977 2047 4981
rect 2080 4977 2084 4981
rect 2118 4977 2122 4981
rect 2138 4977 2142 4981
rect 2175 4977 2179 4981
rect 2212 4977 2216 4981
rect 2250 4977 2254 4981
rect 2270 4977 2274 4981
rect 2307 4977 2311 4981
rect 4572 7954 4576 7960
rect 4593 7959 4597 7965
rect 4635 7950 4639 7963
rect 4678 7952 4682 7965
rect 4711 7954 4717 7963
rect 4601 7352 4605 7358
rect 4620 7359 4624 7368
rect 4667 7353 4676 7374
rect 4745 7353 4754 7374
rect 1190 4502 1196 4506
rect 2117 4502 2123 4506
rect 2426 4502 2432 4506
rect 2735 4502 2741 4506
rect 3044 4502 3050 4506
rect 3353 4502 3359 4506
rect 1197 4483 1206 4487
rect 2124 4483 2133 4487
rect 2433 4483 2442 4487
rect 2742 4483 2751 4487
rect 3051 4483 3060 4487
rect 3360 4483 3369 4487
rect 1191 4431 1212 4440
rect 1191 4353 1212 4362
rect 2118 4431 2139 4440
rect 2118 4353 2139 4362
rect 2427 4431 2448 4440
rect 2427 4353 2448 4362
rect 2736 4431 2757 4440
rect 2736 4353 2757 4362
rect 3045 4431 3066 4440
rect 3045 4353 3066 4362
rect 3354 4431 3375 4440
rect 3354 4353 3375 4362
<< metal1 >>
rect 1060 10290 1320 10293
rect 118 9786 1024 10280
rect 1060 10036 1063 10290
rect 1317 10036 1320 10290
rect 1060 10033 1320 10036
rect 1369 10290 1629 10293
rect 1369 10036 1372 10290
rect 1462 10138 1546 10223
rect 1626 10036 1629 10290
rect 1369 10033 1629 10036
rect 1678 10290 1938 10293
rect 1678 10036 1681 10290
rect 1765 10113 1843 10202
rect 1935 10036 1938 10290
rect 1678 10033 1938 10036
rect 1987 10290 2247 10293
rect 1987 10036 1990 10290
rect 2072 10118 2150 10207
rect 2244 10036 2247 10290
rect 1987 10033 2247 10036
rect 2296 10290 2556 10293
rect 2296 10036 2299 10290
rect 2389 10118 2467 10207
rect 2553 10036 2556 10290
rect 2296 10033 2556 10036
rect 2605 10290 2865 10293
rect 2605 10036 2608 10290
rect 2700 10120 2778 10209
rect 2862 10036 2865 10290
rect 2605 10033 2865 10036
rect 2914 10290 3174 10293
rect 2914 10036 2917 10290
rect 3004 10110 3082 10199
rect 3171 10036 3174 10290
rect 2914 10033 3174 10036
rect 3223 10290 3483 10293
rect 3223 10036 3226 10290
rect 3318 10118 3396 10207
rect 3480 10036 3483 10290
rect 3223 10033 3483 10036
rect 3532 10290 3792 10293
rect 3532 10036 3535 10290
rect 3608 10103 3720 10217
rect 3789 10036 3792 10290
rect 3532 10033 3792 10036
rect 3841 10290 4101 10293
rect 3841 10036 3844 10290
rect 4098 10036 4101 10290
rect 3841 10033 4101 10036
rect 1102 10023 1278 10033
rect 1411 10023 1587 10033
rect 1720 10023 1896 10033
rect 2029 10023 2205 10033
rect 2338 10023 2514 10033
rect 2647 10023 2823 10033
rect 2956 10023 3132 10033
rect 3265 10023 3441 10033
rect 3574 10023 3750 10033
rect 3883 10023 4059 10033
rect 1112 10013 1268 10023
rect 1421 10013 1577 10023
rect 1730 10013 1886 10023
rect 2039 10013 2195 10023
rect 2348 10013 2504 10023
rect 2657 10013 2813 10023
rect 2966 10013 3122 10023
rect 3275 10013 3431 10023
rect 3584 10013 3740 10023
rect 3893 10013 4049 10023
rect 1122 10003 1258 10013
rect 1431 10003 1567 10013
rect 1740 10003 1876 10013
rect 2049 10003 2185 10013
rect 2358 10003 2494 10013
rect 2667 10003 2803 10013
rect 2976 10003 3112 10013
rect 3285 10003 3421 10013
rect 3594 10003 3730 10013
rect 3903 10003 4039 10013
rect 1132 9993 1248 10003
rect 1441 10001 1557 10003
rect 1441 9997 1454 10001
rect 1458 9997 1461 10001
rect 1465 9997 1468 10001
rect 1472 9997 1475 10001
rect 1479 9997 1482 10001
rect 1486 9997 1489 10001
rect 1493 9997 1496 10001
rect 1500 9997 1503 10001
rect 1507 9997 1510 10001
rect 1514 9997 1517 10001
rect 1521 9997 1524 10001
rect 1528 9997 1531 10001
rect 1535 9997 1538 10001
rect 1542 9997 1557 10001
rect 1441 9996 1557 9997
rect 1441 9993 1454 9996
rect 118 9348 593 9786
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 802 9761 821 9762
rect 806 9757 807 9761
rect 811 9757 812 9761
rect 816 9757 817 9761
rect 802 9756 821 9757
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 802 9751 821 9752
rect 806 9747 807 9751
rect 811 9747 812 9751
rect 816 9747 817 9751
rect 802 9746 821 9747
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 802 9741 821 9742
rect 806 9737 807 9741
rect 811 9737 812 9741
rect 816 9737 817 9741
rect 802 9736 821 9737
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 831 9761 850 9762
rect 835 9757 836 9761
rect 840 9757 841 9761
rect 845 9757 846 9761
rect 831 9756 850 9757
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 831 9751 850 9752
rect 835 9747 836 9751
rect 840 9747 841 9751
rect 845 9747 846 9751
rect 831 9746 850 9747
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 831 9741 850 9742
rect 835 9737 836 9741
rect 840 9737 841 9741
rect 845 9737 846 9741
rect 831 9736 850 9737
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 860 9761 879 9762
rect 864 9757 865 9761
rect 869 9757 870 9761
rect 874 9757 875 9761
rect 860 9756 879 9757
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 860 9751 879 9752
rect 864 9747 865 9751
rect 869 9747 870 9751
rect 874 9747 875 9751
rect 860 9746 879 9747
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 860 9741 879 9742
rect 864 9737 865 9741
rect 869 9737 870 9741
rect 874 9737 875 9741
rect 860 9736 879 9737
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 889 9761 908 9762
rect 893 9757 894 9761
rect 898 9757 899 9761
rect 903 9757 904 9761
rect 889 9756 908 9757
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 889 9751 908 9752
rect 893 9747 894 9751
rect 898 9747 899 9751
rect 903 9747 904 9751
rect 889 9746 908 9747
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 889 9741 908 9742
rect 893 9737 894 9741
rect 898 9737 899 9741
rect 903 9737 904 9741
rect 889 9736 908 9737
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 918 9761 937 9762
rect 922 9757 923 9761
rect 927 9757 928 9761
rect 932 9757 933 9761
rect 918 9756 937 9757
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 918 9751 937 9752
rect 922 9747 923 9751
rect 927 9747 928 9751
rect 932 9747 933 9751
rect 918 9746 937 9747
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 918 9741 937 9742
rect 922 9737 923 9741
rect 927 9737 928 9741
rect 932 9737 933 9741
rect 918 9736 937 9737
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 802 9715 821 9716
rect 806 9711 807 9715
rect 811 9711 812 9715
rect 816 9711 817 9715
rect 802 9710 821 9711
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 802 9705 821 9706
rect 806 9701 807 9705
rect 811 9701 812 9705
rect 816 9701 817 9705
rect 802 9700 821 9701
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 802 9695 821 9696
rect 806 9691 807 9695
rect 811 9691 812 9695
rect 816 9691 817 9695
rect 802 9690 821 9691
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 831 9715 850 9716
rect 835 9711 836 9715
rect 840 9711 841 9715
rect 845 9711 846 9715
rect 831 9710 850 9711
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 831 9705 850 9706
rect 835 9701 836 9705
rect 840 9701 841 9705
rect 845 9701 846 9705
rect 831 9700 850 9701
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 831 9695 850 9696
rect 835 9691 836 9695
rect 840 9691 841 9695
rect 845 9691 846 9695
rect 831 9690 850 9691
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 860 9715 879 9716
rect 864 9711 865 9715
rect 869 9711 870 9715
rect 874 9711 875 9715
rect 860 9710 879 9711
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 860 9705 879 9706
rect 864 9701 865 9705
rect 869 9701 870 9705
rect 874 9701 875 9705
rect 860 9700 879 9701
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 860 9695 879 9696
rect 864 9691 865 9695
rect 869 9691 870 9695
rect 874 9691 875 9695
rect 860 9690 879 9691
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 889 9715 908 9716
rect 893 9711 894 9715
rect 898 9711 899 9715
rect 903 9711 904 9715
rect 889 9710 908 9711
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 889 9705 908 9706
rect 893 9701 894 9705
rect 898 9701 899 9705
rect 903 9701 904 9705
rect 889 9700 908 9701
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 889 9695 908 9696
rect 893 9691 894 9695
rect 898 9691 899 9695
rect 903 9691 904 9695
rect 889 9690 908 9691
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 918 9715 937 9716
rect 922 9711 923 9715
rect 927 9711 928 9715
rect 932 9711 933 9715
rect 918 9710 937 9711
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 918 9705 937 9706
rect 922 9701 923 9705
rect 927 9701 928 9705
rect 932 9701 933 9705
rect 918 9700 937 9701
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 918 9695 937 9696
rect 922 9691 923 9695
rect 927 9691 928 9695
rect 932 9691 933 9695
rect 918 9690 937 9691
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 617 9618 618 9622
rect 622 9618 623 9622
rect 627 9618 628 9622
rect 632 9618 633 9622
rect 637 9618 638 9622
rect 642 9618 643 9622
rect 613 9617 647 9618
rect 617 9613 618 9617
rect 622 9613 623 9617
rect 627 9613 628 9617
rect 632 9613 633 9617
rect 637 9613 638 9617
rect 642 9613 643 9617
rect 613 9612 647 9613
rect 617 9608 618 9612
rect 622 9608 623 9612
rect 627 9608 628 9612
rect 632 9608 633 9612
rect 637 9608 638 9612
rect 642 9608 643 9612
rect 613 9607 647 9608
rect 617 9603 618 9607
rect 622 9603 623 9607
rect 627 9603 628 9607
rect 632 9603 633 9607
rect 637 9603 638 9607
rect 642 9603 643 9607
rect 663 9618 664 9622
rect 668 9618 669 9622
rect 673 9618 674 9622
rect 678 9618 679 9622
rect 683 9618 684 9622
rect 688 9618 689 9622
rect 659 9617 693 9618
rect 663 9613 664 9617
rect 668 9613 669 9617
rect 673 9613 674 9617
rect 678 9613 679 9617
rect 683 9613 684 9617
rect 688 9613 689 9617
rect 659 9612 693 9613
rect 663 9608 664 9612
rect 668 9608 669 9612
rect 673 9608 674 9612
rect 678 9608 679 9612
rect 683 9608 684 9612
rect 688 9608 689 9612
rect 1142 9610 1238 9993
rect 1451 9992 1454 9993
rect 1458 9992 1461 9996
rect 1465 9992 1468 9996
rect 1472 9992 1475 9996
rect 1479 9992 1482 9996
rect 1486 9992 1489 9996
rect 1493 9992 1496 9996
rect 1500 9992 1503 9996
rect 1507 9992 1510 9996
rect 1514 9992 1517 9996
rect 1521 9992 1524 9996
rect 1528 9992 1531 9996
rect 1535 9992 1538 9996
rect 1542 9993 1557 9996
rect 1750 10001 1866 10003
rect 1750 9997 1763 10001
rect 1767 9997 1770 10001
rect 1774 9997 1777 10001
rect 1781 9997 1784 10001
rect 1788 9997 1791 10001
rect 1795 9997 1798 10001
rect 1802 9997 1805 10001
rect 1809 9997 1812 10001
rect 1816 9997 1819 10001
rect 1823 9997 1826 10001
rect 1830 9997 1833 10001
rect 1837 9997 1840 10001
rect 1844 9997 1847 10001
rect 1851 9997 1866 10001
rect 1750 9996 1866 9997
rect 1750 9993 1763 9996
rect 1542 9992 1547 9993
rect 1451 9991 1547 9992
rect 1451 9987 1454 9991
rect 1458 9987 1461 9991
rect 1465 9987 1468 9991
rect 1472 9987 1475 9991
rect 1479 9987 1482 9991
rect 1486 9987 1489 9991
rect 1493 9987 1496 9991
rect 1500 9987 1503 9991
rect 1507 9987 1510 9991
rect 1514 9987 1517 9991
rect 1521 9987 1524 9991
rect 1528 9987 1531 9991
rect 1535 9987 1538 9991
rect 1542 9987 1547 9991
rect 1451 9986 1547 9987
rect 1451 9982 1454 9986
rect 1458 9982 1461 9986
rect 1465 9982 1468 9986
rect 1472 9982 1475 9986
rect 1479 9982 1482 9986
rect 1486 9982 1489 9986
rect 1493 9982 1496 9986
rect 1500 9982 1503 9986
rect 1507 9982 1510 9986
rect 1514 9982 1517 9986
rect 1521 9982 1524 9986
rect 1528 9982 1531 9986
rect 1535 9982 1538 9986
rect 1542 9982 1547 9986
rect 1451 9981 1547 9982
rect 1760 9992 1763 9993
rect 1767 9992 1770 9996
rect 1774 9992 1777 9996
rect 1781 9992 1784 9996
rect 1788 9992 1791 9996
rect 1795 9992 1798 9996
rect 1802 9992 1805 9996
rect 1809 9992 1812 9996
rect 1816 9992 1819 9996
rect 1823 9992 1826 9996
rect 1830 9992 1833 9996
rect 1837 9992 1840 9996
rect 1844 9992 1847 9996
rect 1851 9993 1866 9996
rect 2059 10001 2175 10003
rect 2059 9997 2072 10001
rect 2076 9997 2079 10001
rect 2083 9997 2086 10001
rect 2090 9997 2093 10001
rect 2097 9997 2100 10001
rect 2104 9997 2107 10001
rect 2111 9997 2114 10001
rect 2118 9997 2121 10001
rect 2125 9997 2128 10001
rect 2132 9997 2135 10001
rect 2139 9997 2142 10001
rect 2146 9997 2149 10001
rect 2153 9997 2156 10001
rect 2160 9997 2175 10001
rect 2059 9996 2175 9997
rect 2059 9993 2072 9996
rect 1851 9992 1856 9993
rect 1760 9991 1856 9992
rect 1760 9987 1763 9991
rect 1767 9987 1770 9991
rect 1774 9987 1777 9991
rect 1781 9987 1784 9991
rect 1788 9987 1791 9991
rect 1795 9987 1798 9991
rect 1802 9987 1805 9991
rect 1809 9987 1812 9991
rect 1816 9987 1819 9991
rect 1823 9987 1826 9991
rect 1830 9987 1833 9991
rect 1837 9987 1840 9991
rect 1844 9987 1847 9991
rect 1851 9987 1856 9991
rect 1760 9986 1856 9987
rect 1760 9982 1763 9986
rect 1767 9982 1770 9986
rect 1774 9982 1777 9986
rect 1781 9982 1784 9986
rect 1788 9982 1791 9986
rect 1795 9982 1798 9986
rect 1802 9982 1805 9986
rect 1809 9982 1812 9986
rect 1816 9982 1819 9986
rect 1823 9982 1826 9986
rect 1830 9982 1833 9986
rect 1837 9982 1840 9986
rect 1844 9982 1847 9986
rect 1851 9982 1856 9986
rect 1760 9981 1856 9982
rect 2069 9992 2072 9993
rect 2076 9992 2079 9996
rect 2083 9992 2086 9996
rect 2090 9992 2093 9996
rect 2097 9992 2100 9996
rect 2104 9992 2107 9996
rect 2111 9992 2114 9996
rect 2118 9992 2121 9996
rect 2125 9992 2128 9996
rect 2132 9992 2135 9996
rect 2139 9992 2142 9996
rect 2146 9992 2149 9996
rect 2153 9992 2156 9996
rect 2160 9993 2175 9996
rect 2368 10001 2484 10003
rect 2368 9997 2381 10001
rect 2385 9997 2388 10001
rect 2392 9997 2395 10001
rect 2399 9997 2402 10001
rect 2406 9997 2409 10001
rect 2413 9997 2416 10001
rect 2420 9997 2423 10001
rect 2427 9997 2430 10001
rect 2434 9997 2437 10001
rect 2441 9997 2444 10001
rect 2448 9997 2451 10001
rect 2455 9997 2458 10001
rect 2462 9997 2465 10001
rect 2469 9997 2484 10001
rect 2368 9996 2484 9997
rect 2368 9993 2381 9996
rect 2160 9992 2165 9993
rect 2069 9991 2165 9992
rect 2069 9987 2072 9991
rect 2076 9987 2079 9991
rect 2083 9987 2086 9991
rect 2090 9987 2093 9991
rect 2097 9987 2100 9991
rect 2104 9987 2107 9991
rect 2111 9987 2114 9991
rect 2118 9987 2121 9991
rect 2125 9987 2128 9991
rect 2132 9987 2135 9991
rect 2139 9987 2142 9991
rect 2146 9987 2149 9991
rect 2153 9987 2156 9991
rect 2160 9987 2165 9991
rect 2069 9986 2165 9987
rect 2069 9982 2072 9986
rect 2076 9982 2079 9986
rect 2083 9982 2086 9986
rect 2090 9982 2093 9986
rect 2097 9982 2100 9986
rect 2104 9982 2107 9986
rect 2111 9982 2114 9986
rect 2118 9982 2121 9986
rect 2125 9982 2128 9986
rect 2132 9982 2135 9986
rect 2139 9982 2142 9986
rect 2146 9982 2149 9986
rect 2153 9982 2156 9986
rect 2160 9982 2165 9986
rect 2069 9981 2165 9982
rect 2378 9992 2381 9993
rect 2385 9992 2388 9996
rect 2392 9992 2395 9996
rect 2399 9992 2402 9996
rect 2406 9992 2409 9996
rect 2413 9992 2416 9996
rect 2420 9992 2423 9996
rect 2427 9992 2430 9996
rect 2434 9992 2437 9996
rect 2441 9992 2444 9996
rect 2448 9992 2451 9996
rect 2455 9992 2458 9996
rect 2462 9992 2465 9996
rect 2469 9993 2484 9996
rect 2677 10001 2793 10003
rect 2677 9997 2690 10001
rect 2694 9997 2697 10001
rect 2701 9997 2704 10001
rect 2708 9997 2711 10001
rect 2715 9997 2718 10001
rect 2722 9997 2725 10001
rect 2729 9997 2732 10001
rect 2736 9997 2739 10001
rect 2743 9997 2746 10001
rect 2750 9997 2753 10001
rect 2757 9997 2760 10001
rect 2764 9997 2767 10001
rect 2771 9997 2774 10001
rect 2778 9997 2793 10001
rect 2677 9996 2793 9997
rect 2677 9993 2690 9996
rect 2469 9992 2474 9993
rect 2378 9991 2474 9992
rect 2378 9987 2381 9991
rect 2385 9987 2388 9991
rect 2392 9987 2395 9991
rect 2399 9987 2402 9991
rect 2406 9987 2409 9991
rect 2413 9987 2416 9991
rect 2420 9987 2423 9991
rect 2427 9987 2430 9991
rect 2434 9987 2437 9991
rect 2441 9987 2444 9991
rect 2448 9987 2451 9991
rect 2455 9987 2458 9991
rect 2462 9987 2465 9991
rect 2469 9987 2474 9991
rect 2378 9986 2474 9987
rect 2378 9982 2381 9986
rect 2385 9982 2388 9986
rect 2392 9982 2395 9986
rect 2399 9982 2402 9986
rect 2406 9982 2409 9986
rect 2413 9982 2416 9986
rect 2420 9982 2423 9986
rect 2427 9982 2430 9986
rect 2434 9982 2437 9986
rect 2441 9982 2444 9986
rect 2448 9982 2451 9986
rect 2455 9982 2458 9986
rect 2462 9982 2465 9986
rect 2469 9982 2474 9986
rect 2378 9981 2474 9982
rect 2687 9992 2690 9993
rect 2694 9992 2697 9996
rect 2701 9992 2704 9996
rect 2708 9992 2711 9996
rect 2715 9992 2718 9996
rect 2722 9992 2725 9996
rect 2729 9992 2732 9996
rect 2736 9992 2739 9996
rect 2743 9992 2746 9996
rect 2750 9992 2753 9996
rect 2757 9992 2760 9996
rect 2764 9992 2767 9996
rect 2771 9992 2774 9996
rect 2778 9993 2793 9996
rect 2986 10001 3102 10003
rect 2986 9997 2999 10001
rect 3003 9997 3006 10001
rect 3010 9997 3013 10001
rect 3017 9997 3020 10001
rect 3024 9997 3027 10001
rect 3031 9997 3034 10001
rect 3038 9997 3041 10001
rect 3045 9997 3048 10001
rect 3052 9997 3055 10001
rect 3059 9997 3062 10001
rect 3066 9997 3069 10001
rect 3073 9997 3076 10001
rect 3080 9997 3083 10001
rect 3087 9997 3102 10001
rect 2986 9996 3102 9997
rect 2986 9993 2999 9996
rect 2778 9992 2783 9993
rect 2687 9991 2783 9992
rect 2687 9987 2690 9991
rect 2694 9987 2697 9991
rect 2701 9987 2704 9991
rect 2708 9987 2711 9991
rect 2715 9987 2718 9991
rect 2722 9987 2725 9991
rect 2729 9987 2732 9991
rect 2736 9987 2739 9991
rect 2743 9987 2746 9991
rect 2750 9987 2753 9991
rect 2757 9987 2760 9991
rect 2764 9987 2767 9991
rect 2771 9987 2774 9991
rect 2778 9987 2783 9991
rect 2687 9986 2783 9987
rect 2687 9982 2690 9986
rect 2694 9982 2697 9986
rect 2701 9982 2704 9986
rect 2708 9982 2711 9986
rect 2715 9982 2718 9986
rect 2722 9982 2725 9986
rect 2729 9982 2732 9986
rect 2736 9982 2739 9986
rect 2743 9982 2746 9986
rect 2750 9982 2753 9986
rect 2757 9982 2760 9986
rect 2764 9982 2767 9986
rect 2771 9982 2774 9986
rect 2778 9982 2783 9986
rect 2687 9981 2783 9982
rect 2996 9992 2999 9993
rect 3003 9992 3006 9996
rect 3010 9992 3013 9996
rect 3017 9992 3020 9996
rect 3024 9992 3027 9996
rect 3031 9992 3034 9996
rect 3038 9992 3041 9996
rect 3045 9992 3048 9996
rect 3052 9992 3055 9996
rect 3059 9992 3062 9996
rect 3066 9992 3069 9996
rect 3073 9992 3076 9996
rect 3080 9992 3083 9996
rect 3087 9993 3102 9996
rect 3295 10001 3411 10003
rect 3295 9997 3308 10001
rect 3312 9997 3315 10001
rect 3319 9997 3322 10001
rect 3326 9997 3329 10001
rect 3333 9997 3336 10001
rect 3340 9997 3343 10001
rect 3347 9997 3350 10001
rect 3354 9997 3357 10001
rect 3361 9997 3364 10001
rect 3368 9997 3371 10001
rect 3375 9997 3378 10001
rect 3382 9997 3385 10001
rect 3389 9997 3392 10001
rect 3396 9997 3411 10001
rect 3295 9996 3411 9997
rect 3295 9993 3308 9996
rect 3087 9992 3092 9993
rect 2996 9991 3092 9992
rect 2996 9987 2999 9991
rect 3003 9987 3006 9991
rect 3010 9987 3013 9991
rect 3017 9987 3020 9991
rect 3024 9987 3027 9991
rect 3031 9987 3034 9991
rect 3038 9987 3041 9991
rect 3045 9987 3048 9991
rect 3052 9987 3055 9991
rect 3059 9987 3062 9991
rect 3066 9987 3069 9991
rect 3073 9987 3076 9991
rect 3080 9987 3083 9991
rect 3087 9987 3092 9991
rect 2996 9986 3092 9987
rect 2996 9982 2999 9986
rect 3003 9982 3006 9986
rect 3010 9982 3013 9986
rect 3017 9982 3020 9986
rect 3024 9982 3027 9986
rect 3031 9982 3034 9986
rect 3038 9982 3041 9986
rect 3045 9982 3048 9986
rect 3052 9982 3055 9986
rect 3059 9982 3062 9986
rect 3066 9982 3069 9986
rect 3073 9982 3076 9986
rect 3080 9982 3083 9986
rect 3087 9982 3092 9986
rect 2996 9981 3092 9982
rect 3305 9992 3308 9993
rect 3312 9992 3315 9996
rect 3319 9992 3322 9996
rect 3326 9992 3329 9996
rect 3333 9992 3336 9996
rect 3340 9992 3343 9996
rect 3347 9992 3350 9996
rect 3354 9992 3357 9996
rect 3361 9992 3364 9996
rect 3368 9992 3371 9996
rect 3375 9992 3378 9996
rect 3382 9992 3385 9996
rect 3389 9992 3392 9996
rect 3396 9993 3411 9996
rect 3604 10001 3720 10003
rect 3604 9997 3617 10001
rect 3621 9997 3624 10001
rect 3628 9997 3631 10001
rect 3635 9997 3638 10001
rect 3642 9997 3645 10001
rect 3649 9997 3652 10001
rect 3656 9997 3659 10001
rect 3663 9997 3666 10001
rect 3670 9997 3673 10001
rect 3677 9997 3680 10001
rect 3684 9997 3687 10001
rect 3691 9997 3694 10001
rect 3698 9997 3701 10001
rect 3705 9997 3720 10001
rect 3604 9996 3720 9997
rect 3604 9993 3617 9996
rect 3396 9992 3401 9993
rect 3305 9991 3401 9992
rect 3305 9987 3308 9991
rect 3312 9987 3315 9991
rect 3319 9987 3322 9991
rect 3326 9987 3329 9991
rect 3333 9987 3336 9991
rect 3340 9987 3343 9991
rect 3347 9987 3350 9991
rect 3354 9987 3357 9991
rect 3361 9987 3364 9991
rect 3368 9987 3371 9991
rect 3375 9987 3378 9991
rect 3382 9987 3385 9991
rect 3389 9987 3392 9991
rect 3396 9987 3401 9991
rect 3305 9986 3401 9987
rect 3305 9982 3308 9986
rect 3312 9982 3315 9986
rect 3319 9982 3322 9986
rect 3326 9982 3329 9986
rect 3333 9982 3336 9986
rect 3340 9982 3343 9986
rect 3347 9982 3350 9986
rect 3354 9982 3357 9986
rect 3361 9982 3364 9986
rect 3368 9982 3371 9986
rect 3375 9982 3378 9986
rect 3382 9982 3385 9986
rect 3389 9982 3392 9986
rect 3396 9982 3401 9986
rect 3305 9981 3401 9982
rect 3614 9992 3617 9993
rect 3621 9992 3624 9996
rect 3628 9992 3631 9996
rect 3635 9992 3638 9996
rect 3642 9992 3645 9996
rect 3649 9992 3652 9996
rect 3656 9992 3659 9996
rect 3663 9992 3666 9996
rect 3670 9992 3673 9996
rect 3677 9992 3680 9996
rect 3684 9992 3687 9996
rect 3691 9992 3694 9996
rect 3698 9992 3701 9996
rect 3705 9993 3720 9996
rect 3913 10001 4029 10003
rect 3913 9997 3926 10001
rect 3930 9997 3933 10001
rect 3937 9997 3940 10001
rect 3944 9997 3947 10001
rect 3951 9997 3954 10001
rect 3958 9997 3961 10001
rect 3965 9997 3968 10001
rect 3972 9997 3975 10001
rect 3979 9997 3982 10001
rect 3986 9997 3989 10001
rect 3993 9997 3996 10001
rect 4000 9997 4003 10001
rect 4007 9997 4010 10001
rect 4014 9997 4029 10001
rect 3913 9996 4029 9997
rect 3913 9993 3926 9996
rect 3705 9992 3710 9993
rect 3614 9991 3710 9992
rect 3614 9987 3617 9991
rect 3621 9987 3624 9991
rect 3628 9987 3631 9991
rect 3635 9987 3638 9991
rect 3642 9987 3645 9991
rect 3649 9987 3652 9991
rect 3656 9987 3659 9991
rect 3663 9987 3666 9991
rect 3670 9987 3673 9991
rect 3677 9987 3680 9991
rect 3684 9987 3687 9991
rect 3691 9987 3694 9991
rect 3698 9987 3701 9991
rect 3705 9987 3710 9991
rect 3614 9986 3710 9987
rect 3614 9982 3617 9986
rect 3621 9982 3624 9986
rect 3628 9982 3631 9986
rect 3635 9982 3638 9986
rect 3642 9982 3645 9986
rect 3649 9982 3652 9986
rect 3656 9982 3659 9986
rect 3663 9982 3666 9986
rect 3670 9982 3673 9986
rect 3677 9982 3680 9986
rect 3684 9982 3687 9986
rect 3691 9982 3694 9986
rect 3698 9982 3701 9986
rect 3705 9982 3710 9986
rect 3614 9981 3710 9982
rect 3923 9992 3926 9993
rect 3930 9992 3933 9996
rect 3937 9992 3940 9996
rect 3944 9992 3947 9996
rect 3951 9992 3954 9996
rect 3958 9992 3961 9996
rect 3965 9992 3968 9996
rect 3972 9992 3975 9996
rect 3979 9992 3982 9996
rect 3986 9992 3989 9996
rect 3993 9992 3996 9996
rect 4000 9992 4003 9996
rect 4007 9992 4010 9996
rect 4014 9993 4029 9996
rect 4014 9992 4019 9993
rect 3923 9991 4019 9992
rect 3923 9987 3926 9991
rect 3930 9987 3933 9991
rect 3937 9987 3940 9991
rect 3944 9987 3947 9991
rect 3951 9987 3954 9991
rect 3958 9987 3961 9991
rect 3965 9987 3968 9991
rect 3972 9987 3975 9991
rect 3979 9987 3982 9991
rect 3986 9987 3989 9991
rect 3993 9987 3996 9991
rect 4000 9987 4003 9991
rect 4007 9987 4010 9991
rect 4014 9987 4019 9991
rect 3923 9986 4019 9987
rect 3923 9982 3926 9986
rect 3930 9982 3933 9986
rect 3937 9982 3940 9986
rect 3944 9982 3947 9986
rect 3951 9982 3954 9986
rect 3958 9982 3961 9986
rect 3965 9982 3968 9986
rect 3972 9982 3975 9986
rect 3979 9982 3982 9986
rect 3986 9982 3989 9986
rect 3993 9982 3996 9986
rect 4000 9982 4003 9986
rect 4007 9982 4010 9986
rect 4014 9982 4019 9986
rect 3923 9981 4019 9982
rect 1376 9974 1377 9978
rect 1381 9974 1382 9978
rect 1386 9974 1387 9978
rect 1391 9974 1392 9978
rect 1396 9974 1397 9978
rect 1401 9974 1402 9978
rect 1406 9974 1407 9978
rect 1411 9974 1412 9978
rect 1416 9974 1417 9978
rect 1421 9974 1422 9978
rect 1426 9974 1427 9978
rect 1431 9974 1432 9978
rect 1436 9974 1437 9978
rect 1441 9974 1442 9978
rect 1446 9974 1447 9978
rect 1451 9974 1452 9978
rect 1456 9974 1457 9978
rect 1461 9974 1462 9978
rect 1372 9973 1376 9974
rect 1372 9968 1376 9969
rect 1462 9973 1466 9974
rect 1462 9968 1466 9969
rect 1372 9963 1376 9964
rect 1372 9958 1376 9959
rect 1372 9953 1376 9954
rect 1372 9948 1376 9949
rect 1372 9943 1376 9944
rect 1372 9938 1376 9939
rect 1372 9933 1376 9934
rect 1372 9928 1376 9929
rect 1372 9923 1376 9924
rect 1372 9918 1376 9919
rect 1372 9913 1376 9914
rect 1372 9908 1376 9909
rect 1372 9903 1376 9904
rect 1372 9898 1376 9899
rect 1372 9893 1376 9894
rect 1372 9888 1376 9889
rect 1372 9883 1376 9884
rect 1372 9878 1376 9879
rect 1372 9873 1376 9874
rect 1372 9868 1376 9869
rect 1372 9863 1376 9864
rect 1372 9858 1376 9859
rect 1372 9853 1376 9854
rect 1372 9848 1376 9849
rect 1389 9961 1392 9965
rect 1396 9961 1397 9965
rect 1401 9961 1402 9965
rect 1406 9961 1407 9965
rect 1411 9961 1412 9965
rect 1416 9961 1417 9965
rect 1421 9961 1422 9965
rect 1426 9961 1427 9965
rect 1431 9961 1432 9965
rect 1436 9961 1437 9965
rect 1441 9961 1442 9965
rect 1446 9961 1449 9965
rect 1385 9958 1389 9961
rect 1385 9953 1389 9954
rect 1449 9958 1453 9961
rect 1449 9953 1453 9954
rect 1385 9948 1389 9949
rect 1385 9943 1389 9944
rect 1385 9938 1389 9939
rect 1385 9933 1389 9934
rect 1385 9928 1389 9929
rect 1385 9923 1389 9924
rect 1385 9918 1389 9919
rect 1385 9913 1389 9914
rect 1385 9908 1389 9909
rect 1385 9903 1389 9904
rect 1385 9898 1389 9899
rect 1385 9893 1389 9894
rect 1385 9888 1389 9889
rect 1385 9883 1389 9884
rect 1385 9878 1389 9879
rect 1385 9873 1389 9874
rect 1385 9868 1389 9869
rect 1401 9949 1402 9953
rect 1406 9949 1407 9953
rect 1411 9949 1412 9953
rect 1416 9949 1417 9953
rect 1421 9949 1422 9953
rect 1426 9949 1427 9953
rect 1431 9949 1432 9953
rect 1436 9949 1437 9953
rect 1397 9948 1441 9949
rect 1401 9944 1402 9948
rect 1406 9944 1407 9948
rect 1411 9944 1412 9948
rect 1416 9944 1417 9948
rect 1421 9944 1422 9948
rect 1426 9944 1427 9948
rect 1431 9944 1432 9948
rect 1436 9944 1437 9948
rect 1397 9943 1441 9944
rect 1401 9939 1402 9943
rect 1406 9939 1407 9943
rect 1411 9939 1412 9943
rect 1416 9939 1417 9943
rect 1421 9939 1422 9943
rect 1426 9939 1427 9943
rect 1431 9939 1432 9943
rect 1436 9939 1437 9943
rect 1397 9938 1441 9939
rect 1401 9934 1402 9938
rect 1406 9934 1407 9938
rect 1411 9934 1412 9938
rect 1416 9934 1417 9938
rect 1421 9934 1422 9938
rect 1426 9934 1427 9938
rect 1431 9934 1432 9938
rect 1436 9934 1437 9938
rect 1397 9933 1441 9934
rect 1401 9929 1402 9933
rect 1406 9929 1407 9933
rect 1411 9929 1412 9933
rect 1416 9929 1417 9933
rect 1421 9929 1422 9933
rect 1426 9929 1427 9933
rect 1431 9929 1432 9933
rect 1436 9929 1437 9933
rect 1397 9928 1441 9929
rect 1401 9924 1402 9928
rect 1406 9924 1407 9928
rect 1411 9924 1412 9928
rect 1416 9924 1417 9928
rect 1421 9924 1422 9928
rect 1426 9924 1427 9928
rect 1431 9924 1432 9928
rect 1436 9924 1437 9928
rect 1397 9923 1441 9924
rect 1401 9919 1402 9923
rect 1406 9919 1407 9923
rect 1411 9919 1412 9923
rect 1416 9919 1417 9923
rect 1421 9919 1422 9923
rect 1426 9919 1427 9923
rect 1431 9919 1432 9923
rect 1436 9919 1437 9923
rect 1397 9918 1441 9919
rect 1401 9914 1402 9918
rect 1406 9914 1407 9918
rect 1411 9914 1412 9918
rect 1416 9914 1417 9918
rect 1421 9914 1422 9918
rect 1426 9914 1427 9918
rect 1431 9914 1432 9918
rect 1436 9914 1437 9918
rect 1397 9913 1441 9914
rect 1401 9909 1402 9913
rect 1406 9909 1407 9913
rect 1411 9909 1412 9913
rect 1416 9909 1417 9913
rect 1421 9909 1422 9913
rect 1426 9909 1427 9913
rect 1431 9909 1432 9913
rect 1436 9909 1437 9913
rect 1397 9908 1441 9909
rect 1401 9904 1402 9908
rect 1406 9904 1407 9908
rect 1411 9904 1412 9908
rect 1416 9904 1417 9908
rect 1421 9904 1422 9908
rect 1426 9904 1427 9908
rect 1431 9904 1432 9908
rect 1436 9904 1437 9908
rect 1397 9903 1441 9904
rect 1401 9899 1402 9903
rect 1406 9899 1407 9903
rect 1411 9899 1412 9903
rect 1416 9899 1417 9903
rect 1421 9899 1422 9903
rect 1426 9899 1427 9903
rect 1431 9899 1432 9903
rect 1436 9899 1437 9903
rect 1397 9898 1441 9899
rect 1401 9894 1402 9898
rect 1406 9894 1407 9898
rect 1411 9894 1412 9898
rect 1416 9894 1417 9898
rect 1421 9894 1422 9898
rect 1426 9894 1427 9898
rect 1431 9894 1432 9898
rect 1436 9894 1437 9898
rect 1397 9893 1441 9894
rect 1401 9889 1402 9893
rect 1406 9889 1407 9893
rect 1411 9889 1412 9893
rect 1416 9889 1417 9893
rect 1421 9889 1422 9893
rect 1426 9889 1427 9893
rect 1431 9889 1432 9893
rect 1436 9889 1437 9893
rect 1397 9888 1441 9889
rect 1401 9884 1402 9888
rect 1406 9884 1407 9888
rect 1411 9884 1412 9888
rect 1416 9884 1417 9888
rect 1421 9884 1422 9888
rect 1426 9884 1427 9888
rect 1431 9884 1432 9888
rect 1436 9884 1437 9888
rect 1397 9883 1441 9884
rect 1401 9879 1402 9883
rect 1406 9879 1407 9883
rect 1411 9879 1412 9883
rect 1416 9879 1417 9883
rect 1421 9879 1422 9883
rect 1426 9879 1427 9883
rect 1431 9879 1432 9883
rect 1436 9879 1437 9883
rect 1397 9878 1441 9879
rect 1401 9874 1402 9878
rect 1406 9874 1407 9878
rect 1411 9874 1412 9878
rect 1416 9874 1417 9878
rect 1421 9874 1422 9878
rect 1426 9874 1427 9878
rect 1431 9874 1432 9878
rect 1436 9874 1437 9878
rect 1397 9873 1441 9874
rect 1401 9869 1402 9873
rect 1406 9869 1407 9873
rect 1411 9869 1412 9873
rect 1416 9869 1417 9873
rect 1421 9869 1422 9873
rect 1426 9869 1427 9873
rect 1431 9869 1432 9873
rect 1436 9869 1437 9873
rect 1397 9868 1441 9869
rect 1401 9864 1402 9868
rect 1406 9864 1407 9868
rect 1411 9864 1412 9868
rect 1416 9864 1417 9868
rect 1421 9864 1422 9868
rect 1426 9864 1427 9868
rect 1431 9864 1432 9868
rect 1436 9864 1437 9868
rect 1449 9948 1453 9949
rect 1449 9943 1453 9944
rect 1449 9938 1453 9939
rect 1449 9933 1453 9934
rect 1449 9928 1453 9929
rect 1449 9923 1453 9924
rect 1449 9918 1453 9919
rect 1449 9913 1453 9914
rect 1449 9908 1453 9909
rect 1449 9903 1453 9904
rect 1449 9898 1453 9899
rect 1449 9893 1453 9894
rect 1449 9888 1453 9889
rect 1449 9883 1453 9884
rect 1449 9878 1453 9879
rect 1449 9873 1453 9874
rect 1449 9868 1453 9869
rect 1385 9863 1389 9864
rect 1385 9856 1389 9859
rect 1449 9863 1453 9864
rect 1449 9856 1453 9859
rect 1389 9848 1392 9856
rect 1396 9848 1397 9856
rect 1401 9848 1402 9856
rect 1406 9848 1407 9856
rect 1411 9848 1412 9856
rect 1416 9848 1417 9856
rect 1421 9848 1422 9856
rect 1426 9848 1427 9856
rect 1431 9848 1432 9856
rect 1436 9848 1437 9856
rect 1441 9848 1442 9856
rect 1446 9848 1449 9856
rect 1462 9963 1466 9964
rect 1462 9958 1466 9959
rect 1462 9953 1466 9954
rect 1462 9948 1466 9949
rect 1462 9943 1466 9944
rect 1462 9938 1466 9939
rect 1462 9933 1466 9934
rect 1462 9928 1466 9929
rect 1462 9923 1466 9924
rect 1462 9918 1466 9919
rect 1462 9913 1466 9914
rect 1462 9908 1466 9909
rect 1462 9903 1466 9904
rect 1462 9898 1466 9899
rect 1462 9893 1466 9894
rect 1462 9888 1466 9889
rect 1462 9883 1466 9884
rect 1462 9878 1466 9879
rect 1462 9873 1466 9874
rect 1462 9868 1466 9869
rect 1462 9863 1466 9864
rect 1462 9858 1466 9859
rect 1462 9853 1466 9854
rect 1462 9848 1466 9849
rect 1372 9843 1376 9844
rect 1462 9843 1466 9844
rect 1376 9839 1377 9843
rect 1381 9839 1382 9843
rect 1386 9839 1387 9843
rect 1391 9839 1392 9843
rect 1396 9839 1397 9843
rect 1401 9839 1402 9843
rect 1406 9839 1407 9843
rect 1411 9839 1412 9843
rect 1416 9839 1417 9843
rect 1421 9839 1422 9843
rect 1426 9839 1427 9843
rect 1431 9839 1432 9843
rect 1436 9839 1437 9843
rect 1441 9839 1442 9843
rect 1446 9839 1447 9843
rect 1451 9839 1452 9843
rect 1456 9839 1457 9843
rect 1461 9839 1462 9843
rect 1375 9802 1431 9839
rect 1363 9800 1431 9802
rect 1363 9796 1364 9800
rect 1368 9796 1369 9800
rect 1373 9796 1431 9800
rect 1363 9795 1431 9796
rect 1363 9791 1364 9795
rect 1368 9791 1369 9795
rect 1373 9791 1431 9795
rect 1363 9790 1431 9791
rect 1363 9786 1364 9790
rect 1368 9786 1369 9790
rect 1373 9786 1431 9790
rect 1363 9785 1431 9786
rect 1363 9781 1364 9785
rect 1368 9781 1369 9785
rect 1373 9781 1431 9785
rect 1363 9780 1431 9781
rect 1363 9776 1364 9780
rect 1368 9776 1369 9780
rect 1373 9776 1431 9780
rect 1363 9775 1431 9776
rect 1363 9771 1364 9775
rect 1368 9771 1369 9775
rect 1373 9771 1431 9775
rect 1363 9770 1431 9771
rect 1363 9766 1364 9770
rect 1368 9766 1369 9770
rect 1373 9766 1431 9770
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1319 9761 1338 9762
rect 1323 9757 1324 9761
rect 1328 9757 1329 9761
rect 1333 9757 1334 9761
rect 1319 9756 1338 9757
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1319 9751 1338 9752
rect 1323 9747 1324 9751
rect 1328 9747 1329 9751
rect 1333 9747 1334 9751
rect 1319 9746 1338 9747
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1319 9741 1338 9742
rect 1323 9737 1324 9741
rect 1328 9737 1329 9741
rect 1333 9737 1334 9741
rect 1319 9736 1338 9737
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1363 9765 1431 9766
rect 1363 9761 1364 9765
rect 1368 9761 1369 9765
rect 1373 9761 1431 9765
rect 1363 9760 1431 9761
rect 1363 9756 1364 9760
rect 1368 9756 1369 9760
rect 1373 9756 1431 9760
rect 1363 9755 1431 9756
rect 1363 9751 1364 9755
rect 1368 9751 1369 9755
rect 1373 9751 1431 9755
rect 1363 9750 1431 9751
rect 1363 9746 1364 9750
rect 1368 9746 1369 9750
rect 1373 9746 1431 9750
rect 1363 9745 1431 9746
rect 1363 9741 1364 9745
rect 1368 9741 1369 9745
rect 1373 9741 1431 9745
rect 1363 9740 1431 9741
rect 1363 9736 1364 9740
rect 1368 9736 1369 9740
rect 1373 9736 1431 9740
rect 1363 9734 1431 9736
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1319 9715 1338 9716
rect 1323 9711 1324 9715
rect 1328 9711 1329 9715
rect 1333 9711 1334 9715
rect 1319 9710 1338 9711
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1319 9705 1338 9706
rect 1323 9701 1324 9705
rect 1328 9701 1329 9705
rect 1333 9701 1334 9705
rect 1319 9700 1338 9701
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1319 9695 1338 9696
rect 1323 9691 1324 9695
rect 1328 9691 1329 9695
rect 1333 9691 1334 9695
rect 1319 9690 1338 9691
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1473 9715 1525 9981
rect 1536 9974 1537 9978
rect 1541 9974 1542 9978
rect 1546 9974 1547 9978
rect 1551 9974 1552 9978
rect 1556 9974 1557 9978
rect 1561 9974 1562 9978
rect 1566 9974 1567 9978
rect 1571 9974 1572 9978
rect 1576 9974 1577 9978
rect 1581 9974 1582 9978
rect 1586 9974 1587 9978
rect 1591 9974 1592 9978
rect 1596 9974 1597 9978
rect 1601 9974 1602 9978
rect 1606 9974 1607 9978
rect 1611 9974 1612 9978
rect 1616 9974 1617 9978
rect 1621 9974 1622 9978
rect 1532 9973 1536 9974
rect 1532 9968 1536 9969
rect 1622 9973 1626 9974
rect 1622 9968 1626 9969
rect 1532 9963 1536 9964
rect 1532 9958 1536 9959
rect 1532 9953 1536 9954
rect 1532 9948 1536 9949
rect 1532 9943 1536 9944
rect 1532 9938 1536 9939
rect 1532 9933 1536 9934
rect 1532 9928 1536 9929
rect 1532 9923 1536 9924
rect 1532 9918 1536 9919
rect 1532 9913 1536 9914
rect 1532 9908 1536 9909
rect 1532 9903 1536 9904
rect 1532 9898 1536 9899
rect 1532 9893 1536 9894
rect 1532 9888 1536 9889
rect 1532 9883 1536 9884
rect 1532 9878 1536 9879
rect 1532 9873 1536 9874
rect 1532 9868 1536 9869
rect 1532 9863 1536 9864
rect 1532 9858 1536 9859
rect 1532 9853 1536 9854
rect 1532 9848 1536 9849
rect 1549 9961 1552 9965
rect 1556 9961 1557 9965
rect 1561 9961 1562 9965
rect 1566 9961 1567 9965
rect 1571 9961 1572 9965
rect 1576 9961 1577 9965
rect 1581 9961 1582 9965
rect 1586 9961 1587 9965
rect 1591 9961 1592 9965
rect 1596 9961 1597 9965
rect 1601 9961 1602 9965
rect 1606 9961 1609 9965
rect 1545 9958 1549 9961
rect 1545 9953 1549 9954
rect 1609 9958 1613 9961
rect 1609 9953 1613 9954
rect 1545 9948 1549 9949
rect 1545 9943 1549 9944
rect 1545 9938 1549 9939
rect 1545 9933 1549 9934
rect 1545 9928 1549 9929
rect 1545 9923 1549 9924
rect 1545 9918 1549 9919
rect 1545 9913 1549 9914
rect 1545 9908 1549 9909
rect 1545 9903 1549 9904
rect 1545 9898 1549 9899
rect 1545 9893 1549 9894
rect 1545 9888 1549 9889
rect 1545 9883 1549 9884
rect 1545 9878 1549 9879
rect 1545 9873 1549 9874
rect 1545 9868 1549 9869
rect 1556 9949 1557 9953
rect 1561 9949 1562 9953
rect 1566 9949 1567 9953
rect 1571 9949 1572 9953
rect 1576 9949 1577 9953
rect 1581 9949 1582 9953
rect 1586 9949 1587 9953
rect 1591 9949 1592 9953
rect 1596 9949 1597 9953
rect 1556 9948 1601 9949
rect 1556 9944 1557 9948
rect 1561 9944 1562 9948
rect 1566 9944 1567 9948
rect 1571 9944 1572 9948
rect 1576 9944 1577 9948
rect 1581 9944 1582 9948
rect 1586 9944 1587 9948
rect 1591 9944 1592 9948
rect 1596 9944 1597 9948
rect 1556 9943 1601 9944
rect 1556 9939 1557 9943
rect 1561 9939 1562 9943
rect 1566 9939 1567 9943
rect 1571 9939 1572 9943
rect 1576 9939 1577 9943
rect 1581 9939 1582 9943
rect 1586 9939 1587 9943
rect 1591 9939 1592 9943
rect 1596 9939 1597 9943
rect 1556 9938 1601 9939
rect 1556 9934 1557 9938
rect 1561 9934 1562 9938
rect 1566 9934 1567 9938
rect 1571 9934 1572 9938
rect 1576 9934 1577 9938
rect 1581 9934 1582 9938
rect 1586 9934 1587 9938
rect 1591 9934 1592 9938
rect 1596 9934 1597 9938
rect 1556 9933 1601 9934
rect 1556 9929 1557 9933
rect 1561 9929 1562 9933
rect 1566 9929 1567 9933
rect 1571 9929 1572 9933
rect 1576 9929 1577 9933
rect 1581 9929 1582 9933
rect 1586 9929 1587 9933
rect 1591 9929 1592 9933
rect 1596 9929 1597 9933
rect 1556 9928 1601 9929
rect 1556 9924 1557 9928
rect 1561 9924 1562 9928
rect 1566 9924 1567 9928
rect 1571 9924 1572 9928
rect 1576 9924 1577 9928
rect 1581 9924 1582 9928
rect 1586 9924 1587 9928
rect 1591 9924 1592 9928
rect 1596 9924 1597 9928
rect 1556 9923 1601 9924
rect 1556 9919 1557 9923
rect 1561 9919 1562 9923
rect 1566 9919 1567 9923
rect 1571 9919 1572 9923
rect 1576 9919 1577 9923
rect 1581 9919 1582 9923
rect 1586 9919 1587 9923
rect 1591 9919 1592 9923
rect 1596 9919 1597 9923
rect 1556 9918 1601 9919
rect 1556 9914 1557 9918
rect 1561 9914 1562 9918
rect 1566 9914 1567 9918
rect 1571 9914 1572 9918
rect 1576 9914 1577 9918
rect 1581 9914 1582 9918
rect 1586 9914 1587 9918
rect 1591 9914 1592 9918
rect 1596 9914 1597 9918
rect 1556 9913 1601 9914
rect 1556 9909 1557 9913
rect 1561 9909 1562 9913
rect 1566 9909 1567 9913
rect 1571 9909 1572 9913
rect 1576 9909 1577 9913
rect 1581 9909 1582 9913
rect 1586 9909 1587 9913
rect 1591 9909 1592 9913
rect 1596 9909 1597 9913
rect 1556 9908 1601 9909
rect 1556 9904 1557 9908
rect 1561 9904 1562 9908
rect 1566 9904 1567 9908
rect 1571 9904 1572 9908
rect 1576 9904 1577 9908
rect 1581 9904 1582 9908
rect 1586 9904 1587 9908
rect 1591 9904 1592 9908
rect 1596 9904 1597 9908
rect 1556 9903 1601 9904
rect 1556 9899 1557 9903
rect 1561 9899 1562 9903
rect 1566 9899 1567 9903
rect 1571 9899 1572 9903
rect 1576 9899 1577 9903
rect 1581 9899 1582 9903
rect 1586 9899 1587 9903
rect 1591 9899 1592 9903
rect 1596 9899 1597 9903
rect 1556 9898 1601 9899
rect 1556 9894 1557 9898
rect 1561 9894 1562 9898
rect 1566 9894 1567 9898
rect 1571 9894 1572 9898
rect 1576 9894 1577 9898
rect 1581 9894 1582 9898
rect 1586 9894 1587 9898
rect 1591 9894 1592 9898
rect 1596 9894 1597 9898
rect 1556 9893 1601 9894
rect 1556 9889 1557 9893
rect 1561 9889 1562 9893
rect 1566 9889 1567 9893
rect 1571 9889 1572 9893
rect 1576 9889 1577 9893
rect 1581 9889 1582 9893
rect 1586 9889 1587 9893
rect 1591 9889 1592 9893
rect 1596 9889 1597 9893
rect 1556 9888 1601 9889
rect 1556 9884 1557 9888
rect 1561 9884 1562 9888
rect 1566 9884 1567 9888
rect 1571 9884 1572 9888
rect 1576 9884 1577 9888
rect 1581 9884 1582 9888
rect 1586 9884 1587 9888
rect 1591 9884 1592 9888
rect 1596 9884 1597 9888
rect 1556 9883 1601 9884
rect 1556 9879 1557 9883
rect 1561 9879 1562 9883
rect 1566 9879 1567 9883
rect 1571 9879 1572 9883
rect 1576 9879 1577 9883
rect 1581 9879 1582 9883
rect 1586 9879 1587 9883
rect 1591 9879 1592 9883
rect 1596 9879 1597 9883
rect 1556 9878 1601 9879
rect 1556 9874 1557 9878
rect 1561 9874 1562 9878
rect 1566 9874 1567 9878
rect 1571 9874 1572 9878
rect 1576 9874 1577 9878
rect 1581 9874 1582 9878
rect 1586 9874 1587 9878
rect 1591 9874 1592 9878
rect 1596 9874 1597 9878
rect 1556 9873 1601 9874
rect 1556 9869 1557 9873
rect 1561 9869 1562 9873
rect 1566 9869 1567 9873
rect 1571 9869 1572 9873
rect 1576 9869 1577 9873
rect 1581 9869 1582 9873
rect 1586 9869 1587 9873
rect 1591 9869 1592 9873
rect 1596 9869 1597 9873
rect 1556 9868 1601 9869
rect 1556 9864 1557 9868
rect 1561 9864 1562 9868
rect 1566 9864 1567 9868
rect 1571 9864 1572 9868
rect 1576 9864 1577 9868
rect 1581 9864 1582 9868
rect 1586 9864 1587 9868
rect 1591 9864 1592 9868
rect 1596 9864 1597 9868
rect 1609 9948 1613 9949
rect 1609 9943 1613 9944
rect 1609 9938 1613 9939
rect 1609 9933 1613 9934
rect 1609 9928 1613 9929
rect 1609 9923 1613 9924
rect 1609 9918 1613 9919
rect 1609 9913 1613 9914
rect 1609 9908 1613 9909
rect 1609 9903 1613 9904
rect 1609 9898 1613 9899
rect 1609 9893 1613 9894
rect 1609 9888 1613 9889
rect 1609 9883 1613 9884
rect 1609 9878 1613 9879
rect 1609 9873 1613 9874
rect 1609 9868 1613 9869
rect 1545 9863 1549 9864
rect 1545 9856 1549 9859
rect 1609 9863 1613 9864
rect 1609 9856 1613 9859
rect 1549 9848 1552 9856
rect 1556 9848 1557 9856
rect 1561 9848 1562 9856
rect 1566 9848 1567 9856
rect 1571 9848 1572 9856
rect 1576 9848 1577 9856
rect 1581 9848 1582 9856
rect 1586 9848 1587 9856
rect 1591 9848 1592 9856
rect 1596 9848 1597 9856
rect 1601 9848 1602 9856
rect 1606 9848 1609 9856
rect 1622 9963 1626 9964
rect 1622 9958 1626 9959
rect 1622 9953 1626 9954
rect 1622 9948 1626 9949
rect 1622 9943 1626 9944
rect 1622 9938 1626 9939
rect 1622 9933 1626 9934
rect 1622 9928 1626 9929
rect 1622 9923 1626 9924
rect 1622 9918 1626 9919
rect 1622 9913 1626 9914
rect 1622 9908 1626 9909
rect 1622 9903 1626 9904
rect 1622 9898 1626 9899
rect 1622 9893 1626 9894
rect 1622 9888 1626 9889
rect 1622 9883 1626 9884
rect 1622 9878 1626 9879
rect 1622 9873 1626 9874
rect 1622 9868 1626 9869
rect 1622 9863 1626 9864
rect 1622 9858 1626 9859
rect 1622 9853 1626 9854
rect 1622 9848 1626 9849
rect 1532 9843 1536 9844
rect 1622 9843 1626 9844
rect 1536 9839 1537 9843
rect 1541 9839 1542 9843
rect 1546 9839 1547 9843
rect 1551 9839 1552 9843
rect 1556 9839 1557 9843
rect 1561 9839 1562 9843
rect 1566 9839 1567 9843
rect 1571 9839 1572 9843
rect 1576 9839 1577 9843
rect 1581 9839 1582 9843
rect 1586 9839 1587 9843
rect 1591 9839 1592 9843
rect 1596 9839 1597 9843
rect 1601 9839 1602 9843
rect 1606 9839 1607 9843
rect 1611 9839 1612 9843
rect 1616 9839 1617 9843
rect 1621 9839 1622 9843
rect 1685 9974 1686 9978
rect 1690 9974 1691 9978
rect 1695 9974 1696 9978
rect 1700 9974 1701 9978
rect 1705 9974 1706 9978
rect 1710 9974 1711 9978
rect 1715 9974 1716 9978
rect 1720 9974 1721 9978
rect 1725 9974 1726 9978
rect 1730 9974 1731 9978
rect 1735 9974 1736 9978
rect 1740 9974 1741 9978
rect 1745 9974 1746 9978
rect 1750 9974 1751 9978
rect 1755 9974 1756 9978
rect 1760 9974 1761 9978
rect 1765 9974 1766 9978
rect 1770 9974 1771 9978
rect 1681 9973 1685 9974
rect 1681 9968 1685 9969
rect 1771 9973 1775 9974
rect 1771 9968 1775 9969
rect 1681 9963 1685 9964
rect 1681 9958 1685 9959
rect 1681 9953 1685 9954
rect 1681 9948 1685 9949
rect 1681 9943 1685 9944
rect 1681 9938 1685 9939
rect 1681 9933 1685 9934
rect 1681 9928 1685 9929
rect 1681 9923 1685 9924
rect 1681 9918 1685 9919
rect 1681 9913 1685 9914
rect 1681 9908 1685 9909
rect 1681 9903 1685 9904
rect 1681 9898 1685 9899
rect 1681 9893 1685 9894
rect 1681 9888 1685 9889
rect 1681 9883 1685 9884
rect 1681 9878 1685 9879
rect 1681 9873 1685 9874
rect 1681 9868 1685 9869
rect 1681 9863 1685 9864
rect 1681 9858 1685 9859
rect 1681 9853 1685 9854
rect 1681 9848 1685 9849
rect 1698 9961 1701 9965
rect 1705 9961 1706 9965
rect 1710 9961 1711 9965
rect 1715 9961 1716 9965
rect 1720 9961 1721 9965
rect 1725 9961 1726 9965
rect 1730 9961 1731 9965
rect 1735 9961 1736 9965
rect 1740 9961 1741 9965
rect 1745 9961 1746 9965
rect 1750 9961 1751 9965
rect 1755 9961 1758 9965
rect 1694 9958 1698 9961
rect 1694 9953 1698 9954
rect 1758 9958 1762 9961
rect 1758 9953 1762 9954
rect 1694 9948 1698 9949
rect 1694 9943 1698 9944
rect 1694 9938 1698 9939
rect 1694 9933 1698 9934
rect 1694 9928 1698 9929
rect 1694 9923 1698 9924
rect 1694 9918 1698 9919
rect 1694 9913 1698 9914
rect 1694 9908 1698 9909
rect 1694 9903 1698 9904
rect 1694 9898 1698 9899
rect 1694 9893 1698 9894
rect 1694 9888 1698 9889
rect 1694 9883 1698 9884
rect 1694 9878 1698 9879
rect 1694 9873 1698 9874
rect 1694 9868 1698 9869
rect 1710 9949 1711 9953
rect 1715 9949 1716 9953
rect 1720 9949 1721 9953
rect 1725 9949 1726 9953
rect 1730 9949 1731 9953
rect 1735 9949 1736 9953
rect 1740 9949 1741 9953
rect 1745 9949 1746 9953
rect 1706 9948 1750 9949
rect 1710 9944 1711 9948
rect 1715 9944 1716 9948
rect 1720 9944 1721 9948
rect 1725 9944 1726 9948
rect 1730 9944 1731 9948
rect 1735 9944 1736 9948
rect 1740 9944 1741 9948
rect 1745 9944 1746 9948
rect 1706 9943 1750 9944
rect 1710 9939 1711 9943
rect 1715 9939 1716 9943
rect 1720 9939 1721 9943
rect 1725 9939 1726 9943
rect 1730 9939 1731 9943
rect 1735 9939 1736 9943
rect 1740 9939 1741 9943
rect 1745 9939 1746 9943
rect 1706 9938 1750 9939
rect 1710 9934 1711 9938
rect 1715 9934 1716 9938
rect 1720 9934 1721 9938
rect 1725 9934 1726 9938
rect 1730 9934 1731 9938
rect 1735 9934 1736 9938
rect 1740 9934 1741 9938
rect 1745 9934 1746 9938
rect 1706 9933 1750 9934
rect 1710 9929 1711 9933
rect 1715 9929 1716 9933
rect 1720 9929 1721 9933
rect 1725 9929 1726 9933
rect 1730 9929 1731 9933
rect 1735 9929 1736 9933
rect 1740 9929 1741 9933
rect 1745 9929 1746 9933
rect 1706 9928 1750 9929
rect 1710 9924 1711 9928
rect 1715 9924 1716 9928
rect 1720 9924 1721 9928
rect 1725 9924 1726 9928
rect 1730 9924 1731 9928
rect 1735 9924 1736 9928
rect 1740 9924 1741 9928
rect 1745 9924 1746 9928
rect 1706 9923 1750 9924
rect 1710 9919 1711 9923
rect 1715 9919 1716 9923
rect 1720 9919 1721 9923
rect 1725 9919 1726 9923
rect 1730 9919 1731 9923
rect 1735 9919 1736 9923
rect 1740 9919 1741 9923
rect 1745 9919 1746 9923
rect 1706 9918 1750 9919
rect 1710 9914 1711 9918
rect 1715 9914 1716 9918
rect 1720 9914 1721 9918
rect 1725 9914 1726 9918
rect 1730 9914 1731 9918
rect 1735 9914 1736 9918
rect 1740 9914 1741 9918
rect 1745 9914 1746 9918
rect 1706 9913 1750 9914
rect 1710 9909 1711 9913
rect 1715 9909 1716 9913
rect 1720 9909 1721 9913
rect 1725 9909 1726 9913
rect 1730 9909 1731 9913
rect 1735 9909 1736 9913
rect 1740 9909 1741 9913
rect 1745 9909 1746 9913
rect 1706 9908 1750 9909
rect 1710 9904 1711 9908
rect 1715 9904 1716 9908
rect 1720 9904 1721 9908
rect 1725 9904 1726 9908
rect 1730 9904 1731 9908
rect 1735 9904 1736 9908
rect 1740 9904 1741 9908
rect 1745 9904 1746 9908
rect 1706 9903 1750 9904
rect 1710 9899 1711 9903
rect 1715 9899 1716 9903
rect 1720 9899 1721 9903
rect 1725 9899 1726 9903
rect 1730 9899 1731 9903
rect 1735 9899 1736 9903
rect 1740 9899 1741 9903
rect 1745 9899 1746 9903
rect 1706 9898 1750 9899
rect 1710 9894 1711 9898
rect 1715 9894 1716 9898
rect 1720 9894 1721 9898
rect 1725 9894 1726 9898
rect 1730 9894 1731 9898
rect 1735 9894 1736 9898
rect 1740 9894 1741 9898
rect 1745 9894 1746 9898
rect 1706 9893 1750 9894
rect 1710 9889 1711 9893
rect 1715 9889 1716 9893
rect 1720 9889 1721 9893
rect 1725 9889 1726 9893
rect 1730 9889 1731 9893
rect 1735 9889 1736 9893
rect 1740 9889 1741 9893
rect 1745 9889 1746 9893
rect 1706 9888 1750 9889
rect 1710 9884 1711 9888
rect 1715 9884 1716 9888
rect 1720 9884 1721 9888
rect 1725 9884 1726 9888
rect 1730 9884 1731 9888
rect 1735 9884 1736 9888
rect 1740 9884 1741 9888
rect 1745 9884 1746 9888
rect 1706 9883 1750 9884
rect 1710 9879 1711 9883
rect 1715 9879 1716 9883
rect 1720 9879 1721 9883
rect 1725 9879 1726 9883
rect 1730 9879 1731 9883
rect 1735 9879 1736 9883
rect 1740 9879 1741 9883
rect 1745 9879 1746 9883
rect 1706 9878 1750 9879
rect 1710 9874 1711 9878
rect 1715 9874 1716 9878
rect 1720 9874 1721 9878
rect 1725 9874 1726 9878
rect 1730 9874 1731 9878
rect 1735 9874 1736 9878
rect 1740 9874 1741 9878
rect 1745 9874 1746 9878
rect 1706 9873 1750 9874
rect 1710 9869 1711 9873
rect 1715 9869 1716 9873
rect 1720 9869 1721 9873
rect 1725 9869 1726 9873
rect 1730 9869 1731 9873
rect 1735 9869 1736 9873
rect 1740 9869 1741 9873
rect 1745 9869 1746 9873
rect 1706 9868 1750 9869
rect 1710 9864 1711 9868
rect 1715 9864 1716 9868
rect 1720 9864 1721 9868
rect 1725 9864 1726 9868
rect 1730 9864 1731 9868
rect 1735 9864 1736 9868
rect 1740 9864 1741 9868
rect 1745 9864 1746 9868
rect 1758 9948 1762 9949
rect 1758 9943 1762 9944
rect 1758 9938 1762 9939
rect 1758 9933 1762 9934
rect 1758 9928 1762 9929
rect 1758 9923 1762 9924
rect 1758 9918 1762 9919
rect 1758 9913 1762 9914
rect 1758 9908 1762 9909
rect 1758 9903 1762 9904
rect 1758 9898 1762 9899
rect 1758 9893 1762 9894
rect 1758 9888 1762 9889
rect 1758 9883 1762 9884
rect 1758 9878 1762 9879
rect 1758 9873 1762 9874
rect 1758 9868 1762 9869
rect 1694 9863 1698 9864
rect 1694 9856 1698 9859
rect 1758 9863 1762 9864
rect 1758 9856 1762 9859
rect 1698 9848 1701 9856
rect 1705 9848 1706 9856
rect 1710 9848 1711 9856
rect 1715 9848 1716 9856
rect 1720 9848 1721 9856
rect 1725 9848 1726 9856
rect 1730 9848 1731 9856
rect 1735 9848 1736 9856
rect 1740 9848 1741 9856
rect 1745 9848 1746 9856
rect 1750 9848 1751 9856
rect 1755 9848 1758 9856
rect 1771 9963 1775 9964
rect 1771 9958 1775 9959
rect 1771 9953 1775 9954
rect 1797 9961 1818 9981
rect 1845 9974 1846 9978
rect 1850 9974 1851 9978
rect 1855 9974 1856 9978
rect 1860 9974 1861 9978
rect 1865 9974 1866 9978
rect 1870 9974 1871 9978
rect 1875 9974 1876 9978
rect 1880 9974 1881 9978
rect 1885 9974 1886 9978
rect 1890 9974 1891 9978
rect 1895 9974 1896 9978
rect 1900 9974 1901 9978
rect 1905 9974 1906 9978
rect 1910 9974 1911 9978
rect 1915 9974 1916 9978
rect 1920 9974 1921 9978
rect 1925 9974 1926 9978
rect 1930 9974 1931 9978
rect 1841 9973 1845 9974
rect 1841 9968 1845 9969
rect 1931 9973 1935 9974
rect 1931 9968 1935 9969
rect 1841 9963 1845 9964
rect 1841 9958 1845 9959
rect 1841 9953 1845 9954
rect 1771 9948 1775 9949
rect 1771 9943 1775 9944
rect 1771 9938 1775 9939
rect 1771 9933 1775 9934
rect 1771 9928 1775 9929
rect 1771 9923 1775 9924
rect 1771 9918 1775 9919
rect 1771 9913 1775 9914
rect 1771 9908 1775 9909
rect 1771 9903 1775 9904
rect 1771 9898 1775 9899
rect 1771 9893 1775 9894
rect 1771 9888 1775 9889
rect 1771 9883 1775 9884
rect 1841 9948 1845 9949
rect 1841 9943 1845 9944
rect 1841 9938 1845 9939
rect 1841 9933 1845 9934
rect 1841 9928 1845 9929
rect 1841 9923 1845 9924
rect 1841 9918 1845 9919
rect 1841 9913 1845 9914
rect 1841 9908 1845 9909
rect 1841 9903 1845 9904
rect 1841 9898 1845 9899
rect 1841 9893 1845 9894
rect 1841 9888 1845 9889
rect 1841 9883 1845 9884
rect 1771 9878 1775 9879
rect 1771 9873 1775 9874
rect 1771 9868 1775 9869
rect 1771 9863 1775 9864
rect 1771 9858 1775 9859
rect 1771 9853 1775 9854
rect 1771 9848 1775 9849
rect 1681 9843 1685 9844
rect 1797 9846 1818 9874
rect 1841 9878 1845 9879
rect 1841 9873 1845 9874
rect 1841 9868 1845 9869
rect 1841 9863 1845 9864
rect 1841 9858 1845 9859
rect 1841 9853 1845 9854
rect 1841 9848 1845 9849
rect 1858 9961 1861 9965
rect 1865 9961 1866 9965
rect 1870 9961 1871 9965
rect 1875 9961 1876 9965
rect 1880 9961 1881 9965
rect 1885 9961 1886 9965
rect 1890 9961 1891 9965
rect 1895 9961 1896 9965
rect 1900 9961 1901 9965
rect 1905 9961 1906 9965
rect 1910 9961 1911 9965
rect 1915 9961 1918 9965
rect 1854 9958 1858 9961
rect 1854 9953 1858 9954
rect 1918 9958 1922 9961
rect 1918 9953 1922 9954
rect 1854 9948 1858 9949
rect 1854 9943 1858 9944
rect 1854 9938 1858 9939
rect 1854 9933 1858 9934
rect 1854 9928 1858 9929
rect 1854 9923 1858 9924
rect 1854 9918 1858 9919
rect 1854 9913 1858 9914
rect 1854 9908 1858 9909
rect 1854 9903 1858 9904
rect 1854 9898 1858 9899
rect 1854 9893 1858 9894
rect 1854 9888 1858 9889
rect 1854 9883 1858 9884
rect 1854 9878 1858 9879
rect 1854 9873 1858 9874
rect 1854 9868 1858 9869
rect 1865 9949 1866 9953
rect 1870 9949 1871 9953
rect 1875 9949 1876 9953
rect 1880 9949 1881 9953
rect 1885 9949 1886 9953
rect 1890 9949 1891 9953
rect 1895 9949 1896 9953
rect 1900 9949 1901 9953
rect 1905 9949 1906 9953
rect 1865 9948 1910 9949
rect 1865 9944 1866 9948
rect 1870 9944 1871 9948
rect 1875 9944 1876 9948
rect 1880 9944 1881 9948
rect 1885 9944 1886 9948
rect 1890 9944 1891 9948
rect 1895 9944 1896 9948
rect 1900 9944 1901 9948
rect 1905 9944 1906 9948
rect 1865 9943 1910 9944
rect 1865 9939 1866 9943
rect 1870 9939 1871 9943
rect 1875 9939 1876 9943
rect 1880 9939 1881 9943
rect 1885 9939 1886 9943
rect 1890 9939 1891 9943
rect 1895 9939 1896 9943
rect 1900 9939 1901 9943
rect 1905 9939 1906 9943
rect 1865 9938 1910 9939
rect 1865 9934 1866 9938
rect 1870 9934 1871 9938
rect 1875 9934 1876 9938
rect 1880 9934 1881 9938
rect 1885 9934 1886 9938
rect 1890 9934 1891 9938
rect 1895 9934 1896 9938
rect 1900 9934 1901 9938
rect 1905 9934 1906 9938
rect 1865 9933 1910 9934
rect 1865 9929 1866 9933
rect 1870 9929 1871 9933
rect 1875 9929 1876 9933
rect 1880 9929 1881 9933
rect 1885 9929 1886 9933
rect 1890 9929 1891 9933
rect 1895 9929 1896 9933
rect 1900 9929 1901 9933
rect 1905 9929 1906 9933
rect 1865 9928 1910 9929
rect 1865 9924 1866 9928
rect 1870 9924 1871 9928
rect 1875 9924 1876 9928
rect 1880 9924 1881 9928
rect 1885 9924 1886 9928
rect 1890 9924 1891 9928
rect 1895 9924 1896 9928
rect 1900 9924 1901 9928
rect 1905 9924 1906 9928
rect 1865 9923 1910 9924
rect 1865 9919 1866 9923
rect 1870 9919 1871 9923
rect 1875 9919 1876 9923
rect 1880 9919 1881 9923
rect 1885 9919 1886 9923
rect 1890 9919 1891 9923
rect 1895 9919 1896 9923
rect 1900 9919 1901 9923
rect 1905 9919 1906 9923
rect 1865 9918 1910 9919
rect 1865 9914 1866 9918
rect 1870 9914 1871 9918
rect 1875 9914 1876 9918
rect 1880 9914 1881 9918
rect 1885 9914 1886 9918
rect 1890 9914 1891 9918
rect 1895 9914 1896 9918
rect 1900 9914 1901 9918
rect 1905 9914 1906 9918
rect 1865 9913 1910 9914
rect 1865 9909 1866 9913
rect 1870 9909 1871 9913
rect 1875 9909 1876 9913
rect 1880 9909 1881 9913
rect 1885 9909 1886 9913
rect 1890 9909 1891 9913
rect 1895 9909 1896 9913
rect 1900 9909 1901 9913
rect 1905 9909 1906 9913
rect 1865 9908 1910 9909
rect 1865 9904 1866 9908
rect 1870 9904 1871 9908
rect 1875 9904 1876 9908
rect 1880 9904 1881 9908
rect 1885 9904 1886 9908
rect 1890 9904 1891 9908
rect 1895 9904 1896 9908
rect 1900 9904 1901 9908
rect 1905 9904 1906 9908
rect 1865 9903 1910 9904
rect 1865 9899 1866 9903
rect 1870 9899 1871 9903
rect 1875 9899 1876 9903
rect 1880 9899 1881 9903
rect 1885 9899 1886 9903
rect 1890 9899 1891 9903
rect 1895 9899 1896 9903
rect 1900 9899 1901 9903
rect 1905 9899 1906 9903
rect 1865 9898 1910 9899
rect 1865 9894 1866 9898
rect 1870 9894 1871 9898
rect 1875 9894 1876 9898
rect 1880 9894 1881 9898
rect 1885 9894 1886 9898
rect 1890 9894 1891 9898
rect 1895 9894 1896 9898
rect 1900 9894 1901 9898
rect 1905 9894 1906 9898
rect 1865 9893 1910 9894
rect 1865 9889 1866 9893
rect 1870 9889 1871 9893
rect 1875 9889 1876 9893
rect 1880 9889 1881 9893
rect 1885 9889 1886 9893
rect 1890 9889 1891 9893
rect 1895 9889 1896 9893
rect 1900 9889 1901 9893
rect 1905 9889 1906 9893
rect 1865 9888 1910 9889
rect 1865 9884 1866 9888
rect 1870 9884 1871 9888
rect 1875 9884 1876 9888
rect 1880 9884 1881 9888
rect 1885 9884 1886 9888
rect 1890 9884 1891 9888
rect 1895 9884 1896 9888
rect 1900 9884 1901 9888
rect 1905 9884 1906 9888
rect 1865 9883 1910 9884
rect 1865 9879 1866 9883
rect 1870 9879 1871 9883
rect 1875 9879 1876 9883
rect 1880 9879 1881 9883
rect 1885 9879 1886 9883
rect 1890 9879 1891 9883
rect 1895 9879 1896 9883
rect 1900 9879 1901 9883
rect 1905 9879 1906 9883
rect 1865 9878 1910 9879
rect 1865 9874 1866 9878
rect 1870 9874 1871 9878
rect 1875 9874 1876 9878
rect 1880 9874 1881 9878
rect 1885 9874 1886 9878
rect 1890 9874 1891 9878
rect 1895 9874 1896 9878
rect 1900 9874 1901 9878
rect 1905 9874 1906 9878
rect 1865 9873 1910 9874
rect 1865 9869 1866 9873
rect 1870 9869 1871 9873
rect 1875 9869 1876 9873
rect 1880 9869 1881 9873
rect 1885 9869 1886 9873
rect 1890 9869 1891 9873
rect 1895 9869 1896 9873
rect 1900 9869 1901 9873
rect 1905 9869 1906 9873
rect 1865 9868 1910 9869
rect 1865 9864 1866 9868
rect 1870 9864 1871 9868
rect 1875 9864 1876 9868
rect 1880 9864 1881 9868
rect 1885 9864 1886 9868
rect 1890 9864 1891 9868
rect 1895 9864 1896 9868
rect 1900 9864 1901 9868
rect 1905 9864 1906 9868
rect 1918 9948 1922 9949
rect 1918 9943 1922 9944
rect 1918 9938 1922 9939
rect 1918 9933 1922 9934
rect 1918 9928 1922 9929
rect 1918 9923 1922 9924
rect 1918 9918 1922 9919
rect 1918 9913 1922 9914
rect 1918 9908 1922 9909
rect 1918 9903 1922 9904
rect 1918 9898 1922 9899
rect 1918 9893 1922 9894
rect 1918 9888 1922 9889
rect 1918 9883 1922 9884
rect 1918 9878 1922 9879
rect 1918 9873 1922 9874
rect 1918 9868 1922 9869
rect 1854 9863 1858 9864
rect 1854 9856 1858 9859
rect 1918 9863 1922 9864
rect 1918 9856 1922 9859
rect 1858 9848 1861 9856
rect 1865 9848 1866 9856
rect 1870 9848 1871 9856
rect 1875 9848 1876 9856
rect 1880 9848 1881 9856
rect 1885 9848 1886 9856
rect 1890 9848 1891 9856
rect 1895 9848 1896 9856
rect 1900 9848 1901 9856
rect 1905 9848 1906 9856
rect 1910 9848 1911 9856
rect 1915 9848 1918 9856
rect 1931 9963 1935 9964
rect 1931 9958 1935 9959
rect 1931 9953 1935 9954
rect 1931 9948 1935 9949
rect 1931 9943 1935 9944
rect 1931 9938 1935 9939
rect 1931 9933 1935 9934
rect 1931 9928 1935 9929
rect 1931 9923 1935 9924
rect 1931 9918 1935 9919
rect 1931 9913 1935 9914
rect 1931 9908 1935 9909
rect 1931 9903 1935 9904
rect 1931 9898 1935 9899
rect 1931 9893 1935 9894
rect 1931 9888 1935 9889
rect 1931 9883 1935 9884
rect 1931 9878 1935 9879
rect 1931 9873 1935 9874
rect 1931 9868 1935 9869
rect 1931 9863 1935 9864
rect 1931 9858 1935 9859
rect 1931 9853 1935 9854
rect 1931 9848 1935 9849
rect 1799 9844 1816 9846
rect 1771 9843 1775 9844
rect 1685 9839 1686 9843
rect 1690 9839 1691 9843
rect 1695 9839 1696 9843
rect 1700 9839 1701 9843
rect 1705 9839 1706 9843
rect 1710 9839 1711 9843
rect 1715 9839 1716 9843
rect 1720 9839 1721 9843
rect 1725 9839 1726 9843
rect 1730 9839 1731 9843
rect 1735 9839 1736 9843
rect 1740 9839 1741 9843
rect 1745 9839 1746 9843
rect 1750 9839 1751 9843
rect 1755 9839 1756 9843
rect 1760 9839 1761 9843
rect 1765 9839 1766 9843
rect 1770 9839 1771 9843
rect 1801 9842 1814 9844
rect 1841 9843 1845 9844
rect 1931 9843 1935 9844
rect 1473 9711 1499 9715
rect 1503 9711 1504 9715
rect 1508 9711 1525 9715
rect 1569 9722 1625 9839
rect 1684 9831 1740 9839
rect 1803 9831 1812 9842
rect 1845 9839 1846 9843
rect 1850 9839 1851 9843
rect 1855 9839 1856 9843
rect 1860 9839 1861 9843
rect 1865 9839 1866 9843
rect 1870 9839 1871 9843
rect 1875 9839 1876 9843
rect 1880 9839 1881 9843
rect 1885 9839 1886 9843
rect 1890 9839 1891 9843
rect 1895 9839 1896 9843
rect 1900 9839 1901 9843
rect 1905 9839 1906 9843
rect 1910 9839 1911 9843
rect 1915 9839 1916 9843
rect 1920 9839 1921 9843
rect 1925 9839 1926 9843
rect 1930 9839 1931 9843
rect 1994 9974 1995 9978
rect 1999 9974 2000 9978
rect 2004 9974 2005 9978
rect 2009 9974 2010 9978
rect 2014 9974 2015 9978
rect 2019 9974 2020 9978
rect 2024 9974 2025 9978
rect 2029 9974 2030 9978
rect 2034 9974 2035 9978
rect 2039 9974 2040 9978
rect 2044 9974 2045 9978
rect 2049 9974 2050 9978
rect 2054 9974 2055 9978
rect 2059 9974 2060 9978
rect 2064 9974 2065 9978
rect 2069 9974 2070 9978
rect 2074 9974 2075 9978
rect 2079 9974 2080 9978
rect 1990 9973 1994 9974
rect 1990 9968 1994 9969
rect 2080 9973 2084 9974
rect 2080 9968 2084 9969
rect 1990 9963 1994 9964
rect 1990 9958 1994 9959
rect 1990 9953 1994 9954
rect 1990 9948 1994 9949
rect 1990 9943 1994 9944
rect 1990 9938 1994 9939
rect 1990 9933 1994 9934
rect 1990 9928 1994 9929
rect 1990 9923 1994 9924
rect 1990 9918 1994 9919
rect 1990 9913 1994 9914
rect 1990 9908 1994 9909
rect 1990 9903 1994 9904
rect 1990 9898 1994 9899
rect 1990 9893 1994 9894
rect 1990 9888 1994 9889
rect 1990 9883 1994 9884
rect 1990 9878 1994 9879
rect 1990 9873 1994 9874
rect 1990 9868 1994 9869
rect 1990 9863 1994 9864
rect 1990 9858 1994 9859
rect 1990 9853 1994 9854
rect 1990 9848 1994 9849
rect 2007 9961 2010 9965
rect 2014 9961 2015 9965
rect 2019 9961 2020 9965
rect 2024 9961 2025 9965
rect 2029 9961 2030 9965
rect 2034 9961 2035 9965
rect 2039 9961 2040 9965
rect 2044 9961 2045 9965
rect 2049 9961 2050 9965
rect 2054 9961 2055 9965
rect 2059 9961 2060 9965
rect 2064 9961 2067 9965
rect 2003 9958 2007 9961
rect 2003 9953 2007 9954
rect 2067 9958 2071 9961
rect 2067 9953 2071 9954
rect 2003 9948 2007 9949
rect 2003 9943 2007 9944
rect 2003 9938 2007 9939
rect 2003 9933 2007 9934
rect 2003 9928 2007 9929
rect 2003 9923 2007 9924
rect 2003 9918 2007 9919
rect 2003 9913 2007 9914
rect 2003 9908 2007 9909
rect 2003 9903 2007 9904
rect 2003 9898 2007 9899
rect 2003 9893 2007 9894
rect 2003 9888 2007 9889
rect 2003 9883 2007 9884
rect 2003 9878 2007 9879
rect 2003 9873 2007 9874
rect 2003 9868 2007 9869
rect 2019 9949 2020 9953
rect 2024 9949 2025 9953
rect 2029 9949 2030 9953
rect 2034 9949 2035 9953
rect 2039 9949 2040 9953
rect 2044 9949 2045 9953
rect 2049 9949 2050 9953
rect 2054 9949 2055 9953
rect 2015 9948 2059 9949
rect 2019 9944 2020 9948
rect 2024 9944 2025 9948
rect 2029 9944 2030 9948
rect 2034 9944 2035 9948
rect 2039 9944 2040 9948
rect 2044 9944 2045 9948
rect 2049 9944 2050 9948
rect 2054 9944 2055 9948
rect 2015 9943 2059 9944
rect 2019 9939 2020 9943
rect 2024 9939 2025 9943
rect 2029 9939 2030 9943
rect 2034 9939 2035 9943
rect 2039 9939 2040 9943
rect 2044 9939 2045 9943
rect 2049 9939 2050 9943
rect 2054 9939 2055 9943
rect 2015 9938 2059 9939
rect 2019 9934 2020 9938
rect 2024 9934 2025 9938
rect 2029 9934 2030 9938
rect 2034 9934 2035 9938
rect 2039 9934 2040 9938
rect 2044 9934 2045 9938
rect 2049 9934 2050 9938
rect 2054 9934 2055 9938
rect 2015 9933 2059 9934
rect 2019 9929 2020 9933
rect 2024 9929 2025 9933
rect 2029 9929 2030 9933
rect 2034 9929 2035 9933
rect 2039 9929 2040 9933
rect 2044 9929 2045 9933
rect 2049 9929 2050 9933
rect 2054 9929 2055 9933
rect 2015 9928 2059 9929
rect 2019 9924 2020 9928
rect 2024 9924 2025 9928
rect 2029 9924 2030 9928
rect 2034 9924 2035 9928
rect 2039 9924 2040 9928
rect 2044 9924 2045 9928
rect 2049 9924 2050 9928
rect 2054 9924 2055 9928
rect 2015 9923 2059 9924
rect 2019 9919 2020 9923
rect 2024 9919 2025 9923
rect 2029 9919 2030 9923
rect 2034 9919 2035 9923
rect 2039 9919 2040 9923
rect 2044 9919 2045 9923
rect 2049 9919 2050 9923
rect 2054 9919 2055 9923
rect 2015 9918 2059 9919
rect 2019 9914 2020 9918
rect 2024 9914 2025 9918
rect 2029 9914 2030 9918
rect 2034 9914 2035 9918
rect 2039 9914 2040 9918
rect 2044 9914 2045 9918
rect 2049 9914 2050 9918
rect 2054 9914 2055 9918
rect 2015 9913 2059 9914
rect 2019 9909 2020 9913
rect 2024 9909 2025 9913
rect 2029 9909 2030 9913
rect 2034 9909 2035 9913
rect 2039 9909 2040 9913
rect 2044 9909 2045 9913
rect 2049 9909 2050 9913
rect 2054 9909 2055 9913
rect 2015 9908 2059 9909
rect 2019 9904 2020 9908
rect 2024 9904 2025 9908
rect 2029 9904 2030 9908
rect 2034 9904 2035 9908
rect 2039 9904 2040 9908
rect 2044 9904 2045 9908
rect 2049 9904 2050 9908
rect 2054 9904 2055 9908
rect 2015 9903 2059 9904
rect 2019 9899 2020 9903
rect 2024 9899 2025 9903
rect 2029 9899 2030 9903
rect 2034 9899 2035 9903
rect 2039 9899 2040 9903
rect 2044 9899 2045 9903
rect 2049 9899 2050 9903
rect 2054 9899 2055 9903
rect 2015 9898 2059 9899
rect 2019 9894 2020 9898
rect 2024 9894 2025 9898
rect 2029 9894 2030 9898
rect 2034 9894 2035 9898
rect 2039 9894 2040 9898
rect 2044 9894 2045 9898
rect 2049 9894 2050 9898
rect 2054 9894 2055 9898
rect 2015 9893 2059 9894
rect 2019 9889 2020 9893
rect 2024 9889 2025 9893
rect 2029 9889 2030 9893
rect 2034 9889 2035 9893
rect 2039 9889 2040 9893
rect 2044 9889 2045 9893
rect 2049 9889 2050 9893
rect 2054 9889 2055 9893
rect 2015 9888 2059 9889
rect 2019 9884 2020 9888
rect 2024 9884 2025 9888
rect 2029 9884 2030 9888
rect 2034 9884 2035 9888
rect 2039 9884 2040 9888
rect 2044 9884 2045 9888
rect 2049 9884 2050 9888
rect 2054 9884 2055 9888
rect 2015 9883 2059 9884
rect 2019 9879 2020 9883
rect 2024 9879 2025 9883
rect 2029 9879 2030 9883
rect 2034 9879 2035 9883
rect 2039 9879 2040 9883
rect 2044 9879 2045 9883
rect 2049 9879 2050 9883
rect 2054 9879 2055 9883
rect 2015 9878 2059 9879
rect 2019 9874 2020 9878
rect 2024 9874 2025 9878
rect 2029 9874 2030 9878
rect 2034 9874 2035 9878
rect 2039 9874 2040 9878
rect 2044 9874 2045 9878
rect 2049 9874 2050 9878
rect 2054 9874 2055 9878
rect 2015 9873 2059 9874
rect 2019 9869 2020 9873
rect 2024 9869 2025 9873
rect 2029 9869 2030 9873
rect 2034 9869 2035 9873
rect 2039 9869 2040 9873
rect 2044 9869 2045 9873
rect 2049 9869 2050 9873
rect 2054 9869 2055 9873
rect 2015 9868 2059 9869
rect 2019 9864 2020 9868
rect 2024 9864 2025 9868
rect 2029 9864 2030 9868
rect 2034 9864 2035 9868
rect 2039 9864 2040 9868
rect 2044 9864 2045 9868
rect 2049 9864 2050 9868
rect 2054 9864 2055 9868
rect 2067 9948 2071 9949
rect 2067 9943 2071 9944
rect 2067 9938 2071 9939
rect 2067 9933 2071 9934
rect 2067 9928 2071 9929
rect 2067 9923 2071 9924
rect 2067 9918 2071 9919
rect 2067 9913 2071 9914
rect 2067 9908 2071 9909
rect 2067 9903 2071 9904
rect 2067 9898 2071 9899
rect 2067 9893 2071 9894
rect 2067 9888 2071 9889
rect 2067 9883 2071 9884
rect 2067 9878 2071 9879
rect 2067 9873 2071 9874
rect 2067 9868 2071 9869
rect 2003 9863 2007 9864
rect 2003 9856 2007 9859
rect 2067 9863 2071 9864
rect 2067 9856 2071 9859
rect 2007 9848 2010 9856
rect 2014 9848 2015 9856
rect 2019 9848 2020 9856
rect 2024 9848 2025 9856
rect 2029 9848 2030 9856
rect 2034 9848 2035 9856
rect 2039 9848 2040 9856
rect 2044 9848 2045 9856
rect 2049 9848 2050 9856
rect 2054 9848 2055 9856
rect 2059 9848 2060 9856
rect 2064 9848 2067 9856
rect 2080 9963 2084 9964
rect 2080 9958 2084 9959
rect 2080 9953 2084 9954
rect 2106 9961 2127 9981
rect 2154 9974 2155 9978
rect 2159 9974 2160 9978
rect 2164 9974 2165 9978
rect 2169 9974 2170 9978
rect 2174 9974 2175 9978
rect 2179 9974 2180 9978
rect 2184 9974 2185 9978
rect 2189 9974 2190 9978
rect 2194 9974 2195 9978
rect 2199 9974 2200 9978
rect 2204 9974 2205 9978
rect 2209 9974 2210 9978
rect 2214 9974 2215 9978
rect 2219 9974 2220 9978
rect 2224 9974 2225 9978
rect 2229 9974 2230 9978
rect 2234 9974 2235 9978
rect 2239 9974 2240 9978
rect 2150 9973 2154 9974
rect 2150 9968 2154 9969
rect 2240 9973 2244 9974
rect 2240 9968 2244 9969
rect 2150 9963 2154 9964
rect 2150 9958 2154 9959
rect 2150 9953 2154 9954
rect 2080 9948 2084 9949
rect 2080 9943 2084 9944
rect 2080 9938 2084 9939
rect 2080 9933 2084 9934
rect 2080 9928 2084 9929
rect 2080 9923 2084 9924
rect 2080 9918 2084 9919
rect 2080 9913 2084 9914
rect 2080 9908 2084 9909
rect 2080 9903 2084 9904
rect 2080 9898 2084 9899
rect 2080 9893 2084 9894
rect 2080 9888 2084 9889
rect 2080 9883 2084 9884
rect 2150 9948 2154 9949
rect 2150 9943 2154 9944
rect 2150 9938 2154 9939
rect 2150 9933 2154 9934
rect 2150 9928 2154 9929
rect 2150 9923 2154 9924
rect 2150 9918 2154 9919
rect 2150 9913 2154 9914
rect 2150 9908 2154 9909
rect 2150 9903 2154 9904
rect 2150 9898 2154 9899
rect 2150 9893 2154 9894
rect 2150 9888 2154 9889
rect 2150 9883 2154 9884
rect 2080 9878 2084 9879
rect 2080 9873 2084 9874
rect 2080 9868 2084 9869
rect 2080 9863 2084 9864
rect 2080 9858 2084 9859
rect 2080 9853 2084 9854
rect 2080 9848 2084 9849
rect 1990 9843 1994 9844
rect 2106 9846 2127 9874
rect 2150 9878 2154 9879
rect 2150 9873 2154 9874
rect 2150 9868 2154 9869
rect 2150 9863 2154 9864
rect 2150 9858 2154 9859
rect 2150 9853 2154 9854
rect 2150 9848 2154 9849
rect 2167 9961 2170 9965
rect 2174 9961 2175 9965
rect 2179 9961 2180 9965
rect 2184 9961 2185 9965
rect 2189 9961 2190 9965
rect 2194 9961 2195 9965
rect 2199 9961 2200 9965
rect 2204 9961 2205 9965
rect 2209 9961 2210 9965
rect 2214 9961 2215 9965
rect 2219 9961 2220 9965
rect 2224 9961 2227 9965
rect 2163 9958 2167 9961
rect 2163 9953 2167 9954
rect 2227 9958 2231 9961
rect 2227 9953 2231 9954
rect 2163 9948 2167 9949
rect 2163 9943 2167 9944
rect 2163 9938 2167 9939
rect 2163 9933 2167 9934
rect 2163 9928 2167 9929
rect 2163 9923 2167 9924
rect 2163 9918 2167 9919
rect 2163 9913 2167 9914
rect 2163 9908 2167 9909
rect 2163 9903 2167 9904
rect 2163 9898 2167 9899
rect 2163 9893 2167 9894
rect 2163 9888 2167 9889
rect 2163 9883 2167 9884
rect 2163 9878 2167 9879
rect 2163 9873 2167 9874
rect 2163 9868 2167 9869
rect 2174 9949 2175 9953
rect 2179 9949 2180 9953
rect 2184 9949 2185 9953
rect 2189 9949 2190 9953
rect 2194 9949 2195 9953
rect 2199 9949 2200 9953
rect 2204 9949 2205 9953
rect 2209 9949 2210 9953
rect 2214 9949 2215 9953
rect 2174 9948 2219 9949
rect 2174 9944 2175 9948
rect 2179 9944 2180 9948
rect 2184 9944 2185 9948
rect 2189 9944 2190 9948
rect 2194 9944 2195 9948
rect 2199 9944 2200 9948
rect 2204 9944 2205 9948
rect 2209 9944 2210 9948
rect 2214 9944 2215 9948
rect 2174 9943 2219 9944
rect 2174 9939 2175 9943
rect 2179 9939 2180 9943
rect 2184 9939 2185 9943
rect 2189 9939 2190 9943
rect 2194 9939 2195 9943
rect 2199 9939 2200 9943
rect 2204 9939 2205 9943
rect 2209 9939 2210 9943
rect 2214 9939 2215 9943
rect 2174 9938 2219 9939
rect 2174 9934 2175 9938
rect 2179 9934 2180 9938
rect 2184 9934 2185 9938
rect 2189 9934 2190 9938
rect 2194 9934 2195 9938
rect 2199 9934 2200 9938
rect 2204 9934 2205 9938
rect 2209 9934 2210 9938
rect 2214 9934 2215 9938
rect 2174 9933 2219 9934
rect 2174 9929 2175 9933
rect 2179 9929 2180 9933
rect 2184 9929 2185 9933
rect 2189 9929 2190 9933
rect 2194 9929 2195 9933
rect 2199 9929 2200 9933
rect 2204 9929 2205 9933
rect 2209 9929 2210 9933
rect 2214 9929 2215 9933
rect 2174 9928 2219 9929
rect 2174 9924 2175 9928
rect 2179 9924 2180 9928
rect 2184 9924 2185 9928
rect 2189 9924 2190 9928
rect 2194 9924 2195 9928
rect 2199 9924 2200 9928
rect 2204 9924 2205 9928
rect 2209 9924 2210 9928
rect 2214 9924 2215 9928
rect 2174 9923 2219 9924
rect 2174 9919 2175 9923
rect 2179 9919 2180 9923
rect 2184 9919 2185 9923
rect 2189 9919 2190 9923
rect 2194 9919 2195 9923
rect 2199 9919 2200 9923
rect 2204 9919 2205 9923
rect 2209 9919 2210 9923
rect 2214 9919 2215 9923
rect 2174 9918 2219 9919
rect 2174 9914 2175 9918
rect 2179 9914 2180 9918
rect 2184 9914 2185 9918
rect 2189 9914 2190 9918
rect 2194 9914 2195 9918
rect 2199 9914 2200 9918
rect 2204 9914 2205 9918
rect 2209 9914 2210 9918
rect 2214 9914 2215 9918
rect 2174 9913 2219 9914
rect 2174 9909 2175 9913
rect 2179 9909 2180 9913
rect 2184 9909 2185 9913
rect 2189 9909 2190 9913
rect 2194 9909 2195 9913
rect 2199 9909 2200 9913
rect 2204 9909 2205 9913
rect 2209 9909 2210 9913
rect 2214 9909 2215 9913
rect 2174 9908 2219 9909
rect 2174 9904 2175 9908
rect 2179 9904 2180 9908
rect 2184 9904 2185 9908
rect 2189 9904 2190 9908
rect 2194 9904 2195 9908
rect 2199 9904 2200 9908
rect 2204 9904 2205 9908
rect 2209 9904 2210 9908
rect 2214 9904 2215 9908
rect 2174 9903 2219 9904
rect 2174 9899 2175 9903
rect 2179 9899 2180 9903
rect 2184 9899 2185 9903
rect 2189 9899 2190 9903
rect 2194 9899 2195 9903
rect 2199 9899 2200 9903
rect 2204 9899 2205 9903
rect 2209 9899 2210 9903
rect 2214 9899 2215 9903
rect 2174 9898 2219 9899
rect 2174 9894 2175 9898
rect 2179 9894 2180 9898
rect 2184 9894 2185 9898
rect 2189 9894 2190 9898
rect 2194 9894 2195 9898
rect 2199 9894 2200 9898
rect 2204 9894 2205 9898
rect 2209 9894 2210 9898
rect 2214 9894 2215 9898
rect 2174 9893 2219 9894
rect 2174 9889 2175 9893
rect 2179 9889 2180 9893
rect 2184 9889 2185 9893
rect 2189 9889 2190 9893
rect 2194 9889 2195 9893
rect 2199 9889 2200 9893
rect 2204 9889 2205 9893
rect 2209 9889 2210 9893
rect 2214 9889 2215 9893
rect 2174 9888 2219 9889
rect 2174 9884 2175 9888
rect 2179 9884 2180 9888
rect 2184 9884 2185 9888
rect 2189 9884 2190 9888
rect 2194 9884 2195 9888
rect 2199 9884 2200 9888
rect 2204 9884 2205 9888
rect 2209 9884 2210 9888
rect 2214 9884 2215 9888
rect 2174 9883 2219 9884
rect 2174 9879 2175 9883
rect 2179 9879 2180 9883
rect 2184 9879 2185 9883
rect 2189 9879 2190 9883
rect 2194 9879 2195 9883
rect 2199 9879 2200 9883
rect 2204 9879 2205 9883
rect 2209 9879 2210 9883
rect 2214 9879 2215 9883
rect 2174 9878 2219 9879
rect 2174 9874 2175 9878
rect 2179 9874 2180 9878
rect 2184 9874 2185 9878
rect 2189 9874 2190 9878
rect 2194 9874 2195 9878
rect 2199 9874 2200 9878
rect 2204 9874 2205 9878
rect 2209 9874 2210 9878
rect 2214 9874 2215 9878
rect 2174 9873 2219 9874
rect 2174 9869 2175 9873
rect 2179 9869 2180 9873
rect 2184 9869 2185 9873
rect 2189 9869 2190 9873
rect 2194 9869 2195 9873
rect 2199 9869 2200 9873
rect 2204 9869 2205 9873
rect 2209 9869 2210 9873
rect 2214 9869 2215 9873
rect 2174 9868 2219 9869
rect 2174 9864 2175 9868
rect 2179 9864 2180 9868
rect 2184 9864 2185 9868
rect 2189 9864 2190 9868
rect 2194 9864 2195 9868
rect 2199 9864 2200 9868
rect 2204 9864 2205 9868
rect 2209 9864 2210 9868
rect 2214 9864 2215 9868
rect 2227 9948 2231 9949
rect 2227 9943 2231 9944
rect 2227 9938 2231 9939
rect 2227 9933 2231 9934
rect 2227 9928 2231 9929
rect 2227 9923 2231 9924
rect 2227 9918 2231 9919
rect 2227 9913 2231 9914
rect 2227 9908 2231 9909
rect 2227 9903 2231 9904
rect 2227 9898 2231 9899
rect 2227 9893 2231 9894
rect 2227 9888 2231 9889
rect 2227 9883 2231 9884
rect 2227 9878 2231 9879
rect 2227 9873 2231 9874
rect 2227 9868 2231 9869
rect 2163 9863 2167 9864
rect 2163 9856 2167 9859
rect 2227 9863 2231 9864
rect 2227 9856 2231 9859
rect 2167 9848 2170 9856
rect 2174 9848 2175 9856
rect 2179 9848 2180 9856
rect 2184 9848 2185 9856
rect 2189 9848 2190 9856
rect 2194 9848 2195 9856
rect 2199 9848 2200 9856
rect 2204 9848 2205 9856
rect 2209 9848 2210 9856
rect 2214 9848 2215 9856
rect 2219 9848 2220 9856
rect 2224 9848 2227 9856
rect 2240 9963 2244 9964
rect 2240 9958 2244 9959
rect 2240 9953 2244 9954
rect 2240 9948 2244 9949
rect 2240 9943 2244 9944
rect 2240 9938 2244 9939
rect 2240 9933 2244 9934
rect 2240 9928 2244 9929
rect 2240 9923 2244 9924
rect 2240 9918 2244 9919
rect 2240 9913 2244 9914
rect 2240 9908 2244 9909
rect 2240 9903 2244 9904
rect 2240 9898 2244 9899
rect 2240 9893 2244 9894
rect 2240 9888 2244 9889
rect 2240 9883 2244 9884
rect 2240 9878 2244 9879
rect 2240 9873 2244 9874
rect 2240 9868 2244 9869
rect 2240 9863 2244 9864
rect 2240 9858 2244 9859
rect 2240 9853 2244 9854
rect 2240 9848 2244 9849
rect 2108 9844 2125 9846
rect 2080 9843 2084 9844
rect 1994 9839 1995 9843
rect 1999 9839 2000 9843
rect 2004 9839 2005 9843
rect 2009 9839 2010 9843
rect 2014 9839 2015 9843
rect 2019 9839 2020 9843
rect 2024 9839 2025 9843
rect 2029 9839 2030 9843
rect 2034 9839 2035 9843
rect 2039 9839 2040 9843
rect 2044 9839 2045 9843
rect 2049 9839 2050 9843
rect 2054 9839 2055 9843
rect 2059 9839 2060 9843
rect 2064 9839 2065 9843
rect 2069 9839 2070 9843
rect 2074 9839 2075 9843
rect 2079 9839 2080 9843
rect 2110 9842 2123 9844
rect 2150 9843 2154 9844
rect 2240 9843 2244 9844
rect 1878 9831 1934 9839
rect 1684 9827 1743 9831
rect 1869 9827 1934 9831
rect 1684 9815 1740 9827
rect 1799 9819 1829 9823
rect 1684 9811 1743 9815
rect 1813 9812 1817 9819
rect 1878 9815 1934 9827
rect 1684 9802 1740 9811
rect 1869 9811 1934 9815
rect 1799 9803 1810 9807
rect 1672 9800 1740 9802
rect 1672 9796 1673 9800
rect 1677 9796 1678 9800
rect 1682 9799 1740 9800
rect 1803 9800 1810 9803
rect 1822 9803 1829 9807
rect 1822 9800 1826 9803
rect 1682 9796 1743 9799
rect 1672 9795 1743 9796
rect 1672 9791 1673 9795
rect 1677 9791 1678 9795
rect 1682 9791 1740 9795
rect 1803 9791 1826 9800
rect 1878 9799 1934 9811
rect 1993 9831 2049 9839
rect 2112 9831 2121 9842
rect 2154 9839 2155 9843
rect 2159 9839 2160 9843
rect 2164 9839 2165 9843
rect 2169 9839 2170 9843
rect 2174 9839 2175 9843
rect 2179 9839 2180 9843
rect 2184 9839 2185 9843
rect 2189 9839 2190 9843
rect 2194 9839 2195 9843
rect 2199 9839 2200 9843
rect 2204 9839 2205 9843
rect 2209 9839 2210 9843
rect 2214 9839 2215 9843
rect 2219 9839 2220 9843
rect 2224 9839 2225 9843
rect 2229 9839 2230 9843
rect 2234 9839 2235 9843
rect 2239 9839 2240 9843
rect 2303 9974 2304 9978
rect 2308 9974 2309 9978
rect 2313 9974 2314 9978
rect 2318 9974 2319 9978
rect 2323 9974 2324 9978
rect 2328 9974 2329 9978
rect 2333 9974 2334 9978
rect 2338 9974 2339 9978
rect 2343 9974 2344 9978
rect 2348 9974 2349 9978
rect 2353 9974 2354 9978
rect 2358 9974 2359 9978
rect 2363 9974 2364 9978
rect 2368 9974 2369 9978
rect 2373 9974 2374 9978
rect 2378 9974 2379 9978
rect 2383 9974 2384 9978
rect 2388 9974 2389 9978
rect 2299 9973 2303 9974
rect 2299 9968 2303 9969
rect 2389 9973 2393 9974
rect 2389 9968 2393 9969
rect 2299 9963 2303 9964
rect 2299 9958 2303 9959
rect 2299 9953 2303 9954
rect 2299 9948 2303 9949
rect 2299 9943 2303 9944
rect 2299 9938 2303 9939
rect 2299 9933 2303 9934
rect 2299 9928 2303 9929
rect 2299 9923 2303 9924
rect 2299 9918 2303 9919
rect 2299 9913 2303 9914
rect 2299 9908 2303 9909
rect 2299 9903 2303 9904
rect 2299 9898 2303 9899
rect 2299 9893 2303 9894
rect 2299 9888 2303 9889
rect 2299 9883 2303 9884
rect 2299 9878 2303 9879
rect 2299 9873 2303 9874
rect 2299 9868 2303 9869
rect 2299 9863 2303 9864
rect 2299 9858 2303 9859
rect 2299 9853 2303 9854
rect 2299 9848 2303 9849
rect 2316 9961 2319 9965
rect 2323 9961 2324 9965
rect 2328 9961 2329 9965
rect 2333 9961 2334 9965
rect 2338 9961 2339 9965
rect 2343 9961 2344 9965
rect 2348 9961 2349 9965
rect 2353 9961 2354 9965
rect 2358 9961 2359 9965
rect 2363 9961 2364 9965
rect 2368 9961 2369 9965
rect 2373 9961 2376 9965
rect 2312 9958 2316 9961
rect 2312 9953 2316 9954
rect 2376 9958 2380 9961
rect 2376 9953 2380 9954
rect 2312 9948 2316 9949
rect 2312 9943 2316 9944
rect 2312 9938 2316 9939
rect 2312 9933 2316 9934
rect 2312 9928 2316 9929
rect 2312 9923 2316 9924
rect 2312 9918 2316 9919
rect 2312 9913 2316 9914
rect 2312 9908 2316 9909
rect 2312 9903 2316 9904
rect 2312 9898 2316 9899
rect 2312 9893 2316 9894
rect 2312 9888 2316 9889
rect 2312 9883 2316 9884
rect 2312 9878 2316 9879
rect 2312 9873 2316 9874
rect 2312 9868 2316 9869
rect 2328 9949 2329 9953
rect 2333 9949 2334 9953
rect 2338 9949 2339 9953
rect 2343 9949 2344 9953
rect 2348 9949 2349 9953
rect 2353 9949 2354 9953
rect 2358 9949 2359 9953
rect 2363 9949 2364 9953
rect 2324 9948 2368 9949
rect 2328 9944 2329 9948
rect 2333 9944 2334 9948
rect 2338 9944 2339 9948
rect 2343 9944 2344 9948
rect 2348 9944 2349 9948
rect 2353 9944 2354 9948
rect 2358 9944 2359 9948
rect 2363 9944 2364 9948
rect 2324 9943 2368 9944
rect 2328 9939 2329 9943
rect 2333 9939 2334 9943
rect 2338 9939 2339 9943
rect 2343 9939 2344 9943
rect 2348 9939 2349 9943
rect 2353 9939 2354 9943
rect 2358 9939 2359 9943
rect 2363 9939 2364 9943
rect 2324 9938 2368 9939
rect 2328 9934 2329 9938
rect 2333 9934 2334 9938
rect 2338 9934 2339 9938
rect 2343 9934 2344 9938
rect 2348 9934 2349 9938
rect 2353 9934 2354 9938
rect 2358 9934 2359 9938
rect 2363 9934 2364 9938
rect 2324 9933 2368 9934
rect 2328 9929 2329 9933
rect 2333 9929 2334 9933
rect 2338 9929 2339 9933
rect 2343 9929 2344 9933
rect 2348 9929 2349 9933
rect 2353 9929 2354 9933
rect 2358 9929 2359 9933
rect 2363 9929 2364 9933
rect 2324 9928 2368 9929
rect 2328 9924 2329 9928
rect 2333 9924 2334 9928
rect 2338 9924 2339 9928
rect 2343 9924 2344 9928
rect 2348 9924 2349 9928
rect 2353 9924 2354 9928
rect 2358 9924 2359 9928
rect 2363 9924 2364 9928
rect 2324 9923 2368 9924
rect 2328 9919 2329 9923
rect 2333 9919 2334 9923
rect 2338 9919 2339 9923
rect 2343 9919 2344 9923
rect 2348 9919 2349 9923
rect 2353 9919 2354 9923
rect 2358 9919 2359 9923
rect 2363 9919 2364 9923
rect 2324 9918 2368 9919
rect 2328 9914 2329 9918
rect 2333 9914 2334 9918
rect 2338 9914 2339 9918
rect 2343 9914 2344 9918
rect 2348 9914 2349 9918
rect 2353 9914 2354 9918
rect 2358 9914 2359 9918
rect 2363 9914 2364 9918
rect 2324 9913 2368 9914
rect 2328 9909 2329 9913
rect 2333 9909 2334 9913
rect 2338 9909 2339 9913
rect 2343 9909 2344 9913
rect 2348 9909 2349 9913
rect 2353 9909 2354 9913
rect 2358 9909 2359 9913
rect 2363 9909 2364 9913
rect 2324 9908 2368 9909
rect 2328 9904 2329 9908
rect 2333 9904 2334 9908
rect 2338 9904 2339 9908
rect 2343 9904 2344 9908
rect 2348 9904 2349 9908
rect 2353 9904 2354 9908
rect 2358 9904 2359 9908
rect 2363 9904 2364 9908
rect 2324 9903 2368 9904
rect 2328 9899 2329 9903
rect 2333 9899 2334 9903
rect 2338 9899 2339 9903
rect 2343 9899 2344 9903
rect 2348 9899 2349 9903
rect 2353 9899 2354 9903
rect 2358 9899 2359 9903
rect 2363 9899 2364 9903
rect 2324 9898 2368 9899
rect 2328 9894 2329 9898
rect 2333 9894 2334 9898
rect 2338 9894 2339 9898
rect 2343 9894 2344 9898
rect 2348 9894 2349 9898
rect 2353 9894 2354 9898
rect 2358 9894 2359 9898
rect 2363 9894 2364 9898
rect 2324 9893 2368 9894
rect 2328 9889 2329 9893
rect 2333 9889 2334 9893
rect 2338 9889 2339 9893
rect 2343 9889 2344 9893
rect 2348 9889 2349 9893
rect 2353 9889 2354 9893
rect 2358 9889 2359 9893
rect 2363 9889 2364 9893
rect 2324 9888 2368 9889
rect 2328 9884 2329 9888
rect 2333 9884 2334 9888
rect 2338 9884 2339 9888
rect 2343 9884 2344 9888
rect 2348 9884 2349 9888
rect 2353 9884 2354 9888
rect 2358 9884 2359 9888
rect 2363 9884 2364 9888
rect 2324 9883 2368 9884
rect 2328 9879 2329 9883
rect 2333 9879 2334 9883
rect 2338 9879 2339 9883
rect 2343 9879 2344 9883
rect 2348 9879 2349 9883
rect 2353 9879 2354 9883
rect 2358 9879 2359 9883
rect 2363 9879 2364 9883
rect 2324 9878 2368 9879
rect 2328 9874 2329 9878
rect 2333 9874 2334 9878
rect 2338 9874 2339 9878
rect 2343 9874 2344 9878
rect 2348 9874 2349 9878
rect 2353 9874 2354 9878
rect 2358 9874 2359 9878
rect 2363 9874 2364 9878
rect 2324 9873 2368 9874
rect 2328 9869 2329 9873
rect 2333 9869 2334 9873
rect 2338 9869 2339 9873
rect 2343 9869 2344 9873
rect 2348 9869 2349 9873
rect 2353 9869 2354 9873
rect 2358 9869 2359 9873
rect 2363 9869 2364 9873
rect 2324 9868 2368 9869
rect 2328 9864 2329 9868
rect 2333 9864 2334 9868
rect 2338 9864 2339 9868
rect 2343 9864 2344 9868
rect 2348 9864 2349 9868
rect 2353 9864 2354 9868
rect 2358 9864 2359 9868
rect 2363 9864 2364 9868
rect 2376 9948 2380 9949
rect 2376 9943 2380 9944
rect 2376 9938 2380 9939
rect 2376 9933 2380 9934
rect 2376 9928 2380 9929
rect 2376 9923 2380 9924
rect 2376 9918 2380 9919
rect 2376 9913 2380 9914
rect 2376 9908 2380 9909
rect 2376 9903 2380 9904
rect 2376 9898 2380 9899
rect 2376 9893 2380 9894
rect 2376 9888 2380 9889
rect 2376 9883 2380 9884
rect 2376 9878 2380 9879
rect 2376 9873 2380 9874
rect 2376 9868 2380 9869
rect 2312 9863 2316 9864
rect 2312 9856 2316 9859
rect 2376 9863 2380 9864
rect 2376 9856 2380 9859
rect 2316 9848 2319 9856
rect 2323 9848 2324 9856
rect 2328 9848 2329 9856
rect 2333 9848 2334 9856
rect 2338 9848 2339 9856
rect 2343 9848 2344 9856
rect 2348 9848 2349 9856
rect 2353 9848 2354 9856
rect 2358 9848 2359 9856
rect 2363 9848 2364 9856
rect 2368 9848 2369 9856
rect 2373 9848 2376 9856
rect 2389 9963 2393 9964
rect 2389 9958 2393 9959
rect 2389 9953 2393 9954
rect 2415 9961 2436 9981
rect 2463 9974 2464 9978
rect 2468 9974 2469 9978
rect 2473 9974 2474 9978
rect 2478 9974 2479 9978
rect 2483 9974 2484 9978
rect 2488 9974 2489 9978
rect 2493 9974 2494 9978
rect 2498 9974 2499 9978
rect 2503 9974 2504 9978
rect 2508 9974 2509 9978
rect 2513 9974 2514 9978
rect 2518 9974 2519 9978
rect 2523 9974 2524 9978
rect 2528 9974 2529 9978
rect 2533 9974 2534 9978
rect 2538 9974 2539 9978
rect 2543 9974 2544 9978
rect 2548 9974 2549 9978
rect 2459 9973 2463 9974
rect 2459 9968 2463 9969
rect 2549 9973 2553 9974
rect 2549 9968 2553 9969
rect 2459 9963 2463 9964
rect 2459 9958 2463 9959
rect 2459 9953 2463 9954
rect 2389 9948 2393 9949
rect 2389 9943 2393 9944
rect 2389 9938 2393 9939
rect 2389 9933 2393 9934
rect 2389 9928 2393 9929
rect 2389 9923 2393 9924
rect 2389 9918 2393 9919
rect 2389 9913 2393 9914
rect 2389 9908 2393 9909
rect 2389 9903 2393 9904
rect 2389 9898 2393 9899
rect 2389 9893 2393 9894
rect 2389 9888 2393 9889
rect 2389 9883 2393 9884
rect 2459 9948 2463 9949
rect 2459 9943 2463 9944
rect 2459 9938 2463 9939
rect 2459 9933 2463 9934
rect 2459 9928 2463 9929
rect 2459 9923 2463 9924
rect 2459 9918 2463 9919
rect 2459 9913 2463 9914
rect 2459 9908 2463 9909
rect 2459 9903 2463 9904
rect 2459 9898 2463 9899
rect 2459 9893 2463 9894
rect 2459 9888 2463 9889
rect 2459 9883 2463 9884
rect 2389 9878 2393 9879
rect 2389 9873 2393 9874
rect 2389 9868 2393 9869
rect 2389 9863 2393 9864
rect 2389 9858 2393 9859
rect 2389 9853 2393 9854
rect 2389 9848 2393 9849
rect 2299 9843 2303 9844
rect 2415 9846 2436 9874
rect 2459 9878 2463 9879
rect 2459 9873 2463 9874
rect 2459 9868 2463 9869
rect 2459 9863 2463 9864
rect 2459 9858 2463 9859
rect 2459 9853 2463 9854
rect 2459 9848 2463 9849
rect 2476 9961 2479 9965
rect 2483 9961 2484 9965
rect 2488 9961 2489 9965
rect 2493 9961 2494 9965
rect 2498 9961 2499 9965
rect 2503 9961 2504 9965
rect 2508 9961 2509 9965
rect 2513 9961 2514 9965
rect 2518 9961 2519 9965
rect 2523 9961 2524 9965
rect 2528 9961 2529 9965
rect 2533 9961 2536 9965
rect 2472 9958 2476 9961
rect 2472 9953 2476 9954
rect 2536 9958 2540 9961
rect 2536 9953 2540 9954
rect 2472 9948 2476 9949
rect 2472 9943 2476 9944
rect 2472 9938 2476 9939
rect 2472 9933 2476 9934
rect 2472 9928 2476 9929
rect 2472 9923 2476 9924
rect 2472 9918 2476 9919
rect 2472 9913 2476 9914
rect 2472 9908 2476 9909
rect 2472 9903 2476 9904
rect 2472 9898 2476 9899
rect 2472 9893 2476 9894
rect 2472 9888 2476 9889
rect 2472 9883 2476 9884
rect 2472 9878 2476 9879
rect 2472 9873 2476 9874
rect 2472 9868 2476 9869
rect 2483 9949 2484 9953
rect 2488 9949 2489 9953
rect 2493 9949 2494 9953
rect 2498 9949 2499 9953
rect 2503 9949 2504 9953
rect 2508 9949 2509 9953
rect 2513 9949 2514 9953
rect 2518 9949 2519 9953
rect 2523 9949 2524 9953
rect 2483 9948 2528 9949
rect 2483 9944 2484 9948
rect 2488 9944 2489 9948
rect 2493 9944 2494 9948
rect 2498 9944 2499 9948
rect 2503 9944 2504 9948
rect 2508 9944 2509 9948
rect 2513 9944 2514 9948
rect 2518 9944 2519 9948
rect 2523 9944 2524 9948
rect 2483 9943 2528 9944
rect 2483 9939 2484 9943
rect 2488 9939 2489 9943
rect 2493 9939 2494 9943
rect 2498 9939 2499 9943
rect 2503 9939 2504 9943
rect 2508 9939 2509 9943
rect 2513 9939 2514 9943
rect 2518 9939 2519 9943
rect 2523 9939 2524 9943
rect 2483 9938 2528 9939
rect 2483 9934 2484 9938
rect 2488 9934 2489 9938
rect 2493 9934 2494 9938
rect 2498 9934 2499 9938
rect 2503 9934 2504 9938
rect 2508 9934 2509 9938
rect 2513 9934 2514 9938
rect 2518 9934 2519 9938
rect 2523 9934 2524 9938
rect 2483 9933 2528 9934
rect 2483 9929 2484 9933
rect 2488 9929 2489 9933
rect 2493 9929 2494 9933
rect 2498 9929 2499 9933
rect 2503 9929 2504 9933
rect 2508 9929 2509 9933
rect 2513 9929 2514 9933
rect 2518 9929 2519 9933
rect 2523 9929 2524 9933
rect 2483 9928 2528 9929
rect 2483 9924 2484 9928
rect 2488 9924 2489 9928
rect 2493 9924 2494 9928
rect 2498 9924 2499 9928
rect 2503 9924 2504 9928
rect 2508 9924 2509 9928
rect 2513 9924 2514 9928
rect 2518 9924 2519 9928
rect 2523 9924 2524 9928
rect 2483 9923 2528 9924
rect 2483 9919 2484 9923
rect 2488 9919 2489 9923
rect 2493 9919 2494 9923
rect 2498 9919 2499 9923
rect 2503 9919 2504 9923
rect 2508 9919 2509 9923
rect 2513 9919 2514 9923
rect 2518 9919 2519 9923
rect 2523 9919 2524 9923
rect 2483 9918 2528 9919
rect 2483 9914 2484 9918
rect 2488 9914 2489 9918
rect 2493 9914 2494 9918
rect 2498 9914 2499 9918
rect 2503 9914 2504 9918
rect 2508 9914 2509 9918
rect 2513 9914 2514 9918
rect 2518 9914 2519 9918
rect 2523 9914 2524 9918
rect 2483 9913 2528 9914
rect 2483 9909 2484 9913
rect 2488 9909 2489 9913
rect 2493 9909 2494 9913
rect 2498 9909 2499 9913
rect 2503 9909 2504 9913
rect 2508 9909 2509 9913
rect 2513 9909 2514 9913
rect 2518 9909 2519 9913
rect 2523 9909 2524 9913
rect 2483 9908 2528 9909
rect 2483 9904 2484 9908
rect 2488 9904 2489 9908
rect 2493 9904 2494 9908
rect 2498 9904 2499 9908
rect 2503 9904 2504 9908
rect 2508 9904 2509 9908
rect 2513 9904 2514 9908
rect 2518 9904 2519 9908
rect 2523 9904 2524 9908
rect 2483 9903 2528 9904
rect 2483 9899 2484 9903
rect 2488 9899 2489 9903
rect 2493 9899 2494 9903
rect 2498 9899 2499 9903
rect 2503 9899 2504 9903
rect 2508 9899 2509 9903
rect 2513 9899 2514 9903
rect 2518 9899 2519 9903
rect 2523 9899 2524 9903
rect 2483 9898 2528 9899
rect 2483 9894 2484 9898
rect 2488 9894 2489 9898
rect 2493 9894 2494 9898
rect 2498 9894 2499 9898
rect 2503 9894 2504 9898
rect 2508 9894 2509 9898
rect 2513 9894 2514 9898
rect 2518 9894 2519 9898
rect 2523 9894 2524 9898
rect 2483 9893 2528 9894
rect 2483 9889 2484 9893
rect 2488 9889 2489 9893
rect 2493 9889 2494 9893
rect 2498 9889 2499 9893
rect 2503 9889 2504 9893
rect 2508 9889 2509 9893
rect 2513 9889 2514 9893
rect 2518 9889 2519 9893
rect 2523 9889 2524 9893
rect 2483 9888 2528 9889
rect 2483 9884 2484 9888
rect 2488 9884 2489 9888
rect 2493 9884 2494 9888
rect 2498 9884 2499 9888
rect 2503 9884 2504 9888
rect 2508 9884 2509 9888
rect 2513 9884 2514 9888
rect 2518 9884 2519 9888
rect 2523 9884 2524 9888
rect 2483 9883 2528 9884
rect 2483 9879 2484 9883
rect 2488 9879 2489 9883
rect 2493 9879 2494 9883
rect 2498 9879 2499 9883
rect 2503 9879 2504 9883
rect 2508 9879 2509 9883
rect 2513 9879 2514 9883
rect 2518 9879 2519 9883
rect 2523 9879 2524 9883
rect 2483 9878 2528 9879
rect 2483 9874 2484 9878
rect 2488 9874 2489 9878
rect 2493 9874 2494 9878
rect 2498 9874 2499 9878
rect 2503 9874 2504 9878
rect 2508 9874 2509 9878
rect 2513 9874 2514 9878
rect 2518 9874 2519 9878
rect 2523 9874 2524 9878
rect 2483 9873 2528 9874
rect 2483 9869 2484 9873
rect 2488 9869 2489 9873
rect 2493 9869 2494 9873
rect 2498 9869 2499 9873
rect 2503 9869 2504 9873
rect 2508 9869 2509 9873
rect 2513 9869 2514 9873
rect 2518 9869 2519 9873
rect 2523 9869 2524 9873
rect 2483 9868 2528 9869
rect 2483 9864 2484 9868
rect 2488 9864 2489 9868
rect 2493 9864 2494 9868
rect 2498 9864 2499 9868
rect 2503 9864 2504 9868
rect 2508 9864 2509 9868
rect 2513 9864 2514 9868
rect 2518 9864 2519 9868
rect 2523 9864 2524 9868
rect 2536 9948 2540 9949
rect 2536 9943 2540 9944
rect 2536 9938 2540 9939
rect 2536 9933 2540 9934
rect 2536 9928 2540 9929
rect 2536 9923 2540 9924
rect 2536 9918 2540 9919
rect 2536 9913 2540 9914
rect 2536 9908 2540 9909
rect 2536 9903 2540 9904
rect 2536 9898 2540 9899
rect 2536 9893 2540 9894
rect 2536 9888 2540 9889
rect 2536 9883 2540 9884
rect 2536 9878 2540 9879
rect 2536 9873 2540 9874
rect 2536 9868 2540 9869
rect 2472 9863 2476 9864
rect 2472 9856 2476 9859
rect 2536 9863 2540 9864
rect 2536 9856 2540 9859
rect 2476 9848 2479 9856
rect 2483 9848 2484 9856
rect 2488 9848 2489 9856
rect 2493 9848 2494 9856
rect 2498 9848 2499 9856
rect 2503 9848 2504 9856
rect 2508 9848 2509 9856
rect 2513 9848 2514 9856
rect 2518 9848 2519 9856
rect 2523 9848 2524 9856
rect 2528 9848 2529 9856
rect 2533 9848 2536 9856
rect 2549 9963 2553 9964
rect 2549 9958 2553 9959
rect 2549 9953 2553 9954
rect 2549 9948 2553 9949
rect 2549 9943 2553 9944
rect 2549 9938 2553 9939
rect 2549 9933 2553 9934
rect 2549 9928 2553 9929
rect 2549 9923 2553 9924
rect 2549 9918 2553 9919
rect 2549 9913 2553 9914
rect 2549 9908 2553 9909
rect 2549 9903 2553 9904
rect 2549 9898 2553 9899
rect 2549 9893 2553 9894
rect 2549 9888 2553 9889
rect 2549 9883 2553 9884
rect 2549 9878 2553 9879
rect 2549 9873 2553 9874
rect 2549 9868 2553 9869
rect 2549 9863 2553 9864
rect 2549 9858 2553 9859
rect 2549 9853 2553 9854
rect 2549 9848 2553 9849
rect 2417 9844 2434 9846
rect 2389 9843 2393 9844
rect 2303 9839 2304 9843
rect 2308 9839 2309 9843
rect 2313 9839 2314 9843
rect 2318 9839 2319 9843
rect 2323 9839 2324 9843
rect 2328 9839 2329 9843
rect 2333 9839 2334 9843
rect 2338 9839 2339 9843
rect 2343 9839 2344 9843
rect 2348 9839 2349 9843
rect 2353 9839 2354 9843
rect 2358 9839 2359 9843
rect 2363 9839 2364 9843
rect 2368 9839 2369 9843
rect 2373 9839 2374 9843
rect 2378 9839 2379 9843
rect 2383 9839 2384 9843
rect 2388 9839 2389 9843
rect 2419 9842 2432 9844
rect 2459 9843 2463 9844
rect 2549 9843 2553 9844
rect 2187 9831 2243 9839
rect 1993 9827 2052 9831
rect 2178 9827 2243 9831
rect 1993 9815 2049 9827
rect 2108 9819 2138 9823
rect 1993 9811 2052 9815
rect 2122 9812 2126 9819
rect 2187 9815 2243 9827
rect 1993 9802 2049 9811
rect 2178 9811 2243 9815
rect 2108 9803 2119 9807
rect 1869 9795 1934 9799
rect 1672 9790 1740 9791
rect 1672 9786 1673 9790
rect 1677 9786 1678 9790
rect 1682 9786 1740 9790
rect 1799 9787 1829 9791
rect 1672 9785 1740 9786
rect 1672 9781 1673 9785
rect 1677 9781 1678 9785
rect 1682 9783 1740 9785
rect 1682 9781 1743 9783
rect 1672 9780 1743 9781
rect 1672 9776 1673 9780
rect 1677 9776 1678 9780
rect 1682 9779 1743 9780
rect 1682 9776 1740 9779
rect 1672 9775 1740 9776
rect 1672 9771 1673 9775
rect 1677 9771 1678 9775
rect 1682 9771 1740 9775
rect 1672 9770 1740 9771
rect 1672 9766 1673 9770
rect 1677 9766 1678 9770
rect 1682 9766 1740 9770
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1628 9761 1647 9762
rect 1632 9757 1633 9761
rect 1637 9757 1638 9761
rect 1642 9757 1643 9761
rect 1628 9756 1647 9757
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1628 9751 1647 9752
rect 1632 9747 1633 9751
rect 1637 9747 1638 9751
rect 1642 9747 1643 9751
rect 1628 9746 1647 9747
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1628 9741 1647 9742
rect 1632 9737 1633 9741
rect 1637 9737 1638 9741
rect 1642 9737 1643 9741
rect 1628 9736 1647 9737
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1672 9765 1740 9766
rect 1672 9761 1673 9765
rect 1677 9761 1678 9765
rect 1682 9761 1740 9765
rect 1672 9760 1740 9761
rect 1672 9756 1673 9760
rect 1677 9756 1678 9760
rect 1682 9756 1740 9760
rect 1672 9755 1740 9756
rect 1672 9751 1673 9755
rect 1677 9751 1678 9755
rect 1682 9751 1740 9755
rect 1672 9750 1740 9751
rect 1672 9746 1673 9750
rect 1677 9746 1678 9750
rect 1682 9746 1740 9750
rect 1672 9745 1740 9746
rect 1672 9741 1673 9745
rect 1677 9741 1678 9745
rect 1682 9741 1740 9745
rect 1672 9740 1740 9741
rect 1672 9736 1673 9740
rect 1677 9736 1678 9740
rect 1682 9736 1740 9740
rect 1672 9734 1740 9736
rect 1573 9718 1574 9722
rect 1578 9718 1579 9722
rect 1583 9718 1584 9722
rect 1588 9718 1589 9722
rect 1593 9718 1594 9722
rect 1598 9718 1599 9722
rect 1603 9718 1604 9722
rect 1608 9718 1609 9722
rect 1613 9718 1614 9722
rect 1618 9718 1619 9722
rect 1623 9718 1625 9722
rect 1569 9717 1625 9718
rect 1573 9713 1574 9717
rect 1578 9713 1579 9717
rect 1583 9713 1584 9717
rect 1588 9713 1589 9717
rect 1593 9713 1594 9717
rect 1598 9713 1599 9717
rect 1603 9713 1604 9717
rect 1608 9713 1609 9717
rect 1613 9713 1614 9717
rect 1618 9713 1619 9717
rect 1623 9713 1625 9717
rect 1569 9712 1625 9713
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1628 9715 1647 9716
rect 1473 9710 1525 9711
rect 1473 9706 1499 9710
rect 1503 9706 1504 9710
rect 1508 9706 1525 9710
rect 1473 9705 1525 9706
rect 1473 9701 1499 9705
rect 1503 9701 1504 9705
rect 1508 9701 1525 9705
rect 1473 9700 1525 9701
rect 1473 9696 1499 9700
rect 1503 9696 1504 9700
rect 1508 9696 1525 9700
rect 1473 9695 1525 9696
rect 1473 9691 1499 9695
rect 1503 9691 1504 9695
rect 1508 9691 1525 9695
rect 1473 9690 1525 9691
rect 1473 9686 1499 9690
rect 1503 9686 1504 9690
rect 1508 9686 1525 9690
rect 1632 9711 1633 9715
rect 1637 9711 1638 9715
rect 1642 9711 1643 9715
rect 1628 9710 1647 9711
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1628 9705 1647 9706
rect 1632 9701 1633 9705
rect 1637 9701 1638 9705
rect 1642 9701 1643 9705
rect 1628 9700 1647 9701
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1628 9695 1647 9696
rect 1632 9691 1633 9695
rect 1637 9691 1638 9695
rect 1642 9691 1643 9695
rect 1628 9690 1647 9691
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1473 9685 1525 9686
rect 1473 9681 1499 9685
rect 1503 9681 1504 9685
rect 1508 9681 1525 9685
rect 1473 9680 1525 9681
rect 1473 9676 1499 9680
rect 1503 9676 1504 9680
rect 1508 9676 1525 9680
rect 1473 9675 1525 9676
rect 1473 9671 1499 9675
rect 1503 9671 1504 9675
rect 1508 9671 1525 9675
rect 1473 9670 1525 9671
rect 1473 9666 1499 9670
rect 1503 9666 1504 9670
rect 1508 9666 1525 9670
rect 1473 9665 1525 9666
rect 1473 9661 1499 9665
rect 1503 9661 1504 9665
rect 1508 9661 1525 9665
rect 1473 9610 1525 9661
rect 659 9607 693 9608
rect 663 9603 664 9607
rect 668 9603 669 9607
rect 673 9603 674 9607
rect 678 9603 679 9607
rect 683 9603 684 9607
rect 688 9603 689 9607
rect 617 9592 618 9596
rect 622 9592 623 9596
rect 627 9592 628 9596
rect 632 9592 633 9596
rect 637 9592 638 9596
rect 642 9592 643 9596
rect 613 9591 647 9592
rect 617 9587 618 9591
rect 622 9587 623 9591
rect 627 9587 628 9591
rect 632 9587 633 9591
rect 637 9587 638 9591
rect 642 9587 643 9591
rect 613 9586 647 9587
rect 617 9582 618 9586
rect 622 9582 623 9586
rect 627 9582 628 9586
rect 632 9582 633 9586
rect 637 9582 638 9586
rect 642 9582 643 9586
rect 613 9581 647 9582
rect 617 9577 618 9581
rect 622 9577 623 9581
rect 627 9577 628 9581
rect 632 9577 633 9581
rect 637 9577 638 9581
rect 642 9577 643 9581
rect 663 9592 664 9596
rect 668 9592 669 9596
rect 673 9592 674 9596
rect 678 9592 679 9596
rect 683 9592 684 9596
rect 688 9592 689 9596
rect 1804 9593 1817 9787
rect 1878 9783 1934 9795
rect 1869 9779 1934 9783
rect 1878 9722 1934 9779
rect 1981 9800 2049 9802
rect 1981 9796 1982 9800
rect 1986 9796 1987 9800
rect 1991 9799 2049 9800
rect 2112 9800 2119 9803
rect 2131 9803 2138 9807
rect 2131 9800 2135 9803
rect 1991 9796 2052 9799
rect 1981 9795 2052 9796
rect 1981 9791 1982 9795
rect 1986 9791 1987 9795
rect 1991 9791 2049 9795
rect 2112 9791 2135 9800
rect 2187 9799 2243 9811
rect 2302 9831 2358 9839
rect 2421 9831 2430 9842
rect 2463 9839 2464 9843
rect 2468 9839 2469 9843
rect 2473 9839 2474 9843
rect 2478 9839 2479 9843
rect 2483 9839 2484 9843
rect 2488 9839 2489 9843
rect 2493 9839 2494 9843
rect 2498 9839 2499 9843
rect 2503 9839 2504 9843
rect 2508 9839 2509 9843
rect 2513 9839 2514 9843
rect 2518 9839 2519 9843
rect 2523 9839 2524 9843
rect 2528 9839 2529 9843
rect 2533 9839 2534 9843
rect 2538 9839 2539 9843
rect 2543 9839 2544 9843
rect 2548 9839 2549 9843
rect 2612 9974 2613 9978
rect 2617 9974 2618 9978
rect 2622 9974 2623 9978
rect 2627 9974 2628 9978
rect 2632 9974 2633 9978
rect 2637 9974 2638 9978
rect 2642 9974 2643 9978
rect 2647 9974 2648 9978
rect 2652 9974 2653 9978
rect 2657 9974 2658 9978
rect 2662 9974 2663 9978
rect 2667 9974 2668 9978
rect 2672 9974 2673 9978
rect 2677 9974 2678 9978
rect 2682 9974 2683 9978
rect 2687 9974 2688 9978
rect 2692 9974 2693 9978
rect 2697 9974 2698 9978
rect 2608 9973 2612 9974
rect 2608 9968 2612 9969
rect 2698 9973 2702 9974
rect 2698 9968 2702 9969
rect 2608 9963 2612 9964
rect 2608 9958 2612 9959
rect 2608 9953 2612 9954
rect 2608 9948 2612 9949
rect 2608 9943 2612 9944
rect 2608 9938 2612 9939
rect 2608 9933 2612 9934
rect 2608 9928 2612 9929
rect 2608 9923 2612 9924
rect 2608 9918 2612 9919
rect 2608 9913 2612 9914
rect 2608 9908 2612 9909
rect 2608 9903 2612 9904
rect 2608 9898 2612 9899
rect 2608 9893 2612 9894
rect 2608 9888 2612 9889
rect 2608 9883 2612 9884
rect 2608 9878 2612 9879
rect 2608 9873 2612 9874
rect 2608 9868 2612 9869
rect 2608 9863 2612 9864
rect 2608 9858 2612 9859
rect 2608 9853 2612 9854
rect 2608 9848 2612 9849
rect 2625 9961 2628 9965
rect 2632 9961 2633 9965
rect 2637 9961 2638 9965
rect 2642 9961 2643 9965
rect 2647 9961 2648 9965
rect 2652 9961 2653 9965
rect 2657 9961 2658 9965
rect 2662 9961 2663 9965
rect 2667 9961 2668 9965
rect 2672 9961 2673 9965
rect 2677 9961 2678 9965
rect 2682 9961 2685 9965
rect 2621 9958 2625 9961
rect 2621 9953 2625 9954
rect 2685 9958 2689 9961
rect 2685 9953 2689 9954
rect 2621 9948 2625 9949
rect 2621 9943 2625 9944
rect 2621 9938 2625 9939
rect 2621 9933 2625 9934
rect 2621 9928 2625 9929
rect 2621 9923 2625 9924
rect 2621 9918 2625 9919
rect 2621 9913 2625 9914
rect 2621 9908 2625 9909
rect 2621 9903 2625 9904
rect 2621 9898 2625 9899
rect 2621 9893 2625 9894
rect 2621 9888 2625 9889
rect 2621 9883 2625 9884
rect 2621 9878 2625 9879
rect 2621 9873 2625 9874
rect 2621 9868 2625 9869
rect 2637 9949 2638 9953
rect 2642 9949 2643 9953
rect 2647 9949 2648 9953
rect 2652 9949 2653 9953
rect 2657 9949 2658 9953
rect 2662 9949 2663 9953
rect 2667 9949 2668 9953
rect 2672 9949 2673 9953
rect 2633 9948 2677 9949
rect 2637 9944 2638 9948
rect 2642 9944 2643 9948
rect 2647 9944 2648 9948
rect 2652 9944 2653 9948
rect 2657 9944 2658 9948
rect 2662 9944 2663 9948
rect 2667 9944 2668 9948
rect 2672 9944 2673 9948
rect 2633 9943 2677 9944
rect 2637 9939 2638 9943
rect 2642 9939 2643 9943
rect 2647 9939 2648 9943
rect 2652 9939 2653 9943
rect 2657 9939 2658 9943
rect 2662 9939 2663 9943
rect 2667 9939 2668 9943
rect 2672 9939 2673 9943
rect 2633 9938 2677 9939
rect 2637 9934 2638 9938
rect 2642 9934 2643 9938
rect 2647 9934 2648 9938
rect 2652 9934 2653 9938
rect 2657 9934 2658 9938
rect 2662 9934 2663 9938
rect 2667 9934 2668 9938
rect 2672 9934 2673 9938
rect 2633 9933 2677 9934
rect 2637 9929 2638 9933
rect 2642 9929 2643 9933
rect 2647 9929 2648 9933
rect 2652 9929 2653 9933
rect 2657 9929 2658 9933
rect 2662 9929 2663 9933
rect 2667 9929 2668 9933
rect 2672 9929 2673 9933
rect 2633 9928 2677 9929
rect 2637 9924 2638 9928
rect 2642 9924 2643 9928
rect 2647 9924 2648 9928
rect 2652 9924 2653 9928
rect 2657 9924 2658 9928
rect 2662 9924 2663 9928
rect 2667 9924 2668 9928
rect 2672 9924 2673 9928
rect 2633 9923 2677 9924
rect 2637 9919 2638 9923
rect 2642 9919 2643 9923
rect 2647 9919 2648 9923
rect 2652 9919 2653 9923
rect 2657 9919 2658 9923
rect 2662 9919 2663 9923
rect 2667 9919 2668 9923
rect 2672 9919 2673 9923
rect 2633 9918 2677 9919
rect 2637 9914 2638 9918
rect 2642 9914 2643 9918
rect 2647 9914 2648 9918
rect 2652 9914 2653 9918
rect 2657 9914 2658 9918
rect 2662 9914 2663 9918
rect 2667 9914 2668 9918
rect 2672 9914 2673 9918
rect 2633 9913 2677 9914
rect 2637 9909 2638 9913
rect 2642 9909 2643 9913
rect 2647 9909 2648 9913
rect 2652 9909 2653 9913
rect 2657 9909 2658 9913
rect 2662 9909 2663 9913
rect 2667 9909 2668 9913
rect 2672 9909 2673 9913
rect 2633 9908 2677 9909
rect 2637 9904 2638 9908
rect 2642 9904 2643 9908
rect 2647 9904 2648 9908
rect 2652 9904 2653 9908
rect 2657 9904 2658 9908
rect 2662 9904 2663 9908
rect 2667 9904 2668 9908
rect 2672 9904 2673 9908
rect 2633 9903 2677 9904
rect 2637 9899 2638 9903
rect 2642 9899 2643 9903
rect 2647 9899 2648 9903
rect 2652 9899 2653 9903
rect 2657 9899 2658 9903
rect 2662 9899 2663 9903
rect 2667 9899 2668 9903
rect 2672 9899 2673 9903
rect 2633 9898 2677 9899
rect 2637 9894 2638 9898
rect 2642 9894 2643 9898
rect 2647 9894 2648 9898
rect 2652 9894 2653 9898
rect 2657 9894 2658 9898
rect 2662 9894 2663 9898
rect 2667 9894 2668 9898
rect 2672 9894 2673 9898
rect 2633 9893 2677 9894
rect 2637 9889 2638 9893
rect 2642 9889 2643 9893
rect 2647 9889 2648 9893
rect 2652 9889 2653 9893
rect 2657 9889 2658 9893
rect 2662 9889 2663 9893
rect 2667 9889 2668 9893
rect 2672 9889 2673 9893
rect 2633 9888 2677 9889
rect 2637 9884 2638 9888
rect 2642 9884 2643 9888
rect 2647 9884 2648 9888
rect 2652 9884 2653 9888
rect 2657 9884 2658 9888
rect 2662 9884 2663 9888
rect 2667 9884 2668 9888
rect 2672 9884 2673 9888
rect 2633 9883 2677 9884
rect 2637 9879 2638 9883
rect 2642 9879 2643 9883
rect 2647 9879 2648 9883
rect 2652 9879 2653 9883
rect 2657 9879 2658 9883
rect 2662 9879 2663 9883
rect 2667 9879 2668 9883
rect 2672 9879 2673 9883
rect 2633 9878 2677 9879
rect 2637 9874 2638 9878
rect 2642 9874 2643 9878
rect 2647 9874 2648 9878
rect 2652 9874 2653 9878
rect 2657 9874 2658 9878
rect 2662 9874 2663 9878
rect 2667 9874 2668 9878
rect 2672 9874 2673 9878
rect 2633 9873 2677 9874
rect 2637 9869 2638 9873
rect 2642 9869 2643 9873
rect 2647 9869 2648 9873
rect 2652 9869 2653 9873
rect 2657 9869 2658 9873
rect 2662 9869 2663 9873
rect 2667 9869 2668 9873
rect 2672 9869 2673 9873
rect 2633 9868 2677 9869
rect 2637 9864 2638 9868
rect 2642 9864 2643 9868
rect 2647 9864 2648 9868
rect 2652 9864 2653 9868
rect 2657 9864 2658 9868
rect 2662 9864 2663 9868
rect 2667 9864 2668 9868
rect 2672 9864 2673 9868
rect 2685 9948 2689 9949
rect 2685 9943 2689 9944
rect 2685 9938 2689 9939
rect 2685 9933 2689 9934
rect 2685 9928 2689 9929
rect 2685 9923 2689 9924
rect 2685 9918 2689 9919
rect 2685 9913 2689 9914
rect 2685 9908 2689 9909
rect 2685 9903 2689 9904
rect 2685 9898 2689 9899
rect 2685 9893 2689 9894
rect 2685 9888 2689 9889
rect 2685 9883 2689 9884
rect 2685 9878 2689 9879
rect 2685 9873 2689 9874
rect 2685 9868 2689 9869
rect 2621 9863 2625 9864
rect 2621 9856 2625 9859
rect 2685 9863 2689 9864
rect 2685 9856 2689 9859
rect 2625 9848 2628 9856
rect 2632 9848 2633 9856
rect 2637 9848 2638 9856
rect 2642 9848 2643 9856
rect 2647 9848 2648 9856
rect 2652 9848 2653 9856
rect 2657 9848 2658 9856
rect 2662 9848 2663 9856
rect 2667 9848 2668 9856
rect 2672 9848 2673 9856
rect 2677 9848 2678 9856
rect 2682 9848 2685 9856
rect 2698 9963 2702 9964
rect 2698 9958 2702 9959
rect 2698 9953 2702 9954
rect 2724 9961 2745 9981
rect 2772 9974 2773 9978
rect 2777 9974 2778 9978
rect 2782 9974 2783 9978
rect 2787 9974 2788 9978
rect 2792 9974 2793 9978
rect 2797 9974 2798 9978
rect 2802 9974 2803 9978
rect 2807 9974 2808 9978
rect 2812 9974 2813 9978
rect 2817 9974 2818 9978
rect 2822 9974 2823 9978
rect 2827 9974 2828 9978
rect 2832 9974 2833 9978
rect 2837 9974 2838 9978
rect 2842 9974 2843 9978
rect 2847 9974 2848 9978
rect 2852 9974 2853 9978
rect 2857 9974 2858 9978
rect 2768 9973 2772 9974
rect 2768 9968 2772 9969
rect 2858 9973 2862 9974
rect 2858 9968 2862 9969
rect 2768 9963 2772 9964
rect 2768 9958 2772 9959
rect 2768 9953 2772 9954
rect 2698 9948 2702 9949
rect 2698 9943 2702 9944
rect 2698 9938 2702 9939
rect 2698 9933 2702 9934
rect 2698 9928 2702 9929
rect 2698 9923 2702 9924
rect 2698 9918 2702 9919
rect 2698 9913 2702 9914
rect 2698 9908 2702 9909
rect 2698 9903 2702 9904
rect 2698 9898 2702 9899
rect 2698 9893 2702 9894
rect 2698 9888 2702 9889
rect 2698 9883 2702 9884
rect 2768 9948 2772 9949
rect 2768 9943 2772 9944
rect 2768 9938 2772 9939
rect 2768 9933 2772 9934
rect 2768 9928 2772 9929
rect 2768 9923 2772 9924
rect 2768 9918 2772 9919
rect 2768 9913 2772 9914
rect 2768 9908 2772 9909
rect 2768 9903 2772 9904
rect 2768 9898 2772 9899
rect 2768 9893 2772 9894
rect 2768 9888 2772 9889
rect 2768 9883 2772 9884
rect 2698 9878 2702 9879
rect 2698 9873 2702 9874
rect 2698 9868 2702 9869
rect 2698 9863 2702 9864
rect 2698 9858 2702 9859
rect 2698 9853 2702 9854
rect 2698 9848 2702 9849
rect 2608 9843 2612 9844
rect 2724 9846 2745 9874
rect 2768 9878 2772 9879
rect 2768 9873 2772 9874
rect 2768 9868 2772 9869
rect 2768 9863 2772 9864
rect 2768 9858 2772 9859
rect 2768 9853 2772 9854
rect 2768 9848 2772 9849
rect 2785 9961 2788 9965
rect 2792 9961 2793 9965
rect 2797 9961 2798 9965
rect 2802 9961 2803 9965
rect 2807 9961 2808 9965
rect 2812 9961 2813 9965
rect 2817 9961 2818 9965
rect 2822 9961 2823 9965
rect 2827 9961 2828 9965
rect 2832 9961 2833 9965
rect 2837 9961 2838 9965
rect 2842 9961 2845 9965
rect 2781 9958 2785 9961
rect 2781 9953 2785 9954
rect 2845 9958 2849 9961
rect 2845 9953 2849 9954
rect 2781 9948 2785 9949
rect 2781 9943 2785 9944
rect 2781 9938 2785 9939
rect 2781 9933 2785 9934
rect 2781 9928 2785 9929
rect 2781 9923 2785 9924
rect 2781 9918 2785 9919
rect 2781 9913 2785 9914
rect 2781 9908 2785 9909
rect 2781 9903 2785 9904
rect 2781 9898 2785 9899
rect 2781 9893 2785 9894
rect 2781 9888 2785 9889
rect 2781 9883 2785 9884
rect 2781 9878 2785 9879
rect 2781 9873 2785 9874
rect 2781 9868 2785 9869
rect 2792 9949 2793 9953
rect 2797 9949 2798 9953
rect 2802 9949 2803 9953
rect 2807 9949 2808 9953
rect 2812 9949 2813 9953
rect 2817 9949 2818 9953
rect 2822 9949 2823 9953
rect 2827 9949 2828 9953
rect 2832 9949 2833 9953
rect 2792 9948 2837 9949
rect 2792 9944 2793 9948
rect 2797 9944 2798 9948
rect 2802 9944 2803 9948
rect 2807 9944 2808 9948
rect 2812 9944 2813 9948
rect 2817 9944 2818 9948
rect 2822 9944 2823 9948
rect 2827 9944 2828 9948
rect 2832 9944 2833 9948
rect 2792 9943 2837 9944
rect 2792 9939 2793 9943
rect 2797 9939 2798 9943
rect 2802 9939 2803 9943
rect 2807 9939 2808 9943
rect 2812 9939 2813 9943
rect 2817 9939 2818 9943
rect 2822 9939 2823 9943
rect 2827 9939 2828 9943
rect 2832 9939 2833 9943
rect 2792 9938 2837 9939
rect 2792 9934 2793 9938
rect 2797 9934 2798 9938
rect 2802 9934 2803 9938
rect 2807 9934 2808 9938
rect 2812 9934 2813 9938
rect 2817 9934 2818 9938
rect 2822 9934 2823 9938
rect 2827 9934 2828 9938
rect 2832 9934 2833 9938
rect 2792 9933 2837 9934
rect 2792 9929 2793 9933
rect 2797 9929 2798 9933
rect 2802 9929 2803 9933
rect 2807 9929 2808 9933
rect 2812 9929 2813 9933
rect 2817 9929 2818 9933
rect 2822 9929 2823 9933
rect 2827 9929 2828 9933
rect 2832 9929 2833 9933
rect 2792 9928 2837 9929
rect 2792 9924 2793 9928
rect 2797 9924 2798 9928
rect 2802 9924 2803 9928
rect 2807 9924 2808 9928
rect 2812 9924 2813 9928
rect 2817 9924 2818 9928
rect 2822 9924 2823 9928
rect 2827 9924 2828 9928
rect 2832 9924 2833 9928
rect 2792 9923 2837 9924
rect 2792 9919 2793 9923
rect 2797 9919 2798 9923
rect 2802 9919 2803 9923
rect 2807 9919 2808 9923
rect 2812 9919 2813 9923
rect 2817 9919 2818 9923
rect 2822 9919 2823 9923
rect 2827 9919 2828 9923
rect 2832 9919 2833 9923
rect 2792 9918 2837 9919
rect 2792 9914 2793 9918
rect 2797 9914 2798 9918
rect 2802 9914 2803 9918
rect 2807 9914 2808 9918
rect 2812 9914 2813 9918
rect 2817 9914 2818 9918
rect 2822 9914 2823 9918
rect 2827 9914 2828 9918
rect 2832 9914 2833 9918
rect 2792 9913 2837 9914
rect 2792 9909 2793 9913
rect 2797 9909 2798 9913
rect 2802 9909 2803 9913
rect 2807 9909 2808 9913
rect 2812 9909 2813 9913
rect 2817 9909 2818 9913
rect 2822 9909 2823 9913
rect 2827 9909 2828 9913
rect 2832 9909 2833 9913
rect 2792 9908 2837 9909
rect 2792 9904 2793 9908
rect 2797 9904 2798 9908
rect 2802 9904 2803 9908
rect 2807 9904 2808 9908
rect 2812 9904 2813 9908
rect 2817 9904 2818 9908
rect 2822 9904 2823 9908
rect 2827 9904 2828 9908
rect 2832 9904 2833 9908
rect 2792 9903 2837 9904
rect 2792 9899 2793 9903
rect 2797 9899 2798 9903
rect 2802 9899 2803 9903
rect 2807 9899 2808 9903
rect 2812 9899 2813 9903
rect 2817 9899 2818 9903
rect 2822 9899 2823 9903
rect 2827 9899 2828 9903
rect 2832 9899 2833 9903
rect 2792 9898 2837 9899
rect 2792 9894 2793 9898
rect 2797 9894 2798 9898
rect 2802 9894 2803 9898
rect 2807 9894 2808 9898
rect 2812 9894 2813 9898
rect 2817 9894 2818 9898
rect 2822 9894 2823 9898
rect 2827 9894 2828 9898
rect 2832 9894 2833 9898
rect 2792 9893 2837 9894
rect 2792 9889 2793 9893
rect 2797 9889 2798 9893
rect 2802 9889 2803 9893
rect 2807 9889 2808 9893
rect 2812 9889 2813 9893
rect 2817 9889 2818 9893
rect 2822 9889 2823 9893
rect 2827 9889 2828 9893
rect 2832 9889 2833 9893
rect 2792 9888 2837 9889
rect 2792 9884 2793 9888
rect 2797 9884 2798 9888
rect 2802 9884 2803 9888
rect 2807 9884 2808 9888
rect 2812 9884 2813 9888
rect 2817 9884 2818 9888
rect 2822 9884 2823 9888
rect 2827 9884 2828 9888
rect 2832 9884 2833 9888
rect 2792 9883 2837 9884
rect 2792 9879 2793 9883
rect 2797 9879 2798 9883
rect 2802 9879 2803 9883
rect 2807 9879 2808 9883
rect 2812 9879 2813 9883
rect 2817 9879 2818 9883
rect 2822 9879 2823 9883
rect 2827 9879 2828 9883
rect 2832 9879 2833 9883
rect 2792 9878 2837 9879
rect 2792 9874 2793 9878
rect 2797 9874 2798 9878
rect 2802 9874 2803 9878
rect 2807 9874 2808 9878
rect 2812 9874 2813 9878
rect 2817 9874 2818 9878
rect 2822 9874 2823 9878
rect 2827 9874 2828 9878
rect 2832 9874 2833 9878
rect 2792 9873 2837 9874
rect 2792 9869 2793 9873
rect 2797 9869 2798 9873
rect 2802 9869 2803 9873
rect 2807 9869 2808 9873
rect 2812 9869 2813 9873
rect 2817 9869 2818 9873
rect 2822 9869 2823 9873
rect 2827 9869 2828 9873
rect 2832 9869 2833 9873
rect 2792 9868 2837 9869
rect 2792 9864 2793 9868
rect 2797 9864 2798 9868
rect 2802 9864 2803 9868
rect 2807 9864 2808 9868
rect 2812 9864 2813 9868
rect 2817 9864 2818 9868
rect 2822 9864 2823 9868
rect 2827 9864 2828 9868
rect 2832 9864 2833 9868
rect 2845 9948 2849 9949
rect 2845 9943 2849 9944
rect 2845 9938 2849 9939
rect 2845 9933 2849 9934
rect 2845 9928 2849 9929
rect 2845 9923 2849 9924
rect 2845 9918 2849 9919
rect 2845 9913 2849 9914
rect 2845 9908 2849 9909
rect 2845 9903 2849 9904
rect 2845 9898 2849 9899
rect 2845 9893 2849 9894
rect 2845 9888 2849 9889
rect 2845 9883 2849 9884
rect 2845 9878 2849 9879
rect 2845 9873 2849 9874
rect 2845 9868 2849 9869
rect 2781 9863 2785 9864
rect 2781 9856 2785 9859
rect 2845 9863 2849 9864
rect 2845 9856 2849 9859
rect 2785 9848 2788 9856
rect 2792 9848 2793 9856
rect 2797 9848 2798 9856
rect 2802 9848 2803 9856
rect 2807 9848 2808 9856
rect 2812 9848 2813 9856
rect 2817 9848 2818 9856
rect 2822 9848 2823 9856
rect 2827 9848 2828 9856
rect 2832 9848 2833 9856
rect 2837 9848 2838 9856
rect 2842 9848 2845 9856
rect 2858 9963 2862 9964
rect 2858 9958 2862 9959
rect 2858 9953 2862 9954
rect 2858 9948 2862 9949
rect 2858 9943 2862 9944
rect 2858 9938 2862 9939
rect 2858 9933 2862 9934
rect 2858 9928 2862 9929
rect 2858 9923 2862 9924
rect 2858 9918 2862 9919
rect 2858 9913 2862 9914
rect 2858 9908 2862 9909
rect 2858 9903 2862 9904
rect 2858 9898 2862 9899
rect 2858 9893 2862 9894
rect 2858 9888 2862 9889
rect 2858 9883 2862 9884
rect 2858 9878 2862 9879
rect 2858 9873 2862 9874
rect 2858 9868 2862 9869
rect 2858 9863 2862 9864
rect 2858 9858 2862 9859
rect 2858 9853 2862 9854
rect 2858 9848 2862 9849
rect 2726 9844 2743 9846
rect 2698 9843 2702 9844
rect 2612 9839 2613 9843
rect 2617 9839 2618 9843
rect 2622 9839 2623 9843
rect 2627 9839 2628 9843
rect 2632 9839 2633 9843
rect 2637 9839 2638 9843
rect 2642 9839 2643 9843
rect 2647 9839 2648 9843
rect 2652 9839 2653 9843
rect 2657 9839 2658 9843
rect 2662 9839 2663 9843
rect 2667 9839 2668 9843
rect 2672 9839 2673 9843
rect 2677 9839 2678 9843
rect 2682 9839 2683 9843
rect 2687 9839 2688 9843
rect 2692 9839 2693 9843
rect 2697 9839 2698 9843
rect 2728 9842 2741 9844
rect 2768 9843 2772 9844
rect 2858 9843 2862 9844
rect 2496 9831 2552 9839
rect 2302 9827 2361 9831
rect 2487 9827 2552 9831
rect 2302 9815 2358 9827
rect 2417 9819 2447 9823
rect 2302 9811 2361 9815
rect 2431 9812 2435 9819
rect 2496 9815 2552 9827
rect 2302 9802 2358 9811
rect 2487 9811 2552 9815
rect 2417 9803 2428 9807
rect 2178 9795 2243 9799
rect 1981 9790 2049 9791
rect 1981 9786 1982 9790
rect 1986 9786 1987 9790
rect 1991 9786 2049 9790
rect 2108 9787 2138 9791
rect 1981 9785 2049 9786
rect 1981 9781 1982 9785
rect 1986 9781 1987 9785
rect 1991 9783 2049 9785
rect 1991 9781 2052 9783
rect 1981 9780 2052 9781
rect 1981 9776 1982 9780
rect 1986 9776 1987 9780
rect 1991 9779 2052 9780
rect 1991 9776 2049 9779
rect 1981 9775 2049 9776
rect 1981 9771 1982 9775
rect 1986 9771 1987 9775
rect 1991 9771 2049 9775
rect 1981 9770 2049 9771
rect 1981 9766 1982 9770
rect 1986 9766 1987 9770
rect 1991 9766 2049 9770
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1937 9761 1956 9762
rect 1941 9757 1942 9761
rect 1946 9757 1947 9761
rect 1951 9757 1952 9761
rect 1937 9756 1956 9757
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1937 9751 1956 9752
rect 1941 9747 1942 9751
rect 1946 9747 1947 9751
rect 1951 9747 1952 9751
rect 1937 9746 1956 9747
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1937 9741 1956 9742
rect 1941 9737 1942 9741
rect 1946 9737 1947 9741
rect 1951 9737 1952 9741
rect 1937 9736 1956 9737
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1981 9765 2049 9766
rect 1981 9761 1982 9765
rect 1986 9761 1987 9765
rect 1991 9761 2049 9765
rect 1981 9760 2049 9761
rect 1981 9756 1982 9760
rect 1986 9756 1987 9760
rect 1991 9756 2049 9760
rect 1981 9755 2049 9756
rect 1981 9751 1982 9755
rect 1986 9751 1987 9755
rect 1991 9751 2049 9755
rect 1981 9750 2049 9751
rect 1981 9746 1982 9750
rect 1986 9746 1987 9750
rect 1991 9746 2049 9750
rect 1981 9745 2049 9746
rect 1981 9741 1982 9745
rect 1986 9741 1987 9745
rect 1991 9741 2049 9745
rect 1981 9740 2049 9741
rect 1981 9736 1982 9740
rect 1986 9736 1987 9740
rect 1991 9736 2049 9740
rect 1981 9734 2049 9736
rect 1882 9718 1883 9722
rect 1887 9718 1888 9722
rect 1892 9718 1893 9722
rect 1897 9718 1898 9722
rect 1902 9718 1903 9722
rect 1907 9718 1908 9722
rect 1912 9718 1913 9722
rect 1917 9718 1918 9722
rect 1922 9718 1923 9722
rect 1927 9718 1928 9722
rect 1932 9718 1934 9722
rect 1878 9717 1934 9718
rect 1882 9713 1883 9717
rect 1887 9713 1888 9717
rect 1892 9713 1893 9717
rect 1897 9713 1898 9717
rect 1902 9713 1903 9717
rect 1907 9713 1908 9717
rect 1912 9713 1913 9717
rect 1917 9713 1918 9717
rect 1922 9713 1923 9717
rect 1927 9713 1928 9717
rect 1932 9713 1934 9717
rect 1878 9712 1934 9713
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1937 9715 1956 9716
rect 1941 9711 1942 9715
rect 1946 9711 1947 9715
rect 1951 9711 1952 9715
rect 1937 9710 1956 9711
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1937 9705 1956 9706
rect 1941 9701 1942 9705
rect 1946 9701 1947 9705
rect 1951 9701 1952 9705
rect 1937 9700 1956 9701
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1937 9695 1956 9696
rect 1941 9691 1942 9695
rect 1946 9691 1947 9695
rect 1951 9691 1952 9695
rect 1937 9690 1956 9691
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 2113 9597 2126 9787
rect 2187 9783 2243 9795
rect 2178 9779 2243 9783
rect 2187 9722 2243 9779
rect 2290 9800 2358 9802
rect 2290 9796 2291 9800
rect 2295 9796 2296 9800
rect 2300 9799 2358 9800
rect 2421 9800 2428 9803
rect 2440 9803 2447 9807
rect 2440 9800 2444 9803
rect 2300 9796 2361 9799
rect 2290 9795 2361 9796
rect 2290 9791 2291 9795
rect 2295 9791 2296 9795
rect 2300 9791 2358 9795
rect 2421 9791 2444 9800
rect 2496 9799 2552 9811
rect 2611 9831 2667 9839
rect 2730 9831 2739 9842
rect 2772 9839 2773 9843
rect 2777 9839 2778 9843
rect 2782 9839 2783 9843
rect 2787 9839 2788 9843
rect 2792 9839 2793 9843
rect 2797 9839 2798 9843
rect 2802 9839 2803 9843
rect 2807 9839 2808 9843
rect 2812 9839 2813 9843
rect 2817 9839 2818 9843
rect 2822 9839 2823 9843
rect 2827 9839 2828 9843
rect 2832 9839 2833 9843
rect 2837 9839 2838 9843
rect 2842 9839 2843 9843
rect 2847 9839 2848 9843
rect 2852 9839 2853 9843
rect 2857 9839 2858 9843
rect 2921 9974 2922 9978
rect 2926 9974 2927 9978
rect 2931 9974 2932 9978
rect 2936 9974 2937 9978
rect 2941 9974 2942 9978
rect 2946 9974 2947 9978
rect 2951 9974 2952 9978
rect 2956 9974 2957 9978
rect 2961 9974 2962 9978
rect 2966 9974 2967 9978
rect 2971 9974 2972 9978
rect 2976 9974 2977 9978
rect 2981 9974 2982 9978
rect 2986 9974 2987 9978
rect 2991 9974 2992 9978
rect 2996 9974 2997 9978
rect 3001 9974 3002 9978
rect 3006 9974 3007 9978
rect 2917 9973 2921 9974
rect 2917 9968 2921 9969
rect 3007 9973 3011 9974
rect 3007 9968 3011 9969
rect 2917 9963 2921 9964
rect 2917 9958 2921 9959
rect 2917 9953 2921 9954
rect 2917 9948 2921 9949
rect 2917 9943 2921 9944
rect 2917 9938 2921 9939
rect 2917 9933 2921 9934
rect 2917 9928 2921 9929
rect 2917 9923 2921 9924
rect 2917 9918 2921 9919
rect 2917 9913 2921 9914
rect 2917 9908 2921 9909
rect 2917 9903 2921 9904
rect 2917 9898 2921 9899
rect 2917 9893 2921 9894
rect 2917 9888 2921 9889
rect 2917 9883 2921 9884
rect 2917 9878 2921 9879
rect 2917 9873 2921 9874
rect 2917 9868 2921 9869
rect 2917 9863 2921 9864
rect 2917 9858 2921 9859
rect 2917 9853 2921 9854
rect 2917 9848 2921 9849
rect 2934 9961 2937 9965
rect 2941 9961 2942 9965
rect 2946 9961 2947 9965
rect 2951 9961 2952 9965
rect 2956 9961 2957 9965
rect 2961 9961 2962 9965
rect 2966 9961 2967 9965
rect 2971 9961 2972 9965
rect 2976 9961 2977 9965
rect 2981 9961 2982 9965
rect 2986 9961 2987 9965
rect 2991 9961 2994 9965
rect 2930 9958 2934 9961
rect 2930 9953 2934 9954
rect 2994 9958 2998 9961
rect 2994 9953 2998 9954
rect 2930 9948 2934 9949
rect 2930 9943 2934 9944
rect 2930 9938 2934 9939
rect 2930 9933 2934 9934
rect 2930 9928 2934 9929
rect 2930 9923 2934 9924
rect 2930 9918 2934 9919
rect 2930 9913 2934 9914
rect 2930 9908 2934 9909
rect 2930 9903 2934 9904
rect 2930 9898 2934 9899
rect 2930 9893 2934 9894
rect 2930 9888 2934 9889
rect 2930 9883 2934 9884
rect 2930 9878 2934 9879
rect 2930 9873 2934 9874
rect 2930 9868 2934 9869
rect 2946 9949 2947 9953
rect 2951 9949 2952 9953
rect 2956 9949 2957 9953
rect 2961 9949 2962 9953
rect 2966 9949 2967 9953
rect 2971 9949 2972 9953
rect 2976 9949 2977 9953
rect 2981 9949 2982 9953
rect 2942 9948 2986 9949
rect 2946 9944 2947 9948
rect 2951 9944 2952 9948
rect 2956 9944 2957 9948
rect 2961 9944 2962 9948
rect 2966 9944 2967 9948
rect 2971 9944 2972 9948
rect 2976 9944 2977 9948
rect 2981 9944 2982 9948
rect 2942 9943 2986 9944
rect 2946 9939 2947 9943
rect 2951 9939 2952 9943
rect 2956 9939 2957 9943
rect 2961 9939 2962 9943
rect 2966 9939 2967 9943
rect 2971 9939 2972 9943
rect 2976 9939 2977 9943
rect 2981 9939 2982 9943
rect 2942 9938 2986 9939
rect 2946 9934 2947 9938
rect 2951 9934 2952 9938
rect 2956 9934 2957 9938
rect 2961 9934 2962 9938
rect 2966 9934 2967 9938
rect 2971 9934 2972 9938
rect 2976 9934 2977 9938
rect 2981 9934 2982 9938
rect 2942 9933 2986 9934
rect 2946 9929 2947 9933
rect 2951 9929 2952 9933
rect 2956 9929 2957 9933
rect 2961 9929 2962 9933
rect 2966 9929 2967 9933
rect 2971 9929 2972 9933
rect 2976 9929 2977 9933
rect 2981 9929 2982 9933
rect 2942 9928 2986 9929
rect 2946 9924 2947 9928
rect 2951 9924 2952 9928
rect 2956 9924 2957 9928
rect 2961 9924 2962 9928
rect 2966 9924 2967 9928
rect 2971 9924 2972 9928
rect 2976 9924 2977 9928
rect 2981 9924 2982 9928
rect 2942 9923 2986 9924
rect 2946 9919 2947 9923
rect 2951 9919 2952 9923
rect 2956 9919 2957 9923
rect 2961 9919 2962 9923
rect 2966 9919 2967 9923
rect 2971 9919 2972 9923
rect 2976 9919 2977 9923
rect 2981 9919 2982 9923
rect 2942 9918 2986 9919
rect 2946 9914 2947 9918
rect 2951 9914 2952 9918
rect 2956 9914 2957 9918
rect 2961 9914 2962 9918
rect 2966 9914 2967 9918
rect 2971 9914 2972 9918
rect 2976 9914 2977 9918
rect 2981 9914 2982 9918
rect 2942 9913 2986 9914
rect 2946 9909 2947 9913
rect 2951 9909 2952 9913
rect 2956 9909 2957 9913
rect 2961 9909 2962 9913
rect 2966 9909 2967 9913
rect 2971 9909 2972 9913
rect 2976 9909 2977 9913
rect 2981 9909 2982 9913
rect 2942 9908 2986 9909
rect 2946 9904 2947 9908
rect 2951 9904 2952 9908
rect 2956 9904 2957 9908
rect 2961 9904 2962 9908
rect 2966 9904 2967 9908
rect 2971 9904 2972 9908
rect 2976 9904 2977 9908
rect 2981 9904 2982 9908
rect 2942 9903 2986 9904
rect 2946 9899 2947 9903
rect 2951 9899 2952 9903
rect 2956 9899 2957 9903
rect 2961 9899 2962 9903
rect 2966 9899 2967 9903
rect 2971 9899 2972 9903
rect 2976 9899 2977 9903
rect 2981 9899 2982 9903
rect 2942 9898 2986 9899
rect 2946 9894 2947 9898
rect 2951 9894 2952 9898
rect 2956 9894 2957 9898
rect 2961 9894 2962 9898
rect 2966 9894 2967 9898
rect 2971 9894 2972 9898
rect 2976 9894 2977 9898
rect 2981 9894 2982 9898
rect 2942 9893 2986 9894
rect 2946 9889 2947 9893
rect 2951 9889 2952 9893
rect 2956 9889 2957 9893
rect 2961 9889 2962 9893
rect 2966 9889 2967 9893
rect 2971 9889 2972 9893
rect 2976 9889 2977 9893
rect 2981 9889 2982 9893
rect 2942 9888 2986 9889
rect 2946 9884 2947 9888
rect 2951 9884 2952 9888
rect 2956 9884 2957 9888
rect 2961 9884 2962 9888
rect 2966 9884 2967 9888
rect 2971 9884 2972 9888
rect 2976 9884 2977 9888
rect 2981 9884 2982 9888
rect 2942 9883 2986 9884
rect 2946 9879 2947 9883
rect 2951 9879 2952 9883
rect 2956 9879 2957 9883
rect 2961 9879 2962 9883
rect 2966 9879 2967 9883
rect 2971 9879 2972 9883
rect 2976 9879 2977 9883
rect 2981 9879 2982 9883
rect 2942 9878 2986 9879
rect 2946 9874 2947 9878
rect 2951 9874 2952 9878
rect 2956 9874 2957 9878
rect 2961 9874 2962 9878
rect 2966 9874 2967 9878
rect 2971 9874 2972 9878
rect 2976 9874 2977 9878
rect 2981 9874 2982 9878
rect 2942 9873 2986 9874
rect 2946 9869 2947 9873
rect 2951 9869 2952 9873
rect 2956 9869 2957 9873
rect 2961 9869 2962 9873
rect 2966 9869 2967 9873
rect 2971 9869 2972 9873
rect 2976 9869 2977 9873
rect 2981 9869 2982 9873
rect 2942 9868 2986 9869
rect 2946 9864 2947 9868
rect 2951 9864 2952 9868
rect 2956 9864 2957 9868
rect 2961 9864 2962 9868
rect 2966 9864 2967 9868
rect 2971 9864 2972 9868
rect 2976 9864 2977 9868
rect 2981 9864 2982 9868
rect 2994 9948 2998 9949
rect 2994 9943 2998 9944
rect 2994 9938 2998 9939
rect 2994 9933 2998 9934
rect 2994 9928 2998 9929
rect 2994 9923 2998 9924
rect 2994 9918 2998 9919
rect 2994 9913 2998 9914
rect 2994 9908 2998 9909
rect 2994 9903 2998 9904
rect 2994 9898 2998 9899
rect 2994 9893 2998 9894
rect 2994 9888 2998 9889
rect 2994 9883 2998 9884
rect 2994 9878 2998 9879
rect 2994 9873 2998 9874
rect 2994 9868 2998 9869
rect 2930 9863 2934 9864
rect 2930 9856 2934 9859
rect 2994 9863 2998 9864
rect 2994 9856 2998 9859
rect 2934 9848 2937 9856
rect 2941 9848 2942 9856
rect 2946 9848 2947 9856
rect 2951 9848 2952 9856
rect 2956 9848 2957 9856
rect 2961 9848 2962 9856
rect 2966 9848 2967 9856
rect 2971 9848 2972 9856
rect 2976 9848 2977 9856
rect 2981 9848 2982 9856
rect 2986 9848 2987 9856
rect 2991 9848 2994 9856
rect 3007 9963 3011 9964
rect 3007 9958 3011 9959
rect 3007 9953 3011 9954
rect 3033 9961 3054 9981
rect 3081 9974 3082 9978
rect 3086 9974 3087 9978
rect 3091 9974 3092 9978
rect 3096 9974 3097 9978
rect 3101 9974 3102 9978
rect 3106 9974 3107 9978
rect 3111 9974 3112 9978
rect 3116 9974 3117 9978
rect 3121 9974 3122 9978
rect 3126 9974 3127 9978
rect 3131 9974 3132 9978
rect 3136 9974 3137 9978
rect 3141 9974 3142 9978
rect 3146 9974 3147 9978
rect 3151 9974 3152 9978
rect 3156 9974 3157 9978
rect 3161 9974 3162 9978
rect 3166 9974 3167 9978
rect 3077 9973 3081 9974
rect 3077 9968 3081 9969
rect 3167 9973 3171 9974
rect 3167 9968 3171 9969
rect 3077 9963 3081 9964
rect 3077 9958 3081 9959
rect 3077 9953 3081 9954
rect 3007 9948 3011 9949
rect 3007 9943 3011 9944
rect 3007 9938 3011 9939
rect 3007 9933 3011 9934
rect 3007 9928 3011 9929
rect 3007 9923 3011 9924
rect 3007 9918 3011 9919
rect 3007 9913 3011 9914
rect 3007 9908 3011 9909
rect 3007 9903 3011 9904
rect 3007 9898 3011 9899
rect 3007 9893 3011 9894
rect 3007 9888 3011 9889
rect 3007 9883 3011 9884
rect 3077 9948 3081 9949
rect 3077 9943 3081 9944
rect 3077 9938 3081 9939
rect 3077 9933 3081 9934
rect 3077 9928 3081 9929
rect 3077 9923 3081 9924
rect 3077 9918 3081 9919
rect 3077 9913 3081 9914
rect 3077 9908 3081 9909
rect 3077 9903 3081 9904
rect 3077 9898 3081 9899
rect 3077 9893 3081 9894
rect 3077 9888 3081 9889
rect 3077 9883 3081 9884
rect 3007 9878 3011 9879
rect 3007 9873 3011 9874
rect 3007 9868 3011 9869
rect 3007 9863 3011 9864
rect 3007 9858 3011 9859
rect 3007 9853 3011 9854
rect 3007 9848 3011 9849
rect 2917 9843 2921 9844
rect 3033 9846 3054 9874
rect 3077 9878 3081 9879
rect 3077 9873 3081 9874
rect 3077 9868 3081 9869
rect 3077 9863 3081 9864
rect 3077 9858 3081 9859
rect 3077 9853 3081 9854
rect 3077 9848 3081 9849
rect 3094 9961 3097 9965
rect 3101 9961 3102 9965
rect 3106 9961 3107 9965
rect 3111 9961 3112 9965
rect 3116 9961 3117 9965
rect 3121 9961 3122 9965
rect 3126 9961 3127 9965
rect 3131 9961 3132 9965
rect 3136 9961 3137 9965
rect 3141 9961 3142 9965
rect 3146 9961 3147 9965
rect 3151 9961 3154 9965
rect 3090 9958 3094 9961
rect 3090 9953 3094 9954
rect 3154 9958 3158 9961
rect 3154 9953 3158 9954
rect 3090 9948 3094 9949
rect 3090 9943 3094 9944
rect 3090 9938 3094 9939
rect 3090 9933 3094 9934
rect 3090 9928 3094 9929
rect 3090 9923 3094 9924
rect 3090 9918 3094 9919
rect 3090 9913 3094 9914
rect 3090 9908 3094 9909
rect 3090 9903 3094 9904
rect 3090 9898 3094 9899
rect 3090 9893 3094 9894
rect 3090 9888 3094 9889
rect 3090 9883 3094 9884
rect 3090 9878 3094 9879
rect 3090 9873 3094 9874
rect 3090 9868 3094 9869
rect 3101 9949 3102 9953
rect 3106 9949 3107 9953
rect 3111 9949 3112 9953
rect 3116 9949 3117 9953
rect 3121 9949 3122 9953
rect 3126 9949 3127 9953
rect 3131 9949 3132 9953
rect 3136 9949 3137 9953
rect 3141 9949 3142 9953
rect 3101 9948 3146 9949
rect 3101 9944 3102 9948
rect 3106 9944 3107 9948
rect 3111 9944 3112 9948
rect 3116 9944 3117 9948
rect 3121 9944 3122 9948
rect 3126 9944 3127 9948
rect 3131 9944 3132 9948
rect 3136 9944 3137 9948
rect 3141 9944 3142 9948
rect 3101 9943 3146 9944
rect 3101 9939 3102 9943
rect 3106 9939 3107 9943
rect 3111 9939 3112 9943
rect 3116 9939 3117 9943
rect 3121 9939 3122 9943
rect 3126 9939 3127 9943
rect 3131 9939 3132 9943
rect 3136 9939 3137 9943
rect 3141 9939 3142 9943
rect 3101 9938 3146 9939
rect 3101 9934 3102 9938
rect 3106 9934 3107 9938
rect 3111 9934 3112 9938
rect 3116 9934 3117 9938
rect 3121 9934 3122 9938
rect 3126 9934 3127 9938
rect 3131 9934 3132 9938
rect 3136 9934 3137 9938
rect 3141 9934 3142 9938
rect 3101 9933 3146 9934
rect 3101 9929 3102 9933
rect 3106 9929 3107 9933
rect 3111 9929 3112 9933
rect 3116 9929 3117 9933
rect 3121 9929 3122 9933
rect 3126 9929 3127 9933
rect 3131 9929 3132 9933
rect 3136 9929 3137 9933
rect 3141 9929 3142 9933
rect 3101 9928 3146 9929
rect 3101 9924 3102 9928
rect 3106 9924 3107 9928
rect 3111 9924 3112 9928
rect 3116 9924 3117 9928
rect 3121 9924 3122 9928
rect 3126 9924 3127 9928
rect 3131 9924 3132 9928
rect 3136 9924 3137 9928
rect 3141 9924 3142 9928
rect 3101 9923 3146 9924
rect 3101 9919 3102 9923
rect 3106 9919 3107 9923
rect 3111 9919 3112 9923
rect 3116 9919 3117 9923
rect 3121 9919 3122 9923
rect 3126 9919 3127 9923
rect 3131 9919 3132 9923
rect 3136 9919 3137 9923
rect 3141 9919 3142 9923
rect 3101 9918 3146 9919
rect 3101 9914 3102 9918
rect 3106 9914 3107 9918
rect 3111 9914 3112 9918
rect 3116 9914 3117 9918
rect 3121 9914 3122 9918
rect 3126 9914 3127 9918
rect 3131 9914 3132 9918
rect 3136 9914 3137 9918
rect 3141 9914 3142 9918
rect 3101 9913 3146 9914
rect 3101 9909 3102 9913
rect 3106 9909 3107 9913
rect 3111 9909 3112 9913
rect 3116 9909 3117 9913
rect 3121 9909 3122 9913
rect 3126 9909 3127 9913
rect 3131 9909 3132 9913
rect 3136 9909 3137 9913
rect 3141 9909 3142 9913
rect 3101 9908 3146 9909
rect 3101 9904 3102 9908
rect 3106 9904 3107 9908
rect 3111 9904 3112 9908
rect 3116 9904 3117 9908
rect 3121 9904 3122 9908
rect 3126 9904 3127 9908
rect 3131 9904 3132 9908
rect 3136 9904 3137 9908
rect 3141 9904 3142 9908
rect 3101 9903 3146 9904
rect 3101 9899 3102 9903
rect 3106 9899 3107 9903
rect 3111 9899 3112 9903
rect 3116 9899 3117 9903
rect 3121 9899 3122 9903
rect 3126 9899 3127 9903
rect 3131 9899 3132 9903
rect 3136 9899 3137 9903
rect 3141 9899 3142 9903
rect 3101 9898 3146 9899
rect 3101 9894 3102 9898
rect 3106 9894 3107 9898
rect 3111 9894 3112 9898
rect 3116 9894 3117 9898
rect 3121 9894 3122 9898
rect 3126 9894 3127 9898
rect 3131 9894 3132 9898
rect 3136 9894 3137 9898
rect 3141 9894 3142 9898
rect 3101 9893 3146 9894
rect 3101 9889 3102 9893
rect 3106 9889 3107 9893
rect 3111 9889 3112 9893
rect 3116 9889 3117 9893
rect 3121 9889 3122 9893
rect 3126 9889 3127 9893
rect 3131 9889 3132 9893
rect 3136 9889 3137 9893
rect 3141 9889 3142 9893
rect 3101 9888 3146 9889
rect 3101 9884 3102 9888
rect 3106 9884 3107 9888
rect 3111 9884 3112 9888
rect 3116 9884 3117 9888
rect 3121 9884 3122 9888
rect 3126 9884 3127 9888
rect 3131 9884 3132 9888
rect 3136 9884 3137 9888
rect 3141 9884 3142 9888
rect 3101 9883 3146 9884
rect 3101 9879 3102 9883
rect 3106 9879 3107 9883
rect 3111 9879 3112 9883
rect 3116 9879 3117 9883
rect 3121 9879 3122 9883
rect 3126 9879 3127 9883
rect 3131 9879 3132 9883
rect 3136 9879 3137 9883
rect 3141 9879 3142 9883
rect 3101 9878 3146 9879
rect 3101 9874 3102 9878
rect 3106 9874 3107 9878
rect 3111 9874 3112 9878
rect 3116 9874 3117 9878
rect 3121 9874 3122 9878
rect 3126 9874 3127 9878
rect 3131 9874 3132 9878
rect 3136 9874 3137 9878
rect 3141 9874 3142 9878
rect 3101 9873 3146 9874
rect 3101 9869 3102 9873
rect 3106 9869 3107 9873
rect 3111 9869 3112 9873
rect 3116 9869 3117 9873
rect 3121 9869 3122 9873
rect 3126 9869 3127 9873
rect 3131 9869 3132 9873
rect 3136 9869 3137 9873
rect 3141 9869 3142 9873
rect 3101 9868 3146 9869
rect 3101 9864 3102 9868
rect 3106 9864 3107 9868
rect 3111 9864 3112 9868
rect 3116 9864 3117 9868
rect 3121 9864 3122 9868
rect 3126 9864 3127 9868
rect 3131 9864 3132 9868
rect 3136 9864 3137 9868
rect 3141 9864 3142 9868
rect 3154 9948 3158 9949
rect 3154 9943 3158 9944
rect 3154 9938 3158 9939
rect 3154 9933 3158 9934
rect 3154 9928 3158 9929
rect 3154 9923 3158 9924
rect 3154 9918 3158 9919
rect 3154 9913 3158 9914
rect 3154 9908 3158 9909
rect 3154 9903 3158 9904
rect 3154 9898 3158 9899
rect 3154 9893 3158 9894
rect 3154 9888 3158 9889
rect 3154 9883 3158 9884
rect 3154 9878 3158 9879
rect 3154 9873 3158 9874
rect 3154 9868 3158 9869
rect 3090 9863 3094 9864
rect 3090 9856 3094 9859
rect 3154 9863 3158 9864
rect 3154 9856 3158 9859
rect 3094 9848 3097 9856
rect 3101 9848 3102 9856
rect 3106 9848 3107 9856
rect 3111 9848 3112 9856
rect 3116 9848 3117 9856
rect 3121 9848 3122 9856
rect 3126 9848 3127 9856
rect 3131 9848 3132 9856
rect 3136 9848 3137 9856
rect 3141 9848 3142 9856
rect 3146 9848 3147 9856
rect 3151 9848 3154 9856
rect 3167 9963 3171 9964
rect 3167 9958 3171 9959
rect 3167 9953 3171 9954
rect 3167 9948 3171 9949
rect 3167 9943 3171 9944
rect 3167 9938 3171 9939
rect 3167 9933 3171 9934
rect 3167 9928 3171 9929
rect 3167 9923 3171 9924
rect 3167 9918 3171 9919
rect 3167 9913 3171 9914
rect 3167 9908 3171 9909
rect 3167 9903 3171 9904
rect 3167 9898 3171 9899
rect 3167 9893 3171 9894
rect 3167 9888 3171 9889
rect 3167 9883 3171 9884
rect 3167 9878 3171 9879
rect 3167 9873 3171 9874
rect 3167 9868 3171 9869
rect 3167 9863 3171 9864
rect 3167 9858 3171 9859
rect 3167 9853 3171 9854
rect 3167 9848 3171 9849
rect 3035 9844 3052 9846
rect 3007 9843 3011 9844
rect 2921 9839 2922 9843
rect 2926 9839 2927 9843
rect 2931 9839 2932 9843
rect 2936 9839 2937 9843
rect 2941 9839 2942 9843
rect 2946 9839 2947 9843
rect 2951 9839 2952 9843
rect 2956 9839 2957 9843
rect 2961 9839 2962 9843
rect 2966 9839 2967 9843
rect 2971 9839 2972 9843
rect 2976 9839 2977 9843
rect 2981 9839 2982 9843
rect 2986 9839 2987 9843
rect 2991 9839 2992 9843
rect 2996 9839 2997 9843
rect 3001 9839 3002 9843
rect 3006 9839 3007 9843
rect 3037 9842 3050 9844
rect 3077 9843 3081 9844
rect 3167 9843 3171 9844
rect 2805 9831 2861 9839
rect 2611 9827 2670 9831
rect 2796 9827 2861 9831
rect 2611 9815 2667 9827
rect 2726 9819 2756 9823
rect 2611 9811 2670 9815
rect 2740 9812 2744 9819
rect 2805 9815 2861 9827
rect 2611 9802 2667 9811
rect 2796 9811 2861 9815
rect 2726 9803 2737 9807
rect 2487 9795 2552 9799
rect 2290 9790 2358 9791
rect 2290 9786 2291 9790
rect 2295 9786 2296 9790
rect 2300 9786 2358 9790
rect 2417 9787 2447 9791
rect 2290 9785 2358 9786
rect 2290 9781 2291 9785
rect 2295 9781 2296 9785
rect 2300 9783 2358 9785
rect 2300 9781 2361 9783
rect 2290 9780 2361 9781
rect 2290 9776 2291 9780
rect 2295 9776 2296 9780
rect 2300 9779 2361 9780
rect 2300 9776 2358 9779
rect 2290 9775 2358 9776
rect 2290 9771 2291 9775
rect 2295 9771 2296 9775
rect 2300 9771 2358 9775
rect 2290 9770 2358 9771
rect 2290 9766 2291 9770
rect 2295 9766 2296 9770
rect 2300 9766 2358 9770
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2246 9761 2265 9762
rect 2250 9757 2251 9761
rect 2255 9757 2256 9761
rect 2260 9757 2261 9761
rect 2246 9756 2265 9757
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2246 9751 2265 9752
rect 2250 9747 2251 9751
rect 2255 9747 2256 9751
rect 2260 9747 2261 9751
rect 2246 9746 2265 9747
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2246 9741 2265 9742
rect 2250 9737 2251 9741
rect 2255 9737 2256 9741
rect 2260 9737 2261 9741
rect 2246 9736 2265 9737
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2290 9765 2358 9766
rect 2290 9761 2291 9765
rect 2295 9761 2296 9765
rect 2300 9761 2358 9765
rect 2290 9760 2358 9761
rect 2290 9756 2291 9760
rect 2295 9756 2296 9760
rect 2300 9756 2358 9760
rect 2290 9755 2358 9756
rect 2290 9751 2291 9755
rect 2295 9751 2296 9755
rect 2300 9751 2358 9755
rect 2290 9750 2358 9751
rect 2290 9746 2291 9750
rect 2295 9746 2296 9750
rect 2300 9746 2358 9750
rect 2290 9745 2358 9746
rect 2290 9741 2291 9745
rect 2295 9741 2296 9745
rect 2300 9741 2358 9745
rect 2290 9740 2358 9741
rect 2290 9736 2291 9740
rect 2295 9736 2296 9740
rect 2300 9736 2358 9740
rect 2290 9734 2358 9736
rect 2191 9718 2192 9722
rect 2196 9718 2197 9722
rect 2201 9718 2202 9722
rect 2206 9718 2207 9722
rect 2211 9718 2212 9722
rect 2216 9718 2217 9722
rect 2221 9718 2222 9722
rect 2226 9718 2227 9722
rect 2231 9718 2232 9722
rect 2236 9718 2237 9722
rect 2241 9718 2243 9722
rect 2187 9717 2243 9718
rect 2191 9713 2192 9717
rect 2196 9713 2197 9717
rect 2201 9713 2202 9717
rect 2206 9713 2207 9717
rect 2211 9713 2212 9717
rect 2216 9713 2217 9717
rect 2221 9713 2222 9717
rect 2226 9713 2227 9717
rect 2231 9713 2232 9717
rect 2236 9713 2237 9717
rect 2241 9713 2243 9717
rect 2187 9712 2243 9713
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2246 9715 2265 9716
rect 2250 9711 2251 9715
rect 2255 9711 2256 9715
rect 2260 9711 2261 9715
rect 2246 9710 2265 9711
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2246 9705 2265 9706
rect 2250 9701 2251 9705
rect 2255 9701 2256 9705
rect 2260 9701 2261 9705
rect 2246 9700 2265 9701
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2246 9695 2265 9696
rect 2250 9691 2251 9695
rect 2255 9691 2256 9695
rect 2260 9691 2261 9695
rect 2246 9690 2265 9691
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2422 9597 2435 9787
rect 2496 9783 2552 9795
rect 2487 9779 2552 9783
rect 2496 9722 2552 9779
rect 2599 9800 2667 9802
rect 2599 9796 2600 9800
rect 2604 9796 2605 9800
rect 2609 9799 2667 9800
rect 2730 9800 2737 9803
rect 2749 9803 2756 9807
rect 2749 9800 2753 9803
rect 2609 9796 2670 9799
rect 2599 9795 2670 9796
rect 2599 9791 2600 9795
rect 2604 9791 2605 9795
rect 2609 9791 2667 9795
rect 2730 9791 2753 9800
rect 2805 9799 2861 9811
rect 2920 9831 2976 9839
rect 3039 9831 3048 9842
rect 3081 9839 3082 9843
rect 3086 9839 3087 9843
rect 3091 9839 3092 9843
rect 3096 9839 3097 9843
rect 3101 9839 3102 9843
rect 3106 9839 3107 9843
rect 3111 9839 3112 9843
rect 3116 9839 3117 9843
rect 3121 9839 3122 9843
rect 3126 9839 3127 9843
rect 3131 9839 3132 9843
rect 3136 9839 3137 9843
rect 3141 9839 3142 9843
rect 3146 9839 3147 9843
rect 3151 9839 3152 9843
rect 3156 9839 3157 9843
rect 3161 9839 3162 9843
rect 3166 9839 3167 9843
rect 3230 9974 3231 9978
rect 3235 9974 3236 9978
rect 3240 9974 3241 9978
rect 3245 9974 3246 9978
rect 3250 9974 3251 9978
rect 3255 9974 3256 9978
rect 3260 9974 3261 9978
rect 3265 9974 3266 9978
rect 3270 9974 3271 9978
rect 3275 9974 3276 9978
rect 3280 9974 3281 9978
rect 3285 9974 3286 9978
rect 3290 9974 3291 9978
rect 3295 9974 3296 9978
rect 3300 9974 3301 9978
rect 3305 9974 3306 9978
rect 3310 9974 3311 9978
rect 3315 9974 3316 9978
rect 3226 9973 3230 9974
rect 3226 9968 3230 9969
rect 3316 9973 3320 9974
rect 3316 9968 3320 9969
rect 3226 9963 3230 9964
rect 3226 9958 3230 9959
rect 3226 9953 3230 9954
rect 3226 9948 3230 9949
rect 3226 9943 3230 9944
rect 3226 9938 3230 9939
rect 3226 9933 3230 9934
rect 3226 9928 3230 9929
rect 3226 9923 3230 9924
rect 3226 9918 3230 9919
rect 3226 9913 3230 9914
rect 3226 9908 3230 9909
rect 3226 9903 3230 9904
rect 3226 9898 3230 9899
rect 3226 9893 3230 9894
rect 3226 9888 3230 9889
rect 3226 9883 3230 9884
rect 3226 9878 3230 9879
rect 3226 9873 3230 9874
rect 3226 9868 3230 9869
rect 3226 9863 3230 9864
rect 3226 9858 3230 9859
rect 3226 9853 3230 9854
rect 3226 9848 3230 9849
rect 3243 9961 3246 9965
rect 3250 9961 3251 9965
rect 3255 9961 3256 9965
rect 3260 9961 3261 9965
rect 3265 9961 3266 9965
rect 3270 9961 3271 9965
rect 3275 9961 3276 9965
rect 3280 9961 3281 9965
rect 3285 9961 3286 9965
rect 3290 9961 3291 9965
rect 3295 9961 3296 9965
rect 3300 9961 3303 9965
rect 3239 9958 3243 9961
rect 3239 9953 3243 9954
rect 3303 9958 3307 9961
rect 3303 9953 3307 9954
rect 3239 9948 3243 9949
rect 3239 9943 3243 9944
rect 3239 9938 3243 9939
rect 3239 9933 3243 9934
rect 3239 9928 3243 9929
rect 3239 9923 3243 9924
rect 3239 9918 3243 9919
rect 3239 9913 3243 9914
rect 3239 9908 3243 9909
rect 3239 9903 3243 9904
rect 3239 9898 3243 9899
rect 3239 9893 3243 9894
rect 3239 9888 3243 9889
rect 3239 9883 3243 9884
rect 3239 9878 3243 9879
rect 3239 9873 3243 9874
rect 3239 9868 3243 9869
rect 3255 9949 3256 9953
rect 3260 9949 3261 9953
rect 3265 9949 3266 9953
rect 3270 9949 3271 9953
rect 3275 9949 3276 9953
rect 3280 9949 3281 9953
rect 3285 9949 3286 9953
rect 3290 9949 3291 9953
rect 3251 9948 3295 9949
rect 3255 9944 3256 9948
rect 3260 9944 3261 9948
rect 3265 9944 3266 9948
rect 3270 9944 3271 9948
rect 3275 9944 3276 9948
rect 3280 9944 3281 9948
rect 3285 9944 3286 9948
rect 3290 9944 3291 9948
rect 3251 9943 3295 9944
rect 3255 9939 3256 9943
rect 3260 9939 3261 9943
rect 3265 9939 3266 9943
rect 3270 9939 3271 9943
rect 3275 9939 3276 9943
rect 3280 9939 3281 9943
rect 3285 9939 3286 9943
rect 3290 9939 3291 9943
rect 3251 9938 3295 9939
rect 3255 9934 3256 9938
rect 3260 9934 3261 9938
rect 3265 9934 3266 9938
rect 3270 9934 3271 9938
rect 3275 9934 3276 9938
rect 3280 9934 3281 9938
rect 3285 9934 3286 9938
rect 3290 9934 3291 9938
rect 3251 9933 3295 9934
rect 3255 9929 3256 9933
rect 3260 9929 3261 9933
rect 3265 9929 3266 9933
rect 3270 9929 3271 9933
rect 3275 9929 3276 9933
rect 3280 9929 3281 9933
rect 3285 9929 3286 9933
rect 3290 9929 3291 9933
rect 3251 9928 3295 9929
rect 3255 9924 3256 9928
rect 3260 9924 3261 9928
rect 3265 9924 3266 9928
rect 3270 9924 3271 9928
rect 3275 9924 3276 9928
rect 3280 9924 3281 9928
rect 3285 9924 3286 9928
rect 3290 9924 3291 9928
rect 3251 9923 3295 9924
rect 3255 9919 3256 9923
rect 3260 9919 3261 9923
rect 3265 9919 3266 9923
rect 3270 9919 3271 9923
rect 3275 9919 3276 9923
rect 3280 9919 3281 9923
rect 3285 9919 3286 9923
rect 3290 9919 3291 9923
rect 3251 9918 3295 9919
rect 3255 9914 3256 9918
rect 3260 9914 3261 9918
rect 3265 9914 3266 9918
rect 3270 9914 3271 9918
rect 3275 9914 3276 9918
rect 3280 9914 3281 9918
rect 3285 9914 3286 9918
rect 3290 9914 3291 9918
rect 3251 9913 3295 9914
rect 3255 9909 3256 9913
rect 3260 9909 3261 9913
rect 3265 9909 3266 9913
rect 3270 9909 3271 9913
rect 3275 9909 3276 9913
rect 3280 9909 3281 9913
rect 3285 9909 3286 9913
rect 3290 9909 3291 9913
rect 3251 9908 3295 9909
rect 3255 9904 3256 9908
rect 3260 9904 3261 9908
rect 3265 9904 3266 9908
rect 3270 9904 3271 9908
rect 3275 9904 3276 9908
rect 3280 9904 3281 9908
rect 3285 9904 3286 9908
rect 3290 9904 3291 9908
rect 3251 9903 3295 9904
rect 3255 9899 3256 9903
rect 3260 9899 3261 9903
rect 3265 9899 3266 9903
rect 3270 9899 3271 9903
rect 3275 9899 3276 9903
rect 3280 9899 3281 9903
rect 3285 9899 3286 9903
rect 3290 9899 3291 9903
rect 3251 9898 3295 9899
rect 3255 9894 3256 9898
rect 3260 9894 3261 9898
rect 3265 9894 3266 9898
rect 3270 9894 3271 9898
rect 3275 9894 3276 9898
rect 3280 9894 3281 9898
rect 3285 9894 3286 9898
rect 3290 9894 3291 9898
rect 3251 9893 3295 9894
rect 3255 9889 3256 9893
rect 3260 9889 3261 9893
rect 3265 9889 3266 9893
rect 3270 9889 3271 9893
rect 3275 9889 3276 9893
rect 3280 9889 3281 9893
rect 3285 9889 3286 9893
rect 3290 9889 3291 9893
rect 3251 9888 3295 9889
rect 3255 9884 3256 9888
rect 3260 9884 3261 9888
rect 3265 9884 3266 9888
rect 3270 9884 3271 9888
rect 3275 9884 3276 9888
rect 3280 9884 3281 9888
rect 3285 9884 3286 9888
rect 3290 9884 3291 9888
rect 3251 9883 3295 9884
rect 3255 9879 3256 9883
rect 3260 9879 3261 9883
rect 3265 9879 3266 9883
rect 3270 9879 3271 9883
rect 3275 9879 3276 9883
rect 3280 9879 3281 9883
rect 3285 9879 3286 9883
rect 3290 9879 3291 9883
rect 3251 9878 3295 9879
rect 3255 9874 3256 9878
rect 3260 9874 3261 9878
rect 3265 9874 3266 9878
rect 3270 9874 3271 9878
rect 3275 9874 3276 9878
rect 3280 9874 3281 9878
rect 3285 9874 3286 9878
rect 3290 9874 3291 9878
rect 3251 9873 3295 9874
rect 3255 9869 3256 9873
rect 3260 9869 3261 9873
rect 3265 9869 3266 9873
rect 3270 9869 3271 9873
rect 3275 9869 3276 9873
rect 3280 9869 3281 9873
rect 3285 9869 3286 9873
rect 3290 9869 3291 9873
rect 3251 9868 3295 9869
rect 3255 9864 3256 9868
rect 3260 9864 3261 9868
rect 3265 9864 3266 9868
rect 3270 9864 3271 9868
rect 3275 9864 3276 9868
rect 3280 9864 3281 9868
rect 3285 9864 3286 9868
rect 3290 9864 3291 9868
rect 3303 9948 3307 9949
rect 3303 9943 3307 9944
rect 3303 9938 3307 9939
rect 3303 9933 3307 9934
rect 3303 9928 3307 9929
rect 3303 9923 3307 9924
rect 3303 9918 3307 9919
rect 3303 9913 3307 9914
rect 3303 9908 3307 9909
rect 3303 9903 3307 9904
rect 3303 9898 3307 9899
rect 3303 9893 3307 9894
rect 3303 9888 3307 9889
rect 3303 9883 3307 9884
rect 3303 9878 3307 9879
rect 3303 9873 3307 9874
rect 3303 9868 3307 9869
rect 3239 9863 3243 9864
rect 3239 9856 3243 9859
rect 3303 9863 3307 9864
rect 3303 9856 3307 9859
rect 3243 9848 3246 9856
rect 3250 9848 3251 9856
rect 3255 9848 3256 9856
rect 3260 9848 3261 9856
rect 3265 9848 3266 9856
rect 3270 9848 3271 9856
rect 3275 9848 3276 9856
rect 3280 9848 3281 9856
rect 3285 9848 3286 9856
rect 3290 9848 3291 9856
rect 3295 9848 3296 9856
rect 3300 9848 3303 9856
rect 3316 9963 3320 9964
rect 3316 9958 3320 9959
rect 3316 9953 3320 9954
rect 3316 9948 3320 9949
rect 3316 9943 3320 9944
rect 3316 9938 3320 9939
rect 3316 9933 3320 9934
rect 3316 9928 3320 9929
rect 3316 9923 3320 9924
rect 3316 9918 3320 9919
rect 3316 9913 3320 9914
rect 3316 9908 3320 9909
rect 3316 9903 3320 9904
rect 3316 9898 3320 9899
rect 3316 9893 3320 9894
rect 3316 9888 3320 9889
rect 3316 9883 3320 9884
rect 3316 9878 3320 9879
rect 3316 9873 3320 9874
rect 3316 9868 3320 9869
rect 3316 9863 3320 9864
rect 3316 9858 3320 9859
rect 3316 9853 3320 9854
rect 3316 9848 3320 9849
rect 3226 9843 3230 9844
rect 3316 9843 3320 9844
rect 3230 9839 3231 9843
rect 3235 9839 3236 9843
rect 3240 9839 3241 9843
rect 3245 9839 3246 9843
rect 3250 9839 3251 9843
rect 3255 9839 3256 9843
rect 3260 9839 3261 9843
rect 3265 9839 3266 9843
rect 3270 9839 3271 9843
rect 3275 9839 3276 9843
rect 3280 9839 3281 9843
rect 3285 9839 3286 9843
rect 3290 9839 3291 9843
rect 3295 9839 3296 9843
rect 3300 9839 3301 9843
rect 3305 9839 3306 9843
rect 3310 9839 3311 9843
rect 3315 9839 3316 9843
rect 3114 9831 3170 9839
rect 2920 9827 2979 9831
rect 3105 9827 3170 9831
rect 2920 9815 2976 9827
rect 3035 9819 3065 9823
rect 2920 9811 2979 9815
rect 3049 9812 3053 9819
rect 3114 9815 3170 9827
rect 2920 9802 2976 9811
rect 3105 9811 3170 9815
rect 3035 9803 3046 9807
rect 2796 9795 2861 9799
rect 2599 9790 2667 9791
rect 2599 9786 2600 9790
rect 2604 9786 2605 9790
rect 2609 9786 2667 9790
rect 2726 9787 2756 9791
rect 2599 9785 2667 9786
rect 2599 9781 2600 9785
rect 2604 9781 2605 9785
rect 2609 9783 2667 9785
rect 2609 9781 2670 9783
rect 2599 9780 2670 9781
rect 2599 9776 2600 9780
rect 2604 9776 2605 9780
rect 2609 9779 2670 9780
rect 2609 9776 2667 9779
rect 2599 9775 2667 9776
rect 2599 9771 2600 9775
rect 2604 9771 2605 9775
rect 2609 9771 2667 9775
rect 2599 9770 2667 9771
rect 2599 9766 2600 9770
rect 2604 9766 2605 9770
rect 2609 9766 2667 9770
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2555 9761 2574 9762
rect 2559 9757 2560 9761
rect 2564 9757 2565 9761
rect 2569 9757 2570 9761
rect 2555 9756 2574 9757
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2555 9751 2574 9752
rect 2559 9747 2560 9751
rect 2564 9747 2565 9751
rect 2569 9747 2570 9751
rect 2555 9746 2574 9747
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2555 9741 2574 9742
rect 2559 9737 2560 9741
rect 2564 9737 2565 9741
rect 2569 9737 2570 9741
rect 2555 9736 2574 9737
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2599 9765 2667 9766
rect 2599 9761 2600 9765
rect 2604 9761 2605 9765
rect 2609 9761 2667 9765
rect 2599 9760 2667 9761
rect 2599 9756 2600 9760
rect 2604 9756 2605 9760
rect 2609 9756 2667 9760
rect 2599 9755 2667 9756
rect 2599 9751 2600 9755
rect 2604 9751 2605 9755
rect 2609 9751 2667 9755
rect 2599 9750 2667 9751
rect 2599 9746 2600 9750
rect 2604 9746 2605 9750
rect 2609 9746 2667 9750
rect 2599 9745 2667 9746
rect 2599 9741 2600 9745
rect 2604 9741 2605 9745
rect 2609 9741 2667 9745
rect 2599 9740 2667 9741
rect 2599 9736 2600 9740
rect 2604 9736 2605 9740
rect 2609 9736 2667 9740
rect 2599 9734 2667 9736
rect 2500 9718 2501 9722
rect 2505 9718 2506 9722
rect 2510 9718 2511 9722
rect 2515 9718 2516 9722
rect 2520 9718 2521 9722
rect 2525 9718 2526 9722
rect 2530 9718 2531 9722
rect 2535 9718 2536 9722
rect 2540 9718 2541 9722
rect 2545 9718 2546 9722
rect 2550 9718 2552 9722
rect 2496 9717 2552 9718
rect 2500 9713 2501 9717
rect 2505 9713 2506 9717
rect 2510 9713 2511 9717
rect 2515 9713 2516 9717
rect 2520 9713 2521 9717
rect 2525 9713 2526 9717
rect 2530 9713 2531 9717
rect 2535 9713 2536 9717
rect 2540 9713 2541 9717
rect 2545 9713 2546 9717
rect 2550 9713 2552 9717
rect 2496 9712 2552 9713
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2555 9715 2574 9716
rect 2559 9711 2560 9715
rect 2564 9711 2565 9715
rect 2569 9711 2570 9715
rect 2555 9710 2574 9711
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2555 9705 2574 9706
rect 2559 9701 2560 9705
rect 2564 9701 2565 9705
rect 2569 9701 2570 9705
rect 2555 9700 2574 9701
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2555 9695 2574 9696
rect 2559 9691 2560 9695
rect 2564 9691 2565 9695
rect 2569 9691 2570 9695
rect 2555 9690 2574 9691
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2731 9609 2744 9787
rect 2805 9783 2861 9795
rect 2796 9779 2861 9783
rect 2805 9722 2861 9779
rect 2908 9800 2976 9802
rect 2908 9796 2909 9800
rect 2913 9796 2914 9800
rect 2918 9799 2976 9800
rect 3039 9800 3046 9803
rect 3058 9803 3065 9807
rect 3058 9800 3062 9803
rect 2918 9796 2979 9799
rect 2908 9795 2979 9796
rect 2908 9791 2909 9795
rect 2913 9791 2914 9795
rect 2918 9791 2976 9795
rect 3039 9791 3062 9800
rect 3114 9799 3170 9811
rect 3229 9802 3285 9839
rect 3105 9795 3170 9799
rect 2908 9790 2976 9791
rect 2908 9786 2909 9790
rect 2913 9786 2914 9790
rect 2918 9786 2976 9790
rect 3035 9787 3065 9791
rect 2908 9785 2976 9786
rect 2908 9781 2909 9785
rect 2913 9781 2914 9785
rect 2918 9783 2976 9785
rect 2918 9781 2979 9783
rect 2908 9780 2979 9781
rect 2908 9776 2909 9780
rect 2913 9776 2914 9780
rect 2918 9779 2979 9780
rect 2918 9776 2976 9779
rect 2908 9775 2976 9776
rect 2908 9771 2909 9775
rect 2913 9771 2914 9775
rect 2918 9771 2976 9775
rect 2908 9770 2976 9771
rect 2908 9766 2909 9770
rect 2913 9766 2914 9770
rect 2918 9766 2976 9770
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2864 9761 2883 9762
rect 2868 9757 2869 9761
rect 2873 9757 2874 9761
rect 2878 9757 2879 9761
rect 2864 9756 2883 9757
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2864 9751 2883 9752
rect 2868 9747 2869 9751
rect 2873 9747 2874 9751
rect 2878 9747 2879 9751
rect 2864 9746 2883 9747
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2864 9741 2883 9742
rect 2868 9737 2869 9741
rect 2873 9737 2874 9741
rect 2878 9737 2879 9741
rect 2864 9736 2883 9737
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2908 9765 2976 9766
rect 2908 9761 2909 9765
rect 2913 9761 2914 9765
rect 2918 9761 2976 9765
rect 2908 9760 2976 9761
rect 2908 9756 2909 9760
rect 2913 9756 2914 9760
rect 2918 9756 2976 9760
rect 2908 9755 2976 9756
rect 2908 9751 2909 9755
rect 2913 9751 2914 9755
rect 2918 9751 2976 9755
rect 2908 9750 2976 9751
rect 2908 9746 2909 9750
rect 2913 9746 2914 9750
rect 2918 9746 2976 9750
rect 2908 9745 2976 9746
rect 2908 9741 2909 9745
rect 2913 9741 2914 9745
rect 2918 9741 2976 9745
rect 2908 9740 2976 9741
rect 2908 9736 2909 9740
rect 2913 9736 2914 9740
rect 2918 9736 2976 9740
rect 2908 9734 2976 9736
rect 2809 9718 2810 9722
rect 2814 9718 2815 9722
rect 2819 9718 2820 9722
rect 2824 9718 2825 9722
rect 2829 9718 2830 9722
rect 2834 9718 2835 9722
rect 2839 9718 2840 9722
rect 2844 9718 2845 9722
rect 2849 9718 2850 9722
rect 2854 9718 2855 9722
rect 2859 9718 2861 9722
rect 2805 9717 2861 9718
rect 2809 9713 2810 9717
rect 2814 9713 2815 9717
rect 2819 9713 2820 9717
rect 2824 9713 2825 9717
rect 2829 9713 2830 9717
rect 2834 9713 2835 9717
rect 2839 9713 2840 9717
rect 2844 9713 2845 9717
rect 2849 9713 2850 9717
rect 2854 9713 2855 9717
rect 2859 9713 2861 9717
rect 2805 9712 2861 9713
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2864 9715 2883 9716
rect 2868 9711 2869 9715
rect 2873 9711 2874 9715
rect 2878 9711 2879 9715
rect 2864 9710 2883 9711
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2864 9705 2883 9706
rect 2868 9701 2869 9705
rect 2873 9701 2874 9705
rect 2878 9701 2879 9705
rect 2864 9700 2883 9701
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2864 9695 2883 9696
rect 2868 9691 2869 9695
rect 2873 9691 2874 9695
rect 2878 9691 2879 9695
rect 2864 9690 2883 9691
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 3040 9611 3053 9787
rect 3114 9783 3170 9795
rect 3105 9779 3170 9783
rect 3114 9722 3170 9779
rect 3217 9800 3285 9802
rect 3217 9796 3218 9800
rect 3222 9796 3223 9800
rect 3227 9796 3285 9800
rect 3217 9795 3285 9796
rect 3217 9791 3218 9795
rect 3222 9791 3223 9795
rect 3227 9791 3285 9795
rect 3217 9790 3285 9791
rect 3217 9786 3218 9790
rect 3222 9786 3223 9790
rect 3227 9786 3285 9790
rect 3217 9785 3285 9786
rect 3217 9781 3218 9785
rect 3222 9781 3223 9785
rect 3227 9781 3285 9785
rect 3217 9780 3285 9781
rect 3217 9776 3218 9780
rect 3222 9776 3223 9780
rect 3227 9776 3285 9780
rect 3217 9775 3285 9776
rect 3217 9771 3218 9775
rect 3222 9771 3223 9775
rect 3227 9771 3285 9775
rect 3217 9770 3285 9771
rect 3217 9766 3218 9770
rect 3222 9766 3223 9770
rect 3227 9766 3285 9770
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3173 9761 3192 9762
rect 3177 9757 3178 9761
rect 3182 9757 3183 9761
rect 3187 9757 3188 9761
rect 3173 9756 3192 9757
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3173 9751 3192 9752
rect 3177 9747 3178 9751
rect 3182 9747 3183 9751
rect 3187 9747 3188 9751
rect 3173 9746 3192 9747
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3173 9741 3192 9742
rect 3177 9737 3178 9741
rect 3182 9737 3183 9741
rect 3187 9737 3188 9741
rect 3173 9736 3192 9737
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3217 9765 3285 9766
rect 3217 9761 3218 9765
rect 3222 9761 3223 9765
rect 3227 9761 3285 9765
rect 3217 9760 3285 9761
rect 3217 9756 3218 9760
rect 3222 9756 3223 9760
rect 3227 9756 3285 9760
rect 3217 9755 3285 9756
rect 3217 9751 3218 9755
rect 3222 9751 3223 9755
rect 3227 9751 3285 9755
rect 3217 9750 3285 9751
rect 3217 9746 3218 9750
rect 3222 9746 3223 9750
rect 3227 9746 3285 9750
rect 3217 9745 3285 9746
rect 3217 9741 3218 9745
rect 3222 9741 3223 9745
rect 3227 9741 3285 9745
rect 3217 9740 3285 9741
rect 3217 9736 3218 9740
rect 3222 9736 3223 9740
rect 3227 9736 3285 9740
rect 3217 9734 3285 9736
rect 3118 9718 3119 9722
rect 3123 9718 3124 9722
rect 3128 9718 3129 9722
rect 3133 9718 3134 9722
rect 3138 9718 3139 9722
rect 3143 9718 3144 9722
rect 3148 9718 3149 9722
rect 3153 9718 3154 9722
rect 3158 9718 3159 9722
rect 3163 9718 3164 9722
rect 3168 9718 3170 9722
rect 3114 9717 3170 9718
rect 3118 9713 3119 9717
rect 3123 9713 3124 9717
rect 3128 9713 3129 9717
rect 3133 9713 3134 9717
rect 3138 9713 3139 9717
rect 3143 9713 3144 9717
rect 3148 9713 3149 9717
rect 3153 9713 3154 9717
rect 3158 9713 3159 9717
rect 3163 9713 3164 9717
rect 3168 9713 3170 9717
rect 3114 9712 3170 9713
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3173 9715 3192 9716
rect 3177 9711 3178 9715
rect 3182 9711 3183 9715
rect 3187 9711 3188 9715
rect 3173 9710 3192 9711
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3173 9705 3192 9706
rect 3177 9701 3178 9705
rect 3182 9701 3183 9705
rect 3187 9701 3188 9705
rect 3173 9700 3192 9701
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3173 9695 3192 9696
rect 3177 9691 3178 9695
rect 3182 9691 3183 9695
rect 3187 9691 3188 9695
rect 3173 9690 3192 9691
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3327 9715 3379 9981
rect 3390 9974 3391 9978
rect 3395 9974 3396 9978
rect 3400 9974 3401 9978
rect 3405 9974 3406 9978
rect 3410 9974 3411 9978
rect 3415 9974 3416 9978
rect 3420 9974 3421 9978
rect 3425 9974 3426 9978
rect 3430 9974 3431 9978
rect 3435 9974 3436 9978
rect 3440 9974 3441 9978
rect 3445 9974 3446 9978
rect 3450 9974 3451 9978
rect 3455 9974 3456 9978
rect 3460 9974 3461 9978
rect 3465 9974 3466 9978
rect 3470 9974 3471 9978
rect 3475 9974 3476 9978
rect 3386 9973 3390 9974
rect 3386 9968 3390 9969
rect 3476 9973 3480 9974
rect 3476 9968 3480 9969
rect 3386 9963 3390 9964
rect 3386 9958 3390 9959
rect 3386 9953 3390 9954
rect 3386 9948 3390 9949
rect 3386 9943 3390 9944
rect 3386 9938 3390 9939
rect 3386 9933 3390 9934
rect 3386 9928 3390 9929
rect 3386 9923 3390 9924
rect 3386 9918 3390 9919
rect 3386 9913 3390 9914
rect 3386 9908 3390 9909
rect 3386 9903 3390 9904
rect 3386 9898 3390 9899
rect 3386 9893 3390 9894
rect 3386 9888 3390 9889
rect 3386 9883 3390 9884
rect 3386 9878 3390 9879
rect 3386 9873 3390 9874
rect 3386 9868 3390 9869
rect 3386 9863 3390 9864
rect 3386 9858 3390 9859
rect 3386 9853 3390 9854
rect 3386 9848 3390 9849
rect 3403 9961 3406 9965
rect 3410 9961 3411 9965
rect 3415 9961 3416 9965
rect 3420 9961 3421 9965
rect 3425 9961 3426 9965
rect 3430 9961 3431 9965
rect 3435 9961 3436 9965
rect 3440 9961 3441 9965
rect 3445 9961 3446 9965
rect 3450 9961 3451 9965
rect 3455 9961 3456 9965
rect 3460 9961 3463 9965
rect 3399 9958 3403 9961
rect 3399 9953 3403 9954
rect 3463 9958 3467 9961
rect 3463 9953 3467 9954
rect 3399 9948 3403 9949
rect 3399 9943 3403 9944
rect 3399 9938 3403 9939
rect 3399 9933 3403 9934
rect 3399 9928 3403 9929
rect 3399 9923 3403 9924
rect 3399 9918 3403 9919
rect 3399 9913 3403 9914
rect 3399 9908 3403 9909
rect 3399 9903 3403 9904
rect 3399 9898 3403 9899
rect 3399 9893 3403 9894
rect 3399 9888 3403 9889
rect 3399 9883 3403 9884
rect 3399 9878 3403 9879
rect 3399 9873 3403 9874
rect 3399 9868 3403 9869
rect 3410 9949 3411 9953
rect 3415 9949 3416 9953
rect 3420 9949 3421 9953
rect 3425 9949 3426 9953
rect 3430 9949 3431 9953
rect 3435 9949 3436 9953
rect 3440 9949 3441 9953
rect 3445 9949 3446 9953
rect 3450 9949 3451 9953
rect 3410 9948 3455 9949
rect 3410 9944 3411 9948
rect 3415 9944 3416 9948
rect 3420 9944 3421 9948
rect 3425 9944 3426 9948
rect 3430 9944 3431 9948
rect 3435 9944 3436 9948
rect 3440 9944 3441 9948
rect 3445 9944 3446 9948
rect 3450 9944 3451 9948
rect 3410 9943 3455 9944
rect 3410 9939 3411 9943
rect 3415 9939 3416 9943
rect 3420 9939 3421 9943
rect 3425 9939 3426 9943
rect 3430 9939 3431 9943
rect 3435 9939 3436 9943
rect 3440 9939 3441 9943
rect 3445 9939 3446 9943
rect 3450 9939 3451 9943
rect 3410 9938 3455 9939
rect 3410 9934 3411 9938
rect 3415 9934 3416 9938
rect 3420 9934 3421 9938
rect 3425 9934 3426 9938
rect 3430 9934 3431 9938
rect 3435 9934 3436 9938
rect 3440 9934 3441 9938
rect 3445 9934 3446 9938
rect 3450 9934 3451 9938
rect 3410 9933 3455 9934
rect 3410 9929 3411 9933
rect 3415 9929 3416 9933
rect 3420 9929 3421 9933
rect 3425 9929 3426 9933
rect 3430 9929 3431 9933
rect 3435 9929 3436 9933
rect 3440 9929 3441 9933
rect 3445 9929 3446 9933
rect 3450 9929 3451 9933
rect 3410 9928 3455 9929
rect 3410 9924 3411 9928
rect 3415 9924 3416 9928
rect 3420 9924 3421 9928
rect 3425 9924 3426 9928
rect 3430 9924 3431 9928
rect 3435 9924 3436 9928
rect 3440 9924 3441 9928
rect 3445 9924 3446 9928
rect 3450 9924 3451 9928
rect 3410 9923 3455 9924
rect 3410 9919 3411 9923
rect 3415 9919 3416 9923
rect 3420 9919 3421 9923
rect 3425 9919 3426 9923
rect 3430 9919 3431 9923
rect 3435 9919 3436 9923
rect 3440 9919 3441 9923
rect 3445 9919 3446 9923
rect 3450 9919 3451 9923
rect 3410 9918 3455 9919
rect 3410 9914 3411 9918
rect 3415 9914 3416 9918
rect 3420 9914 3421 9918
rect 3425 9914 3426 9918
rect 3430 9914 3431 9918
rect 3435 9914 3436 9918
rect 3440 9914 3441 9918
rect 3445 9914 3446 9918
rect 3450 9914 3451 9918
rect 3410 9913 3455 9914
rect 3410 9909 3411 9913
rect 3415 9909 3416 9913
rect 3420 9909 3421 9913
rect 3425 9909 3426 9913
rect 3430 9909 3431 9913
rect 3435 9909 3436 9913
rect 3440 9909 3441 9913
rect 3445 9909 3446 9913
rect 3450 9909 3451 9913
rect 3410 9908 3455 9909
rect 3410 9904 3411 9908
rect 3415 9904 3416 9908
rect 3420 9904 3421 9908
rect 3425 9904 3426 9908
rect 3430 9904 3431 9908
rect 3435 9904 3436 9908
rect 3440 9904 3441 9908
rect 3445 9904 3446 9908
rect 3450 9904 3451 9908
rect 3410 9903 3455 9904
rect 3410 9899 3411 9903
rect 3415 9899 3416 9903
rect 3420 9899 3421 9903
rect 3425 9899 3426 9903
rect 3430 9899 3431 9903
rect 3435 9899 3436 9903
rect 3440 9899 3441 9903
rect 3445 9899 3446 9903
rect 3450 9899 3451 9903
rect 3410 9898 3455 9899
rect 3410 9894 3411 9898
rect 3415 9894 3416 9898
rect 3420 9894 3421 9898
rect 3425 9894 3426 9898
rect 3430 9894 3431 9898
rect 3435 9894 3436 9898
rect 3440 9894 3441 9898
rect 3445 9894 3446 9898
rect 3450 9894 3451 9898
rect 3410 9893 3455 9894
rect 3410 9889 3411 9893
rect 3415 9889 3416 9893
rect 3420 9889 3421 9893
rect 3425 9889 3426 9893
rect 3430 9889 3431 9893
rect 3435 9889 3436 9893
rect 3440 9889 3441 9893
rect 3445 9889 3446 9893
rect 3450 9889 3451 9893
rect 3410 9888 3455 9889
rect 3410 9884 3411 9888
rect 3415 9884 3416 9888
rect 3420 9884 3421 9888
rect 3425 9884 3426 9888
rect 3430 9884 3431 9888
rect 3435 9884 3436 9888
rect 3440 9884 3441 9888
rect 3445 9884 3446 9888
rect 3450 9884 3451 9888
rect 3410 9883 3455 9884
rect 3410 9879 3411 9883
rect 3415 9879 3416 9883
rect 3420 9879 3421 9883
rect 3425 9879 3426 9883
rect 3430 9879 3431 9883
rect 3435 9879 3436 9883
rect 3440 9879 3441 9883
rect 3445 9879 3446 9883
rect 3450 9879 3451 9883
rect 3410 9878 3455 9879
rect 3410 9874 3411 9878
rect 3415 9874 3416 9878
rect 3420 9874 3421 9878
rect 3425 9874 3426 9878
rect 3430 9874 3431 9878
rect 3435 9874 3436 9878
rect 3440 9874 3441 9878
rect 3445 9874 3446 9878
rect 3450 9874 3451 9878
rect 3410 9873 3455 9874
rect 3410 9869 3411 9873
rect 3415 9869 3416 9873
rect 3420 9869 3421 9873
rect 3425 9869 3426 9873
rect 3430 9869 3431 9873
rect 3435 9869 3436 9873
rect 3440 9869 3441 9873
rect 3445 9869 3446 9873
rect 3450 9869 3451 9873
rect 3410 9868 3455 9869
rect 3410 9864 3411 9868
rect 3415 9864 3416 9868
rect 3420 9864 3421 9868
rect 3425 9864 3426 9868
rect 3430 9864 3431 9868
rect 3435 9864 3436 9868
rect 3440 9864 3441 9868
rect 3445 9864 3446 9868
rect 3450 9864 3451 9868
rect 3463 9948 3467 9949
rect 3463 9943 3467 9944
rect 3463 9938 3467 9939
rect 3463 9933 3467 9934
rect 3463 9928 3467 9929
rect 3463 9923 3467 9924
rect 3463 9918 3467 9919
rect 3463 9913 3467 9914
rect 3463 9908 3467 9909
rect 3463 9903 3467 9904
rect 3463 9898 3467 9899
rect 3463 9893 3467 9894
rect 3463 9888 3467 9889
rect 3463 9883 3467 9884
rect 3463 9878 3467 9879
rect 3463 9873 3467 9874
rect 3463 9868 3467 9869
rect 3399 9863 3403 9864
rect 3399 9856 3403 9859
rect 3463 9863 3467 9864
rect 3463 9856 3467 9859
rect 3403 9848 3406 9856
rect 3410 9848 3411 9856
rect 3415 9848 3416 9856
rect 3420 9848 3421 9856
rect 3425 9848 3426 9856
rect 3430 9848 3431 9856
rect 3435 9848 3436 9856
rect 3440 9848 3441 9856
rect 3445 9848 3446 9856
rect 3450 9848 3451 9856
rect 3455 9848 3456 9856
rect 3460 9848 3463 9856
rect 3476 9963 3480 9964
rect 3476 9958 3480 9959
rect 3476 9953 3480 9954
rect 3476 9948 3480 9949
rect 3476 9943 3480 9944
rect 3476 9938 3480 9939
rect 3476 9933 3480 9934
rect 3476 9928 3480 9929
rect 3476 9923 3480 9924
rect 3476 9918 3480 9919
rect 3476 9913 3480 9914
rect 3476 9908 3480 9909
rect 3476 9903 3480 9904
rect 3476 9898 3480 9899
rect 3476 9893 3480 9894
rect 3476 9888 3480 9889
rect 3476 9883 3480 9884
rect 3476 9878 3480 9879
rect 3476 9873 3480 9874
rect 3476 9868 3480 9869
rect 3476 9863 3480 9864
rect 3476 9858 3480 9859
rect 3476 9853 3480 9854
rect 3476 9848 3480 9849
rect 3386 9843 3390 9844
rect 3476 9843 3480 9844
rect 3390 9839 3391 9843
rect 3395 9839 3396 9843
rect 3400 9839 3401 9843
rect 3405 9839 3406 9843
rect 3410 9839 3411 9843
rect 3415 9839 3416 9843
rect 3420 9839 3421 9843
rect 3425 9839 3426 9843
rect 3430 9839 3431 9843
rect 3435 9839 3436 9843
rect 3440 9839 3441 9843
rect 3445 9839 3446 9843
rect 3450 9839 3451 9843
rect 3455 9839 3456 9843
rect 3460 9839 3461 9843
rect 3465 9839 3466 9843
rect 3470 9839 3471 9843
rect 3475 9839 3476 9843
rect 3539 9974 3540 9978
rect 3544 9974 3545 9978
rect 3549 9974 3550 9978
rect 3554 9974 3555 9978
rect 3559 9974 3560 9978
rect 3564 9974 3565 9978
rect 3569 9974 3570 9978
rect 3574 9974 3575 9978
rect 3579 9974 3580 9978
rect 3584 9974 3585 9978
rect 3589 9974 3590 9978
rect 3594 9974 3595 9978
rect 3599 9974 3600 9978
rect 3604 9974 3605 9978
rect 3609 9974 3610 9978
rect 3614 9974 3615 9978
rect 3619 9974 3620 9978
rect 3624 9974 3625 9978
rect 3535 9973 3539 9974
rect 3535 9968 3539 9969
rect 3625 9973 3629 9974
rect 3625 9968 3629 9969
rect 3535 9963 3539 9964
rect 3535 9958 3539 9959
rect 3535 9953 3539 9954
rect 3535 9948 3539 9949
rect 3535 9943 3539 9944
rect 3535 9938 3539 9939
rect 3535 9933 3539 9934
rect 3535 9928 3539 9929
rect 3535 9923 3539 9924
rect 3535 9918 3539 9919
rect 3535 9913 3539 9914
rect 3535 9908 3539 9909
rect 3535 9903 3539 9904
rect 3535 9898 3539 9899
rect 3535 9893 3539 9894
rect 3535 9888 3539 9889
rect 3535 9883 3539 9884
rect 3535 9878 3539 9879
rect 3535 9873 3539 9874
rect 3535 9868 3539 9869
rect 3535 9863 3539 9864
rect 3535 9858 3539 9859
rect 3535 9853 3539 9854
rect 3535 9848 3539 9849
rect 3552 9961 3555 9965
rect 3559 9961 3560 9965
rect 3564 9961 3565 9965
rect 3569 9961 3570 9965
rect 3574 9961 3575 9965
rect 3579 9961 3580 9965
rect 3584 9961 3585 9965
rect 3589 9961 3590 9965
rect 3594 9961 3595 9965
rect 3599 9961 3600 9965
rect 3604 9961 3605 9965
rect 3609 9961 3612 9965
rect 3548 9958 3552 9961
rect 3548 9953 3552 9954
rect 3612 9958 3616 9961
rect 3612 9953 3616 9954
rect 3548 9948 3552 9949
rect 3548 9943 3552 9944
rect 3548 9938 3552 9939
rect 3548 9933 3552 9934
rect 3548 9928 3552 9929
rect 3548 9923 3552 9924
rect 3548 9918 3552 9919
rect 3548 9913 3552 9914
rect 3548 9908 3552 9909
rect 3548 9903 3552 9904
rect 3548 9898 3552 9899
rect 3548 9893 3552 9894
rect 3548 9888 3552 9889
rect 3548 9883 3552 9884
rect 3548 9878 3552 9879
rect 3548 9873 3552 9874
rect 3548 9868 3552 9869
rect 3564 9949 3565 9953
rect 3569 9949 3570 9953
rect 3574 9949 3575 9953
rect 3579 9949 3580 9953
rect 3584 9949 3585 9953
rect 3589 9949 3590 9953
rect 3594 9949 3595 9953
rect 3599 9949 3600 9953
rect 3560 9948 3604 9949
rect 3564 9944 3565 9948
rect 3569 9944 3570 9948
rect 3574 9944 3575 9948
rect 3579 9944 3580 9948
rect 3584 9944 3585 9948
rect 3589 9944 3590 9948
rect 3594 9944 3595 9948
rect 3599 9944 3600 9948
rect 3560 9943 3604 9944
rect 3564 9939 3565 9943
rect 3569 9939 3570 9943
rect 3574 9939 3575 9943
rect 3579 9939 3580 9943
rect 3584 9939 3585 9943
rect 3589 9939 3590 9943
rect 3594 9939 3595 9943
rect 3599 9939 3600 9943
rect 3560 9938 3604 9939
rect 3564 9934 3565 9938
rect 3569 9934 3570 9938
rect 3574 9934 3575 9938
rect 3579 9934 3580 9938
rect 3584 9934 3585 9938
rect 3589 9934 3590 9938
rect 3594 9934 3595 9938
rect 3599 9934 3600 9938
rect 3560 9933 3604 9934
rect 3564 9929 3565 9933
rect 3569 9929 3570 9933
rect 3574 9929 3575 9933
rect 3579 9929 3580 9933
rect 3584 9929 3585 9933
rect 3589 9929 3590 9933
rect 3594 9929 3595 9933
rect 3599 9929 3600 9933
rect 3560 9928 3604 9929
rect 3564 9924 3565 9928
rect 3569 9924 3570 9928
rect 3574 9924 3575 9928
rect 3579 9924 3580 9928
rect 3584 9924 3585 9928
rect 3589 9924 3590 9928
rect 3594 9924 3595 9928
rect 3599 9924 3600 9928
rect 3560 9923 3604 9924
rect 3564 9919 3565 9923
rect 3569 9919 3570 9923
rect 3574 9919 3575 9923
rect 3579 9919 3580 9923
rect 3584 9919 3585 9923
rect 3589 9919 3590 9923
rect 3594 9919 3595 9923
rect 3599 9919 3600 9923
rect 3560 9918 3604 9919
rect 3564 9914 3565 9918
rect 3569 9914 3570 9918
rect 3574 9914 3575 9918
rect 3579 9914 3580 9918
rect 3584 9914 3585 9918
rect 3589 9914 3590 9918
rect 3594 9914 3595 9918
rect 3599 9914 3600 9918
rect 3560 9913 3604 9914
rect 3564 9909 3565 9913
rect 3569 9909 3570 9913
rect 3574 9909 3575 9913
rect 3579 9909 3580 9913
rect 3584 9909 3585 9913
rect 3589 9909 3590 9913
rect 3594 9909 3595 9913
rect 3599 9909 3600 9913
rect 3560 9908 3604 9909
rect 3564 9904 3565 9908
rect 3569 9904 3570 9908
rect 3574 9904 3575 9908
rect 3579 9904 3580 9908
rect 3584 9904 3585 9908
rect 3589 9904 3590 9908
rect 3594 9904 3595 9908
rect 3599 9904 3600 9908
rect 3560 9903 3604 9904
rect 3564 9899 3565 9903
rect 3569 9899 3570 9903
rect 3574 9899 3575 9903
rect 3579 9899 3580 9903
rect 3584 9899 3585 9903
rect 3589 9899 3590 9903
rect 3594 9899 3595 9903
rect 3599 9899 3600 9903
rect 3560 9898 3604 9899
rect 3564 9894 3565 9898
rect 3569 9894 3570 9898
rect 3574 9894 3575 9898
rect 3579 9894 3580 9898
rect 3584 9894 3585 9898
rect 3589 9894 3590 9898
rect 3594 9894 3595 9898
rect 3599 9894 3600 9898
rect 3560 9893 3604 9894
rect 3564 9889 3565 9893
rect 3569 9889 3570 9893
rect 3574 9889 3575 9893
rect 3579 9889 3580 9893
rect 3584 9889 3585 9893
rect 3589 9889 3590 9893
rect 3594 9889 3595 9893
rect 3599 9889 3600 9893
rect 3560 9888 3604 9889
rect 3564 9884 3565 9888
rect 3569 9884 3570 9888
rect 3574 9884 3575 9888
rect 3579 9884 3580 9888
rect 3584 9884 3585 9888
rect 3589 9884 3590 9888
rect 3594 9884 3595 9888
rect 3599 9884 3600 9888
rect 3560 9883 3604 9884
rect 3564 9879 3565 9883
rect 3569 9879 3570 9883
rect 3574 9879 3575 9883
rect 3579 9879 3580 9883
rect 3584 9879 3585 9883
rect 3589 9879 3590 9883
rect 3594 9879 3595 9883
rect 3599 9879 3600 9883
rect 3560 9878 3604 9879
rect 3564 9874 3565 9878
rect 3569 9874 3570 9878
rect 3574 9874 3575 9878
rect 3579 9874 3580 9878
rect 3584 9874 3585 9878
rect 3589 9874 3590 9878
rect 3594 9874 3595 9878
rect 3599 9874 3600 9878
rect 3560 9873 3604 9874
rect 3564 9869 3565 9873
rect 3569 9869 3570 9873
rect 3574 9869 3575 9873
rect 3579 9869 3580 9873
rect 3584 9869 3585 9873
rect 3589 9869 3590 9873
rect 3594 9869 3595 9873
rect 3599 9869 3600 9873
rect 3560 9868 3604 9869
rect 3564 9864 3565 9868
rect 3569 9864 3570 9868
rect 3574 9864 3575 9868
rect 3579 9864 3580 9868
rect 3584 9864 3585 9868
rect 3589 9864 3590 9868
rect 3594 9864 3595 9868
rect 3599 9864 3600 9868
rect 3612 9948 3616 9949
rect 3612 9943 3616 9944
rect 3612 9938 3616 9939
rect 3612 9933 3616 9934
rect 3612 9928 3616 9929
rect 3612 9923 3616 9924
rect 3612 9918 3616 9919
rect 3612 9913 3616 9914
rect 3612 9908 3616 9909
rect 3612 9903 3616 9904
rect 3612 9898 3616 9899
rect 3612 9893 3616 9894
rect 3612 9888 3616 9889
rect 3612 9883 3616 9884
rect 3612 9878 3616 9879
rect 3612 9873 3616 9874
rect 3612 9868 3616 9869
rect 3548 9863 3552 9864
rect 3548 9856 3552 9859
rect 3612 9863 3616 9864
rect 3612 9856 3616 9859
rect 3552 9848 3555 9856
rect 3559 9848 3560 9856
rect 3564 9848 3565 9856
rect 3569 9848 3570 9856
rect 3574 9848 3575 9856
rect 3579 9848 3580 9856
rect 3584 9848 3585 9856
rect 3589 9848 3590 9856
rect 3594 9848 3595 9856
rect 3599 9848 3600 9856
rect 3604 9848 3605 9856
rect 3609 9848 3612 9856
rect 3625 9963 3629 9964
rect 3625 9958 3629 9959
rect 3625 9953 3629 9954
rect 3625 9948 3629 9949
rect 3625 9943 3629 9944
rect 3625 9938 3629 9939
rect 3625 9933 3629 9934
rect 3625 9928 3629 9929
rect 3625 9923 3629 9924
rect 3625 9918 3629 9919
rect 3625 9913 3629 9914
rect 3625 9908 3629 9909
rect 3625 9903 3629 9904
rect 3625 9898 3629 9899
rect 3625 9893 3629 9894
rect 3625 9888 3629 9889
rect 3625 9883 3629 9884
rect 3625 9878 3629 9879
rect 3625 9873 3629 9874
rect 3625 9868 3629 9869
rect 3625 9863 3629 9864
rect 3625 9858 3629 9859
rect 3625 9853 3629 9854
rect 3625 9848 3629 9849
rect 3535 9843 3539 9844
rect 3625 9843 3629 9844
rect 3539 9839 3540 9843
rect 3544 9839 3545 9843
rect 3549 9839 3550 9843
rect 3554 9839 3555 9843
rect 3559 9839 3560 9843
rect 3564 9839 3565 9843
rect 3569 9839 3570 9843
rect 3574 9839 3575 9843
rect 3579 9839 3580 9843
rect 3584 9839 3585 9843
rect 3589 9839 3590 9843
rect 3594 9839 3595 9843
rect 3599 9839 3600 9843
rect 3604 9839 3605 9843
rect 3609 9839 3610 9843
rect 3614 9839 3615 9843
rect 3619 9839 3620 9843
rect 3624 9839 3625 9843
rect 3327 9711 3353 9715
rect 3357 9711 3358 9715
rect 3362 9711 3379 9715
rect 3423 9722 3479 9839
rect 3538 9802 3594 9839
rect 3526 9800 3594 9802
rect 3526 9796 3527 9800
rect 3531 9796 3532 9800
rect 3536 9796 3594 9800
rect 3526 9795 3594 9796
rect 3526 9791 3527 9795
rect 3531 9791 3532 9795
rect 3536 9791 3594 9795
rect 3526 9790 3594 9791
rect 3526 9786 3527 9790
rect 3531 9786 3532 9790
rect 3536 9786 3594 9790
rect 3526 9785 3594 9786
rect 3526 9781 3527 9785
rect 3531 9781 3532 9785
rect 3536 9781 3594 9785
rect 3526 9780 3594 9781
rect 3526 9776 3527 9780
rect 3531 9776 3532 9780
rect 3536 9776 3594 9780
rect 3526 9775 3594 9776
rect 3526 9771 3527 9775
rect 3531 9771 3532 9775
rect 3536 9771 3594 9775
rect 3526 9770 3594 9771
rect 3526 9766 3527 9770
rect 3531 9766 3532 9770
rect 3536 9766 3594 9770
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3482 9761 3501 9762
rect 3486 9757 3487 9761
rect 3491 9757 3492 9761
rect 3496 9757 3497 9761
rect 3482 9756 3501 9757
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3482 9751 3501 9752
rect 3486 9747 3487 9751
rect 3491 9747 3492 9751
rect 3496 9747 3497 9751
rect 3482 9746 3501 9747
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3482 9741 3501 9742
rect 3486 9737 3487 9741
rect 3491 9737 3492 9741
rect 3496 9737 3497 9741
rect 3482 9736 3501 9737
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3526 9765 3594 9766
rect 3526 9761 3527 9765
rect 3531 9761 3532 9765
rect 3536 9761 3594 9765
rect 3526 9760 3594 9761
rect 3526 9756 3527 9760
rect 3531 9756 3532 9760
rect 3536 9756 3594 9760
rect 3526 9755 3594 9756
rect 3526 9751 3527 9755
rect 3531 9751 3532 9755
rect 3536 9751 3594 9755
rect 3526 9750 3594 9751
rect 3526 9746 3527 9750
rect 3531 9746 3532 9750
rect 3536 9746 3594 9750
rect 3526 9745 3594 9746
rect 3526 9741 3527 9745
rect 3531 9741 3532 9745
rect 3536 9741 3594 9745
rect 3526 9740 3594 9741
rect 3526 9736 3527 9740
rect 3531 9736 3532 9740
rect 3536 9736 3594 9740
rect 3526 9734 3594 9736
rect 3634 9795 3688 9981
rect 3699 9974 3700 9978
rect 3704 9974 3705 9978
rect 3709 9974 3710 9978
rect 3714 9974 3715 9978
rect 3719 9974 3720 9978
rect 3724 9974 3725 9978
rect 3729 9974 3730 9978
rect 3734 9974 3735 9978
rect 3739 9974 3740 9978
rect 3744 9974 3745 9978
rect 3749 9974 3750 9978
rect 3754 9974 3755 9978
rect 3759 9974 3760 9978
rect 3764 9974 3765 9978
rect 3769 9974 3770 9978
rect 3774 9974 3775 9978
rect 3779 9974 3780 9978
rect 3784 9974 3785 9978
rect 3695 9973 3699 9974
rect 3695 9968 3699 9969
rect 3785 9973 3789 9974
rect 3785 9968 3789 9969
rect 3695 9963 3699 9964
rect 3695 9958 3699 9959
rect 3695 9953 3699 9954
rect 3695 9948 3699 9949
rect 3695 9943 3699 9944
rect 3695 9938 3699 9939
rect 3695 9933 3699 9934
rect 3695 9928 3699 9929
rect 3695 9923 3699 9924
rect 3695 9918 3699 9919
rect 3695 9913 3699 9914
rect 3695 9908 3699 9909
rect 3695 9903 3699 9904
rect 3695 9898 3699 9899
rect 3695 9893 3699 9894
rect 3695 9888 3699 9889
rect 3695 9883 3699 9884
rect 3695 9878 3699 9879
rect 3695 9873 3699 9874
rect 3695 9868 3699 9869
rect 3695 9863 3699 9864
rect 3695 9858 3699 9859
rect 3695 9853 3699 9854
rect 3695 9848 3699 9849
rect 3712 9961 3715 9965
rect 3719 9961 3720 9965
rect 3724 9961 3725 9965
rect 3729 9961 3730 9965
rect 3734 9961 3735 9965
rect 3739 9961 3740 9965
rect 3744 9961 3745 9965
rect 3749 9961 3750 9965
rect 3754 9961 3755 9965
rect 3759 9961 3760 9965
rect 3764 9961 3765 9965
rect 3769 9961 3772 9965
rect 3708 9958 3712 9961
rect 3708 9953 3712 9954
rect 3772 9958 3776 9961
rect 3772 9953 3776 9954
rect 3708 9948 3712 9949
rect 3708 9943 3712 9944
rect 3708 9938 3712 9939
rect 3708 9933 3712 9934
rect 3708 9928 3712 9929
rect 3708 9923 3712 9924
rect 3708 9918 3712 9919
rect 3708 9913 3712 9914
rect 3708 9908 3712 9909
rect 3708 9903 3712 9904
rect 3708 9898 3712 9899
rect 3708 9893 3712 9894
rect 3708 9888 3712 9889
rect 3708 9883 3712 9884
rect 3708 9878 3712 9879
rect 3708 9873 3712 9874
rect 3708 9868 3712 9869
rect 3719 9949 3720 9953
rect 3724 9949 3725 9953
rect 3729 9949 3730 9953
rect 3734 9949 3735 9953
rect 3739 9949 3740 9953
rect 3744 9949 3745 9953
rect 3749 9949 3750 9953
rect 3754 9949 3755 9953
rect 3759 9949 3760 9953
rect 3719 9948 3764 9949
rect 3719 9944 3720 9948
rect 3724 9944 3725 9948
rect 3729 9944 3730 9948
rect 3734 9944 3735 9948
rect 3739 9944 3740 9948
rect 3744 9944 3745 9948
rect 3749 9944 3750 9948
rect 3754 9944 3755 9948
rect 3759 9944 3760 9948
rect 3719 9943 3764 9944
rect 3719 9939 3720 9943
rect 3724 9939 3725 9943
rect 3729 9939 3730 9943
rect 3734 9939 3735 9943
rect 3739 9939 3740 9943
rect 3744 9939 3745 9943
rect 3749 9939 3750 9943
rect 3754 9939 3755 9943
rect 3759 9939 3760 9943
rect 3719 9938 3764 9939
rect 3719 9934 3720 9938
rect 3724 9934 3725 9938
rect 3729 9934 3730 9938
rect 3734 9934 3735 9938
rect 3739 9934 3740 9938
rect 3744 9934 3745 9938
rect 3749 9934 3750 9938
rect 3754 9934 3755 9938
rect 3759 9934 3760 9938
rect 3719 9933 3764 9934
rect 3719 9929 3720 9933
rect 3724 9929 3725 9933
rect 3729 9929 3730 9933
rect 3734 9929 3735 9933
rect 3739 9929 3740 9933
rect 3744 9929 3745 9933
rect 3749 9929 3750 9933
rect 3754 9929 3755 9933
rect 3759 9929 3760 9933
rect 3719 9928 3764 9929
rect 3719 9924 3720 9928
rect 3724 9924 3725 9928
rect 3729 9924 3730 9928
rect 3734 9924 3735 9928
rect 3739 9924 3740 9928
rect 3744 9924 3745 9928
rect 3749 9924 3750 9928
rect 3754 9924 3755 9928
rect 3759 9924 3760 9928
rect 3719 9923 3764 9924
rect 3719 9919 3720 9923
rect 3724 9919 3725 9923
rect 3729 9919 3730 9923
rect 3734 9919 3735 9923
rect 3739 9919 3740 9923
rect 3744 9919 3745 9923
rect 3749 9919 3750 9923
rect 3754 9919 3755 9923
rect 3759 9919 3760 9923
rect 3719 9918 3764 9919
rect 3719 9914 3720 9918
rect 3724 9914 3725 9918
rect 3729 9914 3730 9918
rect 3734 9914 3735 9918
rect 3739 9914 3740 9918
rect 3744 9914 3745 9918
rect 3749 9914 3750 9918
rect 3754 9914 3755 9918
rect 3759 9914 3760 9918
rect 3719 9913 3764 9914
rect 3719 9909 3720 9913
rect 3724 9909 3725 9913
rect 3729 9909 3730 9913
rect 3734 9909 3735 9913
rect 3739 9909 3740 9913
rect 3744 9909 3745 9913
rect 3749 9909 3750 9913
rect 3754 9909 3755 9913
rect 3759 9909 3760 9913
rect 3719 9908 3764 9909
rect 3719 9904 3720 9908
rect 3724 9904 3725 9908
rect 3729 9904 3730 9908
rect 3734 9904 3735 9908
rect 3739 9904 3740 9908
rect 3744 9904 3745 9908
rect 3749 9904 3750 9908
rect 3754 9904 3755 9908
rect 3759 9904 3760 9908
rect 3719 9903 3764 9904
rect 3719 9899 3720 9903
rect 3724 9899 3725 9903
rect 3729 9899 3730 9903
rect 3734 9899 3735 9903
rect 3739 9899 3740 9903
rect 3744 9899 3745 9903
rect 3749 9899 3750 9903
rect 3754 9899 3755 9903
rect 3759 9899 3760 9903
rect 3719 9898 3764 9899
rect 3719 9894 3720 9898
rect 3724 9894 3725 9898
rect 3729 9894 3730 9898
rect 3734 9894 3735 9898
rect 3739 9894 3740 9898
rect 3744 9894 3745 9898
rect 3749 9894 3750 9898
rect 3754 9894 3755 9898
rect 3759 9894 3760 9898
rect 3719 9893 3764 9894
rect 3719 9889 3720 9893
rect 3724 9889 3725 9893
rect 3729 9889 3730 9893
rect 3734 9889 3735 9893
rect 3739 9889 3740 9893
rect 3744 9889 3745 9893
rect 3749 9889 3750 9893
rect 3754 9889 3755 9893
rect 3759 9889 3760 9893
rect 3719 9888 3764 9889
rect 3719 9884 3720 9888
rect 3724 9884 3725 9888
rect 3729 9884 3730 9888
rect 3734 9884 3735 9888
rect 3739 9884 3740 9888
rect 3744 9884 3745 9888
rect 3749 9884 3750 9888
rect 3754 9884 3755 9888
rect 3759 9884 3760 9888
rect 3719 9883 3764 9884
rect 3719 9879 3720 9883
rect 3724 9879 3725 9883
rect 3729 9879 3730 9883
rect 3734 9879 3735 9883
rect 3739 9879 3740 9883
rect 3744 9879 3745 9883
rect 3749 9879 3750 9883
rect 3754 9879 3755 9883
rect 3759 9879 3760 9883
rect 3719 9878 3764 9879
rect 3719 9874 3720 9878
rect 3724 9874 3725 9878
rect 3729 9874 3730 9878
rect 3734 9874 3735 9878
rect 3739 9874 3740 9878
rect 3744 9874 3745 9878
rect 3749 9874 3750 9878
rect 3754 9874 3755 9878
rect 3759 9874 3760 9878
rect 3719 9873 3764 9874
rect 3719 9869 3720 9873
rect 3724 9869 3725 9873
rect 3729 9869 3730 9873
rect 3734 9869 3735 9873
rect 3739 9869 3740 9873
rect 3744 9869 3745 9873
rect 3749 9869 3750 9873
rect 3754 9869 3755 9873
rect 3759 9869 3760 9873
rect 3719 9868 3764 9869
rect 3719 9864 3720 9868
rect 3724 9864 3725 9868
rect 3729 9864 3730 9868
rect 3734 9864 3735 9868
rect 3739 9864 3740 9868
rect 3744 9864 3745 9868
rect 3749 9864 3750 9868
rect 3754 9864 3755 9868
rect 3759 9864 3760 9868
rect 3772 9948 3776 9949
rect 3772 9943 3776 9944
rect 3772 9938 3776 9939
rect 3772 9933 3776 9934
rect 3772 9928 3776 9929
rect 3772 9923 3776 9924
rect 3772 9918 3776 9919
rect 3772 9913 3776 9914
rect 3772 9908 3776 9909
rect 3772 9903 3776 9904
rect 3772 9898 3776 9899
rect 3772 9893 3776 9894
rect 3772 9888 3776 9889
rect 3772 9883 3776 9884
rect 3772 9878 3776 9879
rect 3772 9873 3776 9874
rect 3772 9868 3776 9869
rect 3708 9863 3712 9864
rect 3708 9856 3712 9859
rect 3772 9863 3776 9864
rect 3772 9856 3776 9859
rect 3712 9848 3715 9856
rect 3719 9848 3720 9856
rect 3724 9848 3725 9856
rect 3729 9848 3730 9856
rect 3734 9848 3735 9856
rect 3739 9848 3740 9856
rect 3744 9848 3745 9856
rect 3749 9848 3750 9856
rect 3754 9848 3755 9856
rect 3759 9848 3760 9856
rect 3764 9848 3765 9856
rect 3769 9848 3772 9856
rect 3785 9963 3789 9964
rect 3785 9958 3789 9959
rect 3785 9953 3789 9954
rect 3785 9948 3789 9949
rect 3785 9943 3789 9944
rect 3785 9938 3789 9939
rect 3785 9933 3789 9934
rect 3785 9928 3789 9929
rect 3785 9923 3789 9924
rect 3785 9918 3789 9919
rect 3785 9913 3789 9914
rect 3785 9908 3789 9909
rect 3785 9903 3789 9904
rect 3785 9898 3789 9899
rect 3785 9893 3789 9894
rect 3785 9888 3789 9889
rect 3785 9883 3789 9884
rect 3785 9878 3789 9879
rect 3785 9873 3789 9874
rect 3785 9868 3789 9869
rect 3785 9863 3789 9864
rect 3785 9858 3789 9859
rect 3785 9853 3789 9854
rect 3785 9848 3789 9849
rect 3695 9843 3699 9844
rect 3785 9843 3789 9844
rect 3699 9839 3700 9843
rect 3704 9839 3705 9843
rect 3709 9839 3710 9843
rect 3714 9839 3715 9843
rect 3719 9839 3720 9843
rect 3724 9839 3725 9843
rect 3729 9839 3730 9843
rect 3734 9839 3735 9843
rect 3739 9839 3740 9843
rect 3744 9839 3745 9843
rect 3749 9839 3750 9843
rect 3754 9839 3755 9843
rect 3759 9839 3760 9843
rect 3764 9839 3765 9843
rect 3769 9839 3770 9843
rect 3774 9839 3775 9843
rect 3779 9839 3780 9843
rect 3784 9839 3785 9843
rect 3848 9974 3849 9978
rect 3853 9974 3854 9978
rect 3858 9974 3859 9978
rect 3863 9974 3864 9978
rect 3868 9974 3869 9978
rect 3873 9974 3874 9978
rect 3878 9974 3879 9978
rect 3883 9974 3884 9978
rect 3888 9974 3889 9978
rect 3893 9974 3894 9978
rect 3898 9974 3899 9978
rect 3903 9974 3904 9978
rect 3908 9974 3909 9978
rect 3913 9974 3914 9978
rect 3918 9974 3919 9978
rect 3923 9974 3924 9978
rect 3928 9974 3929 9978
rect 3933 9974 3934 9978
rect 3844 9973 3848 9974
rect 3844 9968 3848 9969
rect 3934 9973 3938 9974
rect 3934 9968 3938 9969
rect 3844 9963 3848 9964
rect 3844 9958 3848 9959
rect 3844 9953 3848 9954
rect 3844 9948 3848 9949
rect 3844 9943 3848 9944
rect 3844 9938 3848 9939
rect 3844 9933 3848 9934
rect 3844 9928 3848 9929
rect 3844 9923 3848 9924
rect 3844 9918 3848 9919
rect 3844 9913 3848 9914
rect 3844 9908 3848 9909
rect 3844 9903 3848 9904
rect 3844 9898 3848 9899
rect 3844 9893 3848 9894
rect 3844 9888 3848 9889
rect 3844 9883 3848 9884
rect 3844 9878 3848 9879
rect 3844 9873 3848 9874
rect 3844 9868 3848 9869
rect 3844 9863 3848 9864
rect 3844 9858 3848 9859
rect 3844 9853 3848 9854
rect 3844 9848 3848 9849
rect 3861 9961 3864 9965
rect 3868 9961 3869 9965
rect 3873 9961 3874 9965
rect 3878 9961 3879 9965
rect 3883 9961 3884 9965
rect 3888 9961 3889 9965
rect 3893 9961 3894 9965
rect 3898 9961 3899 9965
rect 3903 9961 3904 9965
rect 3908 9961 3909 9965
rect 3913 9961 3914 9965
rect 3918 9961 3921 9965
rect 3857 9958 3861 9961
rect 3857 9953 3861 9954
rect 3921 9958 3925 9961
rect 3921 9953 3925 9954
rect 3857 9948 3861 9949
rect 3857 9943 3861 9944
rect 3857 9938 3861 9939
rect 3857 9933 3861 9934
rect 3857 9928 3861 9929
rect 3857 9923 3861 9924
rect 3857 9918 3861 9919
rect 3857 9913 3861 9914
rect 3857 9908 3861 9909
rect 3857 9903 3861 9904
rect 3857 9898 3861 9899
rect 3857 9893 3861 9894
rect 3857 9888 3861 9889
rect 3857 9883 3861 9884
rect 3857 9878 3861 9879
rect 3857 9873 3861 9874
rect 3857 9868 3861 9869
rect 3873 9949 3874 9953
rect 3878 9949 3879 9953
rect 3883 9949 3884 9953
rect 3888 9949 3889 9953
rect 3893 9949 3894 9953
rect 3898 9949 3899 9953
rect 3903 9949 3904 9953
rect 3908 9949 3909 9953
rect 3869 9948 3913 9949
rect 3873 9944 3874 9948
rect 3878 9944 3879 9948
rect 3883 9944 3884 9948
rect 3888 9944 3889 9948
rect 3893 9944 3894 9948
rect 3898 9944 3899 9948
rect 3903 9944 3904 9948
rect 3908 9944 3909 9948
rect 3869 9943 3913 9944
rect 3873 9939 3874 9943
rect 3878 9939 3879 9943
rect 3883 9939 3884 9943
rect 3888 9939 3889 9943
rect 3893 9939 3894 9943
rect 3898 9939 3899 9943
rect 3903 9939 3904 9943
rect 3908 9939 3909 9943
rect 3869 9938 3913 9939
rect 3873 9934 3874 9938
rect 3878 9934 3879 9938
rect 3883 9934 3884 9938
rect 3888 9934 3889 9938
rect 3893 9934 3894 9938
rect 3898 9934 3899 9938
rect 3903 9934 3904 9938
rect 3908 9934 3909 9938
rect 3869 9933 3913 9934
rect 3873 9929 3874 9933
rect 3878 9929 3879 9933
rect 3883 9929 3884 9933
rect 3888 9929 3889 9933
rect 3893 9929 3894 9933
rect 3898 9929 3899 9933
rect 3903 9929 3904 9933
rect 3908 9929 3909 9933
rect 3869 9928 3913 9929
rect 3873 9924 3874 9928
rect 3878 9924 3879 9928
rect 3883 9924 3884 9928
rect 3888 9924 3889 9928
rect 3893 9924 3894 9928
rect 3898 9924 3899 9928
rect 3903 9924 3904 9928
rect 3908 9924 3909 9928
rect 3869 9923 3913 9924
rect 3873 9919 3874 9923
rect 3878 9919 3879 9923
rect 3883 9919 3884 9923
rect 3888 9919 3889 9923
rect 3893 9919 3894 9923
rect 3898 9919 3899 9923
rect 3903 9919 3904 9923
rect 3908 9919 3909 9923
rect 3869 9918 3913 9919
rect 3873 9914 3874 9918
rect 3878 9914 3879 9918
rect 3883 9914 3884 9918
rect 3888 9914 3889 9918
rect 3893 9914 3894 9918
rect 3898 9914 3899 9918
rect 3903 9914 3904 9918
rect 3908 9914 3909 9918
rect 3869 9913 3913 9914
rect 3873 9909 3874 9913
rect 3878 9909 3879 9913
rect 3883 9909 3884 9913
rect 3888 9909 3889 9913
rect 3893 9909 3894 9913
rect 3898 9909 3899 9913
rect 3903 9909 3904 9913
rect 3908 9909 3909 9913
rect 3869 9908 3913 9909
rect 3873 9904 3874 9908
rect 3878 9904 3879 9908
rect 3883 9904 3884 9908
rect 3888 9904 3889 9908
rect 3893 9904 3894 9908
rect 3898 9904 3899 9908
rect 3903 9904 3904 9908
rect 3908 9904 3909 9908
rect 3869 9903 3913 9904
rect 3873 9899 3874 9903
rect 3878 9899 3879 9903
rect 3883 9899 3884 9903
rect 3888 9899 3889 9903
rect 3893 9899 3894 9903
rect 3898 9899 3899 9903
rect 3903 9899 3904 9903
rect 3908 9899 3909 9903
rect 3869 9898 3913 9899
rect 3873 9894 3874 9898
rect 3878 9894 3879 9898
rect 3883 9894 3884 9898
rect 3888 9894 3889 9898
rect 3893 9894 3894 9898
rect 3898 9894 3899 9898
rect 3903 9894 3904 9898
rect 3908 9894 3909 9898
rect 3869 9893 3913 9894
rect 3873 9889 3874 9893
rect 3878 9889 3879 9893
rect 3883 9889 3884 9893
rect 3888 9889 3889 9893
rect 3893 9889 3894 9893
rect 3898 9889 3899 9893
rect 3903 9889 3904 9893
rect 3908 9889 3909 9893
rect 3869 9888 3913 9889
rect 3873 9884 3874 9888
rect 3878 9884 3879 9888
rect 3883 9884 3884 9888
rect 3888 9884 3889 9888
rect 3893 9884 3894 9888
rect 3898 9884 3899 9888
rect 3903 9884 3904 9888
rect 3908 9884 3909 9888
rect 3869 9883 3913 9884
rect 3873 9879 3874 9883
rect 3878 9879 3879 9883
rect 3883 9879 3884 9883
rect 3888 9879 3889 9883
rect 3893 9879 3894 9883
rect 3898 9879 3899 9883
rect 3903 9879 3904 9883
rect 3908 9879 3909 9883
rect 3869 9878 3913 9879
rect 3873 9874 3874 9878
rect 3878 9874 3879 9878
rect 3883 9874 3884 9878
rect 3888 9874 3889 9878
rect 3893 9874 3894 9878
rect 3898 9874 3899 9878
rect 3903 9874 3904 9878
rect 3908 9874 3909 9878
rect 3869 9873 3913 9874
rect 3873 9869 3874 9873
rect 3878 9869 3879 9873
rect 3883 9869 3884 9873
rect 3888 9869 3889 9873
rect 3893 9869 3894 9873
rect 3898 9869 3899 9873
rect 3903 9869 3904 9873
rect 3908 9869 3909 9873
rect 3869 9868 3913 9869
rect 3873 9864 3874 9868
rect 3878 9864 3879 9868
rect 3883 9864 3884 9868
rect 3888 9864 3889 9868
rect 3893 9864 3894 9868
rect 3898 9864 3899 9868
rect 3903 9864 3904 9868
rect 3908 9864 3909 9868
rect 3921 9948 3925 9949
rect 3921 9943 3925 9944
rect 3921 9938 3925 9939
rect 3921 9933 3925 9934
rect 3921 9928 3925 9929
rect 3921 9923 3925 9924
rect 3921 9918 3925 9919
rect 3921 9913 3925 9914
rect 3921 9908 3925 9909
rect 3921 9903 3925 9904
rect 3921 9898 3925 9899
rect 3921 9893 3925 9894
rect 3921 9888 3925 9889
rect 3921 9883 3925 9884
rect 3921 9878 3925 9879
rect 3921 9873 3925 9874
rect 3921 9868 3925 9869
rect 3857 9863 3861 9864
rect 3857 9856 3861 9859
rect 3921 9863 3925 9864
rect 3921 9856 3925 9859
rect 3861 9848 3864 9856
rect 3868 9848 3869 9856
rect 3873 9848 3874 9856
rect 3878 9848 3879 9856
rect 3883 9848 3884 9856
rect 3888 9848 3889 9856
rect 3893 9848 3894 9856
rect 3898 9848 3899 9856
rect 3903 9848 3904 9856
rect 3908 9848 3909 9856
rect 3913 9848 3914 9856
rect 3918 9848 3921 9856
rect 3934 9963 3938 9964
rect 3934 9958 3938 9959
rect 3934 9953 3938 9954
rect 3960 9961 3981 9981
rect 4008 9974 4009 9978
rect 4013 9974 4014 9978
rect 4018 9974 4019 9978
rect 4023 9974 4024 9978
rect 4028 9974 4029 9978
rect 4033 9974 4034 9978
rect 4038 9974 4039 9978
rect 4043 9974 4044 9978
rect 4048 9974 4049 9978
rect 4053 9974 4054 9978
rect 4058 9974 4059 9978
rect 4063 9974 4064 9978
rect 4068 9974 4069 9978
rect 4073 9974 4074 9978
rect 4078 9974 4079 9978
rect 4083 9974 4084 9978
rect 4088 9974 4089 9978
rect 4093 9974 4094 9978
rect 4004 9973 4008 9974
rect 4004 9968 4008 9969
rect 4094 9973 4098 9974
rect 4094 9968 4098 9969
rect 4004 9963 4008 9964
rect 4004 9958 4008 9959
rect 4004 9953 4008 9954
rect 3934 9948 3938 9949
rect 3934 9943 3938 9944
rect 3934 9938 3938 9939
rect 3934 9933 3938 9934
rect 3934 9928 3938 9929
rect 3934 9923 3938 9924
rect 3934 9918 3938 9919
rect 3934 9913 3938 9914
rect 3934 9908 3938 9909
rect 3934 9903 3938 9904
rect 3934 9898 3938 9899
rect 3934 9893 3938 9894
rect 3934 9888 3938 9889
rect 3934 9883 3938 9884
rect 4004 9948 4008 9949
rect 4004 9943 4008 9944
rect 4004 9938 4008 9939
rect 4004 9933 4008 9934
rect 4004 9928 4008 9929
rect 4004 9923 4008 9924
rect 4004 9918 4008 9919
rect 4004 9913 4008 9914
rect 4004 9908 4008 9909
rect 4004 9903 4008 9904
rect 4004 9898 4008 9899
rect 4004 9893 4008 9894
rect 4004 9888 4008 9889
rect 4004 9883 4008 9884
rect 3934 9878 3938 9879
rect 3934 9873 3938 9874
rect 3934 9868 3938 9869
rect 3934 9863 3938 9864
rect 3934 9858 3938 9859
rect 3934 9853 3938 9854
rect 3934 9848 3938 9849
rect 3844 9843 3848 9844
rect 3960 9846 3981 9874
rect 4004 9878 4008 9879
rect 4004 9873 4008 9874
rect 4004 9868 4008 9869
rect 4004 9863 4008 9864
rect 4004 9858 4008 9859
rect 4004 9853 4008 9854
rect 4004 9848 4008 9849
rect 4021 9961 4024 9965
rect 4028 9961 4029 9965
rect 4033 9961 4034 9965
rect 4038 9961 4039 9965
rect 4043 9961 4044 9965
rect 4048 9961 4049 9965
rect 4053 9961 4054 9965
rect 4058 9961 4059 9965
rect 4063 9961 4064 9965
rect 4068 9961 4069 9965
rect 4073 9961 4074 9965
rect 4078 9961 4081 9965
rect 4017 9958 4021 9961
rect 4017 9953 4021 9954
rect 4081 9958 4085 9961
rect 4081 9953 4085 9954
rect 4017 9948 4021 9949
rect 4017 9943 4021 9944
rect 4017 9938 4021 9939
rect 4017 9933 4021 9934
rect 4017 9928 4021 9929
rect 4017 9923 4021 9924
rect 4017 9918 4021 9919
rect 4017 9913 4021 9914
rect 4017 9908 4021 9909
rect 4017 9903 4021 9904
rect 4017 9898 4021 9899
rect 4017 9893 4021 9894
rect 4017 9888 4021 9889
rect 4017 9883 4021 9884
rect 4017 9878 4021 9879
rect 4017 9873 4021 9874
rect 4017 9868 4021 9869
rect 4028 9949 4029 9953
rect 4033 9949 4034 9953
rect 4038 9949 4039 9953
rect 4043 9949 4044 9953
rect 4048 9949 4049 9953
rect 4053 9949 4054 9953
rect 4058 9949 4059 9953
rect 4063 9949 4064 9953
rect 4068 9949 4069 9953
rect 4028 9948 4073 9949
rect 4028 9944 4029 9948
rect 4033 9944 4034 9948
rect 4038 9944 4039 9948
rect 4043 9944 4044 9948
rect 4048 9944 4049 9948
rect 4053 9944 4054 9948
rect 4058 9944 4059 9948
rect 4063 9944 4064 9948
rect 4068 9944 4069 9948
rect 4028 9943 4073 9944
rect 4028 9939 4029 9943
rect 4033 9939 4034 9943
rect 4038 9939 4039 9943
rect 4043 9939 4044 9943
rect 4048 9939 4049 9943
rect 4053 9939 4054 9943
rect 4058 9939 4059 9943
rect 4063 9939 4064 9943
rect 4068 9939 4069 9943
rect 4028 9938 4073 9939
rect 4028 9934 4029 9938
rect 4033 9934 4034 9938
rect 4038 9934 4039 9938
rect 4043 9934 4044 9938
rect 4048 9934 4049 9938
rect 4053 9934 4054 9938
rect 4058 9934 4059 9938
rect 4063 9934 4064 9938
rect 4068 9934 4069 9938
rect 4028 9933 4073 9934
rect 4028 9929 4029 9933
rect 4033 9929 4034 9933
rect 4038 9929 4039 9933
rect 4043 9929 4044 9933
rect 4048 9929 4049 9933
rect 4053 9929 4054 9933
rect 4058 9929 4059 9933
rect 4063 9929 4064 9933
rect 4068 9929 4069 9933
rect 4028 9928 4073 9929
rect 4028 9924 4029 9928
rect 4033 9924 4034 9928
rect 4038 9924 4039 9928
rect 4043 9924 4044 9928
rect 4048 9924 4049 9928
rect 4053 9924 4054 9928
rect 4058 9924 4059 9928
rect 4063 9924 4064 9928
rect 4068 9924 4069 9928
rect 4028 9923 4073 9924
rect 4028 9919 4029 9923
rect 4033 9919 4034 9923
rect 4038 9919 4039 9923
rect 4043 9919 4044 9923
rect 4048 9919 4049 9923
rect 4053 9919 4054 9923
rect 4058 9919 4059 9923
rect 4063 9919 4064 9923
rect 4068 9919 4069 9923
rect 4028 9918 4073 9919
rect 4028 9914 4029 9918
rect 4033 9914 4034 9918
rect 4038 9914 4039 9918
rect 4043 9914 4044 9918
rect 4048 9914 4049 9918
rect 4053 9914 4054 9918
rect 4058 9914 4059 9918
rect 4063 9914 4064 9918
rect 4068 9914 4069 9918
rect 4028 9913 4073 9914
rect 4028 9909 4029 9913
rect 4033 9909 4034 9913
rect 4038 9909 4039 9913
rect 4043 9909 4044 9913
rect 4048 9909 4049 9913
rect 4053 9909 4054 9913
rect 4058 9909 4059 9913
rect 4063 9909 4064 9913
rect 4068 9909 4069 9913
rect 4028 9908 4073 9909
rect 4028 9904 4029 9908
rect 4033 9904 4034 9908
rect 4038 9904 4039 9908
rect 4043 9904 4044 9908
rect 4048 9904 4049 9908
rect 4053 9904 4054 9908
rect 4058 9904 4059 9908
rect 4063 9904 4064 9908
rect 4068 9904 4069 9908
rect 4028 9903 4073 9904
rect 4028 9899 4029 9903
rect 4033 9899 4034 9903
rect 4038 9899 4039 9903
rect 4043 9899 4044 9903
rect 4048 9899 4049 9903
rect 4053 9899 4054 9903
rect 4058 9899 4059 9903
rect 4063 9899 4064 9903
rect 4068 9899 4069 9903
rect 4028 9898 4073 9899
rect 4028 9894 4029 9898
rect 4033 9894 4034 9898
rect 4038 9894 4039 9898
rect 4043 9894 4044 9898
rect 4048 9894 4049 9898
rect 4053 9894 4054 9898
rect 4058 9894 4059 9898
rect 4063 9894 4064 9898
rect 4068 9894 4069 9898
rect 4028 9893 4073 9894
rect 4028 9889 4029 9893
rect 4033 9889 4034 9893
rect 4038 9889 4039 9893
rect 4043 9889 4044 9893
rect 4048 9889 4049 9893
rect 4053 9889 4054 9893
rect 4058 9889 4059 9893
rect 4063 9889 4064 9893
rect 4068 9889 4069 9893
rect 4028 9888 4073 9889
rect 4028 9884 4029 9888
rect 4033 9884 4034 9888
rect 4038 9884 4039 9888
rect 4043 9884 4044 9888
rect 4048 9884 4049 9888
rect 4053 9884 4054 9888
rect 4058 9884 4059 9888
rect 4063 9884 4064 9888
rect 4068 9884 4069 9888
rect 4028 9883 4073 9884
rect 4028 9879 4029 9883
rect 4033 9879 4034 9883
rect 4038 9879 4039 9883
rect 4043 9879 4044 9883
rect 4048 9879 4049 9883
rect 4053 9879 4054 9883
rect 4058 9879 4059 9883
rect 4063 9879 4064 9883
rect 4068 9879 4069 9883
rect 4028 9878 4073 9879
rect 4028 9874 4029 9878
rect 4033 9874 4034 9878
rect 4038 9874 4039 9878
rect 4043 9874 4044 9878
rect 4048 9874 4049 9878
rect 4053 9874 4054 9878
rect 4058 9874 4059 9878
rect 4063 9874 4064 9878
rect 4068 9874 4069 9878
rect 4028 9873 4073 9874
rect 4028 9869 4029 9873
rect 4033 9869 4034 9873
rect 4038 9869 4039 9873
rect 4043 9869 4044 9873
rect 4048 9869 4049 9873
rect 4053 9869 4054 9873
rect 4058 9869 4059 9873
rect 4063 9869 4064 9873
rect 4068 9869 4069 9873
rect 4028 9868 4073 9869
rect 4028 9864 4029 9868
rect 4033 9864 4034 9868
rect 4038 9864 4039 9868
rect 4043 9864 4044 9868
rect 4048 9864 4049 9868
rect 4053 9864 4054 9868
rect 4058 9864 4059 9868
rect 4063 9864 4064 9868
rect 4068 9864 4069 9868
rect 4081 9948 4085 9949
rect 4081 9943 4085 9944
rect 4081 9938 4085 9939
rect 4081 9933 4085 9934
rect 4081 9928 4085 9929
rect 4081 9923 4085 9924
rect 4081 9918 4085 9919
rect 4081 9913 4085 9914
rect 4081 9908 4085 9909
rect 4081 9903 4085 9904
rect 4081 9898 4085 9899
rect 4081 9893 4085 9894
rect 4081 9888 4085 9889
rect 4081 9883 4085 9884
rect 4081 9878 4085 9879
rect 4081 9873 4085 9874
rect 4081 9868 4085 9869
rect 4017 9863 4021 9864
rect 4017 9856 4021 9859
rect 4081 9863 4085 9864
rect 4081 9856 4085 9859
rect 4021 9848 4024 9856
rect 4028 9848 4029 9856
rect 4033 9848 4034 9856
rect 4038 9848 4039 9856
rect 4043 9848 4044 9856
rect 4048 9848 4049 9856
rect 4053 9848 4054 9856
rect 4058 9848 4059 9856
rect 4063 9848 4064 9856
rect 4068 9848 4069 9856
rect 4073 9848 4074 9856
rect 4078 9848 4081 9856
rect 4094 9963 4098 9964
rect 4094 9958 4098 9959
rect 4094 9953 4098 9954
rect 4094 9948 4098 9949
rect 4094 9943 4098 9944
rect 4094 9938 4098 9939
rect 4094 9933 4098 9934
rect 4094 9928 4098 9929
rect 4094 9923 4098 9924
rect 4094 9918 4098 9919
rect 4094 9913 4098 9914
rect 4094 9908 4098 9909
rect 4094 9903 4098 9904
rect 4094 9898 4098 9899
rect 4094 9893 4098 9894
rect 4094 9888 4098 9889
rect 4094 9883 4098 9884
rect 4094 9878 4098 9879
rect 4094 9873 4098 9874
rect 4094 9868 4098 9869
rect 4094 9863 4098 9864
rect 4094 9858 4098 9859
rect 4094 9853 4098 9854
rect 4094 9848 4098 9849
rect 3962 9844 3979 9846
rect 3934 9843 3938 9844
rect 3848 9839 3849 9843
rect 3853 9839 3854 9843
rect 3858 9839 3859 9843
rect 3863 9839 3864 9843
rect 3868 9839 3869 9843
rect 3873 9839 3874 9843
rect 3878 9839 3879 9843
rect 3883 9839 3884 9843
rect 3888 9839 3889 9843
rect 3893 9839 3894 9843
rect 3898 9839 3899 9843
rect 3903 9839 3904 9843
rect 3908 9839 3909 9843
rect 3913 9839 3914 9843
rect 3918 9839 3919 9843
rect 3923 9839 3924 9843
rect 3928 9839 3929 9843
rect 3933 9839 3934 9843
rect 3964 9842 3977 9844
rect 4004 9843 4008 9844
rect 4094 9843 4098 9844
rect 3634 9791 3662 9795
rect 3666 9791 3667 9795
rect 3671 9791 3688 9795
rect 3634 9790 3688 9791
rect 3634 9786 3662 9790
rect 3666 9786 3667 9790
rect 3671 9786 3688 9790
rect 3634 9785 3688 9786
rect 3634 9781 3662 9785
rect 3666 9781 3667 9785
rect 3671 9781 3688 9785
rect 3634 9780 3688 9781
rect 3634 9776 3662 9780
rect 3666 9776 3667 9780
rect 3671 9776 3688 9780
rect 3634 9775 3688 9776
rect 3634 9771 3662 9775
rect 3666 9771 3667 9775
rect 3671 9771 3688 9775
rect 3634 9770 3688 9771
rect 3634 9766 3662 9770
rect 3666 9766 3667 9770
rect 3671 9766 3688 9770
rect 3634 9765 3688 9766
rect 3634 9761 3662 9765
rect 3666 9761 3667 9765
rect 3671 9761 3688 9765
rect 3634 9760 3688 9761
rect 3634 9756 3662 9760
rect 3666 9756 3667 9760
rect 3671 9756 3688 9760
rect 3634 9755 3688 9756
rect 3634 9751 3662 9755
rect 3666 9751 3667 9755
rect 3671 9751 3688 9755
rect 3634 9750 3688 9751
rect 3634 9746 3662 9750
rect 3666 9746 3667 9750
rect 3671 9746 3688 9750
rect 3634 9745 3688 9746
rect 3634 9741 3662 9745
rect 3666 9741 3667 9745
rect 3671 9741 3688 9745
rect 3427 9718 3428 9722
rect 3432 9718 3433 9722
rect 3437 9718 3438 9722
rect 3442 9718 3443 9722
rect 3447 9718 3448 9722
rect 3452 9718 3453 9722
rect 3457 9718 3458 9722
rect 3462 9718 3463 9722
rect 3467 9718 3468 9722
rect 3472 9718 3473 9722
rect 3477 9718 3479 9722
rect 3423 9717 3479 9718
rect 3427 9713 3428 9717
rect 3432 9713 3433 9717
rect 3437 9713 3438 9717
rect 3442 9713 3443 9717
rect 3447 9713 3448 9717
rect 3452 9713 3453 9717
rect 3457 9713 3458 9717
rect 3462 9713 3463 9717
rect 3467 9713 3468 9717
rect 3472 9713 3473 9717
rect 3477 9713 3479 9717
rect 3423 9712 3479 9713
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3482 9715 3501 9716
rect 3327 9710 3379 9711
rect 3327 9706 3353 9710
rect 3357 9706 3358 9710
rect 3362 9706 3379 9710
rect 3327 9705 3379 9706
rect 3327 9701 3353 9705
rect 3357 9701 3358 9705
rect 3362 9701 3379 9705
rect 3327 9700 3379 9701
rect 3327 9696 3353 9700
rect 3357 9696 3358 9700
rect 3362 9696 3379 9700
rect 3327 9695 3379 9696
rect 3327 9691 3353 9695
rect 3357 9691 3358 9695
rect 3362 9691 3379 9695
rect 3327 9690 3379 9691
rect 3327 9686 3353 9690
rect 3357 9686 3358 9690
rect 3362 9686 3379 9690
rect 3486 9711 3487 9715
rect 3491 9711 3492 9715
rect 3496 9711 3497 9715
rect 3482 9710 3501 9711
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3482 9705 3501 9706
rect 3486 9701 3487 9705
rect 3491 9701 3492 9705
rect 3496 9701 3497 9705
rect 3482 9700 3501 9701
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3482 9695 3501 9696
rect 3486 9691 3487 9695
rect 3491 9691 3492 9695
rect 3496 9691 3497 9695
rect 3482 9690 3501 9691
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 2731 9605 3021 9609
rect 3327 9685 3379 9686
rect 3327 9681 3353 9685
rect 3357 9681 3358 9685
rect 3362 9681 3379 9685
rect 3327 9680 3379 9681
rect 3327 9676 3353 9680
rect 3357 9676 3358 9680
rect 3362 9676 3379 9680
rect 3327 9675 3379 9676
rect 3327 9671 3353 9675
rect 3357 9671 3358 9675
rect 3362 9671 3379 9675
rect 3327 9670 3379 9671
rect 3327 9666 3353 9670
rect 3357 9666 3358 9670
rect 3362 9666 3379 9670
rect 3327 9665 3379 9666
rect 3327 9661 3353 9665
rect 3357 9661 3358 9665
rect 3362 9661 3379 9665
rect 3327 9610 3379 9661
rect 3634 9629 3688 9741
rect 3732 9722 3788 9839
rect 3847 9831 3903 9839
rect 3966 9831 3975 9842
rect 4008 9839 4009 9843
rect 4013 9839 4014 9843
rect 4018 9839 4019 9843
rect 4023 9839 4024 9843
rect 4028 9839 4029 9843
rect 4033 9839 4034 9843
rect 4038 9839 4039 9843
rect 4043 9839 4044 9843
rect 4048 9839 4049 9843
rect 4053 9839 4054 9843
rect 4058 9839 4059 9843
rect 4063 9839 4064 9843
rect 4068 9839 4069 9843
rect 4073 9839 4074 9843
rect 4078 9839 4079 9843
rect 4083 9839 4084 9843
rect 4088 9839 4089 9843
rect 4093 9839 4094 9843
rect 4041 9831 4097 9839
rect 3847 9827 3906 9831
rect 4032 9827 4097 9831
rect 3847 9815 3903 9827
rect 3962 9819 3992 9823
rect 3847 9811 3906 9815
rect 3976 9812 3980 9819
rect 4041 9815 4097 9827
rect 3847 9802 3903 9811
rect 4032 9811 4097 9815
rect 3962 9803 3973 9807
rect 3835 9800 3903 9802
rect 3835 9796 3836 9800
rect 3840 9796 3841 9800
rect 3845 9799 3903 9800
rect 3966 9800 3973 9803
rect 3985 9803 3992 9807
rect 3985 9800 3989 9803
rect 3845 9796 3906 9799
rect 3835 9795 3906 9796
rect 3835 9791 3836 9795
rect 3840 9791 3841 9795
rect 3845 9791 3903 9795
rect 3966 9791 3989 9800
rect 4041 9799 4097 9811
rect 4032 9795 4097 9799
rect 3835 9790 3903 9791
rect 3835 9786 3836 9790
rect 3840 9786 3841 9790
rect 3845 9786 3903 9790
rect 3962 9787 3992 9791
rect 3835 9785 3903 9786
rect 3835 9781 3836 9785
rect 3840 9781 3841 9785
rect 3845 9783 3903 9785
rect 3845 9781 3906 9783
rect 3835 9780 3906 9781
rect 3835 9776 3836 9780
rect 3840 9776 3841 9780
rect 3845 9779 3906 9780
rect 3845 9776 3903 9779
rect 3835 9775 3903 9776
rect 3835 9771 3836 9775
rect 3840 9771 3841 9775
rect 3845 9771 3903 9775
rect 3835 9770 3903 9771
rect 3835 9766 3836 9770
rect 3840 9766 3841 9770
rect 3845 9766 3903 9770
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3791 9761 3810 9762
rect 3795 9757 3796 9761
rect 3800 9757 3801 9761
rect 3805 9757 3806 9761
rect 3791 9756 3810 9757
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3791 9751 3810 9752
rect 3795 9747 3796 9751
rect 3800 9747 3801 9751
rect 3805 9747 3806 9751
rect 3791 9746 3810 9747
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3791 9741 3810 9742
rect 3795 9737 3796 9741
rect 3800 9737 3801 9741
rect 3805 9737 3806 9741
rect 3791 9736 3810 9737
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3835 9765 3903 9766
rect 3835 9761 3836 9765
rect 3840 9761 3841 9765
rect 3845 9761 3903 9765
rect 3835 9760 3903 9761
rect 3835 9756 3836 9760
rect 3840 9756 3841 9760
rect 3845 9756 3903 9760
rect 3835 9755 3903 9756
rect 3835 9751 3836 9755
rect 3840 9751 3841 9755
rect 3845 9751 3903 9755
rect 3835 9750 3903 9751
rect 3835 9746 3836 9750
rect 3840 9746 3841 9750
rect 3845 9746 3903 9750
rect 3835 9745 3903 9746
rect 3835 9741 3836 9745
rect 3840 9741 3841 9745
rect 3845 9741 3903 9745
rect 3835 9740 3903 9741
rect 3835 9736 3836 9740
rect 3840 9736 3841 9740
rect 3845 9736 3903 9740
rect 3835 9734 3903 9736
rect 3736 9718 3737 9722
rect 3741 9718 3742 9722
rect 3746 9718 3747 9722
rect 3751 9718 3752 9722
rect 3756 9718 3757 9722
rect 3761 9718 3762 9722
rect 3766 9718 3767 9722
rect 3771 9718 3772 9722
rect 3776 9718 3777 9722
rect 3781 9718 3782 9722
rect 3786 9718 3788 9722
rect 3732 9717 3788 9718
rect 3736 9713 3737 9717
rect 3741 9713 3742 9717
rect 3746 9713 3747 9717
rect 3751 9713 3752 9717
rect 3756 9713 3757 9717
rect 3761 9713 3762 9717
rect 3766 9713 3767 9717
rect 3771 9713 3772 9717
rect 3776 9713 3777 9717
rect 3781 9713 3782 9717
rect 3786 9713 3788 9717
rect 3732 9712 3788 9713
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3791 9715 3810 9716
rect 3795 9711 3796 9715
rect 3800 9711 3801 9715
rect 3805 9711 3806 9715
rect 3791 9710 3810 9711
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3791 9705 3810 9706
rect 3795 9701 3796 9705
rect 3800 9701 3801 9705
rect 3805 9701 3806 9705
rect 3791 9700 3810 9701
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3791 9695 3810 9696
rect 3795 9691 3796 9695
rect 3800 9691 3801 9695
rect 3805 9691 3806 9695
rect 3791 9690 3810 9691
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 3634 9609 3690 9629
rect 2731 9604 2997 9605
rect 659 9591 693 9592
rect 663 9587 664 9591
rect 668 9587 669 9591
rect 673 9587 674 9591
rect 678 9587 679 9591
rect 683 9587 684 9591
rect 688 9587 689 9591
rect 659 9586 693 9587
rect 663 9582 664 9586
rect 668 9582 669 9586
rect 673 9582 674 9586
rect 678 9582 679 9586
rect 683 9582 684 9586
rect 688 9582 689 9586
rect 659 9581 693 9582
rect 663 9577 664 9581
rect 668 9577 669 9581
rect 673 9577 674 9581
rect 678 9577 679 9581
rect 683 9577 684 9581
rect 688 9577 689 9581
rect 2435 9575 2497 9597
rect 3967 9574 3980 9787
rect 4041 9783 4097 9795
rect 4141 9786 5073 10261
rect 4032 9779 4097 9783
rect 4041 9722 4097 9779
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4100 9761 4119 9762
rect 4104 9757 4105 9761
rect 4109 9757 4110 9761
rect 4114 9757 4115 9761
rect 4100 9756 4119 9757
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4100 9751 4119 9752
rect 4104 9747 4105 9751
rect 4109 9747 4110 9751
rect 4114 9747 4115 9751
rect 4100 9746 4119 9747
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4100 9741 4119 9742
rect 4104 9737 4105 9741
rect 4109 9737 4110 9741
rect 4114 9737 4115 9741
rect 4100 9736 4119 9737
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4292 9761 4311 9762
rect 4296 9757 4297 9761
rect 4301 9757 4302 9761
rect 4306 9757 4307 9761
rect 4292 9756 4311 9757
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4292 9751 4311 9752
rect 4296 9747 4297 9751
rect 4301 9747 4302 9751
rect 4306 9747 4307 9751
rect 4292 9746 4311 9747
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4292 9741 4311 9742
rect 4296 9737 4297 9741
rect 4301 9737 4302 9741
rect 4306 9737 4307 9741
rect 4292 9736 4311 9737
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4318 9761 4337 9762
rect 4322 9757 4323 9761
rect 4327 9757 4328 9761
rect 4332 9757 4333 9761
rect 4318 9756 4337 9757
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4318 9751 4337 9752
rect 4322 9747 4323 9751
rect 4327 9747 4328 9751
rect 4332 9747 4333 9751
rect 4318 9746 4337 9747
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4318 9741 4337 9742
rect 4322 9737 4323 9741
rect 4327 9737 4328 9741
rect 4332 9737 4333 9741
rect 4318 9736 4337 9737
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4344 9761 4363 9762
rect 4348 9757 4349 9761
rect 4353 9757 4354 9761
rect 4358 9757 4359 9761
rect 4344 9756 4363 9757
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4344 9751 4363 9752
rect 4348 9747 4349 9751
rect 4353 9747 4354 9751
rect 4358 9747 4359 9751
rect 4344 9746 4363 9747
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4344 9741 4363 9742
rect 4348 9737 4349 9741
rect 4353 9737 4354 9741
rect 4358 9737 4359 9741
rect 4344 9736 4363 9737
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4370 9761 4389 9762
rect 4374 9757 4375 9761
rect 4379 9757 4380 9761
rect 4384 9757 4385 9761
rect 4370 9756 4389 9757
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4370 9751 4389 9752
rect 4374 9747 4375 9751
rect 4379 9747 4380 9751
rect 4384 9747 4385 9751
rect 4370 9746 4389 9747
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4370 9741 4389 9742
rect 4374 9737 4375 9741
rect 4379 9737 4380 9741
rect 4384 9737 4385 9741
rect 4370 9736 4389 9737
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4396 9761 4415 9762
rect 4400 9757 4401 9761
rect 4405 9757 4406 9761
rect 4410 9757 4411 9761
rect 4396 9756 4415 9757
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4396 9751 4415 9752
rect 4400 9747 4401 9751
rect 4405 9747 4406 9751
rect 4410 9747 4411 9751
rect 4396 9746 4415 9747
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4396 9741 4415 9742
rect 4400 9737 4401 9741
rect 4405 9737 4406 9741
rect 4410 9737 4411 9741
rect 4396 9736 4415 9737
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 4045 9718 4046 9722
rect 4050 9718 4051 9722
rect 4055 9718 4056 9722
rect 4060 9718 4061 9722
rect 4065 9718 4066 9722
rect 4070 9718 4071 9722
rect 4075 9718 4076 9722
rect 4080 9718 4081 9722
rect 4085 9718 4086 9722
rect 4090 9718 4091 9722
rect 4095 9718 4097 9722
rect 4041 9717 4097 9718
rect 4045 9713 4046 9717
rect 4050 9713 4051 9717
rect 4055 9713 4056 9717
rect 4060 9713 4061 9717
rect 4065 9713 4066 9717
rect 4070 9713 4071 9717
rect 4075 9713 4076 9717
rect 4080 9713 4081 9717
rect 4085 9713 4086 9717
rect 4090 9713 4091 9717
rect 4095 9713 4097 9717
rect 4041 9712 4097 9713
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4100 9715 4119 9716
rect 4104 9711 4105 9715
rect 4109 9711 4110 9715
rect 4114 9711 4115 9715
rect 4100 9710 4119 9711
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4100 9705 4119 9706
rect 4104 9701 4105 9705
rect 4109 9701 4110 9705
rect 4114 9701 4115 9705
rect 4100 9700 4119 9701
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4100 9695 4119 9696
rect 4104 9691 4105 9695
rect 4109 9691 4110 9695
rect 4114 9691 4115 9695
rect 4100 9690 4119 9691
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4292 9715 4311 9716
rect 4296 9711 4297 9715
rect 4301 9711 4302 9715
rect 4306 9711 4307 9715
rect 4292 9710 4311 9711
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4292 9705 4311 9706
rect 4296 9701 4297 9705
rect 4301 9701 4302 9705
rect 4306 9701 4307 9705
rect 4292 9700 4311 9701
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4292 9695 4311 9696
rect 4296 9691 4297 9695
rect 4301 9691 4302 9695
rect 4306 9691 4307 9695
rect 4292 9690 4311 9691
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4318 9715 4337 9716
rect 4322 9711 4323 9715
rect 4327 9711 4328 9715
rect 4332 9711 4333 9715
rect 4318 9710 4337 9711
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4318 9705 4337 9706
rect 4322 9701 4323 9705
rect 4327 9701 4328 9705
rect 4332 9701 4333 9705
rect 4318 9700 4337 9701
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4318 9695 4337 9696
rect 4322 9691 4323 9695
rect 4327 9691 4328 9695
rect 4332 9691 4333 9695
rect 4318 9690 4337 9691
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4344 9715 4363 9716
rect 4348 9711 4349 9715
rect 4353 9711 4354 9715
rect 4358 9711 4359 9715
rect 4344 9710 4363 9711
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4344 9705 4363 9706
rect 4348 9701 4349 9705
rect 4353 9701 4354 9705
rect 4358 9701 4359 9705
rect 4344 9700 4363 9701
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4344 9695 4363 9696
rect 4348 9691 4349 9695
rect 4353 9691 4354 9695
rect 4358 9691 4359 9695
rect 4344 9690 4363 9691
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4370 9715 4389 9716
rect 4374 9711 4375 9715
rect 4379 9711 4380 9715
rect 4384 9711 4385 9715
rect 4370 9710 4389 9711
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4370 9705 4389 9706
rect 4374 9701 4375 9705
rect 4379 9701 4380 9705
rect 4384 9701 4385 9705
rect 4370 9700 4389 9701
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4370 9695 4389 9696
rect 4374 9691 4375 9695
rect 4379 9691 4380 9695
rect 4384 9691 4385 9695
rect 4370 9690 4389 9691
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4396 9715 4415 9716
rect 4400 9711 4401 9715
rect 4405 9711 4406 9715
rect 4410 9711 4411 9715
rect 4396 9710 4415 9711
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4396 9705 4415 9706
rect 4400 9701 4401 9705
rect 4405 9701 4406 9705
rect 4410 9701 4411 9705
rect 4396 9700 4415 9701
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4396 9695 4415 9696
rect 4400 9691 4401 9695
rect 4405 9691 4406 9695
rect 4410 9691 4411 9695
rect 4396 9690 4415 9691
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 617 9566 618 9570
rect 622 9566 623 9570
rect 627 9566 628 9570
rect 632 9566 633 9570
rect 637 9566 638 9570
rect 642 9566 643 9570
rect 613 9565 647 9566
rect 617 9561 618 9565
rect 622 9561 623 9565
rect 627 9561 628 9565
rect 632 9561 633 9565
rect 637 9561 638 9565
rect 642 9561 643 9565
rect 613 9560 647 9561
rect 617 9556 618 9560
rect 622 9556 623 9560
rect 627 9556 628 9560
rect 632 9556 633 9560
rect 637 9556 638 9560
rect 642 9556 643 9560
rect 613 9555 647 9556
rect 617 9551 618 9555
rect 622 9551 623 9555
rect 627 9551 628 9555
rect 632 9551 633 9555
rect 637 9551 638 9555
rect 642 9551 643 9555
rect 663 9566 664 9570
rect 668 9566 669 9570
rect 673 9566 674 9570
rect 678 9566 679 9570
rect 683 9566 684 9570
rect 688 9566 689 9570
rect 659 9565 693 9566
rect 663 9561 664 9565
rect 668 9561 669 9565
rect 673 9561 674 9565
rect 678 9561 679 9565
rect 683 9561 684 9565
rect 688 9561 689 9565
rect 659 9560 693 9561
rect 663 9556 664 9560
rect 668 9556 669 9560
rect 673 9556 674 9560
rect 678 9556 679 9560
rect 683 9556 684 9560
rect 688 9556 689 9560
rect 659 9555 693 9556
rect 663 9551 664 9555
rect 668 9551 669 9555
rect 673 9551 674 9555
rect 678 9551 679 9555
rect 683 9551 684 9555
rect 688 9551 689 9555
rect 2134 9549 2401 9571
rect 2414 9549 2476 9571
rect 2134 9547 2416 9549
rect 617 9540 618 9544
rect 622 9540 623 9544
rect 627 9540 628 9544
rect 632 9540 633 9544
rect 637 9540 638 9544
rect 642 9540 643 9544
rect 613 9539 647 9540
rect 617 9535 618 9539
rect 622 9535 623 9539
rect 627 9535 628 9539
rect 632 9535 633 9539
rect 637 9535 638 9539
rect 642 9535 643 9539
rect 613 9534 647 9535
rect 617 9530 618 9534
rect 622 9530 623 9534
rect 627 9530 628 9534
rect 632 9530 633 9534
rect 637 9530 638 9534
rect 642 9530 643 9534
rect 613 9529 647 9530
rect 617 9525 618 9529
rect 622 9525 623 9529
rect 627 9525 628 9529
rect 632 9525 633 9529
rect 637 9525 638 9529
rect 642 9525 643 9529
rect 663 9540 664 9544
rect 668 9540 669 9544
rect 673 9540 674 9544
rect 678 9540 679 9544
rect 683 9540 684 9544
rect 688 9540 689 9544
rect 659 9539 693 9540
rect 663 9535 664 9539
rect 668 9535 669 9539
rect 673 9535 674 9539
rect 678 9535 679 9539
rect 683 9535 684 9539
rect 688 9535 689 9539
rect 659 9534 693 9535
rect 663 9530 664 9534
rect 668 9530 669 9534
rect 673 9530 674 9534
rect 678 9530 679 9534
rect 683 9530 684 9534
rect 688 9530 689 9534
rect 659 9529 693 9530
rect 663 9525 664 9529
rect 668 9525 669 9529
rect 673 9525 674 9529
rect 678 9525 679 9529
rect 683 9525 684 9529
rect 688 9525 689 9529
rect 617 9514 618 9518
rect 622 9514 623 9518
rect 627 9514 628 9518
rect 632 9514 633 9518
rect 637 9514 638 9518
rect 642 9514 643 9518
rect 613 9513 647 9514
rect 617 9509 618 9513
rect 622 9509 623 9513
rect 627 9509 628 9513
rect 632 9509 633 9513
rect 637 9509 638 9513
rect 642 9509 643 9513
rect 613 9508 647 9509
rect 617 9504 618 9508
rect 622 9504 623 9508
rect 627 9504 628 9508
rect 632 9504 633 9508
rect 637 9504 638 9508
rect 642 9504 643 9508
rect 613 9503 647 9504
rect 617 9499 618 9503
rect 622 9499 623 9503
rect 627 9499 628 9503
rect 632 9499 633 9503
rect 637 9499 638 9503
rect 642 9499 643 9503
rect 663 9514 664 9518
rect 668 9514 669 9518
rect 673 9514 674 9518
rect 678 9514 679 9518
rect 683 9514 684 9518
rect 688 9514 689 9518
rect 659 9513 693 9514
rect 663 9509 664 9513
rect 668 9509 669 9513
rect 673 9509 674 9513
rect 678 9509 679 9513
rect 683 9509 684 9513
rect 688 9509 689 9513
rect 659 9508 693 9509
rect 663 9504 664 9508
rect 668 9504 669 9508
rect 673 9504 674 9508
rect 678 9504 679 9508
rect 683 9504 684 9508
rect 688 9504 689 9508
rect 659 9503 693 9504
rect 663 9499 664 9503
rect 668 9499 669 9503
rect 673 9499 674 9503
rect 678 9499 679 9503
rect 683 9499 684 9503
rect 688 9499 689 9503
rect 2830 9497 3769 9501
rect 2818 9489 3757 9493
rect 2806 9482 3745 9486
rect 2794 9475 3733 9479
rect 2782 9467 3327 9471
rect 3382 9467 3721 9471
rect 3727 9467 3788 9471
rect 3692 9463 3709 9464
rect 2770 9459 3635 9463
rect 3690 9460 3709 9463
rect 3715 9460 3788 9464
rect 3690 9459 3698 9460
rect 3968 9456 3980 9574
rect 4483 9573 4484 9577
rect 4488 9573 4489 9577
rect 4493 9573 4494 9577
rect 4498 9573 4499 9577
rect 4503 9573 4504 9577
rect 4508 9573 4509 9577
rect 4479 9572 4513 9573
rect 4483 9568 4484 9572
rect 4488 9568 4489 9572
rect 4493 9568 4494 9572
rect 4498 9568 4499 9572
rect 4503 9568 4504 9572
rect 4508 9568 4509 9572
rect 4479 9567 4513 9568
rect 4483 9563 4484 9567
rect 4488 9563 4489 9567
rect 4493 9563 4494 9567
rect 4498 9563 4499 9567
rect 4503 9563 4504 9567
rect 4508 9563 4509 9567
rect 4479 9562 4513 9563
rect 4483 9558 4484 9562
rect 4488 9558 4489 9562
rect 4493 9558 4494 9562
rect 4498 9558 4499 9562
rect 4503 9558 4504 9562
rect 4508 9558 4509 9562
rect 4529 9573 4530 9577
rect 4534 9573 4535 9577
rect 4539 9573 4540 9577
rect 4544 9573 4545 9577
rect 4549 9573 4550 9577
rect 4554 9573 4555 9577
rect 4525 9572 4559 9573
rect 4529 9568 4530 9572
rect 4534 9568 4535 9572
rect 4539 9568 4540 9572
rect 4544 9568 4545 9572
rect 4549 9568 4550 9572
rect 4554 9568 4555 9572
rect 4525 9567 4559 9568
rect 4529 9563 4530 9567
rect 4534 9563 4535 9567
rect 4539 9563 4540 9567
rect 4544 9563 4545 9567
rect 4549 9563 4550 9567
rect 4554 9563 4555 9567
rect 4525 9562 4559 9563
rect 4529 9558 4530 9562
rect 4534 9558 4535 9562
rect 4539 9558 4540 9562
rect 4544 9558 4545 9562
rect 4549 9558 4550 9562
rect 4554 9558 4555 9562
rect 4483 9544 4484 9548
rect 4488 9544 4489 9548
rect 4493 9544 4494 9548
rect 4498 9544 4499 9548
rect 4503 9544 4504 9548
rect 4508 9544 4509 9548
rect 4479 9543 4513 9544
rect 4483 9539 4484 9543
rect 4488 9539 4489 9543
rect 4493 9539 4494 9543
rect 4498 9539 4499 9543
rect 4503 9539 4504 9543
rect 4508 9539 4509 9543
rect 4479 9538 4513 9539
rect 4483 9534 4484 9538
rect 4488 9534 4489 9538
rect 4493 9534 4494 9538
rect 4498 9534 4499 9538
rect 4503 9534 4504 9538
rect 4508 9534 4509 9538
rect 4479 9533 4513 9534
rect 4483 9529 4484 9533
rect 4488 9529 4489 9533
rect 4493 9529 4494 9533
rect 4498 9529 4499 9533
rect 4503 9529 4504 9533
rect 4508 9529 4509 9533
rect 4529 9544 4530 9548
rect 4534 9544 4535 9548
rect 4539 9544 4540 9548
rect 4544 9544 4545 9548
rect 4549 9544 4550 9548
rect 4554 9544 4555 9548
rect 4525 9543 4559 9544
rect 4529 9539 4530 9543
rect 4534 9539 4535 9543
rect 4539 9539 4540 9543
rect 4544 9539 4545 9543
rect 4549 9539 4550 9543
rect 4554 9539 4555 9543
rect 4525 9538 4559 9539
rect 4529 9534 4530 9538
rect 4534 9534 4535 9538
rect 4539 9534 4540 9538
rect 4544 9534 4545 9538
rect 4549 9534 4550 9538
rect 4554 9534 4555 9538
rect 4525 9533 4559 9534
rect 4529 9529 4530 9533
rect 4534 9529 4535 9533
rect 4539 9529 4540 9533
rect 4544 9529 4545 9533
rect 4549 9529 4550 9533
rect 4554 9529 4555 9533
rect 4483 9515 4484 9519
rect 4488 9515 4489 9519
rect 4493 9515 4494 9519
rect 4498 9515 4499 9519
rect 4503 9515 4504 9519
rect 4508 9515 4509 9519
rect 4479 9514 4513 9515
rect 4483 9510 4484 9514
rect 4488 9510 4489 9514
rect 4493 9510 4494 9514
rect 4498 9510 4499 9514
rect 4503 9510 4504 9514
rect 4508 9510 4509 9514
rect 4479 9509 4513 9510
rect 4483 9505 4484 9509
rect 4488 9505 4489 9509
rect 4493 9505 4494 9509
rect 4498 9505 4499 9509
rect 4503 9505 4504 9509
rect 4508 9505 4509 9509
rect 4479 9504 4513 9505
rect 4483 9500 4484 9504
rect 4488 9500 4489 9504
rect 4493 9500 4494 9504
rect 4498 9500 4499 9504
rect 4503 9500 4504 9504
rect 4508 9500 4509 9504
rect 4529 9515 4530 9519
rect 4534 9515 4535 9519
rect 4539 9515 4540 9519
rect 4544 9515 4545 9519
rect 4549 9515 4550 9519
rect 4554 9515 4555 9519
rect 4525 9514 4559 9515
rect 4529 9510 4530 9514
rect 4534 9510 4535 9514
rect 4539 9510 4540 9514
rect 4544 9510 4545 9514
rect 4549 9510 4550 9514
rect 4554 9510 4555 9514
rect 4525 9509 4559 9510
rect 4529 9505 4530 9509
rect 4534 9505 4535 9509
rect 4539 9505 4540 9509
rect 4544 9505 4545 9509
rect 4549 9505 4550 9509
rect 4554 9505 4555 9509
rect 4525 9504 4559 9505
rect 4529 9500 4530 9504
rect 4534 9500 4535 9504
rect 4539 9500 4540 9504
rect 4544 9500 4545 9504
rect 4549 9500 4550 9504
rect 4554 9500 4555 9504
rect 4483 9486 4484 9490
rect 4488 9486 4489 9490
rect 4493 9486 4494 9490
rect 4498 9486 4499 9490
rect 4503 9486 4504 9490
rect 4508 9486 4509 9490
rect 4479 9485 4513 9486
rect 4483 9481 4484 9485
rect 4488 9481 4489 9485
rect 4493 9481 4494 9485
rect 4498 9481 4499 9485
rect 4503 9481 4504 9485
rect 4508 9481 4509 9485
rect 4479 9480 4513 9481
rect 4483 9476 4484 9480
rect 4488 9476 4489 9480
rect 4493 9476 4494 9480
rect 4498 9476 4499 9480
rect 4503 9476 4504 9480
rect 4508 9476 4509 9480
rect 4479 9475 4513 9476
rect 4483 9471 4484 9475
rect 4488 9471 4489 9475
rect 4493 9471 4494 9475
rect 4498 9471 4499 9475
rect 4503 9471 4504 9475
rect 4508 9471 4509 9475
rect 4529 9486 4530 9490
rect 4534 9486 4535 9490
rect 4539 9486 4540 9490
rect 4544 9486 4545 9490
rect 4549 9486 4550 9490
rect 4554 9486 4555 9490
rect 4525 9485 4559 9486
rect 4529 9481 4530 9485
rect 4534 9481 4535 9485
rect 4539 9481 4540 9485
rect 4544 9481 4545 9485
rect 4549 9481 4550 9485
rect 4554 9481 4555 9485
rect 4525 9480 4559 9481
rect 4529 9476 4530 9480
rect 4534 9476 4535 9480
rect 4539 9476 4540 9480
rect 4544 9476 4545 9480
rect 4549 9476 4550 9480
rect 4554 9476 4555 9480
rect 4525 9475 4559 9476
rect 4529 9471 4530 9475
rect 4534 9471 4535 9475
rect 4539 9471 4540 9475
rect 4544 9471 4545 9475
rect 4549 9471 4550 9475
rect 4554 9471 4555 9475
rect 2842 9452 3781 9456
rect 3787 9452 3980 9456
rect 4483 9457 4484 9461
rect 4488 9457 4489 9461
rect 4493 9457 4494 9461
rect 4498 9457 4499 9461
rect 4503 9457 4504 9461
rect 4508 9457 4509 9461
rect 4479 9456 4513 9457
rect 4483 9452 4484 9456
rect 4488 9452 4489 9456
rect 4493 9452 4494 9456
rect 4498 9452 4499 9456
rect 4503 9452 4504 9456
rect 4508 9452 4509 9456
rect 4479 9451 4513 9452
rect 3053 9444 3423 9448
rect 4483 9447 4484 9451
rect 4488 9447 4489 9451
rect 4493 9447 4494 9451
rect 4498 9447 4499 9451
rect 4503 9447 4504 9451
rect 4508 9447 4509 9451
rect 4479 9446 4513 9447
rect 4483 9442 4484 9446
rect 4488 9442 4489 9446
rect 4493 9442 4494 9446
rect 4498 9442 4499 9446
rect 4503 9442 4504 9446
rect 4508 9442 4509 9446
rect 4529 9457 4530 9461
rect 4534 9457 4535 9461
rect 4539 9457 4540 9461
rect 4544 9457 4545 9461
rect 4549 9457 4550 9461
rect 4554 9457 4555 9461
rect 4525 9456 4559 9457
rect 4529 9452 4530 9456
rect 4534 9452 4535 9456
rect 4539 9452 4540 9456
rect 4544 9452 4545 9456
rect 4549 9452 4550 9456
rect 4554 9452 4555 9456
rect 4525 9451 4559 9452
rect 4529 9447 4530 9451
rect 4534 9447 4535 9451
rect 4539 9447 4540 9451
rect 4544 9447 4545 9451
rect 4549 9447 4550 9451
rect 4554 9447 4555 9451
rect 4525 9446 4559 9447
rect 4529 9442 4530 9446
rect 4534 9442 4535 9446
rect 4539 9442 4540 9446
rect 4544 9442 4545 9446
rect 4549 9442 4550 9446
rect 4554 9442 4555 9446
rect 3026 9434 3411 9438
rect 4579 9355 5073 9786
rect 2830 9347 2857 9351
rect 2861 9347 2893 9351
rect 2897 9347 2960 9351
rect 2964 9347 2989 9351
rect 2993 9347 3025 9351
rect 3029 9347 3092 9351
rect 3096 9347 3121 9351
rect 3125 9347 3157 9351
rect 3161 9347 3224 9351
rect 3228 9347 3253 9351
rect 3257 9347 3289 9351
rect 3293 9347 3356 9351
rect 3360 9347 3376 9351
rect 3775 9347 3802 9351
rect 3806 9347 3838 9351
rect 3842 9347 3905 9351
rect 3909 9347 3934 9351
rect 3938 9347 3970 9351
rect 3974 9347 4037 9351
rect 4041 9347 4066 9351
rect 4070 9347 4102 9351
rect 4106 9347 4169 9351
rect 4173 9347 4198 9351
rect 4202 9347 4234 9351
rect 4238 9347 4301 9351
rect 4305 9347 4321 9351
rect 2770 9340 2881 9344
rect 2885 9340 2909 9344
rect 2913 9340 2939 9344
rect 2943 9340 2976 9344
rect 2980 9340 3013 9344
rect 3017 9340 3041 9344
rect 3045 9340 3071 9344
rect 3075 9340 3108 9344
rect 3112 9340 3145 9344
rect 3149 9340 3173 9344
rect 3177 9340 3203 9344
rect 3207 9340 3240 9344
rect 3244 9340 3277 9344
rect 3281 9340 3305 9344
rect 3309 9340 3335 9344
rect 3339 9340 3372 9344
rect 3715 9340 3826 9344
rect 3830 9340 3854 9344
rect 3858 9340 3884 9344
rect 3888 9340 3921 9344
rect 3925 9340 3958 9344
rect 3962 9340 3986 9344
rect 3990 9340 4016 9344
rect 4020 9340 4053 9344
rect 4057 9340 4090 9344
rect 4094 9340 4118 9344
rect 4122 9340 4148 9344
rect 4152 9340 4185 9344
rect 4189 9340 4222 9344
rect 4226 9340 4250 9344
rect 4254 9340 4280 9344
rect 4284 9340 4317 9344
rect 2851 9330 2854 9340
rect 2872 9330 2875 9340
rect 2888 9330 2891 9340
rect 2902 9333 2907 9337
rect 2911 9333 2918 9337
rect 2930 9330 2933 9340
rect 2946 9330 2949 9340
rect 2967 9330 2970 9340
rect 2983 9330 2986 9340
rect 3004 9330 3007 9340
rect 3020 9330 3023 9340
rect 3034 9333 3039 9337
rect 3043 9333 3050 9337
rect 3062 9330 3065 9340
rect 3078 9330 3081 9340
rect 3099 9330 3102 9340
rect 3115 9330 3118 9340
rect 3136 9330 3139 9340
rect 3152 9330 3155 9340
rect 3166 9333 3171 9337
rect 3175 9333 3182 9337
rect 3194 9330 3197 9340
rect 3210 9330 3213 9340
rect 3231 9330 3234 9340
rect 3247 9330 3250 9340
rect 3268 9330 3271 9340
rect 3284 9330 3287 9340
rect 3298 9333 3303 9337
rect 3307 9333 3314 9337
rect 3326 9330 3329 9340
rect 3342 9330 3345 9340
rect 3363 9330 3366 9340
rect 3796 9330 3799 9340
rect 3817 9330 3820 9340
rect 3833 9330 3836 9340
rect 3847 9333 3852 9337
rect 3856 9333 3863 9337
rect 3875 9330 3878 9340
rect 3891 9330 3894 9340
rect 3912 9330 3915 9340
rect 3928 9330 3931 9340
rect 3949 9330 3952 9340
rect 3965 9330 3968 9340
rect 3979 9333 3984 9337
rect 3988 9333 3995 9337
rect 4007 9330 4010 9340
rect 4023 9330 4026 9340
rect 4044 9330 4047 9340
rect 4060 9330 4063 9340
rect 4081 9330 4084 9340
rect 4097 9330 4100 9340
rect 4111 9333 4116 9337
rect 4120 9333 4127 9337
rect 4139 9330 4142 9340
rect 4155 9330 4158 9340
rect 4176 9330 4179 9340
rect 4192 9330 4195 9340
rect 4213 9330 4216 9340
rect 4229 9330 4232 9340
rect 4243 9333 4248 9337
rect 4252 9333 4259 9337
rect 4271 9330 4274 9340
rect 4287 9330 4290 9340
rect 4308 9330 4311 9340
rect 617 9321 618 9325
rect 622 9321 623 9325
rect 627 9321 628 9325
rect 632 9321 633 9325
rect 637 9321 638 9325
rect 642 9321 643 9325
rect 613 9320 647 9321
rect 617 9316 618 9320
rect 622 9316 623 9320
rect 627 9316 628 9320
rect 632 9316 633 9320
rect 637 9316 638 9320
rect 642 9316 643 9320
rect 613 9315 647 9316
rect 617 9311 618 9315
rect 622 9311 623 9315
rect 627 9311 628 9315
rect 632 9311 633 9315
rect 637 9311 638 9315
rect 642 9311 643 9315
rect 613 9310 647 9311
rect 86 9304 346 9307
rect 617 9306 618 9310
rect 622 9306 623 9310
rect 627 9306 628 9310
rect 632 9306 633 9310
rect 637 9306 638 9310
rect 642 9306 643 9310
rect 663 9321 664 9325
rect 668 9321 669 9325
rect 673 9321 674 9325
rect 678 9321 679 9325
rect 683 9321 684 9325
rect 688 9321 689 9325
rect 659 9320 693 9321
rect 663 9316 664 9320
rect 668 9316 669 9320
rect 673 9316 674 9320
rect 678 9316 679 9320
rect 683 9316 684 9320
rect 688 9316 689 9320
rect 659 9315 693 9316
rect 663 9311 664 9315
rect 668 9311 669 9315
rect 673 9311 674 9315
rect 678 9311 679 9315
rect 683 9311 684 9315
rect 688 9311 689 9315
rect 2496 9314 2505 9318
rect 2509 9314 2541 9318
rect 2545 9314 2608 9318
rect 2612 9314 2824 9318
rect 2868 9316 2873 9319
rect 2877 9316 2901 9319
rect 2926 9316 2933 9319
rect 2937 9316 2959 9319
rect 659 9310 693 9311
rect 663 9306 664 9310
rect 668 9306 669 9310
rect 673 9306 674 9310
rect 678 9306 679 9310
rect 683 9306 684 9310
rect 688 9306 689 9310
rect 2496 9307 2529 9311
rect 2533 9307 2557 9311
rect 2561 9307 2587 9311
rect 2591 9307 2624 9311
rect 2628 9307 2764 9311
rect 86 9050 89 9304
rect 343 9265 346 9304
rect 2499 9297 2502 9307
rect 2520 9297 2523 9307
rect 2536 9297 2539 9307
rect 2550 9300 2555 9304
rect 2559 9300 2566 9304
rect 2578 9297 2581 9307
rect 2594 9297 2597 9307
rect 2615 9297 2618 9307
rect 2884 9306 2891 9309
rect 2895 9310 2914 9313
rect 2914 9303 2917 9309
rect 2942 9306 2949 9309
rect 2953 9310 2970 9313
rect 3000 9316 3005 9319
rect 3009 9316 3033 9319
rect 3058 9316 3065 9319
rect 3069 9316 3091 9319
rect 3016 9306 3023 9309
rect 3027 9310 3046 9313
rect 3046 9303 3049 9309
rect 3074 9306 3081 9309
rect 3085 9310 3102 9313
rect 3132 9316 3137 9319
rect 3141 9316 3165 9319
rect 3190 9316 3197 9319
rect 3201 9316 3223 9319
rect 3148 9306 3155 9309
rect 3159 9310 3178 9313
rect 3178 9303 3181 9309
rect 3206 9306 3213 9309
rect 3217 9310 3234 9313
rect 3264 9316 3269 9319
rect 3273 9316 3297 9319
rect 3322 9316 3329 9319
rect 3333 9316 3355 9319
rect 3441 9314 3450 9318
rect 3454 9314 3486 9318
rect 3490 9314 3553 9318
rect 3557 9314 3769 9318
rect 3280 9306 3287 9309
rect 3291 9310 3310 9313
rect 2494 9280 2503 9284
rect 2516 9283 2521 9286
rect 2525 9283 2549 9286
rect 2574 9283 2581 9286
rect 2585 9283 2607 9286
rect 2851 9287 2854 9299
rect 2872 9287 2875 9299
rect 2888 9287 2891 9299
rect 2902 9290 2914 9293
rect 2930 9287 2933 9299
rect 2946 9287 2949 9299
rect 2967 9287 2970 9299
rect 2983 9287 2986 9299
rect 3004 9287 3007 9299
rect 3020 9287 3023 9299
rect 3034 9290 3046 9293
rect 3062 9287 3065 9299
rect 3078 9287 3081 9299
rect 3099 9287 3102 9299
rect 3115 9287 3118 9299
rect 3136 9287 3139 9299
rect 3152 9287 3155 9299
rect 3166 9290 3178 9293
rect 3194 9287 3197 9299
rect 3210 9287 3213 9299
rect 3231 9287 3234 9299
rect 3310 9303 3313 9309
rect 3338 9306 3345 9309
rect 3349 9310 3366 9313
rect 3813 9316 3818 9319
rect 3822 9316 3846 9319
rect 3871 9316 3878 9319
rect 3882 9316 3904 9319
rect 3441 9307 3474 9311
rect 3478 9307 3502 9311
rect 3506 9307 3532 9311
rect 3536 9307 3569 9311
rect 3573 9307 3709 9311
rect 3247 9287 3250 9299
rect 3268 9287 3271 9299
rect 3284 9287 3287 9299
rect 3298 9290 3310 9293
rect 3326 9287 3329 9299
rect 3342 9287 3345 9299
rect 3363 9287 3366 9299
rect 3444 9297 3447 9307
rect 3465 9297 3468 9307
rect 3481 9297 3484 9307
rect 3495 9300 3500 9304
rect 3504 9300 3511 9304
rect 3523 9297 3526 9307
rect 3539 9297 3542 9307
rect 3560 9297 3563 9307
rect 3829 9306 3836 9309
rect 3840 9310 3859 9313
rect 3859 9303 3862 9309
rect 3887 9306 3894 9309
rect 3898 9310 3915 9313
rect 3945 9316 3950 9319
rect 3954 9316 3978 9319
rect 4003 9316 4010 9319
rect 4014 9316 4036 9319
rect 3961 9306 3968 9309
rect 3972 9310 3991 9313
rect 3991 9303 3994 9309
rect 4019 9306 4026 9309
rect 4030 9310 4047 9313
rect 4077 9316 4082 9319
rect 4086 9316 4110 9319
rect 4135 9316 4142 9319
rect 4146 9316 4168 9319
rect 4093 9306 4100 9309
rect 4104 9310 4123 9313
rect 4123 9303 4126 9309
rect 4151 9306 4158 9309
rect 4162 9310 4179 9313
rect 4209 9316 4214 9319
rect 4218 9316 4242 9319
rect 4267 9316 4274 9319
rect 4278 9316 4300 9319
rect 4826 9316 5086 9319
rect 4225 9306 4232 9309
rect 4236 9310 4255 9313
rect 2782 9283 2881 9287
rect 2885 9283 2909 9287
rect 2913 9283 2939 9287
rect 2943 9283 3013 9287
rect 3017 9283 3041 9287
rect 3045 9283 3071 9287
rect 3075 9283 3145 9287
rect 3149 9283 3173 9287
rect 3177 9283 3203 9287
rect 3207 9283 3277 9287
rect 3281 9283 3305 9287
rect 3309 9283 3335 9287
rect 3339 9283 3376 9287
rect 2532 9273 2539 9276
rect 2543 9277 2562 9280
rect 2562 9270 2565 9276
rect 2590 9273 2597 9276
rect 2601 9277 2616 9280
rect 3439 9280 3448 9284
rect 3461 9283 3466 9286
rect 3470 9283 3494 9286
rect 3519 9283 3526 9286
rect 3530 9283 3552 9286
rect 3796 9287 3799 9299
rect 3817 9287 3820 9299
rect 3833 9287 3836 9299
rect 3847 9290 3859 9293
rect 3875 9287 3878 9299
rect 3891 9287 3894 9299
rect 3912 9287 3915 9299
rect 3928 9287 3931 9299
rect 3949 9287 3952 9299
rect 3965 9287 3968 9299
rect 3979 9290 3991 9293
rect 4007 9287 4010 9299
rect 4023 9287 4026 9299
rect 4044 9287 4047 9299
rect 4060 9287 4063 9299
rect 4081 9287 4084 9299
rect 4097 9287 4100 9299
rect 4111 9290 4123 9293
rect 4139 9287 4142 9299
rect 4155 9287 4158 9299
rect 4176 9287 4179 9299
rect 4255 9303 4258 9309
rect 4283 9306 4290 9309
rect 4294 9310 4311 9313
rect 4192 9287 4195 9299
rect 4213 9287 4216 9299
rect 4229 9287 4232 9299
rect 4243 9290 4255 9293
rect 4271 9287 4274 9299
rect 4287 9287 4290 9299
rect 4308 9287 4311 9299
rect 3727 9283 3826 9287
rect 3830 9283 3854 9287
rect 3858 9283 3884 9287
rect 3888 9283 3958 9287
rect 3962 9283 3986 9287
rect 3990 9283 4016 9287
rect 4020 9283 4090 9287
rect 4094 9283 4118 9287
rect 4122 9283 4148 9287
rect 4152 9283 4222 9287
rect 4226 9283 4250 9287
rect 4254 9283 4280 9287
rect 4284 9283 4321 9287
rect 2818 9276 2857 9280
rect 2861 9276 2908 9280
rect 2912 9276 2958 9280
rect 2962 9276 2989 9280
rect 2993 9276 3040 9280
rect 3044 9276 3090 9280
rect 3094 9276 3121 9280
rect 3125 9276 3172 9280
rect 3176 9276 3222 9280
rect 3226 9276 3253 9280
rect 3257 9276 3304 9280
rect 3308 9276 3354 9280
rect 3358 9276 3376 9280
rect 3477 9273 3484 9276
rect 3488 9277 3507 9280
rect 343 9255 356 9265
rect 343 9245 366 9255
rect 2499 9254 2502 9266
rect 2520 9254 2523 9266
rect 2536 9254 2539 9266
rect 2550 9257 2562 9260
rect 2578 9254 2581 9266
rect 2594 9254 2597 9266
rect 2615 9254 2618 9266
rect 2770 9263 2855 9267
rect 2859 9263 2871 9267
rect 2875 9263 2889 9267
rect 2893 9263 2900 9267
rect 2904 9263 2906 9267
rect 2910 9263 2925 9267
rect 2929 9263 2962 9267
rect 2966 9263 2967 9267
rect 2971 9263 2979 9267
rect 2983 9263 3007 9267
rect 3011 9263 3023 9267
rect 3027 9263 3047 9267
rect 3051 9263 3101 9267
rect 3105 9263 3128 9267
rect 3132 9263 3182 9267
rect 3186 9263 3205 9267
rect 3507 9270 3510 9276
rect 3535 9273 3542 9276
rect 3546 9277 3561 9280
rect 3763 9276 3802 9280
rect 3806 9276 3853 9280
rect 3857 9276 3903 9280
rect 3907 9276 3934 9280
rect 3938 9276 3985 9280
rect 3989 9276 4035 9280
rect 4039 9276 4066 9280
rect 4070 9276 4117 9280
rect 4121 9276 4167 9280
rect 4171 9276 4198 9280
rect 4202 9276 4249 9280
rect 4253 9276 4299 9280
rect 4303 9276 4321 9280
rect 4826 9277 4829 9316
rect 4816 9267 4829 9277
rect 2806 9256 2882 9260
rect 2886 9256 2913 9260
rect 2917 9256 2935 9260
rect 2939 9256 3000 9260
rect 3004 9256 3018 9260
rect 3030 9259 3033 9263
rect 2496 9250 2529 9254
rect 2533 9250 2557 9254
rect 2561 9250 2587 9254
rect 2591 9250 2776 9254
rect 343 9235 376 9245
rect 2496 9243 2505 9247
rect 2509 9243 2556 9247
rect 2560 9243 2606 9247
rect 2610 9243 2812 9247
rect 2925 9249 2928 9253
rect 2952 9249 2953 9253
rect 2997 9249 2999 9253
rect 3039 9246 3042 9251
rect 3054 9253 3057 9263
rect 3084 9259 3087 9263
rect 3111 9259 3114 9263
rect 343 9225 386 9235
rect 2494 9227 2510 9231
rect 2619 9229 2623 9233
rect 2635 9229 2639 9233
rect 2643 9229 2857 9233
rect 2865 9232 2868 9238
rect 2872 9232 2875 9238
rect 2865 9229 2875 9232
rect 343 9129 769 9225
rect 2865 9224 2868 9229
rect 2502 9220 2506 9224
rect 2518 9220 2639 9224
rect 2872 9224 2875 9229
rect 2881 9234 2884 9238
rect 2881 9230 2883 9234
rect 2887 9230 2889 9234
rect 2897 9233 2900 9238
rect 2925 9235 2928 9238
rect 2897 9231 2908 9233
rect 2881 9224 2884 9230
rect 2897 9229 2903 9231
rect 2897 9224 2900 9229
rect 2907 9229 2908 9231
rect 2926 9231 2928 9235
rect 2925 9224 2928 9231
rect 3028 9242 3031 9245
rect 3070 9242 3073 9245
rect 2941 9234 2944 9238
rect 2951 9234 2954 9238
rect 2951 9230 2960 9234
rect 2972 9233 2975 9238
rect 2997 9234 3000 9238
rect 2941 9224 2944 9230
rect 2951 9224 2954 9230
rect 2972 9229 2973 9233
rect 2977 9229 2980 9232
rect 2999 9230 3000 9234
rect 3015 9233 3018 9238
rect 3039 9237 3042 9242
rect 3047 9238 3058 9241
rect 3070 9239 3078 9242
rect 2972 9224 2975 9229
rect 2997 9224 3000 9230
rect 3015 9224 3018 9229
rect 2489 9212 2505 9216
rect 2509 9212 2572 9216
rect 2576 9212 2608 9216
rect 2612 9212 2824 9216
rect 2917 9211 2918 9215
rect 2942 9212 2943 9216
rect 2989 9211 2990 9215
rect 2493 9205 2526 9209
rect 2530 9205 2556 9209
rect 2560 9205 2584 9209
rect 2588 9205 2764 9209
rect 2499 9195 2502 9205
rect 2520 9195 2523 9205
rect 2536 9195 2539 9205
rect 2551 9198 2558 9202
rect 2562 9198 2567 9202
rect 2578 9195 2581 9205
rect 2594 9195 2597 9205
rect 2615 9195 2618 9205
rect 2794 9204 2870 9208
rect 2874 9204 2929 9208
rect 2933 9204 2954 9208
rect 2958 9204 2985 9208
rect 2989 9204 3018 9208
rect 3030 9201 3033 9233
rect 3047 9232 3050 9238
rect 3070 9233 3073 9239
rect 3082 9234 3085 9237
rect 3093 9237 3096 9251
rect 3120 9246 3123 9251
rect 3135 9253 3138 9263
rect 3165 9259 3168 9263
rect 3104 9242 3105 9245
rect 3109 9242 3112 9245
rect 3151 9242 3154 9245
rect 3093 9234 3101 9237
rect 3120 9237 3123 9242
rect 3093 9229 3096 9234
rect 3101 9230 3105 9234
rect 3128 9238 3139 9241
rect 3151 9239 3159 9242
rect 3045 9223 3050 9228
rect 3054 9201 3057 9229
rect 3084 9201 3087 9225
rect 3111 9201 3114 9233
rect 3128 9232 3131 9238
rect 3151 9233 3154 9239
rect 3163 9234 3166 9237
rect 3174 9237 3177 9251
rect 3328 9250 3411 9258
rect 3444 9254 3447 9266
rect 3465 9254 3468 9266
rect 3481 9254 3484 9266
rect 3495 9257 3507 9260
rect 3523 9254 3526 9266
rect 3539 9254 3542 9266
rect 3560 9254 3563 9266
rect 3715 9263 3800 9267
rect 3804 9263 3816 9267
rect 3820 9263 3834 9267
rect 3838 9263 3845 9267
rect 3849 9263 3851 9267
rect 3855 9263 3870 9267
rect 3874 9263 3907 9267
rect 3911 9263 3912 9267
rect 3916 9263 3924 9267
rect 3928 9263 3952 9267
rect 3956 9263 3968 9267
rect 3972 9263 3992 9267
rect 3996 9263 4046 9267
rect 4050 9263 4073 9267
rect 4077 9263 4127 9267
rect 4131 9263 4150 9267
rect 3751 9256 3827 9260
rect 3831 9256 3858 9260
rect 3862 9256 3880 9260
rect 3884 9256 3945 9260
rect 3949 9256 3963 9260
rect 3975 9259 3978 9263
rect 3441 9250 3474 9254
rect 3478 9250 3502 9254
rect 3506 9250 3532 9254
rect 3536 9250 3721 9254
rect 3365 9241 3423 9245
rect 3441 9243 3450 9247
rect 3454 9243 3501 9247
rect 3505 9243 3551 9247
rect 3555 9243 3757 9247
rect 3870 9249 3873 9253
rect 3897 9249 3898 9253
rect 3942 9249 3944 9253
rect 3984 9246 3987 9251
rect 3999 9253 4002 9263
rect 4029 9259 4032 9263
rect 4056 9259 4059 9263
rect 3174 9234 3186 9237
rect 3174 9229 3177 9234
rect 3126 9223 3131 9228
rect 3135 9201 3138 9229
rect 3439 9227 3455 9231
rect 3564 9229 3568 9233
rect 3580 9229 3584 9233
rect 3588 9229 3802 9233
rect 3810 9232 3813 9238
rect 3817 9232 3820 9238
rect 3810 9229 3820 9232
rect 3165 9201 3168 9225
rect 3810 9224 3813 9229
rect 3447 9220 3451 9224
rect 3463 9220 3584 9224
rect 3817 9224 3820 9229
rect 3826 9234 3829 9238
rect 3826 9230 3828 9234
rect 3832 9230 3834 9234
rect 3842 9233 3845 9238
rect 3870 9235 3873 9238
rect 3842 9231 3853 9233
rect 3826 9224 3829 9230
rect 3842 9229 3848 9231
rect 3842 9224 3845 9229
rect 3852 9229 3853 9231
rect 3871 9231 3873 9235
rect 3870 9224 3873 9231
rect 3973 9242 3976 9245
rect 4015 9242 4018 9245
rect 3886 9234 3889 9238
rect 3896 9234 3899 9238
rect 3896 9230 3905 9234
rect 3917 9233 3920 9238
rect 3942 9234 3945 9238
rect 3886 9224 3889 9230
rect 3896 9224 3899 9230
rect 3917 9229 3918 9233
rect 3922 9229 3925 9232
rect 3944 9230 3945 9234
rect 3960 9233 3963 9238
rect 3984 9237 3987 9242
rect 3992 9238 4003 9241
rect 4015 9239 4023 9242
rect 3917 9224 3920 9229
rect 3942 9224 3945 9230
rect 3960 9224 3963 9229
rect 3434 9212 3450 9216
rect 3454 9212 3517 9216
rect 3521 9212 3553 9216
rect 3557 9212 3769 9216
rect 3862 9211 3863 9215
rect 3887 9212 3888 9216
rect 3934 9211 3935 9215
rect 3438 9205 3471 9209
rect 3475 9205 3501 9209
rect 3505 9205 3529 9209
rect 3533 9205 3709 9209
rect 2782 9197 2856 9201
rect 2860 9197 2862 9201
rect 2866 9197 2870 9201
rect 2874 9197 2888 9201
rect 2892 9197 2897 9201
rect 2901 9197 2906 9201
rect 2910 9197 2929 9201
rect 2933 9197 2963 9201
rect 2967 9197 2978 9201
rect 2982 9197 3006 9201
rect 3010 9197 3023 9201
rect 3027 9197 3047 9201
rect 3051 9197 3101 9201
rect 3108 9197 3128 9201
rect 3132 9197 3182 9201
rect 2510 9181 2532 9184
rect 2536 9181 2543 9184
rect 2794 9190 2870 9194
rect 2874 9190 2929 9194
rect 2933 9190 2954 9194
rect 2958 9190 2985 9194
rect 2989 9190 3018 9194
rect 2568 9181 2592 9184
rect 2596 9181 2601 9184
rect 2917 9183 2918 9187
rect 2942 9182 2943 9186
rect 2989 9183 2990 9187
rect 2614 9178 2623 9182
rect 2501 9175 2516 9178
rect 2555 9175 2574 9178
rect 2520 9171 2527 9174
rect 2552 9168 2555 9174
rect 2578 9171 2585 9174
rect 2865 9169 2868 9174
rect 2872 9169 2875 9174
rect 2855 9166 2857 9169
rect 2865 9166 2875 9169
rect 2499 9152 2502 9164
rect 2520 9152 2523 9164
rect 2536 9152 2539 9164
rect 2555 9155 2567 9158
rect 2578 9152 2581 9164
rect 2594 9152 2597 9164
rect 2615 9152 2618 9164
rect 2865 9160 2868 9166
rect 2872 9160 2875 9166
rect 2881 9168 2884 9174
rect 2897 9169 2900 9174
rect 2881 9164 2883 9168
rect 2887 9164 2889 9168
rect 2897 9167 2903 9169
rect 2907 9167 2908 9169
rect 2897 9165 2908 9167
rect 2925 9167 2928 9174
rect 2881 9160 2884 9164
rect 2897 9160 2900 9165
rect 2926 9163 2928 9167
rect 2925 9160 2928 9163
rect 2941 9168 2944 9174
rect 2951 9168 2954 9174
rect 2972 9169 2975 9174
rect 2951 9164 2960 9168
rect 2972 9165 2973 9169
rect 2977 9166 2980 9169
rect 2997 9168 3000 9174
rect 3015 9169 3018 9174
rect 3054 9177 3057 9197
rect 3135 9177 3138 9197
rect 3444 9195 3447 9205
rect 3465 9195 3468 9205
rect 3481 9195 3484 9205
rect 3496 9198 3503 9202
rect 3507 9198 3512 9202
rect 3523 9195 3526 9205
rect 3539 9195 3542 9205
rect 3560 9195 3563 9205
rect 3739 9204 3815 9208
rect 3819 9204 3874 9208
rect 3878 9204 3899 9208
rect 3903 9204 3930 9208
rect 3934 9204 3963 9208
rect 3975 9201 3978 9233
rect 3992 9232 3995 9238
rect 4015 9233 4018 9239
rect 4027 9234 4030 9237
rect 4038 9237 4041 9251
rect 4065 9246 4068 9251
rect 4080 9253 4083 9263
rect 4110 9259 4113 9263
rect 4049 9242 4050 9245
rect 4054 9242 4057 9245
rect 4806 9257 4829 9267
rect 4096 9242 4099 9245
rect 4038 9234 4046 9237
rect 4065 9237 4068 9242
rect 4038 9229 4041 9234
rect 4046 9230 4050 9234
rect 4073 9238 4084 9241
rect 4096 9239 4104 9242
rect 3990 9223 3995 9228
rect 3999 9201 4002 9229
rect 4029 9201 4032 9225
rect 4056 9201 4059 9233
rect 4073 9232 4076 9238
rect 4096 9233 4099 9239
rect 4108 9234 4111 9237
rect 4119 9237 4122 9251
rect 4796 9247 4829 9257
rect 4119 9234 4131 9237
rect 4786 9237 4829 9247
rect 4119 9229 4122 9234
rect 4071 9223 4076 9228
rect 4080 9201 4083 9229
rect 4110 9201 4113 9225
rect 3727 9197 3801 9201
rect 3805 9197 3807 9201
rect 3811 9197 3815 9201
rect 3819 9197 3833 9201
rect 3837 9197 3842 9201
rect 3846 9197 3851 9201
rect 3855 9197 3874 9201
rect 3878 9197 3908 9201
rect 3912 9197 3923 9201
rect 3927 9197 3951 9201
rect 3955 9197 3968 9201
rect 3972 9197 3992 9201
rect 3996 9197 4046 9201
rect 4053 9197 4073 9201
rect 4077 9197 4127 9201
rect 3455 9181 3477 9184
rect 3481 9181 3488 9184
rect 3739 9190 3815 9194
rect 3819 9190 3874 9194
rect 3878 9190 3899 9194
rect 3903 9190 3930 9194
rect 3934 9190 3963 9194
rect 3513 9181 3537 9184
rect 3541 9181 3546 9184
rect 3862 9183 3863 9187
rect 3887 9182 3888 9186
rect 3934 9183 3935 9187
rect 3559 9178 3568 9182
rect 3446 9175 3461 9178
rect 2941 9160 2944 9164
rect 2951 9160 2954 9164
rect 2972 9160 2975 9165
rect 2999 9164 3000 9168
rect 2997 9160 3000 9164
rect 3015 9160 3018 9165
rect 3045 9164 3050 9169
rect 3054 9165 3055 9168
rect 3070 9167 3073 9173
rect 3070 9164 3078 9167
rect 3125 9164 3130 9169
rect 3134 9165 3136 9168
rect 3151 9167 3154 9173
rect 3500 9175 3519 9178
rect 3465 9171 3472 9174
rect 3497 9168 3500 9174
rect 3151 9164 3159 9167
rect 3523 9171 3530 9174
rect 3810 9169 3813 9174
rect 3817 9169 3820 9174
rect 3800 9166 3802 9169
rect 3810 9166 3820 9169
rect 3070 9161 3073 9164
rect 3151 9161 3154 9164
rect 2489 9148 2526 9152
rect 2530 9148 2556 9152
rect 2560 9148 2584 9152
rect 2588 9148 2776 9152
rect 2925 9145 2928 9149
rect 2952 9145 2953 9149
rect 2997 9145 2999 9149
rect 2489 9141 2507 9145
rect 2511 9141 2557 9145
rect 2561 9141 2608 9145
rect 2612 9141 2812 9145
rect 2870 9138 2882 9142
rect 2886 9138 2913 9142
rect 2917 9138 2935 9142
rect 2939 9138 3000 9142
rect 3004 9138 3018 9142
rect 3054 9135 3057 9153
rect 3135 9135 3138 9153
rect 3444 9152 3447 9164
rect 3465 9152 3468 9164
rect 3481 9152 3484 9164
rect 3500 9155 3512 9158
rect 3523 9152 3526 9164
rect 3539 9152 3542 9164
rect 3560 9152 3563 9164
rect 3810 9160 3813 9166
rect 3817 9160 3820 9166
rect 3826 9168 3829 9174
rect 3842 9169 3845 9174
rect 3826 9164 3828 9168
rect 3832 9164 3834 9168
rect 3842 9167 3848 9169
rect 3852 9167 3853 9169
rect 3842 9165 3853 9167
rect 3870 9167 3873 9174
rect 3826 9160 3829 9164
rect 3842 9160 3845 9165
rect 3871 9163 3873 9167
rect 3870 9160 3873 9163
rect 3886 9168 3889 9174
rect 3896 9168 3899 9174
rect 3917 9169 3920 9174
rect 3896 9164 3905 9168
rect 3917 9165 3918 9169
rect 3922 9166 3925 9169
rect 3942 9168 3945 9174
rect 3960 9169 3963 9174
rect 3999 9177 4002 9197
rect 4080 9177 4083 9197
rect 3886 9160 3889 9164
rect 3896 9160 3899 9164
rect 3917 9160 3920 9165
rect 3944 9164 3945 9168
rect 3942 9160 3945 9164
rect 3960 9160 3963 9165
rect 3990 9164 3995 9169
rect 3999 9165 4000 9168
rect 4015 9167 4018 9173
rect 4015 9164 4023 9167
rect 4070 9164 4075 9169
rect 4079 9165 4081 9168
rect 4096 9167 4099 9173
rect 4096 9164 4104 9167
rect 4015 9161 4018 9164
rect 4096 9161 4099 9164
rect 3434 9148 3471 9152
rect 3475 9148 3501 9152
rect 3505 9148 3529 9152
rect 3533 9148 3721 9152
rect 3870 9145 3873 9149
rect 3897 9145 3898 9149
rect 3942 9145 3944 9149
rect 3434 9141 3452 9145
rect 3456 9141 3502 9145
rect 3506 9141 3553 9145
rect 3557 9141 3757 9145
rect 3815 9138 3827 9142
rect 3831 9138 3858 9142
rect 3862 9138 3880 9142
rect 3884 9138 3945 9142
rect 3949 9138 3963 9142
rect 3999 9135 4002 9153
rect 4080 9135 4083 9153
rect 4403 9141 4829 9237
rect 2770 9131 2855 9135
rect 2859 9131 2871 9135
rect 2875 9131 2889 9135
rect 2893 9131 2900 9135
rect 2904 9131 2906 9135
rect 2910 9131 2925 9135
rect 2929 9131 2962 9135
rect 2966 9131 2967 9135
rect 2971 9131 2979 9135
rect 2983 9131 3007 9135
rect 3011 9131 3023 9135
rect 3027 9131 3047 9135
rect 3051 9131 3101 9135
rect 3105 9131 3128 9135
rect 3132 9131 3190 9135
rect 3194 9131 3205 9135
rect 3715 9131 3800 9135
rect 3804 9131 3816 9135
rect 3820 9131 3834 9135
rect 3838 9131 3845 9135
rect 3849 9131 3851 9135
rect 3855 9131 3870 9135
rect 3874 9131 3907 9135
rect 3911 9131 3912 9135
rect 3916 9131 3924 9135
rect 3928 9131 3952 9135
rect 3956 9131 3968 9135
rect 3972 9131 3992 9135
rect 3996 9131 4046 9135
rect 4050 9131 4073 9135
rect 4077 9131 4135 9135
rect 4139 9131 4150 9135
rect 4786 9131 4829 9141
rect 343 9119 386 9129
rect 2806 9124 2866 9128
rect 2870 9124 2882 9128
rect 2886 9124 2913 9128
rect 2917 9124 2935 9128
rect 2939 9124 3000 9128
rect 3004 9124 3018 9128
rect 3054 9121 3057 9131
rect 3084 9127 3087 9131
rect 3135 9127 3138 9131
rect 343 9109 376 9119
rect 2925 9117 2928 9121
rect 2952 9117 2953 9121
rect 2997 9117 2999 9121
rect 343 9099 366 9109
rect 343 9089 356 9099
rect 2854 9097 2857 9100
rect 2865 9100 2868 9106
rect 2872 9100 2875 9106
rect 2865 9097 2875 9100
rect 2865 9092 2868 9097
rect 343 9050 346 9089
rect 2872 9092 2875 9097
rect 2881 9102 2884 9106
rect 2881 9098 2883 9102
rect 2887 9098 2889 9102
rect 2897 9101 2900 9106
rect 2925 9103 2928 9106
rect 2897 9099 2908 9101
rect 2881 9092 2884 9098
rect 2897 9097 2903 9099
rect 2897 9092 2900 9097
rect 2907 9097 2908 9099
rect 2926 9099 2928 9103
rect 2925 9092 2928 9099
rect 3070 9110 3073 9113
rect 2941 9102 2944 9106
rect 2951 9102 2954 9106
rect 2951 9098 2960 9102
rect 2972 9101 2975 9106
rect 2997 9102 3000 9106
rect 2941 9092 2944 9098
rect 2951 9092 2954 9098
rect 2972 9097 2973 9101
rect 2977 9097 2980 9100
rect 2999 9098 3000 9102
rect 3015 9101 3018 9106
rect 3047 9106 3058 9109
rect 3070 9107 3078 9110
rect 2972 9092 2975 9097
rect 2997 9092 3000 9098
rect 3047 9100 3050 9106
rect 3070 9101 3073 9107
rect 3082 9102 3085 9105
rect 3093 9105 3096 9119
rect 3144 9114 3147 9119
rect 3159 9121 3162 9131
rect 3189 9127 3192 9131
rect 3128 9110 3129 9113
rect 3133 9110 3136 9113
rect 3365 9120 3621 9125
rect 3751 9124 3811 9128
rect 3815 9124 3827 9128
rect 3831 9124 3858 9128
rect 3862 9124 3880 9128
rect 3884 9124 3945 9128
rect 3949 9124 3963 9128
rect 3999 9121 4002 9131
rect 4029 9127 4032 9131
rect 4080 9127 4083 9131
rect 3175 9110 3178 9113
rect 3101 9105 3106 9110
rect 3144 9105 3147 9110
rect 3093 9102 3101 9105
rect 3015 9092 3018 9097
rect 3093 9097 3096 9102
rect 3152 9106 3163 9109
rect 3175 9107 3183 9110
rect 3045 9091 3050 9096
rect 2917 9079 2918 9083
rect 2942 9080 2943 9084
rect 2989 9079 2990 9083
rect 2794 9072 2870 9076
rect 2874 9072 2929 9076
rect 2933 9072 2954 9076
rect 2958 9072 2985 9076
rect 2989 9072 3018 9076
rect 3054 9069 3057 9097
rect 3084 9069 3087 9093
rect 3135 9069 3138 9101
rect 3152 9100 3155 9106
rect 3175 9101 3178 9107
rect 3187 9102 3190 9105
rect 3198 9105 3201 9119
rect 3870 9117 3873 9121
rect 3897 9117 3898 9121
rect 3942 9117 3944 9121
rect 3198 9102 3204 9105
rect 3363 9102 3383 9106
rect 3387 9102 3437 9106
rect 3441 9102 3580 9106
rect 3584 9102 3668 9106
rect 3198 9097 3201 9102
rect 3150 9091 3155 9096
rect 3159 9069 3162 9097
rect 3366 9098 3369 9102
rect 3189 9069 3192 9093
rect 3375 9085 3378 9090
rect 3390 9092 3393 9102
rect 3420 9098 3423 9102
rect 3359 9081 3360 9084
rect 3364 9081 3367 9084
rect 3406 9081 3409 9084
rect 3375 9076 3378 9081
rect 3383 9077 3394 9080
rect 3406 9078 3414 9081
rect 3406 9072 3409 9078
rect 3418 9073 3421 9076
rect 3429 9076 3432 9090
rect 3540 9095 3543 9102
rect 3593 9095 3596 9102
rect 3799 9097 3802 9100
rect 3810 9100 3813 9106
rect 3817 9100 3820 9106
rect 3810 9097 3820 9100
rect 3429 9073 3441 9076
rect 2782 9065 2856 9069
rect 2860 9065 2862 9069
rect 2866 9065 2870 9069
rect 2874 9065 2888 9069
rect 2892 9065 2897 9069
rect 2901 9065 2906 9069
rect 2910 9065 2929 9069
rect 2933 9065 2963 9069
rect 2967 9065 2978 9069
rect 2982 9065 3006 9069
rect 3010 9065 3023 9069
rect 3027 9065 3047 9069
rect 3051 9065 3101 9069
rect 3105 9065 3128 9069
rect 3132 9065 3152 9069
rect 3156 9065 3204 9069
rect 2794 9058 2870 9062
rect 2874 9058 2929 9062
rect 2933 9058 2954 9062
rect 2958 9058 2985 9062
rect 2989 9058 3018 9062
rect 2917 9051 2918 9055
rect 2942 9050 2943 9054
rect 2989 9051 2990 9055
rect 86 9047 346 9050
rect 3054 9046 3057 9065
rect 3159 9046 3162 9065
rect 2865 9037 2868 9042
rect 2872 9037 2875 9042
rect 2855 9034 2857 9037
rect 2865 9034 2875 9037
rect 2865 9028 2868 9034
rect 2872 9028 2875 9034
rect 2881 9036 2884 9042
rect 2897 9037 2900 9042
rect 2881 9032 2883 9036
rect 2887 9032 2889 9036
rect 2897 9035 2903 9037
rect 2907 9035 2908 9037
rect 2897 9033 2908 9035
rect 2925 9035 2928 9042
rect 2881 9028 2884 9032
rect 2897 9028 2900 9033
rect 2926 9031 2928 9035
rect 2925 9028 2928 9031
rect 2941 9036 2944 9042
rect 2951 9036 2954 9042
rect 2972 9037 2975 9042
rect 2951 9032 2960 9036
rect 2972 9033 2973 9037
rect 2977 9034 2980 9037
rect 2997 9036 3000 9042
rect 3015 9037 3018 9042
rect 2941 9028 2944 9032
rect 2951 9028 2954 9032
rect 2972 9028 2975 9033
rect 2999 9032 3000 9036
rect 3044 9033 3049 9038
rect 3053 9034 3055 9037
rect 3070 9036 3073 9042
rect 3070 9033 3078 9036
rect 3150 9033 3155 9038
rect 3159 9034 3160 9037
rect 3175 9036 3178 9042
rect 3175 9033 3183 9036
rect 2997 9028 3000 9032
rect 3015 9028 3018 9033
rect 3070 9030 3073 9033
rect 3175 9030 3178 9033
rect 3366 9026 3369 9072
rect 3429 9068 3432 9073
rect 3390 9026 3393 9068
rect 3420 9026 3423 9064
rect 3438 9058 3441 9073
rect 3810 9092 3813 9097
rect 3817 9092 3820 9097
rect 3826 9102 3829 9106
rect 3826 9098 3828 9102
rect 3832 9098 3834 9102
rect 3842 9101 3845 9106
rect 3870 9103 3873 9106
rect 3842 9099 3853 9101
rect 3826 9092 3829 9098
rect 3842 9097 3848 9099
rect 3842 9092 3845 9097
rect 3852 9097 3853 9099
rect 3871 9099 3873 9103
rect 3870 9092 3873 9099
rect 4015 9110 4018 9113
rect 3886 9102 3889 9106
rect 3896 9102 3899 9106
rect 3896 9098 3905 9102
rect 3917 9101 3920 9106
rect 3942 9102 3945 9106
rect 3886 9092 3889 9098
rect 3896 9092 3899 9098
rect 3917 9097 3918 9101
rect 3922 9097 3925 9100
rect 3944 9098 3945 9102
rect 3960 9101 3963 9106
rect 3992 9106 4003 9109
rect 4015 9107 4023 9110
rect 3917 9092 3920 9097
rect 3942 9092 3945 9098
rect 3992 9100 3995 9106
rect 4015 9101 4018 9107
rect 4027 9102 4030 9105
rect 4038 9105 4041 9119
rect 4089 9114 4092 9119
rect 4104 9121 4107 9131
rect 4134 9127 4137 9131
rect 4073 9110 4074 9113
rect 4078 9110 4081 9113
rect 4796 9121 4829 9131
rect 4120 9110 4123 9113
rect 4046 9105 4051 9110
rect 4089 9105 4092 9110
rect 4038 9102 4046 9105
rect 3960 9092 3963 9097
rect 4038 9097 4041 9102
rect 4097 9106 4108 9109
rect 4120 9107 4128 9110
rect 3990 9091 3995 9096
rect 3862 9079 3863 9083
rect 3887 9080 3888 9084
rect 3934 9079 3935 9083
rect 3739 9072 3815 9076
rect 3819 9072 3874 9076
rect 3878 9072 3899 9076
rect 3903 9072 3930 9076
rect 3934 9072 3963 9076
rect 3999 9069 4002 9097
rect 4029 9069 4032 9093
rect 4080 9069 4083 9101
rect 4097 9100 4100 9106
rect 4120 9101 4123 9107
rect 4132 9102 4135 9105
rect 4143 9105 4146 9119
rect 4806 9111 4829 9121
rect 4143 9102 4149 9105
rect 4143 9097 4146 9102
rect 4816 9101 4829 9111
rect 4095 9091 4100 9096
rect 4104 9069 4107 9097
rect 4134 9069 4137 9093
rect 3727 9065 3801 9069
rect 3805 9065 3807 9069
rect 3811 9065 3815 9069
rect 3819 9065 3833 9069
rect 3837 9065 3842 9069
rect 3846 9065 3851 9069
rect 3855 9065 3874 9069
rect 3878 9065 3908 9069
rect 3912 9065 3923 9069
rect 3927 9065 3951 9069
rect 3955 9065 3968 9069
rect 3972 9065 3992 9069
rect 3996 9065 4046 9069
rect 4050 9065 4073 9069
rect 4077 9065 4097 9069
rect 4101 9065 4149 9069
rect 3438 9053 3555 9058
rect 3573 9057 3576 9065
rect 3573 9053 3593 9057
rect 3597 9053 3608 9057
rect 3573 9045 3576 9053
rect 3626 9049 3629 9065
rect 3739 9058 3815 9062
rect 3819 9058 3874 9062
rect 3878 9058 3899 9062
rect 3903 9058 3930 9062
rect 3934 9058 3963 9062
rect 3862 9051 3863 9055
rect 3887 9050 3888 9054
rect 3934 9051 3935 9055
rect 3630 9045 3745 9049
rect 3999 9046 4002 9065
rect 4104 9046 4107 9065
rect 4826 9062 4829 9101
rect 5083 9062 5086 9316
rect 4483 9056 4484 9060
rect 4488 9056 4489 9060
rect 4493 9056 4494 9060
rect 4498 9056 4499 9060
rect 4503 9056 4504 9060
rect 4508 9056 4509 9060
rect 4479 9055 4513 9056
rect 4483 9051 4484 9055
rect 4488 9051 4489 9055
rect 4493 9051 4494 9055
rect 4498 9051 4499 9055
rect 4503 9051 4504 9055
rect 4508 9051 4509 9055
rect 4479 9050 4513 9051
rect 4483 9046 4484 9050
rect 4488 9046 4489 9050
rect 4493 9046 4494 9050
rect 4498 9046 4499 9050
rect 4503 9046 4504 9050
rect 4508 9046 4509 9050
rect 3672 9033 3709 9037
rect 3810 9037 3813 9042
rect 3817 9037 3820 9042
rect 3800 9034 3802 9037
rect 3810 9034 3820 9037
rect 3540 9026 3543 9033
rect 3593 9026 3596 9033
rect 3660 9026 3721 9030
rect 3810 9028 3813 9034
rect 3363 9022 3383 9026
rect 3387 9022 3437 9026
rect 3441 9022 3580 9026
rect 3584 9022 3660 9026
rect 617 9012 618 9016
rect 622 9012 623 9016
rect 627 9012 628 9016
rect 632 9012 633 9016
rect 637 9012 638 9016
rect 642 9012 643 9016
rect 613 9011 647 9012
rect 617 9007 618 9011
rect 622 9007 623 9011
rect 627 9007 628 9011
rect 632 9007 633 9011
rect 637 9007 638 9011
rect 642 9007 643 9011
rect 613 9006 647 9007
rect 617 9002 618 9006
rect 622 9002 623 9006
rect 627 9002 628 9006
rect 632 9002 633 9006
rect 637 9002 638 9006
rect 642 9002 643 9006
rect 613 9001 647 9002
rect 86 8995 346 8998
rect 617 8997 618 9001
rect 622 8997 623 9001
rect 627 8997 628 9001
rect 632 8997 633 9001
rect 637 8997 638 9001
rect 642 8997 643 9001
rect 663 9012 664 9016
rect 668 9012 669 9016
rect 673 9012 674 9016
rect 678 9012 679 9016
rect 683 9012 684 9016
rect 688 9012 689 9016
rect 2925 9013 2928 9017
rect 2952 9013 2953 9017
rect 2997 9013 2999 9017
rect 659 9011 693 9012
rect 663 9007 664 9011
rect 668 9007 669 9011
rect 673 9007 674 9011
rect 678 9007 679 9011
rect 683 9007 684 9011
rect 688 9007 689 9011
rect 659 9006 693 9007
rect 2806 9006 2882 9010
rect 2886 9006 2913 9010
rect 2917 9006 2935 9010
rect 2939 9006 3000 9010
rect 3004 9006 3018 9010
rect 663 9002 664 9006
rect 668 9002 669 9006
rect 673 9002 674 9006
rect 678 9002 679 9006
rect 683 9002 684 9006
rect 688 9002 689 9006
rect 3054 9003 3057 9022
rect 3159 9003 3162 9022
rect 3390 9012 3393 9022
rect 3680 9017 3781 9021
rect 3817 9028 3820 9034
rect 3826 9036 3829 9042
rect 3842 9037 3845 9042
rect 3826 9032 3828 9036
rect 3832 9032 3834 9036
rect 3842 9035 3848 9037
rect 3852 9035 3853 9037
rect 3842 9033 3853 9035
rect 3870 9035 3873 9042
rect 3826 9028 3829 9032
rect 3842 9028 3845 9033
rect 3871 9031 3873 9035
rect 3870 9028 3873 9031
rect 3886 9036 3889 9042
rect 3896 9036 3899 9042
rect 3917 9037 3920 9042
rect 3896 9032 3905 9036
rect 3917 9033 3918 9037
rect 3922 9034 3925 9037
rect 3942 9036 3945 9042
rect 3960 9037 3963 9042
rect 3886 9028 3889 9032
rect 3896 9028 3899 9032
rect 3917 9028 3920 9033
rect 3944 9032 3945 9036
rect 3989 9033 3994 9038
rect 3998 9034 4000 9037
rect 4015 9036 4018 9042
rect 4015 9033 4023 9036
rect 4095 9033 4100 9038
rect 4104 9034 4105 9037
rect 4120 9036 4123 9042
rect 4479 9045 4513 9046
rect 4483 9041 4484 9045
rect 4488 9041 4489 9045
rect 4493 9041 4494 9045
rect 4498 9041 4499 9045
rect 4503 9041 4504 9045
rect 4508 9041 4509 9045
rect 4529 9056 4530 9060
rect 4534 9056 4535 9060
rect 4539 9056 4540 9060
rect 4544 9056 4545 9060
rect 4549 9056 4550 9060
rect 4554 9056 4555 9060
rect 4826 9059 5086 9062
rect 4525 9055 4559 9056
rect 4529 9051 4530 9055
rect 4534 9051 4535 9055
rect 4539 9051 4540 9055
rect 4544 9051 4545 9055
rect 4549 9051 4550 9055
rect 4554 9051 4555 9055
rect 4525 9050 4559 9051
rect 4529 9046 4530 9050
rect 4534 9046 4535 9050
rect 4539 9046 4540 9050
rect 4544 9046 4545 9050
rect 4549 9046 4550 9050
rect 4554 9046 4555 9050
rect 4525 9045 4559 9046
rect 4529 9041 4530 9045
rect 4534 9041 4535 9045
rect 4539 9041 4540 9045
rect 4544 9041 4545 9045
rect 4549 9041 4550 9045
rect 4554 9041 4555 9045
rect 4120 9033 4128 9036
rect 3942 9028 3945 9032
rect 3960 9028 3963 9033
rect 4015 9030 4018 9033
rect 4120 9030 4123 9033
rect 3870 9013 3873 9017
rect 3897 9013 3898 9017
rect 3942 9013 3944 9017
rect 3598 9008 3733 9012
rect 659 9001 693 9002
rect 663 8997 664 9001
rect 668 8997 669 9001
rect 673 8997 674 9001
rect 678 8997 679 9001
rect 683 8997 684 9001
rect 688 8997 689 9001
rect 2770 8999 2855 9003
rect 2859 8999 2871 9003
rect 2875 8999 2889 9003
rect 2893 8999 2900 9003
rect 2904 8999 2906 9003
rect 2910 8999 2925 9003
rect 2929 8999 2962 9003
rect 2966 8999 2967 9003
rect 2971 8999 2979 9003
rect 2983 8999 3007 9003
rect 3011 8999 3023 9003
rect 3027 8999 3047 9003
rect 3051 8999 3101 9003
rect 3105 8999 3128 9003
rect 3132 8999 3182 9003
rect 3186 8999 3190 9003
rect 3194 8999 3218 9003
rect 3222 8999 3272 9003
rect 3330 9000 3391 9003
rect 3406 9002 3409 9008
rect 3751 9006 3827 9010
rect 3831 9006 3858 9010
rect 3862 9006 3880 9010
rect 3884 9006 3945 9010
rect 3949 9006 3963 9010
rect 3999 9003 4002 9022
rect 4104 9003 4107 9022
rect 4826 9007 5086 9010
rect 3406 8999 3414 9002
rect 3715 8999 3800 9003
rect 3804 8999 3816 9003
rect 3820 8999 3834 9003
rect 3838 8999 3845 9003
rect 3849 8999 3851 9003
rect 3855 8999 3870 9003
rect 3874 8999 3907 9003
rect 3911 8999 3912 9003
rect 3916 8999 3924 9003
rect 3928 8999 3952 9003
rect 3956 8999 3968 9003
rect 3972 8999 3992 9003
rect 3996 8999 4046 9003
rect 4050 8999 4073 9003
rect 4077 8999 4127 9003
rect 4131 8999 4135 9003
rect 4139 8999 4163 9003
rect 4167 8999 4217 9003
rect 86 8741 89 8995
rect 343 8956 346 8995
rect 2806 8992 2882 8996
rect 2886 8992 2913 8996
rect 2917 8992 2935 8996
rect 2939 8992 3000 8996
rect 3004 8992 3018 8996
rect 3054 8989 3057 8999
rect 3084 8995 3087 8999
rect 3111 8995 3114 8999
rect 2925 8985 2928 8989
rect 2952 8985 2953 8989
rect 2997 8985 2999 8989
rect 2854 8965 2857 8968
rect 2865 8968 2868 8974
rect 2872 8968 2875 8974
rect 2865 8965 2875 8968
rect 2865 8960 2868 8965
rect 2872 8960 2875 8965
rect 2881 8970 2884 8974
rect 2881 8966 2883 8970
rect 2887 8966 2889 8970
rect 2897 8969 2900 8974
rect 2925 8971 2928 8974
rect 2897 8967 2908 8969
rect 2881 8960 2884 8966
rect 2897 8965 2903 8967
rect 2897 8960 2900 8965
rect 2907 8965 2908 8967
rect 2926 8967 2928 8971
rect 2925 8960 2928 8967
rect 3070 8978 3073 8981
rect 2941 8970 2944 8974
rect 2951 8970 2954 8974
rect 2951 8966 2960 8970
rect 2972 8969 2975 8974
rect 2997 8970 3000 8974
rect 2941 8960 2944 8966
rect 2951 8960 2954 8966
rect 2972 8965 2973 8969
rect 2977 8965 2980 8968
rect 2999 8966 3000 8970
rect 3015 8969 3018 8974
rect 3047 8974 3058 8977
rect 3070 8975 3078 8978
rect 2972 8960 2975 8965
rect 2997 8960 3000 8966
rect 3047 8968 3050 8974
rect 3070 8969 3073 8975
rect 3082 8970 3085 8973
rect 3093 8973 3096 8987
rect 3120 8982 3123 8987
rect 3135 8989 3138 8999
rect 3165 8995 3168 8999
rect 3201 8995 3204 8999
rect 3104 8978 3105 8981
rect 3109 8978 3112 8981
rect 3151 8978 3154 8981
rect 3093 8970 3101 8973
rect 3120 8973 3123 8978
rect 3015 8960 3018 8965
rect 3093 8965 3096 8970
rect 3101 8966 3105 8970
rect 3128 8974 3139 8977
rect 3151 8975 3159 8978
rect 3045 8959 3050 8964
rect 343 8946 356 8956
rect 2917 8947 2918 8951
rect 2942 8948 2943 8952
rect 2989 8947 2990 8951
rect 343 8936 366 8946
rect 2794 8940 2870 8944
rect 2874 8940 2929 8944
rect 2933 8940 2954 8944
rect 2958 8940 2985 8944
rect 2989 8940 3018 8944
rect 3054 8937 3057 8965
rect 3084 8937 3087 8961
rect 3111 8937 3114 8969
rect 3128 8968 3131 8974
rect 3151 8969 3154 8975
rect 3163 8970 3166 8973
rect 3174 8973 3177 8987
rect 3210 8982 3213 8987
rect 3225 8989 3228 8999
rect 3255 8995 3258 8999
rect 3406 8996 3409 8999
rect 3199 8978 3202 8981
rect 3241 8978 3244 8981
rect 3174 8970 3183 8973
rect 3210 8973 3213 8978
rect 3174 8965 3177 8970
rect 3126 8959 3131 8964
rect 3135 8937 3138 8965
rect 3217 8976 3229 8977
rect 3221 8974 3229 8976
rect 3241 8975 3249 8978
rect 3241 8969 3244 8975
rect 3253 8970 3256 8973
rect 3264 8973 3267 8987
rect 3751 8992 3827 8996
rect 3831 8992 3858 8996
rect 3862 8992 3880 8996
rect 3884 8992 3945 8996
rect 3949 8992 3963 8996
rect 3999 8989 4002 8999
rect 4029 8995 4032 8999
rect 4056 8995 4059 8999
rect 3390 8976 3393 8988
rect 3870 8985 3873 8989
rect 3897 8985 3898 8989
rect 3942 8985 3944 8989
rect 3264 8970 3284 8973
rect 3165 8937 3168 8961
rect 3201 8937 3204 8969
rect 3264 8965 3267 8970
rect 3341 8972 3359 8976
rect 3363 8972 3383 8976
rect 3387 8972 3437 8976
rect 3441 8972 3486 8976
rect 3490 8972 3668 8976
rect 3225 8937 3228 8965
rect 3344 8968 3347 8972
rect 3366 8968 3369 8972
rect 3255 8937 3258 8961
rect 3353 8955 3356 8960
rect 3375 8955 3378 8960
rect 3390 8962 3393 8972
rect 3420 8968 3423 8972
rect 3337 8951 3338 8954
rect 3342 8951 3345 8954
rect 3357 8951 3360 8955
rect 3364 8951 3367 8954
rect 3406 8951 3409 8954
rect 3353 8946 3356 8951
rect 3375 8946 3378 8951
rect 3383 8947 3394 8950
rect 3406 8948 3414 8951
rect 3406 8942 3409 8948
rect 3418 8943 3421 8946
rect 3429 8946 3432 8960
rect 3446 8965 3449 8972
rect 3499 8965 3502 8972
rect 3799 8965 3802 8968
rect 3810 8968 3813 8974
rect 3817 8968 3820 8974
rect 3810 8965 3820 8968
rect 3429 8943 3441 8946
rect 343 8926 376 8936
rect 2782 8933 2856 8937
rect 2860 8933 2862 8937
rect 2866 8933 2870 8937
rect 2874 8933 2888 8937
rect 2892 8933 2897 8937
rect 2901 8933 2906 8937
rect 2910 8933 2929 8937
rect 2933 8933 2963 8937
rect 2967 8933 2978 8937
rect 2982 8933 3006 8937
rect 3010 8933 3023 8937
rect 3027 8933 3047 8937
rect 3051 8933 3101 8937
rect 3108 8933 3128 8937
rect 3132 8933 3182 8937
rect 3186 8933 3218 8937
rect 3222 8933 3272 8937
rect 2794 8926 2870 8930
rect 2874 8926 2929 8930
rect 2933 8926 2954 8930
rect 2958 8926 2985 8930
rect 2989 8926 3018 8930
rect 343 8916 386 8926
rect 2917 8919 2918 8923
rect 2942 8918 2943 8922
rect 2989 8919 2990 8923
rect 343 8820 769 8916
rect 2865 8905 2868 8910
rect 2872 8905 2875 8910
rect 2855 8902 2857 8905
rect 2865 8902 2875 8905
rect 2865 8896 2868 8902
rect 2872 8896 2875 8902
rect 2881 8904 2884 8910
rect 2897 8905 2900 8910
rect 2881 8900 2883 8904
rect 2887 8900 2889 8904
rect 2897 8903 2903 8905
rect 2907 8903 2908 8905
rect 2897 8901 2908 8903
rect 2925 8903 2928 8910
rect 2881 8896 2884 8900
rect 2897 8896 2900 8901
rect 2926 8899 2928 8903
rect 2925 8896 2928 8899
rect 2941 8904 2944 8910
rect 2951 8904 2954 8910
rect 2972 8905 2975 8910
rect 2951 8900 2960 8904
rect 2972 8901 2973 8905
rect 2977 8902 2980 8905
rect 2997 8904 3000 8910
rect 3015 8905 3018 8910
rect 3054 8911 3057 8933
rect 3135 8911 3138 8933
rect 3225 8911 3228 8933
rect 2941 8896 2944 8900
rect 2951 8896 2954 8900
rect 2972 8896 2975 8901
rect 2999 8900 3000 8904
rect 2997 8896 3000 8900
rect 3015 8896 3018 8901
rect 3045 8898 3050 8903
rect 3054 8899 3055 8902
rect 3070 8901 3073 8907
rect 3070 8898 3078 8901
rect 3125 8898 3130 8903
rect 3134 8899 3136 8902
rect 3151 8901 3154 8907
rect 3151 8898 3159 8901
rect 3218 8899 3226 8902
rect 3241 8901 3244 8907
rect 3241 8898 3249 8901
rect 3070 8895 3073 8898
rect 3151 8895 3154 8898
rect 3241 8895 3244 8898
rect 3344 8896 3347 8942
rect 3366 8896 3369 8942
rect 3429 8938 3432 8943
rect 3390 8896 3393 8938
rect 3420 8896 3423 8934
rect 3438 8928 3441 8943
rect 3810 8960 3813 8965
rect 3817 8960 3820 8965
rect 3826 8970 3829 8974
rect 3826 8966 3828 8970
rect 3832 8966 3834 8970
rect 3842 8969 3845 8974
rect 3870 8971 3873 8974
rect 3842 8967 3853 8969
rect 3826 8960 3829 8966
rect 3842 8965 3848 8967
rect 3842 8960 3845 8965
rect 3852 8965 3853 8967
rect 3871 8967 3873 8971
rect 3870 8960 3873 8967
rect 4015 8978 4018 8981
rect 3886 8970 3889 8974
rect 3896 8970 3899 8974
rect 3896 8966 3905 8970
rect 3917 8969 3920 8974
rect 3942 8970 3945 8974
rect 3886 8960 3889 8966
rect 3896 8960 3899 8966
rect 3917 8965 3918 8969
rect 3922 8965 3925 8968
rect 3944 8966 3945 8970
rect 3960 8969 3963 8974
rect 3992 8974 4003 8977
rect 4015 8975 4023 8978
rect 3917 8960 3920 8965
rect 3942 8960 3945 8966
rect 3992 8968 3995 8974
rect 4015 8969 4018 8975
rect 4027 8970 4030 8973
rect 4038 8973 4041 8987
rect 4065 8982 4068 8987
rect 4080 8989 4083 8999
rect 4110 8995 4113 8999
rect 4146 8995 4149 8999
rect 4049 8978 4050 8981
rect 4054 8978 4057 8981
rect 4096 8978 4099 8981
rect 4038 8970 4046 8973
rect 4065 8973 4068 8978
rect 3960 8960 3963 8965
rect 4038 8965 4041 8970
rect 4046 8966 4050 8970
rect 4073 8974 4084 8977
rect 4096 8975 4104 8978
rect 3990 8959 3995 8964
rect 3862 8947 3863 8951
rect 3887 8948 3888 8952
rect 3934 8947 3935 8951
rect 3739 8940 3815 8944
rect 3819 8940 3874 8944
rect 3878 8940 3899 8944
rect 3903 8940 3930 8944
rect 3934 8940 3963 8944
rect 3999 8937 4002 8965
rect 4029 8937 4032 8961
rect 4056 8937 4059 8969
rect 4073 8968 4076 8974
rect 4096 8969 4099 8975
rect 4108 8970 4111 8973
rect 4119 8973 4122 8987
rect 4155 8982 4158 8987
rect 4170 8989 4173 8999
rect 4200 8995 4203 8999
rect 4144 8978 4147 8981
rect 4186 8978 4189 8981
rect 4119 8970 4128 8973
rect 4155 8973 4158 8978
rect 4119 8965 4122 8970
rect 4071 8959 4076 8964
rect 4080 8937 4083 8965
rect 4162 8976 4174 8977
rect 4166 8974 4174 8976
rect 4186 8975 4194 8978
rect 4186 8969 4189 8975
rect 4198 8970 4201 8973
rect 4209 8973 4212 8987
rect 4209 8970 4229 8973
rect 4110 8937 4113 8961
rect 4146 8937 4149 8969
rect 4209 8965 4212 8970
rect 4826 8968 4829 9007
rect 4170 8937 4173 8965
rect 4200 8937 4203 8961
rect 4816 8958 4829 8968
rect 4806 8948 4829 8958
rect 4796 8938 4829 8948
rect 3438 8923 3461 8928
rect 3479 8927 3482 8935
rect 3479 8923 3488 8927
rect 3492 8923 3514 8927
rect 3479 8915 3482 8923
rect 3532 8919 3535 8935
rect 3727 8933 3801 8937
rect 3805 8933 3807 8937
rect 3811 8933 3815 8937
rect 3819 8933 3833 8937
rect 3837 8933 3842 8937
rect 3846 8933 3851 8937
rect 3855 8933 3874 8937
rect 3878 8933 3908 8937
rect 3912 8933 3923 8937
rect 3927 8933 3951 8937
rect 3955 8933 3968 8937
rect 3972 8933 3992 8937
rect 3996 8933 4046 8937
rect 4053 8933 4073 8937
rect 4077 8933 4127 8937
rect 4131 8933 4163 8937
rect 4167 8933 4217 8937
rect 3739 8926 3815 8930
rect 3819 8926 3874 8930
rect 3878 8926 3899 8930
rect 3903 8926 3930 8930
rect 3934 8926 3963 8930
rect 3862 8919 3863 8923
rect 3887 8918 3888 8922
rect 3934 8919 3935 8923
rect 3536 8915 3769 8916
rect 3535 8912 3769 8915
rect 3446 8896 3449 8903
rect 3499 8896 3502 8903
rect 3810 8905 3813 8910
rect 3817 8905 3820 8910
rect 3800 8902 3802 8905
rect 3810 8902 3820 8905
rect 3810 8896 3813 8902
rect 2925 8881 2928 8885
rect 2952 8881 2953 8885
rect 2997 8881 2999 8885
rect 3341 8892 3359 8896
rect 3363 8892 3383 8896
rect 3387 8892 3437 8896
rect 3441 8892 3486 8896
rect 3490 8892 3660 8896
rect 2806 8874 2882 8878
rect 2886 8874 2913 8878
rect 2917 8874 2935 8878
rect 2939 8874 3000 8878
rect 3004 8874 3018 8878
rect 3054 8871 3057 8887
rect 3135 8871 3138 8887
rect 3225 8871 3228 8887
rect 3390 8882 3393 8892
rect 3817 8896 3820 8902
rect 3826 8904 3829 8910
rect 3842 8905 3845 8910
rect 3826 8900 3828 8904
rect 3832 8900 3834 8904
rect 3842 8903 3848 8905
rect 3852 8903 3853 8905
rect 3842 8901 3853 8903
rect 3870 8903 3873 8910
rect 3826 8896 3829 8900
rect 3842 8896 3845 8901
rect 3871 8899 3873 8903
rect 3870 8896 3873 8899
rect 3886 8904 3889 8910
rect 3896 8904 3899 8910
rect 3917 8905 3920 8910
rect 3896 8900 3905 8904
rect 3917 8901 3918 8905
rect 3922 8902 3925 8905
rect 3942 8904 3945 8910
rect 3960 8905 3963 8910
rect 3999 8911 4002 8933
rect 4080 8911 4083 8933
rect 4170 8911 4173 8933
rect 4786 8928 4829 8938
rect 3886 8896 3889 8900
rect 3896 8896 3899 8900
rect 3917 8896 3920 8901
rect 3944 8900 3945 8904
rect 3942 8896 3945 8900
rect 3960 8896 3963 8901
rect 3990 8898 3995 8903
rect 3999 8899 4000 8902
rect 4015 8901 4018 8907
rect 4015 8898 4023 8901
rect 4070 8898 4075 8903
rect 4079 8899 4081 8902
rect 4096 8901 4099 8907
rect 4096 8898 4104 8901
rect 4163 8899 4171 8902
rect 4186 8901 4189 8907
rect 4186 8898 4194 8901
rect 4015 8895 4018 8898
rect 4096 8895 4099 8898
rect 4186 8895 4189 8898
rect 3492 8882 3757 8886
rect 3870 8881 3873 8885
rect 3897 8881 3898 8885
rect 3942 8881 3944 8885
rect 2770 8867 2855 8871
rect 2859 8867 2871 8871
rect 2875 8867 2889 8871
rect 2893 8867 2900 8871
rect 2904 8867 2906 8871
rect 2910 8867 2925 8871
rect 2929 8867 2962 8871
rect 2966 8867 2967 8871
rect 2971 8867 2979 8871
rect 2983 8867 3007 8871
rect 3011 8867 3023 8871
rect 3027 8867 3047 8871
rect 3051 8867 3101 8871
rect 3105 8867 3128 8871
rect 3132 8867 3218 8871
rect 3222 8867 3276 8871
rect 3332 8870 3391 8873
rect 3406 8872 3409 8878
rect 3751 8874 3827 8878
rect 3831 8874 3858 8878
rect 3862 8874 3880 8878
rect 3884 8874 3945 8878
rect 3949 8874 3963 8878
rect 3406 8869 3414 8872
rect 3999 8871 4002 8887
rect 4080 8871 4083 8887
rect 4170 8871 4173 8887
rect 2806 8860 2882 8864
rect 2886 8860 2913 8864
rect 2917 8860 2935 8864
rect 2939 8860 3000 8864
rect 3004 8860 3018 8864
rect 3054 8857 3057 8867
rect 3084 8863 3087 8867
rect 3406 8866 3409 8869
rect 3715 8867 3800 8871
rect 3804 8867 3816 8871
rect 3820 8867 3834 8871
rect 3838 8867 3845 8871
rect 3849 8867 3851 8871
rect 3855 8867 3870 8871
rect 3874 8867 3907 8871
rect 3911 8867 3912 8871
rect 3916 8867 3924 8871
rect 3928 8867 3952 8871
rect 3956 8867 3968 8871
rect 3972 8867 3992 8871
rect 3996 8867 4046 8871
rect 4050 8867 4073 8871
rect 4077 8867 4163 8871
rect 4167 8867 4221 8871
rect 2925 8853 2928 8857
rect 2952 8853 2953 8857
rect 2997 8853 2999 8857
rect 2854 8833 2857 8836
rect 2865 8836 2868 8842
rect 2872 8836 2875 8842
rect 2865 8833 2875 8836
rect 2865 8828 2868 8833
rect 2872 8828 2875 8833
rect 2881 8838 2884 8842
rect 2881 8834 2883 8838
rect 2887 8834 2889 8838
rect 2897 8837 2900 8842
rect 2925 8839 2928 8842
rect 2897 8835 2908 8837
rect 2881 8828 2884 8834
rect 2897 8833 2903 8835
rect 2897 8828 2900 8833
rect 2907 8833 2908 8835
rect 2926 8835 2928 8839
rect 2925 8828 2928 8835
rect 3070 8846 3073 8849
rect 2941 8838 2944 8842
rect 2951 8838 2954 8842
rect 2951 8834 2960 8838
rect 2972 8837 2975 8842
rect 2997 8838 3000 8842
rect 2941 8828 2944 8834
rect 2951 8828 2954 8834
rect 2972 8833 2973 8837
rect 2977 8833 2980 8836
rect 2999 8834 3000 8838
rect 3015 8837 3018 8842
rect 3047 8842 3058 8845
rect 3070 8843 3078 8846
rect 2972 8828 2975 8833
rect 2997 8828 3000 8834
rect 3047 8836 3050 8842
rect 3070 8837 3073 8843
rect 3082 8838 3085 8841
rect 3093 8841 3096 8855
rect 3751 8860 3827 8864
rect 3831 8860 3858 8864
rect 3862 8860 3880 8864
rect 3884 8860 3945 8864
rect 3949 8860 3963 8864
rect 3390 8846 3393 8858
rect 3999 8857 4002 8867
rect 4029 8863 4032 8867
rect 3870 8853 3873 8857
rect 3897 8853 3898 8857
rect 3942 8853 3944 8857
rect 3101 8841 3106 8846
rect 3359 8842 3383 8846
rect 3387 8842 3668 8846
rect 3093 8838 3101 8841
rect 3015 8828 3018 8833
rect 3093 8833 3096 8838
rect 3799 8833 3802 8836
rect 3810 8836 3813 8842
rect 3817 8836 3820 8842
rect 3810 8833 3820 8836
rect 3045 8827 3050 8832
rect 343 8810 386 8820
rect 2355 8819 2476 8823
rect 2364 8812 2373 8816
rect 2377 8812 2409 8816
rect 2413 8812 2476 8816
rect 2480 8812 2505 8816
rect 2509 8812 2541 8816
rect 2545 8812 2608 8816
rect 2612 8812 2637 8816
rect 2641 8812 2673 8816
rect 2677 8812 2740 8816
rect 2744 8812 2824 8816
rect 2917 8815 2918 8819
rect 2942 8816 2943 8820
rect 2989 8815 2990 8819
rect 343 8800 376 8810
rect 2364 8805 2397 8809
rect 2401 8805 2425 8809
rect 2429 8805 2455 8809
rect 2459 8805 2492 8809
rect 2496 8805 2529 8809
rect 2533 8805 2557 8809
rect 2561 8805 2587 8809
rect 2591 8805 2624 8809
rect 2628 8805 2661 8809
rect 2665 8805 2689 8809
rect 2693 8805 2719 8809
rect 2723 8805 2756 8809
rect 2760 8805 2764 8809
rect 2849 8808 2870 8812
rect 2874 8808 2879 8812
rect 2883 8808 2929 8812
rect 2933 8808 2954 8812
rect 2958 8808 2985 8812
rect 2989 8808 3018 8812
rect 3054 8805 3057 8833
rect 3084 8805 3087 8829
rect 3810 8828 3813 8833
rect 3817 8828 3820 8833
rect 3826 8838 3829 8842
rect 3826 8834 3828 8838
rect 3832 8834 3834 8838
rect 3842 8837 3845 8842
rect 3870 8839 3873 8842
rect 3842 8835 3853 8837
rect 3826 8828 3829 8834
rect 3842 8833 3848 8835
rect 3842 8828 3845 8833
rect 3852 8833 3853 8835
rect 3871 8835 3873 8839
rect 3870 8828 3873 8835
rect 4015 8846 4018 8849
rect 3886 8838 3889 8842
rect 3896 8838 3899 8842
rect 3896 8834 3905 8838
rect 3917 8837 3920 8842
rect 3942 8838 3945 8842
rect 3886 8828 3889 8834
rect 3896 8828 3899 8834
rect 3917 8833 3918 8837
rect 3922 8833 3925 8836
rect 3944 8834 3945 8838
rect 3960 8837 3963 8842
rect 3992 8842 4003 8845
rect 4015 8843 4023 8846
rect 3917 8828 3920 8833
rect 3942 8828 3945 8834
rect 3992 8836 3995 8842
rect 4015 8837 4018 8843
rect 4027 8838 4030 8841
rect 4038 8841 4041 8855
rect 4046 8841 4051 8846
rect 4038 8838 4046 8841
rect 3960 8828 3963 8833
rect 4038 8833 4041 8838
rect 3990 8827 3995 8832
rect 3309 8812 3318 8816
rect 3322 8812 3354 8816
rect 3358 8812 3421 8816
rect 3425 8812 3450 8816
rect 3454 8812 3486 8816
rect 3490 8812 3553 8816
rect 3557 8812 3582 8816
rect 3586 8812 3618 8816
rect 3622 8812 3685 8816
rect 3689 8812 3769 8816
rect 3862 8815 3863 8819
rect 3887 8816 3888 8820
rect 3934 8815 3935 8819
rect 3309 8805 3342 8809
rect 3346 8805 3370 8809
rect 3374 8805 3400 8809
rect 3404 8805 3437 8809
rect 3441 8805 3474 8809
rect 3478 8805 3502 8809
rect 3506 8805 3532 8809
rect 3536 8805 3569 8809
rect 3573 8805 3606 8809
rect 3610 8805 3634 8809
rect 3638 8805 3664 8809
rect 3668 8805 3701 8809
rect 3705 8805 3709 8809
rect 3794 8808 3815 8812
rect 3819 8808 3824 8812
rect 3828 8808 3874 8812
rect 3878 8808 3899 8812
rect 3903 8808 3930 8812
rect 3934 8808 3963 8812
rect 3999 8805 4002 8833
rect 4403 8832 4829 8928
rect 4029 8805 4032 8829
rect 4786 8822 4829 8832
rect 4796 8812 4829 8822
rect 343 8790 366 8800
rect 2367 8795 2370 8805
rect 2388 8795 2391 8805
rect 2404 8795 2407 8805
rect 2418 8798 2423 8802
rect 2427 8798 2434 8802
rect 2446 8795 2449 8805
rect 2462 8795 2465 8805
rect 2483 8795 2486 8805
rect 2499 8795 2502 8805
rect 2520 8795 2523 8805
rect 2536 8795 2539 8805
rect 2550 8798 2555 8802
rect 2559 8798 2566 8802
rect 2578 8795 2581 8805
rect 2594 8795 2597 8805
rect 2615 8795 2618 8805
rect 2631 8795 2634 8805
rect 2652 8795 2655 8805
rect 2668 8795 2671 8805
rect 2682 8798 2687 8802
rect 2691 8798 2698 8802
rect 2710 8795 2713 8805
rect 2726 8795 2729 8805
rect 2747 8795 2750 8805
rect 2782 8801 2856 8805
rect 2860 8801 2862 8805
rect 2866 8801 2870 8805
rect 2874 8801 2888 8805
rect 2892 8801 2897 8805
rect 2901 8801 2906 8805
rect 2910 8801 2929 8805
rect 2933 8801 2963 8805
rect 2967 8801 2978 8805
rect 2982 8801 3006 8805
rect 3010 8801 3023 8805
rect 3027 8801 3047 8805
rect 3051 8801 3131 8805
rect 3135 8801 3149 8805
rect 3153 8801 3158 8805
rect 3162 8801 3167 8805
rect 3171 8801 3190 8805
rect 3194 8801 3224 8805
rect 3228 8801 3239 8805
rect 3243 8801 3267 8805
rect 3271 8801 3280 8805
rect 343 8780 356 8790
rect 343 8741 346 8780
rect 2355 8778 2371 8782
rect 2384 8781 2389 8784
rect 2393 8781 2417 8784
rect 2442 8781 2449 8784
rect 2453 8781 2475 8784
rect 2495 8781 2502 8784
rect 2516 8781 2521 8784
rect 2525 8781 2549 8784
rect 2574 8781 2581 8784
rect 2585 8781 2607 8784
rect 2627 8781 2634 8784
rect 2648 8781 2653 8784
rect 2657 8781 2681 8784
rect 2794 8794 2870 8798
rect 2874 8794 2879 8798
rect 2883 8794 2929 8798
rect 2933 8794 2954 8798
rect 2958 8794 2985 8798
rect 2989 8794 3018 8798
rect 2706 8781 2713 8784
rect 2717 8781 2739 8784
rect 2917 8787 2918 8791
rect 2942 8786 2943 8790
rect 2989 8787 2990 8791
rect 2400 8771 2407 8774
rect 2411 8775 2430 8778
rect 2430 8768 2433 8774
rect 2458 8771 2465 8774
rect 2469 8775 2484 8778
rect 2532 8771 2539 8774
rect 2543 8775 2562 8778
rect 2562 8768 2565 8774
rect 2590 8771 2597 8774
rect 2601 8775 2616 8778
rect 2664 8771 2671 8774
rect 2675 8775 2694 8778
rect 2694 8768 2697 8774
rect 2722 8771 2729 8774
rect 2733 8775 2750 8778
rect 2865 8773 2868 8778
rect 2872 8773 2875 8778
rect 2855 8770 2857 8773
rect 2865 8770 2875 8773
rect 2865 8764 2868 8770
rect 2367 8752 2370 8764
rect 2388 8752 2391 8764
rect 2404 8752 2407 8764
rect 2418 8755 2430 8758
rect 2446 8752 2449 8764
rect 2462 8752 2465 8764
rect 2483 8752 2486 8764
rect 2499 8752 2502 8764
rect 2520 8752 2523 8764
rect 2536 8752 2539 8764
rect 2550 8755 2562 8758
rect 2578 8752 2581 8764
rect 2594 8752 2597 8764
rect 2615 8752 2618 8764
rect 2631 8752 2634 8764
rect 2652 8752 2655 8764
rect 2668 8752 2671 8764
rect 2682 8755 2694 8758
rect 2710 8752 2713 8764
rect 2726 8752 2729 8764
rect 2747 8752 2750 8764
rect 2872 8764 2875 8770
rect 2881 8772 2884 8778
rect 2897 8773 2900 8778
rect 2881 8768 2883 8772
rect 2887 8768 2889 8772
rect 2897 8771 2903 8773
rect 2907 8771 2908 8773
rect 2897 8769 2908 8771
rect 2925 8771 2928 8778
rect 2881 8764 2884 8768
rect 2897 8764 2900 8769
rect 2926 8767 2928 8771
rect 2925 8764 2928 8767
rect 2941 8772 2944 8778
rect 2951 8772 2954 8778
rect 2972 8773 2975 8778
rect 2951 8768 2960 8772
rect 2972 8769 2973 8773
rect 2977 8770 2980 8773
rect 2997 8772 3000 8778
rect 3015 8773 3018 8778
rect 3054 8775 3057 8801
rect 3090 8794 3109 8798
rect 3113 8794 3131 8798
rect 3135 8794 3190 8798
rect 3194 8794 3215 8798
rect 3219 8794 3246 8798
rect 3250 8794 3279 8798
rect 3312 8795 3315 8805
rect 3333 8795 3336 8805
rect 3349 8795 3352 8805
rect 3363 8798 3368 8802
rect 3372 8798 3379 8802
rect 3391 8795 3394 8805
rect 3407 8795 3410 8805
rect 3428 8795 3431 8805
rect 3444 8795 3447 8805
rect 3465 8795 3468 8805
rect 3481 8795 3484 8805
rect 3495 8798 3500 8802
rect 3504 8798 3511 8802
rect 3523 8795 3526 8805
rect 3539 8795 3542 8805
rect 3560 8795 3563 8805
rect 3576 8795 3579 8805
rect 3597 8795 3600 8805
rect 3613 8795 3616 8805
rect 3627 8798 3632 8802
rect 3636 8798 3643 8802
rect 3655 8795 3658 8805
rect 3671 8795 3674 8805
rect 3692 8795 3695 8805
rect 3727 8801 3801 8805
rect 3805 8801 3807 8805
rect 3811 8801 3815 8805
rect 3819 8801 3833 8805
rect 3837 8801 3842 8805
rect 3846 8801 3851 8805
rect 3855 8801 3874 8805
rect 3878 8801 3908 8805
rect 3912 8801 3923 8805
rect 3927 8801 3951 8805
rect 3955 8801 3968 8805
rect 3972 8801 3992 8805
rect 3996 8801 4076 8805
rect 4080 8801 4094 8805
rect 4098 8801 4103 8805
rect 4107 8801 4112 8805
rect 4116 8801 4135 8805
rect 4139 8801 4169 8805
rect 4173 8801 4184 8805
rect 4188 8801 4212 8805
rect 4216 8801 4225 8805
rect 4806 8802 4829 8812
rect 3090 8782 3093 8794
rect 3178 8787 3179 8791
rect 3203 8786 3204 8790
rect 3250 8787 3251 8791
rect 2941 8764 2944 8768
rect 2951 8764 2954 8768
rect 2972 8764 2975 8769
rect 2999 8768 3000 8772
rect 3117 8773 3120 8778
rect 3126 8773 3129 8778
rect 3133 8773 3136 8778
rect 2997 8764 3000 8768
rect 3015 8764 3018 8769
rect 3044 8762 3049 8767
rect 3053 8763 3055 8766
rect 3070 8765 3073 8771
rect 3102 8770 3136 8773
rect 3070 8762 3078 8765
rect 3070 8759 3073 8762
rect 2364 8748 2397 8752
rect 2401 8748 2425 8752
rect 2429 8748 2455 8752
rect 2459 8748 2529 8752
rect 2533 8748 2557 8752
rect 2561 8748 2587 8752
rect 2591 8748 2661 8752
rect 2665 8748 2689 8752
rect 2693 8748 2719 8752
rect 2723 8748 2776 8752
rect 2925 8749 2928 8753
rect 2952 8749 2953 8753
rect 2997 8749 2999 8753
rect 3102 8756 3105 8770
rect 3126 8764 3129 8770
rect 3133 8764 3136 8770
rect 3142 8772 3145 8778
rect 3158 8773 3161 8778
rect 3142 8768 3144 8772
rect 3148 8768 3150 8772
rect 3158 8771 3164 8773
rect 3168 8771 3169 8773
rect 3158 8769 3169 8771
rect 3186 8771 3189 8778
rect 3142 8764 3145 8768
rect 3158 8764 3161 8769
rect 3187 8767 3189 8771
rect 3186 8764 3189 8767
rect 3329 8781 3334 8784
rect 3338 8781 3362 8784
rect 3387 8781 3394 8784
rect 3398 8781 3420 8784
rect 3440 8781 3447 8784
rect 3461 8781 3466 8784
rect 3470 8781 3494 8784
rect 3519 8781 3526 8784
rect 3530 8781 3552 8784
rect 3572 8781 3579 8784
rect 3593 8781 3598 8784
rect 3602 8781 3626 8784
rect 3739 8794 3815 8798
rect 3819 8794 3824 8798
rect 3828 8794 3874 8798
rect 3878 8794 3899 8798
rect 3903 8794 3930 8798
rect 3934 8794 3963 8798
rect 3651 8781 3658 8784
rect 3662 8781 3684 8784
rect 3862 8787 3863 8791
rect 3887 8786 3888 8790
rect 3934 8787 3935 8791
rect 3202 8772 3205 8778
rect 3212 8772 3215 8778
rect 3233 8773 3236 8778
rect 3212 8768 3221 8772
rect 3233 8769 3234 8773
rect 3238 8770 3241 8773
rect 3258 8772 3261 8778
rect 3276 8773 3279 8778
rect 3202 8764 3205 8768
rect 3212 8764 3215 8768
rect 3233 8764 3236 8769
rect 3260 8768 3261 8772
rect 3258 8764 3261 8768
rect 3276 8764 3279 8769
rect 3345 8771 3352 8774
rect 3356 8775 3375 8778
rect 3375 8768 3378 8774
rect 3403 8771 3410 8774
rect 3414 8775 3429 8778
rect 3477 8771 3484 8774
rect 3488 8775 3507 8778
rect 3507 8768 3510 8774
rect 3535 8771 3542 8774
rect 3546 8775 3561 8778
rect 3609 8771 3616 8774
rect 3620 8775 3639 8778
rect 3639 8768 3642 8774
rect 3667 8771 3674 8774
rect 3678 8775 3695 8778
rect 3810 8773 3813 8778
rect 3817 8773 3820 8778
rect 3800 8770 3802 8773
rect 3810 8770 3820 8773
rect 3810 8764 3813 8770
rect 2364 8741 2373 8745
rect 2377 8741 2424 8745
rect 2428 8741 2474 8745
rect 2478 8741 2505 8745
rect 2509 8741 2556 8745
rect 2560 8741 2606 8745
rect 2610 8741 2637 8745
rect 2641 8741 2688 8745
rect 2692 8741 2738 8745
rect 2742 8742 2812 8745
rect 2868 8742 2882 8746
rect 2886 8742 2913 8746
rect 2917 8742 2935 8746
rect 2939 8742 3000 8746
rect 3004 8742 3018 8746
rect 86 8738 346 8741
rect 3054 8739 3057 8751
rect 3186 8749 3189 8753
rect 3213 8749 3214 8753
rect 3258 8749 3260 8753
rect 3312 8752 3315 8764
rect 3333 8752 3336 8764
rect 3349 8752 3352 8764
rect 3363 8755 3375 8758
rect 3391 8752 3394 8764
rect 3407 8752 3410 8764
rect 3428 8752 3431 8764
rect 3444 8752 3447 8764
rect 3465 8752 3468 8764
rect 3481 8752 3484 8764
rect 3495 8755 3507 8758
rect 3523 8752 3526 8764
rect 3539 8752 3542 8764
rect 3560 8752 3563 8764
rect 3576 8752 3579 8764
rect 3597 8752 3600 8764
rect 3613 8752 3616 8764
rect 3627 8755 3639 8758
rect 3655 8752 3658 8764
rect 3671 8752 3674 8764
rect 3692 8752 3695 8764
rect 3817 8764 3820 8770
rect 3826 8772 3829 8778
rect 3842 8773 3845 8778
rect 3826 8768 3828 8772
rect 3832 8768 3834 8772
rect 3842 8771 3848 8773
rect 3852 8771 3853 8773
rect 3842 8769 3853 8771
rect 3870 8771 3873 8778
rect 3826 8764 3829 8768
rect 3842 8764 3845 8769
rect 3871 8767 3873 8771
rect 3870 8764 3873 8767
rect 3886 8772 3889 8778
rect 3896 8772 3899 8778
rect 3917 8773 3920 8778
rect 3896 8768 3905 8772
rect 3917 8769 3918 8773
rect 3922 8770 3925 8773
rect 3942 8772 3945 8778
rect 3960 8773 3963 8778
rect 3999 8775 4002 8801
rect 4035 8794 4054 8798
rect 4058 8794 4076 8798
rect 4080 8794 4135 8798
rect 4139 8794 4160 8798
rect 4164 8794 4191 8798
rect 4195 8794 4224 8798
rect 4035 8782 4038 8794
rect 4816 8792 4829 8802
rect 4123 8787 4124 8791
rect 4148 8786 4149 8790
rect 4195 8787 4196 8791
rect 3886 8764 3889 8768
rect 3896 8764 3899 8768
rect 3917 8764 3920 8769
rect 3944 8768 3945 8772
rect 4062 8773 4065 8778
rect 4071 8773 4074 8778
rect 4078 8773 4081 8778
rect 3942 8764 3945 8768
rect 3960 8764 3963 8769
rect 3989 8762 3994 8767
rect 3998 8763 4000 8766
rect 4015 8765 4018 8771
rect 4047 8770 4081 8773
rect 4015 8762 4023 8765
rect 4015 8759 4018 8762
rect 3309 8748 3342 8752
rect 3346 8748 3370 8752
rect 3374 8748 3400 8752
rect 3404 8748 3474 8752
rect 3478 8748 3502 8752
rect 3506 8748 3532 8752
rect 3536 8748 3606 8752
rect 3610 8748 3634 8752
rect 3638 8748 3664 8752
rect 3668 8748 3721 8752
rect 3870 8749 3873 8753
rect 3897 8749 3898 8753
rect 3942 8749 3944 8753
rect 4047 8756 4050 8770
rect 4071 8764 4074 8770
rect 4078 8764 4081 8770
rect 4087 8772 4090 8778
rect 4103 8773 4106 8778
rect 4087 8768 4089 8772
rect 4093 8768 4095 8772
rect 4103 8771 4109 8773
rect 4113 8771 4114 8773
rect 4103 8769 4114 8771
rect 4131 8771 4134 8778
rect 4087 8764 4090 8768
rect 4103 8764 4106 8769
rect 4132 8767 4134 8771
rect 4131 8764 4134 8767
rect 4147 8772 4150 8778
rect 4157 8772 4160 8778
rect 4178 8773 4181 8778
rect 4157 8768 4166 8772
rect 4178 8769 4179 8773
rect 4183 8770 4186 8773
rect 4203 8772 4206 8778
rect 4221 8773 4224 8778
rect 4147 8764 4150 8768
rect 4157 8764 4160 8768
rect 4178 8764 4181 8769
rect 4205 8768 4206 8772
rect 4203 8764 4206 8768
rect 4221 8764 4224 8769
rect 3094 8742 3099 8746
rect 3103 8742 3143 8746
rect 3147 8742 3174 8746
rect 3178 8742 3196 8746
rect 3200 8742 3261 8746
rect 3265 8742 3279 8746
rect 3309 8741 3318 8745
rect 3322 8741 3369 8745
rect 3373 8741 3419 8745
rect 3423 8741 3450 8745
rect 3454 8741 3501 8745
rect 3505 8741 3551 8745
rect 3555 8741 3582 8745
rect 3586 8741 3633 8745
rect 3637 8741 3683 8745
rect 3687 8742 3757 8745
rect 3813 8742 3827 8746
rect 3831 8742 3858 8746
rect 3862 8742 3880 8746
rect 3884 8742 3945 8746
rect 3949 8742 3963 8746
rect 3999 8739 4002 8751
rect 4131 8749 4134 8753
rect 4158 8749 4159 8753
rect 4203 8749 4205 8753
rect 4826 8753 4829 8792
rect 5083 8753 5086 9007
rect 4483 8747 4484 8751
rect 4488 8747 4489 8751
rect 4493 8747 4494 8751
rect 4498 8747 4499 8751
rect 4503 8747 4504 8751
rect 4508 8747 4509 8751
rect 4479 8746 4513 8747
rect 4039 8742 4044 8746
rect 4048 8742 4088 8746
rect 4092 8742 4119 8746
rect 4123 8742 4141 8746
rect 4145 8742 4206 8746
rect 4210 8742 4224 8746
rect 4483 8742 4484 8746
rect 4488 8742 4489 8746
rect 4493 8742 4494 8746
rect 4498 8742 4499 8746
rect 4503 8742 4504 8746
rect 4508 8742 4509 8746
rect 4479 8741 4513 8742
rect 2371 8735 2755 8738
rect 2770 8735 2855 8739
rect 2859 8735 2871 8739
rect 2875 8735 2889 8739
rect 2893 8735 2900 8739
rect 2904 8735 2906 8739
rect 2910 8735 2925 8739
rect 2929 8735 2962 8739
rect 2966 8735 2967 8739
rect 2971 8735 2979 8739
rect 2983 8735 3007 8739
rect 3011 8735 3047 8739
rect 3051 8735 3090 8739
rect 3094 8735 3101 8739
rect 3105 8735 3116 8739
rect 3120 8735 3132 8739
rect 3136 8735 3150 8739
rect 3154 8735 3161 8739
rect 3165 8735 3167 8739
rect 3171 8735 3186 8739
rect 3190 8735 3223 8739
rect 3227 8735 3228 8739
rect 3232 8735 3240 8739
rect 3244 8735 3268 8739
rect 3272 8735 3280 8739
rect 3316 8735 3700 8738
rect 3715 8735 3800 8739
rect 3804 8735 3816 8739
rect 3820 8735 3834 8739
rect 3838 8735 3845 8739
rect 3849 8735 3851 8739
rect 3855 8735 3870 8739
rect 3874 8735 3907 8739
rect 3911 8735 3912 8739
rect 3916 8735 3924 8739
rect 3928 8735 3952 8739
rect 3956 8735 3992 8739
rect 3996 8735 4035 8739
rect 4039 8735 4046 8739
rect 4050 8735 4061 8739
rect 4065 8735 4077 8739
rect 4081 8735 4095 8739
rect 4099 8735 4106 8739
rect 4110 8735 4112 8739
rect 4116 8735 4131 8739
rect 4135 8735 4168 8739
rect 4172 8735 4173 8739
rect 4177 8735 4185 8739
rect 4189 8735 4213 8739
rect 4217 8735 4225 8739
rect 4483 8737 4484 8741
rect 4488 8737 4489 8741
rect 4493 8737 4494 8741
rect 4498 8737 4499 8741
rect 4503 8737 4504 8741
rect 4508 8737 4509 8741
rect 4479 8736 4513 8737
rect 2514 8728 2623 8731
rect 2806 8728 2864 8732
rect 2868 8728 3098 8731
rect 3288 8729 3296 8733
rect 3459 8728 3568 8731
rect 3751 8728 3809 8732
rect 3813 8728 4043 8731
rect 4233 8729 4241 8733
rect 4483 8732 4484 8736
rect 4488 8732 4489 8736
rect 4493 8732 4494 8736
rect 4498 8732 4499 8736
rect 4503 8732 4504 8736
rect 4508 8732 4509 8736
rect 4529 8747 4530 8751
rect 4534 8747 4535 8751
rect 4539 8747 4540 8751
rect 4544 8747 4545 8751
rect 4549 8747 4550 8751
rect 4554 8747 4555 8751
rect 4826 8750 5086 8753
rect 4525 8746 4559 8747
rect 4529 8742 4530 8746
rect 4534 8742 4535 8746
rect 4539 8742 4540 8746
rect 4544 8742 4545 8746
rect 4549 8742 4550 8746
rect 4554 8742 4555 8746
rect 4525 8741 4559 8742
rect 4529 8737 4530 8741
rect 4534 8737 4535 8741
rect 4539 8737 4540 8741
rect 4544 8737 4545 8741
rect 4549 8737 4550 8741
rect 4554 8737 4555 8741
rect 4525 8736 4559 8737
rect 4529 8732 4530 8736
rect 4534 8732 4535 8736
rect 4539 8732 4540 8736
rect 4544 8732 4545 8736
rect 4549 8732 4550 8736
rect 4554 8732 4555 8736
rect 2494 8720 2498 8724
rect 2502 8720 2506 8724
rect 2794 8721 3108 8724
rect 2482 8719 2486 8720
rect 2514 8719 2518 8720
rect 2842 8714 3115 8717
rect 3284 8711 3288 8716
rect 3439 8720 3443 8724
rect 3447 8720 3451 8724
rect 3739 8721 4053 8724
rect 3427 8719 3431 8720
rect 3459 8719 3463 8720
rect 3787 8714 4058 8718
rect 4229 8711 4233 8716
rect 2355 8707 2482 8711
rect 2486 8707 2502 8711
rect 2518 8707 3427 8711
rect 3431 8707 3447 8711
rect 3463 8707 4321 8711
rect 617 8703 618 8707
rect 622 8703 623 8707
rect 627 8703 628 8707
rect 632 8703 633 8707
rect 637 8703 638 8707
rect 642 8703 643 8707
rect 613 8702 647 8703
rect 617 8698 618 8702
rect 622 8698 623 8702
rect 627 8698 628 8702
rect 632 8698 633 8702
rect 637 8698 638 8702
rect 642 8698 643 8702
rect 613 8697 647 8698
rect 617 8693 618 8697
rect 622 8693 623 8697
rect 627 8693 628 8697
rect 632 8693 633 8697
rect 637 8693 638 8697
rect 642 8693 643 8697
rect 613 8692 647 8693
rect 86 8686 346 8689
rect 617 8688 618 8692
rect 622 8688 623 8692
rect 627 8688 628 8692
rect 632 8688 633 8692
rect 637 8688 638 8692
rect 642 8688 643 8692
rect 663 8703 664 8707
rect 668 8703 669 8707
rect 673 8703 674 8707
rect 678 8703 679 8707
rect 683 8703 684 8707
rect 688 8703 689 8707
rect 659 8702 693 8703
rect 663 8698 664 8702
rect 668 8698 669 8702
rect 673 8698 674 8702
rect 678 8698 679 8702
rect 683 8698 684 8702
rect 688 8698 689 8702
rect 659 8697 693 8698
rect 663 8693 664 8697
rect 668 8693 669 8697
rect 673 8693 674 8697
rect 678 8693 679 8697
rect 683 8693 684 8697
rect 688 8693 689 8697
rect 2510 8700 2755 8703
rect 2830 8700 3156 8704
rect 3160 8700 3192 8704
rect 3196 8700 3259 8704
rect 3263 8700 3279 8704
rect 3455 8700 3700 8703
rect 3775 8700 4101 8704
rect 4105 8700 4137 8704
rect 4141 8700 4204 8704
rect 4208 8700 4224 8704
rect 659 8692 693 8693
rect 2525 8693 2755 8696
rect 2770 8693 3142 8697
rect 3146 8693 3180 8697
rect 3184 8693 3208 8697
rect 3212 8693 3238 8697
rect 3242 8693 3275 8697
rect 4826 8698 5086 8701
rect 663 8688 664 8692
rect 668 8688 669 8692
rect 673 8688 674 8692
rect 678 8688 679 8692
rect 683 8688 684 8692
rect 688 8688 689 8692
rect 86 8432 89 8686
rect 343 8647 346 8686
rect 2494 8684 2498 8688
rect 2502 8684 2506 8688
rect 3150 8683 3153 8693
rect 3171 8683 3174 8693
rect 3187 8683 3190 8693
rect 3201 8686 3206 8690
rect 3210 8686 3217 8690
rect 3229 8683 3232 8693
rect 3245 8683 3248 8693
rect 3266 8683 3269 8693
rect 3470 8693 3700 8696
rect 3715 8693 4087 8697
rect 4091 8693 4125 8697
rect 4129 8693 4153 8697
rect 4157 8693 4183 8697
rect 4187 8693 4220 8697
rect 3439 8684 3443 8688
rect 3447 8684 3451 8688
rect 4095 8683 4098 8693
rect 4116 8683 4119 8693
rect 4132 8683 4135 8693
rect 4146 8686 4151 8690
rect 4155 8686 4162 8690
rect 4174 8683 4177 8693
rect 4190 8683 4193 8693
rect 4211 8683 4214 8693
rect 2514 8677 2624 8680
rect 2364 8670 2373 8674
rect 2377 8670 2409 8674
rect 2413 8670 2476 8674
rect 2480 8670 2505 8674
rect 2509 8670 2541 8674
rect 2545 8670 2608 8674
rect 2612 8670 2637 8674
rect 2641 8670 2673 8674
rect 2677 8670 2740 8674
rect 2744 8670 2824 8674
rect 2364 8663 2397 8667
rect 2401 8663 2425 8667
rect 2429 8663 2455 8667
rect 2459 8663 2492 8667
rect 2496 8663 2529 8667
rect 2533 8663 2557 8667
rect 2561 8663 2587 8667
rect 2591 8663 2624 8667
rect 2628 8663 2661 8667
rect 2665 8663 2689 8667
rect 2693 8663 2719 8667
rect 2723 8663 2756 8667
rect 2760 8663 2764 8667
rect 3167 8669 3172 8672
rect 3176 8669 3200 8672
rect 3459 8677 3569 8680
rect 3225 8669 3232 8672
rect 3236 8669 3258 8672
rect 3309 8670 3318 8674
rect 3322 8670 3354 8674
rect 3358 8670 3421 8674
rect 3425 8670 3450 8674
rect 3454 8670 3486 8674
rect 3490 8670 3553 8674
rect 3557 8670 3582 8674
rect 3586 8670 3618 8674
rect 3622 8670 3685 8674
rect 3689 8670 3769 8674
rect 2367 8653 2370 8663
rect 2388 8653 2391 8663
rect 2404 8653 2407 8663
rect 2418 8656 2423 8660
rect 2427 8656 2434 8660
rect 2446 8653 2449 8663
rect 2462 8653 2465 8663
rect 2483 8653 2486 8663
rect 2499 8653 2502 8663
rect 2520 8653 2523 8663
rect 2536 8653 2539 8663
rect 2550 8656 2555 8660
rect 2559 8656 2566 8660
rect 2578 8653 2581 8663
rect 2594 8653 2597 8663
rect 2615 8653 2618 8663
rect 2631 8653 2634 8663
rect 2652 8653 2655 8663
rect 2668 8653 2671 8663
rect 2682 8656 2687 8660
rect 2691 8656 2698 8660
rect 2710 8653 2713 8663
rect 2726 8653 2729 8663
rect 2747 8653 2750 8663
rect 3183 8659 3190 8662
rect 3194 8663 3213 8666
rect 343 8637 356 8647
rect 343 8627 366 8637
rect 2384 8639 2389 8642
rect 2393 8639 2417 8642
rect 2442 8639 2449 8642
rect 2453 8639 2475 8642
rect 2495 8639 2502 8642
rect 2516 8639 2521 8642
rect 2525 8639 2549 8642
rect 2574 8639 2581 8642
rect 2585 8639 2607 8642
rect 2627 8639 2634 8642
rect 2648 8639 2653 8642
rect 2657 8639 2681 8642
rect 2706 8639 2713 8642
rect 2717 8639 2739 8642
rect 3213 8656 3216 8662
rect 3241 8659 3248 8662
rect 3252 8663 3267 8666
rect 3309 8663 3342 8667
rect 3346 8663 3370 8667
rect 3374 8663 3400 8667
rect 3404 8663 3437 8667
rect 3441 8663 3474 8667
rect 3478 8663 3502 8667
rect 3506 8663 3532 8667
rect 3536 8663 3569 8667
rect 3573 8663 3606 8667
rect 3610 8663 3634 8667
rect 3638 8663 3664 8667
rect 3668 8663 3701 8667
rect 3705 8663 3709 8667
rect 4112 8669 4117 8672
rect 4121 8669 4145 8672
rect 4170 8669 4177 8672
rect 4181 8669 4203 8672
rect 3312 8653 3315 8663
rect 3333 8653 3336 8663
rect 3349 8653 3352 8663
rect 3363 8656 3368 8660
rect 3372 8656 3379 8660
rect 3391 8653 3394 8663
rect 3407 8653 3410 8663
rect 3428 8653 3431 8663
rect 3444 8653 3447 8663
rect 3465 8653 3468 8663
rect 3481 8653 3484 8663
rect 3495 8656 3500 8660
rect 3504 8656 3511 8660
rect 3523 8653 3526 8663
rect 3539 8653 3542 8663
rect 3560 8653 3563 8663
rect 3576 8653 3579 8663
rect 3597 8653 3600 8663
rect 3613 8653 3616 8663
rect 3627 8656 3632 8660
rect 3636 8656 3643 8660
rect 3655 8653 3658 8663
rect 3671 8653 3674 8663
rect 3692 8653 3695 8663
rect 4128 8659 4135 8662
rect 4139 8663 4158 8666
rect 3150 8640 3153 8652
rect 3171 8640 3174 8652
rect 3187 8640 3190 8652
rect 3201 8643 3213 8646
rect 3229 8640 3232 8652
rect 3245 8640 3248 8652
rect 3266 8640 3269 8652
rect 343 8617 376 8627
rect 2400 8629 2407 8632
rect 2411 8633 2430 8636
rect 2430 8626 2433 8632
rect 2458 8629 2465 8632
rect 2469 8633 2484 8636
rect 2532 8629 2539 8632
rect 2543 8633 2562 8636
rect 2562 8626 2565 8632
rect 2590 8629 2597 8632
rect 2601 8633 2616 8636
rect 2664 8629 2671 8632
rect 2675 8633 2694 8636
rect 2694 8626 2697 8632
rect 2722 8629 2729 8632
rect 2733 8633 2750 8636
rect 2782 8636 3180 8640
rect 3184 8636 3208 8640
rect 3212 8636 3238 8640
rect 3242 8636 3279 8640
rect 3329 8639 3334 8642
rect 3338 8639 3362 8642
rect 3387 8639 3394 8642
rect 3398 8639 3420 8642
rect 3440 8639 3447 8642
rect 3461 8639 3466 8642
rect 3470 8639 3494 8642
rect 3519 8639 3526 8642
rect 3530 8639 3552 8642
rect 3572 8639 3579 8642
rect 3593 8639 3598 8642
rect 3602 8639 3626 8642
rect 3651 8639 3658 8642
rect 3662 8639 3684 8642
rect 4158 8656 4161 8662
rect 4186 8659 4193 8662
rect 4197 8663 4212 8666
rect 4826 8659 4829 8698
rect 4095 8640 4098 8652
rect 4116 8640 4119 8652
rect 4132 8640 4135 8652
rect 4146 8643 4158 8646
rect 4174 8640 4177 8652
rect 4190 8640 4193 8652
rect 4211 8640 4214 8652
rect 4816 8649 4829 8659
rect 2818 8629 3156 8633
rect 3160 8629 3207 8633
rect 3211 8629 3257 8633
rect 3261 8629 3279 8633
rect 3345 8629 3352 8632
rect 3356 8633 3375 8636
rect 343 8607 386 8617
rect 2367 8610 2370 8622
rect 2388 8610 2391 8622
rect 2404 8610 2407 8622
rect 2418 8613 2430 8616
rect 2446 8610 2449 8622
rect 2462 8610 2465 8622
rect 2483 8610 2486 8622
rect 2499 8610 2502 8622
rect 2520 8610 2523 8622
rect 2536 8610 2539 8622
rect 2550 8613 2562 8616
rect 2578 8610 2581 8622
rect 2594 8610 2597 8622
rect 2615 8610 2618 8622
rect 2631 8610 2634 8622
rect 2652 8610 2655 8622
rect 2668 8610 2671 8622
rect 2682 8613 2694 8616
rect 2710 8610 2713 8622
rect 2726 8610 2729 8622
rect 2747 8610 2750 8622
rect 3153 8622 3274 8625
rect 3375 8626 3378 8632
rect 3403 8629 3410 8632
rect 3414 8633 3429 8636
rect 3477 8629 3484 8632
rect 3488 8633 3507 8636
rect 3507 8626 3510 8632
rect 3535 8629 3542 8632
rect 3546 8633 3561 8636
rect 3609 8629 3616 8632
rect 3620 8633 3639 8636
rect 3639 8626 3642 8632
rect 3667 8629 3674 8632
rect 3678 8633 3695 8636
rect 3727 8636 4125 8640
rect 4129 8636 4153 8640
rect 4157 8636 4183 8640
rect 4187 8636 4224 8640
rect 4806 8639 4829 8649
rect 3763 8629 4101 8633
rect 4105 8629 4152 8633
rect 4156 8629 4202 8633
rect 4206 8629 4224 8633
rect 4796 8629 4829 8639
rect 2830 8614 3156 8618
rect 3160 8614 3192 8618
rect 3196 8614 3259 8618
rect 3263 8614 3279 8618
rect 343 8511 769 8607
rect 2364 8606 2397 8610
rect 2401 8606 2425 8610
rect 2429 8606 2455 8610
rect 2459 8606 2529 8610
rect 2533 8606 2557 8610
rect 2561 8606 2587 8610
rect 2591 8606 2661 8610
rect 2665 8606 2689 8610
rect 2693 8606 2719 8610
rect 2723 8606 2776 8610
rect 3146 8607 3180 8611
rect 3184 8607 3208 8611
rect 3212 8607 3238 8611
rect 3242 8607 3275 8611
rect 3312 8610 3315 8622
rect 3333 8610 3336 8622
rect 3349 8610 3352 8622
rect 3363 8613 3375 8616
rect 3391 8610 3394 8622
rect 3407 8610 3410 8622
rect 3428 8610 3431 8622
rect 3444 8610 3447 8622
rect 3465 8610 3468 8622
rect 3481 8610 3484 8622
rect 3495 8613 3507 8616
rect 3523 8610 3526 8622
rect 3539 8610 3542 8622
rect 3560 8610 3563 8622
rect 3576 8610 3579 8622
rect 3597 8610 3600 8622
rect 3613 8610 3616 8622
rect 3627 8613 3639 8616
rect 3655 8610 3658 8622
rect 3671 8610 3674 8622
rect 3692 8610 3695 8622
rect 4098 8622 4219 8625
rect 4786 8619 4829 8629
rect 3775 8614 4101 8618
rect 4105 8614 4137 8618
rect 4141 8614 4204 8618
rect 4208 8614 4224 8618
rect 2364 8599 2373 8603
rect 2377 8599 2424 8603
rect 2428 8599 2474 8603
rect 2478 8599 2505 8603
rect 2509 8599 2556 8603
rect 2560 8599 2606 8603
rect 2610 8599 2637 8603
rect 2641 8599 2688 8603
rect 2692 8599 2738 8603
rect 2742 8599 2812 8603
rect 3150 8597 3153 8607
rect 3171 8597 3174 8607
rect 3187 8597 3190 8607
rect 3201 8600 3206 8604
rect 3210 8600 3217 8604
rect 3229 8597 3232 8607
rect 3245 8597 3248 8607
rect 3266 8597 3269 8607
rect 3309 8606 3342 8610
rect 3346 8606 3370 8610
rect 3374 8606 3400 8610
rect 3404 8606 3474 8610
rect 3478 8606 3502 8610
rect 3506 8606 3532 8610
rect 3536 8606 3606 8610
rect 3610 8606 3634 8610
rect 3638 8606 3664 8610
rect 3668 8606 3721 8610
rect 4091 8607 4125 8611
rect 4129 8607 4153 8611
rect 4157 8607 4183 8611
rect 4187 8607 4220 8611
rect 3309 8599 3318 8603
rect 3322 8599 3369 8603
rect 3373 8599 3419 8603
rect 3423 8599 3450 8603
rect 3454 8599 3501 8603
rect 3505 8599 3551 8603
rect 3555 8599 3582 8603
rect 3586 8599 3633 8603
rect 3637 8599 3683 8603
rect 3687 8599 3757 8603
rect 4095 8597 4098 8607
rect 4116 8597 4119 8607
rect 4132 8597 4135 8607
rect 4146 8600 4151 8604
rect 4155 8600 4162 8604
rect 4174 8597 4177 8607
rect 4190 8597 4193 8607
rect 4211 8597 4214 8607
rect 2370 8592 2755 8595
rect 2364 8584 2373 8588
rect 2377 8584 2409 8588
rect 2413 8584 2476 8588
rect 2480 8584 2505 8588
rect 2509 8584 2541 8588
rect 2545 8584 2608 8588
rect 2612 8584 2637 8588
rect 2641 8584 2673 8588
rect 2677 8584 2740 8588
rect 2744 8584 2824 8588
rect 2364 8577 2397 8581
rect 2401 8577 2425 8581
rect 2429 8577 2455 8581
rect 2459 8577 2492 8581
rect 2496 8577 2529 8581
rect 2533 8577 2557 8581
rect 2561 8577 2587 8581
rect 2591 8577 2624 8581
rect 2628 8577 2661 8581
rect 2665 8577 2689 8581
rect 2693 8577 2719 8581
rect 2723 8577 2756 8581
rect 2760 8577 2764 8581
rect 3167 8583 3172 8586
rect 3176 8583 3200 8586
rect 3315 8592 3700 8595
rect 3225 8583 3232 8586
rect 3236 8583 3258 8586
rect 3309 8584 3318 8588
rect 3322 8584 3354 8588
rect 3358 8584 3421 8588
rect 3425 8584 3450 8588
rect 3454 8584 3486 8588
rect 3490 8584 3553 8588
rect 3557 8584 3582 8588
rect 3586 8584 3618 8588
rect 3622 8584 3685 8588
rect 3689 8584 3769 8588
rect 2367 8567 2370 8577
rect 2388 8567 2391 8577
rect 2404 8567 2407 8577
rect 2418 8570 2423 8574
rect 2427 8570 2434 8574
rect 2446 8567 2449 8577
rect 2462 8567 2465 8577
rect 2483 8567 2486 8577
rect 2499 8567 2502 8577
rect 2520 8567 2523 8577
rect 2536 8567 2539 8577
rect 2550 8570 2555 8574
rect 2559 8570 2566 8574
rect 2578 8567 2581 8577
rect 2594 8567 2597 8577
rect 2615 8567 2618 8577
rect 2631 8567 2634 8577
rect 2652 8567 2655 8577
rect 2668 8567 2671 8577
rect 2682 8570 2687 8574
rect 2691 8570 2698 8574
rect 2710 8567 2713 8577
rect 2726 8567 2729 8577
rect 2747 8567 2750 8577
rect 3183 8573 3190 8576
rect 3194 8577 3213 8580
rect 2384 8553 2389 8556
rect 2393 8553 2417 8556
rect 2442 8553 2449 8556
rect 2453 8553 2475 8556
rect 2495 8553 2502 8556
rect 2516 8553 2521 8556
rect 2525 8553 2549 8556
rect 2574 8553 2581 8556
rect 2585 8553 2607 8556
rect 2627 8553 2634 8556
rect 2648 8553 2653 8556
rect 2657 8553 2681 8556
rect 2706 8553 2713 8556
rect 2717 8553 2739 8556
rect 3213 8570 3216 8576
rect 3241 8573 3248 8576
rect 3252 8577 3267 8580
rect 3278 8575 3289 8579
rect 3309 8577 3342 8581
rect 3346 8577 3370 8581
rect 3374 8577 3400 8581
rect 3404 8577 3437 8581
rect 3441 8577 3474 8581
rect 3478 8577 3502 8581
rect 3506 8577 3532 8581
rect 3536 8577 3569 8581
rect 3573 8577 3606 8581
rect 3610 8577 3634 8581
rect 3638 8577 3664 8581
rect 3668 8577 3701 8581
rect 3705 8577 3709 8581
rect 4112 8583 4117 8586
rect 4121 8583 4145 8586
rect 4170 8583 4177 8586
rect 4181 8583 4203 8586
rect 3312 8567 3315 8577
rect 3333 8567 3336 8577
rect 3349 8567 3352 8577
rect 3363 8570 3368 8574
rect 3372 8570 3379 8574
rect 3391 8567 3394 8577
rect 3407 8567 3410 8577
rect 3428 8567 3431 8577
rect 3444 8567 3447 8577
rect 3465 8567 3468 8577
rect 3481 8567 3484 8577
rect 3495 8570 3500 8574
rect 3504 8570 3511 8574
rect 3523 8567 3526 8577
rect 3539 8567 3542 8577
rect 3560 8567 3563 8577
rect 3576 8567 3579 8577
rect 3597 8567 3600 8577
rect 3613 8567 3616 8577
rect 3627 8570 3632 8574
rect 3636 8570 3643 8574
rect 3655 8567 3658 8577
rect 3671 8567 3674 8577
rect 3692 8567 3695 8577
rect 4128 8573 4135 8576
rect 4139 8577 4158 8580
rect 3150 8554 3153 8566
rect 3171 8554 3174 8566
rect 3187 8554 3190 8566
rect 3201 8557 3213 8560
rect 3229 8554 3232 8566
rect 3245 8554 3248 8566
rect 3266 8554 3269 8566
rect 2400 8543 2407 8546
rect 2411 8547 2430 8550
rect 2430 8540 2433 8546
rect 2458 8543 2465 8546
rect 2469 8547 2484 8550
rect 2532 8543 2539 8546
rect 2543 8547 2562 8550
rect 2562 8540 2565 8546
rect 2590 8543 2597 8546
rect 2601 8547 2616 8550
rect 2664 8543 2671 8546
rect 2675 8547 2694 8550
rect 2694 8540 2697 8546
rect 2722 8543 2729 8546
rect 2733 8547 2750 8550
rect 2782 8550 3180 8554
rect 3184 8550 3208 8554
rect 3212 8550 3238 8554
rect 3242 8550 3279 8554
rect 3329 8553 3334 8556
rect 3338 8553 3362 8556
rect 3387 8553 3394 8556
rect 3398 8553 3420 8556
rect 3440 8553 3447 8556
rect 3461 8553 3466 8556
rect 3470 8553 3494 8556
rect 3519 8553 3526 8556
rect 3530 8553 3552 8556
rect 3572 8553 3579 8556
rect 3593 8553 3598 8556
rect 3602 8553 3626 8556
rect 3651 8553 3658 8556
rect 3662 8553 3684 8556
rect 4158 8570 4161 8576
rect 4186 8573 4193 8576
rect 4197 8577 4212 8580
rect 4223 8575 4234 8579
rect 4095 8554 4098 8566
rect 4116 8554 4119 8566
rect 4132 8554 4135 8566
rect 4146 8557 4158 8560
rect 4174 8554 4177 8566
rect 4190 8554 4193 8566
rect 4211 8554 4214 8566
rect 2818 8543 3156 8547
rect 3160 8543 3207 8547
rect 3211 8543 3257 8547
rect 3261 8543 3279 8547
rect 3345 8543 3352 8546
rect 3356 8547 3375 8550
rect 3375 8540 3378 8546
rect 3403 8543 3410 8546
rect 3414 8547 3429 8550
rect 3477 8543 3484 8546
rect 3488 8547 3507 8550
rect 3507 8540 3510 8546
rect 3535 8543 3542 8546
rect 3546 8547 3561 8550
rect 3609 8543 3616 8546
rect 3620 8547 3639 8550
rect 3639 8540 3642 8546
rect 3667 8543 3674 8546
rect 3678 8547 3695 8550
rect 3727 8550 4125 8554
rect 4129 8550 4153 8554
rect 4157 8550 4183 8554
rect 4187 8550 4224 8554
rect 3763 8543 4101 8547
rect 4105 8543 4152 8547
rect 4156 8543 4202 8547
rect 4206 8543 4224 8547
rect 2367 8524 2370 8536
rect 2388 8524 2391 8536
rect 2404 8524 2407 8536
rect 2418 8527 2430 8530
rect 2446 8524 2449 8536
rect 2462 8524 2465 8536
rect 2483 8524 2486 8536
rect 2499 8524 2502 8536
rect 2520 8524 2523 8536
rect 2536 8524 2539 8536
rect 2550 8527 2562 8530
rect 2578 8524 2581 8536
rect 2594 8524 2597 8536
rect 2615 8524 2618 8536
rect 2631 8524 2634 8536
rect 2652 8524 2655 8536
rect 2668 8524 2671 8536
rect 2682 8527 2694 8530
rect 2710 8524 2713 8536
rect 2726 8524 2729 8536
rect 2747 8524 2750 8536
rect 3312 8524 3315 8536
rect 3333 8524 3336 8536
rect 3349 8524 3352 8536
rect 3363 8527 3375 8530
rect 3391 8524 3394 8536
rect 3407 8524 3410 8536
rect 3428 8524 3431 8536
rect 3444 8524 3447 8536
rect 3465 8524 3468 8536
rect 3481 8524 3484 8536
rect 3495 8527 3507 8530
rect 3523 8524 3526 8536
rect 3539 8524 3542 8536
rect 3560 8524 3563 8536
rect 3576 8524 3579 8536
rect 3597 8524 3600 8536
rect 3613 8524 3616 8536
rect 3627 8527 3639 8530
rect 3655 8524 3658 8536
rect 3671 8524 3674 8536
rect 3692 8524 3695 8536
rect 2364 8520 2397 8524
rect 2401 8520 2425 8524
rect 2429 8520 2455 8524
rect 2459 8520 2529 8524
rect 2533 8520 2557 8524
rect 2561 8520 2587 8524
rect 2591 8520 2661 8524
rect 2665 8520 2689 8524
rect 2693 8520 2719 8524
rect 2723 8520 2776 8524
rect 3309 8520 3342 8524
rect 3346 8520 3370 8524
rect 3374 8520 3400 8524
rect 3404 8520 3474 8524
rect 3478 8520 3502 8524
rect 3506 8520 3532 8524
rect 3536 8520 3606 8524
rect 3610 8520 3634 8524
rect 3638 8520 3664 8524
rect 3668 8520 3721 8524
rect 4403 8523 4829 8619
rect 2364 8513 2373 8517
rect 2377 8513 2424 8517
rect 2428 8513 2474 8517
rect 2478 8513 2505 8517
rect 2509 8513 2556 8517
rect 2560 8513 2606 8517
rect 2610 8513 2637 8517
rect 2641 8513 2688 8517
rect 2692 8513 2738 8517
rect 2742 8513 2812 8517
rect 3309 8513 3318 8517
rect 3322 8513 3369 8517
rect 3373 8513 3419 8517
rect 3423 8513 3450 8517
rect 3454 8513 3501 8517
rect 3505 8513 3551 8517
rect 3555 8513 3582 8517
rect 3586 8513 3633 8517
rect 3637 8513 3683 8517
rect 3687 8513 3757 8517
rect 4786 8513 4829 8523
rect 343 8501 386 8511
rect 2370 8507 2755 8510
rect 3315 8507 3700 8510
rect 4796 8503 4829 8513
rect 343 8491 376 8501
rect 2495 8500 2599 8503
rect 3440 8500 3544 8503
rect 2611 8492 2615 8496
rect 2619 8492 2623 8496
rect 343 8481 366 8491
rect 3556 8492 3560 8496
rect 3564 8492 3568 8496
rect 4806 8493 4829 8503
rect 2354 8481 2599 8485
rect 2603 8481 2619 8485
rect 2635 8481 3296 8485
rect 3300 8481 3544 8485
rect 3548 8481 3564 8485
rect 3580 8481 4241 8485
rect 4245 8481 4323 8485
rect 4816 8483 4829 8493
rect 343 8471 356 8481
rect 2627 8474 2755 8477
rect 3572 8474 3700 8477
rect 343 8432 346 8471
rect 2642 8467 2755 8470
rect 3587 8467 3700 8470
rect 2611 8458 2615 8462
rect 2619 8458 2623 8462
rect 3556 8458 3560 8462
rect 3564 8458 3568 8462
rect 2495 8451 2599 8454
rect 3440 8451 3544 8454
rect 2364 8444 2373 8448
rect 2377 8444 2409 8448
rect 2413 8444 2476 8448
rect 2480 8444 2505 8448
rect 2509 8444 2541 8448
rect 2545 8444 2608 8448
rect 2612 8444 2637 8448
rect 2641 8444 2673 8448
rect 2677 8444 2740 8448
rect 2744 8444 2824 8448
rect 3309 8444 3318 8448
rect 3322 8444 3354 8448
rect 3358 8444 3421 8448
rect 3425 8444 3450 8448
rect 3454 8444 3486 8448
rect 3490 8444 3553 8448
rect 3557 8444 3582 8448
rect 3586 8444 3618 8448
rect 3622 8444 3685 8448
rect 3689 8444 3769 8448
rect 4826 8444 4829 8483
rect 5083 8444 5086 8698
rect 2364 8437 2397 8441
rect 2401 8437 2425 8441
rect 2429 8437 2455 8441
rect 2459 8437 2492 8441
rect 2496 8437 2529 8441
rect 2533 8437 2557 8441
rect 2561 8437 2587 8441
rect 2591 8437 2624 8441
rect 2628 8437 2661 8441
rect 2665 8437 2689 8441
rect 2693 8437 2719 8441
rect 2723 8437 2756 8441
rect 2760 8437 2764 8441
rect 3309 8437 3342 8441
rect 3346 8437 3370 8441
rect 3374 8437 3400 8441
rect 3404 8437 3437 8441
rect 3441 8437 3474 8441
rect 3478 8437 3502 8441
rect 3506 8437 3532 8441
rect 3536 8437 3569 8441
rect 3573 8437 3606 8441
rect 3610 8437 3634 8441
rect 3638 8437 3664 8441
rect 3668 8437 3701 8441
rect 3705 8437 3709 8441
rect 4483 8438 4484 8442
rect 4488 8438 4489 8442
rect 4493 8438 4494 8442
rect 4498 8438 4499 8442
rect 4503 8438 4504 8442
rect 4508 8438 4509 8442
rect 4479 8437 4513 8438
rect 86 8429 346 8432
rect 2367 8427 2370 8437
rect 2388 8427 2391 8437
rect 2404 8427 2407 8437
rect 2418 8430 2423 8434
rect 2427 8430 2434 8434
rect 2446 8427 2449 8437
rect 2462 8427 2465 8437
rect 2483 8427 2486 8437
rect 2499 8427 2502 8437
rect 2520 8427 2523 8437
rect 2536 8427 2539 8437
rect 2550 8430 2555 8434
rect 2559 8430 2566 8434
rect 2578 8427 2581 8437
rect 2594 8427 2597 8437
rect 2615 8427 2618 8437
rect 2631 8427 2634 8437
rect 2652 8427 2655 8437
rect 2668 8427 2671 8437
rect 2682 8430 2687 8434
rect 2691 8430 2698 8434
rect 2710 8427 2713 8437
rect 2726 8427 2729 8437
rect 2747 8427 2750 8437
rect 3312 8427 3315 8437
rect 3333 8427 3336 8437
rect 3349 8427 3352 8437
rect 3363 8430 3368 8434
rect 3372 8430 3379 8434
rect 3391 8427 3394 8437
rect 3407 8427 3410 8437
rect 3428 8427 3431 8437
rect 3444 8427 3447 8437
rect 3465 8427 3468 8437
rect 3481 8427 3484 8437
rect 3495 8430 3500 8434
rect 3504 8430 3511 8434
rect 3523 8427 3526 8437
rect 3539 8427 3542 8437
rect 3560 8427 3563 8437
rect 3576 8427 3579 8437
rect 3597 8427 3600 8437
rect 3613 8427 3616 8437
rect 3627 8430 3632 8434
rect 3636 8430 3643 8434
rect 3655 8427 3658 8437
rect 3671 8427 3674 8437
rect 3692 8427 3695 8437
rect 4483 8433 4484 8437
rect 4488 8433 4489 8437
rect 4493 8433 4494 8437
rect 4498 8433 4499 8437
rect 4503 8433 4504 8437
rect 4508 8433 4509 8437
rect 4479 8432 4513 8433
rect 4483 8428 4484 8432
rect 4488 8428 4489 8432
rect 4493 8428 4494 8432
rect 4498 8428 4499 8432
rect 4503 8428 4504 8432
rect 4508 8428 4509 8432
rect 4479 8427 4513 8428
rect 2384 8413 2389 8416
rect 2393 8413 2417 8416
rect 2442 8413 2449 8416
rect 2453 8413 2475 8416
rect 2495 8413 2502 8416
rect 2516 8413 2521 8416
rect 2525 8413 2549 8416
rect 2574 8413 2581 8416
rect 2585 8413 2607 8416
rect 2627 8413 2634 8416
rect 2648 8413 2653 8416
rect 2657 8413 2681 8416
rect 2706 8413 2713 8416
rect 2717 8413 2739 8416
rect 2400 8403 2407 8406
rect 2411 8407 2430 8410
rect 617 8394 618 8398
rect 622 8394 623 8398
rect 627 8394 628 8398
rect 632 8394 633 8398
rect 637 8394 638 8398
rect 642 8394 643 8398
rect 613 8393 647 8394
rect 617 8389 618 8393
rect 622 8389 623 8393
rect 627 8389 628 8393
rect 632 8389 633 8393
rect 637 8389 638 8393
rect 642 8389 643 8393
rect 613 8388 647 8389
rect 617 8384 618 8388
rect 622 8384 623 8388
rect 627 8384 628 8388
rect 632 8384 633 8388
rect 637 8384 638 8388
rect 642 8384 643 8388
rect 613 8383 647 8384
rect 86 8377 346 8380
rect 617 8379 618 8383
rect 622 8379 623 8383
rect 627 8379 628 8383
rect 632 8379 633 8383
rect 637 8379 638 8383
rect 642 8379 643 8383
rect 663 8394 664 8398
rect 668 8394 669 8398
rect 673 8394 674 8398
rect 678 8394 679 8398
rect 683 8394 684 8398
rect 688 8394 689 8398
rect 659 8393 693 8394
rect 663 8389 664 8393
rect 668 8389 669 8393
rect 673 8389 674 8393
rect 678 8389 679 8393
rect 683 8389 684 8393
rect 688 8389 689 8393
rect 659 8388 693 8389
rect 663 8384 664 8388
rect 668 8384 669 8388
rect 673 8384 674 8388
rect 678 8384 679 8388
rect 683 8384 684 8388
rect 688 8384 689 8388
rect 2430 8400 2433 8406
rect 2458 8403 2465 8406
rect 2469 8407 2484 8410
rect 2532 8403 2539 8406
rect 2543 8407 2562 8410
rect 2562 8400 2565 8406
rect 2590 8403 2597 8406
rect 2601 8407 2616 8410
rect 2664 8403 2671 8406
rect 2675 8407 2694 8410
rect 2694 8400 2697 8406
rect 2722 8403 2729 8406
rect 2733 8407 2750 8410
rect 3329 8413 3334 8416
rect 3338 8413 3362 8416
rect 3387 8413 3394 8416
rect 3398 8413 3420 8416
rect 3440 8413 3447 8416
rect 3461 8413 3466 8416
rect 3470 8413 3494 8416
rect 3519 8413 3526 8416
rect 3530 8413 3552 8416
rect 3572 8413 3579 8416
rect 3593 8413 3598 8416
rect 3602 8413 3626 8416
rect 4483 8423 4484 8427
rect 4488 8423 4489 8427
rect 4493 8423 4494 8427
rect 4498 8423 4499 8427
rect 4503 8423 4504 8427
rect 4508 8423 4509 8427
rect 4529 8438 4530 8442
rect 4534 8438 4535 8442
rect 4539 8438 4540 8442
rect 4544 8438 4545 8442
rect 4549 8438 4550 8442
rect 4554 8438 4555 8442
rect 4826 8441 5086 8444
rect 4525 8437 4559 8438
rect 4529 8433 4530 8437
rect 4534 8433 4535 8437
rect 4539 8433 4540 8437
rect 4544 8433 4545 8437
rect 4549 8433 4550 8437
rect 4554 8433 4555 8437
rect 4525 8432 4559 8433
rect 4529 8428 4530 8432
rect 4534 8428 4535 8432
rect 4539 8428 4540 8432
rect 4544 8428 4545 8432
rect 4549 8428 4550 8432
rect 4554 8428 4555 8432
rect 4525 8427 4559 8428
rect 4529 8423 4530 8427
rect 4534 8423 4535 8427
rect 4539 8423 4540 8427
rect 4544 8423 4545 8427
rect 4549 8423 4550 8427
rect 4554 8423 4555 8427
rect 3651 8413 3658 8416
rect 3662 8413 3684 8416
rect 3345 8403 3352 8406
rect 3356 8407 3375 8410
rect 3375 8400 3378 8406
rect 3403 8403 3410 8406
rect 3414 8407 3429 8410
rect 3477 8403 3484 8406
rect 3488 8407 3507 8410
rect 3507 8400 3510 8406
rect 3535 8403 3542 8406
rect 3546 8407 3561 8410
rect 3609 8403 3616 8406
rect 3620 8407 3639 8410
rect 3639 8400 3642 8406
rect 3667 8403 3674 8406
rect 3678 8407 3695 8410
rect 2367 8384 2370 8396
rect 2388 8384 2391 8396
rect 2404 8384 2407 8396
rect 2418 8387 2430 8390
rect 2446 8384 2449 8396
rect 2462 8384 2465 8396
rect 2483 8384 2486 8396
rect 2499 8384 2502 8396
rect 2520 8384 2523 8396
rect 2536 8384 2539 8396
rect 2550 8387 2562 8390
rect 2578 8384 2581 8396
rect 2594 8384 2597 8396
rect 2615 8384 2618 8396
rect 2631 8384 2634 8396
rect 2652 8384 2655 8396
rect 2668 8384 2671 8396
rect 2682 8387 2694 8390
rect 2710 8384 2713 8396
rect 2726 8384 2729 8396
rect 2747 8384 2750 8396
rect 3312 8384 3315 8396
rect 3333 8384 3336 8396
rect 3349 8384 3352 8396
rect 3363 8387 3375 8390
rect 3391 8384 3394 8396
rect 3407 8384 3410 8396
rect 3428 8384 3431 8396
rect 3444 8384 3447 8396
rect 3465 8384 3468 8396
rect 3481 8384 3484 8396
rect 3495 8387 3507 8390
rect 3523 8384 3526 8396
rect 3539 8384 3542 8396
rect 3560 8384 3563 8396
rect 3576 8384 3579 8396
rect 3597 8384 3600 8396
rect 3613 8384 3616 8396
rect 3627 8387 3639 8390
rect 3655 8384 3658 8396
rect 3671 8384 3674 8396
rect 3692 8384 3695 8396
rect 4826 8389 5086 8392
rect 659 8383 693 8384
rect 663 8379 664 8383
rect 668 8379 669 8383
rect 673 8379 674 8383
rect 678 8379 679 8383
rect 683 8379 684 8383
rect 688 8379 689 8383
rect 2364 8380 2397 8384
rect 2401 8380 2425 8384
rect 2429 8380 2455 8384
rect 2459 8380 2529 8384
rect 2533 8380 2557 8384
rect 2561 8380 2587 8384
rect 2591 8380 2661 8384
rect 2665 8380 2689 8384
rect 2693 8380 2719 8384
rect 2723 8380 2776 8384
rect 3309 8380 3342 8384
rect 3346 8380 3370 8384
rect 3374 8380 3400 8384
rect 3404 8380 3474 8384
rect 3478 8380 3502 8384
rect 3506 8380 3532 8384
rect 3536 8380 3606 8384
rect 3610 8380 3634 8384
rect 3638 8380 3664 8384
rect 3668 8380 3721 8384
rect 86 8123 89 8377
rect 343 8338 346 8377
rect 2364 8373 2373 8377
rect 2377 8373 2424 8377
rect 2428 8373 2474 8377
rect 2478 8373 2505 8377
rect 2509 8373 2556 8377
rect 2560 8373 2606 8377
rect 2610 8373 2637 8377
rect 2641 8373 2688 8377
rect 2692 8373 2738 8377
rect 2742 8373 2812 8377
rect 3309 8373 3318 8377
rect 3322 8373 3369 8377
rect 3373 8373 3419 8377
rect 3423 8373 3450 8377
rect 3454 8373 3501 8377
rect 3505 8373 3551 8377
rect 3555 8373 3582 8377
rect 3586 8373 3633 8377
rect 3637 8373 3683 8377
rect 3687 8373 3757 8377
rect 2830 8365 2857 8369
rect 2861 8365 2893 8369
rect 2897 8365 2960 8369
rect 2964 8365 2989 8369
rect 2993 8365 3025 8369
rect 3029 8365 3092 8369
rect 3096 8365 3121 8369
rect 3125 8365 3157 8369
rect 3161 8365 3224 8369
rect 3228 8365 3253 8369
rect 3257 8365 3289 8369
rect 3293 8365 3356 8369
rect 3360 8365 3376 8369
rect 3775 8365 3802 8369
rect 3806 8365 3838 8369
rect 3842 8365 3905 8369
rect 3909 8365 3934 8369
rect 3938 8365 3970 8369
rect 3974 8365 4037 8369
rect 4041 8365 4066 8369
rect 4070 8365 4102 8369
rect 4106 8365 4169 8369
rect 4173 8365 4198 8369
rect 4202 8365 4234 8369
rect 4238 8365 4301 8369
rect 4305 8365 4321 8369
rect 2770 8358 2881 8362
rect 2885 8358 2909 8362
rect 2913 8358 2939 8362
rect 2943 8358 2976 8362
rect 2980 8358 3013 8362
rect 3017 8358 3041 8362
rect 3045 8358 3071 8362
rect 3075 8358 3108 8362
rect 3112 8358 3145 8362
rect 3149 8358 3173 8362
rect 3177 8358 3203 8362
rect 3207 8358 3240 8362
rect 3244 8358 3277 8362
rect 3281 8358 3305 8362
rect 3309 8358 3335 8362
rect 3339 8358 3372 8362
rect 3715 8358 3826 8362
rect 3830 8358 3854 8362
rect 3858 8358 3884 8362
rect 3888 8358 3921 8362
rect 3925 8358 3958 8362
rect 3962 8358 3986 8362
rect 3990 8358 4016 8362
rect 4020 8358 4053 8362
rect 4057 8358 4090 8362
rect 4094 8358 4118 8362
rect 4122 8358 4148 8362
rect 4152 8358 4185 8362
rect 4189 8358 4222 8362
rect 4226 8358 4250 8362
rect 4254 8358 4280 8362
rect 4284 8358 4317 8362
rect 2851 8348 2854 8358
rect 2872 8348 2875 8358
rect 2888 8348 2891 8358
rect 2902 8351 2907 8355
rect 2911 8351 2918 8355
rect 2930 8348 2933 8358
rect 2946 8348 2949 8358
rect 2967 8348 2970 8358
rect 2983 8348 2986 8358
rect 3004 8348 3007 8358
rect 3020 8348 3023 8358
rect 3034 8351 3039 8355
rect 3043 8351 3050 8355
rect 3062 8348 3065 8358
rect 3078 8348 3081 8358
rect 3099 8348 3102 8358
rect 3115 8348 3118 8358
rect 3136 8348 3139 8358
rect 3152 8348 3155 8358
rect 3166 8351 3171 8355
rect 3175 8351 3182 8355
rect 3194 8348 3197 8358
rect 3210 8348 3213 8358
rect 3231 8348 3234 8358
rect 3247 8348 3250 8358
rect 3268 8348 3271 8358
rect 3284 8348 3287 8358
rect 3298 8351 3303 8355
rect 3307 8351 3314 8355
rect 3326 8348 3329 8358
rect 3342 8348 3345 8358
rect 3363 8348 3366 8358
rect 3796 8348 3799 8358
rect 3817 8348 3820 8358
rect 3833 8348 3836 8358
rect 3847 8351 3852 8355
rect 3856 8351 3863 8355
rect 3875 8348 3878 8358
rect 3891 8348 3894 8358
rect 3912 8348 3915 8358
rect 3928 8348 3931 8358
rect 3949 8348 3952 8358
rect 3965 8348 3968 8358
rect 3979 8351 3984 8355
rect 3988 8351 3995 8355
rect 4007 8348 4010 8358
rect 4023 8348 4026 8358
rect 4044 8348 4047 8358
rect 4060 8348 4063 8358
rect 4081 8348 4084 8358
rect 4097 8348 4100 8358
rect 4111 8351 4116 8355
rect 4120 8351 4127 8355
rect 4139 8348 4142 8358
rect 4155 8348 4158 8358
rect 4176 8348 4179 8358
rect 4192 8348 4195 8358
rect 4213 8348 4216 8358
rect 4229 8348 4232 8358
rect 4243 8351 4248 8355
rect 4252 8351 4259 8355
rect 4271 8348 4274 8358
rect 4287 8348 4290 8358
rect 4308 8348 4311 8358
rect 4826 8350 4829 8389
rect 343 8328 356 8338
rect 2496 8332 2505 8336
rect 2509 8332 2541 8336
rect 2545 8332 2608 8336
rect 2612 8332 2824 8336
rect 2868 8334 2873 8337
rect 2877 8334 2901 8337
rect 2926 8334 2933 8337
rect 2937 8334 2959 8337
rect 343 8318 366 8328
rect 2496 8325 2529 8329
rect 2533 8325 2557 8329
rect 2561 8325 2587 8329
rect 2591 8325 2624 8329
rect 2628 8325 2764 8329
rect 343 8308 376 8318
rect 2499 8315 2502 8325
rect 2520 8315 2523 8325
rect 2536 8315 2539 8325
rect 2550 8318 2555 8322
rect 2559 8318 2566 8322
rect 2578 8315 2581 8325
rect 2594 8315 2597 8325
rect 2615 8315 2618 8325
rect 2884 8324 2891 8327
rect 2895 8328 2914 8331
rect 2914 8321 2917 8327
rect 2942 8324 2949 8327
rect 2953 8328 2970 8331
rect 3000 8334 3005 8337
rect 3009 8334 3033 8337
rect 3058 8334 3065 8337
rect 3069 8334 3091 8337
rect 3016 8324 3023 8327
rect 3027 8328 3046 8331
rect 3046 8321 3049 8327
rect 3074 8324 3081 8327
rect 3085 8328 3102 8331
rect 3132 8334 3137 8337
rect 3141 8334 3165 8337
rect 3190 8334 3197 8337
rect 3201 8334 3223 8337
rect 3148 8324 3155 8327
rect 3159 8328 3178 8331
rect 3178 8321 3181 8327
rect 3206 8324 3213 8327
rect 3217 8328 3234 8331
rect 3264 8334 3269 8337
rect 3273 8334 3297 8337
rect 3322 8334 3329 8337
rect 3333 8334 3355 8337
rect 3441 8332 3450 8336
rect 3454 8332 3486 8336
rect 3490 8332 3553 8336
rect 3557 8332 3769 8336
rect 3280 8324 3287 8327
rect 3291 8328 3310 8331
rect 343 8298 386 8308
rect 2494 8298 2503 8302
rect 2516 8301 2521 8304
rect 2525 8301 2549 8304
rect 2574 8301 2581 8304
rect 2585 8301 2607 8304
rect 2851 8305 2854 8317
rect 2872 8305 2875 8317
rect 2888 8305 2891 8317
rect 2902 8308 2914 8311
rect 2930 8305 2933 8317
rect 2946 8305 2949 8317
rect 2967 8305 2970 8317
rect 2983 8305 2986 8317
rect 3004 8305 3007 8317
rect 3020 8305 3023 8317
rect 3034 8308 3046 8311
rect 3062 8305 3065 8317
rect 3078 8305 3081 8317
rect 3099 8305 3102 8317
rect 3115 8305 3118 8317
rect 3136 8305 3139 8317
rect 3152 8305 3155 8317
rect 3166 8308 3178 8311
rect 3194 8305 3197 8317
rect 3210 8305 3213 8317
rect 3231 8305 3234 8317
rect 3310 8321 3313 8327
rect 3338 8324 3345 8327
rect 3349 8328 3366 8331
rect 3813 8334 3818 8337
rect 3822 8334 3846 8337
rect 3871 8334 3878 8337
rect 3882 8334 3904 8337
rect 3441 8325 3474 8329
rect 3478 8325 3502 8329
rect 3506 8325 3532 8329
rect 3536 8325 3569 8329
rect 3573 8325 3709 8329
rect 3247 8305 3250 8317
rect 3268 8305 3271 8317
rect 3284 8305 3287 8317
rect 3298 8308 3310 8311
rect 3326 8305 3329 8317
rect 3342 8305 3345 8317
rect 3363 8305 3366 8317
rect 3444 8315 3447 8325
rect 3465 8315 3468 8325
rect 3481 8315 3484 8325
rect 3495 8318 3500 8322
rect 3504 8318 3511 8322
rect 3523 8315 3526 8325
rect 3539 8315 3542 8325
rect 3560 8315 3563 8325
rect 3829 8324 3836 8327
rect 3840 8328 3859 8331
rect 3859 8321 3862 8327
rect 3887 8324 3894 8327
rect 3898 8328 3915 8331
rect 3945 8334 3950 8337
rect 3954 8334 3978 8337
rect 4003 8334 4010 8337
rect 4014 8334 4036 8337
rect 3961 8324 3968 8327
rect 3972 8328 3991 8331
rect 3991 8321 3994 8327
rect 4019 8324 4026 8327
rect 4030 8328 4047 8331
rect 4077 8334 4082 8337
rect 4086 8334 4110 8337
rect 4135 8334 4142 8337
rect 4146 8334 4168 8337
rect 4093 8324 4100 8327
rect 4104 8328 4123 8331
rect 4123 8321 4126 8327
rect 4151 8324 4158 8327
rect 4162 8328 4179 8331
rect 4209 8334 4214 8337
rect 4218 8334 4242 8337
rect 4816 8340 4829 8350
rect 4267 8334 4274 8337
rect 4278 8334 4300 8337
rect 4225 8324 4232 8327
rect 4236 8328 4255 8331
rect 2782 8301 2881 8305
rect 2885 8301 2909 8305
rect 2913 8301 2939 8305
rect 2943 8301 3013 8305
rect 3017 8301 3041 8305
rect 3045 8301 3071 8305
rect 3075 8301 3145 8305
rect 3149 8301 3173 8305
rect 3177 8301 3203 8305
rect 3207 8301 3277 8305
rect 3281 8301 3305 8305
rect 3309 8301 3335 8305
rect 3339 8301 3376 8305
rect 343 8202 769 8298
rect 2532 8291 2539 8294
rect 2543 8295 2562 8298
rect 2562 8288 2565 8294
rect 2590 8291 2597 8294
rect 2601 8295 2616 8298
rect 3439 8298 3448 8302
rect 3461 8301 3466 8304
rect 3470 8301 3494 8304
rect 3519 8301 3526 8304
rect 3530 8301 3552 8304
rect 3796 8305 3799 8317
rect 3817 8305 3820 8317
rect 3833 8305 3836 8317
rect 3847 8308 3859 8311
rect 3875 8305 3878 8317
rect 3891 8305 3894 8317
rect 3912 8305 3915 8317
rect 3928 8305 3931 8317
rect 3949 8305 3952 8317
rect 3965 8305 3968 8317
rect 3979 8308 3991 8311
rect 4007 8305 4010 8317
rect 4023 8305 4026 8317
rect 4044 8305 4047 8317
rect 4060 8305 4063 8317
rect 4081 8305 4084 8317
rect 4097 8305 4100 8317
rect 4111 8308 4123 8311
rect 4139 8305 4142 8317
rect 4155 8305 4158 8317
rect 4176 8305 4179 8317
rect 4255 8321 4258 8327
rect 4283 8324 4290 8327
rect 4294 8328 4311 8331
rect 4806 8330 4829 8340
rect 4796 8320 4829 8330
rect 4192 8305 4195 8317
rect 4213 8305 4216 8317
rect 4229 8305 4232 8317
rect 4243 8308 4255 8311
rect 4271 8305 4274 8317
rect 4287 8305 4290 8317
rect 4308 8305 4311 8317
rect 4786 8310 4829 8320
rect 3727 8301 3826 8305
rect 3830 8301 3854 8305
rect 3858 8301 3884 8305
rect 3888 8301 3958 8305
rect 3962 8301 3986 8305
rect 3990 8301 4016 8305
rect 4020 8301 4090 8305
rect 4094 8301 4118 8305
rect 4122 8301 4148 8305
rect 4152 8301 4222 8305
rect 4226 8301 4250 8305
rect 4254 8301 4280 8305
rect 4284 8301 4321 8305
rect 2818 8294 2857 8298
rect 2861 8294 2908 8298
rect 2912 8294 2958 8298
rect 2962 8294 2989 8298
rect 2993 8294 3040 8298
rect 3044 8294 3090 8298
rect 3094 8294 3121 8298
rect 3125 8294 3172 8298
rect 3176 8294 3222 8298
rect 3226 8294 3253 8298
rect 3257 8294 3304 8298
rect 3308 8294 3354 8298
rect 3358 8294 3376 8298
rect 3477 8291 3484 8294
rect 3488 8295 3507 8298
rect 2499 8272 2502 8284
rect 2520 8272 2523 8284
rect 2536 8272 2539 8284
rect 2550 8275 2562 8278
rect 2578 8272 2581 8284
rect 2594 8272 2597 8284
rect 2615 8272 2618 8284
rect 2770 8281 2855 8285
rect 2859 8281 2871 8285
rect 2875 8281 2889 8285
rect 2893 8281 2900 8285
rect 2904 8281 2906 8285
rect 2910 8281 2925 8285
rect 2929 8281 2962 8285
rect 2966 8281 2967 8285
rect 2971 8281 2979 8285
rect 2983 8281 3007 8285
rect 3011 8281 3023 8285
rect 3027 8281 3047 8285
rect 3051 8281 3101 8285
rect 3105 8281 3128 8285
rect 3132 8281 3182 8285
rect 3186 8281 3205 8285
rect 3507 8288 3510 8294
rect 3535 8291 3542 8294
rect 3546 8295 3561 8298
rect 3763 8294 3802 8298
rect 3806 8294 3853 8298
rect 3857 8294 3903 8298
rect 3907 8294 3934 8298
rect 3938 8294 3985 8298
rect 3989 8294 4035 8298
rect 4039 8294 4066 8298
rect 4070 8294 4117 8298
rect 4121 8294 4167 8298
rect 4171 8294 4198 8298
rect 4202 8294 4249 8298
rect 4253 8294 4299 8298
rect 4303 8294 4321 8298
rect 2806 8274 2882 8278
rect 2886 8274 2913 8278
rect 2917 8274 2935 8278
rect 2939 8274 3000 8278
rect 3004 8274 3018 8278
rect 3030 8277 3033 8281
rect 2496 8268 2529 8272
rect 2533 8268 2557 8272
rect 2561 8268 2587 8272
rect 2591 8268 2776 8272
rect 2496 8261 2505 8265
rect 2509 8261 2556 8265
rect 2560 8261 2606 8265
rect 2610 8261 2812 8265
rect 2925 8267 2928 8271
rect 2952 8267 2953 8271
rect 2997 8267 2999 8271
rect 3039 8264 3042 8269
rect 3054 8271 3057 8281
rect 3084 8277 3087 8281
rect 3111 8277 3114 8281
rect 2494 8245 2510 8249
rect 2619 8247 2623 8251
rect 2635 8247 2639 8251
rect 2643 8247 2857 8251
rect 2865 8250 2868 8256
rect 2872 8250 2875 8256
rect 2865 8247 2875 8250
rect 2865 8242 2868 8247
rect 2502 8238 2506 8242
rect 2518 8238 2639 8242
rect 2872 8242 2875 8247
rect 2881 8252 2884 8256
rect 2881 8248 2883 8252
rect 2887 8248 2889 8252
rect 2897 8251 2900 8256
rect 2925 8253 2928 8256
rect 2897 8249 2908 8251
rect 2881 8242 2884 8248
rect 2897 8247 2903 8249
rect 2897 8242 2900 8247
rect 2907 8247 2908 8249
rect 2926 8249 2928 8253
rect 2925 8242 2928 8249
rect 3028 8260 3031 8263
rect 3070 8260 3073 8263
rect 2941 8252 2944 8256
rect 2951 8252 2954 8256
rect 2951 8248 2960 8252
rect 2972 8251 2975 8256
rect 2997 8252 3000 8256
rect 2941 8242 2944 8248
rect 2951 8242 2954 8248
rect 2972 8247 2973 8251
rect 2977 8247 2980 8250
rect 2999 8248 3000 8252
rect 3015 8251 3018 8256
rect 3039 8255 3042 8260
rect 3047 8256 3058 8259
rect 3070 8257 3078 8260
rect 2972 8242 2975 8247
rect 2997 8242 3000 8248
rect 3015 8242 3018 8247
rect 2489 8230 2505 8234
rect 2509 8230 2572 8234
rect 2576 8230 2608 8234
rect 2612 8230 2824 8234
rect 2917 8229 2918 8233
rect 2942 8230 2943 8234
rect 2989 8229 2990 8233
rect 2493 8223 2526 8227
rect 2530 8223 2556 8227
rect 2560 8223 2584 8227
rect 2588 8223 2764 8227
rect 2499 8213 2502 8223
rect 2520 8213 2523 8223
rect 2536 8213 2539 8223
rect 2551 8216 2558 8220
rect 2562 8216 2567 8220
rect 2578 8213 2581 8223
rect 2594 8213 2597 8223
rect 2615 8213 2618 8223
rect 2794 8222 2870 8226
rect 2874 8222 2929 8226
rect 2933 8222 2954 8226
rect 2958 8222 2985 8226
rect 2989 8222 3018 8226
rect 3030 8219 3033 8251
rect 3047 8250 3050 8256
rect 3070 8251 3073 8257
rect 3082 8252 3085 8255
rect 3093 8255 3096 8269
rect 3120 8264 3123 8269
rect 3135 8271 3138 8281
rect 3165 8277 3168 8281
rect 3104 8260 3105 8263
rect 3109 8260 3112 8263
rect 3444 8272 3447 8284
rect 3465 8272 3468 8284
rect 3481 8272 3484 8284
rect 3495 8275 3507 8278
rect 3523 8272 3526 8284
rect 3539 8272 3542 8284
rect 3560 8272 3563 8284
rect 3715 8281 3800 8285
rect 3804 8281 3816 8285
rect 3820 8281 3834 8285
rect 3838 8281 3845 8285
rect 3849 8281 3851 8285
rect 3855 8281 3870 8285
rect 3874 8281 3907 8285
rect 3911 8281 3912 8285
rect 3916 8281 3924 8285
rect 3928 8281 3952 8285
rect 3956 8281 3968 8285
rect 3972 8281 3992 8285
rect 3996 8281 4046 8285
rect 4050 8281 4073 8285
rect 4077 8281 4127 8285
rect 4131 8281 4150 8285
rect 3751 8274 3827 8278
rect 3831 8274 3858 8278
rect 3862 8274 3880 8278
rect 3884 8274 3945 8278
rect 3949 8274 3963 8278
rect 3975 8277 3978 8281
rect 3151 8260 3154 8263
rect 3093 8252 3101 8255
rect 3120 8255 3123 8260
rect 3093 8247 3096 8252
rect 3101 8248 3105 8252
rect 3128 8256 3139 8259
rect 3151 8257 3159 8260
rect 3045 8241 3050 8246
rect 3054 8219 3057 8247
rect 3084 8219 3087 8243
rect 3111 8219 3114 8251
rect 3128 8250 3131 8256
rect 3151 8251 3154 8257
rect 3163 8252 3166 8255
rect 3174 8255 3177 8269
rect 3441 8268 3474 8272
rect 3478 8268 3502 8272
rect 3506 8268 3532 8272
rect 3536 8268 3721 8272
rect 3441 8261 3450 8265
rect 3454 8261 3501 8265
rect 3505 8261 3551 8265
rect 3555 8261 3757 8265
rect 3870 8267 3873 8271
rect 3897 8267 3898 8271
rect 3942 8267 3944 8271
rect 3984 8264 3987 8269
rect 3999 8271 4002 8281
rect 4029 8277 4032 8281
rect 4056 8277 4059 8281
rect 3174 8252 3186 8255
rect 3174 8247 3177 8252
rect 3126 8241 3131 8246
rect 3135 8219 3138 8247
rect 3439 8245 3455 8249
rect 3564 8247 3568 8251
rect 3580 8247 3584 8251
rect 3588 8247 3802 8251
rect 3810 8250 3813 8256
rect 3817 8250 3820 8256
rect 3810 8247 3820 8250
rect 3165 8219 3168 8243
rect 3810 8242 3813 8247
rect 3447 8238 3451 8242
rect 3463 8238 3584 8242
rect 3817 8242 3820 8247
rect 3826 8252 3829 8256
rect 3826 8248 3828 8252
rect 3832 8248 3834 8252
rect 3842 8251 3845 8256
rect 3870 8253 3873 8256
rect 3842 8249 3853 8251
rect 3826 8242 3829 8248
rect 3842 8247 3848 8249
rect 3842 8242 3845 8247
rect 3852 8247 3853 8249
rect 3871 8249 3873 8253
rect 3870 8242 3873 8249
rect 3973 8260 3976 8263
rect 4015 8260 4018 8263
rect 3886 8252 3889 8256
rect 3896 8252 3899 8256
rect 3896 8248 3905 8252
rect 3917 8251 3920 8256
rect 3942 8252 3945 8256
rect 3886 8242 3889 8248
rect 3896 8242 3899 8248
rect 3917 8247 3918 8251
rect 3922 8247 3925 8250
rect 3944 8248 3945 8252
rect 3960 8251 3963 8256
rect 3984 8255 3987 8260
rect 3992 8256 4003 8259
rect 4015 8257 4023 8260
rect 3917 8242 3920 8247
rect 3942 8242 3945 8248
rect 3960 8242 3963 8247
rect 3434 8230 3450 8234
rect 3454 8230 3517 8234
rect 3521 8230 3553 8234
rect 3557 8230 3769 8234
rect 3862 8229 3863 8233
rect 3887 8230 3888 8234
rect 3934 8229 3935 8233
rect 3438 8223 3471 8227
rect 3475 8223 3501 8227
rect 3505 8223 3529 8227
rect 3533 8223 3709 8227
rect 2782 8215 2856 8219
rect 2860 8215 2862 8219
rect 2866 8215 2870 8219
rect 2874 8215 2888 8219
rect 2892 8215 2897 8219
rect 2901 8215 2906 8219
rect 2910 8215 2929 8219
rect 2933 8215 2963 8219
rect 2967 8215 2978 8219
rect 2982 8215 3006 8219
rect 3010 8215 3023 8219
rect 3027 8215 3047 8219
rect 3051 8215 3101 8219
rect 3108 8215 3128 8219
rect 3132 8215 3182 8219
rect 343 8192 386 8202
rect 2510 8199 2532 8202
rect 2536 8199 2543 8202
rect 2794 8208 2870 8212
rect 2874 8208 2929 8212
rect 2933 8208 2954 8212
rect 2958 8208 2985 8212
rect 2989 8208 3018 8212
rect 2568 8199 2592 8202
rect 2596 8199 2601 8202
rect 2917 8201 2918 8205
rect 2942 8200 2943 8204
rect 2989 8201 2990 8205
rect 2614 8196 2623 8200
rect 2501 8193 2516 8196
rect 343 8182 376 8192
rect 2555 8193 2574 8196
rect 2520 8189 2527 8192
rect 2552 8186 2555 8192
rect 2578 8189 2585 8192
rect 2865 8187 2868 8192
rect 2872 8187 2875 8192
rect 2855 8184 2857 8187
rect 2865 8184 2875 8187
rect 343 8172 366 8182
rect 343 8162 356 8172
rect 2499 8170 2502 8182
rect 2520 8170 2523 8182
rect 2536 8170 2539 8182
rect 2555 8173 2567 8176
rect 2578 8170 2581 8182
rect 2594 8170 2597 8182
rect 2615 8170 2618 8182
rect 2865 8178 2868 8184
rect 2872 8178 2875 8184
rect 2881 8186 2884 8192
rect 2897 8187 2900 8192
rect 2881 8182 2883 8186
rect 2887 8182 2889 8186
rect 2897 8185 2903 8187
rect 2907 8185 2908 8187
rect 2897 8183 2908 8185
rect 2925 8185 2928 8192
rect 2881 8178 2884 8182
rect 2897 8178 2900 8183
rect 2926 8181 2928 8185
rect 2925 8178 2928 8181
rect 2941 8186 2944 8192
rect 2951 8186 2954 8192
rect 2972 8187 2975 8192
rect 2951 8182 2960 8186
rect 2972 8183 2973 8187
rect 2977 8184 2980 8187
rect 2997 8186 3000 8192
rect 3015 8187 3018 8192
rect 3054 8195 3057 8215
rect 3135 8195 3138 8215
rect 3444 8213 3447 8223
rect 3465 8213 3468 8223
rect 3481 8213 3484 8223
rect 3496 8216 3503 8220
rect 3507 8216 3512 8220
rect 3523 8213 3526 8223
rect 3539 8213 3542 8223
rect 3560 8213 3563 8223
rect 3739 8222 3815 8226
rect 3819 8222 3874 8226
rect 3878 8222 3899 8226
rect 3903 8222 3930 8226
rect 3934 8222 3963 8226
rect 3975 8219 3978 8251
rect 3992 8250 3995 8256
rect 4015 8251 4018 8257
rect 4027 8252 4030 8255
rect 4038 8255 4041 8269
rect 4065 8264 4068 8269
rect 4080 8271 4083 8281
rect 4110 8277 4113 8281
rect 4049 8260 4050 8263
rect 4054 8260 4057 8263
rect 4096 8260 4099 8263
rect 4038 8252 4046 8255
rect 4065 8255 4068 8260
rect 4038 8247 4041 8252
rect 4046 8248 4050 8252
rect 4073 8256 4084 8259
rect 4096 8257 4104 8260
rect 3990 8241 3995 8246
rect 3999 8219 4002 8247
rect 4029 8219 4032 8243
rect 4056 8219 4059 8251
rect 4073 8250 4076 8256
rect 4096 8251 4099 8257
rect 4108 8252 4111 8255
rect 4119 8255 4122 8269
rect 4119 8252 4131 8255
rect 4119 8247 4122 8252
rect 4071 8241 4076 8246
rect 4080 8219 4083 8247
rect 4110 8219 4113 8243
rect 3727 8215 3801 8219
rect 3805 8215 3807 8219
rect 3811 8215 3815 8219
rect 3819 8215 3833 8219
rect 3837 8215 3842 8219
rect 3846 8215 3851 8219
rect 3855 8215 3874 8219
rect 3878 8215 3908 8219
rect 3912 8215 3923 8219
rect 3927 8215 3951 8219
rect 3955 8215 3968 8219
rect 3972 8215 3992 8219
rect 3996 8215 4046 8219
rect 4053 8215 4073 8219
rect 4077 8215 4127 8219
rect 3455 8199 3477 8202
rect 3481 8199 3488 8202
rect 3739 8208 3815 8212
rect 3819 8208 3874 8212
rect 3878 8208 3899 8212
rect 3903 8208 3930 8212
rect 3934 8208 3963 8212
rect 3513 8199 3537 8202
rect 3541 8199 3546 8202
rect 3862 8201 3863 8205
rect 3887 8200 3888 8204
rect 3934 8201 3935 8205
rect 3559 8196 3568 8200
rect 3446 8193 3461 8196
rect 2941 8178 2944 8182
rect 2951 8178 2954 8182
rect 2972 8178 2975 8183
rect 2999 8182 3000 8186
rect 2997 8178 3000 8182
rect 3015 8178 3018 8183
rect 3045 8182 3050 8187
rect 3054 8183 3055 8186
rect 3070 8185 3073 8191
rect 3070 8182 3078 8185
rect 3125 8182 3130 8187
rect 3134 8183 3136 8186
rect 3151 8185 3154 8191
rect 3500 8193 3519 8196
rect 3465 8189 3472 8192
rect 3497 8186 3500 8192
rect 3151 8182 3159 8185
rect 3523 8189 3530 8192
rect 3810 8187 3813 8192
rect 3817 8187 3820 8192
rect 3800 8184 3802 8187
rect 3810 8184 3820 8187
rect 3070 8179 3073 8182
rect 3151 8179 3154 8182
rect 2489 8166 2526 8170
rect 2530 8166 2556 8170
rect 2560 8166 2584 8170
rect 2588 8166 2776 8170
rect 2925 8163 2928 8167
rect 2952 8163 2953 8167
rect 2997 8163 2999 8167
rect 343 8123 346 8162
rect 2489 8159 2507 8163
rect 2511 8159 2557 8163
rect 2561 8159 2608 8163
rect 2612 8159 2812 8163
rect 2870 8156 2882 8160
rect 2886 8156 2913 8160
rect 2917 8156 2935 8160
rect 2939 8156 3000 8160
rect 3004 8156 3018 8160
rect 3054 8153 3057 8171
rect 3135 8153 3138 8171
rect 3444 8170 3447 8182
rect 3465 8170 3468 8182
rect 3481 8170 3484 8182
rect 3500 8173 3512 8176
rect 3523 8170 3526 8182
rect 3539 8170 3542 8182
rect 3560 8170 3563 8182
rect 3810 8178 3813 8184
rect 3817 8178 3820 8184
rect 3826 8186 3829 8192
rect 3842 8187 3845 8192
rect 3826 8182 3828 8186
rect 3832 8182 3834 8186
rect 3842 8185 3848 8187
rect 3852 8185 3853 8187
rect 3842 8183 3853 8185
rect 3870 8185 3873 8192
rect 3826 8178 3829 8182
rect 3842 8178 3845 8183
rect 3871 8181 3873 8185
rect 3870 8178 3873 8181
rect 3886 8186 3889 8192
rect 3896 8186 3899 8192
rect 3917 8187 3920 8192
rect 3896 8182 3905 8186
rect 3917 8183 3918 8187
rect 3922 8184 3925 8187
rect 3942 8186 3945 8192
rect 3960 8187 3963 8192
rect 3999 8195 4002 8215
rect 4080 8195 4083 8215
rect 4403 8214 4829 8310
rect 4786 8204 4829 8214
rect 4796 8194 4829 8204
rect 3886 8178 3889 8182
rect 3896 8178 3899 8182
rect 3917 8178 3920 8183
rect 3944 8182 3945 8186
rect 3942 8178 3945 8182
rect 3960 8178 3963 8183
rect 3990 8182 3995 8187
rect 3999 8183 4000 8186
rect 4015 8185 4018 8191
rect 4015 8182 4023 8185
rect 4070 8182 4075 8187
rect 4079 8183 4081 8186
rect 4096 8185 4099 8191
rect 4096 8182 4104 8185
rect 4806 8184 4829 8194
rect 4015 8179 4018 8182
rect 4096 8179 4099 8182
rect 4816 8174 4829 8184
rect 3434 8166 3471 8170
rect 3475 8166 3501 8170
rect 3505 8166 3529 8170
rect 3533 8166 3721 8170
rect 3870 8163 3873 8167
rect 3897 8163 3898 8167
rect 3942 8163 3944 8167
rect 3434 8159 3452 8163
rect 3456 8159 3502 8163
rect 3506 8159 3553 8163
rect 3557 8159 3757 8163
rect 3815 8156 3827 8160
rect 3831 8156 3858 8160
rect 3862 8156 3880 8160
rect 3884 8156 3945 8160
rect 3949 8156 3963 8160
rect 3999 8153 4002 8171
rect 4080 8153 4083 8171
rect 2770 8149 2855 8153
rect 2859 8149 2871 8153
rect 2875 8149 2889 8153
rect 2893 8149 2900 8153
rect 2904 8149 2906 8153
rect 2910 8149 2925 8153
rect 2929 8149 2962 8153
rect 2966 8149 2967 8153
rect 2971 8149 2979 8153
rect 2983 8149 3007 8153
rect 3011 8149 3023 8153
rect 3027 8149 3047 8153
rect 3051 8149 3101 8153
rect 3105 8149 3128 8153
rect 3132 8149 3190 8153
rect 3194 8149 3205 8153
rect 3715 8149 3800 8153
rect 3804 8149 3816 8153
rect 3820 8149 3834 8153
rect 3838 8149 3845 8153
rect 3849 8149 3851 8153
rect 3855 8149 3870 8153
rect 3874 8149 3907 8153
rect 3911 8149 3912 8153
rect 3916 8149 3924 8153
rect 3928 8149 3952 8153
rect 3956 8149 3968 8153
rect 3972 8149 3992 8153
rect 3996 8149 4046 8153
rect 4050 8149 4073 8153
rect 4077 8149 4135 8153
rect 4139 8149 4150 8153
rect 2806 8142 2866 8146
rect 2870 8142 2882 8146
rect 2886 8142 2913 8146
rect 2917 8142 2935 8146
rect 2939 8142 3000 8146
rect 3004 8142 3018 8146
rect 3054 8139 3057 8149
rect 3084 8145 3087 8149
rect 3135 8145 3138 8149
rect 2925 8135 2928 8139
rect 2952 8135 2953 8139
rect 2997 8135 2999 8139
rect 86 8120 346 8123
rect 2854 8115 2857 8118
rect 2865 8118 2868 8124
rect 2872 8118 2875 8124
rect 2865 8115 2875 8118
rect 2865 8110 2868 8115
rect 2872 8110 2875 8115
rect 2881 8120 2884 8124
rect 2881 8116 2883 8120
rect 2887 8116 2889 8120
rect 2897 8119 2900 8124
rect 2925 8121 2928 8124
rect 2897 8117 2908 8119
rect 2881 8110 2884 8116
rect 2897 8115 2903 8117
rect 2897 8110 2900 8115
rect 2907 8115 2908 8117
rect 2926 8117 2928 8121
rect 2925 8110 2928 8117
rect 3070 8128 3073 8131
rect 2941 8120 2944 8124
rect 2951 8120 2954 8124
rect 2951 8116 2960 8120
rect 2972 8119 2975 8124
rect 2997 8120 3000 8124
rect 2941 8110 2944 8116
rect 2951 8110 2954 8116
rect 2972 8115 2973 8119
rect 2977 8115 2980 8118
rect 2999 8116 3000 8120
rect 3015 8119 3018 8124
rect 3047 8124 3058 8127
rect 3070 8125 3078 8128
rect 2972 8110 2975 8115
rect 2997 8110 3000 8116
rect 3047 8118 3050 8124
rect 3070 8119 3073 8125
rect 3082 8120 3085 8123
rect 3093 8123 3096 8137
rect 3144 8132 3147 8137
rect 3159 8139 3162 8149
rect 3189 8145 3192 8149
rect 3128 8128 3129 8131
rect 3133 8128 3136 8131
rect 3751 8142 3811 8146
rect 3815 8142 3827 8146
rect 3831 8142 3858 8146
rect 3862 8142 3880 8146
rect 3884 8142 3945 8146
rect 3949 8142 3963 8146
rect 3999 8139 4002 8149
rect 4029 8145 4032 8149
rect 4080 8145 4083 8149
rect 3175 8128 3178 8131
rect 3101 8123 3106 8128
rect 3144 8123 3147 8128
rect 3093 8120 3101 8123
rect 3015 8110 3018 8115
rect 3093 8115 3096 8120
rect 3152 8124 3163 8127
rect 3175 8125 3183 8128
rect 3045 8109 3050 8114
rect 2917 8097 2918 8101
rect 2942 8098 2943 8102
rect 2989 8097 2990 8101
rect 2794 8090 2870 8094
rect 2874 8090 2929 8094
rect 2933 8090 2954 8094
rect 2958 8090 2985 8094
rect 2989 8090 3018 8094
rect 617 8085 618 8089
rect 622 8085 623 8089
rect 627 8085 628 8089
rect 632 8085 633 8089
rect 637 8085 638 8089
rect 642 8085 643 8089
rect 613 8084 647 8085
rect 617 8080 618 8084
rect 622 8080 623 8084
rect 627 8080 628 8084
rect 632 8080 633 8084
rect 637 8080 638 8084
rect 642 8080 643 8084
rect 613 8079 647 8080
rect 617 8075 618 8079
rect 622 8075 623 8079
rect 627 8075 628 8079
rect 632 8075 633 8079
rect 637 8075 638 8079
rect 642 8075 643 8079
rect 613 8074 647 8075
rect 86 8068 346 8071
rect 617 8070 618 8074
rect 622 8070 623 8074
rect 627 8070 628 8074
rect 632 8070 633 8074
rect 637 8070 638 8074
rect 642 8070 643 8074
rect 663 8085 664 8089
rect 668 8085 669 8089
rect 673 8085 674 8089
rect 678 8085 679 8089
rect 683 8085 684 8089
rect 688 8085 689 8089
rect 3054 8087 3057 8115
rect 3084 8087 3087 8111
rect 3135 8087 3138 8119
rect 3152 8118 3155 8124
rect 3175 8119 3178 8125
rect 3187 8120 3190 8123
rect 3198 8123 3201 8137
rect 3870 8135 3873 8139
rect 3897 8135 3898 8139
rect 3942 8135 3944 8139
rect 3198 8120 3204 8123
rect 3198 8115 3201 8120
rect 3799 8115 3802 8118
rect 3810 8118 3813 8124
rect 3817 8118 3820 8124
rect 3810 8115 3820 8118
rect 3150 8109 3155 8114
rect 3159 8087 3162 8115
rect 3189 8087 3192 8111
rect 3810 8110 3813 8115
rect 3817 8110 3820 8115
rect 3826 8120 3829 8124
rect 3826 8116 3828 8120
rect 3832 8116 3834 8120
rect 3842 8119 3845 8124
rect 3870 8121 3873 8124
rect 3842 8117 3853 8119
rect 3826 8110 3829 8116
rect 3842 8115 3848 8117
rect 3842 8110 3845 8115
rect 3852 8115 3853 8117
rect 3871 8117 3873 8121
rect 3870 8110 3873 8117
rect 4015 8128 4018 8131
rect 3886 8120 3889 8124
rect 3896 8120 3899 8124
rect 3896 8116 3905 8120
rect 3917 8119 3920 8124
rect 3942 8120 3945 8124
rect 3886 8110 3889 8116
rect 3896 8110 3899 8116
rect 3917 8115 3918 8119
rect 3922 8115 3925 8118
rect 3944 8116 3945 8120
rect 3960 8119 3963 8124
rect 3992 8124 4003 8127
rect 4015 8125 4023 8128
rect 3917 8110 3920 8115
rect 3942 8110 3945 8116
rect 3992 8118 3995 8124
rect 4015 8119 4018 8125
rect 4027 8120 4030 8123
rect 4038 8123 4041 8137
rect 4089 8132 4092 8137
rect 4104 8139 4107 8149
rect 4134 8145 4137 8149
rect 4073 8128 4074 8131
rect 4078 8128 4081 8131
rect 4120 8128 4123 8131
rect 4046 8123 4051 8128
rect 4089 8123 4092 8128
rect 4038 8120 4046 8123
rect 3960 8110 3963 8115
rect 4038 8115 4041 8120
rect 4097 8124 4108 8127
rect 4120 8125 4128 8128
rect 3990 8109 3995 8114
rect 3862 8097 3863 8101
rect 3887 8098 3888 8102
rect 3934 8097 3935 8101
rect 3739 8090 3815 8094
rect 3819 8090 3874 8094
rect 3878 8090 3899 8094
rect 3903 8090 3930 8094
rect 3934 8090 3963 8094
rect 3999 8087 4002 8115
rect 4029 8087 4032 8111
rect 4080 8087 4083 8119
rect 4097 8118 4100 8124
rect 4120 8119 4123 8125
rect 4132 8120 4135 8123
rect 4143 8123 4146 8137
rect 4826 8135 4829 8174
rect 5083 8135 5086 8389
rect 4483 8129 4484 8133
rect 4488 8129 4489 8133
rect 4493 8129 4494 8133
rect 4498 8129 4499 8133
rect 4503 8129 4504 8133
rect 4508 8129 4509 8133
rect 4479 8128 4513 8129
rect 4483 8124 4484 8128
rect 4488 8124 4489 8128
rect 4493 8124 4494 8128
rect 4498 8124 4499 8128
rect 4503 8124 4504 8128
rect 4508 8124 4509 8128
rect 4143 8120 4149 8123
rect 4479 8123 4513 8124
rect 4143 8115 4146 8120
rect 4095 8109 4100 8114
rect 4104 8087 4107 8115
rect 4483 8119 4484 8123
rect 4488 8119 4489 8123
rect 4493 8119 4494 8123
rect 4498 8119 4499 8123
rect 4503 8119 4504 8123
rect 4508 8119 4509 8123
rect 4479 8118 4513 8119
rect 4483 8114 4484 8118
rect 4488 8114 4489 8118
rect 4493 8114 4494 8118
rect 4498 8114 4499 8118
rect 4503 8114 4504 8118
rect 4508 8114 4509 8118
rect 4529 8129 4530 8133
rect 4534 8129 4535 8133
rect 4539 8129 4540 8133
rect 4544 8129 4545 8133
rect 4549 8129 4550 8133
rect 4554 8129 4555 8133
rect 4826 8132 5086 8135
rect 4525 8128 4559 8129
rect 4529 8124 4530 8128
rect 4534 8124 4535 8128
rect 4539 8124 4540 8128
rect 4544 8124 4545 8128
rect 4549 8124 4550 8128
rect 4554 8124 4555 8128
rect 4525 8123 4559 8124
rect 4529 8119 4530 8123
rect 4534 8119 4535 8123
rect 4539 8119 4540 8123
rect 4544 8119 4545 8123
rect 4549 8119 4550 8123
rect 4554 8119 4555 8123
rect 4525 8118 4559 8119
rect 4529 8114 4530 8118
rect 4534 8114 4535 8118
rect 4539 8114 4540 8118
rect 4544 8114 4545 8118
rect 4549 8114 4550 8118
rect 4554 8114 4555 8118
rect 4134 8087 4137 8111
rect 4483 8098 4484 8102
rect 4488 8098 4489 8102
rect 4493 8098 4494 8102
rect 4498 8098 4499 8102
rect 4503 8098 4504 8102
rect 4508 8098 4509 8102
rect 4479 8097 4513 8098
rect 4483 8093 4484 8097
rect 4488 8093 4489 8097
rect 4493 8093 4494 8097
rect 4498 8093 4499 8097
rect 4503 8093 4504 8097
rect 4508 8093 4509 8097
rect 4479 8092 4513 8093
rect 4483 8088 4484 8092
rect 4488 8088 4489 8092
rect 4493 8088 4494 8092
rect 4498 8088 4499 8092
rect 4503 8088 4504 8092
rect 4508 8088 4509 8092
rect 4479 8087 4513 8088
rect 659 8084 693 8085
rect 663 8080 664 8084
rect 668 8080 669 8084
rect 673 8080 674 8084
rect 678 8080 679 8084
rect 683 8080 684 8084
rect 688 8080 689 8084
rect 2782 8083 2856 8087
rect 2860 8083 2862 8087
rect 2866 8083 2870 8087
rect 2874 8083 2888 8087
rect 2892 8083 2897 8087
rect 2901 8083 2906 8087
rect 2910 8083 2929 8087
rect 2933 8083 2963 8087
rect 2967 8083 2978 8087
rect 2982 8083 3006 8087
rect 3010 8083 3023 8087
rect 3027 8083 3047 8087
rect 3051 8083 3101 8087
rect 3105 8083 3128 8087
rect 3132 8083 3152 8087
rect 3156 8083 3204 8087
rect 3727 8083 3801 8087
rect 3805 8083 3807 8087
rect 3811 8083 3815 8087
rect 3819 8083 3833 8087
rect 3837 8083 3842 8087
rect 3846 8083 3851 8087
rect 3855 8083 3874 8087
rect 3878 8083 3908 8087
rect 3912 8083 3923 8087
rect 3927 8083 3951 8087
rect 3955 8083 3968 8087
rect 3972 8083 3992 8087
rect 3996 8083 4046 8087
rect 4050 8083 4073 8087
rect 4077 8083 4097 8087
rect 4101 8083 4149 8087
rect 4483 8083 4484 8087
rect 4488 8083 4489 8087
rect 4493 8083 4494 8087
rect 4498 8083 4499 8087
rect 4503 8083 4504 8087
rect 4508 8083 4509 8087
rect 4529 8098 4530 8102
rect 4534 8098 4535 8102
rect 4539 8098 4540 8102
rect 4544 8098 4545 8102
rect 4549 8098 4550 8102
rect 4554 8098 4555 8102
rect 4525 8097 4559 8098
rect 4529 8093 4530 8097
rect 4534 8093 4535 8097
rect 4539 8093 4540 8097
rect 4544 8093 4545 8097
rect 4549 8093 4550 8097
rect 4554 8093 4555 8097
rect 4525 8092 4559 8093
rect 4529 8088 4530 8092
rect 4534 8088 4535 8092
rect 4539 8088 4540 8092
rect 4544 8088 4545 8092
rect 4549 8088 4550 8092
rect 4554 8088 4555 8092
rect 4525 8087 4559 8088
rect 4529 8083 4530 8087
rect 4534 8083 4535 8087
rect 4539 8083 4540 8087
rect 4544 8083 4545 8087
rect 4549 8083 4550 8087
rect 4554 8083 4555 8087
rect 659 8079 693 8080
rect 663 8075 664 8079
rect 668 8075 669 8079
rect 673 8075 674 8079
rect 678 8075 679 8079
rect 683 8075 684 8079
rect 688 8075 689 8079
rect 2794 8076 2870 8080
rect 2874 8076 2929 8080
rect 2933 8076 2954 8080
rect 2958 8076 2985 8080
rect 2989 8076 3018 8080
rect 659 8074 693 8075
rect 663 8070 664 8074
rect 668 8070 669 8074
rect 673 8070 674 8074
rect 678 8070 679 8074
rect 683 8070 684 8074
rect 688 8070 689 8074
rect 2917 8069 2918 8073
rect 2942 8068 2943 8072
rect 2989 8069 2990 8073
rect 86 7814 89 8068
rect 343 8029 346 8068
rect 3054 8064 3057 8083
rect 3159 8064 3162 8083
rect 3739 8076 3815 8080
rect 3819 8076 3874 8080
rect 3878 8076 3899 8080
rect 3903 8076 3930 8080
rect 3934 8076 3963 8080
rect 3862 8069 3863 8073
rect 3887 8068 3888 8072
rect 3934 8069 3935 8073
rect 3999 8064 4002 8083
rect 4104 8064 4107 8083
rect 4826 8081 5086 8084
rect 4505 8078 4754 8080
rect 4505 8074 4506 8078
rect 4510 8074 4511 8078
rect 4515 8074 4754 8078
rect 4505 8073 4754 8074
rect 4505 8069 4506 8073
rect 4510 8069 4511 8073
rect 4515 8069 4754 8073
rect 4505 8068 4754 8069
rect 4505 8064 4506 8068
rect 4510 8064 4511 8068
rect 4515 8064 4754 8068
rect 2865 8055 2868 8060
rect 2872 8055 2875 8060
rect 2855 8052 2857 8055
rect 2865 8052 2875 8055
rect 2865 8046 2868 8052
rect 2872 8046 2875 8052
rect 2881 8054 2884 8060
rect 2897 8055 2900 8060
rect 2881 8050 2883 8054
rect 2887 8050 2889 8054
rect 2897 8053 2903 8055
rect 2907 8053 2908 8055
rect 2897 8051 2908 8053
rect 2925 8053 2928 8060
rect 2881 8046 2884 8050
rect 2897 8046 2900 8051
rect 2926 8049 2928 8053
rect 2925 8046 2928 8049
rect 2941 8054 2944 8060
rect 2951 8054 2954 8060
rect 2972 8055 2975 8060
rect 2951 8050 2960 8054
rect 2972 8051 2973 8055
rect 2977 8052 2980 8055
rect 2997 8054 3000 8060
rect 3015 8055 3018 8060
rect 2941 8046 2944 8050
rect 2951 8046 2954 8050
rect 2972 8046 2975 8051
rect 2999 8050 3000 8054
rect 3044 8051 3049 8056
rect 3053 8052 3055 8055
rect 3070 8054 3073 8060
rect 3070 8051 3078 8054
rect 3150 8051 3155 8056
rect 3159 8052 3160 8055
rect 3175 8054 3178 8060
rect 3175 8051 3183 8054
rect 3810 8055 3813 8060
rect 3817 8055 3820 8060
rect 3800 8052 3802 8055
rect 3810 8052 3820 8055
rect 2997 8046 3000 8050
rect 3015 8046 3018 8051
rect 3070 8048 3073 8051
rect 3175 8048 3178 8051
rect 3810 8046 3813 8052
rect 2925 8031 2928 8035
rect 2952 8031 2953 8035
rect 2997 8031 2999 8035
rect 343 8019 356 8029
rect 2806 8024 2882 8028
rect 2886 8024 2913 8028
rect 2917 8024 2935 8028
rect 2939 8024 3000 8028
rect 3004 8024 3018 8028
rect 3054 8021 3057 8040
rect 3159 8021 3162 8040
rect 3817 8046 3820 8052
rect 3826 8054 3829 8060
rect 3842 8055 3845 8060
rect 3826 8050 3828 8054
rect 3832 8050 3834 8054
rect 3842 8053 3848 8055
rect 3852 8053 3853 8055
rect 3842 8051 3853 8053
rect 3870 8053 3873 8060
rect 3826 8046 3829 8050
rect 3842 8046 3845 8051
rect 3871 8049 3873 8053
rect 3870 8046 3873 8049
rect 3886 8054 3889 8060
rect 3896 8054 3899 8060
rect 3917 8055 3920 8060
rect 3896 8050 3905 8054
rect 3917 8051 3918 8055
rect 3922 8052 3925 8055
rect 3942 8054 3945 8060
rect 3960 8055 3963 8060
rect 3886 8046 3889 8050
rect 3896 8046 3899 8050
rect 3917 8046 3920 8051
rect 3944 8050 3945 8054
rect 3989 8051 3994 8056
rect 3998 8052 4000 8055
rect 4015 8054 4018 8060
rect 4015 8051 4023 8054
rect 4095 8051 4100 8056
rect 4104 8052 4105 8055
rect 4120 8054 4123 8060
rect 4505 8063 4754 8064
rect 4505 8059 4506 8063
rect 4510 8059 4511 8063
rect 4515 8059 4754 8063
rect 4505 8058 4754 8059
rect 4120 8051 4128 8054
rect 4505 8054 4506 8058
rect 4510 8054 4511 8058
rect 4515 8054 4754 8058
rect 4505 8053 4754 8054
rect 3942 8046 3945 8050
rect 3960 8046 3963 8051
rect 4015 8048 4018 8051
rect 4120 8048 4123 8051
rect 4505 8049 4506 8053
rect 4510 8049 4511 8053
rect 4515 8049 4754 8053
rect 4505 8048 4754 8049
rect 4505 8044 4506 8048
rect 4510 8044 4511 8048
rect 4515 8044 4754 8048
rect 4505 8043 4754 8044
rect 3870 8031 3873 8035
rect 3897 8031 3898 8035
rect 3942 8031 3944 8035
rect 3751 8024 3827 8028
rect 3831 8024 3858 8028
rect 3862 8024 3880 8028
rect 3884 8024 3945 8028
rect 3949 8024 3963 8028
rect 3999 8021 4002 8040
rect 4104 8021 4107 8040
rect 4505 8039 4506 8043
rect 4510 8039 4511 8043
rect 4515 8039 4754 8043
rect 4826 8042 4829 8081
rect 4505 8038 4670 8039
rect 4505 8034 4506 8038
rect 4510 8034 4511 8038
rect 4515 8037 4670 8038
rect 4515 8034 4626 8037
rect 4645 8034 4649 8037
rect 4661 8034 4670 8037
rect 4688 8034 4692 8039
rect 4704 8034 4713 8039
rect 4729 8034 4733 8039
rect 4745 8034 4754 8039
rect 4505 8033 4626 8034
rect 4505 8029 4506 8033
rect 4510 8029 4511 8033
rect 4515 8029 4626 8033
rect 4505 8028 4626 8029
rect 4505 8024 4506 8028
rect 4510 8024 4511 8028
rect 4515 8024 4626 8028
rect 343 8009 366 8019
rect 2770 8017 2855 8021
rect 2859 8017 2871 8021
rect 2875 8017 2889 8021
rect 2893 8017 2900 8021
rect 2904 8017 2906 8021
rect 2910 8017 2925 8021
rect 2929 8017 2962 8021
rect 2966 8017 2967 8021
rect 2971 8017 2979 8021
rect 2983 8017 3007 8021
rect 3011 8017 3023 8021
rect 3027 8017 3047 8021
rect 3051 8017 3101 8021
rect 3105 8017 3128 8021
rect 3132 8017 3182 8021
rect 3186 8017 3190 8021
rect 3194 8017 3218 8021
rect 3222 8017 3272 8021
rect 3715 8017 3800 8021
rect 3804 8017 3816 8021
rect 3820 8017 3834 8021
rect 3838 8017 3845 8021
rect 3849 8017 3851 8021
rect 3855 8017 3870 8021
rect 3874 8017 3907 8021
rect 3911 8017 3912 8021
rect 3916 8017 3924 8021
rect 3928 8017 3952 8021
rect 3956 8017 3968 8021
rect 3972 8017 3992 8021
rect 3996 8017 4046 8021
rect 4050 8017 4073 8021
rect 4077 8017 4127 8021
rect 4131 8017 4135 8021
rect 4139 8017 4163 8021
rect 4167 8017 4217 8021
rect 2806 8010 2882 8014
rect 2886 8010 2913 8014
rect 2917 8010 2935 8014
rect 2939 8010 3000 8014
rect 3004 8010 3018 8014
rect 343 7999 376 8009
rect 3054 8007 3057 8017
rect 3084 8013 3087 8017
rect 3111 8013 3114 8017
rect 2925 8003 2928 8007
rect 2952 8003 2953 8007
rect 2997 8003 2999 8007
rect 343 7989 386 7999
rect 343 7893 769 7989
rect 2854 7983 2857 7986
rect 2865 7986 2868 7992
rect 2872 7986 2875 7992
rect 2865 7983 2875 7986
rect 2865 7978 2868 7983
rect 2872 7978 2875 7983
rect 2881 7988 2884 7992
rect 2881 7984 2883 7988
rect 2887 7984 2889 7988
rect 2897 7987 2900 7992
rect 2925 7989 2928 7992
rect 2897 7985 2908 7987
rect 2881 7978 2884 7984
rect 2897 7983 2903 7985
rect 2897 7978 2900 7983
rect 2907 7983 2908 7985
rect 2926 7985 2928 7989
rect 2925 7978 2928 7985
rect 3070 7996 3073 7999
rect 2941 7988 2944 7992
rect 2951 7988 2954 7992
rect 2951 7984 2960 7988
rect 2972 7987 2975 7992
rect 2997 7988 3000 7992
rect 2941 7978 2944 7984
rect 2951 7978 2954 7984
rect 2972 7983 2973 7987
rect 2977 7983 2980 7986
rect 2999 7984 3000 7988
rect 3015 7987 3018 7992
rect 3047 7992 3058 7995
rect 3070 7993 3078 7996
rect 2972 7978 2975 7983
rect 2997 7978 3000 7984
rect 3047 7986 3050 7992
rect 3070 7987 3073 7993
rect 3082 7988 3085 7991
rect 3093 7991 3096 8005
rect 3120 8000 3123 8005
rect 3135 8007 3138 8017
rect 3165 8013 3168 8017
rect 3201 8013 3204 8017
rect 3104 7996 3105 7999
rect 3109 7996 3112 7999
rect 3151 7996 3154 7999
rect 3093 7988 3101 7991
rect 3120 7991 3123 7996
rect 3015 7978 3018 7983
rect 3093 7983 3096 7988
rect 3101 7984 3105 7988
rect 3128 7992 3139 7995
rect 3151 7993 3159 7996
rect 3045 7977 3050 7982
rect 2917 7965 2918 7969
rect 2942 7966 2943 7970
rect 2989 7965 2990 7969
rect 2794 7958 2870 7962
rect 2874 7958 2929 7962
rect 2933 7958 2954 7962
rect 2958 7958 2985 7962
rect 2989 7958 3018 7962
rect 3054 7955 3057 7983
rect 3084 7955 3087 7979
rect 3111 7955 3114 7987
rect 3128 7986 3131 7992
rect 3151 7987 3154 7993
rect 3163 7988 3166 7991
rect 3174 7991 3177 8005
rect 3210 8000 3213 8005
rect 3225 8007 3228 8017
rect 3255 8013 3258 8017
rect 3199 7996 3202 7999
rect 3751 8010 3827 8014
rect 3831 8010 3858 8014
rect 3862 8010 3880 8014
rect 3884 8010 3945 8014
rect 3949 8010 3963 8014
rect 3999 8007 4002 8017
rect 4029 8013 4032 8017
rect 4056 8013 4059 8017
rect 3241 7996 3244 7999
rect 3174 7988 3183 7991
rect 3210 7991 3213 7996
rect 3174 7983 3177 7988
rect 3126 7977 3131 7982
rect 3135 7955 3138 7983
rect 3217 7994 3229 7995
rect 3221 7992 3229 7994
rect 3241 7993 3249 7996
rect 3241 7987 3244 7993
rect 3253 7988 3256 7991
rect 3264 7991 3267 8005
rect 3870 8003 3873 8007
rect 3897 8003 3898 8007
rect 3942 8003 3944 8007
rect 3264 7988 3284 7991
rect 3165 7955 3168 7979
rect 3201 7955 3204 7987
rect 3264 7983 3267 7988
rect 3799 7983 3802 7986
rect 3810 7986 3813 7992
rect 3817 7986 3820 7992
rect 3810 7983 3820 7986
rect 3225 7955 3228 7983
rect 3255 7955 3258 7979
rect 3810 7978 3813 7983
rect 3817 7978 3820 7983
rect 3826 7988 3829 7992
rect 3826 7984 3828 7988
rect 3832 7984 3834 7988
rect 3842 7987 3845 7992
rect 3870 7989 3873 7992
rect 3842 7985 3853 7987
rect 3826 7978 3829 7984
rect 3842 7983 3848 7985
rect 3842 7978 3845 7983
rect 3852 7983 3853 7985
rect 3871 7985 3873 7989
rect 3870 7978 3873 7985
rect 4015 7996 4018 7999
rect 3886 7988 3889 7992
rect 3896 7988 3899 7992
rect 3896 7984 3905 7988
rect 3917 7987 3920 7992
rect 3942 7988 3945 7992
rect 3886 7978 3889 7984
rect 3896 7978 3899 7984
rect 3917 7983 3918 7987
rect 3922 7983 3925 7986
rect 3944 7984 3945 7988
rect 3960 7987 3963 7992
rect 3992 7992 4003 7995
rect 4015 7993 4023 7996
rect 3917 7978 3920 7983
rect 3942 7978 3945 7984
rect 3992 7986 3995 7992
rect 4015 7987 4018 7993
rect 4027 7988 4030 7991
rect 4038 7991 4041 8005
rect 4065 8000 4068 8005
rect 4080 8007 4083 8017
rect 4110 8013 4113 8017
rect 4146 8013 4149 8017
rect 4049 7996 4050 7999
rect 4054 7996 4057 7999
rect 4096 7996 4099 7999
rect 4038 7988 4046 7991
rect 4065 7991 4068 7996
rect 3960 7978 3963 7983
rect 4038 7983 4041 7988
rect 4046 7984 4050 7988
rect 4073 7992 4084 7995
rect 4096 7993 4104 7996
rect 3990 7977 3995 7982
rect 3862 7965 3863 7969
rect 3887 7966 3888 7970
rect 3934 7965 3935 7969
rect 3739 7958 3815 7962
rect 3819 7958 3874 7962
rect 3878 7958 3899 7962
rect 3903 7958 3930 7962
rect 3934 7958 3963 7962
rect 3999 7955 4002 7983
rect 4029 7955 4032 7979
rect 4056 7955 4059 7987
rect 4073 7986 4076 7992
rect 4096 7987 4099 7993
rect 4108 7988 4111 7991
rect 4119 7991 4122 8005
rect 4155 8000 4158 8005
rect 4170 8007 4173 8017
rect 4200 8013 4203 8017
rect 4574 8015 4578 8024
rect 4590 8015 4594 8024
rect 4606 8015 4610 8024
rect 4622 8015 4626 8024
rect 4144 7996 4147 7999
rect 4186 7996 4189 7999
rect 4119 7988 4128 7991
rect 4155 7991 4158 7996
rect 4119 7983 4122 7988
rect 4071 7977 4076 7982
rect 4080 7955 4083 7983
rect 4162 7994 4174 7995
rect 4166 7992 4174 7994
rect 4186 7993 4194 7996
rect 4186 7987 4189 7993
rect 4198 7988 4201 7991
rect 4209 7991 4212 8005
rect 4209 7988 4229 7991
rect 4110 7955 4113 7979
rect 4146 7955 4149 7987
rect 4209 7983 4212 7988
rect 4170 7955 4173 7983
rect 4200 7955 4203 7979
rect 4626 7975 4627 8015
rect 4665 7975 4666 8034
rect 4582 7963 4586 7975
rect 4598 7972 4602 7975
rect 4614 7972 4618 7975
rect 4598 7968 4618 7972
rect 4637 7972 4641 7975
rect 4653 7972 4657 7975
rect 4637 7968 4657 7972
rect 4680 7974 4684 7975
rect 4708 7975 4709 8034
rect 4749 7975 4750 8034
rect 4816 8032 4829 8042
rect 4806 8022 4829 8032
rect 4796 8012 4829 8022
rect 4786 8002 4829 8012
rect 4696 7974 4700 7975
rect 4680 7972 4700 7974
rect 4721 7972 4741 7975
rect 4680 7970 4741 7972
rect 4774 7970 4829 8002
rect 2782 7951 2856 7955
rect 2860 7951 2862 7955
rect 2866 7951 2870 7955
rect 2874 7951 2888 7955
rect 2892 7951 2897 7955
rect 2901 7951 2906 7955
rect 2910 7951 2929 7955
rect 2933 7951 2963 7955
rect 2967 7951 2978 7955
rect 2982 7951 3006 7955
rect 3010 7951 3023 7955
rect 3027 7951 3047 7955
rect 3051 7951 3101 7955
rect 3108 7951 3128 7955
rect 3132 7951 3182 7955
rect 3186 7951 3218 7955
rect 3222 7951 3272 7955
rect 3727 7951 3801 7955
rect 3805 7951 3807 7955
rect 3811 7951 3815 7955
rect 3819 7951 3833 7955
rect 3837 7951 3842 7955
rect 3846 7951 3851 7955
rect 3855 7951 3874 7955
rect 3878 7951 3908 7955
rect 3912 7951 3923 7955
rect 3927 7951 3951 7955
rect 3955 7951 3968 7955
rect 3972 7951 3992 7955
rect 3996 7951 4046 7955
rect 4053 7951 4073 7955
rect 4077 7951 4127 7955
rect 4131 7951 4163 7955
rect 4167 7951 4217 7955
rect 2794 7944 2870 7948
rect 2874 7944 2929 7948
rect 2933 7944 2954 7948
rect 2958 7944 2985 7948
rect 2989 7944 3018 7948
rect 2917 7937 2918 7941
rect 2942 7936 2943 7940
rect 2989 7937 2990 7941
rect 2865 7923 2868 7928
rect 2872 7923 2875 7928
rect 2855 7920 2857 7923
rect 2865 7920 2875 7923
rect 2865 7914 2868 7920
rect 2872 7914 2875 7920
rect 2881 7922 2884 7928
rect 2897 7923 2900 7928
rect 2881 7918 2883 7922
rect 2887 7918 2889 7922
rect 2897 7921 2903 7923
rect 2907 7921 2908 7923
rect 2897 7919 2908 7921
rect 2925 7921 2928 7928
rect 2881 7914 2884 7918
rect 2897 7914 2900 7919
rect 2926 7917 2928 7921
rect 2925 7914 2928 7917
rect 2941 7922 2944 7928
rect 2951 7922 2954 7928
rect 2972 7923 2975 7928
rect 2951 7918 2960 7922
rect 2972 7919 2973 7923
rect 2977 7920 2980 7923
rect 2997 7922 3000 7928
rect 3015 7923 3018 7928
rect 3054 7929 3057 7951
rect 3135 7929 3138 7951
rect 3225 7929 3228 7951
rect 3739 7944 3815 7948
rect 3819 7944 3874 7948
rect 3878 7944 3899 7948
rect 3903 7944 3930 7948
rect 3934 7944 3963 7948
rect 3862 7937 3863 7941
rect 3887 7936 3888 7940
rect 3934 7937 3935 7941
rect 2941 7914 2944 7918
rect 2951 7914 2954 7918
rect 2972 7914 2975 7919
rect 2999 7918 3000 7922
rect 2997 7914 3000 7918
rect 3015 7914 3018 7919
rect 3045 7916 3050 7921
rect 3054 7917 3055 7920
rect 3070 7919 3073 7925
rect 3070 7916 3078 7919
rect 3125 7916 3130 7921
rect 3134 7917 3136 7920
rect 3151 7919 3154 7925
rect 3151 7916 3159 7919
rect 3218 7917 3226 7920
rect 3241 7919 3244 7925
rect 3810 7923 3813 7928
rect 3817 7923 3820 7928
rect 3800 7920 3802 7923
rect 3241 7916 3249 7919
rect 3810 7920 3820 7923
rect 3070 7913 3073 7916
rect 3151 7913 3154 7916
rect 3241 7913 3244 7916
rect 3810 7914 3813 7920
rect 2925 7899 2928 7903
rect 2952 7899 2953 7903
rect 2997 7899 2999 7903
rect 3817 7914 3820 7920
rect 3826 7922 3829 7928
rect 3842 7923 3845 7928
rect 3826 7918 3828 7922
rect 3832 7918 3834 7922
rect 3842 7921 3848 7923
rect 3852 7921 3853 7923
rect 3842 7919 3853 7921
rect 3870 7921 3873 7928
rect 3826 7914 3829 7918
rect 3842 7914 3845 7919
rect 3871 7917 3873 7921
rect 3870 7914 3873 7917
rect 3886 7922 3889 7928
rect 3896 7922 3899 7928
rect 3917 7923 3920 7928
rect 3896 7918 3905 7922
rect 3917 7919 3918 7923
rect 3922 7920 3925 7923
rect 3942 7922 3945 7928
rect 3960 7923 3963 7928
rect 3999 7929 4002 7951
rect 4080 7929 4083 7951
rect 4170 7929 4173 7951
rect 4369 7950 4572 7963
rect 4582 7959 4593 7963
rect 4605 7963 4618 7968
rect 4648 7965 4657 7968
rect 4691 7966 4829 7970
rect 4648 7963 4678 7965
rect 4582 7945 4586 7959
rect 4605 7956 4635 7963
rect 4598 7950 4635 7956
rect 4639 7950 4640 7963
rect 4648 7954 4659 7963
rect 4667 7954 4678 7963
rect 4648 7952 4678 7954
rect 4682 7952 4683 7965
rect 4598 7949 4618 7950
rect 4598 7945 4602 7949
rect 4614 7945 4618 7949
rect 4648 7945 4657 7952
rect 4691 7945 4700 7966
rect 4721 7952 4829 7966
rect 4721 7945 4741 7952
rect 3886 7914 3889 7918
rect 3896 7914 3899 7918
rect 3917 7914 3920 7919
rect 3944 7918 3945 7922
rect 3942 7914 3945 7918
rect 3960 7914 3963 7919
rect 3990 7916 3995 7921
rect 3999 7917 4000 7920
rect 4015 7919 4018 7925
rect 4015 7916 4023 7919
rect 4070 7916 4075 7921
rect 4079 7917 4081 7920
rect 4096 7919 4099 7925
rect 4096 7916 4104 7919
rect 4163 7917 4171 7920
rect 4186 7919 4189 7925
rect 4186 7916 4194 7919
rect 4015 7913 4018 7916
rect 4096 7913 4099 7916
rect 4186 7913 4189 7916
rect 343 7883 386 7893
rect 2806 7892 2882 7896
rect 2886 7892 2913 7896
rect 2917 7892 2935 7896
rect 2939 7892 3000 7896
rect 3004 7892 3018 7896
rect 3054 7889 3057 7905
rect 3135 7889 3138 7905
rect 3225 7889 3228 7905
rect 3870 7899 3873 7903
rect 3897 7899 3898 7903
rect 3942 7899 3944 7903
rect 3751 7892 3827 7896
rect 3831 7892 3858 7896
rect 3862 7892 3880 7896
rect 3884 7892 3945 7896
rect 3949 7892 3963 7896
rect 3999 7889 4002 7905
rect 4080 7889 4083 7905
rect 4170 7889 4173 7905
rect 4626 7889 4627 7945
rect 2770 7885 2855 7889
rect 2859 7885 2871 7889
rect 2875 7885 2889 7889
rect 2893 7885 2900 7889
rect 2904 7885 2906 7889
rect 2910 7885 2925 7889
rect 2929 7885 2962 7889
rect 2966 7885 2967 7889
rect 2971 7885 2979 7889
rect 2983 7885 3007 7889
rect 3011 7885 3023 7889
rect 3027 7885 3047 7889
rect 3051 7885 3101 7889
rect 3105 7885 3128 7889
rect 3132 7885 3218 7889
rect 3222 7885 3276 7889
rect 3715 7885 3800 7889
rect 3804 7885 3816 7889
rect 3820 7885 3834 7889
rect 3838 7885 3845 7889
rect 3849 7885 3851 7889
rect 3855 7885 3870 7889
rect 3874 7885 3907 7889
rect 3911 7885 3912 7889
rect 3916 7885 3924 7889
rect 3928 7885 3952 7889
rect 3956 7885 3968 7889
rect 3972 7885 3992 7889
rect 3996 7885 4046 7889
rect 4050 7885 4073 7889
rect 4077 7885 4163 7889
rect 4167 7885 4221 7889
rect 4574 7886 4578 7889
rect 4590 7886 4594 7889
rect 4606 7886 4610 7889
rect 4622 7886 4626 7889
rect 343 7873 376 7883
rect 2806 7878 2882 7882
rect 2886 7878 2913 7882
rect 2917 7878 2935 7882
rect 2939 7878 3000 7882
rect 3004 7878 3018 7882
rect 3054 7875 3057 7885
rect 3084 7881 3087 7885
rect 343 7863 366 7873
rect 2925 7871 2928 7875
rect 2952 7871 2953 7875
rect 2997 7871 2999 7875
rect 343 7853 356 7863
rect 343 7814 346 7853
rect 2854 7851 2857 7854
rect 2865 7854 2868 7860
rect 2872 7854 2875 7860
rect 2865 7851 2875 7854
rect 2865 7846 2868 7851
rect 2872 7846 2875 7851
rect 2881 7856 2884 7860
rect 2881 7852 2883 7856
rect 2887 7852 2889 7856
rect 2897 7855 2900 7860
rect 2925 7857 2928 7860
rect 2897 7853 2908 7855
rect 2881 7846 2884 7852
rect 2897 7851 2903 7853
rect 2897 7846 2900 7851
rect 2907 7851 2908 7853
rect 2926 7853 2928 7857
rect 2925 7846 2928 7853
rect 3751 7878 3827 7882
rect 3831 7878 3858 7882
rect 3862 7878 3880 7882
rect 3884 7878 3945 7882
rect 3949 7878 3963 7882
rect 3999 7875 4002 7885
rect 4029 7881 4032 7885
rect 3070 7864 3073 7867
rect 2941 7856 2944 7860
rect 2951 7856 2954 7860
rect 2951 7852 2960 7856
rect 2972 7855 2975 7860
rect 2997 7856 3000 7860
rect 2941 7846 2944 7852
rect 2951 7846 2954 7852
rect 2972 7851 2973 7855
rect 2977 7851 2980 7854
rect 2999 7852 3000 7856
rect 3015 7855 3018 7860
rect 3047 7860 3058 7863
rect 3070 7861 3078 7864
rect 2972 7846 2975 7851
rect 2997 7846 3000 7852
rect 3047 7854 3050 7860
rect 3070 7855 3073 7861
rect 3082 7856 3085 7859
rect 3093 7859 3096 7873
rect 3870 7871 3873 7875
rect 3897 7871 3898 7875
rect 3942 7871 3944 7875
rect 3101 7859 3106 7864
rect 3093 7856 3101 7859
rect 3015 7846 3018 7851
rect 3093 7851 3096 7856
rect 3799 7851 3802 7854
rect 3810 7854 3813 7860
rect 3817 7854 3820 7860
rect 3810 7851 3820 7854
rect 3045 7845 3050 7850
rect 2364 7830 2373 7834
rect 2377 7830 2409 7834
rect 2413 7830 2476 7834
rect 2480 7830 2505 7834
rect 2509 7830 2541 7834
rect 2545 7830 2608 7834
rect 2612 7830 2637 7834
rect 2641 7830 2673 7834
rect 2677 7830 2740 7834
rect 2744 7830 2824 7834
rect 2917 7833 2918 7837
rect 2942 7834 2943 7838
rect 2989 7833 2990 7837
rect 2364 7823 2397 7827
rect 2401 7823 2425 7827
rect 2429 7823 2455 7827
rect 2459 7823 2492 7827
rect 2496 7823 2529 7827
rect 2533 7823 2557 7827
rect 2561 7823 2587 7827
rect 2591 7823 2624 7827
rect 2628 7823 2661 7827
rect 2665 7823 2689 7827
rect 2693 7823 2719 7827
rect 2723 7823 2756 7827
rect 2760 7823 2764 7827
rect 2849 7826 2870 7830
rect 2874 7826 2879 7830
rect 2883 7826 2929 7830
rect 2933 7826 2954 7830
rect 2958 7826 2985 7830
rect 2989 7826 3018 7830
rect 3054 7823 3057 7851
rect 3084 7823 3087 7847
rect 3810 7846 3813 7851
rect 3817 7846 3820 7851
rect 3826 7856 3829 7860
rect 3826 7852 3828 7856
rect 3832 7852 3834 7856
rect 3842 7855 3845 7860
rect 3870 7857 3873 7860
rect 3842 7853 3853 7855
rect 3826 7846 3829 7852
rect 3842 7851 3848 7853
rect 3842 7846 3845 7851
rect 3852 7851 3853 7853
rect 3871 7853 3873 7857
rect 3870 7846 3873 7853
rect 4015 7864 4018 7867
rect 3886 7856 3889 7860
rect 3896 7856 3899 7860
rect 3896 7852 3905 7856
rect 3917 7855 3920 7860
rect 3942 7856 3945 7860
rect 3886 7846 3889 7852
rect 3896 7846 3899 7852
rect 3917 7851 3918 7855
rect 3922 7851 3925 7854
rect 3944 7852 3945 7856
rect 3960 7855 3963 7860
rect 3992 7860 4003 7863
rect 4015 7861 4023 7864
rect 3917 7846 3920 7851
rect 3942 7846 3945 7852
rect 3992 7854 3995 7860
rect 4015 7855 4018 7861
rect 4027 7856 4030 7859
rect 4038 7859 4041 7873
rect 4046 7859 4051 7864
rect 4038 7856 4046 7859
rect 3960 7846 3963 7851
rect 4038 7851 4041 7856
rect 3990 7845 3995 7850
rect 3309 7830 3318 7834
rect 3322 7830 3354 7834
rect 3358 7830 3421 7834
rect 3425 7830 3450 7834
rect 3454 7830 3486 7834
rect 3490 7830 3553 7834
rect 3557 7830 3582 7834
rect 3586 7830 3618 7834
rect 3622 7830 3685 7834
rect 3689 7830 3769 7834
rect 3862 7833 3863 7837
rect 3887 7834 3888 7838
rect 3934 7833 3935 7837
rect 3309 7823 3342 7827
rect 3346 7823 3370 7827
rect 3374 7823 3400 7827
rect 3404 7823 3437 7827
rect 3441 7823 3474 7827
rect 3478 7823 3502 7827
rect 3506 7823 3532 7827
rect 3536 7823 3569 7827
rect 3573 7823 3606 7827
rect 3610 7823 3634 7827
rect 3638 7823 3664 7827
rect 3668 7823 3701 7827
rect 3705 7823 3709 7827
rect 3794 7826 3815 7830
rect 3819 7826 3824 7830
rect 3828 7826 3874 7830
rect 3878 7826 3899 7830
rect 3903 7826 3930 7830
rect 3934 7826 3963 7830
rect 3999 7823 4002 7851
rect 4527 7854 4626 7886
rect 4641 7939 4653 7945
rect 4665 7857 4666 7945
rect 4684 7939 4696 7945
rect 4708 7857 4709 7945
rect 4725 7939 4737 7945
rect 4749 7857 4750 7945
rect 4774 7906 4829 7952
rect 4786 7896 4829 7906
rect 4796 7886 4829 7896
rect 4806 7876 4829 7886
rect 4816 7866 4829 7876
rect 4645 7854 4649 7857
rect 4661 7854 4670 7857
rect 4688 7854 4692 7857
rect 4704 7854 4713 7857
rect 4729 7854 4733 7857
rect 4745 7854 4754 7857
rect 4029 7823 4032 7847
rect 4527 7830 4754 7854
rect 4527 7828 4595 7830
rect 4527 7824 4529 7828
rect 4533 7824 4534 7828
rect 4538 7824 4539 7828
rect 4543 7824 4544 7828
rect 4548 7824 4549 7828
rect 4553 7824 4554 7828
rect 4558 7824 4559 7828
rect 4563 7824 4564 7828
rect 4568 7824 4569 7828
rect 4573 7824 4574 7828
rect 4578 7824 4579 7828
rect 4583 7824 4584 7828
rect 4588 7824 4589 7828
rect 4593 7824 4595 7828
rect 4826 7827 4829 7866
rect 5083 7827 5086 8081
rect 4826 7824 5086 7827
rect 4527 7823 4595 7824
rect 86 7811 346 7814
rect 2367 7813 2370 7823
rect 2388 7813 2391 7823
rect 2404 7813 2407 7823
rect 2418 7816 2423 7820
rect 2427 7816 2434 7820
rect 2446 7813 2449 7823
rect 2462 7813 2465 7823
rect 2483 7813 2486 7823
rect 2499 7813 2502 7823
rect 2520 7813 2523 7823
rect 2536 7813 2539 7823
rect 2550 7816 2555 7820
rect 2559 7816 2566 7820
rect 2578 7813 2581 7823
rect 2594 7813 2597 7823
rect 2615 7813 2618 7823
rect 2631 7813 2634 7823
rect 2652 7813 2655 7823
rect 2668 7813 2671 7823
rect 2682 7816 2687 7820
rect 2691 7816 2698 7820
rect 2710 7813 2713 7823
rect 2726 7813 2729 7823
rect 2747 7813 2750 7823
rect 2782 7819 2856 7823
rect 2860 7819 2862 7823
rect 2866 7819 2870 7823
rect 2874 7819 2888 7823
rect 2892 7819 2897 7823
rect 2901 7819 2906 7823
rect 2910 7819 2929 7823
rect 2933 7819 2963 7823
rect 2967 7819 2978 7823
rect 2982 7819 3006 7823
rect 3010 7819 3023 7823
rect 3027 7819 3047 7823
rect 3051 7819 3131 7823
rect 3135 7819 3149 7823
rect 3153 7819 3158 7823
rect 3162 7819 3167 7823
rect 3171 7819 3190 7823
rect 3194 7819 3224 7823
rect 3228 7819 3239 7823
rect 3243 7819 3267 7823
rect 3271 7819 3280 7823
rect 2384 7799 2389 7802
rect 2393 7799 2417 7802
rect 2442 7799 2449 7802
rect 2453 7799 2475 7802
rect 2495 7799 2502 7802
rect 2516 7799 2521 7802
rect 2525 7799 2549 7802
rect 2574 7799 2581 7802
rect 2585 7799 2607 7802
rect 2627 7799 2634 7802
rect 2648 7799 2653 7802
rect 2657 7799 2681 7802
rect 2794 7812 2870 7816
rect 2874 7812 2879 7816
rect 2883 7812 2929 7816
rect 2933 7812 2954 7816
rect 2958 7812 2985 7816
rect 2989 7812 3018 7816
rect 2706 7799 2713 7802
rect 2717 7799 2739 7802
rect 2917 7805 2918 7809
rect 2942 7804 2943 7808
rect 2989 7805 2990 7809
rect 2400 7789 2407 7792
rect 2411 7793 2430 7796
rect 2430 7786 2433 7792
rect 2458 7789 2465 7792
rect 2469 7793 2484 7796
rect 2532 7789 2539 7792
rect 2543 7793 2562 7796
rect 2562 7786 2565 7792
rect 2590 7789 2597 7792
rect 2601 7793 2616 7796
rect 2664 7789 2671 7792
rect 2675 7793 2694 7796
rect 2694 7786 2697 7792
rect 2722 7789 2729 7792
rect 2733 7793 2750 7796
rect 2865 7791 2868 7796
rect 2872 7791 2875 7796
rect 2855 7788 2857 7791
rect 2865 7788 2875 7791
rect 2865 7782 2868 7788
rect 617 7776 618 7780
rect 622 7776 623 7780
rect 627 7776 628 7780
rect 632 7776 633 7780
rect 637 7776 638 7780
rect 642 7776 643 7780
rect 613 7775 647 7776
rect 617 7771 618 7775
rect 622 7771 623 7775
rect 627 7771 628 7775
rect 632 7771 633 7775
rect 637 7771 638 7775
rect 642 7771 643 7775
rect 613 7770 647 7771
rect 617 7766 618 7770
rect 622 7766 623 7770
rect 627 7766 628 7770
rect 632 7766 633 7770
rect 637 7766 638 7770
rect 642 7766 643 7770
rect 613 7765 647 7766
rect 86 7759 346 7762
rect 617 7761 618 7765
rect 622 7761 623 7765
rect 627 7761 628 7765
rect 632 7761 633 7765
rect 637 7761 638 7765
rect 642 7761 643 7765
rect 663 7776 664 7780
rect 668 7776 669 7780
rect 673 7776 674 7780
rect 678 7776 679 7780
rect 683 7776 684 7780
rect 688 7776 689 7780
rect 659 7775 693 7776
rect 663 7771 664 7775
rect 668 7771 669 7775
rect 673 7771 674 7775
rect 678 7771 679 7775
rect 683 7771 684 7775
rect 688 7771 689 7775
rect 659 7770 693 7771
rect 2367 7770 2370 7782
rect 2388 7770 2391 7782
rect 2404 7770 2407 7782
rect 2418 7773 2430 7776
rect 2446 7770 2449 7782
rect 2462 7770 2465 7782
rect 2483 7770 2486 7782
rect 2499 7770 2502 7782
rect 2520 7770 2523 7782
rect 2536 7770 2539 7782
rect 2550 7773 2562 7776
rect 2578 7770 2581 7782
rect 2594 7770 2597 7782
rect 2615 7770 2618 7782
rect 2631 7770 2634 7782
rect 2652 7770 2655 7782
rect 2668 7770 2671 7782
rect 2682 7773 2694 7776
rect 2710 7770 2713 7782
rect 2726 7770 2729 7782
rect 2747 7770 2750 7782
rect 2872 7782 2875 7788
rect 2881 7790 2884 7796
rect 2897 7791 2900 7796
rect 2881 7786 2883 7790
rect 2887 7786 2889 7790
rect 2897 7789 2903 7791
rect 2907 7789 2908 7791
rect 2897 7787 2908 7789
rect 2925 7789 2928 7796
rect 2881 7782 2884 7786
rect 2897 7782 2900 7787
rect 2926 7785 2928 7789
rect 2925 7782 2928 7785
rect 2941 7790 2944 7796
rect 2951 7790 2954 7796
rect 2972 7791 2975 7796
rect 2951 7786 2960 7790
rect 2972 7787 2973 7791
rect 2977 7788 2980 7791
rect 2997 7790 3000 7796
rect 3015 7791 3018 7796
rect 3054 7793 3057 7819
rect 3090 7812 3109 7816
rect 3113 7812 3131 7816
rect 3135 7812 3190 7816
rect 3194 7812 3215 7816
rect 3219 7812 3246 7816
rect 3250 7812 3279 7816
rect 3312 7813 3315 7823
rect 3333 7813 3336 7823
rect 3349 7813 3352 7823
rect 3363 7816 3368 7820
rect 3372 7816 3379 7820
rect 3391 7813 3394 7823
rect 3407 7813 3410 7823
rect 3428 7813 3431 7823
rect 3444 7813 3447 7823
rect 3465 7813 3468 7823
rect 3481 7813 3484 7823
rect 3495 7816 3500 7820
rect 3504 7816 3511 7820
rect 3523 7813 3526 7823
rect 3539 7813 3542 7823
rect 3560 7813 3563 7823
rect 3576 7813 3579 7823
rect 3597 7813 3600 7823
rect 3613 7813 3616 7823
rect 3627 7816 3632 7820
rect 3636 7816 3643 7820
rect 3655 7813 3658 7823
rect 3671 7813 3674 7823
rect 3692 7813 3695 7823
rect 3727 7819 3801 7823
rect 3805 7819 3807 7823
rect 3811 7819 3815 7823
rect 3819 7819 3833 7823
rect 3837 7819 3842 7823
rect 3846 7819 3851 7823
rect 3855 7819 3874 7823
rect 3878 7819 3908 7823
rect 3912 7819 3923 7823
rect 3927 7819 3951 7823
rect 3955 7819 3968 7823
rect 3972 7819 3992 7823
rect 3996 7819 4076 7823
rect 4080 7819 4094 7823
rect 4098 7819 4103 7823
rect 4107 7819 4112 7823
rect 4116 7819 4135 7823
rect 4139 7819 4169 7823
rect 4173 7819 4184 7823
rect 4188 7819 4212 7823
rect 4216 7819 4225 7823
rect 4527 7819 4529 7823
rect 4533 7819 4534 7823
rect 4538 7819 4539 7823
rect 4543 7819 4544 7823
rect 4548 7819 4549 7823
rect 4553 7819 4554 7823
rect 4558 7819 4559 7823
rect 4563 7819 4564 7823
rect 4568 7819 4569 7823
rect 4573 7819 4574 7823
rect 4578 7819 4579 7823
rect 4583 7819 4584 7823
rect 4588 7819 4589 7823
rect 4593 7819 4595 7823
rect 3090 7800 3093 7812
rect 3178 7805 3179 7809
rect 3203 7804 3204 7808
rect 3250 7805 3251 7809
rect 2941 7782 2944 7786
rect 2951 7782 2954 7786
rect 2972 7782 2975 7787
rect 2999 7786 3000 7790
rect 3117 7791 3120 7796
rect 3126 7791 3129 7796
rect 3133 7791 3136 7796
rect 2997 7782 3000 7786
rect 3015 7782 3018 7787
rect 3044 7780 3049 7785
rect 3053 7781 3055 7784
rect 3070 7783 3073 7789
rect 3102 7788 3136 7791
rect 3070 7780 3078 7783
rect 3070 7777 3073 7780
rect 663 7766 664 7770
rect 668 7766 669 7770
rect 673 7766 674 7770
rect 678 7766 679 7770
rect 683 7766 684 7770
rect 688 7766 689 7770
rect 2364 7766 2397 7770
rect 2401 7766 2425 7770
rect 2429 7766 2455 7770
rect 2459 7766 2529 7770
rect 2533 7766 2557 7770
rect 2561 7766 2587 7770
rect 2591 7766 2661 7770
rect 2665 7766 2689 7770
rect 2693 7766 2719 7770
rect 2723 7766 2776 7770
rect 2925 7767 2928 7771
rect 2952 7767 2953 7771
rect 2997 7767 2999 7771
rect 3102 7774 3105 7788
rect 3126 7782 3129 7788
rect 3133 7782 3136 7788
rect 3142 7790 3145 7796
rect 3158 7791 3161 7796
rect 3142 7786 3144 7790
rect 3148 7786 3150 7790
rect 3158 7789 3164 7791
rect 3168 7789 3169 7791
rect 3158 7787 3169 7789
rect 3186 7789 3189 7796
rect 3142 7782 3145 7786
rect 3158 7782 3161 7787
rect 3187 7785 3189 7789
rect 3186 7782 3189 7785
rect 3329 7799 3334 7802
rect 3338 7799 3362 7802
rect 3387 7799 3394 7802
rect 3398 7799 3420 7802
rect 3440 7799 3447 7802
rect 3461 7799 3466 7802
rect 3470 7799 3494 7802
rect 3519 7799 3526 7802
rect 3530 7799 3552 7802
rect 3572 7799 3579 7802
rect 3593 7799 3598 7802
rect 3602 7799 3626 7802
rect 3739 7812 3815 7816
rect 3819 7812 3824 7816
rect 3828 7812 3874 7816
rect 3878 7812 3899 7816
rect 3903 7812 3930 7816
rect 3934 7812 3963 7816
rect 3651 7799 3658 7802
rect 3662 7799 3684 7802
rect 3862 7805 3863 7809
rect 3887 7804 3888 7808
rect 3934 7805 3935 7809
rect 3202 7790 3205 7796
rect 3212 7790 3215 7796
rect 3233 7791 3236 7796
rect 3212 7786 3221 7790
rect 3233 7787 3234 7791
rect 3238 7788 3241 7791
rect 3258 7790 3261 7796
rect 3276 7791 3279 7796
rect 3202 7782 3205 7786
rect 3212 7782 3215 7786
rect 3233 7782 3236 7787
rect 3260 7786 3261 7790
rect 3258 7782 3261 7786
rect 3276 7782 3279 7787
rect 3345 7789 3352 7792
rect 3356 7793 3375 7796
rect 3375 7786 3378 7792
rect 3403 7789 3410 7792
rect 3414 7793 3429 7796
rect 3477 7789 3484 7792
rect 3488 7793 3507 7796
rect 3507 7786 3510 7792
rect 3535 7789 3542 7792
rect 3546 7793 3561 7796
rect 3609 7789 3616 7792
rect 3620 7793 3639 7796
rect 3639 7786 3642 7792
rect 3667 7789 3674 7792
rect 3678 7793 3695 7796
rect 3810 7791 3813 7796
rect 3817 7791 3820 7796
rect 3800 7788 3802 7791
rect 3810 7788 3820 7791
rect 3810 7782 3813 7788
rect 659 7765 693 7766
rect 663 7761 664 7765
rect 668 7761 669 7765
rect 673 7761 674 7765
rect 678 7761 679 7765
rect 683 7761 684 7765
rect 688 7761 689 7765
rect 2364 7759 2373 7763
rect 2377 7759 2424 7763
rect 2428 7759 2474 7763
rect 2478 7759 2505 7763
rect 2509 7759 2556 7763
rect 2560 7759 2606 7763
rect 2610 7759 2637 7763
rect 2641 7759 2688 7763
rect 2692 7759 2738 7763
rect 2742 7760 2812 7763
rect 2868 7760 2882 7764
rect 2886 7760 2913 7764
rect 2917 7760 2935 7764
rect 2939 7760 3000 7764
rect 3004 7760 3018 7764
rect 86 7505 89 7759
rect 343 7720 346 7759
rect 3054 7757 3057 7769
rect 3186 7767 3189 7771
rect 3213 7767 3214 7771
rect 3258 7767 3260 7771
rect 3312 7770 3315 7782
rect 3333 7770 3336 7782
rect 3349 7770 3352 7782
rect 3363 7773 3375 7776
rect 3391 7770 3394 7782
rect 3407 7770 3410 7782
rect 3428 7770 3431 7782
rect 3444 7770 3447 7782
rect 3465 7770 3468 7782
rect 3481 7770 3484 7782
rect 3495 7773 3507 7776
rect 3523 7770 3526 7782
rect 3539 7770 3542 7782
rect 3560 7770 3563 7782
rect 3576 7770 3579 7782
rect 3597 7770 3600 7782
rect 3613 7770 3616 7782
rect 3627 7773 3639 7776
rect 3655 7770 3658 7782
rect 3671 7770 3674 7782
rect 3692 7770 3695 7782
rect 3817 7782 3820 7788
rect 3826 7790 3829 7796
rect 3842 7791 3845 7796
rect 3826 7786 3828 7790
rect 3832 7786 3834 7790
rect 3842 7789 3848 7791
rect 3852 7789 3853 7791
rect 3842 7787 3853 7789
rect 3870 7789 3873 7796
rect 3826 7782 3829 7786
rect 3842 7782 3845 7787
rect 3871 7785 3873 7789
rect 3870 7782 3873 7785
rect 3886 7790 3889 7796
rect 3896 7790 3899 7796
rect 3917 7791 3920 7796
rect 3896 7786 3905 7790
rect 3917 7787 3918 7791
rect 3922 7788 3925 7791
rect 3942 7790 3945 7796
rect 3960 7791 3963 7796
rect 3999 7793 4002 7819
rect 4527 7818 4595 7819
rect 4035 7812 4054 7816
rect 4058 7812 4076 7816
rect 4080 7812 4135 7816
rect 4139 7812 4160 7816
rect 4164 7812 4191 7816
rect 4195 7812 4224 7816
rect 4035 7800 4038 7812
rect 4123 7805 4124 7809
rect 4148 7804 4149 7808
rect 4195 7805 4196 7809
rect 3886 7782 3889 7786
rect 3896 7782 3899 7786
rect 3917 7782 3920 7787
rect 3944 7786 3945 7790
rect 4062 7791 4065 7796
rect 4071 7791 4074 7796
rect 4078 7791 4081 7796
rect 3942 7782 3945 7786
rect 3960 7782 3963 7787
rect 3989 7780 3994 7785
rect 3998 7781 4000 7784
rect 4015 7783 4018 7789
rect 4047 7788 4081 7791
rect 4015 7780 4023 7783
rect 4015 7777 4018 7780
rect 3309 7766 3342 7770
rect 3346 7766 3370 7770
rect 3374 7766 3400 7770
rect 3404 7766 3474 7770
rect 3478 7766 3502 7770
rect 3506 7766 3532 7770
rect 3536 7766 3606 7770
rect 3610 7766 3634 7770
rect 3638 7766 3664 7770
rect 3668 7766 3721 7770
rect 3870 7767 3873 7771
rect 3897 7767 3898 7771
rect 3942 7767 3944 7771
rect 4047 7774 4050 7788
rect 4071 7782 4074 7788
rect 4078 7782 4081 7788
rect 4087 7790 4090 7796
rect 4103 7791 4106 7796
rect 4087 7786 4089 7790
rect 4093 7786 4095 7790
rect 4103 7789 4109 7791
rect 4113 7789 4114 7791
rect 4103 7787 4114 7789
rect 4131 7789 4134 7796
rect 4087 7782 4090 7786
rect 4103 7782 4106 7787
rect 4132 7785 4134 7789
rect 4131 7782 4134 7785
rect 4147 7790 4150 7796
rect 4157 7790 4160 7796
rect 4178 7791 4181 7796
rect 4157 7786 4166 7790
rect 4178 7787 4179 7791
rect 4183 7788 4186 7791
rect 4203 7790 4206 7796
rect 4221 7791 4224 7796
rect 4147 7782 4150 7786
rect 4157 7782 4160 7786
rect 4178 7782 4181 7787
rect 4205 7786 4206 7790
rect 4483 7789 4484 7793
rect 4488 7789 4489 7793
rect 4493 7789 4494 7793
rect 4498 7789 4499 7793
rect 4503 7789 4504 7793
rect 4508 7789 4509 7793
rect 4479 7788 4513 7789
rect 4203 7782 4206 7786
rect 4221 7782 4224 7787
rect 4483 7784 4484 7788
rect 4488 7784 4489 7788
rect 4493 7784 4494 7788
rect 4498 7784 4499 7788
rect 4503 7784 4504 7788
rect 4508 7784 4509 7788
rect 4479 7783 4513 7784
rect 4483 7779 4484 7783
rect 4488 7779 4489 7783
rect 4493 7779 4494 7783
rect 4498 7779 4499 7783
rect 4503 7779 4504 7783
rect 4508 7779 4509 7783
rect 4479 7778 4513 7779
rect 4483 7774 4484 7778
rect 4488 7774 4489 7778
rect 4493 7774 4494 7778
rect 4498 7774 4499 7778
rect 4503 7774 4504 7778
rect 4508 7774 4509 7778
rect 4529 7789 4530 7793
rect 4534 7789 4535 7793
rect 4539 7789 4540 7793
rect 4544 7789 4545 7793
rect 4549 7789 4550 7793
rect 4554 7789 4555 7793
rect 4525 7788 4559 7789
rect 4529 7784 4530 7788
rect 4534 7784 4535 7788
rect 4539 7784 4540 7788
rect 4544 7784 4545 7788
rect 4549 7784 4550 7788
rect 4554 7784 4555 7788
rect 4525 7783 4559 7784
rect 4529 7779 4530 7783
rect 4534 7779 4535 7783
rect 4539 7779 4540 7783
rect 4544 7779 4545 7783
rect 4549 7779 4550 7783
rect 4554 7779 4555 7783
rect 4525 7778 4559 7779
rect 4529 7774 4530 7778
rect 4534 7774 4535 7778
rect 4539 7774 4540 7778
rect 4544 7774 4545 7778
rect 4549 7774 4550 7778
rect 4554 7774 4555 7778
rect 3094 7760 3099 7764
rect 3103 7760 3143 7764
rect 3147 7760 3174 7764
rect 3178 7760 3196 7764
rect 3200 7760 3261 7764
rect 3265 7760 3279 7764
rect 3309 7759 3318 7763
rect 3322 7759 3369 7763
rect 3373 7759 3419 7763
rect 3423 7759 3450 7763
rect 3454 7759 3501 7763
rect 3505 7759 3551 7763
rect 3555 7759 3582 7763
rect 3586 7759 3633 7763
rect 3637 7759 3683 7763
rect 3687 7760 3757 7763
rect 3813 7760 3827 7764
rect 3831 7760 3858 7764
rect 3862 7760 3880 7764
rect 3884 7760 3945 7764
rect 3949 7760 3963 7764
rect 3999 7757 4002 7769
rect 4131 7767 4134 7771
rect 4158 7767 4159 7771
rect 4203 7767 4205 7771
rect 4826 7772 5086 7775
rect 4039 7760 4044 7764
rect 4048 7760 4088 7764
rect 4092 7760 4119 7764
rect 4123 7760 4141 7764
rect 4145 7760 4206 7764
rect 4210 7760 4224 7764
rect 2371 7753 2755 7756
rect 2770 7753 2855 7757
rect 2859 7753 2871 7757
rect 2875 7753 2889 7757
rect 2893 7753 2900 7757
rect 2904 7753 2906 7757
rect 2910 7753 2925 7757
rect 2929 7753 2962 7757
rect 2966 7753 2967 7757
rect 2971 7753 2979 7757
rect 2983 7753 3007 7757
rect 3011 7753 3047 7757
rect 3051 7753 3090 7757
rect 3094 7753 3101 7757
rect 3105 7753 3116 7757
rect 3120 7753 3132 7757
rect 3136 7753 3150 7757
rect 3154 7753 3161 7757
rect 3165 7753 3167 7757
rect 3171 7753 3186 7757
rect 3190 7753 3223 7757
rect 3227 7753 3228 7757
rect 3232 7753 3240 7757
rect 3244 7753 3268 7757
rect 3272 7753 3280 7757
rect 3316 7753 3700 7756
rect 3715 7753 3800 7757
rect 3804 7753 3816 7757
rect 3820 7753 3834 7757
rect 3838 7753 3845 7757
rect 3849 7753 3851 7757
rect 3855 7753 3870 7757
rect 3874 7753 3907 7757
rect 3911 7753 3912 7757
rect 3916 7753 3924 7757
rect 3928 7753 3952 7757
rect 3956 7753 3992 7757
rect 3996 7753 4035 7757
rect 4039 7753 4046 7757
rect 4050 7753 4061 7757
rect 4065 7753 4077 7757
rect 4081 7753 4095 7757
rect 4099 7753 4106 7757
rect 4110 7753 4112 7757
rect 4116 7753 4131 7757
rect 4135 7753 4168 7757
rect 4172 7753 4173 7757
rect 4177 7753 4185 7757
rect 4189 7753 4213 7757
rect 4217 7753 4225 7757
rect 2514 7746 2623 7749
rect 2806 7746 2864 7750
rect 2868 7746 3098 7749
rect 3288 7747 3296 7751
rect 3459 7746 3568 7749
rect 3751 7746 3809 7750
rect 3813 7746 4043 7749
rect 4233 7747 4241 7751
rect 2494 7738 2498 7742
rect 2502 7738 2506 7742
rect 2794 7739 3108 7742
rect 2842 7732 3115 7736
rect 3284 7729 3288 7735
rect 3439 7738 3443 7742
rect 3447 7738 3451 7742
rect 3739 7739 4053 7742
rect 3787 7732 4058 7736
rect 4229 7729 4233 7735
rect 4826 7733 4829 7772
rect 2350 7725 2482 7729
rect 2486 7725 2502 7729
rect 2518 7725 3427 7729
rect 3431 7725 3447 7729
rect 3463 7725 4321 7729
rect 4816 7723 4829 7733
rect 343 7710 356 7720
rect 2510 7718 2755 7721
rect 2830 7718 3156 7722
rect 3160 7718 3192 7722
rect 3196 7718 3259 7722
rect 3263 7718 3279 7722
rect 3455 7718 3700 7721
rect 3775 7718 4101 7722
rect 4105 7718 4137 7722
rect 4141 7718 4204 7722
rect 4208 7718 4224 7722
rect 2525 7711 2755 7714
rect 2770 7711 3142 7715
rect 3146 7711 3180 7715
rect 3184 7711 3208 7715
rect 3212 7711 3238 7715
rect 3242 7711 3275 7715
rect 343 7700 366 7710
rect 2494 7702 2498 7706
rect 2502 7702 2506 7706
rect 3150 7701 3153 7711
rect 3171 7701 3174 7711
rect 3187 7701 3190 7711
rect 3201 7704 3206 7708
rect 3210 7704 3217 7708
rect 3229 7701 3232 7711
rect 3245 7701 3248 7711
rect 3266 7701 3269 7711
rect 3470 7711 3700 7714
rect 3715 7711 4087 7715
rect 4091 7711 4125 7715
rect 4129 7711 4153 7715
rect 4157 7711 4183 7715
rect 4187 7711 4220 7715
rect 4806 7713 4829 7723
rect 3439 7702 3443 7706
rect 3447 7702 3451 7706
rect 4095 7701 4098 7711
rect 4116 7701 4119 7711
rect 4132 7701 4135 7711
rect 4146 7704 4151 7708
rect 4155 7704 4162 7708
rect 4174 7701 4177 7711
rect 4190 7701 4193 7711
rect 4211 7701 4214 7711
rect 4796 7703 4829 7713
rect 343 7690 376 7700
rect 2514 7695 2624 7698
rect 343 7680 386 7690
rect 2364 7688 2373 7692
rect 2377 7688 2409 7692
rect 2413 7688 2476 7692
rect 2480 7688 2505 7692
rect 2509 7688 2541 7692
rect 2545 7688 2608 7692
rect 2612 7688 2637 7692
rect 2641 7688 2673 7692
rect 2677 7688 2740 7692
rect 2744 7688 2824 7692
rect 2364 7681 2397 7685
rect 2401 7681 2425 7685
rect 2429 7681 2455 7685
rect 2459 7681 2492 7685
rect 2496 7681 2529 7685
rect 2533 7681 2557 7685
rect 2561 7681 2587 7685
rect 2591 7681 2624 7685
rect 2628 7681 2661 7685
rect 2665 7681 2689 7685
rect 2693 7681 2719 7685
rect 2723 7681 2756 7685
rect 2760 7681 2764 7685
rect 3167 7687 3172 7690
rect 3176 7687 3200 7690
rect 3459 7695 3569 7698
rect 3225 7687 3232 7690
rect 3236 7687 3258 7690
rect 3309 7688 3318 7692
rect 3322 7688 3354 7692
rect 3358 7688 3421 7692
rect 3425 7688 3450 7692
rect 3454 7688 3486 7692
rect 3490 7688 3553 7692
rect 3557 7688 3582 7692
rect 3586 7688 3618 7692
rect 3622 7688 3685 7692
rect 3689 7688 3769 7692
rect 343 7584 769 7680
rect 2367 7671 2370 7681
rect 2388 7671 2391 7681
rect 2404 7671 2407 7681
rect 2418 7674 2423 7678
rect 2427 7674 2434 7678
rect 2446 7671 2449 7681
rect 2462 7671 2465 7681
rect 2483 7671 2486 7681
rect 2499 7671 2502 7681
rect 2520 7671 2523 7681
rect 2536 7671 2539 7681
rect 2550 7674 2555 7678
rect 2559 7674 2566 7678
rect 2578 7671 2581 7681
rect 2594 7671 2597 7681
rect 2615 7671 2618 7681
rect 2631 7671 2634 7681
rect 2652 7671 2655 7681
rect 2668 7671 2671 7681
rect 2682 7674 2687 7678
rect 2691 7674 2698 7678
rect 2710 7671 2713 7681
rect 2726 7671 2729 7681
rect 2747 7671 2750 7681
rect 3183 7677 3190 7680
rect 3194 7681 3213 7684
rect 2384 7657 2389 7660
rect 2393 7657 2417 7660
rect 2442 7657 2449 7660
rect 2453 7657 2475 7660
rect 2495 7657 2502 7660
rect 2516 7657 2521 7660
rect 2525 7657 2549 7660
rect 2574 7657 2581 7660
rect 2585 7657 2607 7660
rect 2627 7657 2634 7660
rect 2648 7657 2653 7660
rect 2657 7657 2681 7660
rect 2706 7657 2713 7660
rect 2717 7657 2739 7660
rect 3213 7674 3216 7680
rect 3241 7677 3248 7680
rect 3252 7681 3267 7684
rect 3309 7681 3342 7685
rect 3346 7681 3370 7685
rect 3374 7681 3400 7685
rect 3404 7681 3437 7685
rect 3441 7681 3474 7685
rect 3478 7681 3502 7685
rect 3506 7681 3532 7685
rect 3536 7681 3569 7685
rect 3573 7681 3606 7685
rect 3610 7681 3634 7685
rect 3638 7681 3664 7685
rect 3668 7681 3701 7685
rect 3705 7681 3709 7685
rect 4112 7687 4117 7690
rect 4121 7687 4145 7690
rect 4786 7693 4829 7703
rect 4170 7687 4177 7690
rect 4181 7687 4203 7690
rect 3312 7671 3315 7681
rect 3333 7671 3336 7681
rect 3349 7671 3352 7681
rect 3363 7674 3368 7678
rect 3372 7674 3379 7678
rect 3391 7671 3394 7681
rect 3407 7671 3410 7681
rect 3428 7671 3431 7681
rect 3444 7671 3447 7681
rect 3465 7671 3468 7681
rect 3481 7671 3484 7681
rect 3495 7674 3500 7678
rect 3504 7674 3511 7678
rect 3523 7671 3526 7681
rect 3539 7671 3542 7681
rect 3560 7671 3563 7681
rect 3576 7671 3579 7681
rect 3597 7671 3600 7681
rect 3613 7671 3616 7681
rect 3627 7674 3632 7678
rect 3636 7674 3643 7678
rect 3655 7671 3658 7681
rect 3671 7671 3674 7681
rect 3692 7671 3695 7681
rect 4128 7677 4135 7680
rect 4139 7681 4158 7684
rect 3150 7658 3153 7670
rect 3171 7658 3174 7670
rect 3187 7658 3190 7670
rect 3201 7661 3213 7664
rect 3229 7658 3232 7670
rect 3245 7658 3248 7670
rect 3266 7658 3269 7670
rect 2400 7647 2407 7650
rect 2411 7651 2430 7654
rect 2430 7644 2433 7650
rect 2458 7647 2465 7650
rect 2469 7651 2484 7654
rect 2532 7647 2539 7650
rect 2543 7651 2562 7654
rect 2562 7644 2565 7650
rect 2590 7647 2597 7650
rect 2601 7651 2616 7654
rect 2664 7647 2671 7650
rect 2675 7651 2694 7654
rect 2694 7644 2697 7650
rect 2722 7647 2729 7650
rect 2733 7651 2750 7654
rect 2782 7654 3180 7658
rect 3184 7654 3208 7658
rect 3212 7654 3238 7658
rect 3242 7654 3279 7658
rect 3329 7657 3334 7660
rect 3338 7657 3362 7660
rect 3387 7657 3394 7660
rect 3398 7657 3420 7660
rect 3440 7657 3447 7660
rect 3461 7657 3466 7660
rect 3470 7657 3494 7660
rect 3519 7657 3526 7660
rect 3530 7657 3552 7660
rect 3572 7657 3579 7660
rect 3593 7657 3598 7660
rect 3602 7657 3626 7660
rect 3651 7657 3658 7660
rect 3662 7657 3684 7660
rect 4158 7674 4161 7680
rect 4186 7677 4193 7680
rect 4197 7681 4212 7684
rect 4095 7658 4098 7670
rect 4116 7658 4119 7670
rect 4132 7658 4135 7670
rect 4146 7661 4158 7664
rect 4174 7658 4177 7670
rect 4190 7658 4193 7670
rect 4211 7658 4214 7670
rect 2818 7647 3156 7651
rect 3160 7647 3207 7651
rect 3211 7647 3257 7651
rect 3261 7647 3279 7651
rect 3345 7647 3352 7650
rect 3356 7651 3375 7654
rect 2367 7628 2370 7640
rect 2388 7628 2391 7640
rect 2404 7628 2407 7640
rect 2418 7631 2430 7634
rect 2446 7628 2449 7640
rect 2462 7628 2465 7640
rect 2483 7628 2486 7640
rect 2499 7628 2502 7640
rect 2520 7628 2523 7640
rect 2536 7628 2539 7640
rect 2550 7631 2562 7634
rect 2578 7628 2581 7640
rect 2594 7628 2597 7640
rect 2615 7628 2618 7640
rect 2631 7628 2634 7640
rect 2652 7628 2655 7640
rect 2668 7628 2671 7640
rect 2682 7631 2694 7634
rect 2710 7628 2713 7640
rect 2726 7628 2729 7640
rect 2747 7628 2750 7640
rect 3153 7640 3274 7643
rect 3375 7644 3378 7650
rect 3403 7647 3410 7650
rect 3414 7651 3429 7654
rect 3477 7647 3484 7650
rect 3488 7651 3507 7654
rect 3507 7644 3510 7650
rect 3535 7647 3542 7650
rect 3546 7651 3561 7654
rect 3609 7647 3616 7650
rect 3620 7651 3639 7654
rect 3639 7644 3642 7650
rect 3667 7647 3674 7650
rect 3678 7651 3695 7654
rect 3727 7654 4125 7658
rect 4129 7654 4153 7658
rect 4157 7654 4183 7658
rect 4187 7654 4224 7658
rect 3763 7647 4101 7651
rect 4105 7647 4152 7651
rect 4156 7647 4202 7651
rect 4206 7647 4224 7651
rect 4403 7648 4829 7693
rect 2830 7632 3156 7636
rect 3160 7632 3192 7636
rect 3196 7632 3259 7636
rect 3263 7632 3279 7636
rect 2364 7624 2397 7628
rect 2401 7624 2425 7628
rect 2429 7624 2455 7628
rect 2459 7624 2529 7628
rect 2533 7624 2557 7628
rect 2561 7624 2587 7628
rect 2591 7624 2661 7628
rect 2665 7624 2689 7628
rect 2693 7624 2719 7628
rect 2723 7624 2776 7628
rect 3146 7625 3180 7629
rect 3184 7625 3208 7629
rect 3212 7625 3238 7629
rect 3242 7625 3275 7629
rect 3312 7628 3315 7640
rect 3333 7628 3336 7640
rect 3349 7628 3352 7640
rect 3363 7631 3375 7634
rect 3391 7628 3394 7640
rect 3407 7628 3410 7640
rect 3428 7628 3431 7640
rect 3444 7628 3447 7640
rect 3465 7628 3468 7640
rect 3481 7628 3484 7640
rect 3495 7631 3507 7634
rect 3523 7628 3526 7640
rect 3539 7628 3542 7640
rect 3560 7628 3563 7640
rect 3576 7628 3579 7640
rect 3597 7628 3600 7640
rect 3613 7628 3616 7640
rect 3627 7631 3639 7634
rect 3655 7628 3658 7640
rect 3671 7628 3674 7640
rect 3692 7628 3695 7640
rect 4098 7640 4219 7643
rect 3775 7632 4101 7636
rect 4105 7632 4137 7636
rect 4141 7632 4204 7636
rect 4208 7632 4224 7636
rect 4384 7635 4829 7648
rect 2364 7617 2373 7621
rect 2377 7617 2424 7621
rect 2428 7617 2474 7621
rect 2478 7617 2505 7621
rect 2509 7617 2556 7621
rect 2560 7617 2606 7621
rect 2610 7617 2637 7621
rect 2641 7617 2688 7621
rect 2692 7617 2738 7621
rect 2742 7617 2812 7621
rect 3150 7615 3153 7625
rect 3171 7615 3174 7625
rect 3187 7615 3190 7625
rect 3201 7618 3206 7622
rect 3210 7618 3217 7622
rect 3229 7615 3232 7625
rect 3245 7615 3248 7625
rect 3266 7615 3269 7625
rect 3309 7624 3342 7628
rect 3346 7624 3370 7628
rect 3374 7624 3400 7628
rect 3404 7624 3474 7628
rect 3478 7624 3502 7628
rect 3506 7624 3532 7628
rect 3536 7624 3606 7628
rect 3610 7624 3634 7628
rect 3638 7624 3664 7628
rect 3668 7624 3721 7628
rect 4091 7625 4125 7629
rect 4129 7625 4153 7629
rect 4157 7625 4183 7629
rect 4187 7625 4220 7629
rect 3309 7617 3318 7621
rect 3322 7617 3369 7621
rect 3373 7617 3419 7621
rect 3423 7617 3450 7621
rect 3454 7617 3501 7621
rect 3505 7617 3551 7621
rect 3555 7617 3582 7621
rect 3586 7617 3633 7621
rect 3637 7617 3683 7621
rect 3687 7617 3757 7621
rect 4095 7615 4098 7625
rect 4116 7615 4119 7625
rect 4132 7615 4135 7625
rect 4146 7618 4151 7622
rect 4155 7618 4162 7622
rect 4174 7615 4177 7625
rect 4190 7615 4193 7625
rect 4211 7615 4214 7625
rect 2370 7610 2755 7613
rect 2364 7602 2373 7606
rect 2377 7602 2409 7606
rect 2413 7602 2476 7606
rect 2480 7602 2505 7606
rect 2509 7602 2541 7606
rect 2545 7602 2608 7606
rect 2612 7602 2637 7606
rect 2641 7602 2673 7606
rect 2677 7602 2740 7606
rect 2744 7602 2824 7606
rect 2364 7595 2397 7599
rect 2401 7595 2425 7599
rect 2429 7595 2455 7599
rect 2459 7595 2492 7599
rect 2496 7595 2529 7599
rect 2533 7595 2557 7599
rect 2561 7595 2587 7599
rect 2591 7595 2624 7599
rect 2628 7595 2661 7599
rect 2665 7595 2689 7599
rect 2693 7595 2719 7599
rect 2723 7595 2756 7599
rect 2760 7595 2764 7599
rect 3167 7601 3172 7604
rect 3176 7601 3200 7604
rect 3315 7610 3700 7613
rect 3225 7601 3232 7604
rect 3236 7601 3258 7604
rect 3309 7602 3318 7606
rect 3322 7602 3354 7606
rect 3358 7602 3421 7606
rect 3425 7602 3450 7606
rect 3454 7602 3486 7606
rect 3490 7602 3553 7606
rect 3557 7602 3582 7606
rect 3586 7602 3618 7606
rect 3622 7602 3685 7606
rect 3689 7602 3769 7606
rect 2367 7585 2370 7595
rect 2388 7585 2391 7595
rect 2404 7585 2407 7595
rect 2418 7588 2423 7592
rect 2427 7588 2434 7592
rect 2446 7585 2449 7595
rect 2462 7585 2465 7595
rect 2483 7585 2486 7595
rect 2499 7585 2502 7595
rect 2520 7585 2523 7595
rect 2536 7585 2539 7595
rect 2550 7588 2555 7592
rect 2559 7588 2566 7592
rect 2578 7585 2581 7595
rect 2594 7585 2597 7595
rect 2615 7585 2618 7595
rect 2631 7585 2634 7595
rect 2652 7585 2655 7595
rect 2668 7585 2671 7595
rect 2682 7588 2687 7592
rect 2691 7588 2698 7592
rect 2710 7585 2713 7595
rect 2726 7585 2729 7595
rect 2747 7585 2750 7595
rect 3183 7591 3190 7594
rect 3194 7595 3213 7598
rect 343 7574 386 7584
rect 343 7564 376 7574
rect 2384 7571 2389 7574
rect 2393 7571 2417 7574
rect 2442 7571 2449 7574
rect 2453 7571 2475 7574
rect 2495 7571 2502 7574
rect 2516 7571 2521 7574
rect 2525 7571 2549 7574
rect 2574 7571 2581 7574
rect 2585 7571 2607 7574
rect 2627 7571 2634 7574
rect 2648 7571 2653 7574
rect 2657 7571 2681 7574
rect 2706 7571 2713 7574
rect 2717 7571 2739 7574
rect 3213 7588 3216 7594
rect 3241 7591 3248 7594
rect 3252 7595 3267 7598
rect 3278 7593 3289 7597
rect 3309 7595 3342 7599
rect 3346 7595 3370 7599
rect 3374 7595 3400 7599
rect 3404 7595 3437 7599
rect 3441 7595 3474 7599
rect 3478 7595 3502 7599
rect 3506 7595 3532 7599
rect 3536 7595 3569 7599
rect 3573 7595 3606 7599
rect 3610 7595 3634 7599
rect 3638 7595 3664 7599
rect 3668 7595 3701 7599
rect 3705 7595 3709 7599
rect 4112 7601 4117 7604
rect 4121 7601 4145 7604
rect 4170 7601 4177 7604
rect 4181 7601 4203 7604
rect 3312 7585 3315 7595
rect 3333 7585 3336 7595
rect 3349 7585 3352 7595
rect 3363 7588 3368 7592
rect 3372 7588 3379 7592
rect 3391 7585 3394 7595
rect 3407 7585 3410 7595
rect 3428 7585 3431 7595
rect 3444 7585 3447 7595
rect 3465 7585 3468 7595
rect 3481 7585 3484 7595
rect 3495 7588 3500 7592
rect 3504 7588 3511 7592
rect 3523 7585 3526 7595
rect 3539 7585 3542 7595
rect 3560 7585 3563 7595
rect 3576 7585 3579 7595
rect 3597 7585 3600 7595
rect 3613 7585 3616 7595
rect 3627 7588 3632 7592
rect 3636 7588 3643 7592
rect 3655 7585 3658 7595
rect 3671 7585 3674 7595
rect 3692 7585 3695 7595
rect 4128 7591 4135 7594
rect 4139 7595 4158 7598
rect 3150 7572 3153 7584
rect 3171 7572 3174 7584
rect 3187 7572 3190 7584
rect 3201 7575 3213 7578
rect 3229 7572 3232 7584
rect 3245 7572 3248 7584
rect 3266 7572 3269 7584
rect 343 7554 366 7564
rect 2400 7561 2407 7564
rect 2411 7565 2430 7568
rect 2430 7558 2433 7564
rect 2458 7561 2465 7564
rect 2469 7565 2484 7568
rect 2532 7561 2539 7564
rect 2543 7565 2562 7568
rect 2562 7558 2565 7564
rect 2590 7561 2597 7564
rect 2601 7565 2616 7568
rect 2664 7561 2671 7564
rect 2675 7565 2694 7568
rect 2694 7558 2697 7564
rect 2722 7561 2729 7564
rect 2733 7565 2750 7568
rect 2782 7568 3180 7572
rect 3184 7568 3208 7572
rect 3212 7568 3238 7572
rect 3242 7568 3279 7572
rect 3329 7571 3334 7574
rect 3338 7571 3362 7574
rect 3387 7571 3394 7574
rect 3398 7571 3420 7574
rect 3440 7571 3447 7574
rect 3461 7571 3466 7574
rect 3470 7571 3494 7574
rect 3519 7571 3526 7574
rect 3530 7571 3552 7574
rect 3572 7571 3579 7574
rect 3593 7571 3598 7574
rect 3602 7571 3626 7574
rect 3651 7571 3658 7574
rect 3662 7571 3684 7574
rect 4158 7588 4161 7594
rect 4186 7591 4193 7594
rect 4197 7595 4212 7598
rect 4403 7597 4829 7635
rect 4223 7593 4234 7597
rect 4786 7587 4829 7597
rect 4095 7572 4098 7584
rect 4116 7572 4119 7584
rect 4132 7572 4135 7584
rect 4146 7575 4158 7578
rect 4174 7572 4177 7584
rect 4190 7572 4193 7584
rect 4211 7572 4214 7584
rect 4796 7577 4829 7587
rect 2818 7561 3156 7565
rect 3160 7561 3207 7565
rect 3211 7561 3257 7565
rect 3261 7561 3279 7565
rect 3345 7561 3352 7564
rect 3356 7565 3375 7568
rect 3375 7558 3378 7564
rect 3403 7561 3410 7564
rect 3414 7565 3429 7568
rect 3477 7561 3484 7564
rect 3488 7565 3507 7568
rect 3507 7558 3510 7564
rect 3535 7561 3542 7564
rect 3546 7565 3561 7568
rect 3609 7561 3616 7564
rect 3620 7565 3639 7568
rect 3639 7558 3642 7564
rect 3667 7561 3674 7564
rect 3678 7565 3695 7568
rect 3727 7568 4125 7572
rect 4129 7568 4153 7572
rect 4157 7568 4183 7572
rect 4187 7568 4224 7572
rect 4806 7567 4829 7577
rect 3763 7561 4101 7565
rect 4105 7561 4152 7565
rect 4156 7561 4202 7565
rect 4206 7561 4224 7565
rect 4816 7557 4829 7567
rect 343 7544 356 7554
rect 343 7505 346 7544
rect 2367 7542 2370 7554
rect 2388 7542 2391 7554
rect 2404 7542 2407 7554
rect 2418 7545 2430 7548
rect 2446 7542 2449 7554
rect 2462 7542 2465 7554
rect 2483 7542 2486 7554
rect 2499 7542 2502 7554
rect 2520 7542 2523 7554
rect 2536 7542 2539 7554
rect 2550 7545 2562 7548
rect 2578 7542 2581 7554
rect 2594 7542 2597 7554
rect 2615 7542 2618 7554
rect 2631 7542 2634 7554
rect 2652 7542 2655 7554
rect 2668 7542 2671 7554
rect 2682 7545 2694 7548
rect 2710 7542 2713 7554
rect 2726 7542 2729 7554
rect 2747 7542 2750 7554
rect 3312 7542 3315 7554
rect 3333 7542 3336 7554
rect 3349 7542 3352 7554
rect 3363 7545 3375 7548
rect 3391 7542 3394 7554
rect 3407 7542 3410 7554
rect 3428 7542 3431 7554
rect 3444 7542 3447 7554
rect 3465 7542 3468 7554
rect 3481 7542 3484 7554
rect 3495 7545 3507 7548
rect 3523 7542 3526 7554
rect 3539 7542 3542 7554
rect 3560 7542 3563 7554
rect 3576 7542 3579 7554
rect 3597 7542 3600 7554
rect 3613 7542 3616 7554
rect 3627 7545 3639 7548
rect 3655 7542 3658 7554
rect 3671 7542 3674 7554
rect 3692 7542 3695 7554
rect 2364 7538 2397 7542
rect 2401 7538 2425 7542
rect 2429 7538 2455 7542
rect 2459 7538 2529 7542
rect 2533 7538 2557 7542
rect 2561 7538 2587 7542
rect 2591 7538 2661 7542
rect 2665 7538 2689 7542
rect 2693 7538 2719 7542
rect 2723 7538 2776 7542
rect 3309 7538 3342 7542
rect 3346 7538 3370 7542
rect 3374 7538 3400 7542
rect 3404 7538 3474 7542
rect 3478 7538 3502 7542
rect 3506 7538 3532 7542
rect 3536 7538 3606 7542
rect 3610 7538 3634 7542
rect 3638 7538 3664 7542
rect 3668 7538 3721 7542
rect 2364 7531 2373 7535
rect 2377 7531 2424 7535
rect 2428 7531 2474 7535
rect 2478 7531 2505 7535
rect 2509 7531 2556 7535
rect 2560 7531 2606 7535
rect 2610 7531 2637 7535
rect 2641 7531 2688 7535
rect 2692 7531 2738 7535
rect 2742 7531 2812 7535
rect 3309 7531 3318 7535
rect 3322 7531 3369 7535
rect 3373 7531 3419 7535
rect 3423 7531 3450 7535
rect 3454 7531 3501 7535
rect 3505 7531 3551 7535
rect 3555 7531 3582 7535
rect 3586 7531 3633 7535
rect 3637 7531 3683 7535
rect 3687 7531 3757 7535
rect 2370 7525 2755 7528
rect 3315 7525 3700 7528
rect 2495 7518 2599 7521
rect 3440 7518 3544 7521
rect 4826 7518 4829 7557
rect 5083 7518 5086 7772
rect 4826 7515 5086 7518
rect 2611 7510 2615 7514
rect 2619 7510 2623 7514
rect 3556 7510 3560 7514
rect 3564 7510 3568 7514
rect 86 7502 346 7505
rect 2347 7499 2599 7503
rect 2603 7499 2619 7503
rect 2635 7499 3296 7503
rect 3300 7499 3544 7503
rect 3548 7499 3564 7503
rect 3580 7499 3836 7503
rect 3844 7499 4241 7503
rect 4245 7499 4360 7503
rect 4527 7498 4595 7499
rect 2627 7492 2755 7495
rect 3572 7492 3700 7495
rect 4527 7494 4529 7498
rect 4533 7494 4534 7498
rect 4538 7494 4539 7498
rect 4543 7494 4544 7498
rect 4548 7494 4549 7498
rect 4553 7494 4554 7498
rect 4558 7494 4559 7498
rect 4563 7494 4564 7498
rect 4568 7494 4569 7498
rect 4573 7494 4574 7498
rect 4578 7494 4579 7498
rect 4583 7494 4584 7498
rect 4588 7494 4589 7498
rect 4593 7494 4595 7498
rect 4527 7493 4595 7494
rect 4527 7489 4529 7493
rect 4533 7489 4534 7493
rect 4538 7489 4539 7493
rect 4543 7489 4544 7493
rect 4548 7489 4549 7493
rect 4553 7489 4554 7493
rect 4558 7489 4559 7493
rect 4563 7489 4564 7493
rect 4568 7489 4569 7493
rect 4573 7489 4574 7493
rect 4578 7489 4579 7493
rect 4583 7489 4584 7493
rect 4588 7489 4589 7493
rect 4593 7489 4595 7493
rect 4826 7490 5086 7493
rect 2642 7485 2755 7488
rect 3587 7485 3700 7488
rect 4527 7487 4595 7489
rect 4527 7486 4632 7487
rect 4636 7486 4637 7490
rect 4641 7486 4642 7490
rect 4646 7486 4647 7490
rect 4651 7486 4652 7490
rect 4656 7486 4657 7490
rect 4661 7486 4662 7490
rect 4666 7486 4667 7490
rect 4671 7486 4672 7490
rect 4676 7486 4677 7490
rect 4681 7486 4682 7490
rect 4686 7486 4687 7490
rect 4691 7486 4692 7490
rect 4696 7486 4697 7490
rect 4701 7486 4702 7490
rect 4706 7486 4707 7490
rect 4711 7486 4712 7490
rect 4716 7486 4717 7490
rect 4721 7486 4722 7490
rect 4726 7486 4727 7490
rect 4731 7486 4732 7490
rect 4736 7486 4737 7490
rect 4741 7486 4742 7490
rect 4746 7486 4747 7490
rect 4751 7486 4752 7490
rect 4756 7486 4757 7490
rect 4761 7486 4762 7490
rect 4766 7486 4767 7490
rect 4527 7485 4636 7486
rect 2611 7476 2615 7480
rect 2619 7476 2623 7480
rect 3556 7476 3560 7480
rect 3564 7476 3568 7480
rect 4527 7481 4632 7485
rect 4527 7480 4636 7481
rect 4527 7476 4632 7480
rect 4767 7485 4771 7486
rect 4767 7480 4771 7481
rect 617 7467 618 7471
rect 622 7467 623 7471
rect 627 7467 628 7471
rect 632 7467 633 7471
rect 637 7467 638 7471
rect 642 7467 643 7471
rect 613 7466 647 7467
rect 617 7462 618 7466
rect 622 7462 623 7466
rect 627 7462 628 7466
rect 632 7462 633 7466
rect 637 7462 638 7466
rect 642 7462 643 7466
rect 613 7461 647 7462
rect 617 7457 618 7461
rect 622 7457 623 7461
rect 627 7457 628 7461
rect 632 7457 633 7461
rect 637 7457 638 7461
rect 642 7457 643 7461
rect 613 7456 647 7457
rect 86 7450 346 7453
rect 617 7452 618 7456
rect 622 7452 623 7456
rect 627 7452 628 7456
rect 632 7452 633 7456
rect 637 7452 638 7456
rect 642 7452 643 7456
rect 663 7467 664 7471
rect 668 7467 669 7471
rect 673 7467 674 7471
rect 678 7467 679 7471
rect 683 7467 684 7471
rect 688 7467 689 7471
rect 2495 7469 2599 7472
rect 3440 7469 3544 7472
rect 3851 7472 3918 7476
rect 4527 7475 4636 7476
rect 659 7466 693 7467
rect 663 7462 664 7466
rect 668 7462 669 7466
rect 673 7462 674 7466
rect 678 7462 679 7466
rect 683 7462 684 7466
rect 688 7462 689 7466
rect 2364 7462 2373 7466
rect 2377 7462 2409 7466
rect 2413 7462 2476 7466
rect 2480 7462 2505 7466
rect 2509 7462 2541 7466
rect 2545 7462 2608 7466
rect 2612 7462 2637 7466
rect 2641 7462 2673 7466
rect 2677 7462 2740 7466
rect 2744 7462 2824 7466
rect 3309 7462 3318 7466
rect 3322 7462 3354 7466
rect 3358 7462 3421 7466
rect 3425 7462 3450 7466
rect 3454 7462 3486 7466
rect 3490 7462 3553 7466
rect 3557 7462 3582 7466
rect 3586 7462 3618 7466
rect 3622 7462 3685 7466
rect 3689 7462 3769 7466
rect 4527 7471 4632 7475
rect 4527 7470 4636 7471
rect 4527 7466 4632 7470
rect 4527 7465 4636 7466
rect 659 7461 693 7462
rect 663 7457 664 7461
rect 668 7457 669 7461
rect 673 7457 674 7461
rect 678 7457 679 7461
rect 683 7457 684 7461
rect 688 7457 689 7461
rect 4527 7461 4632 7465
rect 4527 7460 4636 7461
rect 659 7456 693 7457
rect 663 7452 664 7456
rect 668 7452 669 7456
rect 673 7452 674 7456
rect 678 7452 679 7456
rect 683 7452 684 7456
rect 688 7452 689 7456
rect 2364 7455 2397 7459
rect 2401 7455 2425 7459
rect 2429 7455 2455 7459
rect 2459 7455 2492 7459
rect 2496 7455 2529 7459
rect 2533 7455 2557 7459
rect 2561 7455 2587 7459
rect 2591 7455 2624 7459
rect 2628 7455 2661 7459
rect 2665 7455 2689 7459
rect 2693 7455 2719 7459
rect 2723 7455 2756 7459
rect 2760 7455 2764 7459
rect 3309 7455 3342 7459
rect 3346 7455 3370 7459
rect 3374 7455 3400 7459
rect 3404 7455 3437 7459
rect 3441 7455 3474 7459
rect 3478 7455 3502 7459
rect 3506 7455 3532 7459
rect 3536 7455 3569 7459
rect 3573 7455 3606 7459
rect 3610 7455 3634 7459
rect 3638 7455 3664 7459
rect 3668 7455 3701 7459
rect 3705 7455 3709 7459
rect 4527 7456 4632 7460
rect 4527 7455 4636 7456
rect 86 7196 89 7450
rect 343 7411 346 7450
rect 2367 7445 2370 7455
rect 2388 7445 2391 7455
rect 2404 7445 2407 7455
rect 2418 7448 2423 7452
rect 2427 7448 2434 7452
rect 2446 7445 2449 7455
rect 2462 7445 2465 7455
rect 2483 7445 2486 7455
rect 2499 7445 2502 7455
rect 2520 7445 2523 7455
rect 2536 7445 2539 7455
rect 2550 7448 2555 7452
rect 2559 7448 2566 7452
rect 2578 7445 2581 7455
rect 2594 7445 2597 7455
rect 2615 7445 2618 7455
rect 2631 7445 2634 7455
rect 2652 7445 2655 7455
rect 2668 7445 2671 7455
rect 2682 7448 2687 7452
rect 2691 7448 2698 7452
rect 2710 7445 2713 7455
rect 2726 7445 2729 7455
rect 2747 7445 2750 7455
rect 3312 7445 3315 7455
rect 3333 7445 3336 7455
rect 3349 7445 3352 7455
rect 3363 7448 3368 7452
rect 3372 7448 3379 7452
rect 3391 7445 3394 7455
rect 3407 7445 3410 7455
rect 3428 7445 3431 7455
rect 3444 7445 3447 7455
rect 3465 7445 3468 7455
rect 3481 7445 3484 7455
rect 3495 7448 3500 7452
rect 3504 7448 3511 7452
rect 3523 7445 3526 7455
rect 3539 7445 3542 7455
rect 3560 7445 3563 7455
rect 3576 7445 3579 7455
rect 3597 7445 3600 7455
rect 3613 7445 3616 7455
rect 3627 7448 3632 7452
rect 3636 7448 3643 7452
rect 3655 7445 3658 7455
rect 3671 7445 3674 7455
rect 3692 7445 3695 7455
rect 4527 7451 4632 7455
rect 4527 7450 4636 7451
rect 4527 7446 4632 7450
rect 4527 7445 4636 7446
rect 2384 7431 2389 7434
rect 2393 7431 2417 7434
rect 2442 7431 2449 7434
rect 2453 7431 2475 7434
rect 2495 7431 2502 7434
rect 2516 7431 2521 7434
rect 2525 7431 2549 7434
rect 2574 7431 2581 7434
rect 2585 7431 2607 7434
rect 2627 7431 2634 7434
rect 2648 7431 2653 7434
rect 2657 7431 2681 7434
rect 2706 7431 2713 7434
rect 2717 7431 2739 7434
rect 2400 7421 2407 7424
rect 2411 7425 2430 7428
rect 2430 7418 2433 7424
rect 2458 7421 2465 7424
rect 2469 7425 2484 7428
rect 2532 7421 2539 7424
rect 2543 7425 2562 7428
rect 2562 7418 2565 7424
rect 2590 7421 2597 7424
rect 2601 7425 2616 7428
rect 2664 7421 2671 7424
rect 2675 7425 2694 7428
rect 2694 7418 2697 7424
rect 2722 7421 2729 7424
rect 2733 7425 2750 7428
rect 3329 7431 3334 7434
rect 3338 7431 3362 7434
rect 3387 7431 3394 7434
rect 3398 7431 3420 7434
rect 3440 7431 3447 7434
rect 3461 7431 3466 7434
rect 3470 7431 3494 7434
rect 3519 7431 3526 7434
rect 3530 7431 3552 7434
rect 3572 7431 3579 7434
rect 3593 7431 3598 7434
rect 3602 7431 3626 7434
rect 3651 7431 3658 7434
rect 3662 7431 3684 7434
rect 4527 7441 4632 7445
rect 4527 7440 4636 7441
rect 4527 7436 4632 7440
rect 4527 7435 4636 7436
rect 4527 7431 4632 7435
rect 3345 7421 3352 7424
rect 3356 7425 3375 7428
rect 3375 7418 3378 7424
rect 3403 7421 3410 7424
rect 3414 7425 3429 7428
rect 3477 7421 3484 7424
rect 3488 7425 3507 7428
rect 3507 7418 3510 7424
rect 3535 7421 3542 7424
rect 3546 7425 3561 7428
rect 3609 7421 3616 7424
rect 3620 7425 3639 7428
rect 3639 7418 3642 7424
rect 3667 7421 3674 7424
rect 3678 7425 3695 7428
rect 4572 7428 4576 7431
rect 4588 7428 4592 7431
rect 4604 7428 4608 7431
rect 4620 7428 4624 7431
rect 343 7401 356 7411
rect 2367 7402 2370 7414
rect 2388 7402 2391 7414
rect 2404 7402 2407 7414
rect 2418 7405 2430 7408
rect 2446 7402 2449 7414
rect 2462 7402 2465 7414
rect 2483 7402 2486 7414
rect 2499 7402 2502 7414
rect 2520 7402 2523 7414
rect 2536 7402 2539 7414
rect 2550 7405 2562 7408
rect 2578 7402 2581 7414
rect 2594 7402 2597 7414
rect 2615 7402 2618 7414
rect 2631 7402 2634 7414
rect 2652 7402 2655 7414
rect 2668 7402 2671 7414
rect 2682 7405 2694 7408
rect 2710 7402 2713 7414
rect 2726 7402 2729 7414
rect 2747 7402 2750 7414
rect 3312 7402 3315 7414
rect 3333 7402 3336 7414
rect 3349 7402 3352 7414
rect 3363 7405 3375 7408
rect 3391 7402 3394 7414
rect 3407 7402 3410 7414
rect 3428 7402 3431 7414
rect 3444 7402 3447 7414
rect 3465 7402 3468 7414
rect 3481 7402 3484 7414
rect 3495 7405 3507 7408
rect 3523 7402 3526 7414
rect 3539 7402 3542 7414
rect 3560 7402 3563 7414
rect 3576 7402 3579 7414
rect 3597 7402 3600 7414
rect 3613 7402 3616 7414
rect 3627 7405 3639 7408
rect 3655 7402 3658 7414
rect 3671 7402 3674 7414
rect 3692 7402 3695 7414
rect 343 7391 366 7401
rect 2364 7398 2397 7402
rect 2401 7398 2425 7402
rect 2429 7398 2455 7402
rect 2459 7398 2529 7402
rect 2533 7398 2557 7402
rect 2561 7398 2587 7402
rect 2591 7398 2661 7402
rect 2665 7398 2689 7402
rect 2693 7398 2719 7402
rect 2723 7398 2776 7402
rect 3309 7398 3342 7402
rect 3346 7398 3370 7402
rect 3374 7398 3400 7402
rect 3404 7398 3474 7402
rect 3478 7398 3502 7402
rect 3506 7398 3532 7402
rect 3536 7398 3606 7402
rect 3610 7398 3634 7402
rect 3638 7398 3664 7402
rect 3668 7398 3721 7402
rect 2364 7391 2373 7395
rect 2377 7391 2424 7395
rect 2428 7391 2474 7395
rect 2478 7391 2505 7395
rect 2509 7391 2556 7395
rect 2560 7391 2606 7395
rect 2610 7391 2637 7395
rect 2641 7391 2688 7395
rect 2692 7391 2738 7395
rect 2742 7391 2812 7395
rect 3309 7391 3318 7395
rect 3322 7391 3369 7395
rect 3373 7391 3419 7395
rect 3423 7391 3450 7395
rect 3454 7391 3501 7395
rect 3505 7391 3551 7395
rect 3555 7391 3582 7395
rect 3586 7391 3633 7395
rect 3637 7391 3683 7395
rect 3687 7391 3757 7395
rect 343 7381 376 7391
rect 343 7371 386 7381
rect 4632 7430 4636 7431
rect 4632 7425 4636 7426
rect 4632 7420 4636 7421
rect 4632 7415 4636 7416
rect 4632 7410 4636 7411
rect 4649 7473 4652 7477
rect 4656 7473 4657 7477
rect 4661 7473 4662 7477
rect 4666 7473 4667 7477
rect 4671 7473 4672 7477
rect 4676 7473 4677 7477
rect 4681 7473 4682 7477
rect 4686 7473 4687 7477
rect 4691 7473 4692 7477
rect 4696 7473 4697 7477
rect 4701 7473 4702 7477
rect 4706 7473 4707 7477
rect 4711 7473 4712 7477
rect 4716 7473 4717 7477
rect 4721 7473 4722 7477
rect 4726 7473 4727 7477
rect 4731 7473 4732 7477
rect 4736 7473 4737 7477
rect 4741 7473 4742 7477
rect 4746 7473 4747 7477
rect 4751 7473 4754 7477
rect 4641 7470 4649 7473
rect 4641 7465 4649 7466
rect 4754 7470 4758 7473
rect 4754 7465 4758 7466
rect 4641 7460 4649 7461
rect 4641 7455 4649 7456
rect 4641 7450 4649 7451
rect 4641 7445 4649 7446
rect 4641 7440 4649 7441
rect 4641 7435 4649 7436
rect 4641 7430 4649 7431
rect 4641 7425 4649 7426
rect 4661 7461 4662 7465
rect 4666 7461 4667 7465
rect 4671 7461 4672 7465
rect 4676 7461 4677 7465
rect 4681 7461 4682 7465
rect 4686 7461 4687 7465
rect 4691 7461 4692 7465
rect 4696 7461 4697 7465
rect 4701 7461 4702 7465
rect 4706 7461 4707 7465
rect 4711 7461 4712 7465
rect 4716 7461 4717 7465
rect 4721 7461 4722 7465
rect 4726 7461 4727 7465
rect 4731 7461 4732 7465
rect 4736 7461 4737 7465
rect 4741 7461 4742 7465
rect 4657 7460 4746 7461
rect 4661 7456 4662 7460
rect 4666 7456 4667 7460
rect 4671 7456 4672 7460
rect 4676 7456 4677 7460
rect 4681 7456 4682 7460
rect 4686 7456 4687 7460
rect 4691 7456 4692 7460
rect 4696 7456 4697 7460
rect 4701 7456 4702 7460
rect 4706 7456 4707 7460
rect 4711 7456 4712 7460
rect 4716 7456 4717 7460
rect 4721 7456 4722 7460
rect 4726 7456 4727 7460
rect 4731 7456 4732 7460
rect 4736 7456 4737 7460
rect 4741 7456 4742 7460
rect 4657 7455 4746 7456
rect 4661 7451 4662 7455
rect 4666 7451 4667 7455
rect 4671 7451 4672 7455
rect 4676 7451 4677 7455
rect 4681 7451 4682 7455
rect 4686 7451 4687 7455
rect 4691 7451 4692 7455
rect 4696 7451 4697 7455
rect 4701 7451 4702 7455
rect 4706 7451 4707 7455
rect 4711 7451 4712 7455
rect 4716 7451 4717 7455
rect 4721 7451 4722 7455
rect 4726 7451 4727 7455
rect 4731 7451 4732 7455
rect 4736 7451 4737 7455
rect 4741 7451 4742 7455
rect 4657 7450 4746 7451
rect 4661 7446 4662 7450
rect 4666 7446 4667 7450
rect 4671 7446 4672 7450
rect 4676 7446 4677 7450
rect 4681 7446 4682 7450
rect 4686 7446 4687 7450
rect 4691 7446 4692 7450
rect 4696 7446 4697 7450
rect 4701 7446 4702 7450
rect 4706 7446 4707 7450
rect 4711 7446 4712 7450
rect 4716 7446 4717 7450
rect 4721 7446 4722 7450
rect 4726 7446 4727 7450
rect 4731 7446 4732 7450
rect 4736 7446 4737 7450
rect 4741 7446 4742 7450
rect 4657 7445 4746 7446
rect 4661 7441 4662 7445
rect 4666 7441 4667 7445
rect 4671 7441 4672 7445
rect 4676 7441 4677 7445
rect 4681 7441 4682 7445
rect 4686 7441 4687 7445
rect 4691 7441 4692 7445
rect 4696 7441 4697 7445
rect 4701 7441 4702 7445
rect 4706 7441 4707 7445
rect 4711 7441 4712 7445
rect 4716 7441 4717 7445
rect 4721 7441 4722 7445
rect 4726 7441 4727 7445
rect 4731 7441 4732 7445
rect 4736 7441 4737 7445
rect 4741 7441 4742 7445
rect 4657 7440 4746 7441
rect 4661 7436 4662 7440
rect 4666 7436 4667 7440
rect 4671 7436 4672 7440
rect 4676 7436 4677 7440
rect 4681 7436 4682 7440
rect 4686 7436 4687 7440
rect 4691 7436 4692 7440
rect 4696 7436 4697 7440
rect 4701 7436 4702 7440
rect 4706 7436 4707 7440
rect 4711 7436 4712 7440
rect 4716 7436 4717 7440
rect 4721 7436 4722 7440
rect 4726 7436 4727 7440
rect 4731 7436 4732 7440
rect 4736 7436 4737 7440
rect 4741 7436 4742 7440
rect 4657 7435 4746 7436
rect 4661 7431 4662 7435
rect 4666 7431 4667 7435
rect 4671 7431 4672 7435
rect 4676 7431 4677 7435
rect 4681 7431 4682 7435
rect 4686 7431 4687 7435
rect 4691 7431 4692 7435
rect 4696 7431 4697 7435
rect 4701 7431 4702 7435
rect 4706 7431 4707 7435
rect 4711 7431 4712 7435
rect 4716 7431 4717 7435
rect 4721 7431 4722 7435
rect 4726 7431 4727 7435
rect 4731 7431 4732 7435
rect 4736 7431 4737 7435
rect 4741 7431 4742 7435
rect 4657 7430 4746 7431
rect 4661 7426 4662 7430
rect 4666 7426 4667 7430
rect 4671 7426 4672 7430
rect 4676 7426 4677 7430
rect 4681 7426 4682 7430
rect 4686 7426 4687 7430
rect 4691 7426 4692 7430
rect 4696 7426 4697 7430
rect 4701 7426 4702 7430
rect 4706 7426 4707 7430
rect 4711 7426 4712 7430
rect 4716 7426 4717 7430
rect 4721 7426 4722 7430
rect 4726 7426 4727 7430
rect 4731 7426 4732 7430
rect 4736 7426 4737 7430
rect 4741 7426 4742 7430
rect 4657 7425 4746 7426
rect 4661 7421 4662 7425
rect 4666 7421 4667 7425
rect 4671 7421 4672 7425
rect 4676 7421 4677 7425
rect 4681 7421 4682 7425
rect 4686 7421 4687 7425
rect 4691 7421 4692 7425
rect 4696 7421 4697 7425
rect 4701 7421 4702 7425
rect 4706 7421 4707 7425
rect 4711 7421 4712 7425
rect 4716 7421 4717 7425
rect 4721 7421 4722 7425
rect 4726 7421 4727 7425
rect 4731 7421 4732 7425
rect 4736 7421 4737 7425
rect 4741 7421 4742 7425
rect 4754 7460 4758 7461
rect 4754 7455 4758 7456
rect 4754 7450 4758 7451
rect 4754 7445 4758 7446
rect 4754 7440 4758 7441
rect 4754 7435 4758 7436
rect 4754 7430 4758 7431
rect 4754 7425 4758 7426
rect 4641 7420 4649 7421
rect 4641 7413 4649 7416
rect 4754 7420 4758 7421
rect 4754 7413 4758 7416
rect 4649 7409 4652 7413
rect 4656 7409 4657 7413
rect 4661 7409 4662 7413
rect 4666 7409 4667 7413
rect 4671 7409 4672 7413
rect 4676 7409 4677 7413
rect 4681 7409 4682 7413
rect 4686 7409 4687 7413
rect 4691 7409 4692 7413
rect 4696 7409 4697 7413
rect 4701 7409 4702 7413
rect 4706 7409 4707 7413
rect 4711 7409 4712 7413
rect 4716 7409 4717 7413
rect 4721 7409 4722 7413
rect 4726 7409 4727 7413
rect 4731 7409 4732 7413
rect 4736 7409 4737 7413
rect 4741 7409 4742 7413
rect 4746 7409 4747 7413
rect 4751 7409 4754 7413
rect 4767 7475 4771 7476
rect 4767 7470 4771 7471
rect 4767 7465 4771 7466
rect 4767 7460 4771 7461
rect 4767 7455 4771 7456
rect 4826 7451 4829 7490
rect 4767 7450 4771 7451
rect 4767 7445 4771 7446
rect 4816 7441 4829 7451
rect 4767 7440 4771 7441
rect 4767 7435 4771 7436
rect 4806 7431 4829 7441
rect 4767 7430 4771 7431
rect 4767 7425 4771 7426
rect 4796 7421 4829 7431
rect 4767 7420 4771 7421
rect 4767 7415 4771 7416
rect 4786 7411 4829 7421
rect 4767 7410 4771 7411
rect 4632 7405 4636 7406
rect 4632 7400 4636 7401
rect 4767 7405 4771 7406
rect 4767 7400 4771 7401
rect 4636 7396 4637 7400
rect 4641 7396 4642 7400
rect 4646 7396 4647 7400
rect 4651 7396 4652 7400
rect 4656 7396 4657 7400
rect 4661 7396 4662 7400
rect 4666 7396 4667 7400
rect 4671 7396 4672 7400
rect 4676 7396 4677 7400
rect 4681 7396 4682 7400
rect 4686 7396 4687 7400
rect 4691 7396 4692 7400
rect 4696 7396 4697 7400
rect 4701 7396 4702 7400
rect 4706 7396 4707 7400
rect 4711 7396 4712 7400
rect 4716 7396 4717 7400
rect 4721 7396 4722 7400
rect 4726 7396 4727 7400
rect 4731 7396 4732 7400
rect 4736 7396 4737 7400
rect 4741 7396 4742 7400
rect 4746 7396 4747 7400
rect 4751 7396 4752 7400
rect 4756 7396 4757 7400
rect 4761 7396 4762 7400
rect 4766 7396 4767 7400
rect 4774 7408 4829 7411
rect 4774 7404 4775 7408
rect 4779 7404 4780 7408
rect 4784 7404 4785 7408
rect 4789 7404 4790 7408
rect 4794 7404 4829 7408
rect 4774 7401 4829 7404
rect 4774 7397 4775 7401
rect 4779 7397 4780 7401
rect 4784 7397 4785 7401
rect 4789 7397 4790 7401
rect 4794 7397 4829 7401
rect 4774 7394 4829 7397
rect 4774 7390 4775 7394
rect 4779 7390 4780 7394
rect 4784 7390 4785 7394
rect 4789 7390 4790 7394
rect 4794 7390 4829 7394
rect 4774 7387 4829 7390
rect 4774 7383 4775 7387
rect 4779 7383 4780 7387
rect 4784 7383 4785 7387
rect 4789 7383 4790 7387
rect 4794 7383 4829 7387
rect 4774 7380 4829 7383
rect 4774 7376 4775 7380
rect 4779 7376 4780 7380
rect 4784 7376 4785 7380
rect 4789 7376 4790 7380
rect 4794 7376 4829 7380
rect 4774 7374 4829 7376
rect 4639 7372 4667 7374
rect 343 7275 769 7371
rect 4580 7368 4584 7372
rect 4596 7368 4600 7372
rect 4580 7367 4600 7368
rect 4406 7366 4600 7367
rect 3922 7362 4600 7366
rect 3918 7361 4600 7362
rect 3918 7354 4593 7361
rect 4612 7358 4616 7372
rect 4637 7370 4667 7372
rect 4635 7368 4667 7370
rect 4624 7359 4667 7368
rect 3918 7349 4414 7354
rect 4203 7348 4414 7349
rect 4580 7349 4593 7354
rect 4605 7354 4616 7358
rect 4635 7357 4667 7359
rect 4637 7355 4667 7357
rect 4580 7345 4600 7349
rect 4580 7342 4584 7345
rect 4596 7342 4600 7345
rect 4612 7342 4616 7354
rect 4639 7353 4667 7355
rect 4754 7373 4829 7374
rect 4754 7369 4775 7373
rect 4779 7369 4780 7373
rect 4784 7369 4785 7373
rect 4789 7369 4790 7373
rect 4794 7369 4829 7373
rect 4754 7366 4829 7369
rect 4754 7362 4775 7366
rect 4779 7362 4780 7366
rect 4784 7362 4785 7366
rect 4789 7362 4790 7366
rect 4794 7362 4829 7366
rect 4754 7359 4829 7362
rect 4754 7355 4775 7359
rect 4779 7355 4780 7359
rect 4784 7355 4785 7359
rect 4789 7355 4790 7359
rect 4794 7355 4829 7359
rect 4754 7353 4829 7355
rect 4774 7352 4829 7353
rect 4774 7348 4775 7352
rect 4779 7348 4780 7352
rect 4784 7348 4785 7352
rect 4789 7348 4790 7352
rect 4794 7348 4829 7352
rect 4774 7345 4829 7348
rect 4774 7341 4775 7345
rect 4779 7341 4780 7345
rect 4784 7341 4785 7345
rect 4789 7341 4790 7345
rect 4794 7341 4829 7345
rect 4774 7338 4829 7341
rect 4774 7334 4775 7338
rect 4779 7334 4780 7338
rect 4784 7334 4785 7338
rect 4789 7334 4790 7338
rect 4794 7334 4829 7338
rect 4774 7331 4829 7334
rect 4572 7293 4576 7302
rect 4588 7293 4592 7302
rect 4604 7293 4608 7302
rect 4620 7293 4624 7302
rect 4636 7326 4637 7330
rect 4641 7326 4642 7330
rect 4646 7326 4647 7330
rect 4651 7326 4652 7330
rect 4656 7326 4657 7330
rect 4661 7326 4662 7330
rect 4666 7326 4667 7330
rect 4671 7326 4672 7330
rect 4676 7326 4677 7330
rect 4681 7326 4682 7330
rect 4686 7326 4687 7330
rect 4691 7326 4692 7330
rect 4696 7326 4697 7330
rect 4701 7326 4702 7330
rect 4706 7326 4707 7330
rect 4711 7326 4712 7330
rect 4716 7326 4717 7330
rect 4721 7326 4722 7330
rect 4726 7326 4727 7330
rect 4731 7326 4732 7330
rect 4736 7326 4737 7330
rect 4741 7326 4742 7330
rect 4746 7326 4747 7330
rect 4751 7326 4752 7330
rect 4756 7326 4757 7330
rect 4761 7326 4762 7330
rect 4766 7326 4767 7330
rect 4632 7325 4636 7326
rect 4632 7320 4636 7321
rect 4767 7325 4771 7326
rect 4767 7320 4771 7321
rect 4632 7315 4636 7316
rect 4632 7310 4636 7311
rect 4632 7305 4636 7306
rect 4632 7300 4636 7301
rect 4632 7295 4636 7296
rect 4505 7289 4506 7293
rect 4510 7289 4511 7293
rect 4515 7291 4632 7293
rect 4515 7290 4636 7291
rect 4515 7289 4632 7290
rect 4505 7288 4632 7289
rect 4505 7284 4506 7288
rect 4510 7284 4511 7288
rect 4515 7286 4632 7288
rect 4515 7285 4636 7286
rect 4515 7284 4632 7285
rect 4505 7283 4632 7284
rect 4505 7279 4506 7283
rect 4510 7279 4511 7283
rect 4515 7281 4632 7283
rect 4515 7280 4636 7281
rect 4515 7279 4632 7280
rect 4505 7278 4632 7279
rect 343 7265 386 7275
rect 4505 7274 4506 7278
rect 4510 7274 4511 7278
rect 4515 7276 4632 7278
rect 4515 7275 4636 7276
rect 4515 7274 4632 7275
rect 4505 7273 4632 7274
rect 4505 7269 4506 7273
rect 4510 7269 4511 7273
rect 4515 7271 4632 7273
rect 4515 7270 4636 7271
rect 4515 7269 4632 7270
rect 4505 7268 4632 7269
rect 343 7255 376 7265
rect 4505 7264 4506 7268
rect 4510 7264 4511 7268
rect 4515 7266 4632 7268
rect 4515 7265 4636 7266
rect 4515 7264 4632 7265
rect 4505 7263 4632 7264
rect 4505 7259 4506 7263
rect 4510 7259 4511 7263
rect 4515 7261 4632 7263
rect 4515 7260 4636 7261
rect 4515 7259 4632 7260
rect 4505 7258 4632 7259
rect 343 7245 366 7255
rect 4505 7254 4506 7258
rect 4510 7254 4511 7258
rect 4515 7256 4632 7258
rect 4515 7255 4636 7256
rect 4515 7254 4632 7255
rect 4505 7253 4632 7254
rect 4505 7249 4506 7253
rect 4510 7249 4511 7253
rect 4515 7251 4632 7253
rect 4515 7250 4636 7251
rect 4515 7249 4632 7250
rect 4505 7248 4632 7249
rect 343 7235 356 7245
rect 4505 7244 4506 7248
rect 4510 7244 4511 7248
rect 4515 7246 4632 7248
rect 4649 7313 4652 7317
rect 4656 7313 4657 7317
rect 4661 7313 4662 7317
rect 4666 7313 4667 7317
rect 4671 7313 4672 7317
rect 4676 7313 4677 7317
rect 4681 7313 4682 7317
rect 4686 7313 4687 7317
rect 4691 7313 4692 7317
rect 4696 7313 4697 7317
rect 4701 7313 4702 7317
rect 4706 7313 4707 7317
rect 4711 7313 4712 7317
rect 4716 7313 4717 7317
rect 4721 7313 4722 7317
rect 4726 7313 4727 7317
rect 4731 7313 4732 7317
rect 4736 7313 4737 7317
rect 4741 7313 4742 7317
rect 4746 7313 4747 7317
rect 4751 7313 4754 7317
rect 4641 7310 4649 7313
rect 4754 7310 4758 7313
rect 4641 7305 4649 7306
rect 4641 7300 4649 7301
rect 4641 7295 4649 7296
rect 4641 7290 4649 7291
rect 4641 7285 4649 7286
rect 4641 7280 4649 7281
rect 4641 7275 4649 7276
rect 4641 7270 4649 7271
rect 4641 7265 4649 7266
rect 4657 7305 4746 7306
rect 4661 7301 4662 7305
rect 4666 7301 4667 7305
rect 4671 7301 4672 7305
rect 4676 7301 4677 7305
rect 4681 7301 4682 7305
rect 4686 7301 4687 7305
rect 4691 7301 4692 7305
rect 4696 7301 4697 7305
rect 4701 7301 4702 7305
rect 4706 7301 4707 7305
rect 4711 7301 4712 7305
rect 4716 7301 4717 7305
rect 4721 7301 4722 7305
rect 4726 7301 4727 7305
rect 4731 7301 4732 7305
rect 4736 7301 4737 7305
rect 4741 7301 4742 7305
rect 4657 7300 4746 7301
rect 4661 7296 4662 7300
rect 4666 7296 4667 7300
rect 4671 7296 4672 7300
rect 4676 7296 4677 7300
rect 4681 7296 4682 7300
rect 4686 7296 4687 7300
rect 4691 7296 4692 7300
rect 4696 7296 4697 7300
rect 4701 7296 4702 7300
rect 4706 7296 4707 7300
rect 4711 7296 4712 7300
rect 4716 7296 4717 7300
rect 4721 7296 4722 7300
rect 4726 7296 4727 7300
rect 4731 7296 4732 7300
rect 4736 7296 4737 7300
rect 4741 7296 4742 7300
rect 4657 7295 4746 7296
rect 4661 7291 4662 7295
rect 4666 7291 4667 7295
rect 4671 7291 4672 7295
rect 4676 7291 4677 7295
rect 4681 7291 4682 7295
rect 4686 7291 4687 7295
rect 4691 7291 4692 7295
rect 4696 7291 4697 7295
rect 4701 7291 4702 7295
rect 4706 7291 4707 7295
rect 4711 7291 4712 7295
rect 4716 7291 4717 7295
rect 4721 7291 4722 7295
rect 4726 7291 4727 7295
rect 4731 7291 4732 7295
rect 4736 7291 4737 7295
rect 4741 7291 4742 7295
rect 4657 7290 4746 7291
rect 4661 7286 4662 7290
rect 4666 7286 4667 7290
rect 4671 7286 4672 7290
rect 4676 7286 4677 7290
rect 4681 7286 4682 7290
rect 4686 7286 4687 7290
rect 4691 7286 4692 7290
rect 4696 7286 4697 7290
rect 4701 7286 4702 7290
rect 4706 7286 4707 7290
rect 4711 7286 4712 7290
rect 4716 7286 4717 7290
rect 4721 7286 4722 7290
rect 4726 7286 4727 7290
rect 4731 7286 4732 7290
rect 4736 7286 4737 7290
rect 4741 7286 4742 7290
rect 4657 7285 4746 7286
rect 4661 7281 4662 7285
rect 4666 7281 4667 7285
rect 4671 7281 4672 7285
rect 4676 7281 4677 7285
rect 4681 7281 4682 7285
rect 4686 7281 4687 7285
rect 4691 7281 4692 7285
rect 4696 7281 4697 7285
rect 4701 7281 4702 7285
rect 4706 7281 4707 7285
rect 4711 7281 4712 7285
rect 4716 7281 4717 7285
rect 4721 7281 4722 7285
rect 4726 7281 4727 7285
rect 4731 7281 4732 7285
rect 4736 7281 4737 7285
rect 4741 7281 4742 7285
rect 4657 7280 4746 7281
rect 4661 7276 4662 7280
rect 4666 7276 4667 7280
rect 4671 7276 4672 7280
rect 4676 7276 4677 7280
rect 4681 7276 4682 7280
rect 4686 7276 4687 7280
rect 4691 7276 4692 7280
rect 4696 7276 4697 7280
rect 4701 7276 4702 7280
rect 4706 7276 4707 7280
rect 4711 7276 4712 7280
rect 4716 7276 4717 7280
rect 4721 7276 4722 7280
rect 4726 7276 4727 7280
rect 4731 7276 4732 7280
rect 4736 7276 4737 7280
rect 4741 7276 4742 7280
rect 4657 7275 4746 7276
rect 4661 7271 4662 7275
rect 4666 7271 4667 7275
rect 4671 7271 4672 7275
rect 4676 7271 4677 7275
rect 4681 7271 4682 7275
rect 4686 7271 4687 7275
rect 4691 7271 4692 7275
rect 4696 7271 4697 7275
rect 4701 7271 4702 7275
rect 4706 7271 4707 7275
rect 4711 7271 4712 7275
rect 4716 7271 4717 7275
rect 4721 7271 4722 7275
rect 4726 7271 4727 7275
rect 4731 7271 4732 7275
rect 4736 7271 4737 7275
rect 4741 7271 4742 7275
rect 4657 7270 4746 7271
rect 4661 7266 4662 7270
rect 4666 7266 4667 7270
rect 4671 7266 4672 7270
rect 4676 7266 4677 7270
rect 4681 7266 4682 7270
rect 4686 7266 4687 7270
rect 4691 7266 4692 7270
rect 4696 7266 4697 7270
rect 4701 7266 4702 7270
rect 4706 7266 4707 7270
rect 4711 7266 4712 7270
rect 4716 7266 4717 7270
rect 4721 7266 4722 7270
rect 4726 7266 4727 7270
rect 4731 7266 4732 7270
rect 4736 7266 4737 7270
rect 4741 7266 4742 7270
rect 4657 7265 4746 7266
rect 4661 7261 4662 7265
rect 4666 7261 4667 7265
rect 4671 7261 4672 7265
rect 4676 7261 4677 7265
rect 4681 7261 4682 7265
rect 4686 7261 4687 7265
rect 4691 7261 4692 7265
rect 4696 7261 4697 7265
rect 4701 7261 4702 7265
rect 4706 7261 4707 7265
rect 4711 7261 4712 7265
rect 4716 7261 4717 7265
rect 4721 7261 4722 7265
rect 4726 7261 4727 7265
rect 4731 7261 4732 7265
rect 4736 7261 4737 7265
rect 4741 7261 4742 7265
rect 4754 7305 4758 7306
rect 4754 7300 4758 7301
rect 4754 7295 4758 7296
rect 4754 7290 4758 7291
rect 4754 7285 4758 7286
rect 4754 7280 4758 7281
rect 4754 7275 4758 7276
rect 4754 7270 4758 7271
rect 4754 7265 4758 7266
rect 4641 7260 4649 7261
rect 4641 7253 4649 7256
rect 4754 7260 4758 7261
rect 4754 7253 4758 7256
rect 4649 7249 4652 7253
rect 4656 7249 4657 7253
rect 4661 7249 4662 7253
rect 4666 7249 4667 7253
rect 4671 7249 4672 7253
rect 4676 7249 4677 7253
rect 4681 7249 4682 7253
rect 4686 7249 4687 7253
rect 4691 7249 4692 7253
rect 4696 7249 4697 7253
rect 4701 7249 4702 7253
rect 4706 7249 4707 7253
rect 4711 7249 4712 7253
rect 4716 7249 4717 7253
rect 4721 7249 4722 7253
rect 4726 7249 4727 7253
rect 4731 7249 4732 7253
rect 4736 7249 4737 7253
rect 4741 7249 4742 7253
rect 4746 7249 4747 7253
rect 4751 7249 4754 7253
rect 4767 7315 4771 7316
rect 4774 7327 4775 7331
rect 4779 7327 4780 7331
rect 4784 7327 4785 7331
rect 4789 7327 4790 7331
rect 4794 7327 4829 7331
rect 4774 7324 4829 7327
rect 4774 7320 4775 7324
rect 4779 7320 4780 7324
rect 4784 7320 4785 7324
rect 4789 7320 4790 7324
rect 4794 7320 4829 7324
rect 4774 7315 4829 7320
rect 4767 7310 4771 7311
rect 4767 7305 4771 7306
rect 4786 7305 4829 7315
rect 4767 7300 4771 7301
rect 4767 7295 4771 7296
rect 4796 7295 4829 7305
rect 4767 7290 4771 7291
rect 4767 7285 4771 7286
rect 4806 7285 4829 7295
rect 4767 7280 4771 7281
rect 4767 7275 4771 7276
rect 4816 7275 4829 7285
rect 4767 7270 4771 7271
rect 4767 7265 4771 7266
rect 4767 7260 4771 7261
rect 4767 7255 4771 7256
rect 4767 7250 4771 7251
rect 4515 7245 4636 7246
rect 4515 7244 4632 7245
rect 4505 7243 4632 7244
rect 4505 7239 4506 7243
rect 4510 7239 4511 7243
rect 4515 7241 4632 7243
rect 4515 7240 4636 7241
rect 4767 7245 4771 7246
rect 4767 7240 4771 7241
rect 4515 7239 4632 7240
rect 4505 7237 4632 7239
rect 4636 7236 4637 7240
rect 4641 7236 4642 7240
rect 4646 7236 4647 7240
rect 4651 7236 4652 7240
rect 4656 7236 4657 7240
rect 4661 7236 4662 7240
rect 4666 7236 4667 7240
rect 4671 7236 4672 7240
rect 4676 7236 4677 7240
rect 4681 7236 4682 7240
rect 4686 7236 4687 7240
rect 4691 7236 4692 7240
rect 4696 7236 4697 7240
rect 4701 7236 4702 7240
rect 4706 7236 4707 7240
rect 4711 7236 4712 7240
rect 4716 7236 4717 7240
rect 4721 7236 4722 7240
rect 4726 7236 4727 7240
rect 4731 7236 4732 7240
rect 4736 7236 4737 7240
rect 4741 7236 4742 7240
rect 4746 7236 4747 7240
rect 4751 7236 4752 7240
rect 4756 7236 4757 7240
rect 4761 7236 4762 7240
rect 4766 7236 4767 7240
rect 4826 7236 4829 7275
rect 5083 7236 5086 7490
rect 343 7196 346 7235
rect 4483 7230 4484 7234
rect 4488 7230 4489 7234
rect 4493 7230 4494 7234
rect 4498 7230 4499 7234
rect 4503 7230 4504 7234
rect 4508 7230 4509 7234
rect 4479 7229 4513 7230
rect 4483 7225 4484 7229
rect 4488 7225 4489 7229
rect 4493 7225 4494 7229
rect 4498 7225 4499 7229
rect 4503 7225 4504 7229
rect 4508 7225 4509 7229
rect 4479 7224 4513 7225
rect 4483 7220 4484 7224
rect 4488 7220 4489 7224
rect 4493 7220 4494 7224
rect 4498 7220 4499 7224
rect 4503 7220 4504 7224
rect 4508 7220 4509 7224
rect 4479 7219 4513 7220
rect 4483 7215 4484 7219
rect 4488 7215 4489 7219
rect 4493 7215 4494 7219
rect 4498 7215 4499 7219
rect 4503 7215 4504 7219
rect 4508 7215 4509 7219
rect 4529 7230 4530 7234
rect 4534 7230 4535 7234
rect 4539 7230 4540 7234
rect 4544 7230 4545 7234
rect 4549 7230 4550 7234
rect 4554 7230 4555 7234
rect 4826 7233 5086 7236
rect 4525 7229 4559 7230
rect 4529 7225 4530 7229
rect 4534 7225 4535 7229
rect 4539 7225 4540 7229
rect 4544 7225 4545 7229
rect 4549 7225 4550 7229
rect 4554 7225 4555 7229
rect 4525 7224 4559 7225
rect 4529 7220 4530 7224
rect 4534 7220 4535 7224
rect 4539 7220 4540 7224
rect 4544 7220 4545 7224
rect 4549 7220 4550 7224
rect 4554 7220 4555 7224
rect 4525 7219 4559 7220
rect 4529 7215 4530 7219
rect 4534 7215 4535 7219
rect 4539 7215 4540 7219
rect 4544 7215 4545 7219
rect 4549 7215 4550 7219
rect 4554 7215 4555 7219
rect 86 7193 346 7196
rect 4483 7202 4484 7206
rect 4488 7202 4489 7206
rect 4493 7202 4494 7206
rect 4498 7202 4499 7206
rect 4503 7202 4504 7206
rect 4508 7202 4509 7206
rect 4479 7201 4513 7202
rect 4483 7197 4484 7201
rect 4488 7197 4489 7201
rect 4493 7197 4494 7201
rect 4498 7197 4499 7201
rect 4503 7197 4504 7201
rect 4508 7197 4509 7201
rect 4479 7196 4513 7197
rect 4483 7192 4484 7196
rect 4488 7192 4489 7196
rect 4493 7192 4494 7196
rect 4498 7192 4499 7196
rect 4503 7192 4504 7196
rect 4508 7192 4509 7196
rect 4479 7191 4513 7192
rect 4483 7187 4484 7191
rect 4488 7187 4489 7191
rect 4493 7187 4494 7191
rect 4498 7187 4499 7191
rect 4503 7187 4504 7191
rect 4508 7187 4509 7191
rect 4529 7202 4530 7206
rect 4534 7202 4535 7206
rect 4539 7202 4540 7206
rect 4544 7202 4545 7206
rect 4549 7202 4550 7206
rect 4554 7202 4555 7206
rect 4525 7201 4559 7202
rect 4529 7197 4530 7201
rect 4534 7197 4535 7201
rect 4539 7197 4540 7201
rect 4544 7197 4545 7201
rect 4549 7197 4550 7201
rect 4554 7197 4555 7201
rect 4525 7196 4559 7197
rect 4529 7192 4530 7196
rect 4534 7192 4535 7196
rect 4539 7192 4540 7196
rect 4544 7192 4545 7196
rect 4549 7192 4550 7196
rect 4554 7192 4555 7196
rect 4525 7191 4559 7192
rect 4529 7187 4530 7191
rect 4534 7187 4535 7191
rect 4539 7187 4540 7191
rect 4544 7187 4545 7191
rect 4549 7187 4550 7191
rect 4554 7187 4555 7191
rect 617 7158 618 7162
rect 622 7158 623 7162
rect 627 7158 628 7162
rect 632 7158 633 7162
rect 637 7158 638 7162
rect 642 7158 643 7162
rect 613 7157 647 7158
rect 663 7158 664 7162
rect 668 7158 669 7162
rect 673 7158 674 7162
rect 678 7158 679 7162
rect 683 7158 684 7162
rect 688 7158 689 7162
rect 659 7157 693 7158
rect 4479 7156 4513 7157
rect 4483 7152 4484 7156
rect 4488 7152 4489 7156
rect 4493 7152 4494 7156
rect 4498 7152 4499 7156
rect 4503 7152 4504 7156
rect 4508 7152 4509 7156
rect 4525 7156 4559 7157
rect 4529 7152 4530 7156
rect 4534 7152 4535 7156
rect 4539 7152 4540 7156
rect 4544 7152 4545 7156
rect 4549 7152 4550 7156
rect 4554 7152 4555 7156
rect 617 7123 618 7127
rect 622 7123 623 7127
rect 627 7123 628 7127
rect 632 7123 633 7127
rect 637 7123 638 7127
rect 642 7123 643 7127
rect 613 7122 647 7123
rect 617 7118 618 7122
rect 622 7118 623 7122
rect 627 7118 628 7122
rect 632 7118 633 7122
rect 637 7118 638 7122
rect 642 7118 643 7122
rect 613 7117 647 7118
rect 617 7113 618 7117
rect 622 7113 623 7117
rect 627 7113 628 7117
rect 632 7113 633 7117
rect 637 7113 638 7117
rect 642 7113 643 7117
rect 613 7112 647 7113
rect 86 7106 346 7109
rect 617 7108 618 7112
rect 622 7108 623 7112
rect 627 7108 628 7112
rect 632 7108 633 7112
rect 637 7108 638 7112
rect 642 7108 643 7112
rect 663 7123 664 7127
rect 668 7123 669 7127
rect 673 7123 674 7127
rect 678 7123 679 7127
rect 683 7123 684 7127
rect 688 7123 689 7127
rect 659 7122 693 7123
rect 663 7118 664 7122
rect 668 7118 669 7122
rect 673 7118 674 7122
rect 678 7118 679 7122
rect 683 7118 684 7122
rect 688 7118 689 7122
rect 659 7117 693 7118
rect 663 7113 664 7117
rect 668 7113 669 7117
rect 673 7113 674 7117
rect 678 7113 679 7117
rect 683 7113 684 7117
rect 688 7113 689 7117
rect 659 7112 693 7113
rect 663 7108 664 7112
rect 668 7108 669 7112
rect 673 7108 674 7112
rect 678 7108 679 7112
rect 683 7108 684 7112
rect 688 7108 689 7112
rect 4826 7118 5086 7121
rect 86 6852 89 7106
rect 343 7067 346 7106
rect 4826 7079 4829 7118
rect 4816 7069 4829 7079
rect 343 7057 356 7067
rect 4806 7059 4829 7069
rect 343 7047 366 7057
rect 4796 7049 4829 7059
rect 343 7037 376 7047
rect 4786 7039 4829 7049
rect 343 7027 386 7037
rect 343 6931 769 7027
rect 4403 6943 4829 7039
rect 4786 6933 4829 6943
rect 343 6921 386 6931
rect 4796 6923 4829 6933
rect 343 6911 376 6921
rect 1415 6919 1485 6923
rect 1489 6919 1535 6923
rect 1539 6919 1586 6923
rect 1590 6919 1617 6923
rect 1621 6919 1667 6923
rect 1671 6919 1718 6923
rect 1722 6919 1749 6923
rect 1753 6919 1799 6923
rect 1803 6919 1850 6923
rect 1854 6919 1863 6923
rect 2360 6919 2430 6923
rect 2434 6919 2480 6923
rect 2484 6919 2531 6923
rect 2535 6919 2562 6923
rect 2566 6919 2612 6923
rect 2616 6919 2663 6923
rect 2667 6919 2694 6923
rect 2698 6919 2744 6923
rect 2748 6919 2795 6923
rect 2799 6919 2808 6923
rect 1451 6912 1504 6916
rect 1508 6912 1534 6916
rect 1538 6912 1562 6916
rect 1566 6912 1636 6916
rect 1640 6912 1666 6916
rect 1670 6912 1694 6916
rect 1698 6912 1768 6916
rect 1772 6912 1798 6916
rect 1802 6912 1826 6916
rect 1830 6912 1863 6916
rect 2396 6912 2449 6916
rect 2453 6912 2479 6916
rect 2483 6912 2507 6916
rect 2511 6912 2581 6916
rect 2585 6912 2611 6916
rect 2615 6912 2639 6916
rect 2643 6912 2713 6916
rect 2717 6912 2743 6916
rect 2747 6912 2771 6916
rect 2775 6912 2808 6916
rect 4806 6913 4829 6923
rect 343 6901 366 6911
rect 343 6891 356 6901
rect 1477 6900 1480 6912
rect 1498 6900 1501 6912
rect 1514 6900 1517 6912
rect 1533 6906 1545 6909
rect 1556 6900 1559 6912
rect 1572 6900 1575 6912
rect 1593 6900 1596 6912
rect 1609 6900 1612 6912
rect 1630 6900 1633 6912
rect 1646 6900 1649 6912
rect 1665 6906 1677 6909
rect 1688 6900 1691 6912
rect 1704 6900 1707 6912
rect 1725 6900 1728 6912
rect 1741 6900 1744 6912
rect 1762 6900 1765 6912
rect 1778 6900 1781 6912
rect 1797 6906 1809 6909
rect 1820 6900 1823 6912
rect 1836 6900 1839 6912
rect 1857 6900 1860 6912
rect 2422 6900 2425 6912
rect 2443 6900 2446 6912
rect 2459 6900 2462 6912
rect 2478 6906 2490 6909
rect 2501 6900 2504 6912
rect 2517 6900 2520 6912
rect 2538 6900 2541 6912
rect 2554 6900 2557 6912
rect 2575 6900 2578 6912
rect 2591 6900 2594 6912
rect 2610 6906 2622 6909
rect 2633 6900 2636 6912
rect 2649 6900 2652 6912
rect 2670 6900 2673 6912
rect 2686 6900 2689 6912
rect 2707 6900 2710 6912
rect 2723 6900 2726 6912
rect 2742 6906 2754 6909
rect 2765 6900 2768 6912
rect 2781 6900 2784 6912
rect 2802 6900 2805 6912
rect 4816 6903 4829 6913
rect 343 6852 346 6891
rect 1477 6886 1494 6889
rect 1498 6890 1505 6893
rect 1530 6890 1533 6896
rect 1533 6886 1552 6889
rect 1556 6890 1563 6893
rect 1611 6886 1626 6889
rect 1630 6890 1637 6893
rect 1662 6890 1665 6896
rect 1665 6886 1684 6889
rect 1688 6890 1695 6893
rect 1743 6886 1758 6889
rect 1762 6890 1769 6893
rect 1794 6890 1797 6896
rect 1797 6886 1816 6889
rect 1820 6890 1827 6893
rect 1488 6880 1510 6883
rect 1514 6880 1521 6883
rect 1546 6880 1570 6883
rect 1574 6880 1579 6883
rect 1593 6880 1600 6883
rect 1620 6880 1642 6883
rect 1646 6880 1653 6883
rect 1678 6880 1702 6883
rect 1706 6880 1711 6883
rect 1725 6880 1732 6883
rect 1752 6880 1774 6883
rect 1778 6880 1785 6883
rect 1810 6880 1834 6883
rect 1838 6880 1843 6883
rect 2422 6886 2439 6889
rect 2443 6890 2450 6893
rect 2475 6890 2478 6896
rect 2478 6886 2497 6889
rect 2501 6890 2508 6893
rect 2556 6886 2571 6889
rect 2575 6890 2582 6893
rect 2607 6890 2610 6896
rect 2610 6886 2629 6889
rect 2633 6890 2640 6893
rect 2688 6886 2703 6889
rect 2707 6890 2714 6893
rect 2739 6890 2742 6896
rect 2742 6886 2761 6889
rect 2765 6890 2772 6893
rect 2433 6880 2455 6883
rect 2459 6880 2466 6883
rect 2491 6880 2515 6883
rect 2519 6880 2524 6883
rect 2538 6880 2545 6883
rect 2565 6880 2587 6883
rect 2591 6880 2598 6883
rect 2623 6880 2647 6883
rect 2651 6880 2656 6883
rect 2670 6880 2677 6883
rect 2697 6880 2719 6883
rect 2723 6880 2730 6883
rect 2755 6880 2779 6883
rect 2783 6880 2788 6883
rect 1477 6859 1480 6869
rect 1498 6859 1501 6869
rect 1514 6859 1517 6869
rect 1529 6862 1536 6866
rect 1540 6862 1545 6866
rect 1556 6859 1559 6869
rect 1572 6859 1575 6869
rect 1593 6859 1596 6869
rect 1609 6859 1612 6869
rect 1630 6859 1633 6869
rect 1646 6859 1649 6869
rect 1661 6862 1668 6866
rect 1672 6862 1677 6866
rect 1688 6859 1691 6869
rect 1704 6859 1707 6869
rect 1725 6859 1728 6869
rect 1741 6859 1744 6869
rect 1762 6859 1765 6869
rect 1778 6859 1781 6869
rect 1793 6862 1800 6866
rect 1804 6862 1809 6866
rect 1820 6859 1823 6869
rect 1836 6859 1839 6869
rect 1857 6859 1860 6869
rect 2422 6859 2425 6869
rect 2443 6859 2446 6869
rect 2459 6859 2462 6869
rect 2474 6862 2481 6866
rect 2485 6862 2490 6866
rect 2501 6859 2504 6869
rect 2517 6859 2520 6869
rect 2538 6859 2541 6869
rect 2554 6859 2557 6869
rect 2575 6859 2578 6869
rect 2591 6859 2594 6869
rect 2606 6862 2613 6866
rect 2617 6862 2622 6866
rect 2633 6859 2636 6869
rect 2649 6859 2652 6869
rect 2670 6859 2673 6869
rect 2686 6859 2689 6869
rect 2707 6859 2710 6869
rect 2723 6859 2726 6869
rect 2738 6862 2745 6866
rect 2749 6862 2754 6866
rect 2765 6859 2768 6869
rect 2781 6859 2784 6869
rect 2802 6859 2805 6869
rect 4826 6864 4829 6903
rect 5083 6864 5086 7118
rect 1463 6855 1467 6859
rect 1471 6855 1504 6859
rect 1508 6855 1534 6859
rect 1538 6855 1562 6859
rect 1566 6855 1599 6859
rect 1603 6855 1636 6859
rect 1640 6855 1666 6859
rect 1670 6855 1694 6859
rect 1698 6855 1731 6859
rect 1735 6855 1768 6859
rect 1772 6855 1798 6859
rect 1802 6855 1826 6859
rect 1830 6855 1863 6859
rect 2408 6855 2412 6859
rect 2416 6855 2449 6859
rect 2453 6855 2479 6859
rect 2483 6855 2507 6859
rect 2511 6855 2544 6859
rect 2548 6855 2581 6859
rect 2585 6855 2611 6859
rect 2615 6855 2639 6859
rect 2643 6855 2676 6859
rect 2680 6855 2713 6859
rect 2717 6855 2743 6859
rect 2747 6855 2771 6859
rect 2775 6855 2808 6859
rect 4483 6858 4484 6862
rect 4488 6858 4489 6862
rect 4493 6858 4494 6862
rect 4498 6858 4499 6862
rect 4503 6858 4504 6862
rect 4508 6858 4509 6862
rect 4479 6857 4513 6858
rect 4483 6853 4484 6857
rect 4488 6853 4489 6857
rect 4493 6853 4494 6857
rect 4498 6853 4499 6857
rect 4503 6853 4504 6857
rect 4508 6853 4509 6857
rect 4479 6852 4513 6853
rect 86 6849 346 6852
rect 1403 6848 1483 6852
rect 1487 6848 1550 6852
rect 1554 6848 1586 6852
rect 1590 6848 1615 6852
rect 1619 6848 1682 6852
rect 1686 6848 1718 6852
rect 1722 6848 1747 6852
rect 1751 6848 1814 6852
rect 1818 6848 1850 6852
rect 1854 6848 1863 6852
rect 2348 6848 2428 6852
rect 2432 6848 2495 6852
rect 2499 6848 2531 6852
rect 2535 6848 2560 6852
rect 2564 6848 2627 6852
rect 2631 6848 2663 6852
rect 2667 6848 2692 6852
rect 2696 6848 2759 6852
rect 2763 6848 2795 6852
rect 2799 6848 2808 6852
rect 4483 6848 4484 6852
rect 4488 6848 4489 6852
rect 4493 6848 4494 6852
rect 4498 6848 4499 6852
rect 4503 6848 4504 6852
rect 4508 6848 4509 6852
rect 4479 6847 4513 6848
rect 1628 6842 1732 6845
rect 2573 6842 2677 6845
rect 4483 6843 4484 6847
rect 4488 6843 4489 6847
rect 4493 6843 4494 6847
rect 4498 6843 4499 6847
rect 4503 6843 4504 6847
rect 4508 6843 4509 6847
rect 4529 6858 4530 6862
rect 4534 6858 4535 6862
rect 4539 6858 4540 6862
rect 4544 6858 4545 6862
rect 4549 6858 4550 6862
rect 4554 6858 4555 6862
rect 4826 6861 5086 6864
rect 4525 6857 4559 6858
rect 4529 6853 4530 6857
rect 4534 6853 4535 6857
rect 4539 6853 4540 6857
rect 4544 6853 4545 6857
rect 4549 6853 4550 6857
rect 4554 6853 4555 6857
rect 4525 6852 4559 6853
rect 4529 6848 4530 6852
rect 4534 6848 4535 6852
rect 4539 6848 4540 6852
rect 4544 6848 4545 6852
rect 4549 6848 4550 6852
rect 4554 6848 4555 6852
rect 4525 6847 4559 6848
rect 4529 6843 4530 6847
rect 4534 6843 4535 6847
rect 4539 6843 4540 6847
rect 4544 6843 4545 6847
rect 4549 6843 4550 6847
rect 4554 6843 4555 6847
rect 1604 6834 1608 6838
rect 1612 6834 1616 6838
rect 2549 6834 2553 6838
rect 2557 6834 2561 6838
rect 1472 6826 1585 6829
rect 2417 6826 2530 6829
rect 1472 6819 1600 6822
rect 2417 6819 2545 6822
rect 812 6811 927 6815
rect 931 6811 1592 6815
rect 1608 6811 1624 6815
rect 1628 6811 1872 6815
rect 1876 6811 2537 6815
rect 2553 6811 2569 6815
rect 2573 6811 2825 6815
rect 4826 6809 5086 6812
rect 1604 6800 1608 6804
rect 1612 6800 1616 6804
rect 2549 6800 2553 6804
rect 2557 6800 2561 6804
rect 86 6796 346 6799
rect 86 6542 89 6796
rect 343 6757 346 6796
rect 1628 6793 1732 6796
rect 2573 6793 2677 6796
rect 1472 6786 1857 6789
rect 2417 6786 2802 6789
rect 1415 6779 1485 6783
rect 1489 6779 1535 6783
rect 1539 6779 1586 6783
rect 1590 6779 1617 6783
rect 1621 6779 1667 6783
rect 1671 6779 1718 6783
rect 1722 6779 1749 6783
rect 1753 6779 1799 6783
rect 1803 6779 1850 6783
rect 1854 6779 1863 6783
rect 2360 6779 2430 6783
rect 2434 6779 2480 6783
rect 2484 6779 2531 6783
rect 2535 6779 2562 6783
rect 2566 6779 2612 6783
rect 2616 6779 2663 6783
rect 2667 6779 2694 6783
rect 2698 6779 2744 6783
rect 2748 6779 2795 6783
rect 2799 6779 2808 6783
rect 1451 6772 1504 6776
rect 1508 6772 1534 6776
rect 1538 6772 1562 6776
rect 1566 6772 1636 6776
rect 1640 6772 1666 6776
rect 1670 6772 1694 6776
rect 1698 6772 1768 6776
rect 1772 6772 1798 6776
rect 1802 6772 1826 6776
rect 1830 6772 1863 6776
rect 2396 6772 2449 6776
rect 2453 6772 2479 6776
rect 2483 6772 2507 6776
rect 2511 6772 2581 6776
rect 2585 6772 2611 6776
rect 2615 6772 2639 6776
rect 2643 6772 2713 6776
rect 2717 6772 2743 6776
rect 2747 6772 2771 6776
rect 2775 6772 2808 6776
rect 1477 6760 1480 6772
rect 1498 6760 1501 6772
rect 1514 6760 1517 6772
rect 1533 6766 1545 6769
rect 1556 6760 1559 6772
rect 1572 6760 1575 6772
rect 1593 6760 1596 6772
rect 1609 6760 1612 6772
rect 1630 6760 1633 6772
rect 1646 6760 1649 6772
rect 1665 6766 1677 6769
rect 1688 6760 1691 6772
rect 1704 6760 1707 6772
rect 1725 6760 1728 6772
rect 1741 6760 1744 6772
rect 1762 6760 1765 6772
rect 1778 6760 1781 6772
rect 1797 6766 1809 6769
rect 1820 6760 1823 6772
rect 1836 6760 1839 6772
rect 1857 6760 1860 6772
rect 2422 6760 2425 6772
rect 2443 6760 2446 6772
rect 2459 6760 2462 6772
rect 2478 6766 2490 6769
rect 2501 6760 2504 6772
rect 2517 6760 2520 6772
rect 2538 6760 2541 6772
rect 2554 6760 2557 6772
rect 2575 6760 2578 6772
rect 2591 6760 2594 6772
rect 2610 6766 2622 6769
rect 2633 6760 2636 6772
rect 2649 6760 2652 6772
rect 2670 6760 2673 6772
rect 2686 6760 2689 6772
rect 2707 6760 2710 6772
rect 2723 6760 2726 6772
rect 2742 6766 2754 6769
rect 2765 6760 2768 6772
rect 2781 6760 2784 6772
rect 2802 6760 2805 6772
rect 4826 6770 4829 6809
rect 4816 6760 4829 6770
rect 343 6747 356 6757
rect 948 6749 966 6753
rect 970 6749 1016 6753
rect 1020 6749 1067 6753
rect 1071 6749 1409 6753
rect 343 6737 366 6747
rect 948 6742 985 6746
rect 989 6742 1015 6746
rect 1019 6742 1043 6746
rect 1047 6742 1445 6746
rect 1477 6746 1494 6749
rect 1498 6750 1505 6753
rect 1530 6750 1533 6756
rect 1533 6746 1552 6749
rect 1556 6750 1563 6753
rect 1611 6746 1626 6749
rect 1630 6750 1637 6753
rect 1662 6750 1665 6756
rect 1665 6746 1684 6749
rect 1688 6750 1695 6753
rect 1743 6746 1758 6749
rect 1762 6750 1769 6753
rect 1794 6750 1797 6756
rect 1797 6746 1816 6749
rect 1820 6750 1827 6753
rect 1893 6749 1911 6753
rect 1915 6749 1961 6753
rect 1965 6749 2012 6753
rect 2016 6749 2354 6753
rect 343 6727 376 6737
rect 958 6730 961 6742
rect 979 6730 982 6742
rect 995 6730 998 6742
rect 1014 6736 1026 6739
rect 1037 6730 1040 6742
rect 1053 6730 1056 6742
rect 1074 6730 1077 6742
rect 343 6717 386 6727
rect 938 6717 949 6721
rect 343 6679 769 6717
rect 960 6716 975 6719
rect 979 6720 986 6723
rect 1011 6720 1014 6726
rect 1488 6740 1510 6743
rect 1514 6740 1521 6743
rect 1546 6740 1570 6743
rect 1574 6740 1579 6743
rect 1593 6740 1600 6743
rect 1620 6740 1642 6743
rect 1646 6740 1653 6743
rect 1678 6740 1702 6743
rect 1706 6740 1711 6743
rect 1725 6740 1732 6743
rect 1752 6740 1774 6743
rect 1778 6740 1785 6743
rect 1810 6740 1834 6743
rect 1838 6740 1843 6743
rect 1893 6742 1930 6746
rect 1934 6742 1960 6746
rect 1964 6742 1988 6746
rect 1992 6742 2390 6746
rect 2422 6746 2439 6749
rect 2443 6750 2450 6753
rect 2475 6750 2478 6756
rect 2478 6746 2497 6749
rect 2501 6750 2508 6753
rect 2556 6746 2571 6749
rect 2575 6750 2582 6753
rect 2607 6750 2610 6756
rect 2610 6746 2629 6749
rect 2633 6750 2640 6753
rect 2688 6746 2703 6749
rect 2707 6750 2714 6753
rect 2739 6750 2742 6756
rect 2742 6746 2761 6749
rect 2765 6750 2772 6753
rect 4806 6750 4829 6760
rect 1903 6730 1906 6742
rect 1924 6730 1927 6742
rect 1940 6730 1943 6742
rect 1959 6736 1971 6739
rect 1982 6730 1985 6742
rect 1998 6730 2001 6742
rect 2019 6730 2022 6742
rect 1014 6716 1033 6719
rect 1037 6720 1044 6723
rect 1477 6719 1480 6729
rect 1498 6719 1501 6729
rect 1514 6719 1517 6729
rect 1529 6722 1536 6726
rect 1540 6722 1545 6726
rect 1556 6719 1559 6729
rect 1572 6719 1575 6729
rect 1593 6719 1596 6729
rect 1609 6719 1612 6729
rect 1630 6719 1633 6729
rect 1646 6719 1649 6729
rect 1661 6722 1668 6726
rect 1672 6722 1677 6726
rect 1688 6719 1691 6729
rect 1704 6719 1707 6729
rect 1725 6719 1728 6729
rect 1741 6719 1744 6729
rect 1762 6719 1765 6729
rect 1778 6719 1781 6729
rect 1793 6722 1800 6726
rect 1804 6722 1809 6726
rect 1820 6719 1823 6729
rect 1836 6719 1839 6729
rect 1857 6719 1860 6729
rect 969 6710 991 6713
rect 995 6710 1002 6713
rect 1027 6710 1051 6713
rect 1055 6710 1060 6713
rect 1463 6715 1467 6719
rect 1471 6715 1504 6719
rect 1508 6715 1534 6719
rect 1538 6715 1562 6719
rect 1566 6715 1599 6719
rect 1603 6715 1636 6719
rect 1640 6715 1666 6719
rect 1670 6715 1694 6719
rect 1698 6715 1731 6719
rect 1735 6715 1768 6719
rect 1772 6715 1798 6719
rect 1802 6715 1826 6719
rect 1830 6715 1863 6719
rect 1883 6717 1894 6721
rect 1905 6716 1920 6719
rect 1924 6720 1931 6723
rect 1956 6720 1959 6726
rect 2433 6740 2455 6743
rect 2459 6740 2466 6743
rect 2491 6740 2515 6743
rect 2519 6740 2524 6743
rect 2538 6740 2545 6743
rect 2565 6740 2587 6743
rect 2591 6740 2598 6743
rect 2623 6740 2647 6743
rect 2651 6740 2656 6743
rect 2670 6740 2677 6743
rect 2697 6740 2719 6743
rect 2723 6740 2730 6743
rect 2755 6740 2779 6743
rect 2783 6740 2788 6743
rect 4796 6740 4829 6750
rect 4786 6730 4829 6740
rect 1959 6716 1978 6719
rect 1982 6720 1989 6723
rect 2422 6719 2425 6729
rect 2443 6719 2446 6729
rect 2459 6719 2462 6729
rect 2474 6722 2481 6726
rect 2485 6722 2490 6726
rect 2501 6719 2504 6729
rect 2517 6719 2520 6729
rect 2538 6719 2541 6729
rect 2554 6719 2557 6729
rect 2575 6719 2578 6729
rect 2591 6719 2594 6729
rect 2606 6722 2613 6726
rect 2617 6722 2622 6726
rect 2633 6719 2636 6729
rect 2649 6719 2652 6729
rect 2670 6719 2673 6729
rect 2686 6719 2689 6729
rect 2707 6719 2710 6729
rect 2723 6719 2726 6729
rect 2738 6722 2745 6726
rect 2749 6722 2754 6726
rect 2765 6719 2768 6729
rect 2781 6719 2784 6729
rect 2802 6719 2805 6729
rect 1403 6708 1483 6712
rect 1487 6708 1550 6712
rect 1554 6708 1586 6712
rect 1590 6708 1615 6712
rect 1619 6708 1682 6712
rect 1686 6708 1718 6712
rect 1722 6708 1747 6712
rect 1751 6708 1814 6712
rect 1818 6708 1850 6712
rect 1854 6708 1863 6712
rect 1914 6710 1936 6713
rect 1940 6710 1947 6713
rect 1472 6701 1857 6704
rect 1972 6710 1996 6713
rect 2000 6710 2005 6713
rect 2408 6715 2412 6719
rect 2416 6715 2449 6719
rect 2453 6715 2479 6719
rect 2483 6715 2507 6719
rect 2511 6715 2544 6719
rect 2548 6715 2581 6719
rect 2585 6715 2611 6719
rect 2615 6715 2639 6719
rect 2643 6715 2676 6719
rect 2680 6715 2713 6719
rect 2717 6715 2743 6719
rect 2747 6715 2771 6719
rect 2775 6715 2808 6719
rect 2348 6708 2428 6712
rect 2432 6708 2495 6712
rect 2499 6708 2531 6712
rect 2535 6708 2560 6712
rect 2564 6708 2627 6712
rect 2631 6708 2663 6712
rect 2667 6708 2692 6712
rect 2696 6708 2759 6712
rect 2763 6708 2795 6712
rect 2799 6708 2808 6712
rect 2417 6701 2802 6704
rect 958 6689 961 6699
rect 979 6689 982 6699
rect 995 6689 998 6699
rect 1010 6692 1017 6696
rect 1021 6692 1026 6696
rect 1037 6689 1040 6699
rect 1053 6689 1056 6699
rect 1074 6689 1077 6699
rect 1415 6693 1485 6697
rect 1489 6693 1535 6697
rect 1539 6693 1586 6697
rect 1590 6693 1617 6697
rect 1621 6693 1667 6697
rect 1671 6693 1718 6697
rect 1722 6693 1749 6697
rect 1753 6693 1799 6697
rect 1803 6693 1850 6697
rect 1854 6693 1863 6697
rect 952 6685 985 6689
rect 989 6685 1015 6689
rect 1019 6685 1043 6689
rect 1047 6685 1081 6689
rect 1451 6686 1504 6690
rect 1508 6686 1534 6690
rect 1538 6686 1562 6690
rect 1566 6686 1636 6690
rect 1640 6686 1666 6690
rect 1670 6686 1694 6690
rect 1698 6686 1768 6690
rect 1772 6686 1798 6690
rect 1802 6686 1826 6690
rect 1830 6686 1863 6690
rect 1903 6689 1906 6699
rect 1924 6689 1927 6699
rect 1940 6689 1943 6699
rect 1955 6692 1962 6696
rect 1966 6692 1971 6696
rect 1982 6689 1985 6699
rect 1998 6689 2001 6699
rect 2019 6689 2022 6699
rect 2360 6693 2430 6697
rect 2434 6693 2480 6697
rect 2484 6693 2531 6697
rect 2535 6693 2562 6697
rect 2566 6693 2612 6697
rect 2616 6693 2663 6697
rect 2667 6693 2694 6697
rect 2698 6693 2744 6697
rect 2748 6693 2795 6697
rect 2799 6693 2808 6697
rect 343 6666 788 6679
rect 948 6678 964 6682
rect 968 6678 1031 6682
rect 1035 6678 1067 6682
rect 1071 6678 1397 6682
rect 953 6671 1074 6674
rect 1477 6674 1480 6686
rect 1498 6674 1501 6686
rect 1514 6674 1517 6686
rect 1533 6680 1545 6683
rect 1556 6674 1559 6686
rect 1572 6674 1575 6686
rect 1593 6674 1596 6686
rect 1609 6674 1612 6686
rect 1630 6674 1633 6686
rect 1646 6674 1649 6686
rect 1665 6680 1677 6683
rect 1688 6674 1691 6686
rect 1704 6674 1707 6686
rect 1725 6674 1728 6686
rect 1741 6674 1744 6686
rect 1762 6674 1765 6686
rect 1778 6674 1781 6686
rect 1797 6680 1809 6683
rect 1820 6674 1823 6686
rect 1836 6674 1839 6686
rect 1857 6674 1860 6686
rect 1897 6685 1930 6689
rect 1934 6685 1960 6689
rect 1964 6685 1988 6689
rect 1992 6685 2026 6689
rect 2396 6686 2449 6690
rect 2453 6686 2479 6690
rect 2483 6686 2507 6690
rect 2511 6686 2581 6690
rect 2585 6686 2611 6690
rect 2615 6686 2639 6690
rect 2643 6686 2713 6690
rect 2717 6686 2743 6690
rect 2747 6686 2771 6690
rect 2775 6686 2808 6690
rect 1893 6678 1909 6682
rect 1913 6678 1976 6682
rect 1980 6678 2012 6682
rect 2016 6678 2342 6682
rect 343 6621 769 6666
rect 948 6663 966 6667
rect 970 6663 1016 6667
rect 1020 6663 1067 6667
rect 1071 6663 1409 6667
rect 948 6656 985 6660
rect 989 6656 1015 6660
rect 1019 6656 1043 6660
rect 1047 6656 1445 6660
rect 1477 6660 1494 6663
rect 1498 6664 1505 6667
rect 1530 6664 1533 6670
rect 1533 6660 1552 6663
rect 1556 6664 1563 6667
rect 1611 6660 1626 6663
rect 1630 6664 1637 6667
rect 1662 6664 1665 6670
rect 1665 6660 1684 6663
rect 1688 6664 1695 6667
rect 1743 6660 1758 6663
rect 1762 6664 1769 6667
rect 1794 6664 1797 6670
rect 1898 6671 2019 6674
rect 2422 6674 2425 6686
rect 2443 6674 2446 6686
rect 2459 6674 2462 6686
rect 2478 6680 2490 6683
rect 2501 6674 2504 6686
rect 2517 6674 2520 6686
rect 2538 6674 2541 6686
rect 2554 6674 2557 6686
rect 2575 6674 2578 6686
rect 2591 6674 2594 6686
rect 2610 6680 2622 6683
rect 2633 6674 2636 6686
rect 2649 6674 2652 6686
rect 2670 6674 2673 6686
rect 2686 6674 2689 6686
rect 2707 6674 2710 6686
rect 2723 6674 2726 6686
rect 2742 6680 2754 6683
rect 2765 6674 2768 6686
rect 2781 6674 2784 6686
rect 2802 6674 2805 6686
rect 1797 6660 1816 6663
rect 1820 6664 1827 6667
rect 1893 6663 1911 6667
rect 1915 6663 1961 6667
rect 1965 6663 2012 6667
rect 2016 6663 2354 6667
rect 958 6644 961 6656
rect 979 6644 982 6656
rect 995 6644 998 6656
rect 1014 6650 1026 6653
rect 1037 6644 1040 6656
rect 1053 6644 1056 6656
rect 1074 6644 1077 6656
rect 960 6630 975 6633
rect 979 6634 986 6637
rect 1011 6634 1014 6640
rect 1488 6654 1510 6657
rect 1514 6654 1521 6657
rect 1546 6654 1570 6657
rect 1574 6654 1579 6657
rect 1593 6654 1600 6657
rect 1620 6654 1642 6657
rect 1646 6654 1653 6657
rect 1678 6654 1702 6657
rect 1706 6654 1711 6657
rect 1725 6654 1732 6657
rect 1752 6654 1774 6657
rect 1778 6654 1785 6657
rect 1810 6654 1834 6657
rect 1838 6654 1843 6657
rect 1893 6656 1930 6660
rect 1934 6656 1960 6660
rect 1964 6656 1988 6660
rect 1992 6656 2390 6660
rect 2422 6660 2439 6663
rect 2443 6664 2450 6667
rect 2475 6664 2478 6670
rect 2478 6660 2497 6663
rect 2501 6664 2508 6667
rect 2556 6660 2571 6663
rect 2575 6664 2582 6667
rect 2607 6664 2610 6670
rect 2610 6660 2629 6663
rect 2633 6664 2640 6667
rect 2688 6660 2703 6663
rect 2707 6664 2714 6667
rect 2739 6664 2742 6670
rect 2742 6660 2761 6663
rect 2765 6664 2772 6667
rect 1903 6644 1906 6656
rect 1924 6644 1927 6656
rect 1940 6644 1943 6656
rect 1959 6650 1971 6653
rect 1982 6644 1985 6656
rect 1998 6644 2001 6656
rect 2019 6644 2022 6656
rect 1014 6630 1033 6633
rect 1037 6634 1044 6637
rect 1477 6633 1480 6643
rect 1498 6633 1501 6643
rect 1514 6633 1517 6643
rect 1529 6636 1536 6640
rect 1540 6636 1545 6640
rect 1556 6633 1559 6643
rect 1572 6633 1575 6643
rect 1593 6633 1596 6643
rect 1609 6633 1612 6643
rect 1630 6633 1633 6643
rect 1646 6633 1649 6643
rect 1661 6636 1668 6640
rect 1672 6636 1677 6640
rect 1688 6633 1691 6643
rect 1704 6633 1707 6643
rect 1725 6633 1728 6643
rect 1741 6633 1744 6643
rect 1762 6633 1765 6643
rect 1778 6633 1781 6643
rect 1793 6636 1800 6640
rect 1804 6636 1809 6640
rect 1820 6633 1823 6643
rect 1836 6633 1839 6643
rect 1857 6633 1860 6643
rect 969 6624 991 6627
rect 995 6624 1002 6627
rect 343 6611 386 6621
rect 1027 6624 1051 6627
rect 1055 6624 1060 6627
rect 1463 6629 1467 6633
rect 1471 6629 1504 6633
rect 1508 6629 1534 6633
rect 1538 6629 1562 6633
rect 1566 6629 1599 6633
rect 1603 6629 1636 6633
rect 1640 6629 1666 6633
rect 1670 6629 1694 6633
rect 1698 6629 1731 6633
rect 1735 6629 1768 6633
rect 1772 6629 1798 6633
rect 1802 6629 1826 6633
rect 1830 6629 1863 6633
rect 1905 6630 1920 6633
rect 1924 6634 1931 6637
rect 1956 6634 1959 6640
rect 2433 6654 2455 6657
rect 2459 6654 2466 6657
rect 2491 6654 2515 6657
rect 2519 6654 2524 6657
rect 2538 6654 2545 6657
rect 2565 6654 2587 6657
rect 2591 6654 2598 6657
rect 2623 6654 2647 6657
rect 2651 6654 2656 6657
rect 2670 6654 2677 6657
rect 2697 6654 2719 6657
rect 2723 6654 2730 6657
rect 2755 6654 2779 6657
rect 2783 6654 2788 6657
rect 1959 6630 1978 6633
rect 1982 6634 1989 6637
rect 2422 6633 2425 6643
rect 2443 6633 2446 6643
rect 2459 6633 2462 6643
rect 2474 6636 2481 6640
rect 2485 6636 2490 6640
rect 2501 6633 2504 6643
rect 2517 6633 2520 6643
rect 2538 6633 2541 6643
rect 2554 6633 2557 6643
rect 2575 6633 2578 6643
rect 2591 6633 2594 6643
rect 2606 6636 2613 6640
rect 2617 6636 2622 6640
rect 2633 6633 2636 6643
rect 2649 6633 2652 6643
rect 2670 6633 2673 6643
rect 2686 6633 2689 6643
rect 2707 6633 2710 6643
rect 2723 6633 2726 6643
rect 2738 6636 2745 6640
rect 2749 6636 2754 6640
rect 2765 6633 2768 6643
rect 2781 6633 2784 6643
rect 2802 6633 2805 6643
rect 4403 6634 4829 6730
rect 1403 6622 1483 6626
rect 1487 6622 1550 6626
rect 1554 6622 1586 6626
rect 1590 6622 1615 6626
rect 1619 6622 1682 6626
rect 1686 6622 1718 6626
rect 1722 6622 1747 6626
rect 1751 6622 1814 6626
rect 1818 6622 1850 6626
rect 1854 6622 1863 6626
rect 1914 6624 1936 6627
rect 1940 6624 1947 6627
rect 1603 6616 1713 6619
rect 1972 6624 1996 6627
rect 2000 6624 2005 6627
rect 2408 6629 2412 6633
rect 2416 6629 2449 6633
rect 2453 6629 2479 6633
rect 2483 6629 2507 6633
rect 2511 6629 2544 6633
rect 2548 6629 2581 6633
rect 2585 6629 2611 6633
rect 2615 6629 2639 6633
rect 2643 6629 2676 6633
rect 2680 6629 2713 6633
rect 2717 6629 2743 6633
rect 2747 6629 2771 6633
rect 2775 6629 2808 6633
rect 2348 6622 2428 6626
rect 2432 6622 2495 6626
rect 2499 6622 2531 6626
rect 2535 6622 2560 6626
rect 2564 6622 2627 6626
rect 2631 6622 2663 6626
rect 2667 6622 2692 6626
rect 2696 6622 2759 6626
rect 2763 6622 2795 6626
rect 2799 6622 2808 6626
rect 4786 6624 4829 6634
rect 2548 6616 2658 6619
rect 4796 6614 4829 6624
rect 343 6601 376 6611
rect 958 6603 961 6613
rect 979 6603 982 6613
rect 995 6603 998 6613
rect 1010 6606 1017 6610
rect 1021 6606 1026 6610
rect 1037 6603 1040 6613
rect 1053 6603 1056 6613
rect 1074 6603 1077 6613
rect 1721 6608 1725 6612
rect 1729 6608 1733 6612
rect 343 6591 366 6601
rect 952 6599 985 6603
rect 989 6599 1015 6603
rect 1019 6599 1043 6603
rect 1047 6599 1081 6603
rect 1085 6599 1457 6603
rect 1472 6600 1702 6603
rect 1903 6603 1906 6613
rect 1924 6603 1927 6613
rect 1940 6603 1943 6613
rect 1955 6606 1962 6610
rect 1966 6606 1971 6610
rect 1982 6603 1985 6613
rect 1998 6603 2001 6613
rect 2019 6603 2022 6613
rect 2666 6608 2670 6612
rect 2674 6608 2678 6612
rect 4806 6604 4829 6614
rect 1897 6599 1930 6603
rect 1934 6599 1960 6603
rect 1964 6599 1988 6603
rect 1992 6599 2026 6603
rect 2030 6599 2402 6603
rect 2417 6600 2647 6603
rect 948 6592 964 6596
rect 968 6592 1031 6596
rect 1035 6592 1067 6596
rect 1071 6592 1397 6596
rect 1472 6593 1717 6596
rect 1893 6592 1909 6596
rect 1913 6592 1976 6596
rect 1980 6592 2012 6596
rect 2016 6592 2342 6596
rect 2417 6593 2662 6596
rect 4816 6594 4829 6604
rect 343 6581 356 6591
rect 851 6585 1709 6589
rect 1725 6585 1741 6589
rect 1745 6585 2654 6589
rect 2670 6585 2686 6589
rect 2690 6585 2822 6589
rect 343 6542 346 6581
rect 939 6579 943 6585
rect 1114 6578 1385 6582
rect 1119 6572 1433 6575
rect 1721 6572 1725 6576
rect 1729 6572 1733 6576
rect 1884 6579 1888 6585
rect 2057 6578 2330 6582
rect 2064 6572 2378 6575
rect 2666 6572 2670 6576
rect 2674 6572 2678 6576
rect 931 6563 939 6567
rect 1129 6565 1359 6568
rect 1363 6564 1421 6568
rect 1604 6565 1713 6568
rect 1876 6563 1884 6567
rect 2074 6565 2304 6568
rect 2308 6564 2366 6568
rect 2549 6565 2658 6568
rect 947 6557 955 6561
rect 959 6557 983 6561
rect 987 6557 995 6561
rect 999 6557 1000 6561
rect 1004 6557 1037 6561
rect 1041 6557 1056 6561
rect 1060 6557 1062 6561
rect 1066 6557 1073 6561
rect 1077 6557 1091 6561
rect 1095 6557 1107 6561
rect 1111 6557 1122 6561
rect 1126 6557 1133 6561
rect 1137 6557 1176 6561
rect 1180 6557 1216 6561
rect 1220 6557 1244 6561
rect 1248 6557 1256 6561
rect 1260 6557 1261 6561
rect 1265 6557 1298 6561
rect 1302 6557 1317 6561
rect 1321 6557 1323 6561
rect 1327 6557 1334 6561
rect 1338 6557 1352 6561
rect 1356 6557 1368 6561
rect 1372 6557 1457 6561
rect 1472 6558 1856 6561
rect 1892 6557 1900 6561
rect 1904 6557 1928 6561
rect 1932 6557 1940 6561
rect 1944 6557 1945 6561
rect 1949 6557 1982 6561
rect 1986 6557 2001 6561
rect 2005 6557 2007 6561
rect 2011 6557 2018 6561
rect 2022 6557 2036 6561
rect 2040 6557 2052 6561
rect 2056 6557 2067 6561
rect 2071 6557 2078 6561
rect 2082 6557 2121 6561
rect 2125 6557 2161 6561
rect 2165 6557 2189 6561
rect 2193 6557 2201 6561
rect 2205 6557 2206 6561
rect 2210 6557 2243 6561
rect 2247 6557 2262 6561
rect 2266 6557 2268 6561
rect 2272 6557 2279 6561
rect 2283 6557 2297 6561
rect 2301 6557 2313 6561
rect 2317 6557 2402 6561
rect 2417 6558 2801 6561
rect 948 6550 962 6554
rect 966 6550 1027 6554
rect 1031 6550 1049 6554
rect 1053 6550 1080 6554
rect 1084 6550 1124 6554
rect 1128 6550 1133 6554
rect 86 6539 346 6542
rect 967 6543 969 6547
rect 1013 6543 1014 6547
rect 1038 6543 1041 6547
rect 1170 6545 1173 6557
rect 1209 6550 1223 6554
rect 1227 6550 1288 6554
rect 1292 6550 1310 6554
rect 1314 6550 1341 6554
rect 1345 6550 1359 6554
rect 1415 6551 1485 6554
rect 1489 6551 1535 6555
rect 1539 6551 1586 6555
rect 1590 6551 1617 6555
rect 1621 6551 1667 6555
rect 1671 6551 1718 6555
rect 1722 6551 1749 6555
rect 1753 6551 1799 6555
rect 1803 6551 1850 6555
rect 1854 6551 1863 6555
rect 1893 6550 1907 6554
rect 1911 6550 1972 6554
rect 1976 6550 1994 6554
rect 1998 6550 2025 6554
rect 2029 6550 2069 6554
rect 2073 6550 2078 6554
rect 617 6536 618 6540
rect 622 6536 623 6540
rect 627 6536 628 6540
rect 632 6536 633 6540
rect 637 6536 638 6540
rect 642 6536 643 6540
rect 613 6535 647 6536
rect 617 6531 618 6535
rect 622 6531 623 6535
rect 627 6531 628 6535
rect 632 6531 633 6535
rect 637 6531 638 6535
rect 642 6531 643 6535
rect 613 6530 647 6531
rect 617 6526 618 6530
rect 622 6526 623 6530
rect 627 6526 628 6530
rect 632 6526 633 6530
rect 637 6526 638 6530
rect 642 6526 643 6530
rect 613 6525 647 6526
rect 617 6521 618 6525
rect 622 6521 623 6525
rect 627 6521 628 6525
rect 632 6521 633 6525
rect 637 6521 638 6525
rect 642 6521 643 6525
rect 663 6536 664 6540
rect 668 6536 669 6540
rect 673 6536 674 6540
rect 678 6536 679 6540
rect 683 6536 684 6540
rect 688 6536 689 6540
rect 659 6535 693 6536
rect 663 6531 664 6535
rect 668 6531 669 6535
rect 673 6531 674 6535
rect 678 6531 679 6535
rect 683 6531 684 6535
rect 688 6531 689 6535
rect 659 6530 693 6531
rect 663 6526 664 6530
rect 668 6526 669 6530
rect 673 6526 674 6530
rect 678 6526 679 6530
rect 683 6526 684 6530
rect 688 6526 689 6530
rect 948 6527 951 6532
rect 966 6528 969 6532
rect 659 6525 693 6526
rect 663 6521 664 6525
rect 668 6521 669 6525
rect 673 6521 674 6525
rect 678 6521 679 6525
rect 683 6521 684 6525
rect 688 6521 689 6525
rect 966 6524 967 6528
rect 991 6527 994 6532
rect 1012 6528 1015 6532
rect 1022 6528 1025 6532
rect 948 6518 951 6523
rect 966 6518 969 6524
rect 986 6523 989 6526
rect 993 6523 994 6527
rect 1006 6524 1015 6528
rect 991 6518 994 6523
rect 1012 6518 1015 6524
rect 1022 6518 1025 6524
rect 1038 6529 1041 6532
rect 1038 6525 1040 6529
rect 1066 6527 1069 6532
rect 1082 6528 1085 6532
rect 1038 6518 1041 6525
rect 1058 6525 1069 6527
rect 1058 6523 1059 6525
rect 1063 6523 1069 6525
rect 1077 6524 1079 6528
rect 1083 6524 1085 6528
rect 1066 6518 1069 6523
rect 1082 6518 1085 6524
rect 1091 6526 1094 6532
rect 1098 6526 1101 6532
rect 1122 6526 1125 6540
rect 1228 6543 1230 6547
rect 1274 6543 1275 6547
rect 1299 6543 1302 6547
rect 1451 6544 1504 6548
rect 1508 6544 1534 6548
rect 1538 6544 1562 6548
rect 1566 6544 1636 6548
rect 1640 6544 1666 6548
rect 1670 6544 1694 6548
rect 1698 6544 1768 6548
rect 1772 6544 1798 6548
rect 1802 6544 1826 6548
rect 1830 6544 1863 6548
rect 1154 6534 1157 6537
rect 1149 6531 1157 6534
rect 1091 6523 1125 6526
rect 1154 6525 1157 6531
rect 1172 6530 1174 6533
rect 1178 6529 1183 6534
rect 1209 6527 1212 6532
rect 1227 6528 1230 6532
rect 1091 6518 1094 6523
rect 1098 6518 1101 6523
rect 1107 6518 1110 6523
rect 1227 6524 1228 6528
rect 1252 6527 1255 6532
rect 1273 6528 1276 6532
rect 1283 6528 1286 6532
rect 976 6505 977 6509
rect 1023 6506 1024 6510
rect 1048 6505 1049 6509
rect 1134 6502 1137 6514
rect 948 6498 977 6502
rect 981 6498 1008 6502
rect 1012 6498 1033 6502
rect 1037 6498 1092 6502
rect 1096 6498 1114 6502
rect 1118 6498 1137 6502
rect 577 6495 645 6496
rect 1170 6495 1173 6521
rect 1209 6518 1212 6523
rect 1227 6518 1230 6524
rect 1247 6523 1250 6526
rect 1254 6523 1255 6527
rect 1267 6524 1276 6528
rect 1252 6518 1255 6523
rect 1273 6518 1276 6524
rect 1283 6518 1286 6524
rect 1299 6529 1302 6532
rect 1299 6525 1301 6529
rect 1327 6527 1330 6532
rect 1343 6528 1346 6532
rect 1299 6518 1302 6525
rect 1319 6525 1330 6527
rect 1319 6523 1320 6525
rect 1324 6523 1330 6525
rect 1338 6524 1340 6528
rect 1344 6524 1346 6528
rect 1327 6518 1330 6523
rect 1343 6518 1346 6524
rect 1352 6526 1355 6532
rect 1477 6532 1480 6544
rect 1498 6532 1501 6544
rect 1514 6532 1517 6544
rect 1533 6538 1545 6541
rect 1556 6532 1559 6544
rect 1572 6532 1575 6544
rect 1593 6532 1596 6544
rect 1609 6532 1612 6544
rect 1630 6532 1633 6544
rect 1646 6532 1649 6544
rect 1665 6538 1677 6541
rect 1688 6532 1691 6544
rect 1704 6532 1707 6544
rect 1725 6532 1728 6544
rect 1741 6532 1744 6544
rect 1762 6532 1765 6544
rect 1778 6532 1781 6544
rect 1797 6538 1809 6541
rect 1820 6532 1823 6544
rect 1836 6532 1839 6544
rect 1857 6532 1860 6544
rect 1912 6543 1914 6547
rect 1958 6543 1959 6547
rect 1983 6543 1986 6547
rect 2115 6545 2118 6557
rect 4826 6555 4829 6594
rect 5083 6555 5086 6809
rect 2154 6550 2168 6554
rect 2172 6550 2233 6554
rect 2237 6550 2255 6554
rect 2259 6550 2286 6554
rect 2290 6550 2304 6554
rect 2360 6551 2430 6554
rect 2434 6551 2480 6555
rect 2484 6551 2531 6555
rect 2535 6551 2562 6555
rect 2566 6551 2612 6555
rect 2616 6551 2663 6555
rect 2667 6551 2694 6555
rect 2698 6551 2744 6555
rect 2748 6551 2795 6555
rect 2799 6551 2808 6555
rect 4483 6549 4484 6553
rect 4488 6549 4489 6553
rect 4493 6549 4494 6553
rect 4498 6549 4499 6553
rect 4503 6549 4504 6553
rect 4508 6549 4509 6553
rect 4479 6548 4513 6549
rect 1359 6526 1362 6532
rect 1352 6523 1362 6526
rect 1370 6523 1372 6526
rect 1352 6518 1355 6523
rect 1359 6518 1362 6523
rect 1477 6518 1494 6521
rect 1498 6522 1505 6525
rect 1530 6522 1533 6528
rect 1533 6518 1552 6521
rect 1556 6522 1563 6525
rect 1611 6518 1626 6521
rect 1630 6522 1637 6525
rect 1662 6522 1665 6528
rect 1665 6518 1684 6521
rect 1688 6522 1695 6525
rect 1743 6518 1758 6521
rect 1762 6522 1769 6525
rect 1794 6522 1797 6528
rect 1797 6518 1816 6521
rect 1820 6522 1827 6525
rect 1893 6527 1896 6532
rect 1911 6528 1914 6532
rect 1911 6524 1912 6528
rect 1936 6527 1939 6532
rect 1957 6528 1960 6532
rect 1967 6528 1970 6532
rect 1893 6518 1896 6523
rect 1911 6518 1914 6524
rect 1931 6523 1934 6526
rect 1938 6523 1939 6527
rect 1951 6524 1960 6528
rect 1936 6518 1939 6523
rect 1957 6518 1960 6524
rect 1967 6518 1970 6524
rect 1237 6505 1238 6509
rect 1284 6506 1285 6510
rect 1309 6505 1310 6509
rect 1488 6512 1510 6515
rect 1514 6512 1521 6515
rect 1209 6498 1238 6502
rect 1242 6498 1269 6502
rect 1273 6498 1294 6502
rect 1298 6498 1344 6502
rect 1348 6498 1353 6502
rect 1357 6498 1433 6502
rect 1546 6512 1570 6515
rect 1574 6512 1579 6515
rect 1593 6512 1600 6515
rect 1620 6512 1642 6515
rect 1646 6512 1653 6515
rect 1678 6512 1702 6515
rect 1706 6512 1711 6515
rect 1725 6512 1732 6515
rect 1752 6512 1774 6515
rect 1778 6512 1785 6515
rect 1810 6512 1834 6515
rect 1838 6512 1843 6515
rect 1983 6529 1986 6532
rect 1983 6525 1985 6529
rect 2011 6527 2014 6532
rect 2027 6528 2030 6532
rect 1983 6518 1986 6525
rect 2003 6525 2014 6527
rect 2003 6523 2004 6525
rect 2008 6523 2014 6525
rect 2022 6524 2024 6528
rect 2028 6524 2030 6528
rect 2011 6518 2014 6523
rect 2027 6518 2030 6524
rect 2036 6526 2039 6532
rect 2043 6526 2046 6532
rect 2067 6526 2070 6540
rect 2173 6543 2175 6547
rect 2219 6543 2220 6547
rect 2244 6543 2247 6547
rect 2396 6544 2449 6548
rect 2453 6544 2479 6548
rect 2483 6544 2507 6548
rect 2511 6544 2581 6548
rect 2585 6544 2611 6548
rect 2615 6544 2639 6548
rect 2643 6544 2713 6548
rect 2717 6544 2743 6548
rect 2747 6544 2771 6548
rect 2775 6544 2808 6548
rect 4483 6544 4484 6548
rect 4488 6544 4489 6548
rect 4493 6544 4494 6548
rect 4498 6544 4499 6548
rect 4503 6544 4504 6548
rect 4508 6544 4509 6548
rect 2099 6534 2102 6537
rect 2094 6531 2102 6534
rect 2036 6523 2070 6526
rect 2099 6525 2102 6531
rect 2117 6530 2119 6533
rect 2123 6529 2128 6534
rect 2154 6527 2157 6532
rect 2172 6528 2175 6532
rect 2036 6518 2039 6523
rect 2043 6518 2046 6523
rect 2052 6518 2055 6523
rect 2172 6524 2173 6528
rect 2197 6527 2200 6532
rect 2218 6528 2221 6532
rect 2228 6528 2231 6532
rect 1921 6505 1922 6509
rect 1968 6506 1969 6510
rect 1993 6505 1994 6509
rect 2079 6502 2082 6514
rect 577 6491 579 6495
rect 583 6491 584 6495
rect 588 6491 589 6495
rect 593 6491 594 6495
rect 598 6491 599 6495
rect 603 6491 604 6495
rect 608 6491 609 6495
rect 613 6491 614 6495
rect 618 6491 619 6495
rect 623 6491 624 6495
rect 628 6491 629 6495
rect 633 6491 634 6495
rect 638 6491 639 6495
rect 643 6491 645 6495
rect 947 6491 956 6495
rect 960 6491 984 6495
rect 988 6491 999 6495
rect 1003 6491 1033 6495
rect 1037 6491 1056 6495
rect 1060 6491 1065 6495
rect 1069 6491 1074 6495
rect 1078 6491 1092 6495
rect 1096 6491 1176 6495
rect 1180 6491 1200 6495
rect 1204 6491 1217 6495
rect 1221 6491 1245 6495
rect 1249 6491 1260 6495
rect 1264 6491 1294 6495
rect 1298 6491 1317 6495
rect 1321 6491 1326 6495
rect 1330 6491 1335 6495
rect 1339 6491 1353 6495
rect 1357 6491 1361 6495
rect 1365 6491 1367 6495
rect 1371 6491 1445 6495
rect 1477 6491 1480 6501
rect 1498 6491 1501 6501
rect 1514 6491 1517 6501
rect 1529 6494 1536 6498
rect 1540 6494 1545 6498
rect 1556 6491 1559 6501
rect 1572 6491 1575 6501
rect 1593 6491 1596 6501
rect 1609 6491 1612 6501
rect 1630 6491 1633 6501
rect 1646 6491 1649 6501
rect 1661 6494 1668 6498
rect 1672 6494 1677 6498
rect 1688 6491 1691 6501
rect 1704 6491 1707 6501
rect 1725 6491 1728 6501
rect 1741 6491 1744 6501
rect 1762 6491 1765 6501
rect 1778 6491 1781 6501
rect 1793 6494 1800 6498
rect 1804 6494 1809 6498
rect 1820 6491 1823 6501
rect 1836 6491 1839 6501
rect 1857 6491 1860 6501
rect 1893 6498 1922 6502
rect 1926 6498 1953 6502
rect 1957 6498 1978 6502
rect 1982 6498 2037 6502
rect 2041 6498 2059 6502
rect 2063 6498 2082 6502
rect 2115 6495 2118 6521
rect 2154 6518 2157 6523
rect 2172 6518 2175 6524
rect 2192 6523 2195 6526
rect 2199 6523 2200 6527
rect 2212 6524 2221 6528
rect 2197 6518 2200 6523
rect 2218 6518 2221 6524
rect 2228 6518 2231 6524
rect 2244 6529 2247 6532
rect 2244 6525 2246 6529
rect 2272 6527 2275 6532
rect 2288 6528 2291 6532
rect 2244 6518 2247 6525
rect 2264 6525 2275 6527
rect 2264 6523 2265 6525
rect 2269 6523 2275 6525
rect 2283 6524 2285 6528
rect 2289 6524 2291 6528
rect 2272 6518 2275 6523
rect 2288 6518 2291 6524
rect 2297 6526 2300 6532
rect 2422 6532 2425 6544
rect 2443 6532 2446 6544
rect 2459 6532 2462 6544
rect 2478 6538 2490 6541
rect 2501 6532 2504 6544
rect 2517 6532 2520 6544
rect 2538 6532 2541 6544
rect 2554 6532 2557 6544
rect 2575 6532 2578 6544
rect 2591 6532 2594 6544
rect 2610 6538 2622 6541
rect 2633 6532 2636 6544
rect 2649 6532 2652 6544
rect 2670 6532 2673 6544
rect 2686 6532 2689 6544
rect 2707 6532 2710 6544
rect 2723 6532 2726 6544
rect 2742 6538 2754 6541
rect 2765 6532 2768 6544
rect 2781 6532 2784 6544
rect 2802 6532 2805 6544
rect 4479 6543 4513 6544
rect 4483 6539 4484 6543
rect 4488 6539 4489 6543
rect 4493 6539 4494 6543
rect 4498 6539 4499 6543
rect 4503 6539 4504 6543
rect 4508 6539 4509 6543
rect 4479 6538 4513 6539
rect 4483 6534 4484 6538
rect 4488 6534 4489 6538
rect 4493 6534 4494 6538
rect 4498 6534 4499 6538
rect 4503 6534 4504 6538
rect 4508 6534 4509 6538
rect 4529 6549 4530 6553
rect 4534 6549 4535 6553
rect 4539 6549 4540 6553
rect 4544 6549 4545 6553
rect 4549 6549 4550 6553
rect 4554 6549 4555 6553
rect 4826 6552 5086 6555
rect 4525 6548 4559 6549
rect 4529 6544 4530 6548
rect 4534 6544 4535 6548
rect 4539 6544 4540 6548
rect 4544 6544 4545 6548
rect 4549 6544 4550 6548
rect 4554 6544 4555 6548
rect 4525 6543 4559 6544
rect 4529 6539 4530 6543
rect 4534 6539 4535 6543
rect 4539 6539 4540 6543
rect 4544 6539 4545 6543
rect 4549 6539 4550 6543
rect 4554 6539 4555 6543
rect 4525 6538 4559 6539
rect 4529 6534 4530 6538
rect 4534 6534 4535 6538
rect 4539 6534 4540 6538
rect 4544 6534 4545 6538
rect 4549 6534 4550 6538
rect 4554 6534 4555 6538
rect 2304 6526 2307 6532
rect 2297 6523 2307 6526
rect 2315 6523 2317 6526
rect 2297 6518 2300 6523
rect 2304 6518 2307 6523
rect 2422 6518 2439 6521
rect 2443 6522 2450 6525
rect 2475 6522 2478 6528
rect 2478 6518 2497 6521
rect 2501 6522 2508 6525
rect 2556 6518 2571 6521
rect 2575 6522 2582 6525
rect 2607 6522 2610 6528
rect 2610 6518 2629 6521
rect 2633 6522 2640 6525
rect 2688 6518 2703 6521
rect 2707 6522 2714 6525
rect 2739 6522 2742 6528
rect 2742 6518 2761 6521
rect 2765 6522 2772 6525
rect 2182 6505 2183 6509
rect 2229 6506 2230 6510
rect 2254 6505 2255 6509
rect 2433 6512 2455 6515
rect 2459 6512 2466 6515
rect 2154 6498 2183 6502
rect 2187 6498 2214 6502
rect 2218 6498 2239 6502
rect 2243 6498 2289 6502
rect 2293 6498 2298 6502
rect 2302 6498 2378 6502
rect 2491 6512 2515 6515
rect 2519 6512 2524 6515
rect 2538 6512 2545 6515
rect 2565 6512 2587 6515
rect 2591 6512 2598 6515
rect 2623 6512 2647 6515
rect 2651 6512 2656 6515
rect 2670 6512 2677 6515
rect 2697 6512 2719 6515
rect 2723 6512 2730 6515
rect 2755 6512 2779 6515
rect 2783 6512 2788 6515
rect 1892 6491 1901 6495
rect 1905 6491 1929 6495
rect 1933 6491 1944 6495
rect 1948 6491 1978 6495
rect 1982 6491 2001 6495
rect 2005 6491 2010 6495
rect 2014 6491 2019 6495
rect 2023 6491 2037 6495
rect 2041 6491 2121 6495
rect 2125 6491 2145 6495
rect 2149 6491 2162 6495
rect 2166 6491 2190 6495
rect 2194 6491 2205 6495
rect 2209 6491 2239 6495
rect 2243 6491 2262 6495
rect 2266 6491 2271 6495
rect 2275 6491 2280 6495
rect 2284 6491 2298 6495
rect 2302 6491 2306 6495
rect 2310 6491 2312 6495
rect 2316 6491 2390 6495
rect 2422 6491 2425 6501
rect 2443 6491 2446 6501
rect 2459 6491 2462 6501
rect 2474 6494 2481 6498
rect 2485 6494 2490 6498
rect 2501 6491 2504 6501
rect 2517 6491 2520 6501
rect 2538 6491 2541 6501
rect 2554 6491 2557 6501
rect 2575 6491 2578 6501
rect 2591 6491 2594 6501
rect 2606 6494 2613 6498
rect 2617 6494 2622 6498
rect 2633 6491 2636 6501
rect 2649 6491 2652 6501
rect 2670 6491 2673 6501
rect 2686 6491 2689 6501
rect 2707 6491 2710 6501
rect 2723 6491 2726 6501
rect 2738 6494 2745 6498
rect 2749 6494 2754 6498
rect 2765 6491 2768 6501
rect 2781 6491 2784 6501
rect 2802 6491 2805 6501
rect 4826 6500 5086 6503
rect 577 6490 645 6491
rect 86 6487 346 6490
rect 86 6233 89 6487
rect 343 6448 346 6487
rect 577 6486 579 6490
rect 583 6486 584 6490
rect 588 6486 589 6490
rect 593 6486 594 6490
rect 598 6486 599 6490
rect 603 6486 604 6490
rect 608 6486 609 6490
rect 613 6486 614 6490
rect 618 6486 619 6490
rect 623 6486 624 6490
rect 628 6486 629 6490
rect 633 6486 634 6490
rect 638 6486 639 6490
rect 643 6486 645 6490
rect 577 6484 645 6486
rect 418 6460 645 6484
rect 1140 6467 1143 6491
rect 418 6457 427 6460
rect 439 6457 443 6460
rect 459 6457 468 6460
rect 480 6457 484 6460
rect 502 6457 511 6460
rect 523 6457 527 6460
rect 343 6438 356 6448
rect 343 6428 366 6438
rect 343 6418 376 6428
rect 343 6408 386 6418
rect 343 6362 398 6408
rect 422 6369 423 6457
rect 435 6369 447 6375
rect 463 6369 464 6457
rect 476 6369 488 6375
rect 506 6369 507 6457
rect 519 6369 531 6375
rect 546 6428 645 6460
rect 1170 6463 1173 6491
rect 1209 6484 1238 6488
rect 1242 6484 1269 6488
rect 1273 6484 1294 6488
rect 1298 6484 1344 6488
rect 1348 6484 1353 6488
rect 1357 6484 1378 6488
rect 1463 6487 1467 6491
rect 1471 6487 1504 6491
rect 1508 6487 1534 6491
rect 1538 6487 1562 6491
rect 1566 6487 1599 6491
rect 1603 6487 1636 6491
rect 1640 6487 1666 6491
rect 1670 6487 1694 6491
rect 1698 6487 1731 6491
rect 1735 6487 1768 6491
rect 1772 6487 1798 6491
rect 1802 6487 1826 6491
rect 1830 6487 1863 6491
rect 1237 6477 1238 6481
rect 1284 6476 1285 6480
rect 1309 6477 1310 6481
rect 1403 6480 1483 6484
rect 1487 6480 1550 6484
rect 1554 6480 1586 6484
rect 1590 6480 1615 6484
rect 1619 6480 1682 6484
rect 1686 6480 1718 6484
rect 1722 6480 1747 6484
rect 1751 6480 1814 6484
rect 1818 6480 1850 6484
rect 1854 6480 1863 6484
rect 1177 6464 1182 6469
rect 1131 6458 1134 6463
rect 1209 6463 1212 6468
rect 1126 6455 1134 6458
rect 1121 6450 1126 6455
rect 1131 6441 1134 6455
rect 1142 6455 1145 6458
rect 1154 6453 1157 6459
rect 1177 6454 1180 6460
rect 1227 6462 1230 6468
rect 1252 6463 1255 6468
rect 1149 6450 1157 6453
rect 1169 6451 1180 6454
rect 1209 6454 1212 6459
rect 1227 6458 1228 6462
rect 1247 6460 1250 6463
rect 1254 6459 1255 6463
rect 1273 6462 1276 6468
rect 1283 6462 1286 6468
rect 1227 6454 1230 6458
rect 1252 6454 1255 6459
rect 1267 6458 1276 6462
rect 1273 6454 1276 6458
rect 1283 6454 1286 6458
rect 1154 6447 1157 6450
rect 1299 6461 1302 6468
rect 1299 6457 1301 6461
rect 1319 6461 1320 6463
rect 1327 6463 1330 6468
rect 1324 6461 1330 6463
rect 1343 6462 1346 6468
rect 1319 6459 1330 6461
rect 1299 6454 1302 6457
rect 1327 6454 1330 6459
rect 1338 6458 1340 6462
rect 1344 6458 1346 6462
rect 1343 6454 1346 6458
rect 1352 6463 1355 6468
rect 1359 6463 1362 6468
rect 2085 6467 2088 6491
rect 2115 6463 2118 6491
rect 2154 6484 2183 6488
rect 2187 6484 2214 6488
rect 2218 6484 2239 6488
rect 2243 6484 2289 6488
rect 2293 6484 2298 6488
rect 2302 6484 2323 6488
rect 2408 6487 2412 6491
rect 2416 6487 2449 6491
rect 2453 6487 2479 6491
rect 2483 6487 2507 6491
rect 2511 6487 2544 6491
rect 2548 6487 2581 6491
rect 2585 6487 2611 6491
rect 2615 6487 2639 6491
rect 2643 6487 2676 6491
rect 2680 6487 2713 6491
rect 2717 6487 2743 6491
rect 2747 6487 2771 6491
rect 2775 6487 2808 6491
rect 2182 6477 2183 6481
rect 2229 6476 2230 6480
rect 2254 6477 2255 6481
rect 2348 6480 2428 6484
rect 2432 6480 2495 6484
rect 2499 6480 2531 6484
rect 2535 6480 2560 6484
rect 2564 6480 2627 6484
rect 2631 6480 2663 6484
rect 2667 6480 2692 6484
rect 2696 6480 2759 6484
rect 2763 6480 2795 6484
rect 2799 6480 2808 6484
rect 2122 6464 2127 6469
rect 1352 6460 1362 6463
rect 1352 6454 1355 6460
rect 1359 6454 1362 6460
rect 1370 6460 1373 6463
rect 2076 6458 2079 6463
rect 2154 6463 2157 6468
rect 2071 6455 2079 6458
rect 2066 6450 2071 6455
rect 1228 6439 1230 6443
rect 1274 6439 1275 6443
rect 1299 6439 1302 6443
rect 2076 6441 2079 6455
rect 2087 6455 2090 6458
rect 2099 6453 2102 6459
rect 2122 6454 2125 6460
rect 2172 6462 2175 6468
rect 2197 6463 2200 6468
rect 2094 6450 2102 6453
rect 2114 6451 2125 6454
rect 2154 6454 2157 6459
rect 2172 6458 2173 6462
rect 2192 6460 2195 6463
rect 2199 6459 2200 6463
rect 2218 6462 2221 6468
rect 2228 6462 2231 6468
rect 2172 6454 2175 6458
rect 2197 6454 2200 6459
rect 2212 6458 2221 6462
rect 2218 6454 2221 6458
rect 2228 6454 2231 6458
rect 2099 6447 2102 6450
rect 1140 6429 1143 6433
rect 1170 6429 1173 6439
rect 1209 6432 1223 6436
rect 1227 6432 1288 6436
rect 1292 6432 1310 6436
rect 1314 6432 1341 6436
rect 1345 6432 1421 6436
rect 2244 6461 2247 6468
rect 2244 6457 2246 6461
rect 2264 6461 2265 6463
rect 2272 6463 2275 6468
rect 2269 6461 2275 6463
rect 2288 6462 2291 6468
rect 2264 6459 2275 6461
rect 2244 6454 2247 6457
rect 2272 6454 2275 6459
rect 2283 6458 2285 6462
rect 2289 6458 2291 6462
rect 2288 6454 2291 6458
rect 2297 6463 2300 6468
rect 2304 6463 2307 6468
rect 2297 6460 2307 6463
rect 2297 6454 2300 6460
rect 2304 6454 2307 6460
rect 2315 6460 2318 6463
rect 4826 6461 4829 6500
rect 4816 6451 4829 6461
rect 2173 6439 2175 6443
rect 2219 6439 2220 6443
rect 2244 6439 2247 6443
rect 4806 6441 4829 6451
rect 2085 6429 2088 6433
rect 2115 6429 2118 6439
rect 2154 6432 2168 6436
rect 2172 6432 2233 6436
rect 2237 6432 2255 6436
rect 2259 6432 2286 6436
rect 2290 6432 2366 6436
rect 4796 6431 4829 6441
rect 546 6425 550 6428
rect 562 6425 566 6428
rect 578 6425 582 6428
rect 594 6425 598 6428
rect 951 6425 1005 6429
rect 1009 6425 1095 6429
rect 1099 6425 1122 6429
rect 1126 6425 1176 6429
rect 1180 6425 1200 6429
rect 1204 6425 1216 6429
rect 1220 6425 1244 6429
rect 1248 6425 1256 6429
rect 1260 6425 1261 6429
rect 1265 6425 1298 6429
rect 1302 6425 1317 6429
rect 1321 6425 1323 6429
rect 1327 6425 1334 6429
rect 1338 6425 1352 6429
rect 1356 6425 1368 6429
rect 1372 6425 1457 6429
rect 1896 6425 1950 6429
rect 1954 6425 2040 6429
rect 2044 6425 2067 6429
rect 2071 6425 2121 6429
rect 2125 6425 2145 6429
rect 2149 6425 2161 6429
rect 2165 6425 2189 6429
rect 2193 6425 2201 6429
rect 2205 6425 2206 6429
rect 2210 6425 2243 6429
rect 2247 6425 2262 6429
rect 2266 6425 2268 6429
rect 2272 6425 2279 6429
rect 2283 6425 2297 6429
rect 2301 6425 2313 6429
rect 2317 6425 2402 6429
rect 545 6369 546 6425
rect 999 6409 1002 6425
rect 1089 6409 1092 6425
rect 1170 6409 1173 6425
rect 1209 6418 1223 6422
rect 1227 6418 1288 6422
rect 1292 6418 1310 6422
rect 1314 6418 1341 6422
rect 1345 6418 1421 6422
rect 1228 6411 1230 6415
rect 1274 6411 1275 6415
rect 1299 6411 1302 6415
rect 1944 6409 1947 6425
rect 2034 6409 2037 6425
rect 2115 6409 2118 6425
rect 2154 6418 2168 6422
rect 2172 6418 2233 6422
rect 2237 6418 2255 6422
rect 2259 6418 2286 6422
rect 2290 6418 2366 6422
rect 4786 6421 4829 6431
rect 983 6398 986 6401
rect 1073 6398 1076 6401
rect 1154 6398 1157 6401
rect 978 6395 986 6398
rect 983 6389 986 6395
rect 1001 6394 1009 6397
rect 1068 6395 1076 6398
rect 1073 6389 1076 6395
rect 1091 6394 1093 6397
rect 1097 6393 1102 6398
rect 1149 6395 1157 6398
rect 1154 6389 1157 6395
rect 1172 6394 1173 6397
rect 1177 6393 1182 6398
rect 1209 6395 1212 6400
rect 1227 6396 1230 6400
rect 1227 6392 1228 6396
rect 1252 6395 1255 6400
rect 1273 6396 1276 6400
rect 1283 6396 1286 6400
rect 431 6362 451 6369
rect 343 6348 451 6362
rect 472 6348 481 6369
rect 515 6362 524 6369
rect 554 6365 558 6369
rect 570 6365 574 6369
rect 554 6364 574 6365
rect 489 6349 490 6362
rect 494 6360 524 6362
rect 494 6351 505 6360
rect 513 6351 524 6360
rect 532 6351 533 6364
rect 537 6358 574 6364
rect 537 6351 567 6358
rect 586 6355 590 6369
rect 494 6349 524 6351
rect 343 6344 481 6348
rect 515 6346 524 6349
rect 554 6346 567 6351
rect 579 6351 590 6355
rect 600 6351 803 6364
rect 999 6363 1002 6385
rect 1089 6363 1092 6385
rect 1170 6363 1173 6385
rect 1209 6386 1212 6391
rect 1227 6386 1230 6392
rect 1247 6391 1250 6394
rect 1254 6391 1255 6395
rect 1267 6392 1276 6396
rect 1252 6386 1255 6391
rect 1273 6386 1276 6392
rect 1283 6386 1286 6392
rect 1299 6397 1302 6400
rect 1299 6393 1301 6397
rect 1327 6395 1330 6400
rect 1343 6396 1346 6400
rect 1299 6386 1302 6393
rect 1319 6393 1330 6395
rect 1319 6391 1320 6393
rect 1324 6391 1330 6393
rect 1338 6392 1340 6396
rect 1344 6392 1346 6396
rect 1327 6386 1330 6391
rect 1343 6386 1346 6392
rect 1352 6394 1355 6400
rect 2173 6411 2175 6415
rect 2219 6411 2220 6415
rect 2244 6411 2247 6415
rect 1359 6394 1362 6400
rect 1928 6398 1931 6401
rect 2018 6398 2021 6401
rect 2099 6398 2102 6401
rect 1352 6391 1362 6394
rect 1923 6395 1931 6398
rect 1370 6391 1372 6394
rect 1352 6386 1355 6391
rect 1359 6386 1362 6391
rect 1928 6389 1931 6395
rect 1946 6394 1954 6397
rect 2013 6395 2021 6398
rect 2018 6389 2021 6395
rect 2036 6394 2038 6397
rect 2042 6393 2047 6398
rect 2094 6395 2102 6398
rect 2099 6389 2102 6395
rect 2117 6394 2118 6397
rect 2122 6393 2127 6398
rect 2154 6395 2157 6400
rect 2172 6396 2175 6400
rect 2172 6392 2173 6396
rect 2197 6395 2200 6400
rect 2218 6396 2221 6400
rect 2228 6396 2231 6400
rect 1237 6373 1238 6377
rect 1284 6374 1285 6378
rect 1309 6373 1310 6377
rect 1209 6366 1238 6370
rect 1242 6366 1269 6370
rect 1273 6366 1294 6370
rect 1298 6366 1353 6370
rect 1357 6366 1433 6370
rect 1944 6363 1947 6385
rect 2034 6363 2037 6385
rect 2115 6363 2118 6385
rect 2154 6386 2157 6391
rect 2172 6386 2175 6392
rect 2192 6391 2195 6394
rect 2199 6391 2200 6395
rect 2212 6392 2221 6396
rect 2197 6386 2200 6391
rect 2218 6386 2221 6392
rect 2228 6386 2231 6392
rect 2244 6397 2247 6400
rect 2244 6393 2246 6397
rect 2272 6395 2275 6400
rect 2288 6396 2291 6400
rect 2244 6386 2247 6393
rect 2264 6393 2275 6395
rect 2264 6391 2265 6393
rect 2269 6391 2275 6393
rect 2283 6392 2285 6396
rect 2289 6392 2291 6396
rect 2272 6386 2275 6391
rect 2288 6386 2291 6392
rect 2297 6394 2300 6400
rect 2304 6394 2307 6400
rect 2297 6391 2307 6394
rect 2315 6391 2317 6394
rect 2297 6386 2300 6391
rect 2304 6386 2307 6391
rect 2182 6373 2183 6377
rect 2229 6374 2230 6378
rect 2254 6373 2255 6377
rect 2154 6366 2183 6370
rect 2187 6366 2214 6370
rect 2218 6366 2239 6370
rect 2243 6366 2298 6370
rect 2302 6366 2378 6370
rect 955 6359 1005 6363
rect 1009 6359 1041 6363
rect 1045 6359 1095 6363
rect 1099 6359 1119 6363
rect 1126 6359 1176 6363
rect 1180 6359 1200 6363
rect 1204 6359 1217 6363
rect 1221 6359 1245 6363
rect 1249 6359 1260 6363
rect 1264 6359 1294 6363
rect 1298 6359 1317 6363
rect 1321 6359 1326 6363
rect 1330 6359 1335 6363
rect 1339 6359 1353 6363
rect 1357 6359 1361 6363
rect 1365 6359 1367 6363
rect 1371 6359 1445 6363
rect 1900 6359 1950 6363
rect 1954 6359 1986 6363
rect 1990 6359 2040 6363
rect 2044 6359 2064 6363
rect 2071 6359 2121 6363
rect 2125 6359 2145 6363
rect 2149 6359 2162 6363
rect 2166 6359 2190 6363
rect 2194 6359 2205 6363
rect 2209 6359 2239 6363
rect 2243 6359 2262 6363
rect 2266 6359 2271 6363
rect 2275 6359 2280 6363
rect 2284 6359 2298 6363
rect 2302 6359 2306 6363
rect 2310 6359 2312 6363
rect 2316 6359 2390 6363
rect 343 6312 398 6344
rect 431 6342 492 6344
rect 431 6339 451 6342
rect 472 6340 492 6342
rect 472 6339 476 6340
rect 343 6302 386 6312
rect 343 6292 376 6302
rect 343 6282 366 6292
rect 343 6272 356 6282
rect 422 6280 423 6339
rect 463 6280 464 6339
rect 488 6339 492 6340
rect 515 6342 535 6346
rect 515 6339 519 6342
rect 531 6339 535 6342
rect 554 6342 574 6346
rect 554 6339 558 6342
rect 570 6339 574 6342
rect 586 6339 590 6351
rect 506 6280 507 6339
rect 545 6299 546 6339
rect 969 6335 972 6359
rect 999 6331 1002 6359
rect 960 6326 963 6331
rect 1023 6327 1026 6359
rect 1059 6335 1062 6359
rect 943 6323 963 6326
rect 960 6309 963 6323
rect 971 6323 974 6326
rect 983 6321 986 6327
rect 978 6318 986 6321
rect 998 6320 1006 6322
rect 998 6319 1010 6320
rect 1089 6331 1092 6359
rect 1096 6332 1101 6337
rect 1050 6326 1053 6331
rect 1014 6318 1017 6323
rect 1044 6323 1053 6326
rect 983 6315 986 6318
rect 1025 6315 1028 6318
rect 546 6290 550 6299
rect 562 6290 566 6299
rect 578 6290 582 6299
rect 594 6290 598 6299
rect 969 6297 972 6301
rect 999 6297 1002 6307
rect 1014 6309 1017 6314
rect 1050 6309 1053 6323
rect 1061 6323 1064 6326
rect 1073 6321 1076 6327
rect 1096 6322 1099 6328
rect 1113 6327 1116 6359
rect 1140 6335 1143 6359
rect 1170 6331 1173 6359
rect 1209 6352 1238 6356
rect 1242 6352 1269 6356
rect 1273 6352 1294 6356
rect 1298 6352 1353 6356
rect 1357 6352 1433 6356
rect 1237 6345 1238 6349
rect 1284 6344 1285 6348
rect 1309 6345 1310 6349
rect 1177 6332 1182 6337
rect 1068 6318 1076 6321
rect 1088 6319 1099 6322
rect 1122 6326 1126 6330
rect 1131 6326 1134 6331
rect 1209 6331 1212 6336
rect 1104 6318 1107 6323
rect 1126 6323 1134 6326
rect 1073 6315 1076 6318
rect 1115 6315 1118 6318
rect 1122 6315 1123 6318
rect 1023 6297 1026 6301
rect 1059 6297 1062 6301
rect 1089 6297 1092 6307
rect 1104 6309 1107 6314
rect 1131 6309 1134 6323
rect 1142 6323 1145 6326
rect 1154 6321 1157 6327
rect 1177 6322 1180 6328
rect 1227 6330 1230 6336
rect 1252 6331 1255 6336
rect 1149 6318 1157 6321
rect 1169 6319 1180 6322
rect 1209 6322 1212 6327
rect 1227 6326 1228 6330
rect 1247 6328 1250 6331
rect 1254 6327 1255 6331
rect 1273 6330 1276 6336
rect 1283 6330 1286 6336
rect 1227 6322 1230 6326
rect 1252 6322 1255 6327
rect 1267 6326 1276 6330
rect 1273 6322 1276 6326
rect 1283 6322 1286 6326
rect 1154 6315 1157 6318
rect 1299 6329 1302 6336
rect 1299 6325 1301 6329
rect 1319 6329 1320 6331
rect 1327 6331 1330 6336
rect 1324 6329 1330 6331
rect 1343 6330 1346 6336
rect 1319 6327 1330 6329
rect 1299 6322 1302 6325
rect 1327 6322 1330 6327
rect 1338 6326 1340 6330
rect 1344 6326 1346 6330
rect 1343 6322 1346 6326
rect 1352 6331 1355 6336
rect 1359 6331 1362 6336
rect 1914 6335 1917 6359
rect 1944 6331 1947 6359
rect 1352 6328 1362 6331
rect 1352 6322 1355 6328
rect 1359 6322 1362 6328
rect 1370 6328 1373 6331
rect 1905 6326 1908 6331
rect 1968 6327 1971 6359
rect 2004 6335 2007 6359
rect 1888 6323 1908 6326
rect 1228 6307 1230 6311
rect 1274 6307 1275 6311
rect 1299 6307 1302 6311
rect 1905 6309 1908 6323
rect 1916 6323 1919 6326
rect 1928 6321 1931 6327
rect 1923 6318 1931 6321
rect 1943 6320 1951 6322
rect 1943 6319 1955 6320
rect 2034 6331 2037 6359
rect 2041 6332 2046 6337
rect 1995 6326 1998 6331
rect 1959 6318 1962 6323
rect 1989 6323 1998 6326
rect 1928 6315 1931 6318
rect 1113 6297 1116 6301
rect 1140 6297 1143 6301
rect 1170 6297 1173 6307
rect 1209 6300 1223 6304
rect 1227 6300 1288 6304
rect 1292 6300 1310 6304
rect 1314 6300 1341 6304
rect 1345 6300 1421 6304
rect 1970 6315 1973 6318
rect 1914 6297 1917 6301
rect 1944 6297 1947 6307
rect 1959 6309 1962 6314
rect 1995 6309 1998 6323
rect 2006 6323 2009 6326
rect 2018 6321 2021 6327
rect 2041 6322 2044 6328
rect 2058 6327 2061 6359
rect 2085 6335 2088 6359
rect 2115 6331 2118 6359
rect 2154 6352 2183 6356
rect 2187 6352 2214 6356
rect 2218 6352 2239 6356
rect 2243 6352 2298 6356
rect 2302 6352 2378 6356
rect 2182 6345 2183 6349
rect 2229 6344 2230 6348
rect 2254 6345 2255 6349
rect 2122 6332 2127 6337
rect 2013 6318 2021 6321
rect 2033 6319 2044 6322
rect 2067 6326 2071 6330
rect 2076 6326 2079 6331
rect 2154 6331 2157 6336
rect 2049 6318 2052 6323
rect 2071 6323 2079 6326
rect 2018 6315 2021 6318
rect 2060 6315 2063 6318
rect 2067 6315 2068 6318
rect 1968 6297 1971 6301
rect 2004 6297 2007 6301
rect 2034 6297 2037 6307
rect 2049 6309 2052 6314
rect 2076 6309 2079 6323
rect 2087 6323 2090 6326
rect 2099 6321 2102 6327
rect 2122 6322 2125 6328
rect 2172 6330 2175 6336
rect 2197 6331 2200 6336
rect 2094 6318 2102 6321
rect 2114 6319 2125 6322
rect 2154 6322 2157 6327
rect 2172 6326 2173 6330
rect 2192 6328 2195 6331
rect 2199 6327 2200 6331
rect 2218 6330 2221 6336
rect 2228 6330 2231 6336
rect 2172 6322 2175 6326
rect 2197 6322 2200 6327
rect 2212 6326 2221 6330
rect 2218 6322 2221 6326
rect 2228 6322 2231 6326
rect 2099 6315 2102 6318
rect 2244 6329 2247 6336
rect 2244 6325 2246 6329
rect 2264 6329 2265 6331
rect 2272 6331 2275 6336
rect 2269 6329 2275 6331
rect 2288 6330 2291 6336
rect 2264 6327 2275 6329
rect 2244 6322 2247 6325
rect 2272 6322 2275 6327
rect 2283 6326 2285 6330
rect 2289 6326 2291 6330
rect 2288 6322 2291 6326
rect 2297 6331 2300 6336
rect 2304 6331 2307 6336
rect 2297 6328 2307 6331
rect 2297 6322 2300 6328
rect 2304 6322 2307 6328
rect 2315 6328 2318 6331
rect 4403 6325 4829 6421
rect 4786 6315 4829 6325
rect 2173 6307 2175 6311
rect 2219 6307 2220 6311
rect 2244 6307 2247 6311
rect 2058 6297 2061 6301
rect 2085 6297 2088 6301
rect 2115 6297 2118 6307
rect 4796 6305 4829 6315
rect 2154 6300 2168 6304
rect 2172 6300 2233 6304
rect 2237 6300 2255 6304
rect 2259 6300 2286 6304
rect 2290 6300 2366 6304
rect 955 6293 1005 6297
rect 1009 6293 1033 6297
rect 1037 6293 1041 6297
rect 1045 6293 1095 6297
rect 1099 6293 1122 6297
rect 1126 6293 1176 6297
rect 1180 6293 1200 6297
rect 1204 6293 1216 6297
rect 1220 6293 1244 6297
rect 1248 6293 1256 6297
rect 1260 6293 1261 6297
rect 1265 6293 1298 6297
rect 1302 6293 1317 6297
rect 1321 6293 1323 6297
rect 1327 6293 1334 6297
rect 1338 6293 1352 6297
rect 1356 6293 1368 6297
rect 1372 6293 1457 6297
rect 1900 6293 1950 6297
rect 1954 6293 1978 6297
rect 1982 6293 1986 6297
rect 1990 6293 2040 6297
rect 2044 6293 2067 6297
rect 2071 6293 2121 6297
rect 2125 6293 2145 6297
rect 2149 6293 2161 6297
rect 2165 6293 2189 6297
rect 2193 6293 2201 6297
rect 2205 6293 2206 6297
rect 2210 6293 2243 6297
rect 2247 6293 2262 6297
rect 2266 6293 2268 6297
rect 2272 6293 2279 6297
rect 2283 6293 2297 6297
rect 2301 6293 2313 6297
rect 2317 6293 2402 6297
rect 4806 6295 4829 6305
rect 546 6286 657 6290
rect 661 6286 662 6290
rect 666 6286 667 6290
rect 546 6285 667 6286
rect 546 6281 657 6285
rect 661 6281 662 6285
rect 666 6281 667 6285
rect 546 6280 667 6281
rect 418 6275 427 6280
rect 439 6275 443 6280
rect 459 6275 468 6280
rect 480 6275 484 6280
rect 502 6277 511 6280
rect 523 6277 527 6280
rect 546 6277 657 6280
rect 502 6276 657 6277
rect 661 6276 662 6280
rect 666 6276 667 6280
rect 502 6275 667 6276
rect 343 6233 346 6272
rect 418 6271 657 6275
rect 661 6271 662 6275
rect 666 6271 667 6275
rect 1065 6274 1068 6293
rect 1170 6274 1173 6293
rect 1209 6286 1223 6290
rect 1227 6286 1288 6290
rect 1292 6286 1310 6290
rect 1314 6286 1341 6290
rect 1345 6286 1421 6290
rect 1228 6279 1230 6283
rect 1274 6279 1275 6283
rect 1299 6279 1302 6283
rect 418 6270 667 6271
rect 418 6266 657 6270
rect 661 6266 662 6270
rect 666 6266 667 6270
rect 418 6265 667 6266
rect 418 6261 657 6265
rect 661 6261 662 6265
rect 666 6261 667 6265
rect 1049 6263 1052 6266
rect 1154 6263 1157 6266
rect 1209 6263 1212 6268
rect 1227 6264 1230 6268
rect 418 6260 667 6261
rect 418 6256 657 6260
rect 661 6256 662 6260
rect 666 6256 667 6260
rect 1044 6260 1052 6263
rect 418 6255 667 6256
rect 418 6251 657 6255
rect 661 6251 662 6255
rect 666 6251 667 6255
rect 418 6250 667 6251
rect 1049 6254 1052 6260
rect 1067 6259 1068 6262
rect 1072 6258 1077 6263
rect 1149 6260 1157 6263
rect 1154 6254 1157 6260
rect 1172 6259 1174 6262
rect 1178 6258 1183 6263
rect 1227 6260 1228 6264
rect 1252 6263 1255 6268
rect 1273 6264 1276 6268
rect 1283 6264 1286 6268
rect 1209 6254 1212 6259
rect 1227 6254 1230 6260
rect 1247 6259 1250 6262
rect 1254 6259 1255 6263
rect 1267 6260 1276 6264
rect 1252 6254 1255 6259
rect 1273 6254 1276 6260
rect 1283 6254 1286 6260
rect 1299 6265 1302 6268
rect 1299 6261 1301 6265
rect 1327 6263 1330 6268
rect 1343 6264 1346 6268
rect 1299 6254 1302 6261
rect 1319 6261 1330 6263
rect 1319 6259 1320 6261
rect 1324 6259 1330 6261
rect 1338 6260 1340 6264
rect 1344 6260 1346 6264
rect 1327 6254 1330 6259
rect 1343 6254 1346 6260
rect 1352 6262 1355 6268
rect 2010 6274 2013 6293
rect 2115 6274 2118 6293
rect 2154 6286 2168 6290
rect 2172 6286 2233 6290
rect 2237 6286 2255 6290
rect 2259 6286 2286 6290
rect 2290 6286 2366 6290
rect 4816 6285 4829 6295
rect 2173 6279 2175 6283
rect 2219 6279 2220 6283
rect 2244 6279 2247 6283
rect 1359 6262 1362 6268
rect 1994 6263 1997 6266
rect 2099 6263 2102 6266
rect 2154 6263 2157 6268
rect 2172 6264 2175 6268
rect 1352 6259 1362 6262
rect 1370 6259 1372 6262
rect 1352 6254 1355 6259
rect 1359 6254 1362 6259
rect 1989 6260 1997 6263
rect 1994 6254 1997 6260
rect 2012 6259 2013 6262
rect 2017 6258 2022 6263
rect 2094 6260 2102 6263
rect 2099 6254 2102 6260
rect 2117 6259 2119 6262
rect 2123 6258 2128 6263
rect 2172 6260 2173 6264
rect 2197 6263 2200 6268
rect 2218 6264 2221 6268
rect 2228 6264 2231 6268
rect 2154 6254 2157 6259
rect 2172 6254 2175 6260
rect 2192 6259 2195 6262
rect 2199 6259 2200 6263
rect 2212 6260 2221 6264
rect 2197 6254 2200 6259
rect 2218 6254 2221 6260
rect 2228 6254 2231 6260
rect 2244 6265 2247 6268
rect 2244 6261 2246 6265
rect 2272 6263 2275 6268
rect 2288 6264 2291 6268
rect 2244 6254 2247 6261
rect 2264 6261 2275 6263
rect 2264 6259 2265 6261
rect 2269 6259 2275 6261
rect 2283 6260 2285 6264
rect 2289 6260 2291 6264
rect 2272 6254 2275 6259
rect 2288 6254 2291 6260
rect 2297 6262 2300 6268
rect 2304 6262 2307 6268
rect 2297 6259 2307 6262
rect 2315 6259 2317 6262
rect 2297 6254 2300 6259
rect 2304 6254 2307 6259
rect 418 6246 657 6250
rect 661 6246 662 6250
rect 666 6246 667 6250
rect 418 6245 667 6246
rect 418 6241 657 6245
rect 661 6241 662 6245
rect 666 6241 667 6245
rect 418 6240 667 6241
rect 418 6236 657 6240
rect 661 6236 662 6240
rect 666 6236 667 6240
rect 418 6234 667 6236
rect 86 6230 346 6233
rect 1065 6231 1068 6250
rect 1170 6231 1173 6250
rect 1237 6241 1238 6245
rect 1284 6242 1285 6246
rect 1309 6241 1310 6245
rect 1209 6234 1238 6238
rect 1242 6234 1269 6238
rect 1273 6234 1294 6238
rect 1298 6234 1353 6238
rect 1357 6234 1433 6238
rect 2010 6231 2013 6250
rect 2115 6231 2118 6250
rect 4826 6246 4829 6285
rect 5083 6246 5086 6500
rect 2182 6241 2183 6245
rect 2229 6242 2230 6246
rect 2254 6241 2255 6245
rect 4483 6240 4484 6244
rect 4488 6240 4489 6244
rect 4493 6240 4494 6244
rect 4498 6240 4499 6244
rect 4503 6240 4504 6244
rect 4508 6240 4509 6244
rect 4479 6239 4513 6240
rect 2154 6234 2183 6238
rect 2187 6234 2214 6238
rect 2218 6234 2239 6238
rect 2243 6234 2298 6238
rect 2302 6234 2378 6238
rect 4483 6235 4484 6239
rect 4488 6235 4489 6239
rect 4493 6235 4494 6239
rect 4498 6235 4499 6239
rect 4503 6235 4504 6239
rect 4508 6235 4509 6239
rect 4479 6234 4513 6235
rect 617 6227 618 6231
rect 622 6227 623 6231
rect 627 6227 628 6231
rect 632 6227 633 6231
rect 637 6227 638 6231
rect 642 6227 643 6231
rect 613 6226 647 6227
rect 617 6222 618 6226
rect 622 6222 623 6226
rect 627 6222 628 6226
rect 632 6222 633 6226
rect 637 6222 638 6226
rect 642 6222 643 6226
rect 613 6221 647 6222
rect 617 6217 618 6221
rect 622 6217 623 6221
rect 627 6217 628 6221
rect 632 6217 633 6221
rect 637 6217 638 6221
rect 642 6217 643 6221
rect 613 6216 647 6217
rect 617 6212 618 6216
rect 622 6212 623 6216
rect 627 6212 628 6216
rect 632 6212 633 6216
rect 637 6212 638 6216
rect 642 6212 643 6216
rect 663 6227 664 6231
rect 668 6227 669 6231
rect 673 6227 674 6231
rect 678 6227 679 6231
rect 683 6227 684 6231
rect 688 6227 689 6231
rect 1023 6227 1071 6231
rect 1075 6227 1095 6231
rect 1099 6227 1122 6231
rect 1126 6227 1176 6231
rect 1180 6227 1200 6231
rect 1204 6227 1217 6231
rect 1221 6227 1245 6231
rect 1249 6227 1260 6231
rect 1264 6227 1294 6231
rect 1298 6227 1317 6231
rect 1321 6227 1326 6231
rect 1330 6227 1335 6231
rect 1339 6227 1353 6231
rect 1357 6227 1361 6231
rect 1365 6227 1367 6231
rect 1371 6227 1445 6231
rect 1968 6227 2016 6231
rect 2020 6227 2040 6231
rect 2044 6227 2067 6231
rect 2071 6227 2121 6231
rect 2125 6227 2145 6231
rect 2149 6227 2162 6231
rect 2166 6227 2190 6231
rect 2194 6227 2205 6231
rect 2209 6227 2239 6231
rect 2243 6227 2262 6231
rect 2266 6227 2271 6231
rect 2275 6227 2280 6231
rect 2284 6227 2298 6231
rect 2302 6227 2306 6231
rect 2310 6227 2312 6231
rect 2316 6227 2390 6231
rect 4483 6230 4484 6234
rect 4488 6230 4489 6234
rect 4493 6230 4494 6234
rect 4498 6230 4499 6234
rect 4503 6230 4504 6234
rect 4508 6230 4509 6234
rect 4479 6229 4513 6230
rect 659 6226 693 6227
rect 663 6222 664 6226
rect 668 6222 669 6226
rect 673 6222 674 6226
rect 678 6222 679 6226
rect 683 6222 684 6226
rect 688 6222 689 6226
rect 659 6221 693 6222
rect 663 6217 664 6221
rect 668 6217 669 6221
rect 673 6217 674 6221
rect 678 6217 679 6221
rect 683 6217 684 6221
rect 688 6217 689 6221
rect 659 6216 693 6217
rect 663 6212 664 6216
rect 668 6212 669 6216
rect 673 6212 674 6216
rect 678 6212 679 6216
rect 683 6212 684 6216
rect 688 6212 689 6216
rect 1035 6203 1038 6227
rect 617 6196 618 6200
rect 622 6196 623 6200
rect 627 6196 628 6200
rect 632 6196 633 6200
rect 637 6196 638 6200
rect 642 6196 643 6200
rect 613 6195 647 6196
rect 617 6191 618 6195
rect 622 6191 623 6195
rect 627 6191 628 6195
rect 632 6191 633 6195
rect 637 6191 638 6195
rect 642 6191 643 6195
rect 613 6190 647 6191
rect 617 6186 618 6190
rect 622 6186 623 6190
rect 627 6186 628 6190
rect 632 6186 633 6190
rect 637 6186 638 6190
rect 642 6186 643 6190
rect 613 6185 647 6186
rect 86 6179 346 6182
rect 617 6181 618 6185
rect 622 6181 623 6185
rect 627 6181 628 6185
rect 632 6181 633 6185
rect 637 6181 638 6185
rect 642 6181 643 6185
rect 663 6196 664 6200
rect 668 6196 669 6200
rect 673 6196 674 6200
rect 678 6196 679 6200
rect 683 6196 684 6200
rect 688 6196 689 6200
rect 659 6195 693 6196
rect 663 6191 664 6195
rect 668 6191 669 6195
rect 673 6191 674 6195
rect 678 6191 679 6195
rect 683 6191 684 6195
rect 688 6191 689 6195
rect 1065 6199 1068 6227
rect 1072 6200 1077 6205
rect 1026 6194 1029 6199
rect 659 6190 693 6191
rect 1023 6191 1029 6194
rect 663 6186 664 6190
rect 668 6186 669 6190
rect 673 6186 674 6190
rect 678 6186 679 6190
rect 683 6186 684 6190
rect 688 6186 689 6190
rect 659 6185 693 6186
rect 663 6181 664 6185
rect 668 6181 669 6185
rect 673 6181 674 6185
rect 678 6181 679 6185
rect 683 6181 684 6185
rect 688 6181 689 6185
rect 86 5925 89 6179
rect 343 6140 346 6179
rect 1026 6177 1029 6191
rect 1037 6191 1040 6194
rect 1049 6189 1052 6195
rect 1072 6190 1075 6196
rect 1089 6195 1092 6227
rect 1140 6203 1143 6227
rect 1170 6199 1173 6227
rect 1209 6220 1238 6224
rect 1242 6220 1269 6224
rect 1273 6220 1294 6224
rect 1298 6220 1353 6224
rect 1357 6220 1433 6224
rect 1237 6213 1238 6217
rect 1284 6212 1285 6216
rect 1309 6213 1310 6217
rect 1177 6200 1182 6205
rect 1044 6186 1052 6189
rect 1064 6187 1075 6190
rect 1131 6194 1134 6199
rect 1209 6199 1212 6204
rect 1126 6191 1134 6194
rect 1080 6186 1083 6191
rect 1121 6186 1126 6191
rect 1049 6183 1052 6186
rect 1091 6183 1094 6186
rect 1098 6183 1099 6186
rect 1035 6165 1038 6169
rect 1065 6165 1068 6175
rect 1080 6177 1083 6182
rect 1131 6177 1134 6191
rect 1142 6191 1145 6194
rect 1154 6189 1157 6195
rect 1177 6190 1180 6196
rect 1227 6198 1230 6204
rect 1252 6199 1255 6204
rect 1149 6186 1157 6189
rect 1169 6187 1180 6190
rect 1209 6190 1212 6195
rect 1227 6194 1228 6198
rect 1247 6196 1250 6199
rect 1254 6195 1255 6199
rect 1273 6198 1276 6204
rect 1283 6198 1286 6204
rect 1227 6190 1230 6194
rect 1252 6190 1255 6195
rect 1267 6194 1276 6198
rect 1273 6190 1276 6194
rect 1283 6190 1286 6194
rect 1154 6183 1157 6186
rect 1299 6197 1302 6204
rect 1299 6193 1301 6197
rect 1319 6197 1320 6199
rect 1327 6199 1330 6204
rect 1324 6197 1330 6199
rect 1343 6198 1346 6204
rect 1319 6195 1330 6197
rect 1299 6190 1302 6193
rect 1327 6190 1330 6195
rect 1338 6194 1340 6198
rect 1344 6194 1346 6198
rect 1343 6190 1346 6194
rect 1352 6199 1355 6204
rect 1359 6199 1362 6204
rect 1980 6203 1983 6227
rect 2010 6199 2013 6227
rect 2017 6200 2022 6205
rect 1352 6196 1362 6199
rect 1352 6190 1355 6196
rect 1359 6190 1362 6196
rect 1370 6196 1373 6199
rect 1971 6194 1974 6199
rect 1968 6191 1974 6194
rect 1228 6175 1230 6179
rect 1274 6175 1275 6179
rect 1299 6175 1302 6179
rect 1971 6177 1974 6191
rect 1982 6191 1985 6194
rect 1994 6189 1997 6195
rect 2017 6190 2020 6196
rect 2034 6195 2037 6227
rect 2085 6203 2088 6227
rect 2115 6199 2118 6227
rect 4483 6225 4484 6229
rect 4488 6225 4489 6229
rect 4493 6225 4494 6229
rect 4498 6225 4499 6229
rect 4503 6225 4504 6229
rect 4508 6225 4509 6229
rect 4529 6240 4530 6244
rect 4534 6240 4535 6244
rect 4539 6240 4540 6244
rect 4544 6240 4545 6244
rect 4549 6240 4550 6244
rect 4554 6240 4555 6244
rect 4826 6243 5086 6246
rect 4525 6239 4559 6240
rect 4529 6235 4530 6239
rect 4534 6235 4535 6239
rect 4539 6235 4540 6239
rect 4544 6235 4545 6239
rect 4549 6235 4550 6239
rect 4554 6235 4555 6239
rect 4525 6234 4559 6235
rect 4529 6230 4530 6234
rect 4534 6230 4535 6234
rect 4539 6230 4540 6234
rect 4544 6230 4545 6234
rect 4549 6230 4550 6234
rect 4554 6230 4555 6234
rect 4525 6229 4559 6230
rect 4529 6225 4530 6229
rect 4534 6225 4535 6229
rect 4539 6225 4540 6229
rect 4544 6225 4545 6229
rect 4549 6225 4550 6229
rect 4554 6225 4555 6229
rect 2154 6220 2183 6224
rect 2187 6220 2214 6224
rect 2218 6220 2239 6224
rect 2243 6220 2298 6224
rect 2302 6220 2378 6224
rect 2182 6213 2183 6217
rect 2229 6212 2230 6216
rect 2254 6213 2255 6217
rect 2122 6200 2127 6205
rect 1989 6186 1997 6189
rect 2009 6187 2020 6190
rect 2076 6194 2079 6199
rect 2154 6199 2157 6204
rect 2071 6191 2079 6194
rect 2025 6186 2028 6191
rect 2066 6186 2071 6191
rect 1994 6183 1997 6186
rect 1089 6165 1092 6169
rect 1140 6165 1143 6169
rect 1170 6165 1173 6175
rect 1209 6168 1223 6172
rect 1227 6168 1288 6172
rect 1292 6168 1310 6172
rect 1314 6168 1341 6172
rect 1345 6168 1357 6172
rect 1361 6168 1421 6172
rect 2036 6183 2039 6186
rect 2043 6183 2044 6186
rect 1980 6165 1983 6169
rect 2010 6165 2013 6175
rect 2025 6177 2028 6182
rect 2076 6177 2079 6191
rect 2087 6191 2090 6194
rect 2099 6189 2102 6195
rect 2122 6190 2125 6196
rect 2172 6198 2175 6204
rect 2197 6199 2200 6204
rect 2094 6186 2102 6189
rect 2114 6187 2125 6190
rect 2154 6190 2157 6195
rect 2172 6194 2173 6198
rect 2192 6196 2195 6199
rect 2199 6195 2200 6199
rect 2218 6198 2221 6204
rect 2228 6198 2231 6204
rect 2172 6190 2175 6194
rect 2197 6190 2200 6195
rect 2212 6194 2221 6198
rect 2218 6190 2221 6194
rect 2228 6190 2231 6194
rect 2099 6183 2102 6186
rect 2244 6197 2247 6204
rect 2244 6193 2246 6197
rect 2264 6197 2265 6199
rect 2272 6199 2275 6204
rect 2269 6197 2275 6199
rect 2288 6198 2291 6204
rect 2264 6195 2275 6197
rect 2244 6190 2247 6193
rect 2272 6190 2275 6195
rect 2283 6194 2285 6198
rect 2289 6194 2291 6198
rect 2288 6190 2291 6194
rect 2297 6199 2300 6204
rect 2304 6199 2307 6204
rect 2297 6196 2307 6199
rect 2297 6190 2300 6196
rect 2304 6190 2307 6196
rect 2315 6196 2318 6199
rect 4826 6191 5086 6194
rect 2173 6175 2175 6179
rect 2219 6175 2220 6179
rect 2244 6175 2247 6179
rect 2034 6165 2037 6169
rect 2085 6165 2088 6169
rect 2115 6165 2118 6175
rect 2154 6168 2168 6172
rect 2172 6168 2233 6172
rect 2237 6168 2255 6172
rect 2259 6168 2286 6172
rect 2290 6168 2302 6172
rect 2306 6168 2366 6172
rect 1022 6161 1033 6165
rect 1037 6161 1095 6165
rect 1099 6161 1122 6165
rect 1126 6161 1176 6165
rect 1180 6161 1200 6165
rect 1204 6161 1216 6165
rect 1220 6161 1244 6165
rect 1248 6161 1256 6165
rect 1260 6161 1261 6165
rect 1265 6161 1298 6165
rect 1302 6161 1317 6165
rect 1321 6161 1323 6165
rect 1327 6161 1334 6165
rect 1338 6161 1352 6165
rect 1356 6161 1368 6165
rect 1372 6161 1457 6165
rect 1967 6161 1978 6165
rect 1982 6161 2040 6165
rect 2044 6161 2067 6165
rect 2071 6161 2121 6165
rect 2125 6161 2145 6165
rect 2149 6161 2161 6165
rect 2165 6161 2189 6165
rect 2193 6161 2201 6165
rect 2205 6161 2206 6165
rect 2210 6161 2243 6165
rect 2247 6161 2262 6165
rect 2266 6161 2268 6165
rect 2272 6161 2279 6165
rect 2283 6161 2297 6165
rect 2301 6161 2313 6165
rect 2317 6161 2402 6165
rect 1089 6143 1092 6161
rect 1170 6143 1173 6161
rect 1209 6154 1223 6158
rect 1227 6154 1288 6158
rect 1292 6154 1310 6158
rect 1314 6154 1341 6158
rect 1345 6154 1357 6158
rect 1415 6151 1615 6155
rect 1619 6151 1666 6155
rect 1670 6151 1716 6155
rect 1720 6151 1738 6155
rect 1228 6147 1230 6151
rect 1274 6147 1275 6151
rect 1299 6147 1302 6151
rect 1451 6144 1639 6148
rect 1643 6144 1667 6148
rect 1671 6144 1697 6148
rect 1701 6144 1738 6148
rect 343 6130 356 6140
rect 1073 6132 1076 6135
rect 1154 6132 1157 6135
rect 343 6120 366 6130
rect 1068 6129 1076 6132
rect 1073 6123 1076 6129
rect 1091 6128 1093 6131
rect 1097 6127 1102 6132
rect 1149 6129 1157 6132
rect 1154 6123 1157 6129
rect 1172 6128 1173 6131
rect 1177 6127 1182 6132
rect 1209 6131 1212 6136
rect 1227 6132 1230 6136
rect 1227 6128 1228 6132
rect 1252 6131 1255 6136
rect 1273 6132 1276 6136
rect 1283 6132 1286 6136
rect 343 6110 376 6120
rect 343 6100 386 6110
rect 343 6004 769 6100
rect 1089 6099 1092 6119
rect 1170 6099 1173 6119
rect 1209 6122 1212 6127
rect 1227 6122 1230 6128
rect 1247 6127 1250 6130
rect 1254 6127 1255 6131
rect 1267 6128 1276 6132
rect 1252 6122 1255 6127
rect 1273 6122 1276 6128
rect 1283 6122 1286 6128
rect 1299 6133 1302 6136
rect 1299 6129 1301 6133
rect 1327 6131 1330 6136
rect 1343 6132 1346 6136
rect 1299 6122 1302 6129
rect 1319 6129 1330 6131
rect 1319 6127 1320 6129
rect 1324 6127 1330 6129
rect 1338 6128 1340 6132
rect 1344 6128 1346 6132
rect 1327 6122 1330 6127
rect 1343 6122 1346 6128
rect 1352 6130 1355 6136
rect 1359 6130 1362 6136
rect 1609 6132 1612 6144
rect 1630 6132 1633 6144
rect 1646 6132 1649 6144
rect 1660 6138 1672 6141
rect 1688 6132 1691 6144
rect 1704 6132 1707 6144
rect 1725 6132 1728 6144
rect 2034 6143 2037 6161
rect 2115 6143 2118 6161
rect 2154 6154 2168 6158
rect 2172 6154 2233 6158
rect 2237 6154 2255 6158
rect 2259 6154 2286 6158
rect 2290 6154 2302 6158
rect 2360 6151 2560 6155
rect 2564 6151 2611 6155
rect 2615 6151 2661 6155
rect 2665 6151 2683 6155
rect 4826 6152 4829 6191
rect 2173 6147 2175 6151
rect 2219 6147 2220 6151
rect 2244 6147 2247 6151
rect 2396 6144 2584 6148
rect 2588 6144 2612 6148
rect 2616 6144 2642 6148
rect 2646 6144 2683 6148
rect 2018 6132 2021 6135
rect 2099 6132 2102 6135
rect 1352 6127 1362 6130
rect 1370 6127 1372 6130
rect 1352 6122 1355 6127
rect 1359 6122 1362 6127
rect 1642 6122 1649 6125
rect 2013 6129 2021 6132
rect 1672 6122 1675 6128
rect 1700 6122 1707 6125
rect 1653 6118 1672 6121
rect 2018 6123 2021 6129
rect 2036 6128 2038 6131
rect 2042 6127 2047 6132
rect 2094 6129 2102 6132
rect 2099 6123 2102 6129
rect 2117 6128 2118 6131
rect 2122 6127 2127 6132
rect 2154 6131 2157 6136
rect 2172 6132 2175 6136
rect 2172 6128 2173 6132
rect 2197 6131 2200 6136
rect 2218 6132 2221 6136
rect 2228 6132 2231 6136
rect 1711 6118 1726 6121
rect 1604 6114 1613 6118
rect 1237 6109 1238 6113
rect 1284 6110 1285 6114
rect 1309 6109 1310 6113
rect 1626 6112 1631 6115
rect 1635 6112 1659 6115
rect 1209 6102 1238 6106
rect 1242 6102 1269 6106
rect 1273 6102 1294 6106
rect 1298 6102 1353 6106
rect 1357 6102 1433 6106
rect 1684 6112 1691 6115
rect 1695 6112 1717 6115
rect 1045 6095 1095 6099
rect 1099 6095 1119 6099
rect 1126 6095 1176 6099
rect 1180 6095 1200 6099
rect 1204 6095 1217 6099
rect 1221 6095 1245 6099
rect 1249 6095 1260 6099
rect 1264 6095 1294 6099
rect 1298 6095 1317 6099
rect 1321 6095 1326 6099
rect 1330 6095 1335 6099
rect 1339 6095 1353 6099
rect 1357 6095 1361 6099
rect 1365 6095 1367 6099
rect 1371 6095 1445 6099
rect 1059 6071 1062 6095
rect 1089 6067 1092 6095
rect 1096 6068 1101 6073
rect 1050 6062 1053 6067
rect 1041 6059 1053 6062
rect 1050 6045 1053 6059
rect 1061 6059 1064 6062
rect 1073 6057 1076 6063
rect 1096 6058 1099 6064
rect 1113 6063 1116 6095
rect 1140 6071 1143 6095
rect 1170 6067 1173 6095
rect 1177 6068 1182 6073
rect 1068 6054 1076 6057
rect 1088 6055 1099 6058
rect 1122 6062 1126 6066
rect 1131 6062 1134 6067
rect 1104 6054 1107 6059
rect 1126 6059 1134 6062
rect 1073 6051 1076 6054
rect 1115 6051 1118 6054
rect 1122 6051 1123 6054
rect 1059 6033 1062 6037
rect 1089 6033 1092 6043
rect 1104 6045 1107 6050
rect 1131 6045 1134 6059
rect 1142 6059 1145 6062
rect 1154 6057 1157 6063
rect 1177 6058 1180 6064
rect 1194 6063 1197 6095
rect 1209 6088 1238 6092
rect 1242 6088 1269 6092
rect 1273 6088 1294 6092
rect 1298 6088 1353 6092
rect 1357 6088 1433 6092
rect 1609 6091 1612 6101
rect 1630 6091 1633 6101
rect 1646 6091 1649 6101
rect 1660 6094 1665 6098
rect 1669 6094 1676 6098
rect 1688 6091 1691 6101
rect 1704 6091 1707 6101
rect 1725 6091 1728 6101
rect 2034 6099 2037 6119
rect 2115 6099 2118 6119
rect 2154 6122 2157 6127
rect 2172 6122 2175 6128
rect 2192 6127 2195 6130
rect 2199 6127 2200 6131
rect 2212 6128 2221 6132
rect 2197 6122 2200 6127
rect 2218 6122 2221 6128
rect 2228 6122 2231 6128
rect 2244 6133 2247 6136
rect 2244 6129 2246 6133
rect 2272 6131 2275 6136
rect 2288 6132 2291 6136
rect 2244 6122 2247 6129
rect 2264 6129 2275 6131
rect 2264 6127 2265 6129
rect 2269 6127 2275 6129
rect 2283 6128 2285 6132
rect 2289 6128 2291 6132
rect 2272 6122 2275 6127
rect 2288 6122 2291 6128
rect 2297 6130 2300 6136
rect 2304 6130 2307 6136
rect 2554 6132 2557 6144
rect 2575 6132 2578 6144
rect 2591 6132 2594 6144
rect 2605 6138 2617 6141
rect 2633 6132 2636 6144
rect 2649 6132 2652 6144
rect 2670 6132 2673 6144
rect 4816 6142 4829 6152
rect 4806 6132 4829 6142
rect 2297 6127 2307 6130
rect 2315 6127 2317 6130
rect 2297 6122 2300 6127
rect 2304 6122 2307 6127
rect 2587 6122 2594 6125
rect 2617 6122 2620 6128
rect 2645 6122 2652 6125
rect 2598 6118 2617 6121
rect 4796 6122 4829 6132
rect 2656 6118 2671 6121
rect 2549 6114 2558 6118
rect 2182 6109 2183 6113
rect 2229 6110 2230 6114
rect 2254 6109 2255 6113
rect 2571 6112 2576 6115
rect 2580 6112 2604 6115
rect 2154 6102 2183 6106
rect 2187 6102 2214 6106
rect 2218 6102 2239 6106
rect 2243 6102 2298 6106
rect 2302 6102 2378 6106
rect 2629 6112 2636 6115
rect 2640 6112 2662 6115
rect 4786 6112 4829 6122
rect 1990 6095 2040 6099
rect 2044 6095 2064 6099
rect 2071 6095 2121 6099
rect 2125 6095 2145 6099
rect 2149 6095 2162 6099
rect 2166 6095 2190 6099
rect 2194 6095 2205 6099
rect 2209 6095 2239 6099
rect 2243 6095 2262 6099
rect 2266 6095 2271 6099
rect 2275 6095 2280 6099
rect 2284 6095 2298 6099
rect 2302 6095 2306 6099
rect 2310 6095 2312 6099
rect 2316 6095 2390 6099
rect 1463 6087 1639 6091
rect 1643 6087 1667 6091
rect 1671 6087 1697 6091
rect 1701 6087 1734 6091
rect 1237 6081 1238 6085
rect 1284 6080 1285 6084
rect 1309 6081 1310 6085
rect 1403 6080 1615 6084
rect 1619 6080 1651 6084
rect 1655 6080 1718 6084
rect 1722 6080 1738 6084
rect 1209 6067 1212 6072
rect 1227 6066 1230 6072
rect 1252 6067 1255 6072
rect 1149 6054 1157 6057
rect 1169 6055 1180 6058
rect 1185 6054 1188 6059
rect 1209 6058 1212 6063
rect 1227 6062 1228 6066
rect 1247 6064 1250 6067
rect 1254 6063 1255 6067
rect 1273 6066 1276 6072
rect 1283 6066 1286 6072
rect 1227 6058 1230 6062
rect 1252 6058 1255 6063
rect 1267 6062 1276 6066
rect 1273 6058 1276 6062
rect 1283 6058 1286 6062
rect 1154 6051 1157 6054
rect 1196 6051 1199 6054
rect 1299 6065 1302 6072
rect 1299 6061 1301 6065
rect 1319 6065 1320 6067
rect 1327 6067 1330 6072
rect 1324 6065 1330 6067
rect 1343 6066 1346 6072
rect 1319 6063 1330 6065
rect 1299 6058 1302 6061
rect 1327 6058 1330 6063
rect 1338 6062 1340 6066
rect 1344 6062 1346 6066
rect 1343 6058 1346 6062
rect 1352 6067 1355 6072
rect 1588 6072 1709 6076
rect 1721 6072 1725 6076
rect 1359 6067 1362 6072
rect 2004 6071 2007 6095
rect 1352 6064 1362 6067
rect 1352 6058 1355 6064
rect 1359 6058 1362 6064
rect 1370 6063 1584 6067
rect 1588 6063 1592 6067
rect 1604 6063 1608 6067
rect 1717 6065 1733 6069
rect 2034 6067 2037 6095
rect 2041 6068 2046 6073
rect 1995 6062 1998 6067
rect 1986 6059 1998 6062
rect 1113 6033 1116 6037
rect 1140 6033 1143 6037
rect 1170 6033 1173 6043
rect 1185 6045 1188 6050
rect 1228 6043 1230 6047
rect 1274 6043 1275 6047
rect 1299 6043 1302 6047
rect 1415 6049 1617 6053
rect 1621 6049 1667 6053
rect 1671 6049 1718 6053
rect 1722 6049 1731 6053
rect 1451 6042 1636 6046
rect 1640 6042 1666 6046
rect 1670 6042 1694 6046
rect 1698 6042 1731 6046
rect 1995 6045 1998 6059
rect 2006 6059 2009 6062
rect 2018 6057 2021 6063
rect 2041 6058 2044 6064
rect 2058 6063 2061 6095
rect 2085 6071 2088 6095
rect 2115 6067 2118 6095
rect 2122 6068 2127 6073
rect 2013 6054 2021 6057
rect 2033 6055 2044 6058
rect 2067 6062 2071 6066
rect 2076 6062 2079 6067
rect 2049 6054 2052 6059
rect 2071 6059 2079 6062
rect 2018 6051 2021 6054
rect 1194 6033 1197 6037
rect 1209 6036 1223 6040
rect 1227 6036 1288 6040
rect 1292 6036 1310 6040
rect 1314 6036 1341 6040
rect 1345 6036 1421 6040
rect 1022 6029 1041 6033
rect 1045 6029 1095 6033
rect 1099 6029 1122 6033
rect 1126 6029 1176 6033
rect 1180 6029 1200 6033
rect 1204 6029 1216 6033
rect 1220 6029 1244 6033
rect 1248 6029 1256 6033
rect 1260 6029 1261 6033
rect 1265 6029 1298 6033
rect 1302 6029 1317 6033
rect 1321 6029 1323 6033
rect 1327 6029 1334 6033
rect 1338 6029 1352 6033
rect 1356 6029 1368 6033
rect 1372 6029 1457 6033
rect 1609 6030 1612 6042
rect 1630 6030 1633 6042
rect 1646 6030 1649 6042
rect 1665 6036 1677 6039
rect 1688 6030 1691 6042
rect 1704 6030 1707 6042
rect 1725 6030 1728 6042
rect 2060 6051 2063 6054
rect 2067 6051 2068 6054
rect 2004 6033 2007 6037
rect 2034 6033 2037 6043
rect 2049 6045 2052 6050
rect 2076 6045 2079 6059
rect 2087 6059 2090 6062
rect 2099 6057 2102 6063
rect 2122 6058 2125 6064
rect 2139 6063 2142 6095
rect 2154 6088 2183 6092
rect 2187 6088 2214 6092
rect 2218 6088 2239 6092
rect 2243 6088 2298 6092
rect 2302 6088 2378 6092
rect 2554 6091 2557 6101
rect 2575 6091 2578 6101
rect 2591 6091 2594 6101
rect 2605 6094 2610 6098
rect 2614 6094 2621 6098
rect 2633 6091 2636 6101
rect 2649 6091 2652 6101
rect 2670 6091 2673 6101
rect 2408 6087 2584 6091
rect 2588 6087 2612 6091
rect 2616 6087 2642 6091
rect 2646 6087 2679 6091
rect 2182 6081 2183 6085
rect 2229 6080 2230 6084
rect 2254 6081 2255 6085
rect 2348 6080 2560 6084
rect 2564 6080 2596 6084
rect 2600 6080 2663 6084
rect 2667 6080 2683 6084
rect 2154 6067 2157 6072
rect 2172 6066 2175 6072
rect 2197 6067 2200 6072
rect 2094 6054 2102 6057
rect 2114 6055 2125 6058
rect 2130 6054 2133 6059
rect 2154 6058 2157 6063
rect 2172 6062 2173 6066
rect 2192 6064 2195 6067
rect 2199 6063 2200 6067
rect 2218 6066 2221 6072
rect 2228 6066 2231 6072
rect 2172 6058 2175 6062
rect 2197 6058 2200 6063
rect 2212 6062 2221 6066
rect 2218 6058 2221 6062
rect 2228 6058 2231 6062
rect 2099 6051 2102 6054
rect 2141 6051 2144 6054
rect 2244 6065 2247 6072
rect 2244 6061 2246 6065
rect 2264 6065 2265 6067
rect 2272 6067 2275 6072
rect 2269 6065 2275 6067
rect 2288 6066 2291 6072
rect 2264 6063 2275 6065
rect 2244 6058 2247 6061
rect 2272 6058 2275 6063
rect 2283 6062 2285 6066
rect 2289 6062 2291 6066
rect 2288 6058 2291 6062
rect 2297 6067 2300 6072
rect 2533 6072 2654 6076
rect 2666 6072 2670 6076
rect 2304 6067 2307 6072
rect 2297 6064 2307 6067
rect 2297 6058 2300 6064
rect 2304 6058 2307 6064
rect 2315 6063 2529 6067
rect 2533 6063 2537 6067
rect 2549 6063 2553 6067
rect 2662 6065 2678 6069
rect 2058 6033 2061 6037
rect 2085 6033 2088 6037
rect 2115 6033 2118 6043
rect 2130 6045 2133 6050
rect 2173 6043 2175 6047
rect 2219 6043 2220 6047
rect 2244 6043 2247 6047
rect 2360 6049 2562 6053
rect 2566 6049 2612 6053
rect 2616 6049 2663 6053
rect 2667 6049 2676 6053
rect 2396 6042 2581 6046
rect 2585 6042 2611 6046
rect 2615 6042 2639 6046
rect 2643 6042 2676 6046
rect 2139 6033 2142 6037
rect 2154 6036 2168 6040
rect 2172 6036 2233 6040
rect 2237 6036 2255 6040
rect 2259 6036 2286 6040
rect 2290 6036 2366 6040
rect 851 6016 869 6020
rect 873 6016 919 6020
rect 923 6016 970 6020
rect 974 6016 1001 6020
rect 1005 6016 1051 6020
rect 1055 6016 1102 6020
rect 1106 6016 1133 6020
rect 1137 6016 1183 6020
rect 1187 6016 1234 6020
rect 1238 6016 1265 6020
rect 1269 6016 1315 6020
rect 1319 6016 1366 6020
rect 1370 6016 1409 6020
rect 1611 6016 1626 6019
rect 1630 6020 1637 6023
rect 1662 6020 1665 6026
rect 1967 6029 1986 6033
rect 1990 6029 2040 6033
rect 2044 6029 2067 6033
rect 2071 6029 2121 6033
rect 2125 6029 2145 6033
rect 2149 6029 2161 6033
rect 2165 6029 2189 6033
rect 2193 6029 2201 6033
rect 2205 6029 2206 6033
rect 2210 6029 2243 6033
rect 2247 6029 2262 6033
rect 2266 6029 2268 6033
rect 2272 6029 2279 6033
rect 2283 6029 2297 6033
rect 2301 6029 2313 6033
rect 2317 6029 2402 6033
rect 2554 6030 2557 6042
rect 2575 6030 2578 6042
rect 2591 6030 2594 6042
rect 2610 6036 2622 6039
rect 2633 6030 2636 6042
rect 2649 6030 2652 6042
rect 2670 6030 2673 6042
rect 1665 6016 1684 6019
rect 1688 6020 1695 6023
rect 1796 6016 1814 6020
rect 1818 6016 1864 6020
rect 1868 6016 1915 6020
rect 1919 6016 1946 6020
rect 1950 6016 1996 6020
rect 2000 6016 2047 6020
rect 2051 6016 2078 6020
rect 2082 6016 2128 6020
rect 2132 6016 2179 6020
rect 2183 6016 2210 6020
rect 2214 6016 2260 6020
rect 2264 6016 2311 6020
rect 2315 6016 2354 6020
rect 851 6009 888 6013
rect 892 6009 918 6013
rect 922 6009 946 6013
rect 950 6009 1020 6013
rect 1024 6009 1050 6013
rect 1054 6009 1078 6013
rect 1082 6009 1152 6013
rect 1156 6009 1182 6013
rect 1186 6009 1210 6013
rect 1214 6009 1284 6013
rect 1288 6009 1314 6013
rect 1318 6009 1342 6013
rect 1346 6009 1445 6013
rect 343 5994 386 6004
rect 861 5997 864 6009
rect 882 5997 885 6009
rect 898 5997 901 6009
rect 917 6003 929 6006
rect 940 5997 943 6009
rect 956 5997 959 6009
rect 977 5997 980 6009
rect 343 5984 376 5994
rect 343 5974 366 5984
rect 861 5983 878 5986
rect 882 5987 889 5990
rect 914 5987 917 5993
rect 993 5997 996 6009
rect 1014 5997 1017 6009
rect 1030 5997 1033 6009
rect 1049 6003 1061 6006
rect 1072 5997 1075 6009
rect 1088 5997 1091 6009
rect 1109 5997 1112 6009
rect 1125 5997 1128 6009
rect 1146 5997 1149 6009
rect 1162 5997 1165 6009
rect 1181 6003 1193 6006
rect 1204 5997 1207 6009
rect 1220 5997 1223 6009
rect 1241 5997 1244 6009
rect 1257 5997 1260 6009
rect 1278 5997 1281 6009
rect 1294 5997 1297 6009
rect 1313 6003 1325 6006
rect 1336 5997 1339 6009
rect 1352 5997 1355 6009
rect 1373 5997 1376 6009
rect 1620 6010 1642 6013
rect 1646 6010 1653 6013
rect 1678 6010 1702 6013
rect 1706 6010 1711 6013
rect 1724 6012 1733 6016
rect 2556 6016 2571 6019
rect 2575 6020 2582 6023
rect 2607 6020 2610 6026
rect 2610 6016 2629 6019
rect 2633 6020 2640 6023
rect 4403 6016 4829 6112
rect 1796 6009 1833 6013
rect 1837 6009 1863 6013
rect 1867 6009 1891 6013
rect 1895 6009 1965 6013
rect 1969 6009 1995 6013
rect 1999 6009 2023 6013
rect 2027 6009 2097 6013
rect 2101 6009 2127 6013
rect 2131 6009 2155 6013
rect 2159 6009 2229 6013
rect 2233 6009 2259 6013
rect 2263 6009 2287 6013
rect 2291 6009 2390 6013
rect 917 5983 936 5986
rect 940 5987 947 5990
rect 872 5977 894 5980
rect 898 5977 905 5980
rect 343 5964 356 5974
rect 930 5977 954 5980
rect 958 5977 963 5980
rect 993 5983 1010 5986
rect 1014 5987 1021 5990
rect 1046 5987 1049 5993
rect 1049 5983 1068 5986
rect 1072 5987 1079 5990
rect 1004 5977 1026 5980
rect 1030 5977 1037 5980
rect 1062 5977 1086 5980
rect 1090 5977 1095 5980
rect 1125 5983 1142 5986
rect 1146 5987 1153 5990
rect 1178 5987 1181 5993
rect 1181 5983 1200 5986
rect 1204 5987 1211 5990
rect 1136 5977 1158 5980
rect 1162 5977 1169 5980
rect 1194 5977 1218 5980
rect 1222 5977 1227 5980
rect 1257 5983 1274 5986
rect 1278 5987 1285 5990
rect 1310 5987 1313 5993
rect 1313 5983 1332 5986
rect 1336 5987 1343 5990
rect 1609 5989 1612 5999
rect 1630 5989 1633 5999
rect 1646 5989 1649 5999
rect 1661 5992 1668 5996
rect 1672 5992 1677 5996
rect 1688 5989 1691 5999
rect 1704 5989 1707 5999
rect 1725 5989 1728 5999
rect 1806 5997 1809 6009
rect 1827 5997 1830 6009
rect 1843 5997 1846 6009
rect 1862 6003 1874 6006
rect 1885 5997 1888 6009
rect 1901 5997 1904 6009
rect 1922 5997 1925 6009
rect 1463 5985 1599 5989
rect 1603 5985 1636 5989
rect 1640 5985 1666 5989
rect 1670 5985 1694 5989
rect 1698 5985 1731 5989
rect 1268 5977 1290 5980
rect 1294 5977 1301 5980
rect 1326 5977 1350 5980
rect 1354 5977 1359 5980
rect 1806 5983 1823 5986
rect 1827 5987 1834 5990
rect 1859 5987 1862 5993
rect 1938 5997 1941 6009
rect 1959 5997 1962 6009
rect 1975 5997 1978 6009
rect 1994 6003 2006 6006
rect 2017 5997 2020 6009
rect 2033 5997 2036 6009
rect 2054 5997 2057 6009
rect 2070 5997 2073 6009
rect 2091 5997 2094 6009
rect 2107 5997 2110 6009
rect 2126 6003 2138 6006
rect 2149 5997 2152 6009
rect 2165 5997 2168 6009
rect 2186 5997 2189 6009
rect 2202 5997 2205 6009
rect 2223 5997 2226 6009
rect 2239 5997 2242 6009
rect 2258 6003 2270 6006
rect 2281 5997 2284 6009
rect 2297 5997 2300 6009
rect 2318 5997 2321 6009
rect 2565 6010 2587 6013
rect 2591 6010 2598 6013
rect 2623 6010 2647 6013
rect 2651 6010 2656 6013
rect 2669 6012 2678 6016
rect 4786 6006 4829 6016
rect 1862 5983 1881 5986
rect 1885 5987 1892 5990
rect 1403 5978 1615 5982
rect 1619 5978 1682 5982
rect 1686 5978 1718 5982
rect 1722 5978 1731 5982
rect 1817 5977 1839 5980
rect 1843 5977 1850 5980
rect 1875 5977 1899 5980
rect 1903 5977 1908 5980
rect 1938 5983 1955 5986
rect 1959 5987 1966 5990
rect 1991 5987 1994 5993
rect 1994 5983 2013 5986
rect 2017 5987 2024 5990
rect 1949 5977 1971 5980
rect 1975 5977 1982 5980
rect 2007 5977 2031 5980
rect 2035 5977 2040 5980
rect 2070 5983 2087 5986
rect 2091 5987 2098 5990
rect 2123 5987 2126 5993
rect 2126 5983 2145 5986
rect 2149 5987 2156 5990
rect 2081 5977 2103 5980
rect 2107 5977 2114 5980
rect 2139 5977 2163 5980
rect 2167 5977 2172 5980
rect 2202 5983 2219 5986
rect 2223 5987 2230 5990
rect 2255 5987 2258 5993
rect 2258 5983 2277 5986
rect 2281 5987 2288 5990
rect 2554 5989 2557 5999
rect 2575 5989 2578 5999
rect 2591 5989 2594 5999
rect 2606 5992 2613 5996
rect 2617 5992 2622 5996
rect 2633 5989 2636 5999
rect 2649 5989 2652 5999
rect 2670 5989 2673 5999
rect 4796 5996 4829 6006
rect 2408 5985 2544 5989
rect 2548 5985 2581 5989
rect 2585 5985 2611 5989
rect 2615 5985 2639 5989
rect 2643 5985 2676 5989
rect 4806 5986 4829 5996
rect 2213 5977 2235 5980
rect 2239 5977 2246 5980
rect 2271 5977 2295 5980
rect 2299 5977 2304 5980
rect 2348 5978 2560 5982
rect 2564 5978 2627 5982
rect 2631 5978 2663 5982
rect 2667 5978 2676 5982
rect 4816 5976 4829 5986
rect 343 5925 346 5964
rect 861 5956 864 5966
rect 882 5956 885 5966
rect 898 5956 901 5966
rect 913 5959 920 5963
rect 924 5959 929 5963
rect 940 5956 943 5966
rect 956 5956 959 5966
rect 977 5956 980 5966
rect 993 5956 996 5966
rect 1014 5956 1017 5966
rect 1030 5956 1033 5966
rect 1045 5959 1052 5963
rect 1056 5959 1061 5963
rect 1072 5956 1075 5966
rect 1088 5956 1091 5966
rect 1109 5956 1112 5966
rect 1125 5956 1128 5966
rect 1146 5956 1149 5966
rect 1162 5956 1165 5966
rect 1177 5959 1184 5963
rect 1188 5959 1193 5963
rect 1204 5956 1207 5966
rect 1220 5956 1223 5966
rect 1241 5956 1244 5966
rect 1257 5956 1260 5966
rect 1278 5956 1281 5966
rect 1294 5956 1297 5966
rect 1309 5959 1316 5963
rect 1320 5959 1325 5963
rect 1336 5956 1339 5966
rect 1352 5956 1355 5966
rect 1373 5956 1376 5966
rect 1806 5956 1809 5966
rect 1827 5956 1830 5966
rect 1843 5956 1846 5966
rect 1858 5959 1865 5963
rect 1869 5959 1874 5963
rect 1885 5956 1888 5966
rect 1901 5956 1904 5966
rect 1922 5956 1925 5966
rect 1938 5956 1941 5966
rect 1959 5956 1962 5966
rect 1975 5956 1978 5966
rect 1990 5959 1997 5963
rect 2001 5959 2006 5963
rect 2017 5956 2020 5966
rect 2033 5956 2036 5966
rect 2054 5956 2057 5966
rect 2070 5956 2073 5966
rect 2091 5956 2094 5966
rect 2107 5956 2110 5966
rect 2122 5959 2129 5963
rect 2133 5959 2138 5963
rect 2149 5956 2152 5966
rect 2165 5956 2168 5966
rect 2186 5956 2189 5966
rect 2202 5956 2205 5966
rect 2223 5956 2226 5966
rect 2239 5956 2242 5966
rect 2254 5959 2261 5963
rect 2265 5959 2270 5963
rect 2281 5956 2284 5966
rect 2297 5956 2300 5966
rect 2318 5956 2321 5966
rect 855 5952 888 5956
rect 892 5952 918 5956
rect 922 5952 946 5956
rect 950 5952 983 5956
rect 987 5952 1020 5956
rect 1024 5952 1050 5956
rect 1054 5952 1078 5956
rect 1082 5952 1115 5956
rect 1119 5952 1152 5956
rect 1156 5952 1182 5956
rect 1186 5952 1210 5956
rect 1214 5952 1247 5956
rect 1251 5952 1284 5956
rect 1288 5952 1314 5956
rect 1318 5952 1342 5956
rect 1346 5952 1457 5956
rect 1800 5952 1833 5956
rect 1837 5952 1863 5956
rect 1867 5952 1891 5956
rect 1895 5952 1928 5956
rect 1932 5952 1965 5956
rect 1969 5952 1995 5956
rect 1999 5952 2023 5956
rect 2027 5952 2060 5956
rect 2064 5952 2097 5956
rect 2101 5952 2127 5956
rect 2131 5952 2155 5956
rect 2159 5952 2192 5956
rect 2196 5952 2229 5956
rect 2233 5952 2259 5956
rect 2263 5952 2287 5956
rect 2291 5952 2402 5956
rect 851 5945 867 5949
rect 871 5945 934 5949
rect 938 5945 970 5949
rect 974 5945 999 5949
rect 1003 5945 1066 5949
rect 1070 5945 1102 5949
rect 1106 5945 1131 5949
rect 1135 5945 1198 5949
rect 1202 5945 1234 5949
rect 1238 5945 1263 5949
rect 1267 5945 1330 5949
rect 1334 5945 1366 5949
rect 1370 5945 1397 5949
rect 1796 5945 1812 5949
rect 1816 5945 1879 5949
rect 1883 5945 1915 5949
rect 1919 5945 1944 5949
rect 1948 5945 2011 5949
rect 2015 5945 2047 5949
rect 2051 5945 2076 5949
rect 2080 5945 2143 5949
rect 2147 5945 2179 5949
rect 2183 5945 2208 5949
rect 2212 5945 2275 5949
rect 2279 5945 2311 5949
rect 2315 5945 2342 5949
rect 1415 5937 1485 5941
rect 1489 5937 1535 5941
rect 1539 5937 1586 5941
rect 1590 5937 1617 5941
rect 1621 5937 1667 5941
rect 1671 5937 1718 5941
rect 1722 5937 1749 5941
rect 1753 5937 1799 5941
rect 1803 5937 1850 5941
rect 1854 5937 1863 5941
rect 2360 5937 2430 5941
rect 2434 5937 2480 5941
rect 2484 5937 2531 5941
rect 2535 5937 2562 5941
rect 2566 5937 2612 5941
rect 2616 5937 2663 5941
rect 2667 5937 2694 5941
rect 2698 5937 2744 5941
rect 2748 5937 2795 5941
rect 2799 5937 2808 5941
rect 4826 5937 4829 5976
rect 5083 5937 5086 6191
rect 1451 5930 1504 5934
rect 1508 5930 1534 5934
rect 1538 5930 1562 5934
rect 1566 5930 1636 5934
rect 1640 5930 1666 5934
rect 1670 5930 1694 5934
rect 1698 5930 1768 5934
rect 1772 5930 1798 5934
rect 1802 5930 1826 5934
rect 1830 5930 1863 5934
rect 2396 5930 2449 5934
rect 2453 5930 2479 5934
rect 2483 5930 2507 5934
rect 2511 5930 2581 5934
rect 2585 5930 2611 5934
rect 2615 5930 2639 5934
rect 2643 5930 2713 5934
rect 2717 5930 2743 5934
rect 2747 5930 2771 5934
rect 2775 5930 2808 5934
rect 4483 5931 4484 5935
rect 4488 5931 4489 5935
rect 4493 5931 4494 5935
rect 4498 5931 4499 5935
rect 4503 5931 4504 5935
rect 4508 5931 4509 5935
rect 4479 5930 4513 5931
rect 86 5922 346 5925
rect 1477 5918 1480 5930
rect 1498 5918 1501 5930
rect 1514 5918 1517 5930
rect 1533 5924 1545 5927
rect 1556 5918 1559 5930
rect 1572 5918 1575 5930
rect 1593 5918 1596 5930
rect 1609 5918 1612 5930
rect 1630 5918 1633 5930
rect 1646 5918 1649 5930
rect 1665 5924 1677 5927
rect 1688 5918 1691 5930
rect 1704 5918 1707 5930
rect 1725 5918 1728 5930
rect 1741 5918 1744 5930
rect 1762 5918 1765 5930
rect 1778 5918 1781 5930
rect 1797 5924 1809 5927
rect 1820 5918 1823 5930
rect 1836 5918 1839 5930
rect 1857 5918 1860 5930
rect 2422 5918 2425 5930
rect 2443 5918 2446 5930
rect 2459 5918 2462 5930
rect 2478 5924 2490 5927
rect 2501 5918 2504 5930
rect 2517 5918 2520 5930
rect 2538 5918 2541 5930
rect 2554 5918 2557 5930
rect 2575 5918 2578 5930
rect 2591 5918 2594 5930
rect 2610 5924 2622 5927
rect 2633 5918 2636 5930
rect 2649 5918 2652 5930
rect 2670 5918 2673 5930
rect 2686 5918 2689 5930
rect 2707 5918 2710 5930
rect 2723 5918 2726 5930
rect 2742 5924 2754 5927
rect 2765 5918 2768 5930
rect 2781 5918 2784 5930
rect 2802 5918 2805 5930
rect 1477 5904 1494 5907
rect 1498 5908 1505 5911
rect 1530 5908 1533 5914
rect 1533 5904 1552 5907
rect 1556 5908 1563 5911
rect 1611 5904 1626 5907
rect 1630 5908 1637 5911
rect 1662 5908 1665 5914
rect 1665 5904 1684 5907
rect 1688 5908 1695 5911
rect 1743 5904 1758 5907
rect 1762 5908 1769 5911
rect 1794 5908 1797 5914
rect 1797 5904 1816 5907
rect 1820 5908 1827 5911
rect 1488 5898 1510 5901
rect 1514 5898 1521 5901
rect 617 5887 618 5891
rect 622 5887 623 5891
rect 627 5887 628 5891
rect 632 5887 633 5891
rect 637 5887 638 5891
rect 642 5887 643 5891
rect 613 5886 647 5887
rect 617 5882 618 5886
rect 622 5882 623 5886
rect 627 5882 628 5886
rect 632 5882 633 5886
rect 637 5882 638 5886
rect 642 5882 643 5886
rect 613 5881 647 5882
rect 617 5877 618 5881
rect 622 5877 623 5881
rect 627 5877 628 5881
rect 632 5877 633 5881
rect 637 5877 638 5881
rect 642 5877 643 5881
rect 613 5876 647 5877
rect 86 5870 346 5873
rect 617 5872 618 5876
rect 622 5872 623 5876
rect 627 5872 628 5876
rect 632 5872 633 5876
rect 637 5872 638 5876
rect 642 5872 643 5876
rect 663 5887 664 5891
rect 668 5887 669 5891
rect 673 5887 674 5891
rect 678 5887 679 5891
rect 683 5887 684 5891
rect 688 5887 689 5891
rect 1546 5898 1570 5901
rect 1574 5898 1579 5901
rect 1593 5898 1600 5901
rect 1620 5898 1642 5901
rect 1646 5898 1653 5901
rect 1678 5898 1702 5901
rect 1706 5898 1711 5901
rect 1725 5898 1732 5901
rect 1752 5898 1774 5901
rect 1778 5898 1785 5901
rect 1810 5898 1834 5901
rect 1838 5898 1843 5901
rect 2422 5904 2439 5907
rect 2443 5908 2450 5911
rect 2475 5908 2478 5914
rect 2478 5904 2497 5907
rect 2501 5908 2508 5911
rect 2556 5904 2571 5907
rect 2575 5908 2582 5911
rect 2607 5908 2610 5914
rect 2610 5904 2629 5907
rect 2633 5908 2640 5911
rect 2688 5904 2703 5907
rect 2707 5908 2714 5911
rect 2739 5908 2742 5914
rect 4483 5926 4484 5930
rect 4488 5926 4489 5930
rect 4493 5926 4494 5930
rect 4498 5926 4499 5930
rect 4503 5926 4504 5930
rect 4508 5926 4509 5930
rect 4479 5925 4513 5926
rect 4483 5921 4484 5925
rect 4488 5921 4489 5925
rect 4493 5921 4494 5925
rect 4498 5921 4499 5925
rect 4503 5921 4504 5925
rect 4508 5921 4509 5925
rect 4479 5920 4513 5921
rect 4483 5916 4484 5920
rect 4488 5916 4489 5920
rect 4493 5916 4494 5920
rect 4498 5916 4499 5920
rect 4503 5916 4504 5920
rect 4508 5916 4509 5920
rect 4529 5931 4530 5935
rect 4534 5931 4535 5935
rect 4539 5931 4540 5935
rect 4544 5931 4545 5935
rect 4549 5931 4550 5935
rect 4554 5931 4555 5935
rect 4826 5934 5086 5937
rect 4525 5930 4559 5931
rect 4529 5926 4530 5930
rect 4534 5926 4535 5930
rect 4539 5926 4540 5930
rect 4544 5926 4545 5930
rect 4549 5926 4550 5930
rect 4554 5926 4555 5930
rect 4525 5925 4559 5926
rect 4529 5921 4530 5925
rect 4534 5921 4535 5925
rect 4539 5921 4540 5925
rect 4544 5921 4545 5925
rect 4549 5921 4550 5925
rect 4554 5921 4555 5925
rect 4525 5920 4559 5921
rect 4529 5916 4530 5920
rect 4534 5916 4535 5920
rect 4539 5916 4540 5920
rect 4544 5916 4545 5920
rect 4549 5916 4550 5920
rect 4554 5916 4555 5920
rect 2742 5904 2761 5907
rect 2765 5908 2772 5911
rect 2433 5898 2455 5901
rect 2459 5898 2466 5901
rect 2491 5898 2515 5901
rect 2519 5898 2524 5901
rect 2538 5898 2545 5901
rect 2565 5898 2587 5901
rect 2591 5898 2598 5901
rect 2623 5898 2647 5901
rect 2651 5898 2656 5901
rect 2670 5898 2677 5901
rect 2697 5898 2719 5901
rect 2723 5898 2730 5901
rect 2755 5898 2779 5901
rect 2783 5898 2788 5901
rect 659 5886 693 5887
rect 663 5882 664 5886
rect 668 5882 669 5886
rect 673 5882 674 5886
rect 678 5882 679 5886
rect 683 5882 684 5886
rect 688 5882 689 5886
rect 659 5881 693 5882
rect 663 5877 664 5881
rect 668 5877 669 5881
rect 673 5877 674 5881
rect 678 5877 679 5881
rect 683 5877 684 5881
rect 688 5877 689 5881
rect 1477 5877 1480 5887
rect 1498 5877 1501 5887
rect 1514 5877 1517 5887
rect 1529 5880 1536 5884
rect 1540 5880 1545 5884
rect 1556 5877 1559 5887
rect 1572 5877 1575 5887
rect 1593 5877 1596 5887
rect 1609 5877 1612 5887
rect 1630 5877 1633 5887
rect 1646 5877 1649 5887
rect 1661 5880 1668 5884
rect 1672 5880 1677 5884
rect 1688 5877 1691 5887
rect 1704 5877 1707 5887
rect 1725 5877 1728 5887
rect 1741 5877 1744 5887
rect 1762 5877 1765 5887
rect 1778 5877 1781 5887
rect 1793 5880 1800 5884
rect 1804 5880 1809 5884
rect 1820 5877 1823 5887
rect 1836 5877 1839 5887
rect 1857 5877 1860 5887
rect 2422 5877 2425 5887
rect 2443 5877 2446 5887
rect 2459 5877 2462 5887
rect 2474 5880 2481 5884
rect 2485 5880 2490 5884
rect 2501 5877 2504 5887
rect 2517 5877 2520 5887
rect 2538 5877 2541 5887
rect 2554 5877 2557 5887
rect 2575 5877 2578 5887
rect 2591 5877 2594 5887
rect 2606 5880 2613 5884
rect 2617 5880 2622 5884
rect 2633 5877 2636 5887
rect 2649 5877 2652 5887
rect 2670 5877 2673 5887
rect 2686 5877 2689 5887
rect 2707 5877 2710 5887
rect 2723 5877 2726 5887
rect 2738 5880 2745 5884
rect 2749 5880 2754 5884
rect 2765 5877 2768 5887
rect 2781 5877 2784 5887
rect 2802 5877 2805 5887
rect 4826 5882 5086 5885
rect 659 5876 693 5877
rect 663 5872 664 5876
rect 668 5872 669 5876
rect 673 5872 674 5876
rect 678 5872 679 5876
rect 683 5872 684 5876
rect 688 5872 689 5876
rect 1463 5873 1467 5877
rect 1471 5873 1504 5877
rect 1508 5873 1534 5877
rect 1538 5873 1562 5877
rect 1566 5873 1599 5877
rect 1603 5873 1636 5877
rect 1640 5873 1666 5877
rect 1670 5873 1694 5877
rect 1698 5873 1731 5877
rect 1735 5873 1768 5877
rect 1772 5873 1798 5877
rect 1802 5873 1826 5877
rect 1830 5873 1863 5877
rect 2408 5873 2412 5877
rect 2416 5873 2449 5877
rect 2453 5873 2479 5877
rect 2483 5873 2507 5877
rect 2511 5873 2544 5877
rect 2548 5873 2581 5877
rect 2585 5873 2611 5877
rect 2615 5873 2639 5877
rect 2643 5873 2676 5877
rect 2680 5873 2713 5877
rect 2717 5873 2743 5877
rect 2747 5873 2771 5877
rect 2775 5873 2808 5877
rect 86 5616 89 5870
rect 343 5831 346 5870
rect 1403 5866 1483 5870
rect 1487 5866 1550 5870
rect 1554 5866 1586 5870
rect 1590 5866 1615 5870
rect 1619 5866 1682 5870
rect 1686 5866 1718 5870
rect 1722 5866 1747 5870
rect 1751 5866 1814 5870
rect 1818 5866 1850 5870
rect 1854 5866 1863 5870
rect 2348 5866 2428 5870
rect 2432 5866 2495 5870
rect 2499 5866 2531 5870
rect 2535 5866 2560 5870
rect 2564 5866 2627 5870
rect 2631 5866 2663 5870
rect 2667 5866 2692 5870
rect 2696 5866 2759 5870
rect 2763 5866 2795 5870
rect 2799 5866 2808 5870
rect 1628 5860 1732 5863
rect 2573 5860 2677 5863
rect 1604 5852 1608 5856
rect 1612 5852 1616 5856
rect 2549 5852 2553 5856
rect 2557 5852 2561 5856
rect 1472 5844 1585 5847
rect 2417 5844 2530 5847
rect 4826 5843 4829 5882
rect 1472 5837 1600 5840
rect 2417 5837 2545 5840
rect 4816 5833 4829 5843
rect 343 5821 356 5831
rect 849 5829 927 5833
rect 931 5829 1592 5833
rect 1608 5829 1624 5833
rect 1628 5829 1872 5833
rect 1876 5829 2537 5833
rect 2553 5829 2569 5833
rect 2573 5829 2818 5833
rect 343 5811 366 5821
rect 1604 5818 1608 5822
rect 1612 5818 1616 5822
rect 4806 5823 4829 5833
rect 2549 5818 2553 5822
rect 2557 5818 2561 5822
rect 1628 5811 1732 5814
rect 2573 5811 2677 5814
rect 4796 5813 4829 5823
rect 343 5801 376 5811
rect 1472 5804 1857 5807
rect 2417 5804 2802 5807
rect 4786 5803 4829 5813
rect 343 5791 386 5801
rect 1415 5797 1485 5801
rect 1489 5797 1535 5801
rect 1539 5797 1586 5801
rect 1590 5797 1617 5801
rect 1621 5797 1667 5801
rect 1671 5797 1718 5801
rect 1722 5797 1749 5801
rect 1753 5797 1799 5801
rect 1803 5797 1850 5801
rect 1854 5797 1863 5801
rect 2360 5797 2430 5801
rect 2434 5797 2480 5801
rect 2484 5797 2531 5801
rect 2535 5797 2562 5801
rect 2566 5797 2612 5801
rect 2616 5797 2663 5801
rect 2667 5797 2694 5801
rect 2698 5797 2744 5801
rect 2748 5797 2795 5801
rect 2799 5797 2808 5801
rect 343 5695 769 5791
rect 1451 5790 1504 5794
rect 1508 5790 1534 5794
rect 1538 5790 1562 5794
rect 1566 5790 1636 5794
rect 1640 5790 1666 5794
rect 1670 5790 1694 5794
rect 1698 5790 1768 5794
rect 1772 5790 1798 5794
rect 1802 5790 1826 5794
rect 1830 5790 1863 5794
rect 2396 5790 2449 5794
rect 2453 5790 2479 5794
rect 2483 5790 2507 5794
rect 2511 5790 2581 5794
rect 2585 5790 2611 5794
rect 2615 5790 2639 5794
rect 2643 5790 2713 5794
rect 2717 5790 2743 5794
rect 2747 5790 2771 5794
rect 2775 5790 2808 5794
rect 1477 5778 1480 5790
rect 1498 5778 1501 5790
rect 1514 5778 1517 5790
rect 1533 5784 1545 5787
rect 1556 5778 1559 5790
rect 1572 5778 1575 5790
rect 1593 5778 1596 5790
rect 1609 5778 1612 5790
rect 1630 5778 1633 5790
rect 1646 5778 1649 5790
rect 1665 5784 1677 5787
rect 1688 5778 1691 5790
rect 1704 5778 1707 5790
rect 1725 5778 1728 5790
rect 1741 5778 1744 5790
rect 1762 5778 1765 5790
rect 1778 5778 1781 5790
rect 1797 5784 1809 5787
rect 1820 5778 1823 5790
rect 1836 5778 1839 5790
rect 1857 5778 1860 5790
rect 2422 5778 2425 5790
rect 2443 5778 2446 5790
rect 2459 5778 2462 5790
rect 2478 5784 2490 5787
rect 2501 5778 2504 5790
rect 2517 5778 2520 5790
rect 2538 5778 2541 5790
rect 2554 5778 2557 5790
rect 2575 5778 2578 5790
rect 2591 5778 2594 5790
rect 2610 5784 2622 5787
rect 2633 5778 2636 5790
rect 2649 5778 2652 5790
rect 2670 5778 2673 5790
rect 2686 5778 2689 5790
rect 2707 5778 2710 5790
rect 2723 5778 2726 5790
rect 2742 5784 2754 5787
rect 2765 5778 2768 5790
rect 2781 5778 2784 5790
rect 2802 5778 2805 5790
rect 948 5767 966 5771
rect 970 5767 1016 5771
rect 1020 5767 1067 5771
rect 1071 5767 1409 5771
rect 948 5760 985 5764
rect 989 5760 1015 5764
rect 1019 5760 1043 5764
rect 1047 5760 1445 5764
rect 1477 5764 1494 5767
rect 1498 5768 1505 5771
rect 1530 5768 1533 5774
rect 1533 5764 1552 5767
rect 1556 5768 1563 5771
rect 1611 5764 1626 5767
rect 1630 5768 1637 5771
rect 1662 5768 1665 5774
rect 1665 5764 1684 5767
rect 1688 5768 1695 5771
rect 1743 5764 1758 5767
rect 1762 5768 1769 5771
rect 1794 5768 1797 5774
rect 1797 5764 1816 5767
rect 1820 5768 1827 5771
rect 1893 5767 1911 5771
rect 1915 5767 1961 5771
rect 1965 5767 2012 5771
rect 2016 5767 2354 5771
rect 958 5748 961 5760
rect 979 5748 982 5760
rect 995 5748 998 5760
rect 1014 5754 1026 5757
rect 1037 5748 1040 5760
rect 1053 5748 1056 5760
rect 1074 5748 1077 5760
rect 938 5735 949 5739
rect 960 5734 975 5737
rect 979 5738 986 5741
rect 1011 5738 1014 5744
rect 1488 5758 1510 5761
rect 1514 5758 1521 5761
rect 1546 5758 1570 5761
rect 1574 5758 1579 5761
rect 1593 5758 1600 5761
rect 1620 5758 1642 5761
rect 1646 5758 1653 5761
rect 1678 5758 1702 5761
rect 1706 5758 1711 5761
rect 1725 5758 1732 5761
rect 1752 5758 1774 5761
rect 1778 5758 1785 5761
rect 1810 5758 1834 5761
rect 1838 5758 1843 5761
rect 1893 5760 1930 5764
rect 1934 5760 1960 5764
rect 1964 5760 1988 5764
rect 1992 5760 2390 5764
rect 2422 5764 2439 5767
rect 2443 5768 2450 5771
rect 2475 5768 2478 5774
rect 2478 5764 2497 5767
rect 2501 5768 2508 5771
rect 2556 5764 2571 5767
rect 2575 5768 2582 5771
rect 2607 5768 2610 5774
rect 2610 5764 2629 5767
rect 2633 5768 2640 5771
rect 2688 5764 2703 5767
rect 2707 5768 2714 5771
rect 2739 5768 2742 5774
rect 2742 5764 2761 5767
rect 2765 5768 2772 5771
rect 1903 5748 1906 5760
rect 1924 5748 1927 5760
rect 1940 5748 1943 5760
rect 1959 5754 1971 5757
rect 1982 5748 1985 5760
rect 1998 5748 2001 5760
rect 2019 5748 2022 5760
rect 1014 5734 1033 5737
rect 1037 5738 1044 5741
rect 1477 5737 1480 5747
rect 1498 5737 1501 5747
rect 1514 5737 1517 5747
rect 1529 5740 1536 5744
rect 1540 5740 1545 5744
rect 1556 5737 1559 5747
rect 1572 5737 1575 5747
rect 1593 5737 1596 5747
rect 1609 5737 1612 5747
rect 1630 5737 1633 5747
rect 1646 5737 1649 5747
rect 1661 5740 1668 5744
rect 1672 5740 1677 5744
rect 1688 5737 1691 5747
rect 1704 5737 1707 5747
rect 1725 5737 1728 5747
rect 1741 5737 1744 5747
rect 1762 5737 1765 5747
rect 1778 5737 1781 5747
rect 1793 5740 1800 5744
rect 1804 5740 1809 5744
rect 1820 5737 1823 5747
rect 1836 5737 1839 5747
rect 1857 5737 1860 5747
rect 969 5728 991 5731
rect 995 5728 1002 5731
rect 1027 5728 1051 5731
rect 1055 5728 1060 5731
rect 1463 5733 1467 5737
rect 1471 5733 1504 5737
rect 1508 5733 1534 5737
rect 1538 5733 1562 5737
rect 1566 5733 1599 5737
rect 1603 5733 1636 5737
rect 1640 5733 1666 5737
rect 1670 5733 1694 5737
rect 1698 5733 1731 5737
rect 1735 5733 1768 5737
rect 1772 5733 1798 5737
rect 1802 5733 1826 5737
rect 1830 5733 1863 5737
rect 1883 5735 1894 5739
rect 1905 5734 1920 5737
rect 1924 5738 1931 5741
rect 1956 5738 1959 5744
rect 2433 5758 2455 5761
rect 2459 5758 2466 5761
rect 2491 5758 2515 5761
rect 2519 5758 2524 5761
rect 2538 5758 2545 5761
rect 2565 5758 2587 5761
rect 2591 5758 2598 5761
rect 2623 5758 2647 5761
rect 2651 5758 2656 5761
rect 2670 5758 2677 5761
rect 2697 5758 2719 5761
rect 2723 5758 2730 5761
rect 2755 5758 2779 5761
rect 2783 5758 2788 5761
rect 1959 5734 1978 5737
rect 1982 5738 1989 5741
rect 2422 5737 2425 5747
rect 2443 5737 2446 5747
rect 2459 5737 2462 5747
rect 2474 5740 2481 5744
rect 2485 5740 2490 5744
rect 2501 5737 2504 5747
rect 2517 5737 2520 5747
rect 2538 5737 2541 5747
rect 2554 5737 2557 5747
rect 2575 5737 2578 5747
rect 2591 5737 2594 5747
rect 2606 5740 2613 5744
rect 2617 5740 2622 5744
rect 2633 5737 2636 5747
rect 2649 5737 2652 5747
rect 2670 5737 2673 5747
rect 2686 5737 2689 5747
rect 2707 5737 2710 5747
rect 2723 5737 2726 5747
rect 2738 5740 2745 5744
rect 2749 5740 2754 5744
rect 2765 5737 2768 5747
rect 2781 5737 2784 5747
rect 2802 5737 2805 5747
rect 1403 5726 1483 5730
rect 1487 5726 1550 5730
rect 1554 5726 1586 5730
rect 1590 5726 1615 5730
rect 1619 5726 1682 5730
rect 1686 5726 1718 5730
rect 1722 5726 1747 5730
rect 1751 5726 1814 5730
rect 1818 5726 1850 5730
rect 1854 5726 1863 5730
rect 1914 5728 1936 5731
rect 1940 5728 1947 5731
rect 1472 5719 1857 5722
rect 1972 5728 1996 5731
rect 2000 5728 2005 5731
rect 2408 5733 2412 5737
rect 2416 5733 2449 5737
rect 2453 5733 2479 5737
rect 2483 5733 2507 5737
rect 2511 5733 2544 5737
rect 2548 5733 2581 5737
rect 2585 5733 2611 5737
rect 2615 5733 2639 5737
rect 2643 5733 2676 5737
rect 2680 5733 2713 5737
rect 2717 5733 2743 5737
rect 2747 5733 2771 5737
rect 2775 5733 2808 5737
rect 2348 5726 2428 5730
rect 2432 5726 2495 5730
rect 2499 5726 2531 5730
rect 2535 5726 2560 5730
rect 2564 5726 2627 5730
rect 2631 5726 2663 5730
rect 2667 5726 2692 5730
rect 2696 5726 2759 5730
rect 2763 5726 2795 5730
rect 2799 5726 2808 5730
rect 2417 5719 2802 5722
rect 958 5707 961 5717
rect 979 5707 982 5717
rect 995 5707 998 5717
rect 1010 5710 1017 5714
rect 1021 5710 1026 5714
rect 1037 5707 1040 5717
rect 1053 5707 1056 5717
rect 1074 5707 1077 5717
rect 1415 5711 1485 5715
rect 1489 5711 1535 5715
rect 1539 5711 1586 5715
rect 1590 5711 1617 5715
rect 1621 5711 1667 5715
rect 1671 5711 1718 5715
rect 1722 5711 1749 5715
rect 1753 5711 1799 5715
rect 1803 5711 1850 5715
rect 1854 5711 1863 5715
rect 952 5703 985 5707
rect 989 5703 1015 5707
rect 1019 5703 1043 5707
rect 1047 5703 1081 5707
rect 1451 5704 1504 5708
rect 1508 5704 1534 5708
rect 1538 5704 1562 5708
rect 1566 5704 1636 5708
rect 1640 5704 1666 5708
rect 1670 5704 1694 5708
rect 1698 5704 1768 5708
rect 1772 5704 1798 5708
rect 1802 5704 1826 5708
rect 1830 5704 1863 5708
rect 1903 5707 1906 5717
rect 1924 5707 1927 5717
rect 1940 5707 1943 5717
rect 1955 5710 1962 5714
rect 1966 5710 1971 5714
rect 1982 5707 1985 5717
rect 1998 5707 2001 5717
rect 2019 5707 2022 5717
rect 2360 5711 2430 5715
rect 2434 5711 2480 5715
rect 2484 5711 2531 5715
rect 2535 5711 2562 5715
rect 2566 5711 2612 5715
rect 2616 5711 2663 5715
rect 2667 5711 2694 5715
rect 2698 5711 2744 5715
rect 2748 5711 2795 5715
rect 2799 5711 2808 5715
rect 948 5696 964 5700
rect 968 5696 1031 5700
rect 1035 5696 1067 5700
rect 1071 5696 1397 5700
rect 343 5685 386 5695
rect 953 5689 1074 5692
rect 1477 5692 1480 5704
rect 1498 5692 1501 5704
rect 1514 5692 1517 5704
rect 1533 5698 1545 5701
rect 1556 5692 1559 5704
rect 1572 5692 1575 5704
rect 1593 5692 1596 5704
rect 1609 5692 1612 5704
rect 1630 5692 1633 5704
rect 1646 5692 1649 5704
rect 1665 5698 1677 5701
rect 1688 5692 1691 5704
rect 1704 5692 1707 5704
rect 1725 5692 1728 5704
rect 1741 5692 1744 5704
rect 1762 5692 1765 5704
rect 1778 5692 1781 5704
rect 1797 5698 1809 5701
rect 1820 5692 1823 5704
rect 1836 5692 1839 5704
rect 1857 5692 1860 5704
rect 1897 5703 1930 5707
rect 1934 5703 1960 5707
rect 1964 5703 1988 5707
rect 1992 5703 2026 5707
rect 2396 5704 2449 5708
rect 2453 5704 2479 5708
rect 2483 5704 2507 5708
rect 2511 5704 2581 5708
rect 2585 5704 2611 5708
rect 2615 5704 2639 5708
rect 2643 5704 2713 5708
rect 2717 5704 2743 5708
rect 2747 5704 2771 5708
rect 2775 5704 2808 5708
rect 4403 5707 4829 5803
rect 1893 5696 1909 5700
rect 1913 5696 1976 5700
rect 1980 5696 2012 5700
rect 2016 5696 2342 5700
rect 343 5675 376 5685
rect 948 5681 966 5685
rect 970 5681 1016 5685
rect 1020 5681 1067 5685
rect 1071 5681 1409 5685
rect 343 5665 366 5675
rect 948 5674 985 5678
rect 989 5674 1015 5678
rect 1019 5674 1043 5678
rect 1047 5674 1445 5678
rect 1477 5678 1494 5681
rect 1498 5682 1505 5685
rect 1530 5682 1533 5688
rect 1533 5678 1552 5681
rect 1556 5682 1563 5685
rect 1611 5678 1626 5681
rect 1630 5682 1637 5685
rect 1662 5682 1665 5688
rect 1665 5678 1684 5681
rect 1688 5682 1695 5685
rect 1743 5678 1758 5681
rect 1762 5682 1769 5685
rect 1794 5682 1797 5688
rect 1898 5689 2019 5692
rect 2422 5692 2425 5704
rect 2443 5692 2446 5704
rect 2459 5692 2462 5704
rect 2478 5698 2490 5701
rect 2501 5692 2504 5704
rect 2517 5692 2520 5704
rect 2538 5692 2541 5704
rect 2554 5692 2557 5704
rect 2575 5692 2578 5704
rect 2591 5692 2594 5704
rect 2610 5698 2622 5701
rect 2633 5692 2636 5704
rect 2649 5692 2652 5704
rect 2670 5692 2673 5704
rect 2686 5692 2689 5704
rect 2707 5692 2710 5704
rect 2723 5692 2726 5704
rect 2742 5698 2754 5701
rect 2765 5692 2768 5704
rect 2781 5692 2784 5704
rect 2802 5692 2805 5704
rect 4786 5697 4829 5707
rect 1797 5678 1816 5681
rect 1820 5682 1827 5685
rect 1893 5681 1911 5685
rect 1915 5681 1961 5685
rect 1965 5681 2012 5685
rect 2016 5681 2354 5685
rect 343 5655 356 5665
rect 958 5662 961 5674
rect 979 5662 982 5674
rect 995 5662 998 5674
rect 1014 5668 1026 5671
rect 1037 5662 1040 5674
rect 1053 5662 1056 5674
rect 1074 5662 1077 5674
rect 343 5616 346 5655
rect 960 5648 975 5651
rect 979 5652 986 5655
rect 1011 5652 1014 5658
rect 1488 5672 1510 5675
rect 1514 5672 1521 5675
rect 1546 5672 1570 5675
rect 1574 5672 1579 5675
rect 1593 5672 1600 5675
rect 1620 5672 1642 5675
rect 1646 5672 1653 5675
rect 1678 5672 1702 5675
rect 1706 5672 1711 5675
rect 1725 5672 1732 5675
rect 1752 5672 1774 5675
rect 1778 5672 1785 5675
rect 1810 5672 1834 5675
rect 1838 5672 1843 5675
rect 1893 5674 1930 5678
rect 1934 5674 1960 5678
rect 1964 5674 1988 5678
rect 1992 5674 2390 5678
rect 2422 5678 2439 5681
rect 2443 5682 2450 5685
rect 2475 5682 2478 5688
rect 2478 5678 2497 5681
rect 2501 5682 2508 5685
rect 2556 5678 2571 5681
rect 2575 5682 2582 5685
rect 2607 5682 2610 5688
rect 2610 5678 2629 5681
rect 2633 5682 2640 5685
rect 2688 5678 2703 5681
rect 2707 5682 2714 5685
rect 2739 5682 2742 5688
rect 2742 5678 2761 5681
rect 2765 5682 2772 5685
rect 4796 5687 4829 5697
rect 1903 5662 1906 5674
rect 1924 5662 1927 5674
rect 1940 5662 1943 5674
rect 1959 5668 1971 5671
rect 1982 5662 1985 5674
rect 1998 5662 2001 5674
rect 2019 5662 2022 5674
rect 1014 5648 1033 5651
rect 1037 5652 1044 5655
rect 1477 5651 1480 5661
rect 1498 5651 1501 5661
rect 1514 5651 1517 5661
rect 1529 5654 1536 5658
rect 1540 5654 1545 5658
rect 1556 5651 1559 5661
rect 1572 5651 1575 5661
rect 1593 5651 1596 5661
rect 1609 5651 1612 5661
rect 1630 5651 1633 5661
rect 1646 5651 1649 5661
rect 1661 5654 1668 5658
rect 1672 5654 1677 5658
rect 1688 5651 1691 5661
rect 1704 5651 1707 5661
rect 1725 5651 1728 5661
rect 1741 5651 1744 5661
rect 1762 5651 1765 5661
rect 1778 5651 1781 5661
rect 1793 5654 1800 5658
rect 1804 5654 1809 5658
rect 1820 5651 1823 5661
rect 1836 5651 1839 5661
rect 1857 5651 1860 5661
rect 969 5642 991 5645
rect 995 5642 1002 5645
rect 1027 5642 1051 5645
rect 1055 5642 1060 5645
rect 1463 5647 1467 5651
rect 1471 5647 1504 5651
rect 1508 5647 1534 5651
rect 1538 5647 1562 5651
rect 1566 5647 1599 5651
rect 1603 5647 1636 5651
rect 1640 5647 1666 5651
rect 1670 5647 1694 5651
rect 1698 5647 1731 5651
rect 1735 5647 1768 5651
rect 1772 5647 1798 5651
rect 1802 5647 1826 5651
rect 1830 5647 1863 5651
rect 1905 5648 1920 5651
rect 1924 5652 1931 5655
rect 1956 5652 1959 5658
rect 2433 5672 2455 5675
rect 2459 5672 2466 5675
rect 2491 5672 2515 5675
rect 2519 5672 2524 5675
rect 2538 5672 2545 5675
rect 2565 5672 2587 5675
rect 2591 5672 2598 5675
rect 2623 5672 2647 5675
rect 2651 5672 2656 5675
rect 2670 5672 2677 5675
rect 2697 5672 2719 5675
rect 2723 5672 2730 5675
rect 2755 5672 2779 5675
rect 2783 5672 2788 5675
rect 4806 5677 4829 5687
rect 4816 5667 4829 5677
rect 1959 5648 1978 5651
rect 1982 5652 1989 5655
rect 2422 5651 2425 5661
rect 2443 5651 2446 5661
rect 2459 5651 2462 5661
rect 2474 5654 2481 5658
rect 2485 5654 2490 5658
rect 2501 5651 2504 5661
rect 2517 5651 2520 5661
rect 2538 5651 2541 5661
rect 2554 5651 2557 5661
rect 2575 5651 2578 5661
rect 2591 5651 2594 5661
rect 2606 5654 2613 5658
rect 2617 5654 2622 5658
rect 2633 5651 2636 5661
rect 2649 5651 2652 5661
rect 2670 5651 2673 5661
rect 2686 5651 2689 5661
rect 2707 5651 2710 5661
rect 2723 5651 2726 5661
rect 2738 5654 2745 5658
rect 2749 5654 2754 5658
rect 2765 5651 2768 5661
rect 2781 5651 2784 5661
rect 2802 5651 2805 5661
rect 1403 5640 1483 5644
rect 1487 5640 1550 5644
rect 1554 5640 1586 5644
rect 1590 5640 1615 5644
rect 1619 5640 1682 5644
rect 1686 5640 1718 5644
rect 1722 5640 1747 5644
rect 1751 5640 1814 5644
rect 1818 5640 1850 5644
rect 1854 5640 1863 5644
rect 1914 5642 1936 5645
rect 1940 5642 1947 5645
rect 1603 5634 1713 5637
rect 1972 5642 1996 5645
rect 2000 5642 2005 5645
rect 2408 5647 2412 5651
rect 2416 5647 2449 5651
rect 2453 5647 2479 5651
rect 2483 5647 2507 5651
rect 2511 5647 2544 5651
rect 2548 5647 2581 5651
rect 2585 5647 2611 5651
rect 2615 5647 2639 5651
rect 2643 5647 2676 5651
rect 2680 5647 2713 5651
rect 2717 5647 2743 5651
rect 2747 5647 2771 5651
rect 2775 5647 2808 5651
rect 2348 5640 2428 5644
rect 2432 5640 2495 5644
rect 2499 5640 2531 5644
rect 2535 5640 2560 5644
rect 2564 5640 2627 5644
rect 2631 5640 2663 5644
rect 2667 5640 2692 5644
rect 2696 5640 2759 5644
rect 2763 5640 2795 5644
rect 2799 5640 2808 5644
rect 2548 5634 2658 5637
rect 958 5621 961 5631
rect 979 5621 982 5631
rect 995 5621 998 5631
rect 1010 5624 1017 5628
rect 1021 5624 1026 5628
rect 1037 5621 1040 5631
rect 1053 5621 1056 5631
rect 1074 5621 1077 5631
rect 1721 5626 1725 5630
rect 1729 5626 1733 5630
rect 952 5617 985 5621
rect 989 5617 1015 5621
rect 1019 5617 1043 5621
rect 1047 5617 1081 5621
rect 1085 5617 1457 5621
rect 1472 5618 1702 5621
rect 1903 5621 1906 5631
rect 1924 5621 1927 5631
rect 1940 5621 1943 5631
rect 1955 5624 1962 5628
rect 1966 5624 1971 5628
rect 1982 5621 1985 5631
rect 1998 5621 2001 5631
rect 2019 5621 2022 5631
rect 2666 5626 2670 5630
rect 2674 5626 2678 5630
rect 4826 5628 4829 5667
rect 5083 5628 5086 5882
rect 4483 5622 4484 5626
rect 4488 5622 4489 5626
rect 4493 5622 4494 5626
rect 4498 5622 4499 5626
rect 4503 5622 4504 5626
rect 4508 5622 4509 5626
rect 86 5613 346 5616
rect 1897 5617 1930 5621
rect 1934 5617 1960 5621
rect 1964 5617 1988 5621
rect 1992 5617 2026 5621
rect 2030 5617 2402 5621
rect 2417 5618 2647 5621
rect 4479 5621 4513 5622
rect 948 5610 964 5614
rect 968 5610 1031 5614
rect 1035 5610 1067 5614
rect 1071 5610 1397 5614
rect 1472 5611 1717 5614
rect 1893 5610 1909 5614
rect 1913 5610 1976 5614
rect 1980 5610 2012 5614
rect 2016 5610 2342 5614
rect 2417 5611 2662 5614
rect 4483 5617 4484 5621
rect 4488 5617 4489 5621
rect 4493 5617 4494 5621
rect 4498 5617 4499 5621
rect 4503 5617 4504 5621
rect 4508 5617 4509 5621
rect 4479 5616 4513 5617
rect 4483 5612 4484 5616
rect 4488 5612 4489 5616
rect 4493 5612 4494 5616
rect 4498 5612 4499 5616
rect 4503 5612 4504 5616
rect 4508 5612 4509 5616
rect 4479 5611 4513 5612
rect 4483 5607 4484 5611
rect 4488 5607 4489 5611
rect 4493 5607 4494 5611
rect 4498 5607 4499 5611
rect 4503 5607 4504 5611
rect 4508 5607 4509 5611
rect 4529 5622 4530 5626
rect 4534 5622 4535 5626
rect 4539 5622 4540 5626
rect 4544 5622 4545 5626
rect 4549 5622 4550 5626
rect 4554 5622 4555 5626
rect 4826 5625 5086 5628
rect 4525 5621 4559 5622
rect 4529 5617 4530 5621
rect 4534 5617 4535 5621
rect 4539 5617 4540 5621
rect 4544 5617 4545 5621
rect 4549 5617 4550 5621
rect 4554 5617 4555 5621
rect 4525 5616 4559 5617
rect 4529 5612 4530 5616
rect 4534 5612 4535 5616
rect 4539 5612 4540 5616
rect 4544 5612 4545 5616
rect 4549 5612 4550 5616
rect 4554 5612 4555 5616
rect 4525 5611 4559 5612
rect 4529 5607 4530 5611
rect 4534 5607 4535 5611
rect 4539 5607 4540 5611
rect 4544 5607 4545 5611
rect 4549 5607 4550 5611
rect 4554 5607 4555 5611
rect 851 5603 1709 5607
rect 1725 5603 1741 5607
rect 1745 5603 2654 5607
rect 2670 5603 2686 5607
rect 2690 5603 2817 5607
rect 939 5598 943 5603
rect 1114 5596 1385 5600
rect 1709 5594 1713 5595
rect 1741 5594 1745 5595
rect 1119 5590 1433 5593
rect 1721 5590 1725 5594
rect 1729 5590 1733 5594
rect 1884 5598 1888 5603
rect 2057 5597 2330 5600
rect 2654 5594 2658 5595
rect 2686 5594 2690 5595
rect 2064 5590 2378 5593
rect 2666 5590 2670 5594
rect 2674 5590 2678 5594
rect 617 5578 618 5582
rect 622 5578 623 5582
rect 627 5578 628 5582
rect 632 5578 633 5582
rect 637 5578 638 5582
rect 642 5578 643 5582
rect 613 5577 647 5578
rect 617 5573 618 5577
rect 622 5573 623 5577
rect 627 5573 628 5577
rect 632 5573 633 5577
rect 637 5573 638 5577
rect 642 5573 643 5577
rect 613 5572 647 5573
rect 617 5568 618 5572
rect 622 5568 623 5572
rect 627 5568 628 5572
rect 632 5568 633 5572
rect 637 5568 638 5572
rect 642 5568 643 5572
rect 613 5567 647 5568
rect 86 5561 346 5564
rect 617 5563 618 5567
rect 622 5563 623 5567
rect 627 5563 628 5567
rect 632 5563 633 5567
rect 637 5563 638 5567
rect 642 5563 643 5567
rect 663 5578 664 5582
rect 668 5578 669 5582
rect 673 5578 674 5582
rect 678 5578 679 5582
rect 683 5578 684 5582
rect 688 5578 689 5582
rect 931 5581 939 5585
rect 1129 5583 1359 5586
rect 1363 5582 1421 5586
rect 1604 5583 1713 5586
rect 1876 5581 1884 5585
rect 2074 5583 2304 5586
rect 2308 5582 2366 5586
rect 2549 5583 2658 5586
rect 659 5577 693 5578
rect 663 5573 664 5577
rect 668 5573 669 5577
rect 673 5573 674 5577
rect 678 5573 679 5577
rect 683 5573 684 5577
rect 688 5573 689 5577
rect 947 5575 955 5579
rect 959 5575 983 5579
rect 987 5575 995 5579
rect 999 5575 1000 5579
rect 1004 5575 1037 5579
rect 1041 5575 1056 5579
rect 1060 5575 1062 5579
rect 1066 5575 1073 5579
rect 1077 5575 1091 5579
rect 1095 5575 1107 5579
rect 1111 5575 1122 5579
rect 1126 5575 1133 5579
rect 1137 5575 1176 5579
rect 1180 5575 1216 5579
rect 1220 5575 1244 5579
rect 1248 5575 1256 5579
rect 1260 5575 1261 5579
rect 1265 5575 1298 5579
rect 1302 5575 1317 5579
rect 1321 5575 1323 5579
rect 1327 5575 1334 5579
rect 1338 5575 1352 5579
rect 1356 5575 1368 5579
rect 1372 5575 1457 5579
rect 1472 5576 1856 5579
rect 1892 5575 1900 5579
rect 1904 5575 1928 5579
rect 1932 5575 1940 5579
rect 1944 5575 1945 5579
rect 1949 5575 1982 5579
rect 1986 5575 2001 5579
rect 2005 5575 2007 5579
rect 2011 5575 2018 5579
rect 2022 5575 2036 5579
rect 2040 5575 2052 5579
rect 2056 5575 2067 5579
rect 2071 5575 2078 5579
rect 2082 5575 2121 5579
rect 2125 5575 2161 5579
rect 2165 5575 2189 5579
rect 2193 5575 2201 5579
rect 2205 5575 2206 5579
rect 2210 5575 2243 5579
rect 2247 5575 2262 5579
rect 2266 5575 2268 5579
rect 2272 5575 2279 5579
rect 2283 5575 2297 5579
rect 2301 5575 2313 5579
rect 2317 5575 2402 5579
rect 2417 5576 2801 5579
rect 659 5572 693 5573
rect 663 5568 664 5572
rect 668 5568 669 5572
rect 673 5568 674 5572
rect 678 5568 679 5572
rect 683 5568 684 5572
rect 688 5568 689 5572
rect 948 5568 962 5572
rect 966 5568 1027 5572
rect 1031 5568 1049 5572
rect 1053 5568 1080 5572
rect 1084 5568 1124 5572
rect 1128 5568 1133 5572
rect 659 5567 693 5568
rect 663 5563 664 5567
rect 668 5563 669 5567
rect 673 5563 674 5567
rect 678 5563 679 5567
rect 683 5563 684 5567
rect 688 5563 689 5567
rect 86 5307 89 5561
rect 343 5522 346 5561
rect 967 5561 969 5565
rect 1013 5561 1014 5565
rect 1038 5561 1041 5565
rect 1170 5563 1173 5575
rect 1209 5568 1223 5572
rect 1227 5568 1288 5572
rect 1292 5568 1310 5572
rect 1314 5568 1341 5572
rect 1345 5568 1359 5572
rect 1415 5569 1485 5572
rect 1489 5569 1535 5573
rect 1539 5569 1586 5573
rect 1590 5569 1617 5573
rect 1621 5569 1667 5573
rect 1671 5569 1718 5573
rect 1722 5569 1749 5573
rect 1753 5569 1799 5573
rect 1803 5569 1850 5573
rect 1854 5569 1863 5573
rect 1893 5568 1907 5572
rect 1911 5568 1972 5572
rect 1976 5568 1994 5572
rect 1998 5568 2025 5572
rect 2029 5568 2069 5572
rect 2073 5568 2078 5572
rect 948 5545 951 5550
rect 966 5546 969 5550
rect 966 5542 967 5546
rect 991 5545 994 5550
rect 1012 5546 1015 5550
rect 1022 5546 1025 5550
rect 948 5536 951 5541
rect 966 5536 969 5542
rect 986 5541 989 5544
rect 993 5541 994 5545
rect 1006 5542 1015 5546
rect 991 5536 994 5541
rect 1012 5536 1015 5542
rect 1022 5536 1025 5542
rect 1038 5547 1041 5550
rect 1038 5543 1040 5547
rect 1066 5545 1069 5550
rect 1082 5546 1085 5550
rect 1038 5536 1041 5543
rect 1058 5543 1069 5545
rect 1058 5541 1059 5543
rect 1063 5541 1069 5543
rect 1077 5542 1079 5546
rect 1083 5542 1085 5546
rect 1066 5536 1069 5541
rect 1082 5536 1085 5542
rect 1091 5544 1094 5550
rect 1098 5544 1101 5550
rect 1122 5544 1125 5558
rect 1228 5561 1230 5565
rect 1274 5561 1275 5565
rect 1299 5561 1302 5565
rect 1451 5562 1504 5566
rect 1508 5562 1534 5566
rect 1538 5562 1562 5566
rect 1566 5562 1636 5566
rect 1640 5562 1666 5566
rect 1670 5562 1694 5566
rect 1698 5562 1768 5566
rect 1772 5562 1798 5566
rect 1802 5562 1826 5566
rect 1830 5562 1863 5566
rect 1154 5552 1157 5555
rect 1149 5549 1157 5552
rect 1091 5541 1125 5544
rect 1154 5543 1157 5549
rect 1172 5548 1174 5551
rect 1178 5547 1183 5552
rect 1209 5545 1212 5550
rect 1227 5546 1230 5550
rect 1091 5536 1094 5541
rect 1098 5536 1101 5541
rect 1107 5536 1110 5541
rect 1227 5542 1228 5546
rect 1252 5545 1255 5550
rect 1273 5546 1276 5550
rect 1283 5546 1286 5550
rect 976 5523 977 5527
rect 1023 5524 1024 5528
rect 1048 5523 1049 5527
rect 343 5512 356 5522
rect 1134 5520 1137 5532
rect 948 5516 977 5520
rect 981 5516 1008 5520
rect 1012 5516 1033 5520
rect 1037 5516 1092 5520
rect 1096 5516 1114 5520
rect 1118 5516 1137 5520
rect 1170 5513 1173 5539
rect 1209 5536 1212 5541
rect 1227 5536 1230 5542
rect 1247 5541 1250 5544
rect 1254 5541 1255 5545
rect 1267 5542 1276 5546
rect 1252 5536 1255 5541
rect 1273 5536 1276 5542
rect 1283 5536 1286 5542
rect 1299 5547 1302 5550
rect 1299 5543 1301 5547
rect 1327 5545 1330 5550
rect 1343 5546 1346 5550
rect 1299 5536 1302 5543
rect 1319 5543 1330 5545
rect 1319 5541 1320 5543
rect 1324 5541 1330 5543
rect 1338 5542 1340 5546
rect 1344 5542 1346 5546
rect 1327 5536 1330 5541
rect 1343 5536 1346 5542
rect 1352 5544 1355 5550
rect 1477 5550 1480 5562
rect 1498 5550 1501 5562
rect 1514 5550 1517 5562
rect 1533 5556 1545 5559
rect 1556 5550 1559 5562
rect 1572 5550 1575 5562
rect 1593 5550 1596 5562
rect 1609 5550 1612 5562
rect 1630 5550 1633 5562
rect 1646 5550 1649 5562
rect 1665 5556 1677 5559
rect 1688 5550 1691 5562
rect 1704 5550 1707 5562
rect 1725 5550 1728 5562
rect 1741 5550 1744 5562
rect 1762 5550 1765 5562
rect 1778 5550 1781 5562
rect 1797 5556 1809 5559
rect 1820 5550 1823 5562
rect 1836 5550 1839 5562
rect 1857 5550 1860 5562
rect 1912 5561 1914 5565
rect 1958 5561 1959 5565
rect 1983 5561 1986 5565
rect 2115 5563 2118 5575
rect 4826 5573 5086 5576
rect 2154 5568 2168 5572
rect 2172 5568 2233 5572
rect 2237 5568 2255 5572
rect 2259 5568 2286 5572
rect 2290 5568 2304 5572
rect 2360 5569 2430 5572
rect 2434 5569 2480 5573
rect 2484 5569 2531 5573
rect 2535 5569 2562 5573
rect 2566 5569 2612 5573
rect 2616 5569 2663 5573
rect 2667 5569 2694 5573
rect 2698 5569 2744 5573
rect 2748 5569 2795 5573
rect 2799 5569 2808 5573
rect 1359 5544 1362 5550
rect 1352 5541 1362 5544
rect 1370 5541 1372 5544
rect 1352 5536 1355 5541
rect 1359 5536 1362 5541
rect 1477 5536 1494 5539
rect 1498 5540 1505 5543
rect 1530 5540 1533 5546
rect 1533 5536 1552 5539
rect 1556 5540 1563 5543
rect 1611 5536 1626 5539
rect 1630 5540 1637 5543
rect 1662 5540 1665 5546
rect 1665 5536 1684 5539
rect 1688 5540 1695 5543
rect 1743 5536 1758 5539
rect 1762 5540 1769 5543
rect 1794 5540 1797 5546
rect 1797 5536 1816 5539
rect 1820 5540 1827 5543
rect 1893 5545 1896 5550
rect 1911 5546 1914 5550
rect 1911 5542 1912 5546
rect 1936 5545 1939 5550
rect 1957 5546 1960 5550
rect 1967 5546 1970 5550
rect 1893 5536 1896 5541
rect 1911 5536 1914 5542
rect 1931 5541 1934 5544
rect 1938 5541 1939 5545
rect 1951 5542 1960 5546
rect 1936 5536 1939 5541
rect 1957 5536 1960 5542
rect 1967 5536 1970 5542
rect 1237 5523 1238 5527
rect 1284 5524 1285 5528
rect 1309 5523 1310 5527
rect 1488 5530 1510 5533
rect 1514 5530 1521 5533
rect 1209 5516 1238 5520
rect 1242 5516 1269 5520
rect 1273 5516 1294 5520
rect 1298 5516 1344 5520
rect 1348 5516 1353 5520
rect 1357 5516 1433 5520
rect 1546 5530 1570 5533
rect 1574 5530 1579 5533
rect 1593 5530 1600 5533
rect 1620 5530 1642 5533
rect 1646 5530 1653 5533
rect 1678 5530 1702 5533
rect 1706 5530 1711 5533
rect 1725 5530 1732 5533
rect 1752 5530 1774 5533
rect 1778 5530 1785 5533
rect 1810 5530 1834 5533
rect 1838 5530 1843 5533
rect 1983 5547 1986 5550
rect 1983 5543 1985 5547
rect 2011 5545 2014 5550
rect 2027 5546 2030 5550
rect 1983 5536 1986 5543
rect 2003 5543 2014 5545
rect 2003 5541 2004 5543
rect 2008 5541 2014 5543
rect 2022 5542 2024 5546
rect 2028 5542 2030 5546
rect 2011 5536 2014 5541
rect 2027 5536 2030 5542
rect 2036 5544 2039 5550
rect 2043 5544 2046 5550
rect 2067 5544 2070 5558
rect 2173 5561 2175 5565
rect 2219 5561 2220 5565
rect 2244 5561 2247 5565
rect 2396 5562 2449 5566
rect 2453 5562 2479 5566
rect 2483 5562 2507 5566
rect 2511 5562 2581 5566
rect 2585 5562 2611 5566
rect 2615 5562 2639 5566
rect 2643 5562 2713 5566
rect 2717 5562 2743 5566
rect 2747 5562 2771 5566
rect 2775 5562 2808 5566
rect 2099 5552 2102 5555
rect 2094 5549 2102 5552
rect 2036 5541 2070 5544
rect 2099 5543 2102 5549
rect 2117 5548 2119 5551
rect 2123 5547 2128 5552
rect 2154 5545 2157 5550
rect 2172 5546 2175 5550
rect 2036 5536 2039 5541
rect 2043 5536 2046 5541
rect 2052 5536 2055 5541
rect 2172 5542 2173 5546
rect 2197 5545 2200 5550
rect 2218 5546 2221 5550
rect 2228 5546 2231 5550
rect 1921 5523 1922 5527
rect 1968 5524 1969 5528
rect 1993 5523 1994 5527
rect 2079 5520 2082 5532
rect 343 5502 366 5512
rect 947 5509 956 5513
rect 960 5509 984 5513
rect 988 5509 999 5513
rect 1003 5509 1033 5513
rect 1037 5509 1056 5513
rect 1060 5509 1065 5513
rect 1069 5509 1074 5513
rect 1078 5509 1092 5513
rect 1096 5509 1176 5513
rect 1180 5509 1200 5513
rect 1204 5509 1217 5513
rect 1221 5509 1245 5513
rect 1249 5509 1260 5513
rect 1264 5509 1294 5513
rect 1298 5509 1317 5513
rect 1321 5509 1326 5513
rect 1330 5509 1335 5513
rect 1339 5509 1353 5513
rect 1357 5509 1361 5513
rect 1365 5509 1367 5513
rect 1371 5509 1445 5513
rect 1477 5509 1480 5519
rect 1498 5509 1501 5519
rect 1514 5509 1517 5519
rect 1529 5512 1536 5516
rect 1540 5512 1545 5516
rect 1556 5509 1559 5519
rect 1572 5509 1575 5519
rect 1593 5509 1596 5519
rect 1609 5509 1612 5519
rect 1630 5509 1633 5519
rect 1646 5509 1649 5519
rect 1661 5512 1668 5516
rect 1672 5512 1677 5516
rect 1688 5509 1691 5519
rect 1704 5509 1707 5519
rect 1725 5509 1728 5519
rect 1741 5509 1744 5519
rect 1762 5509 1765 5519
rect 1778 5509 1781 5519
rect 1793 5512 1800 5516
rect 1804 5512 1809 5516
rect 1820 5509 1823 5519
rect 1836 5509 1839 5519
rect 1857 5509 1860 5519
rect 1893 5516 1922 5520
rect 1926 5516 1953 5520
rect 1957 5516 1978 5520
rect 1982 5516 2037 5520
rect 2041 5516 2059 5520
rect 2063 5516 2082 5520
rect 2115 5513 2118 5539
rect 2154 5536 2157 5541
rect 2172 5536 2175 5542
rect 2192 5541 2195 5544
rect 2199 5541 2200 5545
rect 2212 5542 2221 5546
rect 2197 5536 2200 5541
rect 2218 5536 2221 5542
rect 2228 5536 2231 5542
rect 2244 5547 2247 5550
rect 2244 5543 2246 5547
rect 2272 5545 2275 5550
rect 2288 5546 2291 5550
rect 2244 5536 2247 5543
rect 2264 5543 2275 5545
rect 2264 5541 2265 5543
rect 2269 5541 2275 5543
rect 2283 5542 2285 5546
rect 2289 5542 2291 5546
rect 2272 5536 2275 5541
rect 2288 5536 2291 5542
rect 2297 5544 2300 5550
rect 2422 5550 2425 5562
rect 2443 5550 2446 5562
rect 2459 5550 2462 5562
rect 2478 5556 2490 5559
rect 2501 5550 2504 5562
rect 2517 5550 2520 5562
rect 2538 5550 2541 5562
rect 2554 5550 2557 5562
rect 2575 5550 2578 5562
rect 2591 5550 2594 5562
rect 2610 5556 2622 5559
rect 2633 5550 2636 5562
rect 2649 5550 2652 5562
rect 2670 5550 2673 5562
rect 2686 5550 2689 5562
rect 2707 5550 2710 5562
rect 2723 5550 2726 5562
rect 2742 5556 2754 5559
rect 2765 5550 2768 5562
rect 2781 5550 2784 5562
rect 2802 5550 2805 5562
rect 2304 5544 2307 5550
rect 2297 5541 2307 5544
rect 2315 5541 2317 5544
rect 2297 5536 2300 5541
rect 2304 5536 2307 5541
rect 2422 5536 2439 5539
rect 2443 5540 2450 5543
rect 2475 5540 2478 5546
rect 2478 5536 2497 5539
rect 2501 5540 2508 5543
rect 2556 5536 2571 5539
rect 2575 5540 2582 5543
rect 2607 5540 2610 5546
rect 2610 5536 2629 5539
rect 2633 5540 2640 5543
rect 2688 5536 2703 5539
rect 2707 5540 2714 5543
rect 2739 5540 2742 5546
rect 2742 5536 2761 5539
rect 2765 5540 2772 5543
rect 2182 5523 2183 5527
rect 2229 5524 2230 5528
rect 2254 5523 2255 5527
rect 2433 5530 2455 5533
rect 2459 5530 2466 5533
rect 2154 5516 2183 5520
rect 2187 5516 2214 5520
rect 2218 5516 2239 5520
rect 2243 5516 2289 5520
rect 2293 5516 2298 5520
rect 2302 5516 2378 5520
rect 2491 5530 2515 5533
rect 2519 5530 2524 5533
rect 2538 5530 2545 5533
rect 2565 5530 2587 5533
rect 2591 5530 2598 5533
rect 2623 5530 2647 5533
rect 2651 5530 2656 5533
rect 2670 5530 2677 5533
rect 2697 5530 2719 5533
rect 2723 5530 2730 5533
rect 2755 5530 2779 5533
rect 2783 5530 2788 5533
rect 2801 5532 4246 5536
rect 4251 5532 4255 5536
rect 4826 5534 4829 5573
rect 4816 5524 4829 5534
rect 1892 5509 1901 5513
rect 1905 5509 1929 5513
rect 1933 5509 1944 5513
rect 1948 5509 1978 5513
rect 1982 5509 2001 5513
rect 2005 5509 2010 5513
rect 2014 5509 2019 5513
rect 2023 5509 2037 5513
rect 2041 5509 2121 5513
rect 2125 5509 2145 5513
rect 2149 5509 2162 5513
rect 2166 5509 2190 5513
rect 2194 5509 2205 5513
rect 2209 5509 2239 5513
rect 2243 5509 2262 5513
rect 2266 5509 2271 5513
rect 2275 5509 2280 5513
rect 2284 5509 2298 5513
rect 2302 5509 2306 5513
rect 2310 5509 2312 5513
rect 2316 5509 2390 5513
rect 2422 5509 2425 5519
rect 2443 5509 2446 5519
rect 2459 5509 2462 5519
rect 2474 5512 2481 5516
rect 2485 5512 2490 5516
rect 2501 5509 2504 5519
rect 2517 5509 2520 5519
rect 2538 5509 2541 5519
rect 2554 5509 2557 5519
rect 2575 5509 2578 5519
rect 2591 5509 2594 5519
rect 2606 5512 2613 5516
rect 2617 5512 2622 5516
rect 2633 5509 2636 5519
rect 2649 5509 2652 5519
rect 2670 5509 2673 5519
rect 2686 5509 2689 5519
rect 2707 5509 2710 5519
rect 2723 5509 2726 5519
rect 2738 5512 2745 5516
rect 2749 5512 2754 5516
rect 2765 5509 2768 5519
rect 2781 5509 2784 5519
rect 2802 5509 2805 5519
rect 4806 5514 4829 5524
rect 343 5492 376 5502
rect 343 5482 386 5492
rect 1140 5485 1143 5509
rect 343 5386 769 5482
rect 1170 5481 1173 5509
rect 1209 5502 1238 5506
rect 1242 5502 1269 5506
rect 1273 5502 1294 5506
rect 1298 5502 1344 5506
rect 1348 5502 1353 5506
rect 1357 5502 1378 5506
rect 1463 5505 1467 5509
rect 1471 5505 1504 5509
rect 1508 5505 1534 5509
rect 1538 5505 1562 5509
rect 1566 5505 1599 5509
rect 1603 5505 1636 5509
rect 1640 5505 1666 5509
rect 1670 5505 1694 5509
rect 1698 5505 1731 5509
rect 1735 5505 1768 5509
rect 1772 5505 1798 5509
rect 1802 5505 1826 5509
rect 1830 5505 1863 5509
rect 1237 5495 1238 5499
rect 1284 5494 1285 5498
rect 1309 5495 1310 5499
rect 1403 5498 1483 5502
rect 1487 5498 1550 5502
rect 1554 5498 1586 5502
rect 1590 5498 1615 5502
rect 1619 5498 1682 5502
rect 1686 5498 1718 5502
rect 1722 5498 1747 5502
rect 1751 5498 1814 5502
rect 1818 5498 1850 5502
rect 1854 5498 1863 5502
rect 1177 5482 1182 5487
rect 1131 5476 1134 5481
rect 1209 5481 1212 5486
rect 1126 5473 1134 5476
rect 1121 5468 1126 5473
rect 1131 5459 1134 5473
rect 1142 5473 1145 5476
rect 1154 5471 1157 5477
rect 1177 5472 1180 5478
rect 1227 5480 1230 5486
rect 1252 5481 1255 5486
rect 1149 5468 1157 5471
rect 1169 5469 1180 5472
rect 1209 5472 1212 5477
rect 1227 5476 1228 5480
rect 1247 5478 1250 5481
rect 1254 5477 1255 5481
rect 1273 5480 1276 5486
rect 1283 5480 1286 5486
rect 1227 5472 1230 5476
rect 1252 5472 1255 5477
rect 1267 5476 1276 5480
rect 1273 5472 1276 5476
rect 1283 5472 1286 5476
rect 1154 5465 1157 5468
rect 1299 5479 1302 5486
rect 1299 5475 1301 5479
rect 1319 5479 1320 5481
rect 1327 5481 1330 5486
rect 1324 5479 1330 5481
rect 1343 5480 1346 5486
rect 1319 5477 1330 5479
rect 1299 5472 1302 5475
rect 1327 5472 1330 5477
rect 1338 5476 1340 5480
rect 1344 5476 1346 5480
rect 1343 5472 1346 5476
rect 1352 5481 1355 5486
rect 1359 5481 1362 5486
rect 2085 5485 2088 5509
rect 2115 5481 2118 5509
rect 2154 5502 2183 5506
rect 2187 5502 2214 5506
rect 2218 5502 2239 5506
rect 2243 5502 2289 5506
rect 2293 5502 2298 5506
rect 2302 5502 2323 5506
rect 2408 5505 2412 5509
rect 2416 5505 2449 5509
rect 2453 5505 2479 5509
rect 2483 5505 2507 5509
rect 2511 5505 2544 5509
rect 2548 5505 2581 5509
rect 2585 5505 2611 5509
rect 2615 5505 2639 5509
rect 2643 5505 2676 5509
rect 2680 5505 2713 5509
rect 2717 5505 2743 5509
rect 2747 5505 2771 5509
rect 2775 5505 2808 5509
rect 4796 5504 4829 5514
rect 2182 5495 2183 5499
rect 2229 5494 2230 5498
rect 2254 5495 2255 5499
rect 2348 5498 2428 5502
rect 2432 5498 2495 5502
rect 2499 5498 2531 5502
rect 2535 5498 2560 5502
rect 2564 5498 2627 5502
rect 2631 5498 2663 5502
rect 2667 5498 2692 5502
rect 2696 5498 2759 5502
rect 2763 5498 2795 5502
rect 2799 5498 2808 5502
rect 4786 5494 4829 5504
rect 2122 5482 2127 5487
rect 1352 5478 1362 5481
rect 1352 5472 1355 5478
rect 1359 5472 1362 5478
rect 1370 5478 1373 5481
rect 2076 5476 2079 5481
rect 2154 5481 2157 5486
rect 2071 5473 2079 5476
rect 1504 5468 1785 5472
rect 1789 5468 1813 5472
rect 2066 5468 2071 5473
rect 1228 5457 1230 5461
rect 1274 5457 1275 5461
rect 1299 5457 1302 5461
rect 1140 5447 1143 5451
rect 1170 5447 1173 5457
rect 1779 5456 1782 5468
rect 1209 5450 1223 5454
rect 1227 5450 1288 5454
rect 1292 5450 1310 5454
rect 1314 5450 1341 5454
rect 1345 5450 1421 5454
rect 2076 5459 2079 5473
rect 2087 5473 2090 5476
rect 2099 5471 2102 5477
rect 2122 5472 2125 5478
rect 2172 5480 2175 5486
rect 2197 5481 2200 5486
rect 2094 5468 2102 5471
rect 2114 5469 2125 5472
rect 2154 5472 2157 5477
rect 2172 5476 2173 5480
rect 2192 5478 2195 5481
rect 2199 5477 2200 5481
rect 2218 5480 2221 5486
rect 2228 5480 2231 5486
rect 2172 5472 2175 5476
rect 2197 5472 2200 5477
rect 2212 5476 2221 5480
rect 2218 5472 2221 5476
rect 2228 5472 2231 5476
rect 2099 5465 2102 5468
rect 2244 5479 2247 5486
rect 2244 5475 2246 5479
rect 2264 5479 2265 5481
rect 2272 5481 2275 5486
rect 2269 5479 2275 5481
rect 2288 5480 2291 5486
rect 2264 5477 2275 5479
rect 2244 5472 2247 5475
rect 2272 5472 2275 5477
rect 2283 5476 2285 5480
rect 2289 5476 2291 5480
rect 2288 5472 2291 5476
rect 2297 5481 2300 5486
rect 2304 5481 2307 5486
rect 2297 5478 2307 5481
rect 2297 5472 2300 5478
rect 2304 5472 2307 5478
rect 2315 5478 2318 5481
rect 2173 5457 2175 5461
rect 2219 5457 2220 5461
rect 2244 5457 2247 5461
rect 951 5443 1005 5447
rect 1009 5443 1095 5447
rect 1099 5443 1122 5447
rect 1126 5443 1176 5447
rect 1180 5443 1200 5447
rect 1204 5443 1216 5447
rect 1220 5443 1244 5447
rect 1248 5443 1256 5447
rect 1260 5443 1261 5447
rect 1265 5443 1298 5447
rect 1302 5443 1317 5447
rect 1321 5443 1323 5447
rect 1327 5443 1334 5447
rect 1338 5443 1352 5447
rect 1356 5443 1368 5447
rect 1372 5443 1457 5447
rect 1763 5445 1766 5448
rect 2085 5447 2088 5451
rect 2115 5447 2118 5457
rect 2154 5450 2168 5454
rect 2172 5450 2233 5454
rect 2237 5450 2255 5454
rect 2259 5450 2286 5454
rect 2290 5450 2366 5454
rect 999 5427 1002 5443
rect 1089 5427 1092 5443
rect 1170 5427 1173 5443
rect 1758 5442 1766 5445
rect 1209 5436 1223 5440
rect 1227 5436 1288 5440
rect 1292 5436 1310 5440
rect 1314 5436 1341 5440
rect 1345 5436 1421 5440
rect 1763 5436 1766 5442
rect 1781 5441 1840 5444
rect 1896 5443 1950 5447
rect 1954 5443 2040 5447
rect 2044 5443 2067 5447
rect 2071 5443 2121 5447
rect 2125 5443 2145 5447
rect 2149 5443 2161 5447
rect 2165 5443 2189 5447
rect 2193 5443 2201 5447
rect 2205 5443 2206 5447
rect 2210 5443 2243 5447
rect 2247 5443 2262 5447
rect 2266 5443 2268 5447
rect 2272 5443 2279 5447
rect 2283 5443 2297 5447
rect 2301 5443 2313 5447
rect 2317 5443 2402 5447
rect 1228 5429 1230 5433
rect 1274 5429 1275 5433
rect 1299 5429 1302 5433
rect 1415 5428 1680 5432
rect 983 5416 986 5419
rect 1073 5416 1076 5419
rect 1154 5416 1157 5419
rect 978 5413 986 5416
rect 983 5407 986 5413
rect 1001 5412 1009 5415
rect 1068 5413 1076 5416
rect 1073 5407 1076 5413
rect 1091 5412 1093 5415
rect 1097 5411 1102 5416
rect 1149 5413 1157 5416
rect 1154 5407 1157 5413
rect 1172 5412 1173 5415
rect 1177 5411 1182 5416
rect 1209 5413 1212 5418
rect 1227 5414 1230 5418
rect 1227 5410 1228 5414
rect 1252 5413 1255 5418
rect 1273 5414 1276 5418
rect 1283 5414 1286 5418
rect 343 5376 386 5386
rect 999 5381 1002 5403
rect 1089 5381 1092 5403
rect 1170 5381 1173 5403
rect 1209 5404 1212 5409
rect 1227 5404 1230 5410
rect 1247 5409 1250 5412
rect 1254 5409 1255 5413
rect 1267 5410 1276 5414
rect 1252 5404 1255 5409
rect 1273 5404 1276 5410
rect 1283 5404 1286 5410
rect 1299 5415 1302 5418
rect 1299 5411 1301 5415
rect 1327 5413 1330 5418
rect 1343 5414 1346 5418
rect 1299 5404 1302 5411
rect 1319 5411 1330 5413
rect 1319 5409 1320 5411
rect 1324 5409 1330 5411
rect 1338 5410 1340 5414
rect 1344 5410 1346 5414
rect 1327 5404 1330 5409
rect 1343 5404 1346 5410
rect 1352 5412 1355 5418
rect 1779 5422 1782 5432
rect 1944 5427 1947 5443
rect 2034 5427 2037 5443
rect 2115 5427 2118 5443
rect 2154 5436 2168 5440
rect 2172 5436 2233 5440
rect 2237 5436 2255 5440
rect 2259 5436 2286 5440
rect 2290 5436 2366 5440
rect 1512 5418 1682 5422
rect 1686 5418 1731 5422
rect 1735 5418 1785 5422
rect 1789 5418 1809 5422
rect 1813 5418 1831 5422
rect 2173 5429 2175 5433
rect 2219 5429 2220 5433
rect 2244 5429 2247 5433
rect 1359 5412 1362 5418
rect 1352 5409 1362 5412
rect 1370 5409 1372 5412
rect 1352 5404 1355 5409
rect 1359 5404 1362 5409
rect 1670 5411 1673 5418
rect 1723 5411 1726 5418
rect 1403 5399 1637 5402
rect 1403 5398 1636 5399
rect 1237 5391 1238 5395
rect 1284 5392 1285 5396
rect 1309 5391 1310 5395
rect 1209 5384 1238 5388
rect 1242 5384 1269 5388
rect 1273 5384 1294 5388
rect 1298 5384 1353 5388
rect 1357 5384 1433 5388
rect 955 5377 1005 5381
rect 1009 5377 1041 5381
rect 1045 5377 1095 5381
rect 1099 5377 1119 5381
rect 1126 5377 1176 5381
rect 1180 5377 1200 5381
rect 1204 5377 1217 5381
rect 1221 5377 1245 5381
rect 1249 5377 1260 5381
rect 1264 5377 1294 5381
rect 1298 5377 1317 5381
rect 1321 5377 1326 5381
rect 1330 5377 1335 5381
rect 1339 5377 1353 5381
rect 1357 5377 1361 5381
rect 1365 5377 1367 5381
rect 1371 5377 1445 5381
rect 1637 5379 1640 5395
rect 1690 5391 1693 5399
rect 1658 5387 1680 5391
rect 1684 5387 1693 5391
rect 1690 5379 1693 5387
rect 1711 5386 1734 5391
rect 343 5366 376 5376
rect 343 5356 366 5366
rect 343 5346 356 5356
rect 969 5353 972 5377
rect 999 5349 1002 5377
rect 343 5307 346 5346
rect 960 5344 963 5349
rect 1023 5345 1026 5377
rect 1059 5353 1062 5377
rect 943 5341 963 5344
rect 960 5327 963 5341
rect 971 5341 974 5344
rect 983 5339 986 5345
rect 978 5336 986 5339
rect 998 5338 1006 5340
rect 998 5337 1010 5338
rect 1089 5349 1092 5377
rect 1096 5350 1101 5355
rect 1050 5344 1053 5349
rect 1014 5336 1017 5341
rect 1044 5341 1053 5344
rect 983 5333 986 5336
rect 1025 5333 1028 5336
rect 969 5315 972 5319
rect 999 5315 1002 5325
rect 1014 5327 1017 5332
rect 1050 5327 1053 5341
rect 1061 5341 1064 5344
rect 1073 5339 1076 5345
rect 1096 5340 1099 5346
rect 1113 5345 1116 5377
rect 1140 5353 1143 5377
rect 1170 5349 1173 5377
rect 1209 5370 1238 5374
rect 1242 5370 1269 5374
rect 1273 5370 1294 5374
rect 1298 5370 1353 5374
rect 1357 5370 1433 5374
rect 1237 5363 1238 5367
rect 1284 5362 1285 5366
rect 1309 5363 1310 5367
rect 1177 5350 1182 5355
rect 1068 5336 1076 5339
rect 1088 5337 1099 5340
rect 1122 5344 1126 5348
rect 1131 5344 1134 5349
rect 1209 5349 1212 5354
rect 1104 5336 1107 5341
rect 1126 5341 1134 5344
rect 1073 5333 1076 5336
rect 1115 5333 1118 5336
rect 1122 5333 1123 5336
rect 1023 5315 1026 5319
rect 1059 5315 1062 5319
rect 1089 5315 1092 5325
rect 1104 5327 1107 5332
rect 1131 5327 1134 5341
rect 1142 5341 1145 5344
rect 1154 5339 1157 5345
rect 1177 5340 1180 5346
rect 1227 5348 1230 5354
rect 1252 5349 1255 5354
rect 1149 5336 1157 5339
rect 1169 5337 1180 5340
rect 1209 5340 1212 5345
rect 1227 5344 1228 5348
rect 1247 5346 1250 5349
rect 1254 5345 1255 5349
rect 1273 5348 1276 5354
rect 1283 5348 1286 5354
rect 1227 5340 1230 5344
rect 1252 5340 1255 5345
rect 1267 5344 1276 5348
rect 1273 5340 1276 5344
rect 1283 5340 1286 5344
rect 1154 5333 1157 5336
rect 1299 5347 1302 5354
rect 1299 5343 1301 5347
rect 1319 5347 1320 5349
rect 1327 5349 1330 5354
rect 1324 5347 1330 5349
rect 1343 5348 1346 5354
rect 1319 5345 1330 5347
rect 1299 5340 1302 5343
rect 1327 5340 1330 5345
rect 1338 5344 1340 5348
rect 1344 5344 1346 5348
rect 1343 5340 1346 5344
rect 1352 5349 1355 5354
rect 1359 5349 1362 5354
rect 1731 5371 1734 5386
rect 1749 5380 1752 5418
rect 1779 5376 1782 5418
rect 1740 5371 1743 5376
rect 1803 5372 1806 5418
rect 1825 5372 1828 5418
rect 1928 5416 1931 5419
rect 2018 5416 2021 5419
rect 2099 5416 2102 5419
rect 1923 5413 1931 5416
rect 1928 5407 1931 5413
rect 1946 5412 1954 5415
rect 2013 5413 2021 5416
rect 2018 5407 2021 5413
rect 2036 5412 2038 5415
rect 2042 5411 2047 5416
rect 2094 5413 2102 5416
rect 2099 5407 2102 5413
rect 2117 5412 2118 5415
rect 2122 5411 2127 5416
rect 2154 5413 2157 5418
rect 2172 5414 2175 5418
rect 2172 5410 2173 5414
rect 2197 5413 2200 5418
rect 2218 5414 2221 5418
rect 2228 5414 2231 5418
rect 1944 5381 1947 5403
rect 2034 5381 2037 5403
rect 2115 5381 2118 5403
rect 2154 5404 2157 5409
rect 2172 5404 2175 5410
rect 2192 5409 2195 5412
rect 2199 5409 2200 5413
rect 2212 5410 2221 5414
rect 2197 5404 2200 5409
rect 2218 5404 2221 5410
rect 2228 5404 2231 5410
rect 2244 5415 2247 5418
rect 2244 5411 2246 5415
rect 2272 5413 2275 5418
rect 2288 5414 2291 5418
rect 2244 5404 2247 5411
rect 2264 5411 2275 5413
rect 2264 5409 2265 5411
rect 2269 5409 2275 5411
rect 2283 5410 2285 5414
rect 2289 5410 2291 5414
rect 2272 5404 2275 5409
rect 2288 5404 2291 5410
rect 2297 5412 2300 5418
rect 2304 5412 2307 5418
rect 2297 5409 2307 5412
rect 2315 5409 2317 5412
rect 2297 5404 2300 5409
rect 2304 5404 2307 5409
rect 4403 5398 4829 5494
rect 2182 5391 2183 5395
rect 2229 5392 2230 5396
rect 2254 5391 2255 5395
rect 4786 5388 4829 5398
rect 2154 5384 2183 5388
rect 2187 5384 2214 5388
rect 2218 5384 2239 5388
rect 2243 5384 2298 5388
rect 2302 5384 2378 5388
rect 1900 5377 1950 5381
rect 1954 5377 1986 5381
rect 1990 5377 2040 5381
rect 2044 5377 2064 5381
rect 2071 5377 2121 5381
rect 2125 5377 2145 5381
rect 2149 5377 2162 5381
rect 2166 5377 2190 5381
rect 2194 5377 2205 5381
rect 2209 5377 2239 5381
rect 2243 5377 2262 5381
rect 2266 5377 2271 5381
rect 2275 5377 2280 5381
rect 2284 5377 2298 5381
rect 2302 5377 2306 5381
rect 2310 5377 2312 5381
rect 2316 5377 2390 5381
rect 4796 5378 4829 5388
rect 1731 5368 1743 5371
rect 1352 5346 1362 5349
rect 1352 5340 1355 5346
rect 1359 5340 1362 5346
rect 1370 5346 1373 5349
rect 1670 5342 1673 5349
rect 1723 5342 1726 5349
rect 1740 5354 1743 5368
rect 1751 5368 1754 5371
rect 1763 5366 1766 5372
rect 1758 5363 1766 5366
rect 1778 5364 1789 5367
rect 1794 5363 1797 5368
rect 1816 5363 1819 5368
rect 1763 5360 1766 5363
rect 1805 5360 1808 5363
rect 1812 5359 1815 5363
rect 1827 5360 1830 5363
rect 1834 5360 1835 5363
rect 1749 5342 1752 5346
rect 1779 5342 1782 5352
rect 1794 5354 1797 5359
rect 1816 5354 1819 5359
rect 1914 5353 1917 5377
rect 1803 5342 1806 5346
rect 1825 5342 1828 5346
rect 1944 5349 1947 5377
rect 1504 5338 1682 5342
rect 1686 5338 1731 5342
rect 1735 5338 1785 5342
rect 1789 5338 1809 5342
rect 1813 5338 1831 5342
rect 1905 5344 1908 5349
rect 1968 5345 1971 5377
rect 2004 5353 2007 5377
rect 1888 5341 1908 5344
rect 1228 5325 1230 5329
rect 1274 5325 1275 5329
rect 1299 5325 1302 5329
rect 1779 5326 1782 5338
rect 1113 5315 1116 5319
rect 1140 5315 1143 5319
rect 1170 5315 1173 5325
rect 1209 5318 1223 5322
rect 1227 5318 1288 5322
rect 1292 5318 1310 5322
rect 1314 5318 1341 5322
rect 1345 5318 1421 5322
rect 1905 5327 1908 5341
rect 1916 5341 1919 5344
rect 1928 5339 1931 5345
rect 1923 5336 1931 5339
rect 1943 5338 1951 5340
rect 1943 5337 1955 5338
rect 2034 5349 2037 5377
rect 2041 5350 2046 5355
rect 1995 5344 1998 5349
rect 1959 5336 1962 5341
rect 1989 5341 1998 5344
rect 1928 5333 1931 5336
rect 1970 5333 1973 5336
rect 1763 5315 1766 5318
rect 1914 5315 1917 5319
rect 1944 5315 1947 5325
rect 1959 5327 1962 5332
rect 1995 5327 1998 5341
rect 2006 5341 2009 5344
rect 2018 5339 2021 5345
rect 2041 5340 2044 5346
rect 2058 5345 2061 5377
rect 2085 5353 2088 5377
rect 2115 5349 2118 5377
rect 2154 5370 2183 5374
rect 2187 5370 2214 5374
rect 2218 5370 2239 5374
rect 2243 5370 2298 5374
rect 2302 5370 2378 5374
rect 4806 5368 4829 5378
rect 2182 5363 2183 5367
rect 2229 5362 2230 5366
rect 2254 5363 2255 5367
rect 4816 5358 4829 5368
rect 2122 5350 2127 5355
rect 2013 5336 2021 5339
rect 2033 5337 2044 5340
rect 2067 5344 2071 5348
rect 2076 5344 2079 5349
rect 2154 5349 2157 5354
rect 2049 5336 2052 5341
rect 2071 5341 2079 5344
rect 2018 5333 2021 5336
rect 2060 5333 2063 5336
rect 2067 5333 2068 5336
rect 1968 5315 1971 5319
rect 2004 5315 2007 5319
rect 2034 5315 2037 5325
rect 2049 5327 2052 5332
rect 2076 5327 2079 5341
rect 2087 5341 2090 5344
rect 2099 5339 2102 5345
rect 2122 5340 2125 5346
rect 2172 5348 2175 5354
rect 2197 5349 2200 5354
rect 2094 5336 2102 5339
rect 2114 5337 2125 5340
rect 2154 5340 2157 5345
rect 2172 5344 2173 5348
rect 2192 5346 2195 5349
rect 2199 5345 2200 5349
rect 2218 5348 2221 5354
rect 2228 5348 2231 5354
rect 2172 5340 2175 5344
rect 2197 5340 2200 5345
rect 2212 5344 2221 5348
rect 2218 5340 2221 5344
rect 2228 5340 2231 5344
rect 2099 5333 2102 5336
rect 2244 5347 2247 5354
rect 2244 5343 2246 5347
rect 2264 5347 2265 5349
rect 2272 5349 2275 5354
rect 2269 5347 2275 5349
rect 2288 5348 2291 5354
rect 2264 5345 2275 5347
rect 2244 5340 2247 5343
rect 2272 5340 2275 5345
rect 2283 5344 2285 5348
rect 2289 5344 2291 5348
rect 2288 5340 2291 5344
rect 2297 5349 2300 5354
rect 2304 5349 2307 5354
rect 2297 5346 2307 5349
rect 2297 5340 2300 5346
rect 2304 5340 2307 5346
rect 2315 5346 2318 5349
rect 2173 5325 2175 5329
rect 2219 5325 2220 5329
rect 2244 5325 2247 5329
rect 2058 5315 2061 5319
rect 2085 5315 2088 5319
rect 2115 5315 2118 5325
rect 2154 5318 2168 5322
rect 2172 5318 2233 5322
rect 2237 5318 2255 5322
rect 2259 5318 2286 5322
rect 2290 5318 2366 5322
rect 4826 5319 4829 5358
rect 5083 5319 5086 5573
rect 955 5311 1005 5315
rect 1009 5311 1033 5315
rect 1037 5311 1041 5315
rect 1045 5311 1095 5315
rect 1099 5311 1122 5315
rect 1126 5311 1176 5315
rect 1180 5311 1200 5315
rect 1204 5311 1216 5315
rect 1220 5311 1244 5315
rect 1248 5311 1256 5315
rect 1260 5311 1261 5315
rect 1265 5311 1298 5315
rect 1302 5311 1317 5315
rect 1321 5311 1323 5315
rect 1327 5311 1334 5315
rect 1338 5311 1352 5315
rect 1356 5311 1368 5315
rect 1372 5311 1457 5315
rect 1758 5312 1766 5315
rect 86 5304 346 5307
rect 1065 5292 1068 5311
rect 1170 5292 1173 5311
rect 1209 5304 1223 5308
rect 1227 5304 1288 5308
rect 1292 5304 1310 5308
rect 1314 5304 1341 5308
rect 1345 5304 1421 5308
rect 1763 5306 1766 5312
rect 1781 5311 1842 5314
rect 1900 5311 1950 5315
rect 1954 5311 1978 5315
rect 1982 5311 1986 5315
rect 1990 5311 2040 5315
rect 2044 5311 2067 5315
rect 2071 5311 2121 5315
rect 2125 5311 2145 5315
rect 2149 5311 2161 5315
rect 2165 5311 2189 5315
rect 2193 5311 2201 5315
rect 2205 5311 2206 5315
rect 2210 5311 2243 5315
rect 2247 5311 2262 5315
rect 2266 5311 2268 5315
rect 2272 5311 2279 5315
rect 2283 5311 2297 5315
rect 2301 5311 2313 5315
rect 2317 5311 2402 5315
rect 4483 5313 4484 5317
rect 4488 5313 4489 5317
rect 4493 5313 4494 5317
rect 4498 5313 4499 5317
rect 4503 5313 4504 5317
rect 4508 5313 4509 5317
rect 4479 5312 4513 5313
rect 1439 5302 1574 5306
rect 1228 5297 1230 5301
rect 1274 5297 1275 5301
rect 1299 5297 1302 5301
rect 1049 5281 1052 5284
rect 1154 5281 1157 5284
rect 1209 5281 1212 5286
rect 1227 5282 1230 5286
rect 1044 5278 1052 5281
rect 617 5269 618 5273
rect 622 5269 623 5273
rect 627 5269 628 5273
rect 632 5269 633 5273
rect 637 5269 638 5273
rect 642 5269 643 5273
rect 613 5268 647 5269
rect 617 5264 618 5268
rect 622 5264 623 5268
rect 627 5264 628 5268
rect 632 5264 633 5268
rect 637 5264 638 5268
rect 642 5264 643 5268
rect 613 5263 647 5264
rect 617 5259 618 5263
rect 622 5259 623 5263
rect 627 5259 628 5263
rect 632 5259 633 5263
rect 637 5259 638 5263
rect 642 5259 643 5263
rect 613 5258 647 5259
rect 86 5252 346 5255
rect 617 5254 618 5258
rect 622 5254 623 5258
rect 627 5254 628 5258
rect 632 5254 633 5258
rect 637 5254 638 5258
rect 642 5254 643 5258
rect 663 5269 664 5273
rect 668 5269 669 5273
rect 673 5269 674 5273
rect 678 5269 679 5273
rect 683 5269 684 5273
rect 688 5269 689 5273
rect 659 5268 693 5269
rect 1049 5272 1052 5278
rect 1067 5277 1068 5280
rect 1072 5276 1077 5281
rect 1149 5278 1157 5281
rect 1154 5272 1157 5278
rect 1172 5277 1174 5280
rect 1178 5276 1183 5281
rect 1227 5278 1228 5282
rect 1252 5281 1255 5286
rect 1273 5282 1276 5286
rect 1283 5282 1286 5286
rect 1209 5272 1212 5277
rect 1227 5272 1230 5278
rect 1247 5277 1250 5280
rect 1254 5277 1255 5281
rect 1267 5278 1276 5282
rect 1252 5272 1255 5277
rect 1273 5272 1276 5278
rect 1283 5272 1286 5278
rect 1299 5283 1302 5286
rect 1299 5279 1301 5283
rect 1327 5281 1330 5286
rect 1343 5282 1346 5286
rect 1299 5272 1302 5279
rect 1319 5279 1330 5281
rect 1319 5277 1320 5279
rect 1324 5277 1330 5279
rect 1338 5278 1340 5282
rect 1344 5278 1346 5282
rect 1327 5272 1330 5277
rect 1343 5272 1346 5278
rect 1352 5280 1355 5286
rect 1391 5293 1492 5297
rect 1779 5292 1782 5302
rect 2010 5292 2013 5311
rect 2115 5292 2118 5311
rect 4483 5308 4484 5312
rect 4488 5308 4489 5312
rect 4493 5308 4494 5312
rect 4498 5308 4499 5312
rect 4503 5308 4504 5312
rect 4508 5308 4509 5312
rect 2154 5304 2168 5308
rect 2172 5304 2233 5308
rect 2237 5304 2255 5308
rect 2259 5304 2286 5308
rect 2290 5304 2366 5308
rect 4479 5307 4513 5308
rect 4483 5303 4484 5307
rect 4488 5303 4489 5307
rect 4493 5303 4494 5307
rect 4498 5303 4499 5307
rect 4503 5303 4504 5307
rect 4508 5303 4509 5307
rect 4479 5302 4513 5303
rect 2173 5297 2175 5301
rect 2219 5297 2220 5301
rect 2244 5297 2247 5301
rect 4483 5298 4484 5302
rect 4488 5298 4489 5302
rect 4493 5298 4494 5302
rect 4498 5298 4499 5302
rect 4503 5298 4504 5302
rect 4508 5298 4509 5302
rect 4529 5313 4530 5317
rect 4534 5313 4535 5317
rect 4539 5313 4540 5317
rect 4544 5313 4545 5317
rect 4549 5313 4550 5317
rect 4554 5313 4555 5317
rect 4826 5316 5086 5319
rect 4525 5312 4559 5313
rect 4529 5308 4530 5312
rect 4534 5308 4535 5312
rect 4539 5308 4540 5312
rect 4544 5308 4545 5312
rect 4549 5308 4550 5312
rect 4554 5308 4555 5312
rect 4525 5307 4559 5308
rect 4529 5303 4530 5307
rect 4534 5303 4535 5307
rect 4539 5303 4540 5307
rect 4544 5303 4545 5307
rect 4549 5303 4550 5307
rect 4554 5303 4555 5307
rect 4525 5302 4559 5303
rect 4529 5298 4530 5302
rect 4534 5298 4535 5302
rect 4539 5298 4540 5302
rect 4544 5298 4545 5302
rect 4549 5298 4550 5302
rect 4554 5298 4555 5302
rect 1512 5288 1588 5292
rect 1592 5288 1731 5292
rect 1735 5288 1785 5292
rect 1789 5288 1809 5292
rect 1359 5280 1362 5286
rect 1451 5284 1512 5288
rect 1576 5281 1579 5288
rect 1629 5281 1632 5288
rect 1352 5277 1362 5280
rect 1370 5277 1372 5280
rect 1352 5272 1355 5277
rect 1359 5272 1362 5277
rect 1463 5277 1500 5281
rect 663 5264 664 5268
rect 668 5264 669 5268
rect 673 5264 674 5268
rect 678 5264 679 5268
rect 683 5264 684 5268
rect 688 5264 689 5268
rect 659 5263 693 5264
rect 663 5259 664 5263
rect 668 5259 669 5263
rect 673 5259 674 5263
rect 678 5259 679 5263
rect 683 5259 684 5263
rect 688 5259 689 5263
rect 659 5258 693 5259
rect 663 5254 664 5258
rect 668 5254 669 5258
rect 673 5254 674 5258
rect 678 5254 679 5258
rect 683 5254 684 5258
rect 688 5254 689 5258
rect 86 4998 89 5252
rect 343 5213 346 5252
rect 1065 5249 1068 5268
rect 1170 5249 1173 5268
rect 1427 5265 1542 5269
rect 1237 5259 1238 5263
rect 1284 5260 1285 5264
rect 1309 5259 1310 5263
rect 1209 5252 1238 5256
rect 1242 5252 1269 5256
rect 1273 5252 1294 5256
rect 1298 5252 1353 5256
rect 1357 5252 1433 5256
rect 1543 5249 1546 5265
rect 1596 5261 1599 5269
rect 1564 5257 1575 5261
rect 1579 5257 1599 5261
rect 1596 5249 1599 5257
rect 1617 5256 1734 5261
rect 1023 5245 1071 5249
rect 1075 5245 1095 5249
rect 1099 5245 1122 5249
rect 1126 5245 1176 5249
rect 1180 5245 1200 5249
rect 1204 5245 1217 5249
rect 1221 5245 1245 5249
rect 1249 5245 1260 5249
rect 1264 5245 1294 5249
rect 1298 5245 1317 5249
rect 1321 5245 1326 5249
rect 1330 5245 1335 5249
rect 1339 5245 1353 5249
rect 1357 5245 1361 5249
rect 1365 5245 1367 5249
rect 1371 5245 1445 5249
rect 1035 5221 1038 5245
rect 1065 5217 1068 5245
rect 1072 5218 1077 5223
rect 343 5203 356 5213
rect 1026 5212 1029 5217
rect 1023 5209 1029 5212
rect 343 5193 366 5203
rect 1026 5195 1029 5209
rect 1037 5209 1040 5212
rect 1049 5207 1052 5213
rect 1072 5208 1075 5214
rect 1089 5213 1092 5245
rect 1140 5221 1143 5245
rect 1170 5217 1173 5245
rect 1209 5238 1238 5242
rect 1242 5238 1269 5242
rect 1273 5238 1294 5242
rect 1298 5238 1353 5242
rect 1357 5238 1433 5242
rect 1237 5231 1238 5235
rect 1284 5230 1285 5234
rect 1309 5231 1310 5235
rect 1177 5218 1182 5223
rect 1044 5204 1052 5207
rect 1064 5205 1075 5208
rect 1131 5212 1134 5217
rect 1209 5217 1212 5222
rect 1126 5209 1134 5212
rect 1080 5204 1083 5209
rect 1121 5204 1126 5209
rect 1049 5201 1052 5204
rect 343 5183 376 5193
rect 1091 5201 1094 5204
rect 1098 5201 1099 5204
rect 1035 5183 1038 5187
rect 1065 5183 1068 5193
rect 1080 5195 1083 5200
rect 1131 5195 1134 5209
rect 1142 5209 1145 5212
rect 1154 5207 1157 5213
rect 1177 5208 1180 5214
rect 1227 5216 1230 5222
rect 1252 5217 1255 5222
rect 1149 5204 1157 5207
rect 1169 5205 1180 5208
rect 1209 5208 1212 5213
rect 1227 5212 1228 5216
rect 1247 5214 1250 5217
rect 1254 5213 1255 5217
rect 1273 5216 1276 5222
rect 1283 5216 1286 5222
rect 1227 5208 1230 5212
rect 1252 5208 1255 5213
rect 1267 5212 1276 5216
rect 1273 5208 1276 5212
rect 1283 5208 1286 5212
rect 1154 5201 1157 5204
rect 1299 5215 1302 5222
rect 1299 5211 1301 5215
rect 1319 5215 1320 5217
rect 1327 5217 1330 5222
rect 1324 5215 1330 5217
rect 1343 5216 1346 5222
rect 1319 5213 1330 5215
rect 1299 5208 1302 5211
rect 1327 5208 1330 5213
rect 1338 5212 1340 5216
rect 1344 5212 1346 5216
rect 1343 5208 1346 5212
rect 1352 5217 1355 5222
rect 1359 5217 1362 5222
rect 1731 5241 1734 5256
rect 1749 5250 1752 5288
rect 1779 5246 1782 5288
rect 1740 5241 1743 5246
rect 1803 5242 1806 5288
rect 1994 5281 1997 5284
rect 2099 5281 2102 5284
rect 2154 5281 2157 5286
rect 2172 5282 2175 5286
rect 1989 5278 1997 5281
rect 1994 5272 1997 5278
rect 2012 5277 2013 5280
rect 2017 5276 2022 5281
rect 2094 5278 2102 5281
rect 2099 5272 2102 5278
rect 2117 5277 2119 5280
rect 2123 5276 2128 5281
rect 2172 5278 2173 5282
rect 2197 5281 2200 5286
rect 2218 5282 2221 5286
rect 2228 5282 2231 5286
rect 2154 5272 2157 5277
rect 2172 5272 2175 5278
rect 2192 5277 2195 5280
rect 2199 5277 2200 5281
rect 2212 5278 2221 5282
rect 2197 5272 2200 5277
rect 2218 5272 2221 5278
rect 2228 5272 2231 5278
rect 2244 5283 2247 5286
rect 2244 5279 2246 5283
rect 2272 5281 2275 5286
rect 2288 5282 2291 5286
rect 2244 5272 2247 5279
rect 2264 5279 2275 5281
rect 2264 5277 2265 5279
rect 2269 5277 2275 5279
rect 2283 5278 2285 5282
rect 2289 5278 2291 5282
rect 2272 5272 2275 5277
rect 2288 5272 2291 5278
rect 2297 5280 2300 5286
rect 2304 5280 2307 5286
rect 2297 5277 2307 5280
rect 2315 5277 2317 5280
rect 2297 5272 2300 5277
rect 2304 5272 2307 5277
rect 2010 5249 2013 5268
rect 2115 5249 2118 5268
rect 4826 5264 5086 5267
rect 2182 5259 2183 5263
rect 2229 5260 2230 5264
rect 2254 5259 2255 5263
rect 2154 5252 2183 5256
rect 2187 5252 2214 5256
rect 2218 5252 2239 5256
rect 2243 5252 2298 5256
rect 2302 5252 2378 5256
rect 1968 5245 2016 5249
rect 2020 5245 2040 5249
rect 2044 5245 2067 5249
rect 2071 5245 2121 5249
rect 2125 5245 2145 5249
rect 2149 5245 2162 5249
rect 2166 5245 2190 5249
rect 2194 5245 2205 5249
rect 2209 5245 2239 5249
rect 2243 5245 2262 5249
rect 2266 5245 2271 5249
rect 2275 5245 2280 5249
rect 2284 5245 2298 5249
rect 2302 5245 2306 5249
rect 2310 5245 2312 5249
rect 2316 5245 2390 5249
rect 1731 5238 1743 5241
rect 1352 5214 1362 5217
rect 1352 5208 1355 5214
rect 1359 5208 1362 5214
rect 1370 5214 1373 5217
rect 1576 5212 1579 5219
rect 1629 5212 1632 5219
rect 1740 5224 1743 5238
rect 1751 5238 1754 5241
rect 1763 5236 1766 5242
rect 1758 5233 1766 5236
rect 1778 5234 1789 5237
rect 1794 5233 1797 5238
rect 1763 5230 1766 5233
rect 1805 5230 1808 5233
rect 1812 5230 1813 5233
rect 1749 5212 1752 5216
rect 1779 5212 1782 5222
rect 1794 5224 1797 5229
rect 1980 5221 1983 5245
rect 1803 5212 1806 5216
rect 2010 5217 2013 5245
rect 2017 5218 2022 5223
rect 1971 5212 1974 5217
rect 1504 5208 1588 5212
rect 1592 5208 1731 5212
rect 1735 5208 1785 5212
rect 1789 5208 1809 5212
rect 1968 5209 1974 5212
rect 1228 5193 1230 5197
rect 1274 5193 1275 5197
rect 1299 5193 1302 5197
rect 1971 5195 1974 5209
rect 1982 5209 1985 5212
rect 1994 5207 1997 5213
rect 2017 5208 2020 5214
rect 2034 5213 2037 5245
rect 2085 5221 2088 5245
rect 2115 5217 2118 5245
rect 2154 5238 2183 5242
rect 2187 5238 2214 5242
rect 2218 5238 2239 5242
rect 2243 5238 2298 5242
rect 2302 5238 2378 5242
rect 2182 5231 2183 5235
rect 2229 5230 2230 5234
rect 2254 5231 2255 5235
rect 2122 5218 2127 5223
rect 1989 5204 1997 5207
rect 2009 5205 2020 5208
rect 2076 5212 2079 5217
rect 2154 5217 2157 5222
rect 2071 5209 2079 5212
rect 2025 5204 2028 5209
rect 2066 5204 2071 5209
rect 1994 5201 1997 5204
rect 1089 5183 1092 5187
rect 1140 5183 1143 5187
rect 1170 5183 1173 5193
rect 1209 5186 1223 5190
rect 1227 5186 1288 5190
rect 1292 5186 1310 5190
rect 1314 5186 1341 5190
rect 1345 5186 1357 5190
rect 1361 5186 1421 5190
rect 1551 5189 1807 5194
rect 2036 5201 2039 5204
rect 2043 5201 2044 5204
rect 1980 5183 1983 5187
rect 2010 5183 2013 5193
rect 2025 5195 2028 5200
rect 2076 5195 2079 5209
rect 2087 5209 2090 5212
rect 2099 5207 2102 5213
rect 2122 5208 2125 5214
rect 2172 5216 2175 5222
rect 2197 5217 2200 5222
rect 2094 5204 2102 5207
rect 2114 5205 2125 5208
rect 2154 5208 2157 5213
rect 2172 5212 2173 5216
rect 2192 5214 2195 5217
rect 2199 5213 2200 5217
rect 2218 5216 2221 5222
rect 2228 5216 2231 5222
rect 2172 5208 2175 5212
rect 2197 5208 2200 5213
rect 2212 5212 2221 5216
rect 2218 5208 2221 5212
rect 2228 5208 2231 5212
rect 2099 5201 2102 5204
rect 2244 5215 2247 5222
rect 2244 5211 2246 5215
rect 2264 5215 2265 5217
rect 2272 5217 2275 5222
rect 2269 5215 2275 5217
rect 2288 5216 2291 5222
rect 2264 5213 2275 5215
rect 2244 5208 2247 5211
rect 2272 5208 2275 5213
rect 2283 5212 2285 5216
rect 2289 5212 2291 5216
rect 2288 5208 2291 5212
rect 2297 5217 2300 5222
rect 4826 5225 4829 5264
rect 2304 5217 2307 5222
rect 2297 5214 2307 5217
rect 2297 5208 2300 5214
rect 2304 5208 2307 5214
rect 2315 5214 2318 5217
rect 4816 5215 4829 5225
rect 4806 5205 4829 5215
rect 2173 5193 2175 5197
rect 2219 5193 2220 5197
rect 2244 5193 2247 5197
rect 4796 5195 4829 5205
rect 2034 5183 2037 5187
rect 2085 5183 2088 5187
rect 2115 5183 2118 5193
rect 2154 5186 2168 5190
rect 2172 5186 2233 5190
rect 2237 5186 2255 5190
rect 2259 5186 2286 5190
rect 2290 5186 2302 5190
rect 2306 5186 2366 5190
rect 4786 5185 4829 5195
rect 343 5173 386 5183
rect 1022 5179 1033 5183
rect 1037 5179 1095 5183
rect 1099 5179 1122 5183
rect 1126 5179 1176 5183
rect 1180 5179 1200 5183
rect 1204 5179 1216 5183
rect 1220 5179 1244 5183
rect 1248 5179 1256 5183
rect 1260 5179 1261 5183
rect 1265 5179 1298 5183
rect 1302 5179 1317 5183
rect 1321 5179 1323 5183
rect 1327 5179 1334 5183
rect 1338 5179 1352 5183
rect 1356 5179 1368 5183
rect 1372 5179 1457 5183
rect 1967 5179 1978 5183
rect 1982 5179 2040 5183
rect 2044 5179 2067 5183
rect 2071 5179 2121 5183
rect 2125 5179 2145 5183
rect 2149 5179 2161 5183
rect 2165 5179 2189 5183
rect 2193 5179 2201 5183
rect 2205 5179 2206 5183
rect 2210 5179 2243 5183
rect 2247 5179 2262 5183
rect 2266 5179 2268 5183
rect 2272 5179 2279 5183
rect 2283 5179 2297 5183
rect 2301 5179 2313 5183
rect 2317 5179 2402 5183
rect 343 5077 769 5173
rect 1089 5161 1092 5179
rect 1170 5161 1173 5179
rect 1209 5172 1223 5176
rect 1227 5172 1288 5176
rect 1292 5172 1310 5176
rect 1314 5172 1341 5176
rect 1345 5172 1357 5176
rect 1415 5169 1615 5173
rect 1619 5169 1666 5173
rect 1670 5169 1716 5173
rect 1720 5169 1738 5173
rect 1228 5165 1230 5169
rect 1274 5165 1275 5169
rect 1299 5165 1302 5169
rect 1451 5162 1639 5166
rect 1643 5162 1667 5166
rect 1671 5162 1697 5166
rect 1701 5162 1738 5166
rect 1073 5150 1076 5153
rect 1154 5150 1157 5153
rect 1068 5147 1076 5150
rect 1073 5141 1076 5147
rect 1091 5146 1093 5149
rect 1097 5145 1102 5150
rect 1149 5147 1157 5150
rect 1154 5141 1157 5147
rect 1172 5146 1173 5149
rect 1177 5145 1182 5150
rect 1209 5149 1212 5154
rect 1227 5150 1230 5154
rect 1227 5146 1228 5150
rect 1252 5149 1255 5154
rect 1273 5150 1276 5154
rect 1283 5150 1286 5154
rect 1089 5117 1092 5137
rect 1170 5117 1173 5137
rect 1209 5140 1212 5145
rect 1227 5140 1230 5146
rect 1247 5145 1250 5148
rect 1254 5145 1255 5149
rect 1267 5146 1276 5150
rect 1252 5140 1255 5145
rect 1273 5140 1276 5146
rect 1283 5140 1286 5146
rect 1299 5151 1302 5154
rect 1299 5147 1301 5151
rect 1327 5149 1330 5154
rect 1343 5150 1346 5154
rect 1299 5140 1302 5147
rect 1319 5147 1330 5149
rect 1319 5145 1320 5147
rect 1324 5145 1330 5147
rect 1338 5146 1340 5150
rect 1344 5146 1346 5150
rect 1327 5140 1330 5145
rect 1343 5140 1346 5146
rect 1352 5148 1355 5154
rect 1359 5148 1362 5154
rect 1609 5150 1612 5162
rect 1630 5150 1633 5162
rect 1646 5150 1649 5162
rect 1660 5156 1672 5159
rect 1688 5150 1691 5162
rect 1704 5150 1707 5162
rect 1725 5150 1728 5162
rect 2034 5161 2037 5179
rect 2115 5161 2118 5179
rect 2154 5172 2168 5176
rect 2172 5172 2233 5176
rect 2237 5172 2255 5176
rect 2259 5172 2286 5176
rect 2290 5172 2302 5176
rect 2360 5169 2560 5173
rect 2564 5169 2611 5173
rect 2615 5169 2661 5173
rect 2665 5169 2683 5173
rect 2173 5165 2175 5169
rect 2219 5165 2220 5169
rect 2244 5165 2247 5169
rect 2396 5162 2584 5166
rect 2588 5162 2612 5166
rect 2616 5162 2642 5166
rect 2646 5162 2683 5166
rect 2018 5150 2021 5153
rect 2099 5150 2102 5153
rect 1352 5145 1362 5148
rect 1370 5145 1372 5148
rect 1352 5140 1355 5145
rect 1359 5140 1362 5145
rect 1642 5140 1649 5143
rect 2013 5147 2021 5150
rect 1672 5140 1675 5146
rect 1700 5140 1707 5143
rect 1653 5136 1672 5139
rect 2018 5141 2021 5147
rect 2036 5146 2038 5149
rect 2042 5145 2047 5150
rect 2094 5147 2102 5150
rect 2099 5141 2102 5147
rect 2117 5146 2118 5149
rect 2122 5145 2127 5150
rect 2154 5149 2157 5154
rect 2172 5150 2175 5154
rect 2172 5146 2173 5150
rect 2197 5149 2200 5154
rect 2218 5150 2221 5154
rect 2228 5150 2231 5154
rect 1711 5136 1726 5139
rect 1604 5132 1613 5136
rect 1237 5127 1238 5131
rect 1284 5128 1285 5132
rect 1309 5127 1310 5131
rect 1626 5130 1631 5133
rect 1635 5130 1659 5133
rect 1209 5120 1238 5124
rect 1242 5120 1269 5124
rect 1273 5120 1294 5124
rect 1298 5120 1353 5124
rect 1357 5120 1433 5124
rect 1684 5130 1691 5133
rect 1695 5130 1717 5133
rect 1045 5113 1095 5117
rect 1099 5113 1119 5117
rect 1126 5113 1176 5117
rect 1180 5113 1200 5117
rect 1204 5113 1217 5117
rect 1221 5113 1245 5117
rect 1249 5113 1260 5117
rect 1264 5113 1294 5117
rect 1298 5113 1317 5117
rect 1321 5113 1326 5117
rect 1330 5113 1335 5117
rect 1339 5113 1353 5117
rect 1357 5113 1361 5117
rect 1365 5113 1367 5117
rect 1371 5113 1445 5117
rect 1059 5089 1062 5113
rect 1089 5085 1092 5113
rect 1096 5086 1101 5091
rect 1050 5080 1053 5085
rect 343 5067 386 5077
rect 1041 5077 1053 5080
rect 343 5057 376 5067
rect 1050 5063 1053 5077
rect 1061 5077 1064 5080
rect 1073 5075 1076 5081
rect 1096 5076 1099 5082
rect 1113 5081 1116 5113
rect 1140 5089 1143 5113
rect 1170 5085 1173 5113
rect 1177 5086 1182 5091
rect 1068 5072 1076 5075
rect 1088 5073 1099 5076
rect 1122 5080 1126 5084
rect 1131 5080 1134 5085
rect 1104 5072 1107 5077
rect 1126 5077 1134 5080
rect 1073 5069 1076 5072
rect 343 5047 366 5057
rect 1115 5069 1118 5072
rect 1122 5069 1123 5072
rect 1059 5051 1062 5055
rect 1089 5051 1092 5061
rect 1104 5063 1107 5068
rect 1131 5063 1134 5077
rect 1142 5077 1145 5080
rect 1154 5075 1157 5081
rect 1177 5076 1180 5082
rect 1194 5081 1197 5113
rect 1209 5106 1238 5110
rect 1242 5106 1269 5110
rect 1273 5106 1294 5110
rect 1298 5106 1353 5110
rect 1357 5106 1433 5110
rect 1609 5109 1612 5119
rect 1630 5109 1633 5119
rect 1646 5109 1649 5119
rect 1660 5112 1665 5116
rect 1669 5112 1676 5116
rect 1688 5109 1691 5119
rect 1704 5109 1707 5119
rect 1725 5109 1728 5119
rect 2034 5117 2037 5137
rect 2115 5117 2118 5137
rect 2154 5140 2157 5145
rect 2172 5140 2175 5146
rect 2192 5145 2195 5148
rect 2199 5145 2200 5149
rect 2212 5146 2221 5150
rect 2197 5140 2200 5145
rect 2218 5140 2221 5146
rect 2228 5140 2231 5146
rect 2244 5151 2247 5154
rect 2244 5147 2246 5151
rect 2272 5149 2275 5154
rect 2288 5150 2291 5154
rect 2244 5140 2247 5147
rect 2264 5147 2275 5149
rect 2264 5145 2265 5147
rect 2269 5145 2275 5147
rect 2283 5146 2285 5150
rect 2289 5146 2291 5150
rect 2272 5140 2275 5145
rect 2288 5140 2291 5146
rect 2297 5148 2300 5154
rect 2304 5148 2307 5154
rect 2554 5150 2557 5162
rect 2575 5150 2578 5162
rect 2591 5150 2594 5162
rect 2605 5156 2617 5159
rect 2633 5150 2636 5162
rect 2649 5150 2652 5162
rect 2670 5150 2673 5162
rect 2297 5145 2307 5148
rect 2315 5145 2317 5148
rect 2297 5140 2300 5145
rect 2304 5140 2307 5145
rect 2587 5140 2594 5143
rect 2617 5140 2620 5146
rect 2645 5140 2652 5143
rect 2598 5136 2617 5139
rect 2656 5136 2671 5139
rect 2549 5132 2558 5136
rect 2182 5127 2183 5131
rect 2229 5128 2230 5132
rect 2254 5127 2255 5131
rect 2571 5130 2576 5133
rect 2580 5130 2604 5133
rect 2154 5120 2183 5124
rect 2187 5120 2214 5124
rect 2218 5120 2239 5124
rect 2243 5120 2298 5124
rect 2302 5120 2378 5124
rect 2629 5130 2636 5133
rect 2640 5130 2662 5133
rect 1990 5113 2040 5117
rect 2044 5113 2064 5117
rect 2071 5113 2121 5117
rect 2125 5113 2145 5117
rect 2149 5113 2162 5117
rect 2166 5113 2190 5117
rect 2194 5113 2205 5117
rect 2209 5113 2239 5117
rect 2243 5113 2262 5117
rect 2266 5113 2271 5117
rect 2275 5113 2280 5117
rect 2284 5113 2298 5117
rect 2302 5113 2306 5117
rect 2310 5113 2312 5117
rect 2316 5113 2390 5117
rect 1463 5105 1639 5109
rect 1643 5105 1667 5109
rect 1671 5105 1697 5109
rect 1701 5105 1734 5109
rect 1237 5099 1238 5103
rect 1284 5098 1285 5102
rect 1309 5099 1310 5103
rect 1403 5098 1615 5102
rect 1619 5098 1651 5102
rect 1655 5098 1718 5102
rect 1722 5098 1738 5102
rect 1209 5085 1212 5090
rect 1227 5084 1230 5090
rect 1252 5085 1255 5090
rect 1149 5072 1157 5075
rect 1169 5073 1180 5076
rect 1185 5072 1188 5077
rect 1209 5076 1212 5081
rect 1227 5080 1228 5084
rect 1247 5082 1250 5085
rect 1254 5081 1255 5085
rect 1273 5084 1276 5090
rect 1283 5084 1286 5090
rect 1227 5076 1230 5080
rect 1252 5076 1255 5081
rect 1267 5080 1276 5084
rect 1273 5076 1276 5080
rect 1283 5076 1286 5080
rect 1154 5069 1157 5072
rect 1196 5069 1199 5072
rect 1299 5083 1302 5090
rect 1299 5079 1301 5083
rect 1319 5083 1320 5085
rect 1327 5085 1330 5090
rect 1324 5083 1330 5085
rect 1343 5084 1346 5090
rect 1319 5081 1330 5083
rect 1299 5076 1302 5079
rect 1327 5076 1330 5081
rect 1338 5080 1340 5084
rect 1344 5080 1346 5084
rect 1343 5076 1346 5080
rect 1352 5085 1355 5090
rect 1588 5090 1709 5094
rect 1721 5090 1725 5094
rect 1359 5085 1362 5090
rect 2004 5089 2007 5113
rect 1352 5082 1362 5085
rect 1352 5076 1355 5082
rect 1359 5076 1362 5082
rect 1370 5081 1584 5085
rect 1588 5081 1592 5085
rect 1604 5081 1608 5085
rect 1717 5083 1733 5087
rect 2034 5085 2037 5113
rect 2041 5086 2046 5091
rect 1995 5080 1998 5085
rect 1986 5077 1998 5080
rect 1113 5051 1116 5055
rect 1140 5051 1143 5055
rect 1170 5051 1173 5061
rect 1185 5063 1188 5068
rect 1228 5061 1230 5065
rect 1274 5061 1275 5065
rect 1299 5061 1302 5065
rect 1415 5067 1617 5071
rect 1621 5067 1667 5071
rect 1671 5067 1718 5071
rect 1722 5067 1731 5071
rect 1749 5069 1807 5073
rect 1451 5060 1636 5064
rect 1640 5060 1666 5064
rect 1670 5060 1694 5064
rect 1698 5060 1731 5064
rect 1194 5051 1197 5055
rect 1209 5054 1223 5058
rect 1227 5054 1288 5058
rect 1292 5054 1310 5058
rect 1314 5054 1341 5058
rect 1345 5054 1421 5058
rect 1022 5047 1041 5051
rect 1045 5047 1095 5051
rect 1099 5047 1122 5051
rect 1126 5047 1176 5051
rect 1180 5047 1200 5051
rect 1204 5047 1216 5051
rect 1220 5047 1244 5051
rect 1248 5047 1256 5051
rect 1260 5047 1261 5051
rect 1265 5047 1298 5051
rect 1302 5047 1317 5051
rect 1321 5047 1323 5051
rect 1327 5047 1334 5051
rect 1338 5047 1352 5051
rect 1356 5047 1368 5051
rect 1372 5047 1457 5051
rect 1609 5048 1612 5060
rect 1630 5048 1633 5060
rect 1646 5048 1649 5060
rect 1665 5054 1677 5057
rect 1688 5048 1691 5060
rect 1704 5048 1707 5060
rect 1725 5048 1728 5060
rect 1761 5056 1844 5064
rect 1995 5063 1998 5077
rect 2006 5077 2009 5080
rect 2018 5075 2021 5081
rect 2041 5076 2044 5082
rect 2058 5081 2061 5113
rect 2085 5089 2088 5113
rect 2115 5085 2118 5113
rect 2122 5086 2127 5091
rect 2013 5072 2021 5075
rect 2033 5073 2044 5076
rect 2067 5080 2071 5084
rect 2076 5080 2079 5085
rect 2049 5072 2052 5077
rect 2071 5077 2079 5080
rect 2018 5069 2021 5072
rect 2060 5069 2063 5072
rect 2067 5069 2068 5072
rect 2004 5051 2007 5055
rect 2034 5051 2037 5061
rect 2049 5063 2052 5068
rect 2076 5063 2079 5077
rect 2087 5077 2090 5080
rect 2099 5075 2102 5081
rect 2122 5076 2125 5082
rect 2139 5081 2142 5113
rect 2154 5106 2183 5110
rect 2187 5106 2214 5110
rect 2218 5106 2239 5110
rect 2243 5106 2298 5110
rect 2302 5106 2378 5110
rect 2554 5109 2557 5119
rect 2575 5109 2578 5119
rect 2591 5109 2594 5119
rect 2605 5112 2610 5116
rect 2614 5112 2621 5116
rect 2633 5109 2636 5119
rect 2649 5109 2652 5119
rect 2670 5109 2673 5119
rect 2408 5105 2584 5109
rect 2588 5105 2612 5109
rect 2616 5105 2642 5109
rect 2646 5105 2679 5109
rect 2182 5099 2183 5103
rect 2229 5098 2230 5102
rect 2254 5099 2255 5103
rect 2348 5098 2560 5102
rect 2564 5098 2596 5102
rect 2600 5098 2663 5102
rect 2667 5098 2683 5102
rect 2154 5085 2157 5090
rect 2172 5084 2175 5090
rect 2197 5085 2200 5090
rect 2094 5072 2102 5075
rect 2114 5073 2125 5076
rect 2130 5072 2133 5077
rect 2154 5076 2157 5081
rect 2172 5080 2173 5084
rect 2192 5082 2195 5085
rect 2199 5081 2200 5085
rect 2218 5084 2221 5090
rect 2228 5084 2231 5090
rect 2172 5076 2175 5080
rect 2197 5076 2200 5081
rect 2212 5080 2221 5084
rect 2218 5076 2221 5080
rect 2228 5076 2231 5080
rect 2099 5069 2102 5072
rect 2141 5069 2144 5072
rect 2244 5083 2247 5090
rect 2244 5079 2246 5083
rect 2264 5083 2265 5085
rect 2272 5085 2275 5090
rect 2269 5083 2275 5085
rect 2288 5084 2291 5090
rect 2264 5081 2275 5083
rect 2244 5076 2247 5079
rect 2272 5076 2275 5081
rect 2283 5080 2285 5084
rect 2289 5080 2291 5084
rect 2288 5076 2291 5080
rect 2297 5085 2300 5090
rect 2533 5090 2654 5094
rect 2666 5090 2670 5094
rect 2304 5085 2307 5090
rect 4403 5089 4829 5185
rect 2297 5082 2307 5085
rect 2297 5076 2300 5082
rect 2304 5076 2307 5082
rect 2315 5081 2529 5085
rect 2533 5081 2537 5085
rect 2549 5081 2553 5085
rect 2662 5083 2678 5087
rect 4786 5079 4829 5089
rect 2058 5051 2061 5055
rect 2085 5051 2088 5055
rect 2115 5051 2118 5061
rect 2130 5063 2133 5068
rect 2173 5061 2175 5065
rect 2219 5061 2220 5065
rect 2244 5061 2247 5065
rect 2360 5067 2562 5071
rect 2566 5067 2612 5071
rect 2616 5067 2663 5071
rect 2667 5067 2676 5071
rect 4796 5069 4829 5079
rect 2396 5060 2581 5064
rect 2585 5060 2611 5064
rect 2615 5060 2639 5064
rect 2643 5060 2676 5064
rect 2139 5051 2142 5055
rect 2154 5054 2168 5058
rect 2172 5054 2233 5058
rect 2237 5054 2255 5058
rect 2259 5054 2286 5058
rect 2290 5054 2366 5058
rect 343 5037 356 5047
rect 343 4998 346 5037
rect 851 5034 869 5038
rect 873 5034 919 5038
rect 923 5034 970 5038
rect 974 5034 1001 5038
rect 1005 5034 1051 5038
rect 1055 5034 1102 5038
rect 1106 5034 1133 5038
rect 1137 5034 1183 5038
rect 1187 5034 1234 5038
rect 1238 5034 1265 5038
rect 1269 5034 1315 5038
rect 1319 5034 1366 5038
rect 1370 5034 1409 5038
rect 1611 5034 1626 5037
rect 1630 5038 1637 5041
rect 1662 5038 1665 5044
rect 1967 5047 1986 5051
rect 1990 5047 2040 5051
rect 2044 5047 2067 5051
rect 2071 5047 2121 5051
rect 2125 5047 2145 5051
rect 2149 5047 2161 5051
rect 2165 5047 2189 5051
rect 2193 5047 2201 5051
rect 2205 5047 2206 5051
rect 2210 5047 2243 5051
rect 2247 5047 2262 5051
rect 2266 5047 2268 5051
rect 2272 5047 2279 5051
rect 2283 5047 2297 5051
rect 2301 5047 2313 5051
rect 2317 5047 2402 5051
rect 2554 5048 2557 5060
rect 2575 5048 2578 5060
rect 2591 5048 2594 5060
rect 2610 5054 2622 5057
rect 2633 5048 2636 5060
rect 2649 5048 2652 5060
rect 2670 5048 2673 5060
rect 4806 5059 4829 5069
rect 4816 5049 4829 5059
rect 1665 5034 1684 5037
rect 1688 5038 1695 5041
rect 1796 5034 1814 5038
rect 1818 5034 1864 5038
rect 1868 5034 1915 5038
rect 1919 5034 1946 5038
rect 1950 5034 1996 5038
rect 2000 5034 2047 5038
rect 2051 5034 2078 5038
rect 2082 5034 2128 5038
rect 2132 5034 2179 5038
rect 2183 5034 2210 5038
rect 2214 5034 2260 5038
rect 2264 5034 2311 5038
rect 2315 5034 2354 5038
rect 851 5027 888 5031
rect 892 5027 918 5031
rect 922 5027 946 5031
rect 950 5027 1020 5031
rect 1024 5027 1050 5031
rect 1054 5027 1078 5031
rect 1082 5027 1152 5031
rect 1156 5027 1182 5031
rect 1186 5027 1210 5031
rect 1214 5027 1284 5031
rect 1288 5027 1314 5031
rect 1318 5027 1342 5031
rect 1346 5027 1445 5031
rect 861 5015 864 5027
rect 882 5015 885 5027
rect 898 5015 901 5027
rect 917 5021 929 5024
rect 940 5015 943 5027
rect 956 5015 959 5027
rect 977 5015 980 5027
rect 861 5001 878 5004
rect 882 5005 889 5008
rect 914 5005 917 5011
rect 993 5015 996 5027
rect 1014 5015 1017 5027
rect 1030 5015 1033 5027
rect 1049 5021 1061 5024
rect 1072 5015 1075 5027
rect 1088 5015 1091 5027
rect 1109 5015 1112 5027
rect 1125 5015 1128 5027
rect 1146 5015 1149 5027
rect 1162 5015 1165 5027
rect 1181 5021 1193 5024
rect 1204 5015 1207 5027
rect 1220 5015 1223 5027
rect 1241 5015 1244 5027
rect 1257 5015 1260 5027
rect 1278 5015 1281 5027
rect 1294 5015 1297 5027
rect 1313 5021 1325 5024
rect 1336 5015 1339 5027
rect 1352 5015 1355 5027
rect 1373 5015 1376 5027
rect 1620 5028 1642 5031
rect 1646 5028 1653 5031
rect 1678 5028 1702 5031
rect 1706 5028 1711 5031
rect 1724 5030 1733 5034
rect 2556 5034 2571 5037
rect 2575 5038 2582 5041
rect 2607 5038 2610 5044
rect 2610 5034 2629 5037
rect 2633 5038 2640 5041
rect 1796 5027 1833 5031
rect 1837 5027 1863 5031
rect 1867 5027 1891 5031
rect 1895 5027 1965 5031
rect 1969 5027 1995 5031
rect 1999 5027 2023 5031
rect 2027 5027 2097 5031
rect 2101 5027 2127 5031
rect 2131 5027 2155 5031
rect 2159 5027 2229 5031
rect 2233 5027 2259 5031
rect 2263 5027 2287 5031
rect 2291 5027 2390 5031
rect 917 5001 936 5004
rect 940 5005 947 5008
rect 86 4995 346 4998
rect 872 4995 894 4998
rect 898 4995 905 4998
rect 930 4995 954 4998
rect 958 4995 963 4998
rect 993 5001 1010 5004
rect 1014 5005 1021 5008
rect 1046 5005 1049 5011
rect 1049 5001 1068 5004
rect 1072 5005 1079 5008
rect 1004 4995 1026 4998
rect 1030 4995 1037 4998
rect 1062 4995 1086 4998
rect 1090 4995 1095 4998
rect 1125 5001 1142 5004
rect 1146 5005 1153 5008
rect 1178 5005 1181 5011
rect 1181 5001 1200 5004
rect 1204 5005 1211 5008
rect 1136 4995 1158 4998
rect 1162 4995 1169 4998
rect 1194 4995 1218 4998
rect 1222 4995 1227 4998
rect 1257 5001 1274 5004
rect 1278 5005 1285 5008
rect 1310 5005 1313 5011
rect 1313 5001 1332 5004
rect 1336 5005 1343 5008
rect 1609 5007 1612 5017
rect 1630 5007 1633 5017
rect 1646 5007 1649 5017
rect 1661 5010 1668 5014
rect 1672 5010 1677 5014
rect 1688 5007 1691 5017
rect 1704 5007 1707 5017
rect 1725 5007 1728 5017
rect 1806 5015 1809 5027
rect 1827 5015 1830 5027
rect 1843 5015 1846 5027
rect 1862 5021 1874 5024
rect 1885 5015 1888 5027
rect 1901 5015 1904 5027
rect 1922 5015 1925 5027
rect 1463 5003 1599 5007
rect 1603 5003 1636 5007
rect 1640 5003 1666 5007
rect 1670 5003 1694 5007
rect 1698 5003 1731 5007
rect 1268 4995 1290 4998
rect 1294 4995 1301 4998
rect 1326 4995 1350 4998
rect 1354 4995 1359 4998
rect 1806 5001 1823 5004
rect 1827 5005 1834 5008
rect 1859 5005 1862 5011
rect 1938 5015 1941 5027
rect 1959 5015 1962 5027
rect 1975 5015 1978 5027
rect 1994 5021 2006 5024
rect 2017 5015 2020 5027
rect 2033 5015 2036 5027
rect 2054 5015 2057 5027
rect 2070 5015 2073 5027
rect 2091 5015 2094 5027
rect 2107 5015 2110 5027
rect 2126 5021 2138 5024
rect 2149 5015 2152 5027
rect 2165 5015 2168 5027
rect 2186 5015 2189 5027
rect 2202 5015 2205 5027
rect 2223 5015 2226 5027
rect 2239 5015 2242 5027
rect 2258 5021 2270 5024
rect 2281 5015 2284 5027
rect 2297 5015 2300 5027
rect 2318 5015 2321 5027
rect 2565 5028 2587 5031
rect 2591 5028 2598 5031
rect 2623 5028 2647 5031
rect 2651 5028 2656 5031
rect 2669 5030 2678 5034
rect 1862 5001 1881 5004
rect 1885 5005 1892 5008
rect 1403 4996 1615 5000
rect 1619 4996 1682 5000
rect 1686 4996 1718 5000
rect 1722 4996 1731 5000
rect 1817 4995 1839 4998
rect 1843 4995 1850 4998
rect 1875 4995 1899 4998
rect 1903 4995 1908 4998
rect 1938 5001 1955 5004
rect 1959 5005 1966 5008
rect 1991 5005 1994 5011
rect 1994 5001 2013 5004
rect 2017 5005 2024 5008
rect 1949 4995 1971 4998
rect 1975 4995 1982 4998
rect 2007 4995 2031 4998
rect 2035 4995 2040 4998
rect 2070 5001 2087 5004
rect 2091 5005 2098 5008
rect 2123 5005 2126 5011
rect 2126 5001 2145 5004
rect 2149 5005 2156 5008
rect 2081 4995 2103 4998
rect 2107 4995 2114 4998
rect 2139 4995 2163 4998
rect 2167 4995 2172 4998
rect 2202 5001 2219 5004
rect 2223 5005 2230 5008
rect 2255 5005 2258 5011
rect 2258 5001 2277 5004
rect 2281 5005 2288 5008
rect 2554 5007 2557 5017
rect 2575 5007 2578 5017
rect 2591 5007 2594 5017
rect 2606 5010 2613 5014
rect 2617 5010 2622 5014
rect 2633 5007 2636 5017
rect 2649 5007 2652 5017
rect 2670 5007 2673 5017
rect 4826 5010 4829 5049
rect 5083 5010 5086 5264
rect 2408 5003 2544 5007
rect 2548 5003 2581 5007
rect 2585 5003 2611 5007
rect 2615 5003 2639 5007
rect 2643 5003 2676 5007
rect 4483 5004 4484 5008
rect 4488 5004 4489 5008
rect 4493 5004 4494 5008
rect 4498 5004 4499 5008
rect 4503 5004 4504 5008
rect 4508 5004 4509 5008
rect 4479 5003 4513 5004
rect 2213 4995 2235 4998
rect 2239 4995 2246 4998
rect 2271 4995 2295 4998
rect 2299 4995 2304 4998
rect 2348 4996 2560 5000
rect 2564 4996 2627 5000
rect 2631 4996 2663 5000
rect 2667 4996 2676 5000
rect 4483 4999 4484 5003
rect 4488 4999 4489 5003
rect 4493 4999 4494 5003
rect 4498 4999 4499 5003
rect 4503 4999 4504 5003
rect 4508 4999 4509 5003
rect 4479 4998 4513 4999
rect 4483 4994 4484 4998
rect 4488 4994 4489 4998
rect 4493 4994 4494 4998
rect 4498 4994 4499 4998
rect 4503 4994 4504 4998
rect 4508 4994 4509 4998
rect 4479 4993 4513 4994
rect 4483 4989 4484 4993
rect 4488 4989 4489 4993
rect 4493 4989 4494 4993
rect 4498 4989 4499 4993
rect 4503 4989 4504 4993
rect 4508 4989 4509 4993
rect 4529 5004 4530 5008
rect 4534 5004 4535 5008
rect 4539 5004 4540 5008
rect 4544 5004 4545 5008
rect 4549 5004 4550 5008
rect 4554 5004 4555 5008
rect 4826 5007 5086 5010
rect 4525 5003 4559 5004
rect 4529 4999 4530 5003
rect 4534 4999 4535 5003
rect 4539 4999 4540 5003
rect 4544 4999 4545 5003
rect 4549 4999 4550 5003
rect 4554 4999 4555 5003
rect 4525 4998 4559 4999
rect 4529 4994 4530 4998
rect 4534 4994 4535 4998
rect 4539 4994 4540 4998
rect 4544 4994 4545 4998
rect 4549 4994 4550 4998
rect 4554 4994 4555 4998
rect 4525 4993 4559 4994
rect 4529 4989 4530 4993
rect 4534 4989 4535 4993
rect 4539 4989 4540 4993
rect 4544 4989 4545 4993
rect 4549 4989 4550 4993
rect 4554 4989 4555 4993
rect 861 4974 864 4984
rect 882 4974 885 4984
rect 898 4974 901 4984
rect 913 4977 920 4981
rect 924 4977 929 4981
rect 940 4974 943 4984
rect 956 4974 959 4984
rect 977 4974 980 4984
rect 993 4974 996 4984
rect 1014 4974 1017 4984
rect 1030 4974 1033 4984
rect 1045 4977 1052 4981
rect 1056 4977 1061 4981
rect 1072 4974 1075 4984
rect 1088 4974 1091 4984
rect 1109 4974 1112 4984
rect 1125 4974 1128 4984
rect 1146 4974 1149 4984
rect 1162 4974 1165 4984
rect 1177 4977 1184 4981
rect 1188 4977 1193 4981
rect 1204 4974 1207 4984
rect 1220 4974 1223 4984
rect 1241 4974 1244 4984
rect 1257 4974 1260 4984
rect 1278 4974 1281 4984
rect 1294 4974 1297 4984
rect 1309 4977 1316 4981
rect 1320 4977 1325 4981
rect 1336 4974 1339 4984
rect 1352 4974 1355 4984
rect 1373 4974 1376 4984
rect 1806 4974 1809 4984
rect 1827 4974 1830 4984
rect 1843 4974 1846 4984
rect 1858 4977 1865 4981
rect 1869 4977 1874 4981
rect 1885 4974 1888 4984
rect 1901 4974 1904 4984
rect 1922 4974 1925 4984
rect 1938 4974 1941 4984
rect 1959 4974 1962 4984
rect 1975 4974 1978 4984
rect 1990 4977 1997 4981
rect 2001 4977 2006 4981
rect 2017 4974 2020 4984
rect 2033 4974 2036 4984
rect 2054 4974 2057 4984
rect 2070 4974 2073 4984
rect 2091 4974 2094 4984
rect 2107 4974 2110 4984
rect 2122 4977 2129 4981
rect 2133 4977 2138 4981
rect 2149 4974 2152 4984
rect 2165 4974 2168 4984
rect 2186 4974 2189 4984
rect 2202 4974 2205 4984
rect 2223 4974 2226 4984
rect 2239 4974 2242 4984
rect 2254 4977 2261 4981
rect 2265 4977 2270 4981
rect 2281 4974 2284 4984
rect 2297 4974 2300 4984
rect 2318 4974 2321 4984
rect 855 4970 888 4974
rect 892 4970 918 4974
rect 922 4970 946 4974
rect 950 4970 983 4974
rect 987 4970 1020 4974
rect 1024 4970 1050 4974
rect 1054 4970 1078 4974
rect 1082 4970 1115 4974
rect 1119 4970 1152 4974
rect 1156 4970 1182 4974
rect 1186 4970 1210 4974
rect 1214 4970 1247 4974
rect 1251 4970 1284 4974
rect 1288 4970 1314 4974
rect 1318 4970 1342 4974
rect 1346 4970 1457 4974
rect 1800 4970 1833 4974
rect 1837 4970 1863 4974
rect 1867 4970 1891 4974
rect 1895 4970 1928 4974
rect 1932 4970 1965 4974
rect 1969 4970 1995 4974
rect 1999 4970 2023 4974
rect 2027 4970 2060 4974
rect 2064 4970 2097 4974
rect 2101 4970 2127 4974
rect 2131 4970 2155 4974
rect 2159 4970 2192 4974
rect 2196 4970 2229 4974
rect 2233 4970 2259 4974
rect 2263 4970 2287 4974
rect 2291 4970 2402 4974
rect 851 4963 867 4967
rect 871 4963 934 4967
rect 938 4963 970 4967
rect 974 4963 999 4967
rect 1003 4963 1066 4967
rect 1070 4963 1102 4967
rect 1106 4963 1131 4967
rect 1135 4963 1198 4967
rect 1202 4963 1234 4967
rect 1238 4963 1263 4967
rect 1267 4963 1330 4967
rect 1334 4963 1366 4967
rect 1370 4963 1397 4967
rect 1796 4963 1812 4967
rect 1816 4963 1879 4967
rect 1883 4963 1915 4967
rect 1919 4963 1944 4967
rect 1948 4963 2011 4967
rect 2015 4963 2047 4967
rect 2051 4963 2076 4967
rect 2080 4963 2143 4967
rect 2147 4963 2179 4967
rect 2183 4963 2208 4967
rect 2212 4963 2275 4967
rect 2279 4963 2311 4967
rect 2315 4963 2342 4967
rect 99 4528 593 4959
rect 2674 4932 3836 4936
rect 3844 4932 3847 4936
rect 1761 4876 2146 4880
rect 617 4868 618 4872
rect 622 4868 623 4872
rect 627 4868 628 4872
rect 632 4868 633 4872
rect 637 4868 638 4872
rect 642 4868 643 4872
rect 613 4867 647 4868
rect 617 4863 618 4867
rect 622 4863 623 4867
rect 627 4863 628 4867
rect 632 4863 633 4867
rect 637 4863 638 4867
rect 642 4863 643 4867
rect 613 4862 647 4863
rect 617 4858 618 4862
rect 622 4858 623 4862
rect 627 4858 628 4862
rect 632 4858 633 4862
rect 637 4858 638 4862
rect 642 4858 643 4862
rect 613 4857 647 4858
rect 617 4853 618 4857
rect 622 4853 623 4857
rect 627 4853 628 4857
rect 632 4853 633 4857
rect 637 4853 638 4857
rect 642 4853 643 4857
rect 663 4868 664 4872
rect 668 4868 669 4872
rect 673 4868 674 4872
rect 678 4868 679 4872
rect 683 4868 684 4872
rect 688 4868 689 4872
rect 659 4867 693 4868
rect 663 4863 664 4867
rect 668 4863 669 4867
rect 673 4863 674 4867
rect 678 4863 679 4867
rect 683 4863 684 4867
rect 688 4863 689 4867
rect 1749 4866 2119 4870
rect 659 4862 693 4863
rect 663 4858 664 4862
rect 668 4858 669 4862
rect 673 4858 674 4862
rect 678 4858 679 4862
rect 683 4858 684 4862
rect 688 4858 689 4862
rect 659 4857 693 4858
rect 663 4853 664 4857
rect 668 4853 669 4857
rect 673 4853 674 4857
rect 678 4853 679 4857
rect 683 4853 684 4857
rect 688 4853 689 4857
rect 1192 4858 1385 4862
rect 1391 4858 2330 4862
rect 617 4839 618 4843
rect 622 4839 623 4843
rect 627 4839 628 4843
rect 632 4839 633 4843
rect 637 4839 638 4843
rect 642 4839 643 4843
rect 613 4838 647 4839
rect 617 4834 618 4838
rect 622 4834 623 4838
rect 627 4834 628 4838
rect 632 4834 633 4838
rect 637 4834 638 4838
rect 642 4834 643 4838
rect 613 4833 647 4834
rect 617 4829 618 4833
rect 622 4829 623 4833
rect 627 4829 628 4833
rect 632 4829 633 4833
rect 637 4829 638 4833
rect 642 4829 643 4833
rect 613 4828 647 4829
rect 617 4824 618 4828
rect 622 4824 623 4828
rect 627 4824 628 4828
rect 632 4824 633 4828
rect 637 4824 638 4828
rect 642 4824 643 4828
rect 663 4839 664 4843
rect 668 4839 669 4843
rect 673 4839 674 4843
rect 678 4839 679 4843
rect 683 4839 684 4843
rect 688 4839 689 4843
rect 659 4838 693 4839
rect 663 4834 664 4838
rect 668 4834 669 4838
rect 673 4834 674 4838
rect 678 4834 679 4838
rect 683 4834 684 4838
rect 688 4834 689 4838
rect 659 4833 693 4834
rect 663 4829 664 4833
rect 668 4829 669 4833
rect 673 4829 674 4833
rect 678 4829 679 4833
rect 683 4829 684 4833
rect 688 4829 689 4833
rect 659 4828 693 4829
rect 663 4824 664 4828
rect 668 4824 669 4828
rect 673 4824 674 4828
rect 678 4824 679 4828
rect 683 4824 684 4828
rect 688 4824 689 4828
rect 617 4810 618 4814
rect 622 4810 623 4814
rect 627 4810 628 4814
rect 632 4810 633 4814
rect 637 4810 638 4814
rect 642 4810 643 4814
rect 613 4809 647 4810
rect 617 4805 618 4809
rect 622 4805 623 4809
rect 627 4805 628 4809
rect 632 4805 633 4809
rect 637 4805 638 4809
rect 642 4805 643 4809
rect 613 4804 647 4805
rect 617 4800 618 4804
rect 622 4800 623 4804
rect 627 4800 628 4804
rect 632 4800 633 4804
rect 637 4800 638 4804
rect 642 4800 643 4804
rect 613 4799 647 4800
rect 617 4795 618 4799
rect 622 4795 623 4799
rect 627 4795 628 4799
rect 632 4795 633 4799
rect 637 4795 638 4799
rect 642 4795 643 4799
rect 663 4810 664 4814
rect 668 4810 669 4814
rect 673 4810 674 4814
rect 678 4810 679 4814
rect 683 4810 684 4814
rect 688 4810 689 4814
rect 659 4809 693 4810
rect 663 4805 664 4809
rect 668 4805 669 4809
rect 673 4805 674 4809
rect 678 4805 679 4809
rect 683 4805 684 4809
rect 688 4805 689 4809
rect 659 4804 693 4805
rect 663 4800 664 4804
rect 668 4800 669 4804
rect 673 4800 674 4804
rect 678 4800 679 4804
rect 683 4800 684 4804
rect 688 4800 689 4804
rect 659 4799 693 4800
rect 663 4795 664 4799
rect 668 4795 669 4799
rect 673 4795 674 4799
rect 678 4795 679 4799
rect 683 4795 684 4799
rect 688 4795 689 4799
rect 617 4781 618 4785
rect 622 4781 623 4785
rect 627 4781 628 4785
rect 632 4781 633 4785
rect 637 4781 638 4785
rect 642 4781 643 4785
rect 613 4780 647 4781
rect 617 4776 618 4780
rect 622 4776 623 4780
rect 627 4776 628 4780
rect 632 4776 633 4780
rect 637 4776 638 4780
rect 642 4776 643 4780
rect 613 4775 647 4776
rect 617 4771 618 4775
rect 622 4771 623 4775
rect 627 4771 628 4775
rect 632 4771 633 4775
rect 637 4771 638 4775
rect 642 4771 643 4775
rect 613 4770 647 4771
rect 617 4766 618 4770
rect 622 4766 623 4770
rect 627 4766 628 4770
rect 632 4766 633 4770
rect 637 4766 638 4770
rect 642 4766 643 4770
rect 663 4781 664 4785
rect 668 4781 669 4785
rect 673 4781 674 4785
rect 678 4781 679 4785
rect 683 4781 684 4785
rect 688 4781 689 4785
rect 659 4780 693 4781
rect 663 4776 664 4780
rect 668 4776 669 4780
rect 673 4776 674 4780
rect 678 4776 679 4780
rect 683 4776 684 4780
rect 688 4776 689 4780
rect 659 4775 693 4776
rect 663 4771 664 4775
rect 668 4771 669 4775
rect 673 4771 674 4775
rect 678 4771 679 4775
rect 683 4771 684 4775
rect 688 4771 689 4775
rect 659 4770 693 4771
rect 663 4766 664 4770
rect 668 4766 669 4770
rect 673 4766 674 4770
rect 678 4766 679 4770
rect 683 4766 684 4770
rect 688 4766 689 4770
rect 617 4752 618 4756
rect 622 4752 623 4756
rect 627 4752 628 4756
rect 632 4752 633 4756
rect 637 4752 638 4756
rect 642 4752 643 4756
rect 613 4751 647 4752
rect 617 4747 618 4751
rect 622 4747 623 4751
rect 627 4747 628 4751
rect 632 4747 633 4751
rect 637 4747 638 4751
rect 642 4747 643 4751
rect 613 4746 647 4747
rect 617 4742 618 4746
rect 622 4742 623 4746
rect 627 4742 628 4746
rect 632 4742 633 4746
rect 637 4742 638 4746
rect 642 4742 643 4746
rect 613 4741 647 4742
rect 617 4737 618 4741
rect 622 4737 623 4741
rect 627 4737 628 4741
rect 632 4737 633 4741
rect 637 4737 638 4741
rect 642 4737 643 4741
rect 663 4752 664 4756
rect 668 4752 669 4756
rect 673 4752 674 4756
rect 678 4752 679 4756
rect 683 4752 684 4756
rect 688 4752 689 4756
rect 659 4751 693 4752
rect 663 4747 664 4751
rect 668 4747 669 4751
rect 673 4747 674 4751
rect 678 4747 679 4751
rect 683 4747 684 4751
rect 688 4747 689 4751
rect 659 4746 693 4747
rect 663 4742 664 4746
rect 668 4742 669 4746
rect 673 4742 674 4746
rect 678 4742 679 4746
rect 683 4742 684 4746
rect 688 4742 689 4746
rect 659 4741 693 4742
rect 663 4737 664 4741
rect 668 4737 669 4741
rect 673 4737 674 4741
rect 678 4737 679 4741
rect 683 4737 684 4741
rect 688 4737 689 4741
rect 1192 4740 1204 4858
rect 1474 4854 1482 4855
rect 1384 4850 1457 4854
rect 1463 4851 1482 4854
rect 1537 4851 2402 4855
rect 1463 4850 1480 4851
rect 1384 4843 1445 4847
rect 1451 4843 1790 4847
rect 1845 4843 2390 4847
rect 1439 4835 2378 4839
rect 1427 4828 2366 4832
rect 1415 4821 2354 4825
rect 1403 4813 2342 4817
rect 4483 4811 4484 4815
rect 4488 4811 4489 4815
rect 4493 4811 4494 4815
rect 4498 4811 4499 4815
rect 4503 4811 4504 4815
rect 4508 4811 4509 4815
rect 4479 4810 4513 4811
rect 4483 4806 4484 4810
rect 4488 4806 4489 4810
rect 4493 4806 4494 4810
rect 4498 4806 4499 4810
rect 4503 4806 4504 4810
rect 4508 4806 4509 4810
rect 4479 4805 4513 4806
rect 4483 4801 4484 4805
rect 4488 4801 4489 4805
rect 4493 4801 4494 4805
rect 4498 4801 4499 4805
rect 4503 4801 4504 4805
rect 4508 4801 4509 4805
rect 4479 4800 4513 4801
rect 4483 4796 4484 4800
rect 4488 4796 4489 4800
rect 4493 4796 4494 4800
rect 4498 4796 4499 4800
rect 4503 4796 4504 4800
rect 4508 4796 4509 4800
rect 4529 4811 4530 4815
rect 4534 4811 4535 4815
rect 4539 4811 4540 4815
rect 4544 4811 4545 4815
rect 4549 4811 4550 4815
rect 4554 4811 4555 4815
rect 4525 4810 4559 4811
rect 4529 4806 4530 4810
rect 4534 4806 4535 4810
rect 4539 4806 4540 4810
rect 4544 4806 4545 4810
rect 4549 4806 4550 4810
rect 4554 4806 4555 4810
rect 4525 4805 4559 4806
rect 4529 4801 4530 4805
rect 4534 4801 4535 4805
rect 4539 4801 4540 4805
rect 4544 4801 4545 4805
rect 4549 4801 4550 4805
rect 4554 4801 4555 4805
rect 4525 4800 4559 4801
rect 4529 4796 4530 4800
rect 4534 4796 4535 4800
rect 4539 4796 4540 4800
rect 4544 4796 4545 4800
rect 4549 4796 4550 4800
rect 4554 4796 4555 4800
rect 4483 4785 4484 4789
rect 4488 4785 4489 4789
rect 4493 4785 4494 4789
rect 4498 4785 4499 4789
rect 4503 4785 4504 4789
rect 4508 4785 4509 4789
rect 4479 4784 4513 4785
rect 4483 4780 4484 4784
rect 4488 4780 4489 4784
rect 4493 4780 4494 4784
rect 4498 4780 4499 4784
rect 4503 4780 4504 4784
rect 4508 4780 4509 4784
rect 4479 4779 4513 4780
rect 4483 4775 4484 4779
rect 4488 4775 4489 4779
rect 4493 4775 4494 4779
rect 4498 4775 4499 4779
rect 4503 4775 4504 4779
rect 4508 4775 4509 4779
rect 4479 4774 4513 4775
rect 4483 4770 4484 4774
rect 4488 4770 4489 4774
rect 4493 4770 4494 4774
rect 4498 4770 4499 4774
rect 4503 4770 4504 4774
rect 4508 4770 4509 4774
rect 4529 4785 4530 4789
rect 4534 4785 4535 4789
rect 4539 4785 4540 4789
rect 4544 4785 4545 4789
rect 4549 4785 4550 4789
rect 4554 4785 4555 4789
rect 4525 4784 4559 4785
rect 4529 4780 4530 4784
rect 4534 4780 4535 4784
rect 4539 4780 4540 4784
rect 4544 4780 4545 4784
rect 4549 4780 4550 4784
rect 4554 4780 4555 4784
rect 4525 4779 4559 4780
rect 4529 4775 4530 4779
rect 4534 4775 4535 4779
rect 4539 4775 4540 4779
rect 4544 4775 4545 4779
rect 4549 4775 4550 4779
rect 4554 4775 4555 4779
rect 4525 4774 4559 4775
rect 4529 4770 4530 4774
rect 4534 4770 4535 4774
rect 4539 4770 4540 4774
rect 4544 4770 4545 4774
rect 4549 4770 4550 4774
rect 4554 4770 4555 4774
rect 4483 4759 4484 4763
rect 4488 4759 4489 4763
rect 4493 4759 4494 4763
rect 4498 4759 4499 4763
rect 4503 4759 4504 4763
rect 4508 4759 4509 4763
rect 4479 4758 4513 4759
rect 4483 4754 4484 4758
rect 4488 4754 4489 4758
rect 4493 4754 4494 4758
rect 4498 4754 4499 4758
rect 4503 4754 4504 4758
rect 4508 4754 4509 4758
rect 4479 4753 4513 4754
rect 4483 4749 4484 4753
rect 4488 4749 4489 4753
rect 4493 4749 4494 4753
rect 4498 4749 4499 4753
rect 4503 4749 4504 4753
rect 4508 4749 4509 4753
rect 4479 4748 4513 4749
rect 4483 4744 4484 4748
rect 4488 4744 4489 4748
rect 4493 4744 4494 4748
rect 4498 4744 4499 4748
rect 4503 4744 4504 4748
rect 4508 4744 4509 4748
rect 4529 4759 4530 4763
rect 4534 4759 4535 4763
rect 4539 4759 4540 4763
rect 4544 4759 4545 4763
rect 4549 4759 4550 4763
rect 4554 4759 4555 4763
rect 4525 4758 4559 4759
rect 4529 4754 4530 4758
rect 4534 4754 4535 4758
rect 4539 4754 4540 4758
rect 4544 4754 4545 4758
rect 4549 4754 4550 4758
rect 4554 4754 4555 4758
rect 4525 4753 4559 4754
rect 4529 4749 4530 4753
rect 4534 4749 4535 4753
rect 4539 4749 4540 4753
rect 4544 4749 4545 4753
rect 4549 4749 4550 4753
rect 4554 4749 4555 4753
rect 4525 4748 4559 4749
rect 4529 4744 4530 4748
rect 4534 4744 4535 4748
rect 4539 4744 4540 4748
rect 4544 4744 4545 4748
rect 4549 4744 4550 4748
rect 4554 4744 4555 4748
rect 761 4624 762 4628
rect 766 4624 767 4628
rect 771 4624 772 4628
rect 757 4623 776 4624
rect 761 4619 762 4623
rect 766 4619 767 4623
rect 771 4619 772 4623
rect 757 4618 776 4619
rect 761 4614 762 4618
rect 766 4614 767 4618
rect 771 4614 772 4618
rect 757 4613 776 4614
rect 761 4609 762 4613
rect 766 4609 767 4613
rect 771 4609 772 4613
rect 757 4608 776 4609
rect 761 4604 762 4608
rect 766 4604 767 4608
rect 771 4604 772 4608
rect 757 4603 776 4604
rect 761 4599 762 4603
rect 766 4599 767 4603
rect 771 4599 772 4603
rect 757 4598 776 4599
rect 761 4594 762 4598
rect 766 4594 767 4598
rect 771 4594 772 4598
rect 787 4624 788 4628
rect 792 4624 793 4628
rect 797 4624 798 4628
rect 783 4623 802 4624
rect 787 4619 788 4623
rect 792 4619 793 4623
rect 797 4619 798 4623
rect 783 4618 802 4619
rect 787 4614 788 4618
rect 792 4614 793 4618
rect 797 4614 798 4618
rect 783 4613 802 4614
rect 787 4609 788 4613
rect 792 4609 793 4613
rect 797 4609 798 4613
rect 783 4608 802 4609
rect 787 4604 788 4608
rect 792 4604 793 4608
rect 797 4604 798 4608
rect 783 4603 802 4604
rect 787 4599 788 4603
rect 792 4599 793 4603
rect 797 4599 798 4603
rect 783 4598 802 4599
rect 787 4594 788 4598
rect 792 4594 793 4598
rect 797 4594 798 4598
rect 813 4624 814 4628
rect 818 4624 819 4628
rect 823 4624 824 4628
rect 809 4623 828 4624
rect 813 4619 814 4623
rect 818 4619 819 4623
rect 823 4619 824 4623
rect 809 4618 828 4619
rect 813 4614 814 4618
rect 818 4614 819 4618
rect 823 4614 824 4618
rect 809 4613 828 4614
rect 813 4609 814 4613
rect 818 4609 819 4613
rect 823 4609 824 4613
rect 809 4608 828 4609
rect 813 4604 814 4608
rect 818 4604 819 4608
rect 823 4604 824 4608
rect 809 4603 828 4604
rect 813 4599 814 4603
rect 818 4599 819 4603
rect 823 4599 824 4603
rect 809 4598 828 4599
rect 813 4594 814 4598
rect 818 4594 819 4598
rect 823 4594 824 4598
rect 839 4624 840 4628
rect 844 4624 845 4628
rect 849 4624 850 4628
rect 835 4623 854 4624
rect 839 4619 840 4623
rect 844 4619 845 4623
rect 849 4619 850 4623
rect 835 4618 854 4619
rect 839 4614 840 4618
rect 844 4614 845 4618
rect 849 4614 850 4618
rect 835 4613 854 4614
rect 839 4609 840 4613
rect 844 4609 845 4613
rect 849 4609 850 4613
rect 835 4608 854 4609
rect 839 4604 840 4608
rect 844 4604 845 4608
rect 849 4604 850 4608
rect 835 4603 854 4604
rect 839 4599 840 4603
rect 844 4599 845 4603
rect 849 4599 850 4603
rect 835 4598 854 4599
rect 839 4594 840 4598
rect 844 4594 845 4598
rect 849 4594 850 4598
rect 865 4624 866 4628
rect 870 4624 871 4628
rect 875 4624 876 4628
rect 861 4623 880 4624
rect 865 4619 866 4623
rect 870 4619 871 4623
rect 875 4619 876 4623
rect 861 4618 880 4619
rect 865 4614 866 4618
rect 870 4614 871 4618
rect 875 4614 876 4618
rect 861 4613 880 4614
rect 865 4609 866 4613
rect 870 4609 871 4613
rect 875 4609 876 4613
rect 861 4608 880 4609
rect 865 4604 866 4608
rect 870 4604 871 4608
rect 875 4604 876 4608
rect 861 4603 880 4604
rect 865 4599 866 4603
rect 870 4599 871 4603
rect 875 4599 876 4603
rect 861 4598 880 4599
rect 865 4594 866 4598
rect 870 4594 871 4598
rect 875 4594 876 4598
rect 1057 4624 1058 4628
rect 1062 4624 1063 4628
rect 1067 4624 1068 4628
rect 1053 4623 1072 4624
rect 1057 4619 1058 4623
rect 1062 4619 1063 4623
rect 1067 4619 1068 4623
rect 1053 4618 1072 4619
rect 1057 4614 1058 4618
rect 1062 4614 1063 4618
rect 1067 4614 1068 4618
rect 1053 4613 1072 4614
rect 1057 4609 1058 4613
rect 1062 4609 1063 4613
rect 1067 4609 1068 4613
rect 1053 4608 1072 4609
rect 1057 4604 1058 4608
rect 1062 4604 1063 4608
rect 1067 4604 1068 4608
rect 1053 4603 1072 4604
rect 1057 4599 1058 4603
rect 1062 4599 1063 4603
rect 1067 4599 1068 4603
rect 1053 4598 1072 4599
rect 1057 4594 1058 4598
rect 1062 4594 1063 4598
rect 1067 4594 1068 4598
rect 1075 4601 1131 4602
rect 1075 4597 1077 4601
rect 1081 4597 1082 4601
rect 1086 4597 1087 4601
rect 1091 4597 1092 4601
rect 1096 4597 1097 4601
rect 1101 4597 1102 4601
rect 1106 4597 1107 4601
rect 1111 4597 1112 4601
rect 1116 4597 1117 4601
rect 1121 4597 1122 4601
rect 1126 4597 1127 4601
rect 1075 4596 1131 4597
rect 1075 4592 1077 4596
rect 1081 4592 1082 4596
rect 1086 4592 1087 4596
rect 1091 4592 1092 4596
rect 1096 4592 1097 4596
rect 1101 4592 1102 4596
rect 1106 4592 1107 4596
rect 1111 4592 1112 4596
rect 1116 4592 1117 4596
rect 1121 4592 1122 4596
rect 1126 4592 1127 4596
rect 761 4578 762 4582
rect 766 4578 767 4582
rect 771 4578 772 4582
rect 757 4577 776 4578
rect 761 4573 762 4577
rect 766 4573 767 4577
rect 771 4573 772 4577
rect 757 4572 776 4573
rect 761 4568 762 4572
rect 766 4568 767 4572
rect 771 4568 772 4572
rect 757 4567 776 4568
rect 761 4563 762 4567
rect 766 4563 767 4567
rect 771 4563 772 4567
rect 757 4562 776 4563
rect 761 4558 762 4562
rect 766 4558 767 4562
rect 771 4558 772 4562
rect 757 4557 776 4558
rect 761 4553 762 4557
rect 766 4553 767 4557
rect 771 4553 772 4557
rect 757 4552 776 4553
rect 761 4548 762 4552
rect 766 4548 767 4552
rect 771 4548 772 4552
rect 787 4578 788 4582
rect 792 4578 793 4582
rect 797 4578 798 4582
rect 783 4577 802 4578
rect 787 4573 788 4577
rect 792 4573 793 4577
rect 797 4573 798 4577
rect 783 4572 802 4573
rect 787 4568 788 4572
rect 792 4568 793 4572
rect 797 4568 798 4572
rect 783 4567 802 4568
rect 787 4563 788 4567
rect 792 4563 793 4567
rect 797 4563 798 4567
rect 783 4562 802 4563
rect 787 4558 788 4562
rect 792 4558 793 4562
rect 797 4558 798 4562
rect 783 4557 802 4558
rect 787 4553 788 4557
rect 792 4553 793 4557
rect 797 4553 798 4557
rect 783 4552 802 4553
rect 787 4548 788 4552
rect 792 4548 793 4552
rect 797 4548 798 4552
rect 813 4578 814 4582
rect 818 4578 819 4582
rect 823 4578 824 4582
rect 809 4577 828 4578
rect 813 4573 814 4577
rect 818 4573 819 4577
rect 823 4573 824 4577
rect 809 4572 828 4573
rect 813 4568 814 4572
rect 818 4568 819 4572
rect 823 4568 824 4572
rect 809 4567 828 4568
rect 813 4563 814 4567
rect 818 4563 819 4567
rect 823 4563 824 4567
rect 809 4562 828 4563
rect 813 4558 814 4562
rect 818 4558 819 4562
rect 823 4558 824 4562
rect 809 4557 828 4558
rect 813 4553 814 4557
rect 818 4553 819 4557
rect 823 4553 824 4557
rect 809 4552 828 4553
rect 813 4548 814 4552
rect 818 4548 819 4552
rect 823 4548 824 4552
rect 839 4578 840 4582
rect 844 4578 845 4582
rect 849 4578 850 4582
rect 835 4577 854 4578
rect 839 4573 840 4577
rect 844 4573 845 4577
rect 849 4573 850 4577
rect 835 4572 854 4573
rect 839 4568 840 4572
rect 844 4568 845 4572
rect 849 4568 850 4572
rect 835 4567 854 4568
rect 839 4563 840 4567
rect 844 4563 845 4567
rect 849 4563 850 4567
rect 835 4562 854 4563
rect 839 4558 840 4562
rect 844 4558 845 4562
rect 849 4558 850 4562
rect 835 4557 854 4558
rect 839 4553 840 4557
rect 844 4553 845 4557
rect 849 4553 850 4557
rect 835 4552 854 4553
rect 839 4548 840 4552
rect 844 4548 845 4552
rect 849 4548 850 4552
rect 865 4578 866 4582
rect 870 4578 871 4582
rect 875 4578 876 4582
rect 861 4577 880 4578
rect 865 4573 866 4577
rect 870 4573 871 4577
rect 875 4573 876 4577
rect 861 4572 880 4573
rect 865 4568 866 4572
rect 870 4568 871 4572
rect 875 4568 876 4572
rect 861 4567 880 4568
rect 865 4563 866 4567
rect 870 4563 871 4567
rect 875 4563 876 4567
rect 861 4562 880 4563
rect 865 4558 866 4562
rect 870 4558 871 4562
rect 875 4558 876 4562
rect 861 4557 880 4558
rect 865 4553 866 4557
rect 870 4553 871 4557
rect 875 4553 876 4557
rect 861 4552 880 4553
rect 865 4548 866 4552
rect 870 4548 871 4552
rect 875 4548 876 4552
rect 1057 4578 1058 4582
rect 1062 4578 1063 4582
rect 1067 4578 1068 4582
rect 1053 4577 1072 4578
rect 1057 4573 1058 4577
rect 1062 4573 1063 4577
rect 1067 4573 1068 4577
rect 1053 4572 1072 4573
rect 1057 4568 1058 4572
rect 1062 4568 1063 4572
rect 1067 4568 1068 4572
rect 1053 4567 1072 4568
rect 1057 4563 1058 4567
rect 1062 4563 1063 4567
rect 1067 4563 1068 4567
rect 1053 4562 1072 4563
rect 1057 4558 1058 4562
rect 1062 4558 1063 4562
rect 1067 4558 1068 4562
rect 1053 4557 1072 4558
rect 1057 4553 1058 4557
rect 1062 4553 1063 4557
rect 1067 4553 1068 4557
rect 1053 4552 1072 4553
rect 1057 4548 1058 4552
rect 1062 4548 1063 4552
rect 1067 4548 1068 4552
rect 1075 4535 1131 4592
rect 1075 4531 1140 4535
rect 99 4053 1031 4528
rect 1075 4519 1131 4531
rect 1192 4527 1205 4740
rect 2675 4717 2737 4739
rect 4483 4733 4484 4737
rect 4488 4733 4489 4737
rect 4493 4733 4494 4737
rect 4498 4733 4499 4737
rect 4503 4733 4504 4737
rect 4508 4733 4509 4737
rect 4479 4732 4513 4733
rect 4483 4728 4484 4732
rect 4488 4728 4489 4732
rect 4493 4728 4494 4732
rect 4498 4728 4499 4732
rect 4503 4728 4504 4732
rect 4508 4728 4509 4732
rect 4479 4727 4513 4728
rect 4483 4723 4484 4727
rect 4488 4723 4489 4727
rect 4493 4723 4494 4727
rect 4498 4723 4499 4727
rect 4503 4723 4504 4727
rect 4508 4723 4509 4727
rect 4479 4722 4513 4723
rect 2175 4709 2441 4710
rect 1482 4685 1538 4705
rect 1366 4624 1367 4628
rect 1371 4624 1372 4628
rect 1376 4624 1377 4628
rect 1362 4623 1381 4624
rect 1366 4619 1367 4623
rect 1371 4619 1372 4623
rect 1376 4619 1377 4623
rect 1362 4618 1381 4619
rect 1366 4614 1367 4618
rect 1371 4614 1372 4618
rect 1376 4614 1377 4618
rect 1362 4613 1381 4614
rect 1366 4609 1367 4613
rect 1371 4609 1372 4613
rect 1376 4609 1377 4613
rect 1362 4608 1381 4609
rect 1366 4604 1367 4608
rect 1371 4604 1372 4608
rect 1376 4604 1377 4608
rect 1362 4603 1381 4604
rect 1366 4599 1367 4603
rect 1371 4599 1372 4603
rect 1376 4599 1377 4603
rect 1362 4598 1381 4599
rect 1366 4594 1367 4598
rect 1371 4594 1372 4598
rect 1376 4594 1377 4598
rect 1384 4601 1440 4602
rect 1384 4597 1386 4601
rect 1390 4597 1391 4601
rect 1395 4597 1396 4601
rect 1400 4597 1401 4601
rect 1405 4597 1406 4601
rect 1410 4597 1411 4601
rect 1415 4597 1416 4601
rect 1420 4597 1421 4601
rect 1425 4597 1426 4601
rect 1430 4597 1431 4601
rect 1435 4597 1436 4601
rect 1384 4596 1440 4597
rect 1384 4592 1386 4596
rect 1390 4592 1391 4596
rect 1395 4592 1396 4596
rect 1400 4592 1401 4596
rect 1405 4592 1406 4596
rect 1410 4592 1411 4596
rect 1415 4592 1416 4596
rect 1420 4592 1421 4596
rect 1425 4592 1426 4596
rect 1430 4592 1431 4596
rect 1435 4592 1436 4596
rect 1269 4578 1337 4580
rect 1269 4574 1327 4578
rect 1331 4574 1332 4578
rect 1336 4574 1337 4578
rect 1269 4573 1337 4574
rect 1269 4569 1327 4573
rect 1331 4569 1332 4573
rect 1336 4569 1337 4573
rect 1269 4568 1337 4569
rect 1269 4564 1327 4568
rect 1331 4564 1332 4568
rect 1336 4564 1337 4568
rect 1269 4563 1337 4564
rect 1269 4559 1327 4563
rect 1331 4559 1332 4563
rect 1336 4559 1337 4563
rect 1269 4558 1337 4559
rect 1269 4554 1327 4558
rect 1331 4554 1332 4558
rect 1336 4554 1337 4558
rect 1269 4553 1337 4554
rect 1269 4549 1327 4553
rect 1331 4549 1332 4553
rect 1336 4549 1337 4553
rect 1269 4548 1337 4549
rect 1366 4578 1367 4582
rect 1371 4578 1372 4582
rect 1376 4578 1377 4582
rect 1362 4577 1381 4578
rect 1366 4573 1367 4577
rect 1371 4573 1372 4577
rect 1376 4573 1377 4577
rect 1362 4572 1381 4573
rect 1366 4568 1367 4572
rect 1371 4568 1372 4572
rect 1376 4568 1377 4572
rect 1362 4567 1381 4568
rect 1366 4563 1367 4567
rect 1371 4563 1372 4567
rect 1376 4563 1377 4567
rect 1362 4562 1381 4563
rect 1366 4558 1367 4562
rect 1371 4558 1372 4562
rect 1376 4558 1377 4562
rect 1362 4557 1381 4558
rect 1366 4553 1367 4557
rect 1371 4553 1372 4557
rect 1376 4553 1377 4557
rect 1362 4552 1381 4553
rect 1366 4548 1367 4552
rect 1371 4548 1372 4552
rect 1376 4548 1377 4552
rect 1269 4544 1327 4548
rect 1331 4544 1332 4548
rect 1336 4544 1337 4548
rect 1269 4543 1337 4544
rect 1269 4539 1327 4543
rect 1331 4539 1332 4543
rect 1336 4539 1337 4543
rect 1269 4538 1337 4539
rect 1269 4535 1327 4538
rect 1266 4534 1327 4535
rect 1331 4534 1332 4538
rect 1336 4534 1337 4538
rect 1266 4533 1337 4534
rect 1266 4531 1327 4533
rect 1269 4529 1327 4531
rect 1331 4529 1332 4533
rect 1336 4529 1337 4533
rect 1269 4528 1337 4529
rect 1180 4523 1210 4527
rect 1269 4524 1327 4528
rect 1331 4524 1332 4528
rect 1336 4524 1337 4528
rect 1269 4523 1337 4524
rect 1075 4515 1140 4519
rect 1075 4503 1131 4515
rect 1183 4514 1206 4523
rect 1269 4519 1327 4523
rect 1331 4519 1332 4523
rect 1336 4519 1337 4523
rect 1266 4518 1337 4519
rect 1266 4515 1327 4518
rect 1183 4511 1187 4514
rect 1180 4507 1187 4511
rect 1199 4511 1206 4514
rect 1269 4514 1327 4515
rect 1331 4514 1332 4518
rect 1336 4514 1337 4518
rect 1269 4512 1337 4514
rect 1199 4507 1210 4511
rect 1075 4499 1140 4503
rect 1269 4503 1325 4512
rect 1075 4487 1131 4499
rect 1192 4495 1196 4502
rect 1266 4499 1325 4503
rect 1180 4491 1210 4495
rect 1269 4487 1325 4499
rect 1075 4483 1140 4487
rect 1266 4483 1325 4487
rect 1075 4475 1131 4483
rect 1078 4471 1079 4475
rect 1083 4471 1084 4475
rect 1088 4471 1089 4475
rect 1093 4471 1094 4475
rect 1098 4471 1099 4475
rect 1103 4471 1104 4475
rect 1108 4471 1109 4475
rect 1113 4471 1114 4475
rect 1118 4471 1119 4475
rect 1123 4471 1124 4475
rect 1128 4471 1129 4475
rect 1133 4471 1134 4475
rect 1138 4471 1139 4475
rect 1143 4471 1144 4475
rect 1148 4471 1149 4475
rect 1153 4471 1154 4475
rect 1158 4471 1159 4475
rect 1163 4471 1164 4475
rect 1197 4472 1206 4483
rect 1269 4475 1325 4483
rect 1384 4475 1440 4592
rect 1484 4573 1538 4685
rect 1793 4653 1845 4704
rect 1793 4649 1810 4653
rect 1814 4649 1815 4653
rect 1819 4649 1845 4653
rect 1793 4648 1845 4649
rect 1793 4644 1810 4648
rect 1814 4644 1815 4648
rect 1819 4644 1845 4648
rect 1793 4643 1845 4644
rect 1793 4639 1810 4643
rect 1814 4639 1815 4643
rect 1819 4639 1845 4643
rect 1793 4638 1845 4639
rect 1793 4634 1810 4638
rect 1814 4634 1815 4638
rect 1819 4634 1845 4638
rect 1793 4633 1845 4634
rect 1793 4629 1810 4633
rect 1814 4629 1815 4633
rect 1819 4629 1845 4633
rect 1793 4628 1845 4629
rect 2151 4705 2441 4709
rect 1675 4624 1676 4628
rect 1680 4624 1681 4628
rect 1685 4624 1686 4628
rect 1671 4623 1690 4624
rect 1675 4619 1676 4623
rect 1680 4619 1681 4623
rect 1685 4619 1686 4623
rect 1671 4618 1690 4619
rect 1675 4614 1676 4618
rect 1680 4614 1681 4618
rect 1685 4614 1686 4618
rect 1671 4613 1690 4614
rect 1675 4609 1676 4613
rect 1680 4609 1681 4613
rect 1685 4609 1686 4613
rect 1671 4608 1690 4609
rect 1675 4604 1676 4608
rect 1680 4604 1681 4608
rect 1685 4604 1686 4608
rect 1671 4603 1690 4604
rect 1675 4599 1676 4603
rect 1680 4599 1681 4603
rect 1685 4599 1686 4603
rect 1793 4624 1810 4628
rect 1814 4624 1815 4628
rect 1819 4624 1845 4628
rect 1793 4623 1845 4624
rect 1793 4619 1810 4623
rect 1814 4619 1815 4623
rect 1819 4619 1845 4623
rect 1793 4618 1845 4619
rect 1793 4614 1810 4618
rect 1814 4614 1815 4618
rect 1819 4614 1845 4618
rect 1793 4613 1845 4614
rect 1793 4609 1810 4613
rect 1814 4609 1815 4613
rect 1819 4609 1845 4613
rect 1793 4608 1845 4609
rect 1793 4604 1810 4608
rect 1814 4604 1815 4608
rect 1819 4604 1845 4608
rect 1793 4603 1845 4604
rect 1671 4598 1690 4599
rect 1675 4594 1676 4598
rect 1680 4594 1681 4598
rect 1685 4594 1686 4598
rect 1693 4601 1749 4602
rect 1693 4597 1695 4601
rect 1699 4597 1700 4601
rect 1704 4597 1705 4601
rect 1709 4597 1710 4601
rect 1714 4597 1715 4601
rect 1719 4597 1720 4601
rect 1724 4597 1725 4601
rect 1729 4597 1730 4601
rect 1734 4597 1735 4601
rect 1739 4597 1740 4601
rect 1744 4597 1745 4601
rect 1693 4596 1749 4597
rect 1693 4592 1695 4596
rect 1699 4592 1700 4596
rect 1704 4592 1705 4596
rect 1709 4592 1710 4596
rect 1714 4592 1715 4596
rect 1719 4592 1720 4596
rect 1724 4592 1725 4596
rect 1729 4592 1730 4596
rect 1734 4592 1735 4596
rect 1739 4592 1740 4596
rect 1744 4592 1745 4596
rect 1484 4569 1501 4573
rect 1505 4569 1506 4573
rect 1510 4569 1538 4573
rect 1484 4568 1538 4569
rect 1484 4564 1501 4568
rect 1505 4564 1506 4568
rect 1510 4564 1538 4568
rect 1484 4563 1538 4564
rect 1484 4559 1501 4563
rect 1505 4559 1506 4563
rect 1510 4559 1538 4563
rect 1484 4558 1538 4559
rect 1484 4554 1501 4558
rect 1505 4554 1506 4558
rect 1510 4554 1538 4558
rect 1484 4553 1538 4554
rect 1484 4549 1501 4553
rect 1505 4549 1506 4553
rect 1510 4549 1538 4553
rect 1484 4548 1538 4549
rect 1484 4544 1501 4548
rect 1505 4544 1506 4548
rect 1510 4544 1538 4548
rect 1484 4543 1538 4544
rect 1484 4539 1501 4543
rect 1505 4539 1506 4543
rect 1510 4539 1538 4543
rect 1484 4538 1538 4539
rect 1484 4534 1501 4538
rect 1505 4534 1506 4538
rect 1510 4534 1538 4538
rect 1484 4533 1538 4534
rect 1484 4529 1501 4533
rect 1505 4529 1506 4533
rect 1510 4529 1538 4533
rect 1484 4528 1538 4529
rect 1484 4524 1501 4528
rect 1505 4524 1506 4528
rect 1510 4524 1538 4528
rect 1484 4523 1538 4524
rect 1484 4519 1501 4523
rect 1505 4519 1506 4523
rect 1510 4519 1538 4523
rect 1074 4470 1078 4471
rect 1164 4470 1168 4471
rect 1195 4470 1208 4472
rect 1238 4471 1239 4475
rect 1243 4471 1244 4475
rect 1248 4471 1249 4475
rect 1253 4471 1254 4475
rect 1258 4471 1259 4475
rect 1263 4471 1264 4475
rect 1268 4471 1269 4475
rect 1273 4471 1274 4475
rect 1278 4471 1279 4475
rect 1283 4471 1284 4475
rect 1288 4471 1289 4475
rect 1293 4471 1294 4475
rect 1298 4471 1299 4475
rect 1303 4471 1304 4475
rect 1308 4471 1309 4475
rect 1313 4471 1314 4475
rect 1318 4471 1319 4475
rect 1323 4471 1324 4475
rect 1234 4470 1238 4471
rect 1193 4468 1210 4470
rect 1074 4465 1078 4466
rect 1074 4460 1078 4461
rect 1074 4455 1078 4456
rect 1074 4450 1078 4451
rect 1074 4445 1078 4446
rect 1074 4440 1078 4441
rect 1074 4435 1078 4436
rect 1074 4430 1078 4431
rect 1074 4425 1078 4426
rect 1074 4420 1078 4421
rect 1074 4415 1078 4416
rect 1074 4410 1078 4411
rect 1074 4405 1078 4406
rect 1074 4400 1078 4401
rect 1074 4395 1078 4396
rect 1074 4390 1078 4391
rect 1074 4385 1078 4386
rect 1074 4380 1078 4381
rect 1074 4375 1078 4376
rect 1074 4370 1078 4371
rect 1074 4365 1078 4366
rect 1074 4360 1078 4361
rect 1074 4355 1078 4356
rect 1074 4350 1078 4351
rect 1091 4458 1094 4466
rect 1098 4458 1099 4466
rect 1103 4458 1104 4466
rect 1108 4458 1109 4466
rect 1113 4458 1114 4466
rect 1118 4458 1119 4466
rect 1123 4458 1124 4466
rect 1128 4458 1129 4466
rect 1133 4458 1134 4466
rect 1138 4458 1139 4466
rect 1143 4458 1144 4466
rect 1148 4458 1151 4466
rect 1087 4455 1091 4458
rect 1087 4450 1091 4451
rect 1151 4455 1155 4458
rect 1151 4450 1155 4451
rect 1087 4445 1091 4446
rect 1087 4440 1091 4441
rect 1087 4435 1091 4436
rect 1087 4430 1091 4431
rect 1087 4425 1091 4426
rect 1087 4420 1091 4421
rect 1087 4415 1091 4416
rect 1087 4410 1091 4411
rect 1087 4405 1091 4406
rect 1087 4400 1091 4401
rect 1087 4395 1091 4396
rect 1087 4390 1091 4391
rect 1087 4385 1091 4386
rect 1087 4380 1091 4381
rect 1087 4375 1091 4376
rect 1087 4370 1091 4371
rect 1087 4365 1091 4366
rect 1103 4446 1104 4450
rect 1108 4446 1109 4450
rect 1113 4446 1114 4450
rect 1118 4446 1119 4450
rect 1123 4446 1124 4450
rect 1128 4446 1129 4450
rect 1133 4446 1134 4450
rect 1138 4446 1139 4450
rect 1143 4446 1144 4450
rect 1099 4445 1144 4446
rect 1103 4441 1104 4445
rect 1108 4441 1109 4445
rect 1113 4441 1114 4445
rect 1118 4441 1119 4445
rect 1123 4441 1124 4445
rect 1128 4441 1129 4445
rect 1133 4441 1134 4445
rect 1138 4441 1139 4445
rect 1143 4441 1144 4445
rect 1099 4440 1144 4441
rect 1103 4436 1104 4440
rect 1108 4436 1109 4440
rect 1113 4436 1114 4440
rect 1118 4436 1119 4440
rect 1123 4436 1124 4440
rect 1128 4436 1129 4440
rect 1133 4436 1134 4440
rect 1138 4436 1139 4440
rect 1143 4436 1144 4440
rect 1099 4435 1144 4436
rect 1103 4431 1104 4435
rect 1108 4431 1109 4435
rect 1113 4431 1114 4435
rect 1118 4431 1119 4435
rect 1123 4431 1124 4435
rect 1128 4431 1129 4435
rect 1133 4431 1134 4435
rect 1138 4431 1139 4435
rect 1143 4431 1144 4435
rect 1099 4430 1144 4431
rect 1103 4426 1104 4430
rect 1108 4426 1109 4430
rect 1113 4426 1114 4430
rect 1118 4426 1119 4430
rect 1123 4426 1124 4430
rect 1128 4426 1129 4430
rect 1133 4426 1134 4430
rect 1138 4426 1139 4430
rect 1143 4426 1144 4430
rect 1099 4425 1144 4426
rect 1103 4421 1104 4425
rect 1108 4421 1109 4425
rect 1113 4421 1114 4425
rect 1118 4421 1119 4425
rect 1123 4421 1124 4425
rect 1128 4421 1129 4425
rect 1133 4421 1134 4425
rect 1138 4421 1139 4425
rect 1143 4421 1144 4425
rect 1099 4420 1144 4421
rect 1103 4416 1104 4420
rect 1108 4416 1109 4420
rect 1113 4416 1114 4420
rect 1118 4416 1119 4420
rect 1123 4416 1124 4420
rect 1128 4416 1129 4420
rect 1133 4416 1134 4420
rect 1138 4416 1139 4420
rect 1143 4416 1144 4420
rect 1099 4415 1144 4416
rect 1103 4411 1104 4415
rect 1108 4411 1109 4415
rect 1113 4411 1114 4415
rect 1118 4411 1119 4415
rect 1123 4411 1124 4415
rect 1128 4411 1129 4415
rect 1133 4411 1134 4415
rect 1138 4411 1139 4415
rect 1143 4411 1144 4415
rect 1099 4410 1144 4411
rect 1103 4406 1104 4410
rect 1108 4406 1109 4410
rect 1113 4406 1114 4410
rect 1118 4406 1119 4410
rect 1123 4406 1124 4410
rect 1128 4406 1129 4410
rect 1133 4406 1134 4410
rect 1138 4406 1139 4410
rect 1143 4406 1144 4410
rect 1099 4405 1144 4406
rect 1103 4401 1104 4405
rect 1108 4401 1109 4405
rect 1113 4401 1114 4405
rect 1118 4401 1119 4405
rect 1123 4401 1124 4405
rect 1128 4401 1129 4405
rect 1133 4401 1134 4405
rect 1138 4401 1139 4405
rect 1143 4401 1144 4405
rect 1099 4400 1144 4401
rect 1103 4396 1104 4400
rect 1108 4396 1109 4400
rect 1113 4396 1114 4400
rect 1118 4396 1119 4400
rect 1123 4396 1124 4400
rect 1128 4396 1129 4400
rect 1133 4396 1134 4400
rect 1138 4396 1139 4400
rect 1143 4396 1144 4400
rect 1099 4395 1144 4396
rect 1103 4391 1104 4395
rect 1108 4391 1109 4395
rect 1113 4391 1114 4395
rect 1118 4391 1119 4395
rect 1123 4391 1124 4395
rect 1128 4391 1129 4395
rect 1133 4391 1134 4395
rect 1138 4391 1139 4395
rect 1143 4391 1144 4395
rect 1099 4390 1144 4391
rect 1103 4386 1104 4390
rect 1108 4386 1109 4390
rect 1113 4386 1114 4390
rect 1118 4386 1119 4390
rect 1123 4386 1124 4390
rect 1128 4386 1129 4390
rect 1133 4386 1134 4390
rect 1138 4386 1139 4390
rect 1143 4386 1144 4390
rect 1099 4385 1144 4386
rect 1103 4381 1104 4385
rect 1108 4381 1109 4385
rect 1113 4381 1114 4385
rect 1118 4381 1119 4385
rect 1123 4381 1124 4385
rect 1128 4381 1129 4385
rect 1133 4381 1134 4385
rect 1138 4381 1139 4385
rect 1143 4381 1144 4385
rect 1099 4380 1144 4381
rect 1103 4376 1104 4380
rect 1108 4376 1109 4380
rect 1113 4376 1114 4380
rect 1118 4376 1119 4380
rect 1123 4376 1124 4380
rect 1128 4376 1129 4380
rect 1133 4376 1134 4380
rect 1138 4376 1139 4380
rect 1143 4376 1144 4380
rect 1099 4375 1144 4376
rect 1103 4371 1104 4375
rect 1108 4371 1109 4375
rect 1113 4371 1114 4375
rect 1118 4371 1119 4375
rect 1123 4371 1124 4375
rect 1128 4371 1129 4375
rect 1133 4371 1134 4375
rect 1138 4371 1139 4375
rect 1143 4371 1144 4375
rect 1099 4370 1144 4371
rect 1103 4366 1104 4370
rect 1108 4366 1109 4370
rect 1113 4366 1114 4370
rect 1118 4366 1119 4370
rect 1123 4366 1124 4370
rect 1128 4366 1129 4370
rect 1133 4366 1134 4370
rect 1138 4366 1139 4370
rect 1143 4366 1144 4370
rect 1099 4365 1144 4366
rect 1103 4361 1104 4365
rect 1108 4361 1109 4365
rect 1113 4361 1114 4365
rect 1118 4361 1119 4365
rect 1123 4361 1124 4365
rect 1128 4361 1129 4365
rect 1133 4361 1134 4365
rect 1138 4361 1139 4365
rect 1143 4361 1144 4365
rect 1151 4445 1155 4446
rect 1151 4440 1155 4441
rect 1151 4435 1155 4436
rect 1151 4430 1155 4431
rect 1151 4425 1155 4426
rect 1151 4420 1155 4421
rect 1151 4415 1155 4416
rect 1151 4410 1155 4411
rect 1151 4405 1155 4406
rect 1151 4400 1155 4401
rect 1151 4395 1155 4396
rect 1151 4390 1155 4391
rect 1151 4385 1155 4386
rect 1151 4380 1155 4381
rect 1151 4375 1155 4376
rect 1151 4370 1155 4371
rect 1151 4365 1155 4366
rect 1087 4360 1091 4361
rect 1087 4353 1091 4356
rect 1151 4360 1155 4361
rect 1151 4353 1155 4356
rect 1091 4349 1094 4353
rect 1098 4349 1099 4353
rect 1103 4349 1104 4353
rect 1108 4349 1109 4353
rect 1113 4349 1114 4353
rect 1118 4349 1119 4353
rect 1123 4349 1124 4353
rect 1128 4349 1129 4353
rect 1133 4349 1134 4353
rect 1138 4349 1139 4353
rect 1143 4349 1144 4353
rect 1148 4349 1151 4353
rect 1164 4465 1168 4466
rect 1164 4460 1168 4461
rect 1164 4455 1168 4456
rect 1164 4450 1168 4451
rect 1164 4445 1168 4446
rect 1164 4440 1168 4441
rect 1164 4435 1168 4436
rect 1191 4440 1212 4468
rect 1324 4470 1328 4471
rect 1234 4465 1238 4466
rect 1234 4460 1238 4461
rect 1234 4455 1238 4456
rect 1234 4450 1238 4451
rect 1234 4445 1238 4446
rect 1234 4440 1238 4441
rect 1234 4435 1238 4436
rect 1164 4430 1168 4431
rect 1164 4425 1168 4426
rect 1164 4420 1168 4421
rect 1164 4415 1168 4416
rect 1164 4410 1168 4411
rect 1164 4405 1168 4406
rect 1164 4400 1168 4401
rect 1164 4395 1168 4396
rect 1164 4390 1168 4391
rect 1164 4385 1168 4386
rect 1164 4380 1168 4381
rect 1164 4375 1168 4376
rect 1164 4370 1168 4371
rect 1164 4365 1168 4366
rect 1234 4430 1238 4431
rect 1234 4425 1238 4426
rect 1234 4420 1238 4421
rect 1234 4415 1238 4416
rect 1234 4410 1238 4411
rect 1234 4405 1238 4406
rect 1234 4400 1238 4401
rect 1234 4395 1238 4396
rect 1234 4390 1238 4391
rect 1234 4385 1238 4386
rect 1234 4380 1238 4381
rect 1234 4375 1238 4376
rect 1234 4370 1238 4371
rect 1234 4365 1238 4366
rect 1164 4360 1168 4361
rect 1164 4355 1168 4356
rect 1164 4350 1168 4351
rect 1074 4345 1078 4346
rect 1074 4340 1078 4341
rect 1164 4345 1168 4346
rect 1164 4340 1168 4341
rect 1078 4336 1079 4340
rect 1083 4336 1084 4340
rect 1088 4336 1089 4340
rect 1093 4336 1094 4340
rect 1098 4336 1099 4340
rect 1103 4336 1104 4340
rect 1108 4336 1109 4340
rect 1113 4336 1114 4340
rect 1118 4336 1119 4340
rect 1123 4336 1124 4340
rect 1128 4336 1129 4340
rect 1133 4336 1134 4340
rect 1138 4336 1139 4340
rect 1143 4336 1144 4340
rect 1148 4336 1149 4340
rect 1153 4336 1154 4340
rect 1158 4336 1159 4340
rect 1163 4336 1164 4340
rect 1191 4333 1212 4353
rect 1234 4360 1238 4361
rect 1234 4355 1238 4356
rect 1234 4350 1238 4351
rect 1251 4458 1254 4466
rect 1258 4458 1259 4466
rect 1263 4458 1264 4466
rect 1268 4458 1269 4466
rect 1273 4458 1274 4466
rect 1278 4458 1279 4466
rect 1283 4458 1284 4466
rect 1288 4458 1289 4466
rect 1293 4458 1294 4466
rect 1298 4458 1299 4466
rect 1303 4458 1304 4466
rect 1308 4458 1311 4466
rect 1247 4455 1251 4458
rect 1247 4450 1251 4451
rect 1311 4455 1315 4458
rect 1311 4450 1315 4451
rect 1247 4445 1251 4446
rect 1247 4440 1251 4441
rect 1247 4435 1251 4436
rect 1247 4430 1251 4431
rect 1247 4425 1251 4426
rect 1247 4420 1251 4421
rect 1247 4415 1251 4416
rect 1247 4410 1251 4411
rect 1247 4405 1251 4406
rect 1247 4400 1251 4401
rect 1247 4395 1251 4396
rect 1247 4390 1251 4391
rect 1247 4385 1251 4386
rect 1247 4380 1251 4381
rect 1247 4375 1251 4376
rect 1247 4370 1251 4371
rect 1247 4365 1251 4366
rect 1263 4446 1264 4450
rect 1268 4446 1269 4450
rect 1273 4446 1274 4450
rect 1278 4446 1279 4450
rect 1283 4446 1284 4450
rect 1288 4446 1289 4450
rect 1293 4446 1294 4450
rect 1298 4446 1299 4450
rect 1259 4445 1303 4446
rect 1263 4441 1264 4445
rect 1268 4441 1269 4445
rect 1273 4441 1274 4445
rect 1278 4441 1279 4445
rect 1283 4441 1284 4445
rect 1288 4441 1289 4445
rect 1293 4441 1294 4445
rect 1298 4441 1299 4445
rect 1259 4440 1303 4441
rect 1263 4436 1264 4440
rect 1268 4436 1269 4440
rect 1273 4436 1274 4440
rect 1278 4436 1279 4440
rect 1283 4436 1284 4440
rect 1288 4436 1289 4440
rect 1293 4436 1294 4440
rect 1298 4436 1299 4440
rect 1259 4435 1303 4436
rect 1263 4431 1264 4435
rect 1268 4431 1269 4435
rect 1273 4431 1274 4435
rect 1278 4431 1279 4435
rect 1283 4431 1284 4435
rect 1288 4431 1289 4435
rect 1293 4431 1294 4435
rect 1298 4431 1299 4435
rect 1259 4430 1303 4431
rect 1263 4426 1264 4430
rect 1268 4426 1269 4430
rect 1273 4426 1274 4430
rect 1278 4426 1279 4430
rect 1283 4426 1284 4430
rect 1288 4426 1289 4430
rect 1293 4426 1294 4430
rect 1298 4426 1299 4430
rect 1259 4425 1303 4426
rect 1263 4421 1264 4425
rect 1268 4421 1269 4425
rect 1273 4421 1274 4425
rect 1278 4421 1279 4425
rect 1283 4421 1284 4425
rect 1288 4421 1289 4425
rect 1293 4421 1294 4425
rect 1298 4421 1299 4425
rect 1259 4420 1303 4421
rect 1263 4416 1264 4420
rect 1268 4416 1269 4420
rect 1273 4416 1274 4420
rect 1278 4416 1279 4420
rect 1283 4416 1284 4420
rect 1288 4416 1289 4420
rect 1293 4416 1294 4420
rect 1298 4416 1299 4420
rect 1259 4415 1303 4416
rect 1263 4411 1264 4415
rect 1268 4411 1269 4415
rect 1273 4411 1274 4415
rect 1278 4411 1279 4415
rect 1283 4411 1284 4415
rect 1288 4411 1289 4415
rect 1293 4411 1294 4415
rect 1298 4411 1299 4415
rect 1259 4410 1303 4411
rect 1263 4406 1264 4410
rect 1268 4406 1269 4410
rect 1273 4406 1274 4410
rect 1278 4406 1279 4410
rect 1283 4406 1284 4410
rect 1288 4406 1289 4410
rect 1293 4406 1294 4410
rect 1298 4406 1299 4410
rect 1259 4405 1303 4406
rect 1263 4401 1264 4405
rect 1268 4401 1269 4405
rect 1273 4401 1274 4405
rect 1278 4401 1279 4405
rect 1283 4401 1284 4405
rect 1288 4401 1289 4405
rect 1293 4401 1294 4405
rect 1298 4401 1299 4405
rect 1259 4400 1303 4401
rect 1263 4396 1264 4400
rect 1268 4396 1269 4400
rect 1273 4396 1274 4400
rect 1278 4396 1279 4400
rect 1283 4396 1284 4400
rect 1288 4396 1289 4400
rect 1293 4396 1294 4400
rect 1298 4396 1299 4400
rect 1259 4395 1303 4396
rect 1263 4391 1264 4395
rect 1268 4391 1269 4395
rect 1273 4391 1274 4395
rect 1278 4391 1279 4395
rect 1283 4391 1284 4395
rect 1288 4391 1289 4395
rect 1293 4391 1294 4395
rect 1298 4391 1299 4395
rect 1259 4390 1303 4391
rect 1263 4386 1264 4390
rect 1268 4386 1269 4390
rect 1273 4386 1274 4390
rect 1278 4386 1279 4390
rect 1283 4386 1284 4390
rect 1288 4386 1289 4390
rect 1293 4386 1294 4390
rect 1298 4386 1299 4390
rect 1259 4385 1303 4386
rect 1263 4381 1264 4385
rect 1268 4381 1269 4385
rect 1273 4381 1274 4385
rect 1278 4381 1279 4385
rect 1283 4381 1284 4385
rect 1288 4381 1289 4385
rect 1293 4381 1294 4385
rect 1298 4381 1299 4385
rect 1259 4380 1303 4381
rect 1263 4376 1264 4380
rect 1268 4376 1269 4380
rect 1273 4376 1274 4380
rect 1278 4376 1279 4380
rect 1283 4376 1284 4380
rect 1288 4376 1289 4380
rect 1293 4376 1294 4380
rect 1298 4376 1299 4380
rect 1259 4375 1303 4376
rect 1263 4371 1264 4375
rect 1268 4371 1269 4375
rect 1273 4371 1274 4375
rect 1278 4371 1279 4375
rect 1283 4371 1284 4375
rect 1288 4371 1289 4375
rect 1293 4371 1294 4375
rect 1298 4371 1299 4375
rect 1259 4370 1303 4371
rect 1263 4366 1264 4370
rect 1268 4366 1269 4370
rect 1273 4366 1274 4370
rect 1278 4366 1279 4370
rect 1283 4366 1284 4370
rect 1288 4366 1289 4370
rect 1293 4366 1294 4370
rect 1298 4366 1299 4370
rect 1259 4365 1303 4366
rect 1263 4361 1264 4365
rect 1268 4361 1269 4365
rect 1273 4361 1274 4365
rect 1278 4361 1279 4365
rect 1283 4361 1284 4365
rect 1288 4361 1289 4365
rect 1293 4361 1294 4365
rect 1298 4361 1299 4365
rect 1311 4445 1315 4446
rect 1311 4440 1315 4441
rect 1311 4435 1315 4436
rect 1311 4430 1315 4431
rect 1311 4425 1315 4426
rect 1311 4420 1315 4421
rect 1311 4415 1315 4416
rect 1311 4410 1315 4411
rect 1311 4405 1315 4406
rect 1311 4400 1315 4401
rect 1311 4395 1315 4396
rect 1311 4390 1315 4391
rect 1311 4385 1315 4386
rect 1311 4380 1315 4381
rect 1311 4375 1315 4376
rect 1311 4370 1315 4371
rect 1311 4365 1315 4366
rect 1247 4360 1251 4361
rect 1247 4353 1251 4356
rect 1311 4360 1315 4361
rect 1311 4353 1315 4356
rect 1251 4349 1254 4353
rect 1258 4349 1259 4353
rect 1263 4349 1264 4353
rect 1268 4349 1269 4353
rect 1273 4349 1274 4353
rect 1278 4349 1279 4353
rect 1283 4349 1284 4353
rect 1288 4349 1289 4353
rect 1293 4349 1294 4353
rect 1298 4349 1299 4353
rect 1303 4349 1304 4353
rect 1308 4349 1311 4353
rect 1324 4465 1328 4466
rect 1324 4460 1328 4461
rect 1324 4455 1328 4456
rect 1324 4450 1328 4451
rect 1324 4445 1328 4446
rect 1324 4440 1328 4441
rect 1324 4435 1328 4436
rect 1324 4430 1328 4431
rect 1324 4425 1328 4426
rect 1324 4420 1328 4421
rect 1324 4415 1328 4416
rect 1324 4410 1328 4411
rect 1324 4405 1328 4406
rect 1324 4400 1328 4401
rect 1324 4395 1328 4396
rect 1324 4390 1328 4391
rect 1324 4385 1328 4386
rect 1324 4380 1328 4381
rect 1324 4375 1328 4376
rect 1324 4370 1328 4371
rect 1324 4365 1328 4366
rect 1324 4360 1328 4361
rect 1324 4355 1328 4356
rect 1324 4350 1328 4351
rect 1234 4345 1238 4346
rect 1234 4340 1238 4341
rect 1324 4345 1328 4346
rect 1324 4340 1328 4341
rect 1238 4336 1239 4340
rect 1243 4336 1244 4340
rect 1248 4336 1249 4340
rect 1253 4336 1254 4340
rect 1258 4336 1259 4340
rect 1263 4336 1264 4340
rect 1268 4336 1269 4340
rect 1273 4336 1274 4340
rect 1278 4336 1279 4340
rect 1283 4336 1284 4340
rect 1288 4336 1289 4340
rect 1293 4336 1294 4340
rect 1298 4336 1299 4340
rect 1303 4336 1304 4340
rect 1308 4336 1309 4340
rect 1313 4336 1314 4340
rect 1318 4336 1319 4340
rect 1323 4336 1324 4340
rect 1387 4471 1388 4475
rect 1392 4471 1393 4475
rect 1397 4471 1398 4475
rect 1402 4471 1403 4475
rect 1407 4471 1408 4475
rect 1412 4471 1413 4475
rect 1417 4471 1418 4475
rect 1422 4471 1423 4475
rect 1427 4471 1428 4475
rect 1432 4471 1433 4475
rect 1437 4471 1438 4475
rect 1442 4471 1443 4475
rect 1447 4471 1448 4475
rect 1452 4471 1453 4475
rect 1457 4471 1458 4475
rect 1462 4471 1463 4475
rect 1467 4471 1468 4475
rect 1472 4471 1473 4475
rect 1383 4470 1387 4471
rect 1473 4470 1477 4471
rect 1383 4465 1387 4466
rect 1383 4460 1387 4461
rect 1383 4455 1387 4456
rect 1383 4450 1387 4451
rect 1383 4445 1387 4446
rect 1383 4440 1387 4441
rect 1383 4435 1387 4436
rect 1383 4430 1387 4431
rect 1383 4425 1387 4426
rect 1383 4420 1387 4421
rect 1383 4415 1387 4416
rect 1383 4410 1387 4411
rect 1383 4405 1387 4406
rect 1383 4400 1387 4401
rect 1383 4395 1387 4396
rect 1383 4390 1387 4391
rect 1383 4385 1387 4386
rect 1383 4380 1387 4381
rect 1383 4375 1387 4376
rect 1383 4370 1387 4371
rect 1383 4365 1387 4366
rect 1383 4360 1387 4361
rect 1383 4355 1387 4356
rect 1383 4350 1387 4351
rect 1400 4458 1403 4466
rect 1407 4458 1408 4466
rect 1412 4458 1413 4466
rect 1417 4458 1418 4466
rect 1422 4458 1423 4466
rect 1427 4458 1428 4466
rect 1432 4458 1433 4466
rect 1437 4458 1438 4466
rect 1442 4458 1443 4466
rect 1447 4458 1448 4466
rect 1452 4458 1453 4466
rect 1457 4458 1460 4466
rect 1396 4455 1400 4458
rect 1396 4450 1400 4451
rect 1460 4455 1464 4458
rect 1460 4450 1464 4451
rect 1396 4445 1400 4446
rect 1396 4440 1400 4441
rect 1396 4435 1400 4436
rect 1396 4430 1400 4431
rect 1396 4425 1400 4426
rect 1396 4420 1400 4421
rect 1396 4415 1400 4416
rect 1396 4410 1400 4411
rect 1396 4405 1400 4406
rect 1396 4400 1400 4401
rect 1396 4395 1400 4396
rect 1396 4390 1400 4391
rect 1396 4385 1400 4386
rect 1396 4380 1400 4381
rect 1396 4375 1400 4376
rect 1396 4370 1400 4371
rect 1396 4365 1400 4366
rect 1412 4446 1413 4450
rect 1417 4446 1418 4450
rect 1422 4446 1423 4450
rect 1427 4446 1428 4450
rect 1432 4446 1433 4450
rect 1437 4446 1438 4450
rect 1442 4446 1443 4450
rect 1447 4446 1448 4450
rect 1452 4446 1453 4450
rect 1408 4445 1453 4446
rect 1412 4441 1413 4445
rect 1417 4441 1418 4445
rect 1422 4441 1423 4445
rect 1427 4441 1428 4445
rect 1432 4441 1433 4445
rect 1437 4441 1438 4445
rect 1442 4441 1443 4445
rect 1447 4441 1448 4445
rect 1452 4441 1453 4445
rect 1408 4440 1453 4441
rect 1412 4436 1413 4440
rect 1417 4436 1418 4440
rect 1422 4436 1423 4440
rect 1427 4436 1428 4440
rect 1432 4436 1433 4440
rect 1437 4436 1438 4440
rect 1442 4436 1443 4440
rect 1447 4436 1448 4440
rect 1452 4436 1453 4440
rect 1408 4435 1453 4436
rect 1412 4431 1413 4435
rect 1417 4431 1418 4435
rect 1422 4431 1423 4435
rect 1427 4431 1428 4435
rect 1432 4431 1433 4435
rect 1437 4431 1438 4435
rect 1442 4431 1443 4435
rect 1447 4431 1448 4435
rect 1452 4431 1453 4435
rect 1408 4430 1453 4431
rect 1412 4426 1413 4430
rect 1417 4426 1418 4430
rect 1422 4426 1423 4430
rect 1427 4426 1428 4430
rect 1432 4426 1433 4430
rect 1437 4426 1438 4430
rect 1442 4426 1443 4430
rect 1447 4426 1448 4430
rect 1452 4426 1453 4430
rect 1408 4425 1453 4426
rect 1412 4421 1413 4425
rect 1417 4421 1418 4425
rect 1422 4421 1423 4425
rect 1427 4421 1428 4425
rect 1432 4421 1433 4425
rect 1437 4421 1438 4425
rect 1442 4421 1443 4425
rect 1447 4421 1448 4425
rect 1452 4421 1453 4425
rect 1408 4420 1453 4421
rect 1412 4416 1413 4420
rect 1417 4416 1418 4420
rect 1422 4416 1423 4420
rect 1427 4416 1428 4420
rect 1432 4416 1433 4420
rect 1437 4416 1438 4420
rect 1442 4416 1443 4420
rect 1447 4416 1448 4420
rect 1452 4416 1453 4420
rect 1408 4415 1453 4416
rect 1412 4411 1413 4415
rect 1417 4411 1418 4415
rect 1422 4411 1423 4415
rect 1427 4411 1428 4415
rect 1432 4411 1433 4415
rect 1437 4411 1438 4415
rect 1442 4411 1443 4415
rect 1447 4411 1448 4415
rect 1452 4411 1453 4415
rect 1408 4410 1453 4411
rect 1412 4406 1413 4410
rect 1417 4406 1418 4410
rect 1422 4406 1423 4410
rect 1427 4406 1428 4410
rect 1432 4406 1433 4410
rect 1437 4406 1438 4410
rect 1442 4406 1443 4410
rect 1447 4406 1448 4410
rect 1452 4406 1453 4410
rect 1408 4405 1453 4406
rect 1412 4401 1413 4405
rect 1417 4401 1418 4405
rect 1422 4401 1423 4405
rect 1427 4401 1428 4405
rect 1432 4401 1433 4405
rect 1437 4401 1438 4405
rect 1442 4401 1443 4405
rect 1447 4401 1448 4405
rect 1452 4401 1453 4405
rect 1408 4400 1453 4401
rect 1412 4396 1413 4400
rect 1417 4396 1418 4400
rect 1422 4396 1423 4400
rect 1427 4396 1428 4400
rect 1432 4396 1433 4400
rect 1437 4396 1438 4400
rect 1442 4396 1443 4400
rect 1447 4396 1448 4400
rect 1452 4396 1453 4400
rect 1408 4395 1453 4396
rect 1412 4391 1413 4395
rect 1417 4391 1418 4395
rect 1422 4391 1423 4395
rect 1427 4391 1428 4395
rect 1432 4391 1433 4395
rect 1437 4391 1438 4395
rect 1442 4391 1443 4395
rect 1447 4391 1448 4395
rect 1452 4391 1453 4395
rect 1408 4390 1453 4391
rect 1412 4386 1413 4390
rect 1417 4386 1418 4390
rect 1422 4386 1423 4390
rect 1427 4386 1428 4390
rect 1432 4386 1433 4390
rect 1437 4386 1438 4390
rect 1442 4386 1443 4390
rect 1447 4386 1448 4390
rect 1452 4386 1453 4390
rect 1408 4385 1453 4386
rect 1412 4381 1413 4385
rect 1417 4381 1418 4385
rect 1422 4381 1423 4385
rect 1427 4381 1428 4385
rect 1432 4381 1433 4385
rect 1437 4381 1438 4385
rect 1442 4381 1443 4385
rect 1447 4381 1448 4385
rect 1452 4381 1453 4385
rect 1408 4380 1453 4381
rect 1412 4376 1413 4380
rect 1417 4376 1418 4380
rect 1422 4376 1423 4380
rect 1427 4376 1428 4380
rect 1432 4376 1433 4380
rect 1437 4376 1438 4380
rect 1442 4376 1443 4380
rect 1447 4376 1448 4380
rect 1452 4376 1453 4380
rect 1408 4375 1453 4376
rect 1412 4371 1413 4375
rect 1417 4371 1418 4375
rect 1422 4371 1423 4375
rect 1427 4371 1428 4375
rect 1432 4371 1433 4375
rect 1437 4371 1438 4375
rect 1442 4371 1443 4375
rect 1447 4371 1448 4375
rect 1452 4371 1453 4375
rect 1408 4370 1453 4371
rect 1412 4366 1413 4370
rect 1417 4366 1418 4370
rect 1422 4366 1423 4370
rect 1427 4366 1428 4370
rect 1432 4366 1433 4370
rect 1437 4366 1438 4370
rect 1442 4366 1443 4370
rect 1447 4366 1448 4370
rect 1452 4366 1453 4370
rect 1408 4365 1453 4366
rect 1412 4361 1413 4365
rect 1417 4361 1418 4365
rect 1422 4361 1423 4365
rect 1427 4361 1428 4365
rect 1432 4361 1433 4365
rect 1437 4361 1438 4365
rect 1442 4361 1443 4365
rect 1447 4361 1448 4365
rect 1452 4361 1453 4365
rect 1460 4445 1464 4446
rect 1460 4440 1464 4441
rect 1460 4435 1464 4436
rect 1460 4430 1464 4431
rect 1460 4425 1464 4426
rect 1460 4420 1464 4421
rect 1460 4415 1464 4416
rect 1460 4410 1464 4411
rect 1460 4405 1464 4406
rect 1460 4400 1464 4401
rect 1460 4395 1464 4396
rect 1460 4390 1464 4391
rect 1460 4385 1464 4386
rect 1460 4380 1464 4381
rect 1460 4375 1464 4376
rect 1460 4370 1464 4371
rect 1460 4365 1464 4366
rect 1396 4360 1400 4361
rect 1396 4353 1400 4356
rect 1460 4360 1464 4361
rect 1460 4353 1464 4356
rect 1400 4349 1403 4353
rect 1407 4349 1408 4353
rect 1412 4349 1413 4353
rect 1417 4349 1418 4353
rect 1422 4349 1423 4353
rect 1427 4349 1428 4353
rect 1432 4349 1433 4353
rect 1437 4349 1438 4353
rect 1442 4349 1443 4353
rect 1447 4349 1448 4353
rect 1452 4349 1453 4353
rect 1457 4349 1460 4353
rect 1473 4465 1477 4466
rect 1473 4460 1477 4461
rect 1473 4455 1477 4456
rect 1473 4450 1477 4451
rect 1473 4445 1477 4446
rect 1473 4440 1477 4441
rect 1473 4435 1477 4436
rect 1473 4430 1477 4431
rect 1473 4425 1477 4426
rect 1473 4420 1477 4421
rect 1473 4415 1477 4416
rect 1473 4410 1477 4411
rect 1473 4405 1477 4406
rect 1473 4400 1477 4401
rect 1473 4395 1477 4396
rect 1473 4390 1477 4391
rect 1473 4385 1477 4386
rect 1473 4380 1477 4381
rect 1473 4375 1477 4376
rect 1473 4370 1477 4371
rect 1473 4365 1477 4366
rect 1473 4360 1477 4361
rect 1473 4355 1477 4356
rect 1473 4350 1477 4351
rect 1383 4345 1387 4346
rect 1383 4340 1387 4341
rect 1473 4345 1477 4346
rect 1473 4340 1477 4341
rect 1387 4336 1388 4340
rect 1392 4336 1393 4340
rect 1397 4336 1398 4340
rect 1402 4336 1403 4340
rect 1407 4336 1408 4340
rect 1412 4336 1413 4340
rect 1417 4336 1418 4340
rect 1422 4336 1423 4340
rect 1427 4336 1428 4340
rect 1432 4336 1433 4340
rect 1437 4336 1438 4340
rect 1442 4336 1443 4340
rect 1447 4336 1448 4340
rect 1452 4336 1453 4340
rect 1457 4336 1458 4340
rect 1462 4336 1463 4340
rect 1467 4336 1468 4340
rect 1472 4336 1473 4340
rect 1484 4333 1538 4519
rect 1578 4578 1646 4580
rect 1578 4574 1636 4578
rect 1640 4574 1641 4578
rect 1645 4574 1646 4578
rect 1578 4573 1646 4574
rect 1578 4569 1636 4573
rect 1640 4569 1641 4573
rect 1645 4569 1646 4573
rect 1578 4568 1646 4569
rect 1578 4564 1636 4568
rect 1640 4564 1641 4568
rect 1645 4564 1646 4568
rect 1578 4563 1646 4564
rect 1578 4559 1636 4563
rect 1640 4559 1641 4563
rect 1645 4559 1646 4563
rect 1578 4558 1646 4559
rect 1578 4554 1636 4558
rect 1640 4554 1641 4558
rect 1645 4554 1646 4558
rect 1578 4553 1646 4554
rect 1578 4549 1636 4553
rect 1640 4549 1641 4553
rect 1645 4549 1646 4553
rect 1578 4548 1646 4549
rect 1675 4578 1676 4582
rect 1680 4578 1681 4582
rect 1685 4578 1686 4582
rect 1671 4577 1690 4578
rect 1675 4573 1676 4577
rect 1680 4573 1681 4577
rect 1685 4573 1686 4577
rect 1671 4572 1690 4573
rect 1675 4568 1676 4572
rect 1680 4568 1681 4572
rect 1685 4568 1686 4572
rect 1671 4567 1690 4568
rect 1675 4563 1676 4567
rect 1680 4563 1681 4567
rect 1685 4563 1686 4567
rect 1671 4562 1690 4563
rect 1675 4558 1676 4562
rect 1680 4558 1681 4562
rect 1685 4558 1686 4562
rect 1671 4557 1690 4558
rect 1675 4553 1676 4557
rect 1680 4553 1681 4557
rect 1685 4553 1686 4557
rect 1671 4552 1690 4553
rect 1675 4548 1676 4552
rect 1680 4548 1681 4552
rect 1685 4548 1686 4552
rect 1578 4544 1636 4548
rect 1640 4544 1641 4548
rect 1645 4544 1646 4548
rect 1578 4543 1646 4544
rect 1578 4539 1636 4543
rect 1640 4539 1641 4543
rect 1645 4539 1646 4543
rect 1578 4538 1646 4539
rect 1578 4534 1636 4538
rect 1640 4534 1641 4538
rect 1645 4534 1646 4538
rect 1578 4533 1646 4534
rect 1578 4529 1636 4533
rect 1640 4529 1641 4533
rect 1645 4529 1646 4533
rect 1578 4528 1646 4529
rect 1578 4524 1636 4528
rect 1640 4524 1641 4528
rect 1645 4524 1646 4528
rect 1578 4523 1646 4524
rect 1578 4519 1636 4523
rect 1640 4519 1641 4523
rect 1645 4519 1646 4523
rect 1578 4518 1646 4519
rect 1578 4514 1636 4518
rect 1640 4514 1641 4518
rect 1645 4514 1646 4518
rect 1578 4512 1646 4514
rect 1578 4475 1634 4512
rect 1693 4475 1749 4592
rect 1793 4599 1810 4603
rect 1814 4599 1815 4603
rect 1819 4599 1845 4603
rect 1547 4471 1548 4475
rect 1552 4471 1553 4475
rect 1557 4471 1558 4475
rect 1562 4471 1563 4475
rect 1567 4471 1568 4475
rect 1572 4471 1573 4475
rect 1577 4471 1578 4475
rect 1582 4471 1583 4475
rect 1587 4471 1588 4475
rect 1592 4471 1593 4475
rect 1597 4471 1598 4475
rect 1602 4471 1603 4475
rect 1607 4471 1608 4475
rect 1612 4471 1613 4475
rect 1617 4471 1618 4475
rect 1622 4471 1623 4475
rect 1627 4471 1628 4475
rect 1632 4471 1633 4475
rect 1543 4470 1547 4471
rect 1633 4470 1637 4471
rect 1543 4465 1547 4466
rect 1543 4460 1547 4461
rect 1543 4455 1547 4456
rect 1543 4450 1547 4451
rect 1543 4445 1547 4446
rect 1543 4440 1547 4441
rect 1543 4435 1547 4436
rect 1543 4430 1547 4431
rect 1543 4425 1547 4426
rect 1543 4420 1547 4421
rect 1543 4415 1547 4416
rect 1543 4410 1547 4411
rect 1543 4405 1547 4406
rect 1543 4400 1547 4401
rect 1543 4395 1547 4396
rect 1543 4390 1547 4391
rect 1543 4385 1547 4386
rect 1543 4380 1547 4381
rect 1543 4375 1547 4376
rect 1543 4370 1547 4371
rect 1543 4365 1547 4366
rect 1543 4360 1547 4361
rect 1543 4355 1547 4356
rect 1543 4350 1547 4351
rect 1560 4458 1563 4466
rect 1567 4458 1568 4466
rect 1572 4458 1573 4466
rect 1577 4458 1578 4466
rect 1582 4458 1583 4466
rect 1587 4458 1588 4466
rect 1592 4458 1593 4466
rect 1597 4458 1598 4466
rect 1602 4458 1603 4466
rect 1607 4458 1608 4466
rect 1612 4458 1613 4466
rect 1617 4458 1620 4466
rect 1556 4455 1560 4458
rect 1556 4450 1560 4451
rect 1620 4455 1624 4458
rect 1620 4450 1624 4451
rect 1556 4445 1560 4446
rect 1556 4440 1560 4441
rect 1556 4435 1560 4436
rect 1556 4430 1560 4431
rect 1556 4425 1560 4426
rect 1556 4420 1560 4421
rect 1556 4415 1560 4416
rect 1556 4410 1560 4411
rect 1556 4405 1560 4406
rect 1556 4400 1560 4401
rect 1556 4395 1560 4396
rect 1556 4390 1560 4391
rect 1556 4385 1560 4386
rect 1556 4380 1560 4381
rect 1556 4375 1560 4376
rect 1556 4370 1560 4371
rect 1556 4365 1560 4366
rect 1572 4446 1573 4450
rect 1577 4446 1578 4450
rect 1582 4446 1583 4450
rect 1587 4446 1588 4450
rect 1592 4446 1593 4450
rect 1597 4446 1598 4450
rect 1602 4446 1603 4450
rect 1607 4446 1608 4450
rect 1568 4445 1612 4446
rect 1572 4441 1573 4445
rect 1577 4441 1578 4445
rect 1582 4441 1583 4445
rect 1587 4441 1588 4445
rect 1592 4441 1593 4445
rect 1597 4441 1598 4445
rect 1602 4441 1603 4445
rect 1607 4441 1608 4445
rect 1568 4440 1612 4441
rect 1572 4436 1573 4440
rect 1577 4436 1578 4440
rect 1582 4436 1583 4440
rect 1587 4436 1588 4440
rect 1592 4436 1593 4440
rect 1597 4436 1598 4440
rect 1602 4436 1603 4440
rect 1607 4436 1608 4440
rect 1568 4435 1612 4436
rect 1572 4431 1573 4435
rect 1577 4431 1578 4435
rect 1582 4431 1583 4435
rect 1587 4431 1588 4435
rect 1592 4431 1593 4435
rect 1597 4431 1598 4435
rect 1602 4431 1603 4435
rect 1607 4431 1608 4435
rect 1568 4430 1612 4431
rect 1572 4426 1573 4430
rect 1577 4426 1578 4430
rect 1582 4426 1583 4430
rect 1587 4426 1588 4430
rect 1592 4426 1593 4430
rect 1597 4426 1598 4430
rect 1602 4426 1603 4430
rect 1607 4426 1608 4430
rect 1568 4425 1612 4426
rect 1572 4421 1573 4425
rect 1577 4421 1578 4425
rect 1582 4421 1583 4425
rect 1587 4421 1588 4425
rect 1592 4421 1593 4425
rect 1597 4421 1598 4425
rect 1602 4421 1603 4425
rect 1607 4421 1608 4425
rect 1568 4420 1612 4421
rect 1572 4416 1573 4420
rect 1577 4416 1578 4420
rect 1582 4416 1583 4420
rect 1587 4416 1588 4420
rect 1592 4416 1593 4420
rect 1597 4416 1598 4420
rect 1602 4416 1603 4420
rect 1607 4416 1608 4420
rect 1568 4415 1612 4416
rect 1572 4411 1573 4415
rect 1577 4411 1578 4415
rect 1582 4411 1583 4415
rect 1587 4411 1588 4415
rect 1592 4411 1593 4415
rect 1597 4411 1598 4415
rect 1602 4411 1603 4415
rect 1607 4411 1608 4415
rect 1568 4410 1612 4411
rect 1572 4406 1573 4410
rect 1577 4406 1578 4410
rect 1582 4406 1583 4410
rect 1587 4406 1588 4410
rect 1592 4406 1593 4410
rect 1597 4406 1598 4410
rect 1602 4406 1603 4410
rect 1607 4406 1608 4410
rect 1568 4405 1612 4406
rect 1572 4401 1573 4405
rect 1577 4401 1578 4405
rect 1582 4401 1583 4405
rect 1587 4401 1588 4405
rect 1592 4401 1593 4405
rect 1597 4401 1598 4405
rect 1602 4401 1603 4405
rect 1607 4401 1608 4405
rect 1568 4400 1612 4401
rect 1572 4396 1573 4400
rect 1577 4396 1578 4400
rect 1582 4396 1583 4400
rect 1587 4396 1588 4400
rect 1592 4396 1593 4400
rect 1597 4396 1598 4400
rect 1602 4396 1603 4400
rect 1607 4396 1608 4400
rect 1568 4395 1612 4396
rect 1572 4391 1573 4395
rect 1577 4391 1578 4395
rect 1582 4391 1583 4395
rect 1587 4391 1588 4395
rect 1592 4391 1593 4395
rect 1597 4391 1598 4395
rect 1602 4391 1603 4395
rect 1607 4391 1608 4395
rect 1568 4390 1612 4391
rect 1572 4386 1573 4390
rect 1577 4386 1578 4390
rect 1582 4386 1583 4390
rect 1587 4386 1588 4390
rect 1592 4386 1593 4390
rect 1597 4386 1598 4390
rect 1602 4386 1603 4390
rect 1607 4386 1608 4390
rect 1568 4385 1612 4386
rect 1572 4381 1573 4385
rect 1577 4381 1578 4385
rect 1582 4381 1583 4385
rect 1587 4381 1588 4385
rect 1592 4381 1593 4385
rect 1597 4381 1598 4385
rect 1602 4381 1603 4385
rect 1607 4381 1608 4385
rect 1568 4380 1612 4381
rect 1572 4376 1573 4380
rect 1577 4376 1578 4380
rect 1582 4376 1583 4380
rect 1587 4376 1588 4380
rect 1592 4376 1593 4380
rect 1597 4376 1598 4380
rect 1602 4376 1603 4380
rect 1607 4376 1608 4380
rect 1568 4375 1612 4376
rect 1572 4371 1573 4375
rect 1577 4371 1578 4375
rect 1582 4371 1583 4375
rect 1587 4371 1588 4375
rect 1592 4371 1593 4375
rect 1597 4371 1598 4375
rect 1602 4371 1603 4375
rect 1607 4371 1608 4375
rect 1568 4370 1612 4371
rect 1572 4366 1573 4370
rect 1577 4366 1578 4370
rect 1582 4366 1583 4370
rect 1587 4366 1588 4370
rect 1592 4366 1593 4370
rect 1597 4366 1598 4370
rect 1602 4366 1603 4370
rect 1607 4366 1608 4370
rect 1568 4365 1612 4366
rect 1572 4361 1573 4365
rect 1577 4361 1578 4365
rect 1582 4361 1583 4365
rect 1587 4361 1588 4365
rect 1592 4361 1593 4365
rect 1597 4361 1598 4365
rect 1602 4361 1603 4365
rect 1607 4361 1608 4365
rect 1620 4445 1624 4446
rect 1620 4440 1624 4441
rect 1620 4435 1624 4436
rect 1620 4430 1624 4431
rect 1620 4425 1624 4426
rect 1620 4420 1624 4421
rect 1620 4415 1624 4416
rect 1620 4410 1624 4411
rect 1620 4405 1624 4406
rect 1620 4400 1624 4401
rect 1620 4395 1624 4396
rect 1620 4390 1624 4391
rect 1620 4385 1624 4386
rect 1620 4380 1624 4381
rect 1620 4375 1624 4376
rect 1620 4370 1624 4371
rect 1620 4365 1624 4366
rect 1556 4360 1560 4361
rect 1556 4353 1560 4356
rect 1620 4360 1624 4361
rect 1620 4353 1624 4356
rect 1560 4349 1563 4353
rect 1567 4349 1568 4353
rect 1572 4349 1573 4353
rect 1577 4349 1578 4353
rect 1582 4349 1583 4353
rect 1587 4349 1588 4353
rect 1592 4349 1593 4353
rect 1597 4349 1598 4353
rect 1602 4349 1603 4353
rect 1607 4349 1608 4353
rect 1612 4349 1613 4353
rect 1617 4349 1620 4353
rect 1633 4465 1637 4466
rect 1633 4460 1637 4461
rect 1633 4455 1637 4456
rect 1633 4450 1637 4451
rect 1633 4445 1637 4446
rect 1633 4440 1637 4441
rect 1633 4435 1637 4436
rect 1633 4430 1637 4431
rect 1633 4425 1637 4426
rect 1633 4420 1637 4421
rect 1633 4415 1637 4416
rect 1633 4410 1637 4411
rect 1633 4405 1637 4406
rect 1633 4400 1637 4401
rect 1633 4395 1637 4396
rect 1633 4390 1637 4391
rect 1633 4385 1637 4386
rect 1633 4380 1637 4381
rect 1633 4375 1637 4376
rect 1633 4370 1637 4371
rect 1633 4365 1637 4366
rect 1633 4360 1637 4361
rect 1633 4355 1637 4356
rect 1633 4350 1637 4351
rect 1543 4345 1547 4346
rect 1543 4340 1547 4341
rect 1633 4345 1637 4346
rect 1633 4340 1637 4341
rect 1547 4336 1548 4340
rect 1552 4336 1553 4340
rect 1557 4336 1558 4340
rect 1562 4336 1563 4340
rect 1567 4336 1568 4340
rect 1572 4336 1573 4340
rect 1577 4336 1578 4340
rect 1582 4336 1583 4340
rect 1587 4336 1588 4340
rect 1592 4336 1593 4340
rect 1597 4336 1598 4340
rect 1602 4336 1603 4340
rect 1607 4336 1608 4340
rect 1612 4336 1613 4340
rect 1617 4336 1618 4340
rect 1622 4336 1623 4340
rect 1627 4336 1628 4340
rect 1632 4336 1633 4340
rect 1696 4471 1697 4475
rect 1701 4471 1702 4475
rect 1706 4471 1707 4475
rect 1711 4471 1712 4475
rect 1716 4471 1717 4475
rect 1721 4471 1722 4475
rect 1726 4471 1727 4475
rect 1731 4471 1732 4475
rect 1736 4471 1737 4475
rect 1741 4471 1742 4475
rect 1746 4471 1747 4475
rect 1751 4471 1752 4475
rect 1756 4471 1757 4475
rect 1761 4471 1762 4475
rect 1766 4471 1767 4475
rect 1771 4471 1772 4475
rect 1776 4471 1777 4475
rect 1781 4471 1782 4475
rect 1692 4470 1696 4471
rect 1782 4470 1786 4471
rect 1692 4465 1696 4466
rect 1692 4460 1696 4461
rect 1692 4455 1696 4456
rect 1692 4450 1696 4451
rect 1692 4445 1696 4446
rect 1692 4440 1696 4441
rect 1692 4435 1696 4436
rect 1692 4430 1696 4431
rect 1692 4425 1696 4426
rect 1692 4420 1696 4421
rect 1692 4415 1696 4416
rect 1692 4410 1696 4411
rect 1692 4405 1696 4406
rect 1692 4400 1696 4401
rect 1692 4395 1696 4396
rect 1692 4390 1696 4391
rect 1692 4385 1696 4386
rect 1692 4380 1696 4381
rect 1692 4375 1696 4376
rect 1692 4370 1696 4371
rect 1692 4365 1696 4366
rect 1692 4360 1696 4361
rect 1692 4355 1696 4356
rect 1692 4350 1696 4351
rect 1709 4458 1712 4466
rect 1716 4458 1717 4466
rect 1721 4458 1722 4466
rect 1726 4458 1727 4466
rect 1731 4458 1732 4466
rect 1736 4458 1737 4466
rect 1741 4458 1742 4466
rect 1746 4458 1747 4466
rect 1751 4458 1752 4466
rect 1756 4458 1757 4466
rect 1761 4458 1762 4466
rect 1766 4458 1769 4466
rect 1705 4455 1709 4458
rect 1705 4450 1709 4451
rect 1769 4455 1773 4458
rect 1769 4450 1773 4451
rect 1705 4445 1709 4446
rect 1705 4440 1709 4441
rect 1705 4435 1709 4436
rect 1705 4430 1709 4431
rect 1705 4425 1709 4426
rect 1705 4420 1709 4421
rect 1705 4415 1709 4416
rect 1705 4410 1709 4411
rect 1705 4405 1709 4406
rect 1705 4400 1709 4401
rect 1705 4395 1709 4396
rect 1705 4390 1709 4391
rect 1705 4385 1709 4386
rect 1705 4380 1709 4381
rect 1705 4375 1709 4376
rect 1705 4370 1709 4371
rect 1705 4365 1709 4366
rect 1721 4446 1722 4450
rect 1726 4446 1727 4450
rect 1731 4446 1732 4450
rect 1736 4446 1737 4450
rect 1741 4446 1742 4450
rect 1746 4446 1747 4450
rect 1751 4446 1752 4450
rect 1756 4446 1757 4450
rect 1761 4446 1762 4450
rect 1717 4445 1762 4446
rect 1721 4441 1722 4445
rect 1726 4441 1727 4445
rect 1731 4441 1732 4445
rect 1736 4441 1737 4445
rect 1741 4441 1742 4445
rect 1746 4441 1747 4445
rect 1751 4441 1752 4445
rect 1756 4441 1757 4445
rect 1761 4441 1762 4445
rect 1717 4440 1762 4441
rect 1721 4436 1722 4440
rect 1726 4436 1727 4440
rect 1731 4436 1732 4440
rect 1736 4436 1737 4440
rect 1741 4436 1742 4440
rect 1746 4436 1747 4440
rect 1751 4436 1752 4440
rect 1756 4436 1757 4440
rect 1761 4436 1762 4440
rect 1717 4435 1762 4436
rect 1721 4431 1722 4435
rect 1726 4431 1727 4435
rect 1731 4431 1732 4435
rect 1736 4431 1737 4435
rect 1741 4431 1742 4435
rect 1746 4431 1747 4435
rect 1751 4431 1752 4435
rect 1756 4431 1757 4435
rect 1761 4431 1762 4435
rect 1717 4430 1762 4431
rect 1721 4426 1722 4430
rect 1726 4426 1727 4430
rect 1731 4426 1732 4430
rect 1736 4426 1737 4430
rect 1741 4426 1742 4430
rect 1746 4426 1747 4430
rect 1751 4426 1752 4430
rect 1756 4426 1757 4430
rect 1761 4426 1762 4430
rect 1717 4425 1762 4426
rect 1721 4421 1722 4425
rect 1726 4421 1727 4425
rect 1731 4421 1732 4425
rect 1736 4421 1737 4425
rect 1741 4421 1742 4425
rect 1746 4421 1747 4425
rect 1751 4421 1752 4425
rect 1756 4421 1757 4425
rect 1761 4421 1762 4425
rect 1717 4420 1762 4421
rect 1721 4416 1722 4420
rect 1726 4416 1727 4420
rect 1731 4416 1732 4420
rect 1736 4416 1737 4420
rect 1741 4416 1742 4420
rect 1746 4416 1747 4420
rect 1751 4416 1752 4420
rect 1756 4416 1757 4420
rect 1761 4416 1762 4420
rect 1717 4415 1762 4416
rect 1721 4411 1722 4415
rect 1726 4411 1727 4415
rect 1731 4411 1732 4415
rect 1736 4411 1737 4415
rect 1741 4411 1742 4415
rect 1746 4411 1747 4415
rect 1751 4411 1752 4415
rect 1756 4411 1757 4415
rect 1761 4411 1762 4415
rect 1717 4410 1762 4411
rect 1721 4406 1722 4410
rect 1726 4406 1727 4410
rect 1731 4406 1732 4410
rect 1736 4406 1737 4410
rect 1741 4406 1742 4410
rect 1746 4406 1747 4410
rect 1751 4406 1752 4410
rect 1756 4406 1757 4410
rect 1761 4406 1762 4410
rect 1717 4405 1762 4406
rect 1721 4401 1722 4405
rect 1726 4401 1727 4405
rect 1731 4401 1732 4405
rect 1736 4401 1737 4405
rect 1741 4401 1742 4405
rect 1746 4401 1747 4405
rect 1751 4401 1752 4405
rect 1756 4401 1757 4405
rect 1761 4401 1762 4405
rect 1717 4400 1762 4401
rect 1721 4396 1722 4400
rect 1726 4396 1727 4400
rect 1731 4396 1732 4400
rect 1736 4396 1737 4400
rect 1741 4396 1742 4400
rect 1746 4396 1747 4400
rect 1751 4396 1752 4400
rect 1756 4396 1757 4400
rect 1761 4396 1762 4400
rect 1717 4395 1762 4396
rect 1721 4391 1722 4395
rect 1726 4391 1727 4395
rect 1731 4391 1732 4395
rect 1736 4391 1737 4395
rect 1741 4391 1742 4395
rect 1746 4391 1747 4395
rect 1751 4391 1752 4395
rect 1756 4391 1757 4395
rect 1761 4391 1762 4395
rect 1717 4390 1762 4391
rect 1721 4386 1722 4390
rect 1726 4386 1727 4390
rect 1731 4386 1732 4390
rect 1736 4386 1737 4390
rect 1741 4386 1742 4390
rect 1746 4386 1747 4390
rect 1751 4386 1752 4390
rect 1756 4386 1757 4390
rect 1761 4386 1762 4390
rect 1717 4385 1762 4386
rect 1721 4381 1722 4385
rect 1726 4381 1727 4385
rect 1731 4381 1732 4385
rect 1736 4381 1737 4385
rect 1741 4381 1742 4385
rect 1746 4381 1747 4385
rect 1751 4381 1752 4385
rect 1756 4381 1757 4385
rect 1761 4381 1762 4385
rect 1717 4380 1762 4381
rect 1721 4376 1722 4380
rect 1726 4376 1727 4380
rect 1731 4376 1732 4380
rect 1736 4376 1737 4380
rect 1741 4376 1742 4380
rect 1746 4376 1747 4380
rect 1751 4376 1752 4380
rect 1756 4376 1757 4380
rect 1761 4376 1762 4380
rect 1717 4375 1762 4376
rect 1721 4371 1722 4375
rect 1726 4371 1727 4375
rect 1731 4371 1732 4375
rect 1736 4371 1737 4375
rect 1741 4371 1742 4375
rect 1746 4371 1747 4375
rect 1751 4371 1752 4375
rect 1756 4371 1757 4375
rect 1761 4371 1762 4375
rect 1717 4370 1762 4371
rect 1721 4366 1722 4370
rect 1726 4366 1727 4370
rect 1731 4366 1732 4370
rect 1736 4366 1737 4370
rect 1741 4366 1742 4370
rect 1746 4366 1747 4370
rect 1751 4366 1752 4370
rect 1756 4366 1757 4370
rect 1761 4366 1762 4370
rect 1717 4365 1762 4366
rect 1721 4361 1722 4365
rect 1726 4361 1727 4365
rect 1731 4361 1732 4365
rect 1736 4361 1737 4365
rect 1741 4361 1742 4365
rect 1746 4361 1747 4365
rect 1751 4361 1752 4365
rect 1756 4361 1757 4365
rect 1761 4361 1762 4365
rect 1769 4445 1773 4446
rect 1769 4440 1773 4441
rect 1769 4435 1773 4436
rect 1769 4430 1773 4431
rect 1769 4425 1773 4426
rect 1769 4420 1773 4421
rect 1769 4415 1773 4416
rect 1769 4410 1773 4411
rect 1769 4405 1773 4406
rect 1769 4400 1773 4401
rect 1769 4395 1773 4396
rect 1769 4390 1773 4391
rect 1769 4385 1773 4386
rect 1769 4380 1773 4381
rect 1769 4375 1773 4376
rect 1769 4370 1773 4371
rect 1769 4365 1773 4366
rect 1705 4360 1709 4361
rect 1705 4353 1709 4356
rect 1769 4360 1773 4361
rect 1769 4353 1773 4356
rect 1709 4349 1712 4353
rect 1716 4349 1717 4353
rect 1721 4349 1722 4353
rect 1726 4349 1727 4353
rect 1731 4349 1732 4353
rect 1736 4349 1737 4353
rect 1741 4349 1742 4353
rect 1746 4349 1747 4353
rect 1751 4349 1752 4353
rect 1756 4349 1757 4353
rect 1761 4349 1762 4353
rect 1766 4349 1769 4353
rect 1782 4465 1786 4466
rect 1782 4460 1786 4461
rect 1782 4455 1786 4456
rect 1782 4450 1786 4451
rect 1782 4445 1786 4446
rect 1782 4440 1786 4441
rect 1782 4435 1786 4436
rect 1782 4430 1786 4431
rect 1782 4425 1786 4426
rect 1782 4420 1786 4421
rect 1782 4415 1786 4416
rect 1782 4410 1786 4411
rect 1782 4405 1786 4406
rect 1782 4400 1786 4401
rect 1782 4395 1786 4396
rect 1782 4390 1786 4391
rect 1782 4385 1786 4386
rect 1782 4380 1786 4381
rect 1782 4375 1786 4376
rect 1782 4370 1786 4371
rect 1782 4365 1786 4366
rect 1782 4360 1786 4361
rect 1782 4355 1786 4356
rect 1782 4350 1786 4351
rect 1692 4345 1696 4346
rect 1692 4340 1696 4341
rect 1782 4345 1786 4346
rect 1782 4340 1786 4341
rect 1696 4336 1697 4340
rect 1701 4336 1702 4340
rect 1706 4336 1707 4340
rect 1711 4336 1712 4340
rect 1716 4336 1717 4340
rect 1721 4336 1722 4340
rect 1726 4336 1727 4340
rect 1731 4336 1732 4340
rect 1736 4336 1737 4340
rect 1741 4336 1742 4340
rect 1746 4336 1747 4340
rect 1751 4336 1752 4340
rect 1756 4336 1757 4340
rect 1761 4336 1762 4340
rect 1766 4336 1767 4340
rect 1771 4336 1772 4340
rect 1776 4336 1777 4340
rect 1781 4336 1782 4340
rect 1793 4333 1845 4599
rect 1984 4624 1985 4628
rect 1989 4624 1990 4628
rect 1994 4624 1995 4628
rect 1980 4623 1999 4624
rect 1984 4619 1985 4623
rect 1989 4619 1990 4623
rect 1994 4619 1995 4623
rect 1980 4618 1999 4619
rect 1984 4614 1985 4618
rect 1989 4614 1990 4618
rect 1994 4614 1995 4618
rect 1980 4613 1999 4614
rect 1984 4609 1985 4613
rect 1989 4609 1990 4613
rect 1994 4609 1995 4613
rect 1980 4608 1999 4609
rect 1984 4604 1985 4608
rect 1989 4604 1990 4608
rect 1994 4604 1995 4608
rect 1980 4603 1999 4604
rect 1984 4599 1985 4603
rect 1989 4599 1990 4603
rect 1994 4599 1995 4603
rect 1980 4598 1999 4599
rect 1984 4594 1985 4598
rect 1989 4594 1990 4598
rect 1994 4594 1995 4598
rect 2002 4601 2058 4602
rect 2002 4597 2004 4601
rect 2008 4597 2009 4601
rect 2013 4597 2014 4601
rect 2018 4597 2019 4601
rect 2023 4597 2024 4601
rect 2028 4597 2029 4601
rect 2033 4597 2034 4601
rect 2038 4597 2039 4601
rect 2043 4597 2044 4601
rect 2048 4597 2049 4601
rect 2053 4597 2054 4601
rect 2002 4596 2058 4597
rect 2002 4592 2004 4596
rect 2008 4592 2009 4596
rect 2013 4592 2014 4596
rect 2018 4592 2019 4596
rect 2023 4592 2024 4596
rect 2028 4592 2029 4596
rect 2033 4592 2034 4596
rect 2038 4592 2039 4596
rect 2043 4592 2044 4596
rect 2048 4592 2049 4596
rect 2053 4592 2054 4596
rect 1887 4578 1955 4580
rect 1887 4574 1945 4578
rect 1949 4574 1950 4578
rect 1954 4574 1955 4578
rect 1887 4573 1955 4574
rect 1887 4569 1945 4573
rect 1949 4569 1950 4573
rect 1954 4569 1955 4573
rect 1887 4568 1955 4569
rect 1887 4564 1945 4568
rect 1949 4564 1950 4568
rect 1954 4564 1955 4568
rect 1887 4563 1955 4564
rect 1887 4559 1945 4563
rect 1949 4559 1950 4563
rect 1954 4559 1955 4563
rect 1887 4558 1955 4559
rect 1887 4554 1945 4558
rect 1949 4554 1950 4558
rect 1954 4554 1955 4558
rect 1887 4553 1955 4554
rect 1887 4549 1945 4553
rect 1949 4549 1950 4553
rect 1954 4549 1955 4553
rect 1887 4548 1955 4549
rect 1984 4578 1985 4582
rect 1989 4578 1990 4582
rect 1994 4578 1995 4582
rect 1980 4577 1999 4578
rect 1984 4573 1985 4577
rect 1989 4573 1990 4577
rect 1994 4573 1995 4577
rect 1980 4572 1999 4573
rect 1984 4568 1985 4572
rect 1989 4568 1990 4572
rect 1994 4568 1995 4572
rect 1980 4567 1999 4568
rect 1984 4563 1985 4567
rect 1989 4563 1990 4567
rect 1994 4563 1995 4567
rect 1980 4562 1999 4563
rect 1984 4558 1985 4562
rect 1989 4558 1990 4562
rect 1994 4558 1995 4562
rect 1980 4557 1999 4558
rect 1984 4553 1985 4557
rect 1989 4553 1990 4557
rect 1994 4553 1995 4557
rect 1980 4552 1999 4553
rect 1984 4548 1985 4552
rect 1989 4548 1990 4552
rect 1994 4548 1995 4552
rect 1887 4544 1945 4548
rect 1949 4544 1950 4548
rect 1954 4544 1955 4548
rect 1887 4543 1955 4544
rect 1887 4539 1945 4543
rect 1949 4539 1950 4543
rect 1954 4539 1955 4543
rect 1887 4538 1955 4539
rect 1887 4534 1945 4538
rect 1949 4534 1950 4538
rect 1954 4534 1955 4538
rect 1887 4533 1955 4534
rect 1887 4529 1945 4533
rect 1949 4529 1950 4533
rect 1954 4529 1955 4533
rect 1887 4528 1955 4529
rect 1887 4524 1945 4528
rect 1949 4524 1950 4528
rect 1954 4524 1955 4528
rect 1887 4523 1955 4524
rect 1887 4519 1945 4523
rect 1949 4519 1950 4523
rect 1954 4519 1955 4523
rect 1887 4518 1955 4519
rect 1887 4514 1945 4518
rect 1949 4514 1950 4518
rect 1954 4514 1955 4518
rect 1887 4512 1955 4514
rect 2002 4535 2058 4592
rect 2002 4531 2067 4535
rect 2002 4519 2058 4531
rect 2119 4527 2132 4703
rect 2293 4624 2294 4628
rect 2298 4624 2299 4628
rect 2303 4624 2304 4628
rect 2289 4623 2308 4624
rect 2293 4619 2294 4623
rect 2298 4619 2299 4623
rect 2303 4619 2304 4623
rect 2289 4618 2308 4619
rect 2293 4614 2294 4618
rect 2298 4614 2299 4618
rect 2303 4614 2304 4618
rect 2289 4613 2308 4614
rect 2293 4609 2294 4613
rect 2298 4609 2299 4613
rect 2303 4609 2304 4613
rect 2289 4608 2308 4609
rect 2293 4604 2294 4608
rect 2298 4604 2299 4608
rect 2303 4604 2304 4608
rect 2289 4603 2308 4604
rect 2293 4599 2294 4603
rect 2298 4599 2299 4603
rect 2303 4599 2304 4603
rect 2289 4598 2308 4599
rect 2293 4594 2294 4598
rect 2298 4594 2299 4598
rect 2303 4594 2304 4598
rect 2311 4601 2367 4602
rect 2311 4597 2313 4601
rect 2317 4597 2318 4601
rect 2322 4597 2323 4601
rect 2327 4597 2328 4601
rect 2332 4597 2333 4601
rect 2337 4597 2338 4601
rect 2342 4597 2343 4601
rect 2347 4597 2348 4601
rect 2352 4597 2353 4601
rect 2357 4597 2358 4601
rect 2362 4597 2363 4601
rect 2311 4596 2367 4597
rect 2311 4592 2313 4596
rect 2317 4592 2318 4596
rect 2322 4592 2323 4596
rect 2327 4592 2328 4596
rect 2332 4592 2333 4596
rect 2337 4592 2338 4596
rect 2342 4592 2343 4596
rect 2347 4592 2348 4596
rect 2352 4592 2353 4596
rect 2357 4592 2358 4596
rect 2362 4592 2363 4596
rect 2196 4578 2264 4580
rect 2196 4574 2254 4578
rect 2258 4574 2259 4578
rect 2263 4574 2264 4578
rect 2196 4573 2264 4574
rect 2196 4569 2254 4573
rect 2258 4569 2259 4573
rect 2263 4569 2264 4573
rect 2196 4568 2264 4569
rect 2196 4564 2254 4568
rect 2258 4564 2259 4568
rect 2263 4564 2264 4568
rect 2196 4563 2264 4564
rect 2196 4559 2254 4563
rect 2258 4559 2259 4563
rect 2263 4559 2264 4563
rect 2196 4558 2264 4559
rect 2196 4554 2254 4558
rect 2258 4554 2259 4558
rect 2263 4554 2264 4558
rect 2196 4553 2264 4554
rect 2196 4549 2254 4553
rect 2258 4549 2259 4553
rect 2263 4549 2264 4553
rect 2196 4548 2264 4549
rect 2293 4578 2294 4582
rect 2298 4578 2299 4582
rect 2303 4578 2304 4582
rect 2289 4577 2308 4578
rect 2293 4573 2294 4577
rect 2298 4573 2299 4577
rect 2303 4573 2304 4577
rect 2289 4572 2308 4573
rect 2293 4568 2294 4572
rect 2298 4568 2299 4572
rect 2303 4568 2304 4572
rect 2289 4567 2308 4568
rect 2293 4563 2294 4567
rect 2298 4563 2299 4567
rect 2303 4563 2304 4567
rect 2289 4562 2308 4563
rect 2293 4558 2294 4562
rect 2298 4558 2299 4562
rect 2303 4558 2304 4562
rect 2289 4557 2308 4558
rect 2293 4553 2294 4557
rect 2298 4553 2299 4557
rect 2303 4553 2304 4557
rect 2289 4552 2308 4553
rect 2293 4548 2294 4552
rect 2298 4548 2299 4552
rect 2303 4548 2304 4552
rect 2196 4544 2254 4548
rect 2258 4544 2259 4548
rect 2263 4544 2264 4548
rect 2196 4543 2264 4544
rect 2196 4539 2254 4543
rect 2258 4539 2259 4543
rect 2263 4539 2264 4543
rect 2196 4538 2264 4539
rect 2196 4535 2254 4538
rect 2193 4534 2254 4535
rect 2258 4534 2259 4538
rect 2263 4534 2264 4538
rect 2193 4533 2264 4534
rect 2193 4531 2254 4533
rect 2196 4529 2254 4531
rect 2258 4529 2259 4533
rect 2263 4529 2264 4533
rect 2196 4528 2264 4529
rect 2107 4523 2137 4527
rect 2196 4524 2254 4528
rect 2258 4524 2259 4528
rect 2263 4524 2264 4528
rect 2196 4523 2264 4524
rect 2002 4515 2067 4519
rect 1887 4475 1943 4512
rect 2002 4503 2058 4515
rect 2110 4514 2133 4523
rect 2196 4519 2254 4523
rect 2258 4519 2259 4523
rect 2263 4519 2264 4523
rect 2193 4518 2264 4519
rect 2193 4515 2254 4518
rect 2110 4511 2114 4514
rect 2107 4507 2114 4511
rect 2126 4511 2133 4514
rect 2196 4514 2254 4515
rect 2258 4514 2259 4518
rect 2263 4514 2264 4518
rect 2196 4512 2264 4514
rect 2311 4535 2367 4592
rect 2311 4531 2376 4535
rect 2311 4519 2367 4531
rect 2428 4527 2441 4705
rect 2602 4624 2603 4628
rect 2607 4624 2608 4628
rect 2612 4624 2613 4628
rect 2598 4623 2617 4624
rect 2602 4619 2603 4623
rect 2607 4619 2608 4623
rect 2612 4619 2613 4623
rect 2598 4618 2617 4619
rect 2602 4614 2603 4618
rect 2607 4614 2608 4618
rect 2612 4614 2613 4618
rect 2598 4613 2617 4614
rect 2602 4609 2603 4613
rect 2607 4609 2608 4613
rect 2612 4609 2613 4613
rect 2598 4608 2617 4609
rect 2602 4604 2603 4608
rect 2607 4604 2608 4608
rect 2612 4604 2613 4608
rect 2598 4603 2617 4604
rect 2602 4599 2603 4603
rect 2607 4599 2608 4603
rect 2612 4599 2613 4603
rect 2598 4598 2617 4599
rect 2602 4594 2603 4598
rect 2607 4594 2608 4598
rect 2612 4594 2613 4598
rect 2620 4601 2676 4602
rect 2620 4597 2622 4601
rect 2626 4597 2627 4601
rect 2631 4597 2632 4601
rect 2636 4597 2637 4601
rect 2641 4597 2642 4601
rect 2646 4597 2647 4601
rect 2651 4597 2652 4601
rect 2656 4597 2657 4601
rect 2661 4597 2662 4601
rect 2666 4597 2667 4601
rect 2671 4597 2672 4601
rect 2620 4596 2676 4597
rect 2620 4592 2622 4596
rect 2626 4592 2627 4596
rect 2631 4592 2632 4596
rect 2636 4592 2637 4596
rect 2641 4592 2642 4596
rect 2646 4592 2647 4596
rect 2651 4592 2652 4596
rect 2656 4592 2657 4596
rect 2661 4592 2662 4596
rect 2666 4592 2667 4596
rect 2671 4592 2672 4596
rect 2505 4578 2573 4580
rect 2505 4574 2563 4578
rect 2567 4574 2568 4578
rect 2572 4574 2573 4578
rect 2505 4573 2573 4574
rect 2505 4569 2563 4573
rect 2567 4569 2568 4573
rect 2572 4569 2573 4573
rect 2505 4568 2573 4569
rect 2505 4564 2563 4568
rect 2567 4564 2568 4568
rect 2572 4564 2573 4568
rect 2505 4563 2573 4564
rect 2505 4559 2563 4563
rect 2567 4559 2568 4563
rect 2572 4559 2573 4563
rect 2505 4558 2573 4559
rect 2505 4554 2563 4558
rect 2567 4554 2568 4558
rect 2572 4554 2573 4558
rect 2505 4553 2573 4554
rect 2505 4549 2563 4553
rect 2567 4549 2568 4553
rect 2572 4549 2573 4553
rect 2505 4548 2573 4549
rect 2602 4578 2603 4582
rect 2607 4578 2608 4582
rect 2612 4578 2613 4582
rect 2598 4577 2617 4578
rect 2602 4573 2603 4577
rect 2607 4573 2608 4577
rect 2612 4573 2613 4577
rect 2598 4572 2617 4573
rect 2602 4568 2603 4572
rect 2607 4568 2608 4572
rect 2612 4568 2613 4572
rect 2598 4567 2617 4568
rect 2602 4563 2603 4567
rect 2607 4563 2608 4567
rect 2612 4563 2613 4567
rect 2598 4562 2617 4563
rect 2602 4558 2603 4562
rect 2607 4558 2608 4562
rect 2612 4558 2613 4562
rect 2598 4557 2617 4558
rect 2602 4553 2603 4557
rect 2607 4553 2608 4557
rect 2612 4553 2613 4557
rect 2598 4552 2617 4553
rect 2602 4548 2603 4552
rect 2607 4548 2608 4552
rect 2612 4548 2613 4552
rect 2505 4544 2563 4548
rect 2567 4544 2568 4548
rect 2572 4544 2573 4548
rect 2505 4543 2573 4544
rect 2505 4539 2563 4543
rect 2567 4539 2568 4543
rect 2572 4539 2573 4543
rect 2505 4538 2573 4539
rect 2505 4535 2563 4538
rect 2502 4534 2563 4535
rect 2567 4534 2568 4538
rect 2572 4534 2573 4538
rect 2502 4533 2573 4534
rect 2502 4531 2563 4533
rect 2505 4529 2563 4531
rect 2567 4529 2568 4533
rect 2572 4529 2573 4533
rect 2505 4528 2573 4529
rect 2416 4523 2446 4527
rect 2505 4524 2563 4528
rect 2567 4524 2568 4528
rect 2572 4524 2573 4528
rect 2505 4523 2573 4524
rect 2311 4515 2376 4519
rect 2126 4507 2137 4511
rect 2002 4499 2067 4503
rect 2196 4503 2252 4512
rect 2002 4487 2058 4499
rect 2119 4495 2123 4502
rect 2193 4499 2252 4503
rect 2107 4491 2137 4495
rect 2196 4487 2252 4499
rect 2002 4483 2067 4487
rect 2193 4483 2252 4487
rect 2002 4475 2058 4483
rect 1856 4471 1857 4475
rect 1861 4471 1862 4475
rect 1866 4471 1867 4475
rect 1871 4471 1872 4475
rect 1876 4471 1877 4475
rect 1881 4471 1882 4475
rect 1886 4471 1887 4475
rect 1891 4471 1892 4475
rect 1896 4471 1897 4475
rect 1901 4471 1902 4475
rect 1906 4471 1907 4475
rect 1911 4471 1912 4475
rect 1916 4471 1917 4475
rect 1921 4471 1922 4475
rect 1926 4471 1927 4475
rect 1931 4471 1932 4475
rect 1936 4471 1937 4475
rect 1941 4471 1942 4475
rect 1852 4470 1856 4471
rect 1942 4470 1946 4471
rect 1852 4465 1856 4466
rect 1852 4460 1856 4461
rect 1852 4455 1856 4456
rect 1852 4450 1856 4451
rect 1852 4445 1856 4446
rect 1852 4440 1856 4441
rect 1852 4435 1856 4436
rect 1852 4430 1856 4431
rect 1852 4425 1856 4426
rect 1852 4420 1856 4421
rect 1852 4415 1856 4416
rect 1852 4410 1856 4411
rect 1852 4405 1856 4406
rect 1852 4400 1856 4401
rect 1852 4395 1856 4396
rect 1852 4390 1856 4391
rect 1852 4385 1856 4386
rect 1852 4380 1856 4381
rect 1852 4375 1856 4376
rect 1852 4370 1856 4371
rect 1852 4365 1856 4366
rect 1852 4360 1856 4361
rect 1852 4355 1856 4356
rect 1852 4350 1856 4351
rect 1869 4458 1872 4466
rect 1876 4458 1877 4466
rect 1881 4458 1882 4466
rect 1886 4458 1887 4466
rect 1891 4458 1892 4466
rect 1896 4458 1897 4466
rect 1901 4458 1902 4466
rect 1906 4458 1907 4466
rect 1911 4458 1912 4466
rect 1916 4458 1917 4466
rect 1921 4458 1922 4466
rect 1926 4458 1929 4466
rect 1865 4455 1869 4458
rect 1865 4450 1869 4451
rect 1929 4455 1933 4458
rect 1929 4450 1933 4451
rect 1865 4445 1869 4446
rect 1865 4440 1869 4441
rect 1865 4435 1869 4436
rect 1865 4430 1869 4431
rect 1865 4425 1869 4426
rect 1865 4420 1869 4421
rect 1865 4415 1869 4416
rect 1865 4410 1869 4411
rect 1865 4405 1869 4406
rect 1865 4400 1869 4401
rect 1865 4395 1869 4396
rect 1865 4390 1869 4391
rect 1865 4385 1869 4386
rect 1865 4380 1869 4381
rect 1865 4375 1869 4376
rect 1865 4370 1869 4371
rect 1865 4365 1869 4366
rect 1881 4446 1882 4450
rect 1886 4446 1887 4450
rect 1891 4446 1892 4450
rect 1896 4446 1897 4450
rect 1901 4446 1902 4450
rect 1906 4446 1907 4450
rect 1911 4446 1912 4450
rect 1916 4446 1917 4450
rect 1877 4445 1921 4446
rect 1881 4441 1882 4445
rect 1886 4441 1887 4445
rect 1891 4441 1892 4445
rect 1896 4441 1897 4445
rect 1901 4441 1902 4445
rect 1906 4441 1907 4445
rect 1911 4441 1912 4445
rect 1916 4441 1917 4445
rect 1877 4440 1921 4441
rect 1881 4436 1882 4440
rect 1886 4436 1887 4440
rect 1891 4436 1892 4440
rect 1896 4436 1897 4440
rect 1901 4436 1902 4440
rect 1906 4436 1907 4440
rect 1911 4436 1912 4440
rect 1916 4436 1917 4440
rect 1877 4435 1921 4436
rect 1881 4431 1882 4435
rect 1886 4431 1887 4435
rect 1891 4431 1892 4435
rect 1896 4431 1897 4435
rect 1901 4431 1902 4435
rect 1906 4431 1907 4435
rect 1911 4431 1912 4435
rect 1916 4431 1917 4435
rect 1877 4430 1921 4431
rect 1881 4426 1882 4430
rect 1886 4426 1887 4430
rect 1891 4426 1892 4430
rect 1896 4426 1897 4430
rect 1901 4426 1902 4430
rect 1906 4426 1907 4430
rect 1911 4426 1912 4430
rect 1916 4426 1917 4430
rect 1877 4425 1921 4426
rect 1881 4421 1882 4425
rect 1886 4421 1887 4425
rect 1891 4421 1892 4425
rect 1896 4421 1897 4425
rect 1901 4421 1902 4425
rect 1906 4421 1907 4425
rect 1911 4421 1912 4425
rect 1916 4421 1917 4425
rect 1877 4420 1921 4421
rect 1881 4416 1882 4420
rect 1886 4416 1887 4420
rect 1891 4416 1892 4420
rect 1896 4416 1897 4420
rect 1901 4416 1902 4420
rect 1906 4416 1907 4420
rect 1911 4416 1912 4420
rect 1916 4416 1917 4420
rect 1877 4415 1921 4416
rect 1881 4411 1882 4415
rect 1886 4411 1887 4415
rect 1891 4411 1892 4415
rect 1896 4411 1897 4415
rect 1901 4411 1902 4415
rect 1906 4411 1907 4415
rect 1911 4411 1912 4415
rect 1916 4411 1917 4415
rect 1877 4410 1921 4411
rect 1881 4406 1882 4410
rect 1886 4406 1887 4410
rect 1891 4406 1892 4410
rect 1896 4406 1897 4410
rect 1901 4406 1902 4410
rect 1906 4406 1907 4410
rect 1911 4406 1912 4410
rect 1916 4406 1917 4410
rect 1877 4405 1921 4406
rect 1881 4401 1882 4405
rect 1886 4401 1887 4405
rect 1891 4401 1892 4405
rect 1896 4401 1897 4405
rect 1901 4401 1902 4405
rect 1906 4401 1907 4405
rect 1911 4401 1912 4405
rect 1916 4401 1917 4405
rect 1877 4400 1921 4401
rect 1881 4396 1882 4400
rect 1886 4396 1887 4400
rect 1891 4396 1892 4400
rect 1896 4396 1897 4400
rect 1901 4396 1902 4400
rect 1906 4396 1907 4400
rect 1911 4396 1912 4400
rect 1916 4396 1917 4400
rect 1877 4395 1921 4396
rect 1881 4391 1882 4395
rect 1886 4391 1887 4395
rect 1891 4391 1892 4395
rect 1896 4391 1897 4395
rect 1901 4391 1902 4395
rect 1906 4391 1907 4395
rect 1911 4391 1912 4395
rect 1916 4391 1917 4395
rect 1877 4390 1921 4391
rect 1881 4386 1882 4390
rect 1886 4386 1887 4390
rect 1891 4386 1892 4390
rect 1896 4386 1897 4390
rect 1901 4386 1902 4390
rect 1906 4386 1907 4390
rect 1911 4386 1912 4390
rect 1916 4386 1917 4390
rect 1877 4385 1921 4386
rect 1881 4381 1882 4385
rect 1886 4381 1887 4385
rect 1891 4381 1892 4385
rect 1896 4381 1897 4385
rect 1901 4381 1902 4385
rect 1906 4381 1907 4385
rect 1911 4381 1912 4385
rect 1916 4381 1917 4385
rect 1877 4380 1921 4381
rect 1881 4376 1882 4380
rect 1886 4376 1887 4380
rect 1891 4376 1892 4380
rect 1896 4376 1897 4380
rect 1901 4376 1902 4380
rect 1906 4376 1907 4380
rect 1911 4376 1912 4380
rect 1916 4376 1917 4380
rect 1877 4375 1921 4376
rect 1881 4371 1882 4375
rect 1886 4371 1887 4375
rect 1891 4371 1892 4375
rect 1896 4371 1897 4375
rect 1901 4371 1902 4375
rect 1906 4371 1907 4375
rect 1911 4371 1912 4375
rect 1916 4371 1917 4375
rect 1877 4370 1921 4371
rect 1881 4366 1882 4370
rect 1886 4366 1887 4370
rect 1891 4366 1892 4370
rect 1896 4366 1897 4370
rect 1901 4366 1902 4370
rect 1906 4366 1907 4370
rect 1911 4366 1912 4370
rect 1916 4366 1917 4370
rect 1877 4365 1921 4366
rect 1881 4361 1882 4365
rect 1886 4361 1887 4365
rect 1891 4361 1892 4365
rect 1896 4361 1897 4365
rect 1901 4361 1902 4365
rect 1906 4361 1907 4365
rect 1911 4361 1912 4365
rect 1916 4361 1917 4365
rect 1929 4445 1933 4446
rect 1929 4440 1933 4441
rect 1929 4435 1933 4436
rect 1929 4430 1933 4431
rect 1929 4425 1933 4426
rect 1929 4420 1933 4421
rect 1929 4415 1933 4416
rect 1929 4410 1933 4411
rect 1929 4405 1933 4406
rect 1929 4400 1933 4401
rect 1929 4395 1933 4396
rect 1929 4390 1933 4391
rect 1929 4385 1933 4386
rect 1929 4380 1933 4381
rect 1929 4375 1933 4376
rect 1929 4370 1933 4371
rect 1929 4365 1933 4366
rect 1865 4360 1869 4361
rect 1865 4353 1869 4356
rect 1929 4360 1933 4361
rect 1929 4353 1933 4356
rect 1869 4349 1872 4353
rect 1876 4349 1877 4353
rect 1881 4349 1882 4353
rect 1886 4349 1887 4353
rect 1891 4349 1892 4353
rect 1896 4349 1897 4353
rect 1901 4349 1902 4353
rect 1906 4349 1907 4353
rect 1911 4349 1912 4353
rect 1916 4349 1917 4353
rect 1921 4349 1922 4353
rect 1926 4349 1929 4353
rect 1942 4465 1946 4466
rect 1942 4460 1946 4461
rect 1942 4455 1946 4456
rect 1942 4450 1946 4451
rect 1942 4445 1946 4446
rect 1942 4440 1946 4441
rect 1942 4435 1946 4436
rect 1942 4430 1946 4431
rect 1942 4425 1946 4426
rect 1942 4420 1946 4421
rect 1942 4415 1946 4416
rect 1942 4410 1946 4411
rect 1942 4405 1946 4406
rect 1942 4400 1946 4401
rect 1942 4395 1946 4396
rect 1942 4390 1946 4391
rect 1942 4385 1946 4386
rect 1942 4380 1946 4381
rect 1942 4375 1946 4376
rect 1942 4370 1946 4371
rect 1942 4365 1946 4366
rect 1942 4360 1946 4361
rect 1942 4355 1946 4356
rect 1942 4350 1946 4351
rect 1852 4345 1856 4346
rect 1852 4340 1856 4341
rect 1942 4345 1946 4346
rect 1942 4340 1946 4341
rect 1856 4336 1857 4340
rect 1861 4336 1862 4340
rect 1866 4336 1867 4340
rect 1871 4336 1872 4340
rect 1876 4336 1877 4340
rect 1881 4336 1882 4340
rect 1886 4336 1887 4340
rect 1891 4336 1892 4340
rect 1896 4336 1897 4340
rect 1901 4336 1902 4340
rect 1906 4336 1907 4340
rect 1911 4336 1912 4340
rect 1916 4336 1917 4340
rect 1921 4336 1922 4340
rect 1926 4336 1927 4340
rect 1931 4336 1932 4340
rect 1936 4336 1937 4340
rect 1941 4336 1942 4340
rect 2005 4471 2006 4475
rect 2010 4471 2011 4475
rect 2015 4471 2016 4475
rect 2020 4471 2021 4475
rect 2025 4471 2026 4475
rect 2030 4471 2031 4475
rect 2035 4471 2036 4475
rect 2040 4471 2041 4475
rect 2045 4471 2046 4475
rect 2050 4471 2051 4475
rect 2055 4471 2056 4475
rect 2060 4471 2061 4475
rect 2065 4471 2066 4475
rect 2070 4471 2071 4475
rect 2075 4471 2076 4475
rect 2080 4471 2081 4475
rect 2085 4471 2086 4475
rect 2090 4471 2091 4475
rect 2124 4472 2133 4483
rect 2196 4475 2252 4483
rect 2311 4503 2367 4515
rect 2419 4514 2442 4523
rect 2505 4519 2563 4523
rect 2567 4519 2568 4523
rect 2572 4519 2573 4523
rect 2502 4518 2573 4519
rect 2502 4515 2563 4518
rect 2419 4511 2423 4514
rect 2416 4507 2423 4511
rect 2435 4511 2442 4514
rect 2505 4514 2563 4515
rect 2567 4514 2568 4518
rect 2572 4514 2573 4518
rect 2505 4512 2573 4514
rect 2620 4535 2676 4592
rect 2620 4531 2685 4535
rect 2620 4519 2676 4531
rect 2737 4527 2750 4717
rect 2911 4624 2912 4628
rect 2916 4624 2917 4628
rect 2921 4624 2922 4628
rect 2907 4623 2926 4624
rect 2911 4619 2912 4623
rect 2916 4619 2917 4623
rect 2921 4619 2922 4623
rect 2907 4618 2926 4619
rect 2911 4614 2912 4618
rect 2916 4614 2917 4618
rect 2921 4614 2922 4618
rect 2907 4613 2926 4614
rect 2911 4609 2912 4613
rect 2916 4609 2917 4613
rect 2921 4609 2922 4613
rect 2907 4608 2926 4609
rect 2911 4604 2912 4608
rect 2916 4604 2917 4608
rect 2921 4604 2922 4608
rect 2907 4603 2926 4604
rect 2911 4599 2912 4603
rect 2916 4599 2917 4603
rect 2921 4599 2922 4603
rect 2907 4598 2926 4599
rect 2911 4594 2912 4598
rect 2916 4594 2917 4598
rect 2921 4594 2922 4598
rect 2929 4601 2985 4602
rect 2929 4597 2931 4601
rect 2935 4597 2936 4601
rect 2940 4597 2941 4601
rect 2945 4597 2946 4601
rect 2950 4597 2951 4601
rect 2955 4597 2956 4601
rect 2960 4597 2961 4601
rect 2965 4597 2966 4601
rect 2970 4597 2971 4601
rect 2975 4597 2976 4601
rect 2980 4597 2981 4601
rect 2929 4596 2985 4597
rect 2929 4592 2931 4596
rect 2935 4592 2936 4596
rect 2940 4592 2941 4596
rect 2945 4592 2946 4596
rect 2950 4592 2951 4596
rect 2955 4592 2956 4596
rect 2960 4592 2961 4596
rect 2965 4592 2966 4596
rect 2970 4592 2971 4596
rect 2975 4592 2976 4596
rect 2980 4592 2981 4596
rect 2814 4578 2882 4580
rect 2814 4574 2872 4578
rect 2876 4574 2877 4578
rect 2881 4574 2882 4578
rect 2814 4573 2882 4574
rect 2814 4569 2872 4573
rect 2876 4569 2877 4573
rect 2881 4569 2882 4573
rect 2814 4568 2882 4569
rect 2814 4564 2872 4568
rect 2876 4564 2877 4568
rect 2881 4564 2882 4568
rect 2814 4563 2882 4564
rect 2814 4559 2872 4563
rect 2876 4559 2877 4563
rect 2881 4559 2882 4563
rect 2814 4558 2882 4559
rect 2814 4554 2872 4558
rect 2876 4554 2877 4558
rect 2881 4554 2882 4558
rect 2814 4553 2882 4554
rect 2814 4549 2872 4553
rect 2876 4549 2877 4553
rect 2881 4549 2882 4553
rect 2814 4548 2882 4549
rect 2911 4578 2912 4582
rect 2916 4578 2917 4582
rect 2921 4578 2922 4582
rect 2907 4577 2926 4578
rect 2911 4573 2912 4577
rect 2916 4573 2917 4577
rect 2921 4573 2922 4577
rect 2907 4572 2926 4573
rect 2911 4568 2912 4572
rect 2916 4568 2917 4572
rect 2921 4568 2922 4572
rect 2907 4567 2926 4568
rect 2911 4563 2912 4567
rect 2916 4563 2917 4567
rect 2921 4563 2922 4567
rect 2907 4562 2926 4563
rect 2911 4558 2912 4562
rect 2916 4558 2917 4562
rect 2921 4558 2922 4562
rect 2907 4557 2926 4558
rect 2911 4553 2912 4557
rect 2916 4553 2917 4557
rect 2921 4553 2922 4557
rect 2907 4552 2926 4553
rect 2911 4548 2912 4552
rect 2916 4548 2917 4552
rect 2921 4548 2922 4552
rect 2814 4544 2872 4548
rect 2876 4544 2877 4548
rect 2881 4544 2882 4548
rect 2814 4543 2882 4544
rect 2814 4539 2872 4543
rect 2876 4539 2877 4543
rect 2881 4539 2882 4543
rect 2814 4538 2882 4539
rect 2814 4535 2872 4538
rect 2811 4534 2872 4535
rect 2876 4534 2877 4538
rect 2881 4534 2882 4538
rect 2811 4533 2882 4534
rect 2811 4531 2872 4533
rect 2814 4529 2872 4531
rect 2876 4529 2877 4533
rect 2881 4529 2882 4533
rect 2814 4528 2882 4529
rect 2725 4523 2755 4527
rect 2814 4524 2872 4528
rect 2876 4524 2877 4528
rect 2881 4524 2882 4528
rect 2814 4523 2882 4524
rect 2620 4515 2685 4519
rect 2435 4507 2446 4511
rect 2311 4499 2376 4503
rect 2505 4503 2561 4512
rect 2311 4487 2367 4499
rect 2428 4495 2432 4502
rect 2502 4499 2561 4503
rect 2416 4491 2446 4495
rect 2505 4487 2561 4499
rect 2311 4483 2376 4487
rect 2502 4483 2561 4487
rect 2311 4475 2367 4483
rect 2001 4470 2005 4471
rect 2091 4470 2095 4471
rect 2122 4470 2135 4472
rect 2165 4471 2166 4475
rect 2170 4471 2171 4475
rect 2175 4471 2176 4475
rect 2180 4471 2181 4475
rect 2185 4471 2186 4475
rect 2190 4471 2191 4475
rect 2195 4471 2196 4475
rect 2200 4471 2201 4475
rect 2205 4471 2206 4475
rect 2210 4471 2211 4475
rect 2215 4471 2216 4475
rect 2220 4471 2221 4475
rect 2225 4471 2226 4475
rect 2230 4471 2231 4475
rect 2235 4471 2236 4475
rect 2240 4471 2241 4475
rect 2245 4471 2246 4475
rect 2250 4471 2251 4475
rect 2161 4470 2165 4471
rect 2120 4468 2137 4470
rect 2001 4465 2005 4466
rect 2001 4460 2005 4461
rect 2001 4455 2005 4456
rect 2001 4450 2005 4451
rect 2001 4445 2005 4446
rect 2001 4440 2005 4441
rect 2001 4435 2005 4436
rect 2001 4430 2005 4431
rect 2001 4425 2005 4426
rect 2001 4420 2005 4421
rect 2001 4415 2005 4416
rect 2001 4410 2005 4411
rect 2001 4405 2005 4406
rect 2001 4400 2005 4401
rect 2001 4395 2005 4396
rect 2001 4390 2005 4391
rect 2001 4385 2005 4386
rect 2001 4380 2005 4381
rect 2001 4375 2005 4376
rect 2001 4370 2005 4371
rect 2001 4365 2005 4366
rect 2001 4360 2005 4361
rect 2001 4355 2005 4356
rect 2001 4350 2005 4351
rect 2018 4458 2021 4466
rect 2025 4458 2026 4466
rect 2030 4458 2031 4466
rect 2035 4458 2036 4466
rect 2040 4458 2041 4466
rect 2045 4458 2046 4466
rect 2050 4458 2051 4466
rect 2055 4458 2056 4466
rect 2060 4458 2061 4466
rect 2065 4458 2066 4466
rect 2070 4458 2071 4466
rect 2075 4458 2078 4466
rect 2014 4455 2018 4458
rect 2014 4450 2018 4451
rect 2078 4455 2082 4458
rect 2078 4450 2082 4451
rect 2014 4445 2018 4446
rect 2014 4440 2018 4441
rect 2014 4435 2018 4436
rect 2014 4430 2018 4431
rect 2014 4425 2018 4426
rect 2014 4420 2018 4421
rect 2014 4415 2018 4416
rect 2014 4410 2018 4411
rect 2014 4405 2018 4406
rect 2014 4400 2018 4401
rect 2014 4395 2018 4396
rect 2014 4390 2018 4391
rect 2014 4385 2018 4386
rect 2014 4380 2018 4381
rect 2014 4375 2018 4376
rect 2014 4370 2018 4371
rect 2014 4365 2018 4366
rect 2030 4446 2031 4450
rect 2035 4446 2036 4450
rect 2040 4446 2041 4450
rect 2045 4446 2046 4450
rect 2050 4446 2051 4450
rect 2055 4446 2056 4450
rect 2060 4446 2061 4450
rect 2065 4446 2066 4450
rect 2070 4446 2071 4450
rect 2026 4445 2071 4446
rect 2030 4441 2031 4445
rect 2035 4441 2036 4445
rect 2040 4441 2041 4445
rect 2045 4441 2046 4445
rect 2050 4441 2051 4445
rect 2055 4441 2056 4445
rect 2060 4441 2061 4445
rect 2065 4441 2066 4445
rect 2070 4441 2071 4445
rect 2026 4440 2071 4441
rect 2030 4436 2031 4440
rect 2035 4436 2036 4440
rect 2040 4436 2041 4440
rect 2045 4436 2046 4440
rect 2050 4436 2051 4440
rect 2055 4436 2056 4440
rect 2060 4436 2061 4440
rect 2065 4436 2066 4440
rect 2070 4436 2071 4440
rect 2026 4435 2071 4436
rect 2030 4431 2031 4435
rect 2035 4431 2036 4435
rect 2040 4431 2041 4435
rect 2045 4431 2046 4435
rect 2050 4431 2051 4435
rect 2055 4431 2056 4435
rect 2060 4431 2061 4435
rect 2065 4431 2066 4435
rect 2070 4431 2071 4435
rect 2026 4430 2071 4431
rect 2030 4426 2031 4430
rect 2035 4426 2036 4430
rect 2040 4426 2041 4430
rect 2045 4426 2046 4430
rect 2050 4426 2051 4430
rect 2055 4426 2056 4430
rect 2060 4426 2061 4430
rect 2065 4426 2066 4430
rect 2070 4426 2071 4430
rect 2026 4425 2071 4426
rect 2030 4421 2031 4425
rect 2035 4421 2036 4425
rect 2040 4421 2041 4425
rect 2045 4421 2046 4425
rect 2050 4421 2051 4425
rect 2055 4421 2056 4425
rect 2060 4421 2061 4425
rect 2065 4421 2066 4425
rect 2070 4421 2071 4425
rect 2026 4420 2071 4421
rect 2030 4416 2031 4420
rect 2035 4416 2036 4420
rect 2040 4416 2041 4420
rect 2045 4416 2046 4420
rect 2050 4416 2051 4420
rect 2055 4416 2056 4420
rect 2060 4416 2061 4420
rect 2065 4416 2066 4420
rect 2070 4416 2071 4420
rect 2026 4415 2071 4416
rect 2030 4411 2031 4415
rect 2035 4411 2036 4415
rect 2040 4411 2041 4415
rect 2045 4411 2046 4415
rect 2050 4411 2051 4415
rect 2055 4411 2056 4415
rect 2060 4411 2061 4415
rect 2065 4411 2066 4415
rect 2070 4411 2071 4415
rect 2026 4410 2071 4411
rect 2030 4406 2031 4410
rect 2035 4406 2036 4410
rect 2040 4406 2041 4410
rect 2045 4406 2046 4410
rect 2050 4406 2051 4410
rect 2055 4406 2056 4410
rect 2060 4406 2061 4410
rect 2065 4406 2066 4410
rect 2070 4406 2071 4410
rect 2026 4405 2071 4406
rect 2030 4401 2031 4405
rect 2035 4401 2036 4405
rect 2040 4401 2041 4405
rect 2045 4401 2046 4405
rect 2050 4401 2051 4405
rect 2055 4401 2056 4405
rect 2060 4401 2061 4405
rect 2065 4401 2066 4405
rect 2070 4401 2071 4405
rect 2026 4400 2071 4401
rect 2030 4396 2031 4400
rect 2035 4396 2036 4400
rect 2040 4396 2041 4400
rect 2045 4396 2046 4400
rect 2050 4396 2051 4400
rect 2055 4396 2056 4400
rect 2060 4396 2061 4400
rect 2065 4396 2066 4400
rect 2070 4396 2071 4400
rect 2026 4395 2071 4396
rect 2030 4391 2031 4395
rect 2035 4391 2036 4395
rect 2040 4391 2041 4395
rect 2045 4391 2046 4395
rect 2050 4391 2051 4395
rect 2055 4391 2056 4395
rect 2060 4391 2061 4395
rect 2065 4391 2066 4395
rect 2070 4391 2071 4395
rect 2026 4390 2071 4391
rect 2030 4386 2031 4390
rect 2035 4386 2036 4390
rect 2040 4386 2041 4390
rect 2045 4386 2046 4390
rect 2050 4386 2051 4390
rect 2055 4386 2056 4390
rect 2060 4386 2061 4390
rect 2065 4386 2066 4390
rect 2070 4386 2071 4390
rect 2026 4385 2071 4386
rect 2030 4381 2031 4385
rect 2035 4381 2036 4385
rect 2040 4381 2041 4385
rect 2045 4381 2046 4385
rect 2050 4381 2051 4385
rect 2055 4381 2056 4385
rect 2060 4381 2061 4385
rect 2065 4381 2066 4385
rect 2070 4381 2071 4385
rect 2026 4380 2071 4381
rect 2030 4376 2031 4380
rect 2035 4376 2036 4380
rect 2040 4376 2041 4380
rect 2045 4376 2046 4380
rect 2050 4376 2051 4380
rect 2055 4376 2056 4380
rect 2060 4376 2061 4380
rect 2065 4376 2066 4380
rect 2070 4376 2071 4380
rect 2026 4375 2071 4376
rect 2030 4371 2031 4375
rect 2035 4371 2036 4375
rect 2040 4371 2041 4375
rect 2045 4371 2046 4375
rect 2050 4371 2051 4375
rect 2055 4371 2056 4375
rect 2060 4371 2061 4375
rect 2065 4371 2066 4375
rect 2070 4371 2071 4375
rect 2026 4370 2071 4371
rect 2030 4366 2031 4370
rect 2035 4366 2036 4370
rect 2040 4366 2041 4370
rect 2045 4366 2046 4370
rect 2050 4366 2051 4370
rect 2055 4366 2056 4370
rect 2060 4366 2061 4370
rect 2065 4366 2066 4370
rect 2070 4366 2071 4370
rect 2026 4365 2071 4366
rect 2030 4361 2031 4365
rect 2035 4361 2036 4365
rect 2040 4361 2041 4365
rect 2045 4361 2046 4365
rect 2050 4361 2051 4365
rect 2055 4361 2056 4365
rect 2060 4361 2061 4365
rect 2065 4361 2066 4365
rect 2070 4361 2071 4365
rect 2078 4445 2082 4446
rect 2078 4440 2082 4441
rect 2078 4435 2082 4436
rect 2078 4430 2082 4431
rect 2078 4425 2082 4426
rect 2078 4420 2082 4421
rect 2078 4415 2082 4416
rect 2078 4410 2082 4411
rect 2078 4405 2082 4406
rect 2078 4400 2082 4401
rect 2078 4395 2082 4396
rect 2078 4390 2082 4391
rect 2078 4385 2082 4386
rect 2078 4380 2082 4381
rect 2078 4375 2082 4376
rect 2078 4370 2082 4371
rect 2078 4365 2082 4366
rect 2014 4360 2018 4361
rect 2014 4353 2018 4356
rect 2078 4360 2082 4361
rect 2078 4353 2082 4356
rect 2018 4349 2021 4353
rect 2025 4349 2026 4353
rect 2030 4349 2031 4353
rect 2035 4349 2036 4353
rect 2040 4349 2041 4353
rect 2045 4349 2046 4353
rect 2050 4349 2051 4353
rect 2055 4349 2056 4353
rect 2060 4349 2061 4353
rect 2065 4349 2066 4353
rect 2070 4349 2071 4353
rect 2075 4349 2078 4353
rect 2091 4465 2095 4466
rect 2091 4460 2095 4461
rect 2091 4455 2095 4456
rect 2091 4450 2095 4451
rect 2091 4445 2095 4446
rect 2091 4440 2095 4441
rect 2091 4435 2095 4436
rect 2118 4440 2139 4468
rect 2251 4470 2255 4471
rect 2161 4465 2165 4466
rect 2161 4460 2165 4461
rect 2161 4455 2165 4456
rect 2161 4450 2165 4451
rect 2161 4445 2165 4446
rect 2161 4440 2165 4441
rect 2161 4435 2165 4436
rect 2091 4430 2095 4431
rect 2091 4425 2095 4426
rect 2091 4420 2095 4421
rect 2091 4415 2095 4416
rect 2091 4410 2095 4411
rect 2091 4405 2095 4406
rect 2091 4400 2095 4401
rect 2091 4395 2095 4396
rect 2091 4390 2095 4391
rect 2091 4385 2095 4386
rect 2091 4380 2095 4381
rect 2091 4375 2095 4376
rect 2091 4370 2095 4371
rect 2091 4365 2095 4366
rect 2161 4430 2165 4431
rect 2161 4425 2165 4426
rect 2161 4420 2165 4421
rect 2161 4415 2165 4416
rect 2161 4410 2165 4411
rect 2161 4405 2165 4406
rect 2161 4400 2165 4401
rect 2161 4395 2165 4396
rect 2161 4390 2165 4391
rect 2161 4385 2165 4386
rect 2161 4380 2165 4381
rect 2161 4375 2165 4376
rect 2161 4370 2165 4371
rect 2161 4365 2165 4366
rect 2091 4360 2095 4361
rect 2091 4355 2095 4356
rect 2091 4350 2095 4351
rect 2001 4345 2005 4346
rect 2001 4340 2005 4341
rect 2091 4345 2095 4346
rect 2091 4340 2095 4341
rect 2005 4336 2006 4340
rect 2010 4336 2011 4340
rect 2015 4336 2016 4340
rect 2020 4336 2021 4340
rect 2025 4336 2026 4340
rect 2030 4336 2031 4340
rect 2035 4336 2036 4340
rect 2040 4336 2041 4340
rect 2045 4336 2046 4340
rect 2050 4336 2051 4340
rect 2055 4336 2056 4340
rect 2060 4336 2061 4340
rect 2065 4336 2066 4340
rect 2070 4336 2071 4340
rect 2075 4336 2076 4340
rect 2080 4336 2081 4340
rect 2085 4336 2086 4340
rect 2090 4336 2091 4340
rect 2118 4333 2139 4353
rect 2161 4360 2165 4361
rect 2161 4355 2165 4356
rect 2161 4350 2165 4351
rect 2178 4458 2181 4466
rect 2185 4458 2186 4466
rect 2190 4458 2191 4466
rect 2195 4458 2196 4466
rect 2200 4458 2201 4466
rect 2205 4458 2206 4466
rect 2210 4458 2211 4466
rect 2215 4458 2216 4466
rect 2220 4458 2221 4466
rect 2225 4458 2226 4466
rect 2230 4458 2231 4466
rect 2235 4458 2238 4466
rect 2174 4455 2178 4458
rect 2174 4450 2178 4451
rect 2238 4455 2242 4458
rect 2238 4450 2242 4451
rect 2174 4445 2178 4446
rect 2174 4440 2178 4441
rect 2174 4435 2178 4436
rect 2174 4430 2178 4431
rect 2174 4425 2178 4426
rect 2174 4420 2178 4421
rect 2174 4415 2178 4416
rect 2174 4410 2178 4411
rect 2174 4405 2178 4406
rect 2174 4400 2178 4401
rect 2174 4395 2178 4396
rect 2174 4390 2178 4391
rect 2174 4385 2178 4386
rect 2174 4380 2178 4381
rect 2174 4375 2178 4376
rect 2174 4370 2178 4371
rect 2174 4365 2178 4366
rect 2190 4446 2191 4450
rect 2195 4446 2196 4450
rect 2200 4446 2201 4450
rect 2205 4446 2206 4450
rect 2210 4446 2211 4450
rect 2215 4446 2216 4450
rect 2220 4446 2221 4450
rect 2225 4446 2226 4450
rect 2186 4445 2230 4446
rect 2190 4441 2191 4445
rect 2195 4441 2196 4445
rect 2200 4441 2201 4445
rect 2205 4441 2206 4445
rect 2210 4441 2211 4445
rect 2215 4441 2216 4445
rect 2220 4441 2221 4445
rect 2225 4441 2226 4445
rect 2186 4440 2230 4441
rect 2190 4436 2191 4440
rect 2195 4436 2196 4440
rect 2200 4436 2201 4440
rect 2205 4436 2206 4440
rect 2210 4436 2211 4440
rect 2215 4436 2216 4440
rect 2220 4436 2221 4440
rect 2225 4436 2226 4440
rect 2186 4435 2230 4436
rect 2190 4431 2191 4435
rect 2195 4431 2196 4435
rect 2200 4431 2201 4435
rect 2205 4431 2206 4435
rect 2210 4431 2211 4435
rect 2215 4431 2216 4435
rect 2220 4431 2221 4435
rect 2225 4431 2226 4435
rect 2186 4430 2230 4431
rect 2190 4426 2191 4430
rect 2195 4426 2196 4430
rect 2200 4426 2201 4430
rect 2205 4426 2206 4430
rect 2210 4426 2211 4430
rect 2215 4426 2216 4430
rect 2220 4426 2221 4430
rect 2225 4426 2226 4430
rect 2186 4425 2230 4426
rect 2190 4421 2191 4425
rect 2195 4421 2196 4425
rect 2200 4421 2201 4425
rect 2205 4421 2206 4425
rect 2210 4421 2211 4425
rect 2215 4421 2216 4425
rect 2220 4421 2221 4425
rect 2225 4421 2226 4425
rect 2186 4420 2230 4421
rect 2190 4416 2191 4420
rect 2195 4416 2196 4420
rect 2200 4416 2201 4420
rect 2205 4416 2206 4420
rect 2210 4416 2211 4420
rect 2215 4416 2216 4420
rect 2220 4416 2221 4420
rect 2225 4416 2226 4420
rect 2186 4415 2230 4416
rect 2190 4411 2191 4415
rect 2195 4411 2196 4415
rect 2200 4411 2201 4415
rect 2205 4411 2206 4415
rect 2210 4411 2211 4415
rect 2215 4411 2216 4415
rect 2220 4411 2221 4415
rect 2225 4411 2226 4415
rect 2186 4410 2230 4411
rect 2190 4406 2191 4410
rect 2195 4406 2196 4410
rect 2200 4406 2201 4410
rect 2205 4406 2206 4410
rect 2210 4406 2211 4410
rect 2215 4406 2216 4410
rect 2220 4406 2221 4410
rect 2225 4406 2226 4410
rect 2186 4405 2230 4406
rect 2190 4401 2191 4405
rect 2195 4401 2196 4405
rect 2200 4401 2201 4405
rect 2205 4401 2206 4405
rect 2210 4401 2211 4405
rect 2215 4401 2216 4405
rect 2220 4401 2221 4405
rect 2225 4401 2226 4405
rect 2186 4400 2230 4401
rect 2190 4396 2191 4400
rect 2195 4396 2196 4400
rect 2200 4396 2201 4400
rect 2205 4396 2206 4400
rect 2210 4396 2211 4400
rect 2215 4396 2216 4400
rect 2220 4396 2221 4400
rect 2225 4396 2226 4400
rect 2186 4395 2230 4396
rect 2190 4391 2191 4395
rect 2195 4391 2196 4395
rect 2200 4391 2201 4395
rect 2205 4391 2206 4395
rect 2210 4391 2211 4395
rect 2215 4391 2216 4395
rect 2220 4391 2221 4395
rect 2225 4391 2226 4395
rect 2186 4390 2230 4391
rect 2190 4386 2191 4390
rect 2195 4386 2196 4390
rect 2200 4386 2201 4390
rect 2205 4386 2206 4390
rect 2210 4386 2211 4390
rect 2215 4386 2216 4390
rect 2220 4386 2221 4390
rect 2225 4386 2226 4390
rect 2186 4385 2230 4386
rect 2190 4381 2191 4385
rect 2195 4381 2196 4385
rect 2200 4381 2201 4385
rect 2205 4381 2206 4385
rect 2210 4381 2211 4385
rect 2215 4381 2216 4385
rect 2220 4381 2221 4385
rect 2225 4381 2226 4385
rect 2186 4380 2230 4381
rect 2190 4376 2191 4380
rect 2195 4376 2196 4380
rect 2200 4376 2201 4380
rect 2205 4376 2206 4380
rect 2210 4376 2211 4380
rect 2215 4376 2216 4380
rect 2220 4376 2221 4380
rect 2225 4376 2226 4380
rect 2186 4375 2230 4376
rect 2190 4371 2191 4375
rect 2195 4371 2196 4375
rect 2200 4371 2201 4375
rect 2205 4371 2206 4375
rect 2210 4371 2211 4375
rect 2215 4371 2216 4375
rect 2220 4371 2221 4375
rect 2225 4371 2226 4375
rect 2186 4370 2230 4371
rect 2190 4366 2191 4370
rect 2195 4366 2196 4370
rect 2200 4366 2201 4370
rect 2205 4366 2206 4370
rect 2210 4366 2211 4370
rect 2215 4366 2216 4370
rect 2220 4366 2221 4370
rect 2225 4366 2226 4370
rect 2186 4365 2230 4366
rect 2190 4361 2191 4365
rect 2195 4361 2196 4365
rect 2200 4361 2201 4365
rect 2205 4361 2206 4365
rect 2210 4361 2211 4365
rect 2215 4361 2216 4365
rect 2220 4361 2221 4365
rect 2225 4361 2226 4365
rect 2238 4445 2242 4446
rect 2238 4440 2242 4441
rect 2238 4435 2242 4436
rect 2238 4430 2242 4431
rect 2238 4425 2242 4426
rect 2238 4420 2242 4421
rect 2238 4415 2242 4416
rect 2238 4410 2242 4411
rect 2238 4405 2242 4406
rect 2238 4400 2242 4401
rect 2238 4395 2242 4396
rect 2238 4390 2242 4391
rect 2238 4385 2242 4386
rect 2238 4380 2242 4381
rect 2238 4375 2242 4376
rect 2238 4370 2242 4371
rect 2238 4365 2242 4366
rect 2174 4360 2178 4361
rect 2174 4353 2178 4356
rect 2238 4360 2242 4361
rect 2238 4353 2242 4356
rect 2178 4349 2181 4353
rect 2185 4349 2186 4353
rect 2190 4349 2191 4353
rect 2195 4349 2196 4353
rect 2200 4349 2201 4353
rect 2205 4349 2206 4353
rect 2210 4349 2211 4353
rect 2215 4349 2216 4353
rect 2220 4349 2221 4353
rect 2225 4349 2226 4353
rect 2230 4349 2231 4353
rect 2235 4349 2238 4353
rect 2251 4465 2255 4466
rect 2251 4460 2255 4461
rect 2251 4455 2255 4456
rect 2251 4450 2255 4451
rect 2251 4445 2255 4446
rect 2251 4440 2255 4441
rect 2251 4435 2255 4436
rect 2251 4430 2255 4431
rect 2251 4425 2255 4426
rect 2251 4420 2255 4421
rect 2251 4415 2255 4416
rect 2251 4410 2255 4411
rect 2251 4405 2255 4406
rect 2251 4400 2255 4401
rect 2251 4395 2255 4396
rect 2251 4390 2255 4391
rect 2251 4385 2255 4386
rect 2251 4380 2255 4381
rect 2251 4375 2255 4376
rect 2251 4370 2255 4371
rect 2251 4365 2255 4366
rect 2251 4360 2255 4361
rect 2251 4355 2255 4356
rect 2251 4350 2255 4351
rect 2161 4345 2165 4346
rect 2161 4340 2165 4341
rect 2251 4345 2255 4346
rect 2251 4340 2255 4341
rect 2165 4336 2166 4340
rect 2170 4336 2171 4340
rect 2175 4336 2176 4340
rect 2180 4336 2181 4340
rect 2185 4336 2186 4340
rect 2190 4336 2191 4340
rect 2195 4336 2196 4340
rect 2200 4336 2201 4340
rect 2205 4336 2206 4340
rect 2210 4336 2211 4340
rect 2215 4336 2216 4340
rect 2220 4336 2221 4340
rect 2225 4336 2226 4340
rect 2230 4336 2231 4340
rect 2235 4336 2236 4340
rect 2240 4336 2241 4340
rect 2245 4336 2246 4340
rect 2250 4336 2251 4340
rect 2314 4471 2315 4475
rect 2319 4471 2320 4475
rect 2324 4471 2325 4475
rect 2329 4471 2330 4475
rect 2334 4471 2335 4475
rect 2339 4471 2340 4475
rect 2344 4471 2345 4475
rect 2349 4471 2350 4475
rect 2354 4471 2355 4475
rect 2359 4471 2360 4475
rect 2364 4471 2365 4475
rect 2369 4471 2370 4475
rect 2374 4471 2375 4475
rect 2379 4471 2380 4475
rect 2384 4471 2385 4475
rect 2389 4471 2390 4475
rect 2394 4471 2395 4475
rect 2399 4471 2400 4475
rect 2433 4472 2442 4483
rect 2505 4475 2561 4483
rect 2620 4503 2676 4515
rect 2728 4514 2751 4523
rect 2814 4519 2872 4523
rect 2876 4519 2877 4523
rect 2881 4519 2882 4523
rect 2811 4518 2882 4519
rect 2811 4515 2872 4518
rect 2728 4511 2732 4514
rect 2725 4507 2732 4511
rect 2744 4511 2751 4514
rect 2814 4514 2872 4515
rect 2876 4514 2877 4518
rect 2881 4514 2882 4518
rect 2814 4512 2882 4514
rect 2929 4535 2985 4592
rect 2929 4531 2994 4535
rect 2929 4519 2985 4531
rect 3046 4527 3059 4717
rect 3220 4624 3221 4628
rect 3225 4624 3226 4628
rect 3230 4624 3231 4628
rect 3216 4623 3235 4624
rect 3220 4619 3221 4623
rect 3225 4619 3226 4623
rect 3230 4619 3231 4623
rect 3216 4618 3235 4619
rect 3220 4614 3221 4618
rect 3225 4614 3226 4618
rect 3230 4614 3231 4618
rect 3216 4613 3235 4614
rect 3220 4609 3221 4613
rect 3225 4609 3226 4613
rect 3230 4609 3231 4613
rect 3216 4608 3235 4609
rect 3220 4604 3221 4608
rect 3225 4604 3226 4608
rect 3230 4604 3231 4608
rect 3216 4603 3235 4604
rect 3220 4599 3221 4603
rect 3225 4599 3226 4603
rect 3230 4599 3231 4603
rect 3216 4598 3235 4599
rect 3220 4594 3221 4598
rect 3225 4594 3226 4598
rect 3230 4594 3231 4598
rect 3238 4601 3294 4602
rect 3238 4597 3240 4601
rect 3244 4597 3245 4601
rect 3249 4597 3250 4601
rect 3254 4597 3255 4601
rect 3259 4597 3260 4601
rect 3264 4597 3265 4601
rect 3269 4597 3270 4601
rect 3274 4597 3275 4601
rect 3279 4597 3280 4601
rect 3284 4597 3285 4601
rect 3289 4597 3290 4601
rect 3238 4596 3294 4597
rect 3238 4592 3240 4596
rect 3244 4592 3245 4596
rect 3249 4592 3250 4596
rect 3254 4592 3255 4596
rect 3259 4592 3260 4596
rect 3264 4592 3265 4596
rect 3269 4592 3270 4596
rect 3274 4592 3275 4596
rect 3279 4592 3280 4596
rect 3284 4592 3285 4596
rect 3289 4592 3290 4596
rect 3123 4578 3191 4580
rect 3123 4574 3181 4578
rect 3185 4574 3186 4578
rect 3190 4574 3191 4578
rect 3123 4573 3191 4574
rect 3123 4569 3181 4573
rect 3185 4569 3186 4573
rect 3190 4569 3191 4573
rect 3123 4568 3191 4569
rect 3123 4564 3181 4568
rect 3185 4564 3186 4568
rect 3190 4564 3191 4568
rect 3123 4563 3191 4564
rect 3123 4559 3181 4563
rect 3185 4559 3186 4563
rect 3190 4559 3191 4563
rect 3123 4558 3191 4559
rect 3123 4554 3181 4558
rect 3185 4554 3186 4558
rect 3190 4554 3191 4558
rect 3123 4553 3191 4554
rect 3123 4549 3181 4553
rect 3185 4549 3186 4553
rect 3190 4549 3191 4553
rect 3123 4548 3191 4549
rect 3220 4578 3221 4582
rect 3225 4578 3226 4582
rect 3230 4578 3231 4582
rect 3216 4577 3235 4578
rect 3220 4573 3221 4577
rect 3225 4573 3226 4577
rect 3230 4573 3231 4577
rect 3216 4572 3235 4573
rect 3220 4568 3221 4572
rect 3225 4568 3226 4572
rect 3230 4568 3231 4572
rect 3216 4567 3235 4568
rect 3220 4563 3221 4567
rect 3225 4563 3226 4567
rect 3230 4563 3231 4567
rect 3216 4562 3235 4563
rect 3220 4558 3221 4562
rect 3225 4558 3226 4562
rect 3230 4558 3231 4562
rect 3216 4557 3235 4558
rect 3220 4553 3221 4557
rect 3225 4553 3226 4557
rect 3230 4553 3231 4557
rect 3216 4552 3235 4553
rect 3220 4548 3221 4552
rect 3225 4548 3226 4552
rect 3230 4548 3231 4552
rect 3123 4544 3181 4548
rect 3185 4544 3186 4548
rect 3190 4544 3191 4548
rect 3123 4543 3191 4544
rect 3123 4539 3181 4543
rect 3185 4539 3186 4543
rect 3190 4539 3191 4543
rect 3123 4538 3191 4539
rect 3123 4535 3181 4538
rect 3120 4534 3181 4535
rect 3185 4534 3186 4538
rect 3190 4534 3191 4538
rect 3120 4533 3191 4534
rect 3120 4531 3181 4533
rect 3123 4529 3181 4531
rect 3185 4529 3186 4533
rect 3190 4529 3191 4533
rect 3123 4528 3191 4529
rect 3034 4523 3064 4527
rect 3123 4524 3181 4528
rect 3185 4524 3186 4528
rect 3190 4524 3191 4528
rect 3123 4523 3191 4524
rect 2929 4515 2994 4519
rect 2744 4507 2755 4511
rect 2620 4499 2685 4503
rect 2814 4503 2870 4512
rect 2620 4487 2676 4499
rect 2737 4495 2741 4502
rect 2811 4499 2870 4503
rect 2725 4491 2755 4495
rect 2814 4487 2870 4499
rect 2620 4483 2685 4487
rect 2811 4483 2870 4487
rect 2620 4475 2676 4483
rect 2310 4470 2314 4471
rect 2400 4470 2404 4471
rect 2431 4470 2444 4472
rect 2474 4471 2475 4475
rect 2479 4471 2480 4475
rect 2484 4471 2485 4475
rect 2489 4471 2490 4475
rect 2494 4471 2495 4475
rect 2499 4471 2500 4475
rect 2504 4471 2505 4475
rect 2509 4471 2510 4475
rect 2514 4471 2515 4475
rect 2519 4471 2520 4475
rect 2524 4471 2525 4475
rect 2529 4471 2530 4475
rect 2534 4471 2535 4475
rect 2539 4471 2540 4475
rect 2544 4471 2545 4475
rect 2549 4471 2550 4475
rect 2554 4471 2555 4475
rect 2559 4471 2560 4475
rect 2470 4470 2474 4471
rect 2429 4468 2446 4470
rect 2310 4465 2314 4466
rect 2310 4460 2314 4461
rect 2310 4455 2314 4456
rect 2310 4450 2314 4451
rect 2310 4445 2314 4446
rect 2310 4440 2314 4441
rect 2310 4435 2314 4436
rect 2310 4430 2314 4431
rect 2310 4425 2314 4426
rect 2310 4420 2314 4421
rect 2310 4415 2314 4416
rect 2310 4410 2314 4411
rect 2310 4405 2314 4406
rect 2310 4400 2314 4401
rect 2310 4395 2314 4396
rect 2310 4390 2314 4391
rect 2310 4385 2314 4386
rect 2310 4380 2314 4381
rect 2310 4375 2314 4376
rect 2310 4370 2314 4371
rect 2310 4365 2314 4366
rect 2310 4360 2314 4361
rect 2310 4355 2314 4356
rect 2310 4350 2314 4351
rect 2327 4458 2330 4466
rect 2334 4458 2335 4466
rect 2339 4458 2340 4466
rect 2344 4458 2345 4466
rect 2349 4458 2350 4466
rect 2354 4458 2355 4466
rect 2359 4458 2360 4466
rect 2364 4458 2365 4466
rect 2369 4458 2370 4466
rect 2374 4458 2375 4466
rect 2379 4458 2380 4466
rect 2384 4458 2387 4466
rect 2323 4455 2327 4458
rect 2323 4450 2327 4451
rect 2387 4455 2391 4458
rect 2387 4450 2391 4451
rect 2323 4445 2327 4446
rect 2323 4440 2327 4441
rect 2323 4435 2327 4436
rect 2323 4430 2327 4431
rect 2323 4425 2327 4426
rect 2323 4420 2327 4421
rect 2323 4415 2327 4416
rect 2323 4410 2327 4411
rect 2323 4405 2327 4406
rect 2323 4400 2327 4401
rect 2323 4395 2327 4396
rect 2323 4390 2327 4391
rect 2323 4385 2327 4386
rect 2323 4380 2327 4381
rect 2323 4375 2327 4376
rect 2323 4370 2327 4371
rect 2323 4365 2327 4366
rect 2339 4446 2340 4450
rect 2344 4446 2345 4450
rect 2349 4446 2350 4450
rect 2354 4446 2355 4450
rect 2359 4446 2360 4450
rect 2364 4446 2365 4450
rect 2369 4446 2370 4450
rect 2374 4446 2375 4450
rect 2379 4446 2380 4450
rect 2335 4445 2380 4446
rect 2339 4441 2340 4445
rect 2344 4441 2345 4445
rect 2349 4441 2350 4445
rect 2354 4441 2355 4445
rect 2359 4441 2360 4445
rect 2364 4441 2365 4445
rect 2369 4441 2370 4445
rect 2374 4441 2375 4445
rect 2379 4441 2380 4445
rect 2335 4440 2380 4441
rect 2339 4436 2340 4440
rect 2344 4436 2345 4440
rect 2349 4436 2350 4440
rect 2354 4436 2355 4440
rect 2359 4436 2360 4440
rect 2364 4436 2365 4440
rect 2369 4436 2370 4440
rect 2374 4436 2375 4440
rect 2379 4436 2380 4440
rect 2335 4435 2380 4436
rect 2339 4431 2340 4435
rect 2344 4431 2345 4435
rect 2349 4431 2350 4435
rect 2354 4431 2355 4435
rect 2359 4431 2360 4435
rect 2364 4431 2365 4435
rect 2369 4431 2370 4435
rect 2374 4431 2375 4435
rect 2379 4431 2380 4435
rect 2335 4430 2380 4431
rect 2339 4426 2340 4430
rect 2344 4426 2345 4430
rect 2349 4426 2350 4430
rect 2354 4426 2355 4430
rect 2359 4426 2360 4430
rect 2364 4426 2365 4430
rect 2369 4426 2370 4430
rect 2374 4426 2375 4430
rect 2379 4426 2380 4430
rect 2335 4425 2380 4426
rect 2339 4421 2340 4425
rect 2344 4421 2345 4425
rect 2349 4421 2350 4425
rect 2354 4421 2355 4425
rect 2359 4421 2360 4425
rect 2364 4421 2365 4425
rect 2369 4421 2370 4425
rect 2374 4421 2375 4425
rect 2379 4421 2380 4425
rect 2335 4420 2380 4421
rect 2339 4416 2340 4420
rect 2344 4416 2345 4420
rect 2349 4416 2350 4420
rect 2354 4416 2355 4420
rect 2359 4416 2360 4420
rect 2364 4416 2365 4420
rect 2369 4416 2370 4420
rect 2374 4416 2375 4420
rect 2379 4416 2380 4420
rect 2335 4415 2380 4416
rect 2339 4411 2340 4415
rect 2344 4411 2345 4415
rect 2349 4411 2350 4415
rect 2354 4411 2355 4415
rect 2359 4411 2360 4415
rect 2364 4411 2365 4415
rect 2369 4411 2370 4415
rect 2374 4411 2375 4415
rect 2379 4411 2380 4415
rect 2335 4410 2380 4411
rect 2339 4406 2340 4410
rect 2344 4406 2345 4410
rect 2349 4406 2350 4410
rect 2354 4406 2355 4410
rect 2359 4406 2360 4410
rect 2364 4406 2365 4410
rect 2369 4406 2370 4410
rect 2374 4406 2375 4410
rect 2379 4406 2380 4410
rect 2335 4405 2380 4406
rect 2339 4401 2340 4405
rect 2344 4401 2345 4405
rect 2349 4401 2350 4405
rect 2354 4401 2355 4405
rect 2359 4401 2360 4405
rect 2364 4401 2365 4405
rect 2369 4401 2370 4405
rect 2374 4401 2375 4405
rect 2379 4401 2380 4405
rect 2335 4400 2380 4401
rect 2339 4396 2340 4400
rect 2344 4396 2345 4400
rect 2349 4396 2350 4400
rect 2354 4396 2355 4400
rect 2359 4396 2360 4400
rect 2364 4396 2365 4400
rect 2369 4396 2370 4400
rect 2374 4396 2375 4400
rect 2379 4396 2380 4400
rect 2335 4395 2380 4396
rect 2339 4391 2340 4395
rect 2344 4391 2345 4395
rect 2349 4391 2350 4395
rect 2354 4391 2355 4395
rect 2359 4391 2360 4395
rect 2364 4391 2365 4395
rect 2369 4391 2370 4395
rect 2374 4391 2375 4395
rect 2379 4391 2380 4395
rect 2335 4390 2380 4391
rect 2339 4386 2340 4390
rect 2344 4386 2345 4390
rect 2349 4386 2350 4390
rect 2354 4386 2355 4390
rect 2359 4386 2360 4390
rect 2364 4386 2365 4390
rect 2369 4386 2370 4390
rect 2374 4386 2375 4390
rect 2379 4386 2380 4390
rect 2335 4385 2380 4386
rect 2339 4381 2340 4385
rect 2344 4381 2345 4385
rect 2349 4381 2350 4385
rect 2354 4381 2355 4385
rect 2359 4381 2360 4385
rect 2364 4381 2365 4385
rect 2369 4381 2370 4385
rect 2374 4381 2375 4385
rect 2379 4381 2380 4385
rect 2335 4380 2380 4381
rect 2339 4376 2340 4380
rect 2344 4376 2345 4380
rect 2349 4376 2350 4380
rect 2354 4376 2355 4380
rect 2359 4376 2360 4380
rect 2364 4376 2365 4380
rect 2369 4376 2370 4380
rect 2374 4376 2375 4380
rect 2379 4376 2380 4380
rect 2335 4375 2380 4376
rect 2339 4371 2340 4375
rect 2344 4371 2345 4375
rect 2349 4371 2350 4375
rect 2354 4371 2355 4375
rect 2359 4371 2360 4375
rect 2364 4371 2365 4375
rect 2369 4371 2370 4375
rect 2374 4371 2375 4375
rect 2379 4371 2380 4375
rect 2335 4370 2380 4371
rect 2339 4366 2340 4370
rect 2344 4366 2345 4370
rect 2349 4366 2350 4370
rect 2354 4366 2355 4370
rect 2359 4366 2360 4370
rect 2364 4366 2365 4370
rect 2369 4366 2370 4370
rect 2374 4366 2375 4370
rect 2379 4366 2380 4370
rect 2335 4365 2380 4366
rect 2339 4361 2340 4365
rect 2344 4361 2345 4365
rect 2349 4361 2350 4365
rect 2354 4361 2355 4365
rect 2359 4361 2360 4365
rect 2364 4361 2365 4365
rect 2369 4361 2370 4365
rect 2374 4361 2375 4365
rect 2379 4361 2380 4365
rect 2387 4445 2391 4446
rect 2387 4440 2391 4441
rect 2387 4435 2391 4436
rect 2387 4430 2391 4431
rect 2387 4425 2391 4426
rect 2387 4420 2391 4421
rect 2387 4415 2391 4416
rect 2387 4410 2391 4411
rect 2387 4405 2391 4406
rect 2387 4400 2391 4401
rect 2387 4395 2391 4396
rect 2387 4390 2391 4391
rect 2387 4385 2391 4386
rect 2387 4380 2391 4381
rect 2387 4375 2391 4376
rect 2387 4370 2391 4371
rect 2387 4365 2391 4366
rect 2323 4360 2327 4361
rect 2323 4353 2327 4356
rect 2387 4360 2391 4361
rect 2387 4353 2391 4356
rect 2327 4349 2330 4353
rect 2334 4349 2335 4353
rect 2339 4349 2340 4353
rect 2344 4349 2345 4353
rect 2349 4349 2350 4353
rect 2354 4349 2355 4353
rect 2359 4349 2360 4353
rect 2364 4349 2365 4353
rect 2369 4349 2370 4353
rect 2374 4349 2375 4353
rect 2379 4349 2380 4353
rect 2384 4349 2387 4353
rect 2400 4465 2404 4466
rect 2400 4460 2404 4461
rect 2400 4455 2404 4456
rect 2400 4450 2404 4451
rect 2400 4445 2404 4446
rect 2400 4440 2404 4441
rect 2400 4435 2404 4436
rect 2427 4440 2448 4468
rect 2560 4470 2564 4471
rect 2470 4465 2474 4466
rect 2470 4460 2474 4461
rect 2470 4455 2474 4456
rect 2470 4450 2474 4451
rect 2470 4445 2474 4446
rect 2470 4440 2474 4441
rect 2470 4435 2474 4436
rect 2400 4430 2404 4431
rect 2400 4425 2404 4426
rect 2400 4420 2404 4421
rect 2400 4415 2404 4416
rect 2400 4410 2404 4411
rect 2400 4405 2404 4406
rect 2400 4400 2404 4401
rect 2400 4395 2404 4396
rect 2400 4390 2404 4391
rect 2400 4385 2404 4386
rect 2400 4380 2404 4381
rect 2400 4375 2404 4376
rect 2400 4370 2404 4371
rect 2400 4365 2404 4366
rect 2470 4430 2474 4431
rect 2470 4425 2474 4426
rect 2470 4420 2474 4421
rect 2470 4415 2474 4416
rect 2470 4410 2474 4411
rect 2470 4405 2474 4406
rect 2470 4400 2474 4401
rect 2470 4395 2474 4396
rect 2470 4390 2474 4391
rect 2470 4385 2474 4386
rect 2470 4380 2474 4381
rect 2470 4375 2474 4376
rect 2470 4370 2474 4371
rect 2470 4365 2474 4366
rect 2400 4360 2404 4361
rect 2400 4355 2404 4356
rect 2400 4350 2404 4351
rect 2310 4345 2314 4346
rect 2310 4340 2314 4341
rect 2400 4345 2404 4346
rect 2400 4340 2404 4341
rect 2314 4336 2315 4340
rect 2319 4336 2320 4340
rect 2324 4336 2325 4340
rect 2329 4336 2330 4340
rect 2334 4336 2335 4340
rect 2339 4336 2340 4340
rect 2344 4336 2345 4340
rect 2349 4336 2350 4340
rect 2354 4336 2355 4340
rect 2359 4336 2360 4340
rect 2364 4336 2365 4340
rect 2369 4336 2370 4340
rect 2374 4336 2375 4340
rect 2379 4336 2380 4340
rect 2384 4336 2385 4340
rect 2389 4336 2390 4340
rect 2394 4336 2395 4340
rect 2399 4336 2400 4340
rect 2427 4333 2448 4353
rect 2470 4360 2474 4361
rect 2470 4355 2474 4356
rect 2470 4350 2474 4351
rect 2487 4458 2490 4466
rect 2494 4458 2495 4466
rect 2499 4458 2500 4466
rect 2504 4458 2505 4466
rect 2509 4458 2510 4466
rect 2514 4458 2515 4466
rect 2519 4458 2520 4466
rect 2524 4458 2525 4466
rect 2529 4458 2530 4466
rect 2534 4458 2535 4466
rect 2539 4458 2540 4466
rect 2544 4458 2547 4466
rect 2483 4455 2487 4458
rect 2483 4450 2487 4451
rect 2547 4455 2551 4458
rect 2547 4450 2551 4451
rect 2483 4445 2487 4446
rect 2483 4440 2487 4441
rect 2483 4435 2487 4436
rect 2483 4430 2487 4431
rect 2483 4425 2487 4426
rect 2483 4420 2487 4421
rect 2483 4415 2487 4416
rect 2483 4410 2487 4411
rect 2483 4405 2487 4406
rect 2483 4400 2487 4401
rect 2483 4395 2487 4396
rect 2483 4390 2487 4391
rect 2483 4385 2487 4386
rect 2483 4380 2487 4381
rect 2483 4375 2487 4376
rect 2483 4370 2487 4371
rect 2483 4365 2487 4366
rect 2499 4446 2500 4450
rect 2504 4446 2505 4450
rect 2509 4446 2510 4450
rect 2514 4446 2515 4450
rect 2519 4446 2520 4450
rect 2524 4446 2525 4450
rect 2529 4446 2530 4450
rect 2534 4446 2535 4450
rect 2495 4445 2539 4446
rect 2499 4441 2500 4445
rect 2504 4441 2505 4445
rect 2509 4441 2510 4445
rect 2514 4441 2515 4445
rect 2519 4441 2520 4445
rect 2524 4441 2525 4445
rect 2529 4441 2530 4445
rect 2534 4441 2535 4445
rect 2495 4440 2539 4441
rect 2499 4436 2500 4440
rect 2504 4436 2505 4440
rect 2509 4436 2510 4440
rect 2514 4436 2515 4440
rect 2519 4436 2520 4440
rect 2524 4436 2525 4440
rect 2529 4436 2530 4440
rect 2534 4436 2535 4440
rect 2495 4435 2539 4436
rect 2499 4431 2500 4435
rect 2504 4431 2505 4435
rect 2509 4431 2510 4435
rect 2514 4431 2515 4435
rect 2519 4431 2520 4435
rect 2524 4431 2525 4435
rect 2529 4431 2530 4435
rect 2534 4431 2535 4435
rect 2495 4430 2539 4431
rect 2499 4426 2500 4430
rect 2504 4426 2505 4430
rect 2509 4426 2510 4430
rect 2514 4426 2515 4430
rect 2519 4426 2520 4430
rect 2524 4426 2525 4430
rect 2529 4426 2530 4430
rect 2534 4426 2535 4430
rect 2495 4425 2539 4426
rect 2499 4421 2500 4425
rect 2504 4421 2505 4425
rect 2509 4421 2510 4425
rect 2514 4421 2515 4425
rect 2519 4421 2520 4425
rect 2524 4421 2525 4425
rect 2529 4421 2530 4425
rect 2534 4421 2535 4425
rect 2495 4420 2539 4421
rect 2499 4416 2500 4420
rect 2504 4416 2505 4420
rect 2509 4416 2510 4420
rect 2514 4416 2515 4420
rect 2519 4416 2520 4420
rect 2524 4416 2525 4420
rect 2529 4416 2530 4420
rect 2534 4416 2535 4420
rect 2495 4415 2539 4416
rect 2499 4411 2500 4415
rect 2504 4411 2505 4415
rect 2509 4411 2510 4415
rect 2514 4411 2515 4415
rect 2519 4411 2520 4415
rect 2524 4411 2525 4415
rect 2529 4411 2530 4415
rect 2534 4411 2535 4415
rect 2495 4410 2539 4411
rect 2499 4406 2500 4410
rect 2504 4406 2505 4410
rect 2509 4406 2510 4410
rect 2514 4406 2515 4410
rect 2519 4406 2520 4410
rect 2524 4406 2525 4410
rect 2529 4406 2530 4410
rect 2534 4406 2535 4410
rect 2495 4405 2539 4406
rect 2499 4401 2500 4405
rect 2504 4401 2505 4405
rect 2509 4401 2510 4405
rect 2514 4401 2515 4405
rect 2519 4401 2520 4405
rect 2524 4401 2525 4405
rect 2529 4401 2530 4405
rect 2534 4401 2535 4405
rect 2495 4400 2539 4401
rect 2499 4396 2500 4400
rect 2504 4396 2505 4400
rect 2509 4396 2510 4400
rect 2514 4396 2515 4400
rect 2519 4396 2520 4400
rect 2524 4396 2525 4400
rect 2529 4396 2530 4400
rect 2534 4396 2535 4400
rect 2495 4395 2539 4396
rect 2499 4391 2500 4395
rect 2504 4391 2505 4395
rect 2509 4391 2510 4395
rect 2514 4391 2515 4395
rect 2519 4391 2520 4395
rect 2524 4391 2525 4395
rect 2529 4391 2530 4395
rect 2534 4391 2535 4395
rect 2495 4390 2539 4391
rect 2499 4386 2500 4390
rect 2504 4386 2505 4390
rect 2509 4386 2510 4390
rect 2514 4386 2515 4390
rect 2519 4386 2520 4390
rect 2524 4386 2525 4390
rect 2529 4386 2530 4390
rect 2534 4386 2535 4390
rect 2495 4385 2539 4386
rect 2499 4381 2500 4385
rect 2504 4381 2505 4385
rect 2509 4381 2510 4385
rect 2514 4381 2515 4385
rect 2519 4381 2520 4385
rect 2524 4381 2525 4385
rect 2529 4381 2530 4385
rect 2534 4381 2535 4385
rect 2495 4380 2539 4381
rect 2499 4376 2500 4380
rect 2504 4376 2505 4380
rect 2509 4376 2510 4380
rect 2514 4376 2515 4380
rect 2519 4376 2520 4380
rect 2524 4376 2525 4380
rect 2529 4376 2530 4380
rect 2534 4376 2535 4380
rect 2495 4375 2539 4376
rect 2499 4371 2500 4375
rect 2504 4371 2505 4375
rect 2509 4371 2510 4375
rect 2514 4371 2515 4375
rect 2519 4371 2520 4375
rect 2524 4371 2525 4375
rect 2529 4371 2530 4375
rect 2534 4371 2535 4375
rect 2495 4370 2539 4371
rect 2499 4366 2500 4370
rect 2504 4366 2505 4370
rect 2509 4366 2510 4370
rect 2514 4366 2515 4370
rect 2519 4366 2520 4370
rect 2524 4366 2525 4370
rect 2529 4366 2530 4370
rect 2534 4366 2535 4370
rect 2495 4365 2539 4366
rect 2499 4361 2500 4365
rect 2504 4361 2505 4365
rect 2509 4361 2510 4365
rect 2514 4361 2515 4365
rect 2519 4361 2520 4365
rect 2524 4361 2525 4365
rect 2529 4361 2530 4365
rect 2534 4361 2535 4365
rect 2547 4445 2551 4446
rect 2547 4440 2551 4441
rect 2547 4435 2551 4436
rect 2547 4430 2551 4431
rect 2547 4425 2551 4426
rect 2547 4420 2551 4421
rect 2547 4415 2551 4416
rect 2547 4410 2551 4411
rect 2547 4405 2551 4406
rect 2547 4400 2551 4401
rect 2547 4395 2551 4396
rect 2547 4390 2551 4391
rect 2547 4385 2551 4386
rect 2547 4380 2551 4381
rect 2547 4375 2551 4376
rect 2547 4370 2551 4371
rect 2547 4365 2551 4366
rect 2483 4360 2487 4361
rect 2483 4353 2487 4356
rect 2547 4360 2551 4361
rect 2547 4353 2551 4356
rect 2487 4349 2490 4353
rect 2494 4349 2495 4353
rect 2499 4349 2500 4353
rect 2504 4349 2505 4353
rect 2509 4349 2510 4353
rect 2514 4349 2515 4353
rect 2519 4349 2520 4353
rect 2524 4349 2525 4353
rect 2529 4349 2530 4353
rect 2534 4349 2535 4353
rect 2539 4349 2540 4353
rect 2544 4349 2547 4353
rect 2560 4465 2564 4466
rect 2560 4460 2564 4461
rect 2560 4455 2564 4456
rect 2560 4450 2564 4451
rect 2560 4445 2564 4446
rect 2560 4440 2564 4441
rect 2560 4435 2564 4436
rect 2560 4430 2564 4431
rect 2560 4425 2564 4426
rect 2560 4420 2564 4421
rect 2560 4415 2564 4416
rect 2560 4410 2564 4411
rect 2560 4405 2564 4406
rect 2560 4400 2564 4401
rect 2560 4395 2564 4396
rect 2560 4390 2564 4391
rect 2560 4385 2564 4386
rect 2560 4380 2564 4381
rect 2560 4375 2564 4376
rect 2560 4370 2564 4371
rect 2560 4365 2564 4366
rect 2560 4360 2564 4361
rect 2560 4355 2564 4356
rect 2560 4350 2564 4351
rect 2470 4345 2474 4346
rect 2470 4340 2474 4341
rect 2560 4345 2564 4346
rect 2560 4340 2564 4341
rect 2474 4336 2475 4340
rect 2479 4336 2480 4340
rect 2484 4336 2485 4340
rect 2489 4336 2490 4340
rect 2494 4336 2495 4340
rect 2499 4336 2500 4340
rect 2504 4336 2505 4340
rect 2509 4336 2510 4340
rect 2514 4336 2515 4340
rect 2519 4336 2520 4340
rect 2524 4336 2525 4340
rect 2529 4336 2530 4340
rect 2534 4336 2535 4340
rect 2539 4336 2540 4340
rect 2544 4336 2545 4340
rect 2549 4336 2550 4340
rect 2554 4336 2555 4340
rect 2559 4336 2560 4340
rect 2623 4471 2624 4475
rect 2628 4471 2629 4475
rect 2633 4471 2634 4475
rect 2638 4471 2639 4475
rect 2643 4471 2644 4475
rect 2648 4471 2649 4475
rect 2653 4471 2654 4475
rect 2658 4471 2659 4475
rect 2663 4471 2664 4475
rect 2668 4471 2669 4475
rect 2673 4471 2674 4475
rect 2678 4471 2679 4475
rect 2683 4471 2684 4475
rect 2688 4471 2689 4475
rect 2693 4471 2694 4475
rect 2698 4471 2699 4475
rect 2703 4471 2704 4475
rect 2708 4471 2709 4475
rect 2742 4472 2751 4483
rect 2814 4475 2870 4483
rect 2929 4503 2985 4515
rect 3037 4514 3060 4523
rect 3123 4519 3181 4523
rect 3185 4519 3186 4523
rect 3190 4519 3191 4523
rect 3120 4518 3191 4519
rect 3120 4515 3181 4518
rect 3037 4511 3041 4514
rect 3034 4507 3041 4511
rect 3053 4511 3060 4514
rect 3123 4514 3181 4515
rect 3185 4514 3186 4518
rect 3190 4514 3191 4518
rect 3123 4512 3191 4514
rect 3238 4535 3294 4592
rect 3238 4531 3303 4535
rect 3238 4519 3294 4531
rect 3355 4527 3368 4721
rect 4483 4718 4484 4722
rect 4488 4718 4489 4722
rect 4493 4718 4494 4722
rect 4498 4718 4499 4722
rect 4503 4718 4504 4722
rect 4508 4718 4509 4722
rect 4529 4733 4530 4737
rect 4534 4733 4535 4737
rect 4539 4733 4540 4737
rect 4544 4733 4545 4737
rect 4549 4733 4550 4737
rect 4554 4733 4555 4737
rect 4525 4732 4559 4733
rect 4529 4728 4530 4732
rect 4534 4728 4535 4732
rect 4539 4728 4540 4732
rect 4544 4728 4545 4732
rect 4549 4728 4550 4732
rect 4554 4728 4555 4732
rect 4525 4727 4559 4728
rect 4529 4723 4530 4727
rect 4534 4723 4535 4727
rect 4539 4723 4540 4727
rect 4544 4723 4545 4727
rect 4549 4723 4550 4727
rect 4554 4723 4555 4727
rect 4525 4722 4559 4723
rect 4529 4718 4530 4722
rect 4534 4718 4535 4722
rect 4539 4718 4540 4722
rect 4544 4718 4545 4722
rect 4549 4718 4550 4722
rect 4554 4718 4555 4722
rect 4483 4707 4484 4711
rect 4488 4707 4489 4711
rect 4493 4707 4494 4711
rect 4498 4707 4499 4711
rect 4503 4707 4504 4711
rect 4508 4707 4509 4711
rect 4479 4706 4513 4707
rect 3647 4653 3699 4704
rect 3647 4649 3664 4653
rect 3668 4649 3669 4653
rect 3673 4649 3699 4653
rect 3647 4648 3699 4649
rect 3647 4644 3664 4648
rect 3668 4644 3669 4648
rect 3673 4644 3699 4648
rect 3647 4643 3699 4644
rect 3647 4639 3664 4643
rect 3668 4639 3669 4643
rect 3673 4639 3699 4643
rect 3647 4638 3699 4639
rect 3647 4634 3664 4638
rect 3668 4634 3669 4638
rect 3673 4634 3699 4638
rect 3647 4633 3699 4634
rect 3647 4629 3664 4633
rect 3668 4629 3669 4633
rect 3673 4629 3699 4633
rect 3647 4628 3699 4629
rect 3529 4624 3530 4628
rect 3534 4624 3535 4628
rect 3539 4624 3540 4628
rect 3525 4623 3544 4624
rect 3529 4619 3530 4623
rect 3534 4619 3535 4623
rect 3539 4619 3540 4623
rect 3525 4618 3544 4619
rect 3529 4614 3530 4618
rect 3534 4614 3535 4618
rect 3539 4614 3540 4618
rect 3525 4613 3544 4614
rect 3529 4609 3530 4613
rect 3534 4609 3535 4613
rect 3539 4609 3540 4613
rect 3525 4608 3544 4609
rect 3529 4604 3530 4608
rect 3534 4604 3535 4608
rect 3539 4604 3540 4608
rect 3525 4603 3544 4604
rect 3529 4599 3530 4603
rect 3534 4599 3535 4603
rect 3539 4599 3540 4603
rect 3647 4624 3664 4628
rect 3668 4624 3669 4628
rect 3673 4624 3699 4628
rect 3647 4623 3699 4624
rect 3647 4619 3664 4623
rect 3668 4619 3669 4623
rect 3673 4619 3699 4623
rect 3647 4618 3699 4619
rect 3647 4614 3664 4618
rect 3668 4614 3669 4618
rect 3673 4614 3699 4618
rect 3647 4613 3699 4614
rect 3647 4609 3664 4613
rect 3668 4609 3669 4613
rect 3673 4609 3699 4613
rect 3647 4608 3699 4609
rect 3647 4604 3664 4608
rect 3668 4604 3669 4608
rect 3673 4604 3699 4608
rect 3647 4603 3699 4604
rect 3525 4598 3544 4599
rect 3529 4594 3530 4598
rect 3534 4594 3535 4598
rect 3539 4594 3540 4598
rect 3547 4601 3603 4602
rect 3547 4597 3549 4601
rect 3553 4597 3554 4601
rect 3558 4597 3559 4601
rect 3563 4597 3564 4601
rect 3568 4597 3569 4601
rect 3573 4597 3574 4601
rect 3578 4597 3579 4601
rect 3583 4597 3584 4601
rect 3588 4597 3589 4601
rect 3593 4597 3594 4601
rect 3598 4597 3599 4601
rect 3547 4596 3603 4597
rect 3547 4592 3549 4596
rect 3553 4592 3554 4596
rect 3558 4592 3559 4596
rect 3563 4592 3564 4596
rect 3568 4592 3569 4596
rect 3573 4592 3574 4596
rect 3578 4592 3579 4596
rect 3583 4592 3584 4596
rect 3588 4592 3589 4596
rect 3593 4592 3594 4596
rect 3598 4592 3599 4596
rect 3432 4578 3500 4580
rect 3432 4574 3490 4578
rect 3494 4574 3495 4578
rect 3499 4574 3500 4578
rect 3432 4573 3500 4574
rect 3432 4569 3490 4573
rect 3494 4569 3495 4573
rect 3499 4569 3500 4573
rect 3432 4568 3500 4569
rect 3432 4564 3490 4568
rect 3494 4564 3495 4568
rect 3499 4564 3500 4568
rect 3432 4563 3500 4564
rect 3432 4559 3490 4563
rect 3494 4559 3495 4563
rect 3499 4559 3500 4563
rect 3432 4558 3500 4559
rect 3432 4554 3490 4558
rect 3494 4554 3495 4558
rect 3499 4554 3500 4558
rect 3432 4553 3500 4554
rect 3432 4549 3490 4553
rect 3494 4549 3495 4553
rect 3499 4549 3500 4553
rect 3432 4548 3500 4549
rect 3529 4578 3530 4582
rect 3534 4578 3535 4582
rect 3539 4578 3540 4582
rect 3525 4577 3544 4578
rect 3529 4573 3530 4577
rect 3534 4573 3535 4577
rect 3539 4573 3540 4577
rect 3525 4572 3544 4573
rect 3529 4568 3530 4572
rect 3534 4568 3535 4572
rect 3539 4568 3540 4572
rect 3525 4567 3544 4568
rect 3529 4563 3530 4567
rect 3534 4563 3535 4567
rect 3539 4563 3540 4567
rect 3525 4562 3544 4563
rect 3529 4558 3530 4562
rect 3534 4558 3535 4562
rect 3539 4558 3540 4562
rect 3525 4557 3544 4558
rect 3529 4553 3530 4557
rect 3534 4553 3535 4557
rect 3539 4553 3540 4557
rect 3525 4552 3544 4553
rect 3529 4548 3530 4552
rect 3534 4548 3535 4552
rect 3539 4548 3540 4552
rect 3432 4544 3490 4548
rect 3494 4544 3495 4548
rect 3499 4544 3500 4548
rect 3432 4543 3500 4544
rect 3432 4539 3490 4543
rect 3494 4539 3495 4543
rect 3499 4539 3500 4543
rect 3432 4538 3500 4539
rect 3432 4535 3490 4538
rect 3429 4534 3490 4535
rect 3494 4534 3495 4538
rect 3499 4534 3500 4538
rect 3429 4533 3500 4534
rect 3429 4531 3490 4533
rect 3432 4529 3490 4531
rect 3494 4529 3495 4533
rect 3499 4529 3500 4533
rect 3432 4528 3500 4529
rect 3343 4523 3373 4527
rect 3432 4524 3490 4528
rect 3494 4524 3495 4528
rect 3499 4524 3500 4528
rect 3432 4523 3500 4524
rect 3238 4515 3303 4519
rect 3053 4507 3064 4511
rect 2929 4499 2994 4503
rect 3123 4503 3179 4512
rect 2929 4487 2985 4499
rect 3046 4495 3050 4502
rect 3120 4499 3179 4503
rect 3034 4491 3064 4495
rect 3123 4487 3179 4499
rect 2929 4483 2994 4487
rect 3120 4483 3179 4487
rect 2929 4475 2985 4483
rect 2619 4470 2623 4471
rect 2709 4470 2713 4471
rect 2740 4470 2753 4472
rect 2783 4471 2784 4475
rect 2788 4471 2789 4475
rect 2793 4471 2794 4475
rect 2798 4471 2799 4475
rect 2803 4471 2804 4475
rect 2808 4471 2809 4475
rect 2813 4471 2814 4475
rect 2818 4471 2819 4475
rect 2823 4471 2824 4475
rect 2828 4471 2829 4475
rect 2833 4471 2834 4475
rect 2838 4471 2839 4475
rect 2843 4471 2844 4475
rect 2848 4471 2849 4475
rect 2853 4471 2854 4475
rect 2858 4471 2859 4475
rect 2863 4471 2864 4475
rect 2868 4471 2869 4475
rect 2779 4470 2783 4471
rect 2738 4468 2755 4470
rect 2619 4465 2623 4466
rect 2619 4460 2623 4461
rect 2619 4455 2623 4456
rect 2619 4450 2623 4451
rect 2619 4445 2623 4446
rect 2619 4440 2623 4441
rect 2619 4435 2623 4436
rect 2619 4430 2623 4431
rect 2619 4425 2623 4426
rect 2619 4420 2623 4421
rect 2619 4415 2623 4416
rect 2619 4410 2623 4411
rect 2619 4405 2623 4406
rect 2619 4400 2623 4401
rect 2619 4395 2623 4396
rect 2619 4390 2623 4391
rect 2619 4385 2623 4386
rect 2619 4380 2623 4381
rect 2619 4375 2623 4376
rect 2619 4370 2623 4371
rect 2619 4365 2623 4366
rect 2619 4360 2623 4361
rect 2619 4355 2623 4356
rect 2619 4350 2623 4351
rect 2636 4458 2639 4466
rect 2643 4458 2644 4466
rect 2648 4458 2649 4466
rect 2653 4458 2654 4466
rect 2658 4458 2659 4466
rect 2663 4458 2664 4466
rect 2668 4458 2669 4466
rect 2673 4458 2674 4466
rect 2678 4458 2679 4466
rect 2683 4458 2684 4466
rect 2688 4458 2689 4466
rect 2693 4458 2696 4466
rect 2632 4455 2636 4458
rect 2632 4450 2636 4451
rect 2696 4455 2700 4458
rect 2696 4450 2700 4451
rect 2632 4445 2636 4446
rect 2632 4440 2636 4441
rect 2632 4435 2636 4436
rect 2632 4430 2636 4431
rect 2632 4425 2636 4426
rect 2632 4420 2636 4421
rect 2632 4415 2636 4416
rect 2632 4410 2636 4411
rect 2632 4405 2636 4406
rect 2632 4400 2636 4401
rect 2632 4395 2636 4396
rect 2632 4390 2636 4391
rect 2632 4385 2636 4386
rect 2632 4380 2636 4381
rect 2632 4375 2636 4376
rect 2632 4370 2636 4371
rect 2632 4365 2636 4366
rect 2648 4446 2649 4450
rect 2653 4446 2654 4450
rect 2658 4446 2659 4450
rect 2663 4446 2664 4450
rect 2668 4446 2669 4450
rect 2673 4446 2674 4450
rect 2678 4446 2679 4450
rect 2683 4446 2684 4450
rect 2688 4446 2689 4450
rect 2644 4445 2689 4446
rect 2648 4441 2649 4445
rect 2653 4441 2654 4445
rect 2658 4441 2659 4445
rect 2663 4441 2664 4445
rect 2668 4441 2669 4445
rect 2673 4441 2674 4445
rect 2678 4441 2679 4445
rect 2683 4441 2684 4445
rect 2688 4441 2689 4445
rect 2644 4440 2689 4441
rect 2648 4436 2649 4440
rect 2653 4436 2654 4440
rect 2658 4436 2659 4440
rect 2663 4436 2664 4440
rect 2668 4436 2669 4440
rect 2673 4436 2674 4440
rect 2678 4436 2679 4440
rect 2683 4436 2684 4440
rect 2688 4436 2689 4440
rect 2644 4435 2689 4436
rect 2648 4431 2649 4435
rect 2653 4431 2654 4435
rect 2658 4431 2659 4435
rect 2663 4431 2664 4435
rect 2668 4431 2669 4435
rect 2673 4431 2674 4435
rect 2678 4431 2679 4435
rect 2683 4431 2684 4435
rect 2688 4431 2689 4435
rect 2644 4430 2689 4431
rect 2648 4426 2649 4430
rect 2653 4426 2654 4430
rect 2658 4426 2659 4430
rect 2663 4426 2664 4430
rect 2668 4426 2669 4430
rect 2673 4426 2674 4430
rect 2678 4426 2679 4430
rect 2683 4426 2684 4430
rect 2688 4426 2689 4430
rect 2644 4425 2689 4426
rect 2648 4421 2649 4425
rect 2653 4421 2654 4425
rect 2658 4421 2659 4425
rect 2663 4421 2664 4425
rect 2668 4421 2669 4425
rect 2673 4421 2674 4425
rect 2678 4421 2679 4425
rect 2683 4421 2684 4425
rect 2688 4421 2689 4425
rect 2644 4420 2689 4421
rect 2648 4416 2649 4420
rect 2653 4416 2654 4420
rect 2658 4416 2659 4420
rect 2663 4416 2664 4420
rect 2668 4416 2669 4420
rect 2673 4416 2674 4420
rect 2678 4416 2679 4420
rect 2683 4416 2684 4420
rect 2688 4416 2689 4420
rect 2644 4415 2689 4416
rect 2648 4411 2649 4415
rect 2653 4411 2654 4415
rect 2658 4411 2659 4415
rect 2663 4411 2664 4415
rect 2668 4411 2669 4415
rect 2673 4411 2674 4415
rect 2678 4411 2679 4415
rect 2683 4411 2684 4415
rect 2688 4411 2689 4415
rect 2644 4410 2689 4411
rect 2648 4406 2649 4410
rect 2653 4406 2654 4410
rect 2658 4406 2659 4410
rect 2663 4406 2664 4410
rect 2668 4406 2669 4410
rect 2673 4406 2674 4410
rect 2678 4406 2679 4410
rect 2683 4406 2684 4410
rect 2688 4406 2689 4410
rect 2644 4405 2689 4406
rect 2648 4401 2649 4405
rect 2653 4401 2654 4405
rect 2658 4401 2659 4405
rect 2663 4401 2664 4405
rect 2668 4401 2669 4405
rect 2673 4401 2674 4405
rect 2678 4401 2679 4405
rect 2683 4401 2684 4405
rect 2688 4401 2689 4405
rect 2644 4400 2689 4401
rect 2648 4396 2649 4400
rect 2653 4396 2654 4400
rect 2658 4396 2659 4400
rect 2663 4396 2664 4400
rect 2668 4396 2669 4400
rect 2673 4396 2674 4400
rect 2678 4396 2679 4400
rect 2683 4396 2684 4400
rect 2688 4396 2689 4400
rect 2644 4395 2689 4396
rect 2648 4391 2649 4395
rect 2653 4391 2654 4395
rect 2658 4391 2659 4395
rect 2663 4391 2664 4395
rect 2668 4391 2669 4395
rect 2673 4391 2674 4395
rect 2678 4391 2679 4395
rect 2683 4391 2684 4395
rect 2688 4391 2689 4395
rect 2644 4390 2689 4391
rect 2648 4386 2649 4390
rect 2653 4386 2654 4390
rect 2658 4386 2659 4390
rect 2663 4386 2664 4390
rect 2668 4386 2669 4390
rect 2673 4386 2674 4390
rect 2678 4386 2679 4390
rect 2683 4386 2684 4390
rect 2688 4386 2689 4390
rect 2644 4385 2689 4386
rect 2648 4381 2649 4385
rect 2653 4381 2654 4385
rect 2658 4381 2659 4385
rect 2663 4381 2664 4385
rect 2668 4381 2669 4385
rect 2673 4381 2674 4385
rect 2678 4381 2679 4385
rect 2683 4381 2684 4385
rect 2688 4381 2689 4385
rect 2644 4380 2689 4381
rect 2648 4376 2649 4380
rect 2653 4376 2654 4380
rect 2658 4376 2659 4380
rect 2663 4376 2664 4380
rect 2668 4376 2669 4380
rect 2673 4376 2674 4380
rect 2678 4376 2679 4380
rect 2683 4376 2684 4380
rect 2688 4376 2689 4380
rect 2644 4375 2689 4376
rect 2648 4371 2649 4375
rect 2653 4371 2654 4375
rect 2658 4371 2659 4375
rect 2663 4371 2664 4375
rect 2668 4371 2669 4375
rect 2673 4371 2674 4375
rect 2678 4371 2679 4375
rect 2683 4371 2684 4375
rect 2688 4371 2689 4375
rect 2644 4370 2689 4371
rect 2648 4366 2649 4370
rect 2653 4366 2654 4370
rect 2658 4366 2659 4370
rect 2663 4366 2664 4370
rect 2668 4366 2669 4370
rect 2673 4366 2674 4370
rect 2678 4366 2679 4370
rect 2683 4366 2684 4370
rect 2688 4366 2689 4370
rect 2644 4365 2689 4366
rect 2648 4361 2649 4365
rect 2653 4361 2654 4365
rect 2658 4361 2659 4365
rect 2663 4361 2664 4365
rect 2668 4361 2669 4365
rect 2673 4361 2674 4365
rect 2678 4361 2679 4365
rect 2683 4361 2684 4365
rect 2688 4361 2689 4365
rect 2696 4445 2700 4446
rect 2696 4440 2700 4441
rect 2696 4435 2700 4436
rect 2696 4430 2700 4431
rect 2696 4425 2700 4426
rect 2696 4420 2700 4421
rect 2696 4415 2700 4416
rect 2696 4410 2700 4411
rect 2696 4405 2700 4406
rect 2696 4400 2700 4401
rect 2696 4395 2700 4396
rect 2696 4390 2700 4391
rect 2696 4385 2700 4386
rect 2696 4380 2700 4381
rect 2696 4375 2700 4376
rect 2696 4370 2700 4371
rect 2696 4365 2700 4366
rect 2632 4360 2636 4361
rect 2632 4353 2636 4356
rect 2696 4360 2700 4361
rect 2696 4353 2700 4356
rect 2636 4349 2639 4353
rect 2643 4349 2644 4353
rect 2648 4349 2649 4353
rect 2653 4349 2654 4353
rect 2658 4349 2659 4353
rect 2663 4349 2664 4353
rect 2668 4349 2669 4353
rect 2673 4349 2674 4353
rect 2678 4349 2679 4353
rect 2683 4349 2684 4353
rect 2688 4349 2689 4353
rect 2693 4349 2696 4353
rect 2709 4465 2713 4466
rect 2709 4460 2713 4461
rect 2709 4455 2713 4456
rect 2709 4450 2713 4451
rect 2709 4445 2713 4446
rect 2709 4440 2713 4441
rect 2709 4435 2713 4436
rect 2736 4440 2757 4468
rect 2869 4470 2873 4471
rect 2779 4465 2783 4466
rect 2779 4460 2783 4461
rect 2779 4455 2783 4456
rect 2779 4450 2783 4451
rect 2779 4445 2783 4446
rect 2779 4440 2783 4441
rect 2779 4435 2783 4436
rect 2709 4430 2713 4431
rect 2709 4425 2713 4426
rect 2709 4420 2713 4421
rect 2709 4415 2713 4416
rect 2709 4410 2713 4411
rect 2709 4405 2713 4406
rect 2709 4400 2713 4401
rect 2709 4395 2713 4396
rect 2709 4390 2713 4391
rect 2709 4385 2713 4386
rect 2709 4380 2713 4381
rect 2709 4375 2713 4376
rect 2709 4370 2713 4371
rect 2709 4365 2713 4366
rect 2779 4430 2783 4431
rect 2779 4425 2783 4426
rect 2779 4420 2783 4421
rect 2779 4415 2783 4416
rect 2779 4410 2783 4411
rect 2779 4405 2783 4406
rect 2779 4400 2783 4401
rect 2779 4395 2783 4396
rect 2779 4390 2783 4391
rect 2779 4385 2783 4386
rect 2779 4380 2783 4381
rect 2779 4375 2783 4376
rect 2779 4370 2783 4371
rect 2779 4365 2783 4366
rect 2709 4360 2713 4361
rect 2709 4355 2713 4356
rect 2709 4350 2713 4351
rect 2619 4345 2623 4346
rect 2619 4340 2623 4341
rect 2709 4345 2713 4346
rect 2709 4340 2713 4341
rect 2623 4336 2624 4340
rect 2628 4336 2629 4340
rect 2633 4336 2634 4340
rect 2638 4336 2639 4340
rect 2643 4336 2644 4340
rect 2648 4336 2649 4340
rect 2653 4336 2654 4340
rect 2658 4336 2659 4340
rect 2663 4336 2664 4340
rect 2668 4336 2669 4340
rect 2673 4336 2674 4340
rect 2678 4336 2679 4340
rect 2683 4336 2684 4340
rect 2688 4336 2689 4340
rect 2693 4336 2694 4340
rect 2698 4336 2699 4340
rect 2703 4336 2704 4340
rect 2708 4336 2709 4340
rect 2736 4333 2757 4353
rect 2779 4360 2783 4361
rect 2779 4355 2783 4356
rect 2779 4350 2783 4351
rect 2796 4458 2799 4466
rect 2803 4458 2804 4466
rect 2808 4458 2809 4466
rect 2813 4458 2814 4466
rect 2818 4458 2819 4466
rect 2823 4458 2824 4466
rect 2828 4458 2829 4466
rect 2833 4458 2834 4466
rect 2838 4458 2839 4466
rect 2843 4458 2844 4466
rect 2848 4458 2849 4466
rect 2853 4458 2856 4466
rect 2792 4455 2796 4458
rect 2792 4450 2796 4451
rect 2856 4455 2860 4458
rect 2856 4450 2860 4451
rect 2792 4445 2796 4446
rect 2792 4440 2796 4441
rect 2792 4435 2796 4436
rect 2792 4430 2796 4431
rect 2792 4425 2796 4426
rect 2792 4420 2796 4421
rect 2792 4415 2796 4416
rect 2792 4410 2796 4411
rect 2792 4405 2796 4406
rect 2792 4400 2796 4401
rect 2792 4395 2796 4396
rect 2792 4390 2796 4391
rect 2792 4385 2796 4386
rect 2792 4380 2796 4381
rect 2792 4375 2796 4376
rect 2792 4370 2796 4371
rect 2792 4365 2796 4366
rect 2808 4446 2809 4450
rect 2813 4446 2814 4450
rect 2818 4446 2819 4450
rect 2823 4446 2824 4450
rect 2828 4446 2829 4450
rect 2833 4446 2834 4450
rect 2838 4446 2839 4450
rect 2843 4446 2844 4450
rect 2804 4445 2848 4446
rect 2808 4441 2809 4445
rect 2813 4441 2814 4445
rect 2818 4441 2819 4445
rect 2823 4441 2824 4445
rect 2828 4441 2829 4445
rect 2833 4441 2834 4445
rect 2838 4441 2839 4445
rect 2843 4441 2844 4445
rect 2804 4440 2848 4441
rect 2808 4436 2809 4440
rect 2813 4436 2814 4440
rect 2818 4436 2819 4440
rect 2823 4436 2824 4440
rect 2828 4436 2829 4440
rect 2833 4436 2834 4440
rect 2838 4436 2839 4440
rect 2843 4436 2844 4440
rect 2804 4435 2848 4436
rect 2808 4431 2809 4435
rect 2813 4431 2814 4435
rect 2818 4431 2819 4435
rect 2823 4431 2824 4435
rect 2828 4431 2829 4435
rect 2833 4431 2834 4435
rect 2838 4431 2839 4435
rect 2843 4431 2844 4435
rect 2804 4430 2848 4431
rect 2808 4426 2809 4430
rect 2813 4426 2814 4430
rect 2818 4426 2819 4430
rect 2823 4426 2824 4430
rect 2828 4426 2829 4430
rect 2833 4426 2834 4430
rect 2838 4426 2839 4430
rect 2843 4426 2844 4430
rect 2804 4425 2848 4426
rect 2808 4421 2809 4425
rect 2813 4421 2814 4425
rect 2818 4421 2819 4425
rect 2823 4421 2824 4425
rect 2828 4421 2829 4425
rect 2833 4421 2834 4425
rect 2838 4421 2839 4425
rect 2843 4421 2844 4425
rect 2804 4420 2848 4421
rect 2808 4416 2809 4420
rect 2813 4416 2814 4420
rect 2818 4416 2819 4420
rect 2823 4416 2824 4420
rect 2828 4416 2829 4420
rect 2833 4416 2834 4420
rect 2838 4416 2839 4420
rect 2843 4416 2844 4420
rect 2804 4415 2848 4416
rect 2808 4411 2809 4415
rect 2813 4411 2814 4415
rect 2818 4411 2819 4415
rect 2823 4411 2824 4415
rect 2828 4411 2829 4415
rect 2833 4411 2834 4415
rect 2838 4411 2839 4415
rect 2843 4411 2844 4415
rect 2804 4410 2848 4411
rect 2808 4406 2809 4410
rect 2813 4406 2814 4410
rect 2818 4406 2819 4410
rect 2823 4406 2824 4410
rect 2828 4406 2829 4410
rect 2833 4406 2834 4410
rect 2838 4406 2839 4410
rect 2843 4406 2844 4410
rect 2804 4405 2848 4406
rect 2808 4401 2809 4405
rect 2813 4401 2814 4405
rect 2818 4401 2819 4405
rect 2823 4401 2824 4405
rect 2828 4401 2829 4405
rect 2833 4401 2834 4405
rect 2838 4401 2839 4405
rect 2843 4401 2844 4405
rect 2804 4400 2848 4401
rect 2808 4396 2809 4400
rect 2813 4396 2814 4400
rect 2818 4396 2819 4400
rect 2823 4396 2824 4400
rect 2828 4396 2829 4400
rect 2833 4396 2834 4400
rect 2838 4396 2839 4400
rect 2843 4396 2844 4400
rect 2804 4395 2848 4396
rect 2808 4391 2809 4395
rect 2813 4391 2814 4395
rect 2818 4391 2819 4395
rect 2823 4391 2824 4395
rect 2828 4391 2829 4395
rect 2833 4391 2834 4395
rect 2838 4391 2839 4395
rect 2843 4391 2844 4395
rect 2804 4390 2848 4391
rect 2808 4386 2809 4390
rect 2813 4386 2814 4390
rect 2818 4386 2819 4390
rect 2823 4386 2824 4390
rect 2828 4386 2829 4390
rect 2833 4386 2834 4390
rect 2838 4386 2839 4390
rect 2843 4386 2844 4390
rect 2804 4385 2848 4386
rect 2808 4381 2809 4385
rect 2813 4381 2814 4385
rect 2818 4381 2819 4385
rect 2823 4381 2824 4385
rect 2828 4381 2829 4385
rect 2833 4381 2834 4385
rect 2838 4381 2839 4385
rect 2843 4381 2844 4385
rect 2804 4380 2848 4381
rect 2808 4376 2809 4380
rect 2813 4376 2814 4380
rect 2818 4376 2819 4380
rect 2823 4376 2824 4380
rect 2828 4376 2829 4380
rect 2833 4376 2834 4380
rect 2838 4376 2839 4380
rect 2843 4376 2844 4380
rect 2804 4375 2848 4376
rect 2808 4371 2809 4375
rect 2813 4371 2814 4375
rect 2818 4371 2819 4375
rect 2823 4371 2824 4375
rect 2828 4371 2829 4375
rect 2833 4371 2834 4375
rect 2838 4371 2839 4375
rect 2843 4371 2844 4375
rect 2804 4370 2848 4371
rect 2808 4366 2809 4370
rect 2813 4366 2814 4370
rect 2818 4366 2819 4370
rect 2823 4366 2824 4370
rect 2828 4366 2829 4370
rect 2833 4366 2834 4370
rect 2838 4366 2839 4370
rect 2843 4366 2844 4370
rect 2804 4365 2848 4366
rect 2808 4361 2809 4365
rect 2813 4361 2814 4365
rect 2818 4361 2819 4365
rect 2823 4361 2824 4365
rect 2828 4361 2829 4365
rect 2833 4361 2834 4365
rect 2838 4361 2839 4365
rect 2843 4361 2844 4365
rect 2856 4445 2860 4446
rect 2856 4440 2860 4441
rect 2856 4435 2860 4436
rect 2856 4430 2860 4431
rect 2856 4425 2860 4426
rect 2856 4420 2860 4421
rect 2856 4415 2860 4416
rect 2856 4410 2860 4411
rect 2856 4405 2860 4406
rect 2856 4400 2860 4401
rect 2856 4395 2860 4396
rect 2856 4390 2860 4391
rect 2856 4385 2860 4386
rect 2856 4380 2860 4381
rect 2856 4375 2860 4376
rect 2856 4370 2860 4371
rect 2856 4365 2860 4366
rect 2792 4360 2796 4361
rect 2792 4353 2796 4356
rect 2856 4360 2860 4361
rect 2856 4353 2860 4356
rect 2796 4349 2799 4353
rect 2803 4349 2804 4353
rect 2808 4349 2809 4353
rect 2813 4349 2814 4353
rect 2818 4349 2819 4353
rect 2823 4349 2824 4353
rect 2828 4349 2829 4353
rect 2833 4349 2834 4353
rect 2838 4349 2839 4353
rect 2843 4349 2844 4353
rect 2848 4349 2849 4353
rect 2853 4349 2856 4353
rect 2869 4465 2873 4466
rect 2869 4460 2873 4461
rect 2869 4455 2873 4456
rect 2869 4450 2873 4451
rect 2869 4445 2873 4446
rect 2869 4440 2873 4441
rect 2869 4435 2873 4436
rect 2869 4430 2873 4431
rect 2869 4425 2873 4426
rect 2869 4420 2873 4421
rect 2869 4415 2873 4416
rect 2869 4410 2873 4411
rect 2869 4405 2873 4406
rect 2869 4400 2873 4401
rect 2869 4395 2873 4396
rect 2869 4390 2873 4391
rect 2869 4385 2873 4386
rect 2869 4380 2873 4381
rect 2869 4375 2873 4376
rect 2869 4370 2873 4371
rect 2869 4365 2873 4366
rect 2869 4360 2873 4361
rect 2869 4355 2873 4356
rect 2869 4350 2873 4351
rect 2779 4345 2783 4346
rect 2779 4340 2783 4341
rect 2869 4345 2873 4346
rect 2869 4340 2873 4341
rect 2783 4336 2784 4340
rect 2788 4336 2789 4340
rect 2793 4336 2794 4340
rect 2798 4336 2799 4340
rect 2803 4336 2804 4340
rect 2808 4336 2809 4340
rect 2813 4336 2814 4340
rect 2818 4336 2819 4340
rect 2823 4336 2824 4340
rect 2828 4336 2829 4340
rect 2833 4336 2834 4340
rect 2838 4336 2839 4340
rect 2843 4336 2844 4340
rect 2848 4336 2849 4340
rect 2853 4336 2854 4340
rect 2858 4336 2859 4340
rect 2863 4336 2864 4340
rect 2868 4336 2869 4340
rect 2932 4471 2933 4475
rect 2937 4471 2938 4475
rect 2942 4471 2943 4475
rect 2947 4471 2948 4475
rect 2952 4471 2953 4475
rect 2957 4471 2958 4475
rect 2962 4471 2963 4475
rect 2967 4471 2968 4475
rect 2972 4471 2973 4475
rect 2977 4471 2978 4475
rect 2982 4471 2983 4475
rect 2987 4471 2988 4475
rect 2992 4471 2993 4475
rect 2997 4471 2998 4475
rect 3002 4471 3003 4475
rect 3007 4471 3008 4475
rect 3012 4471 3013 4475
rect 3017 4471 3018 4475
rect 3051 4472 3060 4483
rect 3123 4475 3179 4483
rect 3238 4503 3294 4515
rect 3346 4514 3369 4523
rect 3432 4519 3490 4523
rect 3494 4519 3495 4523
rect 3499 4519 3500 4523
rect 3429 4518 3500 4519
rect 3429 4515 3490 4518
rect 3346 4511 3350 4514
rect 3343 4507 3350 4511
rect 3362 4511 3369 4514
rect 3432 4514 3490 4515
rect 3494 4514 3495 4518
rect 3499 4514 3500 4518
rect 3432 4512 3500 4514
rect 3362 4507 3373 4511
rect 3238 4499 3303 4503
rect 3432 4503 3488 4512
rect 3238 4487 3294 4499
rect 3355 4495 3359 4502
rect 3429 4499 3488 4503
rect 3343 4491 3373 4495
rect 3432 4487 3488 4499
rect 3238 4483 3303 4487
rect 3429 4483 3488 4487
rect 3238 4475 3294 4483
rect 2928 4470 2932 4471
rect 3018 4470 3022 4471
rect 3049 4470 3062 4472
rect 3092 4471 3093 4475
rect 3097 4471 3098 4475
rect 3102 4471 3103 4475
rect 3107 4471 3108 4475
rect 3112 4471 3113 4475
rect 3117 4471 3118 4475
rect 3122 4471 3123 4475
rect 3127 4471 3128 4475
rect 3132 4471 3133 4475
rect 3137 4471 3138 4475
rect 3142 4471 3143 4475
rect 3147 4471 3148 4475
rect 3152 4471 3153 4475
rect 3157 4471 3158 4475
rect 3162 4471 3163 4475
rect 3167 4471 3168 4475
rect 3172 4471 3173 4475
rect 3177 4471 3178 4475
rect 3088 4470 3092 4471
rect 3047 4468 3064 4470
rect 2928 4465 2932 4466
rect 2928 4460 2932 4461
rect 2928 4455 2932 4456
rect 2928 4450 2932 4451
rect 2928 4445 2932 4446
rect 2928 4440 2932 4441
rect 2928 4435 2932 4436
rect 2928 4430 2932 4431
rect 2928 4425 2932 4426
rect 2928 4420 2932 4421
rect 2928 4415 2932 4416
rect 2928 4410 2932 4411
rect 2928 4405 2932 4406
rect 2928 4400 2932 4401
rect 2928 4395 2932 4396
rect 2928 4390 2932 4391
rect 2928 4385 2932 4386
rect 2928 4380 2932 4381
rect 2928 4375 2932 4376
rect 2928 4370 2932 4371
rect 2928 4365 2932 4366
rect 2928 4360 2932 4361
rect 2928 4355 2932 4356
rect 2928 4350 2932 4351
rect 2945 4458 2948 4466
rect 2952 4458 2953 4466
rect 2957 4458 2958 4466
rect 2962 4458 2963 4466
rect 2967 4458 2968 4466
rect 2972 4458 2973 4466
rect 2977 4458 2978 4466
rect 2982 4458 2983 4466
rect 2987 4458 2988 4466
rect 2992 4458 2993 4466
rect 2997 4458 2998 4466
rect 3002 4458 3005 4466
rect 2941 4455 2945 4458
rect 2941 4450 2945 4451
rect 3005 4455 3009 4458
rect 3005 4450 3009 4451
rect 2941 4445 2945 4446
rect 2941 4440 2945 4441
rect 2941 4435 2945 4436
rect 2941 4430 2945 4431
rect 2941 4425 2945 4426
rect 2941 4420 2945 4421
rect 2941 4415 2945 4416
rect 2941 4410 2945 4411
rect 2941 4405 2945 4406
rect 2941 4400 2945 4401
rect 2941 4395 2945 4396
rect 2941 4390 2945 4391
rect 2941 4385 2945 4386
rect 2941 4380 2945 4381
rect 2941 4375 2945 4376
rect 2941 4370 2945 4371
rect 2941 4365 2945 4366
rect 2957 4446 2958 4450
rect 2962 4446 2963 4450
rect 2967 4446 2968 4450
rect 2972 4446 2973 4450
rect 2977 4446 2978 4450
rect 2982 4446 2983 4450
rect 2987 4446 2988 4450
rect 2992 4446 2993 4450
rect 2997 4446 2998 4450
rect 2953 4445 2998 4446
rect 2957 4441 2958 4445
rect 2962 4441 2963 4445
rect 2967 4441 2968 4445
rect 2972 4441 2973 4445
rect 2977 4441 2978 4445
rect 2982 4441 2983 4445
rect 2987 4441 2988 4445
rect 2992 4441 2993 4445
rect 2997 4441 2998 4445
rect 2953 4440 2998 4441
rect 2957 4436 2958 4440
rect 2962 4436 2963 4440
rect 2967 4436 2968 4440
rect 2972 4436 2973 4440
rect 2977 4436 2978 4440
rect 2982 4436 2983 4440
rect 2987 4436 2988 4440
rect 2992 4436 2993 4440
rect 2997 4436 2998 4440
rect 2953 4435 2998 4436
rect 2957 4431 2958 4435
rect 2962 4431 2963 4435
rect 2967 4431 2968 4435
rect 2972 4431 2973 4435
rect 2977 4431 2978 4435
rect 2982 4431 2983 4435
rect 2987 4431 2988 4435
rect 2992 4431 2993 4435
rect 2997 4431 2998 4435
rect 2953 4430 2998 4431
rect 2957 4426 2958 4430
rect 2962 4426 2963 4430
rect 2967 4426 2968 4430
rect 2972 4426 2973 4430
rect 2977 4426 2978 4430
rect 2982 4426 2983 4430
rect 2987 4426 2988 4430
rect 2992 4426 2993 4430
rect 2997 4426 2998 4430
rect 2953 4425 2998 4426
rect 2957 4421 2958 4425
rect 2962 4421 2963 4425
rect 2967 4421 2968 4425
rect 2972 4421 2973 4425
rect 2977 4421 2978 4425
rect 2982 4421 2983 4425
rect 2987 4421 2988 4425
rect 2992 4421 2993 4425
rect 2997 4421 2998 4425
rect 2953 4420 2998 4421
rect 2957 4416 2958 4420
rect 2962 4416 2963 4420
rect 2967 4416 2968 4420
rect 2972 4416 2973 4420
rect 2977 4416 2978 4420
rect 2982 4416 2983 4420
rect 2987 4416 2988 4420
rect 2992 4416 2993 4420
rect 2997 4416 2998 4420
rect 2953 4415 2998 4416
rect 2957 4411 2958 4415
rect 2962 4411 2963 4415
rect 2967 4411 2968 4415
rect 2972 4411 2973 4415
rect 2977 4411 2978 4415
rect 2982 4411 2983 4415
rect 2987 4411 2988 4415
rect 2992 4411 2993 4415
rect 2997 4411 2998 4415
rect 2953 4410 2998 4411
rect 2957 4406 2958 4410
rect 2962 4406 2963 4410
rect 2967 4406 2968 4410
rect 2972 4406 2973 4410
rect 2977 4406 2978 4410
rect 2982 4406 2983 4410
rect 2987 4406 2988 4410
rect 2992 4406 2993 4410
rect 2997 4406 2998 4410
rect 2953 4405 2998 4406
rect 2957 4401 2958 4405
rect 2962 4401 2963 4405
rect 2967 4401 2968 4405
rect 2972 4401 2973 4405
rect 2977 4401 2978 4405
rect 2982 4401 2983 4405
rect 2987 4401 2988 4405
rect 2992 4401 2993 4405
rect 2997 4401 2998 4405
rect 2953 4400 2998 4401
rect 2957 4396 2958 4400
rect 2962 4396 2963 4400
rect 2967 4396 2968 4400
rect 2972 4396 2973 4400
rect 2977 4396 2978 4400
rect 2982 4396 2983 4400
rect 2987 4396 2988 4400
rect 2992 4396 2993 4400
rect 2997 4396 2998 4400
rect 2953 4395 2998 4396
rect 2957 4391 2958 4395
rect 2962 4391 2963 4395
rect 2967 4391 2968 4395
rect 2972 4391 2973 4395
rect 2977 4391 2978 4395
rect 2982 4391 2983 4395
rect 2987 4391 2988 4395
rect 2992 4391 2993 4395
rect 2997 4391 2998 4395
rect 2953 4390 2998 4391
rect 2957 4386 2958 4390
rect 2962 4386 2963 4390
rect 2967 4386 2968 4390
rect 2972 4386 2973 4390
rect 2977 4386 2978 4390
rect 2982 4386 2983 4390
rect 2987 4386 2988 4390
rect 2992 4386 2993 4390
rect 2997 4386 2998 4390
rect 2953 4385 2998 4386
rect 2957 4381 2958 4385
rect 2962 4381 2963 4385
rect 2967 4381 2968 4385
rect 2972 4381 2973 4385
rect 2977 4381 2978 4385
rect 2982 4381 2983 4385
rect 2987 4381 2988 4385
rect 2992 4381 2993 4385
rect 2997 4381 2998 4385
rect 2953 4380 2998 4381
rect 2957 4376 2958 4380
rect 2962 4376 2963 4380
rect 2967 4376 2968 4380
rect 2972 4376 2973 4380
rect 2977 4376 2978 4380
rect 2982 4376 2983 4380
rect 2987 4376 2988 4380
rect 2992 4376 2993 4380
rect 2997 4376 2998 4380
rect 2953 4375 2998 4376
rect 2957 4371 2958 4375
rect 2962 4371 2963 4375
rect 2967 4371 2968 4375
rect 2972 4371 2973 4375
rect 2977 4371 2978 4375
rect 2982 4371 2983 4375
rect 2987 4371 2988 4375
rect 2992 4371 2993 4375
rect 2997 4371 2998 4375
rect 2953 4370 2998 4371
rect 2957 4366 2958 4370
rect 2962 4366 2963 4370
rect 2967 4366 2968 4370
rect 2972 4366 2973 4370
rect 2977 4366 2978 4370
rect 2982 4366 2983 4370
rect 2987 4366 2988 4370
rect 2992 4366 2993 4370
rect 2997 4366 2998 4370
rect 2953 4365 2998 4366
rect 2957 4361 2958 4365
rect 2962 4361 2963 4365
rect 2967 4361 2968 4365
rect 2972 4361 2973 4365
rect 2977 4361 2978 4365
rect 2982 4361 2983 4365
rect 2987 4361 2988 4365
rect 2992 4361 2993 4365
rect 2997 4361 2998 4365
rect 3005 4445 3009 4446
rect 3005 4440 3009 4441
rect 3005 4435 3009 4436
rect 3005 4430 3009 4431
rect 3005 4425 3009 4426
rect 3005 4420 3009 4421
rect 3005 4415 3009 4416
rect 3005 4410 3009 4411
rect 3005 4405 3009 4406
rect 3005 4400 3009 4401
rect 3005 4395 3009 4396
rect 3005 4390 3009 4391
rect 3005 4385 3009 4386
rect 3005 4380 3009 4381
rect 3005 4375 3009 4376
rect 3005 4370 3009 4371
rect 3005 4365 3009 4366
rect 2941 4360 2945 4361
rect 2941 4353 2945 4356
rect 3005 4360 3009 4361
rect 3005 4353 3009 4356
rect 2945 4349 2948 4353
rect 2952 4349 2953 4353
rect 2957 4349 2958 4353
rect 2962 4349 2963 4353
rect 2967 4349 2968 4353
rect 2972 4349 2973 4353
rect 2977 4349 2978 4353
rect 2982 4349 2983 4353
rect 2987 4349 2988 4353
rect 2992 4349 2993 4353
rect 2997 4349 2998 4353
rect 3002 4349 3005 4353
rect 3018 4465 3022 4466
rect 3018 4460 3022 4461
rect 3018 4455 3022 4456
rect 3018 4450 3022 4451
rect 3018 4445 3022 4446
rect 3018 4440 3022 4441
rect 3018 4435 3022 4436
rect 3045 4440 3066 4468
rect 3178 4470 3182 4471
rect 3088 4465 3092 4466
rect 3088 4460 3092 4461
rect 3088 4455 3092 4456
rect 3088 4450 3092 4451
rect 3088 4445 3092 4446
rect 3088 4440 3092 4441
rect 3088 4435 3092 4436
rect 3018 4430 3022 4431
rect 3018 4425 3022 4426
rect 3018 4420 3022 4421
rect 3018 4415 3022 4416
rect 3018 4410 3022 4411
rect 3018 4405 3022 4406
rect 3018 4400 3022 4401
rect 3018 4395 3022 4396
rect 3018 4390 3022 4391
rect 3018 4385 3022 4386
rect 3018 4380 3022 4381
rect 3018 4375 3022 4376
rect 3018 4370 3022 4371
rect 3018 4365 3022 4366
rect 3088 4430 3092 4431
rect 3088 4425 3092 4426
rect 3088 4420 3092 4421
rect 3088 4415 3092 4416
rect 3088 4410 3092 4411
rect 3088 4405 3092 4406
rect 3088 4400 3092 4401
rect 3088 4395 3092 4396
rect 3088 4390 3092 4391
rect 3088 4385 3092 4386
rect 3088 4380 3092 4381
rect 3088 4375 3092 4376
rect 3088 4370 3092 4371
rect 3088 4365 3092 4366
rect 3018 4360 3022 4361
rect 3018 4355 3022 4356
rect 3018 4350 3022 4351
rect 2928 4345 2932 4346
rect 2928 4340 2932 4341
rect 3018 4345 3022 4346
rect 3018 4340 3022 4341
rect 2932 4336 2933 4340
rect 2937 4336 2938 4340
rect 2942 4336 2943 4340
rect 2947 4336 2948 4340
rect 2952 4336 2953 4340
rect 2957 4336 2958 4340
rect 2962 4336 2963 4340
rect 2967 4336 2968 4340
rect 2972 4336 2973 4340
rect 2977 4336 2978 4340
rect 2982 4336 2983 4340
rect 2987 4336 2988 4340
rect 2992 4336 2993 4340
rect 2997 4336 2998 4340
rect 3002 4336 3003 4340
rect 3007 4336 3008 4340
rect 3012 4336 3013 4340
rect 3017 4336 3018 4340
rect 3045 4333 3066 4353
rect 3088 4360 3092 4361
rect 3088 4355 3092 4356
rect 3088 4350 3092 4351
rect 3105 4458 3108 4466
rect 3112 4458 3113 4466
rect 3117 4458 3118 4466
rect 3122 4458 3123 4466
rect 3127 4458 3128 4466
rect 3132 4458 3133 4466
rect 3137 4458 3138 4466
rect 3142 4458 3143 4466
rect 3147 4458 3148 4466
rect 3152 4458 3153 4466
rect 3157 4458 3158 4466
rect 3162 4458 3165 4466
rect 3101 4455 3105 4458
rect 3101 4450 3105 4451
rect 3165 4455 3169 4458
rect 3165 4450 3169 4451
rect 3101 4445 3105 4446
rect 3101 4440 3105 4441
rect 3101 4435 3105 4436
rect 3101 4430 3105 4431
rect 3101 4425 3105 4426
rect 3101 4420 3105 4421
rect 3101 4415 3105 4416
rect 3101 4410 3105 4411
rect 3101 4405 3105 4406
rect 3101 4400 3105 4401
rect 3101 4395 3105 4396
rect 3101 4390 3105 4391
rect 3101 4385 3105 4386
rect 3101 4380 3105 4381
rect 3101 4375 3105 4376
rect 3101 4370 3105 4371
rect 3101 4365 3105 4366
rect 3117 4446 3118 4450
rect 3122 4446 3123 4450
rect 3127 4446 3128 4450
rect 3132 4446 3133 4450
rect 3137 4446 3138 4450
rect 3142 4446 3143 4450
rect 3147 4446 3148 4450
rect 3152 4446 3153 4450
rect 3113 4445 3157 4446
rect 3117 4441 3118 4445
rect 3122 4441 3123 4445
rect 3127 4441 3128 4445
rect 3132 4441 3133 4445
rect 3137 4441 3138 4445
rect 3142 4441 3143 4445
rect 3147 4441 3148 4445
rect 3152 4441 3153 4445
rect 3113 4440 3157 4441
rect 3117 4436 3118 4440
rect 3122 4436 3123 4440
rect 3127 4436 3128 4440
rect 3132 4436 3133 4440
rect 3137 4436 3138 4440
rect 3142 4436 3143 4440
rect 3147 4436 3148 4440
rect 3152 4436 3153 4440
rect 3113 4435 3157 4436
rect 3117 4431 3118 4435
rect 3122 4431 3123 4435
rect 3127 4431 3128 4435
rect 3132 4431 3133 4435
rect 3137 4431 3138 4435
rect 3142 4431 3143 4435
rect 3147 4431 3148 4435
rect 3152 4431 3153 4435
rect 3113 4430 3157 4431
rect 3117 4426 3118 4430
rect 3122 4426 3123 4430
rect 3127 4426 3128 4430
rect 3132 4426 3133 4430
rect 3137 4426 3138 4430
rect 3142 4426 3143 4430
rect 3147 4426 3148 4430
rect 3152 4426 3153 4430
rect 3113 4425 3157 4426
rect 3117 4421 3118 4425
rect 3122 4421 3123 4425
rect 3127 4421 3128 4425
rect 3132 4421 3133 4425
rect 3137 4421 3138 4425
rect 3142 4421 3143 4425
rect 3147 4421 3148 4425
rect 3152 4421 3153 4425
rect 3113 4420 3157 4421
rect 3117 4416 3118 4420
rect 3122 4416 3123 4420
rect 3127 4416 3128 4420
rect 3132 4416 3133 4420
rect 3137 4416 3138 4420
rect 3142 4416 3143 4420
rect 3147 4416 3148 4420
rect 3152 4416 3153 4420
rect 3113 4415 3157 4416
rect 3117 4411 3118 4415
rect 3122 4411 3123 4415
rect 3127 4411 3128 4415
rect 3132 4411 3133 4415
rect 3137 4411 3138 4415
rect 3142 4411 3143 4415
rect 3147 4411 3148 4415
rect 3152 4411 3153 4415
rect 3113 4410 3157 4411
rect 3117 4406 3118 4410
rect 3122 4406 3123 4410
rect 3127 4406 3128 4410
rect 3132 4406 3133 4410
rect 3137 4406 3138 4410
rect 3142 4406 3143 4410
rect 3147 4406 3148 4410
rect 3152 4406 3153 4410
rect 3113 4405 3157 4406
rect 3117 4401 3118 4405
rect 3122 4401 3123 4405
rect 3127 4401 3128 4405
rect 3132 4401 3133 4405
rect 3137 4401 3138 4405
rect 3142 4401 3143 4405
rect 3147 4401 3148 4405
rect 3152 4401 3153 4405
rect 3113 4400 3157 4401
rect 3117 4396 3118 4400
rect 3122 4396 3123 4400
rect 3127 4396 3128 4400
rect 3132 4396 3133 4400
rect 3137 4396 3138 4400
rect 3142 4396 3143 4400
rect 3147 4396 3148 4400
rect 3152 4396 3153 4400
rect 3113 4395 3157 4396
rect 3117 4391 3118 4395
rect 3122 4391 3123 4395
rect 3127 4391 3128 4395
rect 3132 4391 3133 4395
rect 3137 4391 3138 4395
rect 3142 4391 3143 4395
rect 3147 4391 3148 4395
rect 3152 4391 3153 4395
rect 3113 4390 3157 4391
rect 3117 4386 3118 4390
rect 3122 4386 3123 4390
rect 3127 4386 3128 4390
rect 3132 4386 3133 4390
rect 3137 4386 3138 4390
rect 3142 4386 3143 4390
rect 3147 4386 3148 4390
rect 3152 4386 3153 4390
rect 3113 4385 3157 4386
rect 3117 4381 3118 4385
rect 3122 4381 3123 4385
rect 3127 4381 3128 4385
rect 3132 4381 3133 4385
rect 3137 4381 3138 4385
rect 3142 4381 3143 4385
rect 3147 4381 3148 4385
rect 3152 4381 3153 4385
rect 3113 4380 3157 4381
rect 3117 4376 3118 4380
rect 3122 4376 3123 4380
rect 3127 4376 3128 4380
rect 3132 4376 3133 4380
rect 3137 4376 3138 4380
rect 3142 4376 3143 4380
rect 3147 4376 3148 4380
rect 3152 4376 3153 4380
rect 3113 4375 3157 4376
rect 3117 4371 3118 4375
rect 3122 4371 3123 4375
rect 3127 4371 3128 4375
rect 3132 4371 3133 4375
rect 3137 4371 3138 4375
rect 3142 4371 3143 4375
rect 3147 4371 3148 4375
rect 3152 4371 3153 4375
rect 3113 4370 3157 4371
rect 3117 4366 3118 4370
rect 3122 4366 3123 4370
rect 3127 4366 3128 4370
rect 3132 4366 3133 4370
rect 3137 4366 3138 4370
rect 3142 4366 3143 4370
rect 3147 4366 3148 4370
rect 3152 4366 3153 4370
rect 3113 4365 3157 4366
rect 3117 4361 3118 4365
rect 3122 4361 3123 4365
rect 3127 4361 3128 4365
rect 3132 4361 3133 4365
rect 3137 4361 3138 4365
rect 3142 4361 3143 4365
rect 3147 4361 3148 4365
rect 3152 4361 3153 4365
rect 3165 4445 3169 4446
rect 3165 4440 3169 4441
rect 3165 4435 3169 4436
rect 3165 4430 3169 4431
rect 3165 4425 3169 4426
rect 3165 4420 3169 4421
rect 3165 4415 3169 4416
rect 3165 4410 3169 4411
rect 3165 4405 3169 4406
rect 3165 4400 3169 4401
rect 3165 4395 3169 4396
rect 3165 4390 3169 4391
rect 3165 4385 3169 4386
rect 3165 4380 3169 4381
rect 3165 4375 3169 4376
rect 3165 4370 3169 4371
rect 3165 4365 3169 4366
rect 3101 4360 3105 4361
rect 3101 4353 3105 4356
rect 3165 4360 3169 4361
rect 3165 4353 3169 4356
rect 3105 4349 3108 4353
rect 3112 4349 3113 4353
rect 3117 4349 3118 4353
rect 3122 4349 3123 4353
rect 3127 4349 3128 4353
rect 3132 4349 3133 4353
rect 3137 4349 3138 4353
rect 3142 4349 3143 4353
rect 3147 4349 3148 4353
rect 3152 4349 3153 4353
rect 3157 4349 3158 4353
rect 3162 4349 3165 4353
rect 3178 4465 3182 4466
rect 3178 4460 3182 4461
rect 3178 4455 3182 4456
rect 3178 4450 3182 4451
rect 3178 4445 3182 4446
rect 3178 4440 3182 4441
rect 3178 4435 3182 4436
rect 3178 4430 3182 4431
rect 3178 4425 3182 4426
rect 3178 4420 3182 4421
rect 3178 4415 3182 4416
rect 3178 4410 3182 4411
rect 3178 4405 3182 4406
rect 3178 4400 3182 4401
rect 3178 4395 3182 4396
rect 3178 4390 3182 4391
rect 3178 4385 3182 4386
rect 3178 4380 3182 4381
rect 3178 4375 3182 4376
rect 3178 4370 3182 4371
rect 3178 4365 3182 4366
rect 3178 4360 3182 4361
rect 3178 4355 3182 4356
rect 3178 4350 3182 4351
rect 3088 4345 3092 4346
rect 3088 4340 3092 4341
rect 3178 4345 3182 4346
rect 3178 4340 3182 4341
rect 3092 4336 3093 4340
rect 3097 4336 3098 4340
rect 3102 4336 3103 4340
rect 3107 4336 3108 4340
rect 3112 4336 3113 4340
rect 3117 4336 3118 4340
rect 3122 4336 3123 4340
rect 3127 4336 3128 4340
rect 3132 4336 3133 4340
rect 3137 4336 3138 4340
rect 3142 4336 3143 4340
rect 3147 4336 3148 4340
rect 3152 4336 3153 4340
rect 3157 4336 3158 4340
rect 3162 4336 3163 4340
rect 3167 4336 3168 4340
rect 3172 4336 3173 4340
rect 3177 4336 3178 4340
rect 3241 4471 3242 4475
rect 3246 4471 3247 4475
rect 3251 4471 3252 4475
rect 3256 4471 3257 4475
rect 3261 4471 3262 4475
rect 3266 4471 3267 4475
rect 3271 4471 3272 4475
rect 3276 4471 3277 4475
rect 3281 4471 3282 4475
rect 3286 4471 3287 4475
rect 3291 4471 3292 4475
rect 3296 4471 3297 4475
rect 3301 4471 3302 4475
rect 3306 4471 3307 4475
rect 3311 4471 3312 4475
rect 3316 4471 3317 4475
rect 3321 4471 3322 4475
rect 3326 4471 3327 4475
rect 3360 4472 3369 4483
rect 3432 4475 3488 4483
rect 3547 4475 3603 4592
rect 3647 4599 3664 4603
rect 3668 4599 3669 4603
rect 3673 4599 3699 4603
rect 3237 4470 3241 4471
rect 3327 4470 3331 4471
rect 3358 4470 3371 4472
rect 3401 4471 3402 4475
rect 3406 4471 3407 4475
rect 3411 4471 3412 4475
rect 3416 4471 3417 4475
rect 3421 4471 3422 4475
rect 3426 4471 3427 4475
rect 3431 4471 3432 4475
rect 3436 4471 3437 4475
rect 3441 4471 3442 4475
rect 3446 4471 3447 4475
rect 3451 4471 3452 4475
rect 3456 4471 3457 4475
rect 3461 4471 3462 4475
rect 3466 4471 3467 4475
rect 3471 4471 3472 4475
rect 3476 4471 3477 4475
rect 3481 4471 3482 4475
rect 3486 4471 3487 4475
rect 3397 4470 3401 4471
rect 3356 4468 3373 4470
rect 3237 4465 3241 4466
rect 3237 4460 3241 4461
rect 3237 4455 3241 4456
rect 3237 4450 3241 4451
rect 3237 4445 3241 4446
rect 3237 4440 3241 4441
rect 3237 4435 3241 4436
rect 3237 4430 3241 4431
rect 3237 4425 3241 4426
rect 3237 4420 3241 4421
rect 3237 4415 3241 4416
rect 3237 4410 3241 4411
rect 3237 4405 3241 4406
rect 3237 4400 3241 4401
rect 3237 4395 3241 4396
rect 3237 4390 3241 4391
rect 3237 4385 3241 4386
rect 3237 4380 3241 4381
rect 3237 4375 3241 4376
rect 3237 4370 3241 4371
rect 3237 4365 3241 4366
rect 3237 4360 3241 4361
rect 3237 4355 3241 4356
rect 3237 4350 3241 4351
rect 3254 4458 3257 4466
rect 3261 4458 3262 4466
rect 3266 4458 3267 4466
rect 3271 4458 3272 4466
rect 3276 4458 3277 4466
rect 3281 4458 3282 4466
rect 3286 4458 3287 4466
rect 3291 4458 3292 4466
rect 3296 4458 3297 4466
rect 3301 4458 3302 4466
rect 3306 4458 3307 4466
rect 3311 4458 3314 4466
rect 3250 4455 3254 4458
rect 3250 4450 3254 4451
rect 3314 4455 3318 4458
rect 3314 4450 3318 4451
rect 3250 4445 3254 4446
rect 3250 4440 3254 4441
rect 3250 4435 3254 4436
rect 3250 4430 3254 4431
rect 3250 4425 3254 4426
rect 3250 4420 3254 4421
rect 3250 4415 3254 4416
rect 3250 4410 3254 4411
rect 3250 4405 3254 4406
rect 3250 4400 3254 4401
rect 3250 4395 3254 4396
rect 3250 4390 3254 4391
rect 3250 4385 3254 4386
rect 3250 4380 3254 4381
rect 3250 4375 3254 4376
rect 3250 4370 3254 4371
rect 3250 4365 3254 4366
rect 3266 4446 3267 4450
rect 3271 4446 3272 4450
rect 3276 4446 3277 4450
rect 3281 4446 3282 4450
rect 3286 4446 3287 4450
rect 3291 4446 3292 4450
rect 3296 4446 3297 4450
rect 3301 4446 3302 4450
rect 3306 4446 3307 4450
rect 3262 4445 3307 4446
rect 3266 4441 3267 4445
rect 3271 4441 3272 4445
rect 3276 4441 3277 4445
rect 3281 4441 3282 4445
rect 3286 4441 3287 4445
rect 3291 4441 3292 4445
rect 3296 4441 3297 4445
rect 3301 4441 3302 4445
rect 3306 4441 3307 4445
rect 3262 4440 3307 4441
rect 3266 4436 3267 4440
rect 3271 4436 3272 4440
rect 3276 4436 3277 4440
rect 3281 4436 3282 4440
rect 3286 4436 3287 4440
rect 3291 4436 3292 4440
rect 3296 4436 3297 4440
rect 3301 4436 3302 4440
rect 3306 4436 3307 4440
rect 3262 4435 3307 4436
rect 3266 4431 3267 4435
rect 3271 4431 3272 4435
rect 3276 4431 3277 4435
rect 3281 4431 3282 4435
rect 3286 4431 3287 4435
rect 3291 4431 3292 4435
rect 3296 4431 3297 4435
rect 3301 4431 3302 4435
rect 3306 4431 3307 4435
rect 3262 4430 3307 4431
rect 3266 4426 3267 4430
rect 3271 4426 3272 4430
rect 3276 4426 3277 4430
rect 3281 4426 3282 4430
rect 3286 4426 3287 4430
rect 3291 4426 3292 4430
rect 3296 4426 3297 4430
rect 3301 4426 3302 4430
rect 3306 4426 3307 4430
rect 3262 4425 3307 4426
rect 3266 4421 3267 4425
rect 3271 4421 3272 4425
rect 3276 4421 3277 4425
rect 3281 4421 3282 4425
rect 3286 4421 3287 4425
rect 3291 4421 3292 4425
rect 3296 4421 3297 4425
rect 3301 4421 3302 4425
rect 3306 4421 3307 4425
rect 3262 4420 3307 4421
rect 3266 4416 3267 4420
rect 3271 4416 3272 4420
rect 3276 4416 3277 4420
rect 3281 4416 3282 4420
rect 3286 4416 3287 4420
rect 3291 4416 3292 4420
rect 3296 4416 3297 4420
rect 3301 4416 3302 4420
rect 3306 4416 3307 4420
rect 3262 4415 3307 4416
rect 3266 4411 3267 4415
rect 3271 4411 3272 4415
rect 3276 4411 3277 4415
rect 3281 4411 3282 4415
rect 3286 4411 3287 4415
rect 3291 4411 3292 4415
rect 3296 4411 3297 4415
rect 3301 4411 3302 4415
rect 3306 4411 3307 4415
rect 3262 4410 3307 4411
rect 3266 4406 3267 4410
rect 3271 4406 3272 4410
rect 3276 4406 3277 4410
rect 3281 4406 3282 4410
rect 3286 4406 3287 4410
rect 3291 4406 3292 4410
rect 3296 4406 3297 4410
rect 3301 4406 3302 4410
rect 3306 4406 3307 4410
rect 3262 4405 3307 4406
rect 3266 4401 3267 4405
rect 3271 4401 3272 4405
rect 3276 4401 3277 4405
rect 3281 4401 3282 4405
rect 3286 4401 3287 4405
rect 3291 4401 3292 4405
rect 3296 4401 3297 4405
rect 3301 4401 3302 4405
rect 3306 4401 3307 4405
rect 3262 4400 3307 4401
rect 3266 4396 3267 4400
rect 3271 4396 3272 4400
rect 3276 4396 3277 4400
rect 3281 4396 3282 4400
rect 3286 4396 3287 4400
rect 3291 4396 3292 4400
rect 3296 4396 3297 4400
rect 3301 4396 3302 4400
rect 3306 4396 3307 4400
rect 3262 4395 3307 4396
rect 3266 4391 3267 4395
rect 3271 4391 3272 4395
rect 3276 4391 3277 4395
rect 3281 4391 3282 4395
rect 3286 4391 3287 4395
rect 3291 4391 3292 4395
rect 3296 4391 3297 4395
rect 3301 4391 3302 4395
rect 3306 4391 3307 4395
rect 3262 4390 3307 4391
rect 3266 4386 3267 4390
rect 3271 4386 3272 4390
rect 3276 4386 3277 4390
rect 3281 4386 3282 4390
rect 3286 4386 3287 4390
rect 3291 4386 3292 4390
rect 3296 4386 3297 4390
rect 3301 4386 3302 4390
rect 3306 4386 3307 4390
rect 3262 4385 3307 4386
rect 3266 4381 3267 4385
rect 3271 4381 3272 4385
rect 3276 4381 3277 4385
rect 3281 4381 3282 4385
rect 3286 4381 3287 4385
rect 3291 4381 3292 4385
rect 3296 4381 3297 4385
rect 3301 4381 3302 4385
rect 3306 4381 3307 4385
rect 3262 4380 3307 4381
rect 3266 4376 3267 4380
rect 3271 4376 3272 4380
rect 3276 4376 3277 4380
rect 3281 4376 3282 4380
rect 3286 4376 3287 4380
rect 3291 4376 3292 4380
rect 3296 4376 3297 4380
rect 3301 4376 3302 4380
rect 3306 4376 3307 4380
rect 3262 4375 3307 4376
rect 3266 4371 3267 4375
rect 3271 4371 3272 4375
rect 3276 4371 3277 4375
rect 3281 4371 3282 4375
rect 3286 4371 3287 4375
rect 3291 4371 3292 4375
rect 3296 4371 3297 4375
rect 3301 4371 3302 4375
rect 3306 4371 3307 4375
rect 3262 4370 3307 4371
rect 3266 4366 3267 4370
rect 3271 4366 3272 4370
rect 3276 4366 3277 4370
rect 3281 4366 3282 4370
rect 3286 4366 3287 4370
rect 3291 4366 3292 4370
rect 3296 4366 3297 4370
rect 3301 4366 3302 4370
rect 3306 4366 3307 4370
rect 3262 4365 3307 4366
rect 3266 4361 3267 4365
rect 3271 4361 3272 4365
rect 3276 4361 3277 4365
rect 3281 4361 3282 4365
rect 3286 4361 3287 4365
rect 3291 4361 3292 4365
rect 3296 4361 3297 4365
rect 3301 4361 3302 4365
rect 3306 4361 3307 4365
rect 3314 4445 3318 4446
rect 3314 4440 3318 4441
rect 3314 4435 3318 4436
rect 3314 4430 3318 4431
rect 3314 4425 3318 4426
rect 3314 4420 3318 4421
rect 3314 4415 3318 4416
rect 3314 4410 3318 4411
rect 3314 4405 3318 4406
rect 3314 4400 3318 4401
rect 3314 4395 3318 4396
rect 3314 4390 3318 4391
rect 3314 4385 3318 4386
rect 3314 4380 3318 4381
rect 3314 4375 3318 4376
rect 3314 4370 3318 4371
rect 3314 4365 3318 4366
rect 3250 4360 3254 4361
rect 3250 4353 3254 4356
rect 3314 4360 3318 4361
rect 3314 4353 3318 4356
rect 3254 4349 3257 4353
rect 3261 4349 3262 4353
rect 3266 4349 3267 4353
rect 3271 4349 3272 4353
rect 3276 4349 3277 4353
rect 3281 4349 3282 4353
rect 3286 4349 3287 4353
rect 3291 4349 3292 4353
rect 3296 4349 3297 4353
rect 3301 4349 3302 4353
rect 3306 4349 3307 4353
rect 3311 4349 3314 4353
rect 3327 4465 3331 4466
rect 3327 4460 3331 4461
rect 3327 4455 3331 4456
rect 3327 4450 3331 4451
rect 3327 4445 3331 4446
rect 3327 4440 3331 4441
rect 3327 4435 3331 4436
rect 3354 4440 3375 4468
rect 3487 4470 3491 4471
rect 3397 4465 3401 4466
rect 3397 4460 3401 4461
rect 3397 4455 3401 4456
rect 3397 4450 3401 4451
rect 3397 4445 3401 4446
rect 3397 4440 3401 4441
rect 3397 4435 3401 4436
rect 3327 4430 3331 4431
rect 3327 4425 3331 4426
rect 3327 4420 3331 4421
rect 3327 4415 3331 4416
rect 3327 4410 3331 4411
rect 3327 4405 3331 4406
rect 3327 4400 3331 4401
rect 3327 4395 3331 4396
rect 3327 4390 3331 4391
rect 3327 4385 3331 4386
rect 3327 4380 3331 4381
rect 3327 4375 3331 4376
rect 3327 4370 3331 4371
rect 3327 4365 3331 4366
rect 3397 4430 3401 4431
rect 3397 4425 3401 4426
rect 3397 4420 3401 4421
rect 3397 4415 3401 4416
rect 3397 4410 3401 4411
rect 3397 4405 3401 4406
rect 3397 4400 3401 4401
rect 3397 4395 3401 4396
rect 3397 4390 3401 4391
rect 3397 4385 3401 4386
rect 3397 4380 3401 4381
rect 3397 4375 3401 4376
rect 3397 4370 3401 4371
rect 3397 4365 3401 4366
rect 3327 4360 3331 4361
rect 3327 4355 3331 4356
rect 3327 4350 3331 4351
rect 3237 4345 3241 4346
rect 3237 4340 3241 4341
rect 3327 4345 3331 4346
rect 3327 4340 3331 4341
rect 3241 4336 3242 4340
rect 3246 4336 3247 4340
rect 3251 4336 3252 4340
rect 3256 4336 3257 4340
rect 3261 4336 3262 4340
rect 3266 4336 3267 4340
rect 3271 4336 3272 4340
rect 3276 4336 3277 4340
rect 3281 4336 3282 4340
rect 3286 4336 3287 4340
rect 3291 4336 3292 4340
rect 3296 4336 3297 4340
rect 3301 4336 3302 4340
rect 3306 4336 3307 4340
rect 3311 4336 3312 4340
rect 3316 4336 3317 4340
rect 3321 4336 3322 4340
rect 3326 4336 3327 4340
rect 3354 4333 3375 4353
rect 3397 4360 3401 4361
rect 3397 4355 3401 4356
rect 3397 4350 3401 4351
rect 3414 4458 3417 4466
rect 3421 4458 3422 4466
rect 3426 4458 3427 4466
rect 3431 4458 3432 4466
rect 3436 4458 3437 4466
rect 3441 4458 3442 4466
rect 3446 4458 3447 4466
rect 3451 4458 3452 4466
rect 3456 4458 3457 4466
rect 3461 4458 3462 4466
rect 3466 4458 3467 4466
rect 3471 4458 3474 4466
rect 3410 4455 3414 4458
rect 3410 4450 3414 4451
rect 3474 4455 3478 4458
rect 3474 4450 3478 4451
rect 3410 4445 3414 4446
rect 3410 4440 3414 4441
rect 3410 4435 3414 4436
rect 3410 4430 3414 4431
rect 3410 4425 3414 4426
rect 3410 4420 3414 4421
rect 3410 4415 3414 4416
rect 3410 4410 3414 4411
rect 3410 4405 3414 4406
rect 3410 4400 3414 4401
rect 3410 4395 3414 4396
rect 3410 4390 3414 4391
rect 3410 4385 3414 4386
rect 3410 4380 3414 4381
rect 3410 4375 3414 4376
rect 3410 4370 3414 4371
rect 3410 4365 3414 4366
rect 3426 4446 3427 4450
rect 3431 4446 3432 4450
rect 3436 4446 3437 4450
rect 3441 4446 3442 4450
rect 3446 4446 3447 4450
rect 3451 4446 3452 4450
rect 3456 4446 3457 4450
rect 3461 4446 3462 4450
rect 3422 4445 3466 4446
rect 3426 4441 3427 4445
rect 3431 4441 3432 4445
rect 3436 4441 3437 4445
rect 3441 4441 3442 4445
rect 3446 4441 3447 4445
rect 3451 4441 3452 4445
rect 3456 4441 3457 4445
rect 3461 4441 3462 4445
rect 3422 4440 3466 4441
rect 3426 4436 3427 4440
rect 3431 4436 3432 4440
rect 3436 4436 3437 4440
rect 3441 4436 3442 4440
rect 3446 4436 3447 4440
rect 3451 4436 3452 4440
rect 3456 4436 3457 4440
rect 3461 4436 3462 4440
rect 3422 4435 3466 4436
rect 3426 4431 3427 4435
rect 3431 4431 3432 4435
rect 3436 4431 3437 4435
rect 3441 4431 3442 4435
rect 3446 4431 3447 4435
rect 3451 4431 3452 4435
rect 3456 4431 3457 4435
rect 3461 4431 3462 4435
rect 3422 4430 3466 4431
rect 3426 4426 3427 4430
rect 3431 4426 3432 4430
rect 3436 4426 3437 4430
rect 3441 4426 3442 4430
rect 3446 4426 3447 4430
rect 3451 4426 3452 4430
rect 3456 4426 3457 4430
rect 3461 4426 3462 4430
rect 3422 4425 3466 4426
rect 3426 4421 3427 4425
rect 3431 4421 3432 4425
rect 3436 4421 3437 4425
rect 3441 4421 3442 4425
rect 3446 4421 3447 4425
rect 3451 4421 3452 4425
rect 3456 4421 3457 4425
rect 3461 4421 3462 4425
rect 3422 4420 3466 4421
rect 3426 4416 3427 4420
rect 3431 4416 3432 4420
rect 3436 4416 3437 4420
rect 3441 4416 3442 4420
rect 3446 4416 3447 4420
rect 3451 4416 3452 4420
rect 3456 4416 3457 4420
rect 3461 4416 3462 4420
rect 3422 4415 3466 4416
rect 3426 4411 3427 4415
rect 3431 4411 3432 4415
rect 3436 4411 3437 4415
rect 3441 4411 3442 4415
rect 3446 4411 3447 4415
rect 3451 4411 3452 4415
rect 3456 4411 3457 4415
rect 3461 4411 3462 4415
rect 3422 4410 3466 4411
rect 3426 4406 3427 4410
rect 3431 4406 3432 4410
rect 3436 4406 3437 4410
rect 3441 4406 3442 4410
rect 3446 4406 3447 4410
rect 3451 4406 3452 4410
rect 3456 4406 3457 4410
rect 3461 4406 3462 4410
rect 3422 4405 3466 4406
rect 3426 4401 3427 4405
rect 3431 4401 3432 4405
rect 3436 4401 3437 4405
rect 3441 4401 3442 4405
rect 3446 4401 3447 4405
rect 3451 4401 3452 4405
rect 3456 4401 3457 4405
rect 3461 4401 3462 4405
rect 3422 4400 3466 4401
rect 3426 4396 3427 4400
rect 3431 4396 3432 4400
rect 3436 4396 3437 4400
rect 3441 4396 3442 4400
rect 3446 4396 3447 4400
rect 3451 4396 3452 4400
rect 3456 4396 3457 4400
rect 3461 4396 3462 4400
rect 3422 4395 3466 4396
rect 3426 4391 3427 4395
rect 3431 4391 3432 4395
rect 3436 4391 3437 4395
rect 3441 4391 3442 4395
rect 3446 4391 3447 4395
rect 3451 4391 3452 4395
rect 3456 4391 3457 4395
rect 3461 4391 3462 4395
rect 3422 4390 3466 4391
rect 3426 4386 3427 4390
rect 3431 4386 3432 4390
rect 3436 4386 3437 4390
rect 3441 4386 3442 4390
rect 3446 4386 3447 4390
rect 3451 4386 3452 4390
rect 3456 4386 3457 4390
rect 3461 4386 3462 4390
rect 3422 4385 3466 4386
rect 3426 4381 3427 4385
rect 3431 4381 3432 4385
rect 3436 4381 3437 4385
rect 3441 4381 3442 4385
rect 3446 4381 3447 4385
rect 3451 4381 3452 4385
rect 3456 4381 3457 4385
rect 3461 4381 3462 4385
rect 3422 4380 3466 4381
rect 3426 4376 3427 4380
rect 3431 4376 3432 4380
rect 3436 4376 3437 4380
rect 3441 4376 3442 4380
rect 3446 4376 3447 4380
rect 3451 4376 3452 4380
rect 3456 4376 3457 4380
rect 3461 4376 3462 4380
rect 3422 4375 3466 4376
rect 3426 4371 3427 4375
rect 3431 4371 3432 4375
rect 3436 4371 3437 4375
rect 3441 4371 3442 4375
rect 3446 4371 3447 4375
rect 3451 4371 3452 4375
rect 3456 4371 3457 4375
rect 3461 4371 3462 4375
rect 3422 4370 3466 4371
rect 3426 4366 3427 4370
rect 3431 4366 3432 4370
rect 3436 4366 3437 4370
rect 3441 4366 3442 4370
rect 3446 4366 3447 4370
rect 3451 4366 3452 4370
rect 3456 4366 3457 4370
rect 3461 4366 3462 4370
rect 3422 4365 3466 4366
rect 3426 4361 3427 4365
rect 3431 4361 3432 4365
rect 3436 4361 3437 4365
rect 3441 4361 3442 4365
rect 3446 4361 3447 4365
rect 3451 4361 3452 4365
rect 3456 4361 3457 4365
rect 3461 4361 3462 4365
rect 3474 4445 3478 4446
rect 3474 4440 3478 4441
rect 3474 4435 3478 4436
rect 3474 4430 3478 4431
rect 3474 4425 3478 4426
rect 3474 4420 3478 4421
rect 3474 4415 3478 4416
rect 3474 4410 3478 4411
rect 3474 4405 3478 4406
rect 3474 4400 3478 4401
rect 3474 4395 3478 4396
rect 3474 4390 3478 4391
rect 3474 4385 3478 4386
rect 3474 4380 3478 4381
rect 3474 4375 3478 4376
rect 3474 4370 3478 4371
rect 3474 4365 3478 4366
rect 3410 4360 3414 4361
rect 3410 4353 3414 4356
rect 3474 4360 3478 4361
rect 3474 4353 3478 4356
rect 3414 4349 3417 4353
rect 3421 4349 3422 4353
rect 3426 4349 3427 4353
rect 3431 4349 3432 4353
rect 3436 4349 3437 4353
rect 3441 4349 3442 4353
rect 3446 4349 3447 4353
rect 3451 4349 3452 4353
rect 3456 4349 3457 4353
rect 3461 4349 3462 4353
rect 3466 4349 3467 4353
rect 3471 4349 3474 4353
rect 3487 4465 3491 4466
rect 3487 4460 3491 4461
rect 3487 4455 3491 4456
rect 3487 4450 3491 4451
rect 3487 4445 3491 4446
rect 3487 4440 3491 4441
rect 3487 4435 3491 4436
rect 3487 4430 3491 4431
rect 3487 4425 3491 4426
rect 3487 4420 3491 4421
rect 3487 4415 3491 4416
rect 3487 4410 3491 4411
rect 3487 4405 3491 4406
rect 3487 4400 3491 4401
rect 3487 4395 3491 4396
rect 3487 4390 3491 4391
rect 3487 4385 3491 4386
rect 3487 4380 3491 4381
rect 3487 4375 3491 4376
rect 3487 4370 3491 4371
rect 3487 4365 3491 4366
rect 3487 4360 3491 4361
rect 3487 4355 3491 4356
rect 3487 4350 3491 4351
rect 3397 4345 3401 4346
rect 3397 4340 3401 4341
rect 3487 4345 3491 4346
rect 3487 4340 3491 4341
rect 3401 4336 3402 4340
rect 3406 4336 3407 4340
rect 3411 4336 3412 4340
rect 3416 4336 3417 4340
rect 3421 4336 3422 4340
rect 3426 4336 3427 4340
rect 3431 4336 3432 4340
rect 3436 4336 3437 4340
rect 3441 4336 3442 4340
rect 3446 4336 3447 4340
rect 3451 4336 3452 4340
rect 3456 4336 3457 4340
rect 3461 4336 3462 4340
rect 3466 4336 3467 4340
rect 3471 4336 3472 4340
rect 3476 4336 3477 4340
rect 3481 4336 3482 4340
rect 3486 4336 3487 4340
rect 3550 4471 3551 4475
rect 3555 4471 3556 4475
rect 3560 4471 3561 4475
rect 3565 4471 3566 4475
rect 3570 4471 3571 4475
rect 3575 4471 3576 4475
rect 3580 4471 3581 4475
rect 3585 4471 3586 4475
rect 3590 4471 3591 4475
rect 3595 4471 3596 4475
rect 3600 4471 3601 4475
rect 3605 4471 3606 4475
rect 3610 4471 3611 4475
rect 3615 4471 3616 4475
rect 3620 4471 3621 4475
rect 3625 4471 3626 4475
rect 3630 4471 3631 4475
rect 3635 4471 3636 4475
rect 3546 4470 3550 4471
rect 3636 4470 3640 4471
rect 3546 4465 3550 4466
rect 3546 4460 3550 4461
rect 3546 4455 3550 4456
rect 3546 4450 3550 4451
rect 3546 4445 3550 4446
rect 3546 4440 3550 4441
rect 3546 4435 3550 4436
rect 3546 4430 3550 4431
rect 3546 4425 3550 4426
rect 3546 4420 3550 4421
rect 3546 4415 3550 4416
rect 3546 4410 3550 4411
rect 3546 4405 3550 4406
rect 3546 4400 3550 4401
rect 3546 4395 3550 4396
rect 3546 4390 3550 4391
rect 3546 4385 3550 4386
rect 3546 4380 3550 4381
rect 3546 4375 3550 4376
rect 3546 4370 3550 4371
rect 3546 4365 3550 4366
rect 3546 4360 3550 4361
rect 3546 4355 3550 4356
rect 3546 4350 3550 4351
rect 3563 4458 3566 4466
rect 3570 4458 3571 4466
rect 3575 4458 3576 4466
rect 3580 4458 3581 4466
rect 3585 4458 3586 4466
rect 3590 4458 3591 4466
rect 3595 4458 3596 4466
rect 3600 4458 3601 4466
rect 3605 4458 3606 4466
rect 3610 4458 3611 4466
rect 3615 4458 3616 4466
rect 3620 4458 3623 4466
rect 3559 4455 3563 4458
rect 3559 4450 3563 4451
rect 3623 4455 3627 4458
rect 3623 4450 3627 4451
rect 3559 4445 3563 4446
rect 3559 4440 3563 4441
rect 3559 4435 3563 4436
rect 3559 4430 3563 4431
rect 3559 4425 3563 4426
rect 3559 4420 3563 4421
rect 3559 4415 3563 4416
rect 3559 4410 3563 4411
rect 3559 4405 3563 4406
rect 3559 4400 3563 4401
rect 3559 4395 3563 4396
rect 3559 4390 3563 4391
rect 3559 4385 3563 4386
rect 3559 4380 3563 4381
rect 3559 4375 3563 4376
rect 3559 4370 3563 4371
rect 3559 4365 3563 4366
rect 3575 4446 3576 4450
rect 3580 4446 3581 4450
rect 3585 4446 3586 4450
rect 3590 4446 3591 4450
rect 3595 4446 3596 4450
rect 3600 4446 3601 4450
rect 3605 4446 3606 4450
rect 3610 4446 3611 4450
rect 3615 4446 3616 4450
rect 3571 4445 3616 4446
rect 3575 4441 3576 4445
rect 3580 4441 3581 4445
rect 3585 4441 3586 4445
rect 3590 4441 3591 4445
rect 3595 4441 3596 4445
rect 3600 4441 3601 4445
rect 3605 4441 3606 4445
rect 3610 4441 3611 4445
rect 3615 4441 3616 4445
rect 3571 4440 3616 4441
rect 3575 4436 3576 4440
rect 3580 4436 3581 4440
rect 3585 4436 3586 4440
rect 3590 4436 3591 4440
rect 3595 4436 3596 4440
rect 3600 4436 3601 4440
rect 3605 4436 3606 4440
rect 3610 4436 3611 4440
rect 3615 4436 3616 4440
rect 3571 4435 3616 4436
rect 3575 4431 3576 4435
rect 3580 4431 3581 4435
rect 3585 4431 3586 4435
rect 3590 4431 3591 4435
rect 3595 4431 3596 4435
rect 3600 4431 3601 4435
rect 3605 4431 3606 4435
rect 3610 4431 3611 4435
rect 3615 4431 3616 4435
rect 3571 4430 3616 4431
rect 3575 4426 3576 4430
rect 3580 4426 3581 4430
rect 3585 4426 3586 4430
rect 3590 4426 3591 4430
rect 3595 4426 3596 4430
rect 3600 4426 3601 4430
rect 3605 4426 3606 4430
rect 3610 4426 3611 4430
rect 3615 4426 3616 4430
rect 3571 4425 3616 4426
rect 3575 4421 3576 4425
rect 3580 4421 3581 4425
rect 3585 4421 3586 4425
rect 3590 4421 3591 4425
rect 3595 4421 3596 4425
rect 3600 4421 3601 4425
rect 3605 4421 3606 4425
rect 3610 4421 3611 4425
rect 3615 4421 3616 4425
rect 3571 4420 3616 4421
rect 3575 4416 3576 4420
rect 3580 4416 3581 4420
rect 3585 4416 3586 4420
rect 3590 4416 3591 4420
rect 3595 4416 3596 4420
rect 3600 4416 3601 4420
rect 3605 4416 3606 4420
rect 3610 4416 3611 4420
rect 3615 4416 3616 4420
rect 3571 4415 3616 4416
rect 3575 4411 3576 4415
rect 3580 4411 3581 4415
rect 3585 4411 3586 4415
rect 3590 4411 3591 4415
rect 3595 4411 3596 4415
rect 3600 4411 3601 4415
rect 3605 4411 3606 4415
rect 3610 4411 3611 4415
rect 3615 4411 3616 4415
rect 3571 4410 3616 4411
rect 3575 4406 3576 4410
rect 3580 4406 3581 4410
rect 3585 4406 3586 4410
rect 3590 4406 3591 4410
rect 3595 4406 3596 4410
rect 3600 4406 3601 4410
rect 3605 4406 3606 4410
rect 3610 4406 3611 4410
rect 3615 4406 3616 4410
rect 3571 4405 3616 4406
rect 3575 4401 3576 4405
rect 3580 4401 3581 4405
rect 3585 4401 3586 4405
rect 3590 4401 3591 4405
rect 3595 4401 3596 4405
rect 3600 4401 3601 4405
rect 3605 4401 3606 4405
rect 3610 4401 3611 4405
rect 3615 4401 3616 4405
rect 3571 4400 3616 4401
rect 3575 4396 3576 4400
rect 3580 4396 3581 4400
rect 3585 4396 3586 4400
rect 3590 4396 3591 4400
rect 3595 4396 3596 4400
rect 3600 4396 3601 4400
rect 3605 4396 3606 4400
rect 3610 4396 3611 4400
rect 3615 4396 3616 4400
rect 3571 4395 3616 4396
rect 3575 4391 3576 4395
rect 3580 4391 3581 4395
rect 3585 4391 3586 4395
rect 3590 4391 3591 4395
rect 3595 4391 3596 4395
rect 3600 4391 3601 4395
rect 3605 4391 3606 4395
rect 3610 4391 3611 4395
rect 3615 4391 3616 4395
rect 3571 4390 3616 4391
rect 3575 4386 3576 4390
rect 3580 4386 3581 4390
rect 3585 4386 3586 4390
rect 3590 4386 3591 4390
rect 3595 4386 3596 4390
rect 3600 4386 3601 4390
rect 3605 4386 3606 4390
rect 3610 4386 3611 4390
rect 3615 4386 3616 4390
rect 3571 4385 3616 4386
rect 3575 4381 3576 4385
rect 3580 4381 3581 4385
rect 3585 4381 3586 4385
rect 3590 4381 3591 4385
rect 3595 4381 3596 4385
rect 3600 4381 3601 4385
rect 3605 4381 3606 4385
rect 3610 4381 3611 4385
rect 3615 4381 3616 4385
rect 3571 4380 3616 4381
rect 3575 4376 3576 4380
rect 3580 4376 3581 4380
rect 3585 4376 3586 4380
rect 3590 4376 3591 4380
rect 3595 4376 3596 4380
rect 3600 4376 3601 4380
rect 3605 4376 3606 4380
rect 3610 4376 3611 4380
rect 3615 4376 3616 4380
rect 3571 4375 3616 4376
rect 3575 4371 3576 4375
rect 3580 4371 3581 4375
rect 3585 4371 3586 4375
rect 3590 4371 3591 4375
rect 3595 4371 3596 4375
rect 3600 4371 3601 4375
rect 3605 4371 3606 4375
rect 3610 4371 3611 4375
rect 3615 4371 3616 4375
rect 3571 4370 3616 4371
rect 3575 4366 3576 4370
rect 3580 4366 3581 4370
rect 3585 4366 3586 4370
rect 3590 4366 3591 4370
rect 3595 4366 3596 4370
rect 3600 4366 3601 4370
rect 3605 4366 3606 4370
rect 3610 4366 3611 4370
rect 3615 4366 3616 4370
rect 3571 4365 3616 4366
rect 3575 4361 3576 4365
rect 3580 4361 3581 4365
rect 3585 4361 3586 4365
rect 3590 4361 3591 4365
rect 3595 4361 3596 4365
rect 3600 4361 3601 4365
rect 3605 4361 3606 4365
rect 3610 4361 3611 4365
rect 3615 4361 3616 4365
rect 3623 4445 3627 4446
rect 3623 4440 3627 4441
rect 3623 4435 3627 4436
rect 3623 4430 3627 4431
rect 3623 4425 3627 4426
rect 3623 4420 3627 4421
rect 3623 4415 3627 4416
rect 3623 4410 3627 4411
rect 3623 4405 3627 4406
rect 3623 4400 3627 4401
rect 3623 4395 3627 4396
rect 3623 4390 3627 4391
rect 3623 4385 3627 4386
rect 3623 4380 3627 4381
rect 3623 4375 3627 4376
rect 3623 4370 3627 4371
rect 3623 4365 3627 4366
rect 3559 4360 3563 4361
rect 3559 4353 3563 4356
rect 3623 4360 3627 4361
rect 3623 4353 3627 4356
rect 3563 4349 3566 4353
rect 3570 4349 3571 4353
rect 3575 4349 3576 4353
rect 3580 4349 3581 4353
rect 3585 4349 3586 4353
rect 3590 4349 3591 4353
rect 3595 4349 3596 4353
rect 3600 4349 3601 4353
rect 3605 4349 3606 4353
rect 3610 4349 3611 4353
rect 3615 4349 3616 4353
rect 3620 4349 3623 4353
rect 3636 4465 3640 4466
rect 3636 4460 3640 4461
rect 3636 4455 3640 4456
rect 3636 4450 3640 4451
rect 3636 4445 3640 4446
rect 3636 4440 3640 4441
rect 3636 4435 3640 4436
rect 3636 4430 3640 4431
rect 3636 4425 3640 4426
rect 3636 4420 3640 4421
rect 3636 4415 3640 4416
rect 3636 4410 3640 4411
rect 3636 4405 3640 4406
rect 3636 4400 3640 4401
rect 3636 4395 3640 4396
rect 3636 4390 3640 4391
rect 3636 4385 3640 4386
rect 3636 4380 3640 4381
rect 3636 4375 3640 4376
rect 3636 4370 3640 4371
rect 3636 4365 3640 4366
rect 3636 4360 3640 4361
rect 3636 4355 3640 4356
rect 3636 4350 3640 4351
rect 3546 4345 3550 4346
rect 3546 4340 3550 4341
rect 3636 4345 3640 4346
rect 3636 4340 3640 4341
rect 3550 4336 3551 4340
rect 3555 4336 3556 4340
rect 3560 4336 3561 4340
rect 3565 4336 3566 4340
rect 3570 4336 3571 4340
rect 3575 4336 3576 4340
rect 3580 4336 3581 4340
rect 3585 4336 3586 4340
rect 3590 4336 3591 4340
rect 3595 4336 3596 4340
rect 3600 4336 3601 4340
rect 3605 4336 3606 4340
rect 3610 4336 3611 4340
rect 3615 4336 3616 4340
rect 3620 4336 3621 4340
rect 3625 4336 3626 4340
rect 3630 4336 3631 4340
rect 3635 4336 3636 4340
rect 3647 4333 3699 4599
rect 3838 4624 3839 4628
rect 3843 4624 3844 4628
rect 3848 4624 3849 4628
rect 3834 4623 3853 4624
rect 3838 4619 3839 4623
rect 3843 4619 3844 4623
rect 3848 4619 3849 4623
rect 3834 4618 3853 4619
rect 3838 4614 3839 4618
rect 3843 4614 3844 4618
rect 3848 4614 3849 4618
rect 3834 4613 3853 4614
rect 3838 4609 3839 4613
rect 3843 4609 3844 4613
rect 3848 4609 3849 4613
rect 3834 4608 3853 4609
rect 3838 4604 3839 4608
rect 3843 4604 3844 4608
rect 3848 4604 3849 4608
rect 3834 4603 3853 4604
rect 3838 4599 3839 4603
rect 3843 4599 3844 4603
rect 3848 4599 3849 4603
rect 3834 4598 3853 4599
rect 3838 4594 3839 4598
rect 3843 4594 3844 4598
rect 3848 4594 3849 4598
rect 3741 4578 3809 4580
rect 3741 4574 3799 4578
rect 3803 4574 3804 4578
rect 3808 4574 3809 4578
rect 3741 4573 3809 4574
rect 3741 4569 3799 4573
rect 3803 4569 3804 4573
rect 3808 4569 3809 4573
rect 3741 4568 3809 4569
rect 3741 4564 3799 4568
rect 3803 4564 3804 4568
rect 3808 4564 3809 4568
rect 3741 4563 3809 4564
rect 3741 4559 3799 4563
rect 3803 4559 3804 4563
rect 3808 4559 3809 4563
rect 3741 4558 3809 4559
rect 3741 4554 3799 4558
rect 3803 4554 3804 4558
rect 3808 4554 3809 4558
rect 3741 4553 3809 4554
rect 3741 4549 3799 4553
rect 3803 4549 3804 4553
rect 3808 4549 3809 4553
rect 3741 4548 3809 4549
rect 3838 4578 3839 4582
rect 3843 4578 3844 4582
rect 3848 4578 3849 4582
rect 3834 4577 3853 4578
rect 3838 4573 3839 4577
rect 3843 4573 3844 4577
rect 3848 4573 3849 4577
rect 3834 4572 3853 4573
rect 3838 4568 3839 4572
rect 3843 4568 3844 4572
rect 3848 4568 3849 4572
rect 3834 4567 3853 4568
rect 3838 4563 3839 4567
rect 3843 4563 3844 4567
rect 3848 4563 3849 4567
rect 3834 4562 3853 4563
rect 3838 4558 3839 4562
rect 3843 4558 3844 4562
rect 3848 4558 3849 4562
rect 3834 4557 3853 4558
rect 3838 4553 3839 4557
rect 3843 4553 3844 4557
rect 3848 4553 3849 4557
rect 3834 4552 3853 4553
rect 3838 4548 3839 4552
rect 3843 4548 3844 4552
rect 3848 4548 3849 4552
rect 3741 4544 3799 4548
rect 3803 4544 3804 4548
rect 3808 4544 3809 4548
rect 3741 4543 3809 4544
rect 3741 4539 3799 4543
rect 3803 4539 3804 4543
rect 3808 4539 3809 4543
rect 3741 4538 3809 4539
rect 3741 4534 3799 4538
rect 3803 4534 3804 4538
rect 3808 4534 3809 4538
rect 3741 4533 3809 4534
rect 3741 4529 3799 4533
rect 3803 4529 3804 4533
rect 3808 4529 3809 4533
rect 3741 4528 3809 4529
rect 3741 4524 3799 4528
rect 3803 4524 3804 4528
rect 3808 4524 3809 4528
rect 3741 4523 3809 4524
rect 3741 4519 3799 4523
rect 3803 4519 3804 4523
rect 3808 4519 3809 4523
rect 3741 4518 3809 4519
rect 3741 4514 3799 4518
rect 3803 4514 3804 4518
rect 3808 4514 3809 4518
rect 3741 4512 3809 4514
rect 3741 4475 3797 4512
rect 3710 4471 3711 4475
rect 3715 4471 3716 4475
rect 3720 4471 3721 4475
rect 3725 4471 3726 4475
rect 3730 4471 3731 4475
rect 3735 4471 3736 4475
rect 3740 4471 3741 4475
rect 3745 4471 3746 4475
rect 3750 4471 3751 4475
rect 3755 4471 3756 4475
rect 3760 4471 3761 4475
rect 3765 4471 3766 4475
rect 3770 4471 3771 4475
rect 3775 4471 3776 4475
rect 3780 4471 3781 4475
rect 3785 4471 3786 4475
rect 3790 4471 3791 4475
rect 3795 4471 3796 4475
rect 3706 4470 3710 4471
rect 3796 4470 3800 4471
rect 3706 4465 3710 4466
rect 3706 4460 3710 4461
rect 3706 4455 3710 4456
rect 3706 4450 3710 4451
rect 3706 4445 3710 4446
rect 3706 4440 3710 4441
rect 3706 4435 3710 4436
rect 3706 4430 3710 4431
rect 3706 4425 3710 4426
rect 3706 4420 3710 4421
rect 3706 4415 3710 4416
rect 3706 4410 3710 4411
rect 3706 4405 3710 4406
rect 3706 4400 3710 4401
rect 3706 4395 3710 4396
rect 3706 4390 3710 4391
rect 3706 4385 3710 4386
rect 3706 4380 3710 4381
rect 3706 4375 3710 4376
rect 3706 4370 3710 4371
rect 3706 4365 3710 4366
rect 3706 4360 3710 4361
rect 3706 4355 3710 4356
rect 3706 4350 3710 4351
rect 3723 4458 3726 4466
rect 3730 4458 3731 4466
rect 3735 4458 3736 4466
rect 3740 4458 3741 4466
rect 3745 4458 3746 4466
rect 3750 4458 3751 4466
rect 3755 4458 3756 4466
rect 3760 4458 3761 4466
rect 3765 4458 3766 4466
rect 3770 4458 3771 4466
rect 3775 4458 3776 4466
rect 3780 4458 3783 4466
rect 3719 4455 3723 4458
rect 3719 4450 3723 4451
rect 3783 4455 3787 4458
rect 3783 4450 3787 4451
rect 3719 4445 3723 4446
rect 3719 4440 3723 4441
rect 3719 4435 3723 4436
rect 3719 4430 3723 4431
rect 3719 4425 3723 4426
rect 3719 4420 3723 4421
rect 3719 4415 3723 4416
rect 3719 4410 3723 4411
rect 3719 4405 3723 4406
rect 3719 4400 3723 4401
rect 3719 4395 3723 4396
rect 3719 4390 3723 4391
rect 3719 4385 3723 4386
rect 3719 4380 3723 4381
rect 3719 4375 3723 4376
rect 3719 4370 3723 4371
rect 3719 4365 3723 4366
rect 3735 4446 3736 4450
rect 3740 4446 3741 4450
rect 3745 4446 3746 4450
rect 3750 4446 3751 4450
rect 3755 4446 3756 4450
rect 3760 4446 3761 4450
rect 3765 4446 3766 4450
rect 3770 4446 3771 4450
rect 3731 4445 3775 4446
rect 3735 4441 3736 4445
rect 3740 4441 3741 4445
rect 3745 4441 3746 4445
rect 3750 4441 3751 4445
rect 3755 4441 3756 4445
rect 3760 4441 3761 4445
rect 3765 4441 3766 4445
rect 3770 4441 3771 4445
rect 3731 4440 3775 4441
rect 3735 4436 3736 4440
rect 3740 4436 3741 4440
rect 3745 4436 3746 4440
rect 3750 4436 3751 4440
rect 3755 4436 3756 4440
rect 3760 4436 3761 4440
rect 3765 4436 3766 4440
rect 3770 4436 3771 4440
rect 3731 4435 3775 4436
rect 3735 4431 3736 4435
rect 3740 4431 3741 4435
rect 3745 4431 3746 4435
rect 3750 4431 3751 4435
rect 3755 4431 3756 4435
rect 3760 4431 3761 4435
rect 3765 4431 3766 4435
rect 3770 4431 3771 4435
rect 3731 4430 3775 4431
rect 3735 4426 3736 4430
rect 3740 4426 3741 4430
rect 3745 4426 3746 4430
rect 3750 4426 3751 4430
rect 3755 4426 3756 4430
rect 3760 4426 3761 4430
rect 3765 4426 3766 4430
rect 3770 4426 3771 4430
rect 3731 4425 3775 4426
rect 3735 4421 3736 4425
rect 3740 4421 3741 4425
rect 3745 4421 3746 4425
rect 3750 4421 3751 4425
rect 3755 4421 3756 4425
rect 3760 4421 3761 4425
rect 3765 4421 3766 4425
rect 3770 4421 3771 4425
rect 3731 4420 3775 4421
rect 3735 4416 3736 4420
rect 3740 4416 3741 4420
rect 3745 4416 3746 4420
rect 3750 4416 3751 4420
rect 3755 4416 3756 4420
rect 3760 4416 3761 4420
rect 3765 4416 3766 4420
rect 3770 4416 3771 4420
rect 3731 4415 3775 4416
rect 3735 4411 3736 4415
rect 3740 4411 3741 4415
rect 3745 4411 3746 4415
rect 3750 4411 3751 4415
rect 3755 4411 3756 4415
rect 3760 4411 3761 4415
rect 3765 4411 3766 4415
rect 3770 4411 3771 4415
rect 3731 4410 3775 4411
rect 3735 4406 3736 4410
rect 3740 4406 3741 4410
rect 3745 4406 3746 4410
rect 3750 4406 3751 4410
rect 3755 4406 3756 4410
rect 3760 4406 3761 4410
rect 3765 4406 3766 4410
rect 3770 4406 3771 4410
rect 3731 4405 3775 4406
rect 3735 4401 3736 4405
rect 3740 4401 3741 4405
rect 3745 4401 3746 4405
rect 3750 4401 3751 4405
rect 3755 4401 3756 4405
rect 3760 4401 3761 4405
rect 3765 4401 3766 4405
rect 3770 4401 3771 4405
rect 3731 4400 3775 4401
rect 3735 4396 3736 4400
rect 3740 4396 3741 4400
rect 3745 4396 3746 4400
rect 3750 4396 3751 4400
rect 3755 4396 3756 4400
rect 3760 4396 3761 4400
rect 3765 4396 3766 4400
rect 3770 4396 3771 4400
rect 3731 4395 3775 4396
rect 3735 4391 3736 4395
rect 3740 4391 3741 4395
rect 3745 4391 3746 4395
rect 3750 4391 3751 4395
rect 3755 4391 3756 4395
rect 3760 4391 3761 4395
rect 3765 4391 3766 4395
rect 3770 4391 3771 4395
rect 3731 4390 3775 4391
rect 3735 4386 3736 4390
rect 3740 4386 3741 4390
rect 3745 4386 3746 4390
rect 3750 4386 3751 4390
rect 3755 4386 3756 4390
rect 3760 4386 3761 4390
rect 3765 4386 3766 4390
rect 3770 4386 3771 4390
rect 3731 4385 3775 4386
rect 3735 4381 3736 4385
rect 3740 4381 3741 4385
rect 3745 4381 3746 4385
rect 3750 4381 3751 4385
rect 3755 4381 3756 4385
rect 3760 4381 3761 4385
rect 3765 4381 3766 4385
rect 3770 4381 3771 4385
rect 3731 4380 3775 4381
rect 3735 4376 3736 4380
rect 3740 4376 3741 4380
rect 3745 4376 3746 4380
rect 3750 4376 3751 4380
rect 3755 4376 3756 4380
rect 3760 4376 3761 4380
rect 3765 4376 3766 4380
rect 3770 4376 3771 4380
rect 3731 4375 3775 4376
rect 3735 4371 3736 4375
rect 3740 4371 3741 4375
rect 3745 4371 3746 4375
rect 3750 4371 3751 4375
rect 3755 4371 3756 4375
rect 3760 4371 3761 4375
rect 3765 4371 3766 4375
rect 3770 4371 3771 4375
rect 3731 4370 3775 4371
rect 3735 4366 3736 4370
rect 3740 4366 3741 4370
rect 3745 4366 3746 4370
rect 3750 4366 3751 4370
rect 3755 4366 3756 4370
rect 3760 4366 3761 4370
rect 3765 4366 3766 4370
rect 3770 4366 3771 4370
rect 3731 4365 3775 4366
rect 3735 4361 3736 4365
rect 3740 4361 3741 4365
rect 3745 4361 3746 4365
rect 3750 4361 3751 4365
rect 3755 4361 3756 4365
rect 3760 4361 3761 4365
rect 3765 4361 3766 4365
rect 3770 4361 3771 4365
rect 3783 4445 3787 4446
rect 3783 4440 3787 4441
rect 3783 4435 3787 4436
rect 3783 4430 3787 4431
rect 3783 4425 3787 4426
rect 3783 4420 3787 4421
rect 3783 4415 3787 4416
rect 3783 4410 3787 4411
rect 3783 4405 3787 4406
rect 3783 4400 3787 4401
rect 3783 4395 3787 4396
rect 3783 4390 3787 4391
rect 3783 4385 3787 4386
rect 3783 4380 3787 4381
rect 3783 4375 3787 4376
rect 3783 4370 3787 4371
rect 3783 4365 3787 4366
rect 3719 4360 3723 4361
rect 3719 4353 3723 4356
rect 3783 4360 3787 4361
rect 3783 4353 3787 4356
rect 3723 4349 3726 4353
rect 3730 4349 3731 4353
rect 3735 4349 3736 4353
rect 3740 4349 3741 4353
rect 3745 4349 3746 4353
rect 3750 4349 3751 4353
rect 3755 4349 3756 4353
rect 3760 4349 3761 4353
rect 3765 4349 3766 4353
rect 3770 4349 3771 4353
rect 3775 4349 3776 4353
rect 3780 4349 3783 4353
rect 3796 4465 3800 4466
rect 3796 4460 3800 4461
rect 3796 4455 3800 4456
rect 3796 4450 3800 4451
rect 3796 4445 3800 4446
rect 3796 4440 3800 4441
rect 3796 4435 3800 4436
rect 3796 4430 3800 4431
rect 3796 4425 3800 4426
rect 3796 4420 3800 4421
rect 3796 4415 3800 4416
rect 3796 4410 3800 4411
rect 3796 4405 3800 4406
rect 3796 4400 3800 4401
rect 3796 4395 3800 4396
rect 3796 4390 3800 4391
rect 3796 4385 3800 4386
rect 3796 4380 3800 4381
rect 3796 4375 3800 4376
rect 3796 4370 3800 4371
rect 3796 4365 3800 4366
rect 3796 4360 3800 4361
rect 3796 4355 3800 4356
rect 3796 4350 3800 4351
rect 3706 4345 3710 4346
rect 3706 4340 3710 4341
rect 3796 4345 3800 4346
rect 3796 4340 3800 4341
rect 3710 4336 3711 4340
rect 3715 4336 3716 4340
rect 3720 4336 3721 4340
rect 3725 4336 3726 4340
rect 3730 4336 3731 4340
rect 3735 4336 3736 4340
rect 3740 4336 3741 4340
rect 3745 4336 3746 4340
rect 3750 4336 3751 4340
rect 3755 4336 3756 4340
rect 3760 4336 3761 4340
rect 3765 4336 3766 4340
rect 3770 4336 3771 4340
rect 3775 4336 3776 4340
rect 3780 4336 3781 4340
rect 3785 4336 3786 4340
rect 3790 4336 3791 4340
rect 3795 4336 3796 4340
rect 1153 4332 1249 4333
rect 1153 4328 1158 4332
rect 1162 4328 1165 4332
rect 1169 4328 1172 4332
rect 1176 4328 1179 4332
rect 1183 4328 1186 4332
rect 1190 4328 1193 4332
rect 1197 4328 1200 4332
rect 1204 4328 1207 4332
rect 1211 4328 1214 4332
rect 1218 4328 1221 4332
rect 1225 4328 1228 4332
rect 1232 4328 1235 4332
rect 1239 4328 1242 4332
rect 1246 4328 1249 4332
rect 1153 4327 1249 4328
rect 1153 4323 1158 4327
rect 1162 4323 1165 4327
rect 1169 4323 1172 4327
rect 1176 4323 1179 4327
rect 1183 4323 1186 4327
rect 1190 4323 1193 4327
rect 1197 4323 1200 4327
rect 1204 4323 1207 4327
rect 1211 4323 1214 4327
rect 1218 4323 1221 4327
rect 1225 4323 1228 4327
rect 1232 4323 1235 4327
rect 1239 4323 1242 4327
rect 1246 4323 1249 4327
rect 1153 4322 1249 4323
rect 1153 4321 1158 4322
rect 1143 4318 1158 4321
rect 1162 4318 1165 4322
rect 1169 4318 1172 4322
rect 1176 4318 1179 4322
rect 1183 4318 1186 4322
rect 1190 4318 1193 4322
rect 1197 4318 1200 4322
rect 1204 4318 1207 4322
rect 1211 4318 1214 4322
rect 1218 4318 1221 4322
rect 1225 4318 1228 4322
rect 1232 4318 1235 4322
rect 1239 4318 1242 4322
rect 1246 4321 1249 4322
rect 1462 4332 1558 4333
rect 1462 4328 1467 4332
rect 1471 4328 1474 4332
rect 1478 4328 1481 4332
rect 1485 4328 1488 4332
rect 1492 4328 1495 4332
rect 1499 4328 1502 4332
rect 1506 4328 1509 4332
rect 1513 4328 1516 4332
rect 1520 4328 1523 4332
rect 1527 4328 1530 4332
rect 1534 4328 1537 4332
rect 1541 4328 1544 4332
rect 1548 4328 1551 4332
rect 1555 4328 1558 4332
rect 1462 4327 1558 4328
rect 1462 4323 1467 4327
rect 1471 4323 1474 4327
rect 1478 4323 1481 4327
rect 1485 4323 1488 4327
rect 1492 4323 1495 4327
rect 1499 4323 1502 4327
rect 1506 4323 1509 4327
rect 1513 4323 1516 4327
rect 1520 4323 1523 4327
rect 1527 4323 1530 4327
rect 1534 4323 1537 4327
rect 1541 4323 1544 4327
rect 1548 4323 1551 4327
rect 1555 4323 1558 4327
rect 1462 4322 1558 4323
rect 1462 4321 1467 4322
rect 1246 4318 1259 4321
rect 1143 4317 1259 4318
rect 1143 4313 1158 4317
rect 1162 4313 1165 4317
rect 1169 4313 1172 4317
rect 1176 4313 1179 4317
rect 1183 4313 1186 4317
rect 1190 4313 1193 4317
rect 1197 4313 1200 4317
rect 1204 4313 1207 4317
rect 1211 4313 1214 4317
rect 1218 4313 1221 4317
rect 1225 4313 1228 4317
rect 1232 4313 1235 4317
rect 1239 4313 1242 4317
rect 1246 4313 1259 4317
rect 1143 4311 1259 4313
rect 1452 4318 1467 4321
rect 1471 4318 1474 4322
rect 1478 4318 1481 4322
rect 1485 4318 1488 4322
rect 1492 4318 1495 4322
rect 1499 4318 1502 4322
rect 1506 4318 1509 4322
rect 1513 4318 1516 4322
rect 1520 4318 1523 4322
rect 1527 4318 1530 4322
rect 1534 4318 1537 4322
rect 1541 4318 1544 4322
rect 1548 4318 1551 4322
rect 1555 4321 1558 4322
rect 1771 4332 1867 4333
rect 1771 4328 1776 4332
rect 1780 4328 1783 4332
rect 1787 4328 1790 4332
rect 1794 4328 1797 4332
rect 1801 4328 1804 4332
rect 1808 4328 1811 4332
rect 1815 4328 1818 4332
rect 1822 4328 1825 4332
rect 1829 4328 1832 4332
rect 1836 4328 1839 4332
rect 1843 4328 1846 4332
rect 1850 4328 1853 4332
rect 1857 4328 1860 4332
rect 1864 4328 1867 4332
rect 1771 4327 1867 4328
rect 1771 4323 1776 4327
rect 1780 4323 1783 4327
rect 1787 4323 1790 4327
rect 1794 4323 1797 4327
rect 1801 4323 1804 4327
rect 1808 4323 1811 4327
rect 1815 4323 1818 4327
rect 1822 4323 1825 4327
rect 1829 4323 1832 4327
rect 1836 4323 1839 4327
rect 1843 4323 1846 4327
rect 1850 4323 1853 4327
rect 1857 4323 1860 4327
rect 1864 4323 1867 4327
rect 1771 4322 1867 4323
rect 1771 4321 1776 4322
rect 1555 4318 1568 4321
rect 1452 4317 1568 4318
rect 1452 4313 1467 4317
rect 1471 4313 1474 4317
rect 1478 4313 1481 4317
rect 1485 4313 1488 4317
rect 1492 4313 1495 4317
rect 1499 4313 1502 4317
rect 1506 4313 1509 4317
rect 1513 4313 1516 4317
rect 1520 4313 1523 4317
rect 1527 4313 1530 4317
rect 1534 4313 1537 4317
rect 1541 4313 1544 4317
rect 1548 4313 1551 4317
rect 1555 4313 1568 4317
rect 1452 4311 1568 4313
rect 1761 4318 1776 4321
rect 1780 4318 1783 4322
rect 1787 4318 1790 4322
rect 1794 4318 1797 4322
rect 1801 4318 1804 4322
rect 1808 4318 1811 4322
rect 1815 4318 1818 4322
rect 1822 4318 1825 4322
rect 1829 4318 1832 4322
rect 1836 4318 1839 4322
rect 1843 4318 1846 4322
rect 1850 4318 1853 4322
rect 1857 4318 1860 4322
rect 1864 4321 1867 4322
rect 2080 4332 2176 4333
rect 2080 4328 2085 4332
rect 2089 4328 2092 4332
rect 2096 4328 2099 4332
rect 2103 4328 2106 4332
rect 2110 4328 2113 4332
rect 2117 4328 2120 4332
rect 2124 4328 2127 4332
rect 2131 4328 2134 4332
rect 2138 4328 2141 4332
rect 2145 4328 2148 4332
rect 2152 4328 2155 4332
rect 2159 4328 2162 4332
rect 2166 4328 2169 4332
rect 2173 4328 2176 4332
rect 2080 4327 2176 4328
rect 2080 4323 2085 4327
rect 2089 4323 2092 4327
rect 2096 4323 2099 4327
rect 2103 4323 2106 4327
rect 2110 4323 2113 4327
rect 2117 4323 2120 4327
rect 2124 4323 2127 4327
rect 2131 4323 2134 4327
rect 2138 4323 2141 4327
rect 2145 4323 2148 4327
rect 2152 4323 2155 4327
rect 2159 4323 2162 4327
rect 2166 4323 2169 4327
rect 2173 4323 2176 4327
rect 2080 4322 2176 4323
rect 2080 4321 2085 4322
rect 1864 4318 1877 4321
rect 1761 4317 1877 4318
rect 1761 4313 1776 4317
rect 1780 4313 1783 4317
rect 1787 4313 1790 4317
rect 1794 4313 1797 4317
rect 1801 4313 1804 4317
rect 1808 4313 1811 4317
rect 1815 4313 1818 4317
rect 1822 4313 1825 4317
rect 1829 4313 1832 4317
rect 1836 4313 1839 4317
rect 1843 4313 1846 4317
rect 1850 4313 1853 4317
rect 1857 4313 1860 4317
rect 1864 4313 1877 4317
rect 1761 4311 1877 4313
rect 2070 4318 2085 4321
rect 2089 4318 2092 4322
rect 2096 4318 2099 4322
rect 2103 4318 2106 4322
rect 2110 4318 2113 4322
rect 2117 4318 2120 4322
rect 2124 4318 2127 4322
rect 2131 4318 2134 4322
rect 2138 4318 2141 4322
rect 2145 4318 2148 4322
rect 2152 4318 2155 4322
rect 2159 4318 2162 4322
rect 2166 4318 2169 4322
rect 2173 4321 2176 4322
rect 2389 4332 2485 4333
rect 2389 4328 2394 4332
rect 2398 4328 2401 4332
rect 2405 4328 2408 4332
rect 2412 4328 2415 4332
rect 2419 4328 2422 4332
rect 2426 4328 2429 4332
rect 2433 4328 2436 4332
rect 2440 4328 2443 4332
rect 2447 4328 2450 4332
rect 2454 4328 2457 4332
rect 2461 4328 2464 4332
rect 2468 4328 2471 4332
rect 2475 4328 2478 4332
rect 2482 4328 2485 4332
rect 2389 4327 2485 4328
rect 2389 4323 2394 4327
rect 2398 4323 2401 4327
rect 2405 4323 2408 4327
rect 2412 4323 2415 4327
rect 2419 4323 2422 4327
rect 2426 4323 2429 4327
rect 2433 4323 2436 4327
rect 2440 4323 2443 4327
rect 2447 4323 2450 4327
rect 2454 4323 2457 4327
rect 2461 4323 2464 4327
rect 2468 4323 2471 4327
rect 2475 4323 2478 4327
rect 2482 4323 2485 4327
rect 2389 4322 2485 4323
rect 2389 4321 2394 4322
rect 2173 4318 2186 4321
rect 2070 4317 2186 4318
rect 2070 4313 2085 4317
rect 2089 4313 2092 4317
rect 2096 4313 2099 4317
rect 2103 4313 2106 4317
rect 2110 4313 2113 4317
rect 2117 4313 2120 4317
rect 2124 4313 2127 4317
rect 2131 4313 2134 4317
rect 2138 4313 2141 4317
rect 2145 4313 2148 4317
rect 2152 4313 2155 4317
rect 2159 4313 2162 4317
rect 2166 4313 2169 4317
rect 2173 4313 2186 4317
rect 2070 4311 2186 4313
rect 2379 4318 2394 4321
rect 2398 4318 2401 4322
rect 2405 4318 2408 4322
rect 2412 4318 2415 4322
rect 2419 4318 2422 4322
rect 2426 4318 2429 4322
rect 2433 4318 2436 4322
rect 2440 4318 2443 4322
rect 2447 4318 2450 4322
rect 2454 4318 2457 4322
rect 2461 4318 2464 4322
rect 2468 4318 2471 4322
rect 2475 4318 2478 4322
rect 2482 4321 2485 4322
rect 2698 4332 2794 4333
rect 2698 4328 2703 4332
rect 2707 4328 2710 4332
rect 2714 4328 2717 4332
rect 2721 4328 2724 4332
rect 2728 4328 2731 4332
rect 2735 4328 2738 4332
rect 2742 4328 2745 4332
rect 2749 4328 2752 4332
rect 2756 4328 2759 4332
rect 2763 4328 2766 4332
rect 2770 4328 2773 4332
rect 2777 4328 2780 4332
rect 2784 4328 2787 4332
rect 2791 4328 2794 4332
rect 2698 4327 2794 4328
rect 2698 4323 2703 4327
rect 2707 4323 2710 4327
rect 2714 4323 2717 4327
rect 2721 4323 2724 4327
rect 2728 4323 2731 4327
rect 2735 4323 2738 4327
rect 2742 4323 2745 4327
rect 2749 4323 2752 4327
rect 2756 4323 2759 4327
rect 2763 4323 2766 4327
rect 2770 4323 2773 4327
rect 2777 4323 2780 4327
rect 2784 4323 2787 4327
rect 2791 4323 2794 4327
rect 2698 4322 2794 4323
rect 2698 4321 2703 4322
rect 2482 4318 2495 4321
rect 2379 4317 2495 4318
rect 2379 4313 2394 4317
rect 2398 4313 2401 4317
rect 2405 4313 2408 4317
rect 2412 4313 2415 4317
rect 2419 4313 2422 4317
rect 2426 4313 2429 4317
rect 2433 4313 2436 4317
rect 2440 4313 2443 4317
rect 2447 4313 2450 4317
rect 2454 4313 2457 4317
rect 2461 4313 2464 4317
rect 2468 4313 2471 4317
rect 2475 4313 2478 4317
rect 2482 4313 2495 4317
rect 2379 4311 2495 4313
rect 2688 4318 2703 4321
rect 2707 4318 2710 4322
rect 2714 4318 2717 4322
rect 2721 4318 2724 4322
rect 2728 4318 2731 4322
rect 2735 4318 2738 4322
rect 2742 4318 2745 4322
rect 2749 4318 2752 4322
rect 2756 4318 2759 4322
rect 2763 4318 2766 4322
rect 2770 4318 2773 4322
rect 2777 4318 2780 4322
rect 2784 4318 2787 4322
rect 2791 4321 2794 4322
rect 3007 4332 3103 4333
rect 3007 4328 3012 4332
rect 3016 4328 3019 4332
rect 3023 4328 3026 4332
rect 3030 4328 3033 4332
rect 3037 4328 3040 4332
rect 3044 4328 3047 4332
rect 3051 4328 3054 4332
rect 3058 4328 3061 4332
rect 3065 4328 3068 4332
rect 3072 4328 3075 4332
rect 3079 4328 3082 4332
rect 3086 4328 3089 4332
rect 3093 4328 3096 4332
rect 3100 4328 3103 4332
rect 3007 4327 3103 4328
rect 3007 4323 3012 4327
rect 3016 4323 3019 4327
rect 3023 4323 3026 4327
rect 3030 4323 3033 4327
rect 3037 4323 3040 4327
rect 3044 4323 3047 4327
rect 3051 4323 3054 4327
rect 3058 4323 3061 4327
rect 3065 4323 3068 4327
rect 3072 4323 3075 4327
rect 3079 4323 3082 4327
rect 3086 4323 3089 4327
rect 3093 4323 3096 4327
rect 3100 4323 3103 4327
rect 3007 4322 3103 4323
rect 3007 4321 3012 4322
rect 2791 4318 2804 4321
rect 2688 4317 2804 4318
rect 2688 4313 2703 4317
rect 2707 4313 2710 4317
rect 2714 4313 2717 4317
rect 2721 4313 2724 4317
rect 2728 4313 2731 4317
rect 2735 4313 2738 4317
rect 2742 4313 2745 4317
rect 2749 4313 2752 4317
rect 2756 4313 2759 4317
rect 2763 4313 2766 4317
rect 2770 4313 2773 4317
rect 2777 4313 2780 4317
rect 2784 4313 2787 4317
rect 2791 4313 2804 4317
rect 2688 4311 2804 4313
rect 2997 4318 3012 4321
rect 3016 4318 3019 4322
rect 3023 4318 3026 4322
rect 3030 4318 3033 4322
rect 3037 4318 3040 4322
rect 3044 4318 3047 4322
rect 3051 4318 3054 4322
rect 3058 4318 3061 4322
rect 3065 4318 3068 4322
rect 3072 4318 3075 4322
rect 3079 4318 3082 4322
rect 3086 4318 3089 4322
rect 3093 4318 3096 4322
rect 3100 4321 3103 4322
rect 3316 4332 3412 4333
rect 3316 4328 3321 4332
rect 3325 4328 3328 4332
rect 3332 4328 3335 4332
rect 3339 4328 3342 4332
rect 3346 4328 3349 4332
rect 3353 4328 3356 4332
rect 3360 4328 3363 4332
rect 3367 4328 3370 4332
rect 3374 4328 3377 4332
rect 3381 4328 3384 4332
rect 3388 4328 3391 4332
rect 3395 4328 3398 4332
rect 3402 4328 3405 4332
rect 3409 4328 3412 4332
rect 3316 4327 3412 4328
rect 3316 4323 3321 4327
rect 3325 4323 3328 4327
rect 3332 4323 3335 4327
rect 3339 4323 3342 4327
rect 3346 4323 3349 4327
rect 3353 4323 3356 4327
rect 3360 4323 3363 4327
rect 3367 4323 3370 4327
rect 3374 4323 3377 4327
rect 3381 4323 3384 4327
rect 3388 4323 3391 4327
rect 3395 4323 3398 4327
rect 3402 4323 3405 4327
rect 3409 4323 3412 4327
rect 3316 4322 3412 4323
rect 3316 4321 3321 4322
rect 3100 4318 3113 4321
rect 2997 4317 3113 4318
rect 2997 4313 3012 4317
rect 3016 4313 3019 4317
rect 3023 4313 3026 4317
rect 3030 4313 3033 4317
rect 3037 4313 3040 4317
rect 3044 4313 3047 4317
rect 3051 4313 3054 4317
rect 3058 4313 3061 4317
rect 3065 4313 3068 4317
rect 3072 4313 3075 4317
rect 3079 4313 3082 4317
rect 3086 4313 3089 4317
rect 3093 4313 3096 4317
rect 3100 4313 3113 4317
rect 2997 4311 3113 4313
rect 3306 4318 3321 4321
rect 3325 4318 3328 4322
rect 3332 4318 3335 4322
rect 3339 4318 3342 4322
rect 3346 4318 3349 4322
rect 3353 4318 3356 4322
rect 3360 4318 3363 4322
rect 3367 4318 3370 4322
rect 3374 4318 3377 4322
rect 3381 4318 3384 4322
rect 3388 4318 3391 4322
rect 3395 4318 3398 4322
rect 3402 4318 3405 4322
rect 3409 4321 3412 4322
rect 3625 4332 3721 4333
rect 3625 4328 3630 4332
rect 3634 4328 3637 4332
rect 3641 4328 3644 4332
rect 3648 4328 3651 4332
rect 3655 4328 3658 4332
rect 3662 4328 3665 4332
rect 3669 4328 3672 4332
rect 3676 4328 3679 4332
rect 3683 4328 3686 4332
rect 3690 4328 3693 4332
rect 3697 4328 3700 4332
rect 3704 4328 3707 4332
rect 3711 4328 3714 4332
rect 3718 4328 3721 4332
rect 3625 4327 3721 4328
rect 3625 4323 3630 4327
rect 3634 4323 3637 4327
rect 3641 4323 3644 4327
rect 3648 4323 3651 4327
rect 3655 4323 3658 4327
rect 3662 4323 3665 4327
rect 3669 4323 3672 4327
rect 3676 4323 3679 4327
rect 3683 4323 3686 4327
rect 3690 4323 3693 4327
rect 3697 4323 3700 4327
rect 3704 4323 3707 4327
rect 3711 4323 3714 4327
rect 3718 4323 3721 4327
rect 3625 4322 3721 4323
rect 3625 4321 3630 4322
rect 3409 4318 3422 4321
rect 3306 4317 3422 4318
rect 3306 4313 3321 4317
rect 3325 4313 3328 4317
rect 3332 4313 3335 4317
rect 3339 4313 3342 4317
rect 3346 4313 3349 4317
rect 3353 4313 3356 4317
rect 3360 4313 3363 4317
rect 3367 4313 3370 4317
rect 3374 4313 3377 4317
rect 3381 4313 3384 4317
rect 3388 4313 3391 4317
rect 3395 4313 3398 4317
rect 3402 4313 3405 4317
rect 3409 4313 3422 4317
rect 3306 4311 3422 4313
rect 3615 4318 3630 4321
rect 3634 4318 3637 4322
rect 3641 4318 3644 4322
rect 3648 4318 3651 4322
rect 3655 4318 3658 4322
rect 3662 4318 3665 4322
rect 3669 4318 3672 4322
rect 3676 4318 3679 4322
rect 3683 4318 3686 4322
rect 3690 4318 3693 4322
rect 3697 4318 3700 4322
rect 3704 4318 3707 4322
rect 3711 4318 3714 4322
rect 3718 4321 3721 4322
rect 3934 4321 4030 4704
rect 4483 4702 4484 4706
rect 4488 4702 4489 4706
rect 4493 4702 4494 4706
rect 4498 4702 4499 4706
rect 4503 4702 4504 4706
rect 4508 4702 4509 4706
rect 4479 4701 4513 4702
rect 4483 4697 4484 4701
rect 4488 4697 4489 4701
rect 4493 4697 4494 4701
rect 4498 4697 4499 4701
rect 4503 4697 4504 4701
rect 4508 4697 4509 4701
rect 4479 4696 4513 4697
rect 4483 4692 4484 4696
rect 4488 4692 4489 4696
rect 4493 4692 4494 4696
rect 4498 4692 4499 4696
rect 4503 4692 4504 4696
rect 4508 4692 4509 4696
rect 4529 4707 4530 4711
rect 4534 4707 4535 4711
rect 4539 4707 4540 4711
rect 4544 4707 4545 4711
rect 4549 4707 4550 4711
rect 4554 4707 4555 4711
rect 4525 4706 4559 4707
rect 4529 4702 4530 4706
rect 4534 4702 4535 4706
rect 4539 4702 4540 4706
rect 4544 4702 4545 4706
rect 4549 4702 4550 4706
rect 4554 4702 4555 4706
rect 4525 4701 4559 4702
rect 4529 4697 4530 4701
rect 4534 4697 4535 4701
rect 4539 4697 4540 4701
rect 4544 4697 4545 4701
rect 4549 4697 4550 4701
rect 4554 4697 4555 4701
rect 4525 4696 4559 4697
rect 4529 4692 4530 4696
rect 4534 4692 4535 4696
rect 4539 4692 4540 4696
rect 4544 4692 4545 4696
rect 4549 4692 4550 4696
rect 4554 4692 4555 4696
rect 4239 4624 4240 4628
rect 4244 4624 4245 4628
rect 4249 4624 4250 4628
rect 4235 4623 4254 4624
rect 4239 4619 4240 4623
rect 4244 4619 4245 4623
rect 4249 4619 4250 4623
rect 4235 4618 4254 4619
rect 4239 4614 4240 4618
rect 4244 4614 4245 4618
rect 4249 4614 4250 4618
rect 4235 4613 4254 4614
rect 4239 4609 4240 4613
rect 4244 4609 4245 4613
rect 4249 4609 4250 4613
rect 4235 4608 4254 4609
rect 4239 4604 4240 4608
rect 4244 4604 4245 4608
rect 4249 4604 4250 4608
rect 4235 4603 4254 4604
rect 4239 4599 4240 4603
rect 4244 4599 4245 4603
rect 4249 4599 4250 4603
rect 4235 4598 4254 4599
rect 4239 4594 4240 4598
rect 4244 4594 4245 4598
rect 4249 4594 4250 4598
rect 4268 4624 4269 4628
rect 4273 4624 4274 4628
rect 4278 4624 4279 4628
rect 4264 4623 4283 4624
rect 4268 4619 4269 4623
rect 4273 4619 4274 4623
rect 4278 4619 4279 4623
rect 4264 4618 4283 4619
rect 4268 4614 4269 4618
rect 4273 4614 4274 4618
rect 4278 4614 4279 4618
rect 4264 4613 4283 4614
rect 4268 4609 4269 4613
rect 4273 4609 4274 4613
rect 4278 4609 4279 4613
rect 4264 4608 4283 4609
rect 4268 4604 4269 4608
rect 4273 4604 4274 4608
rect 4278 4604 4279 4608
rect 4264 4603 4283 4604
rect 4268 4599 4269 4603
rect 4273 4599 4274 4603
rect 4278 4599 4279 4603
rect 4264 4598 4283 4599
rect 4268 4594 4269 4598
rect 4273 4594 4274 4598
rect 4278 4594 4279 4598
rect 4297 4624 4298 4628
rect 4302 4624 4303 4628
rect 4307 4624 4308 4628
rect 4293 4623 4312 4624
rect 4297 4619 4298 4623
rect 4302 4619 4303 4623
rect 4307 4619 4308 4623
rect 4293 4618 4312 4619
rect 4297 4614 4298 4618
rect 4302 4614 4303 4618
rect 4307 4614 4308 4618
rect 4293 4613 4312 4614
rect 4297 4609 4298 4613
rect 4302 4609 4303 4613
rect 4307 4609 4308 4613
rect 4293 4608 4312 4609
rect 4297 4604 4298 4608
rect 4302 4604 4303 4608
rect 4307 4604 4308 4608
rect 4293 4603 4312 4604
rect 4297 4599 4298 4603
rect 4302 4599 4303 4603
rect 4307 4599 4308 4603
rect 4293 4598 4312 4599
rect 4297 4594 4298 4598
rect 4302 4594 4303 4598
rect 4307 4594 4308 4598
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4336 4624 4337 4628
rect 4322 4623 4341 4624
rect 4326 4619 4327 4623
rect 4331 4619 4332 4623
rect 4336 4619 4337 4623
rect 4322 4618 4341 4619
rect 4326 4614 4327 4618
rect 4331 4614 4332 4618
rect 4336 4614 4337 4618
rect 4322 4613 4341 4614
rect 4326 4609 4327 4613
rect 4331 4609 4332 4613
rect 4336 4609 4337 4613
rect 4322 4608 4341 4609
rect 4326 4604 4327 4608
rect 4331 4604 4332 4608
rect 4336 4604 4337 4608
rect 4322 4603 4341 4604
rect 4326 4599 4327 4603
rect 4331 4599 4332 4603
rect 4336 4599 4337 4603
rect 4322 4598 4341 4599
rect 4326 4594 4327 4598
rect 4331 4594 4332 4598
rect 4336 4594 4337 4598
rect 4355 4624 4356 4628
rect 4360 4624 4361 4628
rect 4365 4624 4366 4628
rect 4351 4623 4370 4624
rect 4355 4619 4356 4623
rect 4360 4619 4361 4623
rect 4365 4619 4366 4623
rect 4351 4618 4370 4619
rect 4355 4614 4356 4618
rect 4360 4614 4361 4618
rect 4365 4614 4366 4618
rect 4351 4613 4370 4614
rect 4355 4609 4356 4613
rect 4360 4609 4361 4613
rect 4365 4609 4366 4613
rect 4351 4608 4370 4609
rect 4355 4604 4356 4608
rect 4360 4604 4361 4608
rect 4365 4604 4366 4608
rect 4351 4603 4370 4604
rect 4355 4599 4356 4603
rect 4360 4599 4361 4603
rect 4365 4599 4366 4603
rect 4351 4598 4370 4599
rect 4355 4594 4356 4598
rect 4360 4594 4361 4598
rect 4365 4594 4366 4598
rect 4239 4578 4240 4582
rect 4244 4578 4245 4582
rect 4249 4578 4250 4582
rect 4235 4577 4254 4578
rect 4239 4573 4240 4577
rect 4244 4573 4245 4577
rect 4249 4573 4250 4577
rect 4235 4572 4254 4573
rect 4239 4568 4240 4572
rect 4244 4568 4245 4572
rect 4249 4568 4250 4572
rect 4235 4567 4254 4568
rect 4239 4563 4240 4567
rect 4244 4563 4245 4567
rect 4249 4563 4250 4567
rect 4235 4562 4254 4563
rect 4239 4558 4240 4562
rect 4244 4558 4245 4562
rect 4249 4558 4250 4562
rect 4235 4557 4254 4558
rect 4239 4553 4240 4557
rect 4244 4553 4245 4557
rect 4249 4553 4250 4557
rect 4235 4552 4254 4553
rect 4239 4548 4240 4552
rect 4244 4548 4245 4552
rect 4249 4548 4250 4552
rect 4268 4578 4269 4582
rect 4273 4578 4274 4582
rect 4278 4578 4279 4582
rect 4264 4577 4283 4578
rect 4268 4573 4269 4577
rect 4273 4573 4274 4577
rect 4278 4573 4279 4577
rect 4264 4572 4283 4573
rect 4268 4568 4269 4572
rect 4273 4568 4274 4572
rect 4278 4568 4279 4572
rect 4264 4567 4283 4568
rect 4268 4563 4269 4567
rect 4273 4563 4274 4567
rect 4278 4563 4279 4567
rect 4264 4562 4283 4563
rect 4268 4558 4269 4562
rect 4273 4558 4274 4562
rect 4278 4558 4279 4562
rect 4264 4557 4283 4558
rect 4268 4553 4269 4557
rect 4273 4553 4274 4557
rect 4278 4553 4279 4557
rect 4264 4552 4283 4553
rect 4268 4548 4269 4552
rect 4273 4548 4274 4552
rect 4278 4548 4279 4552
rect 4297 4578 4298 4582
rect 4302 4578 4303 4582
rect 4307 4578 4308 4582
rect 4293 4577 4312 4578
rect 4297 4573 4298 4577
rect 4302 4573 4303 4577
rect 4307 4573 4308 4577
rect 4293 4572 4312 4573
rect 4297 4568 4298 4572
rect 4302 4568 4303 4572
rect 4307 4568 4308 4572
rect 4293 4567 4312 4568
rect 4297 4563 4298 4567
rect 4302 4563 4303 4567
rect 4307 4563 4308 4567
rect 4293 4562 4312 4563
rect 4297 4558 4298 4562
rect 4302 4558 4303 4562
rect 4307 4558 4308 4562
rect 4293 4557 4312 4558
rect 4297 4553 4298 4557
rect 4302 4553 4303 4557
rect 4307 4553 4308 4557
rect 4293 4552 4312 4553
rect 4297 4548 4298 4552
rect 4302 4548 4303 4552
rect 4307 4548 4308 4552
rect 4326 4578 4327 4582
rect 4331 4578 4332 4582
rect 4336 4578 4337 4582
rect 4322 4577 4341 4578
rect 4326 4573 4327 4577
rect 4331 4573 4332 4577
rect 4336 4573 4337 4577
rect 4322 4572 4341 4573
rect 4326 4568 4327 4572
rect 4331 4568 4332 4572
rect 4336 4568 4337 4572
rect 4322 4567 4341 4568
rect 4326 4563 4327 4567
rect 4331 4563 4332 4567
rect 4336 4563 4337 4567
rect 4322 4562 4341 4563
rect 4326 4558 4327 4562
rect 4331 4558 4332 4562
rect 4336 4558 4337 4562
rect 4322 4557 4341 4558
rect 4326 4553 4327 4557
rect 4331 4553 4332 4557
rect 4336 4553 4337 4557
rect 4322 4552 4341 4553
rect 4326 4548 4327 4552
rect 4331 4548 4332 4552
rect 4336 4548 4337 4552
rect 4355 4578 4356 4582
rect 4360 4578 4361 4582
rect 4365 4578 4366 4582
rect 4351 4577 4370 4578
rect 4355 4573 4356 4577
rect 4360 4573 4361 4577
rect 4365 4573 4366 4577
rect 4351 4572 4370 4573
rect 4355 4568 4356 4572
rect 4360 4568 4361 4572
rect 4365 4568 4366 4572
rect 4351 4567 4370 4568
rect 4355 4563 4356 4567
rect 4360 4563 4361 4567
rect 4365 4563 4366 4567
rect 4351 4562 4370 4563
rect 4355 4558 4356 4562
rect 4360 4558 4361 4562
rect 4365 4558 4366 4562
rect 4351 4557 4370 4558
rect 4355 4553 4356 4557
rect 4360 4553 4361 4557
rect 4365 4553 4366 4557
rect 4351 4552 4370 4553
rect 4355 4548 4356 4552
rect 4360 4548 4361 4552
rect 4365 4548 4366 4552
rect 4579 4528 5054 4966
rect 3718 4318 3731 4321
rect 3615 4317 3731 4318
rect 3615 4313 3630 4317
rect 3634 4313 3637 4317
rect 3641 4313 3644 4317
rect 3648 4313 3651 4317
rect 3655 4313 3658 4317
rect 3662 4313 3665 4317
rect 3669 4313 3672 4317
rect 3676 4313 3679 4317
rect 3683 4313 3686 4317
rect 3690 4313 3693 4317
rect 3697 4313 3700 4317
rect 3704 4313 3707 4317
rect 3711 4313 3714 4317
rect 3718 4313 3731 4317
rect 3615 4311 3731 4313
rect 3924 4311 4040 4321
rect 1133 4301 1269 4311
rect 1442 4301 1578 4311
rect 1751 4301 1887 4311
rect 2060 4301 2196 4311
rect 2369 4301 2505 4311
rect 2678 4301 2814 4311
rect 2987 4301 3123 4311
rect 3296 4301 3432 4311
rect 3605 4301 3741 4311
rect 3914 4301 4050 4311
rect 1123 4291 1279 4301
rect 1432 4291 1588 4301
rect 1741 4291 1897 4301
rect 2050 4291 2206 4301
rect 2359 4291 2515 4301
rect 2668 4291 2824 4301
rect 2977 4291 3133 4301
rect 3286 4291 3442 4301
rect 3595 4291 3751 4301
rect 3904 4291 4060 4301
rect 1113 4281 1289 4291
rect 1422 4281 1598 4291
rect 1731 4281 1907 4291
rect 2040 4281 2216 4291
rect 2349 4281 2525 4291
rect 2658 4281 2834 4291
rect 2967 4281 3143 4291
rect 3276 4281 3452 4291
rect 3585 4281 3761 4291
rect 3894 4281 4070 4291
rect 1071 4278 1331 4281
rect 1071 4024 1074 4278
rect 1328 4024 1331 4278
rect 1071 4021 1331 4024
rect 1380 4278 1640 4281
rect 1380 4024 1383 4278
rect 1452 4097 1564 4211
rect 1637 4024 1640 4278
rect 1380 4021 1640 4024
rect 1689 4278 1949 4281
rect 1689 4024 1692 4278
rect 1776 4107 1854 4196
rect 1946 4024 1949 4278
rect 1689 4021 1949 4024
rect 1998 4278 2258 4281
rect 1998 4024 2001 4278
rect 2090 4115 2168 4204
rect 2255 4024 2258 4278
rect 1998 4021 2258 4024
rect 2307 4278 2567 4281
rect 2307 4024 2310 4278
rect 2394 4105 2472 4194
rect 2564 4024 2567 4278
rect 2307 4021 2567 4024
rect 2616 4278 2876 4281
rect 2616 4024 2619 4278
rect 2705 4107 2783 4196
rect 2873 4024 2876 4278
rect 2616 4021 2876 4024
rect 2925 4278 3185 4281
rect 2925 4024 2928 4278
rect 3022 4107 3100 4196
rect 3182 4024 3185 4278
rect 2925 4021 3185 4024
rect 3234 4278 3494 4281
rect 3234 4024 3237 4278
rect 3329 4112 3407 4201
rect 3491 4024 3494 4278
rect 3234 4021 3494 4024
rect 3543 4278 3803 4281
rect 3543 4024 3546 4278
rect 3626 4091 3710 4176
rect 3800 4024 3803 4278
rect 3543 4021 3803 4024
rect 3852 4278 4112 4281
rect 3852 4024 3855 4278
rect 4109 4024 4112 4278
rect 4148 4034 5054 4528
rect 3852 4021 4112 4024
<< m2contact >>
rect 1454 9997 1458 10001
rect 1461 9997 1465 10001
rect 1468 9997 1472 10001
rect 1475 9997 1479 10001
rect 1482 9997 1486 10001
rect 1489 9997 1493 10001
rect 1496 9997 1500 10001
rect 1503 9997 1507 10001
rect 1510 9997 1514 10001
rect 1517 9997 1521 10001
rect 1524 9997 1528 10001
rect 1531 9997 1535 10001
rect 1538 9997 1542 10001
rect 802 9757 806 9761
rect 807 9757 811 9761
rect 812 9757 816 9761
rect 817 9757 821 9761
rect 802 9747 806 9751
rect 807 9747 811 9751
rect 812 9747 816 9751
rect 817 9747 821 9751
rect 802 9737 806 9741
rect 807 9737 811 9741
rect 812 9737 816 9741
rect 817 9737 821 9741
rect 831 9757 835 9761
rect 836 9757 840 9761
rect 841 9757 845 9761
rect 846 9757 850 9761
rect 831 9747 835 9751
rect 836 9747 840 9751
rect 841 9747 845 9751
rect 846 9747 850 9751
rect 831 9737 835 9741
rect 836 9737 840 9741
rect 841 9737 845 9741
rect 846 9737 850 9741
rect 860 9757 864 9761
rect 865 9757 869 9761
rect 870 9757 874 9761
rect 875 9757 879 9761
rect 860 9747 864 9751
rect 865 9747 869 9751
rect 870 9747 874 9751
rect 875 9747 879 9751
rect 860 9737 864 9741
rect 865 9737 869 9741
rect 870 9737 874 9741
rect 875 9737 879 9741
rect 889 9757 893 9761
rect 894 9757 898 9761
rect 899 9757 903 9761
rect 904 9757 908 9761
rect 889 9747 893 9751
rect 894 9747 898 9751
rect 899 9747 903 9751
rect 904 9747 908 9751
rect 889 9737 893 9741
rect 894 9737 898 9741
rect 899 9737 903 9741
rect 904 9737 908 9741
rect 918 9757 922 9761
rect 923 9757 927 9761
rect 928 9757 932 9761
rect 933 9757 937 9761
rect 918 9747 922 9751
rect 923 9747 927 9751
rect 928 9747 932 9751
rect 933 9747 937 9751
rect 918 9737 922 9741
rect 923 9737 927 9741
rect 928 9737 932 9741
rect 933 9737 937 9741
rect 802 9711 806 9715
rect 807 9711 811 9715
rect 812 9711 816 9715
rect 817 9711 821 9715
rect 802 9701 806 9705
rect 807 9701 811 9705
rect 812 9701 816 9705
rect 817 9701 821 9705
rect 802 9691 806 9695
rect 807 9691 811 9695
rect 812 9691 816 9695
rect 817 9691 821 9695
rect 831 9711 835 9715
rect 836 9711 840 9715
rect 841 9711 845 9715
rect 846 9711 850 9715
rect 831 9701 835 9705
rect 836 9701 840 9705
rect 841 9701 845 9705
rect 846 9701 850 9705
rect 831 9691 835 9695
rect 836 9691 840 9695
rect 841 9691 845 9695
rect 846 9691 850 9695
rect 860 9711 864 9715
rect 865 9711 869 9715
rect 870 9711 874 9715
rect 875 9711 879 9715
rect 860 9701 864 9705
rect 865 9701 869 9705
rect 870 9701 874 9705
rect 875 9701 879 9705
rect 860 9691 864 9695
rect 865 9691 869 9695
rect 870 9691 874 9695
rect 875 9691 879 9695
rect 889 9711 893 9715
rect 894 9711 898 9715
rect 899 9711 903 9715
rect 904 9711 908 9715
rect 889 9701 893 9705
rect 894 9701 898 9705
rect 899 9701 903 9705
rect 904 9701 908 9705
rect 889 9691 893 9695
rect 894 9691 898 9695
rect 899 9691 903 9695
rect 904 9691 908 9695
rect 918 9711 922 9715
rect 923 9711 927 9715
rect 928 9711 932 9715
rect 933 9711 937 9715
rect 918 9701 922 9705
rect 923 9701 927 9705
rect 928 9701 932 9705
rect 933 9701 937 9705
rect 918 9691 922 9695
rect 923 9691 927 9695
rect 928 9691 932 9695
rect 933 9691 937 9695
rect 618 9618 622 9622
rect 628 9618 632 9622
rect 638 9618 642 9622
rect 618 9613 622 9617
rect 628 9613 632 9617
rect 638 9613 642 9617
rect 618 9608 622 9612
rect 628 9608 632 9612
rect 638 9608 642 9612
rect 618 9603 622 9607
rect 628 9603 632 9607
rect 638 9603 642 9607
rect 664 9618 668 9622
rect 674 9618 678 9622
rect 684 9618 688 9622
rect 664 9613 668 9617
rect 674 9613 678 9617
rect 684 9613 688 9617
rect 664 9608 668 9612
rect 674 9608 678 9612
rect 684 9608 688 9612
rect 1454 9992 1458 9996
rect 1461 9992 1465 9996
rect 1468 9992 1472 9996
rect 1475 9992 1479 9996
rect 1482 9992 1486 9996
rect 1489 9992 1493 9996
rect 1496 9992 1500 9996
rect 1503 9992 1507 9996
rect 1510 9992 1514 9996
rect 1517 9992 1521 9996
rect 1524 9992 1528 9996
rect 1531 9992 1535 9996
rect 1538 9992 1542 9996
rect 1763 9997 1767 10001
rect 1770 9997 1774 10001
rect 1777 9997 1781 10001
rect 1784 9997 1788 10001
rect 1791 9997 1795 10001
rect 1798 9997 1802 10001
rect 1805 9997 1809 10001
rect 1812 9997 1816 10001
rect 1819 9997 1823 10001
rect 1826 9997 1830 10001
rect 1833 9997 1837 10001
rect 1840 9997 1844 10001
rect 1847 9997 1851 10001
rect 1454 9987 1458 9991
rect 1461 9987 1465 9991
rect 1468 9987 1472 9991
rect 1475 9987 1479 9991
rect 1482 9987 1486 9991
rect 1489 9987 1493 9991
rect 1496 9987 1500 9991
rect 1503 9987 1507 9991
rect 1510 9987 1514 9991
rect 1517 9987 1521 9991
rect 1524 9987 1528 9991
rect 1531 9987 1535 9991
rect 1538 9987 1542 9991
rect 1454 9982 1458 9986
rect 1461 9982 1465 9986
rect 1468 9982 1472 9986
rect 1475 9982 1479 9986
rect 1482 9982 1486 9986
rect 1489 9982 1493 9986
rect 1496 9982 1500 9986
rect 1503 9982 1507 9986
rect 1510 9982 1514 9986
rect 1517 9982 1521 9986
rect 1524 9982 1528 9986
rect 1531 9982 1535 9986
rect 1538 9982 1542 9986
rect 1763 9992 1767 9996
rect 1770 9992 1774 9996
rect 1777 9992 1781 9996
rect 1784 9992 1788 9996
rect 1791 9992 1795 9996
rect 1798 9992 1802 9996
rect 1805 9992 1809 9996
rect 1812 9992 1816 9996
rect 1819 9992 1823 9996
rect 1826 9992 1830 9996
rect 1833 9992 1837 9996
rect 1840 9992 1844 9996
rect 1847 9992 1851 9996
rect 2072 9997 2076 10001
rect 2079 9997 2083 10001
rect 2086 9997 2090 10001
rect 2093 9997 2097 10001
rect 2100 9997 2104 10001
rect 2107 9997 2111 10001
rect 2114 9997 2118 10001
rect 2121 9997 2125 10001
rect 2128 9997 2132 10001
rect 2135 9997 2139 10001
rect 2142 9997 2146 10001
rect 2149 9997 2153 10001
rect 2156 9997 2160 10001
rect 1763 9987 1767 9991
rect 1770 9987 1774 9991
rect 1777 9987 1781 9991
rect 1784 9987 1788 9991
rect 1791 9987 1795 9991
rect 1798 9987 1802 9991
rect 1805 9987 1809 9991
rect 1812 9987 1816 9991
rect 1819 9987 1823 9991
rect 1826 9987 1830 9991
rect 1833 9987 1837 9991
rect 1840 9987 1844 9991
rect 1847 9987 1851 9991
rect 1763 9982 1767 9986
rect 1770 9982 1774 9986
rect 1777 9982 1781 9986
rect 1784 9982 1788 9986
rect 1791 9982 1795 9986
rect 1798 9982 1802 9986
rect 1805 9982 1809 9986
rect 1812 9982 1816 9986
rect 1819 9982 1823 9986
rect 1826 9982 1830 9986
rect 1833 9982 1837 9986
rect 1840 9982 1844 9986
rect 1847 9982 1851 9986
rect 2072 9992 2076 9996
rect 2079 9992 2083 9996
rect 2086 9992 2090 9996
rect 2093 9992 2097 9996
rect 2100 9992 2104 9996
rect 2107 9992 2111 9996
rect 2114 9992 2118 9996
rect 2121 9992 2125 9996
rect 2128 9992 2132 9996
rect 2135 9992 2139 9996
rect 2142 9992 2146 9996
rect 2149 9992 2153 9996
rect 2156 9992 2160 9996
rect 2381 9997 2385 10001
rect 2388 9997 2392 10001
rect 2395 9997 2399 10001
rect 2402 9997 2406 10001
rect 2409 9997 2413 10001
rect 2416 9997 2420 10001
rect 2423 9997 2427 10001
rect 2430 9997 2434 10001
rect 2437 9997 2441 10001
rect 2444 9997 2448 10001
rect 2451 9997 2455 10001
rect 2458 9997 2462 10001
rect 2465 9997 2469 10001
rect 2072 9987 2076 9991
rect 2079 9987 2083 9991
rect 2086 9987 2090 9991
rect 2093 9987 2097 9991
rect 2100 9987 2104 9991
rect 2107 9987 2111 9991
rect 2114 9987 2118 9991
rect 2121 9987 2125 9991
rect 2128 9987 2132 9991
rect 2135 9987 2139 9991
rect 2142 9987 2146 9991
rect 2149 9987 2153 9991
rect 2156 9987 2160 9991
rect 2072 9982 2076 9986
rect 2079 9982 2083 9986
rect 2086 9982 2090 9986
rect 2093 9982 2097 9986
rect 2100 9982 2104 9986
rect 2107 9982 2111 9986
rect 2114 9982 2118 9986
rect 2121 9982 2125 9986
rect 2128 9982 2132 9986
rect 2135 9982 2139 9986
rect 2142 9982 2146 9986
rect 2149 9982 2153 9986
rect 2156 9982 2160 9986
rect 2381 9992 2385 9996
rect 2388 9992 2392 9996
rect 2395 9992 2399 9996
rect 2402 9992 2406 9996
rect 2409 9992 2413 9996
rect 2416 9992 2420 9996
rect 2423 9992 2427 9996
rect 2430 9992 2434 9996
rect 2437 9992 2441 9996
rect 2444 9992 2448 9996
rect 2451 9992 2455 9996
rect 2458 9992 2462 9996
rect 2465 9992 2469 9996
rect 2690 9997 2694 10001
rect 2697 9997 2701 10001
rect 2704 9997 2708 10001
rect 2711 9997 2715 10001
rect 2718 9997 2722 10001
rect 2725 9997 2729 10001
rect 2732 9997 2736 10001
rect 2739 9997 2743 10001
rect 2746 9997 2750 10001
rect 2753 9997 2757 10001
rect 2760 9997 2764 10001
rect 2767 9997 2771 10001
rect 2774 9997 2778 10001
rect 2381 9987 2385 9991
rect 2388 9987 2392 9991
rect 2395 9987 2399 9991
rect 2402 9987 2406 9991
rect 2409 9987 2413 9991
rect 2416 9987 2420 9991
rect 2423 9987 2427 9991
rect 2430 9987 2434 9991
rect 2437 9987 2441 9991
rect 2444 9987 2448 9991
rect 2451 9987 2455 9991
rect 2458 9987 2462 9991
rect 2465 9987 2469 9991
rect 2381 9982 2385 9986
rect 2388 9982 2392 9986
rect 2395 9982 2399 9986
rect 2402 9982 2406 9986
rect 2409 9982 2413 9986
rect 2416 9982 2420 9986
rect 2423 9982 2427 9986
rect 2430 9982 2434 9986
rect 2437 9982 2441 9986
rect 2444 9982 2448 9986
rect 2451 9982 2455 9986
rect 2458 9982 2462 9986
rect 2465 9982 2469 9986
rect 2690 9992 2694 9996
rect 2697 9992 2701 9996
rect 2704 9992 2708 9996
rect 2711 9992 2715 9996
rect 2718 9992 2722 9996
rect 2725 9992 2729 9996
rect 2732 9992 2736 9996
rect 2739 9992 2743 9996
rect 2746 9992 2750 9996
rect 2753 9992 2757 9996
rect 2760 9992 2764 9996
rect 2767 9992 2771 9996
rect 2774 9992 2778 9996
rect 2999 9997 3003 10001
rect 3006 9997 3010 10001
rect 3013 9997 3017 10001
rect 3020 9997 3024 10001
rect 3027 9997 3031 10001
rect 3034 9997 3038 10001
rect 3041 9997 3045 10001
rect 3048 9997 3052 10001
rect 3055 9997 3059 10001
rect 3062 9997 3066 10001
rect 3069 9997 3073 10001
rect 3076 9997 3080 10001
rect 3083 9997 3087 10001
rect 2690 9987 2694 9991
rect 2697 9987 2701 9991
rect 2704 9987 2708 9991
rect 2711 9987 2715 9991
rect 2718 9987 2722 9991
rect 2725 9987 2729 9991
rect 2732 9987 2736 9991
rect 2739 9987 2743 9991
rect 2746 9987 2750 9991
rect 2753 9987 2757 9991
rect 2760 9987 2764 9991
rect 2767 9987 2771 9991
rect 2774 9987 2778 9991
rect 2690 9982 2694 9986
rect 2697 9982 2701 9986
rect 2704 9982 2708 9986
rect 2711 9982 2715 9986
rect 2718 9982 2722 9986
rect 2725 9982 2729 9986
rect 2732 9982 2736 9986
rect 2739 9982 2743 9986
rect 2746 9982 2750 9986
rect 2753 9982 2757 9986
rect 2760 9982 2764 9986
rect 2767 9982 2771 9986
rect 2774 9982 2778 9986
rect 2999 9992 3003 9996
rect 3006 9992 3010 9996
rect 3013 9992 3017 9996
rect 3020 9992 3024 9996
rect 3027 9992 3031 9996
rect 3034 9992 3038 9996
rect 3041 9992 3045 9996
rect 3048 9992 3052 9996
rect 3055 9992 3059 9996
rect 3062 9992 3066 9996
rect 3069 9992 3073 9996
rect 3076 9992 3080 9996
rect 3083 9992 3087 9996
rect 3308 9997 3312 10001
rect 3315 9997 3319 10001
rect 3322 9997 3326 10001
rect 3329 9997 3333 10001
rect 3336 9997 3340 10001
rect 3343 9997 3347 10001
rect 3350 9997 3354 10001
rect 3357 9997 3361 10001
rect 3364 9997 3368 10001
rect 3371 9997 3375 10001
rect 3378 9997 3382 10001
rect 3385 9997 3389 10001
rect 3392 9997 3396 10001
rect 2999 9987 3003 9991
rect 3006 9987 3010 9991
rect 3013 9987 3017 9991
rect 3020 9987 3024 9991
rect 3027 9987 3031 9991
rect 3034 9987 3038 9991
rect 3041 9987 3045 9991
rect 3048 9987 3052 9991
rect 3055 9987 3059 9991
rect 3062 9987 3066 9991
rect 3069 9987 3073 9991
rect 3076 9987 3080 9991
rect 3083 9987 3087 9991
rect 2999 9982 3003 9986
rect 3006 9982 3010 9986
rect 3013 9982 3017 9986
rect 3020 9982 3024 9986
rect 3027 9982 3031 9986
rect 3034 9982 3038 9986
rect 3041 9982 3045 9986
rect 3048 9982 3052 9986
rect 3055 9982 3059 9986
rect 3062 9982 3066 9986
rect 3069 9982 3073 9986
rect 3076 9982 3080 9986
rect 3083 9982 3087 9986
rect 3308 9992 3312 9996
rect 3315 9992 3319 9996
rect 3322 9992 3326 9996
rect 3329 9992 3333 9996
rect 3336 9992 3340 9996
rect 3343 9992 3347 9996
rect 3350 9992 3354 9996
rect 3357 9992 3361 9996
rect 3364 9992 3368 9996
rect 3371 9992 3375 9996
rect 3378 9992 3382 9996
rect 3385 9992 3389 9996
rect 3392 9992 3396 9996
rect 3617 9997 3621 10001
rect 3624 9997 3628 10001
rect 3631 9997 3635 10001
rect 3638 9997 3642 10001
rect 3645 9997 3649 10001
rect 3652 9997 3656 10001
rect 3659 9997 3663 10001
rect 3666 9997 3670 10001
rect 3673 9997 3677 10001
rect 3680 9997 3684 10001
rect 3687 9997 3691 10001
rect 3694 9997 3698 10001
rect 3701 9997 3705 10001
rect 3308 9987 3312 9991
rect 3315 9987 3319 9991
rect 3322 9987 3326 9991
rect 3329 9987 3333 9991
rect 3336 9987 3340 9991
rect 3343 9987 3347 9991
rect 3350 9987 3354 9991
rect 3357 9987 3361 9991
rect 3364 9987 3368 9991
rect 3371 9987 3375 9991
rect 3378 9987 3382 9991
rect 3385 9987 3389 9991
rect 3392 9987 3396 9991
rect 3308 9982 3312 9986
rect 3315 9982 3319 9986
rect 3322 9982 3326 9986
rect 3329 9982 3333 9986
rect 3336 9982 3340 9986
rect 3343 9982 3347 9986
rect 3350 9982 3354 9986
rect 3357 9982 3361 9986
rect 3364 9982 3368 9986
rect 3371 9982 3375 9986
rect 3378 9982 3382 9986
rect 3385 9982 3389 9986
rect 3392 9982 3396 9986
rect 3617 9992 3621 9996
rect 3624 9992 3628 9996
rect 3631 9992 3635 9996
rect 3638 9992 3642 9996
rect 3645 9992 3649 9996
rect 3652 9992 3656 9996
rect 3659 9992 3663 9996
rect 3666 9992 3670 9996
rect 3673 9992 3677 9996
rect 3680 9992 3684 9996
rect 3687 9992 3691 9996
rect 3694 9992 3698 9996
rect 3701 9992 3705 9996
rect 3926 9997 3930 10001
rect 3933 9997 3937 10001
rect 3940 9997 3944 10001
rect 3947 9997 3951 10001
rect 3954 9997 3958 10001
rect 3961 9997 3965 10001
rect 3968 9997 3972 10001
rect 3975 9997 3979 10001
rect 3982 9997 3986 10001
rect 3989 9997 3993 10001
rect 3996 9997 4000 10001
rect 4003 9997 4007 10001
rect 4010 9997 4014 10001
rect 3617 9987 3621 9991
rect 3624 9987 3628 9991
rect 3631 9987 3635 9991
rect 3638 9987 3642 9991
rect 3645 9987 3649 9991
rect 3652 9987 3656 9991
rect 3659 9987 3663 9991
rect 3666 9987 3670 9991
rect 3673 9987 3677 9991
rect 3680 9987 3684 9991
rect 3687 9987 3691 9991
rect 3694 9987 3698 9991
rect 3701 9987 3705 9991
rect 3617 9982 3621 9986
rect 3624 9982 3628 9986
rect 3631 9982 3635 9986
rect 3638 9982 3642 9986
rect 3645 9982 3649 9986
rect 3652 9982 3656 9986
rect 3659 9982 3663 9986
rect 3666 9982 3670 9986
rect 3673 9982 3677 9986
rect 3680 9982 3684 9986
rect 3687 9982 3691 9986
rect 3694 9982 3698 9986
rect 3701 9982 3705 9986
rect 3926 9992 3930 9996
rect 3933 9992 3937 9996
rect 3940 9992 3944 9996
rect 3947 9992 3951 9996
rect 3954 9992 3958 9996
rect 3961 9992 3965 9996
rect 3968 9992 3972 9996
rect 3975 9992 3979 9996
rect 3982 9992 3986 9996
rect 3989 9992 3993 9996
rect 3996 9992 4000 9996
rect 4003 9992 4007 9996
rect 4010 9992 4014 9996
rect 3926 9987 3930 9991
rect 3933 9987 3937 9991
rect 3940 9987 3944 9991
rect 3947 9987 3951 9991
rect 3954 9987 3958 9991
rect 3961 9987 3965 9991
rect 3968 9987 3972 9991
rect 3975 9987 3979 9991
rect 3982 9987 3986 9991
rect 3989 9987 3993 9991
rect 3996 9987 4000 9991
rect 4003 9987 4007 9991
rect 4010 9987 4014 9991
rect 3926 9982 3930 9986
rect 3933 9982 3937 9986
rect 3940 9982 3944 9986
rect 3947 9982 3951 9986
rect 3954 9982 3958 9986
rect 3961 9982 3965 9986
rect 3968 9982 3972 9986
rect 3975 9982 3979 9986
rect 3982 9982 3986 9986
rect 3989 9982 3993 9986
rect 3996 9982 4000 9986
rect 4003 9982 4007 9986
rect 4010 9982 4014 9986
rect 1397 9949 1401 9953
rect 1407 9949 1411 9953
rect 1417 9949 1421 9953
rect 1427 9949 1431 9953
rect 1437 9949 1441 9953
rect 1402 9944 1406 9948
rect 1412 9944 1416 9948
rect 1422 9944 1426 9948
rect 1432 9944 1436 9948
rect 1397 9939 1401 9943
rect 1407 9939 1411 9943
rect 1417 9939 1421 9943
rect 1427 9939 1431 9943
rect 1437 9939 1441 9943
rect 1402 9934 1406 9938
rect 1412 9934 1416 9938
rect 1422 9934 1426 9938
rect 1432 9934 1436 9938
rect 1397 9929 1401 9933
rect 1407 9929 1411 9933
rect 1417 9929 1421 9933
rect 1427 9929 1431 9933
rect 1437 9929 1441 9933
rect 1402 9924 1406 9928
rect 1412 9924 1416 9928
rect 1422 9924 1426 9928
rect 1432 9924 1436 9928
rect 1397 9919 1401 9923
rect 1407 9919 1411 9923
rect 1417 9919 1421 9923
rect 1427 9919 1431 9923
rect 1437 9919 1441 9923
rect 1402 9914 1406 9918
rect 1412 9914 1416 9918
rect 1422 9914 1426 9918
rect 1432 9914 1436 9918
rect 1397 9909 1401 9913
rect 1407 9909 1411 9913
rect 1417 9909 1421 9913
rect 1427 9909 1431 9913
rect 1437 9909 1441 9913
rect 1402 9904 1406 9908
rect 1412 9904 1416 9908
rect 1422 9904 1426 9908
rect 1432 9904 1436 9908
rect 1397 9899 1401 9903
rect 1407 9899 1411 9903
rect 1417 9899 1421 9903
rect 1427 9899 1431 9903
rect 1437 9899 1441 9903
rect 1402 9894 1406 9898
rect 1412 9894 1416 9898
rect 1422 9894 1426 9898
rect 1432 9894 1436 9898
rect 1397 9889 1401 9893
rect 1407 9889 1411 9893
rect 1417 9889 1421 9893
rect 1427 9889 1431 9893
rect 1437 9889 1441 9893
rect 1402 9884 1406 9888
rect 1412 9884 1416 9888
rect 1422 9884 1426 9888
rect 1432 9884 1436 9888
rect 1397 9879 1401 9883
rect 1407 9879 1411 9883
rect 1417 9879 1421 9883
rect 1427 9879 1431 9883
rect 1437 9879 1441 9883
rect 1402 9874 1406 9878
rect 1412 9874 1416 9878
rect 1422 9874 1426 9878
rect 1432 9874 1436 9878
rect 1397 9869 1401 9873
rect 1407 9869 1411 9873
rect 1417 9869 1421 9873
rect 1427 9869 1431 9873
rect 1437 9869 1441 9873
rect 1402 9864 1406 9868
rect 1412 9864 1416 9868
rect 1422 9864 1426 9868
rect 1432 9864 1436 9868
rect 1385 9848 1389 9852
rect 1392 9848 1396 9852
rect 1397 9848 1401 9852
rect 1402 9848 1406 9852
rect 1407 9848 1411 9852
rect 1412 9848 1416 9852
rect 1417 9848 1421 9852
rect 1422 9848 1426 9852
rect 1427 9848 1431 9852
rect 1432 9848 1436 9852
rect 1437 9848 1441 9852
rect 1442 9848 1446 9852
rect 1449 9848 1453 9852
rect 1364 9796 1368 9800
rect 1369 9796 1373 9800
rect 1364 9791 1368 9795
rect 1369 9791 1373 9795
rect 1364 9786 1368 9790
rect 1369 9786 1373 9790
rect 1364 9781 1368 9785
rect 1369 9781 1373 9785
rect 1364 9776 1368 9780
rect 1369 9776 1373 9780
rect 1364 9771 1368 9775
rect 1369 9771 1373 9775
rect 1364 9766 1368 9770
rect 1369 9766 1373 9770
rect 1319 9757 1323 9761
rect 1324 9757 1328 9761
rect 1329 9757 1333 9761
rect 1334 9757 1338 9761
rect 1319 9747 1323 9751
rect 1324 9747 1328 9751
rect 1329 9747 1333 9751
rect 1334 9747 1338 9751
rect 1319 9737 1323 9741
rect 1324 9737 1328 9741
rect 1329 9737 1333 9741
rect 1334 9737 1338 9741
rect 1364 9761 1368 9765
rect 1369 9761 1373 9765
rect 1364 9756 1368 9760
rect 1369 9756 1373 9760
rect 1364 9751 1368 9755
rect 1369 9751 1373 9755
rect 1364 9746 1368 9750
rect 1369 9746 1373 9750
rect 1364 9741 1368 9745
rect 1369 9741 1373 9745
rect 1364 9736 1368 9740
rect 1369 9736 1373 9740
rect 1319 9711 1323 9715
rect 1324 9711 1328 9715
rect 1329 9711 1333 9715
rect 1334 9711 1338 9715
rect 1319 9701 1323 9705
rect 1324 9701 1328 9705
rect 1329 9701 1333 9705
rect 1334 9701 1338 9705
rect 1319 9691 1323 9695
rect 1324 9691 1328 9695
rect 1329 9691 1333 9695
rect 1334 9691 1338 9695
rect 1557 9949 1561 9953
rect 1567 9949 1571 9953
rect 1577 9949 1581 9953
rect 1587 9949 1591 9953
rect 1597 9949 1601 9953
rect 1562 9944 1566 9948
rect 1572 9944 1576 9948
rect 1582 9944 1586 9948
rect 1592 9944 1596 9948
rect 1557 9939 1561 9943
rect 1567 9939 1571 9943
rect 1577 9939 1581 9943
rect 1587 9939 1591 9943
rect 1597 9939 1601 9943
rect 1562 9934 1566 9938
rect 1572 9934 1576 9938
rect 1582 9934 1586 9938
rect 1592 9934 1596 9938
rect 1557 9929 1561 9933
rect 1567 9929 1571 9933
rect 1577 9929 1581 9933
rect 1587 9929 1591 9933
rect 1597 9929 1601 9933
rect 1562 9924 1566 9928
rect 1572 9924 1576 9928
rect 1582 9924 1586 9928
rect 1592 9924 1596 9928
rect 1557 9919 1561 9923
rect 1567 9919 1571 9923
rect 1577 9919 1581 9923
rect 1587 9919 1591 9923
rect 1597 9919 1601 9923
rect 1562 9914 1566 9918
rect 1572 9914 1576 9918
rect 1582 9914 1586 9918
rect 1592 9914 1596 9918
rect 1557 9909 1561 9913
rect 1567 9909 1571 9913
rect 1577 9909 1581 9913
rect 1587 9909 1591 9913
rect 1597 9909 1601 9913
rect 1562 9904 1566 9908
rect 1572 9904 1576 9908
rect 1582 9904 1586 9908
rect 1592 9904 1596 9908
rect 1557 9899 1561 9903
rect 1567 9899 1571 9903
rect 1577 9899 1581 9903
rect 1587 9899 1591 9903
rect 1597 9899 1601 9903
rect 1562 9894 1566 9898
rect 1572 9894 1576 9898
rect 1582 9894 1586 9898
rect 1592 9894 1596 9898
rect 1557 9889 1561 9893
rect 1567 9889 1571 9893
rect 1577 9889 1581 9893
rect 1587 9889 1591 9893
rect 1597 9889 1601 9893
rect 1562 9884 1566 9888
rect 1572 9884 1576 9888
rect 1582 9884 1586 9888
rect 1592 9884 1596 9888
rect 1557 9879 1561 9883
rect 1567 9879 1571 9883
rect 1577 9879 1581 9883
rect 1587 9879 1591 9883
rect 1597 9879 1601 9883
rect 1562 9874 1566 9878
rect 1572 9874 1576 9878
rect 1582 9874 1586 9878
rect 1592 9874 1596 9878
rect 1557 9869 1561 9873
rect 1567 9869 1571 9873
rect 1577 9869 1581 9873
rect 1587 9869 1591 9873
rect 1597 9869 1601 9873
rect 1562 9864 1566 9868
rect 1572 9864 1576 9868
rect 1582 9864 1586 9868
rect 1592 9864 1596 9868
rect 1545 9848 1549 9852
rect 1552 9848 1556 9852
rect 1557 9848 1561 9852
rect 1562 9848 1566 9852
rect 1567 9848 1571 9852
rect 1572 9848 1576 9852
rect 1577 9848 1581 9852
rect 1582 9848 1586 9852
rect 1587 9848 1591 9852
rect 1592 9848 1596 9852
rect 1597 9848 1601 9852
rect 1602 9848 1606 9852
rect 1609 9848 1613 9852
rect 1706 9949 1710 9953
rect 1716 9949 1720 9953
rect 1726 9949 1730 9953
rect 1736 9949 1740 9953
rect 1746 9949 1750 9953
rect 1711 9944 1715 9948
rect 1721 9944 1725 9948
rect 1731 9944 1735 9948
rect 1741 9944 1745 9948
rect 1706 9939 1710 9943
rect 1716 9939 1720 9943
rect 1726 9939 1730 9943
rect 1736 9939 1740 9943
rect 1746 9939 1750 9943
rect 1711 9934 1715 9938
rect 1721 9934 1725 9938
rect 1731 9934 1735 9938
rect 1741 9934 1745 9938
rect 1706 9929 1710 9933
rect 1716 9929 1720 9933
rect 1726 9929 1730 9933
rect 1736 9929 1740 9933
rect 1746 9929 1750 9933
rect 1711 9924 1715 9928
rect 1721 9924 1725 9928
rect 1731 9924 1735 9928
rect 1741 9924 1745 9928
rect 1706 9919 1710 9923
rect 1716 9919 1720 9923
rect 1726 9919 1730 9923
rect 1736 9919 1740 9923
rect 1746 9919 1750 9923
rect 1711 9914 1715 9918
rect 1721 9914 1725 9918
rect 1731 9914 1735 9918
rect 1741 9914 1745 9918
rect 1706 9909 1710 9913
rect 1716 9909 1720 9913
rect 1726 9909 1730 9913
rect 1736 9909 1740 9913
rect 1746 9909 1750 9913
rect 1711 9904 1715 9908
rect 1721 9904 1725 9908
rect 1731 9904 1735 9908
rect 1741 9904 1745 9908
rect 1706 9899 1710 9903
rect 1716 9899 1720 9903
rect 1726 9899 1730 9903
rect 1736 9899 1740 9903
rect 1746 9899 1750 9903
rect 1711 9894 1715 9898
rect 1721 9894 1725 9898
rect 1731 9894 1735 9898
rect 1741 9894 1745 9898
rect 1706 9889 1710 9893
rect 1716 9889 1720 9893
rect 1726 9889 1730 9893
rect 1736 9889 1740 9893
rect 1746 9889 1750 9893
rect 1711 9884 1715 9888
rect 1721 9884 1725 9888
rect 1731 9884 1735 9888
rect 1741 9884 1745 9888
rect 1706 9879 1710 9883
rect 1716 9879 1720 9883
rect 1726 9879 1730 9883
rect 1736 9879 1740 9883
rect 1746 9879 1750 9883
rect 1711 9874 1715 9878
rect 1721 9874 1725 9878
rect 1731 9874 1735 9878
rect 1741 9874 1745 9878
rect 1706 9869 1710 9873
rect 1716 9869 1720 9873
rect 1726 9869 1730 9873
rect 1736 9869 1740 9873
rect 1746 9869 1750 9873
rect 1711 9864 1715 9868
rect 1721 9864 1725 9868
rect 1731 9864 1735 9868
rect 1741 9864 1745 9868
rect 1694 9848 1698 9852
rect 1701 9848 1705 9852
rect 1706 9848 1710 9852
rect 1711 9848 1715 9852
rect 1716 9848 1720 9852
rect 1721 9848 1725 9852
rect 1726 9848 1730 9852
rect 1731 9848 1735 9852
rect 1736 9848 1740 9852
rect 1741 9848 1745 9852
rect 1746 9848 1750 9852
rect 1751 9848 1755 9852
rect 1758 9848 1762 9852
rect 1866 9949 1870 9953
rect 1876 9949 1880 9953
rect 1886 9949 1890 9953
rect 1896 9949 1900 9953
rect 1906 9949 1910 9953
rect 1871 9944 1875 9948
rect 1881 9944 1885 9948
rect 1891 9944 1895 9948
rect 1901 9944 1905 9948
rect 1866 9939 1870 9943
rect 1876 9939 1880 9943
rect 1886 9939 1890 9943
rect 1896 9939 1900 9943
rect 1906 9939 1910 9943
rect 1871 9934 1875 9938
rect 1881 9934 1885 9938
rect 1891 9934 1895 9938
rect 1901 9934 1905 9938
rect 1866 9929 1870 9933
rect 1876 9929 1880 9933
rect 1886 9929 1890 9933
rect 1896 9929 1900 9933
rect 1906 9929 1910 9933
rect 1871 9924 1875 9928
rect 1881 9924 1885 9928
rect 1891 9924 1895 9928
rect 1901 9924 1905 9928
rect 1866 9919 1870 9923
rect 1876 9919 1880 9923
rect 1886 9919 1890 9923
rect 1896 9919 1900 9923
rect 1906 9919 1910 9923
rect 1871 9914 1875 9918
rect 1881 9914 1885 9918
rect 1891 9914 1895 9918
rect 1901 9914 1905 9918
rect 1866 9909 1870 9913
rect 1876 9909 1880 9913
rect 1886 9909 1890 9913
rect 1896 9909 1900 9913
rect 1906 9909 1910 9913
rect 1871 9904 1875 9908
rect 1881 9904 1885 9908
rect 1891 9904 1895 9908
rect 1901 9904 1905 9908
rect 1866 9899 1870 9903
rect 1876 9899 1880 9903
rect 1886 9899 1890 9903
rect 1896 9899 1900 9903
rect 1906 9899 1910 9903
rect 1871 9894 1875 9898
rect 1881 9894 1885 9898
rect 1891 9894 1895 9898
rect 1901 9894 1905 9898
rect 1866 9889 1870 9893
rect 1876 9889 1880 9893
rect 1886 9889 1890 9893
rect 1896 9889 1900 9893
rect 1906 9889 1910 9893
rect 1871 9884 1875 9888
rect 1881 9884 1885 9888
rect 1891 9884 1895 9888
rect 1901 9884 1905 9888
rect 1866 9879 1870 9883
rect 1876 9879 1880 9883
rect 1886 9879 1890 9883
rect 1896 9879 1900 9883
rect 1906 9879 1910 9883
rect 1871 9874 1875 9878
rect 1881 9874 1885 9878
rect 1891 9874 1895 9878
rect 1901 9874 1905 9878
rect 1866 9869 1870 9873
rect 1876 9869 1880 9873
rect 1886 9869 1890 9873
rect 1896 9869 1900 9873
rect 1906 9869 1910 9873
rect 1871 9864 1875 9868
rect 1881 9864 1885 9868
rect 1891 9864 1895 9868
rect 1901 9864 1905 9868
rect 1854 9848 1858 9852
rect 1861 9848 1865 9852
rect 1866 9848 1870 9852
rect 1871 9848 1875 9852
rect 1876 9848 1880 9852
rect 1881 9848 1885 9852
rect 1886 9848 1890 9852
rect 1891 9848 1895 9852
rect 1896 9848 1900 9852
rect 1901 9848 1905 9852
rect 1906 9848 1910 9852
rect 1911 9848 1915 9852
rect 1918 9848 1922 9852
rect 1499 9711 1503 9715
rect 1504 9711 1508 9715
rect 2015 9949 2019 9953
rect 2025 9949 2029 9953
rect 2035 9949 2039 9953
rect 2045 9949 2049 9953
rect 2055 9949 2059 9953
rect 2020 9944 2024 9948
rect 2030 9944 2034 9948
rect 2040 9944 2044 9948
rect 2050 9944 2054 9948
rect 2015 9939 2019 9943
rect 2025 9939 2029 9943
rect 2035 9939 2039 9943
rect 2045 9939 2049 9943
rect 2055 9939 2059 9943
rect 2020 9934 2024 9938
rect 2030 9934 2034 9938
rect 2040 9934 2044 9938
rect 2050 9934 2054 9938
rect 2015 9929 2019 9933
rect 2025 9929 2029 9933
rect 2035 9929 2039 9933
rect 2045 9929 2049 9933
rect 2055 9929 2059 9933
rect 2020 9924 2024 9928
rect 2030 9924 2034 9928
rect 2040 9924 2044 9928
rect 2050 9924 2054 9928
rect 2015 9919 2019 9923
rect 2025 9919 2029 9923
rect 2035 9919 2039 9923
rect 2045 9919 2049 9923
rect 2055 9919 2059 9923
rect 2020 9914 2024 9918
rect 2030 9914 2034 9918
rect 2040 9914 2044 9918
rect 2050 9914 2054 9918
rect 2015 9909 2019 9913
rect 2025 9909 2029 9913
rect 2035 9909 2039 9913
rect 2045 9909 2049 9913
rect 2055 9909 2059 9913
rect 2020 9904 2024 9908
rect 2030 9904 2034 9908
rect 2040 9904 2044 9908
rect 2050 9904 2054 9908
rect 2015 9899 2019 9903
rect 2025 9899 2029 9903
rect 2035 9899 2039 9903
rect 2045 9899 2049 9903
rect 2055 9899 2059 9903
rect 2020 9894 2024 9898
rect 2030 9894 2034 9898
rect 2040 9894 2044 9898
rect 2050 9894 2054 9898
rect 2015 9889 2019 9893
rect 2025 9889 2029 9893
rect 2035 9889 2039 9893
rect 2045 9889 2049 9893
rect 2055 9889 2059 9893
rect 2020 9884 2024 9888
rect 2030 9884 2034 9888
rect 2040 9884 2044 9888
rect 2050 9884 2054 9888
rect 2015 9879 2019 9883
rect 2025 9879 2029 9883
rect 2035 9879 2039 9883
rect 2045 9879 2049 9883
rect 2055 9879 2059 9883
rect 2020 9874 2024 9878
rect 2030 9874 2034 9878
rect 2040 9874 2044 9878
rect 2050 9874 2054 9878
rect 2015 9869 2019 9873
rect 2025 9869 2029 9873
rect 2035 9869 2039 9873
rect 2045 9869 2049 9873
rect 2055 9869 2059 9873
rect 2020 9864 2024 9868
rect 2030 9864 2034 9868
rect 2040 9864 2044 9868
rect 2050 9864 2054 9868
rect 2003 9848 2007 9852
rect 2010 9848 2014 9852
rect 2015 9848 2019 9852
rect 2020 9848 2024 9852
rect 2025 9848 2029 9852
rect 2030 9848 2034 9852
rect 2035 9848 2039 9852
rect 2040 9848 2044 9852
rect 2045 9848 2049 9852
rect 2050 9848 2054 9852
rect 2055 9848 2059 9852
rect 2060 9848 2064 9852
rect 2067 9848 2071 9852
rect 2175 9949 2179 9953
rect 2185 9949 2189 9953
rect 2195 9949 2199 9953
rect 2205 9949 2209 9953
rect 2215 9949 2219 9953
rect 2180 9944 2184 9948
rect 2190 9944 2194 9948
rect 2200 9944 2204 9948
rect 2210 9944 2214 9948
rect 2175 9939 2179 9943
rect 2185 9939 2189 9943
rect 2195 9939 2199 9943
rect 2205 9939 2209 9943
rect 2215 9939 2219 9943
rect 2180 9934 2184 9938
rect 2190 9934 2194 9938
rect 2200 9934 2204 9938
rect 2210 9934 2214 9938
rect 2175 9929 2179 9933
rect 2185 9929 2189 9933
rect 2195 9929 2199 9933
rect 2205 9929 2209 9933
rect 2215 9929 2219 9933
rect 2180 9924 2184 9928
rect 2190 9924 2194 9928
rect 2200 9924 2204 9928
rect 2210 9924 2214 9928
rect 2175 9919 2179 9923
rect 2185 9919 2189 9923
rect 2195 9919 2199 9923
rect 2205 9919 2209 9923
rect 2215 9919 2219 9923
rect 2180 9914 2184 9918
rect 2190 9914 2194 9918
rect 2200 9914 2204 9918
rect 2210 9914 2214 9918
rect 2175 9909 2179 9913
rect 2185 9909 2189 9913
rect 2195 9909 2199 9913
rect 2205 9909 2209 9913
rect 2215 9909 2219 9913
rect 2180 9904 2184 9908
rect 2190 9904 2194 9908
rect 2200 9904 2204 9908
rect 2210 9904 2214 9908
rect 2175 9899 2179 9903
rect 2185 9899 2189 9903
rect 2195 9899 2199 9903
rect 2205 9899 2209 9903
rect 2215 9899 2219 9903
rect 2180 9894 2184 9898
rect 2190 9894 2194 9898
rect 2200 9894 2204 9898
rect 2210 9894 2214 9898
rect 2175 9889 2179 9893
rect 2185 9889 2189 9893
rect 2195 9889 2199 9893
rect 2205 9889 2209 9893
rect 2215 9889 2219 9893
rect 2180 9884 2184 9888
rect 2190 9884 2194 9888
rect 2200 9884 2204 9888
rect 2210 9884 2214 9888
rect 2175 9879 2179 9883
rect 2185 9879 2189 9883
rect 2195 9879 2199 9883
rect 2205 9879 2209 9883
rect 2215 9879 2219 9883
rect 2180 9874 2184 9878
rect 2190 9874 2194 9878
rect 2200 9874 2204 9878
rect 2210 9874 2214 9878
rect 2175 9869 2179 9873
rect 2185 9869 2189 9873
rect 2195 9869 2199 9873
rect 2205 9869 2209 9873
rect 2215 9869 2219 9873
rect 2180 9864 2184 9868
rect 2190 9864 2194 9868
rect 2200 9864 2204 9868
rect 2210 9864 2214 9868
rect 2163 9848 2167 9852
rect 2170 9848 2174 9852
rect 2175 9848 2179 9852
rect 2180 9848 2184 9852
rect 2185 9848 2189 9852
rect 2190 9848 2194 9852
rect 2195 9848 2199 9852
rect 2200 9848 2204 9852
rect 2205 9848 2209 9852
rect 2210 9848 2214 9852
rect 2215 9848 2219 9852
rect 2220 9848 2224 9852
rect 2227 9848 2231 9852
rect 1778 9827 1782 9831
rect 1836 9827 1840 9831
rect 1778 9811 1782 9815
rect 1836 9811 1840 9815
rect 1673 9796 1677 9800
rect 1678 9796 1682 9800
rect 1778 9795 1782 9799
rect 1673 9791 1677 9795
rect 1678 9791 1682 9795
rect 2324 9949 2328 9953
rect 2334 9949 2338 9953
rect 2344 9949 2348 9953
rect 2354 9949 2358 9953
rect 2364 9949 2368 9953
rect 2329 9944 2333 9948
rect 2339 9944 2343 9948
rect 2349 9944 2353 9948
rect 2359 9944 2363 9948
rect 2324 9939 2328 9943
rect 2334 9939 2338 9943
rect 2344 9939 2348 9943
rect 2354 9939 2358 9943
rect 2364 9939 2368 9943
rect 2329 9934 2333 9938
rect 2339 9934 2343 9938
rect 2349 9934 2353 9938
rect 2359 9934 2363 9938
rect 2324 9929 2328 9933
rect 2334 9929 2338 9933
rect 2344 9929 2348 9933
rect 2354 9929 2358 9933
rect 2364 9929 2368 9933
rect 2329 9924 2333 9928
rect 2339 9924 2343 9928
rect 2349 9924 2353 9928
rect 2359 9924 2363 9928
rect 2324 9919 2328 9923
rect 2334 9919 2338 9923
rect 2344 9919 2348 9923
rect 2354 9919 2358 9923
rect 2364 9919 2368 9923
rect 2329 9914 2333 9918
rect 2339 9914 2343 9918
rect 2349 9914 2353 9918
rect 2359 9914 2363 9918
rect 2324 9909 2328 9913
rect 2334 9909 2338 9913
rect 2344 9909 2348 9913
rect 2354 9909 2358 9913
rect 2364 9909 2368 9913
rect 2329 9904 2333 9908
rect 2339 9904 2343 9908
rect 2349 9904 2353 9908
rect 2359 9904 2363 9908
rect 2324 9899 2328 9903
rect 2334 9899 2338 9903
rect 2344 9899 2348 9903
rect 2354 9899 2358 9903
rect 2364 9899 2368 9903
rect 2329 9894 2333 9898
rect 2339 9894 2343 9898
rect 2349 9894 2353 9898
rect 2359 9894 2363 9898
rect 2324 9889 2328 9893
rect 2334 9889 2338 9893
rect 2344 9889 2348 9893
rect 2354 9889 2358 9893
rect 2364 9889 2368 9893
rect 2329 9884 2333 9888
rect 2339 9884 2343 9888
rect 2349 9884 2353 9888
rect 2359 9884 2363 9888
rect 2324 9879 2328 9883
rect 2334 9879 2338 9883
rect 2344 9879 2348 9883
rect 2354 9879 2358 9883
rect 2364 9879 2368 9883
rect 2329 9874 2333 9878
rect 2339 9874 2343 9878
rect 2349 9874 2353 9878
rect 2359 9874 2363 9878
rect 2324 9869 2328 9873
rect 2334 9869 2338 9873
rect 2344 9869 2348 9873
rect 2354 9869 2358 9873
rect 2364 9869 2368 9873
rect 2329 9864 2333 9868
rect 2339 9864 2343 9868
rect 2349 9864 2353 9868
rect 2359 9864 2363 9868
rect 2312 9848 2316 9852
rect 2319 9848 2323 9852
rect 2324 9848 2328 9852
rect 2329 9848 2333 9852
rect 2334 9848 2338 9852
rect 2339 9848 2343 9852
rect 2344 9848 2348 9852
rect 2349 9848 2353 9852
rect 2354 9848 2358 9852
rect 2359 9848 2363 9852
rect 2364 9848 2368 9852
rect 2369 9848 2373 9852
rect 2376 9848 2380 9852
rect 2484 9949 2488 9953
rect 2494 9949 2498 9953
rect 2504 9949 2508 9953
rect 2514 9949 2518 9953
rect 2524 9949 2528 9953
rect 2489 9944 2493 9948
rect 2499 9944 2503 9948
rect 2509 9944 2513 9948
rect 2519 9944 2523 9948
rect 2484 9939 2488 9943
rect 2494 9939 2498 9943
rect 2504 9939 2508 9943
rect 2514 9939 2518 9943
rect 2524 9939 2528 9943
rect 2489 9934 2493 9938
rect 2499 9934 2503 9938
rect 2509 9934 2513 9938
rect 2519 9934 2523 9938
rect 2484 9929 2488 9933
rect 2494 9929 2498 9933
rect 2504 9929 2508 9933
rect 2514 9929 2518 9933
rect 2524 9929 2528 9933
rect 2489 9924 2493 9928
rect 2499 9924 2503 9928
rect 2509 9924 2513 9928
rect 2519 9924 2523 9928
rect 2484 9919 2488 9923
rect 2494 9919 2498 9923
rect 2504 9919 2508 9923
rect 2514 9919 2518 9923
rect 2524 9919 2528 9923
rect 2489 9914 2493 9918
rect 2499 9914 2503 9918
rect 2509 9914 2513 9918
rect 2519 9914 2523 9918
rect 2484 9909 2488 9913
rect 2494 9909 2498 9913
rect 2504 9909 2508 9913
rect 2514 9909 2518 9913
rect 2524 9909 2528 9913
rect 2489 9904 2493 9908
rect 2499 9904 2503 9908
rect 2509 9904 2513 9908
rect 2519 9904 2523 9908
rect 2484 9899 2488 9903
rect 2494 9899 2498 9903
rect 2504 9899 2508 9903
rect 2514 9899 2518 9903
rect 2524 9899 2528 9903
rect 2489 9894 2493 9898
rect 2499 9894 2503 9898
rect 2509 9894 2513 9898
rect 2519 9894 2523 9898
rect 2484 9889 2488 9893
rect 2494 9889 2498 9893
rect 2504 9889 2508 9893
rect 2514 9889 2518 9893
rect 2524 9889 2528 9893
rect 2489 9884 2493 9888
rect 2499 9884 2503 9888
rect 2509 9884 2513 9888
rect 2519 9884 2523 9888
rect 2484 9879 2488 9883
rect 2494 9879 2498 9883
rect 2504 9879 2508 9883
rect 2514 9879 2518 9883
rect 2524 9879 2528 9883
rect 2489 9874 2493 9878
rect 2499 9874 2503 9878
rect 2509 9874 2513 9878
rect 2519 9874 2523 9878
rect 2484 9869 2488 9873
rect 2494 9869 2498 9873
rect 2504 9869 2508 9873
rect 2514 9869 2518 9873
rect 2524 9869 2528 9873
rect 2489 9864 2493 9868
rect 2499 9864 2503 9868
rect 2509 9864 2513 9868
rect 2519 9864 2523 9868
rect 2472 9848 2476 9852
rect 2479 9848 2483 9852
rect 2484 9848 2488 9852
rect 2489 9848 2493 9852
rect 2494 9848 2498 9852
rect 2499 9848 2503 9852
rect 2504 9848 2508 9852
rect 2509 9848 2513 9852
rect 2514 9848 2518 9852
rect 2519 9848 2523 9852
rect 2524 9848 2528 9852
rect 2529 9848 2533 9852
rect 2536 9848 2540 9852
rect 2087 9827 2091 9831
rect 2145 9827 2149 9831
rect 2087 9811 2091 9815
rect 2145 9811 2149 9815
rect 1836 9795 1840 9799
rect 1673 9786 1677 9790
rect 1678 9786 1682 9790
rect 1673 9781 1677 9785
rect 1678 9781 1682 9785
rect 1673 9776 1677 9780
rect 1678 9776 1682 9780
rect 1778 9779 1782 9783
rect 1673 9771 1677 9775
rect 1678 9771 1682 9775
rect 1673 9766 1677 9770
rect 1678 9766 1682 9770
rect 1628 9757 1632 9761
rect 1633 9757 1637 9761
rect 1638 9757 1642 9761
rect 1643 9757 1647 9761
rect 1628 9747 1632 9751
rect 1633 9747 1637 9751
rect 1638 9747 1642 9751
rect 1643 9747 1647 9751
rect 1628 9737 1632 9741
rect 1633 9737 1637 9741
rect 1638 9737 1642 9741
rect 1643 9737 1647 9741
rect 1673 9761 1677 9765
rect 1678 9761 1682 9765
rect 1673 9756 1677 9760
rect 1678 9756 1682 9760
rect 1673 9751 1677 9755
rect 1678 9751 1682 9755
rect 1673 9746 1677 9750
rect 1678 9746 1682 9750
rect 1673 9741 1677 9745
rect 1678 9741 1682 9745
rect 1673 9736 1677 9740
rect 1678 9736 1682 9740
rect 1569 9718 1573 9722
rect 1574 9718 1578 9722
rect 1579 9718 1583 9722
rect 1584 9718 1588 9722
rect 1589 9718 1593 9722
rect 1594 9718 1598 9722
rect 1599 9718 1603 9722
rect 1604 9718 1608 9722
rect 1609 9718 1613 9722
rect 1614 9718 1618 9722
rect 1619 9718 1623 9722
rect 1569 9713 1573 9717
rect 1574 9713 1578 9717
rect 1579 9713 1583 9717
rect 1584 9713 1588 9717
rect 1589 9713 1593 9717
rect 1594 9713 1598 9717
rect 1599 9713 1603 9717
rect 1604 9713 1608 9717
rect 1609 9713 1613 9717
rect 1614 9713 1618 9717
rect 1619 9713 1623 9717
rect 1499 9706 1503 9710
rect 1504 9706 1508 9710
rect 1499 9701 1503 9705
rect 1504 9701 1508 9705
rect 1499 9696 1503 9700
rect 1504 9696 1508 9700
rect 1499 9691 1503 9695
rect 1504 9691 1508 9695
rect 1499 9686 1503 9690
rect 1504 9686 1508 9690
rect 1628 9711 1632 9715
rect 1633 9711 1637 9715
rect 1638 9711 1642 9715
rect 1643 9711 1647 9715
rect 1628 9701 1632 9705
rect 1633 9701 1637 9705
rect 1638 9701 1642 9705
rect 1643 9701 1647 9705
rect 1628 9691 1632 9695
rect 1633 9691 1637 9695
rect 1638 9691 1642 9695
rect 1643 9691 1647 9695
rect 1499 9681 1503 9685
rect 1504 9681 1508 9685
rect 1499 9676 1503 9680
rect 1504 9676 1508 9680
rect 1499 9671 1503 9675
rect 1504 9671 1508 9675
rect 1499 9666 1503 9670
rect 1504 9666 1508 9670
rect 1499 9661 1503 9665
rect 1504 9661 1508 9665
rect 664 9603 668 9607
rect 674 9603 678 9607
rect 684 9603 688 9607
rect 618 9592 622 9596
rect 628 9592 632 9596
rect 638 9592 642 9596
rect 618 9587 622 9591
rect 628 9587 632 9591
rect 638 9587 642 9591
rect 618 9582 622 9586
rect 628 9582 632 9586
rect 638 9582 642 9586
rect 618 9577 622 9581
rect 628 9577 632 9581
rect 638 9577 642 9581
rect 664 9592 668 9596
rect 674 9592 678 9596
rect 684 9592 688 9596
rect 1836 9779 1840 9783
rect 1982 9796 1986 9800
rect 1987 9796 1991 9800
rect 2087 9795 2091 9799
rect 1982 9791 1986 9795
rect 1987 9791 1991 9795
rect 2633 9949 2637 9953
rect 2643 9949 2647 9953
rect 2653 9949 2657 9953
rect 2663 9949 2667 9953
rect 2673 9949 2677 9953
rect 2638 9944 2642 9948
rect 2648 9944 2652 9948
rect 2658 9944 2662 9948
rect 2668 9944 2672 9948
rect 2633 9939 2637 9943
rect 2643 9939 2647 9943
rect 2653 9939 2657 9943
rect 2663 9939 2667 9943
rect 2673 9939 2677 9943
rect 2638 9934 2642 9938
rect 2648 9934 2652 9938
rect 2658 9934 2662 9938
rect 2668 9934 2672 9938
rect 2633 9929 2637 9933
rect 2643 9929 2647 9933
rect 2653 9929 2657 9933
rect 2663 9929 2667 9933
rect 2673 9929 2677 9933
rect 2638 9924 2642 9928
rect 2648 9924 2652 9928
rect 2658 9924 2662 9928
rect 2668 9924 2672 9928
rect 2633 9919 2637 9923
rect 2643 9919 2647 9923
rect 2653 9919 2657 9923
rect 2663 9919 2667 9923
rect 2673 9919 2677 9923
rect 2638 9914 2642 9918
rect 2648 9914 2652 9918
rect 2658 9914 2662 9918
rect 2668 9914 2672 9918
rect 2633 9909 2637 9913
rect 2643 9909 2647 9913
rect 2653 9909 2657 9913
rect 2663 9909 2667 9913
rect 2673 9909 2677 9913
rect 2638 9904 2642 9908
rect 2648 9904 2652 9908
rect 2658 9904 2662 9908
rect 2668 9904 2672 9908
rect 2633 9899 2637 9903
rect 2643 9899 2647 9903
rect 2653 9899 2657 9903
rect 2663 9899 2667 9903
rect 2673 9899 2677 9903
rect 2638 9894 2642 9898
rect 2648 9894 2652 9898
rect 2658 9894 2662 9898
rect 2668 9894 2672 9898
rect 2633 9889 2637 9893
rect 2643 9889 2647 9893
rect 2653 9889 2657 9893
rect 2663 9889 2667 9893
rect 2673 9889 2677 9893
rect 2638 9884 2642 9888
rect 2648 9884 2652 9888
rect 2658 9884 2662 9888
rect 2668 9884 2672 9888
rect 2633 9879 2637 9883
rect 2643 9879 2647 9883
rect 2653 9879 2657 9883
rect 2663 9879 2667 9883
rect 2673 9879 2677 9883
rect 2638 9874 2642 9878
rect 2648 9874 2652 9878
rect 2658 9874 2662 9878
rect 2668 9874 2672 9878
rect 2633 9869 2637 9873
rect 2643 9869 2647 9873
rect 2653 9869 2657 9873
rect 2663 9869 2667 9873
rect 2673 9869 2677 9873
rect 2638 9864 2642 9868
rect 2648 9864 2652 9868
rect 2658 9864 2662 9868
rect 2668 9864 2672 9868
rect 2621 9848 2625 9852
rect 2628 9848 2632 9852
rect 2633 9848 2637 9852
rect 2638 9848 2642 9852
rect 2643 9848 2647 9852
rect 2648 9848 2652 9852
rect 2653 9848 2657 9852
rect 2658 9848 2662 9852
rect 2663 9848 2667 9852
rect 2668 9848 2672 9852
rect 2673 9848 2677 9852
rect 2678 9848 2682 9852
rect 2685 9848 2689 9852
rect 2793 9949 2797 9953
rect 2803 9949 2807 9953
rect 2813 9949 2817 9953
rect 2823 9949 2827 9953
rect 2833 9949 2837 9953
rect 2798 9944 2802 9948
rect 2808 9944 2812 9948
rect 2818 9944 2822 9948
rect 2828 9944 2832 9948
rect 2793 9939 2797 9943
rect 2803 9939 2807 9943
rect 2813 9939 2817 9943
rect 2823 9939 2827 9943
rect 2833 9939 2837 9943
rect 2798 9934 2802 9938
rect 2808 9934 2812 9938
rect 2818 9934 2822 9938
rect 2828 9934 2832 9938
rect 2793 9929 2797 9933
rect 2803 9929 2807 9933
rect 2813 9929 2817 9933
rect 2823 9929 2827 9933
rect 2833 9929 2837 9933
rect 2798 9924 2802 9928
rect 2808 9924 2812 9928
rect 2818 9924 2822 9928
rect 2828 9924 2832 9928
rect 2793 9919 2797 9923
rect 2803 9919 2807 9923
rect 2813 9919 2817 9923
rect 2823 9919 2827 9923
rect 2833 9919 2837 9923
rect 2798 9914 2802 9918
rect 2808 9914 2812 9918
rect 2818 9914 2822 9918
rect 2828 9914 2832 9918
rect 2793 9909 2797 9913
rect 2803 9909 2807 9913
rect 2813 9909 2817 9913
rect 2823 9909 2827 9913
rect 2833 9909 2837 9913
rect 2798 9904 2802 9908
rect 2808 9904 2812 9908
rect 2818 9904 2822 9908
rect 2828 9904 2832 9908
rect 2793 9899 2797 9903
rect 2803 9899 2807 9903
rect 2813 9899 2817 9903
rect 2823 9899 2827 9903
rect 2833 9899 2837 9903
rect 2798 9894 2802 9898
rect 2808 9894 2812 9898
rect 2818 9894 2822 9898
rect 2828 9894 2832 9898
rect 2793 9889 2797 9893
rect 2803 9889 2807 9893
rect 2813 9889 2817 9893
rect 2823 9889 2827 9893
rect 2833 9889 2837 9893
rect 2798 9884 2802 9888
rect 2808 9884 2812 9888
rect 2818 9884 2822 9888
rect 2828 9884 2832 9888
rect 2793 9879 2797 9883
rect 2803 9879 2807 9883
rect 2813 9879 2817 9883
rect 2823 9879 2827 9883
rect 2833 9879 2837 9883
rect 2798 9874 2802 9878
rect 2808 9874 2812 9878
rect 2818 9874 2822 9878
rect 2828 9874 2832 9878
rect 2793 9869 2797 9873
rect 2803 9869 2807 9873
rect 2813 9869 2817 9873
rect 2823 9869 2827 9873
rect 2833 9869 2837 9873
rect 2798 9864 2802 9868
rect 2808 9864 2812 9868
rect 2818 9864 2822 9868
rect 2828 9864 2832 9868
rect 2781 9848 2785 9852
rect 2788 9848 2792 9852
rect 2793 9848 2797 9852
rect 2798 9848 2802 9852
rect 2803 9848 2807 9852
rect 2808 9848 2812 9852
rect 2813 9848 2817 9852
rect 2818 9848 2822 9852
rect 2823 9848 2827 9852
rect 2828 9848 2832 9852
rect 2833 9848 2837 9852
rect 2838 9848 2842 9852
rect 2845 9848 2849 9852
rect 2396 9827 2400 9831
rect 2454 9827 2458 9831
rect 2396 9811 2400 9815
rect 2454 9811 2458 9815
rect 2145 9795 2149 9799
rect 1982 9786 1986 9790
rect 1987 9786 1991 9790
rect 1982 9781 1986 9785
rect 1987 9781 1991 9785
rect 1982 9776 1986 9780
rect 1987 9776 1991 9780
rect 2087 9779 2091 9783
rect 1982 9771 1986 9775
rect 1987 9771 1991 9775
rect 1982 9766 1986 9770
rect 1987 9766 1991 9770
rect 1937 9757 1941 9761
rect 1942 9757 1946 9761
rect 1947 9757 1951 9761
rect 1952 9757 1956 9761
rect 1937 9747 1941 9751
rect 1942 9747 1946 9751
rect 1947 9747 1951 9751
rect 1952 9747 1956 9751
rect 1937 9737 1941 9741
rect 1942 9737 1946 9741
rect 1947 9737 1951 9741
rect 1952 9737 1956 9741
rect 1982 9761 1986 9765
rect 1987 9761 1991 9765
rect 1982 9756 1986 9760
rect 1987 9756 1991 9760
rect 1982 9751 1986 9755
rect 1987 9751 1991 9755
rect 1982 9746 1986 9750
rect 1987 9746 1991 9750
rect 1982 9741 1986 9745
rect 1987 9741 1991 9745
rect 1982 9736 1986 9740
rect 1987 9736 1991 9740
rect 1878 9718 1882 9722
rect 1883 9718 1887 9722
rect 1888 9718 1892 9722
rect 1893 9718 1897 9722
rect 1898 9718 1902 9722
rect 1903 9718 1907 9722
rect 1908 9718 1912 9722
rect 1913 9718 1917 9722
rect 1918 9718 1922 9722
rect 1923 9718 1927 9722
rect 1928 9718 1932 9722
rect 1878 9713 1882 9717
rect 1883 9713 1887 9717
rect 1888 9713 1892 9717
rect 1893 9713 1897 9717
rect 1898 9713 1902 9717
rect 1903 9713 1907 9717
rect 1908 9713 1912 9717
rect 1913 9713 1917 9717
rect 1918 9713 1922 9717
rect 1923 9713 1927 9717
rect 1928 9713 1932 9717
rect 1937 9711 1941 9715
rect 1942 9711 1946 9715
rect 1947 9711 1951 9715
rect 1952 9711 1956 9715
rect 1937 9701 1941 9705
rect 1942 9701 1946 9705
rect 1947 9701 1951 9705
rect 1952 9701 1956 9705
rect 1937 9691 1941 9695
rect 1942 9691 1946 9695
rect 1947 9691 1951 9695
rect 1952 9691 1956 9695
rect 2145 9779 2149 9783
rect 2291 9796 2295 9800
rect 2296 9796 2300 9800
rect 2396 9795 2400 9799
rect 2291 9791 2295 9795
rect 2296 9791 2300 9795
rect 2942 9949 2946 9953
rect 2952 9949 2956 9953
rect 2962 9949 2966 9953
rect 2972 9949 2976 9953
rect 2982 9949 2986 9953
rect 2947 9944 2951 9948
rect 2957 9944 2961 9948
rect 2967 9944 2971 9948
rect 2977 9944 2981 9948
rect 2942 9939 2946 9943
rect 2952 9939 2956 9943
rect 2962 9939 2966 9943
rect 2972 9939 2976 9943
rect 2982 9939 2986 9943
rect 2947 9934 2951 9938
rect 2957 9934 2961 9938
rect 2967 9934 2971 9938
rect 2977 9934 2981 9938
rect 2942 9929 2946 9933
rect 2952 9929 2956 9933
rect 2962 9929 2966 9933
rect 2972 9929 2976 9933
rect 2982 9929 2986 9933
rect 2947 9924 2951 9928
rect 2957 9924 2961 9928
rect 2967 9924 2971 9928
rect 2977 9924 2981 9928
rect 2942 9919 2946 9923
rect 2952 9919 2956 9923
rect 2962 9919 2966 9923
rect 2972 9919 2976 9923
rect 2982 9919 2986 9923
rect 2947 9914 2951 9918
rect 2957 9914 2961 9918
rect 2967 9914 2971 9918
rect 2977 9914 2981 9918
rect 2942 9909 2946 9913
rect 2952 9909 2956 9913
rect 2962 9909 2966 9913
rect 2972 9909 2976 9913
rect 2982 9909 2986 9913
rect 2947 9904 2951 9908
rect 2957 9904 2961 9908
rect 2967 9904 2971 9908
rect 2977 9904 2981 9908
rect 2942 9899 2946 9903
rect 2952 9899 2956 9903
rect 2962 9899 2966 9903
rect 2972 9899 2976 9903
rect 2982 9899 2986 9903
rect 2947 9894 2951 9898
rect 2957 9894 2961 9898
rect 2967 9894 2971 9898
rect 2977 9894 2981 9898
rect 2942 9889 2946 9893
rect 2952 9889 2956 9893
rect 2962 9889 2966 9893
rect 2972 9889 2976 9893
rect 2982 9889 2986 9893
rect 2947 9884 2951 9888
rect 2957 9884 2961 9888
rect 2967 9884 2971 9888
rect 2977 9884 2981 9888
rect 2942 9879 2946 9883
rect 2952 9879 2956 9883
rect 2962 9879 2966 9883
rect 2972 9879 2976 9883
rect 2982 9879 2986 9883
rect 2947 9874 2951 9878
rect 2957 9874 2961 9878
rect 2967 9874 2971 9878
rect 2977 9874 2981 9878
rect 2942 9869 2946 9873
rect 2952 9869 2956 9873
rect 2962 9869 2966 9873
rect 2972 9869 2976 9873
rect 2982 9869 2986 9873
rect 2947 9864 2951 9868
rect 2957 9864 2961 9868
rect 2967 9864 2971 9868
rect 2977 9864 2981 9868
rect 2930 9848 2934 9852
rect 2937 9848 2941 9852
rect 2942 9848 2946 9852
rect 2947 9848 2951 9852
rect 2952 9848 2956 9852
rect 2957 9848 2961 9852
rect 2962 9848 2966 9852
rect 2967 9848 2971 9852
rect 2972 9848 2976 9852
rect 2977 9848 2981 9852
rect 2982 9848 2986 9852
rect 2987 9848 2991 9852
rect 2994 9848 2998 9852
rect 3102 9949 3106 9953
rect 3112 9949 3116 9953
rect 3122 9949 3126 9953
rect 3132 9949 3136 9953
rect 3142 9949 3146 9953
rect 3107 9944 3111 9948
rect 3117 9944 3121 9948
rect 3127 9944 3131 9948
rect 3137 9944 3141 9948
rect 3102 9939 3106 9943
rect 3112 9939 3116 9943
rect 3122 9939 3126 9943
rect 3132 9939 3136 9943
rect 3142 9939 3146 9943
rect 3107 9934 3111 9938
rect 3117 9934 3121 9938
rect 3127 9934 3131 9938
rect 3137 9934 3141 9938
rect 3102 9929 3106 9933
rect 3112 9929 3116 9933
rect 3122 9929 3126 9933
rect 3132 9929 3136 9933
rect 3142 9929 3146 9933
rect 3107 9924 3111 9928
rect 3117 9924 3121 9928
rect 3127 9924 3131 9928
rect 3137 9924 3141 9928
rect 3102 9919 3106 9923
rect 3112 9919 3116 9923
rect 3122 9919 3126 9923
rect 3132 9919 3136 9923
rect 3142 9919 3146 9923
rect 3107 9914 3111 9918
rect 3117 9914 3121 9918
rect 3127 9914 3131 9918
rect 3137 9914 3141 9918
rect 3102 9909 3106 9913
rect 3112 9909 3116 9913
rect 3122 9909 3126 9913
rect 3132 9909 3136 9913
rect 3142 9909 3146 9913
rect 3107 9904 3111 9908
rect 3117 9904 3121 9908
rect 3127 9904 3131 9908
rect 3137 9904 3141 9908
rect 3102 9899 3106 9903
rect 3112 9899 3116 9903
rect 3122 9899 3126 9903
rect 3132 9899 3136 9903
rect 3142 9899 3146 9903
rect 3107 9894 3111 9898
rect 3117 9894 3121 9898
rect 3127 9894 3131 9898
rect 3137 9894 3141 9898
rect 3102 9889 3106 9893
rect 3112 9889 3116 9893
rect 3122 9889 3126 9893
rect 3132 9889 3136 9893
rect 3142 9889 3146 9893
rect 3107 9884 3111 9888
rect 3117 9884 3121 9888
rect 3127 9884 3131 9888
rect 3137 9884 3141 9888
rect 3102 9879 3106 9883
rect 3112 9879 3116 9883
rect 3122 9879 3126 9883
rect 3132 9879 3136 9883
rect 3142 9879 3146 9883
rect 3107 9874 3111 9878
rect 3117 9874 3121 9878
rect 3127 9874 3131 9878
rect 3137 9874 3141 9878
rect 3102 9869 3106 9873
rect 3112 9869 3116 9873
rect 3122 9869 3126 9873
rect 3132 9869 3136 9873
rect 3142 9869 3146 9873
rect 3107 9864 3111 9868
rect 3117 9864 3121 9868
rect 3127 9864 3131 9868
rect 3137 9864 3141 9868
rect 3090 9848 3094 9852
rect 3097 9848 3101 9852
rect 3102 9848 3106 9852
rect 3107 9848 3111 9852
rect 3112 9848 3116 9852
rect 3117 9848 3121 9852
rect 3122 9848 3126 9852
rect 3127 9848 3131 9852
rect 3132 9848 3136 9852
rect 3137 9848 3141 9852
rect 3142 9848 3146 9852
rect 3147 9848 3151 9852
rect 3154 9848 3158 9852
rect 2705 9827 2709 9831
rect 2763 9827 2767 9831
rect 2705 9811 2709 9815
rect 2763 9811 2767 9815
rect 2454 9795 2458 9799
rect 2291 9786 2295 9790
rect 2296 9786 2300 9790
rect 2291 9781 2295 9785
rect 2296 9781 2300 9785
rect 2291 9776 2295 9780
rect 2296 9776 2300 9780
rect 2396 9779 2400 9783
rect 2291 9771 2295 9775
rect 2296 9771 2300 9775
rect 2291 9766 2295 9770
rect 2296 9766 2300 9770
rect 2246 9757 2250 9761
rect 2251 9757 2255 9761
rect 2256 9757 2260 9761
rect 2261 9757 2265 9761
rect 2246 9747 2250 9751
rect 2251 9747 2255 9751
rect 2256 9747 2260 9751
rect 2261 9747 2265 9751
rect 2246 9737 2250 9741
rect 2251 9737 2255 9741
rect 2256 9737 2260 9741
rect 2261 9737 2265 9741
rect 2291 9761 2295 9765
rect 2296 9761 2300 9765
rect 2291 9756 2295 9760
rect 2296 9756 2300 9760
rect 2291 9751 2295 9755
rect 2296 9751 2300 9755
rect 2291 9746 2295 9750
rect 2296 9746 2300 9750
rect 2291 9741 2295 9745
rect 2296 9741 2300 9745
rect 2291 9736 2295 9740
rect 2296 9736 2300 9740
rect 2187 9718 2191 9722
rect 2192 9718 2196 9722
rect 2197 9718 2201 9722
rect 2202 9718 2206 9722
rect 2207 9718 2211 9722
rect 2212 9718 2216 9722
rect 2217 9718 2221 9722
rect 2222 9718 2226 9722
rect 2227 9718 2231 9722
rect 2232 9718 2236 9722
rect 2237 9718 2241 9722
rect 2187 9713 2191 9717
rect 2192 9713 2196 9717
rect 2197 9713 2201 9717
rect 2202 9713 2206 9717
rect 2207 9713 2211 9717
rect 2212 9713 2216 9717
rect 2217 9713 2221 9717
rect 2222 9713 2226 9717
rect 2227 9713 2231 9717
rect 2232 9713 2236 9717
rect 2237 9713 2241 9717
rect 2246 9711 2250 9715
rect 2251 9711 2255 9715
rect 2256 9711 2260 9715
rect 2261 9711 2265 9715
rect 2246 9701 2250 9705
rect 2251 9701 2255 9705
rect 2256 9701 2260 9705
rect 2261 9701 2265 9705
rect 2246 9691 2250 9695
rect 2251 9691 2255 9695
rect 2256 9691 2260 9695
rect 2261 9691 2265 9695
rect 2113 9593 2126 9597
rect 2454 9779 2458 9783
rect 2600 9796 2604 9800
rect 2605 9796 2609 9800
rect 2705 9795 2709 9799
rect 2600 9791 2604 9795
rect 2605 9791 2609 9795
rect 3251 9949 3255 9953
rect 3261 9949 3265 9953
rect 3271 9949 3275 9953
rect 3281 9949 3285 9953
rect 3291 9949 3295 9953
rect 3256 9944 3260 9948
rect 3266 9944 3270 9948
rect 3276 9944 3280 9948
rect 3286 9944 3290 9948
rect 3251 9939 3255 9943
rect 3261 9939 3265 9943
rect 3271 9939 3275 9943
rect 3281 9939 3285 9943
rect 3291 9939 3295 9943
rect 3256 9934 3260 9938
rect 3266 9934 3270 9938
rect 3276 9934 3280 9938
rect 3286 9934 3290 9938
rect 3251 9929 3255 9933
rect 3261 9929 3265 9933
rect 3271 9929 3275 9933
rect 3281 9929 3285 9933
rect 3291 9929 3295 9933
rect 3256 9924 3260 9928
rect 3266 9924 3270 9928
rect 3276 9924 3280 9928
rect 3286 9924 3290 9928
rect 3251 9919 3255 9923
rect 3261 9919 3265 9923
rect 3271 9919 3275 9923
rect 3281 9919 3285 9923
rect 3291 9919 3295 9923
rect 3256 9914 3260 9918
rect 3266 9914 3270 9918
rect 3276 9914 3280 9918
rect 3286 9914 3290 9918
rect 3251 9909 3255 9913
rect 3261 9909 3265 9913
rect 3271 9909 3275 9913
rect 3281 9909 3285 9913
rect 3291 9909 3295 9913
rect 3256 9904 3260 9908
rect 3266 9904 3270 9908
rect 3276 9904 3280 9908
rect 3286 9904 3290 9908
rect 3251 9899 3255 9903
rect 3261 9899 3265 9903
rect 3271 9899 3275 9903
rect 3281 9899 3285 9903
rect 3291 9899 3295 9903
rect 3256 9894 3260 9898
rect 3266 9894 3270 9898
rect 3276 9894 3280 9898
rect 3286 9894 3290 9898
rect 3251 9889 3255 9893
rect 3261 9889 3265 9893
rect 3271 9889 3275 9893
rect 3281 9889 3285 9893
rect 3291 9889 3295 9893
rect 3256 9884 3260 9888
rect 3266 9884 3270 9888
rect 3276 9884 3280 9888
rect 3286 9884 3290 9888
rect 3251 9879 3255 9883
rect 3261 9879 3265 9883
rect 3271 9879 3275 9883
rect 3281 9879 3285 9883
rect 3291 9879 3295 9883
rect 3256 9874 3260 9878
rect 3266 9874 3270 9878
rect 3276 9874 3280 9878
rect 3286 9874 3290 9878
rect 3251 9869 3255 9873
rect 3261 9869 3265 9873
rect 3271 9869 3275 9873
rect 3281 9869 3285 9873
rect 3291 9869 3295 9873
rect 3256 9864 3260 9868
rect 3266 9864 3270 9868
rect 3276 9864 3280 9868
rect 3286 9864 3290 9868
rect 3239 9848 3243 9852
rect 3246 9848 3250 9852
rect 3251 9848 3255 9852
rect 3256 9848 3260 9852
rect 3261 9848 3265 9852
rect 3266 9848 3270 9852
rect 3271 9848 3275 9852
rect 3276 9848 3280 9852
rect 3281 9848 3285 9852
rect 3286 9848 3290 9852
rect 3291 9848 3295 9852
rect 3296 9848 3300 9852
rect 3303 9848 3307 9852
rect 3014 9827 3018 9831
rect 3072 9827 3076 9831
rect 3014 9811 3018 9815
rect 3072 9811 3076 9815
rect 2763 9795 2767 9799
rect 2600 9786 2604 9790
rect 2605 9786 2609 9790
rect 2600 9781 2604 9785
rect 2605 9781 2609 9785
rect 2600 9776 2604 9780
rect 2605 9776 2609 9780
rect 2705 9779 2709 9783
rect 2600 9771 2604 9775
rect 2605 9771 2609 9775
rect 2600 9766 2604 9770
rect 2605 9766 2609 9770
rect 2555 9757 2559 9761
rect 2560 9757 2564 9761
rect 2565 9757 2569 9761
rect 2570 9757 2574 9761
rect 2555 9747 2559 9751
rect 2560 9747 2564 9751
rect 2565 9747 2569 9751
rect 2570 9747 2574 9751
rect 2555 9737 2559 9741
rect 2560 9737 2564 9741
rect 2565 9737 2569 9741
rect 2570 9737 2574 9741
rect 2600 9761 2604 9765
rect 2605 9761 2609 9765
rect 2600 9756 2604 9760
rect 2605 9756 2609 9760
rect 2600 9751 2604 9755
rect 2605 9751 2609 9755
rect 2600 9746 2604 9750
rect 2605 9746 2609 9750
rect 2600 9741 2604 9745
rect 2605 9741 2609 9745
rect 2600 9736 2604 9740
rect 2605 9736 2609 9740
rect 2496 9718 2500 9722
rect 2501 9718 2505 9722
rect 2506 9718 2510 9722
rect 2511 9718 2515 9722
rect 2516 9718 2520 9722
rect 2521 9718 2525 9722
rect 2526 9718 2530 9722
rect 2531 9718 2535 9722
rect 2536 9718 2540 9722
rect 2541 9718 2545 9722
rect 2546 9718 2550 9722
rect 2496 9713 2500 9717
rect 2501 9713 2505 9717
rect 2506 9713 2510 9717
rect 2511 9713 2515 9717
rect 2516 9713 2520 9717
rect 2521 9713 2525 9717
rect 2526 9713 2530 9717
rect 2531 9713 2535 9717
rect 2536 9713 2540 9717
rect 2541 9713 2545 9717
rect 2546 9713 2550 9717
rect 2555 9711 2559 9715
rect 2560 9711 2564 9715
rect 2565 9711 2569 9715
rect 2570 9711 2574 9715
rect 2555 9701 2559 9705
rect 2560 9701 2564 9705
rect 2565 9701 2569 9705
rect 2570 9701 2574 9705
rect 2555 9691 2559 9695
rect 2560 9691 2564 9695
rect 2565 9691 2569 9695
rect 2570 9691 2574 9695
rect 2763 9779 2767 9783
rect 2909 9796 2913 9800
rect 2914 9796 2918 9800
rect 3014 9795 3018 9799
rect 2909 9791 2913 9795
rect 2914 9791 2918 9795
rect 3072 9795 3076 9799
rect 2909 9786 2913 9790
rect 2914 9786 2918 9790
rect 2909 9781 2913 9785
rect 2914 9781 2918 9785
rect 2909 9776 2913 9780
rect 2914 9776 2918 9780
rect 3014 9779 3018 9783
rect 2909 9771 2913 9775
rect 2914 9771 2918 9775
rect 2909 9766 2913 9770
rect 2914 9766 2918 9770
rect 2864 9757 2868 9761
rect 2869 9757 2873 9761
rect 2874 9757 2878 9761
rect 2879 9757 2883 9761
rect 2864 9747 2868 9751
rect 2869 9747 2873 9751
rect 2874 9747 2878 9751
rect 2879 9747 2883 9751
rect 2864 9737 2868 9741
rect 2869 9737 2873 9741
rect 2874 9737 2878 9741
rect 2879 9737 2883 9741
rect 2909 9761 2913 9765
rect 2914 9761 2918 9765
rect 2909 9756 2913 9760
rect 2914 9756 2918 9760
rect 2909 9751 2913 9755
rect 2914 9751 2918 9755
rect 2909 9746 2913 9750
rect 2914 9746 2918 9750
rect 2909 9741 2913 9745
rect 2914 9741 2918 9745
rect 2909 9736 2913 9740
rect 2914 9736 2918 9740
rect 2805 9718 2809 9722
rect 2810 9718 2814 9722
rect 2815 9718 2819 9722
rect 2820 9718 2824 9722
rect 2825 9718 2829 9722
rect 2830 9718 2834 9722
rect 2835 9718 2839 9722
rect 2840 9718 2844 9722
rect 2845 9718 2849 9722
rect 2850 9718 2854 9722
rect 2855 9718 2859 9722
rect 2805 9713 2809 9717
rect 2810 9713 2814 9717
rect 2815 9713 2819 9717
rect 2820 9713 2824 9717
rect 2825 9713 2829 9717
rect 2830 9713 2834 9717
rect 2835 9713 2839 9717
rect 2840 9713 2844 9717
rect 2845 9713 2849 9717
rect 2850 9713 2854 9717
rect 2855 9713 2859 9717
rect 2864 9711 2868 9715
rect 2869 9711 2873 9715
rect 2874 9711 2878 9715
rect 2879 9711 2883 9715
rect 2864 9701 2868 9705
rect 2869 9701 2873 9705
rect 2874 9701 2878 9705
rect 2879 9701 2883 9705
rect 2864 9691 2868 9695
rect 2869 9691 2873 9695
rect 2874 9691 2878 9695
rect 2879 9691 2883 9695
rect 3072 9779 3076 9783
rect 3218 9796 3222 9800
rect 3223 9796 3227 9800
rect 3218 9791 3222 9795
rect 3223 9791 3227 9795
rect 3218 9786 3222 9790
rect 3223 9786 3227 9790
rect 3218 9781 3222 9785
rect 3223 9781 3227 9785
rect 3218 9776 3222 9780
rect 3223 9776 3227 9780
rect 3218 9771 3222 9775
rect 3223 9771 3227 9775
rect 3218 9766 3222 9770
rect 3223 9766 3227 9770
rect 3173 9757 3177 9761
rect 3178 9757 3182 9761
rect 3183 9757 3187 9761
rect 3188 9757 3192 9761
rect 3173 9747 3177 9751
rect 3178 9747 3182 9751
rect 3183 9747 3187 9751
rect 3188 9747 3192 9751
rect 3173 9737 3177 9741
rect 3178 9737 3182 9741
rect 3183 9737 3187 9741
rect 3188 9737 3192 9741
rect 3218 9761 3222 9765
rect 3223 9761 3227 9765
rect 3218 9756 3222 9760
rect 3223 9756 3227 9760
rect 3218 9751 3222 9755
rect 3223 9751 3227 9755
rect 3218 9746 3222 9750
rect 3223 9746 3227 9750
rect 3218 9741 3222 9745
rect 3223 9741 3227 9745
rect 3218 9736 3222 9740
rect 3223 9736 3227 9740
rect 3114 9718 3118 9722
rect 3119 9718 3123 9722
rect 3124 9718 3128 9722
rect 3129 9718 3133 9722
rect 3134 9718 3138 9722
rect 3139 9718 3143 9722
rect 3144 9718 3148 9722
rect 3149 9718 3153 9722
rect 3154 9718 3158 9722
rect 3159 9718 3163 9722
rect 3164 9718 3168 9722
rect 3114 9713 3118 9717
rect 3119 9713 3123 9717
rect 3124 9713 3128 9717
rect 3129 9713 3133 9717
rect 3134 9713 3138 9717
rect 3139 9713 3143 9717
rect 3144 9713 3148 9717
rect 3149 9713 3153 9717
rect 3154 9713 3158 9717
rect 3159 9713 3163 9717
rect 3164 9713 3168 9717
rect 3173 9711 3177 9715
rect 3178 9711 3182 9715
rect 3183 9711 3187 9715
rect 3188 9711 3192 9715
rect 3173 9701 3177 9705
rect 3178 9701 3182 9705
rect 3183 9701 3187 9705
rect 3188 9701 3192 9705
rect 3173 9691 3177 9695
rect 3178 9691 3182 9695
rect 3183 9691 3187 9695
rect 3188 9691 3192 9695
rect 3411 9949 3415 9953
rect 3421 9949 3425 9953
rect 3431 9949 3435 9953
rect 3441 9949 3445 9953
rect 3451 9949 3455 9953
rect 3416 9944 3420 9948
rect 3426 9944 3430 9948
rect 3436 9944 3440 9948
rect 3446 9944 3450 9948
rect 3411 9939 3415 9943
rect 3421 9939 3425 9943
rect 3431 9939 3435 9943
rect 3441 9939 3445 9943
rect 3451 9939 3455 9943
rect 3416 9934 3420 9938
rect 3426 9934 3430 9938
rect 3436 9934 3440 9938
rect 3446 9934 3450 9938
rect 3411 9929 3415 9933
rect 3421 9929 3425 9933
rect 3431 9929 3435 9933
rect 3441 9929 3445 9933
rect 3451 9929 3455 9933
rect 3416 9924 3420 9928
rect 3426 9924 3430 9928
rect 3436 9924 3440 9928
rect 3446 9924 3450 9928
rect 3411 9919 3415 9923
rect 3421 9919 3425 9923
rect 3431 9919 3435 9923
rect 3441 9919 3445 9923
rect 3451 9919 3455 9923
rect 3416 9914 3420 9918
rect 3426 9914 3430 9918
rect 3436 9914 3440 9918
rect 3446 9914 3450 9918
rect 3411 9909 3415 9913
rect 3421 9909 3425 9913
rect 3431 9909 3435 9913
rect 3441 9909 3445 9913
rect 3451 9909 3455 9913
rect 3416 9904 3420 9908
rect 3426 9904 3430 9908
rect 3436 9904 3440 9908
rect 3446 9904 3450 9908
rect 3411 9899 3415 9903
rect 3421 9899 3425 9903
rect 3431 9899 3435 9903
rect 3441 9899 3445 9903
rect 3451 9899 3455 9903
rect 3416 9894 3420 9898
rect 3426 9894 3430 9898
rect 3436 9894 3440 9898
rect 3446 9894 3450 9898
rect 3411 9889 3415 9893
rect 3421 9889 3425 9893
rect 3431 9889 3435 9893
rect 3441 9889 3445 9893
rect 3451 9889 3455 9893
rect 3416 9884 3420 9888
rect 3426 9884 3430 9888
rect 3436 9884 3440 9888
rect 3446 9884 3450 9888
rect 3411 9879 3415 9883
rect 3421 9879 3425 9883
rect 3431 9879 3435 9883
rect 3441 9879 3445 9883
rect 3451 9879 3455 9883
rect 3416 9874 3420 9878
rect 3426 9874 3430 9878
rect 3436 9874 3440 9878
rect 3446 9874 3450 9878
rect 3411 9869 3415 9873
rect 3421 9869 3425 9873
rect 3431 9869 3435 9873
rect 3441 9869 3445 9873
rect 3451 9869 3455 9873
rect 3416 9864 3420 9868
rect 3426 9864 3430 9868
rect 3436 9864 3440 9868
rect 3446 9864 3450 9868
rect 3399 9848 3403 9852
rect 3406 9848 3410 9852
rect 3411 9848 3415 9852
rect 3416 9848 3420 9852
rect 3421 9848 3425 9852
rect 3426 9848 3430 9852
rect 3431 9848 3435 9852
rect 3436 9848 3440 9852
rect 3441 9848 3445 9852
rect 3446 9848 3450 9852
rect 3451 9848 3455 9852
rect 3456 9848 3460 9852
rect 3463 9848 3467 9852
rect 3560 9949 3564 9953
rect 3570 9949 3574 9953
rect 3580 9949 3584 9953
rect 3590 9949 3594 9953
rect 3600 9949 3604 9953
rect 3565 9944 3569 9948
rect 3575 9944 3579 9948
rect 3585 9944 3589 9948
rect 3595 9944 3599 9948
rect 3560 9939 3564 9943
rect 3570 9939 3574 9943
rect 3580 9939 3584 9943
rect 3590 9939 3594 9943
rect 3600 9939 3604 9943
rect 3565 9934 3569 9938
rect 3575 9934 3579 9938
rect 3585 9934 3589 9938
rect 3595 9934 3599 9938
rect 3560 9929 3564 9933
rect 3570 9929 3574 9933
rect 3580 9929 3584 9933
rect 3590 9929 3594 9933
rect 3600 9929 3604 9933
rect 3565 9924 3569 9928
rect 3575 9924 3579 9928
rect 3585 9924 3589 9928
rect 3595 9924 3599 9928
rect 3560 9919 3564 9923
rect 3570 9919 3574 9923
rect 3580 9919 3584 9923
rect 3590 9919 3594 9923
rect 3600 9919 3604 9923
rect 3565 9914 3569 9918
rect 3575 9914 3579 9918
rect 3585 9914 3589 9918
rect 3595 9914 3599 9918
rect 3560 9909 3564 9913
rect 3570 9909 3574 9913
rect 3580 9909 3584 9913
rect 3590 9909 3594 9913
rect 3600 9909 3604 9913
rect 3565 9904 3569 9908
rect 3575 9904 3579 9908
rect 3585 9904 3589 9908
rect 3595 9904 3599 9908
rect 3560 9899 3564 9903
rect 3570 9899 3574 9903
rect 3580 9899 3584 9903
rect 3590 9899 3594 9903
rect 3600 9899 3604 9903
rect 3565 9894 3569 9898
rect 3575 9894 3579 9898
rect 3585 9894 3589 9898
rect 3595 9894 3599 9898
rect 3560 9889 3564 9893
rect 3570 9889 3574 9893
rect 3580 9889 3584 9893
rect 3590 9889 3594 9893
rect 3600 9889 3604 9893
rect 3565 9884 3569 9888
rect 3575 9884 3579 9888
rect 3585 9884 3589 9888
rect 3595 9884 3599 9888
rect 3560 9879 3564 9883
rect 3570 9879 3574 9883
rect 3580 9879 3584 9883
rect 3590 9879 3594 9883
rect 3600 9879 3604 9883
rect 3565 9874 3569 9878
rect 3575 9874 3579 9878
rect 3585 9874 3589 9878
rect 3595 9874 3599 9878
rect 3560 9869 3564 9873
rect 3570 9869 3574 9873
rect 3580 9869 3584 9873
rect 3590 9869 3594 9873
rect 3600 9869 3604 9873
rect 3565 9864 3569 9868
rect 3575 9864 3579 9868
rect 3585 9864 3589 9868
rect 3595 9864 3599 9868
rect 3548 9848 3552 9852
rect 3555 9848 3559 9852
rect 3560 9848 3564 9852
rect 3565 9848 3569 9852
rect 3570 9848 3574 9852
rect 3575 9848 3579 9852
rect 3580 9848 3584 9852
rect 3585 9848 3589 9852
rect 3590 9848 3594 9852
rect 3595 9848 3599 9852
rect 3600 9848 3604 9852
rect 3605 9848 3609 9852
rect 3612 9848 3616 9852
rect 3353 9711 3357 9715
rect 3358 9711 3362 9715
rect 3527 9796 3531 9800
rect 3532 9796 3536 9800
rect 3527 9791 3531 9795
rect 3532 9791 3536 9795
rect 3527 9786 3531 9790
rect 3532 9786 3536 9790
rect 3527 9781 3531 9785
rect 3532 9781 3536 9785
rect 3527 9776 3531 9780
rect 3532 9776 3536 9780
rect 3527 9771 3531 9775
rect 3532 9771 3536 9775
rect 3527 9766 3531 9770
rect 3532 9766 3536 9770
rect 3482 9757 3486 9761
rect 3487 9757 3491 9761
rect 3492 9757 3496 9761
rect 3497 9757 3501 9761
rect 3482 9747 3486 9751
rect 3487 9747 3491 9751
rect 3492 9747 3496 9751
rect 3497 9747 3501 9751
rect 3482 9737 3486 9741
rect 3487 9737 3491 9741
rect 3492 9737 3496 9741
rect 3497 9737 3501 9741
rect 3527 9761 3531 9765
rect 3532 9761 3536 9765
rect 3527 9756 3531 9760
rect 3532 9756 3536 9760
rect 3527 9751 3531 9755
rect 3532 9751 3536 9755
rect 3527 9746 3531 9750
rect 3532 9746 3536 9750
rect 3527 9741 3531 9745
rect 3532 9741 3536 9745
rect 3527 9736 3531 9740
rect 3532 9736 3536 9740
rect 3720 9949 3724 9953
rect 3730 9949 3734 9953
rect 3740 9949 3744 9953
rect 3750 9949 3754 9953
rect 3760 9949 3764 9953
rect 3725 9944 3729 9948
rect 3735 9944 3739 9948
rect 3745 9944 3749 9948
rect 3755 9944 3759 9948
rect 3720 9939 3724 9943
rect 3730 9939 3734 9943
rect 3740 9939 3744 9943
rect 3750 9939 3754 9943
rect 3760 9939 3764 9943
rect 3725 9934 3729 9938
rect 3735 9934 3739 9938
rect 3745 9934 3749 9938
rect 3755 9934 3759 9938
rect 3720 9929 3724 9933
rect 3730 9929 3734 9933
rect 3740 9929 3744 9933
rect 3750 9929 3754 9933
rect 3760 9929 3764 9933
rect 3725 9924 3729 9928
rect 3735 9924 3739 9928
rect 3745 9924 3749 9928
rect 3755 9924 3759 9928
rect 3720 9919 3724 9923
rect 3730 9919 3734 9923
rect 3740 9919 3744 9923
rect 3750 9919 3754 9923
rect 3760 9919 3764 9923
rect 3725 9914 3729 9918
rect 3735 9914 3739 9918
rect 3745 9914 3749 9918
rect 3755 9914 3759 9918
rect 3720 9909 3724 9913
rect 3730 9909 3734 9913
rect 3740 9909 3744 9913
rect 3750 9909 3754 9913
rect 3760 9909 3764 9913
rect 3725 9904 3729 9908
rect 3735 9904 3739 9908
rect 3745 9904 3749 9908
rect 3755 9904 3759 9908
rect 3720 9899 3724 9903
rect 3730 9899 3734 9903
rect 3740 9899 3744 9903
rect 3750 9899 3754 9903
rect 3760 9899 3764 9903
rect 3725 9894 3729 9898
rect 3735 9894 3739 9898
rect 3745 9894 3749 9898
rect 3755 9894 3759 9898
rect 3720 9889 3724 9893
rect 3730 9889 3734 9893
rect 3740 9889 3744 9893
rect 3750 9889 3754 9893
rect 3760 9889 3764 9893
rect 3725 9884 3729 9888
rect 3735 9884 3739 9888
rect 3745 9884 3749 9888
rect 3755 9884 3759 9888
rect 3720 9879 3724 9883
rect 3730 9879 3734 9883
rect 3740 9879 3744 9883
rect 3750 9879 3754 9883
rect 3760 9879 3764 9883
rect 3725 9874 3729 9878
rect 3735 9874 3739 9878
rect 3745 9874 3749 9878
rect 3755 9874 3759 9878
rect 3720 9869 3724 9873
rect 3730 9869 3734 9873
rect 3740 9869 3744 9873
rect 3750 9869 3754 9873
rect 3760 9869 3764 9873
rect 3725 9864 3729 9868
rect 3735 9864 3739 9868
rect 3745 9864 3749 9868
rect 3755 9864 3759 9868
rect 3708 9848 3712 9852
rect 3715 9848 3719 9852
rect 3720 9848 3724 9852
rect 3725 9848 3729 9852
rect 3730 9848 3734 9852
rect 3735 9848 3739 9852
rect 3740 9848 3744 9852
rect 3745 9848 3749 9852
rect 3750 9848 3754 9852
rect 3755 9848 3759 9852
rect 3760 9848 3764 9852
rect 3765 9848 3769 9852
rect 3772 9848 3776 9852
rect 3869 9949 3873 9953
rect 3879 9949 3883 9953
rect 3889 9949 3893 9953
rect 3899 9949 3903 9953
rect 3909 9949 3913 9953
rect 3874 9944 3878 9948
rect 3884 9944 3888 9948
rect 3894 9944 3898 9948
rect 3904 9944 3908 9948
rect 3869 9939 3873 9943
rect 3879 9939 3883 9943
rect 3889 9939 3893 9943
rect 3899 9939 3903 9943
rect 3909 9939 3913 9943
rect 3874 9934 3878 9938
rect 3884 9934 3888 9938
rect 3894 9934 3898 9938
rect 3904 9934 3908 9938
rect 3869 9929 3873 9933
rect 3879 9929 3883 9933
rect 3889 9929 3893 9933
rect 3899 9929 3903 9933
rect 3909 9929 3913 9933
rect 3874 9924 3878 9928
rect 3884 9924 3888 9928
rect 3894 9924 3898 9928
rect 3904 9924 3908 9928
rect 3869 9919 3873 9923
rect 3879 9919 3883 9923
rect 3889 9919 3893 9923
rect 3899 9919 3903 9923
rect 3909 9919 3913 9923
rect 3874 9914 3878 9918
rect 3884 9914 3888 9918
rect 3894 9914 3898 9918
rect 3904 9914 3908 9918
rect 3869 9909 3873 9913
rect 3879 9909 3883 9913
rect 3889 9909 3893 9913
rect 3899 9909 3903 9913
rect 3909 9909 3913 9913
rect 3874 9904 3878 9908
rect 3884 9904 3888 9908
rect 3894 9904 3898 9908
rect 3904 9904 3908 9908
rect 3869 9899 3873 9903
rect 3879 9899 3883 9903
rect 3889 9899 3893 9903
rect 3899 9899 3903 9903
rect 3909 9899 3913 9903
rect 3874 9894 3878 9898
rect 3884 9894 3888 9898
rect 3894 9894 3898 9898
rect 3904 9894 3908 9898
rect 3869 9889 3873 9893
rect 3879 9889 3883 9893
rect 3889 9889 3893 9893
rect 3899 9889 3903 9893
rect 3909 9889 3913 9893
rect 3874 9884 3878 9888
rect 3884 9884 3888 9888
rect 3894 9884 3898 9888
rect 3904 9884 3908 9888
rect 3869 9879 3873 9883
rect 3879 9879 3883 9883
rect 3889 9879 3893 9883
rect 3899 9879 3903 9883
rect 3909 9879 3913 9883
rect 3874 9874 3878 9878
rect 3884 9874 3888 9878
rect 3894 9874 3898 9878
rect 3904 9874 3908 9878
rect 3869 9869 3873 9873
rect 3879 9869 3883 9873
rect 3889 9869 3893 9873
rect 3899 9869 3903 9873
rect 3909 9869 3913 9873
rect 3874 9864 3878 9868
rect 3884 9864 3888 9868
rect 3894 9864 3898 9868
rect 3904 9864 3908 9868
rect 3857 9848 3861 9852
rect 3864 9848 3868 9852
rect 3869 9848 3873 9852
rect 3874 9848 3878 9852
rect 3879 9848 3883 9852
rect 3884 9848 3888 9852
rect 3889 9848 3893 9852
rect 3894 9848 3898 9852
rect 3899 9848 3903 9852
rect 3904 9848 3908 9852
rect 3909 9848 3913 9852
rect 3914 9848 3918 9852
rect 3921 9848 3925 9852
rect 4029 9949 4033 9953
rect 4039 9949 4043 9953
rect 4049 9949 4053 9953
rect 4059 9949 4063 9953
rect 4069 9949 4073 9953
rect 4034 9944 4038 9948
rect 4044 9944 4048 9948
rect 4054 9944 4058 9948
rect 4064 9944 4068 9948
rect 4029 9939 4033 9943
rect 4039 9939 4043 9943
rect 4049 9939 4053 9943
rect 4059 9939 4063 9943
rect 4069 9939 4073 9943
rect 4034 9934 4038 9938
rect 4044 9934 4048 9938
rect 4054 9934 4058 9938
rect 4064 9934 4068 9938
rect 4029 9929 4033 9933
rect 4039 9929 4043 9933
rect 4049 9929 4053 9933
rect 4059 9929 4063 9933
rect 4069 9929 4073 9933
rect 4034 9924 4038 9928
rect 4044 9924 4048 9928
rect 4054 9924 4058 9928
rect 4064 9924 4068 9928
rect 4029 9919 4033 9923
rect 4039 9919 4043 9923
rect 4049 9919 4053 9923
rect 4059 9919 4063 9923
rect 4069 9919 4073 9923
rect 4034 9914 4038 9918
rect 4044 9914 4048 9918
rect 4054 9914 4058 9918
rect 4064 9914 4068 9918
rect 4029 9909 4033 9913
rect 4039 9909 4043 9913
rect 4049 9909 4053 9913
rect 4059 9909 4063 9913
rect 4069 9909 4073 9913
rect 4034 9904 4038 9908
rect 4044 9904 4048 9908
rect 4054 9904 4058 9908
rect 4064 9904 4068 9908
rect 4029 9899 4033 9903
rect 4039 9899 4043 9903
rect 4049 9899 4053 9903
rect 4059 9899 4063 9903
rect 4069 9899 4073 9903
rect 4034 9894 4038 9898
rect 4044 9894 4048 9898
rect 4054 9894 4058 9898
rect 4064 9894 4068 9898
rect 4029 9889 4033 9893
rect 4039 9889 4043 9893
rect 4049 9889 4053 9893
rect 4059 9889 4063 9893
rect 4069 9889 4073 9893
rect 4034 9884 4038 9888
rect 4044 9884 4048 9888
rect 4054 9884 4058 9888
rect 4064 9884 4068 9888
rect 4029 9879 4033 9883
rect 4039 9879 4043 9883
rect 4049 9879 4053 9883
rect 4059 9879 4063 9883
rect 4069 9879 4073 9883
rect 4034 9874 4038 9878
rect 4044 9874 4048 9878
rect 4054 9874 4058 9878
rect 4064 9874 4068 9878
rect 4029 9869 4033 9873
rect 4039 9869 4043 9873
rect 4049 9869 4053 9873
rect 4059 9869 4063 9873
rect 4069 9869 4073 9873
rect 4034 9864 4038 9868
rect 4044 9864 4048 9868
rect 4054 9864 4058 9868
rect 4064 9864 4068 9868
rect 4017 9848 4021 9852
rect 4024 9848 4028 9852
rect 4029 9848 4033 9852
rect 4034 9848 4038 9852
rect 4039 9848 4043 9852
rect 4044 9848 4048 9852
rect 4049 9848 4053 9852
rect 4054 9848 4058 9852
rect 4059 9848 4063 9852
rect 4064 9848 4068 9852
rect 4069 9848 4073 9852
rect 4074 9848 4078 9852
rect 4081 9848 4085 9852
rect 3662 9791 3666 9795
rect 3667 9791 3671 9795
rect 3662 9786 3666 9790
rect 3667 9786 3671 9790
rect 3662 9781 3666 9785
rect 3667 9781 3671 9785
rect 3662 9776 3666 9780
rect 3667 9776 3671 9780
rect 3662 9771 3666 9775
rect 3667 9771 3671 9775
rect 3662 9766 3666 9770
rect 3667 9766 3671 9770
rect 3662 9761 3666 9765
rect 3667 9761 3671 9765
rect 3662 9756 3666 9760
rect 3667 9756 3671 9760
rect 3662 9751 3666 9755
rect 3667 9751 3671 9755
rect 3662 9746 3666 9750
rect 3667 9746 3671 9750
rect 3662 9741 3666 9745
rect 3667 9741 3671 9745
rect 3423 9718 3427 9722
rect 3428 9718 3432 9722
rect 3433 9718 3437 9722
rect 3438 9718 3442 9722
rect 3443 9718 3447 9722
rect 3448 9718 3452 9722
rect 3453 9718 3457 9722
rect 3458 9718 3462 9722
rect 3463 9718 3467 9722
rect 3468 9718 3472 9722
rect 3473 9718 3477 9722
rect 3423 9713 3427 9717
rect 3428 9713 3432 9717
rect 3433 9713 3437 9717
rect 3438 9713 3442 9717
rect 3443 9713 3447 9717
rect 3448 9713 3452 9717
rect 3453 9713 3457 9717
rect 3458 9713 3462 9717
rect 3463 9713 3467 9717
rect 3468 9713 3472 9717
rect 3473 9713 3477 9717
rect 3353 9706 3357 9710
rect 3358 9706 3362 9710
rect 3353 9701 3357 9705
rect 3358 9701 3362 9705
rect 3353 9696 3357 9700
rect 3358 9696 3362 9700
rect 3353 9691 3357 9695
rect 3358 9691 3362 9695
rect 3353 9686 3357 9690
rect 3358 9686 3362 9690
rect 3482 9711 3486 9715
rect 3487 9711 3491 9715
rect 3492 9711 3496 9715
rect 3497 9711 3501 9715
rect 3482 9701 3486 9705
rect 3487 9701 3491 9705
rect 3492 9701 3496 9705
rect 3497 9701 3501 9705
rect 3482 9691 3486 9695
rect 3487 9691 3491 9695
rect 3492 9691 3496 9695
rect 3497 9691 3501 9695
rect 3021 9605 3026 9609
rect 3040 9607 3053 9611
rect 3353 9681 3357 9685
rect 3358 9681 3362 9685
rect 3353 9676 3357 9680
rect 3358 9676 3362 9680
rect 3353 9671 3357 9675
rect 3358 9671 3362 9675
rect 3353 9666 3357 9670
rect 3358 9666 3362 9670
rect 3353 9661 3357 9665
rect 3358 9661 3362 9665
rect 3327 9606 3379 9610
rect 3941 9827 3945 9831
rect 3999 9827 4003 9831
rect 3941 9811 3945 9815
rect 3999 9811 4003 9815
rect 3836 9796 3840 9800
rect 3841 9796 3845 9800
rect 3941 9795 3945 9799
rect 3836 9791 3840 9795
rect 3841 9791 3845 9795
rect 3999 9795 4003 9799
rect 3836 9786 3840 9790
rect 3841 9786 3845 9790
rect 3836 9781 3840 9785
rect 3841 9781 3845 9785
rect 3836 9776 3840 9780
rect 3841 9776 3845 9780
rect 3941 9779 3945 9783
rect 3836 9771 3840 9775
rect 3841 9771 3845 9775
rect 3836 9766 3840 9770
rect 3841 9766 3845 9770
rect 3791 9757 3795 9761
rect 3796 9757 3800 9761
rect 3801 9757 3805 9761
rect 3806 9757 3810 9761
rect 3791 9747 3795 9751
rect 3796 9747 3800 9751
rect 3801 9747 3805 9751
rect 3806 9747 3810 9751
rect 3791 9737 3795 9741
rect 3796 9737 3800 9741
rect 3801 9737 3805 9741
rect 3806 9737 3810 9741
rect 3836 9761 3840 9765
rect 3841 9761 3845 9765
rect 3836 9756 3840 9760
rect 3841 9756 3845 9760
rect 3836 9751 3840 9755
rect 3841 9751 3845 9755
rect 3836 9746 3840 9750
rect 3841 9746 3845 9750
rect 3836 9741 3840 9745
rect 3841 9741 3845 9745
rect 3836 9736 3840 9740
rect 3841 9736 3845 9740
rect 3732 9718 3736 9722
rect 3737 9718 3741 9722
rect 3742 9718 3746 9722
rect 3747 9718 3751 9722
rect 3752 9718 3756 9722
rect 3757 9718 3761 9722
rect 3762 9718 3766 9722
rect 3767 9718 3771 9722
rect 3772 9718 3776 9722
rect 3777 9718 3781 9722
rect 3782 9718 3786 9722
rect 3732 9713 3736 9717
rect 3737 9713 3741 9717
rect 3742 9713 3746 9717
rect 3747 9713 3751 9717
rect 3752 9713 3756 9717
rect 3757 9713 3761 9717
rect 3762 9713 3766 9717
rect 3767 9713 3771 9717
rect 3772 9713 3776 9717
rect 3777 9713 3781 9717
rect 3782 9713 3786 9717
rect 3791 9711 3795 9715
rect 3796 9711 3800 9715
rect 3801 9711 3805 9715
rect 3806 9711 3810 9715
rect 3791 9701 3795 9705
rect 3796 9701 3800 9705
rect 3801 9701 3805 9705
rect 3806 9701 3810 9705
rect 3791 9691 3795 9695
rect 3796 9691 3800 9695
rect 3801 9691 3805 9695
rect 3806 9691 3810 9695
rect 3634 9604 3690 9609
rect 664 9587 668 9591
rect 674 9587 678 9591
rect 684 9587 688 9591
rect 664 9582 668 9586
rect 674 9582 678 9586
rect 684 9582 688 9586
rect 664 9577 668 9581
rect 674 9577 678 9581
rect 684 9577 688 9581
rect 2422 9575 2435 9597
rect 2497 9575 2502 9597
rect 3999 9779 4003 9783
rect 4100 9757 4104 9761
rect 4105 9757 4109 9761
rect 4110 9757 4114 9761
rect 4115 9757 4119 9761
rect 4100 9747 4104 9751
rect 4105 9747 4109 9751
rect 4110 9747 4114 9751
rect 4115 9747 4119 9751
rect 4100 9737 4104 9741
rect 4105 9737 4109 9741
rect 4110 9737 4114 9741
rect 4115 9737 4119 9741
rect 4292 9757 4296 9761
rect 4297 9757 4301 9761
rect 4302 9757 4306 9761
rect 4307 9757 4311 9761
rect 4292 9747 4296 9751
rect 4297 9747 4301 9751
rect 4302 9747 4306 9751
rect 4307 9747 4311 9751
rect 4292 9737 4296 9741
rect 4297 9737 4301 9741
rect 4302 9737 4306 9741
rect 4307 9737 4311 9741
rect 4318 9757 4322 9761
rect 4323 9757 4327 9761
rect 4328 9757 4332 9761
rect 4333 9757 4337 9761
rect 4318 9747 4322 9751
rect 4323 9747 4327 9751
rect 4328 9747 4332 9751
rect 4333 9747 4337 9751
rect 4318 9737 4322 9741
rect 4323 9737 4327 9741
rect 4328 9737 4332 9741
rect 4333 9737 4337 9741
rect 4344 9757 4348 9761
rect 4349 9757 4353 9761
rect 4354 9757 4358 9761
rect 4359 9757 4363 9761
rect 4344 9747 4348 9751
rect 4349 9747 4353 9751
rect 4354 9747 4358 9751
rect 4359 9747 4363 9751
rect 4344 9737 4348 9741
rect 4349 9737 4353 9741
rect 4354 9737 4358 9741
rect 4359 9737 4363 9741
rect 4370 9757 4374 9761
rect 4375 9757 4379 9761
rect 4380 9757 4384 9761
rect 4385 9757 4389 9761
rect 4370 9747 4374 9751
rect 4375 9747 4379 9751
rect 4380 9747 4384 9751
rect 4385 9747 4389 9751
rect 4370 9737 4374 9741
rect 4375 9737 4379 9741
rect 4380 9737 4384 9741
rect 4385 9737 4389 9741
rect 4396 9757 4400 9761
rect 4401 9757 4405 9761
rect 4406 9757 4410 9761
rect 4411 9757 4415 9761
rect 4396 9747 4400 9751
rect 4401 9747 4405 9751
rect 4406 9747 4410 9751
rect 4411 9747 4415 9751
rect 4396 9737 4400 9741
rect 4401 9737 4405 9741
rect 4406 9737 4410 9741
rect 4411 9737 4415 9741
rect 4041 9718 4045 9722
rect 4046 9718 4050 9722
rect 4051 9718 4055 9722
rect 4056 9718 4060 9722
rect 4061 9718 4065 9722
rect 4066 9718 4070 9722
rect 4071 9718 4075 9722
rect 4076 9718 4080 9722
rect 4081 9718 4085 9722
rect 4086 9718 4090 9722
rect 4091 9718 4095 9722
rect 4041 9713 4045 9717
rect 4046 9713 4050 9717
rect 4051 9713 4055 9717
rect 4056 9713 4060 9717
rect 4061 9713 4065 9717
rect 4066 9713 4070 9717
rect 4071 9713 4075 9717
rect 4076 9713 4080 9717
rect 4081 9713 4085 9717
rect 4086 9713 4090 9717
rect 4091 9713 4095 9717
rect 4100 9711 4104 9715
rect 4105 9711 4109 9715
rect 4110 9711 4114 9715
rect 4115 9711 4119 9715
rect 4100 9701 4104 9705
rect 4105 9701 4109 9705
rect 4110 9701 4114 9705
rect 4115 9701 4119 9705
rect 4100 9691 4104 9695
rect 4105 9691 4109 9695
rect 4110 9691 4114 9695
rect 4115 9691 4119 9695
rect 4292 9711 4296 9715
rect 4297 9711 4301 9715
rect 4302 9711 4306 9715
rect 4307 9711 4311 9715
rect 4292 9701 4296 9705
rect 4297 9701 4301 9705
rect 4302 9701 4306 9705
rect 4307 9701 4311 9705
rect 4292 9691 4296 9695
rect 4297 9691 4301 9695
rect 4302 9691 4306 9695
rect 4307 9691 4311 9695
rect 4318 9711 4322 9715
rect 4323 9711 4327 9715
rect 4328 9711 4332 9715
rect 4333 9711 4337 9715
rect 4318 9701 4322 9705
rect 4323 9701 4327 9705
rect 4328 9701 4332 9705
rect 4333 9701 4337 9705
rect 4318 9691 4322 9695
rect 4323 9691 4327 9695
rect 4328 9691 4332 9695
rect 4333 9691 4337 9695
rect 4344 9711 4348 9715
rect 4349 9711 4353 9715
rect 4354 9711 4358 9715
rect 4359 9711 4363 9715
rect 4344 9701 4348 9705
rect 4349 9701 4353 9705
rect 4354 9701 4358 9705
rect 4359 9701 4363 9705
rect 4344 9691 4348 9695
rect 4349 9691 4353 9695
rect 4354 9691 4358 9695
rect 4359 9691 4363 9695
rect 4370 9711 4374 9715
rect 4375 9711 4379 9715
rect 4380 9711 4384 9715
rect 4385 9711 4389 9715
rect 4370 9701 4374 9705
rect 4375 9701 4379 9705
rect 4380 9701 4384 9705
rect 4385 9701 4389 9705
rect 4370 9691 4374 9695
rect 4375 9691 4379 9695
rect 4380 9691 4384 9695
rect 4385 9691 4389 9695
rect 4396 9711 4400 9715
rect 4401 9711 4405 9715
rect 4406 9711 4410 9715
rect 4411 9711 4415 9715
rect 4396 9701 4400 9705
rect 4401 9701 4405 9705
rect 4406 9701 4410 9705
rect 4411 9701 4415 9705
rect 4396 9691 4400 9695
rect 4401 9691 4405 9695
rect 4406 9691 4410 9695
rect 4411 9691 4415 9695
rect 618 9566 622 9570
rect 628 9566 632 9570
rect 638 9566 642 9570
rect 618 9561 622 9565
rect 628 9561 632 9565
rect 638 9561 642 9565
rect 618 9556 622 9560
rect 628 9556 632 9560
rect 638 9556 642 9560
rect 618 9551 622 9555
rect 628 9551 632 9555
rect 638 9551 642 9555
rect 664 9566 668 9570
rect 674 9566 678 9570
rect 684 9566 688 9570
rect 664 9561 668 9565
rect 674 9561 678 9565
rect 684 9561 688 9565
rect 664 9556 668 9560
rect 674 9556 678 9560
rect 684 9556 688 9560
rect 664 9551 668 9555
rect 674 9551 678 9555
rect 684 9551 688 9555
rect 2113 9547 2134 9572
rect 2401 9549 2414 9571
rect 2476 9549 2481 9571
rect 618 9540 622 9544
rect 628 9540 632 9544
rect 638 9540 642 9544
rect 618 9535 622 9539
rect 628 9535 632 9539
rect 638 9535 642 9539
rect 618 9530 622 9534
rect 628 9530 632 9534
rect 638 9530 642 9534
rect 618 9525 622 9529
rect 628 9525 632 9529
rect 638 9525 642 9529
rect 664 9540 668 9544
rect 674 9540 678 9544
rect 684 9540 688 9544
rect 664 9535 668 9539
rect 674 9535 678 9539
rect 684 9535 688 9539
rect 664 9530 668 9534
rect 674 9530 678 9534
rect 684 9530 688 9534
rect 664 9525 668 9529
rect 674 9525 678 9529
rect 684 9525 688 9529
rect 618 9514 622 9518
rect 628 9514 632 9518
rect 638 9514 642 9518
rect 618 9509 622 9513
rect 628 9509 632 9513
rect 638 9509 642 9513
rect 618 9504 622 9508
rect 628 9504 632 9508
rect 638 9504 642 9508
rect 618 9499 622 9503
rect 628 9499 632 9503
rect 638 9499 642 9503
rect 664 9514 668 9518
rect 674 9514 678 9518
rect 684 9514 688 9518
rect 664 9509 668 9513
rect 674 9509 678 9513
rect 684 9509 688 9513
rect 664 9504 668 9508
rect 674 9504 678 9508
rect 684 9504 688 9508
rect 664 9499 668 9503
rect 674 9499 678 9503
rect 684 9499 688 9503
rect 2824 9497 2830 9501
rect 3769 9497 3775 9501
rect 2812 9489 2818 9493
rect 3757 9489 3763 9493
rect 2800 9482 2806 9486
rect 3745 9482 3751 9486
rect 2788 9475 2794 9479
rect 3733 9475 3739 9479
rect 2776 9466 2782 9471
rect 3327 9467 3382 9471
rect 3721 9467 3727 9471
rect 2764 9459 2770 9463
rect 3635 9459 3690 9463
rect 3709 9460 3715 9464
rect 4484 9573 4488 9577
rect 4494 9573 4498 9577
rect 4504 9573 4508 9577
rect 4484 9568 4488 9572
rect 4494 9568 4498 9572
rect 4504 9568 4508 9572
rect 4484 9563 4488 9567
rect 4494 9563 4498 9567
rect 4504 9563 4508 9567
rect 4484 9558 4488 9562
rect 4494 9558 4498 9562
rect 4504 9558 4508 9562
rect 4530 9573 4534 9577
rect 4540 9573 4544 9577
rect 4550 9573 4554 9577
rect 4530 9568 4534 9572
rect 4540 9568 4544 9572
rect 4550 9568 4554 9572
rect 4530 9563 4534 9567
rect 4540 9563 4544 9567
rect 4550 9563 4554 9567
rect 4530 9558 4534 9562
rect 4540 9558 4544 9562
rect 4550 9558 4554 9562
rect 4484 9544 4488 9548
rect 4494 9544 4498 9548
rect 4504 9544 4508 9548
rect 4484 9539 4488 9543
rect 4494 9539 4498 9543
rect 4504 9539 4508 9543
rect 4484 9534 4488 9538
rect 4494 9534 4498 9538
rect 4504 9534 4508 9538
rect 4484 9529 4488 9533
rect 4494 9529 4498 9533
rect 4504 9529 4508 9533
rect 4530 9544 4534 9548
rect 4540 9544 4544 9548
rect 4550 9544 4554 9548
rect 4530 9539 4534 9543
rect 4540 9539 4544 9543
rect 4550 9539 4554 9543
rect 4530 9534 4534 9538
rect 4540 9534 4544 9538
rect 4550 9534 4554 9538
rect 4530 9529 4534 9533
rect 4540 9529 4544 9533
rect 4550 9529 4554 9533
rect 4484 9515 4488 9519
rect 4494 9515 4498 9519
rect 4504 9515 4508 9519
rect 4484 9510 4488 9514
rect 4494 9510 4498 9514
rect 4504 9510 4508 9514
rect 4484 9505 4488 9509
rect 4494 9505 4498 9509
rect 4504 9505 4508 9509
rect 4484 9500 4488 9504
rect 4494 9500 4498 9504
rect 4504 9500 4508 9504
rect 4530 9515 4534 9519
rect 4540 9515 4544 9519
rect 4550 9515 4554 9519
rect 4530 9510 4534 9514
rect 4540 9510 4544 9514
rect 4550 9510 4554 9514
rect 4530 9505 4534 9509
rect 4540 9505 4544 9509
rect 4550 9505 4554 9509
rect 4530 9500 4534 9504
rect 4540 9500 4544 9504
rect 4550 9500 4554 9504
rect 4484 9486 4488 9490
rect 4494 9486 4498 9490
rect 4504 9486 4508 9490
rect 4484 9481 4488 9485
rect 4494 9481 4498 9485
rect 4504 9481 4508 9485
rect 4484 9476 4488 9480
rect 4494 9476 4498 9480
rect 4504 9476 4508 9480
rect 4484 9471 4488 9475
rect 4494 9471 4498 9475
rect 4504 9471 4508 9475
rect 4530 9486 4534 9490
rect 4540 9486 4544 9490
rect 4550 9486 4554 9490
rect 4530 9481 4534 9485
rect 4540 9481 4544 9485
rect 4550 9481 4554 9485
rect 4530 9476 4534 9480
rect 4540 9476 4544 9480
rect 4550 9476 4554 9480
rect 4530 9471 4534 9475
rect 4540 9471 4544 9475
rect 4550 9471 4554 9475
rect 2836 9452 2842 9456
rect 3781 9452 3787 9456
rect 4484 9457 4488 9461
rect 4494 9457 4498 9461
rect 4504 9457 4508 9461
rect 4484 9452 4488 9456
rect 4494 9452 4498 9456
rect 4504 9452 4508 9456
rect 3040 9444 3053 9448
rect 3423 9444 3427 9448
rect 4484 9447 4488 9451
rect 4494 9447 4498 9451
rect 4504 9447 4508 9451
rect 4484 9442 4488 9446
rect 4494 9442 4498 9446
rect 4504 9442 4508 9446
rect 4530 9457 4534 9461
rect 4540 9457 4544 9461
rect 4550 9457 4554 9461
rect 4530 9452 4534 9456
rect 4540 9452 4544 9456
rect 4550 9452 4554 9456
rect 4530 9447 4534 9451
rect 4540 9447 4544 9451
rect 4550 9447 4554 9451
rect 4530 9442 4534 9446
rect 4540 9442 4544 9446
rect 4550 9442 4554 9446
rect 3021 9434 3026 9438
rect 3411 9434 3416 9438
rect 3757 9412 3763 9416
rect 3745 9404 3751 9408
rect 3733 9396 3739 9400
rect 3721 9388 3727 9392
rect 3709 9380 3715 9384
rect 2824 9347 2830 9351
rect 2857 9347 2861 9351
rect 2893 9347 2897 9351
rect 2960 9347 2964 9351
rect 2989 9347 2993 9351
rect 3025 9347 3029 9351
rect 3092 9347 3096 9351
rect 3121 9347 3125 9351
rect 3157 9347 3161 9351
rect 3224 9347 3228 9351
rect 3253 9347 3257 9351
rect 3289 9347 3293 9351
rect 3356 9347 3360 9351
rect 3769 9347 3775 9351
rect 3802 9347 3806 9351
rect 3838 9347 3842 9351
rect 3905 9347 3909 9351
rect 3934 9347 3938 9351
rect 3970 9347 3974 9351
rect 4037 9347 4041 9351
rect 4066 9347 4070 9351
rect 4102 9347 4106 9351
rect 4169 9347 4173 9351
rect 4198 9347 4202 9351
rect 4234 9347 4238 9351
rect 4301 9347 4305 9351
rect 2764 9340 2770 9344
rect 3709 9340 3715 9344
rect 2857 9333 2861 9337
rect 2907 9333 2911 9337
rect 2960 9333 2964 9337
rect 2989 9333 2993 9337
rect 3039 9333 3043 9337
rect 3092 9333 3096 9337
rect 3121 9333 3125 9337
rect 3171 9333 3175 9337
rect 3224 9333 3228 9337
rect 3253 9333 3257 9337
rect 3303 9333 3307 9337
rect 3356 9333 3360 9337
rect 3802 9333 3806 9337
rect 3852 9333 3856 9337
rect 3905 9333 3909 9337
rect 3934 9333 3938 9337
rect 3984 9333 3988 9337
rect 4037 9333 4041 9337
rect 4066 9333 4070 9337
rect 4116 9333 4120 9337
rect 4169 9333 4173 9337
rect 4198 9333 4202 9337
rect 4248 9333 4252 9337
rect 4301 9333 4305 9337
rect 618 9321 622 9325
rect 628 9321 632 9325
rect 638 9321 642 9325
rect 618 9316 622 9320
rect 628 9316 632 9320
rect 638 9316 642 9320
rect 618 9311 622 9315
rect 628 9311 632 9315
rect 638 9311 642 9315
rect 618 9306 622 9310
rect 628 9306 632 9310
rect 638 9306 642 9310
rect 664 9321 668 9325
rect 674 9321 678 9325
rect 684 9321 688 9325
rect 2880 9322 2884 9326
rect 664 9316 668 9320
rect 674 9316 678 9320
rect 684 9316 688 9320
rect 664 9311 668 9315
rect 674 9311 678 9315
rect 684 9311 688 9315
rect 2505 9314 2509 9318
rect 2541 9314 2545 9318
rect 2608 9314 2612 9318
rect 2824 9314 2830 9318
rect 2851 9313 2855 9317
rect 2864 9316 2868 9322
rect 2901 9316 2905 9322
rect 2914 9318 2918 9322
rect 2938 9322 2942 9326
rect 3012 9322 3016 9326
rect 2922 9316 2926 9322
rect 2959 9316 2963 9322
rect 2975 9318 2979 9322
rect 664 9306 668 9310
rect 674 9306 678 9310
rect 684 9306 688 9310
rect 2764 9307 2770 9311
rect 2505 9300 2509 9304
rect 2555 9300 2559 9304
rect 2608 9300 2612 9304
rect 2864 9303 2868 9307
rect 2880 9303 2884 9309
rect 2914 9309 2918 9313
rect 2901 9303 2905 9307
rect 2922 9303 2926 9307
rect 2938 9303 2942 9309
rect 2983 9313 2987 9317
rect 2996 9316 3000 9322
rect 3033 9316 3037 9322
rect 3046 9318 3050 9322
rect 3070 9322 3074 9326
rect 3144 9322 3148 9326
rect 3054 9316 3058 9322
rect 3091 9316 3095 9322
rect 3107 9318 3111 9322
rect 2959 9303 2963 9307
rect 2975 9303 2979 9307
rect 2996 9303 3000 9307
rect 3012 9303 3016 9309
rect 3046 9309 3050 9313
rect 3033 9303 3037 9307
rect 3054 9303 3058 9307
rect 3070 9303 3074 9309
rect 3115 9313 3119 9317
rect 3128 9316 3132 9322
rect 3165 9316 3169 9322
rect 3178 9318 3182 9322
rect 3202 9322 3206 9326
rect 3276 9322 3280 9326
rect 3186 9316 3190 9322
rect 3223 9316 3227 9322
rect 3239 9318 3243 9322
rect 3091 9303 3095 9307
rect 3107 9303 3111 9307
rect 3128 9303 3132 9307
rect 3144 9303 3148 9309
rect 3178 9309 3182 9313
rect 3165 9303 3169 9307
rect 3186 9303 3190 9307
rect 3202 9303 3206 9309
rect 3247 9313 3251 9317
rect 3260 9316 3264 9322
rect 3297 9316 3301 9322
rect 3310 9318 3314 9322
rect 3334 9322 3338 9326
rect 3825 9322 3829 9326
rect 3318 9316 3322 9322
rect 3355 9316 3359 9322
rect 3371 9318 3375 9322
rect 3450 9314 3454 9318
rect 3486 9314 3490 9318
rect 3553 9314 3557 9318
rect 3769 9314 3775 9318
rect 3223 9303 3227 9307
rect 3239 9303 3243 9307
rect 3260 9303 3264 9307
rect 3276 9303 3280 9309
rect 3310 9309 3314 9313
rect 3297 9303 3301 9307
rect 2528 9289 2532 9293
rect 2490 9280 2494 9284
rect 2512 9283 2516 9289
rect 2549 9283 2553 9289
rect 2562 9285 2566 9289
rect 2586 9289 2590 9293
rect 2570 9283 2574 9289
rect 2607 9283 2611 9289
rect 2623 9283 2627 9289
rect 2857 9292 2861 9296
rect 2894 9290 2898 9294
rect 2914 9290 2918 9294
rect 2958 9290 2962 9294
rect 2989 9292 2993 9296
rect 3026 9290 3030 9294
rect 3046 9290 3050 9294
rect 3090 9290 3094 9294
rect 3121 9292 3125 9296
rect 3158 9290 3162 9294
rect 3178 9290 3182 9294
rect 3222 9290 3226 9294
rect 3239 9295 3243 9299
rect 3318 9303 3322 9307
rect 3334 9303 3338 9309
rect 3796 9313 3800 9317
rect 3809 9316 3813 9322
rect 3846 9316 3850 9322
rect 3859 9318 3863 9322
rect 3883 9322 3887 9326
rect 3957 9322 3961 9326
rect 3867 9316 3871 9322
rect 3904 9316 3908 9322
rect 3920 9318 3924 9322
rect 3709 9307 3715 9311
rect 3355 9303 3359 9307
rect 3371 9303 3375 9307
rect 3253 9292 3257 9296
rect 3290 9290 3294 9294
rect 3310 9290 3314 9294
rect 3354 9290 3358 9294
rect 3371 9295 3375 9299
rect 3450 9300 3454 9304
rect 3500 9300 3504 9304
rect 3553 9300 3557 9304
rect 3809 9303 3813 9307
rect 3825 9303 3829 9309
rect 3859 9309 3863 9313
rect 3846 9303 3850 9307
rect 3867 9303 3871 9307
rect 3883 9303 3887 9309
rect 3928 9313 3932 9317
rect 3941 9316 3945 9322
rect 3978 9316 3982 9322
rect 3991 9318 3995 9322
rect 4015 9322 4019 9326
rect 4089 9322 4093 9326
rect 3999 9316 4003 9322
rect 4036 9316 4040 9322
rect 4052 9318 4056 9322
rect 3904 9303 3908 9307
rect 3920 9303 3924 9307
rect 3941 9303 3945 9307
rect 3957 9303 3961 9309
rect 3991 9309 3995 9313
rect 3978 9303 3982 9307
rect 3999 9303 4003 9307
rect 4015 9303 4019 9309
rect 4060 9313 4064 9317
rect 4073 9316 4077 9322
rect 4110 9316 4114 9322
rect 4123 9318 4127 9322
rect 4147 9322 4151 9326
rect 4221 9322 4225 9326
rect 4131 9316 4135 9322
rect 4168 9316 4172 9322
rect 4184 9318 4188 9322
rect 4036 9303 4040 9307
rect 4052 9303 4056 9307
rect 4073 9303 4077 9307
rect 4089 9303 4093 9309
rect 4123 9309 4127 9313
rect 4110 9303 4114 9307
rect 4131 9303 4135 9307
rect 4147 9303 4151 9309
rect 4192 9313 4196 9317
rect 4205 9316 4209 9322
rect 4242 9316 4246 9322
rect 4255 9318 4259 9322
rect 4279 9322 4283 9326
rect 4263 9316 4267 9322
rect 4300 9316 4304 9322
rect 4316 9318 4320 9322
rect 4168 9303 4172 9307
rect 4184 9303 4188 9307
rect 4205 9303 4209 9307
rect 4221 9303 4225 9309
rect 4255 9309 4259 9313
rect 4242 9303 4246 9307
rect 3473 9289 3477 9293
rect 2776 9283 2782 9287
rect 2512 9270 2516 9274
rect 2528 9270 2532 9276
rect 2562 9276 2566 9280
rect 2549 9270 2553 9274
rect 2570 9270 2574 9274
rect 2586 9270 2590 9276
rect 3435 9280 3439 9284
rect 3457 9283 3461 9289
rect 3494 9283 3498 9289
rect 3507 9285 3511 9289
rect 3531 9289 3535 9293
rect 3515 9283 3519 9289
rect 3552 9283 3556 9289
rect 3568 9283 3572 9289
rect 3802 9292 3806 9296
rect 3839 9290 3843 9294
rect 3859 9290 3863 9294
rect 3903 9290 3907 9294
rect 3934 9292 3938 9296
rect 3971 9290 3975 9294
rect 3991 9290 3995 9294
rect 4035 9290 4039 9294
rect 4066 9292 4070 9296
rect 4103 9290 4107 9294
rect 4123 9290 4127 9294
rect 4167 9290 4171 9294
rect 4184 9295 4188 9299
rect 4263 9303 4267 9307
rect 4279 9303 4283 9309
rect 4300 9303 4304 9307
rect 4316 9303 4320 9307
rect 4198 9292 4202 9296
rect 4235 9290 4239 9294
rect 4255 9290 4259 9294
rect 4299 9290 4303 9294
rect 4316 9295 4320 9299
rect 3721 9283 3727 9287
rect 2812 9276 2818 9280
rect 2857 9276 2861 9280
rect 2908 9276 2912 9280
rect 2958 9276 2962 9280
rect 2989 9276 2993 9280
rect 3040 9276 3044 9280
rect 3090 9276 3094 9280
rect 3121 9276 3125 9280
rect 3172 9276 3176 9280
rect 3222 9276 3226 9280
rect 3253 9276 3257 9280
rect 3304 9276 3308 9280
rect 3354 9276 3358 9280
rect 2607 9270 2611 9274
rect 2623 9270 2627 9274
rect 3457 9270 3461 9274
rect 3473 9270 3477 9276
rect 3507 9276 3511 9280
rect 3494 9270 3498 9274
rect 2505 9259 2509 9263
rect 2542 9257 2546 9261
rect 2562 9257 2566 9261
rect 2606 9257 2610 9261
rect 2764 9263 2770 9267
rect 2855 9263 2859 9267
rect 2889 9263 2893 9267
rect 2906 9263 2910 9267
rect 2962 9263 2966 9267
rect 2979 9263 2983 9267
rect 3007 9263 3011 9267
rect 3515 9270 3519 9274
rect 3531 9270 3535 9276
rect 3757 9276 3763 9280
rect 3802 9276 3806 9280
rect 3853 9276 3857 9280
rect 3903 9276 3907 9280
rect 3934 9276 3938 9280
rect 3985 9276 3989 9280
rect 4035 9276 4039 9280
rect 4066 9276 4070 9280
rect 4117 9276 4121 9280
rect 4167 9276 4171 9280
rect 4198 9276 4202 9280
rect 4249 9276 4253 9280
rect 4299 9276 4303 9280
rect 3552 9270 3556 9274
rect 3568 9270 3572 9274
rect 2800 9256 2806 9260
rect 2882 9256 2886 9260
rect 2913 9256 2917 9260
rect 2935 9256 2939 9260
rect 3000 9256 3004 9260
rect 2776 9250 2782 9254
rect 2505 9243 2509 9247
rect 2556 9243 2560 9247
rect 2606 9243 2610 9247
rect 2812 9243 2818 9247
rect 2856 9246 2860 9250
rect 2881 9249 2885 9253
rect 2888 9246 2892 9250
rect 2906 9246 2910 9250
rect 2928 9249 2932 9253
rect 2953 9249 2957 9253
rect 2963 9246 2967 9250
rect 2979 9246 2983 9250
rect 2999 9249 3003 9253
rect 3006 9246 3010 9250
rect 3070 9256 3074 9260
rect 2623 9236 2627 9240
rect 2490 9227 2494 9231
rect 2615 9229 2619 9233
rect 2639 9229 2643 9233
rect 2498 9220 2502 9224
rect 2639 9220 2643 9224
rect 2883 9230 2887 9234
rect 2903 9227 2907 9231
rect 2922 9231 2926 9235
rect 3024 9242 3028 9246
rect 3039 9242 3043 9246
rect 2941 9230 2945 9234
rect 2960 9230 2964 9234
rect 2973 9229 2977 9233
rect 2995 9230 2999 9234
rect 3003 9229 3007 9233
rect 3015 9229 3019 9233
rect 2856 9216 2860 9220
rect 2888 9216 2892 9220
rect 2906 9216 2910 9220
rect 2963 9216 2967 9220
rect 2978 9216 2982 9220
rect 3006 9216 3010 9220
rect 2505 9212 2509 9216
rect 2572 9212 2576 9216
rect 2608 9212 2612 9216
rect 2824 9212 2830 9216
rect 2870 9212 2874 9216
rect 2913 9211 2917 9215
rect 2935 9212 2942 9216
rect 2985 9211 2989 9215
rect 2764 9205 2770 9209
rect 2505 9198 2509 9202
rect 2558 9198 2562 9202
rect 2608 9198 2612 9202
rect 2788 9204 2794 9208
rect 2870 9204 2874 9208
rect 2929 9204 2933 9208
rect 2954 9204 2958 9208
rect 2985 9204 2989 9208
rect 3078 9234 3082 9242
rect 3151 9256 3155 9260
rect 3105 9242 3109 9246
rect 3120 9242 3124 9246
rect 3101 9234 3105 9238
rect 3047 9228 3051 9232
rect 3060 9220 3064 9224
rect 3159 9234 3163 9242
rect 3321 9250 3328 9258
rect 3411 9250 3416 9258
rect 3450 9259 3454 9263
rect 3487 9257 3491 9261
rect 3507 9257 3511 9261
rect 3551 9257 3555 9261
rect 3709 9263 3715 9267
rect 3800 9263 3804 9267
rect 3834 9263 3838 9267
rect 3851 9263 3855 9267
rect 3907 9263 3911 9267
rect 3924 9263 3928 9267
rect 3952 9263 3956 9267
rect 3745 9256 3751 9260
rect 3827 9256 3831 9260
rect 3858 9256 3862 9260
rect 3880 9256 3884 9260
rect 3945 9256 3949 9260
rect 3721 9250 3727 9254
rect 3361 9241 3365 9245
rect 3423 9241 3427 9245
rect 3450 9243 3454 9247
rect 3501 9243 3505 9247
rect 3551 9243 3555 9247
rect 3757 9243 3763 9247
rect 3801 9246 3805 9250
rect 3826 9249 3830 9253
rect 3833 9246 3837 9250
rect 3851 9246 3855 9250
rect 3873 9249 3877 9253
rect 3898 9249 3902 9253
rect 3908 9246 3912 9250
rect 3924 9246 3928 9250
rect 3944 9249 3948 9253
rect 3951 9246 3955 9250
rect 4015 9256 4019 9260
rect 3186 9234 3190 9238
rect 3568 9236 3572 9240
rect 3128 9228 3132 9232
rect 3435 9227 3439 9231
rect 3560 9229 3564 9233
rect 3584 9229 3588 9233
rect 3141 9220 3145 9224
rect 3443 9220 3447 9224
rect 3584 9220 3588 9224
rect 3828 9230 3832 9234
rect 3848 9227 3852 9231
rect 3867 9231 3871 9235
rect 3969 9242 3973 9246
rect 3984 9242 3988 9246
rect 3886 9230 3890 9234
rect 3905 9230 3909 9234
rect 3918 9229 3922 9233
rect 3940 9230 3944 9234
rect 3948 9229 3952 9233
rect 3960 9229 3964 9233
rect 3801 9216 3805 9220
rect 3833 9216 3837 9220
rect 3851 9216 3855 9220
rect 3908 9216 3912 9220
rect 3923 9216 3927 9220
rect 3951 9216 3955 9220
rect 3450 9212 3454 9216
rect 3517 9212 3521 9216
rect 3553 9212 3557 9216
rect 3769 9212 3775 9216
rect 3815 9212 3819 9216
rect 3858 9211 3862 9215
rect 3880 9212 3887 9216
rect 3930 9211 3934 9215
rect 3709 9205 3715 9209
rect 2776 9197 2782 9201
rect 2856 9197 2860 9201
rect 2870 9197 2874 9201
rect 2888 9197 2892 9201
rect 2906 9197 2910 9201
rect 2929 9197 2933 9201
rect 2963 9197 2967 9201
rect 2978 9197 2982 9201
rect 3006 9197 3010 9201
rect 2527 9187 2531 9191
rect 2490 9181 2494 9187
rect 2506 9181 2510 9187
rect 2543 9181 2547 9187
rect 2551 9183 2555 9187
rect 2585 9187 2589 9191
rect 2788 9190 2794 9194
rect 2870 9190 2874 9194
rect 2929 9190 2933 9194
rect 2954 9190 2958 9194
rect 2985 9190 2989 9194
rect 2564 9181 2568 9187
rect 2601 9181 2605 9187
rect 2870 9182 2874 9186
rect 2913 9183 2917 9187
rect 2935 9182 2942 9186
rect 2985 9183 2989 9187
rect 2623 9178 2627 9182
rect 2856 9178 2860 9182
rect 2888 9178 2892 9182
rect 2906 9178 2910 9182
rect 2963 9178 2967 9182
rect 2978 9178 2982 9182
rect 3006 9178 3010 9182
rect 2490 9168 2494 9172
rect 2506 9168 2510 9172
rect 2551 9174 2555 9178
rect 2527 9168 2531 9174
rect 2543 9168 2547 9172
rect 2564 9168 2568 9172
rect 2585 9168 2589 9174
rect 2601 9168 2605 9172
rect 2851 9166 2855 9170
rect 2507 9155 2511 9159
rect 2551 9155 2555 9159
rect 2571 9155 2575 9159
rect 2608 9157 2612 9161
rect 2883 9164 2887 9168
rect 2903 9167 2907 9171
rect 2922 9163 2926 9167
rect 2941 9164 2945 9168
rect 2960 9164 2964 9168
rect 2973 9165 2977 9169
rect 3070 9180 3074 9184
rect 3450 9198 3454 9202
rect 3503 9198 3507 9202
rect 3553 9198 3557 9202
rect 3733 9204 3739 9208
rect 3815 9204 3819 9208
rect 3874 9204 3878 9208
rect 3899 9204 3903 9208
rect 3930 9204 3934 9208
rect 4023 9234 4027 9242
rect 4096 9256 4100 9260
rect 4050 9242 4054 9246
rect 4065 9242 4069 9246
rect 4046 9234 4050 9238
rect 3992 9228 3996 9232
rect 4005 9220 4009 9224
rect 4104 9234 4108 9242
rect 4131 9234 4135 9238
rect 4073 9228 4077 9232
rect 4086 9220 4090 9224
rect 3721 9197 3727 9201
rect 3801 9197 3805 9201
rect 3815 9197 3819 9201
rect 3833 9197 3837 9201
rect 3851 9197 3855 9201
rect 3874 9197 3878 9201
rect 3908 9197 3912 9201
rect 3923 9197 3927 9201
rect 3951 9197 3955 9201
rect 3472 9187 3476 9191
rect 3151 9180 3155 9184
rect 3435 9181 3439 9187
rect 3451 9181 3455 9187
rect 3488 9181 3492 9187
rect 3496 9183 3500 9187
rect 3530 9187 3534 9191
rect 3733 9190 3739 9194
rect 3815 9190 3819 9194
rect 3874 9190 3878 9194
rect 3899 9190 3903 9194
rect 3930 9190 3934 9194
rect 3509 9181 3513 9187
rect 3546 9181 3550 9187
rect 3815 9182 3819 9186
rect 3858 9183 3862 9187
rect 3880 9182 3887 9186
rect 3930 9183 3934 9187
rect 3568 9178 3572 9182
rect 3801 9178 3805 9182
rect 3833 9178 3837 9182
rect 3851 9178 3855 9182
rect 3908 9178 3912 9182
rect 3923 9178 3927 9182
rect 3951 9178 3955 9182
rect 2995 9164 2999 9168
rect 3003 9165 3007 9169
rect 3015 9165 3019 9169
rect 3050 9165 3054 9169
rect 3078 9164 3082 9168
rect 3130 9165 3134 9169
rect 3435 9168 3439 9172
rect 3451 9168 3455 9172
rect 3496 9174 3500 9178
rect 3472 9168 3476 9174
rect 3488 9168 3492 9172
rect 3159 9164 3163 9168
rect 3509 9168 3513 9172
rect 3530 9168 3534 9174
rect 3546 9168 3550 9172
rect 3796 9166 3800 9170
rect 2776 9148 2782 9152
rect 2856 9148 2860 9152
rect 2881 9145 2885 9149
rect 2888 9148 2892 9152
rect 2906 9148 2910 9152
rect 2928 9145 2932 9149
rect 2953 9145 2957 9149
rect 2963 9148 2967 9152
rect 2979 9148 2983 9152
rect 2999 9145 3003 9149
rect 3006 9148 3010 9152
rect 2507 9141 2511 9145
rect 2557 9141 2561 9145
rect 2608 9141 2612 9145
rect 2812 9141 2818 9145
rect 2866 9138 2870 9142
rect 2882 9138 2886 9142
rect 2913 9138 2917 9142
rect 2935 9138 2939 9142
rect 3000 9138 3004 9142
rect 3060 9144 3064 9148
rect 3452 9155 3456 9159
rect 3496 9155 3500 9159
rect 3516 9155 3520 9159
rect 3553 9157 3557 9161
rect 3828 9164 3832 9168
rect 3848 9167 3852 9171
rect 3867 9163 3871 9167
rect 3886 9164 3890 9168
rect 3905 9164 3909 9168
rect 3918 9165 3922 9169
rect 4015 9180 4019 9184
rect 4096 9180 4100 9184
rect 3940 9164 3944 9168
rect 3948 9165 3952 9169
rect 3960 9165 3964 9169
rect 3995 9165 3999 9169
rect 4023 9164 4027 9168
rect 4075 9165 4079 9169
rect 4104 9164 4108 9168
rect 3721 9148 3727 9152
rect 3801 9148 3805 9152
rect 3141 9144 3145 9148
rect 3826 9145 3830 9149
rect 3833 9148 3837 9152
rect 3851 9148 3855 9152
rect 3873 9145 3877 9149
rect 3898 9145 3902 9149
rect 3908 9148 3912 9152
rect 3924 9148 3928 9152
rect 3944 9145 3948 9149
rect 3951 9148 3955 9152
rect 3452 9141 3456 9145
rect 3502 9141 3506 9145
rect 3553 9141 3557 9145
rect 3757 9141 3763 9145
rect 3811 9138 3815 9142
rect 3827 9138 3831 9142
rect 3858 9138 3862 9142
rect 3880 9138 3884 9142
rect 3945 9138 3949 9142
rect 4005 9144 4009 9148
rect 4086 9144 4090 9148
rect 2764 9131 2770 9135
rect 2855 9131 2859 9135
rect 2889 9131 2893 9135
rect 2906 9131 2910 9135
rect 2962 9131 2966 9135
rect 2979 9131 2983 9135
rect 3007 9131 3011 9135
rect 3709 9131 3715 9135
rect 3800 9131 3804 9135
rect 3834 9131 3838 9135
rect 3851 9131 3855 9135
rect 3907 9131 3911 9135
rect 3924 9131 3928 9135
rect 3952 9131 3956 9135
rect 2800 9124 2806 9128
rect 2866 9124 2870 9128
rect 2882 9124 2886 9128
rect 2913 9124 2917 9128
rect 2935 9124 2939 9128
rect 3000 9124 3004 9128
rect 3070 9124 3074 9128
rect 2856 9114 2860 9118
rect 2881 9117 2885 9121
rect 2888 9114 2892 9118
rect 2906 9114 2910 9118
rect 2928 9117 2932 9121
rect 2953 9117 2957 9121
rect 2963 9114 2967 9118
rect 2979 9114 2983 9118
rect 2999 9117 3003 9121
rect 3006 9114 3010 9118
rect 2850 9097 2854 9101
rect 2883 9098 2887 9102
rect 2903 9095 2907 9099
rect 2922 9099 2926 9103
rect 2941 9098 2945 9102
rect 2960 9098 2964 9102
rect 2973 9097 2977 9101
rect 2995 9098 2999 9102
rect 3003 9097 3007 9101
rect 3015 9097 3019 9101
rect 3078 9102 3082 9110
rect 3175 9124 3179 9128
rect 3129 9110 3133 9114
rect 3144 9110 3148 9114
rect 3361 9120 3365 9124
rect 3745 9124 3751 9128
rect 3811 9124 3815 9128
rect 3827 9124 3831 9128
rect 3858 9124 3862 9128
rect 3880 9124 3884 9128
rect 3945 9124 3949 9128
rect 4015 9124 4019 9128
rect 3047 9096 3051 9100
rect 3101 9101 3105 9105
rect 2856 9084 2860 9088
rect 2888 9084 2892 9088
rect 2906 9084 2910 9088
rect 2963 9084 2967 9088
rect 2978 9084 2982 9088
rect 3006 9084 3010 9088
rect 2870 9080 2874 9084
rect 2913 9079 2917 9083
rect 2935 9080 2942 9084
rect 2985 9079 2989 9083
rect 2788 9072 2794 9076
rect 2870 9072 2874 9076
rect 2929 9072 2933 9076
rect 2954 9072 2958 9076
rect 2985 9072 2989 9076
rect 3060 9088 3064 9092
rect 3183 9102 3187 9110
rect 3801 9114 3805 9118
rect 3826 9117 3830 9121
rect 3833 9114 3837 9118
rect 3851 9114 3855 9118
rect 3873 9117 3877 9121
rect 3898 9117 3902 9121
rect 3908 9114 3912 9118
rect 3924 9114 3928 9118
rect 3944 9117 3948 9121
rect 3951 9114 3955 9118
rect 3204 9102 3208 9106
rect 3668 9102 3672 9106
rect 3152 9096 3156 9100
rect 3165 9088 3169 9092
rect 3406 9095 3410 9099
rect 3360 9081 3364 9085
rect 3375 9081 3379 9085
rect 3383 9073 3387 9077
rect 3414 9073 3418 9081
rect 3795 9097 3799 9101
rect 2776 9065 2782 9069
rect 2856 9065 2860 9069
rect 2870 9065 2874 9069
rect 2888 9065 2892 9069
rect 2906 9065 2910 9069
rect 2929 9065 2933 9069
rect 2963 9065 2967 9069
rect 2978 9065 2982 9069
rect 3006 9065 3010 9069
rect 2788 9058 2794 9062
rect 2870 9058 2874 9062
rect 2929 9058 2933 9062
rect 2954 9058 2958 9062
rect 2985 9058 2989 9062
rect 2870 9050 2874 9054
rect 2913 9051 2917 9055
rect 2935 9050 2942 9054
rect 2985 9051 2989 9055
rect 2856 9046 2860 9050
rect 2888 9046 2892 9050
rect 2906 9046 2910 9050
rect 2963 9046 2967 9050
rect 2978 9046 2982 9050
rect 3006 9046 3010 9050
rect 3070 9049 3074 9053
rect 3175 9049 3179 9053
rect 2851 9034 2855 9038
rect 2883 9032 2887 9036
rect 2903 9035 2907 9039
rect 2922 9031 2926 9035
rect 2941 9032 2945 9036
rect 2960 9032 2964 9036
rect 2973 9033 2977 9037
rect 2995 9032 2999 9036
rect 3003 9033 3007 9037
rect 3015 9033 3019 9037
rect 3049 9034 3053 9038
rect 3078 9033 3082 9037
rect 3155 9034 3159 9038
rect 3183 9033 3187 9037
rect 3396 9059 3400 9063
rect 3828 9098 3832 9102
rect 3848 9095 3852 9099
rect 3867 9099 3871 9103
rect 3886 9098 3890 9102
rect 3905 9098 3909 9102
rect 3918 9097 3922 9101
rect 3940 9098 3944 9102
rect 3948 9097 3952 9101
rect 3960 9097 3964 9101
rect 4023 9102 4027 9110
rect 4120 9124 4124 9128
rect 4074 9110 4078 9114
rect 4089 9110 4093 9114
rect 3992 9096 3996 9100
rect 4046 9101 4050 9105
rect 3801 9084 3805 9088
rect 3833 9084 3837 9088
rect 3851 9084 3855 9088
rect 3908 9084 3912 9088
rect 3923 9084 3927 9088
rect 3951 9084 3955 9088
rect 3815 9080 3819 9084
rect 3858 9079 3862 9083
rect 3880 9080 3887 9084
rect 3930 9079 3934 9083
rect 3733 9072 3739 9076
rect 3815 9072 3819 9076
rect 3874 9072 3878 9076
rect 3899 9072 3903 9076
rect 3930 9072 3934 9076
rect 4005 9088 4009 9092
rect 4128 9102 4132 9110
rect 4149 9102 4153 9106
rect 4097 9096 4101 9100
rect 4110 9088 4114 9092
rect 3721 9065 3727 9069
rect 3801 9065 3805 9069
rect 3815 9065 3819 9069
rect 3833 9065 3837 9069
rect 3851 9065 3855 9069
rect 3874 9065 3878 9069
rect 3908 9065 3912 9069
rect 3923 9065 3927 9069
rect 3951 9065 3955 9069
rect 3593 9053 3597 9057
rect 3733 9058 3739 9062
rect 3815 9058 3819 9062
rect 3874 9058 3878 9062
rect 3899 9058 3903 9062
rect 3930 9058 3934 9062
rect 3815 9050 3819 9054
rect 3858 9051 3862 9055
rect 3880 9050 3887 9054
rect 3930 9051 3934 9055
rect 3626 9045 3630 9049
rect 3745 9045 3751 9049
rect 3801 9046 3805 9050
rect 3833 9046 3837 9050
rect 3851 9046 3855 9050
rect 3908 9046 3912 9050
rect 3923 9046 3927 9050
rect 3951 9046 3955 9050
rect 4015 9049 4019 9053
rect 4484 9056 4488 9060
rect 4494 9056 4498 9060
rect 4504 9056 4508 9060
rect 4120 9049 4124 9053
rect 4484 9051 4488 9055
rect 4494 9051 4498 9055
rect 4504 9051 4508 9055
rect 4484 9046 4488 9050
rect 4494 9046 4498 9050
rect 4504 9046 4508 9050
rect 3668 9033 3672 9037
rect 3709 9033 3715 9037
rect 3796 9034 3800 9038
rect 3721 9026 3727 9030
rect 3660 9022 3665 9026
rect 2856 9016 2860 9020
rect 618 9012 622 9016
rect 628 9012 632 9016
rect 638 9012 642 9016
rect 618 9007 622 9011
rect 628 9007 632 9011
rect 638 9007 642 9011
rect 618 9002 622 9006
rect 628 9002 632 9006
rect 638 9002 642 9006
rect 618 8997 622 9001
rect 628 8997 632 9001
rect 638 8997 642 9001
rect 664 9012 668 9016
rect 674 9012 678 9016
rect 684 9012 688 9016
rect 2881 9013 2885 9017
rect 2888 9016 2892 9020
rect 2906 9016 2910 9020
rect 2928 9013 2932 9017
rect 2953 9013 2957 9017
rect 2963 9016 2967 9020
rect 2979 9016 2983 9020
rect 2999 9013 3003 9017
rect 3006 9016 3010 9020
rect 664 9007 668 9011
rect 674 9007 678 9011
rect 684 9007 688 9011
rect 2800 9006 2806 9010
rect 2882 9006 2886 9010
rect 2913 9006 2917 9010
rect 2935 9006 2939 9010
rect 3000 9006 3004 9010
rect 664 9002 668 9006
rect 674 9002 678 9006
rect 684 9002 688 9006
rect 3060 9013 3064 9017
rect 3165 9013 3169 9017
rect 3406 9015 3410 9019
rect 3676 9017 3680 9021
rect 3781 9017 3787 9021
rect 3828 9032 3832 9036
rect 3848 9035 3852 9039
rect 3867 9031 3871 9035
rect 3886 9032 3890 9036
rect 3905 9032 3909 9036
rect 3918 9033 3922 9037
rect 3940 9032 3944 9036
rect 3948 9033 3952 9037
rect 3960 9033 3964 9037
rect 3994 9034 3998 9038
rect 4023 9033 4027 9037
rect 4100 9034 4104 9038
rect 4484 9041 4488 9045
rect 4494 9041 4498 9045
rect 4504 9041 4508 9045
rect 4530 9056 4534 9060
rect 4540 9056 4544 9060
rect 4550 9056 4554 9060
rect 4530 9051 4534 9055
rect 4540 9051 4544 9055
rect 4550 9051 4554 9055
rect 4530 9046 4534 9050
rect 4540 9046 4544 9050
rect 4550 9046 4554 9050
rect 4530 9041 4534 9045
rect 4540 9041 4544 9045
rect 4550 9041 4554 9045
rect 4128 9033 4132 9037
rect 3801 9016 3805 9020
rect 3826 9013 3830 9017
rect 3833 9016 3837 9020
rect 3851 9016 3855 9020
rect 3873 9013 3877 9017
rect 3898 9013 3902 9017
rect 3908 9016 3912 9020
rect 3924 9016 3928 9020
rect 3944 9013 3948 9017
rect 3951 9016 3955 9020
rect 3593 9008 3598 9012
rect 3733 9008 3739 9012
rect 664 8997 668 9001
rect 674 8997 678 9001
rect 684 8997 688 9001
rect 2764 8999 2770 9003
rect 2855 8999 2859 9003
rect 2889 8999 2893 9003
rect 2906 8999 2910 9003
rect 2962 8999 2966 9003
rect 2979 8999 2983 9003
rect 3007 8999 3011 9003
rect 3326 9000 3330 9004
rect 3745 9006 3751 9010
rect 3827 9006 3831 9010
rect 3858 9006 3862 9010
rect 3880 9006 3884 9010
rect 3945 9006 3949 9010
rect 4005 9013 4009 9017
rect 4110 9013 4114 9017
rect 3414 8999 3418 9003
rect 3709 8999 3715 9003
rect 3800 8999 3804 9003
rect 3834 8999 3838 9003
rect 3851 8999 3855 9003
rect 3907 8999 3911 9003
rect 3924 8999 3928 9003
rect 3952 8999 3956 9003
rect 2800 8992 2806 8996
rect 2882 8992 2886 8996
rect 2913 8992 2917 8996
rect 2935 8992 2939 8996
rect 3000 8992 3004 8996
rect 3070 8992 3074 8996
rect 2856 8982 2860 8986
rect 2881 8985 2885 8989
rect 2888 8982 2892 8986
rect 2906 8982 2910 8986
rect 2928 8985 2932 8989
rect 2953 8985 2957 8989
rect 2963 8982 2967 8986
rect 2979 8982 2983 8986
rect 2999 8985 3003 8989
rect 3006 8982 3010 8986
rect 2850 8965 2854 8969
rect 2883 8966 2887 8970
rect 2903 8963 2907 8967
rect 2922 8967 2926 8971
rect 2941 8966 2945 8970
rect 2960 8966 2964 8970
rect 2973 8965 2977 8969
rect 2995 8966 2999 8970
rect 3003 8965 3007 8969
rect 3015 8965 3019 8969
rect 3078 8970 3082 8978
rect 3151 8992 3155 8996
rect 3105 8978 3109 8982
rect 3120 8978 3124 8982
rect 3101 8970 3105 8974
rect 3047 8964 3051 8968
rect 2856 8952 2860 8956
rect 2888 8952 2892 8956
rect 2906 8952 2910 8956
rect 2963 8952 2967 8956
rect 2978 8952 2982 8956
rect 3006 8952 3010 8956
rect 2870 8948 2874 8952
rect 2913 8947 2917 8951
rect 2935 8948 2942 8952
rect 2985 8947 2989 8951
rect 2788 8940 2794 8944
rect 2870 8940 2874 8944
rect 2929 8940 2933 8944
rect 2954 8940 2958 8944
rect 2985 8940 2989 8944
rect 3060 8956 3064 8960
rect 3159 8970 3163 8978
rect 3241 8992 3245 8996
rect 3195 8978 3199 8982
rect 3210 8978 3214 8982
rect 3183 8970 3187 8974
rect 3128 8964 3132 8968
rect 3217 8972 3221 8976
rect 3249 8970 3253 8978
rect 3745 8992 3751 8996
rect 3827 8992 3831 8996
rect 3858 8992 3862 8996
rect 3880 8992 3884 8996
rect 3945 8992 3949 8996
rect 4015 8992 4019 8996
rect 3396 8979 3400 8983
rect 3801 8982 3805 8986
rect 3826 8985 3830 8989
rect 3833 8982 3837 8986
rect 3851 8982 3855 8986
rect 3873 8985 3877 8989
rect 3898 8985 3902 8989
rect 3908 8982 3912 8986
rect 3924 8982 3928 8986
rect 3944 8985 3948 8989
rect 3951 8982 3955 8986
rect 3141 8956 3145 8960
rect 3284 8969 3288 8973
rect 3668 8972 3672 8976
rect 3231 8956 3235 8960
rect 3406 8965 3410 8969
rect 3338 8951 3342 8955
rect 3353 8951 3357 8955
rect 3360 8951 3364 8955
rect 3375 8951 3379 8955
rect 3383 8943 3387 8947
rect 3414 8943 3418 8951
rect 3795 8965 3799 8969
rect 2776 8933 2782 8937
rect 2856 8933 2860 8937
rect 2870 8933 2874 8937
rect 2888 8933 2892 8937
rect 2906 8933 2910 8937
rect 2929 8933 2933 8937
rect 2963 8933 2967 8937
rect 2978 8933 2982 8937
rect 3006 8933 3010 8937
rect 2788 8926 2794 8930
rect 2870 8926 2874 8930
rect 2929 8926 2933 8930
rect 2954 8926 2958 8930
rect 2985 8926 2989 8930
rect 2870 8918 2874 8922
rect 2913 8919 2917 8923
rect 2935 8918 2942 8922
rect 2985 8919 2989 8923
rect 2856 8914 2860 8918
rect 2888 8914 2892 8918
rect 2906 8914 2910 8918
rect 2963 8914 2967 8918
rect 2978 8914 2982 8918
rect 3006 8914 3010 8918
rect 2851 8902 2855 8906
rect 2883 8900 2887 8904
rect 2903 8903 2907 8907
rect 2922 8899 2926 8903
rect 2941 8900 2945 8904
rect 2960 8900 2964 8904
rect 2973 8901 2977 8905
rect 3070 8914 3074 8918
rect 3151 8914 3155 8918
rect 3241 8914 3245 8918
rect 2995 8900 2999 8904
rect 3003 8901 3007 8905
rect 3015 8901 3019 8905
rect 3050 8899 3054 8903
rect 3078 8898 3082 8902
rect 3130 8899 3134 8903
rect 3159 8898 3163 8902
rect 3214 8899 3218 8903
rect 3249 8898 3253 8902
rect 3396 8929 3400 8933
rect 3828 8966 3832 8970
rect 3848 8963 3852 8967
rect 3867 8967 3871 8971
rect 3886 8966 3890 8970
rect 3905 8966 3909 8970
rect 3918 8965 3922 8969
rect 3940 8966 3944 8970
rect 3948 8965 3952 8969
rect 3960 8965 3964 8969
rect 4023 8970 4027 8978
rect 4096 8992 4100 8996
rect 4050 8978 4054 8982
rect 4065 8978 4069 8982
rect 4046 8970 4050 8974
rect 3992 8964 3996 8968
rect 3801 8952 3805 8956
rect 3833 8952 3837 8956
rect 3851 8952 3855 8956
rect 3908 8952 3912 8956
rect 3923 8952 3927 8956
rect 3951 8952 3955 8956
rect 3815 8948 3819 8952
rect 3858 8947 3862 8951
rect 3880 8948 3887 8952
rect 3930 8947 3934 8951
rect 3733 8940 3739 8944
rect 3815 8940 3819 8944
rect 3874 8940 3878 8944
rect 3899 8940 3903 8944
rect 3930 8940 3934 8944
rect 4005 8956 4009 8960
rect 4104 8970 4108 8978
rect 4186 8992 4190 8996
rect 4140 8978 4144 8982
rect 4155 8978 4159 8982
rect 4128 8970 4132 8974
rect 4073 8964 4077 8968
rect 4162 8972 4166 8976
rect 4194 8970 4198 8978
rect 4086 8956 4090 8960
rect 4229 8969 4233 8973
rect 4176 8956 4180 8960
rect 3488 8923 3492 8927
rect 3721 8933 3727 8937
rect 3801 8933 3805 8937
rect 3815 8933 3819 8937
rect 3833 8933 3837 8937
rect 3851 8933 3855 8937
rect 3874 8933 3878 8937
rect 3908 8933 3912 8937
rect 3923 8933 3927 8937
rect 3951 8933 3955 8937
rect 3733 8926 3739 8930
rect 3815 8926 3819 8930
rect 3874 8926 3878 8930
rect 3899 8926 3903 8930
rect 3930 8926 3934 8930
rect 3532 8915 3536 8919
rect 3815 8918 3819 8922
rect 3858 8919 3862 8923
rect 3880 8918 3887 8922
rect 3930 8919 3934 8923
rect 3769 8912 3775 8916
rect 3801 8914 3805 8918
rect 3833 8914 3837 8918
rect 3851 8914 3855 8918
rect 3908 8914 3912 8918
rect 3923 8914 3927 8918
rect 3951 8914 3955 8918
rect 3796 8902 3800 8906
rect 2856 8884 2860 8888
rect 2881 8881 2885 8885
rect 2888 8884 2892 8888
rect 2906 8884 2910 8888
rect 2928 8881 2932 8885
rect 2953 8881 2957 8885
rect 2963 8884 2967 8888
rect 2979 8884 2983 8888
rect 2999 8881 3003 8885
rect 3006 8884 3010 8888
rect 3660 8892 3665 8896
rect 2800 8874 2806 8878
rect 2882 8874 2886 8878
rect 2913 8874 2917 8878
rect 2935 8874 2939 8878
rect 3000 8874 3004 8878
rect 3060 8878 3064 8882
rect 3141 8878 3145 8882
rect 3406 8885 3410 8889
rect 3828 8900 3832 8904
rect 3848 8903 3852 8907
rect 3867 8899 3871 8903
rect 3886 8900 3890 8904
rect 3905 8900 3909 8904
rect 3918 8901 3922 8905
rect 4015 8914 4019 8918
rect 4096 8914 4100 8918
rect 4186 8914 4190 8918
rect 3940 8900 3944 8904
rect 3948 8901 3952 8905
rect 3960 8901 3964 8905
rect 3995 8899 3999 8903
rect 4023 8898 4027 8902
rect 4075 8899 4079 8903
rect 4104 8898 4108 8902
rect 4159 8899 4163 8903
rect 4194 8898 4198 8902
rect 3488 8882 3492 8886
rect 3757 8882 3763 8886
rect 3801 8884 3805 8888
rect 3231 8878 3235 8882
rect 3826 8881 3830 8885
rect 3833 8884 3837 8888
rect 3851 8884 3855 8888
rect 3873 8881 3877 8885
rect 3898 8881 3902 8885
rect 3908 8884 3912 8888
rect 3924 8884 3928 8888
rect 3944 8881 3948 8885
rect 3951 8884 3955 8888
rect 2764 8867 2770 8871
rect 2855 8867 2859 8871
rect 2889 8867 2893 8871
rect 2906 8867 2910 8871
rect 2962 8867 2966 8871
rect 2979 8867 2983 8871
rect 3007 8867 3011 8871
rect 3328 8870 3332 8874
rect 3745 8874 3751 8878
rect 3827 8874 3831 8878
rect 3858 8874 3862 8878
rect 3880 8874 3884 8878
rect 3945 8874 3949 8878
rect 3414 8869 3418 8873
rect 4005 8878 4009 8882
rect 4086 8878 4090 8882
rect 4176 8878 4180 8882
rect 2800 8860 2806 8864
rect 2882 8860 2886 8864
rect 2913 8860 2917 8864
rect 2935 8860 2939 8864
rect 3000 8860 3004 8864
rect 3070 8860 3074 8864
rect 3709 8867 3715 8871
rect 3800 8867 3804 8871
rect 3834 8867 3838 8871
rect 3851 8867 3855 8871
rect 3907 8867 3911 8871
rect 3924 8867 3928 8871
rect 3952 8867 3956 8871
rect 2856 8850 2860 8854
rect 2881 8853 2885 8857
rect 2888 8850 2892 8854
rect 2906 8850 2910 8854
rect 2928 8853 2932 8857
rect 2953 8853 2957 8857
rect 2963 8850 2967 8854
rect 2979 8850 2983 8854
rect 2999 8853 3003 8857
rect 3006 8850 3010 8854
rect 2850 8833 2854 8837
rect 2883 8834 2887 8838
rect 2903 8831 2907 8835
rect 2922 8835 2926 8839
rect 2941 8834 2945 8838
rect 2960 8834 2964 8838
rect 2973 8833 2977 8837
rect 2995 8834 2999 8838
rect 3003 8833 3007 8837
rect 3015 8833 3019 8837
rect 3078 8838 3082 8846
rect 3745 8860 3751 8864
rect 3827 8860 3831 8864
rect 3858 8860 3862 8864
rect 3880 8860 3884 8864
rect 3945 8860 3949 8864
rect 4015 8860 4019 8864
rect 3396 8849 3400 8853
rect 3801 8850 3805 8854
rect 3826 8853 3830 8857
rect 3833 8850 3837 8854
rect 3851 8850 3855 8854
rect 3873 8853 3877 8857
rect 3898 8853 3902 8857
rect 3908 8850 3912 8854
rect 3924 8850 3928 8854
rect 3944 8853 3948 8857
rect 3951 8850 3955 8854
rect 3668 8842 3672 8846
rect 3047 8832 3051 8836
rect 3101 8837 3105 8841
rect 3795 8833 3799 8837
rect 2351 8819 2355 8823
rect 2476 8819 2480 8823
rect 2856 8820 2860 8824
rect 2888 8820 2892 8824
rect 2906 8820 2910 8824
rect 2963 8820 2967 8824
rect 2978 8820 2982 8824
rect 3006 8820 3010 8824
rect 2870 8816 2874 8820
rect 2373 8812 2377 8816
rect 2409 8812 2413 8816
rect 2476 8812 2480 8816
rect 2505 8812 2509 8816
rect 2541 8812 2545 8816
rect 2608 8812 2612 8816
rect 2637 8812 2641 8816
rect 2673 8812 2677 8816
rect 2740 8812 2744 8816
rect 2824 8812 2830 8816
rect 2913 8815 2917 8819
rect 2935 8816 2942 8820
rect 2985 8815 2989 8819
rect 2764 8805 2770 8809
rect 2870 8808 2874 8812
rect 2879 8808 2883 8812
rect 2929 8808 2933 8812
rect 2954 8808 2958 8812
rect 2985 8808 2989 8812
rect 3060 8824 3064 8828
rect 3828 8834 3832 8838
rect 3848 8831 3852 8835
rect 3867 8835 3871 8839
rect 3886 8834 3890 8838
rect 3905 8834 3909 8838
rect 3918 8833 3922 8837
rect 3940 8834 3944 8838
rect 3948 8833 3952 8837
rect 3960 8833 3964 8837
rect 4023 8838 4027 8846
rect 3992 8832 3996 8836
rect 4046 8837 4050 8841
rect 3801 8820 3805 8824
rect 3833 8820 3837 8824
rect 3851 8820 3855 8824
rect 3908 8820 3912 8824
rect 3923 8820 3927 8824
rect 3951 8820 3955 8824
rect 3815 8816 3819 8820
rect 3318 8812 3322 8816
rect 3354 8812 3358 8816
rect 3421 8812 3425 8816
rect 3450 8812 3454 8816
rect 3486 8812 3490 8816
rect 3553 8812 3557 8816
rect 3582 8812 3586 8816
rect 3618 8812 3622 8816
rect 3685 8812 3689 8816
rect 3769 8812 3775 8816
rect 3858 8815 3862 8819
rect 3880 8816 3887 8820
rect 3930 8815 3934 8819
rect 3709 8805 3715 8809
rect 3815 8808 3819 8812
rect 3824 8808 3828 8812
rect 3874 8808 3878 8812
rect 3899 8808 3903 8812
rect 3930 8808 3934 8812
rect 4005 8824 4009 8828
rect 2373 8798 2377 8802
rect 2423 8798 2427 8802
rect 2476 8798 2480 8802
rect 2505 8798 2509 8802
rect 2555 8798 2559 8802
rect 2608 8798 2612 8802
rect 2637 8798 2641 8802
rect 2687 8798 2691 8802
rect 2740 8798 2744 8802
rect 2776 8801 2782 8805
rect 2856 8801 2860 8805
rect 2870 8801 2874 8805
rect 2888 8801 2892 8805
rect 2906 8801 2910 8805
rect 2929 8801 2933 8805
rect 2963 8801 2967 8805
rect 2978 8801 2982 8805
rect 3006 8801 3010 8805
rect 3131 8801 3135 8805
rect 3149 8801 3153 8805
rect 3167 8801 3171 8805
rect 3190 8801 3194 8805
rect 3224 8801 3228 8805
rect 3239 8801 3243 8805
rect 3267 8801 3271 8805
rect 2396 8787 2400 8791
rect 2351 8778 2355 8782
rect 2380 8781 2384 8787
rect 2417 8781 2421 8787
rect 2430 8783 2434 8787
rect 2454 8787 2458 8791
rect 2528 8787 2532 8791
rect 2438 8781 2442 8787
rect 2475 8781 2479 8787
rect 2491 8781 2495 8787
rect 2512 8781 2516 8787
rect 2549 8781 2553 8787
rect 2562 8783 2566 8787
rect 2586 8787 2590 8791
rect 2660 8787 2664 8791
rect 2570 8781 2574 8787
rect 2607 8781 2611 8787
rect 2623 8781 2627 8787
rect 2644 8781 2648 8787
rect 2681 8781 2685 8787
rect 2694 8783 2698 8787
rect 2718 8787 2722 8791
rect 2788 8794 2794 8798
rect 2870 8794 2874 8798
rect 2879 8794 2883 8798
rect 2929 8794 2933 8798
rect 2954 8794 2958 8798
rect 2985 8794 2989 8798
rect 2702 8781 2706 8787
rect 2739 8781 2743 8787
rect 2755 8783 2759 8787
rect 2870 8786 2874 8790
rect 2913 8787 2917 8791
rect 2935 8786 2942 8790
rect 2985 8787 2989 8791
rect 2856 8782 2860 8786
rect 2888 8782 2892 8786
rect 2906 8782 2910 8786
rect 2963 8782 2967 8786
rect 2978 8782 2982 8786
rect 3006 8782 3010 8786
rect 2380 8768 2384 8772
rect 2396 8768 2400 8774
rect 2430 8774 2434 8778
rect 2417 8768 2421 8772
rect 2438 8768 2442 8772
rect 2454 8768 2458 8774
rect 2475 8768 2479 8772
rect 2491 8768 2495 8772
rect 2512 8768 2516 8772
rect 2528 8768 2532 8774
rect 2562 8774 2566 8778
rect 2549 8768 2553 8772
rect 2570 8768 2574 8772
rect 2586 8768 2590 8774
rect 2607 8768 2611 8772
rect 2623 8768 2627 8772
rect 2644 8768 2648 8772
rect 2660 8768 2664 8774
rect 2694 8774 2698 8778
rect 2681 8768 2685 8772
rect 2702 8768 2706 8772
rect 2718 8768 2722 8774
rect 2739 8768 2743 8772
rect 2755 8768 2759 8772
rect 2851 8770 2855 8774
rect 2373 8757 2377 8761
rect 2410 8755 2414 8759
rect 2430 8755 2434 8759
rect 2474 8755 2478 8759
rect 2505 8757 2509 8761
rect 2542 8755 2546 8759
rect 2562 8755 2566 8759
rect 2606 8755 2610 8759
rect 2637 8757 2641 8761
rect 2674 8755 2678 8759
rect 2694 8755 2698 8759
rect 2738 8755 2742 8759
rect 2883 8768 2887 8772
rect 2903 8771 2907 8775
rect 2922 8767 2926 8771
rect 2941 8768 2945 8772
rect 2960 8768 2964 8772
rect 2973 8769 2977 8773
rect 3109 8794 3113 8798
rect 3131 8794 3135 8798
rect 3190 8794 3194 8798
rect 3215 8794 3219 8798
rect 3246 8794 3250 8798
rect 3318 8798 3322 8802
rect 3368 8798 3372 8802
rect 3421 8798 3425 8802
rect 3450 8798 3454 8802
rect 3500 8798 3504 8802
rect 3553 8798 3557 8802
rect 3582 8798 3586 8802
rect 3632 8798 3636 8802
rect 3685 8798 3689 8802
rect 3721 8801 3727 8805
rect 3801 8801 3805 8805
rect 3815 8801 3819 8805
rect 3833 8801 3837 8805
rect 3851 8801 3855 8805
rect 3874 8801 3878 8805
rect 3908 8801 3912 8805
rect 3923 8801 3927 8805
rect 3951 8801 3955 8805
rect 4076 8801 4080 8805
rect 4094 8801 4098 8805
rect 4112 8801 4116 8805
rect 4135 8801 4139 8805
rect 4169 8801 4173 8805
rect 4184 8801 4188 8805
rect 4212 8801 4216 8805
rect 3131 8786 3135 8790
rect 3174 8787 3178 8791
rect 3196 8786 3203 8790
rect 3246 8787 3250 8791
rect 3341 8787 3345 8791
rect 3149 8782 3153 8786
rect 3167 8782 3171 8786
rect 3224 8782 3228 8786
rect 3239 8782 3243 8786
rect 3267 8782 3271 8786
rect 3070 8778 3074 8782
rect 2995 8768 2999 8772
rect 3003 8769 3007 8773
rect 3015 8769 3019 8773
rect 3049 8763 3053 8767
rect 3089 8769 3093 8773
rect 3078 8762 3082 8766
rect 2856 8752 2860 8756
rect 2776 8748 2782 8752
rect 2881 8749 2885 8753
rect 2888 8752 2892 8756
rect 2906 8752 2910 8756
rect 2928 8749 2932 8753
rect 2953 8749 2957 8753
rect 2963 8752 2967 8756
rect 2979 8752 2983 8756
rect 2999 8749 3003 8753
rect 3006 8752 3010 8756
rect 3144 8768 3148 8772
rect 3164 8771 3168 8775
rect 3183 8767 3187 8771
rect 3312 8778 3316 8782
rect 3325 8781 3329 8787
rect 3362 8781 3366 8787
rect 3375 8783 3379 8787
rect 3399 8787 3403 8791
rect 3473 8787 3477 8791
rect 3383 8781 3387 8787
rect 3420 8781 3424 8787
rect 3436 8781 3440 8787
rect 3457 8781 3461 8787
rect 3494 8781 3498 8787
rect 3507 8783 3511 8787
rect 3531 8787 3535 8791
rect 3605 8787 3609 8791
rect 3515 8781 3519 8787
rect 3552 8781 3556 8787
rect 3568 8781 3572 8787
rect 3589 8781 3593 8787
rect 3626 8781 3630 8787
rect 3639 8783 3643 8787
rect 3663 8787 3667 8791
rect 3733 8794 3739 8798
rect 3815 8794 3819 8798
rect 3824 8794 3828 8798
rect 3874 8794 3878 8798
rect 3899 8794 3903 8798
rect 3930 8794 3934 8798
rect 3647 8781 3651 8787
rect 3684 8781 3688 8787
rect 3700 8783 3704 8787
rect 3815 8786 3819 8790
rect 3858 8787 3862 8791
rect 3880 8786 3887 8790
rect 3930 8787 3934 8791
rect 3801 8782 3805 8786
rect 3833 8782 3837 8786
rect 3851 8782 3855 8786
rect 3908 8782 3912 8786
rect 3923 8782 3927 8786
rect 3951 8782 3955 8786
rect 3202 8768 3206 8772
rect 3221 8768 3225 8772
rect 3234 8769 3238 8773
rect 3256 8768 3260 8772
rect 3264 8769 3268 8773
rect 3276 8769 3280 8773
rect 3325 8768 3329 8772
rect 3341 8768 3345 8774
rect 3375 8774 3379 8778
rect 3362 8768 3366 8772
rect 3383 8768 3387 8772
rect 3399 8768 3403 8774
rect 3420 8768 3424 8772
rect 3436 8768 3440 8772
rect 3457 8768 3461 8772
rect 3473 8768 3477 8774
rect 3507 8774 3511 8778
rect 3494 8768 3498 8772
rect 3515 8768 3519 8772
rect 3531 8768 3535 8774
rect 3552 8768 3556 8772
rect 3568 8768 3572 8772
rect 3589 8768 3593 8772
rect 3605 8768 3609 8774
rect 3639 8774 3643 8778
rect 3626 8768 3630 8772
rect 3647 8768 3651 8772
rect 3663 8768 3667 8774
rect 3684 8768 3688 8772
rect 3700 8768 3704 8772
rect 3796 8770 3800 8774
rect 3090 8752 3094 8756
rect 3116 8752 3120 8756
rect 2373 8741 2377 8745
rect 2424 8741 2428 8745
rect 2474 8741 2478 8745
rect 2505 8741 2509 8745
rect 2556 8741 2560 8745
rect 2606 8741 2610 8745
rect 2637 8741 2641 8745
rect 2688 8741 2692 8745
rect 2738 8741 2742 8745
rect 2812 8742 2818 8746
rect 2864 8742 2868 8746
rect 2882 8742 2886 8746
rect 2913 8742 2917 8746
rect 2935 8742 2939 8746
rect 3000 8742 3004 8746
rect 3142 8749 3146 8753
rect 3149 8752 3153 8756
rect 3167 8752 3171 8756
rect 3189 8749 3193 8753
rect 3214 8749 3218 8753
rect 3224 8752 3228 8756
rect 3240 8752 3244 8756
rect 3260 8749 3264 8753
rect 3267 8752 3271 8756
rect 3318 8757 3322 8761
rect 3355 8755 3359 8759
rect 3375 8755 3379 8759
rect 3419 8755 3423 8759
rect 3450 8757 3454 8761
rect 3487 8755 3491 8759
rect 3507 8755 3511 8759
rect 3551 8755 3555 8759
rect 3582 8757 3586 8761
rect 3619 8755 3623 8759
rect 3639 8755 3643 8759
rect 3683 8755 3687 8759
rect 3828 8768 3832 8772
rect 3848 8771 3852 8775
rect 3867 8767 3871 8771
rect 3886 8768 3890 8772
rect 3905 8768 3909 8772
rect 3918 8769 3922 8773
rect 4054 8794 4058 8798
rect 4076 8794 4080 8798
rect 4135 8794 4139 8798
rect 4160 8794 4164 8798
rect 4191 8794 4195 8798
rect 4076 8786 4080 8790
rect 4119 8787 4123 8791
rect 4141 8786 4148 8790
rect 4191 8787 4195 8791
rect 4094 8782 4098 8786
rect 4112 8782 4116 8786
rect 4169 8782 4173 8786
rect 4184 8782 4188 8786
rect 4212 8782 4216 8786
rect 4015 8778 4019 8782
rect 3940 8768 3944 8772
rect 3948 8769 3952 8773
rect 3960 8769 3964 8773
rect 3994 8763 3998 8767
rect 4034 8769 4038 8773
rect 4023 8762 4027 8766
rect 3801 8752 3805 8756
rect 3721 8748 3727 8752
rect 3826 8749 3830 8753
rect 3833 8752 3837 8756
rect 3851 8752 3855 8756
rect 3873 8749 3877 8753
rect 3898 8749 3902 8753
rect 3908 8752 3912 8756
rect 3924 8752 3928 8756
rect 3944 8749 3948 8753
rect 3951 8752 3955 8756
rect 4089 8768 4093 8772
rect 4109 8771 4113 8775
rect 4128 8767 4132 8771
rect 4147 8768 4151 8772
rect 4166 8768 4170 8772
rect 4179 8769 4183 8773
rect 4201 8768 4205 8772
rect 4209 8769 4213 8773
rect 4221 8769 4225 8773
rect 4035 8752 4039 8756
rect 4061 8752 4065 8756
rect 3060 8742 3064 8746
rect 3099 8742 3103 8746
rect 3143 8742 3147 8746
rect 3174 8742 3178 8746
rect 3196 8742 3200 8746
rect 3261 8742 3265 8746
rect 3318 8741 3322 8745
rect 3369 8741 3373 8745
rect 3419 8741 3423 8745
rect 3450 8741 3454 8745
rect 3501 8741 3505 8745
rect 3551 8741 3555 8745
rect 3582 8741 3586 8745
rect 3633 8741 3637 8745
rect 3683 8741 3687 8745
rect 3757 8742 3763 8746
rect 3809 8742 3813 8746
rect 3827 8742 3831 8746
rect 3858 8742 3862 8746
rect 3880 8742 3884 8746
rect 3945 8742 3949 8746
rect 4087 8749 4091 8753
rect 4094 8752 4098 8756
rect 4112 8752 4116 8756
rect 4134 8749 4138 8753
rect 4159 8749 4163 8753
rect 4169 8752 4173 8756
rect 4185 8752 4189 8756
rect 4205 8749 4209 8753
rect 4212 8752 4216 8756
rect 4484 8747 4488 8751
rect 4494 8747 4498 8751
rect 4504 8747 4508 8751
rect 4005 8742 4009 8746
rect 4044 8742 4048 8746
rect 4088 8742 4092 8746
rect 4119 8742 4123 8746
rect 4141 8742 4145 8746
rect 4206 8742 4210 8746
rect 4484 8742 4488 8746
rect 4494 8742 4498 8746
rect 4504 8742 4508 8746
rect 2367 8734 2371 8738
rect 2755 8734 2759 8738
rect 2764 8735 2770 8739
rect 2855 8735 2859 8739
rect 2889 8735 2893 8739
rect 2906 8735 2910 8739
rect 2962 8735 2966 8739
rect 2979 8735 2983 8739
rect 3007 8735 3011 8739
rect 3090 8735 3094 8739
rect 3116 8735 3120 8739
rect 3150 8735 3154 8739
rect 3167 8735 3171 8739
rect 3223 8735 3227 8739
rect 3240 8735 3244 8739
rect 3268 8735 3272 8739
rect 3312 8734 3316 8738
rect 3700 8734 3704 8738
rect 3709 8735 3715 8739
rect 3800 8735 3804 8739
rect 3834 8735 3838 8739
rect 3851 8735 3855 8739
rect 3907 8735 3911 8739
rect 3924 8735 3928 8739
rect 3952 8735 3956 8739
rect 4035 8735 4039 8739
rect 4061 8735 4065 8739
rect 4095 8735 4099 8739
rect 4112 8735 4116 8739
rect 4168 8735 4172 8739
rect 4185 8735 4189 8739
rect 4213 8735 4217 8739
rect 4484 8737 4488 8741
rect 4494 8737 4498 8741
rect 4504 8737 4508 8741
rect 2490 8727 2495 8731
rect 2623 8727 2627 8731
rect 2800 8728 2806 8732
rect 2864 8728 2868 8732
rect 3098 8728 3102 8732
rect 3284 8729 3288 8733
rect 3296 8729 3300 8733
rect 3435 8727 3440 8731
rect 3568 8727 3572 8731
rect 3745 8728 3751 8732
rect 3809 8728 3813 8732
rect 4043 8728 4047 8732
rect 4229 8729 4233 8733
rect 4241 8729 4245 8733
rect 4484 8732 4488 8736
rect 4494 8732 4498 8736
rect 4504 8732 4508 8736
rect 4530 8747 4534 8751
rect 4540 8747 4544 8751
rect 4550 8747 4554 8751
rect 4530 8742 4534 8746
rect 4540 8742 4544 8746
rect 4550 8742 4554 8746
rect 4530 8737 4534 8741
rect 4540 8737 4544 8741
rect 4550 8737 4554 8741
rect 4530 8732 4534 8736
rect 4540 8732 4544 8736
rect 4550 8732 4554 8736
rect 2498 8720 2502 8724
rect 2788 8720 2794 8724
rect 3108 8721 3112 8725
rect 3273 8721 3277 8725
rect 2482 8715 2486 8719
rect 2514 8715 2518 8719
rect 2836 8714 2842 8718
rect 3443 8720 3447 8724
rect 3733 8720 3739 8724
rect 4053 8721 4057 8725
rect 4218 8721 4222 8725
rect 3427 8715 3431 8719
rect 3459 8715 3463 8719
rect 3781 8714 3787 8718
rect 2482 8707 2486 8711
rect 2514 8707 2518 8711
rect 3427 8707 3431 8711
rect 3459 8707 3463 8711
rect 618 8703 622 8707
rect 628 8703 632 8707
rect 638 8703 642 8707
rect 618 8698 622 8702
rect 628 8698 632 8702
rect 638 8698 642 8702
rect 618 8693 622 8697
rect 628 8693 632 8697
rect 638 8693 642 8697
rect 618 8688 622 8692
rect 628 8688 632 8692
rect 638 8688 642 8692
rect 664 8703 668 8707
rect 674 8703 678 8707
rect 684 8703 688 8707
rect 664 8698 668 8702
rect 674 8698 678 8702
rect 684 8698 688 8702
rect 664 8693 668 8697
rect 674 8693 678 8697
rect 684 8693 688 8697
rect 2498 8700 2502 8704
rect 2755 8700 2759 8704
rect 2824 8700 2830 8704
rect 3156 8700 3160 8704
rect 3192 8700 3196 8704
rect 3259 8700 3263 8704
rect 3443 8700 3447 8704
rect 3700 8700 3704 8704
rect 3769 8700 3775 8704
rect 4101 8700 4105 8704
rect 4137 8700 4141 8704
rect 4204 8700 4208 8704
rect 2755 8692 2759 8696
rect 2764 8693 2770 8697
rect 3142 8693 3146 8697
rect 664 8688 668 8692
rect 674 8688 678 8692
rect 684 8688 688 8692
rect 2482 8688 2486 8692
rect 2514 8688 2518 8692
rect 2498 8684 2502 8688
rect 3156 8686 3160 8690
rect 3206 8686 3210 8690
rect 3259 8686 3263 8690
rect 3700 8692 3704 8696
rect 3709 8693 3715 8697
rect 4087 8693 4091 8697
rect 3427 8688 3431 8692
rect 3459 8688 3463 8692
rect 3443 8684 3447 8688
rect 4101 8686 4105 8690
rect 4151 8686 4155 8690
rect 4204 8686 4208 8690
rect 2490 8677 2495 8681
rect 2624 8677 2628 8681
rect 3179 8675 3183 8679
rect 2373 8670 2377 8674
rect 2409 8670 2413 8674
rect 2476 8670 2480 8674
rect 2505 8670 2509 8674
rect 2541 8670 2545 8674
rect 2608 8670 2612 8674
rect 2637 8670 2641 8674
rect 2673 8670 2677 8674
rect 2740 8670 2744 8674
rect 2824 8670 2830 8674
rect 2764 8663 2770 8667
rect 3150 8666 3154 8670
rect 3163 8669 3167 8675
rect 3200 8669 3204 8675
rect 3213 8671 3217 8675
rect 3237 8675 3241 8679
rect 3435 8677 3440 8681
rect 3569 8677 3573 8681
rect 4124 8675 4128 8679
rect 3221 8669 3225 8675
rect 3258 8669 3262 8675
rect 3274 8669 3278 8675
rect 3318 8670 3322 8674
rect 3354 8670 3358 8674
rect 3421 8670 3425 8674
rect 3450 8670 3454 8674
rect 3486 8670 3490 8674
rect 3553 8670 3557 8674
rect 3582 8670 3586 8674
rect 3618 8670 3622 8674
rect 3685 8670 3689 8674
rect 3769 8670 3775 8674
rect 2373 8656 2377 8660
rect 2423 8656 2427 8660
rect 2476 8656 2480 8660
rect 2505 8656 2509 8660
rect 2555 8656 2559 8660
rect 2608 8656 2612 8660
rect 2637 8656 2641 8660
rect 2687 8656 2691 8660
rect 2740 8656 2744 8660
rect 3163 8656 3167 8660
rect 3179 8656 3183 8662
rect 3213 8662 3217 8666
rect 3200 8656 3204 8660
rect 2396 8645 2400 8649
rect 2367 8636 2371 8640
rect 2380 8639 2384 8645
rect 2417 8639 2421 8645
rect 2430 8641 2434 8645
rect 2454 8645 2458 8649
rect 2528 8645 2532 8649
rect 2438 8639 2442 8645
rect 2475 8639 2479 8645
rect 2491 8639 2495 8645
rect 2512 8639 2516 8645
rect 2549 8639 2553 8645
rect 2562 8641 2566 8645
rect 2586 8645 2590 8649
rect 2660 8645 2664 8649
rect 2570 8639 2574 8645
rect 2607 8639 2611 8645
rect 2623 8639 2627 8645
rect 2644 8639 2648 8645
rect 2681 8639 2685 8645
rect 2694 8641 2698 8645
rect 2718 8645 2722 8649
rect 2702 8639 2706 8645
rect 2739 8639 2743 8645
rect 2755 8641 2759 8645
rect 3221 8656 3225 8660
rect 3237 8656 3241 8662
rect 3709 8663 3715 8667
rect 4095 8666 4099 8670
rect 4108 8669 4112 8675
rect 4145 8669 4149 8675
rect 4158 8671 4162 8675
rect 4182 8675 4186 8679
rect 4166 8669 4170 8675
rect 4203 8669 4207 8675
rect 4219 8669 4223 8675
rect 3258 8656 3262 8660
rect 3274 8656 3278 8660
rect 3318 8656 3322 8660
rect 3368 8656 3372 8660
rect 3421 8656 3425 8660
rect 3450 8656 3454 8660
rect 3500 8656 3504 8660
rect 3553 8656 3557 8660
rect 3582 8656 3586 8660
rect 3632 8656 3636 8660
rect 3685 8656 3689 8660
rect 4108 8656 4112 8660
rect 4124 8656 4128 8662
rect 4158 8662 4162 8666
rect 4145 8656 4149 8660
rect 3156 8645 3160 8649
rect 3193 8643 3197 8647
rect 3213 8643 3217 8647
rect 3257 8643 3261 8647
rect 3341 8645 3345 8649
rect 2380 8626 2384 8630
rect 2396 8626 2400 8632
rect 2430 8632 2434 8636
rect 2417 8626 2421 8630
rect 2438 8626 2442 8630
rect 2454 8626 2458 8632
rect 2475 8626 2479 8630
rect 2491 8626 2495 8630
rect 2512 8626 2516 8630
rect 2528 8626 2532 8632
rect 2562 8632 2566 8636
rect 2549 8626 2553 8630
rect 2570 8626 2574 8630
rect 2586 8626 2590 8632
rect 2607 8626 2611 8630
rect 2623 8626 2627 8630
rect 2644 8626 2648 8630
rect 2660 8626 2664 8632
rect 2694 8632 2698 8636
rect 2681 8626 2685 8630
rect 2702 8626 2706 8630
rect 2718 8626 2722 8632
rect 2776 8636 2782 8640
rect 3312 8636 3316 8640
rect 3325 8639 3329 8645
rect 3362 8639 3366 8645
rect 3375 8641 3379 8645
rect 3399 8645 3403 8649
rect 3473 8645 3477 8649
rect 3383 8639 3387 8645
rect 3420 8639 3424 8645
rect 3436 8639 3440 8645
rect 3457 8639 3461 8645
rect 3494 8639 3498 8645
rect 3507 8641 3511 8645
rect 3531 8645 3535 8649
rect 3605 8645 3609 8649
rect 3515 8639 3519 8645
rect 3552 8639 3556 8645
rect 3568 8639 3572 8645
rect 3589 8639 3593 8645
rect 3626 8639 3630 8645
rect 3639 8641 3643 8645
rect 3663 8645 3667 8649
rect 3647 8639 3651 8645
rect 3684 8639 3688 8645
rect 3700 8641 3704 8645
rect 4166 8656 4170 8660
rect 4182 8656 4186 8662
rect 4203 8656 4207 8660
rect 4219 8656 4223 8660
rect 4101 8645 4105 8649
rect 4138 8643 4142 8647
rect 4158 8643 4162 8647
rect 4202 8643 4206 8647
rect 2739 8626 2743 8630
rect 2755 8626 2759 8630
rect 2812 8629 2818 8633
rect 3156 8629 3160 8633
rect 3207 8629 3211 8633
rect 3257 8629 3261 8633
rect 3325 8626 3329 8630
rect 3341 8626 3345 8632
rect 3375 8632 3379 8636
rect 3362 8626 3366 8630
rect 2373 8615 2377 8619
rect 2410 8613 2414 8617
rect 2430 8613 2434 8617
rect 2474 8613 2478 8617
rect 2505 8615 2509 8619
rect 2542 8613 2546 8617
rect 2562 8613 2566 8617
rect 2606 8613 2610 8617
rect 2637 8615 2641 8619
rect 2674 8613 2678 8617
rect 2694 8613 2698 8617
rect 2738 8613 2742 8617
rect 3149 8621 3153 8625
rect 3274 8622 3278 8626
rect 3383 8626 3387 8630
rect 3399 8626 3403 8632
rect 3420 8626 3424 8630
rect 3436 8626 3440 8630
rect 3457 8626 3461 8630
rect 3473 8626 3477 8632
rect 3507 8632 3511 8636
rect 3494 8626 3498 8630
rect 3515 8626 3519 8630
rect 3531 8626 3535 8632
rect 3552 8626 3556 8630
rect 3568 8626 3572 8630
rect 3589 8626 3593 8630
rect 3605 8626 3609 8632
rect 3639 8632 3643 8636
rect 3626 8626 3630 8630
rect 3647 8626 3651 8630
rect 3663 8626 3667 8632
rect 3721 8636 3727 8640
rect 3684 8626 3688 8630
rect 3700 8626 3704 8630
rect 3757 8629 3763 8633
rect 4101 8629 4105 8633
rect 4152 8629 4156 8633
rect 4202 8629 4206 8633
rect 2824 8614 2830 8618
rect 3156 8614 3160 8618
rect 3192 8614 3196 8618
rect 3259 8614 3263 8618
rect 2776 8606 2782 8610
rect 3142 8607 3146 8611
rect 3318 8615 3322 8619
rect 3355 8613 3359 8617
rect 3375 8613 3379 8617
rect 3419 8613 3423 8617
rect 3450 8615 3454 8619
rect 3487 8613 3491 8617
rect 3507 8613 3511 8617
rect 3551 8613 3555 8617
rect 3582 8615 3586 8619
rect 3619 8613 3623 8617
rect 3639 8613 3643 8617
rect 3683 8613 3687 8617
rect 4094 8621 4098 8625
rect 4219 8622 4223 8626
rect 3769 8614 3775 8618
rect 4101 8614 4105 8618
rect 4137 8614 4141 8618
rect 4204 8614 4208 8618
rect 2373 8599 2377 8603
rect 2424 8599 2428 8603
rect 2474 8599 2478 8603
rect 2505 8599 2509 8603
rect 2556 8599 2560 8603
rect 2606 8599 2610 8603
rect 2637 8599 2641 8603
rect 2688 8599 2692 8603
rect 2738 8599 2742 8603
rect 2812 8599 2818 8603
rect 3156 8600 3160 8604
rect 3206 8600 3210 8604
rect 3259 8600 3263 8604
rect 3721 8606 3727 8610
rect 4087 8607 4091 8611
rect 3318 8599 3322 8603
rect 3369 8599 3373 8603
rect 3419 8599 3423 8603
rect 3450 8599 3454 8603
rect 3501 8599 3505 8603
rect 3551 8599 3555 8603
rect 3582 8599 3586 8603
rect 3633 8599 3637 8603
rect 3683 8599 3687 8603
rect 3757 8599 3763 8603
rect 4101 8600 4105 8604
rect 4151 8600 4155 8604
rect 4204 8600 4208 8604
rect 2366 8592 2370 8596
rect 2755 8592 2759 8596
rect 3179 8589 3183 8593
rect 2373 8584 2377 8588
rect 2409 8584 2413 8588
rect 2476 8584 2480 8588
rect 2505 8584 2509 8588
rect 2541 8584 2545 8588
rect 2608 8584 2612 8588
rect 2637 8584 2641 8588
rect 2673 8584 2677 8588
rect 2740 8584 2744 8588
rect 2824 8584 2830 8588
rect 2764 8577 2770 8581
rect 3150 8580 3154 8584
rect 3163 8583 3167 8589
rect 3200 8583 3204 8589
rect 3213 8585 3217 8589
rect 3237 8589 3241 8593
rect 3311 8592 3315 8596
rect 3700 8592 3704 8596
rect 4124 8589 4128 8593
rect 3221 8583 3225 8589
rect 3258 8583 3262 8589
rect 3274 8585 3278 8589
rect 3296 8583 3300 8587
rect 3318 8584 3322 8588
rect 3354 8584 3358 8588
rect 3421 8584 3425 8588
rect 3450 8584 3454 8588
rect 3486 8584 3490 8588
rect 3553 8584 3557 8588
rect 3582 8584 3586 8588
rect 3618 8584 3622 8588
rect 3685 8584 3689 8588
rect 3769 8584 3775 8588
rect 2373 8570 2377 8574
rect 2423 8570 2427 8574
rect 2476 8570 2480 8574
rect 2505 8570 2509 8574
rect 2555 8570 2559 8574
rect 2608 8570 2612 8574
rect 2637 8570 2641 8574
rect 2687 8570 2691 8574
rect 2740 8570 2744 8574
rect 3163 8570 3167 8574
rect 3179 8570 3183 8576
rect 3213 8576 3217 8580
rect 3200 8570 3204 8574
rect 2396 8559 2400 8563
rect 2367 8550 2371 8554
rect 2380 8553 2384 8559
rect 2417 8553 2421 8559
rect 2430 8555 2434 8559
rect 2454 8559 2458 8563
rect 2528 8559 2532 8563
rect 2438 8553 2442 8559
rect 2475 8553 2479 8559
rect 2491 8553 2495 8559
rect 2512 8553 2516 8559
rect 2549 8553 2553 8559
rect 2562 8555 2566 8559
rect 2586 8559 2590 8563
rect 2660 8559 2664 8563
rect 2570 8553 2574 8559
rect 2607 8553 2611 8559
rect 2623 8553 2627 8559
rect 2644 8553 2648 8559
rect 2681 8553 2685 8559
rect 2694 8555 2698 8559
rect 2718 8559 2722 8563
rect 2702 8553 2706 8559
rect 2739 8553 2743 8559
rect 2755 8555 2759 8559
rect 3221 8570 3225 8574
rect 3237 8570 3241 8576
rect 3258 8570 3262 8574
rect 3274 8570 3278 8579
rect 3709 8577 3715 8581
rect 4095 8580 4099 8584
rect 4108 8583 4112 8589
rect 4145 8583 4149 8589
rect 4158 8585 4162 8589
rect 4182 8589 4186 8593
rect 4166 8583 4170 8589
rect 4203 8583 4207 8589
rect 4219 8585 4223 8589
rect 4241 8583 4245 8587
rect 3296 8567 3300 8571
rect 3318 8570 3322 8574
rect 3368 8570 3372 8574
rect 3421 8570 3425 8574
rect 3450 8570 3454 8574
rect 3500 8570 3504 8574
rect 3553 8570 3557 8574
rect 3582 8570 3586 8574
rect 3632 8570 3636 8574
rect 3685 8570 3689 8574
rect 4108 8570 4112 8574
rect 4124 8570 4128 8576
rect 4158 8576 4162 8580
rect 4145 8570 4149 8574
rect 3156 8559 3160 8563
rect 3193 8557 3197 8561
rect 3213 8557 3217 8561
rect 3257 8557 3261 8561
rect 3341 8559 3345 8563
rect 2380 8540 2384 8544
rect 2396 8540 2400 8546
rect 2430 8546 2434 8550
rect 2417 8540 2421 8544
rect 2438 8540 2442 8544
rect 2454 8540 2458 8546
rect 2475 8540 2479 8544
rect 2491 8540 2495 8544
rect 2512 8540 2516 8544
rect 2528 8540 2532 8546
rect 2562 8546 2566 8550
rect 2549 8540 2553 8544
rect 2570 8540 2574 8544
rect 2586 8540 2590 8546
rect 2607 8540 2611 8544
rect 2623 8540 2627 8544
rect 2644 8540 2648 8544
rect 2660 8540 2664 8546
rect 2694 8546 2698 8550
rect 2681 8540 2685 8544
rect 2702 8540 2706 8544
rect 2718 8540 2722 8546
rect 2776 8550 2782 8554
rect 3312 8550 3316 8554
rect 3325 8553 3329 8559
rect 3362 8553 3366 8559
rect 3375 8555 3379 8559
rect 3399 8559 3403 8563
rect 3473 8559 3477 8563
rect 3383 8553 3387 8559
rect 3420 8553 3424 8559
rect 3436 8553 3440 8559
rect 3457 8553 3461 8559
rect 3494 8553 3498 8559
rect 3507 8555 3511 8559
rect 3531 8559 3535 8563
rect 3605 8559 3609 8563
rect 3515 8553 3519 8559
rect 3552 8553 3556 8559
rect 3568 8553 3572 8559
rect 3589 8553 3593 8559
rect 3626 8553 3630 8559
rect 3639 8555 3643 8559
rect 3663 8559 3667 8563
rect 3647 8553 3651 8559
rect 3684 8553 3688 8559
rect 3700 8555 3704 8559
rect 4166 8570 4170 8574
rect 4182 8570 4186 8576
rect 4203 8570 4207 8574
rect 4219 8570 4223 8579
rect 4241 8567 4245 8571
rect 4101 8559 4105 8563
rect 4138 8557 4142 8561
rect 4158 8557 4162 8561
rect 4202 8557 4206 8561
rect 2739 8540 2743 8544
rect 2755 8540 2759 8544
rect 2812 8543 2818 8547
rect 3156 8543 3160 8547
rect 3207 8543 3211 8547
rect 3257 8543 3261 8547
rect 3325 8540 3329 8544
rect 3341 8540 3345 8546
rect 3375 8546 3379 8550
rect 3362 8540 3366 8544
rect 3383 8540 3387 8544
rect 3399 8540 3403 8546
rect 3420 8540 3424 8544
rect 3436 8540 3440 8544
rect 3457 8540 3461 8544
rect 3473 8540 3477 8546
rect 3507 8546 3511 8550
rect 3494 8540 3498 8544
rect 3515 8540 3519 8544
rect 3531 8540 3535 8546
rect 3552 8540 3556 8544
rect 3568 8540 3572 8544
rect 3589 8540 3593 8544
rect 3605 8540 3609 8546
rect 3639 8546 3643 8550
rect 3626 8540 3630 8544
rect 3647 8540 3651 8544
rect 3663 8540 3667 8546
rect 3721 8550 3727 8554
rect 3684 8540 3688 8544
rect 3700 8540 3704 8544
rect 3757 8543 3763 8547
rect 4101 8543 4105 8547
rect 4152 8543 4156 8547
rect 4202 8543 4206 8547
rect 2373 8529 2377 8533
rect 2410 8527 2414 8531
rect 2430 8527 2434 8531
rect 2474 8527 2478 8531
rect 2505 8529 2509 8533
rect 2542 8527 2546 8531
rect 2562 8527 2566 8531
rect 2606 8527 2610 8531
rect 2637 8529 2641 8533
rect 2674 8527 2678 8531
rect 2694 8527 2698 8531
rect 2738 8527 2742 8531
rect 3318 8529 3322 8533
rect 3355 8527 3359 8531
rect 3375 8527 3379 8531
rect 3419 8527 3423 8531
rect 3450 8529 3454 8533
rect 3487 8527 3491 8531
rect 3507 8527 3511 8531
rect 3551 8527 3555 8531
rect 3582 8529 3586 8533
rect 3619 8527 3623 8531
rect 3639 8527 3643 8531
rect 3683 8527 3687 8531
rect 2776 8520 2782 8524
rect 3721 8520 3727 8524
rect 2373 8513 2377 8517
rect 2424 8513 2428 8517
rect 2474 8513 2478 8517
rect 2505 8513 2509 8517
rect 2556 8513 2560 8517
rect 2606 8513 2610 8517
rect 2637 8513 2641 8517
rect 2688 8513 2692 8517
rect 2738 8513 2742 8517
rect 2812 8513 2818 8517
rect 3318 8513 3322 8517
rect 3369 8513 3373 8517
rect 3419 8513 3423 8517
rect 3450 8513 3454 8517
rect 3501 8513 3505 8517
rect 3551 8513 3555 8517
rect 3582 8513 3586 8517
rect 3633 8513 3637 8517
rect 3683 8513 3687 8517
rect 3757 8513 3763 8517
rect 2366 8506 2370 8510
rect 2755 8506 2759 8510
rect 3311 8506 3315 8510
rect 3700 8506 3704 8510
rect 2491 8499 2495 8503
rect 2599 8499 2603 8503
rect 2623 8499 2627 8503
rect 3436 8499 3440 8503
rect 3544 8499 3548 8503
rect 3568 8499 3572 8503
rect 2615 8492 2619 8496
rect 2599 8488 2603 8492
rect 2631 8488 2635 8492
rect 3560 8492 3564 8496
rect 3544 8488 3548 8492
rect 3576 8488 3580 8492
rect 2599 8481 2603 8485
rect 2631 8481 2635 8485
rect 3296 8481 3300 8485
rect 3544 8481 3548 8485
rect 3576 8481 3580 8485
rect 4241 8481 4245 8485
rect 2615 8474 2619 8478
rect 2755 8474 2759 8478
rect 3560 8474 3564 8478
rect 3700 8474 3704 8478
rect 2755 8466 2759 8470
rect 3700 8466 3704 8470
rect 2599 8462 2603 8466
rect 2631 8462 2635 8466
rect 2615 8458 2619 8462
rect 3544 8462 3548 8466
rect 3576 8462 3580 8466
rect 3560 8458 3564 8462
rect 2491 8451 2495 8455
rect 2599 8451 2603 8455
rect 2623 8451 2627 8455
rect 3436 8451 3440 8455
rect 3544 8451 3548 8455
rect 3568 8451 3572 8455
rect 2373 8444 2377 8448
rect 2409 8444 2413 8448
rect 2476 8444 2480 8448
rect 2505 8444 2509 8448
rect 2541 8444 2545 8448
rect 2608 8444 2612 8448
rect 2637 8444 2641 8448
rect 2673 8444 2677 8448
rect 2740 8444 2744 8448
rect 2824 8444 2830 8448
rect 3318 8444 3322 8448
rect 3354 8444 3358 8448
rect 3421 8444 3425 8448
rect 3450 8444 3454 8448
rect 3486 8444 3490 8448
rect 3553 8444 3557 8448
rect 3582 8444 3586 8448
rect 3618 8444 3622 8448
rect 3685 8444 3689 8448
rect 3769 8444 3775 8448
rect 2764 8437 2770 8441
rect 3709 8437 3715 8441
rect 4484 8438 4488 8442
rect 4494 8438 4498 8442
rect 4504 8438 4508 8442
rect 2373 8430 2377 8434
rect 2423 8430 2427 8434
rect 2476 8430 2480 8434
rect 2505 8430 2509 8434
rect 2555 8430 2559 8434
rect 2608 8430 2612 8434
rect 2637 8430 2641 8434
rect 2687 8430 2691 8434
rect 2740 8430 2744 8434
rect 3318 8430 3322 8434
rect 3368 8430 3372 8434
rect 3421 8430 3425 8434
rect 3450 8430 3454 8434
rect 3500 8430 3504 8434
rect 3553 8430 3557 8434
rect 3582 8430 3586 8434
rect 3632 8430 3636 8434
rect 3685 8430 3689 8434
rect 4484 8433 4488 8437
rect 4494 8433 4498 8437
rect 4504 8433 4508 8437
rect 4484 8428 4488 8432
rect 4494 8428 4498 8432
rect 4504 8428 4508 8432
rect 2396 8419 2400 8423
rect 2367 8410 2371 8414
rect 2380 8413 2384 8419
rect 2417 8413 2421 8419
rect 2430 8415 2434 8419
rect 2454 8419 2458 8423
rect 2528 8419 2532 8423
rect 2438 8413 2442 8419
rect 2475 8413 2479 8419
rect 2491 8413 2495 8419
rect 2512 8413 2516 8419
rect 2549 8413 2553 8419
rect 2562 8415 2566 8419
rect 2586 8419 2590 8423
rect 2660 8419 2664 8423
rect 2570 8413 2574 8419
rect 2607 8413 2611 8419
rect 2623 8413 2627 8419
rect 2644 8413 2648 8419
rect 2681 8413 2685 8419
rect 2694 8415 2698 8419
rect 2718 8419 2722 8423
rect 3341 8419 3345 8423
rect 2702 8413 2706 8419
rect 2739 8413 2743 8419
rect 2755 8415 2759 8419
rect 2380 8400 2384 8404
rect 2396 8400 2400 8406
rect 2430 8406 2434 8410
rect 2417 8400 2421 8404
rect 618 8394 622 8398
rect 628 8394 632 8398
rect 638 8394 642 8398
rect 618 8389 622 8393
rect 628 8389 632 8393
rect 638 8389 642 8393
rect 618 8384 622 8388
rect 628 8384 632 8388
rect 638 8384 642 8388
rect 618 8379 622 8383
rect 628 8379 632 8383
rect 638 8379 642 8383
rect 664 8394 668 8398
rect 674 8394 678 8398
rect 684 8394 688 8398
rect 664 8389 668 8393
rect 674 8389 678 8393
rect 684 8389 688 8393
rect 664 8384 668 8388
rect 674 8384 678 8388
rect 684 8384 688 8388
rect 2438 8400 2442 8404
rect 2454 8400 2458 8406
rect 2475 8400 2479 8404
rect 2491 8400 2495 8404
rect 2512 8400 2516 8404
rect 2528 8400 2532 8406
rect 2562 8406 2566 8410
rect 2549 8400 2553 8404
rect 2570 8400 2574 8404
rect 2586 8400 2590 8406
rect 2607 8400 2611 8404
rect 2623 8400 2627 8404
rect 2644 8400 2648 8404
rect 2660 8400 2664 8406
rect 2694 8406 2698 8410
rect 2681 8400 2685 8404
rect 2702 8400 2706 8404
rect 2718 8400 2722 8406
rect 3312 8410 3316 8414
rect 3325 8413 3329 8419
rect 3362 8413 3366 8419
rect 3375 8415 3379 8419
rect 3399 8419 3403 8423
rect 3473 8419 3477 8423
rect 3383 8413 3387 8419
rect 3420 8413 3424 8419
rect 3436 8413 3440 8419
rect 3457 8413 3461 8419
rect 3494 8413 3498 8419
rect 3507 8415 3511 8419
rect 3531 8419 3535 8423
rect 3605 8419 3609 8423
rect 3515 8413 3519 8419
rect 3552 8413 3556 8419
rect 3568 8413 3572 8419
rect 3589 8413 3593 8419
rect 3626 8413 3630 8419
rect 3639 8415 3643 8419
rect 3663 8419 3667 8423
rect 4484 8423 4488 8427
rect 4494 8423 4498 8427
rect 4504 8423 4508 8427
rect 4530 8438 4534 8442
rect 4540 8438 4544 8442
rect 4550 8438 4554 8442
rect 4530 8433 4534 8437
rect 4540 8433 4544 8437
rect 4550 8433 4554 8437
rect 4530 8428 4534 8432
rect 4540 8428 4544 8432
rect 4550 8428 4554 8432
rect 4530 8423 4534 8427
rect 4540 8423 4544 8427
rect 4550 8423 4554 8427
rect 3647 8413 3651 8419
rect 3684 8413 3688 8419
rect 3700 8415 3704 8419
rect 2739 8400 2743 8404
rect 2755 8400 2759 8404
rect 3325 8400 3329 8404
rect 3341 8400 3345 8406
rect 3375 8406 3379 8410
rect 3362 8400 3366 8404
rect 3383 8400 3387 8404
rect 3399 8400 3403 8406
rect 3420 8400 3424 8404
rect 3436 8400 3440 8404
rect 3457 8400 3461 8404
rect 3473 8400 3477 8406
rect 3507 8406 3511 8410
rect 3494 8400 3498 8404
rect 3515 8400 3519 8404
rect 3531 8400 3535 8406
rect 3552 8400 3556 8404
rect 3568 8400 3572 8404
rect 3589 8400 3593 8404
rect 3605 8400 3609 8406
rect 3639 8406 3643 8410
rect 3626 8400 3630 8404
rect 3647 8400 3651 8404
rect 3663 8400 3667 8406
rect 3684 8400 3688 8404
rect 3700 8400 3704 8404
rect 2373 8389 2377 8393
rect 2410 8387 2414 8391
rect 2430 8387 2434 8391
rect 2474 8387 2478 8391
rect 2505 8389 2509 8393
rect 2542 8387 2546 8391
rect 2562 8387 2566 8391
rect 2606 8387 2610 8391
rect 2637 8389 2641 8393
rect 2674 8387 2678 8391
rect 2694 8387 2698 8391
rect 2738 8387 2742 8391
rect 3318 8389 3322 8393
rect 3355 8387 3359 8391
rect 3375 8387 3379 8391
rect 3419 8387 3423 8391
rect 3450 8389 3454 8393
rect 3487 8387 3491 8391
rect 3507 8387 3511 8391
rect 3551 8387 3555 8391
rect 3582 8389 3586 8393
rect 3619 8387 3623 8391
rect 3639 8387 3643 8391
rect 3683 8387 3687 8391
rect 664 8379 668 8383
rect 674 8379 678 8383
rect 684 8379 688 8383
rect 2776 8380 2782 8384
rect 3721 8380 3727 8384
rect 2373 8373 2377 8377
rect 2424 8373 2428 8377
rect 2474 8373 2478 8377
rect 2505 8373 2509 8377
rect 2556 8373 2560 8377
rect 2606 8373 2610 8377
rect 2637 8373 2641 8377
rect 2688 8373 2692 8377
rect 2738 8373 2742 8377
rect 2812 8373 2818 8377
rect 3318 8373 3322 8377
rect 3369 8373 3373 8377
rect 3419 8373 3423 8377
rect 3450 8373 3454 8377
rect 3501 8373 3505 8377
rect 3551 8373 3555 8377
rect 3582 8373 3586 8377
rect 3633 8373 3637 8377
rect 3683 8373 3687 8377
rect 3757 8373 3763 8377
rect 2824 8365 2830 8369
rect 2857 8365 2861 8369
rect 2893 8365 2897 8369
rect 2960 8365 2964 8369
rect 2989 8365 2993 8369
rect 3025 8365 3029 8369
rect 3092 8365 3096 8369
rect 3121 8365 3125 8369
rect 3157 8365 3161 8369
rect 3224 8365 3228 8369
rect 3253 8365 3257 8369
rect 3289 8365 3293 8369
rect 3356 8365 3360 8369
rect 3769 8365 3775 8369
rect 3802 8365 3806 8369
rect 3838 8365 3842 8369
rect 3905 8365 3909 8369
rect 3934 8365 3938 8369
rect 3970 8365 3974 8369
rect 4037 8365 4041 8369
rect 4066 8365 4070 8369
rect 4102 8365 4106 8369
rect 4169 8365 4173 8369
rect 4198 8365 4202 8369
rect 4234 8365 4238 8369
rect 4301 8365 4305 8369
rect 2764 8358 2770 8362
rect 3709 8358 3715 8362
rect 2857 8351 2861 8355
rect 2907 8351 2911 8355
rect 2960 8351 2964 8355
rect 2989 8351 2993 8355
rect 3039 8351 3043 8355
rect 3092 8351 3096 8355
rect 3121 8351 3125 8355
rect 3171 8351 3175 8355
rect 3224 8351 3228 8355
rect 3253 8351 3257 8355
rect 3303 8351 3307 8355
rect 3356 8351 3360 8355
rect 3802 8351 3806 8355
rect 3852 8351 3856 8355
rect 3905 8351 3909 8355
rect 3934 8351 3938 8355
rect 3984 8351 3988 8355
rect 4037 8351 4041 8355
rect 4066 8351 4070 8355
rect 4116 8351 4120 8355
rect 4169 8351 4173 8355
rect 4198 8351 4202 8355
rect 4248 8351 4252 8355
rect 4301 8351 4305 8355
rect 2880 8340 2884 8344
rect 2505 8332 2509 8336
rect 2541 8332 2545 8336
rect 2608 8332 2612 8336
rect 2824 8332 2830 8336
rect 2851 8331 2855 8335
rect 2864 8334 2868 8340
rect 2901 8334 2905 8340
rect 2914 8336 2918 8340
rect 2938 8340 2942 8344
rect 3012 8340 3016 8344
rect 2922 8334 2926 8340
rect 2959 8334 2963 8340
rect 2975 8336 2979 8340
rect 2764 8325 2770 8329
rect 2505 8318 2509 8322
rect 2555 8318 2559 8322
rect 2608 8318 2612 8322
rect 2864 8321 2868 8325
rect 2880 8321 2884 8327
rect 2914 8327 2918 8331
rect 2901 8321 2905 8325
rect 2922 8321 2926 8325
rect 2938 8321 2942 8327
rect 2983 8331 2987 8335
rect 2996 8334 3000 8340
rect 3033 8334 3037 8340
rect 3046 8336 3050 8340
rect 3070 8340 3074 8344
rect 3144 8340 3148 8344
rect 3054 8334 3058 8340
rect 3091 8334 3095 8340
rect 3107 8336 3111 8340
rect 2959 8321 2963 8325
rect 2975 8321 2979 8325
rect 2996 8321 3000 8325
rect 3012 8321 3016 8327
rect 3046 8327 3050 8331
rect 3033 8321 3037 8325
rect 3054 8321 3058 8325
rect 3070 8321 3074 8327
rect 3115 8331 3119 8335
rect 3128 8334 3132 8340
rect 3165 8334 3169 8340
rect 3178 8336 3182 8340
rect 3202 8340 3206 8344
rect 3276 8340 3280 8344
rect 3186 8334 3190 8340
rect 3223 8334 3227 8340
rect 3239 8336 3243 8340
rect 3091 8321 3095 8325
rect 3107 8321 3111 8325
rect 3128 8321 3132 8325
rect 3144 8321 3148 8327
rect 3178 8327 3182 8331
rect 3165 8321 3169 8325
rect 3186 8321 3190 8325
rect 3202 8321 3206 8327
rect 3247 8331 3251 8335
rect 3260 8334 3264 8340
rect 3297 8334 3301 8340
rect 3310 8336 3314 8340
rect 3334 8340 3338 8344
rect 3825 8340 3829 8344
rect 3318 8334 3322 8340
rect 3355 8334 3359 8340
rect 3371 8336 3375 8340
rect 3450 8332 3454 8336
rect 3486 8332 3490 8336
rect 3553 8332 3557 8336
rect 3769 8332 3775 8336
rect 3223 8321 3227 8325
rect 3239 8321 3243 8325
rect 3260 8321 3264 8325
rect 3276 8321 3280 8327
rect 3310 8327 3314 8331
rect 3297 8321 3301 8325
rect 2528 8307 2532 8311
rect 2490 8298 2494 8302
rect 2512 8301 2516 8307
rect 2549 8301 2553 8307
rect 2562 8303 2566 8307
rect 2586 8307 2590 8311
rect 2570 8301 2574 8307
rect 2607 8301 2611 8307
rect 2623 8301 2627 8307
rect 2857 8310 2861 8314
rect 2894 8308 2898 8312
rect 2914 8308 2918 8312
rect 2958 8308 2962 8312
rect 2989 8310 2993 8314
rect 3026 8308 3030 8312
rect 3046 8308 3050 8312
rect 3090 8308 3094 8312
rect 3121 8310 3125 8314
rect 3158 8308 3162 8312
rect 3178 8308 3182 8312
rect 3222 8308 3226 8312
rect 3239 8313 3243 8317
rect 3318 8321 3322 8325
rect 3334 8321 3338 8327
rect 3796 8331 3800 8335
rect 3809 8334 3813 8340
rect 3846 8334 3850 8340
rect 3859 8336 3863 8340
rect 3883 8340 3887 8344
rect 3957 8340 3961 8344
rect 3867 8334 3871 8340
rect 3904 8334 3908 8340
rect 3920 8336 3924 8340
rect 3709 8325 3715 8329
rect 3355 8321 3359 8325
rect 3371 8321 3375 8325
rect 3253 8310 3257 8314
rect 3290 8308 3294 8312
rect 3310 8308 3314 8312
rect 3354 8308 3358 8312
rect 3371 8313 3375 8317
rect 3450 8318 3454 8322
rect 3500 8318 3504 8322
rect 3553 8318 3557 8322
rect 3809 8321 3813 8325
rect 3825 8321 3829 8327
rect 3859 8327 3863 8331
rect 3846 8321 3850 8325
rect 3867 8321 3871 8325
rect 3883 8321 3887 8327
rect 3928 8331 3932 8335
rect 3941 8334 3945 8340
rect 3978 8334 3982 8340
rect 3991 8336 3995 8340
rect 4015 8340 4019 8344
rect 4089 8340 4093 8344
rect 3999 8334 4003 8340
rect 4036 8334 4040 8340
rect 4052 8336 4056 8340
rect 3904 8321 3908 8325
rect 3920 8321 3924 8325
rect 3941 8321 3945 8325
rect 3957 8321 3961 8327
rect 3991 8327 3995 8331
rect 3978 8321 3982 8325
rect 3999 8321 4003 8325
rect 4015 8321 4019 8327
rect 4060 8331 4064 8335
rect 4073 8334 4077 8340
rect 4110 8334 4114 8340
rect 4123 8336 4127 8340
rect 4147 8340 4151 8344
rect 4221 8340 4225 8344
rect 4131 8334 4135 8340
rect 4168 8334 4172 8340
rect 4184 8336 4188 8340
rect 4036 8321 4040 8325
rect 4052 8321 4056 8325
rect 4073 8321 4077 8325
rect 4089 8321 4093 8327
rect 4123 8327 4127 8331
rect 4110 8321 4114 8325
rect 4131 8321 4135 8325
rect 4147 8321 4151 8327
rect 4192 8331 4196 8335
rect 4205 8334 4209 8340
rect 4242 8334 4246 8340
rect 4255 8336 4259 8340
rect 4279 8340 4283 8344
rect 4263 8334 4267 8340
rect 4300 8334 4304 8340
rect 4316 8336 4320 8340
rect 4168 8321 4172 8325
rect 4184 8321 4188 8325
rect 4205 8321 4209 8325
rect 4221 8321 4225 8327
rect 4255 8327 4259 8331
rect 4242 8321 4246 8325
rect 3473 8307 3477 8311
rect 2776 8301 2782 8305
rect 2512 8288 2516 8292
rect 2528 8288 2532 8294
rect 2562 8294 2566 8298
rect 2549 8288 2553 8292
rect 2570 8288 2574 8292
rect 2586 8288 2590 8294
rect 3435 8298 3439 8302
rect 3457 8301 3461 8307
rect 3494 8301 3498 8307
rect 3507 8303 3511 8307
rect 3531 8307 3535 8311
rect 3515 8301 3519 8307
rect 3552 8301 3556 8307
rect 3568 8301 3572 8307
rect 3802 8310 3806 8314
rect 3839 8308 3843 8312
rect 3859 8308 3863 8312
rect 3903 8308 3907 8312
rect 3934 8310 3938 8314
rect 3971 8308 3975 8312
rect 3991 8308 3995 8312
rect 4035 8308 4039 8312
rect 4066 8310 4070 8314
rect 4103 8308 4107 8312
rect 4123 8308 4127 8312
rect 4167 8308 4171 8312
rect 4184 8313 4188 8317
rect 4263 8321 4267 8325
rect 4279 8321 4283 8327
rect 4300 8321 4304 8325
rect 4316 8321 4320 8325
rect 4198 8310 4202 8314
rect 4235 8308 4239 8312
rect 4255 8308 4259 8312
rect 4299 8308 4303 8312
rect 4316 8313 4320 8317
rect 3721 8301 3727 8305
rect 2812 8294 2818 8298
rect 2857 8294 2861 8298
rect 2908 8294 2912 8298
rect 2958 8294 2962 8298
rect 2989 8294 2993 8298
rect 3040 8294 3044 8298
rect 3090 8294 3094 8298
rect 3121 8294 3125 8298
rect 3172 8294 3176 8298
rect 3222 8294 3226 8298
rect 3253 8294 3257 8298
rect 3304 8294 3308 8298
rect 3354 8294 3358 8298
rect 2607 8288 2611 8292
rect 2623 8288 2627 8292
rect 3457 8288 3461 8292
rect 3473 8288 3477 8294
rect 3507 8294 3511 8298
rect 3494 8288 3498 8292
rect 2505 8277 2509 8281
rect 2542 8275 2546 8279
rect 2562 8275 2566 8279
rect 2606 8275 2610 8279
rect 2764 8281 2770 8285
rect 2855 8281 2859 8285
rect 2889 8281 2893 8285
rect 2906 8281 2910 8285
rect 2962 8281 2966 8285
rect 2979 8281 2983 8285
rect 3007 8281 3011 8285
rect 3515 8288 3519 8292
rect 3531 8288 3535 8294
rect 3757 8294 3763 8298
rect 3802 8294 3806 8298
rect 3853 8294 3857 8298
rect 3903 8294 3907 8298
rect 3934 8294 3938 8298
rect 3985 8294 3989 8298
rect 4035 8294 4039 8298
rect 4066 8294 4070 8298
rect 4117 8294 4121 8298
rect 4167 8294 4171 8298
rect 4198 8294 4202 8298
rect 4249 8294 4253 8298
rect 4299 8294 4303 8298
rect 3552 8288 3556 8292
rect 3568 8288 3572 8292
rect 2800 8274 2806 8278
rect 2882 8274 2886 8278
rect 2913 8274 2917 8278
rect 2935 8274 2939 8278
rect 3000 8274 3004 8278
rect 2776 8268 2782 8272
rect 2505 8261 2509 8265
rect 2556 8261 2560 8265
rect 2606 8261 2610 8265
rect 2812 8261 2818 8265
rect 2856 8264 2860 8268
rect 2881 8267 2885 8271
rect 2888 8264 2892 8268
rect 2906 8264 2910 8268
rect 2928 8267 2932 8271
rect 2953 8267 2957 8271
rect 2963 8264 2967 8268
rect 2979 8264 2983 8268
rect 2999 8267 3003 8271
rect 3006 8264 3010 8268
rect 3070 8274 3074 8278
rect 2623 8254 2627 8258
rect 2490 8245 2494 8249
rect 2615 8247 2619 8251
rect 2639 8247 2643 8251
rect 2498 8238 2502 8242
rect 2639 8238 2643 8242
rect 2883 8248 2887 8252
rect 2903 8245 2907 8249
rect 2922 8249 2926 8253
rect 3024 8260 3028 8264
rect 3039 8260 3043 8264
rect 2941 8248 2945 8252
rect 2960 8248 2964 8252
rect 2973 8247 2977 8251
rect 2995 8248 2999 8252
rect 3003 8247 3007 8251
rect 3015 8247 3019 8251
rect 2856 8234 2860 8238
rect 2888 8234 2892 8238
rect 2906 8234 2910 8238
rect 2963 8234 2967 8238
rect 2978 8234 2982 8238
rect 3006 8234 3010 8238
rect 2505 8230 2509 8234
rect 2572 8230 2576 8234
rect 2608 8230 2612 8234
rect 2824 8230 2830 8234
rect 2870 8230 2874 8234
rect 2913 8229 2917 8233
rect 2935 8230 2942 8234
rect 2985 8229 2989 8233
rect 2764 8223 2770 8227
rect 2505 8216 2509 8220
rect 2558 8216 2562 8220
rect 2608 8216 2612 8220
rect 2788 8222 2794 8226
rect 2870 8222 2874 8226
rect 2929 8222 2933 8226
rect 2954 8222 2958 8226
rect 2985 8222 2989 8226
rect 3078 8252 3082 8260
rect 3151 8274 3155 8278
rect 3105 8260 3109 8264
rect 3120 8260 3124 8264
rect 3450 8277 3454 8281
rect 3487 8275 3491 8279
rect 3507 8275 3511 8279
rect 3551 8275 3555 8279
rect 3709 8281 3715 8285
rect 3800 8281 3804 8285
rect 3834 8281 3838 8285
rect 3851 8281 3855 8285
rect 3907 8281 3911 8285
rect 3924 8281 3928 8285
rect 3952 8281 3956 8285
rect 3745 8274 3751 8278
rect 3827 8274 3831 8278
rect 3858 8274 3862 8278
rect 3880 8274 3884 8278
rect 3945 8274 3949 8278
rect 3101 8252 3105 8256
rect 3047 8246 3051 8250
rect 3060 8238 3064 8242
rect 3159 8252 3163 8260
rect 3721 8268 3727 8272
rect 3450 8261 3454 8265
rect 3501 8261 3505 8265
rect 3551 8261 3555 8265
rect 3757 8261 3763 8265
rect 3801 8264 3805 8268
rect 3826 8267 3830 8271
rect 3833 8264 3837 8268
rect 3851 8264 3855 8268
rect 3873 8267 3877 8271
rect 3898 8267 3902 8271
rect 3908 8264 3912 8268
rect 3924 8264 3928 8268
rect 3944 8267 3948 8271
rect 3951 8264 3955 8268
rect 4015 8274 4019 8278
rect 3186 8252 3190 8256
rect 3568 8254 3572 8258
rect 3128 8246 3132 8250
rect 3435 8245 3439 8249
rect 3560 8247 3564 8251
rect 3584 8247 3588 8251
rect 3141 8238 3145 8242
rect 3443 8238 3447 8242
rect 3584 8238 3588 8242
rect 3828 8248 3832 8252
rect 3848 8245 3852 8249
rect 3867 8249 3871 8253
rect 3969 8260 3973 8264
rect 3984 8260 3988 8264
rect 3886 8248 3890 8252
rect 3905 8248 3909 8252
rect 3918 8247 3922 8251
rect 3940 8248 3944 8252
rect 3948 8247 3952 8251
rect 3960 8247 3964 8251
rect 3801 8234 3805 8238
rect 3833 8234 3837 8238
rect 3851 8234 3855 8238
rect 3908 8234 3912 8238
rect 3923 8234 3927 8238
rect 3951 8234 3955 8238
rect 3450 8230 3454 8234
rect 3517 8230 3521 8234
rect 3553 8230 3557 8234
rect 3769 8230 3775 8234
rect 3815 8230 3819 8234
rect 3858 8229 3862 8233
rect 3880 8230 3887 8234
rect 3930 8229 3934 8233
rect 3709 8223 3715 8227
rect 2776 8215 2782 8219
rect 2856 8215 2860 8219
rect 2870 8215 2874 8219
rect 2888 8215 2892 8219
rect 2906 8215 2910 8219
rect 2929 8215 2933 8219
rect 2963 8215 2967 8219
rect 2978 8215 2982 8219
rect 3006 8215 3010 8219
rect 2527 8205 2531 8209
rect 2490 8199 2494 8205
rect 2506 8199 2510 8205
rect 2543 8199 2547 8205
rect 2551 8201 2555 8205
rect 2585 8205 2589 8209
rect 2788 8208 2794 8212
rect 2870 8208 2874 8212
rect 2929 8208 2933 8212
rect 2954 8208 2958 8212
rect 2985 8208 2989 8212
rect 2564 8199 2568 8205
rect 2601 8199 2605 8205
rect 2870 8200 2874 8204
rect 2913 8201 2917 8205
rect 2935 8200 2942 8204
rect 2985 8201 2989 8205
rect 2623 8196 2627 8200
rect 2856 8196 2860 8200
rect 2888 8196 2892 8200
rect 2906 8196 2910 8200
rect 2963 8196 2967 8200
rect 2978 8196 2982 8200
rect 3006 8196 3010 8200
rect 2490 8186 2494 8190
rect 2506 8186 2510 8190
rect 2551 8192 2555 8196
rect 2527 8186 2531 8192
rect 2543 8186 2547 8190
rect 2564 8186 2568 8190
rect 2585 8186 2589 8192
rect 2601 8186 2605 8190
rect 2851 8184 2855 8188
rect 2507 8173 2511 8177
rect 2551 8173 2555 8177
rect 2571 8173 2575 8177
rect 2608 8175 2612 8179
rect 2883 8182 2887 8186
rect 2903 8185 2907 8189
rect 2922 8181 2926 8185
rect 2941 8182 2945 8186
rect 2960 8182 2964 8186
rect 2973 8183 2977 8187
rect 3070 8198 3074 8202
rect 3450 8216 3454 8220
rect 3503 8216 3507 8220
rect 3553 8216 3557 8220
rect 3733 8222 3739 8226
rect 3815 8222 3819 8226
rect 3874 8222 3878 8226
rect 3899 8222 3903 8226
rect 3930 8222 3934 8226
rect 4023 8252 4027 8260
rect 4096 8274 4100 8278
rect 4050 8260 4054 8264
rect 4065 8260 4069 8264
rect 4046 8252 4050 8256
rect 3992 8246 3996 8250
rect 4005 8238 4009 8242
rect 4104 8252 4108 8260
rect 4131 8252 4135 8256
rect 4073 8246 4077 8250
rect 4086 8238 4090 8242
rect 3721 8215 3727 8219
rect 3801 8215 3805 8219
rect 3815 8215 3819 8219
rect 3833 8215 3837 8219
rect 3851 8215 3855 8219
rect 3874 8215 3878 8219
rect 3908 8215 3912 8219
rect 3923 8215 3927 8219
rect 3951 8215 3955 8219
rect 3472 8205 3476 8209
rect 3151 8198 3155 8202
rect 3435 8199 3439 8205
rect 3451 8199 3455 8205
rect 3488 8199 3492 8205
rect 3496 8201 3500 8205
rect 3530 8205 3534 8209
rect 3733 8208 3739 8212
rect 3815 8208 3819 8212
rect 3874 8208 3878 8212
rect 3899 8208 3903 8212
rect 3930 8208 3934 8212
rect 3509 8199 3513 8205
rect 3546 8199 3550 8205
rect 3815 8200 3819 8204
rect 3858 8201 3862 8205
rect 3880 8200 3887 8204
rect 3930 8201 3934 8205
rect 3568 8196 3572 8200
rect 3801 8196 3805 8200
rect 3833 8196 3837 8200
rect 3851 8196 3855 8200
rect 3908 8196 3912 8200
rect 3923 8196 3927 8200
rect 3951 8196 3955 8200
rect 2995 8182 2999 8186
rect 3003 8183 3007 8187
rect 3015 8183 3019 8187
rect 3050 8183 3054 8187
rect 3078 8182 3082 8186
rect 3130 8183 3134 8187
rect 3435 8186 3439 8190
rect 3451 8186 3455 8190
rect 3496 8192 3500 8196
rect 3472 8186 3476 8192
rect 3488 8186 3492 8190
rect 3159 8182 3163 8186
rect 3509 8186 3513 8190
rect 3530 8186 3534 8192
rect 3546 8186 3550 8190
rect 3796 8184 3800 8188
rect 2776 8166 2782 8170
rect 2856 8166 2860 8170
rect 2881 8163 2885 8167
rect 2888 8166 2892 8170
rect 2906 8166 2910 8170
rect 2928 8163 2932 8167
rect 2953 8163 2957 8167
rect 2963 8166 2967 8170
rect 2979 8166 2983 8170
rect 2999 8163 3003 8167
rect 3006 8166 3010 8170
rect 2507 8159 2511 8163
rect 2557 8159 2561 8163
rect 2608 8159 2612 8163
rect 2812 8159 2818 8163
rect 2866 8156 2870 8160
rect 2882 8156 2886 8160
rect 2913 8156 2917 8160
rect 2935 8156 2939 8160
rect 3000 8156 3004 8160
rect 3060 8162 3064 8166
rect 3452 8173 3456 8177
rect 3496 8173 3500 8177
rect 3516 8173 3520 8177
rect 3553 8175 3557 8179
rect 3828 8182 3832 8186
rect 3848 8185 3852 8189
rect 3867 8181 3871 8185
rect 3886 8182 3890 8186
rect 3905 8182 3909 8186
rect 3918 8183 3922 8187
rect 4015 8198 4019 8202
rect 4096 8198 4100 8202
rect 3940 8182 3944 8186
rect 3948 8183 3952 8187
rect 3960 8183 3964 8187
rect 3995 8183 3999 8187
rect 4023 8182 4027 8186
rect 4075 8183 4079 8187
rect 4104 8182 4108 8186
rect 3721 8166 3727 8170
rect 3801 8166 3805 8170
rect 3141 8162 3145 8166
rect 3826 8163 3830 8167
rect 3833 8166 3837 8170
rect 3851 8166 3855 8170
rect 3873 8163 3877 8167
rect 3898 8163 3902 8167
rect 3908 8166 3912 8170
rect 3924 8166 3928 8170
rect 3944 8163 3948 8167
rect 3951 8166 3955 8170
rect 3452 8159 3456 8163
rect 3502 8159 3506 8163
rect 3553 8159 3557 8163
rect 3757 8159 3763 8163
rect 3811 8156 3815 8160
rect 3827 8156 3831 8160
rect 3858 8156 3862 8160
rect 3880 8156 3884 8160
rect 3945 8156 3949 8160
rect 4005 8162 4009 8166
rect 4086 8162 4090 8166
rect 2764 8149 2770 8153
rect 2855 8149 2859 8153
rect 2889 8149 2893 8153
rect 2906 8149 2910 8153
rect 2962 8149 2966 8153
rect 2979 8149 2983 8153
rect 3007 8149 3011 8153
rect 3709 8149 3715 8153
rect 3800 8149 3804 8153
rect 3834 8149 3838 8153
rect 3851 8149 3855 8153
rect 3907 8149 3911 8153
rect 3924 8149 3928 8153
rect 3952 8149 3956 8153
rect 2800 8142 2806 8146
rect 2866 8142 2870 8146
rect 2882 8142 2886 8146
rect 2913 8142 2917 8146
rect 2935 8142 2939 8146
rect 3000 8142 3004 8146
rect 3070 8142 3074 8146
rect 2856 8132 2860 8136
rect 2881 8135 2885 8139
rect 2888 8132 2892 8136
rect 2906 8132 2910 8136
rect 2928 8135 2932 8139
rect 2953 8135 2957 8139
rect 2963 8132 2967 8136
rect 2979 8132 2983 8136
rect 2999 8135 3003 8139
rect 3006 8132 3010 8136
rect 2850 8115 2854 8119
rect 2883 8116 2887 8120
rect 2903 8113 2907 8117
rect 2922 8117 2926 8121
rect 2941 8116 2945 8120
rect 2960 8116 2964 8120
rect 2973 8115 2977 8119
rect 2995 8116 2999 8120
rect 3003 8115 3007 8119
rect 3015 8115 3019 8119
rect 3078 8120 3082 8128
rect 3175 8142 3179 8146
rect 3129 8128 3133 8132
rect 3144 8128 3148 8132
rect 3745 8142 3751 8146
rect 3811 8142 3815 8146
rect 3827 8142 3831 8146
rect 3858 8142 3862 8146
rect 3880 8142 3884 8146
rect 3945 8142 3949 8146
rect 4015 8142 4019 8146
rect 3047 8114 3051 8118
rect 3101 8119 3105 8123
rect 2856 8102 2860 8106
rect 2888 8102 2892 8106
rect 2906 8102 2910 8106
rect 2963 8102 2967 8106
rect 2978 8102 2982 8106
rect 3006 8102 3010 8106
rect 2870 8098 2874 8102
rect 2913 8097 2917 8101
rect 2935 8098 2942 8102
rect 2985 8097 2989 8101
rect 2788 8090 2794 8094
rect 2870 8090 2874 8094
rect 2929 8090 2933 8094
rect 2954 8090 2958 8094
rect 2985 8090 2989 8094
rect 618 8085 622 8089
rect 628 8085 632 8089
rect 638 8085 642 8089
rect 618 8080 622 8084
rect 628 8080 632 8084
rect 638 8080 642 8084
rect 618 8075 622 8079
rect 628 8075 632 8079
rect 638 8075 642 8079
rect 618 8070 622 8074
rect 628 8070 632 8074
rect 638 8070 642 8074
rect 664 8085 668 8089
rect 674 8085 678 8089
rect 684 8085 688 8089
rect 3060 8106 3064 8110
rect 3183 8120 3187 8128
rect 3801 8132 3805 8136
rect 3826 8135 3830 8139
rect 3833 8132 3837 8136
rect 3851 8132 3855 8136
rect 3873 8135 3877 8139
rect 3898 8135 3902 8139
rect 3908 8132 3912 8136
rect 3924 8132 3928 8136
rect 3944 8135 3948 8139
rect 3951 8132 3955 8136
rect 3204 8120 3208 8124
rect 3152 8114 3156 8118
rect 3795 8115 3799 8119
rect 3165 8106 3169 8110
rect 3828 8116 3832 8120
rect 3848 8113 3852 8117
rect 3867 8117 3871 8121
rect 3886 8116 3890 8120
rect 3905 8116 3909 8120
rect 3918 8115 3922 8119
rect 3940 8116 3944 8120
rect 3948 8115 3952 8119
rect 3960 8115 3964 8119
rect 4023 8120 4027 8128
rect 4120 8142 4124 8146
rect 4074 8128 4078 8132
rect 4089 8128 4093 8132
rect 3992 8114 3996 8118
rect 4046 8119 4050 8123
rect 3801 8102 3805 8106
rect 3833 8102 3837 8106
rect 3851 8102 3855 8106
rect 3908 8102 3912 8106
rect 3923 8102 3927 8106
rect 3951 8102 3955 8106
rect 3815 8098 3819 8102
rect 3858 8097 3862 8101
rect 3880 8098 3887 8102
rect 3930 8097 3934 8101
rect 3733 8090 3739 8094
rect 3815 8090 3819 8094
rect 3874 8090 3878 8094
rect 3899 8090 3903 8094
rect 3930 8090 3934 8094
rect 4005 8106 4009 8110
rect 4128 8120 4132 8128
rect 4484 8129 4488 8133
rect 4494 8129 4498 8133
rect 4504 8129 4508 8133
rect 4484 8124 4488 8128
rect 4494 8124 4498 8128
rect 4504 8124 4508 8128
rect 4149 8120 4153 8124
rect 4097 8114 4101 8118
rect 4484 8119 4488 8123
rect 4494 8119 4498 8123
rect 4504 8119 4508 8123
rect 4484 8114 4488 8118
rect 4494 8114 4498 8118
rect 4504 8114 4508 8118
rect 4530 8129 4534 8133
rect 4540 8129 4544 8133
rect 4550 8129 4554 8133
rect 4530 8124 4534 8128
rect 4540 8124 4544 8128
rect 4550 8124 4554 8128
rect 4530 8119 4534 8123
rect 4540 8119 4544 8123
rect 4550 8119 4554 8123
rect 4530 8114 4534 8118
rect 4540 8114 4544 8118
rect 4550 8114 4554 8118
rect 4110 8106 4114 8110
rect 4484 8098 4488 8102
rect 4494 8098 4498 8102
rect 4504 8098 4508 8102
rect 4484 8093 4488 8097
rect 4494 8093 4498 8097
rect 4504 8093 4508 8097
rect 4484 8088 4488 8092
rect 4494 8088 4498 8092
rect 4504 8088 4508 8092
rect 664 8080 668 8084
rect 674 8080 678 8084
rect 684 8080 688 8084
rect 2776 8083 2782 8087
rect 2856 8083 2860 8087
rect 2870 8083 2874 8087
rect 2888 8083 2892 8087
rect 2906 8083 2910 8087
rect 2929 8083 2933 8087
rect 2963 8083 2967 8087
rect 2978 8083 2982 8087
rect 3006 8083 3010 8087
rect 3721 8083 3727 8087
rect 3801 8083 3805 8087
rect 3815 8083 3819 8087
rect 3833 8083 3837 8087
rect 3851 8083 3855 8087
rect 3874 8083 3878 8087
rect 3908 8083 3912 8087
rect 3923 8083 3927 8087
rect 3951 8083 3955 8087
rect 4484 8083 4488 8087
rect 4494 8083 4498 8087
rect 4504 8083 4508 8087
rect 4530 8098 4534 8102
rect 4540 8098 4544 8102
rect 4550 8098 4554 8102
rect 4530 8093 4534 8097
rect 4540 8093 4544 8097
rect 4550 8093 4554 8097
rect 4530 8088 4534 8092
rect 4540 8088 4544 8092
rect 4550 8088 4554 8092
rect 4530 8083 4534 8087
rect 4540 8083 4544 8087
rect 4550 8083 4554 8087
rect 664 8075 668 8079
rect 674 8075 678 8079
rect 684 8075 688 8079
rect 2788 8076 2794 8080
rect 2870 8076 2874 8080
rect 2929 8076 2933 8080
rect 2954 8076 2958 8080
rect 2985 8076 2989 8080
rect 664 8070 668 8074
rect 674 8070 678 8074
rect 684 8070 688 8074
rect 2870 8068 2874 8072
rect 2913 8069 2917 8073
rect 2935 8068 2942 8072
rect 2985 8069 2989 8073
rect 2856 8064 2860 8068
rect 2888 8064 2892 8068
rect 2906 8064 2910 8068
rect 2963 8064 2967 8068
rect 2978 8064 2982 8068
rect 3006 8064 3010 8068
rect 3070 8067 3074 8071
rect 3733 8076 3739 8080
rect 3815 8076 3819 8080
rect 3874 8076 3878 8080
rect 3899 8076 3903 8080
rect 3930 8076 3934 8080
rect 3175 8067 3179 8071
rect 3815 8068 3819 8072
rect 3858 8069 3862 8073
rect 3880 8068 3887 8072
rect 3930 8069 3934 8073
rect 3801 8064 3805 8068
rect 3833 8064 3837 8068
rect 3851 8064 3855 8068
rect 3908 8064 3912 8068
rect 3923 8064 3927 8068
rect 3951 8064 3955 8068
rect 4015 8067 4019 8071
rect 4506 8074 4510 8078
rect 4511 8074 4515 8078
rect 4120 8067 4124 8071
rect 4506 8069 4510 8073
rect 4511 8069 4515 8073
rect 4506 8064 4510 8068
rect 4511 8064 4515 8068
rect 2851 8052 2855 8056
rect 2883 8050 2887 8054
rect 2903 8053 2907 8057
rect 2922 8049 2926 8053
rect 2941 8050 2945 8054
rect 2960 8050 2964 8054
rect 2973 8051 2977 8055
rect 2995 8050 2999 8054
rect 3003 8051 3007 8055
rect 3015 8051 3019 8055
rect 3049 8052 3053 8056
rect 3078 8051 3082 8055
rect 3155 8052 3159 8056
rect 3183 8051 3187 8055
rect 3796 8052 3800 8056
rect 2856 8034 2860 8038
rect 2881 8031 2885 8035
rect 2888 8034 2892 8038
rect 2906 8034 2910 8038
rect 2928 8031 2932 8035
rect 2953 8031 2957 8035
rect 2963 8034 2967 8038
rect 2979 8034 2983 8038
rect 2999 8031 3003 8035
rect 3006 8034 3010 8038
rect 2800 8024 2806 8028
rect 2882 8024 2886 8028
rect 2913 8024 2917 8028
rect 2935 8024 2939 8028
rect 3000 8024 3004 8028
rect 3060 8031 3064 8035
rect 3828 8050 3832 8054
rect 3848 8053 3852 8057
rect 3867 8049 3871 8053
rect 3886 8050 3890 8054
rect 3905 8050 3909 8054
rect 3918 8051 3922 8055
rect 3940 8050 3944 8054
rect 3948 8051 3952 8055
rect 3960 8051 3964 8055
rect 3994 8052 3998 8056
rect 4023 8051 4027 8055
rect 4100 8052 4104 8056
rect 4506 8059 4510 8063
rect 4511 8059 4515 8063
rect 4128 8051 4132 8055
rect 4506 8054 4510 8058
rect 4511 8054 4515 8058
rect 4506 8049 4510 8053
rect 4511 8049 4515 8053
rect 4506 8044 4510 8048
rect 4511 8044 4515 8048
rect 3165 8031 3169 8035
rect 3801 8034 3805 8038
rect 3826 8031 3830 8035
rect 3833 8034 3837 8038
rect 3851 8034 3855 8038
rect 3873 8031 3877 8035
rect 3898 8031 3902 8035
rect 3908 8034 3912 8038
rect 3924 8034 3928 8038
rect 3944 8031 3948 8035
rect 3951 8034 3955 8038
rect 3745 8024 3751 8028
rect 3827 8024 3831 8028
rect 3858 8024 3862 8028
rect 3880 8024 3884 8028
rect 3945 8024 3949 8028
rect 4005 8031 4009 8035
rect 4506 8039 4510 8043
rect 4511 8039 4515 8043
rect 4110 8031 4114 8035
rect 4506 8034 4510 8038
rect 4511 8034 4515 8038
rect 4506 8029 4510 8033
rect 4511 8029 4515 8033
rect 4506 8024 4510 8028
rect 4511 8024 4515 8028
rect 2764 8017 2770 8021
rect 2855 8017 2859 8021
rect 2889 8017 2893 8021
rect 2906 8017 2910 8021
rect 2962 8017 2966 8021
rect 2979 8017 2983 8021
rect 3007 8017 3011 8021
rect 3709 8017 3715 8021
rect 3800 8017 3804 8021
rect 3834 8017 3838 8021
rect 3851 8017 3855 8021
rect 3907 8017 3911 8021
rect 3924 8017 3928 8021
rect 3952 8017 3956 8021
rect 2800 8010 2806 8014
rect 2882 8010 2886 8014
rect 2913 8010 2917 8014
rect 2935 8010 2939 8014
rect 3000 8010 3004 8014
rect 3070 8010 3074 8014
rect 2856 8000 2860 8004
rect 2881 8003 2885 8007
rect 2888 8000 2892 8004
rect 2906 8000 2910 8004
rect 2928 8003 2932 8007
rect 2953 8003 2957 8007
rect 2963 8000 2967 8004
rect 2979 8000 2983 8004
rect 2999 8003 3003 8007
rect 3006 8000 3010 8004
rect 2850 7983 2854 7987
rect 2883 7984 2887 7988
rect 2903 7981 2907 7985
rect 2922 7985 2926 7989
rect 2941 7984 2945 7988
rect 2960 7984 2964 7988
rect 2973 7983 2977 7987
rect 2995 7984 2999 7988
rect 3003 7983 3007 7987
rect 3015 7983 3019 7987
rect 3078 7988 3082 7996
rect 3151 8010 3155 8014
rect 3105 7996 3109 8000
rect 3120 7996 3124 8000
rect 3101 7988 3105 7992
rect 3047 7982 3051 7986
rect 2856 7970 2860 7974
rect 2888 7970 2892 7974
rect 2906 7970 2910 7974
rect 2963 7970 2967 7974
rect 2978 7970 2982 7974
rect 3006 7970 3010 7974
rect 2870 7966 2874 7970
rect 2913 7965 2917 7969
rect 2935 7966 2942 7970
rect 2985 7965 2989 7969
rect 2788 7958 2794 7962
rect 2870 7958 2874 7962
rect 2929 7958 2933 7962
rect 2954 7958 2958 7962
rect 2985 7958 2989 7962
rect 3060 7974 3064 7978
rect 3159 7988 3163 7996
rect 3241 8010 3245 8014
rect 3195 7996 3199 8000
rect 3210 7996 3214 8000
rect 3745 8010 3751 8014
rect 3827 8010 3831 8014
rect 3858 8010 3862 8014
rect 3880 8010 3884 8014
rect 3945 8010 3949 8014
rect 4015 8010 4019 8014
rect 3183 7988 3187 7992
rect 3128 7982 3132 7986
rect 3217 7990 3221 7994
rect 3249 7988 3253 7996
rect 3801 8000 3805 8004
rect 3826 8003 3830 8007
rect 3833 8000 3837 8004
rect 3851 8000 3855 8004
rect 3873 8003 3877 8007
rect 3898 8003 3902 8007
rect 3908 8000 3912 8004
rect 3924 8000 3928 8004
rect 3944 8003 3948 8007
rect 3951 8000 3955 8004
rect 3141 7974 3145 7978
rect 3284 7987 3288 7991
rect 3795 7983 3799 7987
rect 3231 7974 3235 7978
rect 3828 7984 3832 7988
rect 3848 7981 3852 7985
rect 3867 7985 3871 7989
rect 3886 7984 3890 7988
rect 3905 7984 3909 7988
rect 3918 7983 3922 7987
rect 3940 7984 3944 7988
rect 3948 7983 3952 7987
rect 3960 7983 3964 7987
rect 4023 7988 4027 7996
rect 4096 8010 4100 8014
rect 4050 7996 4054 8000
rect 4065 7996 4069 8000
rect 4046 7988 4050 7992
rect 3992 7982 3996 7986
rect 3801 7970 3805 7974
rect 3833 7970 3837 7974
rect 3851 7970 3855 7974
rect 3908 7970 3912 7974
rect 3923 7970 3927 7974
rect 3951 7970 3955 7974
rect 3815 7966 3819 7970
rect 3858 7965 3862 7969
rect 3880 7966 3887 7970
rect 3930 7965 3934 7969
rect 3733 7958 3739 7962
rect 3815 7958 3819 7962
rect 3874 7958 3878 7962
rect 3899 7958 3903 7962
rect 3930 7958 3934 7962
rect 4005 7974 4009 7978
rect 4104 7988 4108 7996
rect 4186 8010 4190 8014
rect 4140 7996 4144 8000
rect 4155 7996 4159 8000
rect 4128 7988 4132 7992
rect 4073 7982 4077 7986
rect 4162 7990 4166 7994
rect 4194 7988 4198 7996
rect 4086 7974 4090 7978
rect 4229 7987 4233 7991
rect 4574 7982 4578 7986
rect 4176 7974 4180 7978
rect 4590 7982 4594 7986
rect 4606 7982 4610 7986
rect 4622 7982 4626 7986
rect 4645 7982 4649 7986
rect 4661 7982 4665 7986
rect 4688 7982 4692 7986
rect 4704 7982 4708 7986
rect 4729 7982 4733 7986
rect 4745 7982 4749 7986
rect 2776 7951 2782 7955
rect 2856 7951 2860 7955
rect 2870 7951 2874 7955
rect 2888 7951 2892 7955
rect 2906 7951 2910 7955
rect 2929 7951 2933 7955
rect 2963 7951 2967 7955
rect 2978 7951 2982 7955
rect 3006 7951 3010 7955
rect 3721 7951 3727 7955
rect 3801 7951 3805 7955
rect 3815 7951 3819 7955
rect 3833 7951 3837 7955
rect 3851 7951 3855 7955
rect 3874 7951 3878 7955
rect 3908 7951 3912 7955
rect 3923 7951 3927 7955
rect 3951 7951 3955 7955
rect 2788 7944 2794 7948
rect 2870 7944 2874 7948
rect 2929 7944 2933 7948
rect 2954 7944 2958 7948
rect 2985 7944 2989 7948
rect 2870 7936 2874 7940
rect 2913 7937 2917 7941
rect 2935 7936 2942 7940
rect 2985 7937 2989 7941
rect 2856 7932 2860 7936
rect 2888 7932 2892 7936
rect 2906 7932 2910 7936
rect 2963 7932 2967 7936
rect 2978 7932 2982 7936
rect 3006 7932 3010 7936
rect 2851 7920 2855 7924
rect 2883 7918 2887 7922
rect 2903 7921 2907 7925
rect 2922 7917 2926 7921
rect 2941 7918 2945 7922
rect 2960 7918 2964 7922
rect 2973 7919 2977 7923
rect 3070 7932 3074 7936
rect 3151 7932 3155 7936
rect 3733 7944 3739 7948
rect 3815 7944 3819 7948
rect 3874 7944 3878 7948
rect 3899 7944 3903 7948
rect 3930 7944 3934 7948
rect 3815 7936 3819 7940
rect 3858 7937 3862 7941
rect 3880 7936 3887 7940
rect 3930 7937 3934 7941
rect 3241 7932 3245 7936
rect 3801 7932 3805 7936
rect 3833 7932 3837 7936
rect 3851 7932 3855 7936
rect 3908 7932 3912 7936
rect 3923 7932 3927 7936
rect 3951 7932 3955 7936
rect 2995 7918 2999 7922
rect 3003 7919 3007 7923
rect 3015 7919 3019 7923
rect 3050 7917 3054 7921
rect 3078 7916 3082 7920
rect 3130 7917 3134 7921
rect 3159 7916 3163 7920
rect 3214 7917 3218 7921
rect 3796 7920 3800 7924
rect 3249 7916 3253 7920
rect 2856 7902 2860 7906
rect 2881 7899 2885 7903
rect 2888 7902 2892 7906
rect 2906 7902 2910 7906
rect 2928 7899 2932 7903
rect 2953 7899 2957 7903
rect 2963 7902 2967 7906
rect 2979 7902 2983 7906
rect 2999 7899 3003 7903
rect 3006 7902 3010 7906
rect 3828 7918 3832 7922
rect 3848 7921 3852 7925
rect 3867 7917 3871 7921
rect 3886 7918 3890 7922
rect 3905 7918 3909 7922
rect 3918 7919 3922 7923
rect 4015 7932 4019 7936
rect 4096 7932 4100 7936
rect 4360 7950 4369 7963
rect 4659 7954 4667 7963
rect 4703 7954 4711 7963
rect 4186 7932 4190 7936
rect 3940 7918 3944 7922
rect 3948 7919 3952 7923
rect 3960 7919 3964 7923
rect 3995 7917 3999 7921
rect 4023 7916 4027 7920
rect 4075 7917 4079 7921
rect 4104 7916 4108 7920
rect 4159 7917 4163 7921
rect 4574 7924 4578 7928
rect 4194 7916 4198 7920
rect 2800 7892 2806 7896
rect 2882 7892 2886 7896
rect 2913 7892 2917 7896
rect 2935 7892 2939 7896
rect 3000 7892 3004 7896
rect 3060 7896 3064 7900
rect 3141 7896 3145 7900
rect 3801 7902 3805 7906
rect 3231 7896 3235 7900
rect 3826 7899 3830 7903
rect 3833 7902 3837 7906
rect 3851 7902 3855 7906
rect 3873 7899 3877 7903
rect 3898 7899 3902 7903
rect 3908 7902 3912 7906
rect 3924 7902 3928 7906
rect 3944 7899 3948 7903
rect 3951 7902 3955 7906
rect 3745 7892 3751 7896
rect 3827 7892 3831 7896
rect 3858 7892 3862 7896
rect 3880 7892 3884 7896
rect 3945 7892 3949 7896
rect 4005 7896 4009 7900
rect 4086 7896 4090 7900
rect 4176 7896 4180 7900
rect 4590 7924 4594 7928
rect 4606 7924 4610 7928
rect 4622 7924 4626 7928
rect 2764 7885 2770 7889
rect 2855 7885 2859 7889
rect 2889 7885 2893 7889
rect 2906 7885 2910 7889
rect 2962 7885 2966 7889
rect 2979 7885 2983 7889
rect 3007 7885 3011 7889
rect 3709 7885 3715 7889
rect 3800 7885 3804 7889
rect 3834 7885 3838 7889
rect 3851 7885 3855 7889
rect 3907 7885 3911 7889
rect 3924 7885 3928 7889
rect 3952 7885 3956 7889
rect 2800 7878 2806 7882
rect 2882 7878 2886 7882
rect 2913 7878 2917 7882
rect 2935 7878 2939 7882
rect 3000 7878 3004 7882
rect 3070 7878 3074 7882
rect 2856 7868 2860 7872
rect 2881 7871 2885 7875
rect 2888 7868 2892 7872
rect 2906 7868 2910 7872
rect 2928 7871 2932 7875
rect 2953 7871 2957 7875
rect 2963 7868 2967 7872
rect 2979 7868 2983 7872
rect 2999 7871 3003 7875
rect 3006 7868 3010 7872
rect 2850 7851 2854 7855
rect 2883 7852 2887 7856
rect 2903 7849 2907 7853
rect 2922 7853 2926 7857
rect 3745 7878 3751 7882
rect 3827 7878 3831 7882
rect 3858 7878 3862 7882
rect 3880 7878 3884 7882
rect 3945 7878 3949 7882
rect 4015 7878 4019 7882
rect 2941 7852 2945 7856
rect 2960 7852 2964 7856
rect 2973 7851 2977 7855
rect 2995 7852 2999 7856
rect 3003 7851 3007 7855
rect 3015 7851 3019 7855
rect 3078 7856 3082 7864
rect 3801 7868 3805 7872
rect 3826 7871 3830 7875
rect 3833 7868 3837 7872
rect 3851 7868 3855 7872
rect 3873 7871 3877 7875
rect 3898 7871 3902 7875
rect 3908 7868 3912 7872
rect 3924 7868 3928 7872
rect 3944 7871 3948 7875
rect 3951 7868 3955 7872
rect 3047 7850 3051 7854
rect 3101 7855 3105 7859
rect 3795 7851 3799 7855
rect 2856 7838 2860 7842
rect 2888 7838 2892 7842
rect 2906 7838 2910 7842
rect 2963 7838 2967 7842
rect 2978 7838 2982 7842
rect 3006 7838 3010 7842
rect 2870 7834 2874 7838
rect 2373 7830 2377 7834
rect 2409 7830 2413 7834
rect 2476 7830 2480 7834
rect 2505 7830 2509 7834
rect 2541 7830 2545 7834
rect 2608 7830 2612 7834
rect 2637 7830 2641 7834
rect 2673 7830 2677 7834
rect 2740 7830 2744 7834
rect 2824 7830 2830 7834
rect 2913 7833 2917 7837
rect 2935 7834 2942 7838
rect 2985 7833 2989 7837
rect 2764 7823 2770 7827
rect 2870 7826 2874 7830
rect 2879 7826 2883 7830
rect 2929 7826 2933 7830
rect 2954 7826 2958 7830
rect 2985 7826 2989 7830
rect 3060 7842 3064 7846
rect 3828 7852 3832 7856
rect 3848 7849 3852 7853
rect 3867 7853 3871 7857
rect 3886 7852 3890 7856
rect 3905 7852 3909 7856
rect 3918 7851 3922 7855
rect 3940 7852 3944 7856
rect 3948 7851 3952 7855
rect 3960 7851 3964 7855
rect 4023 7856 4027 7864
rect 3992 7850 3996 7854
rect 4046 7855 4050 7859
rect 3801 7838 3805 7842
rect 3833 7838 3837 7842
rect 3851 7838 3855 7842
rect 3908 7838 3912 7842
rect 3923 7838 3927 7842
rect 3951 7838 3955 7842
rect 3815 7834 3819 7838
rect 3318 7830 3322 7834
rect 3354 7830 3358 7834
rect 3421 7830 3425 7834
rect 3450 7830 3454 7834
rect 3486 7830 3490 7834
rect 3553 7830 3557 7834
rect 3582 7830 3586 7834
rect 3618 7830 3622 7834
rect 3685 7830 3689 7834
rect 3769 7830 3775 7834
rect 3858 7833 3862 7837
rect 3880 7834 3887 7838
rect 3930 7833 3934 7837
rect 3709 7823 3715 7827
rect 3815 7826 3819 7830
rect 3824 7826 3828 7830
rect 3874 7826 3878 7830
rect 3899 7826 3903 7830
rect 3930 7826 3934 7830
rect 4645 7924 4649 7928
rect 4661 7924 4665 7928
rect 4688 7924 4692 7928
rect 4704 7924 4708 7928
rect 4729 7924 4733 7928
rect 4745 7924 4749 7928
rect 4005 7842 4009 7846
rect 4529 7824 4533 7828
rect 4534 7824 4538 7828
rect 4539 7824 4543 7828
rect 4544 7824 4548 7828
rect 4549 7824 4553 7828
rect 4554 7824 4558 7828
rect 4559 7824 4563 7828
rect 4564 7824 4568 7828
rect 4569 7824 4573 7828
rect 4574 7824 4578 7828
rect 4579 7824 4583 7828
rect 4584 7824 4588 7828
rect 4589 7824 4593 7828
rect 2373 7816 2377 7820
rect 2423 7816 2427 7820
rect 2476 7816 2480 7820
rect 2505 7816 2509 7820
rect 2555 7816 2559 7820
rect 2608 7816 2612 7820
rect 2637 7816 2641 7820
rect 2687 7816 2691 7820
rect 2740 7816 2744 7820
rect 2776 7819 2782 7823
rect 2856 7819 2860 7823
rect 2870 7819 2874 7823
rect 2888 7819 2892 7823
rect 2906 7819 2910 7823
rect 2929 7819 2933 7823
rect 2963 7819 2967 7823
rect 2978 7819 2982 7823
rect 3006 7819 3010 7823
rect 3131 7819 3135 7823
rect 3149 7819 3153 7823
rect 3167 7819 3171 7823
rect 3190 7819 3194 7823
rect 3224 7819 3228 7823
rect 3239 7819 3243 7823
rect 3267 7819 3271 7823
rect 2396 7805 2400 7809
rect 2367 7796 2371 7800
rect 2380 7799 2384 7805
rect 2417 7799 2421 7805
rect 2430 7801 2434 7805
rect 2454 7805 2458 7809
rect 2528 7805 2532 7809
rect 2438 7799 2442 7805
rect 2475 7799 2479 7805
rect 2491 7799 2495 7805
rect 2512 7799 2516 7805
rect 2549 7799 2553 7805
rect 2562 7801 2566 7805
rect 2586 7805 2590 7809
rect 2660 7805 2664 7809
rect 2570 7799 2574 7805
rect 2607 7799 2611 7805
rect 2623 7799 2627 7805
rect 2644 7799 2648 7805
rect 2681 7799 2685 7805
rect 2694 7801 2698 7805
rect 2718 7805 2722 7809
rect 2788 7812 2794 7816
rect 2870 7812 2874 7816
rect 2879 7812 2883 7816
rect 2929 7812 2933 7816
rect 2954 7812 2958 7816
rect 2985 7812 2989 7816
rect 2702 7799 2706 7805
rect 2739 7799 2743 7805
rect 2755 7801 2759 7805
rect 2870 7804 2874 7808
rect 2913 7805 2917 7809
rect 2935 7804 2942 7808
rect 2985 7805 2989 7809
rect 2856 7800 2860 7804
rect 2888 7800 2892 7804
rect 2906 7800 2910 7804
rect 2963 7800 2967 7804
rect 2978 7800 2982 7804
rect 3006 7800 3010 7804
rect 2380 7786 2384 7790
rect 2396 7786 2400 7792
rect 2430 7792 2434 7796
rect 2417 7786 2421 7790
rect 2438 7786 2442 7790
rect 2454 7786 2458 7792
rect 2475 7786 2479 7790
rect 2491 7786 2495 7790
rect 2512 7786 2516 7790
rect 2528 7786 2532 7792
rect 2562 7792 2566 7796
rect 2549 7786 2553 7790
rect 2570 7786 2574 7790
rect 2586 7786 2590 7792
rect 2607 7786 2611 7790
rect 2623 7786 2627 7790
rect 2644 7786 2648 7790
rect 2660 7786 2664 7792
rect 2694 7792 2698 7796
rect 2681 7786 2685 7790
rect 2702 7786 2706 7790
rect 2718 7786 2722 7792
rect 2739 7786 2743 7790
rect 2755 7786 2759 7790
rect 2851 7788 2855 7792
rect 618 7776 622 7780
rect 628 7776 632 7780
rect 638 7776 642 7780
rect 618 7771 622 7775
rect 628 7771 632 7775
rect 638 7771 642 7775
rect 618 7766 622 7770
rect 628 7766 632 7770
rect 638 7766 642 7770
rect 618 7761 622 7765
rect 628 7761 632 7765
rect 638 7761 642 7765
rect 664 7776 668 7780
rect 674 7776 678 7780
rect 684 7776 688 7780
rect 664 7771 668 7775
rect 674 7771 678 7775
rect 684 7771 688 7775
rect 2373 7775 2377 7779
rect 2410 7773 2414 7777
rect 2430 7773 2434 7777
rect 2474 7773 2478 7777
rect 2505 7775 2509 7779
rect 2542 7773 2546 7777
rect 2562 7773 2566 7777
rect 2606 7773 2610 7777
rect 2637 7775 2641 7779
rect 2674 7773 2678 7777
rect 2694 7773 2698 7777
rect 2738 7773 2742 7777
rect 2883 7786 2887 7790
rect 2903 7789 2907 7793
rect 2922 7785 2926 7789
rect 2941 7786 2945 7790
rect 2960 7786 2964 7790
rect 2973 7787 2977 7791
rect 3109 7812 3113 7816
rect 3131 7812 3135 7816
rect 3190 7812 3194 7816
rect 3215 7812 3219 7816
rect 3246 7812 3250 7816
rect 3318 7816 3322 7820
rect 3368 7816 3372 7820
rect 3421 7816 3425 7820
rect 3450 7816 3454 7820
rect 3500 7816 3504 7820
rect 3553 7816 3557 7820
rect 3582 7816 3586 7820
rect 3632 7816 3636 7820
rect 3685 7816 3689 7820
rect 3721 7819 3727 7823
rect 3801 7819 3805 7823
rect 3815 7819 3819 7823
rect 3833 7819 3837 7823
rect 3851 7819 3855 7823
rect 3874 7819 3878 7823
rect 3908 7819 3912 7823
rect 3923 7819 3927 7823
rect 3951 7819 3955 7823
rect 4076 7819 4080 7823
rect 4094 7819 4098 7823
rect 4112 7819 4116 7823
rect 4135 7819 4139 7823
rect 4169 7819 4173 7823
rect 4184 7819 4188 7823
rect 4212 7819 4216 7823
rect 4529 7819 4533 7823
rect 4534 7819 4538 7823
rect 4539 7819 4543 7823
rect 4544 7819 4548 7823
rect 4549 7819 4553 7823
rect 4554 7819 4558 7823
rect 4559 7819 4563 7823
rect 4564 7819 4568 7823
rect 4569 7819 4573 7823
rect 4574 7819 4578 7823
rect 4579 7819 4583 7823
rect 4584 7819 4588 7823
rect 4589 7819 4593 7823
rect 3131 7804 3135 7808
rect 3174 7805 3178 7809
rect 3196 7804 3203 7808
rect 3246 7805 3250 7809
rect 3341 7805 3345 7809
rect 3149 7800 3153 7804
rect 3167 7800 3171 7804
rect 3224 7800 3228 7804
rect 3239 7800 3243 7804
rect 3267 7800 3271 7804
rect 3070 7796 3074 7800
rect 2995 7786 2999 7790
rect 3003 7787 3007 7791
rect 3015 7787 3019 7791
rect 3049 7781 3053 7785
rect 3089 7787 3093 7791
rect 3078 7780 3082 7784
rect 2856 7770 2860 7774
rect 664 7766 668 7770
rect 674 7766 678 7770
rect 684 7766 688 7770
rect 2776 7766 2782 7770
rect 2881 7767 2885 7771
rect 2888 7770 2892 7774
rect 2906 7770 2910 7774
rect 2928 7767 2932 7771
rect 2953 7767 2957 7771
rect 2963 7770 2967 7774
rect 2979 7770 2983 7774
rect 2999 7767 3003 7771
rect 3006 7770 3010 7774
rect 3144 7786 3148 7790
rect 3164 7789 3168 7793
rect 3183 7785 3187 7789
rect 3312 7796 3316 7800
rect 3325 7799 3329 7805
rect 3362 7799 3366 7805
rect 3375 7801 3379 7805
rect 3399 7805 3403 7809
rect 3473 7805 3477 7809
rect 3383 7799 3387 7805
rect 3420 7799 3424 7805
rect 3436 7799 3440 7805
rect 3457 7799 3461 7805
rect 3494 7799 3498 7805
rect 3507 7801 3511 7805
rect 3531 7805 3535 7809
rect 3605 7805 3609 7809
rect 3515 7799 3519 7805
rect 3552 7799 3556 7805
rect 3568 7799 3572 7805
rect 3589 7799 3593 7805
rect 3626 7799 3630 7805
rect 3639 7801 3643 7805
rect 3663 7805 3667 7809
rect 3733 7812 3739 7816
rect 3815 7812 3819 7816
rect 3824 7812 3828 7816
rect 3874 7812 3878 7816
rect 3899 7812 3903 7816
rect 3930 7812 3934 7816
rect 3647 7799 3651 7805
rect 3684 7799 3688 7805
rect 3700 7801 3704 7805
rect 3815 7804 3819 7808
rect 3858 7805 3862 7809
rect 3880 7804 3887 7808
rect 3930 7805 3934 7809
rect 3801 7800 3805 7804
rect 3833 7800 3837 7804
rect 3851 7800 3855 7804
rect 3908 7800 3912 7804
rect 3923 7800 3927 7804
rect 3951 7800 3955 7804
rect 3202 7786 3206 7790
rect 3221 7786 3225 7790
rect 3234 7787 3238 7791
rect 3256 7786 3260 7790
rect 3264 7787 3268 7791
rect 3276 7787 3280 7791
rect 3325 7786 3329 7790
rect 3341 7786 3345 7792
rect 3375 7792 3379 7796
rect 3362 7786 3366 7790
rect 3383 7786 3387 7790
rect 3399 7786 3403 7792
rect 3420 7786 3424 7790
rect 3436 7786 3440 7790
rect 3457 7786 3461 7790
rect 3473 7786 3477 7792
rect 3507 7792 3511 7796
rect 3494 7786 3498 7790
rect 3515 7786 3519 7790
rect 3531 7786 3535 7792
rect 3552 7786 3556 7790
rect 3568 7786 3572 7790
rect 3589 7786 3593 7790
rect 3605 7786 3609 7792
rect 3639 7792 3643 7796
rect 3626 7786 3630 7790
rect 3647 7786 3651 7790
rect 3663 7786 3667 7792
rect 3684 7786 3688 7790
rect 3700 7786 3704 7790
rect 3796 7788 3800 7792
rect 3090 7770 3094 7774
rect 3116 7770 3120 7774
rect 664 7761 668 7765
rect 674 7761 678 7765
rect 684 7761 688 7765
rect 2373 7759 2377 7763
rect 2424 7759 2428 7763
rect 2474 7759 2478 7763
rect 2505 7759 2509 7763
rect 2556 7759 2560 7763
rect 2606 7759 2610 7763
rect 2637 7759 2641 7763
rect 2688 7759 2692 7763
rect 2738 7759 2742 7763
rect 2812 7760 2818 7764
rect 2864 7760 2868 7764
rect 2882 7760 2886 7764
rect 2913 7760 2917 7764
rect 2935 7760 2939 7764
rect 3000 7760 3004 7764
rect 3142 7767 3146 7771
rect 3149 7770 3153 7774
rect 3167 7770 3171 7774
rect 3189 7767 3193 7771
rect 3214 7767 3218 7771
rect 3224 7770 3228 7774
rect 3240 7770 3244 7774
rect 3260 7767 3264 7771
rect 3267 7770 3271 7774
rect 3318 7775 3322 7779
rect 3355 7773 3359 7777
rect 3375 7773 3379 7777
rect 3419 7773 3423 7777
rect 3450 7775 3454 7779
rect 3487 7773 3491 7777
rect 3507 7773 3511 7777
rect 3551 7773 3555 7777
rect 3582 7775 3586 7779
rect 3619 7773 3623 7777
rect 3639 7773 3643 7777
rect 3683 7773 3687 7777
rect 3828 7786 3832 7790
rect 3848 7789 3852 7793
rect 3867 7785 3871 7789
rect 3886 7786 3890 7790
rect 3905 7786 3909 7790
rect 3918 7787 3922 7791
rect 4054 7812 4058 7816
rect 4076 7812 4080 7816
rect 4135 7812 4139 7816
rect 4160 7812 4164 7816
rect 4191 7812 4195 7816
rect 4076 7804 4080 7808
rect 4119 7805 4123 7809
rect 4141 7804 4148 7808
rect 4191 7805 4195 7809
rect 4094 7800 4098 7804
rect 4112 7800 4116 7804
rect 4169 7800 4173 7804
rect 4184 7800 4188 7804
rect 4212 7800 4216 7804
rect 4015 7796 4019 7800
rect 3940 7786 3944 7790
rect 3948 7787 3952 7791
rect 3960 7787 3964 7791
rect 3994 7781 3998 7785
rect 4034 7787 4038 7791
rect 4023 7780 4027 7784
rect 3801 7770 3805 7774
rect 3721 7766 3727 7770
rect 3826 7767 3830 7771
rect 3833 7770 3837 7774
rect 3851 7770 3855 7774
rect 3873 7767 3877 7771
rect 3898 7767 3902 7771
rect 3908 7770 3912 7774
rect 3924 7770 3928 7774
rect 3944 7767 3948 7771
rect 3951 7770 3955 7774
rect 4089 7786 4093 7790
rect 4109 7789 4113 7793
rect 4128 7785 4132 7789
rect 4147 7786 4151 7790
rect 4166 7786 4170 7790
rect 4179 7787 4183 7791
rect 4201 7786 4205 7790
rect 4209 7787 4213 7791
rect 4221 7787 4225 7791
rect 4484 7789 4488 7793
rect 4494 7789 4498 7793
rect 4504 7789 4508 7793
rect 4484 7784 4488 7788
rect 4494 7784 4498 7788
rect 4504 7784 4508 7788
rect 4484 7779 4488 7783
rect 4494 7779 4498 7783
rect 4504 7779 4508 7783
rect 4484 7774 4488 7778
rect 4494 7774 4498 7778
rect 4504 7774 4508 7778
rect 4530 7789 4534 7793
rect 4540 7789 4544 7793
rect 4550 7789 4554 7793
rect 4530 7784 4534 7788
rect 4540 7784 4544 7788
rect 4550 7784 4554 7788
rect 4530 7779 4534 7783
rect 4540 7779 4544 7783
rect 4550 7779 4554 7783
rect 4530 7774 4534 7778
rect 4540 7774 4544 7778
rect 4550 7774 4554 7778
rect 4035 7770 4039 7774
rect 4061 7770 4065 7774
rect 3060 7760 3064 7764
rect 3099 7760 3103 7764
rect 3143 7760 3147 7764
rect 3174 7760 3178 7764
rect 3196 7760 3200 7764
rect 3261 7760 3265 7764
rect 3318 7759 3322 7763
rect 3369 7759 3373 7763
rect 3419 7759 3423 7763
rect 3450 7759 3454 7763
rect 3501 7759 3505 7763
rect 3551 7759 3555 7763
rect 3582 7759 3586 7763
rect 3633 7759 3637 7763
rect 3683 7759 3687 7763
rect 3757 7760 3763 7764
rect 3809 7760 3813 7764
rect 3827 7760 3831 7764
rect 3858 7760 3862 7764
rect 3880 7760 3884 7764
rect 3945 7760 3949 7764
rect 4087 7767 4091 7771
rect 4094 7770 4098 7774
rect 4112 7770 4116 7774
rect 4134 7767 4138 7771
rect 4159 7767 4163 7771
rect 4169 7770 4173 7774
rect 4185 7770 4189 7774
rect 4205 7767 4209 7771
rect 4212 7770 4216 7774
rect 4005 7760 4009 7764
rect 4044 7760 4048 7764
rect 4088 7760 4092 7764
rect 4119 7760 4123 7764
rect 4141 7760 4145 7764
rect 4206 7760 4210 7764
rect 2367 7752 2371 7756
rect 2755 7752 2759 7756
rect 2764 7753 2770 7757
rect 2855 7753 2859 7757
rect 2889 7753 2893 7757
rect 2906 7753 2910 7757
rect 2962 7753 2966 7757
rect 2979 7753 2983 7757
rect 3007 7753 3011 7757
rect 3090 7753 3094 7757
rect 3116 7753 3120 7757
rect 3150 7753 3154 7757
rect 3167 7753 3171 7757
rect 3223 7753 3227 7757
rect 3240 7753 3244 7757
rect 3268 7753 3272 7757
rect 3312 7752 3316 7756
rect 3700 7752 3704 7756
rect 3709 7753 3715 7757
rect 3800 7753 3804 7757
rect 3834 7753 3838 7757
rect 3851 7753 3855 7757
rect 3907 7753 3911 7757
rect 3924 7753 3928 7757
rect 3952 7753 3956 7757
rect 4035 7753 4039 7757
rect 4061 7753 4065 7757
rect 4095 7753 4099 7757
rect 4112 7753 4116 7757
rect 4168 7753 4172 7757
rect 4185 7753 4189 7757
rect 4213 7753 4217 7757
rect 2490 7745 2495 7749
rect 2623 7745 2627 7749
rect 2800 7746 2806 7750
rect 2864 7746 2868 7750
rect 3098 7746 3102 7750
rect 3284 7747 3288 7751
rect 3296 7747 3300 7751
rect 3435 7745 3440 7749
rect 3568 7745 3572 7749
rect 3745 7746 3751 7750
rect 3809 7746 3813 7750
rect 4043 7746 4047 7750
rect 4229 7747 4233 7751
rect 4241 7747 4245 7751
rect 2498 7738 2502 7742
rect 2788 7738 2794 7742
rect 3108 7739 3112 7743
rect 3273 7739 3277 7743
rect 2482 7734 2486 7738
rect 2514 7734 2518 7738
rect 2836 7732 2842 7736
rect 3443 7738 3447 7742
rect 3733 7738 3739 7742
rect 4053 7739 4057 7743
rect 4218 7739 4222 7743
rect 3427 7734 3431 7738
rect 3459 7734 3463 7738
rect 3781 7732 3787 7736
rect 2482 7725 2486 7729
rect 2514 7725 2518 7729
rect 3427 7725 3431 7729
rect 3459 7725 3463 7729
rect 2498 7718 2502 7722
rect 2755 7718 2759 7722
rect 2824 7718 2830 7722
rect 3156 7718 3160 7722
rect 3192 7718 3196 7722
rect 3259 7718 3263 7722
rect 3443 7718 3447 7722
rect 3700 7718 3704 7722
rect 3769 7718 3775 7722
rect 4101 7718 4105 7722
rect 4137 7718 4141 7722
rect 4204 7718 4208 7722
rect 2755 7710 2759 7714
rect 2764 7711 2770 7715
rect 3142 7711 3146 7715
rect 2482 7706 2486 7710
rect 2514 7706 2518 7710
rect 2498 7702 2502 7706
rect 3156 7704 3160 7708
rect 3206 7704 3210 7708
rect 3259 7704 3263 7708
rect 3700 7710 3704 7714
rect 3709 7711 3715 7715
rect 4087 7711 4091 7715
rect 3427 7706 3431 7710
rect 3459 7706 3463 7710
rect 3443 7702 3447 7706
rect 4101 7704 4105 7708
rect 4151 7704 4155 7708
rect 4204 7704 4208 7708
rect 2490 7695 2495 7699
rect 2624 7695 2628 7699
rect 3179 7693 3183 7697
rect 2373 7688 2377 7692
rect 2409 7688 2413 7692
rect 2476 7688 2480 7692
rect 2505 7688 2509 7692
rect 2541 7688 2545 7692
rect 2608 7688 2612 7692
rect 2637 7688 2641 7692
rect 2673 7688 2677 7692
rect 2740 7688 2744 7692
rect 2824 7688 2830 7692
rect 2764 7681 2770 7685
rect 3150 7684 3154 7688
rect 3163 7687 3167 7693
rect 3200 7687 3204 7693
rect 3213 7689 3217 7693
rect 3237 7693 3241 7697
rect 3435 7695 3440 7699
rect 3569 7695 3573 7699
rect 4124 7693 4128 7697
rect 3221 7687 3225 7693
rect 3258 7687 3262 7693
rect 3274 7687 3278 7693
rect 3318 7688 3322 7692
rect 3354 7688 3358 7692
rect 3421 7688 3425 7692
rect 3450 7688 3454 7692
rect 3486 7688 3490 7692
rect 3553 7688 3557 7692
rect 3582 7688 3586 7692
rect 3618 7688 3622 7692
rect 3685 7688 3689 7692
rect 3769 7688 3775 7692
rect 2373 7674 2377 7678
rect 2423 7674 2427 7678
rect 2476 7674 2480 7678
rect 2505 7674 2509 7678
rect 2555 7674 2559 7678
rect 2608 7674 2612 7678
rect 2637 7674 2641 7678
rect 2687 7674 2691 7678
rect 2740 7674 2744 7678
rect 3163 7674 3167 7678
rect 3179 7674 3183 7680
rect 3213 7680 3217 7684
rect 3200 7674 3204 7678
rect 2396 7663 2400 7667
rect 2367 7654 2371 7658
rect 2380 7657 2384 7663
rect 2417 7657 2421 7663
rect 2430 7659 2434 7663
rect 2454 7663 2458 7667
rect 2528 7663 2532 7667
rect 2438 7657 2442 7663
rect 2475 7657 2479 7663
rect 2491 7657 2495 7663
rect 2512 7657 2516 7663
rect 2549 7657 2553 7663
rect 2562 7659 2566 7663
rect 2586 7663 2590 7667
rect 2660 7663 2664 7667
rect 2570 7657 2574 7663
rect 2607 7657 2611 7663
rect 2623 7657 2627 7663
rect 2644 7657 2648 7663
rect 2681 7657 2685 7663
rect 2694 7659 2698 7663
rect 2718 7663 2722 7667
rect 2702 7657 2706 7663
rect 2739 7657 2743 7663
rect 2755 7659 2759 7663
rect 3221 7674 3225 7678
rect 3237 7674 3241 7680
rect 3709 7681 3715 7685
rect 4095 7684 4099 7688
rect 4108 7687 4112 7693
rect 4145 7687 4149 7693
rect 4158 7689 4162 7693
rect 4182 7693 4186 7697
rect 4166 7687 4170 7693
rect 4203 7687 4207 7693
rect 4219 7687 4223 7693
rect 3258 7674 3262 7678
rect 3274 7674 3278 7678
rect 3318 7674 3322 7678
rect 3368 7674 3372 7678
rect 3421 7674 3425 7678
rect 3450 7674 3454 7678
rect 3500 7674 3504 7678
rect 3553 7674 3557 7678
rect 3582 7674 3586 7678
rect 3632 7674 3636 7678
rect 3685 7674 3689 7678
rect 4108 7674 4112 7678
rect 4124 7674 4128 7680
rect 4158 7680 4162 7684
rect 4145 7674 4149 7678
rect 3156 7663 3160 7667
rect 3193 7661 3197 7665
rect 3213 7661 3217 7665
rect 3257 7661 3261 7665
rect 3341 7663 3345 7667
rect 2380 7644 2384 7648
rect 2396 7644 2400 7650
rect 2430 7650 2434 7654
rect 2417 7644 2421 7648
rect 2438 7644 2442 7648
rect 2454 7644 2458 7650
rect 2475 7644 2479 7648
rect 2491 7644 2495 7648
rect 2512 7644 2516 7648
rect 2528 7644 2532 7650
rect 2562 7650 2566 7654
rect 2549 7644 2553 7648
rect 2570 7644 2574 7648
rect 2586 7644 2590 7650
rect 2607 7644 2611 7648
rect 2623 7644 2627 7648
rect 2644 7644 2648 7648
rect 2660 7644 2664 7650
rect 2694 7650 2698 7654
rect 2681 7644 2685 7648
rect 2702 7644 2706 7648
rect 2718 7644 2722 7650
rect 2776 7654 2782 7658
rect 3312 7654 3316 7658
rect 3325 7657 3329 7663
rect 3362 7657 3366 7663
rect 3375 7659 3379 7663
rect 3399 7663 3403 7667
rect 3473 7663 3477 7667
rect 3383 7657 3387 7663
rect 3420 7657 3424 7663
rect 3436 7657 3440 7663
rect 3457 7657 3461 7663
rect 3494 7657 3498 7663
rect 3507 7659 3511 7663
rect 3531 7663 3535 7667
rect 3605 7663 3609 7667
rect 3515 7657 3519 7663
rect 3552 7657 3556 7663
rect 3568 7657 3572 7663
rect 3589 7657 3593 7663
rect 3626 7657 3630 7663
rect 3639 7659 3643 7663
rect 3663 7663 3667 7667
rect 3647 7657 3651 7663
rect 3684 7657 3688 7663
rect 3700 7659 3704 7663
rect 4166 7674 4170 7678
rect 4182 7674 4186 7680
rect 4203 7674 4207 7678
rect 4219 7674 4223 7678
rect 4101 7663 4105 7667
rect 4138 7661 4142 7665
rect 4158 7661 4162 7665
rect 4202 7661 4206 7665
rect 2739 7644 2743 7648
rect 2755 7644 2759 7648
rect 2812 7647 2818 7651
rect 3156 7647 3160 7651
rect 3207 7647 3211 7651
rect 3257 7647 3261 7651
rect 3325 7644 3329 7648
rect 3341 7644 3345 7650
rect 3375 7650 3379 7654
rect 3362 7644 3366 7648
rect 2373 7633 2377 7637
rect 2410 7631 2414 7635
rect 2430 7631 2434 7635
rect 2474 7631 2478 7635
rect 2505 7633 2509 7637
rect 2542 7631 2546 7635
rect 2562 7631 2566 7635
rect 2606 7631 2610 7635
rect 2637 7633 2641 7637
rect 2674 7631 2678 7635
rect 2694 7631 2698 7635
rect 2738 7631 2742 7635
rect 3149 7639 3153 7643
rect 3274 7640 3278 7644
rect 3383 7644 3387 7648
rect 3399 7644 3403 7650
rect 3420 7644 3424 7648
rect 3436 7644 3440 7648
rect 3457 7644 3461 7648
rect 3473 7644 3477 7650
rect 3507 7650 3511 7654
rect 3494 7644 3498 7648
rect 3515 7644 3519 7648
rect 3531 7644 3535 7650
rect 3552 7644 3556 7648
rect 3568 7644 3572 7648
rect 3589 7644 3593 7648
rect 3605 7644 3609 7650
rect 3639 7650 3643 7654
rect 3626 7644 3630 7648
rect 3647 7644 3651 7648
rect 3663 7644 3667 7650
rect 3721 7654 3727 7658
rect 3684 7644 3688 7648
rect 3700 7644 3704 7648
rect 3757 7647 3763 7651
rect 4101 7647 4105 7651
rect 4152 7647 4156 7651
rect 4202 7647 4206 7651
rect 2824 7632 2830 7636
rect 3156 7632 3160 7636
rect 3192 7632 3196 7636
rect 3259 7632 3263 7636
rect 2776 7624 2782 7628
rect 3142 7625 3146 7629
rect 3318 7633 3322 7637
rect 3355 7631 3359 7635
rect 3375 7631 3379 7635
rect 3419 7631 3423 7635
rect 3450 7633 3454 7637
rect 3487 7631 3491 7635
rect 3507 7631 3511 7635
rect 3551 7631 3555 7635
rect 3582 7633 3586 7637
rect 3619 7631 3623 7635
rect 3639 7631 3643 7635
rect 3683 7631 3687 7635
rect 4094 7639 4098 7643
rect 4219 7640 4223 7644
rect 3769 7632 3775 7636
rect 4101 7632 4105 7636
rect 4137 7632 4141 7636
rect 4204 7632 4208 7636
rect 2373 7617 2377 7621
rect 2424 7617 2428 7621
rect 2474 7617 2478 7621
rect 2505 7617 2509 7621
rect 2556 7617 2560 7621
rect 2606 7617 2610 7621
rect 2637 7617 2641 7621
rect 2688 7617 2692 7621
rect 2738 7617 2742 7621
rect 2812 7617 2818 7621
rect 3156 7618 3160 7622
rect 3206 7618 3210 7622
rect 3259 7618 3263 7622
rect 3721 7624 3727 7628
rect 4087 7625 4091 7629
rect 3318 7617 3322 7621
rect 3369 7617 3373 7621
rect 3419 7617 3423 7621
rect 3450 7617 3454 7621
rect 3501 7617 3505 7621
rect 3551 7617 3555 7621
rect 3582 7617 3586 7621
rect 3633 7617 3637 7621
rect 3683 7617 3687 7621
rect 3757 7617 3763 7621
rect 4101 7618 4105 7622
rect 4151 7618 4155 7622
rect 4204 7618 4208 7622
rect 2366 7610 2370 7614
rect 2755 7610 2759 7614
rect 3179 7607 3183 7611
rect 2373 7602 2377 7606
rect 2409 7602 2413 7606
rect 2476 7602 2480 7606
rect 2505 7602 2509 7606
rect 2541 7602 2545 7606
rect 2608 7602 2612 7606
rect 2637 7602 2641 7606
rect 2673 7602 2677 7606
rect 2740 7602 2744 7606
rect 2824 7602 2830 7606
rect 2764 7595 2770 7599
rect 3150 7598 3154 7602
rect 3163 7601 3167 7607
rect 3200 7601 3204 7607
rect 3213 7603 3217 7607
rect 3237 7607 3241 7611
rect 3311 7610 3315 7614
rect 3700 7610 3704 7614
rect 4124 7607 4128 7611
rect 3221 7601 3225 7607
rect 3258 7601 3262 7607
rect 3274 7603 3278 7607
rect 3296 7601 3300 7605
rect 3318 7602 3322 7606
rect 3354 7602 3358 7606
rect 3421 7602 3425 7606
rect 3450 7602 3454 7606
rect 3486 7602 3490 7606
rect 3553 7602 3557 7606
rect 3582 7602 3586 7606
rect 3618 7602 3622 7606
rect 3685 7602 3689 7606
rect 3769 7602 3775 7606
rect 2373 7588 2377 7592
rect 2423 7588 2427 7592
rect 2476 7588 2480 7592
rect 2505 7588 2509 7592
rect 2555 7588 2559 7592
rect 2608 7588 2612 7592
rect 2637 7588 2641 7592
rect 2687 7588 2691 7592
rect 2740 7588 2744 7592
rect 3163 7588 3167 7592
rect 3179 7588 3183 7594
rect 3213 7594 3217 7598
rect 3200 7588 3204 7592
rect 2396 7577 2400 7581
rect 2367 7568 2371 7572
rect 2380 7571 2384 7577
rect 2417 7571 2421 7577
rect 2430 7573 2434 7577
rect 2454 7577 2458 7581
rect 2528 7577 2532 7581
rect 2438 7571 2442 7577
rect 2475 7571 2479 7577
rect 2491 7571 2495 7577
rect 2512 7571 2516 7577
rect 2549 7571 2553 7577
rect 2562 7573 2566 7577
rect 2586 7577 2590 7581
rect 2660 7577 2664 7581
rect 2570 7571 2574 7577
rect 2607 7571 2611 7577
rect 2623 7571 2627 7577
rect 2644 7571 2648 7577
rect 2681 7571 2685 7577
rect 2694 7573 2698 7577
rect 2718 7577 2722 7581
rect 2702 7571 2706 7577
rect 2739 7571 2743 7577
rect 2755 7573 2759 7577
rect 3221 7588 3225 7592
rect 3237 7588 3241 7594
rect 3258 7588 3262 7592
rect 3274 7588 3278 7597
rect 3709 7595 3715 7599
rect 4095 7598 4099 7602
rect 4108 7601 4112 7607
rect 4145 7601 4149 7607
rect 4158 7603 4162 7607
rect 4182 7607 4186 7611
rect 4166 7601 4170 7607
rect 4203 7601 4207 7607
rect 4219 7603 4223 7607
rect 4241 7601 4245 7605
rect 3296 7585 3300 7589
rect 3318 7588 3322 7592
rect 3368 7588 3372 7592
rect 3421 7588 3425 7592
rect 3450 7588 3454 7592
rect 3500 7588 3504 7592
rect 3553 7588 3557 7592
rect 3582 7588 3586 7592
rect 3632 7588 3636 7592
rect 3685 7588 3689 7592
rect 4108 7588 4112 7592
rect 4124 7588 4128 7594
rect 4158 7594 4162 7598
rect 4145 7588 4149 7592
rect 3156 7577 3160 7581
rect 3193 7575 3197 7579
rect 3213 7575 3217 7579
rect 3257 7575 3261 7579
rect 3341 7577 3345 7581
rect 2380 7558 2384 7562
rect 2396 7558 2400 7564
rect 2430 7564 2434 7568
rect 2417 7558 2421 7562
rect 2438 7558 2442 7562
rect 2454 7558 2458 7564
rect 2475 7558 2479 7562
rect 2491 7558 2495 7562
rect 2512 7558 2516 7562
rect 2528 7558 2532 7564
rect 2562 7564 2566 7568
rect 2549 7558 2553 7562
rect 2570 7558 2574 7562
rect 2586 7558 2590 7564
rect 2607 7558 2611 7562
rect 2623 7558 2627 7562
rect 2644 7558 2648 7562
rect 2660 7558 2664 7564
rect 2694 7564 2698 7568
rect 2681 7558 2685 7562
rect 2702 7558 2706 7562
rect 2718 7558 2722 7564
rect 2776 7568 2782 7572
rect 3312 7568 3316 7572
rect 3325 7571 3329 7577
rect 3362 7571 3366 7577
rect 3375 7573 3379 7577
rect 3399 7577 3403 7581
rect 3473 7577 3477 7581
rect 3383 7571 3387 7577
rect 3420 7571 3424 7577
rect 3436 7571 3440 7577
rect 3457 7571 3461 7577
rect 3494 7571 3498 7577
rect 3507 7573 3511 7577
rect 3531 7577 3535 7581
rect 3605 7577 3609 7581
rect 3515 7571 3519 7577
rect 3552 7571 3556 7577
rect 3568 7571 3572 7577
rect 3589 7571 3593 7577
rect 3626 7571 3630 7577
rect 3639 7573 3643 7577
rect 3663 7577 3667 7581
rect 3647 7571 3651 7577
rect 3684 7571 3688 7577
rect 3700 7573 3704 7577
rect 4166 7588 4170 7592
rect 4182 7588 4186 7594
rect 4203 7588 4207 7592
rect 4219 7588 4223 7597
rect 4241 7585 4245 7589
rect 4101 7577 4105 7581
rect 4138 7575 4142 7579
rect 4158 7575 4162 7579
rect 4202 7575 4206 7579
rect 2739 7558 2743 7562
rect 2755 7558 2759 7562
rect 2812 7561 2818 7565
rect 3156 7561 3160 7565
rect 3207 7561 3211 7565
rect 3257 7561 3261 7565
rect 3325 7558 3329 7562
rect 3341 7558 3345 7564
rect 3375 7564 3379 7568
rect 3362 7558 3366 7562
rect 3383 7558 3387 7562
rect 3399 7558 3403 7564
rect 3420 7558 3424 7562
rect 3436 7558 3440 7562
rect 3457 7558 3461 7562
rect 3473 7558 3477 7564
rect 3507 7564 3511 7568
rect 3494 7558 3498 7562
rect 3515 7558 3519 7562
rect 3531 7558 3535 7564
rect 3552 7558 3556 7562
rect 3568 7558 3572 7562
rect 3589 7558 3593 7562
rect 3605 7558 3609 7564
rect 3639 7564 3643 7568
rect 3626 7558 3630 7562
rect 3647 7558 3651 7562
rect 3663 7558 3667 7564
rect 3721 7568 3727 7572
rect 3684 7558 3688 7562
rect 3700 7558 3704 7562
rect 3757 7561 3763 7565
rect 4101 7561 4105 7565
rect 4152 7561 4156 7565
rect 4202 7561 4206 7565
rect 2373 7547 2377 7551
rect 2410 7545 2414 7549
rect 2430 7545 2434 7549
rect 2474 7545 2478 7549
rect 2505 7547 2509 7551
rect 2542 7545 2546 7549
rect 2562 7545 2566 7549
rect 2606 7545 2610 7549
rect 2637 7547 2641 7551
rect 2674 7545 2678 7549
rect 2694 7545 2698 7549
rect 2738 7545 2742 7549
rect 3318 7547 3322 7551
rect 3355 7545 3359 7549
rect 3375 7545 3379 7549
rect 3419 7545 3423 7549
rect 3450 7547 3454 7551
rect 3487 7545 3491 7549
rect 3507 7545 3511 7549
rect 3551 7545 3555 7549
rect 3582 7547 3586 7551
rect 3619 7545 3623 7549
rect 3639 7545 3643 7549
rect 3683 7545 3687 7549
rect 2776 7538 2782 7542
rect 3721 7538 3727 7542
rect 2373 7531 2377 7535
rect 2424 7531 2428 7535
rect 2474 7531 2478 7535
rect 2505 7531 2509 7535
rect 2556 7531 2560 7535
rect 2606 7531 2610 7535
rect 2637 7531 2641 7535
rect 2688 7531 2692 7535
rect 2738 7531 2742 7535
rect 2812 7531 2818 7535
rect 3318 7531 3322 7535
rect 3369 7531 3373 7535
rect 3419 7531 3423 7535
rect 3450 7531 3454 7535
rect 3501 7531 3505 7535
rect 3551 7531 3555 7535
rect 3582 7531 3586 7535
rect 3633 7531 3637 7535
rect 3683 7531 3687 7535
rect 3757 7531 3763 7535
rect 2366 7524 2370 7528
rect 2755 7524 2759 7528
rect 3311 7524 3315 7528
rect 3700 7524 3704 7528
rect 2491 7517 2495 7521
rect 2599 7517 2603 7521
rect 2623 7517 2627 7521
rect 3436 7517 3440 7521
rect 3544 7517 3548 7521
rect 3568 7517 3572 7521
rect 2615 7510 2619 7514
rect 2599 7506 2603 7510
rect 2631 7506 2635 7510
rect 3560 7510 3564 7514
rect 3544 7506 3548 7510
rect 3576 7506 3580 7510
rect 2599 7499 2603 7503
rect 2631 7499 2635 7503
rect 3296 7499 3300 7503
rect 3544 7499 3548 7503
rect 3576 7499 3580 7503
rect 3836 7499 3844 7503
rect 4241 7499 4245 7503
rect 4360 7499 4369 7503
rect 2615 7492 2619 7496
rect 2755 7492 2759 7496
rect 3560 7492 3564 7496
rect 3700 7492 3704 7496
rect 4529 7494 4533 7498
rect 4534 7494 4538 7498
rect 4539 7494 4543 7498
rect 4544 7494 4548 7498
rect 4549 7494 4553 7498
rect 4554 7494 4558 7498
rect 4559 7494 4563 7498
rect 4564 7494 4568 7498
rect 4569 7494 4573 7498
rect 4574 7494 4578 7498
rect 4579 7494 4583 7498
rect 4584 7494 4588 7498
rect 4589 7494 4593 7498
rect 4529 7489 4533 7493
rect 4534 7489 4538 7493
rect 4539 7489 4543 7493
rect 4544 7489 4548 7493
rect 4549 7489 4553 7493
rect 4554 7489 4558 7493
rect 4559 7489 4563 7493
rect 4564 7489 4568 7493
rect 4569 7489 4573 7493
rect 4574 7489 4578 7493
rect 4579 7489 4583 7493
rect 4584 7489 4588 7493
rect 4589 7489 4593 7493
rect 2755 7484 2759 7488
rect 3700 7484 3704 7488
rect 2599 7480 2603 7484
rect 2631 7480 2635 7484
rect 2615 7476 2619 7480
rect 3544 7480 3548 7484
rect 3576 7480 3580 7484
rect 3560 7476 3564 7480
rect 3836 7480 3844 7484
rect 618 7467 622 7471
rect 628 7467 632 7471
rect 638 7467 642 7471
rect 618 7462 622 7466
rect 628 7462 632 7466
rect 638 7462 642 7466
rect 618 7457 622 7461
rect 628 7457 632 7461
rect 638 7457 642 7461
rect 618 7452 622 7456
rect 628 7452 632 7456
rect 638 7452 642 7456
rect 664 7467 668 7471
rect 674 7467 678 7471
rect 684 7467 688 7471
rect 2491 7469 2495 7473
rect 2599 7469 2603 7473
rect 2623 7469 2627 7473
rect 3436 7469 3440 7473
rect 3544 7469 3548 7473
rect 3568 7469 3572 7473
rect 3918 7472 3922 7476
rect 664 7462 668 7466
rect 674 7462 678 7466
rect 684 7462 688 7466
rect 2373 7462 2377 7466
rect 2409 7462 2413 7466
rect 2476 7462 2480 7466
rect 2505 7462 2509 7466
rect 2541 7462 2545 7466
rect 2608 7462 2612 7466
rect 2637 7462 2641 7466
rect 2673 7462 2677 7466
rect 2740 7462 2744 7466
rect 2824 7462 2830 7466
rect 3318 7462 3322 7466
rect 3354 7462 3358 7466
rect 3421 7462 3425 7466
rect 3450 7462 3454 7466
rect 3486 7462 3490 7466
rect 3553 7462 3557 7466
rect 3582 7462 3586 7466
rect 3618 7462 3622 7466
rect 3685 7462 3689 7466
rect 3769 7462 3775 7466
rect 3836 7464 3844 7468
rect 664 7457 668 7461
rect 674 7457 678 7461
rect 684 7457 688 7461
rect 664 7452 668 7456
rect 674 7452 678 7456
rect 684 7452 688 7456
rect 2764 7455 2770 7459
rect 3709 7455 3715 7459
rect 2373 7448 2377 7452
rect 2423 7448 2427 7452
rect 2476 7448 2480 7452
rect 2505 7448 2509 7452
rect 2555 7448 2559 7452
rect 2608 7448 2612 7452
rect 2637 7448 2641 7452
rect 2687 7448 2691 7452
rect 2740 7448 2744 7452
rect 3318 7448 3322 7452
rect 3368 7448 3372 7452
rect 3421 7448 3425 7452
rect 3450 7448 3454 7452
rect 3500 7448 3504 7452
rect 3553 7448 3557 7452
rect 3582 7448 3586 7452
rect 3632 7448 3636 7452
rect 3685 7448 3689 7452
rect 2396 7437 2400 7441
rect 2367 7428 2371 7432
rect 2380 7431 2384 7437
rect 2417 7431 2421 7437
rect 2430 7433 2434 7437
rect 2454 7437 2458 7441
rect 2528 7437 2532 7441
rect 2438 7431 2442 7437
rect 2475 7431 2479 7437
rect 2491 7431 2495 7437
rect 2512 7431 2516 7437
rect 2549 7431 2553 7437
rect 2562 7433 2566 7437
rect 2586 7437 2590 7441
rect 2660 7437 2664 7441
rect 2570 7431 2574 7437
rect 2607 7431 2611 7437
rect 2623 7431 2627 7437
rect 2644 7431 2648 7437
rect 2681 7431 2685 7437
rect 2694 7433 2698 7437
rect 2718 7437 2722 7441
rect 3341 7437 3345 7441
rect 2702 7431 2706 7437
rect 2739 7431 2743 7437
rect 2755 7433 2759 7437
rect 2380 7418 2384 7422
rect 2396 7418 2400 7424
rect 2430 7424 2434 7428
rect 2417 7418 2421 7422
rect 2438 7418 2442 7422
rect 2454 7418 2458 7424
rect 2475 7418 2479 7422
rect 2491 7418 2495 7422
rect 2512 7418 2516 7422
rect 2528 7418 2532 7424
rect 2562 7424 2566 7428
rect 2549 7418 2553 7422
rect 2570 7418 2574 7422
rect 2586 7418 2590 7424
rect 2607 7418 2611 7422
rect 2623 7418 2627 7422
rect 2644 7418 2648 7422
rect 2660 7418 2664 7424
rect 2694 7424 2698 7428
rect 2681 7418 2685 7422
rect 2702 7418 2706 7422
rect 2718 7418 2722 7424
rect 3312 7428 3316 7432
rect 3325 7431 3329 7437
rect 3362 7431 3366 7437
rect 3375 7433 3379 7437
rect 3399 7437 3403 7441
rect 3473 7437 3477 7441
rect 3383 7431 3387 7437
rect 3420 7431 3424 7437
rect 3436 7431 3440 7437
rect 3457 7431 3461 7437
rect 3494 7431 3498 7437
rect 3507 7433 3511 7437
rect 3531 7437 3535 7441
rect 3605 7437 3609 7441
rect 3515 7431 3519 7437
rect 3552 7431 3556 7437
rect 3568 7431 3572 7437
rect 3589 7431 3593 7437
rect 3626 7431 3630 7437
rect 3639 7433 3643 7437
rect 3663 7437 3667 7441
rect 3647 7431 3651 7437
rect 3684 7431 3688 7437
rect 3700 7433 3704 7437
rect 2739 7418 2743 7422
rect 2755 7418 2759 7422
rect 3325 7418 3329 7422
rect 3341 7418 3345 7424
rect 3375 7424 3379 7428
rect 3362 7418 3366 7422
rect 3383 7418 3387 7422
rect 3399 7418 3403 7424
rect 3420 7418 3424 7422
rect 3436 7418 3440 7422
rect 3457 7418 3461 7422
rect 3473 7418 3477 7424
rect 3507 7424 3511 7428
rect 3494 7418 3498 7422
rect 3515 7418 3519 7422
rect 3531 7418 3535 7424
rect 3552 7418 3556 7422
rect 3568 7418 3572 7422
rect 3589 7418 3593 7422
rect 3605 7418 3609 7424
rect 3639 7424 3643 7428
rect 3626 7418 3630 7422
rect 3647 7418 3651 7422
rect 3663 7418 3667 7424
rect 3684 7418 3688 7422
rect 3700 7418 3704 7422
rect 2373 7407 2377 7411
rect 2410 7405 2414 7409
rect 2430 7405 2434 7409
rect 2474 7405 2478 7409
rect 2505 7407 2509 7411
rect 2542 7405 2546 7409
rect 2562 7405 2566 7409
rect 2606 7405 2610 7409
rect 2637 7407 2641 7411
rect 2674 7405 2678 7409
rect 2694 7405 2698 7409
rect 2738 7405 2742 7409
rect 3318 7407 3322 7411
rect 3355 7405 3359 7409
rect 3375 7405 3379 7409
rect 3419 7405 3423 7409
rect 3450 7407 3454 7411
rect 3487 7405 3491 7409
rect 3507 7405 3511 7409
rect 3551 7405 3555 7409
rect 3582 7407 3586 7411
rect 3619 7405 3623 7409
rect 3639 7405 3643 7409
rect 3683 7405 3687 7409
rect 2776 7398 2782 7402
rect 3721 7398 3727 7402
rect 2373 7391 2377 7395
rect 2424 7391 2428 7395
rect 2474 7391 2478 7395
rect 2505 7391 2509 7395
rect 2556 7391 2560 7395
rect 2606 7391 2610 7395
rect 2637 7391 2641 7395
rect 2688 7391 2692 7395
rect 2738 7391 2742 7395
rect 2812 7391 2818 7395
rect 3318 7391 3322 7395
rect 3369 7391 3373 7395
rect 3419 7391 3423 7395
rect 3450 7391 3454 7395
rect 3501 7391 3505 7395
rect 3551 7391 3555 7395
rect 3582 7391 3586 7395
rect 3633 7391 3637 7395
rect 3683 7391 3687 7395
rect 3757 7391 3763 7395
rect 4572 7389 4576 7393
rect 4588 7389 4592 7393
rect 4604 7389 4608 7393
rect 4641 7473 4645 7477
rect 4641 7466 4645 7470
rect 4641 7461 4645 7465
rect 4641 7456 4645 7460
rect 4641 7451 4645 7455
rect 4641 7446 4645 7450
rect 4641 7441 4645 7445
rect 4641 7436 4645 7440
rect 4641 7431 4645 7435
rect 4641 7426 4645 7430
rect 4641 7421 4645 7425
rect 4662 7461 4666 7465
rect 4672 7461 4676 7465
rect 4682 7461 4686 7465
rect 4692 7461 4696 7465
rect 4702 7461 4706 7465
rect 4712 7461 4716 7465
rect 4722 7461 4726 7465
rect 4732 7461 4736 7465
rect 4742 7461 4746 7465
rect 4657 7456 4661 7460
rect 4667 7456 4671 7460
rect 4677 7456 4681 7460
rect 4687 7456 4691 7460
rect 4697 7456 4701 7460
rect 4707 7456 4711 7460
rect 4717 7456 4721 7460
rect 4727 7456 4731 7460
rect 4737 7456 4741 7460
rect 4662 7451 4666 7455
rect 4672 7451 4676 7455
rect 4682 7451 4686 7455
rect 4692 7451 4696 7455
rect 4702 7451 4706 7455
rect 4712 7451 4716 7455
rect 4722 7451 4726 7455
rect 4732 7451 4736 7455
rect 4742 7451 4746 7455
rect 4657 7446 4661 7450
rect 4667 7446 4671 7450
rect 4677 7446 4681 7450
rect 4687 7446 4691 7450
rect 4697 7446 4701 7450
rect 4707 7446 4711 7450
rect 4717 7446 4721 7450
rect 4727 7446 4731 7450
rect 4737 7446 4741 7450
rect 4662 7441 4666 7445
rect 4672 7441 4676 7445
rect 4682 7441 4686 7445
rect 4692 7441 4696 7445
rect 4702 7441 4706 7445
rect 4712 7441 4716 7445
rect 4722 7441 4726 7445
rect 4732 7441 4736 7445
rect 4742 7441 4746 7445
rect 4657 7436 4661 7440
rect 4667 7436 4671 7440
rect 4677 7436 4681 7440
rect 4687 7436 4691 7440
rect 4697 7436 4701 7440
rect 4707 7436 4711 7440
rect 4717 7436 4721 7440
rect 4727 7436 4731 7440
rect 4737 7436 4741 7440
rect 4662 7431 4666 7435
rect 4672 7431 4676 7435
rect 4682 7431 4686 7435
rect 4692 7431 4696 7435
rect 4702 7431 4706 7435
rect 4712 7431 4716 7435
rect 4722 7431 4726 7435
rect 4732 7431 4736 7435
rect 4742 7431 4746 7435
rect 4657 7426 4661 7430
rect 4667 7426 4671 7430
rect 4677 7426 4681 7430
rect 4687 7426 4691 7430
rect 4697 7426 4701 7430
rect 4707 7426 4711 7430
rect 4717 7426 4721 7430
rect 4727 7426 4731 7430
rect 4737 7426 4741 7430
rect 4662 7421 4666 7425
rect 4672 7421 4676 7425
rect 4682 7421 4686 7425
rect 4692 7421 4696 7425
rect 4702 7421 4706 7425
rect 4712 7421 4716 7425
rect 4722 7421 4726 7425
rect 4732 7421 4736 7425
rect 4742 7421 4746 7425
rect 4641 7416 4645 7420
rect 4641 7409 4645 7413
rect 4775 7404 4779 7408
rect 4780 7404 4784 7408
rect 4785 7404 4789 7408
rect 4790 7404 4794 7408
rect 4775 7397 4779 7401
rect 4780 7397 4784 7401
rect 4785 7397 4789 7401
rect 4790 7397 4794 7401
rect 4620 7389 4624 7393
rect 4775 7390 4779 7394
rect 4780 7390 4784 7394
rect 4785 7390 4789 7394
rect 4790 7390 4794 7394
rect 4775 7383 4779 7387
rect 4780 7383 4784 7387
rect 4785 7383 4789 7387
rect 4790 7383 4794 7387
rect 4775 7376 4779 7380
rect 4780 7376 4784 7380
rect 4785 7376 4789 7380
rect 4790 7376 4794 7380
rect 3918 7362 3922 7366
rect 4775 7369 4779 7373
rect 4780 7369 4784 7373
rect 4785 7369 4789 7373
rect 4790 7369 4794 7373
rect 4775 7362 4779 7366
rect 4780 7362 4784 7366
rect 4785 7362 4789 7366
rect 4790 7362 4794 7366
rect 4775 7355 4779 7359
rect 4780 7355 4784 7359
rect 4785 7355 4789 7359
rect 4790 7355 4794 7359
rect 4775 7348 4779 7352
rect 4780 7348 4784 7352
rect 4785 7348 4789 7352
rect 4790 7348 4794 7352
rect 4572 7331 4576 7335
rect 4588 7331 4592 7335
rect 4604 7331 4608 7335
rect 4620 7331 4624 7335
rect 4775 7341 4779 7345
rect 4780 7341 4784 7345
rect 4785 7341 4789 7345
rect 4790 7341 4794 7345
rect 4775 7334 4779 7338
rect 4780 7334 4784 7338
rect 4785 7334 4789 7338
rect 4790 7334 4794 7338
rect 4506 7289 4510 7293
rect 4511 7289 4515 7293
rect 4506 7284 4510 7288
rect 4511 7284 4515 7288
rect 4506 7279 4510 7283
rect 4511 7279 4515 7283
rect 4506 7274 4510 7278
rect 4511 7274 4515 7278
rect 4506 7269 4510 7273
rect 4511 7269 4515 7273
rect 4506 7264 4510 7268
rect 4511 7264 4515 7268
rect 4506 7259 4510 7263
rect 4511 7259 4515 7263
rect 4506 7254 4510 7258
rect 4511 7254 4515 7258
rect 4506 7249 4510 7253
rect 4511 7249 4515 7253
rect 4506 7244 4510 7248
rect 4511 7244 4515 7248
rect 4641 7313 4645 7317
rect 4641 7306 4645 7310
rect 4641 7301 4645 7305
rect 4641 7296 4645 7300
rect 4641 7291 4645 7295
rect 4641 7286 4645 7290
rect 4641 7281 4645 7285
rect 4641 7276 4645 7280
rect 4641 7271 4645 7275
rect 4641 7266 4645 7270
rect 4641 7261 4645 7265
rect 4662 7301 4666 7305
rect 4672 7301 4676 7305
rect 4682 7301 4686 7305
rect 4692 7301 4696 7305
rect 4702 7301 4706 7305
rect 4712 7301 4716 7305
rect 4722 7301 4726 7305
rect 4732 7301 4736 7305
rect 4742 7301 4746 7305
rect 4657 7296 4661 7300
rect 4667 7296 4671 7300
rect 4677 7296 4681 7300
rect 4687 7296 4691 7300
rect 4697 7296 4701 7300
rect 4707 7296 4711 7300
rect 4717 7296 4721 7300
rect 4727 7296 4731 7300
rect 4737 7296 4741 7300
rect 4662 7291 4666 7295
rect 4672 7291 4676 7295
rect 4682 7291 4686 7295
rect 4692 7291 4696 7295
rect 4702 7291 4706 7295
rect 4712 7291 4716 7295
rect 4722 7291 4726 7295
rect 4732 7291 4736 7295
rect 4742 7291 4746 7295
rect 4657 7286 4661 7290
rect 4667 7286 4671 7290
rect 4677 7286 4681 7290
rect 4687 7286 4691 7290
rect 4697 7286 4701 7290
rect 4707 7286 4711 7290
rect 4717 7286 4721 7290
rect 4727 7286 4731 7290
rect 4737 7286 4741 7290
rect 4662 7281 4666 7285
rect 4672 7281 4676 7285
rect 4682 7281 4686 7285
rect 4692 7281 4696 7285
rect 4702 7281 4706 7285
rect 4712 7281 4716 7285
rect 4722 7281 4726 7285
rect 4732 7281 4736 7285
rect 4742 7281 4746 7285
rect 4657 7276 4661 7280
rect 4667 7276 4671 7280
rect 4677 7276 4681 7280
rect 4687 7276 4691 7280
rect 4697 7276 4701 7280
rect 4707 7276 4711 7280
rect 4717 7276 4721 7280
rect 4727 7276 4731 7280
rect 4737 7276 4741 7280
rect 4662 7271 4666 7275
rect 4672 7271 4676 7275
rect 4682 7271 4686 7275
rect 4692 7271 4696 7275
rect 4702 7271 4706 7275
rect 4712 7271 4716 7275
rect 4722 7271 4726 7275
rect 4732 7271 4736 7275
rect 4742 7271 4746 7275
rect 4657 7266 4661 7270
rect 4667 7266 4671 7270
rect 4677 7266 4681 7270
rect 4687 7266 4691 7270
rect 4697 7266 4701 7270
rect 4707 7266 4711 7270
rect 4717 7266 4721 7270
rect 4727 7266 4731 7270
rect 4737 7266 4741 7270
rect 4662 7261 4666 7265
rect 4672 7261 4676 7265
rect 4682 7261 4686 7265
rect 4692 7261 4696 7265
rect 4702 7261 4706 7265
rect 4712 7261 4716 7265
rect 4722 7261 4726 7265
rect 4732 7261 4736 7265
rect 4742 7261 4746 7265
rect 4641 7256 4645 7260
rect 4641 7249 4645 7253
rect 4775 7327 4779 7331
rect 4780 7327 4784 7331
rect 4785 7327 4789 7331
rect 4790 7327 4794 7331
rect 4775 7320 4779 7324
rect 4780 7320 4784 7324
rect 4785 7320 4789 7324
rect 4790 7320 4794 7324
rect 4506 7239 4510 7243
rect 4511 7239 4515 7243
rect 4484 7230 4488 7234
rect 4494 7230 4498 7234
rect 4504 7230 4508 7234
rect 4484 7225 4488 7229
rect 4494 7225 4498 7229
rect 4504 7225 4508 7229
rect 4484 7220 4488 7224
rect 4494 7220 4498 7224
rect 4504 7220 4508 7224
rect 4484 7215 4488 7219
rect 4494 7215 4498 7219
rect 4504 7215 4508 7219
rect 4530 7230 4534 7234
rect 4540 7230 4544 7234
rect 4550 7230 4554 7234
rect 4530 7225 4534 7229
rect 4540 7225 4544 7229
rect 4550 7225 4554 7229
rect 4530 7220 4534 7224
rect 4540 7220 4544 7224
rect 4550 7220 4554 7224
rect 4530 7215 4534 7219
rect 4540 7215 4544 7219
rect 4550 7215 4554 7219
rect 4484 7202 4488 7206
rect 4494 7202 4498 7206
rect 4504 7202 4508 7206
rect 4484 7197 4488 7201
rect 4494 7197 4498 7201
rect 4504 7197 4508 7201
rect 4484 7192 4488 7196
rect 4494 7192 4498 7196
rect 4504 7192 4508 7196
rect 4484 7187 4488 7191
rect 4494 7187 4498 7191
rect 4504 7187 4508 7191
rect 4530 7202 4534 7206
rect 4540 7202 4544 7206
rect 4550 7202 4554 7206
rect 4530 7197 4534 7201
rect 4540 7197 4544 7201
rect 4550 7197 4554 7201
rect 4530 7192 4534 7196
rect 4540 7192 4544 7196
rect 4550 7192 4554 7196
rect 4530 7187 4534 7191
rect 4540 7187 4544 7191
rect 4550 7187 4554 7191
rect 618 7158 622 7162
rect 628 7158 632 7162
rect 638 7158 642 7162
rect 664 7158 668 7162
rect 674 7158 678 7162
rect 684 7158 688 7162
rect 4484 7152 4488 7156
rect 4494 7152 4498 7156
rect 4504 7152 4508 7156
rect 4530 7152 4534 7156
rect 4540 7152 4544 7156
rect 4550 7152 4554 7156
rect 618 7123 622 7127
rect 628 7123 632 7127
rect 638 7123 642 7127
rect 618 7118 622 7122
rect 628 7118 632 7122
rect 638 7118 642 7122
rect 618 7113 622 7117
rect 628 7113 632 7117
rect 638 7113 642 7117
rect 618 7108 622 7112
rect 628 7108 632 7112
rect 638 7108 642 7112
rect 664 7123 668 7127
rect 674 7123 678 7127
rect 684 7123 688 7127
rect 664 7118 668 7122
rect 674 7118 678 7122
rect 684 7118 688 7122
rect 664 7113 668 7117
rect 674 7113 678 7117
rect 684 7113 688 7117
rect 664 7108 668 7112
rect 674 7108 678 7112
rect 684 7108 688 7112
rect 1409 6919 1415 6923
rect 1485 6919 1489 6923
rect 1535 6919 1539 6923
rect 1586 6919 1590 6923
rect 1617 6919 1621 6923
rect 1667 6919 1671 6923
rect 1718 6919 1722 6923
rect 1749 6919 1753 6923
rect 1799 6919 1803 6923
rect 1850 6919 1854 6923
rect 2354 6919 2360 6923
rect 2430 6919 2434 6923
rect 2480 6919 2484 6923
rect 2531 6919 2535 6923
rect 2562 6919 2566 6923
rect 2612 6919 2616 6923
rect 2663 6919 2667 6923
rect 2694 6919 2698 6923
rect 2744 6919 2748 6923
rect 2795 6919 2799 6923
rect 1445 6912 1451 6916
rect 2390 6912 2396 6916
rect 1485 6905 1489 6909
rect 1529 6905 1533 6909
rect 1549 6905 1553 6909
rect 1586 6903 1590 6907
rect 1617 6905 1621 6909
rect 1661 6905 1665 6909
rect 1681 6905 1685 6909
rect 1718 6903 1722 6907
rect 1749 6905 1753 6909
rect 1793 6905 1797 6909
rect 1813 6905 1817 6909
rect 1850 6903 1854 6907
rect 2430 6905 2434 6909
rect 2474 6905 2478 6909
rect 2494 6905 2498 6909
rect 2531 6903 2535 6907
rect 2562 6905 2566 6909
rect 2606 6905 2610 6909
rect 2626 6905 2630 6909
rect 2663 6903 2667 6907
rect 2694 6905 2698 6909
rect 2738 6905 2742 6909
rect 2758 6905 2762 6909
rect 2795 6903 2799 6907
rect 1468 6892 1472 6896
rect 1484 6892 1488 6896
rect 1505 6890 1509 6896
rect 1521 6892 1525 6896
rect 1542 6892 1546 6896
rect 1529 6886 1533 6890
rect 1563 6890 1567 6896
rect 1579 6892 1583 6896
rect 1600 6892 1604 6896
rect 1616 6892 1620 6896
rect 1637 6890 1641 6896
rect 1653 6892 1657 6896
rect 1674 6892 1678 6896
rect 1661 6886 1665 6890
rect 1695 6890 1699 6896
rect 1711 6892 1715 6896
rect 1732 6892 1736 6896
rect 1748 6892 1752 6896
rect 1769 6890 1773 6896
rect 1785 6892 1789 6896
rect 1806 6892 1810 6896
rect 1793 6886 1797 6890
rect 1827 6890 1831 6896
rect 1843 6892 1847 6896
rect 2413 6892 2417 6896
rect 2429 6892 2433 6896
rect 1468 6877 1472 6881
rect 1484 6877 1488 6883
rect 1521 6877 1525 6883
rect 1505 6873 1509 6877
rect 1529 6877 1533 6881
rect 1542 6877 1546 6883
rect 1579 6877 1583 6883
rect 1600 6877 1604 6883
rect 1616 6877 1620 6883
rect 1653 6877 1657 6883
rect 1563 6873 1567 6877
rect 1637 6873 1641 6877
rect 1661 6877 1665 6881
rect 1674 6877 1678 6883
rect 1711 6877 1715 6883
rect 1732 6877 1736 6883
rect 1748 6877 1752 6883
rect 1785 6877 1789 6883
rect 1695 6873 1699 6877
rect 1769 6873 1773 6877
rect 1793 6877 1797 6881
rect 1806 6877 1810 6883
rect 1843 6877 1847 6883
rect 1856 6882 1860 6886
rect 2450 6890 2454 6896
rect 2466 6892 2470 6896
rect 2487 6892 2491 6896
rect 2474 6886 2478 6890
rect 2508 6890 2512 6896
rect 2524 6892 2528 6896
rect 2545 6892 2549 6896
rect 2561 6892 2565 6896
rect 2582 6890 2586 6896
rect 2598 6892 2602 6896
rect 2619 6892 2623 6896
rect 2606 6886 2610 6890
rect 2640 6890 2644 6896
rect 2656 6892 2660 6896
rect 2677 6892 2681 6896
rect 2693 6892 2697 6896
rect 2714 6890 2718 6896
rect 2730 6892 2734 6896
rect 2751 6892 2755 6896
rect 2738 6886 2742 6890
rect 2772 6890 2776 6896
rect 2788 6892 2792 6896
rect 2413 6877 2417 6881
rect 2429 6877 2433 6883
rect 2466 6877 2470 6883
rect 1827 6873 1831 6877
rect 2450 6873 2454 6877
rect 2474 6877 2478 6881
rect 2487 6877 2491 6883
rect 2524 6877 2528 6883
rect 2545 6877 2549 6883
rect 2561 6877 2565 6883
rect 2598 6877 2602 6883
rect 2508 6873 2512 6877
rect 2582 6873 2586 6877
rect 2606 6877 2610 6881
rect 2619 6877 2623 6883
rect 2656 6877 2660 6883
rect 2677 6877 2681 6883
rect 2693 6877 2697 6883
rect 2730 6877 2734 6883
rect 2640 6873 2644 6877
rect 2714 6873 2718 6877
rect 2738 6877 2742 6881
rect 2751 6877 2755 6883
rect 2788 6877 2792 6883
rect 2801 6882 2805 6886
rect 2772 6873 2776 6877
rect 1483 6862 1487 6866
rect 1536 6862 1540 6866
rect 1586 6862 1590 6866
rect 1615 6862 1619 6866
rect 1668 6862 1672 6866
rect 1718 6862 1722 6866
rect 1747 6862 1751 6866
rect 1800 6862 1804 6866
rect 1850 6862 1854 6866
rect 2428 6862 2432 6866
rect 2481 6862 2485 6866
rect 2531 6862 2535 6866
rect 2560 6862 2564 6866
rect 2613 6862 2617 6866
rect 2663 6862 2667 6866
rect 2692 6862 2696 6866
rect 2745 6862 2749 6866
rect 2795 6862 2799 6866
rect 1457 6855 1463 6859
rect 2402 6855 2408 6859
rect 4484 6858 4488 6862
rect 4494 6858 4498 6862
rect 4504 6858 4508 6862
rect 4484 6853 4488 6857
rect 4494 6853 4498 6857
rect 4504 6853 4508 6857
rect 1397 6848 1403 6852
rect 1483 6848 1487 6852
rect 1550 6848 1554 6852
rect 1586 6848 1590 6852
rect 1615 6848 1619 6852
rect 1682 6848 1686 6852
rect 1718 6848 1722 6852
rect 1747 6848 1751 6852
rect 1814 6848 1818 6852
rect 1850 6848 1854 6852
rect 2342 6848 2348 6852
rect 2428 6848 2432 6852
rect 2495 6848 2499 6852
rect 2531 6848 2535 6852
rect 2560 6848 2564 6852
rect 2627 6848 2631 6852
rect 2663 6848 2667 6852
rect 2692 6848 2696 6852
rect 2759 6848 2763 6852
rect 2795 6848 2799 6852
rect 4484 6848 4488 6852
rect 4494 6848 4498 6852
rect 4504 6848 4508 6852
rect 1600 6841 1604 6845
rect 1624 6841 1628 6845
rect 1732 6841 1736 6845
rect 2545 6841 2549 6845
rect 2569 6841 2573 6845
rect 2677 6841 2681 6845
rect 4484 6843 4488 6847
rect 4494 6843 4498 6847
rect 4504 6843 4508 6847
rect 4530 6858 4534 6862
rect 4540 6858 4544 6862
rect 4550 6858 4554 6862
rect 4530 6853 4534 6857
rect 4540 6853 4544 6857
rect 4550 6853 4554 6857
rect 4530 6848 4534 6852
rect 4540 6848 4544 6852
rect 4550 6848 4554 6852
rect 4530 6843 4534 6847
rect 4540 6843 4544 6847
rect 4550 6843 4554 6847
rect 1608 6834 1612 6838
rect 1592 6830 1596 6834
rect 1624 6830 1628 6834
rect 2553 6834 2557 6838
rect 2537 6830 2541 6834
rect 2569 6830 2573 6834
rect 1468 6826 1472 6830
rect 2413 6826 2417 6830
rect 1468 6818 1472 6822
rect 1608 6818 1612 6822
rect 2413 6818 2417 6822
rect 2553 6818 2557 6822
rect 803 6811 812 6815
rect 927 6811 931 6815
rect 1592 6811 1596 6815
rect 1624 6811 1628 6815
rect 1872 6811 1876 6815
rect 2537 6811 2541 6815
rect 2569 6811 2573 6815
rect 1592 6804 1596 6808
rect 1624 6804 1628 6808
rect 1608 6800 1612 6804
rect 2537 6804 2541 6808
rect 2569 6804 2573 6808
rect 2553 6800 2557 6804
rect 1600 6793 1604 6797
rect 1624 6793 1628 6797
rect 1732 6793 1736 6797
rect 2545 6793 2549 6797
rect 2569 6793 2573 6797
rect 2677 6793 2681 6797
rect 1468 6786 1472 6790
rect 1857 6786 1861 6790
rect 2413 6786 2417 6790
rect 2802 6786 2806 6790
rect 1409 6779 1415 6783
rect 1485 6779 1489 6783
rect 1535 6779 1539 6783
rect 1586 6779 1590 6783
rect 1617 6779 1621 6783
rect 1667 6779 1671 6783
rect 1718 6779 1722 6783
rect 1749 6779 1753 6783
rect 1799 6779 1803 6783
rect 1850 6779 1854 6783
rect 2354 6779 2360 6783
rect 2430 6779 2434 6783
rect 2480 6779 2484 6783
rect 2531 6779 2535 6783
rect 2562 6779 2566 6783
rect 2612 6779 2616 6783
rect 2663 6779 2667 6783
rect 2694 6779 2698 6783
rect 2744 6779 2748 6783
rect 2795 6779 2799 6783
rect 1445 6772 1451 6776
rect 2390 6772 2396 6776
rect 1485 6765 1489 6769
rect 1529 6765 1533 6769
rect 1549 6765 1553 6769
rect 1586 6763 1590 6767
rect 1617 6765 1621 6769
rect 1661 6765 1665 6769
rect 1681 6765 1685 6769
rect 1718 6763 1722 6767
rect 1749 6765 1753 6769
rect 1793 6765 1797 6769
rect 1813 6765 1817 6769
rect 1850 6763 1854 6767
rect 2430 6765 2434 6769
rect 2474 6765 2478 6769
rect 2494 6765 2498 6769
rect 2531 6763 2535 6767
rect 2562 6765 2566 6769
rect 2606 6765 2610 6769
rect 2626 6765 2630 6769
rect 2663 6763 2667 6767
rect 2694 6765 2698 6769
rect 2738 6765 2742 6769
rect 2758 6765 2762 6769
rect 2795 6763 2799 6767
rect 966 6749 970 6753
rect 1016 6749 1020 6753
rect 1067 6749 1071 6753
rect 1409 6749 1415 6753
rect 1468 6752 1472 6756
rect 1484 6752 1488 6756
rect 1445 6742 1451 6746
rect 1505 6750 1509 6756
rect 1521 6752 1525 6756
rect 1542 6752 1546 6756
rect 1529 6746 1533 6750
rect 1563 6750 1567 6756
rect 1579 6752 1583 6756
rect 1600 6752 1604 6756
rect 1616 6752 1620 6756
rect 1637 6750 1641 6756
rect 1653 6752 1657 6756
rect 1674 6752 1678 6756
rect 1661 6746 1665 6750
rect 1695 6750 1699 6756
rect 1711 6752 1715 6756
rect 1732 6752 1736 6756
rect 1748 6752 1752 6756
rect 1769 6750 1773 6756
rect 1785 6752 1789 6756
rect 1806 6752 1810 6756
rect 1793 6746 1797 6750
rect 1827 6750 1831 6756
rect 1843 6752 1847 6756
rect 1911 6749 1915 6753
rect 1961 6749 1965 6753
rect 2012 6749 2016 6753
rect 2354 6749 2360 6753
rect 2413 6752 2417 6756
rect 2429 6752 2433 6756
rect 966 6735 970 6739
rect 1010 6735 1014 6739
rect 1030 6735 1034 6739
rect 1067 6733 1071 6737
rect 927 6725 931 6729
rect 949 6717 953 6726
rect 965 6722 969 6726
rect 986 6720 990 6726
rect 1002 6722 1006 6726
rect 1468 6737 1472 6741
rect 1484 6737 1488 6743
rect 1521 6737 1525 6743
rect 1505 6733 1509 6737
rect 1529 6737 1533 6741
rect 1542 6737 1546 6743
rect 1579 6737 1583 6743
rect 1600 6737 1604 6743
rect 1616 6737 1620 6743
rect 1653 6737 1657 6743
rect 1563 6733 1567 6737
rect 1637 6733 1641 6737
rect 1661 6737 1665 6741
rect 1674 6737 1678 6743
rect 1711 6737 1715 6743
rect 1732 6737 1736 6743
rect 1748 6737 1752 6743
rect 1785 6737 1789 6743
rect 1695 6733 1699 6737
rect 1769 6733 1773 6737
rect 1793 6737 1797 6741
rect 1806 6737 1810 6743
rect 1843 6737 1847 6743
rect 1856 6742 1860 6746
rect 2390 6742 2396 6746
rect 2450 6750 2454 6756
rect 2466 6752 2470 6756
rect 2487 6752 2491 6756
rect 2474 6746 2478 6750
rect 2508 6750 2512 6756
rect 2524 6752 2528 6756
rect 2545 6752 2549 6756
rect 2561 6752 2565 6756
rect 2582 6750 2586 6756
rect 2598 6752 2602 6756
rect 2619 6752 2623 6756
rect 2606 6746 2610 6750
rect 2640 6750 2644 6756
rect 2656 6752 2660 6756
rect 2677 6752 2681 6756
rect 2693 6752 2697 6756
rect 2714 6750 2718 6756
rect 2730 6752 2734 6756
rect 2751 6752 2755 6756
rect 2738 6746 2742 6750
rect 2772 6750 2776 6756
rect 2788 6752 2792 6756
rect 1827 6733 1831 6737
rect 1911 6735 1915 6739
rect 1955 6735 1959 6739
rect 1975 6735 1979 6739
rect 2012 6733 2016 6737
rect 1023 6722 1027 6726
rect 1010 6716 1014 6720
rect 1044 6720 1048 6726
rect 1060 6722 1064 6726
rect 1483 6722 1487 6726
rect 1536 6722 1540 6726
rect 1586 6722 1590 6726
rect 1615 6722 1619 6726
rect 1668 6722 1672 6726
rect 1718 6722 1722 6726
rect 1747 6722 1751 6726
rect 1800 6722 1804 6726
rect 1850 6722 1854 6726
rect 1872 6725 1876 6729
rect 927 6709 931 6713
rect 949 6707 953 6711
rect 965 6707 969 6713
rect 1002 6707 1006 6713
rect 986 6703 990 6707
rect 1010 6707 1014 6711
rect 1023 6707 1027 6713
rect 1060 6707 1064 6713
rect 1073 6712 1077 6716
rect 1457 6715 1463 6719
rect 1894 6717 1898 6726
rect 1910 6722 1914 6726
rect 1931 6720 1935 6726
rect 1947 6722 1951 6726
rect 2413 6737 2417 6741
rect 2429 6737 2433 6743
rect 2466 6737 2470 6743
rect 2450 6733 2454 6737
rect 2474 6737 2478 6741
rect 2487 6737 2491 6743
rect 2524 6737 2528 6743
rect 2545 6737 2549 6743
rect 2561 6737 2565 6743
rect 2598 6737 2602 6743
rect 2508 6733 2512 6737
rect 2582 6733 2586 6737
rect 2606 6737 2610 6741
rect 2619 6737 2623 6743
rect 2656 6737 2660 6743
rect 2677 6737 2681 6743
rect 2693 6737 2697 6743
rect 2730 6737 2734 6743
rect 2640 6733 2644 6737
rect 2714 6733 2718 6737
rect 2738 6737 2742 6741
rect 2751 6737 2755 6743
rect 2788 6737 2792 6743
rect 2801 6742 2805 6746
rect 2772 6733 2776 6737
rect 1968 6722 1972 6726
rect 1955 6716 1959 6720
rect 1989 6720 1993 6726
rect 2005 6722 2009 6726
rect 2428 6722 2432 6726
rect 2481 6722 2485 6726
rect 2531 6722 2535 6726
rect 2560 6722 2564 6726
rect 2613 6722 2617 6726
rect 2663 6722 2667 6726
rect 2692 6722 2696 6726
rect 2745 6722 2749 6726
rect 2795 6722 2799 6726
rect 1397 6708 1403 6712
rect 1483 6708 1487 6712
rect 1550 6708 1554 6712
rect 1586 6708 1590 6712
rect 1615 6708 1619 6712
rect 1682 6708 1686 6712
rect 1718 6708 1722 6712
rect 1747 6708 1751 6712
rect 1814 6708 1818 6712
rect 1850 6708 1854 6712
rect 1872 6709 1876 6713
rect 1894 6707 1898 6711
rect 1910 6707 1914 6713
rect 1947 6707 1951 6713
rect 1044 6703 1048 6707
rect 1468 6700 1472 6704
rect 1857 6700 1861 6704
rect 1931 6703 1935 6707
rect 1955 6707 1959 6711
rect 1968 6707 1972 6713
rect 2005 6707 2009 6713
rect 2018 6712 2022 6716
rect 2402 6715 2408 6719
rect 2342 6708 2348 6712
rect 2428 6708 2432 6712
rect 2495 6708 2499 6712
rect 2531 6708 2535 6712
rect 2560 6708 2564 6712
rect 2627 6708 2631 6712
rect 2663 6708 2667 6712
rect 2692 6708 2696 6712
rect 2759 6708 2763 6712
rect 2795 6708 2799 6712
rect 1989 6703 1993 6707
rect 2413 6700 2417 6704
rect 2802 6700 2806 6704
rect 964 6692 968 6696
rect 1017 6692 1021 6696
rect 1067 6692 1071 6696
rect 1409 6693 1415 6697
rect 1485 6693 1489 6697
rect 1535 6693 1539 6697
rect 1586 6693 1590 6697
rect 1617 6693 1621 6697
rect 1667 6693 1671 6697
rect 1718 6693 1722 6697
rect 1749 6693 1753 6697
rect 1799 6693 1803 6697
rect 1850 6693 1854 6697
rect 1081 6685 1085 6689
rect 1445 6686 1451 6690
rect 1909 6692 1913 6696
rect 1962 6692 1966 6696
rect 2012 6692 2016 6696
rect 2354 6693 2360 6697
rect 2430 6693 2434 6697
rect 2480 6693 2484 6697
rect 2531 6693 2535 6697
rect 2562 6693 2566 6697
rect 2612 6693 2616 6697
rect 2663 6693 2667 6697
rect 2694 6693 2698 6697
rect 2744 6693 2748 6697
rect 2795 6693 2799 6697
rect 964 6678 968 6682
rect 1031 6678 1035 6682
rect 1067 6678 1071 6682
rect 1397 6678 1403 6682
rect 949 6670 953 6674
rect 1074 6671 1078 6675
rect 1485 6679 1489 6683
rect 1529 6679 1533 6683
rect 1549 6679 1553 6683
rect 1586 6677 1590 6681
rect 1617 6679 1621 6683
rect 1661 6679 1665 6683
rect 1681 6679 1685 6683
rect 1718 6677 1722 6681
rect 1749 6679 1753 6683
rect 1793 6679 1797 6683
rect 1813 6679 1817 6683
rect 1850 6677 1854 6681
rect 2026 6685 2030 6689
rect 2390 6686 2396 6690
rect 1909 6678 1913 6682
rect 1976 6678 1980 6682
rect 2012 6678 2016 6682
rect 2342 6678 2348 6682
rect 966 6663 970 6667
rect 1016 6663 1020 6667
rect 1067 6663 1071 6667
rect 1409 6663 1415 6667
rect 1468 6666 1472 6670
rect 1484 6666 1488 6670
rect 1445 6656 1451 6660
rect 1505 6664 1509 6670
rect 1521 6666 1525 6670
rect 1542 6666 1546 6670
rect 1529 6660 1533 6664
rect 1563 6664 1567 6670
rect 1579 6666 1583 6670
rect 1600 6666 1604 6670
rect 1616 6666 1620 6670
rect 1637 6664 1641 6670
rect 1653 6666 1657 6670
rect 1674 6666 1678 6670
rect 1661 6660 1665 6664
rect 1695 6664 1699 6670
rect 1711 6666 1715 6670
rect 1732 6666 1736 6670
rect 1748 6666 1752 6670
rect 1769 6664 1773 6670
rect 1785 6666 1789 6670
rect 1894 6670 1898 6674
rect 2019 6671 2023 6675
rect 2430 6679 2434 6683
rect 2474 6679 2478 6683
rect 2494 6679 2498 6683
rect 2531 6677 2535 6681
rect 2562 6679 2566 6683
rect 2606 6679 2610 6683
rect 2626 6679 2630 6683
rect 2663 6677 2667 6681
rect 2694 6679 2698 6683
rect 2738 6679 2742 6683
rect 2758 6679 2762 6683
rect 2795 6677 2799 6681
rect 1806 6666 1810 6670
rect 1793 6660 1797 6664
rect 1827 6664 1831 6670
rect 1843 6666 1847 6670
rect 1911 6663 1915 6667
rect 1961 6663 1965 6667
rect 2012 6663 2016 6667
rect 2354 6663 2360 6667
rect 2413 6666 2417 6670
rect 2429 6666 2433 6670
rect 966 6649 970 6653
rect 1010 6649 1014 6653
rect 1030 6649 1034 6653
rect 1067 6647 1071 6651
rect 949 6636 953 6640
rect 965 6636 969 6640
rect 986 6634 990 6640
rect 1002 6636 1006 6640
rect 1468 6651 1472 6655
rect 1484 6651 1488 6657
rect 1521 6651 1525 6657
rect 1505 6647 1509 6651
rect 1529 6651 1533 6655
rect 1542 6651 1546 6657
rect 1579 6651 1583 6657
rect 1600 6651 1604 6657
rect 1616 6651 1620 6657
rect 1653 6651 1657 6657
rect 1563 6647 1567 6651
rect 1637 6647 1641 6651
rect 1661 6651 1665 6655
rect 1674 6651 1678 6657
rect 1711 6651 1715 6657
rect 1732 6651 1736 6657
rect 1748 6651 1752 6657
rect 1785 6651 1789 6657
rect 1695 6647 1699 6651
rect 1769 6647 1773 6651
rect 1793 6651 1797 6655
rect 1806 6651 1810 6657
rect 1843 6651 1847 6657
rect 1856 6656 1860 6660
rect 2390 6656 2396 6660
rect 2450 6664 2454 6670
rect 2466 6666 2470 6670
rect 2487 6666 2491 6670
rect 2474 6660 2478 6664
rect 2508 6664 2512 6670
rect 2524 6666 2528 6670
rect 2545 6666 2549 6670
rect 2561 6666 2565 6670
rect 2582 6664 2586 6670
rect 2598 6666 2602 6670
rect 2619 6666 2623 6670
rect 2606 6660 2610 6664
rect 2640 6664 2644 6670
rect 2656 6666 2660 6670
rect 2677 6666 2681 6670
rect 2693 6666 2697 6670
rect 2714 6664 2718 6670
rect 2730 6666 2734 6670
rect 2751 6666 2755 6670
rect 2738 6660 2742 6664
rect 2772 6664 2776 6670
rect 2788 6666 2792 6670
rect 1827 6647 1831 6651
rect 1911 6649 1915 6653
rect 1955 6649 1959 6653
rect 1975 6649 1979 6653
rect 2012 6647 2016 6651
rect 1023 6636 1027 6640
rect 1010 6630 1014 6634
rect 1044 6634 1048 6640
rect 1060 6636 1064 6640
rect 1483 6636 1487 6640
rect 1536 6636 1540 6640
rect 1586 6636 1590 6640
rect 1615 6636 1619 6640
rect 1668 6636 1672 6640
rect 1718 6636 1722 6640
rect 1747 6636 1751 6640
rect 1800 6636 1804 6640
rect 1850 6636 1854 6640
rect 1894 6636 1898 6640
rect 1910 6636 1914 6640
rect 949 6621 953 6627
rect 965 6621 969 6627
rect 1002 6621 1006 6627
rect 986 6617 990 6621
rect 1010 6621 1014 6625
rect 1023 6621 1027 6627
rect 1060 6621 1064 6627
rect 1073 6626 1077 6630
rect 1457 6629 1463 6633
rect 1931 6634 1935 6640
rect 1947 6636 1951 6640
rect 2413 6651 2417 6655
rect 2429 6651 2433 6657
rect 2466 6651 2470 6657
rect 2450 6647 2454 6651
rect 2474 6651 2478 6655
rect 2487 6651 2491 6657
rect 2524 6651 2528 6657
rect 2545 6651 2549 6657
rect 2561 6651 2565 6657
rect 2598 6651 2602 6657
rect 2508 6647 2512 6651
rect 2582 6647 2586 6651
rect 2606 6651 2610 6655
rect 2619 6651 2623 6657
rect 2656 6651 2660 6657
rect 2677 6651 2681 6657
rect 2693 6651 2697 6657
rect 2730 6651 2734 6657
rect 2640 6647 2644 6651
rect 2714 6647 2718 6651
rect 2738 6651 2742 6655
rect 2751 6651 2755 6657
rect 2788 6651 2792 6657
rect 2801 6656 2805 6660
rect 2772 6647 2776 6651
rect 1968 6636 1972 6640
rect 1955 6630 1959 6634
rect 1989 6634 1993 6640
rect 2005 6636 2009 6640
rect 2428 6636 2432 6640
rect 2481 6636 2485 6640
rect 2531 6636 2535 6640
rect 2560 6636 2564 6640
rect 2613 6636 2617 6640
rect 2663 6636 2667 6640
rect 2692 6636 2696 6640
rect 2745 6636 2749 6640
rect 2795 6636 2799 6640
rect 1397 6622 1403 6626
rect 1483 6622 1487 6626
rect 1550 6622 1554 6626
rect 1586 6622 1590 6626
rect 1615 6622 1619 6626
rect 1682 6622 1686 6626
rect 1718 6622 1722 6626
rect 1747 6622 1751 6626
rect 1814 6622 1818 6626
rect 1850 6622 1854 6626
rect 1894 6621 1898 6627
rect 1910 6621 1914 6627
rect 1947 6621 1951 6627
rect 1044 6617 1048 6621
rect 1599 6615 1603 6619
rect 1732 6615 1737 6619
rect 1931 6617 1935 6621
rect 1955 6621 1959 6625
rect 1968 6621 1972 6627
rect 2005 6621 2009 6627
rect 2018 6626 2022 6630
rect 2402 6629 2408 6633
rect 2342 6622 2348 6626
rect 2428 6622 2432 6626
rect 2495 6622 2499 6626
rect 2531 6622 2535 6626
rect 2560 6622 2564 6626
rect 2627 6622 2631 6626
rect 2663 6622 2667 6626
rect 2692 6622 2696 6626
rect 2759 6622 2763 6626
rect 2795 6622 2799 6626
rect 1989 6617 1993 6621
rect 2544 6615 2548 6619
rect 2677 6615 2682 6619
rect 964 6606 968 6610
rect 1017 6606 1021 6610
rect 1067 6606 1071 6610
rect 1725 6608 1729 6612
rect 1709 6604 1713 6608
rect 1741 6604 1745 6608
rect 1081 6599 1085 6603
rect 1457 6599 1463 6603
rect 1468 6600 1472 6604
rect 1909 6606 1913 6610
rect 1962 6606 1966 6610
rect 2012 6606 2016 6610
rect 2670 6608 2674 6612
rect 2654 6604 2658 6608
rect 2686 6604 2690 6608
rect 2026 6599 2030 6603
rect 2402 6599 2408 6603
rect 2413 6600 2417 6604
rect 964 6592 968 6596
rect 1031 6592 1035 6596
rect 1067 6592 1071 6596
rect 1397 6592 1403 6596
rect 1468 6592 1472 6596
rect 1725 6592 1729 6596
rect 1909 6592 1913 6596
rect 1976 6592 1980 6596
rect 2012 6592 2016 6596
rect 2342 6592 2348 6596
rect 2413 6592 2417 6596
rect 2670 6592 2674 6596
rect 1709 6585 1713 6589
rect 1741 6585 1745 6589
rect 2654 6585 2658 6589
rect 2686 6585 2690 6589
rect 1385 6578 1391 6582
rect 1709 6576 1713 6580
rect 1741 6576 1745 6580
rect 950 6571 954 6575
rect 1115 6571 1119 6575
rect 1433 6572 1439 6576
rect 1725 6572 1729 6576
rect 2330 6578 2336 6582
rect 2654 6576 2658 6580
rect 2686 6576 2690 6580
rect 1895 6571 1899 6575
rect 2060 6571 2064 6575
rect 2378 6572 2384 6576
rect 2670 6572 2674 6576
rect 927 6563 931 6567
rect 939 6563 943 6567
rect 1125 6564 1129 6568
rect 1359 6564 1363 6568
rect 1421 6564 1427 6568
rect 1600 6565 1604 6569
rect 1732 6565 1737 6569
rect 1872 6563 1876 6567
rect 1884 6563 1888 6567
rect 2070 6564 2074 6568
rect 2304 6564 2308 6568
rect 2366 6564 2372 6568
rect 2545 6565 2549 6569
rect 2677 6565 2682 6569
rect 955 6557 959 6561
rect 983 6557 987 6561
rect 1000 6557 1004 6561
rect 1056 6557 1060 6561
rect 1073 6557 1077 6561
rect 1107 6557 1111 6561
rect 1133 6557 1137 6561
rect 1216 6557 1220 6561
rect 1244 6557 1248 6561
rect 1261 6557 1265 6561
rect 1317 6557 1321 6561
rect 1334 6557 1338 6561
rect 1368 6557 1372 6561
rect 1457 6557 1463 6561
rect 1468 6558 1472 6562
rect 1856 6558 1860 6562
rect 1900 6557 1904 6561
rect 1928 6557 1932 6561
rect 1945 6557 1949 6561
rect 2001 6557 2005 6561
rect 2018 6557 2022 6561
rect 2052 6557 2056 6561
rect 2078 6557 2082 6561
rect 2161 6557 2165 6561
rect 2189 6557 2193 6561
rect 2206 6557 2210 6561
rect 2262 6557 2266 6561
rect 2279 6557 2283 6561
rect 2313 6557 2317 6561
rect 2402 6557 2408 6561
rect 2413 6558 2417 6562
rect 2801 6558 2805 6562
rect 962 6550 966 6554
rect 1027 6550 1031 6554
rect 1049 6550 1053 6554
rect 1080 6550 1084 6554
rect 1124 6550 1128 6554
rect 1163 6550 1167 6554
rect 956 6540 960 6544
rect 963 6543 967 6547
rect 983 6540 987 6544
rect 999 6540 1003 6544
rect 1009 6543 1013 6547
rect 1034 6543 1038 6547
rect 1056 6540 1060 6544
rect 1074 6540 1078 6544
rect 1081 6543 1085 6547
rect 1223 6550 1227 6554
rect 1288 6550 1292 6554
rect 1310 6550 1314 6554
rect 1341 6550 1345 6554
rect 1359 6550 1363 6554
rect 1409 6550 1415 6554
rect 1485 6551 1489 6555
rect 1535 6551 1539 6555
rect 1586 6551 1590 6555
rect 1617 6551 1621 6555
rect 1667 6551 1671 6555
rect 1718 6551 1722 6555
rect 1749 6551 1753 6555
rect 1799 6551 1803 6555
rect 1850 6551 1854 6555
rect 1907 6550 1911 6554
rect 1972 6550 1976 6554
rect 1994 6550 1998 6554
rect 2025 6550 2029 6554
rect 2069 6550 2073 6554
rect 2108 6550 2112 6554
rect 1107 6540 1111 6544
rect 1133 6540 1137 6544
rect 618 6536 622 6540
rect 628 6536 632 6540
rect 638 6536 642 6540
rect 618 6531 622 6535
rect 628 6531 632 6535
rect 638 6531 642 6535
rect 618 6526 622 6530
rect 628 6526 632 6530
rect 638 6526 642 6530
rect 618 6521 622 6525
rect 628 6521 632 6525
rect 638 6521 642 6525
rect 664 6536 668 6540
rect 674 6536 678 6540
rect 684 6536 688 6540
rect 664 6531 668 6535
rect 674 6531 678 6535
rect 684 6531 688 6535
rect 664 6526 668 6530
rect 674 6526 678 6530
rect 684 6526 688 6530
rect 664 6521 668 6525
rect 674 6521 678 6525
rect 684 6521 688 6525
rect 947 6523 951 6527
rect 959 6523 963 6527
rect 967 6524 971 6528
rect 989 6523 993 6527
rect 1002 6524 1006 6528
rect 1021 6524 1025 6528
rect 1040 6525 1044 6529
rect 1059 6521 1063 6525
rect 1079 6524 1083 6528
rect 1217 6540 1221 6544
rect 1224 6543 1228 6547
rect 1244 6540 1248 6544
rect 1260 6540 1264 6544
rect 1270 6543 1274 6547
rect 1295 6543 1299 6547
rect 1317 6540 1321 6544
rect 1335 6540 1339 6544
rect 1342 6543 1346 6547
rect 1445 6544 1451 6548
rect 1367 6540 1371 6544
rect 1145 6530 1149 6534
rect 1134 6523 1138 6527
rect 1174 6529 1178 6533
rect 1208 6523 1212 6527
rect 1220 6523 1224 6527
rect 1228 6524 1232 6528
rect 1153 6514 1157 6518
rect 956 6510 960 6514
rect 984 6510 988 6514
rect 999 6510 1003 6514
rect 1056 6510 1060 6514
rect 1074 6510 1078 6514
rect 977 6505 981 6509
rect 1024 6506 1031 6510
rect 1049 6505 1053 6509
rect 1092 6506 1096 6510
rect 977 6498 981 6502
rect 1008 6498 1012 6502
rect 1033 6498 1037 6502
rect 1092 6498 1096 6502
rect 1114 6498 1118 6502
rect 1250 6523 1254 6527
rect 1263 6524 1267 6528
rect 1282 6524 1286 6528
rect 1301 6525 1305 6529
rect 1320 6521 1324 6525
rect 1340 6524 1344 6528
rect 1485 6537 1489 6541
rect 1529 6537 1533 6541
rect 1549 6537 1553 6541
rect 1586 6535 1590 6539
rect 1617 6537 1621 6541
rect 1661 6537 1665 6541
rect 1681 6537 1685 6541
rect 1718 6535 1722 6539
rect 1749 6537 1753 6541
rect 1793 6537 1797 6541
rect 1813 6537 1817 6541
rect 1850 6535 1854 6539
rect 1901 6540 1905 6544
rect 1908 6543 1912 6547
rect 1928 6540 1932 6544
rect 1944 6540 1948 6544
rect 1954 6543 1958 6547
rect 1979 6543 1983 6547
rect 2001 6540 2005 6544
rect 2019 6540 2023 6544
rect 2026 6543 2030 6547
rect 2168 6550 2172 6554
rect 2233 6550 2237 6554
rect 2255 6550 2259 6554
rect 2286 6550 2290 6554
rect 2304 6550 2308 6554
rect 2354 6550 2360 6554
rect 2430 6551 2434 6555
rect 2480 6551 2484 6555
rect 2531 6551 2535 6555
rect 2562 6551 2566 6555
rect 2612 6551 2616 6555
rect 2663 6551 2667 6555
rect 2694 6551 2698 6555
rect 2744 6551 2748 6555
rect 2795 6551 2799 6555
rect 4484 6549 4488 6553
rect 4494 6549 4498 6553
rect 4504 6549 4508 6553
rect 2052 6540 2056 6544
rect 2078 6540 2082 6544
rect 1372 6522 1376 6526
rect 1468 6524 1472 6528
rect 1484 6524 1488 6528
rect 1505 6522 1509 6528
rect 1521 6524 1525 6528
rect 1542 6524 1546 6528
rect 1529 6518 1533 6522
rect 1563 6522 1567 6528
rect 1579 6524 1583 6528
rect 1600 6524 1604 6528
rect 1616 6524 1620 6528
rect 1637 6522 1641 6528
rect 1653 6524 1657 6528
rect 1674 6524 1678 6528
rect 1661 6518 1665 6522
rect 1695 6522 1699 6528
rect 1711 6524 1715 6528
rect 1732 6524 1736 6528
rect 1748 6524 1752 6528
rect 1769 6522 1773 6528
rect 1785 6524 1789 6528
rect 1806 6524 1810 6528
rect 1793 6518 1797 6522
rect 1827 6522 1831 6528
rect 1843 6524 1847 6528
rect 1892 6523 1896 6527
rect 1904 6523 1908 6527
rect 1912 6524 1916 6528
rect 1934 6523 1938 6527
rect 1947 6524 1951 6528
rect 1966 6524 1970 6528
rect 1217 6510 1221 6514
rect 1245 6510 1249 6514
rect 1260 6510 1264 6514
rect 1317 6510 1321 6514
rect 1335 6510 1339 6514
rect 1367 6510 1371 6514
rect 1238 6505 1242 6509
rect 1285 6506 1292 6510
rect 1310 6505 1314 6509
rect 1353 6506 1357 6510
rect 1468 6509 1472 6513
rect 1484 6509 1488 6515
rect 1521 6509 1525 6515
rect 1238 6498 1242 6502
rect 1269 6498 1273 6502
rect 1294 6498 1298 6502
rect 1344 6498 1348 6502
rect 1353 6498 1357 6502
rect 1433 6498 1439 6502
rect 1505 6505 1509 6509
rect 1529 6509 1533 6513
rect 1542 6509 1546 6515
rect 1579 6509 1583 6515
rect 1600 6509 1604 6515
rect 1616 6509 1620 6515
rect 1653 6509 1657 6515
rect 1563 6505 1567 6509
rect 1637 6505 1641 6509
rect 1661 6509 1665 6513
rect 1674 6509 1678 6515
rect 1711 6509 1715 6515
rect 1732 6509 1736 6515
rect 1748 6509 1752 6515
rect 1785 6509 1789 6515
rect 1695 6505 1699 6509
rect 1769 6505 1773 6509
rect 1793 6509 1797 6513
rect 1806 6509 1810 6515
rect 1843 6509 1847 6515
rect 1856 6514 1860 6518
rect 1985 6525 1989 6529
rect 2004 6521 2008 6525
rect 2024 6524 2028 6528
rect 2162 6540 2166 6544
rect 2169 6543 2173 6547
rect 2189 6540 2193 6544
rect 2205 6540 2209 6544
rect 2215 6543 2219 6547
rect 2240 6543 2244 6547
rect 2262 6540 2266 6544
rect 2280 6540 2284 6544
rect 2287 6543 2291 6547
rect 2390 6544 2396 6548
rect 4484 6544 4488 6548
rect 4494 6544 4498 6548
rect 4504 6544 4508 6548
rect 2312 6540 2316 6544
rect 2090 6530 2094 6534
rect 2079 6523 2083 6527
rect 2119 6529 2123 6533
rect 2153 6523 2157 6527
rect 2165 6523 2169 6527
rect 2173 6524 2177 6528
rect 2098 6514 2102 6518
rect 1901 6510 1905 6514
rect 1929 6510 1933 6514
rect 1944 6510 1948 6514
rect 2001 6510 2005 6514
rect 2019 6510 2023 6514
rect 1827 6505 1831 6509
rect 1922 6505 1926 6509
rect 1969 6506 1976 6510
rect 1994 6505 1998 6509
rect 2037 6506 2041 6510
rect 579 6491 583 6495
rect 584 6491 588 6495
rect 589 6491 593 6495
rect 594 6491 598 6495
rect 599 6491 603 6495
rect 604 6491 608 6495
rect 609 6491 613 6495
rect 614 6491 618 6495
rect 619 6491 623 6495
rect 624 6491 628 6495
rect 629 6491 633 6495
rect 634 6491 638 6495
rect 639 6491 643 6495
rect 956 6491 960 6495
rect 984 6491 988 6495
rect 999 6491 1003 6495
rect 1033 6491 1037 6495
rect 1056 6491 1060 6495
rect 1074 6491 1078 6495
rect 1092 6491 1096 6495
rect 1217 6491 1221 6495
rect 1245 6491 1249 6495
rect 1260 6491 1264 6495
rect 1294 6491 1298 6495
rect 1317 6491 1321 6495
rect 1335 6491 1339 6495
rect 1353 6491 1357 6495
rect 1367 6491 1371 6495
rect 1445 6491 1451 6495
rect 1483 6494 1487 6498
rect 1536 6494 1540 6498
rect 1586 6494 1590 6498
rect 1615 6494 1619 6498
rect 1668 6494 1672 6498
rect 1718 6494 1722 6498
rect 1747 6494 1751 6498
rect 1800 6494 1804 6498
rect 1850 6494 1854 6498
rect 1922 6498 1926 6502
rect 1953 6498 1957 6502
rect 1978 6498 1982 6502
rect 2037 6498 2041 6502
rect 2059 6498 2063 6502
rect 2195 6523 2199 6527
rect 2208 6524 2212 6528
rect 2227 6524 2231 6528
rect 2246 6525 2250 6529
rect 2265 6521 2269 6525
rect 2285 6524 2289 6528
rect 2430 6537 2434 6541
rect 2474 6537 2478 6541
rect 2494 6537 2498 6541
rect 2531 6535 2535 6539
rect 2562 6537 2566 6541
rect 2606 6537 2610 6541
rect 2626 6537 2630 6541
rect 2663 6535 2667 6539
rect 2694 6537 2698 6541
rect 2738 6537 2742 6541
rect 2758 6537 2762 6541
rect 2795 6535 2799 6539
rect 4484 6539 4488 6543
rect 4494 6539 4498 6543
rect 4504 6539 4508 6543
rect 4484 6534 4488 6538
rect 4494 6534 4498 6538
rect 4504 6534 4508 6538
rect 4530 6549 4534 6553
rect 4540 6549 4544 6553
rect 4550 6549 4554 6553
rect 4530 6544 4534 6548
rect 4540 6544 4544 6548
rect 4550 6544 4554 6548
rect 4530 6539 4534 6543
rect 4540 6539 4544 6543
rect 4550 6539 4554 6543
rect 4530 6534 4534 6538
rect 4540 6534 4544 6538
rect 4550 6534 4554 6538
rect 2317 6522 2321 6526
rect 2413 6524 2417 6528
rect 2429 6524 2433 6528
rect 2450 6522 2454 6528
rect 2466 6524 2470 6528
rect 2487 6524 2491 6528
rect 2474 6518 2478 6522
rect 2508 6522 2512 6528
rect 2524 6524 2528 6528
rect 2545 6524 2549 6528
rect 2561 6524 2565 6528
rect 2582 6522 2586 6528
rect 2598 6524 2602 6528
rect 2619 6524 2623 6528
rect 2606 6518 2610 6522
rect 2640 6522 2644 6528
rect 2656 6524 2660 6528
rect 2677 6524 2681 6528
rect 2693 6524 2697 6528
rect 2714 6522 2718 6528
rect 2730 6524 2734 6528
rect 2751 6524 2755 6528
rect 2738 6518 2742 6522
rect 2772 6522 2776 6528
rect 2788 6524 2792 6528
rect 2162 6510 2166 6514
rect 2190 6510 2194 6514
rect 2205 6510 2209 6514
rect 2262 6510 2266 6514
rect 2280 6510 2284 6514
rect 2312 6510 2316 6514
rect 2183 6505 2187 6509
rect 2230 6506 2237 6510
rect 2255 6505 2259 6509
rect 2298 6506 2302 6510
rect 2413 6509 2417 6513
rect 2429 6509 2433 6515
rect 2466 6509 2470 6515
rect 2183 6498 2187 6502
rect 2214 6498 2218 6502
rect 2239 6498 2243 6502
rect 2289 6498 2293 6502
rect 2298 6498 2302 6502
rect 2378 6498 2384 6502
rect 2450 6505 2454 6509
rect 2474 6509 2478 6513
rect 2487 6509 2491 6515
rect 2524 6509 2528 6515
rect 2545 6509 2549 6515
rect 2561 6509 2565 6515
rect 2598 6509 2602 6515
rect 2508 6505 2512 6509
rect 2582 6505 2586 6509
rect 2606 6509 2610 6513
rect 2619 6509 2623 6515
rect 2656 6509 2660 6515
rect 2677 6509 2681 6515
rect 2693 6509 2697 6515
rect 2730 6509 2734 6515
rect 2640 6505 2644 6509
rect 2714 6505 2718 6509
rect 2738 6509 2742 6513
rect 2751 6509 2755 6515
rect 2788 6509 2792 6515
rect 2801 6514 2805 6518
rect 2772 6505 2776 6509
rect 1901 6491 1905 6495
rect 1929 6491 1933 6495
rect 1944 6491 1948 6495
rect 1978 6491 1982 6495
rect 2001 6491 2005 6495
rect 2019 6491 2023 6495
rect 2037 6491 2041 6495
rect 2162 6491 2166 6495
rect 2190 6491 2194 6495
rect 2205 6491 2209 6495
rect 2239 6491 2243 6495
rect 2262 6491 2266 6495
rect 2280 6491 2284 6495
rect 2298 6491 2302 6495
rect 2312 6491 2316 6495
rect 2390 6491 2396 6495
rect 2428 6494 2432 6498
rect 2481 6494 2485 6498
rect 2531 6494 2535 6498
rect 2560 6494 2564 6498
rect 2613 6494 2617 6498
rect 2663 6494 2667 6498
rect 2692 6494 2696 6498
rect 2745 6494 2749 6498
rect 2795 6494 2799 6498
rect 579 6486 583 6490
rect 584 6486 588 6490
rect 589 6486 593 6490
rect 594 6486 598 6490
rect 599 6486 603 6490
rect 604 6486 608 6490
rect 609 6486 613 6490
rect 614 6486 618 6490
rect 619 6486 623 6490
rect 624 6486 628 6490
rect 629 6486 633 6490
rect 634 6486 638 6490
rect 639 6486 643 6490
rect 1163 6468 1167 6472
rect 423 6386 427 6390
rect 439 6386 443 6390
rect 464 6386 468 6390
rect 480 6386 484 6390
rect 507 6386 511 6390
rect 523 6386 527 6390
rect 1238 6484 1242 6488
rect 1269 6484 1273 6488
rect 1294 6484 1298 6488
rect 1344 6484 1348 6488
rect 1353 6484 1357 6488
rect 1457 6487 1463 6491
rect 1238 6477 1242 6481
rect 1285 6476 1292 6480
rect 1310 6477 1314 6481
rect 1397 6480 1403 6484
rect 1483 6480 1487 6484
rect 1550 6480 1554 6484
rect 1586 6480 1590 6484
rect 1615 6480 1619 6484
rect 1682 6480 1686 6484
rect 1718 6480 1722 6484
rect 1747 6480 1751 6484
rect 1814 6480 1818 6484
rect 1850 6480 1854 6484
rect 1353 6476 1357 6480
rect 1217 6472 1221 6476
rect 1245 6472 1249 6476
rect 1260 6472 1264 6476
rect 1317 6472 1321 6476
rect 1335 6472 1339 6476
rect 1367 6472 1371 6476
rect 1122 6455 1126 6459
rect 1176 6460 1180 6464
rect 1145 6450 1149 6458
rect 1208 6459 1212 6463
rect 1220 6459 1224 6463
rect 1228 6458 1232 6462
rect 1250 6459 1254 6463
rect 1263 6458 1267 6462
rect 1282 6458 1286 6462
rect 1301 6457 1305 6461
rect 1320 6461 1324 6465
rect 1340 6458 1344 6462
rect 2108 6468 2112 6472
rect 2183 6484 2187 6488
rect 2214 6484 2218 6488
rect 2239 6484 2243 6488
rect 2289 6484 2293 6488
rect 2298 6484 2302 6488
rect 2402 6487 2408 6491
rect 2183 6477 2187 6481
rect 2230 6476 2237 6480
rect 2255 6477 2259 6481
rect 2342 6480 2348 6484
rect 2428 6480 2432 6484
rect 2495 6480 2499 6484
rect 2531 6480 2535 6484
rect 2560 6480 2564 6484
rect 2627 6480 2631 6484
rect 2663 6480 2667 6484
rect 2692 6480 2696 6484
rect 2759 6480 2763 6484
rect 2795 6480 2799 6484
rect 2298 6476 2302 6480
rect 2162 6472 2166 6476
rect 2190 6472 2194 6476
rect 2205 6472 2209 6476
rect 2262 6472 2266 6476
rect 2280 6472 2284 6476
rect 2312 6472 2316 6476
rect 1373 6459 1377 6463
rect 2067 6455 2071 6459
rect 2121 6460 2125 6464
rect 1217 6442 1221 6446
rect 1224 6439 1228 6443
rect 1244 6442 1248 6446
rect 1260 6442 1264 6446
rect 1270 6439 1274 6443
rect 1295 6439 1299 6443
rect 1317 6442 1321 6446
rect 1335 6442 1339 6446
rect 1342 6439 1346 6443
rect 1367 6442 1371 6446
rect 2090 6450 2094 6458
rect 2153 6459 2157 6463
rect 2165 6459 2169 6463
rect 2173 6458 2177 6462
rect 2195 6459 2199 6463
rect 2208 6458 2212 6462
rect 2227 6458 2231 6462
rect 1153 6432 1157 6436
rect 1223 6432 1227 6436
rect 1288 6432 1292 6436
rect 1310 6432 1314 6436
rect 1341 6432 1345 6436
rect 1421 6432 1427 6436
rect 2246 6457 2250 6461
rect 2265 6461 2269 6465
rect 2285 6458 2289 6462
rect 2318 6459 2322 6463
rect 2162 6442 2166 6446
rect 2169 6439 2173 6443
rect 2189 6442 2193 6446
rect 2205 6442 2209 6446
rect 2215 6439 2219 6443
rect 2240 6439 2244 6443
rect 2262 6442 2266 6446
rect 2280 6442 2284 6446
rect 2287 6439 2291 6443
rect 2312 6442 2316 6446
rect 2098 6432 2102 6436
rect 2168 6432 2172 6436
rect 2233 6432 2237 6436
rect 2255 6432 2259 6436
rect 2286 6432 2290 6436
rect 2366 6432 2372 6436
rect 1216 6425 1220 6429
rect 1244 6425 1248 6429
rect 1261 6425 1265 6429
rect 1317 6425 1321 6429
rect 1334 6425 1338 6429
rect 1368 6425 1372 6429
rect 1457 6425 1463 6429
rect 2161 6425 2165 6429
rect 2189 6425 2193 6429
rect 2206 6425 2210 6429
rect 2262 6425 2266 6429
rect 2279 6425 2283 6429
rect 2313 6425 2317 6429
rect 2402 6425 2408 6429
rect 546 6386 550 6390
rect 562 6386 566 6390
rect 578 6386 582 6390
rect 992 6414 996 6418
rect 1082 6414 1086 6418
rect 1163 6414 1167 6418
rect 1223 6418 1227 6422
rect 1288 6418 1292 6422
rect 1310 6418 1314 6422
rect 1341 6418 1345 6422
rect 1421 6418 1427 6422
rect 1217 6408 1221 6412
rect 1224 6411 1228 6415
rect 1244 6408 1248 6412
rect 1260 6408 1264 6412
rect 1270 6411 1274 6415
rect 1295 6411 1299 6415
rect 1317 6408 1321 6412
rect 1335 6408 1339 6412
rect 1342 6411 1346 6415
rect 1937 6414 1941 6418
rect 1367 6408 1371 6412
rect 2027 6414 2031 6418
rect 2108 6414 2112 6418
rect 2168 6418 2172 6422
rect 2233 6418 2237 6422
rect 2255 6418 2259 6422
rect 2286 6418 2290 6422
rect 2366 6418 2372 6422
rect 974 6394 978 6398
rect 594 6386 598 6390
rect 1009 6393 1013 6397
rect 1064 6394 1068 6398
rect 1093 6393 1097 6397
rect 1145 6394 1149 6398
rect 1173 6393 1177 6397
rect 1208 6391 1212 6395
rect 1220 6391 1224 6395
rect 1228 6392 1232 6396
rect 982 6378 986 6382
rect 461 6351 469 6360
rect 505 6351 513 6360
rect 803 6351 812 6364
rect 1072 6378 1076 6382
rect 1153 6378 1157 6382
rect 1250 6391 1254 6395
rect 1263 6392 1267 6396
rect 1282 6392 1286 6396
rect 1301 6393 1305 6397
rect 1320 6389 1324 6393
rect 1340 6392 1344 6396
rect 2162 6408 2166 6412
rect 2169 6411 2173 6415
rect 2189 6408 2193 6412
rect 2205 6408 2209 6412
rect 2215 6411 2219 6415
rect 2240 6411 2244 6415
rect 2262 6408 2266 6412
rect 2280 6408 2284 6412
rect 2287 6411 2291 6415
rect 2312 6408 2316 6412
rect 1919 6394 1923 6398
rect 1372 6390 1376 6394
rect 1954 6393 1958 6397
rect 2009 6394 2013 6398
rect 2038 6393 2042 6397
rect 2090 6394 2094 6398
rect 2118 6393 2122 6397
rect 2153 6391 2157 6395
rect 2165 6391 2169 6395
rect 2173 6392 2177 6396
rect 1217 6378 1221 6382
rect 1245 6378 1249 6382
rect 1260 6378 1264 6382
rect 1317 6378 1321 6382
rect 1335 6378 1339 6382
rect 1367 6378 1371 6382
rect 1927 6378 1931 6382
rect 1238 6373 1242 6377
rect 1285 6374 1292 6378
rect 1310 6373 1314 6377
rect 1353 6374 1357 6378
rect 1238 6366 1242 6370
rect 1269 6366 1273 6370
rect 1294 6366 1298 6370
rect 1353 6366 1357 6370
rect 1433 6366 1439 6370
rect 2017 6378 2021 6382
rect 2098 6378 2102 6382
rect 2195 6391 2199 6395
rect 2208 6392 2212 6396
rect 2227 6392 2231 6396
rect 2246 6393 2250 6397
rect 2265 6389 2269 6393
rect 2285 6392 2289 6396
rect 2317 6390 2321 6394
rect 2162 6378 2166 6382
rect 2190 6378 2194 6382
rect 2205 6378 2209 6382
rect 2262 6378 2266 6382
rect 2280 6378 2284 6382
rect 2312 6378 2316 6382
rect 2183 6373 2187 6377
rect 2230 6374 2237 6378
rect 2255 6373 2259 6377
rect 2298 6374 2302 6378
rect 2183 6366 2187 6370
rect 2214 6366 2218 6370
rect 2239 6366 2243 6370
rect 2298 6366 2302 6370
rect 2378 6366 2384 6370
rect 1217 6359 1221 6363
rect 1245 6359 1249 6363
rect 1260 6359 1264 6363
rect 1294 6359 1298 6363
rect 1317 6359 1321 6363
rect 1335 6359 1339 6363
rect 1353 6359 1357 6363
rect 1367 6359 1371 6363
rect 1445 6359 1451 6363
rect 2162 6359 2166 6363
rect 2190 6359 2194 6363
rect 2205 6359 2209 6363
rect 2239 6359 2243 6363
rect 2262 6359 2266 6363
rect 2280 6359 2284 6363
rect 2298 6359 2302 6363
rect 2312 6359 2316 6363
rect 2390 6359 2396 6363
rect 423 6328 427 6332
rect 439 6328 443 6332
rect 464 6328 468 6332
rect 480 6328 484 6332
rect 507 6328 511 6332
rect 523 6328 527 6332
rect 546 6328 550 6332
rect 562 6328 566 6332
rect 578 6328 582 6332
rect 992 6336 996 6340
rect 594 6328 598 6332
rect 939 6323 943 6327
rect 1082 6336 1086 6340
rect 974 6318 978 6326
rect 1006 6320 1010 6324
rect 1095 6328 1099 6332
rect 1040 6322 1044 6326
rect 1013 6314 1017 6318
rect 1028 6314 1032 6318
rect 982 6300 986 6304
rect 1064 6318 1068 6326
rect 1163 6336 1167 6340
rect 1238 6352 1242 6356
rect 1269 6352 1273 6356
rect 1294 6352 1298 6356
rect 1353 6352 1357 6356
rect 1433 6352 1439 6356
rect 1238 6345 1242 6349
rect 1285 6344 1292 6348
rect 1310 6345 1314 6349
rect 1353 6344 1357 6348
rect 1217 6340 1221 6344
rect 1245 6340 1249 6344
rect 1260 6340 1264 6344
rect 1317 6340 1321 6344
rect 1335 6340 1339 6344
rect 1367 6340 1371 6344
rect 1176 6328 1180 6332
rect 1122 6322 1126 6326
rect 1103 6314 1107 6318
rect 1118 6314 1122 6318
rect 1072 6300 1076 6304
rect 1145 6318 1149 6326
rect 1208 6327 1212 6331
rect 1220 6327 1224 6331
rect 1228 6326 1232 6330
rect 1250 6327 1254 6331
rect 1263 6326 1267 6330
rect 1282 6326 1286 6330
rect 1301 6325 1305 6329
rect 1320 6329 1324 6333
rect 1340 6326 1344 6330
rect 1937 6336 1941 6340
rect 1373 6327 1377 6331
rect 1884 6323 1888 6327
rect 2027 6336 2031 6340
rect 1217 6310 1221 6314
rect 1224 6307 1228 6311
rect 1244 6310 1248 6314
rect 1260 6310 1264 6314
rect 1270 6307 1274 6311
rect 1295 6307 1299 6311
rect 1317 6310 1321 6314
rect 1335 6310 1339 6314
rect 1342 6307 1346 6311
rect 1367 6310 1371 6314
rect 1919 6318 1923 6326
rect 1951 6320 1955 6324
rect 2040 6328 2044 6332
rect 1985 6322 1989 6326
rect 1153 6300 1157 6304
rect 1223 6300 1227 6304
rect 1288 6300 1292 6304
rect 1310 6300 1314 6304
rect 1341 6300 1345 6304
rect 1421 6300 1427 6304
rect 1958 6314 1962 6318
rect 1973 6314 1977 6318
rect 1927 6300 1931 6304
rect 2009 6318 2013 6326
rect 2108 6336 2112 6340
rect 2183 6352 2187 6356
rect 2214 6352 2218 6356
rect 2239 6352 2243 6356
rect 2298 6352 2302 6356
rect 2378 6352 2384 6356
rect 2183 6345 2187 6349
rect 2230 6344 2237 6348
rect 2255 6345 2259 6349
rect 2298 6344 2302 6348
rect 2162 6340 2166 6344
rect 2190 6340 2194 6344
rect 2205 6340 2209 6344
rect 2262 6340 2266 6344
rect 2280 6340 2284 6344
rect 2312 6340 2316 6344
rect 2121 6328 2125 6332
rect 2067 6322 2071 6326
rect 2048 6314 2052 6318
rect 2063 6314 2067 6318
rect 2017 6300 2021 6304
rect 2090 6318 2094 6326
rect 2153 6327 2157 6331
rect 2165 6327 2169 6331
rect 2173 6326 2177 6330
rect 2195 6327 2199 6331
rect 2208 6326 2212 6330
rect 2227 6326 2231 6330
rect 2246 6325 2250 6329
rect 2265 6329 2269 6333
rect 2285 6326 2289 6330
rect 2318 6327 2322 6331
rect 2162 6310 2166 6314
rect 2169 6307 2173 6311
rect 2189 6310 2193 6314
rect 2205 6310 2209 6314
rect 2215 6307 2219 6311
rect 2240 6307 2244 6311
rect 2262 6310 2266 6314
rect 2280 6310 2284 6314
rect 2287 6307 2291 6311
rect 2312 6310 2316 6314
rect 2098 6300 2102 6304
rect 2168 6300 2172 6304
rect 2233 6300 2237 6304
rect 2255 6300 2259 6304
rect 2286 6300 2290 6304
rect 2366 6300 2372 6304
rect 1216 6293 1220 6297
rect 1244 6293 1248 6297
rect 1261 6293 1265 6297
rect 1317 6293 1321 6297
rect 1334 6293 1338 6297
rect 1368 6293 1372 6297
rect 1457 6293 1463 6297
rect 2161 6293 2165 6297
rect 2189 6293 2193 6297
rect 2206 6293 2210 6297
rect 2262 6293 2266 6297
rect 2279 6293 2283 6297
rect 2313 6293 2317 6297
rect 2402 6293 2408 6297
rect 657 6286 661 6290
rect 662 6286 666 6290
rect 657 6281 661 6285
rect 662 6281 666 6285
rect 657 6276 661 6280
rect 662 6276 666 6280
rect 1058 6279 1062 6283
rect 657 6271 661 6275
rect 662 6271 666 6275
rect 1163 6279 1167 6283
rect 1223 6286 1227 6290
rect 1288 6286 1292 6290
rect 1310 6286 1314 6290
rect 1341 6286 1345 6290
rect 1421 6286 1427 6290
rect 1217 6276 1221 6280
rect 1224 6279 1228 6283
rect 1244 6276 1248 6280
rect 1260 6276 1264 6280
rect 1270 6279 1274 6283
rect 1295 6279 1299 6283
rect 1317 6276 1321 6280
rect 1335 6276 1339 6280
rect 1342 6279 1346 6283
rect 1367 6276 1371 6280
rect 2003 6279 2007 6283
rect 657 6266 661 6270
rect 662 6266 666 6270
rect 657 6261 661 6265
rect 662 6261 666 6265
rect 657 6256 661 6260
rect 662 6256 666 6260
rect 1040 6259 1044 6263
rect 657 6251 661 6255
rect 662 6251 666 6255
rect 1068 6258 1072 6262
rect 1145 6259 1149 6263
rect 1174 6258 1178 6262
rect 1208 6259 1212 6263
rect 1220 6259 1224 6263
rect 1228 6260 1232 6264
rect 1250 6259 1254 6263
rect 1263 6260 1267 6264
rect 1282 6260 1286 6264
rect 1301 6261 1305 6265
rect 1320 6257 1324 6261
rect 1340 6260 1344 6264
rect 2108 6279 2112 6283
rect 2168 6286 2172 6290
rect 2233 6286 2237 6290
rect 2255 6286 2259 6290
rect 2286 6286 2290 6290
rect 2366 6286 2372 6290
rect 2162 6276 2166 6280
rect 2169 6279 2173 6283
rect 2189 6276 2193 6280
rect 2205 6276 2209 6280
rect 2215 6279 2219 6283
rect 2240 6279 2244 6283
rect 2262 6276 2266 6280
rect 2280 6276 2284 6280
rect 2287 6279 2291 6283
rect 2312 6276 2316 6280
rect 1372 6258 1376 6262
rect 1985 6259 1989 6263
rect 2013 6258 2017 6262
rect 2090 6259 2094 6263
rect 2119 6258 2123 6262
rect 2153 6259 2157 6263
rect 2165 6259 2169 6263
rect 2173 6260 2177 6264
rect 2195 6259 2199 6263
rect 2208 6260 2212 6264
rect 2227 6260 2231 6264
rect 2246 6261 2250 6265
rect 2265 6257 2269 6261
rect 2285 6260 2289 6264
rect 2317 6258 2321 6262
rect 657 6246 661 6250
rect 662 6246 666 6250
rect 657 6241 661 6245
rect 662 6241 666 6245
rect 1048 6243 1052 6247
rect 657 6236 661 6240
rect 662 6236 666 6240
rect 1153 6243 1157 6247
rect 1217 6246 1221 6250
rect 1245 6246 1249 6250
rect 1260 6246 1264 6250
rect 1317 6246 1321 6250
rect 1335 6246 1339 6250
rect 1367 6246 1371 6250
rect 1238 6241 1242 6245
rect 1285 6242 1292 6246
rect 1310 6241 1314 6245
rect 1353 6242 1357 6246
rect 1993 6243 1997 6247
rect 1238 6234 1242 6238
rect 1269 6234 1273 6238
rect 1294 6234 1298 6238
rect 1353 6234 1357 6238
rect 1433 6234 1439 6238
rect 2098 6243 2102 6247
rect 2162 6246 2166 6250
rect 2190 6246 2194 6250
rect 2205 6246 2209 6250
rect 2262 6246 2266 6250
rect 2280 6246 2284 6250
rect 2312 6246 2316 6250
rect 2183 6241 2187 6245
rect 2230 6242 2237 6246
rect 2255 6241 2259 6245
rect 2298 6242 2302 6246
rect 4484 6240 4488 6244
rect 4494 6240 4498 6244
rect 4504 6240 4508 6244
rect 2183 6234 2187 6238
rect 2214 6234 2218 6238
rect 2239 6234 2243 6238
rect 2298 6234 2302 6238
rect 2378 6234 2384 6238
rect 4484 6235 4488 6239
rect 4494 6235 4498 6239
rect 4504 6235 4508 6239
rect 618 6227 622 6231
rect 628 6227 632 6231
rect 638 6227 642 6231
rect 618 6222 622 6226
rect 628 6222 632 6226
rect 638 6222 642 6226
rect 618 6217 622 6221
rect 628 6217 632 6221
rect 638 6217 642 6221
rect 618 6212 622 6216
rect 628 6212 632 6216
rect 638 6212 642 6216
rect 664 6227 668 6231
rect 674 6227 678 6231
rect 684 6227 688 6231
rect 1217 6227 1221 6231
rect 1245 6227 1249 6231
rect 1260 6227 1264 6231
rect 1294 6227 1298 6231
rect 1317 6227 1321 6231
rect 1335 6227 1339 6231
rect 1353 6227 1357 6231
rect 1367 6227 1371 6231
rect 1445 6227 1451 6231
rect 2162 6227 2166 6231
rect 2190 6227 2194 6231
rect 2205 6227 2209 6231
rect 2239 6227 2243 6231
rect 2262 6227 2266 6231
rect 2280 6227 2284 6231
rect 2298 6227 2302 6231
rect 2312 6227 2316 6231
rect 2390 6227 2396 6231
rect 4484 6230 4488 6234
rect 4494 6230 4498 6234
rect 4504 6230 4508 6234
rect 664 6222 668 6226
rect 674 6222 678 6226
rect 684 6222 688 6226
rect 664 6217 668 6221
rect 674 6217 678 6221
rect 684 6217 688 6221
rect 664 6212 668 6216
rect 674 6212 678 6216
rect 684 6212 688 6216
rect 1058 6204 1062 6208
rect 618 6196 622 6200
rect 628 6196 632 6200
rect 638 6196 642 6200
rect 618 6191 622 6195
rect 628 6191 632 6195
rect 638 6191 642 6195
rect 618 6186 622 6190
rect 628 6186 632 6190
rect 638 6186 642 6190
rect 618 6181 622 6185
rect 628 6181 632 6185
rect 638 6181 642 6185
rect 664 6196 668 6200
rect 674 6196 678 6200
rect 684 6196 688 6200
rect 664 6191 668 6195
rect 674 6191 678 6195
rect 684 6191 688 6195
rect 1071 6196 1075 6200
rect 1019 6190 1023 6194
rect 664 6186 668 6190
rect 674 6186 678 6190
rect 684 6186 688 6190
rect 664 6181 668 6185
rect 674 6181 678 6185
rect 684 6181 688 6185
rect 1040 6186 1044 6194
rect 1163 6204 1167 6208
rect 1238 6220 1242 6224
rect 1269 6220 1273 6224
rect 1294 6220 1298 6224
rect 1353 6220 1357 6224
rect 1433 6220 1439 6224
rect 1238 6213 1242 6217
rect 1285 6212 1292 6216
rect 1310 6213 1314 6217
rect 1353 6212 1357 6216
rect 1217 6208 1221 6212
rect 1245 6208 1249 6212
rect 1260 6208 1264 6212
rect 1317 6208 1321 6212
rect 1335 6208 1339 6212
rect 1367 6208 1371 6212
rect 1122 6191 1126 6195
rect 1176 6196 1180 6200
rect 1079 6182 1083 6186
rect 1094 6182 1098 6186
rect 1048 6168 1052 6172
rect 1145 6186 1149 6194
rect 1208 6195 1212 6199
rect 1220 6195 1224 6199
rect 1228 6194 1232 6198
rect 1250 6195 1254 6199
rect 1263 6194 1267 6198
rect 1282 6194 1286 6198
rect 1301 6193 1305 6197
rect 1320 6197 1324 6201
rect 1340 6194 1344 6198
rect 2003 6204 2007 6208
rect 1373 6195 1377 6199
rect 2016 6196 2020 6200
rect 1964 6190 1968 6194
rect 1217 6178 1221 6182
rect 1224 6175 1228 6179
rect 1244 6178 1248 6182
rect 1260 6178 1264 6182
rect 1270 6175 1274 6179
rect 1295 6175 1299 6179
rect 1317 6178 1321 6182
rect 1335 6178 1339 6182
rect 1342 6175 1346 6179
rect 1367 6178 1371 6182
rect 1985 6186 1989 6194
rect 2108 6204 2112 6208
rect 4484 6225 4488 6229
rect 4494 6225 4498 6229
rect 4504 6225 4508 6229
rect 4530 6240 4534 6244
rect 4540 6240 4544 6244
rect 4550 6240 4554 6244
rect 4530 6235 4534 6239
rect 4540 6235 4544 6239
rect 4550 6235 4554 6239
rect 4530 6230 4534 6234
rect 4540 6230 4544 6234
rect 4550 6230 4554 6234
rect 4530 6225 4534 6229
rect 4540 6225 4544 6229
rect 4550 6225 4554 6229
rect 2183 6220 2187 6224
rect 2214 6220 2218 6224
rect 2239 6220 2243 6224
rect 2298 6220 2302 6224
rect 2378 6220 2384 6224
rect 2183 6213 2187 6217
rect 2230 6212 2237 6216
rect 2255 6213 2259 6217
rect 2298 6212 2302 6216
rect 2162 6208 2166 6212
rect 2190 6208 2194 6212
rect 2205 6208 2209 6212
rect 2262 6208 2266 6212
rect 2280 6208 2284 6212
rect 2312 6208 2316 6212
rect 2067 6191 2071 6195
rect 2121 6196 2125 6200
rect 1153 6168 1157 6172
rect 1223 6168 1227 6172
rect 1288 6168 1292 6172
rect 1310 6168 1314 6172
rect 1341 6168 1345 6172
rect 1357 6168 1361 6172
rect 1421 6168 1427 6172
rect 2024 6182 2028 6186
rect 2039 6182 2043 6186
rect 1993 6168 1997 6172
rect 2090 6186 2094 6194
rect 2153 6195 2157 6199
rect 2165 6195 2169 6199
rect 2173 6194 2177 6198
rect 2195 6195 2199 6199
rect 2208 6194 2212 6198
rect 2227 6194 2231 6198
rect 2246 6193 2250 6197
rect 2265 6197 2269 6201
rect 2285 6194 2289 6198
rect 2318 6195 2322 6199
rect 2162 6178 2166 6182
rect 2169 6175 2173 6179
rect 2189 6178 2193 6182
rect 2205 6178 2209 6182
rect 2215 6175 2219 6179
rect 2240 6175 2244 6179
rect 2262 6178 2266 6182
rect 2280 6178 2284 6182
rect 2287 6175 2291 6179
rect 2312 6178 2316 6182
rect 2098 6168 2102 6172
rect 2168 6168 2172 6172
rect 2233 6168 2237 6172
rect 2255 6168 2259 6172
rect 2286 6168 2290 6172
rect 2302 6168 2306 6172
rect 2366 6168 2372 6172
rect 1216 6161 1220 6165
rect 1244 6161 1248 6165
rect 1261 6161 1265 6165
rect 1317 6161 1321 6165
rect 1334 6161 1338 6165
rect 1368 6161 1372 6165
rect 1457 6161 1463 6165
rect 2161 6161 2165 6165
rect 2189 6161 2193 6165
rect 2206 6161 2210 6165
rect 2262 6161 2266 6165
rect 2279 6161 2283 6165
rect 2313 6161 2317 6165
rect 2402 6161 2408 6165
rect 1082 6148 1086 6152
rect 1163 6148 1167 6152
rect 1223 6154 1227 6158
rect 1288 6154 1292 6158
rect 1310 6154 1314 6158
rect 1341 6154 1345 6158
rect 1357 6154 1361 6158
rect 1409 6151 1415 6155
rect 1615 6151 1619 6155
rect 1666 6151 1670 6155
rect 1716 6151 1720 6155
rect 1217 6144 1221 6148
rect 1224 6147 1228 6151
rect 1244 6144 1248 6148
rect 1260 6144 1264 6148
rect 1270 6147 1274 6151
rect 1295 6147 1299 6151
rect 1317 6144 1321 6148
rect 1335 6144 1339 6148
rect 1342 6147 1346 6151
rect 2027 6148 2031 6152
rect 1367 6144 1371 6148
rect 1445 6144 1451 6148
rect 1064 6128 1068 6132
rect 1093 6127 1097 6131
rect 1145 6128 1149 6132
rect 1173 6127 1177 6131
rect 1208 6127 1212 6131
rect 1220 6127 1224 6131
rect 1228 6128 1232 6132
rect 1072 6112 1076 6116
rect 1153 6112 1157 6116
rect 1250 6127 1254 6131
rect 1263 6128 1267 6132
rect 1282 6128 1286 6132
rect 1301 6129 1305 6133
rect 1320 6125 1324 6129
rect 1340 6128 1344 6132
rect 1615 6135 1619 6139
rect 1652 6137 1656 6141
rect 1672 6137 1676 6141
rect 1716 6137 1720 6141
rect 2108 6148 2112 6152
rect 2168 6154 2172 6158
rect 2233 6154 2237 6158
rect 2255 6154 2259 6158
rect 2286 6154 2290 6158
rect 2302 6154 2306 6158
rect 2354 6151 2360 6155
rect 2560 6151 2564 6155
rect 2611 6151 2615 6155
rect 2661 6151 2665 6155
rect 2162 6144 2166 6148
rect 2169 6147 2173 6151
rect 2189 6144 2193 6148
rect 2205 6144 2209 6148
rect 2215 6147 2219 6151
rect 2240 6147 2244 6151
rect 2262 6144 2266 6148
rect 2280 6144 2284 6148
rect 2287 6147 2291 6151
rect 2312 6144 2316 6148
rect 2390 6144 2396 6148
rect 1372 6126 1376 6130
rect 1622 6124 1626 6128
rect 1638 6122 1642 6128
rect 1659 6124 1663 6128
rect 2009 6128 2013 6132
rect 1680 6124 1684 6128
rect 1696 6122 1700 6128
rect 1672 6118 1676 6122
rect 1717 6124 1721 6128
rect 1733 6124 1737 6128
rect 2038 6127 2042 6131
rect 2090 6128 2094 6132
rect 2118 6127 2122 6131
rect 2153 6127 2157 6131
rect 2165 6127 2169 6131
rect 2173 6128 2177 6132
rect 1217 6114 1221 6118
rect 1245 6114 1249 6118
rect 1260 6114 1264 6118
rect 1317 6114 1321 6118
rect 1335 6114 1339 6118
rect 1367 6114 1371 6118
rect 1600 6114 1604 6118
rect 1238 6109 1242 6113
rect 1285 6110 1292 6114
rect 1310 6109 1314 6113
rect 1353 6110 1357 6114
rect 1622 6109 1626 6115
rect 1659 6109 1663 6115
rect 1238 6102 1242 6106
rect 1269 6102 1273 6106
rect 1294 6102 1298 6106
rect 1353 6102 1357 6106
rect 1433 6102 1439 6106
rect 1638 6105 1642 6109
rect 1672 6109 1676 6113
rect 1680 6109 1684 6115
rect 1717 6109 1721 6115
rect 1733 6109 1737 6115
rect 2017 6112 2021 6116
rect 1696 6105 1700 6109
rect 1217 6095 1221 6099
rect 1245 6095 1249 6099
rect 1260 6095 1264 6099
rect 1294 6095 1298 6099
rect 1317 6095 1321 6099
rect 1335 6095 1339 6099
rect 1353 6095 1357 6099
rect 1367 6095 1371 6099
rect 1445 6095 1451 6099
rect 1082 6072 1086 6076
rect 1095 6064 1099 6068
rect 1037 6058 1041 6062
rect 1064 6054 1068 6062
rect 1163 6072 1167 6076
rect 1176 6064 1180 6068
rect 1122 6058 1126 6062
rect 1103 6050 1107 6054
rect 1118 6050 1122 6054
rect 1072 6036 1076 6040
rect 1145 6054 1149 6062
rect 1238 6088 1242 6092
rect 1269 6088 1273 6092
rect 1294 6088 1298 6092
rect 1353 6088 1357 6092
rect 1433 6088 1439 6092
rect 1615 6094 1619 6098
rect 1665 6094 1669 6098
rect 1718 6094 1722 6098
rect 2098 6112 2102 6116
rect 2195 6127 2199 6131
rect 2208 6128 2212 6132
rect 2227 6128 2231 6132
rect 2246 6129 2250 6133
rect 2265 6125 2269 6129
rect 2285 6128 2289 6132
rect 2560 6135 2564 6139
rect 2597 6137 2601 6141
rect 2617 6137 2621 6141
rect 2661 6137 2665 6141
rect 2317 6126 2321 6130
rect 2567 6124 2571 6128
rect 2583 6122 2587 6128
rect 2604 6124 2608 6128
rect 2625 6124 2629 6128
rect 2641 6122 2645 6128
rect 2617 6118 2621 6122
rect 2662 6124 2666 6128
rect 2678 6124 2682 6128
rect 2162 6114 2166 6118
rect 2190 6114 2194 6118
rect 2205 6114 2209 6118
rect 2262 6114 2266 6118
rect 2280 6114 2284 6118
rect 2312 6114 2316 6118
rect 2545 6114 2549 6118
rect 2183 6109 2187 6113
rect 2230 6110 2237 6114
rect 2255 6109 2259 6113
rect 2298 6110 2302 6114
rect 2567 6109 2571 6115
rect 2604 6109 2608 6115
rect 2183 6102 2187 6106
rect 2214 6102 2218 6106
rect 2239 6102 2243 6106
rect 2298 6102 2302 6106
rect 2378 6102 2384 6106
rect 2583 6105 2587 6109
rect 2617 6109 2621 6113
rect 2625 6109 2629 6115
rect 2662 6109 2666 6115
rect 2678 6109 2682 6115
rect 2641 6105 2645 6109
rect 2162 6095 2166 6099
rect 2190 6095 2194 6099
rect 2205 6095 2209 6099
rect 2239 6095 2243 6099
rect 2262 6095 2266 6099
rect 2280 6095 2284 6099
rect 2298 6095 2302 6099
rect 2312 6095 2316 6099
rect 2390 6095 2396 6099
rect 1457 6087 1463 6091
rect 1238 6081 1242 6085
rect 1285 6080 1292 6084
rect 1310 6081 1314 6085
rect 1353 6080 1357 6084
rect 1397 6080 1403 6084
rect 1615 6080 1619 6084
rect 1651 6080 1655 6084
rect 1718 6080 1722 6084
rect 1217 6076 1221 6080
rect 1245 6076 1249 6080
rect 1260 6076 1264 6080
rect 1317 6076 1321 6080
rect 1335 6076 1339 6080
rect 1367 6076 1371 6080
rect 1208 6063 1212 6067
rect 1220 6063 1224 6067
rect 1228 6062 1232 6066
rect 1250 6063 1254 6067
rect 1263 6062 1267 6066
rect 1282 6062 1286 6066
rect 1184 6050 1188 6054
rect 1199 6050 1203 6054
rect 1301 6061 1305 6065
rect 1320 6065 1324 6069
rect 1340 6062 1344 6066
rect 1584 6072 1588 6076
rect 1725 6072 1729 6076
rect 2027 6072 2031 6076
rect 1584 6063 1588 6067
rect 1608 6063 1612 6067
rect 1733 6065 1737 6069
rect 2040 6064 2044 6068
rect 1600 6056 1604 6060
rect 1982 6058 1986 6062
rect 1153 6036 1157 6040
rect 1217 6046 1221 6050
rect 1224 6043 1228 6047
rect 1244 6046 1248 6050
rect 1260 6046 1264 6050
rect 1270 6043 1274 6047
rect 1295 6043 1299 6047
rect 1317 6046 1321 6050
rect 1335 6046 1339 6050
rect 1342 6043 1346 6047
rect 1367 6046 1371 6050
rect 1409 6049 1415 6053
rect 1617 6049 1621 6053
rect 1667 6049 1671 6053
rect 1718 6049 1722 6053
rect 1445 6042 1451 6046
rect 2009 6054 2013 6062
rect 2108 6072 2112 6076
rect 2121 6064 2125 6068
rect 2067 6058 2071 6062
rect 1223 6036 1227 6040
rect 1288 6036 1292 6040
rect 1310 6036 1314 6040
rect 1341 6036 1345 6040
rect 1421 6036 1427 6040
rect 1216 6029 1220 6033
rect 1244 6029 1248 6033
rect 1261 6029 1265 6033
rect 1317 6029 1321 6033
rect 1334 6029 1338 6033
rect 1368 6029 1372 6033
rect 1457 6029 1463 6033
rect 1617 6035 1621 6039
rect 1661 6035 1665 6039
rect 1681 6035 1685 6039
rect 1718 6033 1722 6037
rect 2048 6050 2052 6054
rect 2063 6050 2067 6054
rect 2017 6036 2021 6040
rect 2090 6054 2094 6062
rect 2183 6088 2187 6092
rect 2214 6088 2218 6092
rect 2239 6088 2243 6092
rect 2298 6088 2302 6092
rect 2378 6088 2384 6092
rect 2560 6094 2564 6098
rect 2610 6094 2614 6098
rect 2663 6094 2667 6098
rect 2402 6087 2408 6091
rect 2183 6081 2187 6085
rect 2230 6080 2237 6084
rect 2255 6081 2259 6085
rect 2298 6080 2302 6084
rect 2342 6080 2348 6084
rect 2560 6080 2564 6084
rect 2596 6080 2600 6084
rect 2663 6080 2667 6084
rect 2162 6076 2166 6080
rect 2190 6076 2194 6080
rect 2205 6076 2209 6080
rect 2262 6076 2266 6080
rect 2280 6076 2284 6080
rect 2312 6076 2316 6080
rect 2153 6063 2157 6067
rect 2165 6063 2169 6067
rect 2173 6062 2177 6066
rect 2195 6063 2199 6067
rect 2208 6062 2212 6066
rect 2227 6062 2231 6066
rect 2129 6050 2133 6054
rect 2144 6050 2148 6054
rect 2246 6061 2250 6065
rect 2265 6065 2269 6069
rect 2285 6062 2289 6066
rect 2529 6072 2533 6076
rect 2670 6072 2674 6076
rect 2529 6063 2533 6067
rect 2553 6063 2557 6067
rect 2678 6065 2682 6069
rect 2545 6056 2549 6060
rect 2098 6036 2102 6040
rect 2162 6046 2166 6050
rect 2169 6043 2173 6047
rect 2189 6046 2193 6050
rect 2205 6046 2209 6050
rect 2215 6043 2219 6047
rect 2240 6043 2244 6047
rect 2262 6046 2266 6050
rect 2280 6046 2284 6050
rect 2287 6043 2291 6047
rect 2312 6046 2316 6050
rect 2354 6049 2360 6053
rect 2562 6049 2566 6053
rect 2612 6049 2616 6053
rect 2663 6049 2667 6053
rect 2390 6042 2396 6046
rect 2168 6036 2172 6040
rect 2233 6036 2237 6040
rect 2255 6036 2259 6040
rect 2286 6036 2290 6040
rect 2366 6036 2372 6040
rect 1600 6022 1604 6026
rect 1616 6022 1620 6026
rect 869 6016 873 6020
rect 919 6016 923 6020
rect 970 6016 974 6020
rect 1001 6016 1005 6020
rect 1051 6016 1055 6020
rect 1102 6016 1106 6020
rect 1133 6016 1137 6020
rect 1183 6016 1187 6020
rect 1234 6016 1238 6020
rect 1265 6016 1269 6020
rect 1315 6016 1319 6020
rect 1366 6016 1370 6020
rect 1409 6016 1415 6020
rect 1637 6020 1641 6026
rect 1653 6022 1657 6026
rect 2161 6029 2165 6033
rect 2189 6029 2193 6033
rect 2206 6029 2210 6033
rect 2262 6029 2266 6033
rect 2279 6029 2283 6033
rect 2313 6029 2317 6033
rect 2402 6029 2408 6033
rect 2562 6035 2566 6039
rect 2606 6035 2610 6039
rect 2626 6035 2630 6039
rect 2663 6033 2667 6037
rect 1674 6022 1678 6026
rect 1661 6016 1665 6020
rect 1695 6020 1699 6026
rect 1711 6022 1715 6026
rect 2545 6022 2549 6026
rect 2561 6022 2565 6026
rect 1814 6016 1818 6020
rect 1864 6016 1868 6020
rect 1915 6016 1919 6020
rect 1946 6016 1950 6020
rect 1996 6016 2000 6020
rect 2047 6016 2051 6020
rect 2078 6016 2082 6020
rect 2128 6016 2132 6020
rect 2179 6016 2183 6020
rect 2210 6016 2214 6020
rect 2260 6016 2264 6020
rect 2311 6016 2315 6020
rect 2354 6016 2360 6020
rect 1445 6009 1451 6013
rect 852 5997 856 6001
rect 869 6002 873 6006
rect 913 6002 917 6006
rect 933 6002 937 6006
rect 970 6000 974 6004
rect 852 5989 856 5993
rect 868 5989 872 5993
rect 889 5987 893 5993
rect 905 5989 909 5993
rect 984 5997 988 6001
rect 1001 6002 1005 6006
rect 1045 6002 1049 6006
rect 1065 6002 1069 6006
rect 1102 6000 1106 6004
rect 1133 6002 1137 6006
rect 1177 6002 1181 6006
rect 1197 6002 1201 6006
rect 1234 6000 1238 6004
rect 1265 6002 1269 6006
rect 1309 6002 1313 6006
rect 1329 6002 1333 6006
rect 1366 6000 1370 6004
rect 1600 6007 1604 6013
rect 1616 6007 1620 6013
rect 1653 6007 1657 6013
rect 1637 6003 1641 6007
rect 1661 6007 1665 6011
rect 1674 6007 1678 6013
rect 1711 6007 1715 6013
rect 1733 6012 1737 6016
rect 2582 6020 2586 6026
rect 2598 6022 2602 6026
rect 2619 6022 2623 6026
rect 2606 6016 2610 6020
rect 2640 6020 2644 6026
rect 2656 6022 2660 6026
rect 2390 6009 2396 6013
rect 1695 6003 1699 6007
rect 926 5989 930 5993
rect 913 5983 917 5987
rect 947 5987 951 5993
rect 963 5989 967 5993
rect 984 5989 988 5993
rect 1000 5989 1004 5993
rect 852 5974 856 5978
rect 868 5974 872 5980
rect 905 5974 909 5980
rect 889 5970 893 5974
rect 913 5974 917 5978
rect 926 5974 930 5980
rect 963 5974 967 5980
rect 976 5979 980 5983
rect 1021 5987 1025 5993
rect 1037 5989 1041 5993
rect 1058 5989 1062 5993
rect 1045 5983 1049 5987
rect 1079 5987 1083 5993
rect 1095 5989 1099 5993
rect 1116 5989 1120 5993
rect 1132 5989 1136 5993
rect 984 5974 988 5978
rect 1000 5974 1004 5980
rect 1037 5974 1041 5980
rect 947 5970 951 5974
rect 1021 5970 1025 5974
rect 1045 5974 1049 5978
rect 1058 5974 1062 5980
rect 1095 5974 1099 5980
rect 1108 5979 1112 5983
rect 1153 5987 1157 5993
rect 1169 5989 1173 5993
rect 1190 5989 1194 5993
rect 1177 5983 1181 5987
rect 1211 5987 1215 5993
rect 1227 5989 1231 5993
rect 1248 5989 1252 5993
rect 1264 5989 1268 5993
rect 1116 5974 1120 5978
rect 1132 5974 1136 5980
rect 1169 5974 1173 5980
rect 1079 5970 1083 5974
rect 1153 5970 1157 5974
rect 1177 5974 1181 5978
rect 1190 5974 1194 5980
rect 1227 5974 1231 5980
rect 1240 5979 1244 5983
rect 1285 5987 1289 5993
rect 1301 5989 1305 5993
rect 1322 5989 1326 5993
rect 1309 5983 1313 5987
rect 1343 5987 1347 5993
rect 1359 5989 1363 5993
rect 1615 5992 1619 5996
rect 1668 5992 1672 5996
rect 1718 5992 1722 5996
rect 1797 5997 1801 6001
rect 1814 6002 1818 6006
rect 1858 6002 1862 6006
rect 1878 6002 1882 6006
rect 1915 6000 1919 6004
rect 1797 5989 1801 5993
rect 1813 5989 1817 5993
rect 1457 5985 1463 5989
rect 1248 5974 1252 5978
rect 1264 5974 1268 5980
rect 1301 5974 1305 5980
rect 1211 5970 1215 5974
rect 1285 5970 1289 5974
rect 1309 5974 1313 5978
rect 1322 5974 1326 5980
rect 1359 5974 1363 5980
rect 1372 5979 1376 5983
rect 1834 5987 1838 5993
rect 1850 5989 1854 5993
rect 1929 5997 1933 6001
rect 1946 6002 1950 6006
rect 1990 6002 1994 6006
rect 2010 6002 2014 6006
rect 2047 6000 2051 6004
rect 2078 6002 2082 6006
rect 2122 6002 2126 6006
rect 2142 6002 2146 6006
rect 2179 6000 2183 6004
rect 2210 6002 2214 6006
rect 2254 6002 2258 6006
rect 2274 6002 2278 6006
rect 2311 6000 2315 6004
rect 2545 6007 2549 6013
rect 2561 6007 2565 6013
rect 2598 6007 2602 6013
rect 2582 6003 2586 6007
rect 2606 6007 2610 6011
rect 2619 6007 2623 6013
rect 2656 6007 2660 6013
rect 2678 6012 2682 6016
rect 2640 6003 2644 6007
rect 1871 5989 1875 5993
rect 1858 5983 1862 5987
rect 1892 5987 1896 5993
rect 1908 5989 1912 5993
rect 1929 5989 1933 5993
rect 1945 5989 1949 5993
rect 1397 5978 1403 5982
rect 1615 5978 1619 5982
rect 1682 5978 1686 5982
rect 1718 5978 1722 5982
rect 1797 5974 1801 5978
rect 1813 5974 1817 5980
rect 1850 5974 1854 5980
rect 1343 5970 1347 5974
rect 1834 5970 1838 5974
rect 1858 5974 1862 5978
rect 1871 5974 1875 5980
rect 1908 5974 1912 5980
rect 1921 5979 1925 5983
rect 1966 5987 1970 5993
rect 1982 5989 1986 5993
rect 2003 5989 2007 5993
rect 1990 5983 1994 5987
rect 2024 5987 2028 5993
rect 2040 5989 2044 5993
rect 2061 5989 2065 5993
rect 2077 5989 2081 5993
rect 1929 5974 1933 5978
rect 1945 5974 1949 5980
rect 1982 5974 1986 5980
rect 1892 5970 1896 5974
rect 1966 5970 1970 5974
rect 1990 5974 1994 5978
rect 2003 5974 2007 5980
rect 2040 5974 2044 5980
rect 2053 5979 2057 5983
rect 2098 5987 2102 5993
rect 2114 5989 2118 5993
rect 2135 5989 2139 5993
rect 2122 5983 2126 5987
rect 2156 5987 2160 5993
rect 2172 5989 2176 5993
rect 2193 5989 2197 5993
rect 2209 5989 2213 5993
rect 2061 5974 2065 5978
rect 2077 5974 2081 5980
rect 2114 5974 2118 5980
rect 2024 5970 2028 5974
rect 2098 5970 2102 5974
rect 2122 5974 2126 5978
rect 2135 5974 2139 5980
rect 2172 5974 2176 5980
rect 2185 5979 2189 5983
rect 2230 5987 2234 5993
rect 2246 5989 2250 5993
rect 2267 5989 2271 5993
rect 2254 5983 2258 5987
rect 2288 5987 2292 5993
rect 2304 5989 2308 5993
rect 2560 5992 2564 5996
rect 2613 5992 2617 5996
rect 2663 5992 2667 5996
rect 2402 5985 2408 5989
rect 2193 5974 2197 5978
rect 2209 5974 2213 5980
rect 2246 5974 2250 5980
rect 2156 5970 2160 5974
rect 2230 5970 2234 5974
rect 2254 5974 2258 5978
rect 2267 5974 2271 5980
rect 2304 5974 2308 5980
rect 2317 5979 2321 5983
rect 2342 5978 2348 5982
rect 2560 5978 2564 5982
rect 2627 5978 2631 5982
rect 2663 5978 2667 5982
rect 2288 5970 2292 5974
rect 867 5959 871 5963
rect 920 5959 924 5963
rect 970 5959 974 5963
rect 999 5959 1003 5963
rect 1052 5959 1056 5963
rect 1102 5959 1106 5963
rect 1131 5959 1135 5963
rect 1184 5959 1188 5963
rect 1234 5959 1238 5963
rect 1263 5959 1267 5963
rect 1316 5959 1320 5963
rect 1366 5959 1370 5963
rect 1812 5959 1816 5963
rect 1865 5959 1869 5963
rect 1915 5959 1919 5963
rect 1944 5959 1948 5963
rect 1997 5959 2001 5963
rect 2047 5959 2051 5963
rect 2076 5959 2080 5963
rect 2129 5959 2133 5963
rect 2179 5959 2183 5963
rect 2208 5959 2212 5963
rect 2261 5959 2265 5963
rect 2311 5959 2315 5963
rect 1457 5952 1463 5956
rect 2402 5952 2408 5956
rect 867 5945 871 5949
rect 934 5945 938 5949
rect 970 5945 974 5949
rect 999 5945 1003 5949
rect 1066 5945 1070 5949
rect 1102 5945 1106 5949
rect 1131 5945 1135 5949
rect 1198 5945 1202 5949
rect 1234 5945 1238 5949
rect 1263 5945 1267 5949
rect 1330 5945 1334 5949
rect 1366 5945 1370 5949
rect 1397 5945 1403 5949
rect 1812 5945 1816 5949
rect 1879 5945 1883 5949
rect 1915 5945 1919 5949
rect 1944 5945 1948 5949
rect 2011 5945 2015 5949
rect 2047 5945 2051 5949
rect 2076 5945 2080 5949
rect 2143 5945 2147 5949
rect 2179 5945 2183 5949
rect 2208 5945 2212 5949
rect 2275 5945 2279 5949
rect 2311 5945 2315 5949
rect 2342 5945 2348 5949
rect 1409 5937 1415 5941
rect 1485 5937 1489 5941
rect 1535 5937 1539 5941
rect 1586 5937 1590 5941
rect 1617 5937 1621 5941
rect 1667 5937 1671 5941
rect 1718 5937 1722 5941
rect 1749 5937 1753 5941
rect 1799 5937 1803 5941
rect 1850 5937 1854 5941
rect 2354 5937 2360 5941
rect 2430 5937 2434 5941
rect 2480 5937 2484 5941
rect 2531 5937 2535 5941
rect 2562 5937 2566 5941
rect 2612 5937 2616 5941
rect 2663 5937 2667 5941
rect 2694 5937 2698 5941
rect 2744 5937 2748 5941
rect 2795 5937 2799 5941
rect 1445 5930 1451 5934
rect 2390 5930 2396 5934
rect 4484 5931 4488 5935
rect 4494 5931 4498 5935
rect 4504 5931 4508 5935
rect 1485 5923 1489 5927
rect 1529 5923 1533 5927
rect 1549 5923 1553 5927
rect 1586 5921 1590 5925
rect 1617 5923 1621 5927
rect 1661 5923 1665 5927
rect 1681 5923 1685 5927
rect 1718 5921 1722 5925
rect 1749 5923 1753 5927
rect 1793 5923 1797 5927
rect 1813 5923 1817 5927
rect 1850 5921 1854 5925
rect 2430 5923 2434 5927
rect 2474 5923 2478 5927
rect 2494 5923 2498 5927
rect 2531 5921 2535 5925
rect 2562 5923 2566 5927
rect 2606 5923 2610 5927
rect 2626 5923 2630 5927
rect 2663 5921 2667 5925
rect 2694 5923 2698 5927
rect 2738 5923 2742 5927
rect 2758 5923 2762 5927
rect 2795 5921 2799 5925
rect 1468 5910 1472 5914
rect 1484 5910 1488 5914
rect 1505 5908 1509 5914
rect 1521 5910 1525 5914
rect 1542 5910 1546 5914
rect 1529 5904 1533 5908
rect 1563 5908 1567 5914
rect 1579 5910 1583 5914
rect 1600 5910 1604 5914
rect 1616 5910 1620 5914
rect 1637 5908 1641 5914
rect 1653 5910 1657 5914
rect 1674 5910 1678 5914
rect 1661 5904 1665 5908
rect 1695 5908 1699 5914
rect 1711 5910 1715 5914
rect 1732 5910 1736 5914
rect 1748 5910 1752 5914
rect 1769 5908 1773 5914
rect 1785 5910 1789 5914
rect 1806 5910 1810 5914
rect 1793 5904 1797 5908
rect 1827 5908 1831 5914
rect 1843 5910 1847 5914
rect 2413 5910 2417 5914
rect 2429 5910 2433 5914
rect 1468 5895 1472 5899
rect 1484 5895 1488 5901
rect 1521 5895 1525 5901
rect 618 5887 622 5891
rect 628 5887 632 5891
rect 638 5887 642 5891
rect 618 5882 622 5886
rect 628 5882 632 5886
rect 638 5882 642 5886
rect 618 5877 622 5881
rect 628 5877 632 5881
rect 638 5877 642 5881
rect 618 5872 622 5876
rect 628 5872 632 5876
rect 638 5872 642 5876
rect 664 5887 668 5891
rect 674 5887 678 5891
rect 684 5887 688 5891
rect 1505 5891 1509 5895
rect 1529 5895 1533 5899
rect 1542 5895 1546 5901
rect 1579 5895 1583 5901
rect 1600 5895 1604 5901
rect 1616 5895 1620 5901
rect 1653 5895 1657 5901
rect 1563 5891 1567 5895
rect 1637 5891 1641 5895
rect 1661 5895 1665 5899
rect 1674 5895 1678 5901
rect 1711 5895 1715 5901
rect 1732 5895 1736 5901
rect 1748 5895 1752 5901
rect 1785 5895 1789 5901
rect 1695 5891 1699 5895
rect 1769 5891 1773 5895
rect 1793 5895 1797 5899
rect 1806 5895 1810 5901
rect 1843 5895 1847 5901
rect 1856 5900 1860 5904
rect 2450 5908 2454 5914
rect 2466 5910 2470 5914
rect 2487 5910 2491 5914
rect 2474 5904 2478 5908
rect 2508 5908 2512 5914
rect 2524 5910 2528 5914
rect 2545 5910 2549 5914
rect 2561 5910 2565 5914
rect 2582 5908 2586 5914
rect 2598 5910 2602 5914
rect 2619 5910 2623 5914
rect 2606 5904 2610 5908
rect 2640 5908 2644 5914
rect 2656 5910 2660 5914
rect 2677 5910 2681 5914
rect 2693 5910 2697 5914
rect 2714 5908 2718 5914
rect 2730 5910 2734 5914
rect 4484 5926 4488 5930
rect 4494 5926 4498 5930
rect 4504 5926 4508 5930
rect 4484 5921 4488 5925
rect 4494 5921 4498 5925
rect 4504 5921 4508 5925
rect 4484 5916 4488 5920
rect 4494 5916 4498 5920
rect 4504 5916 4508 5920
rect 4530 5931 4534 5935
rect 4540 5931 4544 5935
rect 4550 5931 4554 5935
rect 4530 5926 4534 5930
rect 4540 5926 4544 5930
rect 4550 5926 4554 5930
rect 4530 5921 4534 5925
rect 4540 5921 4544 5925
rect 4550 5921 4554 5925
rect 4530 5916 4534 5920
rect 4540 5916 4544 5920
rect 4550 5916 4554 5920
rect 2751 5910 2755 5914
rect 2738 5904 2742 5908
rect 2772 5908 2776 5914
rect 2788 5910 2792 5914
rect 2413 5895 2417 5899
rect 2429 5895 2433 5901
rect 2466 5895 2470 5901
rect 1827 5891 1831 5895
rect 2450 5891 2454 5895
rect 2474 5895 2478 5899
rect 2487 5895 2491 5901
rect 2524 5895 2528 5901
rect 2545 5895 2549 5901
rect 2561 5895 2565 5901
rect 2598 5895 2602 5901
rect 2508 5891 2512 5895
rect 2582 5891 2586 5895
rect 2606 5895 2610 5899
rect 2619 5895 2623 5901
rect 2656 5895 2660 5901
rect 2677 5895 2681 5901
rect 2693 5895 2697 5901
rect 2730 5895 2734 5901
rect 2640 5891 2644 5895
rect 2714 5891 2718 5895
rect 2738 5895 2742 5899
rect 2751 5895 2755 5901
rect 2788 5895 2792 5901
rect 2801 5900 2805 5904
rect 2772 5891 2776 5895
rect 664 5882 668 5886
rect 674 5882 678 5886
rect 684 5882 688 5886
rect 664 5877 668 5881
rect 674 5877 678 5881
rect 684 5877 688 5881
rect 1483 5880 1487 5884
rect 1536 5880 1540 5884
rect 1586 5880 1590 5884
rect 1615 5880 1619 5884
rect 1668 5880 1672 5884
rect 1718 5880 1722 5884
rect 1747 5880 1751 5884
rect 1800 5880 1804 5884
rect 1850 5880 1854 5884
rect 2428 5880 2432 5884
rect 2481 5880 2485 5884
rect 2531 5880 2535 5884
rect 2560 5880 2564 5884
rect 2613 5880 2617 5884
rect 2663 5880 2667 5884
rect 2692 5880 2696 5884
rect 2745 5880 2749 5884
rect 2795 5880 2799 5884
rect 664 5872 668 5876
rect 674 5872 678 5876
rect 684 5872 688 5876
rect 1457 5873 1463 5877
rect 2402 5873 2408 5877
rect 1397 5866 1403 5870
rect 1483 5866 1487 5870
rect 1550 5866 1554 5870
rect 1586 5866 1590 5870
rect 1615 5866 1619 5870
rect 1682 5866 1686 5870
rect 1718 5866 1722 5870
rect 1747 5866 1751 5870
rect 1814 5866 1818 5870
rect 1850 5866 1854 5870
rect 2342 5866 2348 5870
rect 2428 5866 2432 5870
rect 2495 5866 2499 5870
rect 2531 5866 2535 5870
rect 2560 5866 2564 5870
rect 2627 5866 2631 5870
rect 2663 5866 2667 5870
rect 2692 5866 2696 5870
rect 2759 5866 2763 5870
rect 2795 5866 2799 5870
rect 1600 5859 1604 5863
rect 1624 5859 1628 5863
rect 1732 5859 1736 5863
rect 2545 5859 2549 5863
rect 2569 5859 2573 5863
rect 2677 5859 2681 5863
rect 1608 5852 1612 5856
rect 1592 5848 1596 5852
rect 1624 5848 1628 5852
rect 2553 5852 2557 5856
rect 2537 5848 2541 5852
rect 2569 5848 2573 5852
rect 1468 5844 1472 5848
rect 2413 5844 2417 5848
rect 1468 5836 1472 5840
rect 1608 5836 1612 5840
rect 2413 5836 2417 5840
rect 2553 5836 2557 5840
rect 927 5829 931 5833
rect 1592 5829 1596 5833
rect 1624 5829 1628 5833
rect 1872 5829 1876 5833
rect 2537 5829 2541 5833
rect 2569 5829 2573 5833
rect 1592 5822 1596 5826
rect 1624 5822 1628 5826
rect 1608 5818 1612 5822
rect 2537 5822 2541 5826
rect 2569 5822 2573 5826
rect 2553 5818 2557 5822
rect 1600 5811 1604 5815
rect 1624 5811 1628 5815
rect 1732 5811 1736 5815
rect 2545 5811 2549 5815
rect 2569 5811 2573 5815
rect 2677 5811 2681 5815
rect 1468 5804 1472 5808
rect 1857 5804 1861 5808
rect 2413 5804 2417 5808
rect 2802 5804 2806 5808
rect 1409 5797 1415 5801
rect 1485 5797 1489 5801
rect 1535 5797 1539 5801
rect 1586 5797 1590 5801
rect 1617 5797 1621 5801
rect 1667 5797 1671 5801
rect 1718 5797 1722 5801
rect 1749 5797 1753 5801
rect 1799 5797 1803 5801
rect 1850 5797 1854 5801
rect 2354 5797 2360 5801
rect 2430 5797 2434 5801
rect 2480 5797 2484 5801
rect 2531 5797 2535 5801
rect 2562 5797 2566 5801
rect 2612 5797 2616 5801
rect 2663 5797 2667 5801
rect 2694 5797 2698 5801
rect 2744 5797 2748 5801
rect 2795 5797 2799 5801
rect 1445 5790 1451 5794
rect 2390 5790 2396 5794
rect 1485 5783 1489 5787
rect 1529 5783 1533 5787
rect 1549 5783 1553 5787
rect 1586 5781 1590 5785
rect 1617 5783 1621 5787
rect 1661 5783 1665 5787
rect 1681 5783 1685 5787
rect 1718 5781 1722 5785
rect 1749 5783 1753 5787
rect 1793 5783 1797 5787
rect 1813 5783 1817 5787
rect 1850 5781 1854 5785
rect 2430 5783 2434 5787
rect 2474 5783 2478 5787
rect 2494 5783 2498 5787
rect 2531 5781 2535 5785
rect 2562 5783 2566 5787
rect 2606 5783 2610 5787
rect 2626 5783 2630 5787
rect 2663 5781 2667 5785
rect 2694 5783 2698 5787
rect 2738 5783 2742 5787
rect 2758 5783 2762 5787
rect 2795 5781 2799 5785
rect 966 5767 970 5771
rect 1016 5767 1020 5771
rect 1067 5767 1071 5771
rect 1409 5767 1415 5771
rect 1468 5770 1472 5774
rect 1484 5770 1488 5774
rect 1445 5760 1451 5764
rect 1505 5768 1509 5774
rect 1521 5770 1525 5774
rect 1542 5770 1546 5774
rect 1529 5764 1533 5768
rect 1563 5768 1567 5774
rect 1579 5770 1583 5774
rect 1600 5770 1604 5774
rect 1616 5770 1620 5774
rect 1637 5768 1641 5774
rect 1653 5770 1657 5774
rect 1674 5770 1678 5774
rect 1661 5764 1665 5768
rect 1695 5768 1699 5774
rect 1711 5770 1715 5774
rect 1732 5770 1736 5774
rect 1748 5770 1752 5774
rect 1769 5768 1773 5774
rect 1785 5770 1789 5774
rect 1806 5770 1810 5774
rect 1793 5764 1797 5768
rect 1827 5768 1831 5774
rect 1843 5770 1847 5774
rect 1911 5767 1915 5771
rect 1961 5767 1965 5771
rect 2012 5767 2016 5771
rect 2354 5767 2360 5771
rect 2413 5770 2417 5774
rect 2429 5770 2433 5774
rect 966 5753 970 5757
rect 1010 5753 1014 5757
rect 1030 5753 1034 5757
rect 1067 5751 1071 5755
rect 927 5743 931 5747
rect 949 5735 953 5744
rect 965 5740 969 5744
rect 986 5738 990 5744
rect 1002 5740 1006 5744
rect 1468 5755 1472 5759
rect 1484 5755 1488 5761
rect 1521 5755 1525 5761
rect 1505 5751 1509 5755
rect 1529 5755 1533 5759
rect 1542 5755 1546 5761
rect 1579 5755 1583 5761
rect 1600 5755 1604 5761
rect 1616 5755 1620 5761
rect 1653 5755 1657 5761
rect 1563 5751 1567 5755
rect 1637 5751 1641 5755
rect 1661 5755 1665 5759
rect 1674 5755 1678 5761
rect 1711 5755 1715 5761
rect 1732 5755 1736 5761
rect 1748 5755 1752 5761
rect 1785 5755 1789 5761
rect 1695 5751 1699 5755
rect 1769 5751 1773 5755
rect 1793 5755 1797 5759
rect 1806 5755 1810 5761
rect 1843 5755 1847 5761
rect 1856 5760 1860 5764
rect 2390 5760 2396 5764
rect 2450 5768 2454 5774
rect 2466 5770 2470 5774
rect 2487 5770 2491 5774
rect 2474 5764 2478 5768
rect 2508 5768 2512 5774
rect 2524 5770 2528 5774
rect 2545 5770 2549 5774
rect 2561 5770 2565 5774
rect 2582 5768 2586 5774
rect 2598 5770 2602 5774
rect 2619 5770 2623 5774
rect 2606 5764 2610 5768
rect 2640 5768 2644 5774
rect 2656 5770 2660 5774
rect 2677 5770 2681 5774
rect 2693 5770 2697 5774
rect 2714 5768 2718 5774
rect 2730 5770 2734 5774
rect 2751 5770 2755 5774
rect 2738 5764 2742 5768
rect 2772 5768 2776 5774
rect 2788 5770 2792 5774
rect 1827 5751 1831 5755
rect 1911 5753 1915 5757
rect 1955 5753 1959 5757
rect 1975 5753 1979 5757
rect 2012 5751 2016 5755
rect 1023 5740 1027 5744
rect 1010 5734 1014 5738
rect 1044 5738 1048 5744
rect 1060 5740 1064 5744
rect 1483 5740 1487 5744
rect 1536 5740 1540 5744
rect 1586 5740 1590 5744
rect 1615 5740 1619 5744
rect 1668 5740 1672 5744
rect 1718 5740 1722 5744
rect 1747 5740 1751 5744
rect 1800 5740 1804 5744
rect 1850 5740 1854 5744
rect 1872 5743 1876 5747
rect 927 5727 931 5731
rect 949 5725 953 5729
rect 965 5725 969 5731
rect 1002 5725 1006 5731
rect 986 5721 990 5725
rect 1010 5725 1014 5729
rect 1023 5725 1027 5731
rect 1060 5725 1064 5731
rect 1073 5730 1077 5734
rect 1457 5733 1463 5737
rect 1894 5735 1898 5744
rect 1910 5740 1914 5744
rect 1931 5738 1935 5744
rect 1947 5740 1951 5744
rect 2413 5755 2417 5759
rect 2429 5755 2433 5761
rect 2466 5755 2470 5761
rect 2450 5751 2454 5755
rect 2474 5755 2478 5759
rect 2487 5755 2491 5761
rect 2524 5755 2528 5761
rect 2545 5755 2549 5761
rect 2561 5755 2565 5761
rect 2598 5755 2602 5761
rect 2508 5751 2512 5755
rect 2582 5751 2586 5755
rect 2606 5755 2610 5759
rect 2619 5755 2623 5761
rect 2656 5755 2660 5761
rect 2677 5755 2681 5761
rect 2693 5755 2697 5761
rect 2730 5755 2734 5761
rect 2640 5751 2644 5755
rect 2714 5751 2718 5755
rect 2738 5755 2742 5759
rect 2751 5755 2755 5761
rect 2788 5755 2792 5761
rect 2801 5760 2805 5764
rect 2772 5751 2776 5755
rect 1968 5740 1972 5744
rect 1955 5734 1959 5738
rect 1989 5738 1993 5744
rect 2005 5740 2009 5744
rect 2428 5740 2432 5744
rect 2481 5740 2485 5744
rect 2531 5740 2535 5744
rect 2560 5740 2564 5744
rect 2613 5740 2617 5744
rect 2663 5740 2667 5744
rect 2692 5740 2696 5744
rect 2745 5740 2749 5744
rect 2795 5740 2799 5744
rect 1397 5726 1403 5730
rect 1483 5726 1487 5730
rect 1550 5726 1554 5730
rect 1586 5726 1590 5730
rect 1615 5726 1619 5730
rect 1682 5726 1686 5730
rect 1718 5726 1722 5730
rect 1747 5726 1751 5730
rect 1814 5726 1818 5730
rect 1850 5726 1854 5730
rect 1872 5727 1876 5731
rect 1894 5725 1898 5729
rect 1910 5725 1914 5731
rect 1947 5725 1951 5731
rect 1044 5721 1048 5725
rect 1468 5718 1472 5722
rect 1857 5718 1861 5722
rect 1931 5721 1935 5725
rect 1955 5725 1959 5729
rect 1968 5725 1972 5731
rect 2005 5725 2009 5731
rect 2018 5730 2022 5734
rect 2402 5733 2408 5737
rect 2342 5726 2348 5730
rect 2428 5726 2432 5730
rect 2495 5726 2499 5730
rect 2531 5726 2535 5730
rect 2560 5726 2564 5730
rect 2627 5726 2631 5730
rect 2663 5726 2667 5730
rect 2692 5726 2696 5730
rect 2759 5726 2763 5730
rect 2795 5726 2799 5730
rect 1989 5721 1993 5725
rect 2413 5718 2417 5722
rect 2802 5718 2806 5722
rect 964 5710 968 5714
rect 1017 5710 1021 5714
rect 1067 5710 1071 5714
rect 1409 5711 1415 5715
rect 1485 5711 1489 5715
rect 1535 5711 1539 5715
rect 1586 5711 1590 5715
rect 1617 5711 1621 5715
rect 1667 5711 1671 5715
rect 1718 5711 1722 5715
rect 1749 5711 1753 5715
rect 1799 5711 1803 5715
rect 1850 5711 1854 5715
rect 1081 5703 1085 5707
rect 1445 5704 1451 5708
rect 1909 5710 1913 5714
rect 1962 5710 1966 5714
rect 2012 5710 2016 5714
rect 2354 5711 2360 5715
rect 2430 5711 2434 5715
rect 2480 5711 2484 5715
rect 2531 5711 2535 5715
rect 2562 5711 2566 5715
rect 2612 5711 2616 5715
rect 2663 5711 2667 5715
rect 2694 5711 2698 5715
rect 2744 5711 2748 5715
rect 2795 5711 2799 5715
rect 964 5696 968 5700
rect 1031 5696 1035 5700
rect 1067 5696 1071 5700
rect 1397 5696 1403 5700
rect 949 5688 953 5692
rect 1074 5689 1078 5693
rect 1485 5697 1489 5701
rect 1529 5697 1533 5701
rect 1549 5697 1553 5701
rect 1586 5695 1590 5699
rect 1617 5697 1621 5701
rect 1661 5697 1665 5701
rect 1681 5697 1685 5701
rect 1718 5695 1722 5699
rect 1749 5697 1753 5701
rect 1793 5697 1797 5701
rect 1813 5697 1817 5701
rect 1850 5695 1854 5699
rect 2026 5703 2030 5707
rect 2390 5704 2396 5708
rect 1909 5696 1913 5700
rect 1976 5696 1980 5700
rect 2012 5696 2016 5700
rect 2342 5696 2348 5700
rect 966 5681 970 5685
rect 1016 5681 1020 5685
rect 1067 5681 1071 5685
rect 1409 5681 1415 5685
rect 1468 5684 1472 5688
rect 1484 5684 1488 5688
rect 1445 5674 1451 5678
rect 1505 5682 1509 5688
rect 1521 5684 1525 5688
rect 1542 5684 1546 5688
rect 1529 5678 1533 5682
rect 1563 5682 1567 5688
rect 1579 5684 1583 5688
rect 1600 5684 1604 5688
rect 1616 5684 1620 5688
rect 1637 5682 1641 5688
rect 1653 5684 1657 5688
rect 1674 5684 1678 5688
rect 1661 5678 1665 5682
rect 1695 5682 1699 5688
rect 1711 5684 1715 5688
rect 1732 5684 1736 5688
rect 1748 5684 1752 5688
rect 1769 5682 1773 5688
rect 1785 5684 1789 5688
rect 1894 5688 1898 5692
rect 2019 5689 2023 5693
rect 2430 5697 2434 5701
rect 2474 5697 2478 5701
rect 2494 5697 2498 5701
rect 2531 5695 2535 5699
rect 2562 5697 2566 5701
rect 2606 5697 2610 5701
rect 2626 5697 2630 5701
rect 2663 5695 2667 5699
rect 2694 5697 2698 5701
rect 2738 5697 2742 5701
rect 2758 5697 2762 5701
rect 2795 5695 2799 5699
rect 1806 5684 1810 5688
rect 1793 5678 1797 5682
rect 1827 5682 1831 5688
rect 1843 5684 1847 5688
rect 1911 5681 1915 5685
rect 1961 5681 1965 5685
rect 2012 5681 2016 5685
rect 2354 5681 2360 5685
rect 2413 5684 2417 5688
rect 2429 5684 2433 5688
rect 966 5667 970 5671
rect 1010 5667 1014 5671
rect 1030 5667 1034 5671
rect 1067 5665 1071 5669
rect 949 5654 953 5658
rect 965 5654 969 5658
rect 986 5652 990 5658
rect 1002 5654 1006 5658
rect 1468 5669 1472 5673
rect 1484 5669 1488 5675
rect 1521 5669 1525 5675
rect 1505 5665 1509 5669
rect 1529 5669 1533 5673
rect 1542 5669 1546 5675
rect 1579 5669 1583 5675
rect 1600 5669 1604 5675
rect 1616 5669 1620 5675
rect 1653 5669 1657 5675
rect 1563 5665 1567 5669
rect 1637 5665 1641 5669
rect 1661 5669 1665 5673
rect 1674 5669 1678 5675
rect 1711 5669 1715 5675
rect 1732 5669 1736 5675
rect 1748 5669 1752 5675
rect 1785 5669 1789 5675
rect 1695 5665 1699 5669
rect 1769 5665 1773 5669
rect 1793 5669 1797 5673
rect 1806 5669 1810 5675
rect 1843 5669 1847 5675
rect 1856 5674 1860 5678
rect 2390 5674 2396 5678
rect 2450 5682 2454 5688
rect 2466 5684 2470 5688
rect 2487 5684 2491 5688
rect 2474 5678 2478 5682
rect 2508 5682 2512 5688
rect 2524 5684 2528 5688
rect 2545 5684 2549 5688
rect 2561 5684 2565 5688
rect 2582 5682 2586 5688
rect 2598 5684 2602 5688
rect 2619 5684 2623 5688
rect 2606 5678 2610 5682
rect 2640 5682 2644 5688
rect 2656 5684 2660 5688
rect 2677 5684 2681 5688
rect 2693 5684 2697 5688
rect 2714 5682 2718 5688
rect 2730 5684 2734 5688
rect 2751 5684 2755 5688
rect 2738 5678 2742 5682
rect 2772 5682 2776 5688
rect 2788 5684 2792 5688
rect 1827 5665 1831 5669
rect 1911 5667 1915 5671
rect 1955 5667 1959 5671
rect 1975 5667 1979 5671
rect 2012 5665 2016 5669
rect 1023 5654 1027 5658
rect 1010 5648 1014 5652
rect 1044 5652 1048 5658
rect 1060 5654 1064 5658
rect 1483 5654 1487 5658
rect 1536 5654 1540 5658
rect 1586 5654 1590 5658
rect 1615 5654 1619 5658
rect 1668 5654 1672 5658
rect 1718 5654 1722 5658
rect 1747 5654 1751 5658
rect 1800 5654 1804 5658
rect 1850 5654 1854 5658
rect 1894 5654 1898 5658
rect 1910 5654 1914 5658
rect 949 5639 953 5645
rect 965 5639 969 5645
rect 1002 5639 1006 5645
rect 986 5635 990 5639
rect 1010 5639 1014 5643
rect 1023 5639 1027 5645
rect 1060 5639 1064 5645
rect 1073 5644 1077 5648
rect 1457 5647 1463 5651
rect 1931 5652 1935 5658
rect 1947 5654 1951 5658
rect 2413 5669 2417 5673
rect 2429 5669 2433 5675
rect 2466 5669 2470 5675
rect 2450 5665 2454 5669
rect 2474 5669 2478 5673
rect 2487 5669 2491 5675
rect 2524 5669 2528 5675
rect 2545 5669 2549 5675
rect 2561 5669 2565 5675
rect 2598 5669 2602 5675
rect 2508 5665 2512 5669
rect 2582 5665 2586 5669
rect 2606 5669 2610 5673
rect 2619 5669 2623 5675
rect 2656 5669 2660 5675
rect 2677 5669 2681 5675
rect 2693 5669 2697 5675
rect 2730 5669 2734 5675
rect 2640 5665 2644 5669
rect 2714 5665 2718 5669
rect 2738 5669 2742 5673
rect 2751 5669 2755 5675
rect 2788 5669 2792 5675
rect 2801 5674 2805 5678
rect 2772 5665 2776 5669
rect 1968 5654 1972 5658
rect 1955 5648 1959 5652
rect 1989 5652 1993 5658
rect 2005 5654 2009 5658
rect 2428 5654 2432 5658
rect 2481 5654 2485 5658
rect 2531 5654 2535 5658
rect 2560 5654 2564 5658
rect 2613 5654 2617 5658
rect 2663 5654 2667 5658
rect 2692 5654 2696 5658
rect 2745 5654 2749 5658
rect 2795 5654 2799 5658
rect 1397 5640 1403 5644
rect 1483 5640 1487 5644
rect 1550 5640 1554 5644
rect 1586 5640 1590 5644
rect 1615 5640 1619 5644
rect 1682 5640 1686 5644
rect 1718 5640 1722 5644
rect 1747 5640 1751 5644
rect 1814 5640 1818 5644
rect 1850 5640 1854 5644
rect 1894 5639 1898 5645
rect 1910 5639 1914 5645
rect 1947 5639 1951 5645
rect 1044 5635 1048 5639
rect 1599 5633 1603 5637
rect 1732 5633 1737 5637
rect 1931 5635 1935 5639
rect 1955 5639 1959 5643
rect 1968 5639 1972 5645
rect 2005 5639 2009 5645
rect 2018 5644 2022 5648
rect 2402 5647 2408 5651
rect 2342 5640 2348 5644
rect 2428 5640 2432 5644
rect 2495 5640 2499 5644
rect 2531 5640 2535 5644
rect 2560 5640 2564 5644
rect 2627 5640 2631 5644
rect 2663 5640 2667 5644
rect 2692 5640 2696 5644
rect 2759 5640 2763 5644
rect 2795 5640 2799 5644
rect 1989 5635 1993 5639
rect 2544 5633 2548 5637
rect 2677 5633 2682 5637
rect 964 5624 968 5628
rect 1017 5624 1021 5628
rect 1067 5624 1071 5628
rect 1725 5626 1729 5630
rect 1709 5622 1713 5626
rect 1741 5622 1745 5626
rect 1081 5617 1085 5621
rect 1457 5617 1463 5621
rect 1468 5618 1472 5622
rect 1909 5624 1913 5628
rect 1962 5624 1966 5628
rect 2012 5624 2016 5628
rect 2670 5626 2674 5630
rect 2654 5622 2658 5626
rect 2686 5622 2690 5626
rect 4484 5622 4488 5626
rect 4494 5622 4498 5626
rect 4504 5622 4508 5626
rect 2026 5617 2030 5621
rect 2402 5617 2408 5621
rect 2413 5618 2417 5622
rect 964 5610 968 5614
rect 1031 5610 1035 5614
rect 1067 5610 1071 5614
rect 1397 5610 1403 5614
rect 1468 5610 1472 5614
rect 1725 5610 1729 5614
rect 1909 5610 1913 5614
rect 1976 5610 1980 5614
rect 2012 5610 2016 5614
rect 2342 5610 2348 5614
rect 2413 5610 2417 5614
rect 2670 5610 2674 5614
rect 4484 5617 4488 5621
rect 4494 5617 4498 5621
rect 4504 5617 4508 5621
rect 4484 5612 4488 5616
rect 4494 5612 4498 5616
rect 4504 5612 4508 5616
rect 4484 5607 4488 5611
rect 4494 5607 4498 5611
rect 4504 5607 4508 5611
rect 4530 5622 4534 5626
rect 4540 5622 4544 5626
rect 4550 5622 4554 5626
rect 4530 5617 4534 5621
rect 4540 5617 4544 5621
rect 4550 5617 4554 5621
rect 4530 5612 4534 5616
rect 4540 5612 4544 5616
rect 4550 5612 4554 5616
rect 4530 5607 4534 5611
rect 4540 5607 4544 5611
rect 4550 5607 4554 5611
rect 1709 5603 1713 5607
rect 1741 5603 1745 5607
rect 2654 5603 2658 5607
rect 2686 5603 2690 5607
rect 1385 5596 1391 5600
rect 1709 5595 1713 5599
rect 1741 5595 1745 5599
rect 950 5589 954 5593
rect 1115 5589 1119 5593
rect 1433 5590 1439 5594
rect 1725 5590 1729 5594
rect 2330 5596 2336 5600
rect 2654 5595 2658 5599
rect 2686 5595 2690 5599
rect 1895 5589 1899 5593
rect 2060 5589 2064 5593
rect 2378 5590 2384 5594
rect 2670 5590 2674 5594
rect 618 5578 622 5582
rect 628 5578 632 5582
rect 638 5578 642 5582
rect 618 5573 622 5577
rect 628 5573 632 5577
rect 638 5573 642 5577
rect 618 5568 622 5572
rect 628 5568 632 5572
rect 638 5568 642 5572
rect 618 5563 622 5567
rect 628 5563 632 5567
rect 638 5563 642 5567
rect 664 5578 668 5582
rect 674 5578 678 5582
rect 684 5578 688 5582
rect 927 5581 931 5585
rect 939 5581 943 5585
rect 1125 5582 1129 5586
rect 1359 5582 1363 5586
rect 1421 5582 1427 5586
rect 1600 5583 1604 5587
rect 1732 5583 1737 5587
rect 1872 5581 1876 5585
rect 1884 5581 1888 5585
rect 2070 5582 2074 5586
rect 2304 5582 2308 5586
rect 2366 5582 2372 5586
rect 2545 5583 2549 5587
rect 2677 5583 2682 5587
rect 664 5573 668 5577
rect 674 5573 678 5577
rect 684 5573 688 5577
rect 955 5575 959 5579
rect 983 5575 987 5579
rect 1000 5575 1004 5579
rect 1056 5575 1060 5579
rect 1073 5575 1077 5579
rect 1107 5575 1111 5579
rect 1133 5575 1137 5579
rect 1216 5575 1220 5579
rect 1244 5575 1248 5579
rect 1261 5575 1265 5579
rect 1317 5575 1321 5579
rect 1334 5575 1338 5579
rect 1368 5575 1372 5579
rect 1457 5575 1463 5579
rect 1468 5576 1472 5580
rect 1856 5576 1860 5580
rect 1900 5575 1904 5579
rect 1928 5575 1932 5579
rect 1945 5575 1949 5579
rect 2001 5575 2005 5579
rect 2018 5575 2022 5579
rect 2052 5575 2056 5579
rect 2078 5575 2082 5579
rect 2161 5575 2165 5579
rect 2189 5575 2193 5579
rect 2206 5575 2210 5579
rect 2262 5575 2266 5579
rect 2279 5575 2283 5579
rect 2313 5575 2317 5579
rect 2402 5575 2408 5579
rect 2413 5576 2417 5580
rect 2801 5576 2805 5580
rect 664 5568 668 5572
rect 674 5568 678 5572
rect 684 5568 688 5572
rect 962 5568 966 5572
rect 1027 5568 1031 5572
rect 1049 5568 1053 5572
rect 1080 5568 1084 5572
rect 1124 5568 1128 5572
rect 1163 5568 1167 5572
rect 664 5563 668 5567
rect 674 5563 678 5567
rect 684 5563 688 5567
rect 956 5558 960 5562
rect 963 5561 967 5565
rect 983 5558 987 5562
rect 999 5558 1003 5562
rect 1009 5561 1013 5565
rect 1034 5561 1038 5565
rect 1056 5558 1060 5562
rect 1074 5558 1078 5562
rect 1081 5561 1085 5565
rect 1223 5568 1227 5572
rect 1288 5568 1292 5572
rect 1310 5568 1314 5572
rect 1341 5568 1345 5572
rect 1359 5568 1363 5572
rect 1409 5568 1415 5572
rect 1485 5569 1489 5573
rect 1535 5569 1539 5573
rect 1586 5569 1590 5573
rect 1617 5569 1621 5573
rect 1667 5569 1671 5573
rect 1718 5569 1722 5573
rect 1749 5569 1753 5573
rect 1799 5569 1803 5573
rect 1850 5569 1854 5573
rect 1907 5568 1911 5572
rect 1972 5568 1976 5572
rect 1994 5568 1998 5572
rect 2025 5568 2029 5572
rect 2069 5568 2073 5572
rect 2108 5568 2112 5572
rect 1107 5558 1111 5562
rect 1133 5558 1137 5562
rect 947 5541 951 5545
rect 959 5541 963 5545
rect 967 5542 971 5546
rect 989 5541 993 5545
rect 1002 5542 1006 5546
rect 1021 5542 1025 5546
rect 1040 5543 1044 5547
rect 1059 5539 1063 5543
rect 1079 5542 1083 5546
rect 1217 5558 1221 5562
rect 1224 5561 1228 5565
rect 1244 5558 1248 5562
rect 1260 5558 1264 5562
rect 1270 5561 1274 5565
rect 1295 5561 1299 5565
rect 1317 5558 1321 5562
rect 1335 5558 1339 5562
rect 1342 5561 1346 5565
rect 1445 5562 1451 5566
rect 1367 5558 1371 5562
rect 1145 5548 1149 5552
rect 1134 5541 1138 5545
rect 1174 5547 1178 5551
rect 1208 5541 1212 5545
rect 1220 5541 1224 5545
rect 1228 5542 1232 5546
rect 1153 5532 1157 5536
rect 956 5528 960 5532
rect 984 5528 988 5532
rect 999 5528 1003 5532
rect 1056 5528 1060 5532
rect 1074 5528 1078 5532
rect 977 5523 981 5527
rect 1024 5524 1031 5528
rect 1049 5523 1053 5527
rect 1092 5524 1096 5528
rect 977 5516 981 5520
rect 1008 5516 1012 5520
rect 1033 5516 1037 5520
rect 1092 5516 1096 5520
rect 1114 5516 1118 5520
rect 1250 5541 1254 5545
rect 1263 5542 1267 5546
rect 1282 5542 1286 5546
rect 1301 5543 1305 5547
rect 1320 5539 1324 5543
rect 1340 5542 1344 5546
rect 1485 5555 1489 5559
rect 1529 5555 1533 5559
rect 1549 5555 1553 5559
rect 1586 5553 1590 5557
rect 1617 5555 1621 5559
rect 1661 5555 1665 5559
rect 1681 5555 1685 5559
rect 1718 5553 1722 5557
rect 1749 5555 1753 5559
rect 1793 5555 1797 5559
rect 1813 5555 1817 5559
rect 1850 5553 1854 5557
rect 1901 5558 1905 5562
rect 1908 5561 1912 5565
rect 1928 5558 1932 5562
rect 1944 5558 1948 5562
rect 1954 5561 1958 5565
rect 1979 5561 1983 5565
rect 2001 5558 2005 5562
rect 2019 5558 2023 5562
rect 2026 5561 2030 5565
rect 2168 5568 2172 5572
rect 2233 5568 2237 5572
rect 2255 5568 2259 5572
rect 2286 5568 2290 5572
rect 2304 5568 2308 5572
rect 2354 5568 2360 5572
rect 2430 5569 2434 5573
rect 2480 5569 2484 5573
rect 2531 5569 2535 5573
rect 2562 5569 2566 5573
rect 2612 5569 2616 5573
rect 2663 5569 2667 5573
rect 2694 5569 2698 5573
rect 2744 5569 2748 5573
rect 2795 5569 2799 5573
rect 2052 5558 2056 5562
rect 2078 5558 2082 5562
rect 1372 5540 1376 5544
rect 1468 5542 1472 5546
rect 1484 5542 1488 5546
rect 1505 5540 1509 5546
rect 1521 5542 1525 5546
rect 1542 5542 1546 5546
rect 1529 5536 1533 5540
rect 1563 5540 1567 5546
rect 1579 5542 1583 5546
rect 1600 5542 1604 5546
rect 1616 5542 1620 5546
rect 1637 5540 1641 5546
rect 1653 5542 1657 5546
rect 1674 5542 1678 5546
rect 1661 5536 1665 5540
rect 1695 5540 1699 5546
rect 1711 5542 1715 5546
rect 1732 5542 1736 5546
rect 1748 5542 1752 5546
rect 1769 5540 1773 5546
rect 1785 5542 1789 5546
rect 1806 5542 1810 5546
rect 1793 5536 1797 5540
rect 1827 5540 1831 5546
rect 1843 5542 1847 5546
rect 1892 5541 1896 5545
rect 1904 5541 1908 5545
rect 1912 5542 1916 5546
rect 1934 5541 1938 5545
rect 1947 5542 1951 5546
rect 1966 5542 1970 5546
rect 1217 5528 1221 5532
rect 1245 5528 1249 5532
rect 1260 5528 1264 5532
rect 1317 5528 1321 5532
rect 1335 5528 1339 5532
rect 1367 5528 1371 5532
rect 1238 5523 1242 5527
rect 1285 5524 1292 5528
rect 1310 5523 1314 5527
rect 1353 5524 1357 5528
rect 1468 5527 1472 5531
rect 1484 5527 1488 5533
rect 1521 5527 1525 5533
rect 1238 5516 1242 5520
rect 1269 5516 1273 5520
rect 1294 5516 1298 5520
rect 1344 5516 1348 5520
rect 1353 5516 1357 5520
rect 1433 5516 1439 5520
rect 1505 5523 1509 5527
rect 1529 5527 1533 5531
rect 1542 5527 1546 5533
rect 1579 5527 1583 5533
rect 1600 5527 1604 5533
rect 1616 5527 1620 5533
rect 1653 5527 1657 5533
rect 1563 5523 1567 5527
rect 1637 5523 1641 5527
rect 1661 5527 1665 5531
rect 1674 5527 1678 5533
rect 1711 5527 1715 5533
rect 1732 5527 1736 5533
rect 1748 5527 1752 5533
rect 1785 5527 1789 5533
rect 1695 5523 1699 5527
rect 1769 5523 1773 5527
rect 1793 5527 1797 5531
rect 1806 5527 1810 5533
rect 1843 5527 1847 5533
rect 1856 5532 1860 5536
rect 1985 5543 1989 5547
rect 2004 5539 2008 5543
rect 2024 5542 2028 5546
rect 2162 5558 2166 5562
rect 2169 5561 2173 5565
rect 2189 5558 2193 5562
rect 2205 5558 2209 5562
rect 2215 5561 2219 5565
rect 2240 5561 2244 5565
rect 2262 5558 2266 5562
rect 2280 5558 2284 5562
rect 2287 5561 2291 5565
rect 2390 5562 2396 5566
rect 2312 5558 2316 5562
rect 2090 5548 2094 5552
rect 2079 5541 2083 5545
rect 2119 5547 2123 5551
rect 2153 5541 2157 5545
rect 2165 5541 2169 5545
rect 2173 5542 2177 5546
rect 2098 5532 2102 5536
rect 1901 5528 1905 5532
rect 1929 5528 1933 5532
rect 1944 5528 1948 5532
rect 2001 5528 2005 5532
rect 2019 5528 2023 5532
rect 1827 5523 1831 5527
rect 1922 5523 1926 5527
rect 1969 5524 1976 5528
rect 1994 5523 1998 5527
rect 2037 5524 2041 5528
rect 956 5509 960 5513
rect 984 5509 988 5513
rect 999 5509 1003 5513
rect 1033 5509 1037 5513
rect 1056 5509 1060 5513
rect 1074 5509 1078 5513
rect 1092 5509 1096 5513
rect 1217 5509 1221 5513
rect 1245 5509 1249 5513
rect 1260 5509 1264 5513
rect 1294 5509 1298 5513
rect 1317 5509 1321 5513
rect 1335 5509 1339 5513
rect 1353 5509 1357 5513
rect 1367 5509 1371 5513
rect 1445 5509 1451 5513
rect 1483 5512 1487 5516
rect 1536 5512 1540 5516
rect 1586 5512 1590 5516
rect 1615 5512 1619 5516
rect 1668 5512 1672 5516
rect 1718 5512 1722 5516
rect 1747 5512 1751 5516
rect 1800 5512 1804 5516
rect 1850 5512 1854 5516
rect 1922 5516 1926 5520
rect 1953 5516 1957 5520
rect 1978 5516 1982 5520
rect 2037 5516 2041 5520
rect 2059 5516 2063 5520
rect 2195 5541 2199 5545
rect 2208 5542 2212 5546
rect 2227 5542 2231 5546
rect 2246 5543 2250 5547
rect 2265 5539 2269 5543
rect 2285 5542 2289 5546
rect 2430 5555 2434 5559
rect 2474 5555 2478 5559
rect 2494 5555 2498 5559
rect 2531 5553 2535 5557
rect 2562 5555 2566 5559
rect 2606 5555 2610 5559
rect 2626 5555 2630 5559
rect 2663 5553 2667 5557
rect 2694 5555 2698 5559
rect 2738 5555 2742 5559
rect 2758 5555 2762 5559
rect 2795 5553 2799 5557
rect 2317 5540 2321 5544
rect 2413 5542 2417 5546
rect 2429 5542 2433 5546
rect 2450 5540 2454 5546
rect 2466 5542 2470 5546
rect 2487 5542 2491 5546
rect 2474 5536 2478 5540
rect 2508 5540 2512 5546
rect 2524 5542 2528 5546
rect 2545 5542 2549 5546
rect 2561 5542 2565 5546
rect 2582 5540 2586 5546
rect 2598 5542 2602 5546
rect 2619 5542 2623 5546
rect 2606 5536 2610 5540
rect 2640 5540 2644 5546
rect 2656 5542 2660 5546
rect 2677 5542 2681 5546
rect 2693 5542 2697 5546
rect 2714 5540 2718 5546
rect 2730 5542 2734 5546
rect 2751 5542 2755 5546
rect 2738 5536 2742 5540
rect 2772 5540 2776 5546
rect 2788 5542 2792 5546
rect 2162 5528 2166 5532
rect 2190 5528 2194 5532
rect 2205 5528 2209 5532
rect 2262 5528 2266 5532
rect 2280 5528 2284 5532
rect 2312 5528 2316 5532
rect 2183 5523 2187 5527
rect 2230 5524 2237 5528
rect 2255 5523 2259 5527
rect 2298 5524 2302 5528
rect 2413 5527 2417 5531
rect 2429 5527 2433 5533
rect 2466 5527 2470 5533
rect 2183 5516 2187 5520
rect 2214 5516 2218 5520
rect 2239 5516 2243 5520
rect 2289 5516 2293 5520
rect 2298 5516 2302 5520
rect 2378 5516 2384 5520
rect 2450 5523 2454 5527
rect 2474 5527 2478 5531
rect 2487 5527 2491 5533
rect 2524 5527 2528 5533
rect 2545 5527 2549 5533
rect 2561 5527 2565 5533
rect 2598 5527 2602 5533
rect 2508 5523 2512 5527
rect 2582 5523 2586 5527
rect 2606 5527 2610 5531
rect 2619 5527 2623 5533
rect 2656 5527 2660 5533
rect 2677 5527 2681 5533
rect 2693 5527 2697 5533
rect 2730 5527 2734 5533
rect 2640 5523 2644 5527
rect 2714 5523 2718 5527
rect 2738 5527 2742 5531
rect 2751 5527 2755 5533
rect 2788 5527 2792 5533
rect 4246 5532 4251 5536
rect 2772 5523 2776 5527
rect 1901 5509 1905 5513
rect 1929 5509 1933 5513
rect 1944 5509 1948 5513
rect 1978 5509 1982 5513
rect 2001 5509 2005 5513
rect 2019 5509 2023 5513
rect 2037 5509 2041 5513
rect 2162 5509 2166 5513
rect 2190 5509 2194 5513
rect 2205 5509 2209 5513
rect 2239 5509 2243 5513
rect 2262 5509 2266 5513
rect 2280 5509 2284 5513
rect 2298 5509 2302 5513
rect 2312 5509 2316 5513
rect 2390 5509 2396 5513
rect 2428 5512 2432 5516
rect 2481 5512 2485 5516
rect 2531 5512 2535 5516
rect 2560 5512 2564 5516
rect 2613 5512 2617 5516
rect 2663 5512 2667 5516
rect 2692 5512 2696 5516
rect 2745 5512 2749 5516
rect 2795 5512 2799 5516
rect 1163 5486 1167 5490
rect 1238 5502 1242 5506
rect 1269 5502 1273 5506
rect 1294 5502 1298 5506
rect 1344 5502 1348 5506
rect 1353 5502 1357 5506
rect 1457 5505 1463 5509
rect 1238 5495 1242 5499
rect 1285 5494 1292 5498
rect 1310 5495 1314 5499
rect 1397 5498 1403 5502
rect 1483 5498 1487 5502
rect 1550 5498 1554 5502
rect 1586 5498 1590 5502
rect 1615 5498 1619 5502
rect 1682 5498 1686 5502
rect 1718 5498 1722 5502
rect 1747 5498 1751 5502
rect 1814 5498 1818 5502
rect 1850 5498 1854 5502
rect 1353 5494 1357 5498
rect 1217 5490 1221 5494
rect 1245 5490 1249 5494
rect 1260 5490 1264 5494
rect 1317 5490 1321 5494
rect 1335 5490 1339 5494
rect 1367 5490 1371 5494
rect 1122 5473 1126 5477
rect 1176 5478 1180 5482
rect 1145 5468 1149 5476
rect 1208 5477 1212 5481
rect 1220 5477 1224 5481
rect 1228 5476 1232 5480
rect 1250 5477 1254 5481
rect 1263 5476 1267 5480
rect 1282 5476 1286 5480
rect 1301 5475 1305 5479
rect 1320 5479 1324 5483
rect 1340 5476 1344 5480
rect 2108 5486 2112 5490
rect 2183 5502 2187 5506
rect 2214 5502 2218 5506
rect 2239 5502 2243 5506
rect 2289 5502 2293 5506
rect 2298 5502 2302 5506
rect 2402 5505 2408 5509
rect 2183 5495 2187 5499
rect 2230 5494 2237 5498
rect 2255 5495 2259 5499
rect 2342 5498 2348 5502
rect 2428 5498 2432 5502
rect 2495 5498 2499 5502
rect 2531 5498 2535 5502
rect 2560 5498 2564 5502
rect 2627 5498 2631 5502
rect 2663 5498 2667 5502
rect 2692 5498 2696 5502
rect 2759 5498 2763 5502
rect 2795 5498 2799 5502
rect 2298 5494 2302 5498
rect 2162 5490 2166 5494
rect 2190 5490 2194 5494
rect 2205 5490 2209 5494
rect 2262 5490 2266 5494
rect 2280 5490 2284 5494
rect 2312 5490 2316 5494
rect 1373 5477 1377 5481
rect 2067 5473 2071 5477
rect 2121 5478 2125 5482
rect 1500 5468 1504 5472
rect 1217 5460 1221 5464
rect 1224 5457 1228 5461
rect 1244 5460 1248 5464
rect 1260 5460 1264 5464
rect 1270 5457 1274 5461
rect 1295 5457 1299 5461
rect 1317 5460 1321 5464
rect 1335 5460 1339 5464
rect 1342 5457 1346 5461
rect 1367 5460 1371 5464
rect 1772 5461 1776 5465
rect 1153 5450 1157 5454
rect 1223 5450 1227 5454
rect 1288 5450 1292 5454
rect 1310 5450 1314 5454
rect 1341 5450 1345 5454
rect 1421 5450 1427 5454
rect 2090 5468 2094 5476
rect 2153 5477 2157 5481
rect 2165 5477 2169 5481
rect 2173 5476 2177 5480
rect 2195 5477 2199 5481
rect 2208 5476 2212 5480
rect 2227 5476 2231 5480
rect 2246 5475 2250 5479
rect 2265 5479 2269 5483
rect 2285 5476 2289 5480
rect 2318 5477 2322 5481
rect 2162 5460 2166 5464
rect 2169 5457 2173 5461
rect 2189 5460 2193 5464
rect 2205 5460 2209 5464
rect 2215 5457 2219 5461
rect 2240 5457 2244 5461
rect 2262 5460 2266 5464
rect 2280 5460 2284 5464
rect 2287 5457 2291 5461
rect 2312 5460 2316 5464
rect 1216 5443 1220 5447
rect 1244 5443 1248 5447
rect 1261 5443 1265 5447
rect 1317 5443 1321 5447
rect 1334 5443 1338 5447
rect 1368 5443 1372 5447
rect 1457 5443 1463 5447
rect 2098 5450 2102 5454
rect 2168 5450 2172 5454
rect 2233 5450 2237 5454
rect 2255 5450 2259 5454
rect 2286 5450 2290 5454
rect 2366 5450 2372 5454
rect 992 5432 996 5436
rect 1082 5432 1086 5436
rect 1163 5432 1167 5436
rect 1754 5441 1758 5445
rect 1223 5436 1227 5440
rect 1288 5436 1292 5440
rect 1310 5436 1314 5440
rect 1341 5436 1345 5440
rect 1421 5436 1427 5440
rect 1840 5440 1844 5444
rect 2161 5443 2165 5447
rect 2189 5443 2193 5447
rect 2206 5443 2210 5447
rect 2262 5443 2266 5447
rect 2279 5443 2283 5447
rect 2313 5443 2317 5447
rect 2402 5443 2408 5447
rect 1217 5426 1221 5430
rect 1224 5429 1228 5433
rect 1244 5426 1248 5430
rect 1260 5426 1264 5430
rect 1270 5429 1274 5433
rect 1295 5429 1299 5433
rect 1317 5426 1321 5430
rect 1335 5426 1339 5430
rect 1342 5429 1346 5433
rect 1937 5432 1941 5436
rect 1367 5426 1371 5430
rect 1409 5428 1415 5432
rect 1680 5428 1684 5432
rect 974 5412 978 5416
rect 1009 5411 1013 5415
rect 1064 5412 1068 5416
rect 1093 5411 1097 5415
rect 1145 5412 1149 5416
rect 1173 5411 1177 5415
rect 1208 5409 1212 5413
rect 1220 5409 1224 5413
rect 1228 5410 1232 5414
rect 982 5396 986 5400
rect 1072 5396 1076 5400
rect 1153 5396 1157 5400
rect 1250 5409 1254 5413
rect 1263 5410 1267 5414
rect 1282 5410 1286 5414
rect 1301 5411 1305 5415
rect 1320 5407 1324 5411
rect 1340 5410 1344 5414
rect 1762 5425 1766 5429
rect 2027 5432 2031 5436
rect 2108 5432 2112 5436
rect 2168 5436 2172 5440
rect 2233 5436 2237 5440
rect 2255 5436 2259 5440
rect 2286 5436 2290 5440
rect 2366 5436 2372 5440
rect 1507 5418 1512 5422
rect 2162 5426 2166 5430
rect 2169 5429 2173 5433
rect 2189 5426 2193 5430
rect 2205 5426 2209 5430
rect 2215 5429 2219 5433
rect 2240 5429 2244 5433
rect 2262 5426 2266 5430
rect 2280 5426 2284 5430
rect 2287 5429 2291 5433
rect 2312 5426 2316 5430
rect 1372 5408 1376 5412
rect 1217 5396 1221 5400
rect 1245 5396 1249 5400
rect 1260 5396 1264 5400
rect 1317 5396 1321 5400
rect 1335 5396 1339 5400
rect 1367 5396 1371 5400
rect 1397 5398 1403 5402
rect 1238 5391 1242 5395
rect 1285 5392 1292 5396
rect 1310 5391 1314 5395
rect 1353 5392 1357 5396
rect 1636 5395 1640 5399
rect 1238 5384 1242 5388
rect 1269 5384 1273 5388
rect 1294 5384 1298 5388
rect 1353 5384 1357 5388
rect 1433 5384 1439 5388
rect 1217 5377 1221 5381
rect 1245 5377 1249 5381
rect 1260 5377 1264 5381
rect 1294 5377 1298 5381
rect 1317 5377 1321 5381
rect 1335 5377 1339 5381
rect 1353 5377 1357 5381
rect 1367 5377 1371 5381
rect 1445 5377 1451 5381
rect 1680 5387 1684 5391
rect 992 5354 996 5358
rect 939 5341 943 5345
rect 1082 5354 1086 5358
rect 974 5336 978 5344
rect 1006 5338 1010 5342
rect 1095 5346 1099 5350
rect 1040 5340 1044 5344
rect 1013 5332 1017 5336
rect 1028 5332 1032 5336
rect 982 5318 986 5322
rect 1064 5336 1068 5344
rect 1163 5354 1167 5358
rect 1238 5370 1242 5374
rect 1269 5370 1273 5374
rect 1294 5370 1298 5374
rect 1353 5370 1357 5374
rect 1433 5370 1439 5374
rect 1238 5363 1242 5367
rect 1285 5362 1292 5366
rect 1310 5363 1314 5367
rect 1353 5362 1357 5366
rect 1217 5358 1221 5362
rect 1245 5358 1249 5362
rect 1260 5358 1264 5362
rect 1317 5358 1321 5362
rect 1335 5358 1339 5362
rect 1367 5358 1371 5362
rect 1176 5346 1180 5350
rect 1122 5340 1126 5344
rect 1103 5332 1107 5336
rect 1118 5332 1122 5336
rect 1072 5318 1076 5322
rect 1145 5336 1149 5344
rect 1208 5345 1212 5349
rect 1220 5345 1224 5349
rect 1228 5344 1232 5348
rect 1250 5345 1254 5349
rect 1263 5344 1267 5348
rect 1282 5344 1286 5348
rect 1301 5343 1305 5347
rect 1320 5347 1324 5351
rect 1340 5344 1344 5348
rect 1772 5381 1776 5385
rect 1919 5412 1923 5416
rect 1954 5411 1958 5415
rect 2009 5412 2013 5416
rect 2038 5411 2042 5415
rect 2090 5412 2094 5416
rect 2118 5411 2122 5415
rect 2153 5409 2157 5413
rect 2165 5409 2169 5413
rect 2173 5410 2177 5414
rect 1927 5396 1931 5400
rect 2017 5396 2021 5400
rect 2098 5396 2102 5400
rect 2195 5409 2199 5413
rect 2208 5410 2212 5414
rect 2227 5410 2231 5414
rect 2246 5411 2250 5415
rect 2265 5407 2269 5411
rect 2285 5410 2289 5414
rect 2317 5408 2321 5412
rect 2162 5396 2166 5400
rect 2190 5396 2194 5400
rect 2205 5396 2209 5400
rect 2262 5396 2266 5400
rect 2280 5396 2284 5400
rect 2312 5396 2316 5400
rect 2183 5391 2187 5395
rect 2230 5392 2237 5396
rect 2255 5391 2259 5395
rect 2298 5392 2302 5396
rect 2183 5384 2187 5388
rect 2214 5384 2218 5388
rect 2239 5384 2243 5388
rect 2298 5384 2302 5388
rect 2378 5384 2384 5388
rect 2162 5377 2166 5381
rect 2190 5377 2194 5381
rect 2205 5377 2209 5381
rect 2239 5377 2243 5381
rect 2262 5377 2266 5381
rect 2280 5377 2284 5381
rect 2298 5377 2302 5381
rect 2312 5377 2316 5381
rect 2390 5377 2396 5381
rect 1373 5345 1377 5349
rect 1754 5363 1758 5371
rect 1785 5367 1789 5371
rect 1793 5359 1797 5363
rect 1808 5359 1812 5363
rect 1815 5359 1819 5363
rect 1830 5359 1834 5363
rect 1762 5345 1766 5349
rect 1937 5354 1941 5358
rect 1500 5338 1504 5342
rect 1884 5341 1888 5345
rect 2027 5354 2031 5358
rect 1217 5328 1221 5332
rect 1224 5325 1228 5329
rect 1244 5328 1248 5332
rect 1260 5328 1264 5332
rect 1270 5325 1274 5329
rect 1295 5325 1299 5329
rect 1317 5328 1321 5332
rect 1335 5328 1339 5332
rect 1342 5325 1346 5329
rect 1367 5328 1371 5332
rect 1772 5331 1776 5335
rect 1153 5318 1157 5322
rect 1223 5318 1227 5322
rect 1288 5318 1292 5322
rect 1310 5318 1314 5322
rect 1341 5318 1345 5322
rect 1421 5318 1427 5322
rect 1919 5336 1923 5344
rect 1951 5338 1955 5342
rect 2040 5346 2044 5350
rect 1985 5340 1989 5344
rect 1958 5332 1962 5336
rect 1973 5332 1977 5336
rect 1927 5318 1931 5322
rect 2009 5336 2013 5344
rect 2108 5354 2112 5358
rect 2183 5370 2187 5374
rect 2214 5370 2218 5374
rect 2239 5370 2243 5374
rect 2298 5370 2302 5374
rect 2378 5370 2384 5374
rect 2183 5363 2187 5367
rect 2230 5362 2237 5366
rect 2255 5363 2259 5367
rect 2298 5362 2302 5366
rect 2162 5358 2166 5362
rect 2190 5358 2194 5362
rect 2205 5358 2209 5362
rect 2262 5358 2266 5362
rect 2280 5358 2284 5362
rect 2312 5358 2316 5362
rect 2121 5346 2125 5350
rect 2067 5340 2071 5344
rect 2048 5332 2052 5336
rect 2063 5332 2067 5336
rect 2017 5318 2021 5322
rect 2090 5336 2094 5344
rect 2153 5345 2157 5349
rect 2165 5345 2169 5349
rect 2173 5344 2177 5348
rect 2195 5345 2199 5349
rect 2208 5344 2212 5348
rect 2227 5344 2231 5348
rect 2246 5343 2250 5347
rect 2265 5347 2269 5351
rect 2285 5344 2289 5348
rect 2318 5345 2322 5349
rect 2162 5328 2166 5332
rect 2169 5325 2173 5329
rect 2189 5328 2193 5332
rect 2205 5328 2209 5332
rect 2215 5325 2219 5329
rect 2240 5325 2244 5329
rect 2262 5328 2266 5332
rect 2280 5328 2284 5332
rect 2287 5325 2291 5329
rect 2312 5328 2316 5332
rect 2098 5318 2102 5322
rect 2168 5318 2172 5322
rect 2233 5318 2237 5322
rect 2255 5318 2259 5322
rect 2286 5318 2290 5322
rect 2366 5318 2372 5322
rect 1216 5311 1220 5315
rect 1244 5311 1248 5315
rect 1261 5311 1265 5315
rect 1317 5311 1321 5315
rect 1334 5311 1338 5315
rect 1368 5311 1372 5315
rect 1457 5311 1463 5315
rect 1754 5311 1758 5315
rect 1058 5297 1062 5301
rect 1163 5297 1167 5301
rect 1223 5304 1227 5308
rect 1288 5304 1292 5308
rect 1310 5304 1314 5308
rect 1341 5304 1345 5308
rect 1421 5304 1427 5308
rect 1842 5310 1846 5314
rect 2161 5311 2165 5315
rect 2189 5311 2193 5315
rect 2206 5311 2210 5315
rect 2262 5311 2266 5315
rect 2279 5311 2283 5315
rect 2313 5311 2317 5315
rect 2402 5311 2408 5315
rect 4484 5313 4488 5317
rect 4494 5313 4498 5317
rect 4504 5313 4508 5317
rect 1433 5302 1439 5306
rect 1574 5302 1579 5306
rect 1217 5294 1221 5298
rect 1224 5297 1228 5301
rect 1244 5294 1248 5298
rect 1260 5294 1264 5298
rect 1270 5297 1274 5301
rect 1295 5297 1299 5301
rect 1317 5294 1321 5298
rect 1335 5294 1339 5298
rect 1342 5297 1346 5301
rect 1367 5294 1371 5298
rect 1040 5277 1044 5281
rect 618 5269 622 5273
rect 628 5269 632 5273
rect 638 5269 642 5273
rect 618 5264 622 5268
rect 628 5264 632 5268
rect 638 5264 642 5268
rect 618 5259 622 5263
rect 628 5259 632 5263
rect 638 5259 642 5263
rect 618 5254 622 5258
rect 628 5254 632 5258
rect 638 5254 642 5258
rect 664 5269 668 5273
rect 674 5269 678 5273
rect 684 5269 688 5273
rect 1068 5276 1072 5280
rect 1145 5277 1149 5281
rect 1174 5276 1178 5280
rect 1208 5277 1212 5281
rect 1220 5277 1224 5281
rect 1228 5278 1232 5282
rect 1250 5277 1254 5281
rect 1263 5278 1267 5282
rect 1282 5278 1286 5282
rect 1301 5279 1305 5283
rect 1320 5275 1324 5279
rect 1340 5278 1344 5282
rect 1385 5293 1391 5297
rect 1492 5293 1496 5297
rect 1762 5295 1766 5299
rect 2003 5297 2007 5301
rect 2108 5297 2112 5301
rect 4484 5308 4488 5312
rect 4494 5308 4498 5312
rect 4504 5308 4508 5312
rect 2168 5304 2172 5308
rect 2233 5304 2237 5308
rect 2255 5304 2259 5308
rect 2286 5304 2290 5308
rect 2366 5304 2372 5308
rect 4484 5303 4488 5307
rect 4494 5303 4498 5307
rect 4504 5303 4508 5307
rect 2162 5294 2166 5298
rect 2169 5297 2173 5301
rect 2189 5294 2193 5298
rect 2205 5294 2209 5298
rect 2215 5297 2219 5301
rect 2240 5297 2244 5301
rect 2262 5294 2266 5298
rect 2280 5294 2284 5298
rect 2287 5297 2291 5301
rect 4484 5298 4488 5302
rect 4494 5298 4498 5302
rect 4504 5298 4508 5302
rect 4530 5313 4534 5317
rect 4540 5313 4544 5317
rect 4550 5313 4554 5317
rect 4530 5308 4534 5312
rect 4540 5308 4544 5312
rect 4550 5308 4554 5312
rect 4530 5303 4534 5307
rect 4540 5303 4544 5307
rect 4550 5303 4554 5307
rect 4530 5298 4534 5302
rect 4540 5298 4544 5302
rect 4550 5298 4554 5302
rect 2312 5294 2316 5298
rect 1507 5288 1512 5292
rect 1445 5284 1451 5288
rect 1372 5276 1376 5280
rect 1457 5277 1463 5281
rect 1500 5277 1504 5281
rect 664 5264 668 5268
rect 674 5264 678 5268
rect 684 5264 688 5268
rect 664 5259 668 5263
rect 674 5259 678 5263
rect 684 5259 688 5263
rect 1048 5261 1052 5265
rect 664 5254 668 5258
rect 674 5254 678 5258
rect 684 5254 688 5258
rect 1153 5261 1157 5265
rect 1217 5264 1221 5268
rect 1245 5264 1249 5268
rect 1260 5264 1264 5268
rect 1317 5264 1321 5268
rect 1335 5264 1339 5268
rect 1367 5264 1371 5268
rect 1421 5265 1427 5269
rect 1542 5265 1546 5269
rect 1238 5259 1242 5263
rect 1285 5260 1292 5264
rect 1310 5259 1314 5263
rect 1353 5260 1357 5264
rect 1238 5252 1242 5256
rect 1269 5252 1273 5256
rect 1294 5252 1298 5256
rect 1353 5252 1357 5256
rect 1433 5252 1439 5256
rect 1575 5257 1579 5261
rect 1217 5245 1221 5249
rect 1245 5245 1249 5249
rect 1260 5245 1264 5249
rect 1294 5245 1298 5249
rect 1317 5245 1321 5249
rect 1335 5245 1339 5249
rect 1353 5245 1357 5249
rect 1367 5245 1371 5249
rect 1445 5245 1451 5249
rect 1058 5222 1062 5226
rect 1071 5214 1075 5218
rect 1019 5208 1023 5212
rect 1040 5204 1044 5212
rect 1163 5222 1167 5226
rect 1238 5238 1242 5242
rect 1269 5238 1273 5242
rect 1294 5238 1298 5242
rect 1353 5238 1357 5242
rect 1433 5238 1439 5242
rect 1238 5231 1242 5235
rect 1285 5230 1292 5234
rect 1310 5231 1314 5235
rect 1353 5230 1357 5234
rect 1217 5226 1221 5230
rect 1245 5226 1249 5230
rect 1260 5226 1264 5230
rect 1317 5226 1321 5230
rect 1335 5226 1339 5230
rect 1367 5226 1371 5230
rect 1122 5209 1126 5213
rect 1176 5214 1180 5218
rect 1079 5200 1083 5204
rect 1094 5200 1098 5204
rect 1048 5186 1052 5190
rect 1145 5204 1149 5212
rect 1208 5213 1212 5217
rect 1220 5213 1224 5217
rect 1228 5212 1232 5216
rect 1250 5213 1254 5217
rect 1263 5212 1267 5216
rect 1282 5212 1286 5216
rect 1301 5211 1305 5215
rect 1320 5215 1324 5219
rect 1340 5212 1344 5216
rect 1772 5251 1776 5255
rect 1985 5277 1989 5281
rect 2013 5276 2017 5280
rect 2090 5277 2094 5281
rect 2119 5276 2123 5280
rect 2153 5277 2157 5281
rect 2165 5277 2169 5281
rect 2173 5278 2177 5282
rect 2195 5277 2199 5281
rect 2208 5278 2212 5282
rect 2227 5278 2231 5282
rect 2246 5279 2250 5283
rect 2265 5275 2269 5279
rect 2285 5278 2289 5282
rect 2317 5276 2321 5280
rect 1993 5261 1997 5265
rect 2098 5261 2102 5265
rect 2162 5264 2166 5268
rect 2190 5264 2194 5268
rect 2205 5264 2209 5268
rect 2262 5264 2266 5268
rect 2280 5264 2284 5268
rect 2312 5264 2316 5268
rect 2183 5259 2187 5263
rect 2230 5260 2237 5264
rect 2255 5259 2259 5263
rect 2298 5260 2302 5264
rect 2183 5252 2187 5256
rect 2214 5252 2218 5256
rect 2239 5252 2243 5256
rect 2298 5252 2302 5256
rect 2378 5252 2384 5256
rect 2162 5245 2166 5249
rect 2190 5245 2194 5249
rect 2205 5245 2209 5249
rect 2239 5245 2243 5249
rect 2262 5245 2266 5249
rect 2280 5245 2284 5249
rect 2298 5245 2302 5249
rect 2312 5245 2316 5249
rect 2390 5245 2396 5249
rect 1373 5213 1377 5217
rect 1754 5233 1758 5241
rect 1785 5237 1789 5241
rect 1793 5229 1797 5233
rect 1808 5229 1812 5233
rect 1762 5215 1766 5219
rect 2003 5222 2007 5226
rect 2016 5214 2020 5218
rect 1500 5208 1504 5212
rect 1964 5208 1968 5212
rect 1217 5196 1221 5200
rect 1224 5193 1228 5197
rect 1244 5196 1248 5200
rect 1260 5196 1264 5200
rect 1270 5193 1274 5197
rect 1295 5193 1299 5197
rect 1317 5196 1321 5200
rect 1335 5196 1339 5200
rect 1342 5193 1346 5197
rect 1367 5196 1371 5200
rect 1985 5204 1989 5212
rect 2108 5222 2112 5226
rect 2183 5238 2187 5242
rect 2214 5238 2218 5242
rect 2239 5238 2243 5242
rect 2298 5238 2302 5242
rect 2378 5238 2384 5242
rect 2183 5231 2187 5235
rect 2230 5230 2237 5234
rect 2255 5231 2259 5235
rect 2298 5230 2302 5234
rect 2162 5226 2166 5230
rect 2190 5226 2194 5230
rect 2205 5226 2209 5230
rect 2262 5226 2266 5230
rect 2280 5226 2284 5230
rect 2312 5226 2316 5230
rect 2067 5209 2071 5213
rect 2121 5214 2125 5218
rect 1153 5186 1157 5190
rect 1223 5186 1227 5190
rect 1288 5186 1292 5190
rect 1310 5186 1314 5190
rect 1341 5186 1345 5190
rect 1357 5186 1361 5190
rect 1421 5186 1427 5190
rect 1807 5190 1811 5194
rect 2024 5200 2028 5204
rect 2039 5200 2043 5204
rect 1993 5186 1997 5190
rect 2090 5204 2094 5212
rect 2153 5213 2157 5217
rect 2165 5213 2169 5217
rect 2173 5212 2177 5216
rect 2195 5213 2199 5217
rect 2208 5212 2212 5216
rect 2227 5212 2231 5216
rect 2246 5211 2250 5215
rect 2265 5215 2269 5219
rect 2285 5212 2289 5216
rect 2318 5213 2322 5217
rect 2162 5196 2166 5200
rect 2169 5193 2173 5197
rect 2189 5196 2193 5200
rect 2205 5196 2209 5200
rect 2215 5193 2219 5197
rect 2240 5193 2244 5197
rect 2262 5196 2266 5200
rect 2280 5196 2284 5200
rect 2287 5193 2291 5197
rect 2312 5196 2316 5200
rect 2098 5186 2102 5190
rect 2168 5186 2172 5190
rect 2233 5186 2237 5190
rect 2255 5186 2259 5190
rect 2286 5186 2290 5190
rect 2302 5186 2306 5190
rect 2366 5186 2372 5190
rect 1216 5179 1220 5183
rect 1244 5179 1248 5183
rect 1261 5179 1265 5183
rect 1317 5179 1321 5183
rect 1334 5179 1338 5183
rect 1368 5179 1372 5183
rect 1457 5179 1463 5183
rect 2161 5179 2165 5183
rect 2189 5179 2193 5183
rect 2206 5179 2210 5183
rect 2262 5179 2266 5183
rect 2279 5179 2283 5183
rect 2313 5179 2317 5183
rect 2402 5179 2408 5183
rect 1082 5166 1086 5170
rect 1163 5166 1167 5170
rect 1223 5172 1227 5176
rect 1288 5172 1292 5176
rect 1310 5172 1314 5176
rect 1341 5172 1345 5176
rect 1357 5172 1361 5176
rect 1409 5169 1415 5173
rect 1615 5169 1619 5173
rect 1666 5169 1670 5173
rect 1716 5169 1720 5173
rect 1217 5162 1221 5166
rect 1224 5165 1228 5169
rect 1244 5162 1248 5166
rect 1260 5162 1264 5166
rect 1270 5165 1274 5169
rect 1295 5165 1299 5169
rect 1317 5162 1321 5166
rect 1335 5162 1339 5166
rect 1342 5165 1346 5169
rect 2027 5166 2031 5170
rect 1367 5162 1371 5166
rect 1445 5162 1451 5166
rect 1064 5146 1068 5150
rect 1093 5145 1097 5149
rect 1145 5146 1149 5150
rect 1173 5145 1177 5149
rect 1208 5145 1212 5149
rect 1220 5145 1224 5149
rect 1228 5146 1232 5150
rect 1072 5130 1076 5134
rect 1153 5130 1157 5134
rect 1250 5145 1254 5149
rect 1263 5146 1267 5150
rect 1282 5146 1286 5150
rect 1301 5147 1305 5151
rect 1320 5143 1324 5147
rect 1340 5146 1344 5150
rect 1615 5153 1619 5157
rect 1652 5155 1656 5159
rect 1672 5155 1676 5159
rect 1716 5155 1720 5159
rect 2108 5166 2112 5170
rect 2168 5172 2172 5176
rect 2233 5172 2237 5176
rect 2255 5172 2259 5176
rect 2286 5172 2290 5176
rect 2302 5172 2306 5176
rect 2354 5169 2360 5173
rect 2560 5169 2564 5173
rect 2611 5169 2615 5173
rect 2661 5169 2665 5173
rect 2162 5162 2166 5166
rect 2169 5165 2173 5169
rect 2189 5162 2193 5166
rect 2205 5162 2209 5166
rect 2215 5165 2219 5169
rect 2240 5165 2244 5169
rect 2262 5162 2266 5166
rect 2280 5162 2284 5166
rect 2287 5165 2291 5169
rect 2312 5162 2316 5166
rect 2390 5162 2396 5166
rect 1372 5144 1376 5148
rect 1622 5142 1626 5146
rect 1638 5140 1642 5146
rect 1659 5142 1663 5146
rect 2009 5146 2013 5150
rect 1680 5142 1684 5146
rect 1696 5140 1700 5146
rect 1672 5136 1676 5140
rect 1717 5142 1721 5146
rect 1733 5142 1737 5146
rect 2038 5145 2042 5149
rect 2090 5146 2094 5150
rect 2118 5145 2122 5149
rect 2153 5145 2157 5149
rect 2165 5145 2169 5149
rect 2173 5146 2177 5150
rect 1217 5132 1221 5136
rect 1245 5132 1249 5136
rect 1260 5132 1264 5136
rect 1317 5132 1321 5136
rect 1335 5132 1339 5136
rect 1367 5132 1371 5136
rect 1600 5132 1604 5136
rect 1238 5127 1242 5131
rect 1285 5128 1292 5132
rect 1310 5127 1314 5131
rect 1353 5128 1357 5132
rect 1622 5127 1626 5133
rect 1659 5127 1663 5133
rect 1238 5120 1242 5124
rect 1269 5120 1273 5124
rect 1294 5120 1298 5124
rect 1353 5120 1357 5124
rect 1433 5120 1439 5124
rect 1638 5123 1642 5127
rect 1672 5127 1676 5131
rect 1680 5127 1684 5133
rect 1717 5127 1721 5133
rect 1733 5127 1737 5133
rect 2017 5130 2021 5134
rect 1696 5123 1700 5127
rect 1217 5113 1221 5117
rect 1245 5113 1249 5117
rect 1260 5113 1264 5117
rect 1294 5113 1298 5117
rect 1317 5113 1321 5117
rect 1335 5113 1339 5117
rect 1353 5113 1357 5117
rect 1367 5113 1371 5117
rect 1445 5113 1451 5117
rect 1082 5090 1086 5094
rect 1095 5082 1099 5086
rect 1037 5076 1041 5080
rect 1064 5072 1068 5080
rect 1163 5090 1167 5094
rect 1176 5082 1180 5086
rect 1122 5076 1126 5080
rect 1103 5068 1107 5072
rect 1118 5068 1122 5072
rect 1072 5054 1076 5058
rect 1145 5072 1149 5080
rect 1238 5106 1242 5110
rect 1269 5106 1273 5110
rect 1294 5106 1298 5110
rect 1353 5106 1357 5110
rect 1433 5106 1439 5110
rect 1615 5112 1619 5116
rect 1665 5112 1669 5116
rect 1718 5112 1722 5116
rect 2098 5130 2102 5134
rect 2195 5145 2199 5149
rect 2208 5146 2212 5150
rect 2227 5146 2231 5150
rect 2246 5147 2250 5151
rect 2265 5143 2269 5147
rect 2285 5146 2289 5150
rect 2560 5153 2564 5157
rect 2597 5155 2601 5159
rect 2617 5155 2621 5159
rect 2661 5155 2665 5159
rect 2317 5144 2321 5148
rect 2567 5142 2571 5146
rect 2583 5140 2587 5146
rect 2604 5142 2608 5146
rect 2625 5142 2629 5146
rect 2641 5140 2645 5146
rect 2617 5136 2621 5140
rect 2662 5142 2666 5146
rect 2678 5142 2682 5146
rect 2162 5132 2166 5136
rect 2190 5132 2194 5136
rect 2205 5132 2209 5136
rect 2262 5132 2266 5136
rect 2280 5132 2284 5136
rect 2312 5132 2316 5136
rect 2545 5132 2549 5136
rect 2183 5127 2187 5131
rect 2230 5128 2237 5132
rect 2255 5127 2259 5131
rect 2298 5128 2302 5132
rect 2567 5127 2571 5133
rect 2604 5127 2608 5133
rect 2183 5120 2187 5124
rect 2214 5120 2218 5124
rect 2239 5120 2243 5124
rect 2298 5120 2302 5124
rect 2378 5120 2384 5124
rect 2583 5123 2587 5127
rect 2617 5127 2621 5131
rect 2625 5127 2629 5133
rect 2662 5127 2666 5133
rect 2678 5127 2682 5133
rect 2641 5123 2645 5127
rect 2162 5113 2166 5117
rect 2190 5113 2194 5117
rect 2205 5113 2209 5117
rect 2239 5113 2243 5117
rect 2262 5113 2266 5117
rect 2280 5113 2284 5117
rect 2298 5113 2302 5117
rect 2312 5113 2316 5117
rect 2390 5113 2396 5117
rect 1457 5105 1463 5109
rect 1238 5099 1242 5103
rect 1285 5098 1292 5102
rect 1310 5099 1314 5103
rect 1353 5098 1357 5102
rect 1397 5098 1403 5102
rect 1615 5098 1619 5102
rect 1651 5098 1655 5102
rect 1718 5098 1722 5102
rect 1217 5094 1221 5098
rect 1245 5094 1249 5098
rect 1260 5094 1264 5098
rect 1317 5094 1321 5098
rect 1335 5094 1339 5098
rect 1367 5094 1371 5098
rect 1208 5081 1212 5085
rect 1220 5081 1224 5085
rect 1228 5080 1232 5084
rect 1250 5081 1254 5085
rect 1263 5080 1267 5084
rect 1282 5080 1286 5084
rect 1184 5068 1188 5072
rect 1199 5068 1203 5072
rect 1301 5079 1305 5083
rect 1320 5083 1324 5087
rect 1340 5080 1344 5084
rect 1584 5090 1588 5094
rect 1725 5090 1729 5094
rect 2027 5090 2031 5094
rect 1584 5081 1588 5085
rect 1608 5081 1612 5085
rect 1733 5083 1737 5087
rect 2040 5082 2044 5086
rect 1600 5074 1604 5078
rect 1982 5076 1986 5080
rect 1153 5054 1157 5058
rect 1217 5064 1221 5068
rect 1224 5061 1228 5065
rect 1244 5064 1248 5068
rect 1260 5064 1264 5068
rect 1270 5061 1274 5065
rect 1295 5061 1299 5065
rect 1317 5064 1321 5068
rect 1335 5064 1339 5068
rect 1342 5061 1346 5065
rect 1367 5064 1371 5068
rect 1409 5067 1415 5071
rect 1617 5067 1621 5071
rect 1667 5067 1671 5071
rect 1718 5067 1722 5071
rect 1745 5069 1749 5073
rect 1807 5069 1811 5073
rect 1445 5060 1451 5064
rect 1223 5054 1227 5058
rect 1288 5054 1292 5058
rect 1310 5054 1314 5058
rect 1341 5054 1345 5058
rect 1421 5054 1427 5058
rect 1216 5047 1220 5051
rect 1244 5047 1248 5051
rect 1261 5047 1265 5051
rect 1317 5047 1321 5051
rect 1334 5047 1338 5051
rect 1368 5047 1372 5051
rect 1457 5047 1463 5051
rect 1617 5053 1621 5057
rect 1661 5053 1665 5057
rect 1681 5053 1685 5057
rect 1718 5051 1722 5055
rect 1756 5056 1761 5064
rect 1844 5056 1857 5064
rect 2009 5072 2013 5080
rect 2108 5090 2112 5094
rect 2121 5082 2125 5086
rect 2067 5076 2071 5080
rect 2048 5068 2052 5072
rect 2063 5068 2067 5072
rect 2017 5054 2021 5058
rect 2090 5072 2094 5080
rect 2183 5106 2187 5110
rect 2214 5106 2218 5110
rect 2239 5106 2243 5110
rect 2298 5106 2302 5110
rect 2378 5106 2384 5110
rect 2560 5112 2564 5116
rect 2610 5112 2614 5116
rect 2663 5112 2667 5116
rect 2402 5105 2408 5109
rect 2183 5099 2187 5103
rect 2230 5098 2237 5102
rect 2255 5099 2259 5103
rect 2298 5098 2302 5102
rect 2342 5098 2348 5102
rect 2560 5098 2564 5102
rect 2596 5098 2600 5102
rect 2663 5098 2667 5102
rect 2162 5094 2166 5098
rect 2190 5094 2194 5098
rect 2205 5094 2209 5098
rect 2262 5094 2266 5098
rect 2280 5094 2284 5098
rect 2312 5094 2316 5098
rect 2153 5081 2157 5085
rect 2165 5081 2169 5085
rect 2173 5080 2177 5084
rect 2195 5081 2199 5085
rect 2208 5080 2212 5084
rect 2227 5080 2231 5084
rect 2129 5068 2133 5072
rect 2144 5068 2148 5072
rect 2246 5079 2250 5083
rect 2265 5083 2269 5087
rect 2285 5080 2289 5084
rect 2529 5090 2533 5094
rect 2670 5090 2674 5094
rect 2529 5081 2533 5085
rect 2553 5081 2557 5085
rect 2678 5083 2682 5087
rect 2545 5074 2549 5078
rect 2098 5054 2102 5058
rect 2162 5064 2166 5068
rect 2169 5061 2173 5065
rect 2189 5064 2193 5068
rect 2205 5064 2209 5068
rect 2215 5061 2219 5065
rect 2240 5061 2244 5065
rect 2262 5064 2266 5068
rect 2280 5064 2284 5068
rect 2287 5061 2291 5065
rect 2312 5064 2316 5068
rect 2354 5067 2360 5071
rect 2562 5067 2566 5071
rect 2612 5067 2616 5071
rect 2663 5067 2667 5071
rect 2390 5060 2396 5064
rect 2168 5054 2172 5058
rect 2233 5054 2237 5058
rect 2255 5054 2259 5058
rect 2286 5054 2290 5058
rect 2366 5054 2372 5058
rect 1600 5040 1604 5044
rect 1616 5040 1620 5044
rect 869 5034 873 5038
rect 919 5034 923 5038
rect 970 5034 974 5038
rect 1001 5034 1005 5038
rect 1051 5034 1055 5038
rect 1102 5034 1106 5038
rect 1133 5034 1137 5038
rect 1183 5034 1187 5038
rect 1234 5034 1238 5038
rect 1265 5034 1269 5038
rect 1315 5034 1319 5038
rect 1366 5034 1370 5038
rect 1409 5034 1415 5038
rect 1637 5038 1641 5044
rect 1653 5040 1657 5044
rect 2161 5047 2165 5051
rect 2189 5047 2193 5051
rect 2206 5047 2210 5051
rect 2262 5047 2266 5051
rect 2279 5047 2283 5051
rect 2313 5047 2317 5051
rect 2402 5047 2408 5051
rect 2562 5053 2566 5057
rect 2606 5053 2610 5057
rect 2626 5053 2630 5057
rect 2663 5051 2667 5055
rect 1674 5040 1678 5044
rect 1661 5034 1665 5038
rect 1695 5038 1699 5044
rect 1711 5040 1715 5044
rect 2545 5040 2549 5044
rect 2561 5040 2565 5044
rect 1814 5034 1818 5038
rect 1864 5034 1868 5038
rect 1915 5034 1919 5038
rect 1946 5034 1950 5038
rect 1996 5034 2000 5038
rect 2047 5034 2051 5038
rect 2078 5034 2082 5038
rect 2128 5034 2132 5038
rect 2179 5034 2183 5038
rect 2210 5034 2214 5038
rect 2260 5034 2264 5038
rect 2311 5034 2315 5038
rect 2354 5034 2360 5038
rect 1445 5027 1451 5031
rect 852 5015 856 5019
rect 869 5020 873 5024
rect 913 5020 917 5024
rect 933 5020 937 5024
rect 970 5018 974 5022
rect 852 5007 856 5011
rect 868 5007 872 5011
rect 889 5005 893 5011
rect 905 5007 909 5011
rect 984 5015 988 5019
rect 1001 5020 1005 5024
rect 1045 5020 1049 5024
rect 1065 5020 1069 5024
rect 1102 5018 1106 5022
rect 1133 5020 1137 5024
rect 1177 5020 1181 5024
rect 1197 5020 1201 5024
rect 1234 5018 1238 5022
rect 1265 5020 1269 5024
rect 1309 5020 1313 5024
rect 1329 5020 1333 5024
rect 1366 5018 1370 5022
rect 1600 5025 1604 5031
rect 1616 5025 1620 5031
rect 1653 5025 1657 5031
rect 1637 5021 1641 5025
rect 1661 5025 1665 5029
rect 1674 5025 1678 5031
rect 1711 5025 1715 5031
rect 1733 5030 1737 5034
rect 2582 5038 2586 5044
rect 2598 5040 2602 5044
rect 2619 5040 2623 5044
rect 2606 5034 2610 5038
rect 2640 5038 2644 5044
rect 2656 5040 2660 5044
rect 2390 5027 2396 5031
rect 1695 5021 1699 5025
rect 926 5007 930 5011
rect 913 5001 917 5005
rect 947 5005 951 5011
rect 963 5007 967 5011
rect 984 5007 988 5011
rect 1000 5007 1004 5011
rect 852 4992 856 4996
rect 868 4992 872 4998
rect 905 4992 909 4998
rect 889 4988 893 4992
rect 913 4992 917 4996
rect 926 4992 930 4998
rect 963 4992 967 4998
rect 976 4997 980 5001
rect 1021 5005 1025 5011
rect 1037 5007 1041 5011
rect 1058 5007 1062 5011
rect 1045 5001 1049 5005
rect 1079 5005 1083 5011
rect 1095 5007 1099 5011
rect 1116 5007 1120 5011
rect 1132 5007 1136 5011
rect 984 4992 988 4996
rect 1000 4992 1004 4998
rect 1037 4992 1041 4998
rect 947 4988 951 4992
rect 1021 4988 1025 4992
rect 1045 4992 1049 4996
rect 1058 4992 1062 4998
rect 1095 4992 1099 4998
rect 1108 4997 1112 5001
rect 1153 5005 1157 5011
rect 1169 5007 1173 5011
rect 1190 5007 1194 5011
rect 1177 5001 1181 5005
rect 1211 5005 1215 5011
rect 1227 5007 1231 5011
rect 1248 5007 1252 5011
rect 1264 5007 1268 5011
rect 1116 4992 1120 4996
rect 1132 4992 1136 4998
rect 1169 4992 1173 4998
rect 1079 4988 1083 4992
rect 1153 4988 1157 4992
rect 1177 4992 1181 4996
rect 1190 4992 1194 4998
rect 1227 4992 1231 4998
rect 1240 4997 1244 5001
rect 1285 5005 1289 5011
rect 1301 5007 1305 5011
rect 1322 5007 1326 5011
rect 1309 5001 1313 5005
rect 1343 5005 1347 5011
rect 1359 5007 1363 5011
rect 1615 5010 1619 5014
rect 1668 5010 1672 5014
rect 1718 5010 1722 5014
rect 1797 5015 1801 5019
rect 1814 5020 1818 5024
rect 1858 5020 1862 5024
rect 1878 5020 1882 5024
rect 1915 5018 1919 5022
rect 1797 5007 1801 5011
rect 1813 5007 1817 5011
rect 1457 5003 1463 5007
rect 1248 4992 1252 4996
rect 1264 4992 1268 4998
rect 1301 4992 1305 4998
rect 1211 4988 1215 4992
rect 1285 4988 1289 4992
rect 1309 4992 1313 4996
rect 1322 4992 1326 4998
rect 1359 4992 1363 4998
rect 1372 4997 1376 5001
rect 1834 5005 1838 5011
rect 1850 5007 1854 5011
rect 1929 5015 1933 5019
rect 1946 5020 1950 5024
rect 1990 5020 1994 5024
rect 2010 5020 2014 5024
rect 2047 5018 2051 5022
rect 2078 5020 2082 5024
rect 2122 5020 2126 5024
rect 2142 5020 2146 5024
rect 2179 5018 2183 5022
rect 2210 5020 2214 5024
rect 2254 5020 2258 5024
rect 2274 5020 2278 5024
rect 2311 5018 2315 5022
rect 2545 5025 2549 5031
rect 2561 5025 2565 5031
rect 2598 5025 2602 5031
rect 2582 5021 2586 5025
rect 2606 5025 2610 5029
rect 2619 5025 2623 5031
rect 2656 5025 2660 5031
rect 2678 5030 2682 5034
rect 2640 5021 2644 5025
rect 1871 5007 1875 5011
rect 1858 5001 1862 5005
rect 1892 5005 1896 5011
rect 1908 5007 1912 5011
rect 1929 5007 1933 5011
rect 1945 5007 1949 5011
rect 1397 4996 1403 5000
rect 1615 4996 1619 5000
rect 1682 4996 1686 5000
rect 1718 4996 1722 5000
rect 1797 4992 1801 4996
rect 1813 4992 1817 4998
rect 1850 4992 1854 4998
rect 1343 4988 1347 4992
rect 1834 4988 1838 4992
rect 1858 4992 1862 4996
rect 1871 4992 1875 4998
rect 1908 4992 1912 4998
rect 1921 4997 1925 5001
rect 1966 5005 1970 5011
rect 1982 5007 1986 5011
rect 2003 5007 2007 5011
rect 1990 5001 1994 5005
rect 2024 5005 2028 5011
rect 2040 5007 2044 5011
rect 2061 5007 2065 5011
rect 2077 5007 2081 5011
rect 1929 4992 1933 4996
rect 1945 4992 1949 4998
rect 1982 4992 1986 4998
rect 1892 4988 1896 4992
rect 1966 4988 1970 4992
rect 1990 4992 1994 4996
rect 2003 4992 2007 4998
rect 2040 4992 2044 4998
rect 2053 4997 2057 5001
rect 2098 5005 2102 5011
rect 2114 5007 2118 5011
rect 2135 5007 2139 5011
rect 2122 5001 2126 5005
rect 2156 5005 2160 5011
rect 2172 5007 2176 5011
rect 2193 5007 2197 5011
rect 2209 5007 2213 5011
rect 2061 4992 2065 4996
rect 2077 4992 2081 4998
rect 2114 4992 2118 4998
rect 2024 4988 2028 4992
rect 2098 4988 2102 4992
rect 2122 4992 2126 4996
rect 2135 4992 2139 4998
rect 2172 4992 2176 4998
rect 2185 4997 2189 5001
rect 2230 5005 2234 5011
rect 2246 5007 2250 5011
rect 2267 5007 2271 5011
rect 2254 5001 2258 5005
rect 2288 5005 2292 5011
rect 2304 5007 2308 5011
rect 2560 5010 2564 5014
rect 2613 5010 2617 5014
rect 2663 5010 2667 5014
rect 2402 5003 2408 5007
rect 4484 5004 4488 5008
rect 4494 5004 4498 5008
rect 4504 5004 4508 5008
rect 2193 4992 2197 4996
rect 2209 4992 2213 4998
rect 2246 4992 2250 4998
rect 2156 4988 2160 4992
rect 2230 4988 2234 4992
rect 2254 4992 2258 4996
rect 2267 4992 2271 4998
rect 2304 4992 2308 4998
rect 2317 4997 2321 5001
rect 2342 4996 2348 5000
rect 2560 4996 2564 5000
rect 2627 4996 2631 5000
rect 2663 4996 2667 5000
rect 4484 4999 4488 5003
rect 4494 4999 4498 5003
rect 4504 4999 4508 5003
rect 4484 4994 4488 4998
rect 4494 4994 4498 4998
rect 4504 4994 4508 4998
rect 2288 4988 2292 4992
rect 4484 4989 4488 4993
rect 4494 4989 4498 4993
rect 4504 4989 4508 4993
rect 4530 5004 4534 5008
rect 4540 5004 4544 5008
rect 4550 5004 4554 5008
rect 4530 4999 4534 5003
rect 4540 4999 4544 5003
rect 4550 4999 4554 5003
rect 4530 4994 4534 4998
rect 4540 4994 4544 4998
rect 4550 4994 4554 4998
rect 4530 4989 4534 4993
rect 4540 4989 4544 4993
rect 4550 4989 4554 4993
rect 867 4977 871 4981
rect 920 4977 924 4981
rect 970 4977 974 4981
rect 999 4977 1003 4981
rect 1052 4977 1056 4981
rect 1102 4977 1106 4981
rect 1131 4977 1135 4981
rect 1184 4977 1188 4981
rect 1234 4977 1238 4981
rect 1263 4977 1267 4981
rect 1316 4977 1320 4981
rect 1366 4977 1370 4981
rect 1812 4977 1816 4981
rect 1865 4977 1869 4981
rect 1915 4977 1919 4981
rect 1944 4977 1948 4981
rect 1997 4977 2001 4981
rect 2047 4977 2051 4981
rect 2076 4977 2080 4981
rect 2129 4977 2133 4981
rect 2179 4977 2183 4981
rect 2208 4977 2212 4981
rect 2261 4977 2265 4981
rect 2311 4977 2315 4981
rect 1457 4970 1463 4974
rect 2402 4970 2408 4974
rect 867 4963 871 4967
rect 934 4963 938 4967
rect 970 4963 974 4967
rect 999 4963 1003 4967
rect 1066 4963 1070 4967
rect 1102 4963 1106 4967
rect 1131 4963 1135 4967
rect 1198 4963 1202 4967
rect 1234 4963 1238 4967
rect 1263 4963 1267 4967
rect 1330 4963 1334 4967
rect 1366 4963 1370 4967
rect 1397 4963 1403 4967
rect 1812 4963 1816 4967
rect 1879 4963 1883 4967
rect 1915 4963 1919 4967
rect 1944 4963 1948 4967
rect 2011 4963 2015 4967
rect 2047 4963 2051 4967
rect 2076 4963 2080 4967
rect 2143 4963 2147 4967
rect 2179 4963 2183 4967
rect 2208 4963 2212 4967
rect 2275 4963 2279 4967
rect 2311 4963 2315 4967
rect 2342 4963 2348 4967
rect 1457 4930 1463 4934
rect 2670 4932 2674 4936
rect 3836 4932 3844 4936
rect 1445 4922 1451 4926
rect 1433 4914 1439 4918
rect 1421 4906 1427 4910
rect 1409 4898 1415 4902
rect 1756 4876 1761 4880
rect 2146 4876 2151 4880
rect 618 4868 622 4872
rect 628 4868 632 4872
rect 638 4868 642 4872
rect 618 4863 622 4867
rect 628 4863 632 4867
rect 638 4863 642 4867
rect 618 4858 622 4862
rect 628 4858 632 4862
rect 638 4858 642 4862
rect 618 4853 622 4857
rect 628 4853 632 4857
rect 638 4853 642 4857
rect 664 4868 668 4872
rect 674 4868 678 4872
rect 684 4868 688 4872
rect 664 4863 668 4867
rect 674 4863 678 4867
rect 684 4863 688 4867
rect 1745 4866 1749 4870
rect 2119 4866 2132 4870
rect 664 4858 668 4862
rect 674 4858 678 4862
rect 684 4858 688 4862
rect 664 4853 668 4857
rect 674 4853 678 4857
rect 684 4853 688 4857
rect 1385 4858 1391 4862
rect 2330 4858 2336 4862
rect 618 4839 622 4843
rect 628 4839 632 4843
rect 638 4839 642 4843
rect 618 4834 622 4838
rect 628 4834 632 4838
rect 638 4834 642 4838
rect 618 4829 622 4833
rect 628 4829 632 4833
rect 638 4829 642 4833
rect 618 4824 622 4828
rect 628 4824 632 4828
rect 638 4824 642 4828
rect 664 4839 668 4843
rect 674 4839 678 4843
rect 684 4839 688 4843
rect 664 4834 668 4838
rect 674 4834 678 4838
rect 684 4834 688 4838
rect 664 4829 668 4833
rect 674 4829 678 4833
rect 684 4829 688 4833
rect 664 4824 668 4828
rect 674 4824 678 4828
rect 684 4824 688 4828
rect 618 4810 622 4814
rect 628 4810 632 4814
rect 638 4810 642 4814
rect 618 4805 622 4809
rect 628 4805 632 4809
rect 638 4805 642 4809
rect 618 4800 622 4804
rect 628 4800 632 4804
rect 638 4800 642 4804
rect 618 4795 622 4799
rect 628 4795 632 4799
rect 638 4795 642 4799
rect 664 4810 668 4814
rect 674 4810 678 4814
rect 684 4810 688 4814
rect 664 4805 668 4809
rect 674 4805 678 4809
rect 684 4805 688 4809
rect 664 4800 668 4804
rect 674 4800 678 4804
rect 684 4800 688 4804
rect 664 4795 668 4799
rect 674 4795 678 4799
rect 684 4795 688 4799
rect 618 4781 622 4785
rect 628 4781 632 4785
rect 638 4781 642 4785
rect 618 4776 622 4780
rect 628 4776 632 4780
rect 638 4776 642 4780
rect 618 4771 622 4775
rect 628 4771 632 4775
rect 638 4771 642 4775
rect 618 4766 622 4770
rect 628 4766 632 4770
rect 638 4766 642 4770
rect 664 4781 668 4785
rect 674 4781 678 4785
rect 684 4781 688 4785
rect 664 4776 668 4780
rect 674 4776 678 4780
rect 684 4776 688 4780
rect 664 4771 668 4775
rect 674 4771 678 4775
rect 684 4771 688 4775
rect 664 4766 668 4770
rect 674 4766 678 4770
rect 684 4766 688 4770
rect 618 4752 622 4756
rect 628 4752 632 4756
rect 638 4752 642 4756
rect 618 4747 622 4751
rect 628 4747 632 4751
rect 638 4747 642 4751
rect 618 4742 622 4746
rect 628 4742 632 4746
rect 638 4742 642 4746
rect 618 4737 622 4741
rect 628 4737 632 4741
rect 638 4737 642 4741
rect 664 4752 668 4756
rect 674 4752 678 4756
rect 684 4752 688 4756
rect 664 4747 668 4751
rect 674 4747 678 4751
rect 684 4747 688 4751
rect 664 4742 668 4746
rect 674 4742 678 4746
rect 684 4742 688 4746
rect 664 4737 668 4741
rect 674 4737 678 4741
rect 684 4737 688 4741
rect 1457 4850 1463 4854
rect 1482 4851 1537 4855
rect 2402 4851 2408 4855
rect 1445 4843 1451 4847
rect 1790 4843 1845 4847
rect 2390 4843 2396 4848
rect 1433 4835 1439 4839
rect 2378 4835 2384 4839
rect 1421 4828 1427 4832
rect 2366 4828 2372 4832
rect 1409 4821 1415 4825
rect 2354 4821 2360 4825
rect 1397 4813 1403 4817
rect 2342 4813 2348 4817
rect 4484 4811 4488 4815
rect 4494 4811 4498 4815
rect 4504 4811 4508 4815
rect 4484 4806 4488 4810
rect 4494 4806 4498 4810
rect 4504 4806 4508 4810
rect 4484 4801 4488 4805
rect 4494 4801 4498 4805
rect 4504 4801 4508 4805
rect 4484 4796 4488 4800
rect 4494 4796 4498 4800
rect 4504 4796 4508 4800
rect 4530 4811 4534 4815
rect 4540 4811 4544 4815
rect 4550 4811 4554 4815
rect 4530 4806 4534 4810
rect 4540 4806 4544 4810
rect 4550 4806 4554 4810
rect 4530 4801 4534 4805
rect 4540 4801 4544 4805
rect 4550 4801 4554 4805
rect 4530 4796 4534 4800
rect 4540 4796 4544 4800
rect 4550 4796 4554 4800
rect 4484 4785 4488 4789
rect 4494 4785 4498 4789
rect 4504 4785 4508 4789
rect 4484 4780 4488 4784
rect 4494 4780 4498 4784
rect 4504 4780 4508 4784
rect 4484 4775 4488 4779
rect 4494 4775 4498 4779
rect 4504 4775 4508 4779
rect 4484 4770 4488 4774
rect 4494 4770 4498 4774
rect 4504 4770 4508 4774
rect 4530 4785 4534 4789
rect 4540 4785 4544 4789
rect 4550 4785 4554 4789
rect 4530 4780 4534 4784
rect 4540 4780 4544 4784
rect 4550 4780 4554 4784
rect 4530 4775 4534 4779
rect 4540 4775 4544 4779
rect 4550 4775 4554 4779
rect 4530 4770 4534 4774
rect 4540 4770 4544 4774
rect 4550 4770 4554 4774
rect 4484 4759 4488 4763
rect 4494 4759 4498 4763
rect 4504 4759 4508 4763
rect 4484 4754 4488 4758
rect 4494 4754 4498 4758
rect 4504 4754 4508 4758
rect 4484 4749 4488 4753
rect 4494 4749 4498 4753
rect 4504 4749 4508 4753
rect 4484 4744 4488 4748
rect 4494 4744 4498 4748
rect 4504 4744 4508 4748
rect 4530 4759 4534 4763
rect 4540 4759 4544 4763
rect 4550 4759 4554 4763
rect 4530 4754 4534 4758
rect 4540 4754 4544 4758
rect 4550 4754 4554 4758
rect 4530 4749 4534 4753
rect 4540 4749 4544 4753
rect 4550 4749 4554 4753
rect 4530 4744 4534 4748
rect 4540 4744 4544 4748
rect 4550 4744 4554 4748
rect 757 4619 761 4623
rect 762 4619 766 4623
rect 767 4619 771 4623
rect 772 4619 776 4623
rect 757 4609 761 4613
rect 762 4609 766 4613
rect 767 4609 771 4613
rect 772 4609 776 4613
rect 757 4599 761 4603
rect 762 4599 766 4603
rect 767 4599 771 4603
rect 772 4599 776 4603
rect 783 4619 787 4623
rect 788 4619 792 4623
rect 793 4619 797 4623
rect 798 4619 802 4623
rect 783 4609 787 4613
rect 788 4609 792 4613
rect 793 4609 797 4613
rect 798 4609 802 4613
rect 783 4599 787 4603
rect 788 4599 792 4603
rect 793 4599 797 4603
rect 798 4599 802 4603
rect 809 4619 813 4623
rect 814 4619 818 4623
rect 819 4619 823 4623
rect 824 4619 828 4623
rect 809 4609 813 4613
rect 814 4609 818 4613
rect 819 4609 823 4613
rect 824 4609 828 4613
rect 809 4599 813 4603
rect 814 4599 818 4603
rect 819 4599 823 4603
rect 824 4599 828 4603
rect 835 4619 839 4623
rect 840 4619 844 4623
rect 845 4619 849 4623
rect 850 4619 854 4623
rect 835 4609 839 4613
rect 840 4609 844 4613
rect 845 4609 849 4613
rect 850 4609 854 4613
rect 835 4599 839 4603
rect 840 4599 844 4603
rect 845 4599 849 4603
rect 850 4599 854 4603
rect 861 4619 865 4623
rect 866 4619 870 4623
rect 871 4619 875 4623
rect 876 4619 880 4623
rect 861 4609 865 4613
rect 866 4609 870 4613
rect 871 4609 875 4613
rect 876 4609 880 4613
rect 861 4599 865 4603
rect 866 4599 870 4603
rect 871 4599 875 4603
rect 876 4599 880 4603
rect 1053 4619 1057 4623
rect 1058 4619 1062 4623
rect 1063 4619 1067 4623
rect 1068 4619 1072 4623
rect 1053 4609 1057 4613
rect 1058 4609 1062 4613
rect 1063 4609 1067 4613
rect 1068 4609 1072 4613
rect 1053 4599 1057 4603
rect 1058 4599 1062 4603
rect 1063 4599 1067 4603
rect 1068 4599 1072 4603
rect 1077 4597 1081 4601
rect 1082 4597 1086 4601
rect 1087 4597 1091 4601
rect 1092 4597 1096 4601
rect 1097 4597 1101 4601
rect 1102 4597 1106 4601
rect 1107 4597 1111 4601
rect 1112 4597 1116 4601
rect 1117 4597 1121 4601
rect 1122 4597 1126 4601
rect 1127 4597 1131 4601
rect 1077 4592 1081 4596
rect 1082 4592 1086 4596
rect 1087 4592 1091 4596
rect 1092 4592 1096 4596
rect 1097 4592 1101 4596
rect 1102 4592 1106 4596
rect 1107 4592 1111 4596
rect 1112 4592 1116 4596
rect 1117 4592 1121 4596
rect 1122 4592 1126 4596
rect 1127 4592 1131 4596
rect 757 4573 761 4577
rect 762 4573 766 4577
rect 767 4573 771 4577
rect 772 4573 776 4577
rect 757 4563 761 4567
rect 762 4563 766 4567
rect 767 4563 771 4567
rect 772 4563 776 4567
rect 757 4553 761 4557
rect 762 4553 766 4557
rect 767 4553 771 4557
rect 772 4553 776 4557
rect 783 4573 787 4577
rect 788 4573 792 4577
rect 793 4573 797 4577
rect 798 4573 802 4577
rect 783 4563 787 4567
rect 788 4563 792 4567
rect 793 4563 797 4567
rect 798 4563 802 4567
rect 783 4553 787 4557
rect 788 4553 792 4557
rect 793 4553 797 4557
rect 798 4553 802 4557
rect 809 4573 813 4577
rect 814 4573 818 4577
rect 819 4573 823 4577
rect 824 4573 828 4577
rect 809 4563 813 4567
rect 814 4563 818 4567
rect 819 4563 823 4567
rect 824 4563 828 4567
rect 809 4553 813 4557
rect 814 4553 818 4557
rect 819 4553 823 4557
rect 824 4553 828 4557
rect 835 4573 839 4577
rect 840 4573 844 4577
rect 845 4573 849 4577
rect 850 4573 854 4577
rect 835 4563 839 4567
rect 840 4563 844 4567
rect 845 4563 849 4567
rect 850 4563 854 4567
rect 835 4553 839 4557
rect 840 4553 844 4557
rect 845 4553 849 4557
rect 850 4553 854 4557
rect 861 4573 865 4577
rect 866 4573 870 4577
rect 871 4573 875 4577
rect 876 4573 880 4577
rect 861 4563 865 4567
rect 866 4563 870 4567
rect 871 4563 875 4567
rect 876 4563 880 4567
rect 861 4553 865 4557
rect 866 4553 870 4557
rect 871 4553 875 4557
rect 876 4553 880 4557
rect 1053 4573 1057 4577
rect 1058 4573 1062 4577
rect 1063 4573 1067 4577
rect 1068 4573 1072 4577
rect 1053 4563 1057 4567
rect 1058 4563 1062 4567
rect 1063 4563 1067 4567
rect 1068 4563 1072 4567
rect 1053 4553 1057 4557
rect 1058 4553 1062 4557
rect 1063 4553 1067 4557
rect 1068 4553 1072 4557
rect 1169 4531 1173 4535
rect 2670 4717 2675 4739
rect 2737 4717 2750 4739
rect 4484 4733 4488 4737
rect 4494 4733 4498 4737
rect 4504 4733 4508 4737
rect 4484 4728 4488 4732
rect 4494 4728 4498 4732
rect 4504 4728 4508 4732
rect 4484 4723 4488 4727
rect 4494 4723 4498 4727
rect 4504 4723 4508 4727
rect 1482 4705 1538 4710
rect 1362 4619 1366 4623
rect 1367 4619 1371 4623
rect 1372 4619 1376 4623
rect 1377 4619 1381 4623
rect 1362 4609 1366 4613
rect 1367 4609 1371 4613
rect 1372 4609 1376 4613
rect 1377 4609 1381 4613
rect 1362 4599 1366 4603
rect 1367 4599 1371 4603
rect 1372 4599 1376 4603
rect 1377 4599 1381 4603
rect 1386 4597 1390 4601
rect 1391 4597 1395 4601
rect 1396 4597 1400 4601
rect 1401 4597 1405 4601
rect 1406 4597 1410 4601
rect 1411 4597 1415 4601
rect 1416 4597 1420 4601
rect 1421 4597 1425 4601
rect 1426 4597 1430 4601
rect 1431 4597 1435 4601
rect 1436 4597 1440 4601
rect 1386 4592 1390 4596
rect 1391 4592 1395 4596
rect 1396 4592 1400 4596
rect 1401 4592 1405 4596
rect 1406 4592 1410 4596
rect 1411 4592 1415 4596
rect 1416 4592 1420 4596
rect 1421 4592 1425 4596
rect 1426 4592 1430 4596
rect 1431 4592 1435 4596
rect 1436 4592 1440 4596
rect 1327 4574 1331 4578
rect 1332 4574 1336 4578
rect 1327 4569 1331 4573
rect 1332 4569 1336 4573
rect 1327 4564 1331 4568
rect 1332 4564 1336 4568
rect 1327 4559 1331 4563
rect 1332 4559 1336 4563
rect 1327 4554 1331 4558
rect 1332 4554 1336 4558
rect 1327 4549 1331 4553
rect 1332 4549 1336 4553
rect 1362 4573 1366 4577
rect 1367 4573 1371 4577
rect 1372 4573 1376 4577
rect 1377 4573 1381 4577
rect 1362 4563 1366 4567
rect 1367 4563 1371 4567
rect 1372 4563 1376 4567
rect 1377 4563 1381 4567
rect 1362 4553 1366 4557
rect 1367 4553 1371 4557
rect 1372 4553 1376 4557
rect 1377 4553 1381 4557
rect 1327 4544 1331 4548
rect 1332 4544 1336 4548
rect 1327 4539 1331 4543
rect 1332 4539 1336 4543
rect 1227 4531 1231 4535
rect 1327 4534 1331 4538
rect 1332 4534 1336 4538
rect 1327 4529 1331 4533
rect 1332 4529 1336 4533
rect 1327 4524 1331 4528
rect 1332 4524 1336 4528
rect 1169 4515 1173 4519
rect 1327 4519 1331 4523
rect 1332 4519 1336 4523
rect 1227 4515 1231 4519
rect 1327 4514 1331 4518
rect 1332 4514 1336 4518
rect 1169 4499 1173 4503
rect 1227 4499 1231 4503
rect 1169 4483 1173 4487
rect 1227 4483 1231 4487
rect 1793 4704 1845 4708
rect 1810 4649 1814 4653
rect 1815 4649 1819 4653
rect 1810 4644 1814 4648
rect 1815 4644 1819 4648
rect 1810 4639 1814 4643
rect 1815 4639 1819 4643
rect 1810 4634 1814 4638
rect 1815 4634 1819 4638
rect 1810 4629 1814 4633
rect 1815 4629 1819 4633
rect 2119 4703 2132 4707
rect 2146 4705 2151 4709
rect 1671 4619 1675 4623
rect 1676 4619 1680 4623
rect 1681 4619 1685 4623
rect 1686 4619 1690 4623
rect 1671 4609 1675 4613
rect 1676 4609 1680 4613
rect 1681 4609 1685 4613
rect 1686 4609 1690 4613
rect 1671 4599 1675 4603
rect 1676 4599 1680 4603
rect 1681 4599 1685 4603
rect 1686 4599 1690 4603
rect 1810 4624 1814 4628
rect 1815 4624 1819 4628
rect 1810 4619 1814 4623
rect 1815 4619 1819 4623
rect 1810 4614 1814 4618
rect 1815 4614 1819 4618
rect 1810 4609 1814 4613
rect 1815 4609 1819 4613
rect 1810 4604 1814 4608
rect 1815 4604 1819 4608
rect 1695 4597 1699 4601
rect 1700 4597 1704 4601
rect 1705 4597 1709 4601
rect 1710 4597 1714 4601
rect 1715 4597 1719 4601
rect 1720 4597 1724 4601
rect 1725 4597 1729 4601
rect 1730 4597 1734 4601
rect 1735 4597 1739 4601
rect 1740 4597 1744 4601
rect 1745 4597 1749 4601
rect 1695 4592 1699 4596
rect 1700 4592 1704 4596
rect 1705 4592 1709 4596
rect 1710 4592 1714 4596
rect 1715 4592 1719 4596
rect 1720 4592 1724 4596
rect 1725 4592 1729 4596
rect 1730 4592 1734 4596
rect 1735 4592 1739 4596
rect 1740 4592 1744 4596
rect 1745 4592 1749 4596
rect 1501 4569 1505 4573
rect 1506 4569 1510 4573
rect 1501 4564 1505 4568
rect 1506 4564 1510 4568
rect 1501 4559 1505 4563
rect 1506 4559 1510 4563
rect 1501 4554 1505 4558
rect 1506 4554 1510 4558
rect 1501 4549 1505 4553
rect 1506 4549 1510 4553
rect 1501 4544 1505 4548
rect 1506 4544 1510 4548
rect 1501 4539 1505 4543
rect 1506 4539 1510 4543
rect 1501 4534 1505 4538
rect 1506 4534 1510 4538
rect 1501 4529 1505 4533
rect 1506 4529 1510 4533
rect 1501 4524 1505 4528
rect 1506 4524 1510 4528
rect 1501 4519 1505 4523
rect 1506 4519 1510 4523
rect 1087 4462 1091 4466
rect 1094 4462 1098 4466
rect 1099 4462 1103 4466
rect 1104 4462 1108 4466
rect 1109 4462 1113 4466
rect 1114 4462 1118 4466
rect 1119 4462 1123 4466
rect 1124 4462 1128 4466
rect 1129 4462 1133 4466
rect 1134 4462 1138 4466
rect 1139 4462 1143 4466
rect 1144 4462 1148 4466
rect 1151 4462 1155 4466
rect 1104 4446 1108 4450
rect 1114 4446 1118 4450
rect 1124 4446 1128 4450
rect 1134 4446 1138 4450
rect 1099 4441 1103 4445
rect 1109 4441 1113 4445
rect 1119 4441 1123 4445
rect 1129 4441 1133 4445
rect 1139 4441 1143 4445
rect 1104 4436 1108 4440
rect 1114 4436 1118 4440
rect 1124 4436 1128 4440
rect 1134 4436 1138 4440
rect 1099 4431 1103 4435
rect 1109 4431 1113 4435
rect 1119 4431 1123 4435
rect 1129 4431 1133 4435
rect 1139 4431 1143 4435
rect 1104 4426 1108 4430
rect 1114 4426 1118 4430
rect 1124 4426 1128 4430
rect 1134 4426 1138 4430
rect 1099 4421 1103 4425
rect 1109 4421 1113 4425
rect 1119 4421 1123 4425
rect 1129 4421 1133 4425
rect 1139 4421 1143 4425
rect 1104 4416 1108 4420
rect 1114 4416 1118 4420
rect 1124 4416 1128 4420
rect 1134 4416 1138 4420
rect 1099 4411 1103 4415
rect 1109 4411 1113 4415
rect 1119 4411 1123 4415
rect 1129 4411 1133 4415
rect 1139 4411 1143 4415
rect 1104 4406 1108 4410
rect 1114 4406 1118 4410
rect 1124 4406 1128 4410
rect 1134 4406 1138 4410
rect 1099 4401 1103 4405
rect 1109 4401 1113 4405
rect 1119 4401 1123 4405
rect 1129 4401 1133 4405
rect 1139 4401 1143 4405
rect 1104 4396 1108 4400
rect 1114 4396 1118 4400
rect 1124 4396 1128 4400
rect 1134 4396 1138 4400
rect 1099 4391 1103 4395
rect 1109 4391 1113 4395
rect 1119 4391 1123 4395
rect 1129 4391 1133 4395
rect 1139 4391 1143 4395
rect 1104 4386 1108 4390
rect 1114 4386 1118 4390
rect 1124 4386 1128 4390
rect 1134 4386 1138 4390
rect 1099 4381 1103 4385
rect 1109 4381 1113 4385
rect 1119 4381 1123 4385
rect 1129 4381 1133 4385
rect 1139 4381 1143 4385
rect 1104 4376 1108 4380
rect 1114 4376 1118 4380
rect 1124 4376 1128 4380
rect 1134 4376 1138 4380
rect 1099 4371 1103 4375
rect 1109 4371 1113 4375
rect 1119 4371 1123 4375
rect 1129 4371 1133 4375
rect 1139 4371 1143 4375
rect 1104 4366 1108 4370
rect 1114 4366 1118 4370
rect 1124 4366 1128 4370
rect 1134 4366 1138 4370
rect 1099 4361 1103 4365
rect 1109 4361 1113 4365
rect 1119 4361 1123 4365
rect 1129 4361 1133 4365
rect 1139 4361 1143 4365
rect 1247 4462 1251 4466
rect 1254 4462 1258 4466
rect 1259 4462 1263 4466
rect 1264 4462 1268 4466
rect 1269 4462 1273 4466
rect 1274 4462 1278 4466
rect 1279 4462 1283 4466
rect 1284 4462 1288 4466
rect 1289 4462 1293 4466
rect 1294 4462 1298 4466
rect 1299 4462 1303 4466
rect 1304 4462 1308 4466
rect 1311 4462 1315 4466
rect 1264 4446 1268 4450
rect 1274 4446 1278 4450
rect 1284 4446 1288 4450
rect 1294 4446 1298 4450
rect 1259 4441 1263 4445
rect 1269 4441 1273 4445
rect 1279 4441 1283 4445
rect 1289 4441 1293 4445
rect 1299 4441 1303 4445
rect 1264 4436 1268 4440
rect 1274 4436 1278 4440
rect 1284 4436 1288 4440
rect 1294 4436 1298 4440
rect 1259 4431 1263 4435
rect 1269 4431 1273 4435
rect 1279 4431 1283 4435
rect 1289 4431 1293 4435
rect 1299 4431 1303 4435
rect 1264 4426 1268 4430
rect 1274 4426 1278 4430
rect 1284 4426 1288 4430
rect 1294 4426 1298 4430
rect 1259 4421 1263 4425
rect 1269 4421 1273 4425
rect 1279 4421 1283 4425
rect 1289 4421 1293 4425
rect 1299 4421 1303 4425
rect 1264 4416 1268 4420
rect 1274 4416 1278 4420
rect 1284 4416 1288 4420
rect 1294 4416 1298 4420
rect 1259 4411 1263 4415
rect 1269 4411 1273 4415
rect 1279 4411 1283 4415
rect 1289 4411 1293 4415
rect 1299 4411 1303 4415
rect 1264 4406 1268 4410
rect 1274 4406 1278 4410
rect 1284 4406 1288 4410
rect 1294 4406 1298 4410
rect 1259 4401 1263 4405
rect 1269 4401 1273 4405
rect 1279 4401 1283 4405
rect 1289 4401 1293 4405
rect 1299 4401 1303 4405
rect 1264 4396 1268 4400
rect 1274 4396 1278 4400
rect 1284 4396 1288 4400
rect 1294 4396 1298 4400
rect 1259 4391 1263 4395
rect 1269 4391 1273 4395
rect 1279 4391 1283 4395
rect 1289 4391 1293 4395
rect 1299 4391 1303 4395
rect 1264 4386 1268 4390
rect 1274 4386 1278 4390
rect 1284 4386 1288 4390
rect 1294 4386 1298 4390
rect 1259 4381 1263 4385
rect 1269 4381 1273 4385
rect 1279 4381 1283 4385
rect 1289 4381 1293 4385
rect 1299 4381 1303 4385
rect 1264 4376 1268 4380
rect 1274 4376 1278 4380
rect 1284 4376 1288 4380
rect 1294 4376 1298 4380
rect 1259 4371 1263 4375
rect 1269 4371 1273 4375
rect 1279 4371 1283 4375
rect 1289 4371 1293 4375
rect 1299 4371 1303 4375
rect 1264 4366 1268 4370
rect 1274 4366 1278 4370
rect 1284 4366 1288 4370
rect 1294 4366 1298 4370
rect 1259 4361 1263 4365
rect 1269 4361 1273 4365
rect 1279 4361 1283 4365
rect 1289 4361 1293 4365
rect 1299 4361 1303 4365
rect 1396 4462 1400 4466
rect 1403 4462 1407 4466
rect 1408 4462 1412 4466
rect 1413 4462 1417 4466
rect 1418 4462 1422 4466
rect 1423 4462 1427 4466
rect 1428 4462 1432 4466
rect 1433 4462 1437 4466
rect 1438 4462 1442 4466
rect 1443 4462 1447 4466
rect 1448 4462 1452 4466
rect 1453 4462 1457 4466
rect 1460 4462 1464 4466
rect 1413 4446 1417 4450
rect 1423 4446 1427 4450
rect 1433 4446 1437 4450
rect 1443 4446 1447 4450
rect 1408 4441 1412 4445
rect 1418 4441 1422 4445
rect 1428 4441 1432 4445
rect 1438 4441 1442 4445
rect 1448 4441 1452 4445
rect 1413 4436 1417 4440
rect 1423 4436 1427 4440
rect 1433 4436 1437 4440
rect 1443 4436 1447 4440
rect 1408 4431 1412 4435
rect 1418 4431 1422 4435
rect 1428 4431 1432 4435
rect 1438 4431 1442 4435
rect 1448 4431 1452 4435
rect 1413 4426 1417 4430
rect 1423 4426 1427 4430
rect 1433 4426 1437 4430
rect 1443 4426 1447 4430
rect 1408 4421 1412 4425
rect 1418 4421 1422 4425
rect 1428 4421 1432 4425
rect 1438 4421 1442 4425
rect 1448 4421 1452 4425
rect 1413 4416 1417 4420
rect 1423 4416 1427 4420
rect 1433 4416 1437 4420
rect 1443 4416 1447 4420
rect 1408 4411 1412 4415
rect 1418 4411 1422 4415
rect 1428 4411 1432 4415
rect 1438 4411 1442 4415
rect 1448 4411 1452 4415
rect 1413 4406 1417 4410
rect 1423 4406 1427 4410
rect 1433 4406 1437 4410
rect 1443 4406 1447 4410
rect 1408 4401 1412 4405
rect 1418 4401 1422 4405
rect 1428 4401 1432 4405
rect 1438 4401 1442 4405
rect 1448 4401 1452 4405
rect 1413 4396 1417 4400
rect 1423 4396 1427 4400
rect 1433 4396 1437 4400
rect 1443 4396 1447 4400
rect 1408 4391 1412 4395
rect 1418 4391 1422 4395
rect 1428 4391 1432 4395
rect 1438 4391 1442 4395
rect 1448 4391 1452 4395
rect 1413 4386 1417 4390
rect 1423 4386 1427 4390
rect 1433 4386 1437 4390
rect 1443 4386 1447 4390
rect 1408 4381 1412 4385
rect 1418 4381 1422 4385
rect 1428 4381 1432 4385
rect 1438 4381 1442 4385
rect 1448 4381 1452 4385
rect 1413 4376 1417 4380
rect 1423 4376 1427 4380
rect 1433 4376 1437 4380
rect 1443 4376 1447 4380
rect 1408 4371 1412 4375
rect 1418 4371 1422 4375
rect 1428 4371 1432 4375
rect 1438 4371 1442 4375
rect 1448 4371 1452 4375
rect 1413 4366 1417 4370
rect 1423 4366 1427 4370
rect 1433 4366 1437 4370
rect 1443 4366 1447 4370
rect 1408 4361 1412 4365
rect 1418 4361 1422 4365
rect 1428 4361 1432 4365
rect 1438 4361 1442 4365
rect 1448 4361 1452 4365
rect 1636 4574 1640 4578
rect 1641 4574 1645 4578
rect 1636 4569 1640 4573
rect 1641 4569 1645 4573
rect 1636 4564 1640 4568
rect 1641 4564 1645 4568
rect 1636 4559 1640 4563
rect 1641 4559 1645 4563
rect 1636 4554 1640 4558
rect 1641 4554 1645 4558
rect 1636 4549 1640 4553
rect 1641 4549 1645 4553
rect 1671 4573 1675 4577
rect 1676 4573 1680 4577
rect 1681 4573 1685 4577
rect 1686 4573 1690 4577
rect 1671 4563 1675 4567
rect 1676 4563 1680 4567
rect 1681 4563 1685 4567
rect 1686 4563 1690 4567
rect 1671 4553 1675 4557
rect 1676 4553 1680 4557
rect 1681 4553 1685 4557
rect 1686 4553 1690 4557
rect 1636 4544 1640 4548
rect 1641 4544 1645 4548
rect 1636 4539 1640 4543
rect 1641 4539 1645 4543
rect 1636 4534 1640 4538
rect 1641 4534 1645 4538
rect 1636 4529 1640 4533
rect 1641 4529 1645 4533
rect 1636 4524 1640 4528
rect 1641 4524 1645 4528
rect 1636 4519 1640 4523
rect 1641 4519 1645 4523
rect 1636 4514 1640 4518
rect 1641 4514 1645 4518
rect 1810 4599 1814 4603
rect 1815 4599 1819 4603
rect 1556 4462 1560 4466
rect 1563 4462 1567 4466
rect 1568 4462 1572 4466
rect 1573 4462 1577 4466
rect 1578 4462 1582 4466
rect 1583 4462 1587 4466
rect 1588 4462 1592 4466
rect 1593 4462 1597 4466
rect 1598 4462 1602 4466
rect 1603 4462 1607 4466
rect 1608 4462 1612 4466
rect 1613 4462 1617 4466
rect 1620 4462 1624 4466
rect 1573 4446 1577 4450
rect 1583 4446 1587 4450
rect 1593 4446 1597 4450
rect 1603 4446 1607 4450
rect 1568 4441 1572 4445
rect 1578 4441 1582 4445
rect 1588 4441 1592 4445
rect 1598 4441 1602 4445
rect 1608 4441 1612 4445
rect 1573 4436 1577 4440
rect 1583 4436 1587 4440
rect 1593 4436 1597 4440
rect 1603 4436 1607 4440
rect 1568 4431 1572 4435
rect 1578 4431 1582 4435
rect 1588 4431 1592 4435
rect 1598 4431 1602 4435
rect 1608 4431 1612 4435
rect 1573 4426 1577 4430
rect 1583 4426 1587 4430
rect 1593 4426 1597 4430
rect 1603 4426 1607 4430
rect 1568 4421 1572 4425
rect 1578 4421 1582 4425
rect 1588 4421 1592 4425
rect 1598 4421 1602 4425
rect 1608 4421 1612 4425
rect 1573 4416 1577 4420
rect 1583 4416 1587 4420
rect 1593 4416 1597 4420
rect 1603 4416 1607 4420
rect 1568 4411 1572 4415
rect 1578 4411 1582 4415
rect 1588 4411 1592 4415
rect 1598 4411 1602 4415
rect 1608 4411 1612 4415
rect 1573 4406 1577 4410
rect 1583 4406 1587 4410
rect 1593 4406 1597 4410
rect 1603 4406 1607 4410
rect 1568 4401 1572 4405
rect 1578 4401 1582 4405
rect 1588 4401 1592 4405
rect 1598 4401 1602 4405
rect 1608 4401 1612 4405
rect 1573 4396 1577 4400
rect 1583 4396 1587 4400
rect 1593 4396 1597 4400
rect 1603 4396 1607 4400
rect 1568 4391 1572 4395
rect 1578 4391 1582 4395
rect 1588 4391 1592 4395
rect 1598 4391 1602 4395
rect 1608 4391 1612 4395
rect 1573 4386 1577 4390
rect 1583 4386 1587 4390
rect 1593 4386 1597 4390
rect 1603 4386 1607 4390
rect 1568 4381 1572 4385
rect 1578 4381 1582 4385
rect 1588 4381 1592 4385
rect 1598 4381 1602 4385
rect 1608 4381 1612 4385
rect 1573 4376 1577 4380
rect 1583 4376 1587 4380
rect 1593 4376 1597 4380
rect 1603 4376 1607 4380
rect 1568 4371 1572 4375
rect 1578 4371 1582 4375
rect 1588 4371 1592 4375
rect 1598 4371 1602 4375
rect 1608 4371 1612 4375
rect 1573 4366 1577 4370
rect 1583 4366 1587 4370
rect 1593 4366 1597 4370
rect 1603 4366 1607 4370
rect 1568 4361 1572 4365
rect 1578 4361 1582 4365
rect 1588 4361 1592 4365
rect 1598 4361 1602 4365
rect 1608 4361 1612 4365
rect 1705 4462 1709 4466
rect 1712 4462 1716 4466
rect 1717 4462 1721 4466
rect 1722 4462 1726 4466
rect 1727 4462 1731 4466
rect 1732 4462 1736 4466
rect 1737 4462 1741 4466
rect 1742 4462 1746 4466
rect 1747 4462 1751 4466
rect 1752 4462 1756 4466
rect 1757 4462 1761 4466
rect 1762 4462 1766 4466
rect 1769 4462 1773 4466
rect 1722 4446 1726 4450
rect 1732 4446 1736 4450
rect 1742 4446 1746 4450
rect 1752 4446 1756 4450
rect 1717 4441 1721 4445
rect 1727 4441 1731 4445
rect 1737 4441 1741 4445
rect 1747 4441 1751 4445
rect 1757 4441 1761 4445
rect 1722 4436 1726 4440
rect 1732 4436 1736 4440
rect 1742 4436 1746 4440
rect 1752 4436 1756 4440
rect 1717 4431 1721 4435
rect 1727 4431 1731 4435
rect 1737 4431 1741 4435
rect 1747 4431 1751 4435
rect 1757 4431 1761 4435
rect 1722 4426 1726 4430
rect 1732 4426 1736 4430
rect 1742 4426 1746 4430
rect 1752 4426 1756 4430
rect 1717 4421 1721 4425
rect 1727 4421 1731 4425
rect 1737 4421 1741 4425
rect 1747 4421 1751 4425
rect 1757 4421 1761 4425
rect 1722 4416 1726 4420
rect 1732 4416 1736 4420
rect 1742 4416 1746 4420
rect 1752 4416 1756 4420
rect 1717 4411 1721 4415
rect 1727 4411 1731 4415
rect 1737 4411 1741 4415
rect 1747 4411 1751 4415
rect 1757 4411 1761 4415
rect 1722 4406 1726 4410
rect 1732 4406 1736 4410
rect 1742 4406 1746 4410
rect 1752 4406 1756 4410
rect 1717 4401 1721 4405
rect 1727 4401 1731 4405
rect 1737 4401 1741 4405
rect 1747 4401 1751 4405
rect 1757 4401 1761 4405
rect 1722 4396 1726 4400
rect 1732 4396 1736 4400
rect 1742 4396 1746 4400
rect 1752 4396 1756 4400
rect 1717 4391 1721 4395
rect 1727 4391 1731 4395
rect 1737 4391 1741 4395
rect 1747 4391 1751 4395
rect 1757 4391 1761 4395
rect 1722 4386 1726 4390
rect 1732 4386 1736 4390
rect 1742 4386 1746 4390
rect 1752 4386 1756 4390
rect 1717 4381 1721 4385
rect 1727 4381 1731 4385
rect 1737 4381 1741 4385
rect 1747 4381 1751 4385
rect 1757 4381 1761 4385
rect 1722 4376 1726 4380
rect 1732 4376 1736 4380
rect 1742 4376 1746 4380
rect 1752 4376 1756 4380
rect 1717 4371 1721 4375
rect 1727 4371 1731 4375
rect 1737 4371 1741 4375
rect 1747 4371 1751 4375
rect 1757 4371 1761 4375
rect 1722 4366 1726 4370
rect 1732 4366 1736 4370
rect 1742 4366 1746 4370
rect 1752 4366 1756 4370
rect 1717 4361 1721 4365
rect 1727 4361 1731 4365
rect 1737 4361 1741 4365
rect 1747 4361 1751 4365
rect 1757 4361 1761 4365
rect 1980 4619 1984 4623
rect 1985 4619 1989 4623
rect 1990 4619 1994 4623
rect 1995 4619 1999 4623
rect 1980 4609 1984 4613
rect 1985 4609 1989 4613
rect 1990 4609 1994 4613
rect 1995 4609 1999 4613
rect 1980 4599 1984 4603
rect 1985 4599 1989 4603
rect 1990 4599 1994 4603
rect 1995 4599 1999 4603
rect 2004 4597 2008 4601
rect 2009 4597 2013 4601
rect 2014 4597 2018 4601
rect 2019 4597 2023 4601
rect 2024 4597 2028 4601
rect 2029 4597 2033 4601
rect 2034 4597 2038 4601
rect 2039 4597 2043 4601
rect 2044 4597 2048 4601
rect 2049 4597 2053 4601
rect 2054 4597 2058 4601
rect 2004 4592 2008 4596
rect 2009 4592 2013 4596
rect 2014 4592 2018 4596
rect 2019 4592 2023 4596
rect 2024 4592 2028 4596
rect 2029 4592 2033 4596
rect 2034 4592 2038 4596
rect 2039 4592 2043 4596
rect 2044 4592 2048 4596
rect 2049 4592 2053 4596
rect 2054 4592 2058 4596
rect 1945 4574 1949 4578
rect 1950 4574 1954 4578
rect 1945 4569 1949 4573
rect 1950 4569 1954 4573
rect 1945 4564 1949 4568
rect 1950 4564 1954 4568
rect 1945 4559 1949 4563
rect 1950 4559 1954 4563
rect 1945 4554 1949 4558
rect 1950 4554 1954 4558
rect 1945 4549 1949 4553
rect 1950 4549 1954 4553
rect 1980 4573 1984 4577
rect 1985 4573 1989 4577
rect 1990 4573 1994 4577
rect 1995 4573 1999 4577
rect 1980 4563 1984 4567
rect 1985 4563 1989 4567
rect 1990 4563 1994 4567
rect 1995 4563 1999 4567
rect 1980 4553 1984 4557
rect 1985 4553 1989 4557
rect 1990 4553 1994 4557
rect 1995 4553 1999 4557
rect 1945 4544 1949 4548
rect 1950 4544 1954 4548
rect 1945 4539 1949 4543
rect 1950 4539 1954 4543
rect 1945 4534 1949 4538
rect 1950 4534 1954 4538
rect 1945 4529 1949 4533
rect 1950 4529 1954 4533
rect 1945 4524 1949 4528
rect 1950 4524 1954 4528
rect 1945 4519 1949 4523
rect 1950 4519 1954 4523
rect 1945 4514 1949 4518
rect 1950 4514 1954 4518
rect 2096 4531 2100 4535
rect 2289 4619 2293 4623
rect 2294 4619 2298 4623
rect 2299 4619 2303 4623
rect 2304 4619 2308 4623
rect 2289 4609 2293 4613
rect 2294 4609 2298 4613
rect 2299 4609 2303 4613
rect 2304 4609 2308 4613
rect 2289 4599 2293 4603
rect 2294 4599 2298 4603
rect 2299 4599 2303 4603
rect 2304 4599 2308 4603
rect 2313 4597 2317 4601
rect 2318 4597 2322 4601
rect 2323 4597 2327 4601
rect 2328 4597 2332 4601
rect 2333 4597 2337 4601
rect 2338 4597 2342 4601
rect 2343 4597 2347 4601
rect 2348 4597 2352 4601
rect 2353 4597 2357 4601
rect 2358 4597 2362 4601
rect 2363 4597 2367 4601
rect 2313 4592 2317 4596
rect 2318 4592 2322 4596
rect 2323 4592 2327 4596
rect 2328 4592 2332 4596
rect 2333 4592 2337 4596
rect 2338 4592 2342 4596
rect 2343 4592 2347 4596
rect 2348 4592 2352 4596
rect 2353 4592 2357 4596
rect 2358 4592 2362 4596
rect 2363 4592 2367 4596
rect 2254 4574 2258 4578
rect 2259 4574 2263 4578
rect 2254 4569 2258 4573
rect 2259 4569 2263 4573
rect 2254 4564 2258 4568
rect 2259 4564 2263 4568
rect 2254 4559 2258 4563
rect 2259 4559 2263 4563
rect 2254 4554 2258 4558
rect 2259 4554 2263 4558
rect 2254 4549 2258 4553
rect 2259 4549 2263 4553
rect 2289 4573 2293 4577
rect 2294 4573 2298 4577
rect 2299 4573 2303 4577
rect 2304 4573 2308 4577
rect 2289 4563 2293 4567
rect 2294 4563 2298 4567
rect 2299 4563 2303 4567
rect 2304 4563 2308 4567
rect 2289 4553 2293 4557
rect 2294 4553 2298 4557
rect 2299 4553 2303 4557
rect 2304 4553 2308 4557
rect 2254 4544 2258 4548
rect 2259 4544 2263 4548
rect 2254 4539 2258 4543
rect 2259 4539 2263 4543
rect 2154 4531 2158 4535
rect 2254 4534 2258 4538
rect 2259 4534 2263 4538
rect 2254 4529 2258 4533
rect 2259 4529 2263 4533
rect 2254 4524 2258 4528
rect 2259 4524 2263 4528
rect 2096 4515 2100 4519
rect 2254 4519 2258 4523
rect 2259 4519 2263 4523
rect 2154 4515 2158 4519
rect 2254 4514 2258 4518
rect 2259 4514 2263 4518
rect 2405 4531 2409 4535
rect 2598 4619 2602 4623
rect 2603 4619 2607 4623
rect 2608 4619 2612 4623
rect 2613 4619 2617 4623
rect 2598 4609 2602 4613
rect 2603 4609 2607 4613
rect 2608 4609 2612 4613
rect 2613 4609 2617 4613
rect 2598 4599 2602 4603
rect 2603 4599 2607 4603
rect 2608 4599 2612 4603
rect 2613 4599 2617 4603
rect 2622 4597 2626 4601
rect 2627 4597 2631 4601
rect 2632 4597 2636 4601
rect 2637 4597 2641 4601
rect 2642 4597 2646 4601
rect 2647 4597 2651 4601
rect 2652 4597 2656 4601
rect 2657 4597 2661 4601
rect 2662 4597 2666 4601
rect 2667 4597 2671 4601
rect 2672 4597 2676 4601
rect 2622 4592 2626 4596
rect 2627 4592 2631 4596
rect 2632 4592 2636 4596
rect 2637 4592 2641 4596
rect 2642 4592 2646 4596
rect 2647 4592 2651 4596
rect 2652 4592 2656 4596
rect 2657 4592 2661 4596
rect 2662 4592 2666 4596
rect 2667 4592 2671 4596
rect 2672 4592 2676 4596
rect 2563 4574 2567 4578
rect 2568 4574 2572 4578
rect 2563 4569 2567 4573
rect 2568 4569 2572 4573
rect 2563 4564 2567 4568
rect 2568 4564 2572 4568
rect 2563 4559 2567 4563
rect 2568 4559 2572 4563
rect 2563 4554 2567 4558
rect 2568 4554 2572 4558
rect 2563 4549 2567 4553
rect 2568 4549 2572 4553
rect 2598 4573 2602 4577
rect 2603 4573 2607 4577
rect 2608 4573 2612 4577
rect 2613 4573 2617 4577
rect 2598 4563 2602 4567
rect 2603 4563 2607 4567
rect 2608 4563 2612 4567
rect 2613 4563 2617 4567
rect 2598 4553 2602 4557
rect 2603 4553 2607 4557
rect 2608 4553 2612 4557
rect 2613 4553 2617 4557
rect 2563 4544 2567 4548
rect 2568 4544 2572 4548
rect 2563 4539 2567 4543
rect 2568 4539 2572 4543
rect 2463 4531 2467 4535
rect 2563 4534 2567 4538
rect 2568 4534 2572 4538
rect 2563 4529 2567 4533
rect 2568 4529 2572 4533
rect 2563 4524 2567 4528
rect 2568 4524 2572 4528
rect 2405 4515 2409 4519
rect 2096 4499 2100 4503
rect 2154 4499 2158 4503
rect 2096 4483 2100 4487
rect 2154 4483 2158 4487
rect 1865 4462 1869 4466
rect 1872 4462 1876 4466
rect 1877 4462 1881 4466
rect 1882 4462 1886 4466
rect 1887 4462 1891 4466
rect 1892 4462 1896 4466
rect 1897 4462 1901 4466
rect 1902 4462 1906 4466
rect 1907 4462 1911 4466
rect 1912 4462 1916 4466
rect 1917 4462 1921 4466
rect 1922 4462 1926 4466
rect 1929 4462 1933 4466
rect 1882 4446 1886 4450
rect 1892 4446 1896 4450
rect 1902 4446 1906 4450
rect 1912 4446 1916 4450
rect 1877 4441 1881 4445
rect 1887 4441 1891 4445
rect 1897 4441 1901 4445
rect 1907 4441 1911 4445
rect 1917 4441 1921 4445
rect 1882 4436 1886 4440
rect 1892 4436 1896 4440
rect 1902 4436 1906 4440
rect 1912 4436 1916 4440
rect 1877 4431 1881 4435
rect 1887 4431 1891 4435
rect 1897 4431 1901 4435
rect 1907 4431 1911 4435
rect 1917 4431 1921 4435
rect 1882 4426 1886 4430
rect 1892 4426 1896 4430
rect 1902 4426 1906 4430
rect 1912 4426 1916 4430
rect 1877 4421 1881 4425
rect 1887 4421 1891 4425
rect 1897 4421 1901 4425
rect 1907 4421 1911 4425
rect 1917 4421 1921 4425
rect 1882 4416 1886 4420
rect 1892 4416 1896 4420
rect 1902 4416 1906 4420
rect 1912 4416 1916 4420
rect 1877 4411 1881 4415
rect 1887 4411 1891 4415
rect 1897 4411 1901 4415
rect 1907 4411 1911 4415
rect 1917 4411 1921 4415
rect 1882 4406 1886 4410
rect 1892 4406 1896 4410
rect 1902 4406 1906 4410
rect 1912 4406 1916 4410
rect 1877 4401 1881 4405
rect 1887 4401 1891 4405
rect 1897 4401 1901 4405
rect 1907 4401 1911 4405
rect 1917 4401 1921 4405
rect 1882 4396 1886 4400
rect 1892 4396 1896 4400
rect 1902 4396 1906 4400
rect 1912 4396 1916 4400
rect 1877 4391 1881 4395
rect 1887 4391 1891 4395
rect 1897 4391 1901 4395
rect 1907 4391 1911 4395
rect 1917 4391 1921 4395
rect 1882 4386 1886 4390
rect 1892 4386 1896 4390
rect 1902 4386 1906 4390
rect 1912 4386 1916 4390
rect 1877 4381 1881 4385
rect 1887 4381 1891 4385
rect 1897 4381 1901 4385
rect 1907 4381 1911 4385
rect 1917 4381 1921 4385
rect 1882 4376 1886 4380
rect 1892 4376 1896 4380
rect 1902 4376 1906 4380
rect 1912 4376 1916 4380
rect 1877 4371 1881 4375
rect 1887 4371 1891 4375
rect 1897 4371 1901 4375
rect 1907 4371 1911 4375
rect 1917 4371 1921 4375
rect 1882 4366 1886 4370
rect 1892 4366 1896 4370
rect 1902 4366 1906 4370
rect 1912 4366 1916 4370
rect 1877 4361 1881 4365
rect 1887 4361 1891 4365
rect 1897 4361 1901 4365
rect 1907 4361 1911 4365
rect 1917 4361 1921 4365
rect 2563 4519 2567 4523
rect 2568 4519 2572 4523
rect 2463 4515 2467 4519
rect 2563 4514 2567 4518
rect 2568 4514 2572 4518
rect 2714 4531 2718 4535
rect 2907 4619 2911 4623
rect 2912 4619 2916 4623
rect 2917 4619 2921 4623
rect 2922 4619 2926 4623
rect 2907 4609 2911 4613
rect 2912 4609 2916 4613
rect 2917 4609 2921 4613
rect 2922 4609 2926 4613
rect 2907 4599 2911 4603
rect 2912 4599 2916 4603
rect 2917 4599 2921 4603
rect 2922 4599 2926 4603
rect 2931 4597 2935 4601
rect 2936 4597 2940 4601
rect 2941 4597 2945 4601
rect 2946 4597 2950 4601
rect 2951 4597 2955 4601
rect 2956 4597 2960 4601
rect 2961 4597 2965 4601
rect 2966 4597 2970 4601
rect 2971 4597 2975 4601
rect 2976 4597 2980 4601
rect 2981 4597 2985 4601
rect 2931 4592 2935 4596
rect 2936 4592 2940 4596
rect 2941 4592 2945 4596
rect 2946 4592 2950 4596
rect 2951 4592 2955 4596
rect 2956 4592 2960 4596
rect 2961 4592 2965 4596
rect 2966 4592 2970 4596
rect 2971 4592 2975 4596
rect 2976 4592 2980 4596
rect 2981 4592 2985 4596
rect 2872 4574 2876 4578
rect 2877 4574 2881 4578
rect 2872 4569 2876 4573
rect 2877 4569 2881 4573
rect 2872 4564 2876 4568
rect 2877 4564 2881 4568
rect 2872 4559 2876 4563
rect 2877 4559 2881 4563
rect 2872 4554 2876 4558
rect 2877 4554 2881 4558
rect 2872 4549 2876 4553
rect 2877 4549 2881 4553
rect 2907 4573 2911 4577
rect 2912 4573 2916 4577
rect 2917 4573 2921 4577
rect 2922 4573 2926 4577
rect 2907 4563 2911 4567
rect 2912 4563 2916 4567
rect 2917 4563 2921 4567
rect 2922 4563 2926 4567
rect 2907 4553 2911 4557
rect 2912 4553 2916 4557
rect 2917 4553 2921 4557
rect 2922 4553 2926 4557
rect 2872 4544 2876 4548
rect 2877 4544 2881 4548
rect 2872 4539 2876 4543
rect 2877 4539 2881 4543
rect 2772 4531 2776 4535
rect 2872 4534 2876 4538
rect 2877 4534 2881 4538
rect 2872 4529 2876 4533
rect 2877 4529 2881 4533
rect 2872 4524 2876 4528
rect 2877 4524 2881 4528
rect 2714 4515 2718 4519
rect 2405 4499 2409 4503
rect 2463 4499 2467 4503
rect 2405 4483 2409 4487
rect 2463 4483 2467 4487
rect 2014 4462 2018 4466
rect 2021 4462 2025 4466
rect 2026 4462 2030 4466
rect 2031 4462 2035 4466
rect 2036 4462 2040 4466
rect 2041 4462 2045 4466
rect 2046 4462 2050 4466
rect 2051 4462 2055 4466
rect 2056 4462 2060 4466
rect 2061 4462 2065 4466
rect 2066 4462 2070 4466
rect 2071 4462 2075 4466
rect 2078 4462 2082 4466
rect 2031 4446 2035 4450
rect 2041 4446 2045 4450
rect 2051 4446 2055 4450
rect 2061 4446 2065 4450
rect 2026 4441 2030 4445
rect 2036 4441 2040 4445
rect 2046 4441 2050 4445
rect 2056 4441 2060 4445
rect 2066 4441 2070 4445
rect 2031 4436 2035 4440
rect 2041 4436 2045 4440
rect 2051 4436 2055 4440
rect 2061 4436 2065 4440
rect 2026 4431 2030 4435
rect 2036 4431 2040 4435
rect 2046 4431 2050 4435
rect 2056 4431 2060 4435
rect 2066 4431 2070 4435
rect 2031 4426 2035 4430
rect 2041 4426 2045 4430
rect 2051 4426 2055 4430
rect 2061 4426 2065 4430
rect 2026 4421 2030 4425
rect 2036 4421 2040 4425
rect 2046 4421 2050 4425
rect 2056 4421 2060 4425
rect 2066 4421 2070 4425
rect 2031 4416 2035 4420
rect 2041 4416 2045 4420
rect 2051 4416 2055 4420
rect 2061 4416 2065 4420
rect 2026 4411 2030 4415
rect 2036 4411 2040 4415
rect 2046 4411 2050 4415
rect 2056 4411 2060 4415
rect 2066 4411 2070 4415
rect 2031 4406 2035 4410
rect 2041 4406 2045 4410
rect 2051 4406 2055 4410
rect 2061 4406 2065 4410
rect 2026 4401 2030 4405
rect 2036 4401 2040 4405
rect 2046 4401 2050 4405
rect 2056 4401 2060 4405
rect 2066 4401 2070 4405
rect 2031 4396 2035 4400
rect 2041 4396 2045 4400
rect 2051 4396 2055 4400
rect 2061 4396 2065 4400
rect 2026 4391 2030 4395
rect 2036 4391 2040 4395
rect 2046 4391 2050 4395
rect 2056 4391 2060 4395
rect 2066 4391 2070 4395
rect 2031 4386 2035 4390
rect 2041 4386 2045 4390
rect 2051 4386 2055 4390
rect 2061 4386 2065 4390
rect 2026 4381 2030 4385
rect 2036 4381 2040 4385
rect 2046 4381 2050 4385
rect 2056 4381 2060 4385
rect 2066 4381 2070 4385
rect 2031 4376 2035 4380
rect 2041 4376 2045 4380
rect 2051 4376 2055 4380
rect 2061 4376 2065 4380
rect 2026 4371 2030 4375
rect 2036 4371 2040 4375
rect 2046 4371 2050 4375
rect 2056 4371 2060 4375
rect 2066 4371 2070 4375
rect 2031 4366 2035 4370
rect 2041 4366 2045 4370
rect 2051 4366 2055 4370
rect 2061 4366 2065 4370
rect 2026 4361 2030 4365
rect 2036 4361 2040 4365
rect 2046 4361 2050 4365
rect 2056 4361 2060 4365
rect 2066 4361 2070 4365
rect 2174 4462 2178 4466
rect 2181 4462 2185 4466
rect 2186 4462 2190 4466
rect 2191 4462 2195 4466
rect 2196 4462 2200 4466
rect 2201 4462 2205 4466
rect 2206 4462 2210 4466
rect 2211 4462 2215 4466
rect 2216 4462 2220 4466
rect 2221 4462 2225 4466
rect 2226 4462 2230 4466
rect 2231 4462 2235 4466
rect 2238 4462 2242 4466
rect 2191 4446 2195 4450
rect 2201 4446 2205 4450
rect 2211 4446 2215 4450
rect 2221 4446 2225 4450
rect 2186 4441 2190 4445
rect 2196 4441 2200 4445
rect 2206 4441 2210 4445
rect 2216 4441 2220 4445
rect 2226 4441 2230 4445
rect 2191 4436 2195 4440
rect 2201 4436 2205 4440
rect 2211 4436 2215 4440
rect 2221 4436 2225 4440
rect 2186 4431 2190 4435
rect 2196 4431 2200 4435
rect 2206 4431 2210 4435
rect 2216 4431 2220 4435
rect 2226 4431 2230 4435
rect 2191 4426 2195 4430
rect 2201 4426 2205 4430
rect 2211 4426 2215 4430
rect 2221 4426 2225 4430
rect 2186 4421 2190 4425
rect 2196 4421 2200 4425
rect 2206 4421 2210 4425
rect 2216 4421 2220 4425
rect 2226 4421 2230 4425
rect 2191 4416 2195 4420
rect 2201 4416 2205 4420
rect 2211 4416 2215 4420
rect 2221 4416 2225 4420
rect 2186 4411 2190 4415
rect 2196 4411 2200 4415
rect 2206 4411 2210 4415
rect 2216 4411 2220 4415
rect 2226 4411 2230 4415
rect 2191 4406 2195 4410
rect 2201 4406 2205 4410
rect 2211 4406 2215 4410
rect 2221 4406 2225 4410
rect 2186 4401 2190 4405
rect 2196 4401 2200 4405
rect 2206 4401 2210 4405
rect 2216 4401 2220 4405
rect 2226 4401 2230 4405
rect 2191 4396 2195 4400
rect 2201 4396 2205 4400
rect 2211 4396 2215 4400
rect 2221 4396 2225 4400
rect 2186 4391 2190 4395
rect 2196 4391 2200 4395
rect 2206 4391 2210 4395
rect 2216 4391 2220 4395
rect 2226 4391 2230 4395
rect 2191 4386 2195 4390
rect 2201 4386 2205 4390
rect 2211 4386 2215 4390
rect 2221 4386 2225 4390
rect 2186 4381 2190 4385
rect 2196 4381 2200 4385
rect 2206 4381 2210 4385
rect 2216 4381 2220 4385
rect 2226 4381 2230 4385
rect 2191 4376 2195 4380
rect 2201 4376 2205 4380
rect 2211 4376 2215 4380
rect 2221 4376 2225 4380
rect 2186 4371 2190 4375
rect 2196 4371 2200 4375
rect 2206 4371 2210 4375
rect 2216 4371 2220 4375
rect 2226 4371 2230 4375
rect 2191 4366 2195 4370
rect 2201 4366 2205 4370
rect 2211 4366 2215 4370
rect 2221 4366 2225 4370
rect 2186 4361 2190 4365
rect 2196 4361 2200 4365
rect 2206 4361 2210 4365
rect 2216 4361 2220 4365
rect 2226 4361 2230 4365
rect 2872 4519 2876 4523
rect 2877 4519 2881 4523
rect 2772 4515 2776 4519
rect 2872 4514 2876 4518
rect 2877 4514 2881 4518
rect 3023 4531 3027 4535
rect 3216 4619 3220 4623
rect 3221 4619 3225 4623
rect 3226 4619 3230 4623
rect 3231 4619 3235 4623
rect 3216 4609 3220 4613
rect 3221 4609 3225 4613
rect 3226 4609 3230 4613
rect 3231 4609 3235 4613
rect 3216 4599 3220 4603
rect 3221 4599 3225 4603
rect 3226 4599 3230 4603
rect 3231 4599 3235 4603
rect 3240 4597 3244 4601
rect 3245 4597 3249 4601
rect 3250 4597 3254 4601
rect 3255 4597 3259 4601
rect 3260 4597 3264 4601
rect 3265 4597 3269 4601
rect 3270 4597 3274 4601
rect 3275 4597 3279 4601
rect 3280 4597 3284 4601
rect 3285 4597 3289 4601
rect 3290 4597 3294 4601
rect 3240 4592 3244 4596
rect 3245 4592 3249 4596
rect 3250 4592 3254 4596
rect 3255 4592 3259 4596
rect 3260 4592 3264 4596
rect 3265 4592 3269 4596
rect 3270 4592 3274 4596
rect 3275 4592 3279 4596
rect 3280 4592 3284 4596
rect 3285 4592 3289 4596
rect 3290 4592 3294 4596
rect 3181 4574 3185 4578
rect 3186 4574 3190 4578
rect 3181 4569 3185 4573
rect 3186 4569 3190 4573
rect 3181 4564 3185 4568
rect 3186 4564 3190 4568
rect 3181 4559 3185 4563
rect 3186 4559 3190 4563
rect 3181 4554 3185 4558
rect 3186 4554 3190 4558
rect 3181 4549 3185 4553
rect 3186 4549 3190 4553
rect 3216 4573 3220 4577
rect 3221 4573 3225 4577
rect 3226 4573 3230 4577
rect 3231 4573 3235 4577
rect 3216 4563 3220 4567
rect 3221 4563 3225 4567
rect 3226 4563 3230 4567
rect 3231 4563 3235 4567
rect 3216 4553 3220 4557
rect 3221 4553 3225 4557
rect 3226 4553 3230 4557
rect 3231 4553 3235 4557
rect 3181 4544 3185 4548
rect 3186 4544 3190 4548
rect 3181 4539 3185 4543
rect 3186 4539 3190 4543
rect 3081 4531 3085 4535
rect 3181 4534 3185 4538
rect 3186 4534 3190 4538
rect 3181 4529 3185 4533
rect 3186 4529 3190 4533
rect 3181 4524 3185 4528
rect 3186 4524 3190 4528
rect 3023 4515 3027 4519
rect 2714 4499 2718 4503
rect 2772 4499 2776 4503
rect 2714 4483 2718 4487
rect 2772 4483 2776 4487
rect 2323 4462 2327 4466
rect 2330 4462 2334 4466
rect 2335 4462 2339 4466
rect 2340 4462 2344 4466
rect 2345 4462 2349 4466
rect 2350 4462 2354 4466
rect 2355 4462 2359 4466
rect 2360 4462 2364 4466
rect 2365 4462 2369 4466
rect 2370 4462 2374 4466
rect 2375 4462 2379 4466
rect 2380 4462 2384 4466
rect 2387 4462 2391 4466
rect 2340 4446 2344 4450
rect 2350 4446 2354 4450
rect 2360 4446 2364 4450
rect 2370 4446 2374 4450
rect 2335 4441 2339 4445
rect 2345 4441 2349 4445
rect 2355 4441 2359 4445
rect 2365 4441 2369 4445
rect 2375 4441 2379 4445
rect 2340 4436 2344 4440
rect 2350 4436 2354 4440
rect 2360 4436 2364 4440
rect 2370 4436 2374 4440
rect 2335 4431 2339 4435
rect 2345 4431 2349 4435
rect 2355 4431 2359 4435
rect 2365 4431 2369 4435
rect 2375 4431 2379 4435
rect 2340 4426 2344 4430
rect 2350 4426 2354 4430
rect 2360 4426 2364 4430
rect 2370 4426 2374 4430
rect 2335 4421 2339 4425
rect 2345 4421 2349 4425
rect 2355 4421 2359 4425
rect 2365 4421 2369 4425
rect 2375 4421 2379 4425
rect 2340 4416 2344 4420
rect 2350 4416 2354 4420
rect 2360 4416 2364 4420
rect 2370 4416 2374 4420
rect 2335 4411 2339 4415
rect 2345 4411 2349 4415
rect 2355 4411 2359 4415
rect 2365 4411 2369 4415
rect 2375 4411 2379 4415
rect 2340 4406 2344 4410
rect 2350 4406 2354 4410
rect 2360 4406 2364 4410
rect 2370 4406 2374 4410
rect 2335 4401 2339 4405
rect 2345 4401 2349 4405
rect 2355 4401 2359 4405
rect 2365 4401 2369 4405
rect 2375 4401 2379 4405
rect 2340 4396 2344 4400
rect 2350 4396 2354 4400
rect 2360 4396 2364 4400
rect 2370 4396 2374 4400
rect 2335 4391 2339 4395
rect 2345 4391 2349 4395
rect 2355 4391 2359 4395
rect 2365 4391 2369 4395
rect 2375 4391 2379 4395
rect 2340 4386 2344 4390
rect 2350 4386 2354 4390
rect 2360 4386 2364 4390
rect 2370 4386 2374 4390
rect 2335 4381 2339 4385
rect 2345 4381 2349 4385
rect 2355 4381 2359 4385
rect 2365 4381 2369 4385
rect 2375 4381 2379 4385
rect 2340 4376 2344 4380
rect 2350 4376 2354 4380
rect 2360 4376 2364 4380
rect 2370 4376 2374 4380
rect 2335 4371 2339 4375
rect 2345 4371 2349 4375
rect 2355 4371 2359 4375
rect 2365 4371 2369 4375
rect 2375 4371 2379 4375
rect 2340 4366 2344 4370
rect 2350 4366 2354 4370
rect 2360 4366 2364 4370
rect 2370 4366 2374 4370
rect 2335 4361 2339 4365
rect 2345 4361 2349 4365
rect 2355 4361 2359 4365
rect 2365 4361 2369 4365
rect 2375 4361 2379 4365
rect 2483 4462 2487 4466
rect 2490 4462 2494 4466
rect 2495 4462 2499 4466
rect 2500 4462 2504 4466
rect 2505 4462 2509 4466
rect 2510 4462 2514 4466
rect 2515 4462 2519 4466
rect 2520 4462 2524 4466
rect 2525 4462 2529 4466
rect 2530 4462 2534 4466
rect 2535 4462 2539 4466
rect 2540 4462 2544 4466
rect 2547 4462 2551 4466
rect 2500 4446 2504 4450
rect 2510 4446 2514 4450
rect 2520 4446 2524 4450
rect 2530 4446 2534 4450
rect 2495 4441 2499 4445
rect 2505 4441 2509 4445
rect 2515 4441 2519 4445
rect 2525 4441 2529 4445
rect 2535 4441 2539 4445
rect 2500 4436 2504 4440
rect 2510 4436 2514 4440
rect 2520 4436 2524 4440
rect 2530 4436 2534 4440
rect 2495 4431 2499 4435
rect 2505 4431 2509 4435
rect 2515 4431 2519 4435
rect 2525 4431 2529 4435
rect 2535 4431 2539 4435
rect 2500 4426 2504 4430
rect 2510 4426 2514 4430
rect 2520 4426 2524 4430
rect 2530 4426 2534 4430
rect 2495 4421 2499 4425
rect 2505 4421 2509 4425
rect 2515 4421 2519 4425
rect 2525 4421 2529 4425
rect 2535 4421 2539 4425
rect 2500 4416 2504 4420
rect 2510 4416 2514 4420
rect 2520 4416 2524 4420
rect 2530 4416 2534 4420
rect 2495 4411 2499 4415
rect 2505 4411 2509 4415
rect 2515 4411 2519 4415
rect 2525 4411 2529 4415
rect 2535 4411 2539 4415
rect 2500 4406 2504 4410
rect 2510 4406 2514 4410
rect 2520 4406 2524 4410
rect 2530 4406 2534 4410
rect 2495 4401 2499 4405
rect 2505 4401 2509 4405
rect 2515 4401 2519 4405
rect 2525 4401 2529 4405
rect 2535 4401 2539 4405
rect 2500 4396 2504 4400
rect 2510 4396 2514 4400
rect 2520 4396 2524 4400
rect 2530 4396 2534 4400
rect 2495 4391 2499 4395
rect 2505 4391 2509 4395
rect 2515 4391 2519 4395
rect 2525 4391 2529 4395
rect 2535 4391 2539 4395
rect 2500 4386 2504 4390
rect 2510 4386 2514 4390
rect 2520 4386 2524 4390
rect 2530 4386 2534 4390
rect 2495 4381 2499 4385
rect 2505 4381 2509 4385
rect 2515 4381 2519 4385
rect 2525 4381 2529 4385
rect 2535 4381 2539 4385
rect 2500 4376 2504 4380
rect 2510 4376 2514 4380
rect 2520 4376 2524 4380
rect 2530 4376 2534 4380
rect 2495 4371 2499 4375
rect 2505 4371 2509 4375
rect 2515 4371 2519 4375
rect 2525 4371 2529 4375
rect 2535 4371 2539 4375
rect 2500 4366 2504 4370
rect 2510 4366 2514 4370
rect 2520 4366 2524 4370
rect 2530 4366 2534 4370
rect 2495 4361 2499 4365
rect 2505 4361 2509 4365
rect 2515 4361 2519 4365
rect 2525 4361 2529 4365
rect 2535 4361 2539 4365
rect 3181 4519 3185 4523
rect 3186 4519 3190 4523
rect 3081 4515 3085 4519
rect 3181 4514 3185 4518
rect 3186 4514 3190 4518
rect 3332 4531 3336 4535
rect 4484 4718 4488 4722
rect 4494 4718 4498 4722
rect 4504 4718 4508 4722
rect 4530 4733 4534 4737
rect 4540 4733 4544 4737
rect 4550 4733 4554 4737
rect 4530 4728 4534 4732
rect 4540 4728 4544 4732
rect 4550 4728 4554 4732
rect 4530 4723 4534 4727
rect 4540 4723 4544 4727
rect 4550 4723 4554 4727
rect 4530 4718 4534 4722
rect 4540 4718 4544 4722
rect 4550 4718 4554 4722
rect 4484 4707 4488 4711
rect 4494 4707 4498 4711
rect 4504 4707 4508 4711
rect 3664 4649 3668 4653
rect 3669 4649 3673 4653
rect 3664 4644 3668 4648
rect 3669 4644 3673 4648
rect 3664 4639 3668 4643
rect 3669 4639 3673 4643
rect 3664 4634 3668 4638
rect 3669 4634 3673 4638
rect 3664 4629 3668 4633
rect 3669 4629 3673 4633
rect 3525 4619 3529 4623
rect 3530 4619 3534 4623
rect 3535 4619 3539 4623
rect 3540 4619 3544 4623
rect 3525 4609 3529 4613
rect 3530 4609 3534 4613
rect 3535 4609 3539 4613
rect 3540 4609 3544 4613
rect 3525 4599 3529 4603
rect 3530 4599 3534 4603
rect 3535 4599 3539 4603
rect 3540 4599 3544 4603
rect 3664 4624 3668 4628
rect 3669 4624 3673 4628
rect 3664 4619 3668 4623
rect 3669 4619 3673 4623
rect 3664 4614 3668 4618
rect 3669 4614 3673 4618
rect 3664 4609 3668 4613
rect 3669 4609 3673 4613
rect 3664 4604 3668 4608
rect 3669 4604 3673 4608
rect 3549 4597 3553 4601
rect 3554 4597 3558 4601
rect 3559 4597 3563 4601
rect 3564 4597 3568 4601
rect 3569 4597 3573 4601
rect 3574 4597 3578 4601
rect 3579 4597 3583 4601
rect 3584 4597 3588 4601
rect 3589 4597 3593 4601
rect 3594 4597 3598 4601
rect 3599 4597 3603 4601
rect 3549 4592 3553 4596
rect 3554 4592 3558 4596
rect 3559 4592 3563 4596
rect 3564 4592 3568 4596
rect 3569 4592 3573 4596
rect 3574 4592 3578 4596
rect 3579 4592 3583 4596
rect 3584 4592 3588 4596
rect 3589 4592 3593 4596
rect 3594 4592 3598 4596
rect 3599 4592 3603 4596
rect 3490 4574 3494 4578
rect 3495 4574 3499 4578
rect 3490 4569 3494 4573
rect 3495 4569 3499 4573
rect 3490 4564 3494 4568
rect 3495 4564 3499 4568
rect 3490 4559 3494 4563
rect 3495 4559 3499 4563
rect 3490 4554 3494 4558
rect 3495 4554 3499 4558
rect 3490 4549 3494 4553
rect 3495 4549 3499 4553
rect 3525 4573 3529 4577
rect 3530 4573 3534 4577
rect 3535 4573 3539 4577
rect 3540 4573 3544 4577
rect 3525 4563 3529 4567
rect 3530 4563 3534 4567
rect 3535 4563 3539 4567
rect 3540 4563 3544 4567
rect 3525 4553 3529 4557
rect 3530 4553 3534 4557
rect 3535 4553 3539 4557
rect 3540 4553 3544 4557
rect 3490 4544 3494 4548
rect 3495 4544 3499 4548
rect 3490 4539 3494 4543
rect 3495 4539 3499 4543
rect 3390 4531 3394 4535
rect 3490 4534 3494 4538
rect 3495 4534 3499 4538
rect 3490 4529 3494 4533
rect 3495 4529 3499 4533
rect 3490 4524 3494 4528
rect 3495 4524 3499 4528
rect 3332 4515 3336 4519
rect 3023 4499 3027 4503
rect 3081 4499 3085 4503
rect 3023 4483 3027 4487
rect 3081 4483 3085 4487
rect 2632 4462 2636 4466
rect 2639 4462 2643 4466
rect 2644 4462 2648 4466
rect 2649 4462 2653 4466
rect 2654 4462 2658 4466
rect 2659 4462 2663 4466
rect 2664 4462 2668 4466
rect 2669 4462 2673 4466
rect 2674 4462 2678 4466
rect 2679 4462 2683 4466
rect 2684 4462 2688 4466
rect 2689 4462 2693 4466
rect 2696 4462 2700 4466
rect 2649 4446 2653 4450
rect 2659 4446 2663 4450
rect 2669 4446 2673 4450
rect 2679 4446 2683 4450
rect 2644 4441 2648 4445
rect 2654 4441 2658 4445
rect 2664 4441 2668 4445
rect 2674 4441 2678 4445
rect 2684 4441 2688 4445
rect 2649 4436 2653 4440
rect 2659 4436 2663 4440
rect 2669 4436 2673 4440
rect 2679 4436 2683 4440
rect 2644 4431 2648 4435
rect 2654 4431 2658 4435
rect 2664 4431 2668 4435
rect 2674 4431 2678 4435
rect 2684 4431 2688 4435
rect 2649 4426 2653 4430
rect 2659 4426 2663 4430
rect 2669 4426 2673 4430
rect 2679 4426 2683 4430
rect 2644 4421 2648 4425
rect 2654 4421 2658 4425
rect 2664 4421 2668 4425
rect 2674 4421 2678 4425
rect 2684 4421 2688 4425
rect 2649 4416 2653 4420
rect 2659 4416 2663 4420
rect 2669 4416 2673 4420
rect 2679 4416 2683 4420
rect 2644 4411 2648 4415
rect 2654 4411 2658 4415
rect 2664 4411 2668 4415
rect 2674 4411 2678 4415
rect 2684 4411 2688 4415
rect 2649 4406 2653 4410
rect 2659 4406 2663 4410
rect 2669 4406 2673 4410
rect 2679 4406 2683 4410
rect 2644 4401 2648 4405
rect 2654 4401 2658 4405
rect 2664 4401 2668 4405
rect 2674 4401 2678 4405
rect 2684 4401 2688 4405
rect 2649 4396 2653 4400
rect 2659 4396 2663 4400
rect 2669 4396 2673 4400
rect 2679 4396 2683 4400
rect 2644 4391 2648 4395
rect 2654 4391 2658 4395
rect 2664 4391 2668 4395
rect 2674 4391 2678 4395
rect 2684 4391 2688 4395
rect 2649 4386 2653 4390
rect 2659 4386 2663 4390
rect 2669 4386 2673 4390
rect 2679 4386 2683 4390
rect 2644 4381 2648 4385
rect 2654 4381 2658 4385
rect 2664 4381 2668 4385
rect 2674 4381 2678 4385
rect 2684 4381 2688 4385
rect 2649 4376 2653 4380
rect 2659 4376 2663 4380
rect 2669 4376 2673 4380
rect 2679 4376 2683 4380
rect 2644 4371 2648 4375
rect 2654 4371 2658 4375
rect 2664 4371 2668 4375
rect 2674 4371 2678 4375
rect 2684 4371 2688 4375
rect 2649 4366 2653 4370
rect 2659 4366 2663 4370
rect 2669 4366 2673 4370
rect 2679 4366 2683 4370
rect 2644 4361 2648 4365
rect 2654 4361 2658 4365
rect 2664 4361 2668 4365
rect 2674 4361 2678 4365
rect 2684 4361 2688 4365
rect 2792 4462 2796 4466
rect 2799 4462 2803 4466
rect 2804 4462 2808 4466
rect 2809 4462 2813 4466
rect 2814 4462 2818 4466
rect 2819 4462 2823 4466
rect 2824 4462 2828 4466
rect 2829 4462 2833 4466
rect 2834 4462 2838 4466
rect 2839 4462 2843 4466
rect 2844 4462 2848 4466
rect 2849 4462 2853 4466
rect 2856 4462 2860 4466
rect 2809 4446 2813 4450
rect 2819 4446 2823 4450
rect 2829 4446 2833 4450
rect 2839 4446 2843 4450
rect 2804 4441 2808 4445
rect 2814 4441 2818 4445
rect 2824 4441 2828 4445
rect 2834 4441 2838 4445
rect 2844 4441 2848 4445
rect 2809 4436 2813 4440
rect 2819 4436 2823 4440
rect 2829 4436 2833 4440
rect 2839 4436 2843 4440
rect 2804 4431 2808 4435
rect 2814 4431 2818 4435
rect 2824 4431 2828 4435
rect 2834 4431 2838 4435
rect 2844 4431 2848 4435
rect 2809 4426 2813 4430
rect 2819 4426 2823 4430
rect 2829 4426 2833 4430
rect 2839 4426 2843 4430
rect 2804 4421 2808 4425
rect 2814 4421 2818 4425
rect 2824 4421 2828 4425
rect 2834 4421 2838 4425
rect 2844 4421 2848 4425
rect 2809 4416 2813 4420
rect 2819 4416 2823 4420
rect 2829 4416 2833 4420
rect 2839 4416 2843 4420
rect 2804 4411 2808 4415
rect 2814 4411 2818 4415
rect 2824 4411 2828 4415
rect 2834 4411 2838 4415
rect 2844 4411 2848 4415
rect 2809 4406 2813 4410
rect 2819 4406 2823 4410
rect 2829 4406 2833 4410
rect 2839 4406 2843 4410
rect 2804 4401 2808 4405
rect 2814 4401 2818 4405
rect 2824 4401 2828 4405
rect 2834 4401 2838 4405
rect 2844 4401 2848 4405
rect 2809 4396 2813 4400
rect 2819 4396 2823 4400
rect 2829 4396 2833 4400
rect 2839 4396 2843 4400
rect 2804 4391 2808 4395
rect 2814 4391 2818 4395
rect 2824 4391 2828 4395
rect 2834 4391 2838 4395
rect 2844 4391 2848 4395
rect 2809 4386 2813 4390
rect 2819 4386 2823 4390
rect 2829 4386 2833 4390
rect 2839 4386 2843 4390
rect 2804 4381 2808 4385
rect 2814 4381 2818 4385
rect 2824 4381 2828 4385
rect 2834 4381 2838 4385
rect 2844 4381 2848 4385
rect 2809 4376 2813 4380
rect 2819 4376 2823 4380
rect 2829 4376 2833 4380
rect 2839 4376 2843 4380
rect 2804 4371 2808 4375
rect 2814 4371 2818 4375
rect 2824 4371 2828 4375
rect 2834 4371 2838 4375
rect 2844 4371 2848 4375
rect 2809 4366 2813 4370
rect 2819 4366 2823 4370
rect 2829 4366 2833 4370
rect 2839 4366 2843 4370
rect 2804 4361 2808 4365
rect 2814 4361 2818 4365
rect 2824 4361 2828 4365
rect 2834 4361 2838 4365
rect 2844 4361 2848 4365
rect 3490 4519 3494 4523
rect 3495 4519 3499 4523
rect 3390 4515 3394 4519
rect 3490 4514 3494 4518
rect 3495 4514 3499 4518
rect 3332 4499 3336 4503
rect 3390 4499 3394 4503
rect 3332 4483 3336 4487
rect 3390 4483 3394 4487
rect 2941 4462 2945 4466
rect 2948 4462 2952 4466
rect 2953 4462 2957 4466
rect 2958 4462 2962 4466
rect 2963 4462 2967 4466
rect 2968 4462 2972 4466
rect 2973 4462 2977 4466
rect 2978 4462 2982 4466
rect 2983 4462 2987 4466
rect 2988 4462 2992 4466
rect 2993 4462 2997 4466
rect 2998 4462 3002 4466
rect 3005 4462 3009 4466
rect 2958 4446 2962 4450
rect 2968 4446 2972 4450
rect 2978 4446 2982 4450
rect 2988 4446 2992 4450
rect 2953 4441 2957 4445
rect 2963 4441 2967 4445
rect 2973 4441 2977 4445
rect 2983 4441 2987 4445
rect 2993 4441 2997 4445
rect 2958 4436 2962 4440
rect 2968 4436 2972 4440
rect 2978 4436 2982 4440
rect 2988 4436 2992 4440
rect 2953 4431 2957 4435
rect 2963 4431 2967 4435
rect 2973 4431 2977 4435
rect 2983 4431 2987 4435
rect 2993 4431 2997 4435
rect 2958 4426 2962 4430
rect 2968 4426 2972 4430
rect 2978 4426 2982 4430
rect 2988 4426 2992 4430
rect 2953 4421 2957 4425
rect 2963 4421 2967 4425
rect 2973 4421 2977 4425
rect 2983 4421 2987 4425
rect 2993 4421 2997 4425
rect 2958 4416 2962 4420
rect 2968 4416 2972 4420
rect 2978 4416 2982 4420
rect 2988 4416 2992 4420
rect 2953 4411 2957 4415
rect 2963 4411 2967 4415
rect 2973 4411 2977 4415
rect 2983 4411 2987 4415
rect 2993 4411 2997 4415
rect 2958 4406 2962 4410
rect 2968 4406 2972 4410
rect 2978 4406 2982 4410
rect 2988 4406 2992 4410
rect 2953 4401 2957 4405
rect 2963 4401 2967 4405
rect 2973 4401 2977 4405
rect 2983 4401 2987 4405
rect 2993 4401 2997 4405
rect 2958 4396 2962 4400
rect 2968 4396 2972 4400
rect 2978 4396 2982 4400
rect 2988 4396 2992 4400
rect 2953 4391 2957 4395
rect 2963 4391 2967 4395
rect 2973 4391 2977 4395
rect 2983 4391 2987 4395
rect 2993 4391 2997 4395
rect 2958 4386 2962 4390
rect 2968 4386 2972 4390
rect 2978 4386 2982 4390
rect 2988 4386 2992 4390
rect 2953 4381 2957 4385
rect 2963 4381 2967 4385
rect 2973 4381 2977 4385
rect 2983 4381 2987 4385
rect 2993 4381 2997 4385
rect 2958 4376 2962 4380
rect 2968 4376 2972 4380
rect 2978 4376 2982 4380
rect 2988 4376 2992 4380
rect 2953 4371 2957 4375
rect 2963 4371 2967 4375
rect 2973 4371 2977 4375
rect 2983 4371 2987 4375
rect 2993 4371 2997 4375
rect 2958 4366 2962 4370
rect 2968 4366 2972 4370
rect 2978 4366 2982 4370
rect 2988 4366 2992 4370
rect 2953 4361 2957 4365
rect 2963 4361 2967 4365
rect 2973 4361 2977 4365
rect 2983 4361 2987 4365
rect 2993 4361 2997 4365
rect 3101 4462 3105 4466
rect 3108 4462 3112 4466
rect 3113 4462 3117 4466
rect 3118 4462 3122 4466
rect 3123 4462 3127 4466
rect 3128 4462 3132 4466
rect 3133 4462 3137 4466
rect 3138 4462 3142 4466
rect 3143 4462 3147 4466
rect 3148 4462 3152 4466
rect 3153 4462 3157 4466
rect 3158 4462 3162 4466
rect 3165 4462 3169 4466
rect 3118 4446 3122 4450
rect 3128 4446 3132 4450
rect 3138 4446 3142 4450
rect 3148 4446 3152 4450
rect 3113 4441 3117 4445
rect 3123 4441 3127 4445
rect 3133 4441 3137 4445
rect 3143 4441 3147 4445
rect 3153 4441 3157 4445
rect 3118 4436 3122 4440
rect 3128 4436 3132 4440
rect 3138 4436 3142 4440
rect 3148 4436 3152 4440
rect 3113 4431 3117 4435
rect 3123 4431 3127 4435
rect 3133 4431 3137 4435
rect 3143 4431 3147 4435
rect 3153 4431 3157 4435
rect 3118 4426 3122 4430
rect 3128 4426 3132 4430
rect 3138 4426 3142 4430
rect 3148 4426 3152 4430
rect 3113 4421 3117 4425
rect 3123 4421 3127 4425
rect 3133 4421 3137 4425
rect 3143 4421 3147 4425
rect 3153 4421 3157 4425
rect 3118 4416 3122 4420
rect 3128 4416 3132 4420
rect 3138 4416 3142 4420
rect 3148 4416 3152 4420
rect 3113 4411 3117 4415
rect 3123 4411 3127 4415
rect 3133 4411 3137 4415
rect 3143 4411 3147 4415
rect 3153 4411 3157 4415
rect 3118 4406 3122 4410
rect 3128 4406 3132 4410
rect 3138 4406 3142 4410
rect 3148 4406 3152 4410
rect 3113 4401 3117 4405
rect 3123 4401 3127 4405
rect 3133 4401 3137 4405
rect 3143 4401 3147 4405
rect 3153 4401 3157 4405
rect 3118 4396 3122 4400
rect 3128 4396 3132 4400
rect 3138 4396 3142 4400
rect 3148 4396 3152 4400
rect 3113 4391 3117 4395
rect 3123 4391 3127 4395
rect 3133 4391 3137 4395
rect 3143 4391 3147 4395
rect 3153 4391 3157 4395
rect 3118 4386 3122 4390
rect 3128 4386 3132 4390
rect 3138 4386 3142 4390
rect 3148 4386 3152 4390
rect 3113 4381 3117 4385
rect 3123 4381 3127 4385
rect 3133 4381 3137 4385
rect 3143 4381 3147 4385
rect 3153 4381 3157 4385
rect 3118 4376 3122 4380
rect 3128 4376 3132 4380
rect 3138 4376 3142 4380
rect 3148 4376 3152 4380
rect 3113 4371 3117 4375
rect 3123 4371 3127 4375
rect 3133 4371 3137 4375
rect 3143 4371 3147 4375
rect 3153 4371 3157 4375
rect 3118 4366 3122 4370
rect 3128 4366 3132 4370
rect 3138 4366 3142 4370
rect 3148 4366 3152 4370
rect 3113 4361 3117 4365
rect 3123 4361 3127 4365
rect 3133 4361 3137 4365
rect 3143 4361 3147 4365
rect 3153 4361 3157 4365
rect 3664 4599 3668 4603
rect 3669 4599 3673 4603
rect 3250 4462 3254 4466
rect 3257 4462 3261 4466
rect 3262 4462 3266 4466
rect 3267 4462 3271 4466
rect 3272 4462 3276 4466
rect 3277 4462 3281 4466
rect 3282 4462 3286 4466
rect 3287 4462 3291 4466
rect 3292 4462 3296 4466
rect 3297 4462 3301 4466
rect 3302 4462 3306 4466
rect 3307 4462 3311 4466
rect 3314 4462 3318 4466
rect 3267 4446 3271 4450
rect 3277 4446 3281 4450
rect 3287 4446 3291 4450
rect 3297 4446 3301 4450
rect 3262 4441 3266 4445
rect 3272 4441 3276 4445
rect 3282 4441 3286 4445
rect 3292 4441 3296 4445
rect 3302 4441 3306 4445
rect 3267 4436 3271 4440
rect 3277 4436 3281 4440
rect 3287 4436 3291 4440
rect 3297 4436 3301 4440
rect 3262 4431 3266 4435
rect 3272 4431 3276 4435
rect 3282 4431 3286 4435
rect 3292 4431 3296 4435
rect 3302 4431 3306 4435
rect 3267 4426 3271 4430
rect 3277 4426 3281 4430
rect 3287 4426 3291 4430
rect 3297 4426 3301 4430
rect 3262 4421 3266 4425
rect 3272 4421 3276 4425
rect 3282 4421 3286 4425
rect 3292 4421 3296 4425
rect 3302 4421 3306 4425
rect 3267 4416 3271 4420
rect 3277 4416 3281 4420
rect 3287 4416 3291 4420
rect 3297 4416 3301 4420
rect 3262 4411 3266 4415
rect 3272 4411 3276 4415
rect 3282 4411 3286 4415
rect 3292 4411 3296 4415
rect 3302 4411 3306 4415
rect 3267 4406 3271 4410
rect 3277 4406 3281 4410
rect 3287 4406 3291 4410
rect 3297 4406 3301 4410
rect 3262 4401 3266 4405
rect 3272 4401 3276 4405
rect 3282 4401 3286 4405
rect 3292 4401 3296 4405
rect 3302 4401 3306 4405
rect 3267 4396 3271 4400
rect 3277 4396 3281 4400
rect 3287 4396 3291 4400
rect 3297 4396 3301 4400
rect 3262 4391 3266 4395
rect 3272 4391 3276 4395
rect 3282 4391 3286 4395
rect 3292 4391 3296 4395
rect 3302 4391 3306 4395
rect 3267 4386 3271 4390
rect 3277 4386 3281 4390
rect 3287 4386 3291 4390
rect 3297 4386 3301 4390
rect 3262 4381 3266 4385
rect 3272 4381 3276 4385
rect 3282 4381 3286 4385
rect 3292 4381 3296 4385
rect 3302 4381 3306 4385
rect 3267 4376 3271 4380
rect 3277 4376 3281 4380
rect 3287 4376 3291 4380
rect 3297 4376 3301 4380
rect 3262 4371 3266 4375
rect 3272 4371 3276 4375
rect 3282 4371 3286 4375
rect 3292 4371 3296 4375
rect 3302 4371 3306 4375
rect 3267 4366 3271 4370
rect 3277 4366 3281 4370
rect 3287 4366 3291 4370
rect 3297 4366 3301 4370
rect 3262 4361 3266 4365
rect 3272 4361 3276 4365
rect 3282 4361 3286 4365
rect 3292 4361 3296 4365
rect 3302 4361 3306 4365
rect 3410 4462 3414 4466
rect 3417 4462 3421 4466
rect 3422 4462 3426 4466
rect 3427 4462 3431 4466
rect 3432 4462 3436 4466
rect 3437 4462 3441 4466
rect 3442 4462 3446 4466
rect 3447 4462 3451 4466
rect 3452 4462 3456 4466
rect 3457 4462 3461 4466
rect 3462 4462 3466 4466
rect 3467 4462 3471 4466
rect 3474 4462 3478 4466
rect 3427 4446 3431 4450
rect 3437 4446 3441 4450
rect 3447 4446 3451 4450
rect 3457 4446 3461 4450
rect 3422 4441 3426 4445
rect 3432 4441 3436 4445
rect 3442 4441 3446 4445
rect 3452 4441 3456 4445
rect 3462 4441 3466 4445
rect 3427 4436 3431 4440
rect 3437 4436 3441 4440
rect 3447 4436 3451 4440
rect 3457 4436 3461 4440
rect 3422 4431 3426 4435
rect 3432 4431 3436 4435
rect 3442 4431 3446 4435
rect 3452 4431 3456 4435
rect 3462 4431 3466 4435
rect 3427 4426 3431 4430
rect 3437 4426 3441 4430
rect 3447 4426 3451 4430
rect 3457 4426 3461 4430
rect 3422 4421 3426 4425
rect 3432 4421 3436 4425
rect 3442 4421 3446 4425
rect 3452 4421 3456 4425
rect 3462 4421 3466 4425
rect 3427 4416 3431 4420
rect 3437 4416 3441 4420
rect 3447 4416 3451 4420
rect 3457 4416 3461 4420
rect 3422 4411 3426 4415
rect 3432 4411 3436 4415
rect 3442 4411 3446 4415
rect 3452 4411 3456 4415
rect 3462 4411 3466 4415
rect 3427 4406 3431 4410
rect 3437 4406 3441 4410
rect 3447 4406 3451 4410
rect 3457 4406 3461 4410
rect 3422 4401 3426 4405
rect 3432 4401 3436 4405
rect 3442 4401 3446 4405
rect 3452 4401 3456 4405
rect 3462 4401 3466 4405
rect 3427 4396 3431 4400
rect 3437 4396 3441 4400
rect 3447 4396 3451 4400
rect 3457 4396 3461 4400
rect 3422 4391 3426 4395
rect 3432 4391 3436 4395
rect 3442 4391 3446 4395
rect 3452 4391 3456 4395
rect 3462 4391 3466 4395
rect 3427 4386 3431 4390
rect 3437 4386 3441 4390
rect 3447 4386 3451 4390
rect 3457 4386 3461 4390
rect 3422 4381 3426 4385
rect 3432 4381 3436 4385
rect 3442 4381 3446 4385
rect 3452 4381 3456 4385
rect 3462 4381 3466 4385
rect 3427 4376 3431 4380
rect 3437 4376 3441 4380
rect 3447 4376 3451 4380
rect 3457 4376 3461 4380
rect 3422 4371 3426 4375
rect 3432 4371 3436 4375
rect 3442 4371 3446 4375
rect 3452 4371 3456 4375
rect 3462 4371 3466 4375
rect 3427 4366 3431 4370
rect 3437 4366 3441 4370
rect 3447 4366 3451 4370
rect 3457 4366 3461 4370
rect 3422 4361 3426 4365
rect 3432 4361 3436 4365
rect 3442 4361 3446 4365
rect 3452 4361 3456 4365
rect 3462 4361 3466 4365
rect 3559 4462 3563 4466
rect 3566 4462 3570 4466
rect 3571 4462 3575 4466
rect 3576 4462 3580 4466
rect 3581 4462 3585 4466
rect 3586 4462 3590 4466
rect 3591 4462 3595 4466
rect 3596 4462 3600 4466
rect 3601 4462 3605 4466
rect 3606 4462 3610 4466
rect 3611 4462 3615 4466
rect 3616 4462 3620 4466
rect 3623 4462 3627 4466
rect 3576 4446 3580 4450
rect 3586 4446 3590 4450
rect 3596 4446 3600 4450
rect 3606 4446 3610 4450
rect 3571 4441 3575 4445
rect 3581 4441 3585 4445
rect 3591 4441 3595 4445
rect 3601 4441 3605 4445
rect 3611 4441 3615 4445
rect 3576 4436 3580 4440
rect 3586 4436 3590 4440
rect 3596 4436 3600 4440
rect 3606 4436 3610 4440
rect 3571 4431 3575 4435
rect 3581 4431 3585 4435
rect 3591 4431 3595 4435
rect 3601 4431 3605 4435
rect 3611 4431 3615 4435
rect 3576 4426 3580 4430
rect 3586 4426 3590 4430
rect 3596 4426 3600 4430
rect 3606 4426 3610 4430
rect 3571 4421 3575 4425
rect 3581 4421 3585 4425
rect 3591 4421 3595 4425
rect 3601 4421 3605 4425
rect 3611 4421 3615 4425
rect 3576 4416 3580 4420
rect 3586 4416 3590 4420
rect 3596 4416 3600 4420
rect 3606 4416 3610 4420
rect 3571 4411 3575 4415
rect 3581 4411 3585 4415
rect 3591 4411 3595 4415
rect 3601 4411 3605 4415
rect 3611 4411 3615 4415
rect 3576 4406 3580 4410
rect 3586 4406 3590 4410
rect 3596 4406 3600 4410
rect 3606 4406 3610 4410
rect 3571 4401 3575 4405
rect 3581 4401 3585 4405
rect 3591 4401 3595 4405
rect 3601 4401 3605 4405
rect 3611 4401 3615 4405
rect 3576 4396 3580 4400
rect 3586 4396 3590 4400
rect 3596 4396 3600 4400
rect 3606 4396 3610 4400
rect 3571 4391 3575 4395
rect 3581 4391 3585 4395
rect 3591 4391 3595 4395
rect 3601 4391 3605 4395
rect 3611 4391 3615 4395
rect 3576 4386 3580 4390
rect 3586 4386 3590 4390
rect 3596 4386 3600 4390
rect 3606 4386 3610 4390
rect 3571 4381 3575 4385
rect 3581 4381 3585 4385
rect 3591 4381 3595 4385
rect 3601 4381 3605 4385
rect 3611 4381 3615 4385
rect 3576 4376 3580 4380
rect 3586 4376 3590 4380
rect 3596 4376 3600 4380
rect 3606 4376 3610 4380
rect 3571 4371 3575 4375
rect 3581 4371 3585 4375
rect 3591 4371 3595 4375
rect 3601 4371 3605 4375
rect 3611 4371 3615 4375
rect 3576 4366 3580 4370
rect 3586 4366 3590 4370
rect 3596 4366 3600 4370
rect 3606 4366 3610 4370
rect 3571 4361 3575 4365
rect 3581 4361 3585 4365
rect 3591 4361 3595 4365
rect 3601 4361 3605 4365
rect 3611 4361 3615 4365
rect 3834 4619 3838 4623
rect 3839 4619 3843 4623
rect 3844 4619 3848 4623
rect 3849 4619 3853 4623
rect 3834 4609 3838 4613
rect 3839 4609 3843 4613
rect 3844 4609 3848 4613
rect 3849 4609 3853 4613
rect 3834 4599 3838 4603
rect 3839 4599 3843 4603
rect 3844 4599 3848 4603
rect 3849 4599 3853 4603
rect 3799 4574 3803 4578
rect 3804 4574 3808 4578
rect 3799 4569 3803 4573
rect 3804 4569 3808 4573
rect 3799 4564 3803 4568
rect 3804 4564 3808 4568
rect 3799 4559 3803 4563
rect 3804 4559 3808 4563
rect 3799 4554 3803 4558
rect 3804 4554 3808 4558
rect 3799 4549 3803 4553
rect 3804 4549 3808 4553
rect 3834 4573 3838 4577
rect 3839 4573 3843 4577
rect 3844 4573 3848 4577
rect 3849 4573 3853 4577
rect 3834 4563 3838 4567
rect 3839 4563 3843 4567
rect 3844 4563 3848 4567
rect 3849 4563 3853 4567
rect 3834 4553 3838 4557
rect 3839 4553 3843 4557
rect 3844 4553 3848 4557
rect 3849 4553 3853 4557
rect 3799 4544 3803 4548
rect 3804 4544 3808 4548
rect 3799 4539 3803 4543
rect 3804 4539 3808 4543
rect 3799 4534 3803 4538
rect 3804 4534 3808 4538
rect 3799 4529 3803 4533
rect 3804 4529 3808 4533
rect 3799 4524 3803 4528
rect 3804 4524 3808 4528
rect 3799 4519 3803 4523
rect 3804 4519 3808 4523
rect 3799 4514 3803 4518
rect 3804 4514 3808 4518
rect 3719 4462 3723 4466
rect 3726 4462 3730 4466
rect 3731 4462 3735 4466
rect 3736 4462 3740 4466
rect 3741 4462 3745 4466
rect 3746 4462 3750 4466
rect 3751 4462 3755 4466
rect 3756 4462 3760 4466
rect 3761 4462 3765 4466
rect 3766 4462 3770 4466
rect 3771 4462 3775 4466
rect 3776 4462 3780 4466
rect 3783 4462 3787 4466
rect 3736 4446 3740 4450
rect 3746 4446 3750 4450
rect 3756 4446 3760 4450
rect 3766 4446 3770 4450
rect 3731 4441 3735 4445
rect 3741 4441 3745 4445
rect 3751 4441 3755 4445
rect 3761 4441 3765 4445
rect 3771 4441 3775 4445
rect 3736 4436 3740 4440
rect 3746 4436 3750 4440
rect 3756 4436 3760 4440
rect 3766 4436 3770 4440
rect 3731 4431 3735 4435
rect 3741 4431 3745 4435
rect 3751 4431 3755 4435
rect 3761 4431 3765 4435
rect 3771 4431 3775 4435
rect 3736 4426 3740 4430
rect 3746 4426 3750 4430
rect 3756 4426 3760 4430
rect 3766 4426 3770 4430
rect 3731 4421 3735 4425
rect 3741 4421 3745 4425
rect 3751 4421 3755 4425
rect 3761 4421 3765 4425
rect 3771 4421 3775 4425
rect 3736 4416 3740 4420
rect 3746 4416 3750 4420
rect 3756 4416 3760 4420
rect 3766 4416 3770 4420
rect 3731 4411 3735 4415
rect 3741 4411 3745 4415
rect 3751 4411 3755 4415
rect 3761 4411 3765 4415
rect 3771 4411 3775 4415
rect 3736 4406 3740 4410
rect 3746 4406 3750 4410
rect 3756 4406 3760 4410
rect 3766 4406 3770 4410
rect 3731 4401 3735 4405
rect 3741 4401 3745 4405
rect 3751 4401 3755 4405
rect 3761 4401 3765 4405
rect 3771 4401 3775 4405
rect 3736 4396 3740 4400
rect 3746 4396 3750 4400
rect 3756 4396 3760 4400
rect 3766 4396 3770 4400
rect 3731 4391 3735 4395
rect 3741 4391 3745 4395
rect 3751 4391 3755 4395
rect 3761 4391 3765 4395
rect 3771 4391 3775 4395
rect 3736 4386 3740 4390
rect 3746 4386 3750 4390
rect 3756 4386 3760 4390
rect 3766 4386 3770 4390
rect 3731 4381 3735 4385
rect 3741 4381 3745 4385
rect 3751 4381 3755 4385
rect 3761 4381 3765 4385
rect 3771 4381 3775 4385
rect 3736 4376 3740 4380
rect 3746 4376 3750 4380
rect 3756 4376 3760 4380
rect 3766 4376 3770 4380
rect 3731 4371 3735 4375
rect 3741 4371 3745 4375
rect 3751 4371 3755 4375
rect 3761 4371 3765 4375
rect 3771 4371 3775 4375
rect 3736 4366 3740 4370
rect 3746 4366 3750 4370
rect 3756 4366 3760 4370
rect 3766 4366 3770 4370
rect 3731 4361 3735 4365
rect 3741 4361 3745 4365
rect 3751 4361 3755 4365
rect 3761 4361 3765 4365
rect 3771 4361 3775 4365
rect 1158 4328 1162 4332
rect 1165 4328 1169 4332
rect 1172 4328 1176 4332
rect 1179 4328 1183 4332
rect 1186 4328 1190 4332
rect 1193 4328 1197 4332
rect 1200 4328 1204 4332
rect 1207 4328 1211 4332
rect 1214 4328 1218 4332
rect 1221 4328 1225 4332
rect 1228 4328 1232 4332
rect 1235 4328 1239 4332
rect 1242 4328 1246 4332
rect 1158 4323 1162 4327
rect 1165 4323 1169 4327
rect 1172 4323 1176 4327
rect 1179 4323 1183 4327
rect 1186 4323 1190 4327
rect 1193 4323 1197 4327
rect 1200 4323 1204 4327
rect 1207 4323 1211 4327
rect 1214 4323 1218 4327
rect 1221 4323 1225 4327
rect 1228 4323 1232 4327
rect 1235 4323 1239 4327
rect 1242 4323 1246 4327
rect 1158 4318 1162 4322
rect 1165 4318 1169 4322
rect 1172 4318 1176 4322
rect 1179 4318 1183 4322
rect 1186 4318 1190 4322
rect 1193 4318 1197 4322
rect 1200 4318 1204 4322
rect 1207 4318 1211 4322
rect 1214 4318 1218 4322
rect 1221 4318 1225 4322
rect 1228 4318 1232 4322
rect 1235 4318 1239 4322
rect 1242 4318 1246 4322
rect 1467 4328 1471 4332
rect 1474 4328 1478 4332
rect 1481 4328 1485 4332
rect 1488 4328 1492 4332
rect 1495 4328 1499 4332
rect 1502 4328 1506 4332
rect 1509 4328 1513 4332
rect 1516 4328 1520 4332
rect 1523 4328 1527 4332
rect 1530 4328 1534 4332
rect 1537 4328 1541 4332
rect 1544 4328 1548 4332
rect 1551 4328 1555 4332
rect 1467 4323 1471 4327
rect 1474 4323 1478 4327
rect 1481 4323 1485 4327
rect 1488 4323 1492 4327
rect 1495 4323 1499 4327
rect 1502 4323 1506 4327
rect 1509 4323 1513 4327
rect 1516 4323 1520 4327
rect 1523 4323 1527 4327
rect 1530 4323 1534 4327
rect 1537 4323 1541 4327
rect 1544 4323 1548 4327
rect 1551 4323 1555 4327
rect 1158 4313 1162 4317
rect 1165 4313 1169 4317
rect 1172 4313 1176 4317
rect 1179 4313 1183 4317
rect 1186 4313 1190 4317
rect 1193 4313 1197 4317
rect 1200 4313 1204 4317
rect 1207 4313 1211 4317
rect 1214 4313 1218 4317
rect 1221 4313 1225 4317
rect 1228 4313 1232 4317
rect 1235 4313 1239 4317
rect 1242 4313 1246 4317
rect 1467 4318 1471 4322
rect 1474 4318 1478 4322
rect 1481 4318 1485 4322
rect 1488 4318 1492 4322
rect 1495 4318 1499 4322
rect 1502 4318 1506 4322
rect 1509 4318 1513 4322
rect 1516 4318 1520 4322
rect 1523 4318 1527 4322
rect 1530 4318 1534 4322
rect 1537 4318 1541 4322
rect 1544 4318 1548 4322
rect 1551 4318 1555 4322
rect 1776 4328 1780 4332
rect 1783 4328 1787 4332
rect 1790 4328 1794 4332
rect 1797 4328 1801 4332
rect 1804 4328 1808 4332
rect 1811 4328 1815 4332
rect 1818 4328 1822 4332
rect 1825 4328 1829 4332
rect 1832 4328 1836 4332
rect 1839 4328 1843 4332
rect 1846 4328 1850 4332
rect 1853 4328 1857 4332
rect 1860 4328 1864 4332
rect 1776 4323 1780 4327
rect 1783 4323 1787 4327
rect 1790 4323 1794 4327
rect 1797 4323 1801 4327
rect 1804 4323 1808 4327
rect 1811 4323 1815 4327
rect 1818 4323 1822 4327
rect 1825 4323 1829 4327
rect 1832 4323 1836 4327
rect 1839 4323 1843 4327
rect 1846 4323 1850 4327
rect 1853 4323 1857 4327
rect 1860 4323 1864 4327
rect 1467 4313 1471 4317
rect 1474 4313 1478 4317
rect 1481 4313 1485 4317
rect 1488 4313 1492 4317
rect 1495 4313 1499 4317
rect 1502 4313 1506 4317
rect 1509 4313 1513 4317
rect 1516 4313 1520 4317
rect 1523 4313 1527 4317
rect 1530 4313 1534 4317
rect 1537 4313 1541 4317
rect 1544 4313 1548 4317
rect 1551 4313 1555 4317
rect 1776 4318 1780 4322
rect 1783 4318 1787 4322
rect 1790 4318 1794 4322
rect 1797 4318 1801 4322
rect 1804 4318 1808 4322
rect 1811 4318 1815 4322
rect 1818 4318 1822 4322
rect 1825 4318 1829 4322
rect 1832 4318 1836 4322
rect 1839 4318 1843 4322
rect 1846 4318 1850 4322
rect 1853 4318 1857 4322
rect 1860 4318 1864 4322
rect 2085 4328 2089 4332
rect 2092 4328 2096 4332
rect 2099 4328 2103 4332
rect 2106 4328 2110 4332
rect 2113 4328 2117 4332
rect 2120 4328 2124 4332
rect 2127 4328 2131 4332
rect 2134 4328 2138 4332
rect 2141 4328 2145 4332
rect 2148 4328 2152 4332
rect 2155 4328 2159 4332
rect 2162 4328 2166 4332
rect 2169 4328 2173 4332
rect 2085 4323 2089 4327
rect 2092 4323 2096 4327
rect 2099 4323 2103 4327
rect 2106 4323 2110 4327
rect 2113 4323 2117 4327
rect 2120 4323 2124 4327
rect 2127 4323 2131 4327
rect 2134 4323 2138 4327
rect 2141 4323 2145 4327
rect 2148 4323 2152 4327
rect 2155 4323 2159 4327
rect 2162 4323 2166 4327
rect 2169 4323 2173 4327
rect 1776 4313 1780 4317
rect 1783 4313 1787 4317
rect 1790 4313 1794 4317
rect 1797 4313 1801 4317
rect 1804 4313 1808 4317
rect 1811 4313 1815 4317
rect 1818 4313 1822 4317
rect 1825 4313 1829 4317
rect 1832 4313 1836 4317
rect 1839 4313 1843 4317
rect 1846 4313 1850 4317
rect 1853 4313 1857 4317
rect 1860 4313 1864 4317
rect 2085 4318 2089 4322
rect 2092 4318 2096 4322
rect 2099 4318 2103 4322
rect 2106 4318 2110 4322
rect 2113 4318 2117 4322
rect 2120 4318 2124 4322
rect 2127 4318 2131 4322
rect 2134 4318 2138 4322
rect 2141 4318 2145 4322
rect 2148 4318 2152 4322
rect 2155 4318 2159 4322
rect 2162 4318 2166 4322
rect 2169 4318 2173 4322
rect 2394 4328 2398 4332
rect 2401 4328 2405 4332
rect 2408 4328 2412 4332
rect 2415 4328 2419 4332
rect 2422 4328 2426 4332
rect 2429 4328 2433 4332
rect 2436 4328 2440 4332
rect 2443 4328 2447 4332
rect 2450 4328 2454 4332
rect 2457 4328 2461 4332
rect 2464 4328 2468 4332
rect 2471 4328 2475 4332
rect 2478 4328 2482 4332
rect 2394 4323 2398 4327
rect 2401 4323 2405 4327
rect 2408 4323 2412 4327
rect 2415 4323 2419 4327
rect 2422 4323 2426 4327
rect 2429 4323 2433 4327
rect 2436 4323 2440 4327
rect 2443 4323 2447 4327
rect 2450 4323 2454 4327
rect 2457 4323 2461 4327
rect 2464 4323 2468 4327
rect 2471 4323 2475 4327
rect 2478 4323 2482 4327
rect 2085 4313 2089 4317
rect 2092 4313 2096 4317
rect 2099 4313 2103 4317
rect 2106 4313 2110 4317
rect 2113 4313 2117 4317
rect 2120 4313 2124 4317
rect 2127 4313 2131 4317
rect 2134 4313 2138 4317
rect 2141 4313 2145 4317
rect 2148 4313 2152 4317
rect 2155 4313 2159 4317
rect 2162 4313 2166 4317
rect 2169 4313 2173 4317
rect 2394 4318 2398 4322
rect 2401 4318 2405 4322
rect 2408 4318 2412 4322
rect 2415 4318 2419 4322
rect 2422 4318 2426 4322
rect 2429 4318 2433 4322
rect 2436 4318 2440 4322
rect 2443 4318 2447 4322
rect 2450 4318 2454 4322
rect 2457 4318 2461 4322
rect 2464 4318 2468 4322
rect 2471 4318 2475 4322
rect 2478 4318 2482 4322
rect 2703 4328 2707 4332
rect 2710 4328 2714 4332
rect 2717 4328 2721 4332
rect 2724 4328 2728 4332
rect 2731 4328 2735 4332
rect 2738 4328 2742 4332
rect 2745 4328 2749 4332
rect 2752 4328 2756 4332
rect 2759 4328 2763 4332
rect 2766 4328 2770 4332
rect 2773 4328 2777 4332
rect 2780 4328 2784 4332
rect 2787 4328 2791 4332
rect 2703 4323 2707 4327
rect 2710 4323 2714 4327
rect 2717 4323 2721 4327
rect 2724 4323 2728 4327
rect 2731 4323 2735 4327
rect 2738 4323 2742 4327
rect 2745 4323 2749 4327
rect 2752 4323 2756 4327
rect 2759 4323 2763 4327
rect 2766 4323 2770 4327
rect 2773 4323 2777 4327
rect 2780 4323 2784 4327
rect 2787 4323 2791 4327
rect 2394 4313 2398 4317
rect 2401 4313 2405 4317
rect 2408 4313 2412 4317
rect 2415 4313 2419 4317
rect 2422 4313 2426 4317
rect 2429 4313 2433 4317
rect 2436 4313 2440 4317
rect 2443 4313 2447 4317
rect 2450 4313 2454 4317
rect 2457 4313 2461 4317
rect 2464 4313 2468 4317
rect 2471 4313 2475 4317
rect 2478 4313 2482 4317
rect 2703 4318 2707 4322
rect 2710 4318 2714 4322
rect 2717 4318 2721 4322
rect 2724 4318 2728 4322
rect 2731 4318 2735 4322
rect 2738 4318 2742 4322
rect 2745 4318 2749 4322
rect 2752 4318 2756 4322
rect 2759 4318 2763 4322
rect 2766 4318 2770 4322
rect 2773 4318 2777 4322
rect 2780 4318 2784 4322
rect 2787 4318 2791 4322
rect 3012 4328 3016 4332
rect 3019 4328 3023 4332
rect 3026 4328 3030 4332
rect 3033 4328 3037 4332
rect 3040 4328 3044 4332
rect 3047 4328 3051 4332
rect 3054 4328 3058 4332
rect 3061 4328 3065 4332
rect 3068 4328 3072 4332
rect 3075 4328 3079 4332
rect 3082 4328 3086 4332
rect 3089 4328 3093 4332
rect 3096 4328 3100 4332
rect 3012 4323 3016 4327
rect 3019 4323 3023 4327
rect 3026 4323 3030 4327
rect 3033 4323 3037 4327
rect 3040 4323 3044 4327
rect 3047 4323 3051 4327
rect 3054 4323 3058 4327
rect 3061 4323 3065 4327
rect 3068 4323 3072 4327
rect 3075 4323 3079 4327
rect 3082 4323 3086 4327
rect 3089 4323 3093 4327
rect 3096 4323 3100 4327
rect 2703 4313 2707 4317
rect 2710 4313 2714 4317
rect 2717 4313 2721 4317
rect 2724 4313 2728 4317
rect 2731 4313 2735 4317
rect 2738 4313 2742 4317
rect 2745 4313 2749 4317
rect 2752 4313 2756 4317
rect 2759 4313 2763 4317
rect 2766 4313 2770 4317
rect 2773 4313 2777 4317
rect 2780 4313 2784 4317
rect 2787 4313 2791 4317
rect 3012 4318 3016 4322
rect 3019 4318 3023 4322
rect 3026 4318 3030 4322
rect 3033 4318 3037 4322
rect 3040 4318 3044 4322
rect 3047 4318 3051 4322
rect 3054 4318 3058 4322
rect 3061 4318 3065 4322
rect 3068 4318 3072 4322
rect 3075 4318 3079 4322
rect 3082 4318 3086 4322
rect 3089 4318 3093 4322
rect 3096 4318 3100 4322
rect 3321 4328 3325 4332
rect 3328 4328 3332 4332
rect 3335 4328 3339 4332
rect 3342 4328 3346 4332
rect 3349 4328 3353 4332
rect 3356 4328 3360 4332
rect 3363 4328 3367 4332
rect 3370 4328 3374 4332
rect 3377 4328 3381 4332
rect 3384 4328 3388 4332
rect 3391 4328 3395 4332
rect 3398 4328 3402 4332
rect 3405 4328 3409 4332
rect 3321 4323 3325 4327
rect 3328 4323 3332 4327
rect 3335 4323 3339 4327
rect 3342 4323 3346 4327
rect 3349 4323 3353 4327
rect 3356 4323 3360 4327
rect 3363 4323 3367 4327
rect 3370 4323 3374 4327
rect 3377 4323 3381 4327
rect 3384 4323 3388 4327
rect 3391 4323 3395 4327
rect 3398 4323 3402 4327
rect 3405 4323 3409 4327
rect 3012 4313 3016 4317
rect 3019 4313 3023 4317
rect 3026 4313 3030 4317
rect 3033 4313 3037 4317
rect 3040 4313 3044 4317
rect 3047 4313 3051 4317
rect 3054 4313 3058 4317
rect 3061 4313 3065 4317
rect 3068 4313 3072 4317
rect 3075 4313 3079 4317
rect 3082 4313 3086 4317
rect 3089 4313 3093 4317
rect 3096 4313 3100 4317
rect 3321 4318 3325 4322
rect 3328 4318 3332 4322
rect 3335 4318 3339 4322
rect 3342 4318 3346 4322
rect 3349 4318 3353 4322
rect 3356 4318 3360 4322
rect 3363 4318 3367 4322
rect 3370 4318 3374 4322
rect 3377 4318 3381 4322
rect 3384 4318 3388 4322
rect 3391 4318 3395 4322
rect 3398 4318 3402 4322
rect 3405 4318 3409 4322
rect 3630 4328 3634 4332
rect 3637 4328 3641 4332
rect 3644 4328 3648 4332
rect 3651 4328 3655 4332
rect 3658 4328 3662 4332
rect 3665 4328 3669 4332
rect 3672 4328 3676 4332
rect 3679 4328 3683 4332
rect 3686 4328 3690 4332
rect 3693 4328 3697 4332
rect 3700 4328 3704 4332
rect 3707 4328 3711 4332
rect 3714 4328 3718 4332
rect 3630 4323 3634 4327
rect 3637 4323 3641 4327
rect 3644 4323 3648 4327
rect 3651 4323 3655 4327
rect 3658 4323 3662 4327
rect 3665 4323 3669 4327
rect 3672 4323 3676 4327
rect 3679 4323 3683 4327
rect 3686 4323 3690 4327
rect 3693 4323 3697 4327
rect 3700 4323 3704 4327
rect 3707 4323 3711 4327
rect 3714 4323 3718 4327
rect 3321 4313 3325 4317
rect 3328 4313 3332 4317
rect 3335 4313 3339 4317
rect 3342 4313 3346 4317
rect 3349 4313 3353 4317
rect 3356 4313 3360 4317
rect 3363 4313 3367 4317
rect 3370 4313 3374 4317
rect 3377 4313 3381 4317
rect 3384 4313 3388 4317
rect 3391 4313 3395 4317
rect 3398 4313 3402 4317
rect 3405 4313 3409 4317
rect 3630 4318 3634 4322
rect 3637 4318 3641 4322
rect 3644 4318 3648 4322
rect 3651 4318 3655 4322
rect 3658 4318 3662 4322
rect 3665 4318 3669 4322
rect 3672 4318 3676 4322
rect 3679 4318 3683 4322
rect 3686 4318 3690 4322
rect 3693 4318 3697 4322
rect 3700 4318 3704 4322
rect 3707 4318 3711 4322
rect 3714 4318 3718 4322
rect 4484 4702 4488 4706
rect 4494 4702 4498 4706
rect 4504 4702 4508 4706
rect 4484 4697 4488 4701
rect 4494 4697 4498 4701
rect 4504 4697 4508 4701
rect 4484 4692 4488 4696
rect 4494 4692 4498 4696
rect 4504 4692 4508 4696
rect 4530 4707 4534 4711
rect 4540 4707 4544 4711
rect 4550 4707 4554 4711
rect 4530 4702 4534 4706
rect 4540 4702 4544 4706
rect 4550 4702 4554 4706
rect 4530 4697 4534 4701
rect 4540 4697 4544 4701
rect 4550 4697 4554 4701
rect 4530 4692 4534 4696
rect 4540 4692 4544 4696
rect 4550 4692 4554 4696
rect 4235 4619 4239 4623
rect 4240 4619 4244 4623
rect 4245 4619 4249 4623
rect 4250 4619 4254 4623
rect 4235 4609 4239 4613
rect 4240 4609 4244 4613
rect 4245 4609 4249 4613
rect 4250 4609 4254 4613
rect 4235 4599 4239 4603
rect 4240 4599 4244 4603
rect 4245 4599 4249 4603
rect 4250 4599 4254 4603
rect 4264 4619 4268 4623
rect 4269 4619 4273 4623
rect 4274 4619 4278 4623
rect 4279 4619 4283 4623
rect 4264 4609 4268 4613
rect 4269 4609 4273 4613
rect 4274 4609 4278 4613
rect 4279 4609 4283 4613
rect 4264 4599 4268 4603
rect 4269 4599 4273 4603
rect 4274 4599 4278 4603
rect 4279 4599 4283 4603
rect 4293 4619 4297 4623
rect 4298 4619 4302 4623
rect 4303 4619 4307 4623
rect 4308 4619 4312 4623
rect 4293 4609 4297 4613
rect 4298 4609 4302 4613
rect 4303 4609 4307 4613
rect 4308 4609 4312 4613
rect 4293 4599 4297 4603
rect 4298 4599 4302 4603
rect 4303 4599 4307 4603
rect 4308 4599 4312 4603
rect 4322 4619 4326 4623
rect 4327 4619 4331 4623
rect 4332 4619 4336 4623
rect 4337 4619 4341 4623
rect 4322 4609 4326 4613
rect 4327 4609 4331 4613
rect 4332 4609 4336 4613
rect 4337 4609 4341 4613
rect 4322 4599 4326 4603
rect 4327 4599 4331 4603
rect 4332 4599 4336 4603
rect 4337 4599 4341 4603
rect 4351 4619 4355 4623
rect 4356 4619 4360 4623
rect 4361 4619 4365 4623
rect 4366 4619 4370 4623
rect 4351 4609 4355 4613
rect 4356 4609 4360 4613
rect 4361 4609 4365 4613
rect 4366 4609 4370 4613
rect 4351 4599 4355 4603
rect 4356 4599 4360 4603
rect 4361 4599 4365 4603
rect 4366 4599 4370 4603
rect 4235 4573 4239 4577
rect 4240 4573 4244 4577
rect 4245 4573 4249 4577
rect 4250 4573 4254 4577
rect 4235 4563 4239 4567
rect 4240 4563 4244 4567
rect 4245 4563 4249 4567
rect 4250 4563 4254 4567
rect 4235 4553 4239 4557
rect 4240 4553 4244 4557
rect 4245 4553 4249 4557
rect 4250 4553 4254 4557
rect 4264 4573 4268 4577
rect 4269 4573 4273 4577
rect 4274 4573 4278 4577
rect 4279 4573 4283 4577
rect 4264 4563 4268 4567
rect 4269 4563 4273 4567
rect 4274 4563 4278 4567
rect 4279 4563 4283 4567
rect 4264 4553 4268 4557
rect 4269 4553 4273 4557
rect 4274 4553 4278 4557
rect 4279 4553 4283 4557
rect 4293 4573 4297 4577
rect 4298 4573 4302 4577
rect 4303 4573 4307 4577
rect 4308 4573 4312 4577
rect 4293 4563 4297 4567
rect 4298 4563 4302 4567
rect 4303 4563 4307 4567
rect 4308 4563 4312 4567
rect 4293 4553 4297 4557
rect 4298 4553 4302 4557
rect 4303 4553 4307 4557
rect 4308 4553 4312 4557
rect 4322 4573 4326 4577
rect 4327 4573 4331 4577
rect 4332 4573 4336 4577
rect 4337 4573 4341 4577
rect 4322 4563 4326 4567
rect 4327 4563 4331 4567
rect 4332 4563 4336 4567
rect 4337 4563 4341 4567
rect 4322 4553 4326 4557
rect 4327 4553 4331 4557
rect 4332 4553 4336 4557
rect 4337 4553 4341 4557
rect 4351 4573 4355 4577
rect 4356 4573 4360 4577
rect 4361 4573 4365 4577
rect 4366 4573 4370 4577
rect 4351 4563 4355 4567
rect 4356 4563 4360 4567
rect 4361 4563 4365 4567
rect 4366 4563 4370 4567
rect 4351 4553 4355 4557
rect 4356 4553 4360 4557
rect 4361 4553 4365 4557
rect 4366 4553 4370 4557
rect 3630 4313 3634 4317
rect 3637 4313 3641 4317
rect 3644 4313 3648 4317
rect 3651 4313 3655 4317
rect 3658 4313 3662 4317
rect 3665 4313 3669 4317
rect 3672 4313 3676 4317
rect 3679 4313 3683 4317
rect 3686 4313 3690 4317
rect 3693 4313 3697 4317
rect 3700 4313 3704 4317
rect 3707 4313 3711 4317
rect 3714 4313 3718 4317
<< metal2 >>
rect 1060 10290 1320 10293
rect 118 9786 1024 10280
rect 1060 10036 1063 10290
rect 1317 10036 1320 10290
rect 1060 10033 1320 10036
rect 1369 10290 1629 10293
rect 1369 10036 1372 10290
rect 1626 10036 1629 10290
rect 1369 10033 1629 10036
rect 1678 10290 1938 10293
rect 1678 10036 1681 10290
rect 1935 10036 1938 10290
rect 1678 10033 1938 10036
rect 1987 10290 2247 10293
rect 1987 10036 1990 10290
rect 2244 10036 2247 10290
rect 1987 10033 2247 10036
rect 2296 10290 2556 10293
rect 2296 10036 2299 10290
rect 2553 10036 2556 10290
rect 2296 10033 2556 10036
rect 2605 10290 2865 10293
rect 2605 10036 2608 10290
rect 2862 10036 2865 10290
rect 2605 10033 2865 10036
rect 2914 10290 3174 10293
rect 2914 10036 2917 10290
rect 3171 10036 3174 10290
rect 2914 10033 3174 10036
rect 3223 10290 3483 10293
rect 3223 10036 3226 10290
rect 3480 10036 3483 10290
rect 3223 10033 3483 10036
rect 3532 10290 3792 10293
rect 3532 10036 3535 10290
rect 3789 10036 3792 10290
rect 3532 10033 3792 10036
rect 3841 10290 4101 10293
rect 3841 10036 3844 10290
rect 4098 10036 4101 10290
rect 3841 10033 4101 10036
rect 1441 10001 1557 10002
rect 1441 9997 1454 10001
rect 1458 9997 1461 10001
rect 1465 9997 1468 10001
rect 1472 9997 1475 10001
rect 1479 9997 1482 10001
rect 1486 9997 1489 10001
rect 1493 9997 1496 10001
rect 1500 9997 1503 10001
rect 1507 9997 1510 10001
rect 1514 9997 1517 10001
rect 1521 9997 1524 10001
rect 1528 9997 1531 10001
rect 1535 9997 1538 10001
rect 1542 9997 1557 10001
rect 1441 9996 1557 9997
rect 1441 9993 1454 9996
rect 1451 9992 1454 9993
rect 1458 9992 1461 9996
rect 1465 9992 1468 9996
rect 1472 9992 1475 9996
rect 1479 9992 1482 9996
rect 1486 9992 1489 9996
rect 1493 9992 1496 9996
rect 1500 9992 1503 9996
rect 1507 9992 1510 9996
rect 1514 9992 1517 9996
rect 1521 9992 1524 9996
rect 1528 9992 1531 9996
rect 1535 9992 1538 9996
rect 1542 9993 1557 9996
rect 1750 10001 1866 10002
rect 1750 9997 1763 10001
rect 1767 9997 1770 10001
rect 1774 9997 1777 10001
rect 1781 9997 1784 10001
rect 1788 9997 1791 10001
rect 1795 9997 1798 10001
rect 1802 9997 1805 10001
rect 1809 9997 1812 10001
rect 1816 9997 1819 10001
rect 1823 9997 1826 10001
rect 1830 9997 1833 10001
rect 1837 9997 1840 10001
rect 1844 9997 1847 10001
rect 1851 9997 1866 10001
rect 1750 9996 1866 9997
rect 1750 9993 1763 9996
rect 1542 9992 1547 9993
rect 1451 9991 1547 9992
rect 1451 9987 1454 9991
rect 1458 9987 1461 9991
rect 1465 9987 1468 9991
rect 1472 9987 1475 9991
rect 1479 9987 1482 9991
rect 1486 9987 1489 9991
rect 1493 9987 1496 9991
rect 1500 9987 1503 9991
rect 1507 9987 1510 9991
rect 1514 9987 1517 9991
rect 1521 9987 1524 9991
rect 1528 9987 1531 9991
rect 1535 9987 1538 9991
rect 1542 9987 1547 9991
rect 1451 9986 1547 9987
rect 1451 9982 1454 9986
rect 1458 9982 1461 9986
rect 1465 9982 1468 9986
rect 1472 9982 1475 9986
rect 1479 9982 1482 9986
rect 1486 9982 1489 9986
rect 1493 9982 1496 9986
rect 1500 9982 1503 9986
rect 1507 9982 1510 9986
rect 1514 9982 1517 9986
rect 1521 9982 1524 9986
rect 1528 9982 1531 9986
rect 1535 9982 1538 9986
rect 1542 9982 1547 9986
rect 1451 9953 1547 9982
rect 1760 9992 1763 9993
rect 1767 9992 1770 9996
rect 1774 9992 1777 9996
rect 1781 9992 1784 9996
rect 1788 9992 1791 9996
rect 1795 9992 1798 9996
rect 1802 9992 1805 9996
rect 1809 9992 1812 9996
rect 1816 9992 1819 9996
rect 1823 9992 1826 9996
rect 1830 9992 1833 9996
rect 1837 9992 1840 9996
rect 1844 9992 1847 9996
rect 1851 9993 1866 9996
rect 2059 10001 2175 10002
rect 2059 9997 2072 10001
rect 2076 9997 2079 10001
rect 2083 9997 2086 10001
rect 2090 9997 2093 10001
rect 2097 9997 2100 10001
rect 2104 9997 2107 10001
rect 2111 9997 2114 10001
rect 2118 9997 2121 10001
rect 2125 9997 2128 10001
rect 2132 9997 2135 10001
rect 2139 9997 2142 10001
rect 2146 9997 2149 10001
rect 2153 9997 2156 10001
rect 2160 9997 2175 10001
rect 2059 9996 2175 9997
rect 2059 9993 2072 9996
rect 1851 9992 1856 9993
rect 1760 9991 1856 9992
rect 1760 9987 1763 9991
rect 1767 9987 1770 9991
rect 1774 9987 1777 9991
rect 1781 9987 1784 9991
rect 1788 9987 1791 9991
rect 1795 9987 1798 9991
rect 1802 9987 1805 9991
rect 1809 9987 1812 9991
rect 1816 9987 1819 9991
rect 1823 9987 1826 9991
rect 1830 9987 1833 9991
rect 1837 9987 1840 9991
rect 1844 9987 1847 9991
rect 1851 9987 1856 9991
rect 1760 9986 1856 9987
rect 1760 9982 1763 9986
rect 1767 9982 1770 9986
rect 1774 9982 1777 9986
rect 1781 9982 1784 9986
rect 1788 9982 1791 9986
rect 1795 9982 1798 9986
rect 1802 9982 1805 9986
rect 1809 9982 1812 9986
rect 1816 9982 1819 9986
rect 1823 9982 1826 9986
rect 1830 9982 1833 9986
rect 1837 9982 1840 9986
rect 1844 9982 1847 9986
rect 1851 9982 1856 9986
rect 1760 9953 1856 9982
rect 2069 9992 2072 9993
rect 2076 9992 2079 9996
rect 2083 9992 2086 9996
rect 2090 9992 2093 9996
rect 2097 9992 2100 9996
rect 2104 9992 2107 9996
rect 2111 9992 2114 9996
rect 2118 9992 2121 9996
rect 2125 9992 2128 9996
rect 2132 9992 2135 9996
rect 2139 9992 2142 9996
rect 2146 9992 2149 9996
rect 2153 9992 2156 9996
rect 2160 9993 2175 9996
rect 2368 10001 2484 10002
rect 2368 9997 2381 10001
rect 2385 9997 2388 10001
rect 2392 9997 2395 10001
rect 2399 9997 2402 10001
rect 2406 9997 2409 10001
rect 2413 9997 2416 10001
rect 2420 9997 2423 10001
rect 2427 9997 2430 10001
rect 2434 9997 2437 10001
rect 2441 9997 2444 10001
rect 2448 9997 2451 10001
rect 2455 9997 2458 10001
rect 2462 9997 2465 10001
rect 2469 9997 2484 10001
rect 2368 9996 2484 9997
rect 2368 9993 2381 9996
rect 2160 9992 2165 9993
rect 2069 9991 2165 9992
rect 2069 9987 2072 9991
rect 2076 9987 2079 9991
rect 2083 9987 2086 9991
rect 2090 9987 2093 9991
rect 2097 9987 2100 9991
rect 2104 9987 2107 9991
rect 2111 9987 2114 9991
rect 2118 9987 2121 9991
rect 2125 9987 2128 9991
rect 2132 9987 2135 9991
rect 2139 9987 2142 9991
rect 2146 9987 2149 9991
rect 2153 9987 2156 9991
rect 2160 9987 2165 9991
rect 2069 9986 2165 9987
rect 2069 9982 2072 9986
rect 2076 9982 2079 9986
rect 2083 9982 2086 9986
rect 2090 9982 2093 9986
rect 2097 9982 2100 9986
rect 2104 9982 2107 9986
rect 2111 9982 2114 9986
rect 2118 9982 2121 9986
rect 2125 9982 2128 9986
rect 2132 9982 2135 9986
rect 2139 9982 2142 9986
rect 2146 9982 2149 9986
rect 2153 9982 2156 9986
rect 2160 9982 2165 9986
rect 2069 9953 2165 9982
rect 2378 9992 2381 9993
rect 2385 9992 2388 9996
rect 2392 9992 2395 9996
rect 2399 9992 2402 9996
rect 2406 9992 2409 9996
rect 2413 9992 2416 9996
rect 2420 9992 2423 9996
rect 2427 9992 2430 9996
rect 2434 9992 2437 9996
rect 2441 9992 2444 9996
rect 2448 9992 2451 9996
rect 2455 9992 2458 9996
rect 2462 9992 2465 9996
rect 2469 9993 2484 9996
rect 2677 10001 2793 10002
rect 2677 9997 2690 10001
rect 2694 9997 2697 10001
rect 2701 9997 2704 10001
rect 2708 9997 2711 10001
rect 2715 9997 2718 10001
rect 2722 9997 2725 10001
rect 2729 9997 2732 10001
rect 2736 9997 2739 10001
rect 2743 9997 2746 10001
rect 2750 9997 2753 10001
rect 2757 9997 2760 10001
rect 2764 9997 2767 10001
rect 2771 9997 2774 10001
rect 2778 9997 2793 10001
rect 2677 9996 2793 9997
rect 2677 9993 2690 9996
rect 2469 9992 2474 9993
rect 2378 9991 2474 9992
rect 2378 9987 2381 9991
rect 2385 9987 2388 9991
rect 2392 9987 2395 9991
rect 2399 9987 2402 9991
rect 2406 9987 2409 9991
rect 2413 9987 2416 9991
rect 2420 9987 2423 9991
rect 2427 9987 2430 9991
rect 2434 9987 2437 9991
rect 2441 9987 2444 9991
rect 2448 9987 2451 9991
rect 2455 9987 2458 9991
rect 2462 9987 2465 9991
rect 2469 9987 2474 9991
rect 2378 9986 2474 9987
rect 2378 9982 2381 9986
rect 2385 9982 2388 9986
rect 2392 9982 2395 9986
rect 2399 9982 2402 9986
rect 2406 9982 2409 9986
rect 2413 9982 2416 9986
rect 2420 9982 2423 9986
rect 2427 9982 2430 9986
rect 2434 9982 2437 9986
rect 2441 9982 2444 9986
rect 2448 9982 2451 9986
rect 2455 9982 2458 9986
rect 2462 9982 2465 9986
rect 2469 9982 2474 9986
rect 2378 9953 2474 9982
rect 2687 9992 2690 9993
rect 2694 9992 2697 9996
rect 2701 9992 2704 9996
rect 2708 9992 2711 9996
rect 2715 9992 2718 9996
rect 2722 9992 2725 9996
rect 2729 9992 2732 9996
rect 2736 9992 2739 9996
rect 2743 9992 2746 9996
rect 2750 9992 2753 9996
rect 2757 9992 2760 9996
rect 2764 9992 2767 9996
rect 2771 9992 2774 9996
rect 2778 9993 2793 9996
rect 2986 10001 3102 10002
rect 2986 9997 2999 10001
rect 3003 9997 3006 10001
rect 3010 9997 3013 10001
rect 3017 9997 3020 10001
rect 3024 9997 3027 10001
rect 3031 9997 3034 10001
rect 3038 9997 3041 10001
rect 3045 9997 3048 10001
rect 3052 9997 3055 10001
rect 3059 9997 3062 10001
rect 3066 9997 3069 10001
rect 3073 9997 3076 10001
rect 3080 9997 3083 10001
rect 3087 9997 3102 10001
rect 2986 9996 3102 9997
rect 2986 9993 2999 9996
rect 2778 9992 2783 9993
rect 2687 9991 2783 9992
rect 2687 9987 2690 9991
rect 2694 9987 2697 9991
rect 2701 9987 2704 9991
rect 2708 9987 2711 9991
rect 2715 9987 2718 9991
rect 2722 9987 2725 9991
rect 2729 9987 2732 9991
rect 2736 9987 2739 9991
rect 2743 9987 2746 9991
rect 2750 9987 2753 9991
rect 2757 9987 2760 9991
rect 2764 9987 2767 9991
rect 2771 9987 2774 9991
rect 2778 9987 2783 9991
rect 2687 9986 2783 9987
rect 2687 9982 2690 9986
rect 2694 9982 2697 9986
rect 2701 9982 2704 9986
rect 2708 9982 2711 9986
rect 2715 9982 2718 9986
rect 2722 9982 2725 9986
rect 2729 9982 2732 9986
rect 2736 9982 2739 9986
rect 2743 9982 2746 9986
rect 2750 9982 2753 9986
rect 2757 9982 2760 9986
rect 2764 9982 2767 9986
rect 2771 9982 2774 9986
rect 2778 9982 2783 9986
rect 2687 9953 2783 9982
rect 2996 9992 2999 9993
rect 3003 9992 3006 9996
rect 3010 9992 3013 9996
rect 3017 9992 3020 9996
rect 3024 9992 3027 9996
rect 3031 9992 3034 9996
rect 3038 9992 3041 9996
rect 3045 9992 3048 9996
rect 3052 9992 3055 9996
rect 3059 9992 3062 9996
rect 3066 9992 3069 9996
rect 3073 9992 3076 9996
rect 3080 9992 3083 9996
rect 3087 9993 3102 9996
rect 3295 10001 3411 10002
rect 3295 9997 3308 10001
rect 3312 9997 3315 10001
rect 3319 9997 3322 10001
rect 3326 9997 3329 10001
rect 3333 9997 3336 10001
rect 3340 9997 3343 10001
rect 3347 9997 3350 10001
rect 3354 9997 3357 10001
rect 3361 9997 3364 10001
rect 3368 9997 3371 10001
rect 3375 9997 3378 10001
rect 3382 9997 3385 10001
rect 3389 9997 3392 10001
rect 3396 9997 3411 10001
rect 3295 9996 3411 9997
rect 3295 9993 3308 9996
rect 3087 9992 3092 9993
rect 2996 9991 3092 9992
rect 2996 9987 2999 9991
rect 3003 9987 3006 9991
rect 3010 9987 3013 9991
rect 3017 9987 3020 9991
rect 3024 9987 3027 9991
rect 3031 9987 3034 9991
rect 3038 9987 3041 9991
rect 3045 9987 3048 9991
rect 3052 9987 3055 9991
rect 3059 9987 3062 9991
rect 3066 9987 3069 9991
rect 3073 9987 3076 9991
rect 3080 9987 3083 9991
rect 3087 9987 3092 9991
rect 2996 9986 3092 9987
rect 2996 9982 2999 9986
rect 3003 9982 3006 9986
rect 3010 9982 3013 9986
rect 3017 9982 3020 9986
rect 3024 9982 3027 9986
rect 3031 9982 3034 9986
rect 3038 9982 3041 9986
rect 3045 9982 3048 9986
rect 3052 9982 3055 9986
rect 3059 9982 3062 9986
rect 3066 9982 3069 9986
rect 3073 9982 3076 9986
rect 3080 9982 3083 9986
rect 3087 9982 3092 9986
rect 2996 9953 3092 9982
rect 3305 9992 3308 9993
rect 3312 9992 3315 9996
rect 3319 9992 3322 9996
rect 3326 9992 3329 9996
rect 3333 9992 3336 9996
rect 3340 9992 3343 9996
rect 3347 9992 3350 9996
rect 3354 9992 3357 9996
rect 3361 9992 3364 9996
rect 3368 9992 3371 9996
rect 3375 9992 3378 9996
rect 3382 9992 3385 9996
rect 3389 9992 3392 9996
rect 3396 9993 3411 9996
rect 3604 10001 3720 10002
rect 3604 9997 3617 10001
rect 3621 9997 3624 10001
rect 3628 9997 3631 10001
rect 3635 9997 3638 10001
rect 3642 9997 3645 10001
rect 3649 9997 3652 10001
rect 3656 9997 3659 10001
rect 3663 9997 3666 10001
rect 3670 9997 3673 10001
rect 3677 9997 3680 10001
rect 3684 9997 3687 10001
rect 3691 9997 3694 10001
rect 3698 9997 3701 10001
rect 3705 9997 3720 10001
rect 3604 9996 3720 9997
rect 3604 9993 3617 9996
rect 3396 9992 3401 9993
rect 3305 9991 3401 9992
rect 3305 9987 3308 9991
rect 3312 9987 3315 9991
rect 3319 9987 3322 9991
rect 3326 9987 3329 9991
rect 3333 9987 3336 9991
rect 3340 9987 3343 9991
rect 3347 9987 3350 9991
rect 3354 9987 3357 9991
rect 3361 9987 3364 9991
rect 3368 9987 3371 9991
rect 3375 9987 3378 9991
rect 3382 9987 3385 9991
rect 3389 9987 3392 9991
rect 3396 9987 3401 9991
rect 3305 9986 3401 9987
rect 3305 9982 3308 9986
rect 3312 9982 3315 9986
rect 3319 9982 3322 9986
rect 3326 9982 3329 9986
rect 3333 9982 3336 9986
rect 3340 9982 3343 9986
rect 3347 9982 3350 9986
rect 3354 9982 3357 9986
rect 3361 9982 3364 9986
rect 3368 9982 3371 9986
rect 3375 9982 3378 9986
rect 3382 9982 3385 9986
rect 3389 9982 3392 9986
rect 3396 9982 3401 9986
rect 3305 9953 3401 9982
rect 3614 9992 3617 9993
rect 3621 9992 3624 9996
rect 3628 9992 3631 9996
rect 3635 9992 3638 9996
rect 3642 9992 3645 9996
rect 3649 9992 3652 9996
rect 3656 9992 3659 9996
rect 3663 9992 3666 9996
rect 3670 9992 3673 9996
rect 3677 9992 3680 9996
rect 3684 9992 3687 9996
rect 3691 9992 3694 9996
rect 3698 9992 3701 9996
rect 3705 9993 3720 9996
rect 3913 10001 4029 10002
rect 3913 9997 3926 10001
rect 3930 9997 3933 10001
rect 3937 9997 3940 10001
rect 3944 9997 3947 10001
rect 3951 9997 3954 10001
rect 3958 9997 3961 10001
rect 3965 9997 3968 10001
rect 3972 9997 3975 10001
rect 3979 9997 3982 10001
rect 3986 9997 3989 10001
rect 3993 9997 3996 10001
rect 4000 9997 4003 10001
rect 4007 9997 4010 10001
rect 4014 9997 4029 10001
rect 3913 9996 4029 9997
rect 3913 9993 3926 9996
rect 3705 9992 3710 9993
rect 3614 9991 3710 9992
rect 3614 9987 3617 9991
rect 3621 9987 3624 9991
rect 3628 9987 3631 9991
rect 3635 9987 3638 9991
rect 3642 9987 3645 9991
rect 3649 9987 3652 9991
rect 3656 9987 3659 9991
rect 3663 9987 3666 9991
rect 3670 9987 3673 9991
rect 3677 9987 3680 9991
rect 3684 9987 3687 9991
rect 3691 9987 3694 9991
rect 3698 9987 3701 9991
rect 3705 9987 3710 9991
rect 3614 9986 3710 9987
rect 3614 9982 3617 9986
rect 3621 9982 3624 9986
rect 3628 9982 3631 9986
rect 3635 9982 3638 9986
rect 3642 9982 3645 9986
rect 3649 9982 3652 9986
rect 3656 9982 3659 9986
rect 3663 9982 3666 9986
rect 3670 9982 3673 9986
rect 3677 9982 3680 9986
rect 3684 9982 3687 9986
rect 3691 9982 3694 9986
rect 3698 9982 3701 9986
rect 3705 9982 3710 9986
rect 3614 9953 3710 9982
rect 3923 9992 3926 9993
rect 3930 9992 3933 9996
rect 3937 9992 3940 9996
rect 3944 9992 3947 9996
rect 3951 9992 3954 9996
rect 3958 9992 3961 9996
rect 3965 9992 3968 9996
rect 3972 9992 3975 9996
rect 3979 9992 3982 9996
rect 3986 9992 3989 9996
rect 3993 9992 3996 9996
rect 4000 9992 4003 9996
rect 4007 9992 4010 9996
rect 4014 9993 4029 9996
rect 4014 9992 4019 9993
rect 3923 9991 4019 9992
rect 3923 9987 3926 9991
rect 3930 9987 3933 9991
rect 3937 9987 3940 9991
rect 3944 9987 3947 9991
rect 3951 9987 3954 9991
rect 3958 9987 3961 9991
rect 3965 9987 3968 9991
rect 3972 9987 3975 9991
rect 3979 9987 3982 9991
rect 3986 9987 3989 9991
rect 3993 9987 3996 9991
rect 4000 9987 4003 9991
rect 4007 9987 4010 9991
rect 4014 9987 4019 9991
rect 3923 9986 4019 9987
rect 3923 9982 3926 9986
rect 3930 9982 3933 9986
rect 3937 9982 3940 9986
rect 3944 9982 3947 9986
rect 3951 9982 3954 9986
rect 3958 9982 3961 9986
rect 3965 9982 3968 9986
rect 3972 9982 3975 9986
rect 3979 9982 3982 9986
rect 3986 9982 3989 9986
rect 3993 9982 3996 9986
rect 4000 9982 4003 9986
rect 4007 9982 4010 9986
rect 4014 9982 4019 9986
rect 3923 9953 4019 9982
rect 1401 9949 1407 9953
rect 1411 9949 1417 9953
rect 1421 9949 1427 9953
rect 1431 9949 1437 9953
rect 1441 9949 1557 9953
rect 1561 9949 1567 9953
rect 1571 9949 1577 9953
rect 1581 9949 1587 9953
rect 1591 9949 1597 9953
rect 1397 9948 1601 9949
rect 1397 9944 1402 9948
rect 1406 9944 1412 9948
rect 1416 9944 1422 9948
rect 1426 9944 1432 9948
rect 1436 9944 1562 9948
rect 1566 9944 1572 9948
rect 1576 9944 1582 9948
rect 1586 9944 1592 9948
rect 1596 9944 1601 9948
rect 1397 9943 1601 9944
rect 1401 9939 1407 9943
rect 1411 9939 1417 9943
rect 1421 9939 1427 9943
rect 1431 9939 1437 9943
rect 1441 9939 1557 9943
rect 1561 9939 1567 9943
rect 1571 9939 1577 9943
rect 1581 9939 1587 9943
rect 1591 9939 1597 9943
rect 1397 9938 1601 9939
rect 1397 9934 1402 9938
rect 1406 9934 1412 9938
rect 1416 9934 1422 9938
rect 1426 9934 1432 9938
rect 1436 9934 1562 9938
rect 1566 9934 1572 9938
rect 1576 9934 1582 9938
rect 1586 9934 1592 9938
rect 1596 9934 1601 9938
rect 1397 9933 1601 9934
rect 1401 9929 1407 9933
rect 1411 9929 1417 9933
rect 1421 9929 1427 9933
rect 1431 9929 1437 9933
rect 1441 9929 1557 9933
rect 1561 9929 1567 9933
rect 1571 9929 1577 9933
rect 1581 9929 1587 9933
rect 1591 9929 1597 9933
rect 1397 9928 1601 9929
rect 1397 9924 1402 9928
rect 1406 9924 1412 9928
rect 1416 9924 1422 9928
rect 1426 9924 1432 9928
rect 1436 9924 1562 9928
rect 1566 9924 1572 9928
rect 1576 9924 1582 9928
rect 1586 9924 1592 9928
rect 1596 9924 1601 9928
rect 1397 9923 1601 9924
rect 1401 9919 1407 9923
rect 1411 9919 1417 9923
rect 1421 9919 1427 9923
rect 1431 9919 1437 9923
rect 1441 9919 1557 9923
rect 1561 9919 1567 9923
rect 1571 9919 1577 9923
rect 1581 9919 1587 9923
rect 1591 9919 1597 9923
rect 1397 9918 1601 9919
rect 1397 9914 1402 9918
rect 1406 9914 1412 9918
rect 1416 9914 1422 9918
rect 1426 9914 1432 9918
rect 1436 9914 1562 9918
rect 1566 9914 1572 9918
rect 1576 9914 1582 9918
rect 1586 9914 1592 9918
rect 1596 9914 1601 9918
rect 1397 9913 1601 9914
rect 1401 9909 1407 9913
rect 1411 9909 1417 9913
rect 1421 9909 1427 9913
rect 1431 9909 1437 9913
rect 1441 9909 1557 9913
rect 1561 9909 1567 9913
rect 1571 9909 1577 9913
rect 1581 9909 1587 9913
rect 1591 9909 1597 9913
rect 1397 9908 1601 9909
rect 1397 9904 1402 9908
rect 1406 9904 1412 9908
rect 1416 9904 1422 9908
rect 1426 9904 1432 9908
rect 1436 9904 1562 9908
rect 1566 9904 1572 9908
rect 1576 9904 1582 9908
rect 1586 9904 1592 9908
rect 1596 9904 1601 9908
rect 1397 9903 1601 9904
rect 1401 9899 1407 9903
rect 1411 9899 1417 9903
rect 1421 9899 1427 9903
rect 1431 9899 1437 9903
rect 1441 9899 1557 9903
rect 1561 9899 1567 9903
rect 1571 9899 1577 9903
rect 1581 9899 1587 9903
rect 1591 9899 1597 9903
rect 1397 9898 1601 9899
rect 1397 9894 1402 9898
rect 1406 9894 1412 9898
rect 1416 9894 1422 9898
rect 1426 9894 1432 9898
rect 1436 9894 1562 9898
rect 1566 9894 1572 9898
rect 1576 9894 1582 9898
rect 1586 9894 1592 9898
rect 1596 9894 1601 9898
rect 1397 9893 1601 9894
rect 1401 9889 1407 9893
rect 1411 9889 1417 9893
rect 1421 9889 1427 9893
rect 1431 9889 1437 9893
rect 1441 9889 1557 9893
rect 1561 9889 1567 9893
rect 1571 9889 1577 9893
rect 1581 9889 1587 9893
rect 1591 9889 1597 9893
rect 1397 9888 1601 9889
rect 1397 9884 1402 9888
rect 1406 9884 1412 9888
rect 1416 9884 1422 9888
rect 1426 9884 1432 9888
rect 1436 9884 1562 9888
rect 1566 9884 1572 9888
rect 1576 9884 1582 9888
rect 1586 9884 1592 9888
rect 1596 9884 1601 9888
rect 1397 9883 1601 9884
rect 1401 9879 1407 9883
rect 1411 9879 1417 9883
rect 1421 9879 1427 9883
rect 1431 9879 1437 9883
rect 1441 9879 1557 9883
rect 1561 9879 1567 9883
rect 1571 9879 1577 9883
rect 1581 9879 1587 9883
rect 1591 9879 1597 9883
rect 1397 9878 1601 9879
rect 1397 9874 1402 9878
rect 1406 9874 1412 9878
rect 1416 9874 1422 9878
rect 1426 9874 1432 9878
rect 1436 9874 1562 9878
rect 1566 9874 1572 9878
rect 1576 9874 1582 9878
rect 1586 9874 1592 9878
rect 1596 9874 1601 9878
rect 1397 9873 1601 9874
rect 1401 9869 1407 9873
rect 1411 9869 1417 9873
rect 1421 9869 1427 9873
rect 1431 9869 1437 9873
rect 1441 9869 1557 9873
rect 1561 9869 1567 9873
rect 1571 9869 1577 9873
rect 1581 9869 1587 9873
rect 1591 9869 1597 9873
rect 1397 9868 1601 9869
rect 1397 9864 1402 9868
rect 1406 9864 1412 9868
rect 1416 9864 1422 9868
rect 1426 9864 1432 9868
rect 1436 9864 1562 9868
rect 1566 9864 1572 9868
rect 1576 9864 1582 9868
rect 1586 9864 1592 9868
rect 1596 9864 1601 9868
rect 1710 9949 1716 9953
rect 1720 9949 1726 9953
rect 1730 9949 1736 9953
rect 1740 9949 1746 9953
rect 1750 9949 1866 9953
rect 1870 9949 1876 9953
rect 1880 9949 1886 9953
rect 1890 9949 1896 9953
rect 1900 9949 1906 9953
rect 1706 9948 1910 9949
rect 1706 9944 1711 9948
rect 1715 9944 1721 9948
rect 1725 9944 1731 9948
rect 1735 9944 1741 9948
rect 1745 9944 1871 9948
rect 1875 9944 1881 9948
rect 1885 9944 1891 9948
rect 1895 9944 1901 9948
rect 1905 9944 1910 9948
rect 1706 9943 1910 9944
rect 1710 9939 1716 9943
rect 1720 9939 1726 9943
rect 1730 9939 1736 9943
rect 1740 9939 1746 9943
rect 1750 9939 1866 9943
rect 1870 9939 1876 9943
rect 1880 9939 1886 9943
rect 1890 9939 1896 9943
rect 1900 9939 1906 9943
rect 1706 9938 1910 9939
rect 1706 9934 1711 9938
rect 1715 9934 1721 9938
rect 1725 9934 1731 9938
rect 1735 9934 1741 9938
rect 1745 9934 1871 9938
rect 1875 9934 1881 9938
rect 1885 9934 1891 9938
rect 1895 9934 1901 9938
rect 1905 9934 1910 9938
rect 1706 9933 1910 9934
rect 1710 9929 1716 9933
rect 1720 9929 1726 9933
rect 1730 9929 1736 9933
rect 1740 9929 1746 9933
rect 1750 9929 1866 9933
rect 1870 9929 1876 9933
rect 1880 9929 1886 9933
rect 1890 9929 1896 9933
rect 1900 9929 1906 9933
rect 1706 9928 1910 9929
rect 1706 9924 1711 9928
rect 1715 9924 1721 9928
rect 1725 9924 1731 9928
rect 1735 9924 1741 9928
rect 1745 9924 1871 9928
rect 1875 9924 1881 9928
rect 1885 9924 1891 9928
rect 1895 9924 1901 9928
rect 1905 9924 1910 9928
rect 1706 9923 1910 9924
rect 1710 9919 1716 9923
rect 1720 9919 1726 9923
rect 1730 9919 1736 9923
rect 1740 9919 1746 9923
rect 1750 9919 1866 9923
rect 1870 9919 1876 9923
rect 1880 9919 1886 9923
rect 1890 9919 1896 9923
rect 1900 9919 1906 9923
rect 1706 9918 1910 9919
rect 1706 9914 1711 9918
rect 1715 9914 1721 9918
rect 1725 9914 1731 9918
rect 1735 9914 1741 9918
rect 1745 9914 1871 9918
rect 1875 9914 1881 9918
rect 1885 9914 1891 9918
rect 1895 9914 1901 9918
rect 1905 9914 1910 9918
rect 1706 9913 1910 9914
rect 1710 9909 1716 9913
rect 1720 9909 1726 9913
rect 1730 9909 1736 9913
rect 1740 9909 1746 9913
rect 1750 9909 1866 9913
rect 1870 9909 1876 9913
rect 1880 9909 1886 9913
rect 1890 9909 1896 9913
rect 1900 9909 1906 9913
rect 1706 9908 1910 9909
rect 1706 9904 1711 9908
rect 1715 9904 1721 9908
rect 1725 9904 1731 9908
rect 1735 9904 1741 9908
rect 1745 9904 1871 9908
rect 1875 9904 1881 9908
rect 1885 9904 1891 9908
rect 1895 9904 1901 9908
rect 1905 9904 1910 9908
rect 1706 9903 1910 9904
rect 1710 9899 1716 9903
rect 1720 9899 1726 9903
rect 1730 9899 1736 9903
rect 1740 9899 1746 9903
rect 1750 9899 1866 9903
rect 1870 9899 1876 9903
rect 1880 9899 1886 9903
rect 1890 9899 1896 9903
rect 1900 9899 1906 9903
rect 1706 9898 1910 9899
rect 1706 9894 1711 9898
rect 1715 9894 1721 9898
rect 1725 9894 1731 9898
rect 1735 9894 1741 9898
rect 1745 9894 1871 9898
rect 1875 9894 1881 9898
rect 1885 9894 1891 9898
rect 1895 9894 1901 9898
rect 1905 9894 1910 9898
rect 1706 9893 1910 9894
rect 1710 9889 1716 9893
rect 1720 9889 1726 9893
rect 1730 9889 1736 9893
rect 1740 9889 1746 9893
rect 1750 9889 1866 9893
rect 1870 9889 1876 9893
rect 1880 9889 1886 9893
rect 1890 9889 1896 9893
rect 1900 9889 1906 9893
rect 1706 9888 1910 9889
rect 1706 9884 1711 9888
rect 1715 9884 1721 9888
rect 1725 9884 1731 9888
rect 1735 9884 1741 9888
rect 1745 9884 1871 9888
rect 1875 9884 1881 9888
rect 1885 9884 1891 9888
rect 1895 9884 1901 9888
rect 1905 9884 1910 9888
rect 1706 9883 1910 9884
rect 1710 9879 1716 9883
rect 1720 9879 1726 9883
rect 1730 9879 1736 9883
rect 1740 9879 1746 9883
rect 1750 9879 1866 9883
rect 1870 9879 1876 9883
rect 1880 9879 1886 9883
rect 1890 9879 1896 9883
rect 1900 9879 1906 9883
rect 1706 9878 1910 9879
rect 1706 9874 1711 9878
rect 1715 9874 1721 9878
rect 1725 9874 1731 9878
rect 1735 9874 1741 9878
rect 1745 9874 1871 9878
rect 1875 9874 1881 9878
rect 1885 9874 1891 9878
rect 1895 9874 1901 9878
rect 1905 9874 1910 9878
rect 1706 9873 1910 9874
rect 1710 9869 1716 9873
rect 1720 9869 1726 9873
rect 1730 9869 1736 9873
rect 1740 9869 1746 9873
rect 1750 9869 1866 9873
rect 1870 9869 1876 9873
rect 1880 9869 1886 9873
rect 1890 9869 1896 9873
rect 1900 9869 1906 9873
rect 1706 9868 1910 9869
rect 1706 9864 1711 9868
rect 1715 9864 1721 9868
rect 1725 9864 1731 9868
rect 1735 9864 1741 9868
rect 1745 9864 1871 9868
rect 1875 9864 1881 9868
rect 1885 9864 1891 9868
rect 1895 9864 1901 9868
rect 1905 9864 1910 9868
rect 2019 9949 2025 9953
rect 2029 9949 2035 9953
rect 2039 9949 2045 9953
rect 2049 9949 2055 9953
rect 2059 9949 2175 9953
rect 2179 9949 2185 9953
rect 2189 9949 2195 9953
rect 2199 9949 2205 9953
rect 2209 9949 2215 9953
rect 2015 9948 2219 9949
rect 2015 9944 2020 9948
rect 2024 9944 2030 9948
rect 2034 9944 2040 9948
rect 2044 9944 2050 9948
rect 2054 9944 2180 9948
rect 2184 9944 2190 9948
rect 2194 9944 2200 9948
rect 2204 9944 2210 9948
rect 2214 9944 2219 9948
rect 2015 9943 2219 9944
rect 2019 9939 2025 9943
rect 2029 9939 2035 9943
rect 2039 9939 2045 9943
rect 2049 9939 2055 9943
rect 2059 9939 2175 9943
rect 2179 9939 2185 9943
rect 2189 9939 2195 9943
rect 2199 9939 2205 9943
rect 2209 9939 2215 9943
rect 2015 9938 2219 9939
rect 2015 9934 2020 9938
rect 2024 9934 2030 9938
rect 2034 9934 2040 9938
rect 2044 9934 2050 9938
rect 2054 9934 2180 9938
rect 2184 9934 2190 9938
rect 2194 9934 2200 9938
rect 2204 9934 2210 9938
rect 2214 9934 2219 9938
rect 2015 9933 2219 9934
rect 2019 9929 2025 9933
rect 2029 9929 2035 9933
rect 2039 9929 2045 9933
rect 2049 9929 2055 9933
rect 2059 9929 2175 9933
rect 2179 9929 2185 9933
rect 2189 9929 2195 9933
rect 2199 9929 2205 9933
rect 2209 9929 2215 9933
rect 2015 9928 2219 9929
rect 2015 9924 2020 9928
rect 2024 9924 2030 9928
rect 2034 9924 2040 9928
rect 2044 9924 2050 9928
rect 2054 9924 2180 9928
rect 2184 9924 2190 9928
rect 2194 9924 2200 9928
rect 2204 9924 2210 9928
rect 2214 9924 2219 9928
rect 2015 9923 2219 9924
rect 2019 9919 2025 9923
rect 2029 9919 2035 9923
rect 2039 9919 2045 9923
rect 2049 9919 2055 9923
rect 2059 9919 2175 9923
rect 2179 9919 2185 9923
rect 2189 9919 2195 9923
rect 2199 9919 2205 9923
rect 2209 9919 2215 9923
rect 2015 9918 2219 9919
rect 2015 9914 2020 9918
rect 2024 9914 2030 9918
rect 2034 9914 2040 9918
rect 2044 9914 2050 9918
rect 2054 9914 2180 9918
rect 2184 9914 2190 9918
rect 2194 9914 2200 9918
rect 2204 9914 2210 9918
rect 2214 9914 2219 9918
rect 2015 9913 2219 9914
rect 2019 9909 2025 9913
rect 2029 9909 2035 9913
rect 2039 9909 2045 9913
rect 2049 9909 2055 9913
rect 2059 9909 2175 9913
rect 2179 9909 2185 9913
rect 2189 9909 2195 9913
rect 2199 9909 2205 9913
rect 2209 9909 2215 9913
rect 2015 9908 2219 9909
rect 2015 9904 2020 9908
rect 2024 9904 2030 9908
rect 2034 9904 2040 9908
rect 2044 9904 2050 9908
rect 2054 9904 2180 9908
rect 2184 9904 2190 9908
rect 2194 9904 2200 9908
rect 2204 9904 2210 9908
rect 2214 9904 2219 9908
rect 2015 9903 2219 9904
rect 2019 9899 2025 9903
rect 2029 9899 2035 9903
rect 2039 9899 2045 9903
rect 2049 9899 2055 9903
rect 2059 9899 2175 9903
rect 2179 9899 2185 9903
rect 2189 9899 2195 9903
rect 2199 9899 2205 9903
rect 2209 9899 2215 9903
rect 2015 9898 2219 9899
rect 2015 9894 2020 9898
rect 2024 9894 2030 9898
rect 2034 9894 2040 9898
rect 2044 9894 2050 9898
rect 2054 9894 2180 9898
rect 2184 9894 2190 9898
rect 2194 9894 2200 9898
rect 2204 9894 2210 9898
rect 2214 9894 2219 9898
rect 2015 9893 2219 9894
rect 2019 9889 2025 9893
rect 2029 9889 2035 9893
rect 2039 9889 2045 9893
rect 2049 9889 2055 9893
rect 2059 9889 2175 9893
rect 2179 9889 2185 9893
rect 2189 9889 2195 9893
rect 2199 9889 2205 9893
rect 2209 9889 2215 9893
rect 2015 9888 2219 9889
rect 2015 9884 2020 9888
rect 2024 9884 2030 9888
rect 2034 9884 2040 9888
rect 2044 9884 2050 9888
rect 2054 9884 2180 9888
rect 2184 9884 2190 9888
rect 2194 9884 2200 9888
rect 2204 9884 2210 9888
rect 2214 9884 2219 9888
rect 2015 9883 2219 9884
rect 2019 9879 2025 9883
rect 2029 9879 2035 9883
rect 2039 9879 2045 9883
rect 2049 9879 2055 9883
rect 2059 9879 2175 9883
rect 2179 9879 2185 9883
rect 2189 9879 2195 9883
rect 2199 9879 2205 9883
rect 2209 9879 2215 9883
rect 2015 9878 2219 9879
rect 2015 9874 2020 9878
rect 2024 9874 2030 9878
rect 2034 9874 2040 9878
rect 2044 9874 2050 9878
rect 2054 9874 2180 9878
rect 2184 9874 2190 9878
rect 2194 9874 2200 9878
rect 2204 9874 2210 9878
rect 2214 9874 2219 9878
rect 2015 9873 2219 9874
rect 2019 9869 2025 9873
rect 2029 9869 2035 9873
rect 2039 9869 2045 9873
rect 2049 9869 2055 9873
rect 2059 9869 2175 9873
rect 2179 9869 2185 9873
rect 2189 9869 2195 9873
rect 2199 9869 2205 9873
rect 2209 9869 2215 9873
rect 2015 9868 2219 9869
rect 2015 9864 2020 9868
rect 2024 9864 2030 9868
rect 2034 9864 2040 9868
rect 2044 9864 2050 9868
rect 2054 9864 2180 9868
rect 2184 9864 2190 9868
rect 2194 9864 2200 9868
rect 2204 9864 2210 9868
rect 2214 9864 2219 9868
rect 2328 9949 2334 9953
rect 2338 9949 2344 9953
rect 2348 9949 2354 9953
rect 2358 9949 2364 9953
rect 2368 9949 2484 9953
rect 2488 9949 2494 9953
rect 2498 9949 2504 9953
rect 2508 9949 2514 9953
rect 2518 9949 2524 9953
rect 2324 9948 2528 9949
rect 2324 9944 2329 9948
rect 2333 9944 2339 9948
rect 2343 9944 2349 9948
rect 2353 9944 2359 9948
rect 2363 9944 2489 9948
rect 2493 9944 2499 9948
rect 2503 9944 2509 9948
rect 2513 9944 2519 9948
rect 2523 9944 2528 9948
rect 2324 9943 2528 9944
rect 2328 9939 2334 9943
rect 2338 9939 2344 9943
rect 2348 9939 2354 9943
rect 2358 9939 2364 9943
rect 2368 9939 2484 9943
rect 2488 9939 2494 9943
rect 2498 9939 2504 9943
rect 2508 9939 2514 9943
rect 2518 9939 2524 9943
rect 2324 9938 2528 9939
rect 2324 9934 2329 9938
rect 2333 9934 2339 9938
rect 2343 9934 2349 9938
rect 2353 9934 2359 9938
rect 2363 9934 2489 9938
rect 2493 9934 2499 9938
rect 2503 9934 2509 9938
rect 2513 9934 2519 9938
rect 2523 9934 2528 9938
rect 2324 9933 2528 9934
rect 2328 9929 2334 9933
rect 2338 9929 2344 9933
rect 2348 9929 2354 9933
rect 2358 9929 2364 9933
rect 2368 9929 2484 9933
rect 2488 9929 2494 9933
rect 2498 9929 2504 9933
rect 2508 9929 2514 9933
rect 2518 9929 2524 9933
rect 2324 9928 2528 9929
rect 2324 9924 2329 9928
rect 2333 9924 2339 9928
rect 2343 9924 2349 9928
rect 2353 9924 2359 9928
rect 2363 9924 2489 9928
rect 2493 9924 2499 9928
rect 2503 9924 2509 9928
rect 2513 9924 2519 9928
rect 2523 9924 2528 9928
rect 2324 9923 2528 9924
rect 2328 9919 2334 9923
rect 2338 9919 2344 9923
rect 2348 9919 2354 9923
rect 2358 9919 2364 9923
rect 2368 9919 2484 9923
rect 2488 9919 2494 9923
rect 2498 9919 2504 9923
rect 2508 9919 2514 9923
rect 2518 9919 2524 9923
rect 2324 9918 2528 9919
rect 2324 9914 2329 9918
rect 2333 9914 2339 9918
rect 2343 9914 2349 9918
rect 2353 9914 2359 9918
rect 2363 9914 2489 9918
rect 2493 9914 2499 9918
rect 2503 9914 2509 9918
rect 2513 9914 2519 9918
rect 2523 9914 2528 9918
rect 2324 9913 2528 9914
rect 2328 9909 2334 9913
rect 2338 9909 2344 9913
rect 2348 9909 2354 9913
rect 2358 9909 2364 9913
rect 2368 9909 2484 9913
rect 2488 9909 2494 9913
rect 2498 9909 2504 9913
rect 2508 9909 2514 9913
rect 2518 9909 2524 9913
rect 2324 9908 2528 9909
rect 2324 9904 2329 9908
rect 2333 9904 2339 9908
rect 2343 9904 2349 9908
rect 2353 9904 2359 9908
rect 2363 9904 2489 9908
rect 2493 9904 2499 9908
rect 2503 9904 2509 9908
rect 2513 9904 2519 9908
rect 2523 9904 2528 9908
rect 2324 9903 2528 9904
rect 2328 9899 2334 9903
rect 2338 9899 2344 9903
rect 2348 9899 2354 9903
rect 2358 9899 2364 9903
rect 2368 9899 2484 9903
rect 2488 9899 2494 9903
rect 2498 9899 2504 9903
rect 2508 9899 2514 9903
rect 2518 9899 2524 9903
rect 2324 9898 2528 9899
rect 2324 9894 2329 9898
rect 2333 9894 2339 9898
rect 2343 9894 2349 9898
rect 2353 9894 2359 9898
rect 2363 9894 2489 9898
rect 2493 9894 2499 9898
rect 2503 9894 2509 9898
rect 2513 9894 2519 9898
rect 2523 9894 2528 9898
rect 2324 9893 2528 9894
rect 2328 9889 2334 9893
rect 2338 9889 2344 9893
rect 2348 9889 2354 9893
rect 2358 9889 2364 9893
rect 2368 9889 2484 9893
rect 2488 9889 2494 9893
rect 2498 9889 2504 9893
rect 2508 9889 2514 9893
rect 2518 9889 2524 9893
rect 2324 9888 2528 9889
rect 2324 9884 2329 9888
rect 2333 9884 2339 9888
rect 2343 9884 2349 9888
rect 2353 9884 2359 9888
rect 2363 9884 2489 9888
rect 2493 9884 2499 9888
rect 2503 9884 2509 9888
rect 2513 9884 2519 9888
rect 2523 9884 2528 9888
rect 2324 9883 2528 9884
rect 2328 9879 2334 9883
rect 2338 9879 2344 9883
rect 2348 9879 2354 9883
rect 2358 9879 2364 9883
rect 2368 9879 2484 9883
rect 2488 9879 2494 9883
rect 2498 9879 2504 9883
rect 2508 9879 2514 9883
rect 2518 9879 2524 9883
rect 2324 9878 2528 9879
rect 2324 9874 2329 9878
rect 2333 9874 2339 9878
rect 2343 9874 2349 9878
rect 2353 9874 2359 9878
rect 2363 9874 2489 9878
rect 2493 9874 2499 9878
rect 2503 9874 2509 9878
rect 2513 9874 2519 9878
rect 2523 9874 2528 9878
rect 2324 9873 2528 9874
rect 2328 9869 2334 9873
rect 2338 9869 2344 9873
rect 2348 9869 2354 9873
rect 2358 9869 2364 9873
rect 2368 9869 2484 9873
rect 2488 9869 2494 9873
rect 2498 9869 2504 9873
rect 2508 9869 2514 9873
rect 2518 9869 2524 9873
rect 2324 9868 2528 9869
rect 2324 9864 2329 9868
rect 2333 9864 2339 9868
rect 2343 9864 2349 9868
rect 2353 9864 2359 9868
rect 2363 9864 2489 9868
rect 2493 9864 2499 9868
rect 2503 9864 2509 9868
rect 2513 9864 2519 9868
rect 2523 9864 2528 9868
rect 2637 9949 2643 9953
rect 2647 9949 2653 9953
rect 2657 9949 2663 9953
rect 2667 9949 2673 9953
rect 2677 9949 2793 9953
rect 2797 9949 2803 9953
rect 2807 9949 2813 9953
rect 2817 9949 2823 9953
rect 2827 9949 2833 9953
rect 2633 9948 2837 9949
rect 2633 9944 2638 9948
rect 2642 9944 2648 9948
rect 2652 9944 2658 9948
rect 2662 9944 2668 9948
rect 2672 9944 2798 9948
rect 2802 9944 2808 9948
rect 2812 9944 2818 9948
rect 2822 9944 2828 9948
rect 2832 9944 2837 9948
rect 2633 9943 2837 9944
rect 2637 9939 2643 9943
rect 2647 9939 2653 9943
rect 2657 9939 2663 9943
rect 2667 9939 2673 9943
rect 2677 9939 2793 9943
rect 2797 9939 2803 9943
rect 2807 9939 2813 9943
rect 2817 9939 2823 9943
rect 2827 9939 2833 9943
rect 2633 9938 2837 9939
rect 2633 9934 2638 9938
rect 2642 9934 2648 9938
rect 2652 9934 2658 9938
rect 2662 9934 2668 9938
rect 2672 9934 2798 9938
rect 2802 9934 2808 9938
rect 2812 9934 2818 9938
rect 2822 9934 2828 9938
rect 2832 9934 2837 9938
rect 2633 9933 2837 9934
rect 2637 9929 2643 9933
rect 2647 9929 2653 9933
rect 2657 9929 2663 9933
rect 2667 9929 2673 9933
rect 2677 9929 2793 9933
rect 2797 9929 2803 9933
rect 2807 9929 2813 9933
rect 2817 9929 2823 9933
rect 2827 9929 2833 9933
rect 2633 9928 2837 9929
rect 2633 9924 2638 9928
rect 2642 9924 2648 9928
rect 2652 9924 2658 9928
rect 2662 9924 2668 9928
rect 2672 9924 2798 9928
rect 2802 9924 2808 9928
rect 2812 9924 2818 9928
rect 2822 9924 2828 9928
rect 2832 9924 2837 9928
rect 2633 9923 2837 9924
rect 2637 9919 2643 9923
rect 2647 9919 2653 9923
rect 2657 9919 2663 9923
rect 2667 9919 2673 9923
rect 2677 9919 2793 9923
rect 2797 9919 2803 9923
rect 2807 9919 2813 9923
rect 2817 9919 2823 9923
rect 2827 9919 2833 9923
rect 2633 9918 2837 9919
rect 2633 9914 2638 9918
rect 2642 9914 2648 9918
rect 2652 9914 2658 9918
rect 2662 9914 2668 9918
rect 2672 9914 2798 9918
rect 2802 9914 2808 9918
rect 2812 9914 2818 9918
rect 2822 9914 2828 9918
rect 2832 9914 2837 9918
rect 2633 9913 2837 9914
rect 2637 9909 2643 9913
rect 2647 9909 2653 9913
rect 2657 9909 2663 9913
rect 2667 9909 2673 9913
rect 2677 9909 2793 9913
rect 2797 9909 2803 9913
rect 2807 9909 2813 9913
rect 2817 9909 2823 9913
rect 2827 9909 2833 9913
rect 2633 9908 2837 9909
rect 2633 9904 2638 9908
rect 2642 9904 2648 9908
rect 2652 9904 2658 9908
rect 2662 9904 2668 9908
rect 2672 9904 2798 9908
rect 2802 9904 2808 9908
rect 2812 9904 2818 9908
rect 2822 9904 2828 9908
rect 2832 9904 2837 9908
rect 2633 9903 2837 9904
rect 2637 9899 2643 9903
rect 2647 9899 2653 9903
rect 2657 9899 2663 9903
rect 2667 9899 2673 9903
rect 2677 9899 2793 9903
rect 2797 9899 2803 9903
rect 2807 9899 2813 9903
rect 2817 9899 2823 9903
rect 2827 9899 2833 9903
rect 2633 9898 2837 9899
rect 2633 9894 2638 9898
rect 2642 9894 2648 9898
rect 2652 9894 2658 9898
rect 2662 9894 2668 9898
rect 2672 9894 2798 9898
rect 2802 9894 2808 9898
rect 2812 9894 2818 9898
rect 2822 9894 2828 9898
rect 2832 9894 2837 9898
rect 2633 9893 2837 9894
rect 2637 9889 2643 9893
rect 2647 9889 2653 9893
rect 2657 9889 2663 9893
rect 2667 9889 2673 9893
rect 2677 9889 2793 9893
rect 2797 9889 2803 9893
rect 2807 9889 2813 9893
rect 2817 9889 2823 9893
rect 2827 9889 2833 9893
rect 2633 9888 2837 9889
rect 2633 9884 2638 9888
rect 2642 9884 2648 9888
rect 2652 9884 2658 9888
rect 2662 9884 2668 9888
rect 2672 9884 2798 9888
rect 2802 9884 2808 9888
rect 2812 9884 2818 9888
rect 2822 9884 2828 9888
rect 2832 9884 2837 9888
rect 2633 9883 2837 9884
rect 2637 9879 2643 9883
rect 2647 9879 2653 9883
rect 2657 9879 2663 9883
rect 2667 9879 2673 9883
rect 2677 9879 2793 9883
rect 2797 9879 2803 9883
rect 2807 9879 2813 9883
rect 2817 9879 2823 9883
rect 2827 9879 2833 9883
rect 2633 9878 2837 9879
rect 2633 9874 2638 9878
rect 2642 9874 2648 9878
rect 2652 9874 2658 9878
rect 2662 9874 2668 9878
rect 2672 9874 2798 9878
rect 2802 9874 2808 9878
rect 2812 9874 2818 9878
rect 2822 9874 2828 9878
rect 2832 9874 2837 9878
rect 2633 9873 2837 9874
rect 2637 9869 2643 9873
rect 2647 9869 2653 9873
rect 2657 9869 2663 9873
rect 2667 9869 2673 9873
rect 2677 9869 2793 9873
rect 2797 9869 2803 9873
rect 2807 9869 2813 9873
rect 2817 9869 2823 9873
rect 2827 9869 2833 9873
rect 2633 9868 2837 9869
rect 2633 9864 2638 9868
rect 2642 9864 2648 9868
rect 2652 9864 2658 9868
rect 2662 9864 2668 9868
rect 2672 9864 2798 9868
rect 2802 9864 2808 9868
rect 2812 9864 2818 9868
rect 2822 9864 2828 9868
rect 2832 9864 2837 9868
rect 2946 9949 2952 9953
rect 2956 9949 2962 9953
rect 2966 9949 2972 9953
rect 2976 9949 2982 9953
rect 2986 9949 3102 9953
rect 3106 9949 3112 9953
rect 3116 9949 3122 9953
rect 3126 9949 3132 9953
rect 3136 9949 3142 9953
rect 2942 9948 3146 9949
rect 2942 9944 2947 9948
rect 2951 9944 2957 9948
rect 2961 9944 2967 9948
rect 2971 9944 2977 9948
rect 2981 9944 3107 9948
rect 3111 9944 3117 9948
rect 3121 9944 3127 9948
rect 3131 9944 3137 9948
rect 3141 9944 3146 9948
rect 2942 9943 3146 9944
rect 2946 9939 2952 9943
rect 2956 9939 2962 9943
rect 2966 9939 2972 9943
rect 2976 9939 2982 9943
rect 2986 9939 3102 9943
rect 3106 9939 3112 9943
rect 3116 9939 3122 9943
rect 3126 9939 3132 9943
rect 3136 9939 3142 9943
rect 2942 9938 3146 9939
rect 2942 9934 2947 9938
rect 2951 9934 2957 9938
rect 2961 9934 2967 9938
rect 2971 9934 2977 9938
rect 2981 9934 3107 9938
rect 3111 9934 3117 9938
rect 3121 9934 3127 9938
rect 3131 9934 3137 9938
rect 3141 9934 3146 9938
rect 2942 9933 3146 9934
rect 2946 9929 2952 9933
rect 2956 9929 2962 9933
rect 2966 9929 2972 9933
rect 2976 9929 2982 9933
rect 2986 9929 3102 9933
rect 3106 9929 3112 9933
rect 3116 9929 3122 9933
rect 3126 9929 3132 9933
rect 3136 9929 3142 9933
rect 2942 9928 3146 9929
rect 2942 9924 2947 9928
rect 2951 9924 2957 9928
rect 2961 9924 2967 9928
rect 2971 9924 2977 9928
rect 2981 9924 3107 9928
rect 3111 9924 3117 9928
rect 3121 9924 3127 9928
rect 3131 9924 3137 9928
rect 3141 9924 3146 9928
rect 2942 9923 3146 9924
rect 2946 9919 2952 9923
rect 2956 9919 2962 9923
rect 2966 9919 2972 9923
rect 2976 9919 2982 9923
rect 2986 9919 3102 9923
rect 3106 9919 3112 9923
rect 3116 9919 3122 9923
rect 3126 9919 3132 9923
rect 3136 9919 3142 9923
rect 2942 9918 3146 9919
rect 2942 9914 2947 9918
rect 2951 9914 2957 9918
rect 2961 9914 2967 9918
rect 2971 9914 2977 9918
rect 2981 9914 3107 9918
rect 3111 9914 3117 9918
rect 3121 9914 3127 9918
rect 3131 9914 3137 9918
rect 3141 9914 3146 9918
rect 2942 9913 3146 9914
rect 2946 9909 2952 9913
rect 2956 9909 2962 9913
rect 2966 9909 2972 9913
rect 2976 9909 2982 9913
rect 2986 9909 3102 9913
rect 3106 9909 3112 9913
rect 3116 9909 3122 9913
rect 3126 9909 3132 9913
rect 3136 9909 3142 9913
rect 2942 9908 3146 9909
rect 2942 9904 2947 9908
rect 2951 9904 2957 9908
rect 2961 9904 2967 9908
rect 2971 9904 2977 9908
rect 2981 9904 3107 9908
rect 3111 9904 3117 9908
rect 3121 9904 3127 9908
rect 3131 9904 3137 9908
rect 3141 9904 3146 9908
rect 2942 9903 3146 9904
rect 2946 9899 2952 9903
rect 2956 9899 2962 9903
rect 2966 9899 2972 9903
rect 2976 9899 2982 9903
rect 2986 9899 3102 9903
rect 3106 9899 3112 9903
rect 3116 9899 3122 9903
rect 3126 9899 3132 9903
rect 3136 9899 3142 9903
rect 2942 9898 3146 9899
rect 2942 9894 2947 9898
rect 2951 9894 2957 9898
rect 2961 9894 2967 9898
rect 2971 9894 2977 9898
rect 2981 9894 3107 9898
rect 3111 9894 3117 9898
rect 3121 9894 3127 9898
rect 3131 9894 3137 9898
rect 3141 9894 3146 9898
rect 2942 9893 3146 9894
rect 2946 9889 2952 9893
rect 2956 9889 2962 9893
rect 2966 9889 2972 9893
rect 2976 9889 2982 9893
rect 2986 9889 3102 9893
rect 3106 9889 3112 9893
rect 3116 9889 3122 9893
rect 3126 9889 3132 9893
rect 3136 9889 3142 9893
rect 2942 9888 3146 9889
rect 2942 9884 2947 9888
rect 2951 9884 2957 9888
rect 2961 9884 2967 9888
rect 2971 9884 2977 9888
rect 2981 9884 3107 9888
rect 3111 9884 3117 9888
rect 3121 9884 3127 9888
rect 3131 9884 3137 9888
rect 3141 9884 3146 9888
rect 2942 9883 3146 9884
rect 2946 9879 2952 9883
rect 2956 9879 2962 9883
rect 2966 9879 2972 9883
rect 2976 9879 2982 9883
rect 2986 9879 3102 9883
rect 3106 9879 3112 9883
rect 3116 9879 3122 9883
rect 3126 9879 3132 9883
rect 3136 9879 3142 9883
rect 2942 9878 3146 9879
rect 2942 9874 2947 9878
rect 2951 9874 2957 9878
rect 2961 9874 2967 9878
rect 2971 9874 2977 9878
rect 2981 9874 3107 9878
rect 3111 9874 3117 9878
rect 3121 9874 3127 9878
rect 3131 9874 3137 9878
rect 3141 9874 3146 9878
rect 2942 9873 3146 9874
rect 2946 9869 2952 9873
rect 2956 9869 2962 9873
rect 2966 9869 2972 9873
rect 2976 9869 2982 9873
rect 2986 9869 3102 9873
rect 3106 9869 3112 9873
rect 3116 9869 3122 9873
rect 3126 9869 3132 9873
rect 3136 9869 3142 9873
rect 2942 9868 3146 9869
rect 2942 9864 2947 9868
rect 2951 9864 2957 9868
rect 2961 9864 2967 9868
rect 2971 9864 2977 9868
rect 2981 9864 3107 9868
rect 3111 9864 3117 9868
rect 3121 9864 3127 9868
rect 3131 9864 3137 9868
rect 3141 9864 3146 9868
rect 3255 9949 3261 9953
rect 3265 9949 3271 9953
rect 3275 9949 3281 9953
rect 3285 9949 3291 9953
rect 3295 9949 3411 9953
rect 3415 9949 3421 9953
rect 3425 9949 3431 9953
rect 3435 9949 3441 9953
rect 3445 9949 3451 9953
rect 3251 9948 3455 9949
rect 3251 9944 3256 9948
rect 3260 9944 3266 9948
rect 3270 9944 3276 9948
rect 3280 9944 3286 9948
rect 3290 9944 3416 9948
rect 3420 9944 3426 9948
rect 3430 9944 3436 9948
rect 3440 9944 3446 9948
rect 3450 9944 3455 9948
rect 3251 9943 3455 9944
rect 3255 9939 3261 9943
rect 3265 9939 3271 9943
rect 3275 9939 3281 9943
rect 3285 9939 3291 9943
rect 3295 9939 3411 9943
rect 3415 9939 3421 9943
rect 3425 9939 3431 9943
rect 3435 9939 3441 9943
rect 3445 9939 3451 9943
rect 3251 9938 3455 9939
rect 3251 9934 3256 9938
rect 3260 9934 3266 9938
rect 3270 9934 3276 9938
rect 3280 9934 3286 9938
rect 3290 9934 3416 9938
rect 3420 9934 3426 9938
rect 3430 9934 3436 9938
rect 3440 9934 3446 9938
rect 3450 9934 3455 9938
rect 3251 9933 3455 9934
rect 3255 9929 3261 9933
rect 3265 9929 3271 9933
rect 3275 9929 3281 9933
rect 3285 9929 3291 9933
rect 3295 9929 3411 9933
rect 3415 9929 3421 9933
rect 3425 9929 3431 9933
rect 3435 9929 3441 9933
rect 3445 9929 3451 9933
rect 3251 9928 3455 9929
rect 3251 9924 3256 9928
rect 3260 9924 3266 9928
rect 3270 9924 3276 9928
rect 3280 9924 3286 9928
rect 3290 9924 3416 9928
rect 3420 9924 3426 9928
rect 3430 9924 3436 9928
rect 3440 9924 3446 9928
rect 3450 9924 3455 9928
rect 3251 9923 3455 9924
rect 3255 9919 3261 9923
rect 3265 9919 3271 9923
rect 3275 9919 3281 9923
rect 3285 9919 3291 9923
rect 3295 9919 3411 9923
rect 3415 9919 3421 9923
rect 3425 9919 3431 9923
rect 3435 9919 3441 9923
rect 3445 9919 3451 9923
rect 3251 9918 3455 9919
rect 3251 9914 3256 9918
rect 3260 9914 3266 9918
rect 3270 9914 3276 9918
rect 3280 9914 3286 9918
rect 3290 9914 3416 9918
rect 3420 9914 3426 9918
rect 3430 9914 3436 9918
rect 3440 9914 3446 9918
rect 3450 9914 3455 9918
rect 3251 9913 3455 9914
rect 3255 9909 3261 9913
rect 3265 9909 3271 9913
rect 3275 9909 3281 9913
rect 3285 9909 3291 9913
rect 3295 9909 3411 9913
rect 3415 9909 3421 9913
rect 3425 9909 3431 9913
rect 3435 9909 3441 9913
rect 3445 9909 3451 9913
rect 3251 9908 3455 9909
rect 3251 9904 3256 9908
rect 3260 9904 3266 9908
rect 3270 9904 3276 9908
rect 3280 9904 3286 9908
rect 3290 9904 3416 9908
rect 3420 9904 3426 9908
rect 3430 9904 3436 9908
rect 3440 9904 3446 9908
rect 3450 9904 3455 9908
rect 3251 9903 3455 9904
rect 3255 9899 3261 9903
rect 3265 9899 3271 9903
rect 3275 9899 3281 9903
rect 3285 9899 3291 9903
rect 3295 9899 3411 9903
rect 3415 9899 3421 9903
rect 3425 9899 3431 9903
rect 3435 9899 3441 9903
rect 3445 9899 3451 9903
rect 3251 9898 3455 9899
rect 3251 9894 3256 9898
rect 3260 9894 3266 9898
rect 3270 9894 3276 9898
rect 3280 9894 3286 9898
rect 3290 9894 3416 9898
rect 3420 9894 3426 9898
rect 3430 9894 3436 9898
rect 3440 9894 3446 9898
rect 3450 9894 3455 9898
rect 3251 9893 3455 9894
rect 3255 9889 3261 9893
rect 3265 9889 3271 9893
rect 3275 9889 3281 9893
rect 3285 9889 3291 9893
rect 3295 9889 3411 9893
rect 3415 9889 3421 9893
rect 3425 9889 3431 9893
rect 3435 9889 3441 9893
rect 3445 9889 3451 9893
rect 3251 9888 3455 9889
rect 3251 9884 3256 9888
rect 3260 9884 3266 9888
rect 3270 9884 3276 9888
rect 3280 9884 3286 9888
rect 3290 9884 3416 9888
rect 3420 9884 3426 9888
rect 3430 9884 3436 9888
rect 3440 9884 3446 9888
rect 3450 9884 3455 9888
rect 3251 9883 3455 9884
rect 3255 9879 3261 9883
rect 3265 9879 3271 9883
rect 3275 9879 3281 9883
rect 3285 9879 3291 9883
rect 3295 9879 3411 9883
rect 3415 9879 3421 9883
rect 3425 9879 3431 9883
rect 3435 9879 3441 9883
rect 3445 9879 3451 9883
rect 3251 9878 3455 9879
rect 3251 9874 3256 9878
rect 3260 9874 3266 9878
rect 3270 9874 3276 9878
rect 3280 9874 3286 9878
rect 3290 9874 3416 9878
rect 3420 9874 3426 9878
rect 3430 9874 3436 9878
rect 3440 9874 3446 9878
rect 3450 9874 3455 9878
rect 3251 9873 3455 9874
rect 3255 9869 3261 9873
rect 3265 9869 3271 9873
rect 3275 9869 3281 9873
rect 3285 9869 3291 9873
rect 3295 9869 3411 9873
rect 3415 9869 3421 9873
rect 3425 9869 3431 9873
rect 3435 9869 3441 9873
rect 3445 9869 3451 9873
rect 3251 9868 3455 9869
rect 3251 9864 3256 9868
rect 3260 9864 3266 9868
rect 3270 9864 3276 9868
rect 3280 9864 3286 9868
rect 3290 9864 3416 9868
rect 3420 9864 3426 9868
rect 3430 9864 3436 9868
rect 3440 9864 3446 9868
rect 3450 9864 3455 9868
rect 3564 9949 3570 9953
rect 3574 9949 3580 9953
rect 3584 9949 3590 9953
rect 3594 9949 3600 9953
rect 3604 9949 3720 9953
rect 3724 9949 3730 9953
rect 3734 9949 3740 9953
rect 3744 9949 3750 9953
rect 3754 9949 3760 9953
rect 3560 9948 3764 9949
rect 3560 9944 3565 9948
rect 3569 9944 3575 9948
rect 3579 9944 3585 9948
rect 3589 9944 3595 9948
rect 3599 9944 3725 9948
rect 3729 9944 3735 9948
rect 3739 9944 3745 9948
rect 3749 9944 3755 9948
rect 3759 9944 3764 9948
rect 3560 9943 3764 9944
rect 3564 9939 3570 9943
rect 3574 9939 3580 9943
rect 3584 9939 3590 9943
rect 3594 9939 3600 9943
rect 3604 9939 3720 9943
rect 3724 9939 3730 9943
rect 3734 9939 3740 9943
rect 3744 9939 3750 9943
rect 3754 9939 3760 9943
rect 3560 9938 3764 9939
rect 3560 9934 3565 9938
rect 3569 9934 3575 9938
rect 3579 9934 3585 9938
rect 3589 9934 3595 9938
rect 3599 9934 3725 9938
rect 3729 9934 3735 9938
rect 3739 9934 3745 9938
rect 3749 9934 3755 9938
rect 3759 9934 3764 9938
rect 3560 9933 3764 9934
rect 3564 9929 3570 9933
rect 3574 9929 3580 9933
rect 3584 9929 3590 9933
rect 3594 9929 3600 9933
rect 3604 9929 3720 9933
rect 3724 9929 3730 9933
rect 3734 9929 3740 9933
rect 3744 9929 3750 9933
rect 3754 9929 3760 9933
rect 3560 9928 3764 9929
rect 3560 9924 3565 9928
rect 3569 9924 3575 9928
rect 3579 9924 3585 9928
rect 3589 9924 3595 9928
rect 3599 9924 3725 9928
rect 3729 9924 3735 9928
rect 3739 9924 3745 9928
rect 3749 9924 3755 9928
rect 3759 9924 3764 9928
rect 3560 9923 3764 9924
rect 3564 9919 3570 9923
rect 3574 9919 3580 9923
rect 3584 9919 3590 9923
rect 3594 9919 3600 9923
rect 3604 9919 3720 9923
rect 3724 9919 3730 9923
rect 3734 9919 3740 9923
rect 3744 9919 3750 9923
rect 3754 9919 3760 9923
rect 3560 9918 3764 9919
rect 3560 9914 3565 9918
rect 3569 9914 3575 9918
rect 3579 9914 3585 9918
rect 3589 9914 3595 9918
rect 3599 9914 3725 9918
rect 3729 9914 3735 9918
rect 3739 9914 3745 9918
rect 3749 9914 3755 9918
rect 3759 9914 3764 9918
rect 3560 9913 3764 9914
rect 3564 9909 3570 9913
rect 3574 9909 3580 9913
rect 3584 9909 3590 9913
rect 3594 9909 3600 9913
rect 3604 9909 3720 9913
rect 3724 9909 3730 9913
rect 3734 9909 3740 9913
rect 3744 9909 3750 9913
rect 3754 9909 3760 9913
rect 3560 9908 3764 9909
rect 3560 9904 3565 9908
rect 3569 9904 3575 9908
rect 3579 9904 3585 9908
rect 3589 9904 3595 9908
rect 3599 9904 3725 9908
rect 3729 9904 3735 9908
rect 3739 9904 3745 9908
rect 3749 9904 3755 9908
rect 3759 9904 3764 9908
rect 3560 9903 3764 9904
rect 3564 9899 3570 9903
rect 3574 9899 3580 9903
rect 3584 9899 3590 9903
rect 3594 9899 3600 9903
rect 3604 9899 3720 9903
rect 3724 9899 3730 9903
rect 3734 9899 3740 9903
rect 3744 9899 3750 9903
rect 3754 9899 3760 9903
rect 3560 9898 3764 9899
rect 3560 9894 3565 9898
rect 3569 9894 3575 9898
rect 3579 9894 3585 9898
rect 3589 9894 3595 9898
rect 3599 9894 3725 9898
rect 3729 9894 3735 9898
rect 3739 9894 3745 9898
rect 3749 9894 3755 9898
rect 3759 9894 3764 9898
rect 3560 9893 3764 9894
rect 3564 9889 3570 9893
rect 3574 9889 3580 9893
rect 3584 9889 3590 9893
rect 3594 9889 3600 9893
rect 3604 9889 3720 9893
rect 3724 9889 3730 9893
rect 3734 9889 3740 9893
rect 3744 9889 3750 9893
rect 3754 9889 3760 9893
rect 3560 9888 3764 9889
rect 3560 9884 3565 9888
rect 3569 9884 3575 9888
rect 3579 9884 3585 9888
rect 3589 9884 3595 9888
rect 3599 9884 3725 9888
rect 3729 9884 3735 9888
rect 3739 9884 3745 9888
rect 3749 9884 3755 9888
rect 3759 9884 3764 9888
rect 3560 9883 3764 9884
rect 3564 9879 3570 9883
rect 3574 9879 3580 9883
rect 3584 9879 3590 9883
rect 3594 9879 3600 9883
rect 3604 9879 3720 9883
rect 3724 9879 3730 9883
rect 3734 9879 3740 9883
rect 3744 9879 3750 9883
rect 3754 9879 3760 9883
rect 3560 9878 3764 9879
rect 3560 9874 3565 9878
rect 3569 9874 3575 9878
rect 3579 9874 3585 9878
rect 3589 9874 3595 9878
rect 3599 9874 3725 9878
rect 3729 9874 3735 9878
rect 3739 9874 3745 9878
rect 3749 9874 3755 9878
rect 3759 9874 3764 9878
rect 3560 9873 3764 9874
rect 3564 9869 3570 9873
rect 3574 9869 3580 9873
rect 3584 9869 3590 9873
rect 3594 9869 3600 9873
rect 3604 9869 3720 9873
rect 3724 9869 3730 9873
rect 3734 9869 3740 9873
rect 3744 9869 3750 9873
rect 3754 9869 3760 9873
rect 3560 9868 3764 9869
rect 3560 9864 3565 9868
rect 3569 9864 3575 9868
rect 3579 9864 3585 9868
rect 3589 9864 3595 9868
rect 3599 9864 3725 9868
rect 3729 9864 3735 9868
rect 3739 9864 3745 9868
rect 3749 9864 3755 9868
rect 3759 9864 3764 9868
rect 3873 9949 3879 9953
rect 3883 9949 3889 9953
rect 3893 9949 3899 9953
rect 3903 9949 3909 9953
rect 3913 9949 4029 9953
rect 4033 9949 4039 9953
rect 4043 9949 4049 9953
rect 4053 9949 4059 9953
rect 4063 9949 4069 9953
rect 3869 9948 4073 9949
rect 3869 9944 3874 9948
rect 3878 9944 3884 9948
rect 3888 9944 3894 9948
rect 3898 9944 3904 9948
rect 3908 9944 4034 9948
rect 4038 9944 4044 9948
rect 4048 9944 4054 9948
rect 4058 9944 4064 9948
rect 4068 9944 4073 9948
rect 3869 9943 4073 9944
rect 3873 9939 3879 9943
rect 3883 9939 3889 9943
rect 3893 9939 3899 9943
rect 3903 9939 3909 9943
rect 3913 9939 4029 9943
rect 4033 9939 4039 9943
rect 4043 9939 4049 9943
rect 4053 9939 4059 9943
rect 4063 9939 4069 9943
rect 3869 9938 4073 9939
rect 3869 9934 3874 9938
rect 3878 9934 3884 9938
rect 3888 9934 3894 9938
rect 3898 9934 3904 9938
rect 3908 9934 4034 9938
rect 4038 9934 4044 9938
rect 4048 9934 4054 9938
rect 4058 9934 4064 9938
rect 4068 9934 4073 9938
rect 3869 9933 4073 9934
rect 3873 9929 3879 9933
rect 3883 9929 3889 9933
rect 3893 9929 3899 9933
rect 3903 9929 3909 9933
rect 3913 9929 4029 9933
rect 4033 9929 4039 9933
rect 4043 9929 4049 9933
rect 4053 9929 4059 9933
rect 4063 9929 4069 9933
rect 3869 9928 4073 9929
rect 3869 9924 3874 9928
rect 3878 9924 3884 9928
rect 3888 9924 3894 9928
rect 3898 9924 3904 9928
rect 3908 9924 4034 9928
rect 4038 9924 4044 9928
rect 4048 9924 4054 9928
rect 4058 9924 4064 9928
rect 4068 9924 4073 9928
rect 3869 9923 4073 9924
rect 3873 9919 3879 9923
rect 3883 9919 3889 9923
rect 3893 9919 3899 9923
rect 3903 9919 3909 9923
rect 3913 9919 4029 9923
rect 4033 9919 4039 9923
rect 4043 9919 4049 9923
rect 4053 9919 4059 9923
rect 4063 9919 4069 9923
rect 3869 9918 4073 9919
rect 3869 9914 3874 9918
rect 3878 9914 3884 9918
rect 3888 9914 3894 9918
rect 3898 9914 3904 9918
rect 3908 9914 4034 9918
rect 4038 9914 4044 9918
rect 4048 9914 4054 9918
rect 4058 9914 4064 9918
rect 4068 9914 4073 9918
rect 3869 9913 4073 9914
rect 3873 9909 3879 9913
rect 3883 9909 3889 9913
rect 3893 9909 3899 9913
rect 3903 9909 3909 9913
rect 3913 9909 4029 9913
rect 4033 9909 4039 9913
rect 4043 9909 4049 9913
rect 4053 9909 4059 9913
rect 4063 9909 4069 9913
rect 3869 9908 4073 9909
rect 3869 9904 3874 9908
rect 3878 9904 3884 9908
rect 3888 9904 3894 9908
rect 3898 9904 3904 9908
rect 3908 9904 4034 9908
rect 4038 9904 4044 9908
rect 4048 9904 4054 9908
rect 4058 9904 4064 9908
rect 4068 9904 4073 9908
rect 3869 9903 4073 9904
rect 3873 9899 3879 9903
rect 3883 9899 3889 9903
rect 3893 9899 3899 9903
rect 3903 9899 3909 9903
rect 3913 9899 4029 9903
rect 4033 9899 4039 9903
rect 4043 9899 4049 9903
rect 4053 9899 4059 9903
rect 4063 9899 4069 9903
rect 3869 9898 4073 9899
rect 3869 9894 3874 9898
rect 3878 9894 3884 9898
rect 3888 9894 3894 9898
rect 3898 9894 3904 9898
rect 3908 9894 4034 9898
rect 4038 9894 4044 9898
rect 4048 9894 4054 9898
rect 4058 9894 4064 9898
rect 4068 9894 4073 9898
rect 3869 9893 4073 9894
rect 3873 9889 3879 9893
rect 3883 9889 3889 9893
rect 3893 9889 3899 9893
rect 3903 9889 3909 9893
rect 3913 9889 4029 9893
rect 4033 9889 4039 9893
rect 4043 9889 4049 9893
rect 4053 9889 4059 9893
rect 4063 9889 4069 9893
rect 3869 9888 4073 9889
rect 3869 9884 3874 9888
rect 3878 9884 3884 9888
rect 3888 9884 3894 9888
rect 3898 9884 3904 9888
rect 3908 9884 4034 9888
rect 4038 9884 4044 9888
rect 4048 9884 4054 9888
rect 4058 9884 4064 9888
rect 4068 9884 4073 9888
rect 3869 9883 4073 9884
rect 3873 9879 3879 9883
rect 3883 9879 3889 9883
rect 3893 9879 3899 9883
rect 3903 9879 3909 9883
rect 3913 9879 4029 9883
rect 4033 9879 4039 9883
rect 4043 9879 4049 9883
rect 4053 9879 4059 9883
rect 4063 9879 4069 9883
rect 3869 9878 4073 9879
rect 3869 9874 3874 9878
rect 3878 9874 3884 9878
rect 3888 9874 3894 9878
rect 3898 9874 3904 9878
rect 3908 9874 4034 9878
rect 4038 9874 4044 9878
rect 4048 9874 4054 9878
rect 4058 9874 4064 9878
rect 4068 9874 4073 9878
rect 3869 9873 4073 9874
rect 3873 9869 3879 9873
rect 3883 9869 3889 9873
rect 3893 9869 3899 9873
rect 3903 9869 3909 9873
rect 3913 9869 4029 9873
rect 4033 9869 4039 9873
rect 4043 9869 4049 9873
rect 4053 9869 4059 9873
rect 4063 9869 4069 9873
rect 3869 9868 4073 9869
rect 3869 9864 3874 9868
rect 3878 9864 3884 9868
rect 3888 9864 3894 9868
rect 3898 9864 3904 9868
rect 3908 9864 4034 9868
rect 4038 9864 4044 9868
rect 4048 9864 4054 9868
rect 4058 9864 4064 9868
rect 4068 9864 4073 9868
rect 1389 9848 1392 9852
rect 1396 9848 1397 9852
rect 1401 9848 1402 9852
rect 1406 9848 1407 9852
rect 1411 9848 1412 9852
rect 1416 9848 1417 9852
rect 1421 9848 1422 9852
rect 1426 9848 1427 9852
rect 1431 9848 1432 9852
rect 1436 9848 1437 9852
rect 1441 9848 1442 9852
rect 1446 9848 1449 9852
rect 1352 9800 1373 9802
rect 1352 9796 1354 9800
rect 1358 9796 1359 9800
rect 1363 9796 1364 9800
rect 1368 9796 1369 9800
rect 1352 9795 1373 9796
rect 1352 9791 1354 9795
rect 1358 9791 1359 9795
rect 1363 9791 1364 9795
rect 1368 9791 1369 9795
rect 1352 9790 1373 9791
rect 1352 9786 1354 9790
rect 1358 9786 1359 9790
rect 1363 9786 1364 9790
rect 1368 9786 1369 9790
rect 118 9348 593 9786
rect 1352 9785 1373 9786
rect 1352 9781 1354 9785
rect 1358 9781 1359 9785
rect 1363 9781 1364 9785
rect 1368 9781 1369 9785
rect 1352 9780 1373 9781
rect 1352 9776 1354 9780
rect 1358 9776 1359 9780
rect 1363 9776 1364 9780
rect 1368 9776 1369 9780
rect 1352 9775 1373 9776
rect 1352 9771 1354 9775
rect 1358 9771 1359 9775
rect 1363 9771 1364 9775
rect 1368 9771 1369 9775
rect 1352 9770 1373 9771
rect 1352 9766 1354 9770
rect 1358 9766 1359 9770
rect 1363 9766 1364 9770
rect 1368 9766 1369 9770
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 802 9761 821 9762
rect 806 9757 807 9761
rect 811 9757 812 9761
rect 816 9757 817 9761
rect 802 9756 821 9757
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 802 9751 821 9752
rect 806 9747 807 9751
rect 811 9747 812 9751
rect 816 9747 817 9751
rect 802 9746 821 9747
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 802 9741 821 9742
rect 806 9737 807 9741
rect 811 9737 812 9741
rect 816 9737 817 9741
rect 802 9736 821 9737
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 831 9761 850 9762
rect 835 9757 836 9761
rect 840 9757 841 9761
rect 845 9757 846 9761
rect 831 9756 850 9757
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 831 9751 850 9752
rect 835 9747 836 9751
rect 840 9747 841 9751
rect 845 9747 846 9751
rect 831 9746 850 9747
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 831 9741 850 9742
rect 835 9737 836 9741
rect 840 9737 841 9741
rect 845 9737 846 9741
rect 831 9736 850 9737
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 860 9761 879 9762
rect 864 9757 865 9761
rect 869 9757 870 9761
rect 874 9757 875 9761
rect 860 9756 879 9757
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 860 9751 879 9752
rect 864 9747 865 9751
rect 869 9747 870 9751
rect 874 9747 875 9751
rect 860 9746 879 9747
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 860 9741 879 9742
rect 864 9737 865 9741
rect 869 9737 870 9741
rect 874 9737 875 9741
rect 860 9736 879 9737
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 889 9761 908 9762
rect 893 9757 894 9761
rect 898 9757 899 9761
rect 903 9757 904 9761
rect 889 9756 908 9757
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 889 9751 908 9752
rect 893 9747 894 9751
rect 898 9747 899 9751
rect 903 9747 904 9751
rect 889 9746 908 9747
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 889 9741 908 9742
rect 893 9737 894 9741
rect 898 9737 899 9741
rect 903 9737 904 9741
rect 889 9736 908 9737
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 918 9761 937 9762
rect 922 9757 923 9761
rect 927 9757 928 9761
rect 932 9757 933 9761
rect 918 9756 937 9757
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 918 9751 937 9752
rect 922 9747 923 9751
rect 927 9747 928 9751
rect 932 9747 933 9751
rect 918 9746 937 9747
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 918 9741 937 9742
rect 922 9737 923 9741
rect 927 9737 928 9741
rect 932 9737 933 9741
rect 918 9736 937 9737
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1319 9761 1338 9762
rect 1323 9757 1324 9761
rect 1328 9757 1329 9761
rect 1333 9757 1334 9761
rect 1319 9756 1338 9757
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1319 9751 1338 9752
rect 1323 9747 1324 9751
rect 1328 9747 1329 9751
rect 1333 9747 1334 9751
rect 1319 9746 1338 9747
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1319 9741 1338 9742
rect 1323 9737 1324 9741
rect 1328 9737 1329 9741
rect 1333 9737 1334 9741
rect 1319 9736 1338 9737
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1352 9765 1373 9766
rect 1352 9761 1354 9765
rect 1358 9761 1359 9765
rect 1363 9761 1364 9765
rect 1368 9761 1369 9765
rect 1352 9760 1373 9761
rect 1352 9756 1354 9760
rect 1358 9756 1359 9760
rect 1363 9756 1364 9760
rect 1368 9756 1369 9760
rect 1352 9755 1373 9756
rect 1352 9751 1354 9755
rect 1358 9751 1359 9755
rect 1363 9751 1364 9755
rect 1368 9751 1369 9755
rect 1352 9750 1373 9751
rect 1352 9746 1354 9750
rect 1358 9746 1359 9750
rect 1363 9746 1364 9750
rect 1368 9746 1369 9750
rect 1352 9745 1373 9746
rect 1352 9741 1354 9745
rect 1358 9741 1359 9745
rect 1363 9741 1364 9745
rect 1368 9741 1369 9745
rect 1352 9740 1373 9741
rect 1352 9736 1354 9740
rect 1358 9736 1359 9740
rect 1363 9736 1364 9740
rect 1368 9736 1369 9740
rect 1352 9734 1373 9736
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 802 9715 821 9716
rect 806 9711 807 9715
rect 811 9711 812 9715
rect 816 9711 817 9715
rect 802 9710 821 9711
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 802 9705 821 9706
rect 806 9701 807 9705
rect 811 9701 812 9705
rect 816 9701 817 9705
rect 802 9700 821 9701
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 802 9695 821 9696
rect 806 9691 807 9695
rect 811 9691 812 9695
rect 816 9691 817 9695
rect 802 9690 821 9691
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 831 9715 850 9716
rect 835 9711 836 9715
rect 840 9711 841 9715
rect 845 9711 846 9715
rect 831 9710 850 9711
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 831 9705 850 9706
rect 835 9701 836 9705
rect 840 9701 841 9705
rect 845 9701 846 9705
rect 831 9700 850 9701
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 831 9695 850 9696
rect 835 9691 836 9695
rect 840 9691 841 9695
rect 845 9691 846 9695
rect 831 9690 850 9691
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 860 9715 879 9716
rect 864 9711 865 9715
rect 869 9711 870 9715
rect 874 9711 875 9715
rect 860 9710 879 9711
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 860 9705 879 9706
rect 864 9701 865 9705
rect 869 9701 870 9705
rect 874 9701 875 9705
rect 860 9700 879 9701
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 860 9695 879 9696
rect 864 9691 865 9695
rect 869 9691 870 9695
rect 874 9691 875 9695
rect 860 9690 879 9691
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 889 9715 908 9716
rect 893 9711 894 9715
rect 898 9711 899 9715
rect 903 9711 904 9715
rect 889 9710 908 9711
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 889 9705 908 9706
rect 893 9701 894 9705
rect 898 9701 899 9705
rect 903 9701 904 9705
rect 889 9700 908 9701
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 889 9695 908 9696
rect 893 9691 894 9695
rect 898 9691 899 9695
rect 903 9691 904 9695
rect 889 9690 908 9691
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 918 9715 937 9716
rect 922 9711 923 9715
rect 927 9711 928 9715
rect 932 9711 933 9715
rect 918 9710 937 9711
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 918 9705 937 9706
rect 922 9701 923 9705
rect 927 9701 928 9705
rect 932 9701 933 9705
rect 918 9700 937 9701
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 918 9695 937 9696
rect 922 9691 923 9695
rect 927 9691 928 9695
rect 932 9691 933 9695
rect 918 9690 937 9691
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1319 9715 1338 9716
rect 1323 9711 1324 9715
rect 1328 9711 1329 9715
rect 1333 9711 1334 9715
rect 1319 9710 1338 9711
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1319 9705 1338 9706
rect 1323 9701 1324 9705
rect 1328 9701 1329 9705
rect 1333 9701 1334 9705
rect 1319 9700 1338 9701
rect 1385 9712 1453 9848
rect 1549 9848 1552 9852
rect 1556 9848 1557 9852
rect 1561 9848 1562 9852
rect 1566 9848 1567 9852
rect 1571 9848 1572 9852
rect 1576 9848 1577 9852
rect 1581 9848 1582 9852
rect 1586 9848 1587 9852
rect 1591 9848 1592 9852
rect 1596 9848 1597 9852
rect 1601 9848 1602 9852
rect 1606 9848 1609 9852
rect 1545 9769 1613 9848
rect 1698 9848 1701 9852
rect 1705 9848 1706 9852
rect 1710 9848 1711 9852
rect 1715 9848 1716 9852
rect 1720 9848 1721 9852
rect 1725 9848 1726 9852
rect 1730 9848 1731 9852
rect 1735 9848 1736 9852
rect 1740 9848 1741 9852
rect 1745 9848 1746 9852
rect 1750 9848 1751 9852
rect 1755 9848 1758 9852
rect 1545 9765 1547 9769
rect 1551 9765 1552 9769
rect 1556 9765 1557 9769
rect 1561 9765 1562 9769
rect 1566 9765 1567 9769
rect 1571 9765 1572 9769
rect 1576 9765 1577 9769
rect 1581 9765 1582 9769
rect 1586 9765 1587 9769
rect 1591 9765 1592 9769
rect 1596 9765 1597 9769
rect 1601 9765 1602 9769
rect 1606 9765 1607 9769
rect 1611 9765 1613 9769
rect 1661 9800 1682 9802
rect 1661 9796 1663 9800
rect 1667 9796 1668 9800
rect 1672 9796 1673 9800
rect 1677 9796 1678 9800
rect 1661 9795 1682 9796
rect 1661 9791 1663 9795
rect 1667 9791 1668 9795
rect 1672 9791 1673 9795
rect 1677 9791 1678 9795
rect 1661 9790 1682 9791
rect 1661 9786 1663 9790
rect 1667 9786 1668 9790
rect 1672 9786 1673 9790
rect 1677 9786 1678 9790
rect 1661 9785 1682 9786
rect 1661 9781 1663 9785
rect 1667 9781 1668 9785
rect 1672 9781 1673 9785
rect 1677 9781 1678 9785
rect 1661 9780 1682 9781
rect 1661 9776 1663 9780
rect 1667 9776 1668 9780
rect 1672 9776 1673 9780
rect 1677 9776 1678 9780
rect 1661 9775 1682 9776
rect 1661 9771 1663 9775
rect 1667 9771 1668 9775
rect 1672 9771 1673 9775
rect 1677 9771 1678 9775
rect 1661 9770 1682 9771
rect 1661 9766 1663 9770
rect 1667 9766 1668 9770
rect 1672 9766 1673 9770
rect 1677 9766 1678 9770
rect 1545 9764 1613 9765
rect 1545 9760 1547 9764
rect 1551 9760 1552 9764
rect 1556 9760 1557 9764
rect 1561 9760 1562 9764
rect 1566 9760 1567 9764
rect 1571 9760 1572 9764
rect 1576 9760 1577 9764
rect 1581 9760 1582 9764
rect 1586 9760 1587 9764
rect 1591 9760 1592 9764
rect 1596 9760 1597 9764
rect 1601 9760 1602 9764
rect 1606 9760 1607 9764
rect 1611 9760 1613 9764
rect 1545 9757 1613 9760
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1628 9761 1647 9762
rect 1632 9757 1633 9761
rect 1637 9757 1638 9761
rect 1642 9757 1643 9761
rect 1628 9756 1647 9757
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1628 9751 1647 9752
rect 1632 9747 1633 9751
rect 1637 9747 1638 9751
rect 1642 9747 1643 9751
rect 1628 9746 1647 9747
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1628 9741 1647 9742
rect 1632 9737 1633 9741
rect 1637 9737 1638 9741
rect 1642 9737 1643 9741
rect 1628 9736 1647 9737
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1661 9765 1682 9766
rect 1661 9761 1663 9765
rect 1667 9761 1668 9765
rect 1672 9761 1673 9765
rect 1677 9761 1678 9765
rect 1661 9760 1682 9761
rect 1661 9756 1663 9760
rect 1667 9756 1668 9760
rect 1672 9756 1673 9760
rect 1677 9756 1678 9760
rect 1661 9755 1682 9756
rect 1661 9751 1663 9755
rect 1667 9751 1668 9755
rect 1672 9751 1673 9755
rect 1677 9751 1678 9755
rect 1661 9750 1682 9751
rect 1661 9746 1663 9750
rect 1667 9746 1668 9750
rect 1672 9746 1673 9750
rect 1677 9746 1678 9750
rect 1661 9745 1682 9746
rect 1661 9741 1663 9745
rect 1667 9741 1668 9745
rect 1672 9741 1673 9745
rect 1677 9741 1678 9745
rect 1661 9740 1682 9741
rect 1661 9736 1663 9740
rect 1667 9736 1668 9740
rect 1672 9736 1673 9740
rect 1677 9736 1678 9740
rect 1661 9734 1682 9736
rect 1573 9718 1574 9722
rect 1578 9718 1579 9722
rect 1583 9718 1584 9722
rect 1588 9718 1589 9722
rect 1593 9718 1594 9722
rect 1598 9718 1599 9722
rect 1603 9718 1604 9722
rect 1608 9718 1609 9722
rect 1613 9718 1614 9722
rect 1618 9718 1619 9722
rect 1623 9718 1625 9722
rect 1569 9717 1625 9718
rect 1385 9708 1387 9712
rect 1391 9708 1392 9712
rect 1396 9708 1397 9712
rect 1401 9708 1402 9712
rect 1406 9708 1407 9712
rect 1411 9708 1412 9712
rect 1416 9708 1417 9712
rect 1421 9708 1422 9712
rect 1426 9708 1427 9712
rect 1431 9708 1432 9712
rect 1436 9708 1437 9712
rect 1441 9708 1442 9712
rect 1446 9708 1447 9712
rect 1451 9708 1453 9712
rect 1385 9707 1453 9708
rect 1385 9703 1387 9707
rect 1391 9703 1392 9707
rect 1396 9703 1397 9707
rect 1401 9703 1402 9707
rect 1406 9703 1407 9707
rect 1411 9703 1412 9707
rect 1416 9703 1417 9707
rect 1421 9703 1422 9707
rect 1426 9703 1427 9707
rect 1431 9703 1432 9707
rect 1436 9703 1437 9707
rect 1441 9703 1442 9707
rect 1446 9703 1447 9707
rect 1451 9703 1453 9707
rect 1385 9700 1453 9703
rect 1488 9711 1489 9715
rect 1493 9711 1494 9715
rect 1498 9711 1499 9715
rect 1503 9711 1504 9715
rect 1488 9710 1508 9711
rect 1488 9706 1489 9710
rect 1493 9706 1494 9710
rect 1498 9706 1499 9710
rect 1503 9706 1504 9710
rect 1488 9705 1508 9706
rect 1488 9701 1489 9705
rect 1493 9701 1494 9705
rect 1498 9701 1499 9705
rect 1503 9701 1504 9705
rect 1573 9713 1574 9717
rect 1578 9713 1579 9717
rect 1583 9713 1584 9717
rect 1588 9713 1589 9717
rect 1593 9713 1594 9717
rect 1598 9713 1599 9717
rect 1603 9713 1604 9717
rect 1608 9713 1609 9717
rect 1613 9713 1614 9717
rect 1618 9713 1619 9717
rect 1623 9713 1625 9717
rect 1569 9712 1625 9713
rect 1573 9708 1574 9712
rect 1578 9708 1579 9712
rect 1583 9708 1584 9712
rect 1588 9708 1589 9712
rect 1593 9708 1594 9712
rect 1598 9708 1599 9712
rect 1603 9708 1604 9712
rect 1608 9708 1609 9712
rect 1613 9708 1614 9712
rect 1618 9708 1619 9712
rect 1623 9708 1625 9712
rect 1569 9707 1625 9708
rect 1573 9703 1574 9707
rect 1578 9703 1579 9707
rect 1583 9703 1584 9707
rect 1588 9703 1589 9707
rect 1593 9703 1594 9707
rect 1598 9703 1599 9707
rect 1603 9703 1604 9707
rect 1608 9703 1609 9707
rect 1613 9703 1614 9707
rect 1618 9703 1619 9707
rect 1623 9703 1625 9707
rect 1569 9701 1625 9703
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1628 9715 1647 9716
rect 1632 9711 1633 9715
rect 1637 9711 1638 9715
rect 1642 9711 1643 9715
rect 1628 9710 1647 9711
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1628 9705 1647 9706
rect 1632 9701 1633 9705
rect 1637 9701 1638 9705
rect 1642 9701 1643 9705
rect 1488 9700 1508 9701
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1319 9695 1338 9696
rect 1323 9691 1324 9695
rect 1328 9691 1329 9695
rect 1333 9691 1334 9695
rect 1319 9690 1338 9691
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1488 9696 1489 9700
rect 1493 9696 1494 9700
rect 1498 9696 1499 9700
rect 1503 9696 1504 9700
rect 1488 9695 1508 9696
rect 1488 9691 1489 9695
rect 1493 9691 1494 9695
rect 1498 9691 1499 9695
rect 1503 9691 1504 9695
rect 1488 9690 1508 9691
rect 1488 9686 1489 9690
rect 1493 9686 1494 9690
rect 1498 9686 1499 9690
rect 1503 9686 1504 9690
rect 1628 9700 1647 9701
rect 1694 9712 1762 9848
rect 1858 9848 1861 9852
rect 1865 9848 1866 9852
rect 1870 9848 1871 9852
rect 1875 9848 1876 9852
rect 1880 9848 1881 9852
rect 1885 9848 1886 9852
rect 1890 9848 1891 9852
rect 1895 9848 1896 9852
rect 1900 9848 1901 9852
rect 1905 9848 1906 9852
rect 1910 9848 1911 9852
rect 1915 9848 1918 9852
rect 1778 9815 1782 9827
rect 1778 9799 1782 9811
rect 1778 9783 1782 9795
rect 1836 9815 1840 9827
rect 1836 9799 1840 9811
rect 1836 9783 1840 9795
rect 1854 9769 1922 9848
rect 2007 9848 2010 9852
rect 2014 9848 2015 9852
rect 2019 9848 2020 9852
rect 2024 9848 2025 9852
rect 2029 9848 2030 9852
rect 2034 9848 2035 9852
rect 2039 9848 2040 9852
rect 2044 9848 2045 9852
rect 2049 9848 2050 9852
rect 2054 9848 2055 9852
rect 2059 9848 2060 9852
rect 2064 9848 2067 9852
rect 1854 9765 1856 9769
rect 1860 9765 1861 9769
rect 1865 9765 1866 9769
rect 1870 9765 1871 9769
rect 1875 9765 1876 9769
rect 1880 9765 1881 9769
rect 1885 9765 1886 9769
rect 1890 9765 1891 9769
rect 1895 9765 1896 9769
rect 1900 9765 1901 9769
rect 1905 9765 1906 9769
rect 1910 9765 1911 9769
rect 1915 9765 1916 9769
rect 1920 9765 1922 9769
rect 1970 9800 1991 9802
rect 1970 9796 1972 9800
rect 1976 9796 1977 9800
rect 1981 9796 1982 9800
rect 1986 9796 1987 9800
rect 1970 9795 1991 9796
rect 1970 9791 1972 9795
rect 1976 9791 1977 9795
rect 1981 9791 1982 9795
rect 1986 9791 1987 9795
rect 1970 9790 1991 9791
rect 1970 9786 1972 9790
rect 1976 9786 1977 9790
rect 1981 9786 1982 9790
rect 1986 9786 1987 9790
rect 1970 9785 1991 9786
rect 1970 9781 1972 9785
rect 1976 9781 1977 9785
rect 1981 9781 1982 9785
rect 1986 9781 1987 9785
rect 1970 9780 1991 9781
rect 1970 9776 1972 9780
rect 1976 9776 1977 9780
rect 1981 9776 1982 9780
rect 1986 9776 1987 9780
rect 1970 9775 1991 9776
rect 1970 9771 1972 9775
rect 1976 9771 1977 9775
rect 1981 9771 1982 9775
rect 1986 9771 1987 9775
rect 1970 9770 1991 9771
rect 1970 9766 1972 9770
rect 1976 9766 1977 9770
rect 1981 9766 1982 9770
rect 1986 9766 1987 9770
rect 1854 9764 1922 9765
rect 1854 9760 1856 9764
rect 1860 9760 1861 9764
rect 1865 9760 1866 9764
rect 1870 9760 1871 9764
rect 1875 9760 1876 9764
rect 1880 9760 1881 9764
rect 1885 9760 1886 9764
rect 1890 9760 1891 9764
rect 1895 9760 1896 9764
rect 1900 9760 1901 9764
rect 1905 9760 1906 9764
rect 1910 9760 1911 9764
rect 1915 9760 1916 9764
rect 1920 9760 1922 9764
rect 1854 9757 1922 9760
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1937 9761 1956 9762
rect 1941 9757 1942 9761
rect 1946 9757 1947 9761
rect 1951 9757 1952 9761
rect 1937 9756 1956 9757
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1937 9751 1956 9752
rect 1941 9747 1942 9751
rect 1946 9747 1947 9751
rect 1951 9747 1952 9751
rect 1937 9746 1956 9747
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1937 9741 1956 9742
rect 1941 9737 1942 9741
rect 1946 9737 1947 9741
rect 1951 9737 1952 9741
rect 1937 9736 1956 9737
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1970 9765 1991 9766
rect 1970 9761 1972 9765
rect 1976 9761 1977 9765
rect 1981 9761 1982 9765
rect 1986 9761 1987 9765
rect 1970 9760 1991 9761
rect 1970 9756 1972 9760
rect 1976 9756 1977 9760
rect 1981 9756 1982 9760
rect 1986 9756 1987 9760
rect 1970 9755 1991 9756
rect 1970 9751 1972 9755
rect 1976 9751 1977 9755
rect 1981 9751 1982 9755
rect 1986 9751 1987 9755
rect 1970 9750 1991 9751
rect 1970 9746 1972 9750
rect 1976 9746 1977 9750
rect 1981 9746 1982 9750
rect 1986 9746 1987 9750
rect 1970 9745 1991 9746
rect 1970 9741 1972 9745
rect 1976 9741 1977 9745
rect 1981 9741 1982 9745
rect 1986 9741 1987 9745
rect 1970 9740 1991 9741
rect 1970 9736 1972 9740
rect 1976 9736 1977 9740
rect 1981 9736 1982 9740
rect 1986 9736 1987 9740
rect 1970 9734 1991 9736
rect 1694 9708 1696 9712
rect 1700 9708 1701 9712
rect 1705 9708 1706 9712
rect 1710 9708 1711 9712
rect 1715 9708 1716 9712
rect 1720 9708 1721 9712
rect 1725 9708 1726 9712
rect 1730 9708 1731 9712
rect 1735 9708 1736 9712
rect 1740 9708 1741 9712
rect 1745 9708 1746 9712
rect 1750 9708 1751 9712
rect 1755 9708 1756 9712
rect 1760 9708 1762 9712
rect 1694 9707 1762 9708
rect 1694 9703 1696 9707
rect 1700 9703 1701 9707
rect 1705 9703 1706 9707
rect 1710 9703 1711 9707
rect 1715 9703 1716 9707
rect 1720 9703 1721 9707
rect 1725 9703 1726 9707
rect 1730 9703 1731 9707
rect 1735 9703 1736 9707
rect 1740 9703 1741 9707
rect 1745 9703 1746 9707
rect 1750 9703 1751 9707
rect 1755 9703 1756 9707
rect 1760 9703 1762 9707
rect 1694 9700 1762 9703
rect 1882 9718 1883 9722
rect 1887 9718 1888 9722
rect 1892 9718 1893 9722
rect 1897 9718 1898 9722
rect 1902 9718 1903 9722
rect 1907 9718 1908 9722
rect 1912 9718 1913 9722
rect 1917 9718 1918 9722
rect 1922 9718 1923 9722
rect 1927 9718 1928 9722
rect 1932 9718 1934 9722
rect 1878 9717 1934 9718
rect 1882 9713 1883 9717
rect 1887 9713 1888 9717
rect 1892 9713 1893 9717
rect 1897 9713 1898 9717
rect 1902 9713 1903 9717
rect 1907 9713 1908 9717
rect 1912 9713 1913 9717
rect 1917 9713 1918 9717
rect 1922 9713 1923 9717
rect 1927 9713 1928 9717
rect 1932 9713 1934 9717
rect 1878 9712 1934 9713
rect 1882 9708 1883 9712
rect 1887 9708 1888 9712
rect 1892 9708 1893 9712
rect 1897 9708 1898 9712
rect 1902 9708 1903 9712
rect 1907 9708 1908 9712
rect 1912 9708 1913 9712
rect 1917 9708 1918 9712
rect 1922 9708 1923 9712
rect 1927 9708 1928 9712
rect 1932 9708 1934 9712
rect 1878 9707 1934 9708
rect 1882 9703 1883 9707
rect 1887 9703 1888 9707
rect 1892 9703 1893 9707
rect 1897 9703 1898 9707
rect 1902 9703 1903 9707
rect 1907 9703 1908 9707
rect 1912 9703 1913 9707
rect 1917 9703 1918 9707
rect 1922 9703 1923 9707
rect 1927 9703 1928 9707
rect 1932 9703 1934 9707
rect 1878 9701 1934 9703
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1937 9715 1956 9716
rect 1941 9711 1942 9715
rect 1946 9711 1947 9715
rect 1951 9711 1952 9715
rect 1937 9710 1956 9711
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1937 9705 1956 9706
rect 1941 9701 1942 9705
rect 1946 9701 1947 9705
rect 1951 9701 1952 9705
rect 1937 9700 1956 9701
rect 2003 9712 2071 9848
rect 2167 9848 2170 9852
rect 2174 9848 2175 9852
rect 2179 9848 2180 9852
rect 2184 9848 2185 9852
rect 2189 9848 2190 9852
rect 2194 9848 2195 9852
rect 2199 9848 2200 9852
rect 2204 9848 2205 9852
rect 2209 9848 2210 9852
rect 2214 9848 2215 9852
rect 2219 9848 2220 9852
rect 2224 9848 2227 9852
rect 2087 9815 2091 9827
rect 2087 9799 2091 9811
rect 2087 9783 2091 9795
rect 2145 9815 2149 9827
rect 2145 9799 2149 9811
rect 2145 9783 2149 9795
rect 2163 9769 2231 9848
rect 2316 9848 2319 9852
rect 2323 9848 2324 9852
rect 2328 9848 2329 9852
rect 2333 9848 2334 9852
rect 2338 9848 2339 9852
rect 2343 9848 2344 9852
rect 2348 9848 2349 9852
rect 2353 9848 2354 9852
rect 2358 9848 2359 9852
rect 2363 9848 2364 9852
rect 2368 9848 2369 9852
rect 2373 9848 2376 9852
rect 2163 9765 2165 9769
rect 2169 9765 2170 9769
rect 2174 9765 2175 9769
rect 2179 9765 2180 9769
rect 2184 9765 2185 9769
rect 2189 9765 2190 9769
rect 2194 9765 2195 9769
rect 2199 9765 2200 9769
rect 2204 9765 2205 9769
rect 2209 9765 2210 9769
rect 2214 9765 2215 9769
rect 2219 9765 2220 9769
rect 2224 9765 2225 9769
rect 2229 9765 2231 9769
rect 2279 9800 2300 9802
rect 2279 9796 2281 9800
rect 2285 9796 2286 9800
rect 2290 9796 2291 9800
rect 2295 9796 2296 9800
rect 2279 9795 2300 9796
rect 2279 9791 2281 9795
rect 2285 9791 2286 9795
rect 2290 9791 2291 9795
rect 2295 9791 2296 9795
rect 2279 9790 2300 9791
rect 2279 9786 2281 9790
rect 2285 9786 2286 9790
rect 2290 9786 2291 9790
rect 2295 9786 2296 9790
rect 2279 9785 2300 9786
rect 2279 9781 2281 9785
rect 2285 9781 2286 9785
rect 2290 9781 2291 9785
rect 2295 9781 2296 9785
rect 2279 9780 2300 9781
rect 2279 9776 2281 9780
rect 2285 9776 2286 9780
rect 2290 9776 2291 9780
rect 2295 9776 2296 9780
rect 2279 9775 2300 9776
rect 2279 9771 2281 9775
rect 2285 9771 2286 9775
rect 2290 9771 2291 9775
rect 2295 9771 2296 9775
rect 2279 9770 2300 9771
rect 2279 9766 2281 9770
rect 2285 9766 2286 9770
rect 2290 9766 2291 9770
rect 2295 9766 2296 9770
rect 2163 9764 2231 9765
rect 2163 9760 2165 9764
rect 2169 9760 2170 9764
rect 2174 9760 2175 9764
rect 2179 9760 2180 9764
rect 2184 9760 2185 9764
rect 2189 9760 2190 9764
rect 2194 9760 2195 9764
rect 2199 9760 2200 9764
rect 2204 9760 2205 9764
rect 2209 9760 2210 9764
rect 2214 9760 2215 9764
rect 2219 9760 2220 9764
rect 2224 9760 2225 9764
rect 2229 9760 2231 9764
rect 2163 9757 2231 9760
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2246 9761 2265 9762
rect 2250 9757 2251 9761
rect 2255 9757 2256 9761
rect 2260 9757 2261 9761
rect 2246 9756 2265 9757
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2246 9751 2265 9752
rect 2250 9747 2251 9751
rect 2255 9747 2256 9751
rect 2260 9747 2261 9751
rect 2246 9746 2265 9747
rect 2003 9708 2005 9712
rect 2009 9708 2010 9712
rect 2014 9708 2015 9712
rect 2019 9708 2020 9712
rect 2024 9708 2025 9712
rect 2029 9708 2030 9712
rect 2034 9708 2035 9712
rect 2039 9708 2040 9712
rect 2044 9708 2045 9712
rect 2049 9708 2050 9712
rect 2054 9708 2055 9712
rect 2059 9708 2060 9712
rect 2064 9708 2065 9712
rect 2069 9708 2071 9712
rect 2003 9707 2071 9708
rect 2003 9703 2005 9707
rect 2009 9703 2010 9707
rect 2014 9703 2015 9707
rect 2019 9703 2020 9707
rect 2024 9703 2025 9707
rect 2029 9703 2030 9707
rect 2034 9703 2035 9707
rect 2039 9703 2040 9707
rect 2044 9703 2045 9707
rect 2049 9703 2050 9707
rect 2054 9703 2055 9707
rect 2059 9703 2060 9707
rect 2064 9703 2065 9707
rect 2069 9703 2071 9707
rect 2003 9700 2071 9703
rect 2166 9741 2174 9743
rect 2166 9736 2167 9741
rect 2172 9736 2174 9741
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1628 9695 1647 9696
rect 1632 9691 1633 9695
rect 1637 9691 1638 9695
rect 1642 9691 1643 9695
rect 1628 9690 1647 9691
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1937 9695 1956 9696
rect 1941 9691 1942 9695
rect 1946 9691 1947 9695
rect 1951 9691 1952 9695
rect 1937 9690 1956 9691
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 1488 9685 1508 9686
rect 1488 9681 1489 9685
rect 1493 9681 1494 9685
rect 1498 9681 1499 9685
rect 1503 9681 1504 9685
rect 1488 9680 1508 9681
rect 1488 9676 1489 9680
rect 1493 9676 1494 9680
rect 1498 9676 1499 9680
rect 1503 9676 1504 9680
rect 1488 9675 1508 9676
rect 1488 9671 1489 9675
rect 1493 9671 1494 9675
rect 1498 9671 1499 9675
rect 1503 9671 1504 9675
rect 1488 9670 1508 9671
rect 1488 9666 1489 9670
rect 1493 9666 1494 9670
rect 1498 9666 1499 9670
rect 1503 9666 1504 9670
rect 1488 9665 1508 9666
rect 1488 9661 1489 9665
rect 1493 9661 1494 9665
rect 1498 9661 1499 9665
rect 1503 9661 1504 9665
rect 1488 9659 1508 9661
rect 2166 9623 2174 9736
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2246 9741 2265 9742
rect 2250 9737 2251 9741
rect 2255 9737 2256 9741
rect 2260 9737 2261 9741
rect 2246 9736 2265 9737
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2279 9765 2300 9766
rect 2279 9761 2281 9765
rect 2285 9761 2286 9765
rect 2290 9761 2291 9765
rect 2295 9761 2296 9765
rect 2279 9760 2300 9761
rect 2279 9756 2281 9760
rect 2285 9756 2286 9760
rect 2290 9756 2291 9760
rect 2295 9756 2296 9760
rect 2279 9755 2300 9756
rect 2279 9751 2281 9755
rect 2285 9751 2286 9755
rect 2290 9751 2291 9755
rect 2295 9751 2296 9755
rect 2279 9750 2300 9751
rect 2279 9746 2281 9750
rect 2285 9746 2286 9750
rect 2290 9746 2291 9750
rect 2295 9746 2296 9750
rect 2279 9745 2300 9746
rect 2279 9741 2281 9745
rect 2285 9741 2286 9745
rect 2290 9741 2291 9745
rect 2295 9741 2296 9745
rect 2279 9740 2300 9741
rect 2279 9736 2281 9740
rect 2285 9736 2286 9740
rect 2290 9736 2291 9740
rect 2295 9736 2296 9740
rect 2279 9734 2300 9736
rect 2191 9718 2192 9722
rect 2196 9718 2197 9722
rect 2201 9718 2202 9722
rect 2206 9718 2207 9722
rect 2211 9718 2212 9722
rect 2216 9718 2217 9722
rect 2221 9718 2222 9722
rect 2226 9718 2227 9722
rect 2231 9718 2232 9722
rect 2236 9718 2237 9722
rect 2241 9718 2243 9722
rect 2187 9717 2243 9718
rect 2191 9713 2192 9717
rect 2196 9713 2197 9717
rect 2201 9713 2202 9717
rect 2206 9713 2207 9717
rect 2211 9713 2212 9717
rect 2216 9713 2217 9717
rect 2221 9713 2222 9717
rect 2226 9713 2227 9717
rect 2231 9713 2232 9717
rect 2236 9713 2237 9717
rect 2241 9713 2243 9717
rect 2187 9712 2243 9713
rect 2191 9708 2192 9712
rect 2196 9708 2197 9712
rect 2201 9708 2202 9712
rect 2206 9708 2207 9712
rect 2211 9708 2212 9712
rect 2216 9708 2217 9712
rect 2221 9708 2222 9712
rect 2226 9708 2227 9712
rect 2231 9708 2232 9712
rect 2236 9708 2237 9712
rect 2241 9708 2243 9712
rect 2187 9707 2243 9708
rect 2191 9703 2192 9707
rect 2196 9703 2197 9707
rect 2201 9703 2202 9707
rect 2206 9703 2207 9707
rect 2211 9703 2212 9707
rect 2216 9703 2217 9707
rect 2221 9703 2222 9707
rect 2226 9703 2227 9707
rect 2231 9703 2232 9707
rect 2236 9703 2237 9707
rect 2241 9703 2243 9707
rect 2187 9701 2243 9703
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2246 9715 2265 9716
rect 2250 9711 2251 9715
rect 2255 9711 2256 9715
rect 2260 9711 2261 9715
rect 2246 9710 2265 9711
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2246 9705 2265 9706
rect 2250 9701 2251 9705
rect 2255 9701 2256 9705
rect 2260 9701 2261 9705
rect 2246 9700 2265 9701
rect 2312 9712 2380 9848
rect 2476 9848 2479 9852
rect 2483 9848 2484 9852
rect 2488 9848 2489 9852
rect 2493 9848 2494 9852
rect 2498 9848 2499 9852
rect 2503 9848 2504 9852
rect 2508 9848 2509 9852
rect 2513 9848 2514 9852
rect 2518 9848 2519 9852
rect 2523 9848 2524 9852
rect 2528 9848 2529 9852
rect 2533 9848 2536 9852
rect 2396 9815 2400 9827
rect 2396 9799 2400 9811
rect 2396 9783 2400 9795
rect 2454 9815 2458 9827
rect 2454 9799 2458 9811
rect 2454 9783 2458 9795
rect 2472 9769 2540 9848
rect 2625 9848 2628 9852
rect 2632 9848 2633 9852
rect 2637 9848 2638 9852
rect 2642 9848 2643 9852
rect 2647 9848 2648 9852
rect 2652 9848 2653 9852
rect 2657 9848 2658 9852
rect 2662 9848 2663 9852
rect 2667 9848 2668 9852
rect 2672 9848 2673 9852
rect 2677 9848 2678 9852
rect 2682 9848 2685 9852
rect 2472 9765 2474 9769
rect 2478 9765 2479 9769
rect 2483 9765 2484 9769
rect 2488 9765 2489 9769
rect 2493 9765 2494 9769
rect 2498 9765 2499 9769
rect 2503 9765 2504 9769
rect 2508 9765 2509 9769
rect 2513 9765 2514 9769
rect 2518 9765 2519 9769
rect 2523 9765 2524 9769
rect 2528 9765 2529 9769
rect 2533 9765 2534 9769
rect 2538 9765 2540 9769
rect 2588 9800 2609 9802
rect 2588 9796 2590 9800
rect 2594 9796 2595 9800
rect 2599 9796 2600 9800
rect 2604 9796 2605 9800
rect 2588 9795 2609 9796
rect 2588 9791 2590 9795
rect 2594 9791 2595 9795
rect 2599 9791 2600 9795
rect 2604 9791 2605 9795
rect 2588 9790 2609 9791
rect 2588 9786 2590 9790
rect 2594 9786 2595 9790
rect 2599 9786 2600 9790
rect 2604 9786 2605 9790
rect 2588 9785 2609 9786
rect 2588 9781 2590 9785
rect 2594 9781 2595 9785
rect 2599 9781 2600 9785
rect 2604 9781 2605 9785
rect 2588 9780 2609 9781
rect 2588 9776 2590 9780
rect 2594 9776 2595 9780
rect 2599 9776 2600 9780
rect 2604 9776 2605 9780
rect 2588 9775 2609 9776
rect 2588 9771 2590 9775
rect 2594 9771 2595 9775
rect 2599 9771 2600 9775
rect 2604 9771 2605 9775
rect 2588 9770 2609 9771
rect 2588 9766 2590 9770
rect 2594 9766 2595 9770
rect 2599 9766 2600 9770
rect 2604 9766 2605 9770
rect 2472 9764 2540 9765
rect 2472 9760 2474 9764
rect 2478 9760 2479 9764
rect 2483 9760 2484 9764
rect 2488 9760 2489 9764
rect 2493 9760 2494 9764
rect 2498 9760 2499 9764
rect 2503 9760 2504 9764
rect 2508 9760 2509 9764
rect 2513 9760 2514 9764
rect 2518 9760 2519 9764
rect 2523 9760 2524 9764
rect 2528 9760 2529 9764
rect 2533 9760 2534 9764
rect 2538 9760 2540 9764
rect 2472 9757 2540 9760
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2555 9761 2574 9762
rect 2559 9757 2560 9761
rect 2564 9757 2565 9761
rect 2569 9757 2570 9761
rect 2555 9756 2574 9757
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2555 9751 2574 9752
rect 2559 9747 2560 9751
rect 2564 9747 2565 9751
rect 2569 9747 2570 9751
rect 2555 9746 2574 9747
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2555 9741 2574 9742
rect 2559 9737 2560 9741
rect 2564 9737 2565 9741
rect 2569 9737 2570 9741
rect 2555 9736 2574 9737
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2588 9765 2609 9766
rect 2588 9761 2590 9765
rect 2594 9761 2595 9765
rect 2599 9761 2600 9765
rect 2604 9761 2605 9765
rect 2588 9760 2609 9761
rect 2588 9756 2590 9760
rect 2594 9756 2595 9760
rect 2599 9756 2600 9760
rect 2604 9756 2605 9760
rect 2588 9755 2609 9756
rect 2588 9751 2590 9755
rect 2594 9751 2595 9755
rect 2599 9751 2600 9755
rect 2604 9751 2605 9755
rect 2588 9750 2609 9751
rect 2588 9746 2590 9750
rect 2594 9746 2595 9750
rect 2599 9746 2600 9750
rect 2604 9746 2605 9750
rect 2588 9745 2609 9746
rect 2588 9741 2590 9745
rect 2594 9741 2595 9745
rect 2599 9741 2600 9745
rect 2604 9741 2605 9745
rect 2588 9740 2609 9741
rect 2588 9736 2590 9740
rect 2594 9736 2595 9740
rect 2599 9736 2600 9740
rect 2604 9736 2605 9740
rect 2588 9734 2609 9736
rect 2312 9708 2314 9712
rect 2318 9708 2319 9712
rect 2323 9708 2324 9712
rect 2328 9708 2329 9712
rect 2333 9708 2334 9712
rect 2338 9708 2339 9712
rect 2343 9708 2344 9712
rect 2348 9708 2349 9712
rect 2353 9708 2354 9712
rect 2358 9708 2359 9712
rect 2363 9708 2364 9712
rect 2368 9708 2369 9712
rect 2373 9708 2374 9712
rect 2378 9708 2380 9712
rect 2312 9707 2380 9708
rect 2312 9703 2314 9707
rect 2318 9703 2319 9707
rect 2323 9703 2324 9707
rect 2328 9703 2329 9707
rect 2333 9703 2334 9707
rect 2338 9703 2339 9707
rect 2343 9703 2344 9707
rect 2348 9703 2349 9707
rect 2353 9703 2354 9707
rect 2358 9703 2359 9707
rect 2363 9703 2364 9707
rect 2368 9703 2369 9707
rect 2373 9703 2374 9707
rect 2378 9703 2380 9707
rect 2312 9700 2380 9703
rect 2500 9718 2501 9722
rect 2505 9718 2506 9722
rect 2510 9718 2511 9722
rect 2515 9718 2516 9722
rect 2520 9718 2521 9722
rect 2525 9718 2526 9722
rect 2530 9718 2531 9722
rect 2535 9718 2536 9722
rect 2540 9718 2541 9722
rect 2545 9718 2546 9722
rect 2550 9718 2552 9722
rect 2496 9717 2552 9718
rect 2500 9713 2501 9717
rect 2505 9713 2506 9717
rect 2510 9713 2511 9717
rect 2515 9713 2516 9717
rect 2520 9713 2521 9717
rect 2525 9713 2526 9717
rect 2530 9713 2531 9717
rect 2535 9713 2536 9717
rect 2540 9713 2541 9717
rect 2545 9713 2546 9717
rect 2550 9713 2552 9717
rect 2496 9712 2552 9713
rect 2500 9708 2501 9712
rect 2505 9708 2506 9712
rect 2510 9708 2511 9712
rect 2515 9708 2516 9712
rect 2520 9708 2521 9712
rect 2525 9708 2526 9712
rect 2530 9708 2531 9712
rect 2535 9708 2536 9712
rect 2540 9708 2541 9712
rect 2545 9708 2546 9712
rect 2550 9708 2552 9712
rect 2496 9707 2552 9708
rect 2500 9703 2501 9707
rect 2505 9703 2506 9707
rect 2510 9703 2511 9707
rect 2515 9703 2516 9707
rect 2520 9703 2521 9707
rect 2525 9703 2526 9707
rect 2530 9703 2531 9707
rect 2535 9703 2536 9707
rect 2540 9703 2541 9707
rect 2545 9703 2546 9707
rect 2550 9703 2552 9707
rect 2496 9701 2552 9703
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2555 9715 2574 9716
rect 2559 9711 2560 9715
rect 2564 9711 2565 9715
rect 2569 9711 2570 9715
rect 2555 9710 2574 9711
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2555 9705 2574 9706
rect 2559 9701 2560 9705
rect 2564 9701 2565 9705
rect 2569 9701 2570 9705
rect 2555 9700 2574 9701
rect 2621 9712 2689 9848
rect 2785 9848 2788 9852
rect 2792 9848 2793 9852
rect 2797 9848 2798 9852
rect 2802 9848 2803 9852
rect 2807 9848 2808 9852
rect 2812 9848 2813 9852
rect 2817 9848 2818 9852
rect 2822 9848 2823 9852
rect 2827 9848 2828 9852
rect 2832 9848 2833 9852
rect 2837 9848 2838 9852
rect 2842 9848 2845 9852
rect 2705 9815 2709 9827
rect 2705 9799 2709 9811
rect 2705 9783 2709 9795
rect 2763 9815 2767 9827
rect 2763 9799 2767 9811
rect 2763 9783 2767 9795
rect 2781 9769 2849 9848
rect 2934 9848 2937 9852
rect 2941 9848 2942 9852
rect 2946 9848 2947 9852
rect 2951 9848 2952 9852
rect 2956 9848 2957 9852
rect 2961 9848 2962 9852
rect 2966 9848 2967 9852
rect 2971 9848 2972 9852
rect 2976 9848 2977 9852
rect 2981 9848 2982 9852
rect 2986 9848 2987 9852
rect 2991 9848 2994 9852
rect 2781 9765 2783 9769
rect 2787 9765 2788 9769
rect 2792 9765 2793 9769
rect 2797 9765 2798 9769
rect 2802 9765 2803 9769
rect 2807 9765 2808 9769
rect 2812 9765 2813 9769
rect 2817 9765 2818 9769
rect 2822 9765 2823 9769
rect 2827 9765 2828 9769
rect 2832 9765 2833 9769
rect 2837 9765 2838 9769
rect 2842 9765 2843 9769
rect 2847 9765 2849 9769
rect 2897 9800 2918 9802
rect 2897 9796 2899 9800
rect 2903 9796 2904 9800
rect 2908 9796 2909 9800
rect 2913 9796 2914 9800
rect 2897 9795 2918 9796
rect 2897 9791 2899 9795
rect 2903 9791 2904 9795
rect 2908 9791 2909 9795
rect 2913 9791 2914 9795
rect 2897 9790 2918 9791
rect 2897 9786 2899 9790
rect 2903 9786 2904 9790
rect 2908 9786 2909 9790
rect 2913 9786 2914 9790
rect 2897 9785 2918 9786
rect 2897 9781 2899 9785
rect 2903 9781 2904 9785
rect 2908 9781 2909 9785
rect 2913 9781 2914 9785
rect 2897 9780 2918 9781
rect 2897 9776 2899 9780
rect 2903 9776 2904 9780
rect 2908 9776 2909 9780
rect 2913 9776 2914 9780
rect 2897 9775 2918 9776
rect 2897 9771 2899 9775
rect 2903 9771 2904 9775
rect 2908 9771 2909 9775
rect 2913 9771 2914 9775
rect 2897 9770 2918 9771
rect 2897 9766 2899 9770
rect 2903 9766 2904 9770
rect 2908 9766 2909 9770
rect 2913 9766 2914 9770
rect 2781 9764 2849 9765
rect 2781 9760 2783 9764
rect 2787 9760 2788 9764
rect 2792 9760 2793 9764
rect 2797 9760 2798 9764
rect 2802 9760 2803 9764
rect 2807 9760 2808 9764
rect 2812 9760 2813 9764
rect 2817 9760 2818 9764
rect 2822 9760 2823 9764
rect 2827 9760 2828 9764
rect 2832 9760 2833 9764
rect 2837 9760 2838 9764
rect 2842 9760 2843 9764
rect 2847 9760 2849 9764
rect 2781 9757 2849 9760
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2864 9761 2883 9762
rect 2868 9757 2869 9761
rect 2873 9757 2874 9761
rect 2878 9757 2879 9761
rect 2864 9756 2883 9757
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2864 9751 2883 9752
rect 2868 9747 2869 9751
rect 2873 9747 2874 9751
rect 2878 9747 2879 9751
rect 2864 9746 2883 9747
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2864 9741 2883 9742
rect 2868 9737 2869 9741
rect 2873 9737 2874 9741
rect 2878 9737 2879 9741
rect 2864 9736 2883 9737
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2897 9765 2918 9766
rect 2897 9761 2899 9765
rect 2903 9761 2904 9765
rect 2908 9761 2909 9765
rect 2913 9761 2914 9765
rect 2897 9760 2918 9761
rect 2897 9756 2899 9760
rect 2903 9756 2904 9760
rect 2908 9756 2909 9760
rect 2913 9756 2914 9760
rect 2897 9755 2918 9756
rect 2897 9751 2899 9755
rect 2903 9751 2904 9755
rect 2908 9751 2909 9755
rect 2913 9751 2914 9755
rect 2897 9750 2918 9751
rect 2897 9746 2899 9750
rect 2903 9746 2904 9750
rect 2908 9746 2909 9750
rect 2913 9746 2914 9750
rect 2897 9745 2918 9746
rect 2897 9741 2899 9745
rect 2903 9741 2904 9745
rect 2908 9741 2909 9745
rect 2913 9741 2914 9745
rect 2897 9740 2918 9741
rect 2897 9736 2899 9740
rect 2903 9736 2904 9740
rect 2908 9736 2909 9740
rect 2913 9736 2914 9740
rect 2897 9734 2918 9736
rect 2621 9708 2623 9712
rect 2627 9708 2628 9712
rect 2632 9708 2633 9712
rect 2637 9708 2638 9712
rect 2642 9708 2643 9712
rect 2647 9708 2648 9712
rect 2652 9708 2653 9712
rect 2657 9708 2658 9712
rect 2662 9708 2663 9712
rect 2667 9708 2668 9712
rect 2672 9708 2673 9712
rect 2677 9708 2678 9712
rect 2682 9708 2683 9712
rect 2687 9708 2689 9712
rect 2621 9707 2689 9708
rect 2621 9703 2623 9707
rect 2627 9703 2628 9707
rect 2632 9703 2633 9707
rect 2637 9703 2638 9707
rect 2642 9703 2643 9707
rect 2647 9703 2648 9707
rect 2652 9703 2653 9707
rect 2657 9703 2658 9707
rect 2662 9703 2663 9707
rect 2667 9703 2668 9707
rect 2672 9703 2673 9707
rect 2677 9703 2678 9707
rect 2682 9703 2683 9707
rect 2687 9703 2689 9707
rect 2621 9700 2689 9703
rect 2809 9718 2810 9722
rect 2814 9718 2815 9722
rect 2819 9718 2820 9722
rect 2824 9718 2825 9722
rect 2829 9718 2830 9722
rect 2834 9718 2835 9722
rect 2839 9718 2840 9722
rect 2844 9718 2845 9722
rect 2849 9718 2850 9722
rect 2854 9718 2855 9722
rect 2859 9718 2861 9722
rect 2805 9717 2861 9718
rect 2809 9713 2810 9717
rect 2814 9713 2815 9717
rect 2819 9713 2820 9717
rect 2824 9713 2825 9717
rect 2829 9713 2830 9717
rect 2834 9713 2835 9717
rect 2839 9713 2840 9717
rect 2844 9713 2845 9717
rect 2849 9713 2850 9717
rect 2854 9713 2855 9717
rect 2859 9713 2861 9717
rect 2805 9712 2861 9713
rect 2809 9708 2810 9712
rect 2814 9708 2815 9712
rect 2819 9708 2820 9712
rect 2824 9708 2825 9712
rect 2829 9708 2830 9712
rect 2834 9708 2835 9712
rect 2839 9708 2840 9712
rect 2844 9708 2845 9712
rect 2849 9708 2850 9712
rect 2854 9708 2855 9712
rect 2859 9708 2861 9712
rect 2805 9707 2861 9708
rect 2809 9703 2810 9707
rect 2814 9703 2815 9707
rect 2819 9703 2820 9707
rect 2824 9703 2825 9707
rect 2829 9703 2830 9707
rect 2834 9703 2835 9707
rect 2839 9703 2840 9707
rect 2844 9703 2845 9707
rect 2849 9703 2850 9707
rect 2854 9703 2855 9707
rect 2859 9703 2861 9707
rect 2805 9701 2861 9703
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2864 9715 2883 9716
rect 2868 9711 2869 9715
rect 2873 9711 2874 9715
rect 2878 9711 2879 9715
rect 2864 9710 2883 9711
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2864 9705 2883 9706
rect 2868 9701 2869 9705
rect 2873 9701 2874 9705
rect 2878 9701 2879 9705
rect 2864 9700 2883 9701
rect 2930 9712 2998 9848
rect 3094 9848 3097 9852
rect 3101 9848 3102 9852
rect 3106 9848 3107 9852
rect 3111 9848 3112 9852
rect 3116 9848 3117 9852
rect 3121 9848 3122 9852
rect 3126 9848 3127 9852
rect 3131 9848 3132 9852
rect 3136 9848 3137 9852
rect 3141 9848 3142 9852
rect 3146 9848 3147 9852
rect 3151 9848 3154 9852
rect 3014 9815 3018 9827
rect 3014 9799 3018 9811
rect 3014 9783 3018 9795
rect 3072 9815 3076 9827
rect 3072 9799 3076 9811
rect 3072 9783 3076 9795
rect 3090 9769 3158 9848
rect 3243 9848 3246 9852
rect 3250 9848 3251 9852
rect 3255 9848 3256 9852
rect 3260 9848 3261 9852
rect 3265 9848 3266 9852
rect 3270 9848 3271 9852
rect 3275 9848 3276 9852
rect 3280 9848 3281 9852
rect 3285 9848 3286 9852
rect 3290 9848 3291 9852
rect 3295 9848 3296 9852
rect 3300 9848 3303 9852
rect 3090 9765 3092 9769
rect 3096 9765 3097 9769
rect 3101 9765 3102 9769
rect 3106 9765 3107 9769
rect 3111 9765 3112 9769
rect 3116 9765 3117 9769
rect 3121 9765 3122 9769
rect 3126 9765 3127 9769
rect 3131 9765 3132 9769
rect 3136 9765 3137 9769
rect 3141 9765 3142 9769
rect 3146 9765 3147 9769
rect 3151 9765 3152 9769
rect 3156 9765 3158 9769
rect 3206 9800 3227 9802
rect 3206 9796 3208 9800
rect 3212 9796 3213 9800
rect 3217 9796 3218 9800
rect 3222 9796 3223 9800
rect 3206 9795 3227 9796
rect 3206 9791 3208 9795
rect 3212 9791 3213 9795
rect 3217 9791 3218 9795
rect 3222 9791 3223 9795
rect 3206 9790 3227 9791
rect 3206 9786 3208 9790
rect 3212 9786 3213 9790
rect 3217 9786 3218 9790
rect 3222 9786 3223 9790
rect 3206 9785 3227 9786
rect 3206 9781 3208 9785
rect 3212 9781 3213 9785
rect 3217 9781 3218 9785
rect 3222 9781 3223 9785
rect 3206 9780 3227 9781
rect 3206 9776 3208 9780
rect 3212 9776 3213 9780
rect 3217 9776 3218 9780
rect 3222 9776 3223 9780
rect 3206 9775 3227 9776
rect 3206 9771 3208 9775
rect 3212 9771 3213 9775
rect 3217 9771 3218 9775
rect 3222 9771 3223 9775
rect 3206 9770 3227 9771
rect 3206 9766 3208 9770
rect 3212 9766 3213 9770
rect 3217 9766 3218 9770
rect 3222 9766 3223 9770
rect 3090 9764 3158 9765
rect 3090 9760 3092 9764
rect 3096 9760 3097 9764
rect 3101 9760 3102 9764
rect 3106 9760 3107 9764
rect 3111 9760 3112 9764
rect 3116 9760 3117 9764
rect 3121 9760 3122 9764
rect 3126 9760 3127 9764
rect 3131 9760 3132 9764
rect 3136 9760 3137 9764
rect 3141 9760 3142 9764
rect 3146 9760 3147 9764
rect 3151 9760 3152 9764
rect 3156 9760 3158 9764
rect 3090 9757 3158 9760
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3173 9761 3192 9762
rect 3177 9757 3178 9761
rect 3182 9757 3183 9761
rect 3187 9757 3188 9761
rect 3173 9756 3192 9757
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3173 9751 3192 9752
rect 3177 9747 3178 9751
rect 3182 9747 3183 9751
rect 3187 9747 3188 9751
rect 3173 9746 3192 9747
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3173 9741 3192 9742
rect 3177 9737 3178 9741
rect 3182 9737 3183 9741
rect 3187 9737 3188 9741
rect 3173 9736 3192 9737
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3206 9765 3227 9766
rect 3206 9761 3208 9765
rect 3212 9761 3213 9765
rect 3217 9761 3218 9765
rect 3222 9761 3223 9765
rect 3206 9760 3227 9761
rect 3206 9756 3208 9760
rect 3212 9756 3213 9760
rect 3217 9756 3218 9760
rect 3222 9756 3223 9760
rect 3206 9755 3227 9756
rect 3206 9751 3208 9755
rect 3212 9751 3213 9755
rect 3217 9751 3218 9755
rect 3222 9751 3223 9755
rect 3206 9750 3227 9751
rect 3206 9746 3208 9750
rect 3212 9746 3213 9750
rect 3217 9746 3218 9750
rect 3222 9746 3223 9750
rect 3206 9745 3227 9746
rect 3206 9741 3208 9745
rect 3212 9741 3213 9745
rect 3217 9741 3218 9745
rect 3222 9741 3223 9745
rect 3206 9740 3227 9741
rect 3206 9736 3208 9740
rect 3212 9736 3213 9740
rect 3217 9736 3218 9740
rect 3222 9736 3223 9740
rect 3206 9734 3227 9736
rect 2930 9708 2932 9712
rect 2936 9708 2937 9712
rect 2941 9708 2942 9712
rect 2946 9708 2947 9712
rect 2951 9708 2952 9712
rect 2956 9708 2957 9712
rect 2961 9708 2962 9712
rect 2966 9708 2967 9712
rect 2971 9708 2972 9712
rect 2976 9708 2977 9712
rect 2981 9708 2982 9712
rect 2986 9708 2987 9712
rect 2991 9708 2992 9712
rect 2996 9708 2998 9712
rect 2930 9707 2998 9708
rect 2930 9703 2932 9707
rect 2936 9703 2937 9707
rect 2941 9703 2942 9707
rect 2946 9703 2947 9707
rect 2951 9703 2952 9707
rect 2956 9703 2957 9707
rect 2961 9703 2962 9707
rect 2966 9703 2967 9707
rect 2971 9703 2972 9707
rect 2976 9703 2977 9707
rect 2981 9703 2982 9707
rect 2986 9703 2987 9707
rect 2991 9703 2992 9707
rect 2996 9703 2998 9707
rect 2930 9700 2998 9703
rect 3118 9718 3119 9722
rect 3123 9718 3124 9722
rect 3128 9718 3129 9722
rect 3133 9718 3134 9722
rect 3138 9718 3139 9722
rect 3143 9718 3144 9722
rect 3148 9718 3149 9722
rect 3153 9718 3154 9722
rect 3158 9718 3159 9722
rect 3163 9718 3164 9722
rect 3168 9718 3170 9722
rect 3114 9717 3170 9718
rect 3118 9713 3119 9717
rect 3123 9713 3124 9717
rect 3128 9713 3129 9717
rect 3133 9713 3134 9717
rect 3138 9713 3139 9717
rect 3143 9713 3144 9717
rect 3148 9713 3149 9717
rect 3153 9713 3154 9717
rect 3158 9713 3159 9717
rect 3163 9713 3164 9717
rect 3168 9713 3170 9717
rect 3114 9712 3170 9713
rect 3118 9708 3119 9712
rect 3123 9708 3124 9712
rect 3128 9708 3129 9712
rect 3133 9708 3134 9712
rect 3138 9708 3139 9712
rect 3143 9708 3144 9712
rect 3148 9708 3149 9712
rect 3153 9708 3154 9712
rect 3158 9708 3159 9712
rect 3163 9708 3164 9712
rect 3168 9708 3170 9712
rect 3114 9707 3170 9708
rect 3118 9703 3119 9707
rect 3123 9703 3124 9707
rect 3128 9703 3129 9707
rect 3133 9703 3134 9707
rect 3138 9703 3139 9707
rect 3143 9703 3144 9707
rect 3148 9703 3149 9707
rect 3153 9703 3154 9707
rect 3158 9703 3159 9707
rect 3163 9703 3164 9707
rect 3168 9703 3170 9707
rect 3114 9701 3170 9703
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3173 9715 3192 9716
rect 3177 9711 3178 9715
rect 3182 9711 3183 9715
rect 3187 9711 3188 9715
rect 3173 9710 3192 9711
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3173 9705 3192 9706
rect 3177 9701 3178 9705
rect 3182 9701 3183 9705
rect 3187 9701 3188 9705
rect 3173 9700 3192 9701
rect 3239 9712 3307 9848
rect 3403 9848 3406 9852
rect 3410 9848 3411 9852
rect 3415 9848 3416 9852
rect 3420 9848 3421 9852
rect 3425 9848 3426 9852
rect 3430 9848 3431 9852
rect 3435 9848 3436 9852
rect 3440 9848 3441 9852
rect 3445 9848 3446 9852
rect 3450 9848 3451 9852
rect 3455 9848 3456 9852
rect 3460 9848 3463 9852
rect 3399 9769 3467 9848
rect 3552 9848 3555 9852
rect 3559 9848 3560 9852
rect 3564 9848 3565 9852
rect 3569 9848 3570 9852
rect 3574 9848 3575 9852
rect 3579 9848 3580 9852
rect 3584 9848 3585 9852
rect 3589 9848 3590 9852
rect 3594 9848 3595 9852
rect 3599 9848 3600 9852
rect 3604 9848 3605 9852
rect 3609 9848 3612 9852
rect 3399 9765 3401 9769
rect 3405 9765 3406 9769
rect 3410 9765 3411 9769
rect 3415 9765 3416 9769
rect 3420 9765 3421 9769
rect 3425 9765 3426 9769
rect 3430 9765 3431 9769
rect 3435 9765 3436 9769
rect 3440 9765 3441 9769
rect 3445 9765 3446 9769
rect 3450 9765 3451 9769
rect 3455 9765 3456 9769
rect 3460 9765 3461 9769
rect 3465 9765 3467 9769
rect 3515 9800 3536 9802
rect 3515 9796 3517 9800
rect 3521 9796 3522 9800
rect 3526 9796 3527 9800
rect 3531 9796 3532 9800
rect 3515 9795 3536 9796
rect 3515 9791 3517 9795
rect 3521 9791 3522 9795
rect 3526 9791 3527 9795
rect 3531 9791 3532 9795
rect 3515 9790 3536 9791
rect 3515 9786 3517 9790
rect 3521 9786 3522 9790
rect 3526 9786 3527 9790
rect 3531 9786 3532 9790
rect 3515 9785 3536 9786
rect 3515 9781 3517 9785
rect 3521 9781 3522 9785
rect 3526 9781 3527 9785
rect 3531 9781 3532 9785
rect 3515 9780 3536 9781
rect 3515 9776 3517 9780
rect 3521 9776 3522 9780
rect 3526 9776 3527 9780
rect 3531 9776 3532 9780
rect 3515 9775 3536 9776
rect 3515 9771 3517 9775
rect 3521 9771 3522 9775
rect 3526 9771 3527 9775
rect 3531 9771 3532 9775
rect 3515 9770 3536 9771
rect 3515 9766 3517 9770
rect 3521 9766 3522 9770
rect 3526 9766 3527 9770
rect 3531 9766 3532 9770
rect 3399 9764 3467 9765
rect 3399 9760 3401 9764
rect 3405 9760 3406 9764
rect 3410 9760 3411 9764
rect 3415 9760 3416 9764
rect 3420 9760 3421 9764
rect 3425 9760 3426 9764
rect 3430 9760 3431 9764
rect 3435 9760 3436 9764
rect 3440 9760 3441 9764
rect 3445 9760 3446 9764
rect 3450 9760 3451 9764
rect 3455 9760 3456 9764
rect 3460 9760 3461 9764
rect 3465 9760 3467 9764
rect 3399 9757 3467 9760
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3482 9761 3501 9762
rect 3486 9757 3487 9761
rect 3491 9757 3492 9761
rect 3496 9757 3497 9761
rect 3482 9756 3501 9757
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3482 9751 3501 9752
rect 3486 9747 3487 9751
rect 3491 9747 3492 9751
rect 3496 9747 3497 9751
rect 3482 9746 3501 9747
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3482 9741 3501 9742
rect 3486 9737 3487 9741
rect 3491 9737 3492 9741
rect 3496 9737 3497 9741
rect 3482 9736 3501 9737
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3515 9765 3536 9766
rect 3515 9761 3517 9765
rect 3521 9761 3522 9765
rect 3526 9761 3527 9765
rect 3531 9761 3532 9765
rect 3515 9760 3536 9761
rect 3515 9756 3517 9760
rect 3521 9756 3522 9760
rect 3526 9756 3527 9760
rect 3531 9756 3532 9760
rect 3515 9755 3536 9756
rect 3515 9751 3517 9755
rect 3521 9751 3522 9755
rect 3526 9751 3527 9755
rect 3531 9751 3532 9755
rect 3515 9750 3536 9751
rect 3515 9746 3517 9750
rect 3521 9746 3522 9750
rect 3526 9746 3527 9750
rect 3531 9746 3532 9750
rect 3515 9745 3536 9746
rect 3515 9741 3517 9745
rect 3521 9741 3522 9745
rect 3526 9741 3527 9745
rect 3531 9741 3532 9745
rect 3515 9740 3536 9741
rect 3515 9736 3517 9740
rect 3521 9736 3522 9740
rect 3526 9736 3527 9740
rect 3531 9736 3532 9740
rect 3515 9734 3536 9736
rect 3427 9718 3428 9722
rect 3432 9718 3433 9722
rect 3437 9718 3438 9722
rect 3442 9718 3443 9722
rect 3447 9718 3448 9722
rect 3452 9718 3453 9722
rect 3457 9718 3458 9722
rect 3462 9718 3463 9722
rect 3467 9718 3468 9722
rect 3472 9718 3473 9722
rect 3477 9718 3479 9722
rect 3423 9717 3479 9718
rect 3239 9708 3241 9712
rect 3245 9708 3246 9712
rect 3250 9708 3251 9712
rect 3255 9708 3256 9712
rect 3260 9708 3261 9712
rect 3265 9708 3266 9712
rect 3270 9708 3271 9712
rect 3275 9708 3276 9712
rect 3280 9708 3281 9712
rect 3285 9708 3286 9712
rect 3290 9708 3291 9712
rect 3295 9708 3296 9712
rect 3300 9708 3301 9712
rect 3305 9708 3307 9712
rect 3239 9707 3307 9708
rect 3239 9703 3241 9707
rect 3245 9703 3246 9707
rect 3250 9703 3251 9707
rect 3255 9703 3256 9707
rect 3260 9703 3261 9707
rect 3265 9703 3266 9707
rect 3270 9703 3271 9707
rect 3275 9703 3276 9707
rect 3280 9703 3281 9707
rect 3285 9703 3286 9707
rect 3290 9703 3291 9707
rect 3295 9703 3296 9707
rect 3300 9703 3301 9707
rect 3305 9703 3307 9707
rect 3239 9700 3307 9703
rect 3342 9711 3343 9715
rect 3347 9711 3348 9715
rect 3352 9711 3353 9715
rect 3357 9711 3358 9715
rect 3342 9710 3362 9711
rect 3342 9706 3343 9710
rect 3347 9706 3348 9710
rect 3352 9706 3353 9710
rect 3357 9706 3358 9710
rect 3342 9705 3362 9706
rect 3342 9701 3343 9705
rect 3347 9701 3348 9705
rect 3352 9701 3353 9705
rect 3357 9701 3358 9705
rect 3427 9713 3428 9717
rect 3432 9713 3433 9717
rect 3437 9713 3438 9717
rect 3442 9713 3443 9717
rect 3447 9713 3448 9717
rect 3452 9713 3453 9717
rect 3457 9713 3458 9717
rect 3462 9713 3463 9717
rect 3467 9713 3468 9717
rect 3472 9713 3473 9717
rect 3477 9713 3479 9717
rect 3423 9712 3479 9713
rect 3427 9708 3428 9712
rect 3432 9708 3433 9712
rect 3437 9708 3438 9712
rect 3442 9708 3443 9712
rect 3447 9708 3448 9712
rect 3452 9708 3453 9712
rect 3457 9708 3458 9712
rect 3462 9708 3463 9712
rect 3467 9708 3468 9712
rect 3472 9708 3473 9712
rect 3477 9708 3479 9712
rect 3423 9707 3479 9708
rect 3427 9703 3428 9707
rect 3432 9703 3433 9707
rect 3437 9703 3438 9707
rect 3442 9703 3443 9707
rect 3447 9703 3448 9707
rect 3452 9703 3453 9707
rect 3457 9703 3458 9707
rect 3462 9703 3463 9707
rect 3467 9703 3468 9707
rect 3472 9703 3473 9707
rect 3477 9703 3479 9707
rect 3423 9701 3479 9703
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3482 9715 3501 9716
rect 3486 9711 3487 9715
rect 3491 9711 3492 9715
rect 3496 9711 3497 9715
rect 3482 9710 3501 9711
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3482 9705 3501 9706
rect 3486 9701 3487 9705
rect 3491 9701 3492 9705
rect 3496 9701 3497 9705
rect 3342 9700 3362 9701
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2246 9695 2265 9696
rect 2250 9691 2251 9695
rect 2255 9691 2256 9695
rect 2260 9691 2261 9695
rect 2246 9690 2265 9691
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2555 9695 2574 9696
rect 2559 9691 2560 9695
rect 2564 9691 2565 9695
rect 2569 9691 2570 9695
rect 2555 9690 2574 9691
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2864 9695 2883 9696
rect 2868 9691 2869 9695
rect 2873 9691 2874 9695
rect 2878 9691 2879 9695
rect 2864 9690 2883 9691
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3173 9695 3192 9696
rect 3177 9691 3178 9695
rect 3182 9691 3183 9695
rect 3187 9691 3188 9695
rect 3173 9690 3192 9691
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3342 9696 3343 9700
rect 3347 9696 3348 9700
rect 3352 9696 3353 9700
rect 3357 9696 3358 9700
rect 3342 9695 3362 9696
rect 3342 9691 3343 9695
rect 3347 9691 3348 9695
rect 3352 9691 3353 9695
rect 3357 9691 3358 9695
rect 3342 9690 3362 9691
rect 3342 9686 3343 9690
rect 3347 9686 3348 9690
rect 3352 9686 3353 9690
rect 3357 9686 3358 9690
rect 3482 9700 3501 9701
rect 3548 9712 3616 9848
rect 3712 9848 3715 9852
rect 3719 9848 3720 9852
rect 3724 9848 3725 9852
rect 3729 9848 3730 9852
rect 3734 9848 3735 9852
rect 3739 9848 3740 9852
rect 3744 9848 3745 9852
rect 3749 9848 3750 9852
rect 3754 9848 3755 9852
rect 3759 9848 3760 9852
rect 3764 9848 3765 9852
rect 3769 9848 3772 9852
rect 3651 9791 3652 9795
rect 3656 9791 3657 9795
rect 3661 9791 3662 9795
rect 3666 9791 3667 9795
rect 3651 9790 3671 9791
rect 3651 9786 3652 9790
rect 3656 9786 3657 9790
rect 3661 9786 3662 9790
rect 3666 9786 3667 9790
rect 3651 9785 3671 9786
rect 3651 9781 3652 9785
rect 3656 9781 3657 9785
rect 3661 9781 3662 9785
rect 3666 9781 3667 9785
rect 3651 9780 3671 9781
rect 3651 9776 3652 9780
rect 3656 9776 3657 9780
rect 3661 9776 3662 9780
rect 3666 9776 3667 9780
rect 3651 9775 3671 9776
rect 3651 9771 3652 9775
rect 3656 9771 3657 9775
rect 3661 9771 3662 9775
rect 3666 9771 3667 9775
rect 3651 9770 3671 9771
rect 3651 9766 3652 9770
rect 3656 9766 3657 9770
rect 3661 9766 3662 9770
rect 3666 9766 3667 9770
rect 3651 9765 3671 9766
rect 3651 9761 3652 9765
rect 3656 9761 3657 9765
rect 3661 9761 3662 9765
rect 3666 9761 3667 9765
rect 3651 9760 3671 9761
rect 3651 9756 3652 9760
rect 3656 9756 3657 9760
rect 3661 9756 3662 9760
rect 3666 9756 3667 9760
rect 3708 9769 3776 9848
rect 3861 9848 3864 9852
rect 3868 9848 3869 9852
rect 3873 9848 3874 9852
rect 3878 9848 3879 9852
rect 3883 9848 3884 9852
rect 3888 9848 3889 9852
rect 3893 9848 3894 9852
rect 3898 9848 3899 9852
rect 3903 9848 3904 9852
rect 3908 9848 3909 9852
rect 3913 9848 3914 9852
rect 3918 9848 3921 9852
rect 3708 9765 3710 9769
rect 3714 9765 3715 9769
rect 3719 9765 3720 9769
rect 3724 9765 3725 9769
rect 3729 9765 3730 9769
rect 3734 9765 3735 9769
rect 3739 9765 3740 9769
rect 3744 9765 3745 9769
rect 3749 9765 3750 9769
rect 3754 9765 3755 9769
rect 3759 9765 3760 9769
rect 3764 9765 3765 9769
rect 3769 9765 3770 9769
rect 3774 9765 3776 9769
rect 3824 9800 3845 9802
rect 3824 9796 3826 9800
rect 3830 9796 3831 9800
rect 3835 9796 3836 9800
rect 3840 9796 3841 9800
rect 3824 9795 3845 9796
rect 3824 9791 3826 9795
rect 3830 9791 3831 9795
rect 3835 9791 3836 9795
rect 3840 9791 3841 9795
rect 3824 9790 3845 9791
rect 3824 9786 3826 9790
rect 3830 9786 3831 9790
rect 3835 9786 3836 9790
rect 3840 9786 3841 9790
rect 3824 9785 3845 9786
rect 3824 9781 3826 9785
rect 3830 9781 3831 9785
rect 3835 9781 3836 9785
rect 3840 9781 3841 9785
rect 3824 9780 3845 9781
rect 3824 9776 3826 9780
rect 3830 9776 3831 9780
rect 3835 9776 3836 9780
rect 3840 9776 3841 9780
rect 3824 9775 3845 9776
rect 3824 9771 3826 9775
rect 3830 9771 3831 9775
rect 3835 9771 3836 9775
rect 3840 9771 3841 9775
rect 3824 9770 3845 9771
rect 3824 9766 3826 9770
rect 3830 9766 3831 9770
rect 3835 9766 3836 9770
rect 3840 9766 3841 9770
rect 3708 9764 3776 9765
rect 3708 9760 3710 9764
rect 3714 9760 3715 9764
rect 3719 9760 3720 9764
rect 3724 9760 3725 9764
rect 3729 9760 3730 9764
rect 3734 9760 3735 9764
rect 3739 9760 3740 9764
rect 3744 9760 3745 9764
rect 3749 9760 3750 9764
rect 3754 9760 3755 9764
rect 3759 9760 3760 9764
rect 3764 9760 3765 9764
rect 3769 9760 3770 9764
rect 3774 9760 3776 9764
rect 3708 9757 3776 9760
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3791 9761 3810 9762
rect 3795 9757 3796 9761
rect 3800 9757 3801 9761
rect 3805 9757 3806 9761
rect 3651 9755 3671 9756
rect 3651 9751 3652 9755
rect 3656 9751 3657 9755
rect 3661 9751 3662 9755
rect 3666 9751 3667 9755
rect 3651 9750 3671 9751
rect 3651 9746 3652 9750
rect 3656 9746 3657 9750
rect 3661 9746 3662 9750
rect 3666 9746 3667 9750
rect 3651 9745 3671 9746
rect 3651 9741 3652 9745
rect 3656 9741 3657 9745
rect 3661 9741 3662 9745
rect 3666 9741 3667 9745
rect 3651 9739 3671 9741
rect 3791 9756 3810 9757
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3791 9751 3810 9752
rect 3795 9747 3796 9751
rect 3800 9747 3801 9751
rect 3805 9747 3806 9751
rect 3791 9746 3810 9747
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3791 9741 3810 9742
rect 3795 9737 3796 9741
rect 3800 9737 3801 9741
rect 3805 9737 3806 9741
rect 3791 9736 3810 9737
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3824 9765 3845 9766
rect 3824 9761 3826 9765
rect 3830 9761 3831 9765
rect 3835 9761 3836 9765
rect 3840 9761 3841 9765
rect 3824 9760 3845 9761
rect 3824 9756 3826 9760
rect 3830 9756 3831 9760
rect 3835 9756 3836 9760
rect 3840 9756 3841 9760
rect 3824 9755 3845 9756
rect 3824 9751 3826 9755
rect 3830 9751 3831 9755
rect 3835 9751 3836 9755
rect 3840 9751 3841 9755
rect 3824 9750 3845 9751
rect 3824 9746 3826 9750
rect 3830 9746 3831 9750
rect 3835 9746 3836 9750
rect 3840 9746 3841 9750
rect 3824 9745 3845 9746
rect 3824 9741 3826 9745
rect 3830 9741 3831 9745
rect 3835 9741 3836 9745
rect 3840 9741 3841 9745
rect 3824 9740 3845 9741
rect 3824 9736 3826 9740
rect 3830 9736 3831 9740
rect 3835 9736 3836 9740
rect 3840 9736 3841 9740
rect 3824 9734 3845 9736
rect 3548 9708 3550 9712
rect 3554 9708 3555 9712
rect 3559 9708 3560 9712
rect 3564 9708 3565 9712
rect 3569 9708 3570 9712
rect 3574 9708 3575 9712
rect 3579 9708 3580 9712
rect 3584 9708 3585 9712
rect 3589 9708 3590 9712
rect 3594 9708 3595 9712
rect 3599 9708 3600 9712
rect 3604 9708 3605 9712
rect 3609 9708 3610 9712
rect 3614 9708 3616 9712
rect 3548 9707 3616 9708
rect 3548 9703 3550 9707
rect 3554 9703 3555 9707
rect 3559 9703 3560 9707
rect 3564 9703 3565 9707
rect 3569 9703 3570 9707
rect 3574 9703 3575 9707
rect 3579 9703 3580 9707
rect 3584 9703 3585 9707
rect 3589 9703 3590 9707
rect 3594 9703 3595 9707
rect 3599 9703 3600 9707
rect 3604 9703 3605 9707
rect 3609 9703 3610 9707
rect 3614 9703 3616 9707
rect 3548 9700 3616 9703
rect 3736 9718 3737 9722
rect 3741 9718 3742 9722
rect 3746 9718 3747 9722
rect 3751 9718 3752 9722
rect 3756 9718 3757 9722
rect 3761 9718 3762 9722
rect 3766 9718 3767 9722
rect 3771 9718 3772 9722
rect 3776 9718 3777 9722
rect 3781 9718 3782 9722
rect 3786 9718 3788 9722
rect 3732 9717 3788 9718
rect 3736 9713 3737 9717
rect 3741 9713 3742 9717
rect 3746 9713 3747 9717
rect 3751 9713 3752 9717
rect 3756 9713 3757 9717
rect 3761 9713 3762 9717
rect 3766 9713 3767 9717
rect 3771 9713 3772 9717
rect 3776 9713 3777 9717
rect 3781 9713 3782 9717
rect 3786 9713 3788 9717
rect 3732 9712 3788 9713
rect 3736 9708 3737 9712
rect 3741 9708 3742 9712
rect 3746 9708 3747 9712
rect 3751 9708 3752 9712
rect 3756 9708 3757 9712
rect 3761 9708 3762 9712
rect 3766 9708 3767 9712
rect 3771 9708 3772 9712
rect 3776 9708 3777 9712
rect 3781 9708 3782 9712
rect 3786 9708 3788 9712
rect 3732 9707 3788 9708
rect 3736 9703 3737 9707
rect 3741 9703 3742 9707
rect 3746 9703 3747 9707
rect 3751 9703 3752 9707
rect 3756 9703 3757 9707
rect 3761 9703 3762 9707
rect 3766 9703 3767 9707
rect 3771 9703 3772 9707
rect 3776 9703 3777 9707
rect 3781 9703 3782 9707
rect 3786 9703 3788 9707
rect 3732 9701 3788 9703
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3791 9715 3810 9716
rect 3795 9711 3796 9715
rect 3800 9711 3801 9715
rect 3805 9711 3806 9715
rect 3791 9710 3810 9711
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3791 9705 3810 9706
rect 3795 9701 3796 9705
rect 3800 9701 3801 9705
rect 3805 9701 3806 9705
rect 3791 9700 3810 9701
rect 3857 9712 3925 9848
rect 4021 9848 4024 9852
rect 4028 9848 4029 9852
rect 4033 9848 4034 9852
rect 4038 9848 4039 9852
rect 4043 9848 4044 9852
rect 4048 9848 4049 9852
rect 4053 9848 4054 9852
rect 4058 9848 4059 9852
rect 4063 9848 4064 9852
rect 4068 9848 4069 9852
rect 4073 9848 4074 9852
rect 4078 9848 4081 9852
rect 3941 9815 3945 9827
rect 3941 9799 3945 9811
rect 3941 9783 3945 9795
rect 3999 9815 4003 9827
rect 3999 9799 4003 9811
rect 3999 9783 4003 9795
rect 4017 9769 4085 9848
rect 4141 9786 5073 10261
rect 4017 9765 4019 9769
rect 4023 9765 4024 9769
rect 4028 9765 4029 9769
rect 4033 9765 4034 9769
rect 4038 9765 4039 9769
rect 4043 9765 4044 9769
rect 4048 9765 4049 9769
rect 4053 9765 4054 9769
rect 4058 9765 4059 9769
rect 4063 9765 4064 9769
rect 4068 9765 4069 9769
rect 4073 9765 4074 9769
rect 4078 9765 4079 9769
rect 4083 9765 4085 9769
rect 4017 9764 4085 9765
rect 4017 9760 4019 9764
rect 4023 9760 4024 9764
rect 4028 9760 4029 9764
rect 4033 9760 4034 9764
rect 4038 9760 4039 9764
rect 4043 9760 4044 9764
rect 4048 9760 4049 9764
rect 4053 9760 4054 9764
rect 4058 9760 4059 9764
rect 4063 9760 4064 9764
rect 4068 9760 4069 9764
rect 4073 9760 4074 9764
rect 4078 9760 4079 9764
rect 4083 9760 4085 9764
rect 4017 9757 4085 9760
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4100 9761 4119 9762
rect 4104 9757 4105 9761
rect 4109 9757 4110 9761
rect 4114 9757 4115 9761
rect 4100 9756 4119 9757
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4100 9751 4119 9752
rect 4104 9747 4105 9751
rect 4109 9747 4110 9751
rect 4114 9747 4115 9751
rect 4100 9746 4119 9747
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4100 9741 4119 9742
rect 4104 9737 4105 9741
rect 4109 9737 4110 9741
rect 4114 9737 4115 9741
rect 4100 9736 4119 9737
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4292 9761 4311 9762
rect 4296 9757 4297 9761
rect 4301 9757 4302 9761
rect 4306 9757 4307 9761
rect 4292 9756 4311 9757
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4292 9751 4311 9752
rect 4296 9747 4297 9751
rect 4301 9747 4302 9751
rect 4306 9747 4307 9751
rect 4292 9746 4311 9747
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4292 9741 4311 9742
rect 4296 9737 4297 9741
rect 4301 9737 4302 9741
rect 4306 9737 4307 9741
rect 4292 9736 4311 9737
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4318 9761 4337 9762
rect 4322 9757 4323 9761
rect 4327 9757 4328 9761
rect 4332 9757 4333 9761
rect 4318 9756 4337 9757
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4318 9751 4337 9752
rect 4322 9747 4323 9751
rect 4327 9747 4328 9751
rect 4332 9747 4333 9751
rect 4318 9746 4337 9747
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4318 9741 4337 9742
rect 4322 9737 4323 9741
rect 4327 9737 4328 9741
rect 4332 9737 4333 9741
rect 4318 9736 4337 9737
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4344 9761 4363 9762
rect 4348 9757 4349 9761
rect 4353 9757 4354 9761
rect 4358 9757 4359 9761
rect 4344 9756 4363 9757
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4344 9751 4363 9752
rect 4348 9747 4349 9751
rect 4353 9747 4354 9751
rect 4358 9747 4359 9751
rect 4344 9746 4363 9747
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4344 9741 4363 9742
rect 4348 9737 4349 9741
rect 4353 9737 4354 9741
rect 4358 9737 4359 9741
rect 4344 9736 4363 9737
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4370 9761 4389 9762
rect 4374 9757 4375 9761
rect 4379 9757 4380 9761
rect 4384 9757 4385 9761
rect 4370 9756 4389 9757
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4370 9751 4389 9752
rect 4374 9747 4375 9751
rect 4379 9747 4380 9751
rect 4384 9747 4385 9751
rect 4370 9746 4389 9747
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4370 9741 4389 9742
rect 4374 9737 4375 9741
rect 4379 9737 4380 9741
rect 4384 9737 4385 9741
rect 4370 9736 4389 9737
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4396 9761 4415 9762
rect 4400 9757 4401 9761
rect 4405 9757 4406 9761
rect 4410 9757 4411 9761
rect 4396 9756 4415 9757
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4396 9751 4415 9752
rect 4400 9747 4401 9751
rect 4405 9747 4406 9751
rect 4410 9747 4411 9751
rect 4396 9746 4415 9747
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4396 9741 4415 9742
rect 4400 9737 4401 9741
rect 4405 9737 4406 9741
rect 4410 9737 4411 9741
rect 4396 9736 4415 9737
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 3857 9708 3859 9712
rect 3863 9708 3864 9712
rect 3868 9708 3869 9712
rect 3873 9708 3874 9712
rect 3878 9708 3879 9712
rect 3883 9708 3884 9712
rect 3888 9708 3889 9712
rect 3893 9708 3894 9712
rect 3898 9708 3899 9712
rect 3903 9708 3904 9712
rect 3908 9708 3909 9712
rect 3913 9708 3914 9712
rect 3918 9708 3919 9712
rect 3923 9708 3925 9712
rect 3857 9707 3925 9708
rect 3857 9703 3859 9707
rect 3863 9703 3864 9707
rect 3868 9703 3869 9707
rect 3873 9703 3874 9707
rect 3878 9703 3879 9707
rect 3883 9703 3884 9707
rect 3888 9703 3889 9707
rect 3893 9703 3894 9707
rect 3898 9703 3899 9707
rect 3903 9703 3904 9707
rect 3908 9703 3909 9707
rect 3913 9703 3914 9707
rect 3918 9703 3919 9707
rect 3923 9703 3925 9707
rect 3857 9700 3925 9703
rect 4045 9718 4046 9722
rect 4050 9718 4051 9722
rect 4055 9718 4056 9722
rect 4060 9718 4061 9722
rect 4065 9718 4066 9722
rect 4070 9718 4071 9722
rect 4075 9718 4076 9722
rect 4080 9718 4081 9722
rect 4085 9718 4086 9722
rect 4090 9718 4091 9722
rect 4095 9718 4097 9722
rect 4041 9717 4097 9718
rect 4045 9713 4046 9717
rect 4050 9713 4051 9717
rect 4055 9713 4056 9717
rect 4060 9713 4061 9717
rect 4065 9713 4066 9717
rect 4070 9713 4071 9717
rect 4075 9713 4076 9717
rect 4080 9713 4081 9717
rect 4085 9713 4086 9717
rect 4090 9713 4091 9717
rect 4095 9713 4097 9717
rect 4041 9712 4097 9713
rect 4045 9708 4046 9712
rect 4050 9708 4051 9712
rect 4055 9708 4056 9712
rect 4060 9708 4061 9712
rect 4065 9708 4066 9712
rect 4070 9708 4071 9712
rect 4075 9708 4076 9712
rect 4080 9708 4081 9712
rect 4085 9708 4086 9712
rect 4090 9708 4091 9712
rect 4095 9708 4097 9712
rect 4041 9707 4097 9708
rect 4045 9703 4046 9707
rect 4050 9703 4051 9707
rect 4055 9703 4056 9707
rect 4060 9703 4061 9707
rect 4065 9703 4066 9707
rect 4070 9703 4071 9707
rect 4075 9703 4076 9707
rect 4080 9703 4081 9707
rect 4085 9703 4086 9707
rect 4090 9703 4091 9707
rect 4095 9703 4097 9707
rect 4041 9701 4097 9703
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4100 9715 4119 9716
rect 4104 9711 4105 9715
rect 4109 9711 4110 9715
rect 4114 9711 4115 9715
rect 4100 9710 4119 9711
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4100 9705 4119 9706
rect 4104 9701 4105 9705
rect 4109 9701 4110 9705
rect 4114 9701 4115 9705
rect 4100 9700 4119 9701
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3482 9695 3501 9696
rect 3486 9691 3487 9695
rect 3491 9691 3492 9695
rect 3496 9691 3497 9695
rect 3482 9690 3501 9691
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3791 9695 3810 9696
rect 3795 9691 3796 9695
rect 3800 9691 3801 9695
rect 3805 9691 3806 9695
rect 3791 9690 3810 9691
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4100 9695 4119 9696
rect 4104 9691 4105 9695
rect 4109 9691 4110 9695
rect 4114 9691 4115 9695
rect 4100 9690 4119 9691
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4292 9715 4311 9716
rect 4296 9711 4297 9715
rect 4301 9711 4302 9715
rect 4306 9711 4307 9715
rect 4292 9710 4311 9711
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4292 9705 4311 9706
rect 4296 9701 4297 9705
rect 4301 9701 4302 9705
rect 4306 9701 4307 9705
rect 4292 9700 4311 9701
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4292 9695 4311 9696
rect 4296 9691 4297 9695
rect 4301 9691 4302 9695
rect 4306 9691 4307 9695
rect 4292 9690 4311 9691
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4318 9715 4337 9716
rect 4322 9711 4323 9715
rect 4327 9711 4328 9715
rect 4332 9711 4333 9715
rect 4318 9710 4337 9711
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4318 9705 4337 9706
rect 4322 9701 4323 9705
rect 4327 9701 4328 9705
rect 4332 9701 4333 9705
rect 4318 9700 4337 9701
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4318 9695 4337 9696
rect 4322 9691 4323 9695
rect 4327 9691 4328 9695
rect 4332 9691 4333 9695
rect 4318 9690 4337 9691
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4344 9715 4363 9716
rect 4348 9711 4349 9715
rect 4353 9711 4354 9715
rect 4358 9711 4359 9715
rect 4344 9710 4363 9711
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4344 9705 4363 9706
rect 4348 9701 4349 9705
rect 4353 9701 4354 9705
rect 4358 9701 4359 9705
rect 4344 9700 4363 9701
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4344 9695 4363 9696
rect 4348 9691 4349 9695
rect 4353 9691 4354 9695
rect 4358 9691 4359 9695
rect 4344 9690 4363 9691
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4370 9715 4389 9716
rect 4374 9711 4375 9715
rect 4379 9711 4380 9715
rect 4384 9711 4385 9715
rect 4370 9710 4389 9711
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4370 9705 4389 9706
rect 4374 9701 4375 9705
rect 4379 9701 4380 9705
rect 4384 9701 4385 9705
rect 4370 9700 4389 9701
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4370 9695 4389 9696
rect 4374 9691 4375 9695
rect 4379 9691 4380 9695
rect 4384 9691 4385 9695
rect 4370 9690 4389 9691
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4396 9715 4415 9716
rect 4400 9711 4401 9715
rect 4405 9711 4406 9715
rect 4410 9711 4411 9715
rect 4396 9710 4415 9711
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4396 9705 4415 9706
rect 4400 9701 4401 9705
rect 4405 9701 4406 9705
rect 4410 9701 4411 9705
rect 4396 9700 4415 9701
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4396 9695 4415 9696
rect 4400 9691 4401 9695
rect 4405 9691 4406 9695
rect 4410 9691 4411 9695
rect 4396 9690 4415 9691
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 3342 9685 3362 9686
rect 3342 9681 3343 9685
rect 3347 9681 3348 9685
rect 3352 9681 3353 9685
rect 3357 9681 3358 9685
rect 3342 9680 3362 9681
rect 3342 9676 3343 9680
rect 3347 9676 3348 9680
rect 3352 9676 3353 9680
rect 3357 9676 3358 9680
rect 3342 9675 3362 9676
rect 3342 9671 3343 9675
rect 3347 9671 3348 9675
rect 3352 9671 3353 9675
rect 3357 9671 3358 9675
rect 3342 9670 3362 9671
rect 3342 9666 3343 9670
rect 3347 9666 3348 9670
rect 3352 9666 3353 9670
rect 3357 9666 3358 9670
rect 3342 9665 3362 9666
rect 3342 9661 3343 9665
rect 3347 9661 3348 9665
rect 3352 9661 3353 9665
rect 3357 9661 3358 9665
rect 3342 9659 3362 9661
rect 617 9618 618 9622
rect 622 9618 623 9622
rect 627 9618 628 9622
rect 632 9618 633 9622
rect 637 9618 638 9622
rect 642 9618 643 9622
rect 613 9617 647 9618
rect 617 9613 618 9617
rect 622 9613 623 9617
rect 627 9613 628 9617
rect 632 9613 633 9617
rect 637 9613 638 9617
rect 642 9613 643 9617
rect 613 9612 647 9613
rect 617 9608 618 9612
rect 622 9608 623 9612
rect 627 9608 628 9612
rect 632 9608 633 9612
rect 637 9608 638 9612
rect 642 9608 643 9612
rect 613 9607 647 9608
rect 617 9603 618 9607
rect 622 9603 623 9607
rect 627 9603 628 9607
rect 632 9603 633 9607
rect 637 9603 638 9607
rect 642 9603 643 9607
rect 663 9618 664 9622
rect 668 9618 669 9622
rect 673 9618 674 9622
rect 678 9618 679 9622
rect 683 9618 684 9622
rect 688 9618 689 9622
rect 659 9617 693 9618
rect 663 9613 664 9617
rect 668 9613 669 9617
rect 673 9613 674 9617
rect 678 9613 679 9617
rect 683 9613 684 9617
rect 688 9613 689 9617
rect 2166 9616 2179 9623
rect 659 9612 693 9613
rect 663 9608 664 9612
rect 668 9608 669 9612
rect 673 9608 674 9612
rect 678 9608 679 9612
rect 683 9608 684 9612
rect 688 9608 689 9612
rect 659 9607 693 9608
rect 663 9603 664 9607
rect 668 9603 669 9607
rect 673 9603 674 9607
rect 678 9603 679 9607
rect 683 9603 684 9607
rect 688 9603 689 9607
rect 617 9592 618 9596
rect 622 9592 623 9596
rect 627 9592 628 9596
rect 632 9592 633 9596
rect 637 9592 638 9596
rect 642 9592 643 9596
rect 613 9591 647 9592
rect 617 9587 618 9591
rect 622 9587 623 9591
rect 627 9587 628 9591
rect 632 9587 633 9591
rect 637 9587 638 9591
rect 642 9587 643 9591
rect 613 9586 647 9587
rect 617 9582 618 9586
rect 622 9582 623 9586
rect 627 9582 628 9586
rect 632 9582 633 9586
rect 637 9582 638 9586
rect 642 9582 643 9586
rect 613 9581 647 9582
rect 617 9577 618 9581
rect 622 9577 623 9581
rect 627 9577 628 9581
rect 632 9577 633 9581
rect 637 9577 638 9581
rect 642 9577 643 9581
rect 663 9592 664 9596
rect 668 9592 669 9596
rect 673 9592 674 9596
rect 678 9592 679 9596
rect 683 9592 684 9596
rect 688 9592 689 9596
rect 659 9591 693 9592
rect 663 9587 664 9591
rect 668 9587 669 9591
rect 673 9587 674 9591
rect 678 9587 679 9591
rect 683 9587 684 9591
rect 688 9587 689 9591
rect 659 9586 693 9587
rect 663 9582 664 9586
rect 668 9582 669 9586
rect 673 9582 674 9586
rect 678 9582 679 9586
rect 683 9582 684 9586
rect 688 9582 689 9586
rect 659 9581 693 9582
rect 663 9577 664 9581
rect 668 9577 669 9581
rect 673 9577 674 9581
rect 678 9577 679 9581
rect 683 9577 684 9581
rect 688 9577 689 9581
rect 2173 9593 2179 9616
rect 2257 9619 2258 9623
rect 2257 9593 2261 9619
rect 2113 9572 2126 9593
rect 617 9566 618 9570
rect 622 9566 623 9570
rect 627 9566 628 9570
rect 632 9566 633 9570
rect 637 9566 638 9570
rect 642 9566 643 9570
rect 613 9565 647 9566
rect 617 9561 618 9565
rect 622 9561 623 9565
rect 627 9561 628 9565
rect 632 9561 633 9565
rect 637 9561 638 9565
rect 642 9561 643 9565
rect 613 9560 647 9561
rect 617 9556 618 9560
rect 622 9556 623 9560
rect 627 9556 628 9560
rect 632 9556 633 9560
rect 637 9556 638 9560
rect 642 9556 643 9560
rect 613 9555 647 9556
rect 617 9551 618 9555
rect 622 9551 623 9555
rect 627 9551 628 9555
rect 632 9551 633 9555
rect 637 9551 638 9555
rect 642 9551 643 9555
rect 663 9566 664 9570
rect 668 9566 669 9570
rect 673 9566 674 9570
rect 678 9566 679 9570
rect 683 9566 684 9570
rect 688 9566 689 9570
rect 659 9565 693 9566
rect 663 9561 664 9565
rect 668 9561 669 9565
rect 673 9561 674 9565
rect 678 9561 679 9565
rect 683 9561 684 9565
rect 688 9561 689 9565
rect 659 9560 693 9561
rect 663 9556 664 9560
rect 668 9556 669 9560
rect 673 9556 674 9560
rect 678 9556 679 9560
rect 683 9556 684 9560
rect 688 9556 689 9560
rect 659 9555 693 9556
rect 663 9551 664 9555
rect 668 9551 669 9555
rect 673 9551 674 9555
rect 678 9551 679 9555
rect 683 9551 684 9555
rect 688 9551 689 9555
rect 2476 9548 2481 9549
rect 617 9540 618 9544
rect 622 9540 623 9544
rect 627 9540 628 9544
rect 632 9540 633 9544
rect 637 9540 638 9544
rect 642 9540 643 9544
rect 613 9539 647 9540
rect 617 9535 618 9539
rect 622 9535 623 9539
rect 627 9535 628 9539
rect 632 9535 633 9539
rect 637 9535 638 9539
rect 642 9535 643 9539
rect 613 9534 647 9535
rect 617 9530 618 9534
rect 622 9530 623 9534
rect 627 9530 628 9534
rect 632 9530 633 9534
rect 637 9530 638 9534
rect 642 9530 643 9534
rect 613 9529 647 9530
rect 617 9525 618 9529
rect 622 9525 623 9529
rect 627 9525 628 9529
rect 632 9525 633 9529
rect 637 9525 638 9529
rect 642 9525 643 9529
rect 663 9540 664 9544
rect 668 9540 669 9544
rect 673 9540 674 9544
rect 678 9540 679 9544
rect 683 9540 684 9544
rect 688 9540 689 9544
rect 659 9539 693 9540
rect 663 9535 664 9539
rect 668 9535 669 9539
rect 673 9535 674 9539
rect 678 9535 679 9539
rect 683 9535 684 9539
rect 688 9535 689 9539
rect 659 9534 693 9535
rect 663 9530 664 9534
rect 668 9530 669 9534
rect 673 9530 674 9534
rect 678 9530 679 9534
rect 683 9530 684 9534
rect 688 9530 689 9534
rect 659 9529 693 9530
rect 663 9525 664 9529
rect 668 9525 669 9529
rect 673 9525 674 9529
rect 678 9525 679 9529
rect 683 9525 684 9529
rect 688 9525 689 9529
rect 617 9514 618 9518
rect 622 9514 623 9518
rect 627 9514 628 9518
rect 632 9514 633 9518
rect 637 9514 638 9518
rect 642 9514 643 9518
rect 613 9513 647 9514
rect 617 9509 618 9513
rect 622 9509 623 9513
rect 627 9509 628 9513
rect 632 9509 633 9513
rect 637 9509 638 9513
rect 642 9509 643 9513
rect 613 9508 647 9509
rect 617 9504 618 9508
rect 622 9504 623 9508
rect 627 9504 628 9508
rect 632 9504 633 9508
rect 637 9504 638 9508
rect 642 9504 643 9508
rect 613 9503 647 9504
rect 617 9499 618 9503
rect 622 9499 623 9503
rect 627 9499 628 9503
rect 632 9499 633 9503
rect 637 9499 638 9503
rect 642 9499 643 9503
rect 663 9514 664 9518
rect 668 9514 669 9518
rect 673 9514 674 9518
rect 678 9514 679 9518
rect 683 9514 684 9518
rect 688 9514 689 9518
rect 659 9513 693 9514
rect 663 9509 664 9513
rect 668 9509 669 9513
rect 673 9509 674 9513
rect 678 9509 679 9513
rect 683 9509 684 9513
rect 688 9509 689 9513
rect 659 9508 693 9509
rect 663 9504 664 9508
rect 668 9504 669 9508
rect 673 9504 674 9508
rect 678 9504 679 9508
rect 683 9504 684 9508
rect 688 9504 689 9508
rect 659 9503 693 9504
rect 663 9499 664 9503
rect 668 9499 669 9503
rect 673 9499 674 9503
rect 678 9499 679 9503
rect 683 9499 684 9503
rect 688 9499 689 9503
rect 617 9321 618 9325
rect 622 9321 623 9325
rect 627 9321 628 9325
rect 632 9321 633 9325
rect 637 9321 638 9325
rect 642 9321 643 9325
rect 613 9320 647 9321
rect 617 9316 618 9320
rect 622 9316 623 9320
rect 627 9316 628 9320
rect 632 9316 633 9320
rect 637 9316 638 9320
rect 642 9316 643 9320
rect 613 9315 647 9316
rect 617 9311 618 9315
rect 622 9311 623 9315
rect 627 9311 628 9315
rect 632 9311 633 9315
rect 637 9311 638 9315
rect 642 9311 643 9315
rect 613 9310 647 9311
rect 86 9304 346 9307
rect 617 9306 618 9310
rect 622 9306 623 9310
rect 627 9306 628 9310
rect 632 9306 633 9310
rect 637 9306 638 9310
rect 642 9306 643 9310
rect 663 9321 664 9325
rect 668 9321 669 9325
rect 673 9321 674 9325
rect 678 9321 679 9325
rect 683 9321 684 9325
rect 688 9321 689 9325
rect 659 9320 693 9321
rect 663 9316 664 9320
rect 668 9316 669 9320
rect 673 9316 674 9320
rect 678 9316 679 9320
rect 683 9316 684 9320
rect 688 9316 689 9320
rect 659 9315 693 9316
rect 663 9311 664 9315
rect 668 9311 669 9315
rect 673 9311 674 9315
rect 678 9311 679 9315
rect 683 9311 684 9315
rect 688 9311 689 9315
rect 659 9310 693 9311
rect 663 9306 664 9310
rect 668 9306 669 9310
rect 673 9306 674 9310
rect 678 9306 679 9310
rect 683 9306 684 9310
rect 688 9306 689 9310
rect 86 9050 89 9304
rect 343 9050 346 9304
rect 86 9047 346 9050
rect 617 9012 618 9016
rect 622 9012 623 9016
rect 627 9012 628 9016
rect 632 9012 633 9016
rect 637 9012 638 9016
rect 642 9012 643 9016
rect 613 9011 647 9012
rect 617 9007 618 9011
rect 622 9007 623 9011
rect 627 9007 628 9011
rect 632 9007 633 9011
rect 637 9007 638 9011
rect 642 9007 643 9011
rect 613 9006 647 9007
rect 617 9002 618 9006
rect 622 9002 623 9006
rect 627 9002 628 9006
rect 632 9002 633 9006
rect 637 9002 638 9006
rect 642 9002 643 9006
rect 613 9001 647 9002
rect 86 8995 346 8998
rect 617 8997 618 9001
rect 622 8997 623 9001
rect 627 8997 628 9001
rect 632 8997 633 9001
rect 637 8997 638 9001
rect 642 8997 643 9001
rect 663 9012 664 9016
rect 668 9012 669 9016
rect 673 9012 674 9016
rect 678 9012 679 9016
rect 683 9012 684 9016
rect 688 9012 689 9016
rect 659 9011 693 9012
rect 663 9007 664 9011
rect 668 9007 669 9011
rect 673 9007 674 9011
rect 678 9007 679 9011
rect 683 9007 684 9011
rect 688 9007 689 9011
rect 659 9006 693 9007
rect 663 9002 664 9006
rect 668 9002 669 9006
rect 673 9002 674 9006
rect 678 9002 679 9006
rect 683 9002 684 9006
rect 688 9002 689 9006
rect 659 9001 693 9002
rect 663 8997 664 9001
rect 668 8997 669 9001
rect 673 8997 674 9001
rect 678 8997 679 9001
rect 683 8997 684 9001
rect 688 8997 689 9001
rect 86 8741 89 8995
rect 343 8741 346 8995
rect 2476 8823 2480 9548
rect 2497 9386 2502 9575
rect 2788 9479 2794 9501
rect 2490 9231 2493 9280
rect 2490 9187 2493 9227
rect 2498 9224 2502 9386
rect 2506 9304 2509 9314
rect 2513 9274 2516 9283
rect 2529 9276 2532 9289
rect 2542 9261 2545 9314
rect 2609 9304 2612 9314
rect 2549 9289 2553 9293
rect 2550 9274 2553 9283
rect 2505 9247 2508 9259
rect 2546 9257 2547 9261
rect 2556 9247 2559 9300
rect 2562 9280 2565 9285
rect 2571 9274 2574 9283
rect 2587 9276 2590 9289
rect 2608 9274 2611 9283
rect 2607 9247 2610 9257
rect 2490 9172 2493 9181
rect 2351 8782 2355 8819
rect 2374 8802 2377 8812
rect 2381 8772 2384 8781
rect 2397 8774 2400 8787
rect 2410 8759 2413 8812
rect 2477 8802 2480 8812
rect 2417 8787 2421 8791
rect 2418 8772 2421 8781
rect 2373 8745 2376 8757
rect 2414 8755 2415 8759
rect 2424 8745 2427 8798
rect 2430 8778 2433 8783
rect 2439 8772 2442 8781
rect 2455 8774 2458 8787
rect 2476 8772 2479 8781
rect 2492 8772 2495 8781
rect 2475 8745 2478 8755
rect 86 8738 346 8741
rect 617 8703 618 8707
rect 622 8703 623 8707
rect 627 8703 628 8707
rect 632 8703 633 8707
rect 637 8703 638 8707
rect 642 8703 643 8707
rect 613 8702 647 8703
rect 617 8698 618 8702
rect 622 8698 623 8702
rect 627 8698 628 8702
rect 632 8698 633 8702
rect 637 8698 638 8702
rect 642 8698 643 8702
rect 613 8697 647 8698
rect 617 8693 618 8697
rect 622 8693 623 8697
rect 627 8693 628 8697
rect 632 8693 633 8697
rect 637 8693 638 8697
rect 642 8693 643 8697
rect 613 8692 647 8693
rect 86 8686 346 8689
rect 617 8688 618 8692
rect 622 8688 623 8692
rect 627 8688 628 8692
rect 632 8688 633 8692
rect 637 8688 638 8692
rect 642 8688 643 8692
rect 663 8703 664 8707
rect 668 8703 669 8707
rect 673 8703 674 8707
rect 678 8703 679 8707
rect 683 8703 684 8707
rect 688 8703 689 8707
rect 659 8702 693 8703
rect 663 8698 664 8702
rect 668 8698 669 8702
rect 673 8698 674 8702
rect 678 8698 679 8702
rect 683 8698 684 8702
rect 688 8698 689 8702
rect 659 8697 693 8698
rect 663 8693 664 8697
rect 668 8693 669 8697
rect 673 8693 674 8697
rect 678 8693 679 8697
rect 683 8693 684 8697
rect 688 8693 689 8697
rect 659 8692 693 8693
rect 663 8688 664 8692
rect 668 8688 669 8692
rect 673 8688 674 8692
rect 678 8688 679 8692
rect 683 8688 684 8692
rect 688 8688 689 8692
rect 86 8432 89 8686
rect 343 8432 346 8686
rect 2367 8640 2370 8734
rect 2492 8731 2495 8768
rect 2498 8724 2502 9220
rect 2615 9233 2619 9367
rect 2764 9344 2770 9459
rect 2764 9311 2770 9340
rect 2624 9281 2627 9283
rect 2624 9274 2627 9277
rect 2624 9240 2627 9270
rect 2764 9267 2770 9307
rect 2505 9202 2508 9212
rect 2506 9172 2509 9181
rect 2527 9174 2530 9187
rect 2543 9172 2546 9181
rect 2552 9178 2555 9183
rect 2507 9145 2510 9155
rect 2558 9145 2561 9198
rect 2564 9187 2568 9191
rect 2564 9172 2567 9181
rect 2572 9159 2575 9212
rect 2608 9202 2611 9212
rect 2585 9174 2588 9187
rect 2601 9172 2604 9181
rect 2570 9155 2571 9159
rect 2609 9145 2612 9157
rect 2506 8802 2509 8812
rect 2513 8772 2516 8781
rect 2529 8774 2532 8787
rect 2542 8759 2545 8812
rect 2609 8802 2612 8812
rect 2549 8787 2553 8791
rect 2550 8772 2553 8781
rect 2505 8745 2508 8757
rect 2546 8755 2547 8759
rect 2556 8745 2559 8798
rect 2562 8778 2565 8783
rect 2571 8772 2574 8781
rect 2587 8774 2590 8787
rect 2608 8772 2611 8781
rect 2607 8745 2610 8755
rect 2482 8711 2486 8715
rect 2482 8692 2486 8707
rect 2498 8704 2502 8720
rect 2514 8719 2518 8724
rect 2514 8711 2518 8715
rect 2514 8692 2518 8707
rect 2498 8688 2502 8689
rect 2514 8684 2518 8688
rect 2374 8660 2377 8670
rect 2381 8630 2384 8639
rect 2397 8632 2400 8645
rect 2410 8617 2413 8670
rect 2477 8660 2480 8670
rect 2417 8645 2421 8649
rect 2418 8630 2421 8639
rect 2373 8603 2376 8615
rect 2414 8613 2415 8617
rect 2424 8603 2427 8656
rect 2492 8645 2495 8677
rect 2430 8636 2433 8641
rect 2439 8630 2442 8639
rect 2455 8632 2458 8645
rect 2476 8630 2479 8639
rect 2492 8630 2495 8639
rect 2475 8603 2478 8613
rect 2367 8554 2370 8592
rect 2374 8574 2377 8584
rect 2381 8544 2384 8553
rect 2397 8546 2400 8559
rect 2410 8531 2413 8584
rect 2477 8574 2480 8584
rect 2417 8559 2421 8563
rect 2418 8544 2421 8553
rect 2373 8517 2376 8529
rect 2414 8527 2415 8531
rect 2424 8517 2427 8570
rect 2430 8550 2433 8555
rect 2439 8544 2442 8553
rect 2455 8546 2458 8559
rect 2476 8544 2479 8553
rect 2492 8544 2495 8553
rect 2475 8517 2478 8527
rect 86 8429 346 8432
rect 2367 8414 2370 8506
rect 2492 8503 2495 8540
rect 2374 8434 2377 8444
rect 2381 8404 2384 8413
rect 2397 8406 2400 8419
rect 617 8394 618 8398
rect 622 8394 623 8398
rect 627 8394 628 8398
rect 632 8394 633 8398
rect 637 8394 638 8398
rect 642 8394 643 8398
rect 613 8393 647 8394
rect 617 8389 618 8393
rect 622 8389 623 8393
rect 627 8389 628 8393
rect 632 8389 633 8393
rect 637 8389 638 8393
rect 642 8389 643 8393
rect 613 8388 647 8389
rect 617 8384 618 8388
rect 622 8384 623 8388
rect 627 8384 628 8388
rect 632 8384 633 8388
rect 637 8384 638 8388
rect 642 8384 643 8388
rect 613 8383 647 8384
rect 86 8377 346 8380
rect 617 8379 618 8383
rect 622 8379 623 8383
rect 627 8379 628 8383
rect 632 8379 633 8383
rect 637 8379 638 8383
rect 642 8379 643 8383
rect 663 8394 664 8398
rect 668 8394 669 8398
rect 673 8394 674 8398
rect 678 8394 679 8398
rect 683 8394 684 8398
rect 688 8394 689 8398
rect 659 8393 693 8394
rect 663 8389 664 8393
rect 668 8389 669 8393
rect 673 8389 674 8393
rect 678 8389 679 8393
rect 683 8389 684 8393
rect 688 8389 689 8393
rect 659 8388 693 8389
rect 663 8384 664 8388
rect 668 8384 669 8388
rect 673 8384 674 8388
rect 678 8384 679 8388
rect 683 8384 684 8388
rect 688 8384 689 8388
rect 659 8383 693 8384
rect 663 8379 664 8383
rect 668 8379 669 8383
rect 673 8379 674 8383
rect 678 8379 679 8383
rect 683 8379 684 8383
rect 688 8379 689 8383
rect 2410 8391 2413 8444
rect 2477 8434 2480 8444
rect 2417 8419 2421 8423
rect 2418 8404 2421 8413
rect 86 8123 89 8377
rect 343 8123 346 8377
rect 2373 8377 2376 8389
rect 2414 8387 2415 8391
rect 2424 8377 2427 8430
rect 2492 8419 2495 8451
rect 2430 8410 2433 8415
rect 2439 8404 2442 8413
rect 2455 8406 2458 8419
rect 2476 8404 2479 8413
rect 2492 8404 2495 8413
rect 2475 8377 2478 8387
rect 2490 8249 2493 8298
rect 2490 8205 2493 8245
rect 2498 8242 2502 8684
rect 2506 8660 2509 8670
rect 2513 8630 2516 8639
rect 2529 8632 2532 8645
rect 2542 8617 2545 8670
rect 2609 8660 2612 8670
rect 2549 8645 2553 8649
rect 2550 8630 2553 8639
rect 2505 8603 2508 8615
rect 2546 8613 2547 8617
rect 2556 8603 2559 8656
rect 2562 8636 2565 8641
rect 2571 8630 2574 8639
rect 2587 8632 2590 8645
rect 2608 8630 2611 8639
rect 2607 8603 2610 8613
rect 2506 8574 2509 8584
rect 2513 8544 2516 8553
rect 2529 8546 2532 8559
rect 2542 8531 2545 8584
rect 2609 8574 2612 8584
rect 2549 8559 2553 8563
rect 2550 8544 2553 8553
rect 2505 8517 2508 8529
rect 2546 8527 2547 8531
rect 2556 8517 2559 8570
rect 2562 8550 2565 8555
rect 2571 8544 2574 8553
rect 2587 8546 2590 8559
rect 2608 8544 2611 8553
rect 2607 8517 2610 8527
rect 2615 8496 2619 9229
rect 2639 9224 2643 9229
rect 2764 9209 2770 9263
rect 2764 9135 2770 9205
rect 2764 9003 2770 9131
rect 2764 8871 2770 8999
rect 2638 8802 2641 8812
rect 2624 8772 2627 8781
rect 2645 8772 2648 8781
rect 2661 8774 2664 8787
rect 2624 8731 2627 8768
rect 2674 8759 2677 8812
rect 2741 8802 2744 8812
rect 2764 8809 2770 8867
rect 2681 8787 2685 8791
rect 2682 8772 2685 8781
rect 2637 8745 2640 8757
rect 2678 8755 2679 8759
rect 2688 8745 2691 8798
rect 2694 8778 2697 8783
rect 2703 8772 2706 8781
rect 2719 8774 2722 8787
rect 2740 8772 2743 8781
rect 2756 8772 2759 8783
rect 2739 8745 2742 8755
rect 2756 8738 2759 8768
rect 2756 8704 2759 8734
rect 2764 8739 2770 8805
rect 2764 8697 2770 8735
rect 2624 8645 2627 8677
rect 2638 8660 2641 8670
rect 2624 8630 2627 8639
rect 2645 8630 2648 8639
rect 2661 8632 2664 8645
rect 2674 8617 2677 8670
rect 2741 8660 2744 8670
rect 2681 8645 2685 8649
rect 2682 8630 2685 8639
rect 2637 8603 2640 8615
rect 2678 8613 2679 8617
rect 2688 8603 2691 8656
rect 2756 8645 2759 8692
rect 2694 8636 2697 8641
rect 2703 8630 2706 8639
rect 2719 8632 2722 8645
rect 2740 8630 2743 8639
rect 2756 8630 2759 8641
rect 2739 8603 2742 8613
rect 2756 8596 2759 8626
rect 2764 8667 2770 8693
rect 2638 8574 2641 8584
rect 2624 8544 2627 8553
rect 2645 8544 2648 8553
rect 2661 8546 2664 8559
rect 2624 8503 2627 8540
rect 2674 8531 2677 8584
rect 2741 8574 2744 8584
rect 2764 8581 2770 8663
rect 2681 8559 2685 8563
rect 2682 8544 2685 8553
rect 2637 8517 2640 8529
rect 2678 8527 2679 8531
rect 2688 8517 2691 8570
rect 2694 8550 2697 8555
rect 2703 8544 2706 8553
rect 2719 8546 2722 8559
rect 2740 8544 2743 8553
rect 2756 8544 2759 8555
rect 2739 8517 2742 8527
rect 2756 8510 2759 8540
rect 2599 8485 2603 8488
rect 2599 8466 2603 8481
rect 2615 8478 2619 8492
rect 2631 8492 2635 8496
rect 2631 8485 2635 8488
rect 2631 8466 2635 8481
rect 2756 8478 2759 8506
rect 2615 8462 2619 8463
rect 2631 8458 2635 8462
rect 2506 8434 2509 8444
rect 2513 8404 2516 8413
rect 2529 8406 2532 8419
rect 2542 8391 2545 8444
rect 2609 8434 2612 8444
rect 2549 8419 2553 8423
rect 2550 8404 2553 8413
rect 2505 8377 2508 8389
rect 2546 8387 2547 8391
rect 2556 8377 2559 8430
rect 2562 8410 2565 8415
rect 2571 8404 2574 8413
rect 2587 8406 2590 8419
rect 2608 8404 2611 8413
rect 2607 8377 2610 8387
rect 2506 8322 2509 8332
rect 2513 8292 2516 8301
rect 2529 8294 2532 8307
rect 2542 8279 2545 8332
rect 2609 8322 2612 8332
rect 2549 8307 2553 8311
rect 2550 8292 2553 8301
rect 2505 8265 2508 8277
rect 2546 8275 2547 8279
rect 2556 8265 2559 8318
rect 2562 8298 2565 8303
rect 2571 8292 2574 8301
rect 2587 8294 2590 8307
rect 2608 8292 2611 8301
rect 2607 8265 2610 8275
rect 2490 8190 2493 8199
rect 86 8120 346 8123
rect 617 8085 618 8089
rect 622 8085 623 8089
rect 627 8085 628 8089
rect 632 8085 633 8089
rect 637 8085 638 8089
rect 642 8085 643 8089
rect 613 8084 647 8085
rect 617 8080 618 8084
rect 622 8080 623 8084
rect 627 8080 628 8084
rect 632 8080 633 8084
rect 637 8080 638 8084
rect 642 8080 643 8084
rect 613 8079 647 8080
rect 617 8075 618 8079
rect 622 8075 623 8079
rect 627 8075 628 8079
rect 632 8075 633 8079
rect 637 8075 638 8079
rect 642 8075 643 8079
rect 613 8074 647 8075
rect 86 8068 346 8071
rect 617 8070 618 8074
rect 622 8070 623 8074
rect 627 8070 628 8074
rect 632 8070 633 8074
rect 637 8070 638 8074
rect 642 8070 643 8074
rect 663 8085 664 8089
rect 668 8085 669 8089
rect 673 8085 674 8089
rect 678 8085 679 8089
rect 683 8085 684 8089
rect 688 8085 689 8089
rect 659 8084 693 8085
rect 663 8080 664 8084
rect 668 8080 669 8084
rect 673 8080 674 8084
rect 678 8080 679 8084
rect 683 8080 684 8084
rect 688 8080 689 8084
rect 659 8079 693 8080
rect 663 8075 664 8079
rect 668 8075 669 8079
rect 673 8075 674 8079
rect 678 8075 679 8079
rect 683 8075 684 8079
rect 688 8075 689 8079
rect 659 8074 693 8075
rect 663 8070 664 8074
rect 668 8070 669 8074
rect 673 8070 674 8074
rect 678 8070 679 8074
rect 683 8070 684 8074
rect 688 8070 689 8074
rect 86 7814 89 8068
rect 343 7814 346 8068
rect 2374 7820 2377 7830
rect 86 7811 346 7814
rect 2381 7790 2384 7799
rect 2397 7792 2400 7805
rect 617 7776 618 7780
rect 622 7776 623 7780
rect 627 7776 628 7780
rect 632 7776 633 7780
rect 637 7776 638 7780
rect 642 7776 643 7780
rect 613 7775 647 7776
rect 617 7771 618 7775
rect 622 7771 623 7775
rect 627 7771 628 7775
rect 632 7771 633 7775
rect 637 7771 638 7775
rect 642 7771 643 7775
rect 613 7770 647 7771
rect 617 7766 618 7770
rect 622 7766 623 7770
rect 627 7766 628 7770
rect 632 7766 633 7770
rect 637 7766 638 7770
rect 642 7766 643 7770
rect 613 7765 647 7766
rect 86 7759 346 7762
rect 617 7761 618 7765
rect 622 7761 623 7765
rect 627 7761 628 7765
rect 632 7761 633 7765
rect 637 7761 638 7765
rect 642 7761 643 7765
rect 663 7776 664 7780
rect 668 7776 669 7780
rect 673 7776 674 7780
rect 678 7776 679 7780
rect 683 7776 684 7780
rect 688 7776 689 7780
rect 659 7775 693 7776
rect 663 7771 664 7775
rect 668 7771 669 7775
rect 673 7771 674 7775
rect 678 7771 679 7775
rect 683 7771 684 7775
rect 688 7771 689 7775
rect 659 7770 693 7771
rect 663 7766 664 7770
rect 668 7766 669 7770
rect 673 7766 674 7770
rect 678 7766 679 7770
rect 683 7766 684 7770
rect 688 7766 689 7770
rect 659 7765 693 7766
rect 663 7761 664 7765
rect 668 7761 669 7765
rect 673 7761 674 7765
rect 678 7761 679 7765
rect 683 7761 684 7765
rect 688 7761 689 7765
rect 2410 7777 2413 7830
rect 2477 7820 2480 7830
rect 2417 7805 2421 7809
rect 2418 7790 2421 7799
rect 2373 7763 2376 7775
rect 2414 7773 2415 7777
rect 2424 7763 2427 7816
rect 2430 7796 2433 7801
rect 2439 7790 2442 7799
rect 2455 7792 2458 7805
rect 2476 7790 2479 7799
rect 2492 7790 2495 7799
rect 2475 7763 2478 7773
rect 86 7505 89 7759
rect 343 7505 346 7759
rect 2367 7658 2370 7752
rect 2492 7749 2495 7786
rect 2498 7742 2502 8238
rect 2615 8251 2619 8458
rect 2624 8419 2627 8451
rect 2638 8434 2641 8444
rect 2624 8404 2627 8413
rect 2645 8404 2648 8413
rect 2661 8406 2664 8419
rect 2674 8391 2677 8444
rect 2741 8434 2744 8444
rect 2681 8419 2685 8423
rect 2682 8404 2685 8413
rect 2637 8377 2640 8389
rect 2678 8387 2679 8391
rect 2688 8377 2691 8430
rect 2756 8419 2759 8466
rect 2694 8410 2697 8415
rect 2703 8404 2706 8413
rect 2719 8406 2722 8419
rect 2740 8404 2743 8413
rect 2756 8411 2759 8415
rect 2764 8441 2770 8577
rect 2756 8404 2759 8407
rect 2739 8377 2742 8387
rect 2764 8362 2770 8437
rect 2764 8329 2770 8358
rect 2624 8299 2627 8301
rect 2624 8292 2627 8295
rect 2624 8258 2627 8288
rect 2764 8285 2770 8325
rect 2505 8220 2508 8230
rect 2506 8190 2509 8199
rect 2527 8192 2530 8205
rect 2543 8190 2546 8199
rect 2552 8196 2555 8201
rect 2507 8163 2510 8173
rect 2558 8163 2561 8216
rect 2564 8205 2568 8209
rect 2564 8190 2567 8199
rect 2572 8177 2575 8230
rect 2608 8220 2611 8230
rect 2585 8192 2588 8205
rect 2601 8190 2604 8199
rect 2570 8173 2571 8177
rect 2609 8163 2612 8175
rect 2506 7820 2509 7830
rect 2513 7790 2516 7799
rect 2529 7792 2532 7805
rect 2542 7777 2545 7830
rect 2609 7820 2612 7830
rect 2549 7805 2553 7809
rect 2550 7790 2553 7799
rect 2505 7763 2508 7775
rect 2546 7773 2547 7777
rect 2556 7763 2559 7816
rect 2562 7796 2565 7801
rect 2571 7790 2574 7799
rect 2587 7792 2590 7805
rect 2608 7790 2611 7799
rect 2607 7763 2610 7773
rect 2482 7729 2486 7734
rect 2482 7710 2486 7725
rect 2498 7722 2502 7738
rect 2514 7738 2518 7742
rect 2514 7729 2518 7734
rect 2514 7710 2518 7725
rect 2498 7706 2502 7707
rect 2514 7702 2518 7706
rect 2374 7678 2377 7688
rect 2381 7648 2384 7657
rect 2397 7650 2400 7663
rect 2410 7635 2413 7688
rect 2477 7678 2480 7688
rect 2417 7663 2421 7667
rect 2418 7648 2421 7657
rect 2373 7621 2376 7633
rect 2414 7631 2415 7635
rect 2424 7621 2427 7674
rect 2492 7663 2495 7695
rect 2430 7654 2433 7659
rect 2439 7648 2442 7657
rect 2455 7650 2458 7663
rect 2476 7648 2479 7657
rect 2492 7648 2495 7657
rect 2475 7621 2478 7631
rect 2367 7572 2370 7610
rect 2374 7592 2377 7602
rect 2381 7562 2384 7571
rect 2397 7564 2400 7577
rect 2410 7549 2413 7602
rect 2477 7592 2480 7602
rect 2417 7577 2421 7581
rect 2418 7562 2421 7571
rect 2373 7535 2376 7547
rect 2414 7545 2415 7549
rect 2424 7535 2427 7588
rect 2430 7568 2433 7573
rect 2439 7562 2442 7571
rect 2455 7564 2458 7577
rect 2476 7562 2479 7571
rect 2492 7562 2495 7571
rect 2475 7535 2478 7545
rect 86 7502 346 7505
rect 617 7467 618 7471
rect 622 7467 623 7471
rect 627 7467 628 7471
rect 632 7467 633 7471
rect 637 7467 638 7471
rect 642 7467 643 7471
rect 613 7466 647 7467
rect 617 7462 618 7466
rect 622 7462 623 7466
rect 627 7462 628 7466
rect 632 7462 633 7466
rect 637 7462 638 7466
rect 642 7462 643 7466
rect 613 7461 647 7462
rect 617 7457 618 7461
rect 622 7457 623 7461
rect 627 7457 628 7461
rect 632 7457 633 7461
rect 637 7457 638 7461
rect 642 7457 643 7461
rect 613 7456 647 7457
rect 86 7450 346 7453
rect 617 7452 618 7456
rect 622 7452 623 7456
rect 627 7452 628 7456
rect 632 7452 633 7456
rect 637 7452 638 7456
rect 642 7452 643 7456
rect 663 7467 664 7471
rect 668 7467 669 7471
rect 673 7467 674 7471
rect 678 7467 679 7471
rect 683 7467 684 7471
rect 688 7467 689 7471
rect 659 7466 693 7467
rect 663 7462 664 7466
rect 668 7462 669 7466
rect 673 7462 674 7466
rect 678 7462 679 7466
rect 683 7462 684 7466
rect 688 7462 689 7466
rect 659 7461 693 7462
rect 663 7457 664 7461
rect 668 7457 669 7461
rect 673 7457 674 7461
rect 678 7457 679 7461
rect 683 7457 684 7461
rect 688 7457 689 7461
rect 659 7456 693 7457
rect 663 7452 664 7456
rect 668 7452 669 7456
rect 673 7452 674 7456
rect 678 7452 679 7456
rect 683 7452 684 7456
rect 688 7452 689 7456
rect 86 7196 89 7450
rect 343 7196 346 7450
rect 2367 7432 2370 7524
rect 2492 7521 2495 7558
rect 2374 7452 2377 7462
rect 2381 7422 2384 7431
rect 2397 7424 2400 7437
rect 2410 7409 2413 7462
rect 2477 7452 2480 7462
rect 2417 7437 2421 7441
rect 2418 7422 2421 7431
rect 2373 7395 2376 7407
rect 2414 7405 2415 7409
rect 2424 7395 2427 7448
rect 2492 7437 2495 7469
rect 2430 7428 2433 7433
rect 2439 7422 2442 7431
rect 2455 7424 2458 7437
rect 2476 7422 2479 7431
rect 2492 7422 2495 7431
rect 2475 7395 2478 7405
rect 2498 7381 2502 7702
rect 2506 7678 2509 7688
rect 2513 7648 2516 7657
rect 2529 7650 2532 7663
rect 2542 7635 2545 7688
rect 2609 7678 2612 7688
rect 2549 7663 2553 7667
rect 2550 7648 2553 7657
rect 2505 7621 2508 7633
rect 2546 7631 2547 7635
rect 2556 7621 2559 7674
rect 2562 7654 2565 7659
rect 2571 7648 2574 7657
rect 2587 7650 2590 7663
rect 2608 7648 2611 7657
rect 2607 7621 2610 7631
rect 2506 7592 2509 7602
rect 2513 7562 2516 7571
rect 2529 7564 2532 7577
rect 2542 7549 2545 7602
rect 2609 7592 2612 7602
rect 2549 7577 2553 7581
rect 2550 7562 2553 7571
rect 2505 7535 2508 7547
rect 2546 7545 2547 7549
rect 2556 7535 2559 7588
rect 2562 7568 2565 7573
rect 2571 7562 2574 7571
rect 2587 7564 2590 7577
rect 2608 7562 2611 7571
rect 2607 7535 2610 7545
rect 2615 7514 2619 8247
rect 2639 8242 2643 8247
rect 2764 8227 2770 8281
rect 2764 8153 2770 8223
rect 2764 8021 2770 8149
rect 2764 7889 2770 8017
rect 2638 7820 2641 7830
rect 2624 7790 2627 7799
rect 2645 7790 2648 7799
rect 2661 7792 2664 7805
rect 2624 7749 2627 7786
rect 2674 7777 2677 7830
rect 2741 7820 2744 7830
rect 2764 7827 2770 7885
rect 2681 7805 2685 7809
rect 2682 7790 2685 7799
rect 2637 7763 2640 7775
rect 2678 7773 2679 7777
rect 2688 7763 2691 7816
rect 2694 7796 2697 7801
rect 2703 7790 2706 7799
rect 2719 7792 2722 7805
rect 2740 7790 2743 7799
rect 2756 7790 2759 7801
rect 2739 7763 2742 7773
rect 2756 7756 2759 7786
rect 2756 7722 2759 7752
rect 2764 7757 2770 7823
rect 2764 7715 2770 7753
rect 2624 7663 2627 7695
rect 2638 7678 2641 7688
rect 2624 7648 2627 7657
rect 2645 7648 2648 7657
rect 2661 7650 2664 7663
rect 2674 7635 2677 7688
rect 2741 7678 2744 7688
rect 2681 7663 2685 7667
rect 2682 7648 2685 7657
rect 2637 7621 2640 7633
rect 2678 7631 2679 7635
rect 2688 7621 2691 7674
rect 2756 7663 2759 7710
rect 2694 7654 2697 7659
rect 2703 7648 2706 7657
rect 2719 7650 2722 7663
rect 2740 7648 2743 7657
rect 2756 7648 2759 7659
rect 2739 7621 2742 7631
rect 2756 7614 2759 7644
rect 2764 7685 2770 7711
rect 2638 7592 2641 7602
rect 2624 7562 2627 7571
rect 2645 7562 2648 7571
rect 2661 7564 2664 7577
rect 2624 7521 2627 7558
rect 2674 7549 2677 7602
rect 2741 7592 2744 7602
rect 2764 7599 2770 7681
rect 2681 7577 2685 7581
rect 2682 7562 2685 7571
rect 2637 7535 2640 7547
rect 2678 7545 2679 7549
rect 2688 7535 2691 7588
rect 2694 7568 2697 7573
rect 2703 7562 2706 7571
rect 2719 7564 2722 7577
rect 2740 7562 2743 7571
rect 2756 7562 2759 7573
rect 2739 7535 2742 7545
rect 2756 7528 2759 7558
rect 2599 7503 2603 7506
rect 2599 7484 2603 7499
rect 2615 7496 2619 7510
rect 2631 7510 2635 7514
rect 2631 7503 2635 7506
rect 2631 7484 2635 7499
rect 2756 7496 2759 7524
rect 2615 7480 2619 7481
rect 2631 7476 2635 7480
rect 2506 7452 2509 7462
rect 2513 7422 2516 7431
rect 2529 7424 2532 7437
rect 2542 7409 2545 7462
rect 2609 7452 2612 7462
rect 2549 7437 2553 7441
rect 2550 7422 2553 7431
rect 2505 7395 2508 7407
rect 2546 7405 2547 7409
rect 2556 7395 2559 7448
rect 2562 7428 2565 7433
rect 2571 7422 2574 7431
rect 2587 7424 2590 7437
rect 2608 7422 2611 7431
rect 2607 7395 2610 7405
rect 2615 7381 2619 7476
rect 2624 7437 2627 7469
rect 2638 7452 2641 7462
rect 2624 7422 2627 7431
rect 2645 7422 2648 7431
rect 2661 7424 2664 7437
rect 2674 7409 2677 7462
rect 2741 7452 2744 7462
rect 2681 7437 2685 7441
rect 2682 7422 2685 7431
rect 2637 7395 2640 7407
rect 2678 7405 2679 7409
rect 2688 7395 2691 7448
rect 2756 7437 2759 7484
rect 2694 7428 2697 7433
rect 2703 7422 2706 7431
rect 2719 7424 2722 7437
rect 2740 7422 2743 7431
rect 2756 7429 2759 7433
rect 2764 7459 2770 7595
rect 2756 7422 2759 7425
rect 2739 7395 2742 7405
rect 2764 7381 2770 7455
rect 2776 9287 2782 9466
rect 2776 9254 2782 9283
rect 2776 9201 2782 9250
rect 2776 9152 2782 9197
rect 2776 9069 2782 9148
rect 2776 8937 2782 9065
rect 2776 8805 2782 8933
rect 2776 8752 2782 8801
rect 2776 8640 2782 8748
rect 2776 8610 2782 8636
rect 2776 8554 2782 8606
rect 2776 8524 2782 8550
rect 2776 8384 2782 8520
rect 2776 8305 2782 8380
rect 2776 8272 2782 8301
rect 2776 8219 2782 8268
rect 2776 8170 2782 8215
rect 2776 8087 2782 8166
rect 2776 7955 2782 8083
rect 2776 7823 2782 7951
rect 2776 7770 2782 7819
rect 2776 7658 2782 7766
rect 2776 7628 2782 7654
rect 2776 7572 2782 7624
rect 2776 7542 2782 7568
rect 2776 7402 2782 7538
rect 2776 7381 2782 7398
rect 2788 9208 2794 9475
rect 2788 9194 2794 9204
rect 2788 9076 2794 9190
rect 2788 9062 2794 9072
rect 2788 8944 2794 9058
rect 2788 8930 2794 8940
rect 2788 8798 2794 8926
rect 2788 8724 2794 8794
rect 2788 8226 2794 8720
rect 2788 8212 2794 8222
rect 2788 8094 2794 8208
rect 2788 8080 2794 8090
rect 2788 7962 2794 8076
rect 2788 7948 2794 7958
rect 2788 7816 2794 7944
rect 2788 7742 2794 7812
rect 2788 7381 2794 7738
rect 2800 9486 2806 9501
rect 2800 9260 2806 9482
rect 2800 9128 2806 9256
rect 2800 9010 2806 9124
rect 2800 8996 2806 9006
rect 2800 8878 2806 8992
rect 2800 8864 2806 8874
rect 2800 8732 2806 8860
rect 2800 8278 2806 8728
rect 2800 8146 2806 8274
rect 2800 8028 2806 8142
rect 2800 8014 2806 8024
rect 2800 7896 2806 8010
rect 2800 7882 2806 7892
rect 2800 7750 2806 7878
rect 2800 7381 2806 7746
rect 2812 9493 2818 9501
rect 2812 9280 2818 9489
rect 2812 9247 2818 9276
rect 2812 9145 2818 9243
rect 2812 8746 2818 9141
rect 2812 8633 2818 8742
rect 2812 8603 2818 8629
rect 2812 8547 2818 8599
rect 2812 8517 2818 8543
rect 2812 8377 2818 8513
rect 2812 8298 2818 8373
rect 2812 8265 2818 8294
rect 2812 8163 2818 8261
rect 2812 7764 2818 8159
rect 2812 7651 2818 7760
rect 2812 7621 2818 7647
rect 2812 7565 2818 7617
rect 2812 7535 2818 7561
rect 2812 7395 2818 7531
rect 2812 7381 2818 7391
rect 2824 9351 2830 9497
rect 2824 9318 2830 9347
rect 2824 9216 2830 9314
rect 2824 8816 2830 9212
rect 2824 8704 2830 8812
rect 2824 8674 2830 8700
rect 2824 8618 2830 8670
rect 2824 8588 2830 8614
rect 2824 8448 2830 8584
rect 2824 8369 2830 8444
rect 2824 8336 2830 8365
rect 2824 8234 2830 8332
rect 2824 7834 2830 8230
rect 2824 7722 2830 7830
rect 2824 7692 2830 7718
rect 2824 7636 2830 7688
rect 2824 7606 2830 7632
rect 2824 7466 2830 7602
rect 2824 7381 2830 7462
rect 2836 8718 2842 9452
rect 3021 9438 3026 9605
rect 3040 9448 3053 9607
rect 3379 9606 3382 9608
rect 3327 9471 3382 9606
rect 3634 9469 3690 9604
rect 4483 9573 4484 9577
rect 4488 9573 4489 9577
rect 4493 9573 4494 9577
rect 4498 9573 4499 9577
rect 4503 9573 4504 9577
rect 4508 9573 4509 9577
rect 4479 9572 4513 9573
rect 4483 9568 4484 9572
rect 4488 9568 4489 9572
rect 4493 9568 4494 9572
rect 4498 9568 4499 9572
rect 4503 9568 4504 9572
rect 4508 9568 4509 9572
rect 4479 9567 4513 9568
rect 4483 9563 4484 9567
rect 4488 9563 4489 9567
rect 4493 9563 4494 9567
rect 4498 9563 4499 9567
rect 4503 9563 4504 9567
rect 4508 9563 4509 9567
rect 4479 9562 4513 9563
rect 4483 9558 4484 9562
rect 4488 9558 4489 9562
rect 4493 9558 4494 9562
rect 4498 9558 4499 9562
rect 4503 9558 4504 9562
rect 4508 9558 4509 9562
rect 4529 9573 4530 9577
rect 4534 9573 4535 9577
rect 4539 9573 4540 9577
rect 4544 9573 4545 9577
rect 4549 9573 4550 9577
rect 4554 9573 4555 9577
rect 4525 9572 4559 9573
rect 4529 9568 4530 9572
rect 4534 9568 4535 9572
rect 4539 9568 4540 9572
rect 4544 9568 4545 9572
rect 4549 9568 4550 9572
rect 4554 9568 4555 9572
rect 4525 9567 4559 9568
rect 4529 9563 4530 9567
rect 4534 9563 4535 9567
rect 4539 9563 4540 9567
rect 4544 9563 4545 9567
rect 4549 9563 4550 9567
rect 4554 9563 4555 9567
rect 4525 9562 4559 9563
rect 4529 9558 4530 9562
rect 4534 9558 4535 9562
rect 4539 9558 4540 9562
rect 4544 9558 4545 9562
rect 4549 9558 4550 9562
rect 4554 9558 4555 9562
rect 4483 9544 4484 9548
rect 4488 9544 4489 9548
rect 4493 9544 4494 9548
rect 4498 9544 4499 9548
rect 4503 9544 4504 9548
rect 4508 9544 4509 9548
rect 4479 9543 4513 9544
rect 4483 9539 4484 9543
rect 4488 9539 4489 9543
rect 4493 9539 4494 9543
rect 4498 9539 4499 9543
rect 4503 9539 4504 9543
rect 4508 9539 4509 9543
rect 4479 9538 4513 9539
rect 4483 9534 4484 9538
rect 4488 9534 4489 9538
rect 4493 9534 4494 9538
rect 4498 9534 4499 9538
rect 4503 9534 4504 9538
rect 4508 9534 4509 9538
rect 4479 9533 4513 9534
rect 4483 9529 4484 9533
rect 4488 9529 4489 9533
rect 4493 9529 4494 9533
rect 4498 9529 4499 9533
rect 4503 9529 4504 9533
rect 4508 9529 4509 9533
rect 4529 9544 4530 9548
rect 4534 9544 4535 9548
rect 4539 9544 4540 9548
rect 4544 9544 4545 9548
rect 4549 9544 4550 9548
rect 4554 9544 4555 9548
rect 4525 9543 4559 9544
rect 4529 9539 4530 9543
rect 4534 9539 4535 9543
rect 4539 9539 4540 9543
rect 4544 9539 4545 9543
rect 4549 9539 4550 9543
rect 4554 9539 4555 9543
rect 4525 9538 4559 9539
rect 4529 9534 4530 9538
rect 4534 9534 4535 9538
rect 4539 9534 4540 9538
rect 4544 9534 4545 9538
rect 4549 9534 4550 9538
rect 4554 9534 4555 9538
rect 4525 9533 4559 9534
rect 4529 9529 4530 9533
rect 4534 9529 4535 9533
rect 4539 9529 4540 9533
rect 4544 9529 4545 9533
rect 4549 9529 4550 9533
rect 4554 9529 4555 9533
rect 4483 9515 4484 9519
rect 4488 9515 4489 9519
rect 4493 9515 4494 9519
rect 4498 9515 4499 9519
rect 4503 9515 4504 9519
rect 4508 9515 4509 9519
rect 4479 9514 4513 9515
rect 4483 9510 4484 9514
rect 4488 9510 4489 9514
rect 4493 9510 4494 9514
rect 4498 9510 4499 9514
rect 4503 9510 4504 9514
rect 4508 9510 4509 9514
rect 4479 9509 4513 9510
rect 4483 9505 4484 9509
rect 4488 9505 4489 9509
rect 4493 9505 4494 9509
rect 4498 9505 4499 9509
rect 4503 9505 4504 9509
rect 4508 9505 4509 9509
rect 4479 9504 4513 9505
rect 4483 9500 4484 9504
rect 4488 9500 4489 9504
rect 4493 9500 4494 9504
rect 4498 9500 4499 9504
rect 4503 9500 4504 9504
rect 4508 9500 4509 9504
rect 4529 9515 4530 9519
rect 4534 9515 4535 9519
rect 4539 9515 4540 9519
rect 4544 9515 4545 9519
rect 4549 9515 4550 9519
rect 4554 9515 4555 9519
rect 4525 9514 4559 9515
rect 4529 9510 4530 9514
rect 4534 9510 4535 9514
rect 4539 9510 4540 9514
rect 4544 9510 4545 9514
rect 4549 9510 4550 9514
rect 4554 9510 4555 9514
rect 4525 9509 4559 9510
rect 4529 9505 4530 9509
rect 4534 9505 4535 9509
rect 4539 9505 4540 9509
rect 4544 9505 4545 9509
rect 4549 9505 4550 9509
rect 4554 9505 4555 9509
rect 4525 9504 4559 9505
rect 4529 9500 4530 9504
rect 4534 9500 4535 9504
rect 4539 9500 4540 9504
rect 4544 9500 4545 9504
rect 4549 9500 4550 9504
rect 4554 9500 4555 9504
rect 3327 9466 3382 9467
rect 3635 9463 3690 9469
rect 2858 9337 2861 9347
rect 2847 9317 2851 9318
rect 2865 9307 2868 9316
rect 2881 9309 2884 9322
rect 2894 9294 2897 9347
rect 2961 9337 2964 9347
rect 2990 9337 2993 9347
rect 2901 9322 2905 9326
rect 2902 9307 2905 9316
rect 2857 9280 2860 9292
rect 2898 9290 2899 9294
rect 2908 9280 2911 9333
rect 2914 9313 2917 9318
rect 2923 9307 2926 9316
rect 2939 9309 2942 9322
rect 2960 9307 2963 9316
rect 2976 9316 2979 9318
rect 2976 9313 2983 9316
rect 2976 9307 2979 9313
rect 2997 9307 3000 9316
rect 3013 9309 3016 9322
rect 2959 9280 2962 9290
rect 2976 9273 2979 9303
rect 3026 9294 3029 9347
rect 3093 9337 3096 9347
rect 3122 9337 3125 9347
rect 3033 9322 3037 9326
rect 3034 9307 3037 9316
rect 2989 9280 2992 9292
rect 3030 9290 3031 9294
rect 3040 9280 3043 9333
rect 3046 9313 3049 9318
rect 3055 9307 3058 9316
rect 3071 9309 3074 9322
rect 3092 9307 3095 9316
rect 3108 9316 3111 9318
rect 3108 9313 3115 9316
rect 3108 9307 3111 9313
rect 3129 9307 3132 9316
rect 3145 9309 3148 9322
rect 3091 9280 3094 9290
rect 2976 9270 3028 9273
rect 2856 9250 2859 9263
rect 2882 9253 2885 9256
rect 2889 9250 2892 9263
rect 2906 9250 2909 9263
rect 2856 9201 2859 9216
rect 2870 9208 2873 9212
rect 2888 9201 2891 9216
rect 2907 9201 2910 9216
rect 2913 9215 2916 9256
rect 2929 9208 2932 9249
rect 2935 9216 2938 9256
rect 2954 9208 2957 9249
rect 2963 9250 2966 9263
rect 2979 9250 2982 9263
rect 3000 9253 3003 9256
rect 3007 9250 3010 9263
rect 3025 9259 3028 9270
rect 3108 9267 3111 9303
rect 3158 9294 3161 9347
rect 3225 9337 3228 9347
rect 3254 9337 3257 9347
rect 3165 9322 3169 9326
rect 3166 9307 3169 9316
rect 3121 9280 3124 9292
rect 3162 9290 3163 9294
rect 3172 9280 3175 9333
rect 3178 9313 3181 9318
rect 3187 9307 3190 9316
rect 3203 9309 3206 9322
rect 3224 9307 3227 9316
rect 3240 9316 3243 9318
rect 3240 9313 3247 9316
rect 3240 9307 3243 9313
rect 3261 9307 3264 9316
rect 3277 9309 3280 9322
rect 3223 9280 3226 9290
rect 3240 9273 3243 9295
rect 3290 9294 3293 9347
rect 3357 9337 3360 9347
rect 3297 9322 3301 9326
rect 3298 9307 3301 9316
rect 3253 9280 3256 9292
rect 3294 9290 3295 9294
rect 3304 9280 3307 9333
rect 3310 9313 3313 9318
rect 3319 9307 3322 9316
rect 3335 9309 3338 9322
rect 3356 9307 3359 9316
rect 3372 9316 3375 9318
rect 3372 9313 3376 9316
rect 3372 9307 3375 9313
rect 3372 9299 3375 9303
rect 3355 9280 3358 9290
rect 3106 9262 3111 9267
rect 3168 9269 3243 9273
rect 3025 9256 3070 9259
rect 3025 9246 3028 9256
rect 3043 9243 3063 9246
rect 3060 9224 3063 9243
rect 2963 9201 2966 9216
rect 2978 9201 2981 9216
rect 2985 9208 2989 9211
rect 3006 9201 3009 9216
rect 2856 9182 2859 9197
rect 2870 9186 2873 9190
rect 2888 9182 2891 9197
rect 2907 9182 2910 9197
rect 2856 9135 2859 9148
rect 2882 9142 2885 9145
rect 2856 9118 2859 9131
rect 2866 9128 2870 9138
rect 2889 9135 2892 9148
rect 2906 9135 2909 9148
rect 2913 9142 2916 9183
rect 2929 9149 2932 9190
rect 2935 9142 2938 9182
rect 2954 9149 2957 9190
rect 2963 9182 2966 9197
rect 2978 9182 2981 9197
rect 2985 9187 2989 9190
rect 3006 9182 3009 9197
rect 2963 9135 2966 9148
rect 2882 9121 2885 9124
rect 2889 9118 2892 9131
rect 2906 9118 2909 9131
rect 2856 9069 2859 9084
rect 2870 9076 2873 9080
rect 2888 9069 2891 9084
rect 2907 9069 2910 9084
rect 2913 9083 2916 9124
rect 2929 9076 2932 9117
rect 2935 9084 2938 9124
rect 2954 9076 2957 9117
rect 2963 9118 2966 9131
rect 2979 9135 2982 9148
rect 3000 9142 3003 9145
rect 3007 9135 3010 9148
rect 3060 9148 3063 9220
rect 3071 9184 3074 9256
rect 3106 9259 3109 9262
rect 3106 9256 3151 9259
rect 3106 9246 3109 9256
rect 2979 9118 2982 9131
rect 3000 9121 3003 9124
rect 3007 9118 3010 9131
rect 3060 9114 3063 9144
rect 3071 9128 3074 9180
rect 3078 9168 3082 9234
rect 3066 9124 3070 9127
rect 3059 9111 3063 9114
rect 3060 9092 3063 9111
rect 2963 9069 2966 9084
rect 2978 9069 2981 9084
rect 2985 9076 2989 9079
rect 3006 9069 3009 9084
rect 2856 9050 2859 9065
rect 2870 9054 2873 9058
rect 2888 9050 2891 9065
rect 2907 9050 2910 9065
rect 2856 9003 2859 9016
rect 2882 9010 2885 9013
rect 2856 8986 2859 8999
rect 2889 9003 2892 9016
rect 2906 9003 2909 9016
rect 2913 9010 2916 9051
rect 2929 9017 2932 9058
rect 2935 9010 2938 9050
rect 2954 9017 2957 9058
rect 2963 9050 2966 9065
rect 2978 9050 2981 9065
rect 2985 9055 2989 9058
rect 3006 9050 3009 9065
rect 2963 9003 2966 9016
rect 2882 8989 2885 8992
rect 2889 8986 2892 8999
rect 2906 8986 2909 8999
rect 2856 8937 2859 8952
rect 2870 8944 2873 8948
rect 2888 8937 2891 8952
rect 2907 8937 2910 8952
rect 2913 8951 2916 8992
rect 2929 8944 2932 8985
rect 2935 8952 2938 8992
rect 2954 8944 2957 8985
rect 2963 8986 2966 8999
rect 2979 9003 2982 9016
rect 3000 9010 3003 9013
rect 3007 9003 3010 9016
rect 3060 9017 3063 9088
rect 3071 9053 3074 9124
rect 2979 8986 2982 8999
rect 3000 8989 3003 8992
rect 3007 8986 3010 8999
rect 3060 8960 3063 9013
rect 3071 8996 3074 9049
rect 3078 9037 3082 9102
rect 3066 8992 3070 8995
rect 3109 8995 3112 9246
rect 3124 9243 3144 9246
rect 3141 9224 3144 9243
rect 3141 9148 3144 9220
rect 3152 9184 3155 9256
rect 3159 9168 3163 9234
rect 3168 9135 3171 9269
rect 3372 9266 3375 9295
rect 3196 9263 3303 9266
rect 3130 9131 3171 9135
rect 3130 9127 3133 9131
rect 3130 9124 3175 9127
rect 3130 9114 3133 9124
rect 3148 9111 3168 9114
rect 3130 9109 3133 9110
rect 3165 9092 3168 9111
rect 3165 9017 3168 9088
rect 3176 9053 3179 9124
rect 3183 9037 3187 9102
rect 2963 8937 2966 8952
rect 2978 8937 2981 8952
rect 2985 8944 2989 8947
rect 3006 8937 3009 8952
rect 2856 8918 2859 8933
rect 2870 8922 2873 8926
rect 2888 8918 2891 8933
rect 2907 8918 2910 8933
rect 2856 8871 2859 8884
rect 2882 8878 2885 8881
rect 2856 8854 2859 8867
rect 2889 8871 2892 8884
rect 2906 8871 2909 8884
rect 2913 8878 2916 8919
rect 2929 8885 2932 8926
rect 2935 8878 2938 8918
rect 2954 8885 2957 8926
rect 2963 8918 2966 8933
rect 2978 8918 2981 8933
rect 2985 8923 2989 8926
rect 3006 8918 3009 8933
rect 2963 8871 2966 8884
rect 2882 8857 2885 8860
rect 2889 8854 2892 8867
rect 2906 8854 2909 8867
rect 2856 8805 2859 8820
rect 2870 8812 2873 8816
rect 2856 8786 2859 8801
rect 2879 8798 2883 8808
rect 2888 8805 2891 8820
rect 2907 8805 2910 8820
rect 2913 8819 2916 8860
rect 2929 8812 2932 8853
rect 2935 8820 2938 8860
rect 2954 8812 2957 8853
rect 2963 8854 2966 8867
rect 2979 8871 2982 8884
rect 3000 8878 3003 8881
rect 3007 8871 3010 8884
rect 3060 8882 3063 8956
rect 3071 8918 3074 8992
rect 3106 8992 3151 8995
rect 3106 8982 3109 8992
rect 3124 8979 3144 8982
rect 2979 8854 2982 8867
rect 3000 8857 3003 8860
rect 3007 8854 3010 8867
rect 3060 8828 3063 8878
rect 3071 8864 3074 8914
rect 3078 8902 3082 8970
rect 3141 8960 3144 8979
rect 3141 8882 3144 8956
rect 3152 8918 3155 8992
rect 3196 8995 3199 9263
rect 3307 9263 3375 9266
rect 3411 9258 3416 9434
rect 3321 9018 3328 9250
rect 3423 9245 3427 9444
rect 3709 9384 3715 9460
rect 3709 9344 3715 9380
rect 3361 9124 3365 9241
rect 3435 9231 3438 9280
rect 3435 9187 3438 9227
rect 3443 9224 3447 9333
rect 3451 9304 3454 9314
rect 3458 9274 3461 9283
rect 3474 9276 3477 9289
rect 3487 9261 3490 9314
rect 3554 9304 3557 9314
rect 3494 9289 3498 9293
rect 3495 9274 3498 9283
rect 3450 9247 3453 9259
rect 3491 9257 3492 9261
rect 3501 9247 3504 9300
rect 3507 9280 3510 9285
rect 3516 9274 3519 9283
rect 3532 9276 3535 9289
rect 3553 9274 3556 9283
rect 3552 9247 3555 9257
rect 3435 9172 3438 9181
rect 3443 9140 3447 9220
rect 3560 9233 3564 9333
rect 3709 9311 3715 9340
rect 3569 9281 3572 9283
rect 3569 9274 3572 9277
rect 3569 9240 3572 9270
rect 3709 9267 3715 9307
rect 3450 9202 3453 9212
rect 3451 9172 3454 9181
rect 3472 9174 3475 9187
rect 3488 9172 3491 9181
rect 3497 9178 3500 9183
rect 3452 9145 3455 9155
rect 3503 9145 3506 9198
rect 3509 9187 3513 9191
rect 3509 9172 3512 9181
rect 3517 9159 3520 9212
rect 3553 9202 3556 9212
rect 3530 9174 3533 9187
rect 3546 9172 3549 9181
rect 3515 9155 3516 9159
rect 3554 9145 3557 9157
rect 3560 9141 3564 9229
rect 3584 9224 3588 9229
rect 3709 9209 3715 9263
rect 3709 9135 3715 9205
rect 3361 9098 3364 9120
rect 3361 9095 3406 9098
rect 3361 9085 3364 9095
rect 3339 9081 3360 9085
rect 3379 9082 3399 9085
rect 3321 9004 3330 9018
rect 3321 9000 3326 9004
rect 3196 8992 3241 8995
rect 3196 8982 3199 8992
rect 3214 8979 3234 8982
rect 3159 8902 3163 8970
rect 3231 8960 3234 8979
rect 3231 8882 3234 8956
rect 3242 8918 3245 8992
rect 3249 8902 3253 8970
rect 3066 8860 3070 8863
rect 2963 8805 2966 8820
rect 2978 8805 2981 8820
rect 2985 8812 2989 8815
rect 3006 8805 3009 8820
rect 2870 8790 2873 8794
rect 2888 8786 2891 8801
rect 2907 8786 2910 8801
rect 2856 8739 2859 8752
rect 2882 8746 2885 8749
rect 2864 8732 2868 8742
rect 2889 8739 2892 8752
rect 2906 8739 2909 8752
rect 2913 8746 2916 8787
rect 2929 8753 2932 8794
rect 2935 8746 2938 8786
rect 2954 8753 2957 8794
rect 2963 8786 2966 8801
rect 2978 8786 2981 8801
rect 2985 8791 2989 8794
rect 3006 8786 3009 8801
rect 2963 8739 2966 8752
rect 2979 8739 2982 8752
rect 3000 8746 3003 8749
rect 3007 8739 3010 8752
rect 3060 8746 3063 8824
rect 3071 8782 3074 8860
rect 3078 8766 3082 8838
rect 3090 8739 3094 8752
rect 3099 8732 3102 8742
rect 3109 8725 3112 8794
rect 3131 8790 3134 8794
rect 3149 8786 3152 8801
rect 3168 8786 3171 8801
rect 3116 8739 3120 8752
rect 3143 8746 3146 8749
rect 3150 8739 3153 8752
rect 3167 8739 3170 8752
rect 3174 8746 3177 8787
rect 3190 8753 3193 8794
rect 3196 8746 3199 8786
rect 3215 8753 3218 8794
rect 3224 8786 3227 8801
rect 3239 8786 3242 8801
rect 3246 8791 3250 8794
rect 3267 8786 3270 8801
rect 3224 8739 3227 8752
rect 3240 8739 3243 8752
rect 3261 8746 3264 8749
rect 3268 8739 3271 8752
rect 3284 8733 3288 8969
rect 3326 8874 3330 9000
rect 3339 8955 3342 9081
rect 3361 9076 3364 9081
rect 3361 9073 3383 9076
rect 3396 9063 3399 9082
rect 3396 8983 3399 9059
rect 3407 9019 3410 9095
rect 3414 9003 3418 9073
rect 3593 9012 3597 9053
rect 3660 9026 3665 9065
rect 3361 8965 3406 8968
rect 3361 8955 3364 8965
rect 3379 8952 3399 8955
rect 3339 8946 3342 8951
rect 3339 8943 3383 8946
rect 3396 8933 3399 8952
rect 3326 8870 3328 8874
rect 3396 8853 3399 8929
rect 3407 8889 3410 8965
rect 3414 8873 3418 8943
rect 3488 8886 3492 8923
rect 3660 8896 3665 9022
rect 3660 8833 3665 8892
rect 3668 9037 3672 9102
rect 3668 8976 3672 9033
rect 3668 8846 3672 8972
rect 3668 8833 3672 8842
rect 3676 9021 3680 9065
rect 3676 8833 3680 9017
rect 3709 9037 3715 9131
rect 3709 9003 3715 9033
rect 3709 8871 3715 8999
rect 3443 8824 3447 8825
rect 3560 8823 3564 8824
rect 3319 8802 3322 8812
rect 3326 8772 3329 8781
rect 3342 8774 3345 8787
rect 3355 8759 3358 8812
rect 3422 8802 3425 8812
rect 3362 8787 3366 8791
rect 3363 8772 3366 8781
rect 3318 8745 3321 8757
rect 3359 8755 3360 8759
rect 3369 8745 3372 8798
rect 3375 8778 3378 8783
rect 3384 8772 3387 8781
rect 3400 8774 3403 8787
rect 3421 8772 3424 8781
rect 3437 8772 3440 8781
rect 3420 8745 3423 8755
rect 3277 8721 3278 8724
rect 2836 7736 2842 8714
rect 3142 8611 3146 8693
rect 3157 8690 3160 8700
rect 3164 8660 3167 8669
rect 3180 8662 3183 8675
rect 3193 8647 3196 8700
rect 3260 8690 3263 8700
rect 3200 8675 3204 8679
rect 3201 8660 3204 8669
rect 3156 8633 3159 8645
rect 3197 8643 3198 8647
rect 3207 8633 3210 8686
rect 3275 8675 3278 8721
rect 3213 8666 3216 8671
rect 3222 8660 3225 8669
rect 3238 8662 3241 8675
rect 3259 8660 3262 8669
rect 3275 8660 3278 8669
rect 3258 8633 3261 8643
rect 3275 8626 3278 8656
rect 3150 8584 3153 8621
rect 3157 8604 3160 8614
rect 3164 8574 3167 8583
rect 3180 8576 3183 8589
rect 3193 8561 3196 8614
rect 3260 8604 3263 8614
rect 3200 8589 3204 8593
rect 3201 8574 3204 8583
rect 3156 8547 3159 8559
rect 3197 8557 3198 8561
rect 3207 8547 3210 8600
rect 3213 8580 3216 8585
rect 3222 8574 3225 8583
rect 3238 8576 3241 8589
rect 3259 8574 3262 8583
rect 3275 8584 3278 8585
rect 3296 8587 3300 8729
rect 3312 8640 3315 8734
rect 3437 8731 3440 8768
rect 3443 8724 3447 8819
rect 3451 8802 3454 8812
rect 3458 8772 3461 8781
rect 3474 8774 3477 8787
rect 3487 8759 3490 8812
rect 3554 8802 3557 8812
rect 3494 8787 3498 8791
rect 3495 8772 3498 8781
rect 3450 8745 3453 8757
rect 3491 8755 3492 8759
rect 3501 8745 3504 8798
rect 3507 8778 3510 8783
rect 3516 8772 3519 8781
rect 3532 8774 3535 8787
rect 3553 8772 3556 8781
rect 3552 8745 3555 8755
rect 3427 8711 3431 8715
rect 3427 8692 3431 8707
rect 3443 8704 3447 8720
rect 3459 8719 3463 8724
rect 3459 8711 3463 8715
rect 3459 8692 3463 8707
rect 3443 8688 3447 8689
rect 3459 8684 3463 8688
rect 3319 8660 3322 8670
rect 3326 8630 3329 8639
rect 3342 8632 3345 8645
rect 3355 8617 3358 8670
rect 3422 8660 3425 8670
rect 3362 8645 3366 8649
rect 3363 8630 3366 8639
rect 3318 8603 3321 8615
rect 3359 8613 3360 8617
rect 3369 8603 3372 8656
rect 3437 8645 3440 8677
rect 3375 8636 3378 8641
rect 3384 8630 3387 8639
rect 3400 8632 3403 8645
rect 3421 8630 3424 8639
rect 3437 8630 3440 8639
rect 3420 8603 3423 8613
rect 3275 8579 3278 8580
rect 3258 8547 3261 8557
rect 3296 8485 3300 8567
rect 3312 8554 3315 8592
rect 3319 8574 3322 8584
rect 3326 8544 3329 8553
rect 3342 8546 3345 8559
rect 3355 8531 3358 8584
rect 3422 8574 3425 8584
rect 3362 8559 3366 8563
rect 3363 8544 3366 8553
rect 3318 8517 3321 8529
rect 3359 8527 3360 8531
rect 3369 8517 3372 8570
rect 3375 8550 3378 8555
rect 3384 8544 3387 8553
rect 3400 8546 3403 8559
rect 3421 8544 3424 8553
rect 3437 8544 3440 8553
rect 3420 8517 3423 8527
rect 3312 8414 3315 8506
rect 3437 8503 3440 8540
rect 3319 8434 3322 8444
rect 3326 8404 3329 8413
rect 3342 8406 3345 8419
rect 3355 8391 3358 8444
rect 3422 8434 3425 8444
rect 3362 8419 3366 8423
rect 3363 8404 3366 8413
rect 3318 8377 3321 8389
rect 3359 8387 3360 8391
rect 3369 8377 3372 8430
rect 3437 8419 3440 8451
rect 3375 8410 3378 8415
rect 3384 8404 3387 8413
rect 3400 8406 3403 8419
rect 3421 8404 3424 8413
rect 3437 8404 3440 8413
rect 3420 8377 3423 8387
rect 2858 8355 2861 8365
rect 2865 8325 2868 8334
rect 2881 8327 2884 8340
rect 2894 8312 2897 8365
rect 2961 8355 2964 8365
rect 2990 8355 2993 8365
rect 2901 8340 2905 8344
rect 2902 8325 2905 8334
rect 2857 8298 2860 8310
rect 2898 8308 2899 8312
rect 2908 8298 2911 8351
rect 2914 8331 2917 8336
rect 2923 8325 2926 8334
rect 2939 8327 2942 8340
rect 2960 8325 2963 8334
rect 2976 8334 2979 8336
rect 2976 8331 2983 8334
rect 2976 8325 2979 8331
rect 2997 8325 3000 8334
rect 3013 8327 3016 8340
rect 2959 8298 2962 8308
rect 2976 8291 2979 8321
rect 3026 8312 3029 8365
rect 3093 8355 3096 8365
rect 3122 8355 3125 8365
rect 3033 8340 3037 8344
rect 3034 8325 3037 8334
rect 2989 8298 2992 8310
rect 3030 8308 3031 8312
rect 3040 8298 3043 8351
rect 3046 8331 3049 8336
rect 3055 8325 3058 8334
rect 3071 8327 3074 8340
rect 3092 8325 3095 8334
rect 3108 8334 3111 8336
rect 3108 8331 3115 8334
rect 3108 8325 3111 8331
rect 3129 8325 3132 8334
rect 3145 8327 3148 8340
rect 3091 8298 3094 8308
rect 2976 8288 3028 8291
rect 2856 8268 2859 8281
rect 2882 8271 2885 8274
rect 2889 8268 2892 8281
rect 2906 8268 2909 8281
rect 2856 8219 2859 8234
rect 2870 8226 2873 8230
rect 2888 8219 2891 8234
rect 2907 8219 2910 8234
rect 2913 8233 2916 8274
rect 2929 8226 2932 8267
rect 2935 8234 2938 8274
rect 2954 8226 2957 8267
rect 2963 8268 2966 8281
rect 2979 8268 2982 8281
rect 3000 8271 3003 8274
rect 3007 8268 3010 8281
rect 3025 8277 3028 8288
rect 3108 8285 3111 8321
rect 3158 8312 3161 8365
rect 3225 8355 3228 8365
rect 3254 8355 3257 8365
rect 3165 8340 3169 8344
rect 3166 8325 3169 8334
rect 3121 8298 3124 8310
rect 3162 8308 3163 8312
rect 3172 8298 3175 8351
rect 3178 8331 3181 8336
rect 3187 8325 3190 8334
rect 3203 8327 3206 8340
rect 3224 8325 3227 8334
rect 3240 8334 3243 8336
rect 3240 8331 3247 8334
rect 3240 8325 3243 8331
rect 3261 8325 3264 8334
rect 3277 8327 3280 8340
rect 3223 8298 3226 8308
rect 3240 8291 3243 8313
rect 3290 8312 3293 8365
rect 3357 8355 3360 8365
rect 3297 8340 3301 8344
rect 3298 8325 3301 8334
rect 3253 8298 3256 8310
rect 3294 8308 3295 8312
rect 3304 8298 3307 8351
rect 3310 8331 3313 8336
rect 3319 8325 3322 8334
rect 3335 8327 3338 8340
rect 3356 8325 3359 8334
rect 3372 8334 3375 8336
rect 3372 8331 3376 8334
rect 3372 8325 3375 8331
rect 3372 8317 3375 8321
rect 3355 8298 3358 8308
rect 3106 8280 3111 8285
rect 3168 8287 3243 8291
rect 3025 8274 3070 8277
rect 3025 8264 3028 8274
rect 3043 8261 3063 8264
rect 3060 8242 3063 8261
rect 2963 8219 2966 8234
rect 2978 8219 2981 8234
rect 2985 8226 2989 8229
rect 3006 8219 3009 8234
rect 2856 8200 2859 8215
rect 2870 8204 2873 8208
rect 2888 8200 2891 8215
rect 2907 8200 2910 8215
rect 2856 8153 2859 8166
rect 2882 8160 2885 8163
rect 2856 8136 2859 8149
rect 2866 8146 2870 8156
rect 2889 8153 2892 8166
rect 2906 8153 2909 8166
rect 2913 8160 2916 8201
rect 2929 8167 2932 8208
rect 2935 8160 2938 8200
rect 2954 8167 2957 8208
rect 2963 8200 2966 8215
rect 2978 8200 2981 8215
rect 2985 8205 2989 8208
rect 3006 8200 3009 8215
rect 2963 8153 2966 8166
rect 2882 8139 2885 8142
rect 2889 8136 2892 8149
rect 2906 8136 2909 8149
rect 2856 8087 2859 8102
rect 2870 8094 2873 8098
rect 2888 8087 2891 8102
rect 2907 8087 2910 8102
rect 2913 8101 2916 8142
rect 2929 8094 2932 8135
rect 2935 8102 2938 8142
rect 2954 8094 2957 8135
rect 2963 8136 2966 8149
rect 2979 8153 2982 8166
rect 3000 8160 3003 8163
rect 3007 8153 3010 8166
rect 3060 8166 3063 8238
rect 3071 8202 3074 8274
rect 3106 8277 3109 8280
rect 3106 8274 3151 8277
rect 3106 8264 3109 8274
rect 2979 8136 2982 8149
rect 3000 8139 3003 8142
rect 3007 8136 3010 8149
rect 3060 8132 3063 8162
rect 3071 8146 3074 8198
rect 3078 8186 3082 8252
rect 3066 8142 3070 8145
rect 3059 8129 3063 8132
rect 3060 8110 3063 8129
rect 2963 8087 2966 8102
rect 2978 8087 2981 8102
rect 2985 8094 2989 8097
rect 3006 8087 3009 8102
rect 2856 8068 2859 8083
rect 2870 8072 2873 8076
rect 2888 8068 2891 8083
rect 2907 8068 2910 8083
rect 2856 8021 2859 8034
rect 2882 8028 2885 8031
rect 2856 8004 2859 8017
rect 2889 8021 2892 8034
rect 2906 8021 2909 8034
rect 2913 8028 2916 8069
rect 2929 8035 2932 8076
rect 2935 8028 2938 8068
rect 2954 8035 2957 8076
rect 2963 8068 2966 8083
rect 2978 8068 2981 8083
rect 2985 8073 2989 8076
rect 3006 8068 3009 8083
rect 2963 8021 2966 8034
rect 2882 8007 2885 8010
rect 2889 8004 2892 8017
rect 2906 8004 2909 8017
rect 2856 7955 2859 7970
rect 2870 7962 2873 7966
rect 2888 7955 2891 7970
rect 2907 7955 2910 7970
rect 2913 7969 2916 8010
rect 2929 7962 2932 8003
rect 2935 7970 2938 8010
rect 2954 7962 2957 8003
rect 2963 8004 2966 8017
rect 2979 8021 2982 8034
rect 3000 8028 3003 8031
rect 3007 8021 3010 8034
rect 3060 8035 3063 8106
rect 3071 8071 3074 8142
rect 2979 8004 2982 8017
rect 3000 8007 3003 8010
rect 3007 8004 3010 8017
rect 3060 7978 3063 8031
rect 3071 8014 3074 8067
rect 3078 8055 3082 8120
rect 3066 8010 3070 8013
rect 3109 8013 3112 8264
rect 3124 8261 3144 8264
rect 3141 8242 3144 8261
rect 3141 8166 3144 8238
rect 3152 8202 3155 8274
rect 3159 8186 3163 8252
rect 3168 8153 3171 8287
rect 3372 8284 3375 8313
rect 3196 8281 3303 8284
rect 3130 8149 3171 8153
rect 3130 8145 3133 8149
rect 3130 8142 3175 8145
rect 3130 8132 3133 8142
rect 3148 8129 3168 8132
rect 3130 8127 3133 8128
rect 3165 8110 3168 8129
rect 3165 8035 3168 8106
rect 3176 8071 3179 8142
rect 3183 8055 3187 8120
rect 2963 7955 2966 7970
rect 2978 7955 2981 7970
rect 2985 7962 2989 7965
rect 3006 7955 3009 7970
rect 2856 7936 2859 7951
rect 2870 7940 2873 7944
rect 2888 7936 2891 7951
rect 2907 7936 2910 7951
rect 2856 7889 2859 7902
rect 2882 7896 2885 7899
rect 2856 7872 2859 7885
rect 2889 7889 2892 7902
rect 2906 7889 2909 7902
rect 2913 7896 2916 7937
rect 2929 7903 2932 7944
rect 2935 7896 2938 7936
rect 2954 7903 2957 7944
rect 2963 7936 2966 7951
rect 2978 7936 2981 7951
rect 2985 7941 2989 7944
rect 3006 7936 3009 7951
rect 2963 7889 2966 7902
rect 2882 7875 2885 7878
rect 2889 7872 2892 7885
rect 2906 7872 2909 7885
rect 2856 7823 2859 7838
rect 2870 7830 2873 7834
rect 2856 7804 2859 7819
rect 2879 7816 2883 7826
rect 2888 7823 2891 7838
rect 2907 7823 2910 7838
rect 2913 7837 2916 7878
rect 2929 7830 2932 7871
rect 2935 7838 2938 7878
rect 2954 7830 2957 7871
rect 2963 7872 2966 7885
rect 2979 7889 2982 7902
rect 3000 7896 3003 7899
rect 3007 7889 3010 7902
rect 3060 7900 3063 7974
rect 3071 7936 3074 8010
rect 3106 8010 3151 8013
rect 3106 8000 3109 8010
rect 3124 7997 3144 8000
rect 2979 7872 2982 7885
rect 3000 7875 3003 7878
rect 3007 7872 3010 7885
rect 3060 7846 3063 7896
rect 3071 7882 3074 7932
rect 3078 7920 3082 7988
rect 3141 7978 3144 7997
rect 3141 7900 3144 7974
rect 3152 7936 3155 8010
rect 3196 8013 3199 8281
rect 3307 8281 3375 8284
rect 3435 8249 3438 8298
rect 3435 8205 3438 8245
rect 3443 8242 3447 8684
rect 3451 8660 3454 8670
rect 3458 8630 3461 8639
rect 3474 8632 3477 8645
rect 3487 8617 3490 8670
rect 3554 8660 3557 8670
rect 3494 8645 3498 8649
rect 3495 8630 3498 8639
rect 3450 8603 3453 8615
rect 3491 8613 3492 8617
rect 3501 8603 3504 8656
rect 3507 8636 3510 8641
rect 3516 8630 3519 8639
rect 3532 8632 3535 8645
rect 3553 8630 3556 8639
rect 3552 8603 3555 8613
rect 3451 8574 3454 8584
rect 3458 8544 3461 8553
rect 3474 8546 3477 8559
rect 3487 8531 3490 8584
rect 3554 8574 3557 8584
rect 3494 8559 3498 8563
rect 3495 8544 3498 8553
rect 3450 8517 3453 8529
rect 3491 8527 3492 8531
rect 3501 8517 3504 8570
rect 3507 8550 3510 8555
rect 3516 8544 3519 8553
rect 3532 8546 3535 8559
rect 3553 8544 3556 8553
rect 3552 8517 3555 8527
rect 3560 8496 3564 8818
rect 3583 8802 3586 8812
rect 3569 8772 3572 8781
rect 3590 8772 3593 8781
rect 3606 8774 3609 8787
rect 3569 8731 3572 8768
rect 3619 8759 3622 8812
rect 3686 8802 3689 8812
rect 3709 8809 3715 8867
rect 3626 8787 3630 8791
rect 3627 8772 3630 8781
rect 3582 8745 3585 8757
rect 3623 8755 3624 8759
rect 3633 8745 3636 8798
rect 3639 8778 3642 8783
rect 3648 8772 3651 8781
rect 3664 8774 3667 8787
rect 3685 8772 3688 8781
rect 3701 8772 3704 8783
rect 3684 8745 3687 8755
rect 3701 8738 3704 8768
rect 3701 8704 3704 8734
rect 3709 8739 3715 8805
rect 3709 8697 3715 8735
rect 3569 8645 3572 8677
rect 3583 8660 3586 8670
rect 3569 8630 3572 8639
rect 3590 8630 3593 8639
rect 3606 8632 3609 8645
rect 3619 8617 3622 8670
rect 3686 8660 3689 8670
rect 3626 8645 3630 8649
rect 3627 8630 3630 8639
rect 3582 8603 3585 8615
rect 3623 8613 3624 8617
rect 3633 8603 3636 8656
rect 3701 8645 3704 8692
rect 3639 8636 3642 8641
rect 3648 8630 3651 8639
rect 3664 8632 3667 8645
rect 3685 8630 3688 8639
rect 3701 8630 3704 8641
rect 3684 8603 3687 8613
rect 3701 8596 3704 8626
rect 3709 8667 3715 8693
rect 3583 8574 3586 8584
rect 3569 8544 3572 8553
rect 3590 8544 3593 8553
rect 3606 8546 3609 8559
rect 3569 8503 3572 8540
rect 3619 8531 3622 8584
rect 3686 8574 3689 8584
rect 3709 8581 3715 8663
rect 3626 8559 3630 8563
rect 3627 8544 3630 8553
rect 3582 8517 3585 8529
rect 3623 8527 3624 8531
rect 3633 8517 3636 8570
rect 3639 8550 3642 8555
rect 3648 8544 3651 8553
rect 3664 8546 3667 8559
rect 3685 8544 3688 8553
rect 3701 8544 3704 8555
rect 3684 8517 3687 8527
rect 3701 8510 3704 8540
rect 3544 8485 3548 8488
rect 3544 8466 3548 8481
rect 3560 8478 3564 8492
rect 3576 8492 3580 8496
rect 3576 8485 3580 8488
rect 3576 8466 3580 8481
rect 3701 8478 3704 8506
rect 3560 8462 3564 8463
rect 3576 8458 3580 8462
rect 3451 8434 3454 8444
rect 3458 8404 3461 8413
rect 3474 8406 3477 8419
rect 3487 8391 3490 8444
rect 3554 8434 3557 8444
rect 3494 8419 3498 8423
rect 3495 8404 3498 8413
rect 3450 8377 3453 8389
rect 3491 8387 3492 8391
rect 3501 8377 3504 8430
rect 3507 8410 3510 8415
rect 3516 8404 3519 8413
rect 3532 8406 3535 8419
rect 3553 8404 3556 8413
rect 3552 8377 3555 8387
rect 3451 8322 3454 8332
rect 3458 8292 3461 8301
rect 3474 8294 3477 8307
rect 3487 8279 3490 8332
rect 3554 8322 3557 8332
rect 3494 8307 3498 8311
rect 3495 8292 3498 8301
rect 3450 8265 3453 8277
rect 3491 8275 3492 8279
rect 3501 8265 3504 8318
rect 3507 8298 3510 8303
rect 3516 8292 3519 8301
rect 3532 8294 3535 8307
rect 3553 8292 3556 8301
rect 3552 8265 3555 8275
rect 3435 8190 3438 8199
rect 3196 8010 3241 8013
rect 3196 8000 3199 8010
rect 3214 7997 3234 8000
rect 3159 7920 3163 7988
rect 3231 7978 3234 7997
rect 3231 7900 3234 7974
rect 3242 7936 3245 8010
rect 3249 7920 3253 7988
rect 3066 7878 3070 7881
rect 2963 7823 2966 7838
rect 2978 7823 2981 7838
rect 2985 7830 2989 7833
rect 3006 7823 3009 7838
rect 2870 7808 2873 7812
rect 2888 7804 2891 7819
rect 2907 7804 2910 7819
rect 2856 7757 2859 7770
rect 2882 7764 2885 7767
rect 2864 7750 2868 7760
rect 2889 7757 2892 7770
rect 2906 7757 2909 7770
rect 2913 7764 2916 7805
rect 2929 7771 2932 7812
rect 2935 7764 2938 7804
rect 2954 7771 2957 7812
rect 2963 7804 2966 7819
rect 2978 7804 2981 7819
rect 2985 7809 2989 7812
rect 3006 7804 3009 7819
rect 2963 7757 2966 7770
rect 2979 7757 2982 7770
rect 3000 7764 3003 7767
rect 3007 7757 3010 7770
rect 3060 7764 3063 7842
rect 3071 7800 3074 7878
rect 3078 7784 3082 7856
rect 3090 7757 3094 7770
rect 3099 7750 3102 7760
rect 3109 7743 3112 7812
rect 3131 7808 3134 7812
rect 3149 7804 3152 7819
rect 3168 7804 3171 7819
rect 3116 7757 3120 7770
rect 3143 7764 3146 7767
rect 3150 7757 3153 7770
rect 3167 7757 3170 7770
rect 3174 7764 3177 7805
rect 3190 7771 3193 7812
rect 3196 7764 3199 7804
rect 3215 7771 3218 7812
rect 3224 7804 3227 7819
rect 3239 7804 3242 7819
rect 3246 7809 3250 7812
rect 3267 7804 3270 7819
rect 3224 7757 3227 7770
rect 3240 7757 3243 7770
rect 3261 7764 3264 7767
rect 3268 7757 3271 7770
rect 3284 7751 3288 7987
rect 3319 7820 3322 7830
rect 3326 7790 3329 7799
rect 3342 7792 3345 7805
rect 3355 7777 3358 7830
rect 3422 7820 3425 7830
rect 3362 7805 3366 7809
rect 3363 7790 3366 7799
rect 3318 7763 3321 7775
rect 3359 7773 3360 7777
rect 3369 7763 3372 7816
rect 3375 7796 3378 7801
rect 3384 7790 3387 7799
rect 3400 7792 3403 7805
rect 3421 7790 3424 7799
rect 3437 7790 3440 7799
rect 3420 7763 3423 7773
rect 3277 7739 3278 7742
rect 2836 7381 2842 7732
rect 3142 7629 3146 7711
rect 3157 7708 3160 7718
rect 3164 7678 3167 7687
rect 3180 7680 3183 7693
rect 3193 7665 3196 7718
rect 3260 7708 3263 7718
rect 3200 7693 3204 7697
rect 3201 7678 3204 7687
rect 3156 7651 3159 7663
rect 3197 7661 3198 7665
rect 3207 7651 3210 7704
rect 3275 7693 3278 7739
rect 3213 7684 3216 7689
rect 3222 7678 3225 7687
rect 3238 7680 3241 7693
rect 3259 7678 3262 7687
rect 3275 7678 3278 7687
rect 3258 7651 3261 7661
rect 3275 7644 3278 7674
rect 3150 7602 3153 7639
rect 3157 7622 3160 7632
rect 3164 7592 3167 7601
rect 3180 7594 3183 7607
rect 3193 7579 3196 7632
rect 3260 7622 3263 7632
rect 3200 7607 3204 7611
rect 3201 7592 3204 7601
rect 3156 7565 3159 7577
rect 3197 7575 3198 7579
rect 3207 7565 3210 7618
rect 3213 7598 3216 7603
rect 3222 7592 3225 7601
rect 3238 7594 3241 7607
rect 3259 7592 3262 7601
rect 3275 7602 3278 7603
rect 3296 7605 3300 7747
rect 3312 7658 3315 7752
rect 3437 7749 3440 7786
rect 3443 7742 3447 8238
rect 3560 8251 3564 8458
rect 3569 8419 3572 8451
rect 3583 8434 3586 8444
rect 3569 8404 3572 8413
rect 3590 8404 3593 8413
rect 3606 8406 3609 8419
rect 3619 8391 3622 8444
rect 3686 8434 3689 8444
rect 3626 8419 3630 8423
rect 3627 8404 3630 8413
rect 3582 8377 3585 8389
rect 3623 8387 3624 8391
rect 3633 8377 3636 8430
rect 3701 8419 3704 8466
rect 3639 8410 3642 8415
rect 3648 8404 3651 8413
rect 3664 8406 3667 8419
rect 3685 8404 3688 8413
rect 3701 8411 3704 8415
rect 3709 8441 3715 8577
rect 3701 8404 3704 8407
rect 3684 8377 3687 8387
rect 3709 8362 3715 8437
rect 3709 8329 3715 8358
rect 3569 8300 3572 8301
rect 3569 8295 3573 8296
rect 3569 8292 3572 8295
rect 3569 8258 3572 8288
rect 3709 8285 3715 8325
rect 3450 8220 3453 8230
rect 3451 8190 3454 8199
rect 3472 8192 3475 8205
rect 3488 8190 3491 8199
rect 3497 8196 3500 8201
rect 3452 8163 3455 8173
rect 3503 8163 3506 8216
rect 3509 8205 3513 8209
rect 3509 8190 3512 8199
rect 3517 8177 3520 8230
rect 3553 8220 3556 8230
rect 3530 8192 3533 8205
rect 3546 8190 3549 8199
rect 3515 8173 3516 8177
rect 3554 8163 3557 8175
rect 3451 7820 3454 7830
rect 3458 7790 3461 7799
rect 3474 7792 3477 7805
rect 3487 7777 3490 7830
rect 3554 7820 3557 7830
rect 3494 7805 3498 7809
rect 3495 7790 3498 7799
rect 3450 7763 3453 7775
rect 3491 7773 3492 7777
rect 3501 7763 3504 7816
rect 3507 7796 3510 7801
rect 3516 7790 3519 7799
rect 3532 7792 3535 7805
rect 3553 7790 3556 7799
rect 3552 7763 3555 7773
rect 3427 7729 3431 7734
rect 3427 7710 3431 7725
rect 3443 7722 3447 7738
rect 3459 7738 3463 7742
rect 3459 7729 3463 7734
rect 3459 7710 3463 7725
rect 3443 7706 3447 7707
rect 3459 7702 3463 7706
rect 3319 7678 3322 7688
rect 3326 7648 3329 7657
rect 3342 7650 3345 7663
rect 3355 7635 3358 7688
rect 3422 7678 3425 7688
rect 3362 7663 3366 7667
rect 3363 7648 3366 7657
rect 3318 7621 3321 7633
rect 3359 7631 3360 7635
rect 3369 7621 3372 7674
rect 3437 7663 3440 7695
rect 3375 7654 3378 7659
rect 3384 7648 3387 7657
rect 3400 7650 3403 7663
rect 3421 7648 3424 7657
rect 3437 7648 3440 7657
rect 3420 7621 3423 7631
rect 3275 7597 3278 7598
rect 3258 7565 3261 7575
rect 3296 7503 3300 7585
rect 3312 7572 3315 7610
rect 3319 7592 3322 7602
rect 3326 7562 3329 7571
rect 3342 7564 3345 7577
rect 3355 7549 3358 7602
rect 3422 7592 3425 7602
rect 3362 7577 3366 7581
rect 3363 7562 3366 7571
rect 3318 7535 3321 7547
rect 3359 7545 3360 7549
rect 3369 7535 3372 7588
rect 3375 7568 3378 7573
rect 3384 7562 3387 7571
rect 3400 7564 3403 7577
rect 3421 7562 3424 7571
rect 3437 7562 3440 7571
rect 3420 7535 3423 7545
rect 3312 7432 3315 7524
rect 3437 7521 3440 7558
rect 3319 7452 3322 7462
rect 3326 7422 3329 7431
rect 3342 7424 3345 7437
rect 3355 7409 3358 7462
rect 3422 7452 3425 7462
rect 3362 7437 3366 7441
rect 3363 7422 3366 7431
rect 3318 7395 3321 7407
rect 3359 7405 3360 7409
rect 3369 7395 3372 7448
rect 3437 7437 3440 7469
rect 3375 7428 3378 7433
rect 3384 7422 3387 7431
rect 3400 7424 3403 7437
rect 3421 7422 3424 7431
rect 3437 7422 3440 7431
rect 3420 7395 3423 7405
rect 3443 7381 3447 7702
rect 3451 7678 3454 7688
rect 3458 7648 3461 7657
rect 3474 7650 3477 7663
rect 3487 7635 3490 7688
rect 3554 7678 3557 7688
rect 3494 7663 3498 7667
rect 3495 7648 3498 7657
rect 3450 7621 3453 7633
rect 3491 7631 3492 7635
rect 3501 7621 3504 7674
rect 3507 7654 3510 7659
rect 3516 7648 3519 7657
rect 3532 7650 3535 7663
rect 3553 7648 3556 7657
rect 3552 7621 3555 7631
rect 3451 7592 3454 7602
rect 3458 7562 3461 7571
rect 3474 7564 3477 7577
rect 3487 7549 3490 7602
rect 3554 7592 3557 7602
rect 3494 7577 3498 7581
rect 3495 7562 3498 7571
rect 3450 7535 3453 7547
rect 3491 7545 3492 7549
rect 3501 7535 3504 7588
rect 3507 7568 3510 7573
rect 3516 7562 3519 7571
rect 3532 7564 3535 7577
rect 3553 7562 3556 7571
rect 3552 7535 3555 7545
rect 3560 7514 3564 8247
rect 3584 8242 3588 8247
rect 3709 8227 3715 8281
rect 3709 8153 3715 8223
rect 3709 8021 3715 8149
rect 3709 7889 3715 8017
rect 3583 7820 3586 7830
rect 3569 7790 3572 7799
rect 3590 7790 3593 7799
rect 3606 7792 3609 7805
rect 3569 7749 3572 7786
rect 3619 7777 3622 7830
rect 3686 7820 3689 7830
rect 3709 7827 3715 7885
rect 3626 7805 3630 7809
rect 3627 7790 3630 7799
rect 3582 7763 3585 7775
rect 3623 7773 3624 7777
rect 3633 7763 3636 7816
rect 3639 7796 3642 7801
rect 3648 7790 3651 7799
rect 3664 7792 3667 7805
rect 3685 7790 3688 7799
rect 3701 7790 3704 7801
rect 3684 7763 3687 7773
rect 3701 7756 3704 7786
rect 3701 7722 3704 7752
rect 3709 7757 3715 7823
rect 3709 7715 3715 7753
rect 3569 7663 3572 7695
rect 3583 7678 3586 7688
rect 3569 7648 3572 7657
rect 3590 7648 3593 7657
rect 3606 7650 3609 7663
rect 3619 7635 3622 7688
rect 3686 7678 3689 7688
rect 3626 7663 3630 7667
rect 3627 7648 3630 7657
rect 3582 7621 3585 7633
rect 3623 7631 3624 7635
rect 3633 7621 3636 7674
rect 3701 7663 3704 7710
rect 3639 7654 3642 7659
rect 3648 7648 3651 7657
rect 3664 7650 3667 7663
rect 3685 7648 3688 7657
rect 3701 7648 3704 7659
rect 3684 7621 3687 7631
rect 3701 7614 3704 7644
rect 3709 7685 3715 7711
rect 3583 7592 3586 7602
rect 3569 7562 3572 7571
rect 3590 7562 3593 7571
rect 3606 7564 3609 7577
rect 3569 7521 3572 7558
rect 3619 7549 3622 7602
rect 3686 7592 3689 7602
rect 3709 7599 3715 7681
rect 3626 7577 3630 7581
rect 3627 7562 3630 7571
rect 3582 7535 3585 7547
rect 3623 7545 3624 7549
rect 3633 7535 3636 7588
rect 3639 7568 3642 7573
rect 3648 7562 3651 7571
rect 3664 7564 3667 7577
rect 3685 7562 3688 7571
rect 3701 7562 3704 7573
rect 3684 7535 3687 7545
rect 3701 7528 3704 7558
rect 3544 7503 3548 7506
rect 3544 7484 3548 7499
rect 3560 7496 3564 7510
rect 3576 7510 3580 7514
rect 3576 7503 3580 7506
rect 3576 7484 3580 7499
rect 3701 7496 3704 7524
rect 3560 7480 3564 7481
rect 3576 7476 3580 7480
rect 3451 7452 3454 7462
rect 3458 7422 3461 7431
rect 3474 7424 3477 7437
rect 3487 7409 3490 7462
rect 3554 7452 3557 7462
rect 3494 7437 3498 7441
rect 3495 7422 3498 7431
rect 3450 7395 3453 7407
rect 3491 7405 3492 7409
rect 3501 7395 3504 7448
rect 3507 7428 3510 7433
rect 3516 7422 3519 7431
rect 3532 7424 3535 7437
rect 3553 7422 3556 7431
rect 3552 7395 3555 7405
rect 3560 7381 3564 7476
rect 3569 7437 3572 7469
rect 3583 7452 3586 7462
rect 3569 7422 3572 7431
rect 3590 7422 3593 7431
rect 3606 7424 3609 7437
rect 3619 7409 3622 7462
rect 3686 7452 3689 7462
rect 3626 7437 3630 7441
rect 3627 7422 3630 7431
rect 3582 7395 3585 7407
rect 3623 7405 3624 7409
rect 3633 7395 3636 7448
rect 3701 7437 3704 7484
rect 3639 7428 3642 7433
rect 3648 7422 3651 7431
rect 3664 7424 3667 7437
rect 3685 7422 3688 7431
rect 3701 7429 3704 7433
rect 3709 7459 3715 7595
rect 3701 7422 3704 7425
rect 3684 7395 3687 7405
rect 3709 7381 3715 7455
rect 3721 9392 3727 9467
rect 3721 9287 3727 9388
rect 3721 9254 3727 9283
rect 3721 9201 3727 9250
rect 3721 9152 3727 9197
rect 3721 9069 3727 9148
rect 3721 9030 3727 9065
rect 3721 8937 3727 9026
rect 3721 8805 3727 8933
rect 3721 8752 3727 8801
rect 3721 8640 3727 8748
rect 3721 8610 3727 8636
rect 3721 8554 3727 8606
rect 3721 8524 3727 8550
rect 3721 8384 3727 8520
rect 3721 8305 3727 8380
rect 3721 8272 3727 8301
rect 3721 8219 3727 8268
rect 3721 8170 3727 8215
rect 3721 8087 3727 8166
rect 3721 7955 3727 8083
rect 3721 7823 3727 7951
rect 3721 7770 3727 7819
rect 3721 7658 3727 7766
rect 3721 7628 3727 7654
rect 3721 7572 3727 7624
rect 3721 7542 3727 7568
rect 3721 7402 3727 7538
rect 3721 7381 3727 7398
rect 3733 9400 3739 9475
rect 3733 9208 3739 9396
rect 3733 9194 3739 9204
rect 3733 9076 3739 9190
rect 3733 9062 3739 9072
rect 3733 9012 3739 9058
rect 3733 8944 3739 9008
rect 3733 8930 3739 8940
rect 3733 8798 3739 8926
rect 3733 8724 3739 8794
rect 3733 8226 3739 8720
rect 3733 8212 3739 8222
rect 3733 8094 3739 8208
rect 3733 8080 3739 8090
rect 3733 7962 3739 8076
rect 3733 7948 3739 7958
rect 3733 7816 3739 7944
rect 3733 7742 3739 7812
rect 3733 7381 3739 7738
rect 3745 9408 3751 9482
rect 3745 9260 3751 9404
rect 3745 9128 3751 9256
rect 3745 9049 3751 9124
rect 3745 9010 3751 9045
rect 3745 8996 3751 9006
rect 3745 8878 3751 8992
rect 3745 8864 3751 8874
rect 3745 8732 3751 8860
rect 3745 8278 3751 8728
rect 3745 8146 3751 8274
rect 3745 8028 3751 8142
rect 3745 8014 3751 8024
rect 3745 7896 3751 8010
rect 3745 7882 3751 7892
rect 3745 7750 3751 7878
rect 3745 7381 3751 7746
rect 3757 9416 3763 9489
rect 3757 9280 3763 9412
rect 3757 9247 3763 9276
rect 3757 9145 3763 9243
rect 3757 8886 3763 9141
rect 3757 8746 3763 8882
rect 3757 8633 3763 8742
rect 3757 8603 3763 8629
rect 3757 8547 3763 8599
rect 3757 8517 3763 8543
rect 3757 8377 3763 8513
rect 3757 8298 3763 8373
rect 3757 8265 3763 8294
rect 3757 8163 3763 8261
rect 3757 7764 3763 8159
rect 3757 7651 3763 7760
rect 3757 7621 3763 7647
rect 3757 7565 3763 7617
rect 3757 7535 3763 7561
rect 3757 7395 3763 7531
rect 3757 7381 3763 7391
rect 3769 9351 3775 9497
rect 4483 9486 4484 9490
rect 4488 9486 4489 9490
rect 4493 9486 4494 9490
rect 4498 9486 4499 9490
rect 4503 9486 4504 9490
rect 4508 9486 4509 9490
rect 4479 9485 4513 9486
rect 4483 9481 4484 9485
rect 4488 9481 4489 9485
rect 4493 9481 4494 9485
rect 4498 9481 4499 9485
rect 4503 9481 4504 9485
rect 4508 9481 4509 9485
rect 4479 9480 4513 9481
rect 4483 9476 4484 9480
rect 4488 9476 4489 9480
rect 4493 9476 4494 9480
rect 4498 9476 4499 9480
rect 4503 9476 4504 9480
rect 4508 9476 4509 9480
rect 4479 9475 4513 9476
rect 4483 9471 4484 9475
rect 4488 9471 4489 9475
rect 4493 9471 4494 9475
rect 4498 9471 4499 9475
rect 4503 9471 4504 9475
rect 4508 9471 4509 9475
rect 4529 9486 4530 9490
rect 4534 9486 4535 9490
rect 4539 9486 4540 9490
rect 4544 9486 4545 9490
rect 4549 9486 4550 9490
rect 4554 9486 4555 9490
rect 4525 9485 4559 9486
rect 4529 9481 4530 9485
rect 4534 9481 4535 9485
rect 4539 9481 4540 9485
rect 4544 9481 4545 9485
rect 4549 9481 4550 9485
rect 4554 9481 4555 9485
rect 4525 9480 4559 9481
rect 4529 9476 4530 9480
rect 4534 9476 4535 9480
rect 4539 9476 4540 9480
rect 4544 9476 4545 9480
rect 4549 9476 4550 9480
rect 4554 9476 4555 9480
rect 4525 9475 4559 9476
rect 4529 9471 4530 9475
rect 4534 9471 4535 9475
rect 4539 9471 4540 9475
rect 4544 9471 4545 9475
rect 4549 9471 4550 9475
rect 4554 9471 4555 9475
rect 4483 9457 4484 9461
rect 4488 9457 4489 9461
rect 4493 9457 4494 9461
rect 4498 9457 4499 9461
rect 4503 9457 4504 9461
rect 4508 9457 4509 9461
rect 4479 9456 4513 9457
rect 3769 9318 3775 9347
rect 3769 9216 3775 9314
rect 3769 8916 3775 9212
rect 3769 8816 3775 8912
rect 3769 8704 3775 8812
rect 3769 8674 3775 8700
rect 3769 8618 3775 8670
rect 3769 8588 3775 8614
rect 3769 8448 3775 8584
rect 3769 8369 3775 8444
rect 3769 8336 3775 8365
rect 3769 8234 3775 8332
rect 3769 7834 3775 8230
rect 3769 7722 3775 7830
rect 3769 7692 3775 7718
rect 3769 7636 3775 7688
rect 3769 7606 3775 7632
rect 3769 7466 3775 7602
rect 3769 7381 3775 7462
rect 3781 9021 3787 9452
rect 4483 9452 4484 9456
rect 4488 9452 4489 9456
rect 4493 9452 4494 9456
rect 4498 9452 4499 9456
rect 4503 9452 4504 9456
rect 4508 9452 4509 9456
rect 4479 9451 4513 9452
rect 4483 9447 4484 9451
rect 4488 9447 4489 9451
rect 4493 9447 4494 9451
rect 4498 9447 4499 9451
rect 4503 9447 4504 9451
rect 4508 9447 4509 9451
rect 4479 9446 4513 9447
rect 4483 9442 4484 9446
rect 4488 9442 4489 9446
rect 4493 9442 4494 9446
rect 4498 9442 4499 9446
rect 4503 9442 4504 9446
rect 4508 9442 4509 9446
rect 4529 9457 4530 9461
rect 4534 9457 4535 9461
rect 4539 9457 4540 9461
rect 4544 9457 4545 9461
rect 4549 9457 4550 9461
rect 4554 9457 4555 9461
rect 4525 9456 4559 9457
rect 4529 9452 4530 9456
rect 4534 9452 4535 9456
rect 4539 9452 4540 9456
rect 4544 9452 4545 9456
rect 4549 9452 4550 9456
rect 4554 9452 4555 9456
rect 4525 9451 4559 9452
rect 4529 9447 4530 9451
rect 4534 9447 4535 9451
rect 4539 9447 4540 9451
rect 4544 9447 4545 9451
rect 4549 9447 4550 9451
rect 4554 9447 4555 9451
rect 4525 9446 4559 9447
rect 4529 9442 4530 9446
rect 4534 9442 4535 9446
rect 4539 9442 4540 9446
rect 4544 9442 4545 9446
rect 4549 9442 4550 9446
rect 4554 9442 4555 9446
rect 4579 9355 5073 9786
rect 3803 9337 3806 9347
rect 3810 9307 3813 9316
rect 3826 9309 3829 9322
rect 3839 9294 3842 9347
rect 3906 9337 3909 9347
rect 3935 9337 3938 9347
rect 3846 9322 3850 9326
rect 3847 9307 3850 9316
rect 3802 9280 3805 9292
rect 3843 9290 3844 9294
rect 3853 9280 3856 9333
rect 3859 9313 3862 9318
rect 3868 9307 3871 9316
rect 3884 9309 3887 9322
rect 3905 9307 3908 9316
rect 3921 9316 3924 9318
rect 3921 9313 3928 9316
rect 3921 9307 3924 9313
rect 3942 9307 3945 9316
rect 3958 9309 3961 9322
rect 3904 9280 3907 9290
rect 3921 9273 3924 9303
rect 3971 9294 3974 9347
rect 4038 9337 4041 9347
rect 4067 9337 4070 9347
rect 3978 9322 3982 9326
rect 3979 9307 3982 9316
rect 3934 9280 3937 9292
rect 3975 9290 3976 9294
rect 3985 9280 3988 9333
rect 3991 9313 3994 9318
rect 4000 9307 4003 9316
rect 4016 9309 4019 9322
rect 4037 9307 4040 9316
rect 4053 9316 4056 9318
rect 4053 9313 4060 9316
rect 4053 9307 4056 9313
rect 4074 9307 4077 9316
rect 4090 9309 4093 9322
rect 4036 9280 4039 9290
rect 3921 9270 3973 9273
rect 3801 9250 3804 9263
rect 3827 9253 3830 9256
rect 3834 9250 3837 9263
rect 3851 9250 3854 9263
rect 3801 9201 3804 9216
rect 3815 9208 3818 9212
rect 3833 9201 3836 9216
rect 3852 9201 3855 9216
rect 3858 9215 3861 9256
rect 3874 9208 3877 9249
rect 3880 9216 3883 9256
rect 3899 9208 3902 9249
rect 3908 9250 3911 9263
rect 3924 9250 3927 9263
rect 3945 9253 3948 9256
rect 3952 9250 3955 9263
rect 3970 9259 3973 9270
rect 4053 9267 4056 9303
rect 4103 9294 4106 9347
rect 4170 9337 4173 9347
rect 4199 9337 4202 9347
rect 4110 9322 4114 9326
rect 4111 9307 4114 9316
rect 4066 9280 4069 9292
rect 4107 9290 4108 9294
rect 4117 9280 4120 9333
rect 4123 9313 4126 9318
rect 4132 9307 4135 9316
rect 4148 9309 4151 9322
rect 4169 9307 4172 9316
rect 4185 9316 4188 9318
rect 4185 9313 4192 9316
rect 4185 9307 4188 9313
rect 4206 9307 4209 9316
rect 4222 9309 4225 9322
rect 4168 9280 4171 9290
rect 4185 9273 4188 9295
rect 4235 9294 4238 9347
rect 4302 9337 4305 9347
rect 4242 9322 4246 9326
rect 4243 9307 4246 9316
rect 4198 9280 4201 9292
rect 4239 9290 4240 9294
rect 4249 9280 4252 9333
rect 4255 9313 4258 9318
rect 4264 9307 4267 9316
rect 4280 9309 4283 9322
rect 4301 9307 4304 9316
rect 4317 9316 4320 9318
rect 4826 9316 5086 9319
rect 4317 9313 4321 9316
rect 4317 9307 4320 9313
rect 4317 9299 4320 9303
rect 4300 9280 4303 9290
rect 4051 9262 4056 9267
rect 4113 9269 4188 9273
rect 3970 9256 4015 9259
rect 3970 9246 3973 9256
rect 3988 9243 4008 9246
rect 4005 9224 4008 9243
rect 3908 9201 3911 9216
rect 3923 9201 3926 9216
rect 3930 9208 3934 9211
rect 3951 9201 3954 9216
rect 3801 9182 3804 9197
rect 3815 9186 3818 9190
rect 3833 9182 3836 9197
rect 3852 9182 3855 9197
rect 3801 9135 3804 9148
rect 3827 9142 3830 9145
rect 3801 9118 3804 9131
rect 3811 9128 3815 9138
rect 3834 9135 3837 9148
rect 3851 9135 3854 9148
rect 3858 9142 3861 9183
rect 3874 9149 3877 9190
rect 3880 9142 3883 9182
rect 3899 9149 3902 9190
rect 3908 9182 3911 9197
rect 3923 9182 3926 9197
rect 3930 9187 3934 9190
rect 3951 9182 3954 9197
rect 3908 9135 3911 9148
rect 3827 9121 3830 9124
rect 3834 9118 3837 9131
rect 3851 9118 3854 9131
rect 3801 9069 3804 9084
rect 3815 9076 3818 9080
rect 3833 9069 3836 9084
rect 3852 9069 3855 9084
rect 3858 9083 3861 9124
rect 3874 9076 3877 9117
rect 3880 9084 3883 9124
rect 3899 9076 3902 9117
rect 3908 9118 3911 9131
rect 3924 9135 3927 9148
rect 3945 9142 3948 9145
rect 3952 9135 3955 9148
rect 4005 9148 4008 9220
rect 4016 9184 4019 9256
rect 4051 9259 4054 9262
rect 4051 9256 4096 9259
rect 4051 9246 4054 9256
rect 3924 9118 3927 9131
rect 3945 9121 3948 9124
rect 3952 9118 3955 9131
rect 4005 9114 4008 9144
rect 4016 9128 4019 9180
rect 4023 9168 4027 9234
rect 4011 9124 4015 9127
rect 4004 9111 4008 9114
rect 4005 9092 4008 9111
rect 3908 9069 3911 9084
rect 3923 9069 3926 9084
rect 3930 9076 3934 9079
rect 3951 9069 3954 9084
rect 3801 9050 3804 9065
rect 3815 9054 3818 9058
rect 3833 9050 3836 9065
rect 3852 9050 3855 9065
rect 3781 8718 3787 9017
rect 3801 9003 3804 9016
rect 3827 9010 3830 9013
rect 3801 8986 3804 8999
rect 3834 9003 3837 9016
rect 3851 9003 3854 9016
rect 3858 9010 3861 9051
rect 3874 9017 3877 9058
rect 3880 9010 3883 9050
rect 3899 9017 3902 9058
rect 3908 9050 3911 9065
rect 3923 9050 3926 9065
rect 3930 9055 3934 9058
rect 3951 9050 3954 9065
rect 3908 9003 3911 9016
rect 3827 8989 3830 8992
rect 3834 8986 3837 8999
rect 3851 8986 3854 8999
rect 3801 8937 3804 8952
rect 3815 8944 3818 8948
rect 3833 8937 3836 8952
rect 3852 8937 3855 8952
rect 3858 8951 3861 8992
rect 3874 8944 3877 8985
rect 3880 8952 3883 8992
rect 3899 8944 3902 8985
rect 3908 8986 3911 8999
rect 3924 9003 3927 9016
rect 3945 9010 3948 9013
rect 3952 9003 3955 9016
rect 4005 9017 4008 9088
rect 4016 9053 4019 9124
rect 3924 8986 3927 8999
rect 3945 8989 3948 8992
rect 3952 8986 3955 8999
rect 4005 8960 4008 9013
rect 4016 8996 4019 9049
rect 4023 9037 4027 9102
rect 4011 8992 4015 8995
rect 4054 8995 4057 9246
rect 4069 9243 4089 9246
rect 4086 9224 4089 9243
rect 4086 9148 4089 9220
rect 4097 9184 4100 9256
rect 4104 9168 4108 9234
rect 4113 9135 4116 9269
rect 4317 9266 4320 9295
rect 4141 9263 4248 9266
rect 4075 9131 4116 9135
rect 4075 9127 4078 9131
rect 4075 9124 4120 9127
rect 4075 9114 4078 9124
rect 4093 9111 4113 9114
rect 4075 9109 4078 9110
rect 4110 9092 4113 9111
rect 4110 9017 4113 9088
rect 4121 9053 4124 9124
rect 4128 9037 4132 9102
rect 3908 8937 3911 8952
rect 3923 8937 3926 8952
rect 3930 8944 3934 8947
rect 3951 8937 3954 8952
rect 3801 8918 3804 8933
rect 3815 8922 3818 8926
rect 3833 8918 3836 8933
rect 3852 8918 3855 8933
rect 3801 8871 3804 8884
rect 3827 8878 3830 8881
rect 3801 8854 3804 8867
rect 3834 8871 3837 8884
rect 3851 8871 3854 8884
rect 3858 8878 3861 8919
rect 3874 8885 3877 8926
rect 3880 8878 3883 8918
rect 3899 8885 3902 8926
rect 3908 8918 3911 8933
rect 3923 8918 3926 8933
rect 3930 8923 3934 8926
rect 3951 8918 3954 8933
rect 3908 8871 3911 8884
rect 3827 8857 3830 8860
rect 3834 8854 3837 8867
rect 3851 8854 3854 8867
rect 3801 8805 3804 8820
rect 3815 8812 3818 8816
rect 3801 8786 3804 8801
rect 3824 8798 3828 8808
rect 3833 8805 3836 8820
rect 3852 8805 3855 8820
rect 3858 8819 3861 8860
rect 3874 8812 3877 8853
rect 3880 8820 3883 8860
rect 3899 8812 3902 8853
rect 3908 8854 3911 8867
rect 3924 8871 3927 8884
rect 3945 8878 3948 8881
rect 3952 8871 3955 8884
rect 4005 8882 4008 8956
rect 4016 8918 4019 8992
rect 4051 8992 4096 8995
rect 4051 8982 4054 8992
rect 4069 8979 4089 8982
rect 3924 8854 3927 8867
rect 3945 8857 3948 8860
rect 3952 8854 3955 8867
rect 4005 8828 4008 8878
rect 4016 8864 4019 8914
rect 4023 8902 4027 8970
rect 4086 8960 4089 8979
rect 4086 8882 4089 8956
rect 4097 8918 4100 8992
rect 4141 8995 4144 9263
rect 4252 9263 4320 9266
rect 4826 9062 4829 9316
rect 5083 9062 5086 9316
rect 4483 9056 4484 9060
rect 4488 9056 4489 9060
rect 4493 9056 4494 9060
rect 4498 9056 4499 9060
rect 4503 9056 4504 9060
rect 4508 9056 4509 9060
rect 4479 9055 4513 9056
rect 4483 9051 4484 9055
rect 4488 9051 4489 9055
rect 4493 9051 4494 9055
rect 4498 9051 4499 9055
rect 4503 9051 4504 9055
rect 4508 9051 4509 9055
rect 4479 9050 4513 9051
rect 4483 9046 4484 9050
rect 4488 9046 4489 9050
rect 4493 9046 4494 9050
rect 4498 9046 4499 9050
rect 4503 9046 4504 9050
rect 4508 9046 4509 9050
rect 4479 9045 4513 9046
rect 4483 9041 4484 9045
rect 4488 9041 4489 9045
rect 4493 9041 4494 9045
rect 4498 9041 4499 9045
rect 4503 9041 4504 9045
rect 4508 9041 4509 9045
rect 4529 9056 4530 9060
rect 4534 9056 4535 9060
rect 4539 9056 4540 9060
rect 4544 9056 4545 9060
rect 4549 9056 4550 9060
rect 4554 9056 4555 9060
rect 4826 9059 5086 9062
rect 4525 9055 4559 9056
rect 4529 9051 4530 9055
rect 4534 9051 4535 9055
rect 4539 9051 4540 9055
rect 4544 9051 4545 9055
rect 4549 9051 4550 9055
rect 4554 9051 4555 9055
rect 4525 9050 4559 9051
rect 4529 9046 4530 9050
rect 4534 9046 4535 9050
rect 4539 9046 4540 9050
rect 4544 9046 4545 9050
rect 4549 9046 4550 9050
rect 4554 9046 4555 9050
rect 4525 9045 4559 9046
rect 4529 9041 4530 9045
rect 4534 9041 4535 9045
rect 4539 9041 4540 9045
rect 4544 9041 4545 9045
rect 4549 9041 4550 9045
rect 4554 9041 4555 9045
rect 4826 9007 5086 9010
rect 4141 8992 4186 8995
rect 4141 8982 4144 8992
rect 4159 8979 4179 8982
rect 4104 8902 4108 8970
rect 4176 8960 4179 8979
rect 4176 8882 4179 8956
rect 4187 8918 4190 8992
rect 4194 8902 4198 8970
rect 4011 8860 4015 8863
rect 3908 8805 3911 8820
rect 3923 8805 3926 8820
rect 3930 8812 3934 8815
rect 3951 8805 3954 8820
rect 3815 8790 3818 8794
rect 3833 8786 3836 8801
rect 3852 8786 3855 8801
rect 3801 8739 3804 8752
rect 3827 8746 3830 8749
rect 3809 8732 3813 8742
rect 3834 8739 3837 8752
rect 3851 8739 3854 8752
rect 3858 8746 3861 8787
rect 3874 8753 3877 8794
rect 3880 8746 3883 8786
rect 3899 8753 3902 8794
rect 3908 8786 3911 8801
rect 3923 8786 3926 8801
rect 3930 8791 3934 8794
rect 3951 8786 3954 8801
rect 3908 8739 3911 8752
rect 3924 8739 3927 8752
rect 3945 8746 3948 8749
rect 3952 8739 3955 8752
rect 4005 8746 4008 8824
rect 4016 8782 4019 8860
rect 4023 8766 4027 8838
rect 4035 8739 4039 8752
rect 4044 8732 4047 8742
rect 4054 8725 4057 8794
rect 4076 8790 4079 8794
rect 4094 8786 4097 8801
rect 4113 8786 4116 8801
rect 4061 8739 4065 8752
rect 4088 8746 4091 8749
rect 4095 8739 4098 8752
rect 4112 8739 4115 8752
rect 4119 8746 4122 8787
rect 4135 8753 4138 8794
rect 4141 8746 4144 8786
rect 4160 8753 4163 8794
rect 4169 8786 4172 8801
rect 4184 8786 4187 8801
rect 4191 8791 4195 8794
rect 4212 8786 4215 8801
rect 4169 8739 4172 8752
rect 4185 8739 4188 8752
rect 4206 8746 4209 8749
rect 4213 8739 4216 8752
rect 4229 8733 4233 8969
rect 4826 8753 4829 9007
rect 5083 8753 5086 9007
rect 4483 8747 4484 8751
rect 4488 8747 4489 8751
rect 4493 8747 4494 8751
rect 4498 8747 4499 8751
rect 4503 8747 4504 8751
rect 4508 8747 4509 8751
rect 4479 8746 4513 8747
rect 4483 8742 4484 8746
rect 4488 8742 4489 8746
rect 4493 8742 4494 8746
rect 4498 8742 4499 8746
rect 4503 8742 4504 8746
rect 4508 8742 4509 8746
rect 4479 8741 4513 8742
rect 4483 8737 4484 8741
rect 4488 8737 4489 8741
rect 4493 8737 4494 8741
rect 4498 8737 4499 8741
rect 4503 8737 4504 8741
rect 4508 8737 4509 8741
rect 4479 8736 4513 8737
rect 4483 8732 4484 8736
rect 4488 8732 4489 8736
rect 4493 8732 4494 8736
rect 4498 8732 4499 8736
rect 4503 8732 4504 8736
rect 4508 8732 4509 8736
rect 4529 8747 4530 8751
rect 4534 8747 4535 8751
rect 4539 8747 4540 8751
rect 4544 8747 4545 8751
rect 4549 8747 4550 8751
rect 4554 8747 4555 8751
rect 4826 8750 5086 8753
rect 4525 8746 4559 8747
rect 4529 8742 4530 8746
rect 4534 8742 4535 8746
rect 4539 8742 4540 8746
rect 4544 8742 4545 8746
rect 4549 8742 4550 8746
rect 4554 8742 4555 8746
rect 4525 8741 4559 8742
rect 4529 8737 4530 8741
rect 4534 8737 4535 8741
rect 4539 8737 4540 8741
rect 4544 8737 4545 8741
rect 4549 8737 4550 8741
rect 4554 8737 4555 8741
rect 4525 8736 4559 8737
rect 4529 8732 4530 8736
rect 4534 8732 4535 8736
rect 4539 8732 4540 8736
rect 4544 8732 4545 8736
rect 4549 8732 4550 8736
rect 4554 8732 4555 8736
rect 4222 8721 4223 8724
rect 3781 7736 3787 8714
rect 4087 8611 4091 8693
rect 4102 8690 4105 8700
rect 4109 8660 4112 8669
rect 4125 8662 4128 8675
rect 4138 8647 4141 8700
rect 4205 8690 4208 8700
rect 4145 8675 4149 8679
rect 4146 8660 4149 8669
rect 4101 8633 4104 8645
rect 4142 8643 4143 8647
rect 4152 8633 4155 8686
rect 4220 8675 4223 8721
rect 4158 8666 4161 8671
rect 4167 8660 4170 8669
rect 4183 8662 4186 8675
rect 4204 8660 4207 8669
rect 4220 8660 4223 8669
rect 4203 8633 4206 8643
rect 4220 8626 4223 8656
rect 4095 8584 4098 8621
rect 4102 8604 4105 8614
rect 4109 8574 4112 8583
rect 4125 8576 4128 8589
rect 4138 8561 4141 8614
rect 4205 8604 4208 8614
rect 4145 8589 4149 8593
rect 4146 8574 4149 8583
rect 4101 8547 4104 8559
rect 4142 8557 4143 8561
rect 4152 8547 4155 8600
rect 4158 8580 4161 8585
rect 4167 8574 4170 8583
rect 4183 8576 4186 8589
rect 4204 8574 4207 8583
rect 4220 8584 4223 8585
rect 4241 8587 4245 8729
rect 4826 8698 5086 8701
rect 4220 8579 4223 8580
rect 4203 8547 4206 8557
rect 4241 8485 4245 8567
rect 4826 8444 4829 8698
rect 5083 8444 5086 8698
rect 4483 8438 4484 8442
rect 4488 8438 4489 8442
rect 4493 8438 4494 8442
rect 4498 8438 4499 8442
rect 4503 8438 4504 8442
rect 4508 8438 4509 8442
rect 4479 8437 4513 8438
rect 4483 8433 4484 8437
rect 4488 8433 4489 8437
rect 4493 8433 4494 8437
rect 4498 8433 4499 8437
rect 4503 8433 4504 8437
rect 4508 8433 4509 8437
rect 4479 8432 4513 8433
rect 4483 8428 4484 8432
rect 4488 8428 4489 8432
rect 4493 8428 4494 8432
rect 4498 8428 4499 8432
rect 4503 8428 4504 8432
rect 4508 8428 4509 8432
rect 4479 8427 4513 8428
rect 4483 8423 4484 8427
rect 4488 8423 4489 8427
rect 4493 8423 4494 8427
rect 4498 8423 4499 8427
rect 4503 8423 4504 8427
rect 4508 8423 4509 8427
rect 4529 8438 4530 8442
rect 4534 8438 4535 8442
rect 4539 8438 4540 8442
rect 4544 8438 4545 8442
rect 4549 8438 4550 8442
rect 4554 8438 4555 8442
rect 4826 8441 5086 8444
rect 4525 8437 4559 8438
rect 4529 8433 4530 8437
rect 4534 8433 4535 8437
rect 4539 8433 4540 8437
rect 4544 8433 4545 8437
rect 4549 8433 4550 8437
rect 4554 8433 4555 8437
rect 4525 8432 4559 8433
rect 4529 8428 4530 8432
rect 4534 8428 4535 8432
rect 4539 8428 4540 8432
rect 4544 8428 4545 8432
rect 4549 8428 4550 8432
rect 4554 8428 4555 8432
rect 4525 8427 4559 8428
rect 4529 8423 4530 8427
rect 4534 8423 4535 8427
rect 4539 8423 4540 8427
rect 4544 8423 4545 8427
rect 4549 8423 4550 8427
rect 4554 8423 4555 8427
rect 4826 8389 5086 8392
rect 3803 8355 3806 8365
rect 3810 8325 3813 8334
rect 3826 8327 3829 8340
rect 3839 8312 3842 8365
rect 3906 8355 3909 8365
rect 3935 8355 3938 8365
rect 3846 8340 3850 8344
rect 3847 8325 3850 8334
rect 3802 8298 3805 8310
rect 3843 8308 3844 8312
rect 3853 8298 3856 8351
rect 3859 8331 3862 8336
rect 3868 8325 3871 8334
rect 3884 8327 3887 8340
rect 3905 8325 3908 8334
rect 3921 8334 3924 8336
rect 3921 8331 3928 8334
rect 3921 8325 3924 8331
rect 3942 8325 3945 8334
rect 3958 8327 3961 8340
rect 3904 8298 3907 8308
rect 3921 8291 3924 8321
rect 3971 8312 3974 8365
rect 4038 8355 4041 8365
rect 4067 8355 4070 8365
rect 3978 8340 3982 8344
rect 3979 8325 3982 8334
rect 3934 8298 3937 8310
rect 3975 8308 3976 8312
rect 3985 8298 3988 8351
rect 3991 8331 3994 8336
rect 4000 8325 4003 8334
rect 4016 8327 4019 8340
rect 4037 8325 4040 8334
rect 4053 8334 4056 8336
rect 4053 8331 4060 8334
rect 4053 8325 4056 8331
rect 4074 8325 4077 8334
rect 4090 8327 4093 8340
rect 4036 8298 4039 8308
rect 3921 8288 3973 8291
rect 3801 8268 3804 8281
rect 3827 8271 3830 8274
rect 3834 8268 3837 8281
rect 3851 8268 3854 8281
rect 3801 8219 3804 8234
rect 3815 8226 3818 8230
rect 3833 8219 3836 8234
rect 3852 8219 3855 8234
rect 3858 8233 3861 8274
rect 3874 8226 3877 8267
rect 3880 8234 3883 8274
rect 3899 8226 3902 8267
rect 3908 8268 3911 8281
rect 3924 8268 3927 8281
rect 3945 8271 3948 8274
rect 3952 8268 3955 8281
rect 3970 8277 3973 8288
rect 4053 8285 4056 8321
rect 4103 8312 4106 8365
rect 4170 8355 4173 8365
rect 4199 8355 4202 8365
rect 4110 8340 4114 8344
rect 4111 8325 4114 8334
rect 4066 8298 4069 8310
rect 4107 8308 4108 8312
rect 4117 8298 4120 8351
rect 4123 8331 4126 8336
rect 4132 8325 4135 8334
rect 4148 8327 4151 8340
rect 4169 8325 4172 8334
rect 4185 8334 4188 8336
rect 4185 8331 4192 8334
rect 4185 8325 4188 8331
rect 4206 8325 4209 8334
rect 4222 8327 4225 8340
rect 4168 8298 4171 8308
rect 4185 8291 4188 8313
rect 4235 8312 4238 8365
rect 4302 8355 4305 8365
rect 4242 8340 4246 8344
rect 4243 8325 4246 8334
rect 4198 8298 4201 8310
rect 4239 8308 4240 8312
rect 4249 8298 4252 8351
rect 4255 8331 4258 8336
rect 4264 8325 4267 8334
rect 4280 8327 4283 8340
rect 4301 8325 4304 8334
rect 4317 8334 4320 8336
rect 4317 8331 4321 8334
rect 4317 8325 4320 8331
rect 4317 8317 4320 8321
rect 4300 8298 4303 8308
rect 4051 8280 4056 8285
rect 4113 8287 4188 8291
rect 3970 8274 4015 8277
rect 3970 8264 3973 8274
rect 3988 8261 4008 8264
rect 4005 8242 4008 8261
rect 3908 8219 3911 8234
rect 3923 8219 3926 8234
rect 3930 8226 3934 8229
rect 3951 8219 3954 8234
rect 3801 8200 3804 8215
rect 3815 8204 3818 8208
rect 3833 8200 3836 8215
rect 3852 8200 3855 8215
rect 3801 8153 3804 8166
rect 3827 8160 3830 8163
rect 3801 8136 3804 8149
rect 3811 8146 3815 8156
rect 3834 8153 3837 8166
rect 3851 8153 3854 8166
rect 3858 8160 3861 8201
rect 3874 8167 3877 8208
rect 3880 8160 3883 8200
rect 3899 8167 3902 8208
rect 3908 8200 3911 8215
rect 3923 8200 3926 8215
rect 3930 8205 3934 8208
rect 3951 8200 3954 8215
rect 3908 8153 3911 8166
rect 3827 8139 3830 8142
rect 3834 8136 3837 8149
rect 3851 8136 3854 8149
rect 3801 8087 3804 8102
rect 3815 8094 3818 8098
rect 3833 8087 3836 8102
rect 3852 8087 3855 8102
rect 3858 8101 3861 8142
rect 3874 8094 3877 8135
rect 3880 8102 3883 8142
rect 3899 8094 3902 8135
rect 3908 8136 3911 8149
rect 3924 8153 3927 8166
rect 3945 8160 3948 8163
rect 3952 8153 3955 8166
rect 4005 8166 4008 8238
rect 4016 8202 4019 8274
rect 4051 8277 4054 8280
rect 4051 8274 4096 8277
rect 4051 8264 4054 8274
rect 3924 8136 3927 8149
rect 3945 8139 3948 8142
rect 3952 8136 3955 8149
rect 4005 8132 4008 8162
rect 4016 8146 4019 8198
rect 4023 8186 4027 8252
rect 4011 8142 4015 8145
rect 4004 8129 4008 8132
rect 4005 8110 4008 8129
rect 3908 8087 3911 8102
rect 3923 8087 3926 8102
rect 3930 8094 3934 8097
rect 3951 8087 3954 8102
rect 3801 8068 3804 8083
rect 3815 8072 3818 8076
rect 3833 8068 3836 8083
rect 3852 8068 3855 8083
rect 3801 8021 3804 8034
rect 3827 8028 3830 8031
rect 3801 8004 3804 8017
rect 3834 8021 3837 8034
rect 3851 8021 3854 8034
rect 3858 8028 3861 8069
rect 3874 8035 3877 8076
rect 3880 8028 3883 8068
rect 3899 8035 3902 8076
rect 3908 8068 3911 8083
rect 3923 8068 3926 8083
rect 3930 8073 3934 8076
rect 3951 8068 3954 8083
rect 3908 8021 3911 8034
rect 3827 8007 3830 8010
rect 3834 8004 3837 8017
rect 3851 8004 3854 8017
rect 3801 7955 3804 7970
rect 3815 7962 3818 7966
rect 3833 7955 3836 7970
rect 3852 7955 3855 7970
rect 3858 7969 3861 8010
rect 3874 7962 3877 8003
rect 3880 7970 3883 8010
rect 3899 7962 3902 8003
rect 3908 8004 3911 8017
rect 3924 8021 3927 8034
rect 3945 8028 3948 8031
rect 3952 8021 3955 8034
rect 4005 8035 4008 8106
rect 4016 8071 4019 8142
rect 3924 8004 3927 8017
rect 3945 8007 3948 8010
rect 3952 8004 3955 8017
rect 4005 7978 4008 8031
rect 4016 8014 4019 8067
rect 4023 8055 4027 8120
rect 4011 8010 4015 8013
rect 4054 8013 4057 8264
rect 4069 8261 4089 8264
rect 4086 8242 4089 8261
rect 4086 8166 4089 8238
rect 4097 8202 4100 8274
rect 4104 8186 4108 8252
rect 4113 8153 4116 8287
rect 4317 8284 4320 8313
rect 4141 8281 4248 8284
rect 4075 8149 4116 8153
rect 4075 8145 4078 8149
rect 4075 8142 4120 8145
rect 4075 8132 4078 8142
rect 4093 8129 4113 8132
rect 4075 8127 4078 8128
rect 4110 8110 4113 8129
rect 4110 8035 4113 8106
rect 4121 8071 4124 8142
rect 4128 8055 4132 8120
rect 3908 7955 3911 7970
rect 3923 7955 3926 7970
rect 3930 7962 3934 7965
rect 3951 7955 3954 7970
rect 3801 7936 3804 7951
rect 3815 7940 3818 7944
rect 3833 7936 3836 7951
rect 3852 7936 3855 7951
rect 3801 7889 3804 7902
rect 3827 7896 3830 7899
rect 3801 7872 3804 7885
rect 3834 7889 3837 7902
rect 3851 7889 3854 7902
rect 3858 7896 3861 7937
rect 3874 7903 3877 7944
rect 3880 7896 3883 7936
rect 3899 7903 3902 7944
rect 3908 7936 3911 7951
rect 3923 7936 3926 7951
rect 3930 7941 3934 7944
rect 3951 7936 3954 7951
rect 3908 7889 3911 7902
rect 3827 7875 3830 7878
rect 3834 7872 3837 7885
rect 3851 7872 3854 7885
rect 3801 7823 3804 7838
rect 3815 7830 3818 7834
rect 3801 7804 3804 7819
rect 3824 7816 3828 7826
rect 3833 7823 3836 7838
rect 3852 7823 3855 7838
rect 3858 7837 3861 7878
rect 3874 7830 3877 7871
rect 3880 7838 3883 7878
rect 3899 7830 3902 7871
rect 3908 7872 3911 7885
rect 3924 7889 3927 7902
rect 3945 7896 3948 7899
rect 3952 7889 3955 7902
rect 4005 7900 4008 7974
rect 4016 7936 4019 8010
rect 4051 8010 4096 8013
rect 4051 8000 4054 8010
rect 4069 7997 4089 8000
rect 3924 7872 3927 7885
rect 3945 7875 3948 7878
rect 3952 7872 3955 7885
rect 4005 7846 4008 7896
rect 4016 7882 4019 7932
rect 4023 7920 4027 7988
rect 4086 7978 4089 7997
rect 4086 7900 4089 7974
rect 4097 7936 4100 8010
rect 4141 8013 4144 8281
rect 4252 8281 4320 8284
rect 4826 8135 4829 8389
rect 5083 8135 5086 8389
rect 4483 8129 4484 8133
rect 4488 8129 4489 8133
rect 4493 8129 4494 8133
rect 4498 8129 4499 8133
rect 4503 8129 4504 8133
rect 4508 8129 4509 8133
rect 4479 8128 4513 8129
rect 4483 8124 4484 8128
rect 4488 8124 4489 8128
rect 4493 8124 4494 8128
rect 4498 8124 4499 8128
rect 4503 8124 4504 8128
rect 4508 8124 4509 8128
rect 4479 8123 4513 8124
rect 4483 8119 4484 8123
rect 4488 8119 4489 8123
rect 4493 8119 4494 8123
rect 4498 8119 4499 8123
rect 4503 8119 4504 8123
rect 4508 8119 4509 8123
rect 4479 8118 4513 8119
rect 4483 8114 4484 8118
rect 4488 8114 4489 8118
rect 4493 8114 4494 8118
rect 4498 8114 4499 8118
rect 4503 8114 4504 8118
rect 4508 8114 4509 8118
rect 4529 8129 4530 8133
rect 4534 8129 4535 8133
rect 4539 8129 4540 8133
rect 4544 8129 4545 8133
rect 4549 8129 4550 8133
rect 4554 8129 4555 8133
rect 4826 8132 5086 8135
rect 4525 8128 4559 8129
rect 4529 8124 4530 8128
rect 4534 8124 4535 8128
rect 4539 8124 4540 8128
rect 4544 8124 4545 8128
rect 4549 8124 4550 8128
rect 4554 8124 4555 8128
rect 4525 8123 4559 8124
rect 4529 8119 4530 8123
rect 4534 8119 4535 8123
rect 4539 8119 4540 8123
rect 4544 8119 4545 8123
rect 4549 8119 4550 8123
rect 4554 8119 4555 8123
rect 4525 8118 4559 8119
rect 4529 8114 4530 8118
rect 4534 8114 4535 8118
rect 4539 8114 4540 8118
rect 4544 8114 4545 8118
rect 4549 8114 4550 8118
rect 4554 8114 4555 8118
rect 4483 8098 4484 8102
rect 4488 8098 4489 8102
rect 4493 8098 4494 8102
rect 4498 8098 4499 8102
rect 4503 8098 4504 8102
rect 4508 8098 4509 8102
rect 4479 8097 4513 8098
rect 4483 8093 4484 8097
rect 4488 8093 4489 8097
rect 4493 8093 4494 8097
rect 4498 8093 4499 8097
rect 4503 8093 4504 8097
rect 4508 8093 4509 8097
rect 4479 8092 4513 8093
rect 4483 8088 4484 8092
rect 4488 8088 4489 8092
rect 4493 8088 4494 8092
rect 4498 8088 4499 8092
rect 4503 8088 4504 8092
rect 4508 8088 4509 8092
rect 4479 8087 4513 8088
rect 4483 8083 4484 8087
rect 4488 8083 4489 8087
rect 4493 8083 4494 8087
rect 4498 8083 4499 8087
rect 4503 8083 4504 8087
rect 4508 8083 4509 8087
rect 4529 8098 4530 8102
rect 4534 8098 4535 8102
rect 4539 8098 4540 8102
rect 4544 8098 4545 8102
rect 4549 8098 4550 8102
rect 4554 8098 4555 8102
rect 4525 8097 4559 8098
rect 4529 8093 4530 8097
rect 4534 8093 4535 8097
rect 4539 8093 4540 8097
rect 4544 8093 4545 8097
rect 4549 8093 4550 8097
rect 4554 8093 4555 8097
rect 4525 8092 4559 8093
rect 4529 8088 4530 8092
rect 4534 8088 4535 8092
rect 4539 8088 4540 8092
rect 4544 8088 4545 8092
rect 4549 8088 4550 8092
rect 4554 8088 4555 8092
rect 4525 8087 4559 8088
rect 4529 8083 4530 8087
rect 4534 8083 4535 8087
rect 4539 8083 4540 8087
rect 4544 8083 4545 8087
rect 4549 8083 4550 8087
rect 4554 8083 4555 8087
rect 4826 8081 5086 8084
rect 4494 8078 4515 8080
rect 4494 8074 4496 8078
rect 4500 8074 4501 8078
rect 4505 8074 4506 8078
rect 4510 8074 4511 8078
rect 4494 8073 4515 8074
rect 4494 8069 4496 8073
rect 4500 8069 4501 8073
rect 4505 8069 4506 8073
rect 4510 8069 4511 8073
rect 4494 8068 4515 8069
rect 4494 8064 4496 8068
rect 4500 8064 4501 8068
rect 4505 8064 4506 8068
rect 4510 8064 4511 8068
rect 4494 8063 4515 8064
rect 4494 8059 4496 8063
rect 4500 8059 4501 8063
rect 4505 8059 4506 8063
rect 4510 8059 4511 8063
rect 4494 8058 4515 8059
rect 4494 8054 4496 8058
rect 4500 8054 4501 8058
rect 4505 8054 4506 8058
rect 4510 8054 4511 8058
rect 4494 8053 4515 8054
rect 4494 8049 4496 8053
rect 4500 8049 4501 8053
rect 4505 8049 4506 8053
rect 4510 8049 4511 8053
rect 4494 8048 4515 8049
rect 4494 8044 4496 8048
rect 4500 8044 4501 8048
rect 4505 8044 4506 8048
rect 4510 8044 4511 8048
rect 4494 8043 4515 8044
rect 4494 8039 4496 8043
rect 4500 8039 4501 8043
rect 4505 8039 4506 8043
rect 4510 8039 4511 8043
rect 4494 8038 4515 8039
rect 4494 8034 4496 8038
rect 4500 8034 4501 8038
rect 4505 8034 4506 8038
rect 4510 8034 4511 8038
rect 4494 8033 4515 8034
rect 4494 8029 4496 8033
rect 4500 8029 4501 8033
rect 4505 8029 4506 8033
rect 4510 8029 4511 8033
rect 4494 8028 4515 8029
rect 4494 8024 4496 8028
rect 4500 8024 4501 8028
rect 4505 8024 4506 8028
rect 4510 8024 4511 8028
rect 4141 8010 4186 8013
rect 4141 8000 4144 8010
rect 4159 7997 4179 8000
rect 4104 7920 4108 7988
rect 4176 7978 4179 7997
rect 4176 7900 4179 7974
rect 4187 7936 4190 8010
rect 4194 7920 4198 7988
rect 4229 7959 4233 7987
rect 4578 7982 4590 7986
rect 4594 7982 4606 7986
rect 4610 7982 4622 7986
rect 4626 7982 4645 7986
rect 4649 7982 4661 7986
rect 4665 7982 4688 7986
rect 4692 7982 4704 7986
rect 4708 7982 4729 7986
rect 4733 7982 4745 7986
rect 4657 7963 4717 7965
rect 4229 7948 4236 7959
rect 4657 7954 4659 7963
rect 4667 7954 4703 7963
rect 4711 7954 4717 7963
rect 4657 7952 4717 7954
rect 4011 7878 4015 7881
rect 3908 7823 3911 7838
rect 3923 7823 3926 7838
rect 3930 7830 3934 7833
rect 3951 7823 3954 7838
rect 3815 7808 3818 7812
rect 3833 7804 3836 7819
rect 3852 7804 3855 7819
rect 3801 7757 3804 7770
rect 3827 7764 3830 7767
rect 3809 7750 3813 7760
rect 3834 7757 3837 7770
rect 3851 7757 3854 7770
rect 3858 7764 3861 7805
rect 3874 7771 3877 7812
rect 3880 7764 3883 7804
rect 3899 7771 3902 7812
rect 3908 7804 3911 7819
rect 3923 7804 3926 7819
rect 3930 7809 3934 7812
rect 3951 7804 3954 7819
rect 3908 7757 3911 7770
rect 3924 7757 3927 7770
rect 3945 7764 3948 7767
rect 3952 7757 3955 7770
rect 4005 7764 4008 7842
rect 4016 7800 4019 7878
rect 4023 7784 4027 7856
rect 4035 7757 4039 7770
rect 4044 7750 4047 7760
rect 4054 7743 4057 7812
rect 4076 7808 4079 7812
rect 4094 7804 4097 7819
rect 4113 7804 4116 7819
rect 4061 7757 4065 7770
rect 4088 7764 4091 7767
rect 4095 7757 4098 7770
rect 4112 7757 4115 7770
rect 4119 7764 4122 7805
rect 4135 7771 4138 7812
rect 4141 7764 4144 7804
rect 4160 7771 4163 7812
rect 4169 7804 4172 7819
rect 4184 7804 4187 7819
rect 4191 7809 4195 7812
rect 4212 7804 4215 7819
rect 4169 7757 4172 7770
rect 4185 7757 4188 7770
rect 4206 7764 4209 7767
rect 4213 7757 4216 7770
rect 4229 7751 4233 7948
rect 4222 7739 4223 7742
rect 3781 7381 3787 7732
rect 4087 7629 4091 7711
rect 4102 7708 4105 7718
rect 4109 7678 4112 7687
rect 4125 7680 4128 7693
rect 4138 7665 4141 7718
rect 4205 7708 4208 7718
rect 4145 7693 4149 7697
rect 4146 7678 4149 7687
rect 4101 7651 4104 7663
rect 4142 7661 4143 7665
rect 4152 7651 4155 7704
rect 4220 7693 4223 7739
rect 4158 7684 4161 7689
rect 4167 7678 4170 7687
rect 4183 7680 4186 7693
rect 4204 7678 4207 7687
rect 4220 7678 4223 7687
rect 4203 7651 4206 7661
rect 4220 7644 4223 7674
rect 4095 7602 4098 7639
rect 4102 7622 4105 7632
rect 4109 7592 4112 7601
rect 4125 7594 4128 7607
rect 4138 7579 4141 7632
rect 4205 7622 4208 7632
rect 4145 7607 4149 7611
rect 4146 7592 4149 7601
rect 4101 7565 4104 7577
rect 4142 7575 4143 7579
rect 4152 7565 4155 7618
rect 4158 7598 4161 7603
rect 4167 7592 4170 7601
rect 4183 7594 4186 7607
rect 4204 7592 4207 7601
rect 4220 7602 4223 7603
rect 4241 7605 4245 7747
rect 4220 7597 4223 7598
rect 4203 7565 4206 7575
rect 4241 7503 4245 7585
rect 4360 7503 4369 7950
rect 4578 7924 4590 7928
rect 4594 7924 4606 7928
rect 4610 7924 4622 7928
rect 4626 7924 4645 7928
rect 4649 7924 4661 7928
rect 4665 7924 4688 7928
rect 4692 7924 4704 7928
rect 4708 7924 4729 7928
rect 4733 7924 4745 7928
rect 4527 7824 4529 7828
rect 4533 7824 4534 7828
rect 4538 7824 4539 7828
rect 4543 7824 4544 7828
rect 4548 7824 4549 7828
rect 4553 7824 4554 7828
rect 4558 7824 4559 7828
rect 4563 7824 4564 7828
rect 4568 7824 4569 7828
rect 4573 7824 4574 7828
rect 4578 7824 4579 7828
rect 4583 7824 4584 7828
rect 4588 7824 4589 7828
rect 4593 7824 4595 7828
rect 4826 7827 4829 8081
rect 5083 7827 5086 8081
rect 4826 7824 5086 7827
rect 4527 7823 4595 7824
rect 4527 7819 4529 7823
rect 4533 7819 4534 7823
rect 4538 7819 4539 7823
rect 4543 7819 4544 7823
rect 4548 7819 4549 7823
rect 4553 7819 4554 7823
rect 4558 7819 4559 7823
rect 4563 7819 4564 7823
rect 4568 7819 4569 7823
rect 4573 7819 4574 7823
rect 4578 7819 4579 7823
rect 4583 7819 4584 7823
rect 4588 7819 4589 7823
rect 4593 7819 4595 7823
rect 4527 7818 4595 7819
rect 4527 7814 4529 7818
rect 4533 7814 4534 7818
rect 4538 7814 4539 7818
rect 4543 7814 4544 7818
rect 4548 7814 4549 7818
rect 4553 7814 4554 7818
rect 4558 7814 4559 7818
rect 4563 7814 4564 7818
rect 4568 7814 4569 7818
rect 4573 7814 4574 7818
rect 4578 7814 4579 7818
rect 4583 7814 4584 7818
rect 4588 7814 4589 7818
rect 4593 7814 4595 7818
rect 4527 7813 4595 7814
rect 4527 7809 4529 7813
rect 4533 7809 4534 7813
rect 4538 7809 4539 7813
rect 4543 7809 4544 7813
rect 4548 7809 4549 7813
rect 4553 7809 4554 7813
rect 4558 7809 4559 7813
rect 4563 7809 4564 7813
rect 4568 7809 4569 7813
rect 4573 7809 4574 7813
rect 4578 7809 4579 7813
rect 4583 7809 4584 7813
rect 4588 7809 4589 7813
rect 4593 7809 4595 7813
rect 4527 7807 4595 7809
rect 4483 7789 4484 7793
rect 4488 7789 4489 7793
rect 4493 7789 4494 7793
rect 4498 7789 4499 7793
rect 4503 7789 4504 7793
rect 4508 7789 4509 7793
rect 4479 7788 4513 7789
rect 4483 7784 4484 7788
rect 4488 7784 4489 7788
rect 4493 7784 4494 7788
rect 4498 7784 4499 7788
rect 4503 7784 4504 7788
rect 4508 7784 4509 7788
rect 4479 7783 4513 7784
rect 4483 7779 4484 7783
rect 4488 7779 4489 7783
rect 4493 7779 4494 7783
rect 4498 7779 4499 7783
rect 4503 7779 4504 7783
rect 4508 7779 4509 7783
rect 4479 7778 4513 7779
rect 4483 7774 4484 7778
rect 4488 7774 4489 7778
rect 4493 7774 4494 7778
rect 4498 7774 4499 7778
rect 4503 7774 4504 7778
rect 4508 7774 4509 7778
rect 4529 7789 4530 7793
rect 4534 7789 4535 7793
rect 4539 7789 4540 7793
rect 4544 7789 4545 7793
rect 4549 7789 4550 7793
rect 4554 7789 4555 7793
rect 4525 7788 4559 7789
rect 4529 7784 4530 7788
rect 4534 7784 4535 7788
rect 4539 7784 4540 7788
rect 4544 7784 4545 7788
rect 4549 7784 4550 7788
rect 4554 7784 4555 7788
rect 4525 7783 4559 7784
rect 4529 7779 4530 7783
rect 4534 7779 4535 7783
rect 4539 7779 4540 7783
rect 4544 7779 4545 7783
rect 4549 7779 4550 7783
rect 4554 7779 4555 7783
rect 4525 7778 4559 7779
rect 4529 7774 4530 7778
rect 4534 7774 4535 7778
rect 4539 7774 4540 7778
rect 4544 7774 4545 7778
rect 4549 7774 4550 7778
rect 4554 7774 4555 7778
rect 4826 7772 5086 7775
rect 4826 7518 4829 7772
rect 5083 7518 5086 7772
rect 4826 7515 5086 7518
rect 4527 7503 4595 7504
rect 4527 7499 4529 7503
rect 4533 7499 4534 7503
rect 4538 7499 4539 7503
rect 4543 7499 4544 7503
rect 4548 7499 4549 7503
rect 4553 7499 4554 7503
rect 4558 7499 4559 7503
rect 4563 7499 4564 7503
rect 4568 7499 4569 7503
rect 4573 7499 4574 7503
rect 4578 7499 4579 7503
rect 4583 7499 4584 7503
rect 4588 7499 4589 7503
rect 4593 7499 4595 7503
rect 3836 7484 3844 7499
rect 4527 7498 4595 7499
rect 4527 7494 4529 7498
rect 4533 7494 4534 7498
rect 4538 7494 4539 7498
rect 4543 7494 4544 7498
rect 4548 7494 4549 7498
rect 4553 7494 4554 7498
rect 4558 7494 4559 7498
rect 4563 7494 4564 7498
rect 4568 7494 4569 7498
rect 4573 7494 4574 7498
rect 4578 7494 4579 7498
rect 4583 7494 4584 7498
rect 4588 7494 4589 7498
rect 4593 7494 4595 7498
rect 4527 7493 4595 7494
rect 4527 7489 4529 7493
rect 4533 7489 4534 7493
rect 4538 7489 4539 7493
rect 4543 7489 4544 7493
rect 4548 7489 4549 7493
rect 4553 7489 4554 7493
rect 4558 7489 4559 7493
rect 4563 7489 4564 7493
rect 4568 7489 4569 7493
rect 4573 7489 4574 7493
rect 4578 7489 4579 7493
rect 4583 7489 4584 7493
rect 4588 7489 4589 7493
rect 4593 7489 4595 7493
rect 4826 7490 5086 7493
rect 86 7193 346 7196
rect 617 7158 618 7162
rect 622 7158 623 7162
rect 627 7158 628 7162
rect 632 7158 633 7162
rect 637 7158 638 7162
rect 642 7158 643 7162
rect 613 7157 647 7158
rect 663 7158 664 7162
rect 668 7158 669 7162
rect 673 7158 674 7162
rect 678 7158 679 7162
rect 683 7158 684 7162
rect 688 7158 689 7162
rect 659 7157 693 7158
rect 617 7123 618 7127
rect 622 7123 623 7127
rect 627 7123 628 7127
rect 632 7123 633 7127
rect 637 7123 638 7127
rect 642 7123 643 7127
rect 613 7122 647 7123
rect 617 7118 618 7122
rect 622 7118 623 7122
rect 627 7118 628 7122
rect 632 7118 633 7122
rect 637 7118 638 7122
rect 642 7118 643 7122
rect 613 7117 647 7118
rect 617 7113 618 7117
rect 622 7113 623 7117
rect 627 7113 628 7117
rect 632 7113 633 7117
rect 637 7113 638 7117
rect 642 7113 643 7117
rect 613 7112 647 7113
rect 86 7106 346 7109
rect 617 7108 618 7112
rect 622 7108 623 7112
rect 627 7108 628 7112
rect 632 7108 633 7112
rect 637 7108 638 7112
rect 642 7108 643 7112
rect 663 7123 664 7127
rect 668 7123 669 7127
rect 673 7123 674 7127
rect 678 7123 679 7127
rect 683 7123 684 7127
rect 688 7123 689 7127
rect 659 7122 693 7123
rect 663 7118 664 7122
rect 668 7118 669 7122
rect 673 7118 674 7122
rect 678 7118 679 7122
rect 683 7118 684 7122
rect 688 7118 689 7122
rect 659 7117 693 7118
rect 663 7113 664 7117
rect 668 7113 669 7117
rect 673 7113 674 7117
rect 678 7113 679 7117
rect 683 7113 684 7117
rect 688 7113 689 7117
rect 659 7112 693 7113
rect 663 7108 664 7112
rect 668 7108 669 7112
rect 673 7108 674 7112
rect 678 7108 679 7112
rect 683 7108 684 7112
rect 688 7108 689 7112
rect 86 6852 89 7106
rect 343 6852 346 7106
rect 86 6849 346 6852
rect 86 6796 346 6799
rect 86 6542 89 6796
rect 343 6542 346 6796
rect 86 6539 346 6542
rect 617 6536 618 6540
rect 622 6536 623 6540
rect 627 6536 628 6540
rect 632 6536 633 6540
rect 637 6536 638 6540
rect 642 6536 643 6540
rect 613 6535 647 6536
rect 617 6531 618 6535
rect 622 6531 623 6535
rect 627 6531 628 6535
rect 632 6531 633 6535
rect 637 6531 638 6535
rect 642 6531 643 6535
rect 613 6530 647 6531
rect 617 6526 618 6530
rect 622 6526 623 6530
rect 627 6526 628 6530
rect 632 6526 633 6530
rect 637 6526 638 6530
rect 642 6526 643 6530
rect 613 6525 647 6526
rect 617 6521 618 6525
rect 622 6521 623 6525
rect 627 6521 628 6525
rect 632 6521 633 6525
rect 637 6521 638 6525
rect 642 6521 643 6525
rect 663 6536 664 6540
rect 668 6536 669 6540
rect 673 6536 674 6540
rect 678 6536 679 6540
rect 683 6536 684 6540
rect 688 6536 689 6540
rect 659 6535 693 6536
rect 663 6531 664 6535
rect 668 6531 669 6535
rect 673 6531 674 6535
rect 678 6531 679 6535
rect 683 6531 684 6535
rect 688 6531 689 6535
rect 659 6530 693 6531
rect 663 6526 664 6530
rect 668 6526 669 6530
rect 673 6526 674 6530
rect 678 6526 679 6530
rect 683 6526 684 6530
rect 688 6526 689 6530
rect 659 6525 693 6526
rect 663 6521 664 6525
rect 668 6521 669 6525
rect 673 6521 674 6525
rect 678 6521 679 6525
rect 683 6521 684 6525
rect 688 6521 689 6525
rect 577 6505 645 6507
rect 577 6501 579 6505
rect 583 6501 584 6505
rect 588 6501 589 6505
rect 593 6501 594 6505
rect 598 6501 599 6505
rect 603 6501 604 6505
rect 608 6501 609 6505
rect 613 6501 614 6505
rect 618 6501 619 6505
rect 623 6501 624 6505
rect 628 6501 629 6505
rect 633 6501 634 6505
rect 638 6501 639 6505
rect 643 6501 645 6505
rect 577 6500 645 6501
rect 577 6496 579 6500
rect 583 6496 584 6500
rect 588 6496 589 6500
rect 593 6496 594 6500
rect 598 6496 599 6500
rect 603 6496 604 6500
rect 608 6496 609 6500
rect 613 6496 614 6500
rect 618 6496 619 6500
rect 623 6496 624 6500
rect 628 6496 629 6500
rect 633 6496 634 6500
rect 638 6496 639 6500
rect 643 6496 645 6500
rect 577 6495 645 6496
rect 577 6491 579 6495
rect 583 6491 584 6495
rect 588 6491 589 6495
rect 593 6491 594 6495
rect 598 6491 599 6495
rect 603 6491 604 6495
rect 608 6491 609 6495
rect 613 6491 614 6495
rect 618 6491 619 6495
rect 623 6491 624 6495
rect 628 6491 629 6495
rect 633 6491 634 6495
rect 638 6491 639 6495
rect 643 6491 645 6495
rect 577 6490 645 6491
rect 86 6487 346 6490
rect 86 6233 89 6487
rect 343 6233 346 6487
rect 577 6486 579 6490
rect 583 6486 584 6490
rect 588 6486 589 6490
rect 593 6486 594 6490
rect 598 6486 599 6490
rect 603 6486 604 6490
rect 608 6486 609 6490
rect 613 6486 614 6490
rect 618 6486 619 6490
rect 623 6486 624 6490
rect 628 6486 629 6490
rect 633 6486 634 6490
rect 638 6486 639 6490
rect 643 6486 645 6490
rect 427 6386 439 6390
rect 443 6386 464 6390
rect 468 6386 480 6390
rect 484 6386 507 6390
rect 511 6386 523 6390
rect 527 6386 546 6390
rect 550 6386 562 6390
rect 566 6386 578 6390
rect 582 6386 594 6390
rect 803 6364 812 6811
rect 927 6729 931 6811
rect 966 6739 969 6749
rect 949 6716 952 6717
rect 927 6567 931 6709
rect 949 6711 952 6712
rect 965 6713 968 6722
rect 986 6707 989 6720
rect 1002 6713 1005 6722
rect 1011 6711 1014 6716
rect 1017 6696 1020 6749
rect 1029 6735 1030 6739
rect 1068 6737 1071 6749
rect 1023 6713 1026 6722
rect 1023 6703 1027 6707
rect 964 6682 967 6692
rect 1031 6682 1034 6735
rect 1044 6707 1047 6720
rect 1060 6713 1063 6722
rect 1067 6682 1070 6692
rect 1074 6675 1077 6712
rect 949 6640 952 6670
rect 966 6653 969 6663
rect 949 6627 952 6636
rect 965 6627 968 6636
rect 986 6621 989 6634
rect 1002 6627 1005 6636
rect 1011 6625 1014 6630
rect 949 6575 952 6621
rect 1017 6610 1020 6663
rect 1029 6649 1030 6653
rect 1068 6651 1071 6663
rect 1023 6627 1026 6636
rect 1023 6617 1027 6621
rect 964 6596 967 6606
rect 1031 6596 1034 6649
rect 1044 6621 1047 6634
rect 1060 6627 1063 6636
rect 1067 6596 1070 6606
rect 1081 6603 1085 6685
rect 1385 6582 1391 6933
rect 949 6572 950 6575
rect 455 6360 515 6362
rect 455 6351 461 6360
rect 469 6351 505 6360
rect 513 6351 515 6360
rect 455 6349 515 6351
rect 427 6328 439 6332
rect 443 6328 464 6332
rect 468 6328 480 6332
rect 484 6328 507 6332
rect 511 6328 523 6332
rect 527 6328 546 6332
rect 550 6328 562 6332
rect 566 6328 578 6332
rect 582 6328 594 6332
rect 939 6327 943 6563
rect 956 6544 959 6557
rect 963 6547 966 6550
rect 984 6544 987 6557
rect 1000 6544 1003 6557
rect 957 6495 960 6510
rect 977 6502 981 6505
rect 985 6495 988 6510
rect 1000 6495 1003 6510
rect 1009 6502 1012 6543
rect 1028 6510 1031 6550
rect 1034 6502 1037 6543
rect 1050 6509 1053 6550
rect 1057 6544 1060 6557
rect 1074 6544 1077 6557
rect 1081 6547 1084 6550
rect 1107 6544 1111 6557
rect 1056 6495 1059 6510
rect 1075 6495 1078 6510
rect 1093 6502 1096 6506
rect 1115 6502 1118 6571
rect 1125 6554 1128 6564
rect 1133 6544 1137 6557
rect 1145 6458 1149 6530
rect 1153 6436 1156 6514
rect 1164 6472 1167 6550
rect 1217 6544 1220 6557
rect 1224 6547 1227 6550
rect 1245 6544 1248 6557
rect 1261 6544 1264 6557
rect 1218 6495 1221 6510
rect 1238 6502 1242 6505
rect 1246 6495 1249 6510
rect 1261 6495 1264 6510
rect 1270 6502 1273 6543
rect 1289 6510 1292 6550
rect 1295 6502 1298 6543
rect 1311 6509 1314 6550
rect 1318 6544 1321 6557
rect 1335 6544 1338 6557
rect 1359 6554 1363 6564
rect 1342 6547 1345 6550
rect 1368 6544 1371 6557
rect 1317 6495 1320 6510
rect 1336 6495 1339 6510
rect 1354 6502 1357 6506
rect 1218 6476 1221 6491
rect 1238 6481 1242 6484
rect 1246 6476 1249 6491
rect 1261 6476 1264 6491
rect 1157 6433 1161 6436
rect 974 6326 978 6394
rect 982 6304 985 6378
rect 993 6340 996 6414
rect 993 6317 996 6336
rect 1064 6326 1068 6394
rect 993 6314 1013 6317
rect 1028 6304 1031 6314
rect 986 6301 1031 6304
rect 661 6286 662 6290
rect 666 6286 667 6290
rect 671 6286 672 6290
rect 676 6286 678 6290
rect 657 6285 678 6286
rect 661 6281 662 6285
rect 666 6281 667 6285
rect 671 6281 672 6285
rect 676 6281 678 6285
rect 657 6280 678 6281
rect 661 6276 662 6280
rect 666 6276 667 6280
rect 671 6276 672 6280
rect 676 6276 678 6280
rect 657 6275 678 6276
rect 661 6271 662 6275
rect 666 6271 667 6275
rect 671 6271 672 6275
rect 676 6271 678 6275
rect 657 6270 678 6271
rect 661 6266 662 6270
rect 666 6266 667 6270
rect 671 6266 672 6270
rect 676 6266 678 6270
rect 657 6265 678 6266
rect 661 6261 662 6265
rect 666 6261 667 6265
rect 671 6261 672 6265
rect 676 6261 678 6265
rect 657 6260 678 6261
rect 661 6256 662 6260
rect 666 6256 667 6260
rect 671 6256 672 6260
rect 676 6256 678 6260
rect 657 6255 678 6256
rect 661 6251 662 6255
rect 666 6251 667 6255
rect 671 6251 672 6255
rect 676 6251 678 6255
rect 657 6250 678 6251
rect 661 6246 662 6250
rect 666 6246 667 6250
rect 671 6246 672 6250
rect 676 6246 678 6250
rect 657 6245 678 6246
rect 661 6241 662 6245
rect 666 6241 667 6245
rect 671 6241 672 6245
rect 676 6241 678 6245
rect 657 6240 678 6241
rect 661 6236 662 6240
rect 666 6236 667 6240
rect 671 6236 672 6240
rect 676 6236 678 6240
rect 657 6234 678 6236
rect 86 6230 346 6233
rect 617 6227 618 6231
rect 622 6227 623 6231
rect 627 6227 628 6231
rect 632 6227 633 6231
rect 637 6227 638 6231
rect 642 6227 643 6231
rect 613 6226 647 6227
rect 617 6222 618 6226
rect 622 6222 623 6226
rect 627 6222 628 6226
rect 632 6222 633 6226
rect 637 6222 638 6226
rect 642 6222 643 6226
rect 613 6221 647 6222
rect 617 6217 618 6221
rect 622 6217 623 6221
rect 627 6217 628 6221
rect 632 6217 633 6221
rect 637 6217 638 6221
rect 642 6217 643 6221
rect 613 6216 647 6217
rect 617 6212 618 6216
rect 622 6212 623 6216
rect 627 6212 628 6216
rect 632 6212 633 6216
rect 637 6212 638 6216
rect 642 6212 643 6216
rect 663 6227 664 6231
rect 668 6227 669 6231
rect 673 6227 674 6231
rect 678 6227 679 6231
rect 683 6227 684 6231
rect 688 6227 689 6231
rect 659 6226 693 6227
rect 663 6222 664 6226
rect 668 6222 669 6226
rect 673 6222 674 6226
rect 678 6222 679 6226
rect 683 6222 684 6226
rect 688 6222 689 6226
rect 659 6221 693 6222
rect 663 6217 664 6221
rect 668 6217 669 6221
rect 673 6217 674 6221
rect 678 6217 679 6221
rect 683 6217 684 6221
rect 688 6217 689 6221
rect 659 6216 693 6217
rect 663 6212 664 6216
rect 668 6212 669 6216
rect 673 6212 674 6216
rect 678 6212 679 6216
rect 683 6212 684 6216
rect 688 6212 689 6216
rect 617 6196 618 6200
rect 622 6196 623 6200
rect 627 6196 628 6200
rect 632 6196 633 6200
rect 637 6196 638 6200
rect 642 6196 643 6200
rect 613 6195 647 6196
rect 617 6191 618 6195
rect 622 6191 623 6195
rect 627 6191 628 6195
rect 632 6191 633 6195
rect 637 6191 638 6195
rect 642 6191 643 6195
rect 613 6190 647 6191
rect 617 6186 618 6190
rect 622 6186 623 6190
rect 627 6186 628 6190
rect 632 6186 633 6190
rect 637 6186 638 6190
rect 642 6186 643 6190
rect 613 6185 647 6186
rect 86 6179 346 6182
rect 617 6181 618 6185
rect 622 6181 623 6185
rect 627 6181 628 6185
rect 632 6181 633 6185
rect 637 6181 638 6185
rect 642 6181 643 6185
rect 663 6196 664 6200
rect 668 6196 669 6200
rect 673 6196 674 6200
rect 678 6196 679 6200
rect 683 6196 684 6200
rect 688 6196 689 6200
rect 659 6195 693 6196
rect 663 6191 664 6195
rect 668 6191 669 6195
rect 673 6191 674 6195
rect 678 6191 679 6195
rect 683 6191 684 6195
rect 688 6191 689 6195
rect 659 6190 693 6191
rect 663 6186 664 6190
rect 668 6186 669 6190
rect 673 6186 674 6190
rect 678 6186 679 6190
rect 683 6186 684 6190
rect 688 6186 689 6190
rect 659 6185 693 6186
rect 663 6181 664 6185
rect 668 6181 669 6185
rect 673 6181 674 6185
rect 678 6181 679 6185
rect 683 6181 684 6185
rect 688 6181 689 6185
rect 86 5925 89 6179
rect 343 5925 346 6179
rect 852 6030 920 6033
rect 1028 6033 1031 6301
rect 1072 6304 1075 6378
rect 1083 6340 1086 6414
rect 1083 6317 1086 6336
rect 1145 6326 1149 6394
rect 1153 6382 1156 6432
rect 1164 6418 1167 6468
rect 1217 6429 1220 6442
rect 1224 6436 1227 6439
rect 1245 6429 1248 6442
rect 1083 6314 1103 6317
rect 1118 6304 1121 6314
rect 1076 6301 1121 6304
rect 1153 6304 1156 6378
rect 1164 6340 1167 6414
rect 1217 6412 1220 6425
rect 1224 6415 1227 6418
rect 1245 6412 1248 6425
rect 1261 6429 1264 6442
rect 1270 6443 1273 6484
rect 1289 6436 1292 6476
rect 1295 6443 1298 6484
rect 1311 6436 1314 6477
rect 1317 6476 1320 6491
rect 1336 6476 1339 6491
rect 1344 6488 1348 6498
rect 1368 6495 1371 6510
rect 1354 6480 1357 6484
rect 1368 6476 1371 6491
rect 1318 6429 1321 6442
rect 1335 6429 1338 6442
rect 1342 6436 1345 6439
rect 1261 6412 1264 6425
rect 1218 6363 1221 6378
rect 1238 6370 1242 6373
rect 1246 6363 1249 6378
rect 1261 6363 1264 6378
rect 1270 6370 1273 6411
rect 1289 6378 1292 6418
rect 1295 6370 1298 6411
rect 1311 6377 1314 6418
rect 1318 6412 1321 6425
rect 1335 6412 1338 6425
rect 1368 6429 1371 6442
rect 1342 6415 1345 6418
rect 1368 6412 1371 6425
rect 1317 6363 1320 6378
rect 1336 6363 1339 6378
rect 1354 6370 1357 6374
rect 1368 6363 1371 6378
rect 1218 6344 1221 6359
rect 1238 6349 1242 6352
rect 1246 6344 1249 6359
rect 1261 6344 1264 6359
rect 1040 6194 1044 6259
rect 1048 6172 1051 6243
rect 1059 6208 1062 6279
rect 1059 6185 1062 6204
rect 1094 6186 1097 6187
rect 1059 6182 1079 6185
rect 1094 6172 1097 6182
rect 1052 6169 1097 6172
rect 1094 6165 1097 6169
rect 1056 6161 1097 6165
rect 924 6030 1031 6033
rect 852 6001 855 6030
rect 1056 6027 1059 6161
rect 1064 6062 1068 6128
rect 1072 6040 1075 6112
rect 1083 6076 1086 6148
rect 1083 6053 1086 6072
rect 1083 6050 1103 6053
rect 1115 6050 1118 6301
rect 1157 6301 1161 6304
rect 1145 6194 1149 6259
rect 1153 6247 1156 6300
rect 1164 6283 1167 6336
rect 1217 6297 1220 6310
rect 1224 6304 1227 6307
rect 1245 6297 1248 6310
rect 1153 6172 1156 6243
rect 1164 6208 1167 6279
rect 1217 6280 1220 6293
rect 1224 6283 1227 6286
rect 1245 6280 1248 6293
rect 1261 6297 1264 6310
rect 1270 6311 1273 6352
rect 1289 6304 1292 6344
rect 1295 6311 1298 6352
rect 1311 6304 1314 6345
rect 1317 6344 1320 6359
rect 1336 6344 1339 6359
rect 1354 6348 1357 6352
rect 1368 6344 1371 6359
rect 1318 6297 1321 6310
rect 1335 6297 1338 6310
rect 1342 6304 1345 6307
rect 1261 6280 1264 6293
rect 1218 6231 1221 6246
rect 1238 6238 1242 6241
rect 1246 6231 1249 6246
rect 1261 6231 1264 6246
rect 1270 6238 1273 6279
rect 1289 6246 1292 6286
rect 1295 6238 1298 6279
rect 1311 6245 1314 6286
rect 1318 6280 1321 6293
rect 1335 6280 1338 6293
rect 1368 6297 1371 6310
rect 1342 6283 1345 6286
rect 1368 6280 1371 6293
rect 1317 6231 1320 6246
rect 1336 6231 1339 6246
rect 1354 6238 1357 6242
rect 1368 6231 1371 6246
rect 1218 6212 1221 6227
rect 1238 6217 1242 6220
rect 1246 6212 1249 6227
rect 1261 6212 1264 6227
rect 1164 6185 1167 6204
rect 1164 6182 1168 6185
rect 1157 6169 1161 6172
rect 1145 6062 1149 6128
rect 1153 6116 1156 6168
rect 1164 6152 1167 6182
rect 1217 6165 1220 6178
rect 1224 6172 1227 6175
rect 1245 6165 1248 6178
rect 1118 6040 1121 6050
rect 1076 6037 1121 6040
rect 1118 6034 1121 6037
rect 1153 6040 1156 6112
rect 1164 6076 1167 6148
rect 1217 6148 1220 6161
rect 1224 6151 1227 6154
rect 1245 6148 1248 6161
rect 1261 6165 1264 6178
rect 1270 6179 1273 6220
rect 1289 6172 1292 6212
rect 1295 6179 1298 6220
rect 1311 6172 1314 6213
rect 1317 6212 1320 6227
rect 1336 6212 1339 6227
rect 1354 6216 1357 6220
rect 1368 6212 1371 6227
rect 1318 6165 1321 6178
rect 1335 6165 1338 6178
rect 1342 6172 1345 6175
rect 1261 6148 1264 6161
rect 1218 6099 1221 6114
rect 1238 6106 1242 6109
rect 1246 6099 1249 6114
rect 1261 6099 1264 6114
rect 1270 6106 1273 6147
rect 1289 6114 1292 6154
rect 1295 6106 1298 6147
rect 1311 6113 1314 6154
rect 1318 6148 1321 6161
rect 1335 6148 1338 6161
rect 1357 6158 1361 6168
rect 1368 6165 1371 6178
rect 1342 6151 1345 6154
rect 1368 6148 1371 6161
rect 1317 6099 1320 6114
rect 1336 6099 1339 6114
rect 1354 6106 1357 6110
rect 1368 6099 1371 6114
rect 1218 6080 1221 6095
rect 1238 6085 1242 6088
rect 1246 6080 1249 6095
rect 1261 6080 1264 6095
rect 1164 6053 1167 6072
rect 1164 6050 1184 6053
rect 1199 6040 1202 6050
rect 1157 6037 1202 6040
rect 984 6023 1059 6027
rect 1116 6029 1121 6034
rect 869 6006 872 6016
rect 852 5993 855 5997
rect 852 5983 855 5989
rect 851 5980 855 5983
rect 852 5978 855 5980
rect 868 5980 871 5989
rect 889 5974 892 5987
rect 905 5980 908 5989
rect 914 5978 917 5983
rect 920 5963 923 6016
rect 932 6002 933 6006
rect 971 6004 974 6016
rect 926 5980 929 5989
rect 926 5970 930 5974
rect 867 5949 870 5959
rect 934 5949 937 6002
rect 984 6001 987 6023
rect 1001 6006 1004 6016
rect 947 5974 950 5987
rect 963 5980 966 5989
rect 984 5983 987 5989
rect 980 5980 987 5983
rect 984 5978 987 5980
rect 1000 5980 1003 5989
rect 1021 5974 1024 5987
rect 1037 5980 1040 5989
rect 1046 5978 1049 5983
rect 1052 5963 1055 6016
rect 1064 6002 1065 6006
rect 1103 6004 1106 6016
rect 1058 5980 1061 5989
rect 1058 5970 1062 5974
rect 970 5949 973 5959
rect 999 5949 1002 5959
rect 1066 5949 1069 6002
rect 1116 5993 1119 6029
rect 1199 6026 1202 6037
rect 1217 6033 1220 6046
rect 1224 6040 1227 6043
rect 1245 6033 1248 6046
rect 1261 6033 1264 6046
rect 1270 6047 1273 6088
rect 1289 6040 1292 6080
rect 1295 6047 1298 6088
rect 1311 6040 1314 6081
rect 1317 6080 1320 6095
rect 1336 6080 1339 6095
rect 1354 6084 1357 6088
rect 1368 6080 1371 6095
rect 1318 6033 1321 6046
rect 1335 6033 1338 6046
rect 1342 6040 1345 6043
rect 1368 6033 1371 6046
rect 1199 6023 1251 6026
rect 1133 6006 1136 6016
rect 1079 5974 1082 5987
rect 1095 5980 1098 5989
rect 1116 5983 1119 5989
rect 1112 5980 1119 5983
rect 1116 5978 1119 5980
rect 1132 5980 1135 5989
rect 1153 5974 1156 5987
rect 1169 5980 1172 5989
rect 1178 5978 1181 5983
rect 1184 5963 1187 6016
rect 1196 6002 1197 6006
rect 1235 6004 1238 6016
rect 1190 5980 1193 5989
rect 1190 5970 1194 5974
rect 1102 5949 1105 5959
rect 1131 5949 1134 5959
rect 1198 5949 1201 6002
rect 1248 5993 1251 6023
rect 1265 6006 1268 6016
rect 1211 5974 1214 5987
rect 1227 5980 1230 5989
rect 1248 5983 1251 5989
rect 1244 5980 1251 5983
rect 1248 5978 1251 5980
rect 1264 5980 1267 5989
rect 1285 5974 1288 5987
rect 1301 5980 1304 5989
rect 1310 5978 1313 5983
rect 1316 5963 1319 6016
rect 1328 6002 1329 6006
rect 1367 6004 1370 6016
rect 1322 5980 1325 5989
rect 1322 5970 1326 5974
rect 1234 5949 1237 5959
rect 1263 5949 1266 5959
rect 1330 5949 1333 6002
rect 1343 5974 1346 5987
rect 1359 5980 1362 5989
rect 1366 5949 1369 5959
rect 86 5922 346 5925
rect 617 5887 618 5891
rect 622 5887 623 5891
rect 627 5887 628 5891
rect 632 5887 633 5891
rect 637 5887 638 5891
rect 642 5887 643 5891
rect 613 5886 647 5887
rect 617 5882 618 5886
rect 622 5882 623 5886
rect 627 5882 628 5886
rect 632 5882 633 5886
rect 637 5882 638 5886
rect 642 5882 643 5886
rect 613 5881 647 5882
rect 617 5877 618 5881
rect 622 5877 623 5881
rect 627 5877 628 5881
rect 632 5877 633 5881
rect 637 5877 638 5881
rect 642 5877 643 5881
rect 613 5876 647 5877
rect 86 5870 346 5873
rect 617 5872 618 5876
rect 622 5872 623 5876
rect 627 5872 628 5876
rect 632 5872 633 5876
rect 637 5872 638 5876
rect 642 5872 643 5876
rect 663 5887 664 5891
rect 668 5887 669 5891
rect 673 5887 674 5891
rect 678 5887 679 5891
rect 683 5887 684 5891
rect 688 5887 689 5891
rect 659 5886 693 5887
rect 663 5882 664 5886
rect 668 5882 669 5886
rect 673 5882 674 5886
rect 678 5882 679 5886
rect 683 5882 684 5886
rect 688 5882 689 5886
rect 659 5881 693 5882
rect 663 5877 664 5881
rect 668 5877 669 5881
rect 673 5877 674 5881
rect 678 5877 679 5881
rect 683 5877 684 5881
rect 688 5877 689 5881
rect 659 5876 693 5877
rect 663 5872 664 5876
rect 668 5872 669 5876
rect 673 5872 674 5876
rect 678 5872 679 5876
rect 683 5872 684 5876
rect 688 5872 689 5876
rect 86 5616 89 5870
rect 343 5616 346 5870
rect 927 5747 931 5829
rect 966 5757 969 5767
rect 949 5734 952 5735
rect 86 5613 346 5616
rect 927 5585 931 5727
rect 949 5729 952 5730
rect 965 5731 968 5740
rect 986 5725 989 5738
rect 1002 5731 1005 5740
rect 1011 5729 1014 5734
rect 1017 5714 1020 5767
rect 1029 5753 1030 5757
rect 1068 5755 1071 5767
rect 1023 5731 1026 5740
rect 1023 5721 1027 5725
rect 964 5700 967 5710
rect 1031 5700 1034 5753
rect 1044 5725 1047 5738
rect 1060 5731 1063 5740
rect 1067 5700 1070 5710
rect 1074 5693 1077 5730
rect 949 5658 952 5688
rect 966 5671 969 5681
rect 949 5645 952 5654
rect 965 5645 968 5654
rect 986 5639 989 5652
rect 1002 5645 1005 5654
rect 1011 5643 1014 5648
rect 949 5593 952 5639
rect 1017 5628 1020 5681
rect 1029 5667 1030 5671
rect 1068 5669 1071 5681
rect 1023 5645 1026 5654
rect 1023 5635 1027 5639
rect 964 5614 967 5624
rect 1031 5614 1034 5667
rect 1044 5639 1047 5652
rect 1060 5645 1063 5654
rect 1067 5614 1070 5624
rect 1081 5621 1085 5703
rect 1385 5600 1391 6578
rect 949 5590 950 5593
rect 617 5578 618 5582
rect 622 5578 623 5582
rect 627 5578 628 5582
rect 632 5578 633 5582
rect 637 5578 638 5582
rect 642 5578 643 5582
rect 613 5577 647 5578
rect 617 5573 618 5577
rect 622 5573 623 5577
rect 627 5573 628 5577
rect 632 5573 633 5577
rect 637 5573 638 5577
rect 642 5573 643 5577
rect 613 5572 647 5573
rect 617 5568 618 5572
rect 622 5568 623 5572
rect 627 5568 628 5572
rect 632 5568 633 5572
rect 637 5568 638 5572
rect 642 5568 643 5572
rect 613 5567 647 5568
rect 86 5561 346 5564
rect 617 5563 618 5567
rect 622 5563 623 5567
rect 627 5563 628 5567
rect 632 5563 633 5567
rect 637 5563 638 5567
rect 642 5563 643 5567
rect 663 5578 664 5582
rect 668 5578 669 5582
rect 673 5578 674 5582
rect 678 5578 679 5582
rect 683 5578 684 5582
rect 688 5578 689 5582
rect 659 5577 693 5578
rect 663 5573 664 5577
rect 668 5573 669 5577
rect 673 5573 674 5577
rect 678 5573 679 5577
rect 683 5573 684 5577
rect 688 5573 689 5577
rect 659 5572 693 5573
rect 663 5568 664 5572
rect 668 5568 669 5572
rect 673 5568 674 5572
rect 678 5568 679 5572
rect 683 5568 684 5572
rect 688 5568 689 5572
rect 659 5567 693 5568
rect 663 5563 664 5567
rect 668 5563 669 5567
rect 673 5563 674 5567
rect 678 5563 679 5567
rect 683 5563 684 5567
rect 688 5563 689 5567
rect 86 5307 89 5561
rect 343 5307 346 5561
rect 939 5345 943 5581
rect 956 5562 959 5575
rect 963 5565 966 5568
rect 984 5562 987 5575
rect 1000 5562 1003 5575
rect 957 5513 960 5528
rect 977 5520 981 5523
rect 985 5513 988 5528
rect 1000 5513 1003 5528
rect 1009 5520 1012 5561
rect 1028 5528 1031 5568
rect 1034 5520 1037 5561
rect 1050 5527 1053 5568
rect 1057 5562 1060 5575
rect 1074 5562 1077 5575
rect 1081 5565 1084 5568
rect 1107 5562 1111 5575
rect 1056 5513 1059 5528
rect 1075 5513 1078 5528
rect 1093 5520 1096 5524
rect 1115 5520 1118 5589
rect 1125 5572 1128 5582
rect 1133 5562 1137 5575
rect 1145 5476 1149 5548
rect 1153 5454 1156 5532
rect 1164 5490 1167 5568
rect 1217 5562 1220 5575
rect 1224 5565 1227 5568
rect 1245 5562 1248 5575
rect 1261 5562 1264 5575
rect 1218 5513 1221 5528
rect 1238 5520 1242 5523
rect 1246 5513 1249 5528
rect 1261 5513 1264 5528
rect 1270 5520 1273 5561
rect 1289 5528 1292 5568
rect 1295 5520 1298 5561
rect 1311 5527 1314 5568
rect 1318 5562 1321 5575
rect 1335 5562 1338 5575
rect 1359 5572 1363 5582
rect 1342 5565 1345 5568
rect 1368 5562 1371 5575
rect 1317 5513 1320 5528
rect 1336 5513 1339 5528
rect 1354 5520 1357 5524
rect 1218 5494 1221 5509
rect 1238 5499 1242 5502
rect 1246 5494 1249 5509
rect 1261 5494 1264 5509
rect 1157 5451 1161 5454
rect 974 5344 978 5412
rect 982 5322 985 5396
rect 993 5358 996 5432
rect 993 5335 996 5354
rect 1064 5344 1068 5412
rect 993 5332 1013 5335
rect 1028 5322 1031 5332
rect 986 5319 1031 5322
rect 86 5304 346 5307
rect 617 5269 618 5273
rect 622 5269 623 5273
rect 627 5269 628 5273
rect 632 5269 633 5273
rect 637 5269 638 5273
rect 642 5269 643 5273
rect 613 5268 647 5269
rect 617 5264 618 5268
rect 622 5264 623 5268
rect 627 5264 628 5268
rect 632 5264 633 5268
rect 637 5264 638 5268
rect 642 5264 643 5268
rect 613 5263 647 5264
rect 617 5259 618 5263
rect 622 5259 623 5263
rect 627 5259 628 5263
rect 632 5259 633 5263
rect 637 5259 638 5263
rect 642 5259 643 5263
rect 613 5258 647 5259
rect 86 5252 346 5255
rect 617 5254 618 5258
rect 622 5254 623 5258
rect 627 5254 628 5258
rect 632 5254 633 5258
rect 637 5254 638 5258
rect 642 5254 643 5258
rect 663 5269 664 5273
rect 668 5269 669 5273
rect 673 5269 674 5273
rect 678 5269 679 5273
rect 683 5269 684 5273
rect 688 5269 689 5273
rect 659 5268 693 5269
rect 663 5264 664 5268
rect 668 5264 669 5268
rect 673 5264 674 5268
rect 678 5264 679 5268
rect 683 5264 684 5268
rect 688 5264 689 5268
rect 659 5263 693 5264
rect 663 5259 664 5263
rect 668 5259 669 5263
rect 673 5259 674 5263
rect 678 5259 679 5263
rect 683 5259 684 5263
rect 688 5259 689 5263
rect 659 5258 693 5259
rect 663 5254 664 5258
rect 668 5254 669 5258
rect 673 5254 674 5258
rect 678 5254 679 5258
rect 683 5254 684 5258
rect 688 5254 689 5258
rect 86 4998 89 5252
rect 343 4998 346 5252
rect 852 5048 920 5051
rect 1028 5051 1031 5319
rect 1072 5322 1075 5396
rect 1083 5358 1086 5432
rect 1083 5335 1086 5354
rect 1145 5344 1149 5412
rect 1153 5400 1156 5450
rect 1164 5436 1167 5486
rect 1217 5447 1220 5460
rect 1224 5454 1227 5457
rect 1245 5447 1248 5460
rect 1083 5332 1103 5335
rect 1118 5322 1121 5332
rect 1076 5319 1121 5322
rect 1153 5322 1156 5396
rect 1164 5358 1167 5432
rect 1217 5430 1220 5443
rect 1224 5433 1227 5436
rect 1245 5430 1248 5443
rect 1261 5447 1264 5460
rect 1270 5461 1273 5502
rect 1289 5454 1292 5494
rect 1295 5461 1298 5502
rect 1311 5454 1314 5495
rect 1317 5494 1320 5509
rect 1336 5494 1339 5509
rect 1344 5506 1348 5516
rect 1368 5513 1371 5528
rect 1354 5498 1357 5502
rect 1368 5494 1371 5509
rect 1318 5447 1321 5460
rect 1335 5447 1338 5460
rect 1342 5454 1345 5457
rect 1261 5430 1264 5443
rect 1218 5381 1221 5396
rect 1238 5388 1242 5391
rect 1246 5381 1249 5396
rect 1261 5381 1264 5396
rect 1270 5388 1273 5429
rect 1289 5396 1292 5436
rect 1295 5388 1298 5429
rect 1311 5395 1314 5436
rect 1318 5430 1321 5443
rect 1335 5430 1338 5443
rect 1368 5447 1371 5460
rect 1342 5433 1345 5436
rect 1368 5430 1371 5443
rect 1317 5381 1320 5396
rect 1336 5381 1339 5396
rect 1354 5388 1357 5392
rect 1368 5381 1371 5396
rect 1218 5362 1221 5377
rect 1238 5367 1242 5370
rect 1246 5362 1249 5377
rect 1261 5362 1264 5377
rect 1040 5212 1044 5277
rect 1048 5190 1051 5261
rect 1059 5226 1062 5297
rect 1059 5203 1062 5222
rect 1094 5204 1097 5205
rect 1059 5200 1079 5203
rect 1094 5190 1097 5200
rect 1052 5187 1097 5190
rect 1094 5183 1097 5187
rect 1056 5179 1097 5183
rect 924 5048 1031 5051
rect 852 5019 855 5048
rect 1056 5045 1059 5179
rect 1064 5080 1068 5146
rect 1072 5058 1075 5130
rect 1083 5094 1086 5166
rect 1083 5071 1086 5090
rect 1083 5068 1103 5071
rect 1115 5068 1118 5319
rect 1157 5319 1161 5322
rect 1145 5212 1149 5277
rect 1153 5265 1156 5318
rect 1164 5301 1167 5354
rect 1217 5315 1220 5328
rect 1224 5322 1227 5325
rect 1245 5315 1248 5328
rect 1153 5190 1156 5261
rect 1164 5226 1167 5297
rect 1217 5298 1220 5311
rect 1224 5301 1227 5304
rect 1245 5298 1248 5311
rect 1261 5315 1264 5328
rect 1270 5329 1273 5370
rect 1289 5322 1292 5362
rect 1295 5329 1298 5370
rect 1311 5322 1314 5363
rect 1317 5362 1320 5377
rect 1336 5362 1339 5377
rect 1354 5366 1357 5370
rect 1368 5362 1371 5377
rect 1318 5315 1321 5328
rect 1335 5315 1338 5328
rect 1342 5322 1345 5325
rect 1261 5298 1264 5311
rect 1218 5249 1221 5264
rect 1238 5256 1242 5259
rect 1246 5249 1249 5264
rect 1261 5249 1264 5264
rect 1270 5256 1273 5297
rect 1289 5264 1292 5304
rect 1295 5256 1298 5297
rect 1311 5263 1314 5304
rect 1318 5298 1321 5311
rect 1335 5298 1338 5311
rect 1368 5315 1371 5328
rect 1342 5301 1345 5304
rect 1368 5298 1371 5311
rect 1385 5297 1391 5596
rect 1317 5249 1320 5264
rect 1336 5249 1339 5264
rect 1354 5256 1357 5260
rect 1368 5249 1371 5264
rect 1218 5230 1221 5245
rect 1238 5235 1242 5238
rect 1246 5230 1249 5245
rect 1261 5230 1264 5245
rect 1164 5203 1167 5222
rect 1164 5200 1168 5203
rect 1157 5187 1161 5190
rect 1145 5080 1149 5146
rect 1153 5134 1156 5186
rect 1164 5170 1167 5200
rect 1217 5183 1220 5196
rect 1224 5190 1227 5193
rect 1245 5183 1248 5196
rect 1118 5058 1121 5068
rect 1076 5055 1121 5058
rect 1118 5052 1121 5055
rect 1153 5058 1156 5130
rect 1164 5094 1167 5166
rect 1217 5166 1220 5179
rect 1224 5169 1227 5172
rect 1245 5166 1248 5179
rect 1261 5183 1264 5196
rect 1270 5197 1273 5238
rect 1289 5190 1292 5230
rect 1295 5197 1298 5238
rect 1311 5190 1314 5231
rect 1317 5230 1320 5245
rect 1336 5230 1339 5245
rect 1354 5234 1357 5238
rect 1368 5230 1371 5245
rect 1318 5183 1321 5196
rect 1335 5183 1338 5196
rect 1342 5190 1345 5193
rect 1261 5166 1264 5179
rect 1218 5117 1221 5132
rect 1238 5124 1242 5127
rect 1246 5117 1249 5132
rect 1261 5117 1264 5132
rect 1270 5124 1273 5165
rect 1289 5132 1292 5172
rect 1295 5124 1298 5165
rect 1311 5131 1314 5172
rect 1318 5166 1321 5179
rect 1335 5166 1338 5179
rect 1357 5176 1361 5186
rect 1368 5183 1371 5196
rect 1342 5169 1345 5172
rect 1368 5166 1371 5179
rect 1317 5117 1320 5132
rect 1336 5117 1339 5132
rect 1354 5124 1357 5128
rect 1368 5117 1371 5132
rect 1218 5098 1221 5113
rect 1238 5103 1242 5106
rect 1246 5098 1249 5113
rect 1261 5098 1264 5113
rect 1164 5071 1167 5090
rect 1164 5068 1184 5071
rect 1199 5058 1202 5068
rect 1157 5055 1202 5058
rect 984 5041 1059 5045
rect 1116 5047 1121 5052
rect 869 5024 872 5034
rect 852 5011 855 5015
rect 852 5001 855 5007
rect 851 4998 855 5001
rect 86 4995 346 4998
rect 852 4996 855 4998
rect 868 4998 871 5007
rect 889 4992 892 5005
rect 905 4998 908 5007
rect 914 4996 917 5001
rect 920 4981 923 5034
rect 932 5020 933 5024
rect 971 5022 974 5034
rect 926 4998 929 5007
rect 926 4988 930 4992
rect 867 4967 870 4977
rect 934 4967 937 5020
rect 984 5019 987 5041
rect 1001 5024 1004 5034
rect 947 4992 950 5005
rect 963 4998 966 5007
rect 984 5001 987 5007
rect 980 4998 987 5001
rect 984 4996 987 4998
rect 1000 4998 1003 5007
rect 1021 4992 1024 5005
rect 1037 4998 1040 5007
rect 1046 4996 1049 5001
rect 1052 4981 1055 5034
rect 1064 5020 1065 5024
rect 1103 5022 1106 5034
rect 1058 4998 1061 5007
rect 1058 4988 1062 4992
rect 970 4967 973 4977
rect 999 4967 1002 4977
rect 1066 4967 1069 5020
rect 1116 5011 1119 5047
rect 1199 5044 1202 5055
rect 1217 5051 1220 5064
rect 1224 5058 1227 5061
rect 1245 5051 1248 5064
rect 1261 5051 1264 5064
rect 1270 5065 1273 5106
rect 1289 5058 1292 5098
rect 1295 5065 1298 5106
rect 1311 5058 1314 5099
rect 1317 5098 1320 5113
rect 1336 5098 1339 5113
rect 1354 5102 1357 5106
rect 1368 5098 1371 5113
rect 1318 5051 1321 5064
rect 1335 5051 1338 5064
rect 1342 5058 1345 5061
rect 1368 5051 1371 5064
rect 1199 5041 1251 5044
rect 1133 5024 1136 5034
rect 1079 4992 1082 5005
rect 1095 4998 1098 5007
rect 1116 5001 1119 5007
rect 1112 4998 1119 5001
rect 1116 4996 1119 4998
rect 1132 4998 1135 5007
rect 1153 4992 1156 5005
rect 1169 4998 1172 5007
rect 1178 4996 1181 5001
rect 1184 4981 1187 5034
rect 1196 5020 1197 5024
rect 1235 5022 1238 5034
rect 1190 4998 1193 5007
rect 1190 4988 1194 4992
rect 1102 4967 1105 4977
rect 1131 4967 1134 4977
rect 1198 4967 1201 5020
rect 1248 5011 1251 5041
rect 1265 5024 1268 5034
rect 1211 4992 1214 5005
rect 1227 4998 1230 5007
rect 1248 5001 1251 5007
rect 1244 4998 1251 5001
rect 1248 4996 1251 4998
rect 1264 4998 1267 5007
rect 1285 4992 1288 5005
rect 1301 4998 1304 5007
rect 1310 4996 1313 5001
rect 1316 4981 1319 5034
rect 1328 5020 1329 5024
rect 1367 5022 1370 5034
rect 1322 4998 1325 5007
rect 1322 4988 1326 4992
rect 1234 4967 1237 4977
rect 1263 4967 1266 4977
rect 1330 4967 1333 5020
rect 1343 4992 1346 5005
rect 1359 4998 1362 5007
rect 1366 4967 1369 4977
rect 99 4528 593 4959
rect 617 4868 618 4872
rect 622 4868 623 4872
rect 627 4868 628 4872
rect 632 4868 633 4872
rect 637 4868 638 4872
rect 642 4868 643 4872
rect 613 4867 647 4868
rect 617 4863 618 4867
rect 622 4863 623 4867
rect 627 4863 628 4867
rect 632 4863 633 4867
rect 637 4863 638 4867
rect 642 4863 643 4867
rect 613 4862 647 4863
rect 617 4858 618 4862
rect 622 4858 623 4862
rect 627 4858 628 4862
rect 632 4858 633 4862
rect 637 4858 638 4862
rect 642 4858 643 4862
rect 613 4857 647 4858
rect 617 4853 618 4857
rect 622 4853 623 4857
rect 627 4853 628 4857
rect 632 4853 633 4857
rect 637 4853 638 4857
rect 642 4853 643 4857
rect 663 4868 664 4872
rect 668 4868 669 4872
rect 673 4868 674 4872
rect 678 4868 679 4872
rect 683 4868 684 4872
rect 688 4868 689 4872
rect 659 4867 693 4868
rect 663 4863 664 4867
rect 668 4863 669 4867
rect 673 4863 674 4867
rect 678 4863 679 4867
rect 683 4863 684 4867
rect 688 4863 689 4867
rect 659 4862 693 4863
rect 663 4858 664 4862
rect 668 4858 669 4862
rect 673 4858 674 4862
rect 678 4858 679 4862
rect 683 4858 684 4862
rect 688 4858 689 4862
rect 1385 4862 1391 5293
rect 1397 6852 1403 6933
rect 1397 6712 1403 6848
rect 1397 6682 1403 6708
rect 1397 6626 1403 6678
rect 1397 6596 1403 6622
rect 1397 6484 1403 6592
rect 1397 6084 1403 6480
rect 1397 5982 1403 6080
rect 1397 5949 1403 5978
rect 1397 5870 1403 5945
rect 1397 5730 1403 5866
rect 1397 5700 1403 5726
rect 1397 5644 1403 5696
rect 1397 5614 1403 5640
rect 1397 5502 1403 5610
rect 1397 5402 1403 5498
rect 1397 5102 1403 5398
rect 1397 5000 1403 5098
rect 1397 4967 1403 4996
rect 659 4857 693 4858
rect 663 4853 664 4857
rect 668 4853 669 4857
rect 673 4853 674 4857
rect 678 4853 679 4857
rect 683 4853 684 4857
rect 688 4853 689 4857
rect 617 4839 618 4843
rect 622 4839 623 4843
rect 627 4839 628 4843
rect 632 4839 633 4843
rect 637 4839 638 4843
rect 642 4839 643 4843
rect 613 4838 647 4839
rect 617 4834 618 4838
rect 622 4834 623 4838
rect 627 4834 628 4838
rect 632 4834 633 4838
rect 637 4834 638 4838
rect 642 4834 643 4838
rect 613 4833 647 4834
rect 617 4829 618 4833
rect 622 4829 623 4833
rect 627 4829 628 4833
rect 632 4829 633 4833
rect 637 4829 638 4833
rect 642 4829 643 4833
rect 613 4828 647 4829
rect 617 4824 618 4828
rect 622 4824 623 4828
rect 627 4824 628 4828
rect 632 4824 633 4828
rect 637 4824 638 4828
rect 642 4824 643 4828
rect 663 4839 664 4843
rect 668 4839 669 4843
rect 673 4839 674 4843
rect 678 4839 679 4843
rect 683 4839 684 4843
rect 688 4839 689 4843
rect 659 4838 693 4839
rect 663 4834 664 4838
rect 668 4834 669 4838
rect 673 4834 674 4838
rect 678 4834 679 4838
rect 683 4834 684 4838
rect 688 4834 689 4838
rect 659 4833 693 4834
rect 663 4829 664 4833
rect 668 4829 669 4833
rect 673 4829 674 4833
rect 678 4829 679 4833
rect 683 4829 684 4833
rect 688 4829 689 4833
rect 659 4828 693 4829
rect 663 4824 664 4828
rect 668 4824 669 4828
rect 673 4824 674 4828
rect 678 4824 679 4828
rect 683 4824 684 4828
rect 688 4824 689 4828
rect 1397 4817 1403 4963
rect 1409 6923 1415 6933
rect 1409 6783 1415 6919
rect 1409 6753 1415 6779
rect 1409 6697 1415 6749
rect 1409 6667 1415 6693
rect 1409 6554 1415 6663
rect 1409 6155 1415 6550
rect 1409 6053 1415 6151
rect 1409 6020 1415 6049
rect 1409 5941 1415 6016
rect 1409 5801 1415 5937
rect 1409 5771 1415 5797
rect 1409 5715 1415 5767
rect 1409 5685 1415 5711
rect 1409 5572 1415 5681
rect 1409 5432 1415 5568
rect 1409 5173 1415 5428
rect 1409 5071 1415 5169
rect 1409 5038 1415 5067
rect 1409 4902 1415 5034
rect 1409 4825 1415 4898
rect 1421 6568 1427 6933
rect 1421 6436 1427 6564
rect 1421 6422 1427 6432
rect 1421 6304 1427 6418
rect 1421 6290 1427 6300
rect 1421 6172 1427 6286
rect 1421 6040 1427 6168
rect 1421 5586 1427 6036
rect 1421 5454 1427 5582
rect 1421 5440 1427 5450
rect 1421 5322 1427 5436
rect 1421 5308 1427 5318
rect 1421 5269 1427 5304
rect 1421 5190 1427 5265
rect 1421 5058 1427 5186
rect 1421 4910 1427 5054
rect 1421 4832 1427 4906
rect 1433 6576 1439 6933
rect 1433 6502 1439 6572
rect 1433 6370 1439 6498
rect 1433 6356 1439 6366
rect 1433 6238 1439 6352
rect 1433 6224 1439 6234
rect 1433 6106 1439 6220
rect 1433 6092 1439 6102
rect 1433 5594 1439 6088
rect 1433 5520 1439 5590
rect 1433 5388 1439 5516
rect 1433 5374 1439 5384
rect 1433 5306 1439 5370
rect 1433 5256 1439 5302
rect 1433 5242 1439 5252
rect 1433 5124 1439 5238
rect 1433 5110 1439 5120
rect 1433 4918 1439 5106
rect 1433 4839 1439 4914
rect 1445 6916 1451 6933
rect 1445 6776 1451 6912
rect 1445 6746 1451 6772
rect 1445 6690 1451 6742
rect 1445 6660 1451 6686
rect 1445 6548 1451 6656
rect 1445 6495 1451 6544
rect 1445 6363 1451 6491
rect 1445 6231 1451 6359
rect 1445 6148 1451 6227
rect 1445 6099 1451 6144
rect 1445 6046 1451 6095
rect 1445 6013 1451 6042
rect 1445 5934 1451 6009
rect 1445 5794 1451 5930
rect 1445 5764 1451 5790
rect 1445 5708 1451 5760
rect 1445 5678 1451 5704
rect 1445 5566 1451 5674
rect 1445 5513 1451 5562
rect 1445 5381 1451 5509
rect 1445 5288 1451 5377
rect 1445 5249 1451 5284
rect 1445 5166 1451 5245
rect 1445 5117 1451 5162
rect 1445 5064 1451 5113
rect 1445 5031 1451 5060
rect 1445 4926 1451 5027
rect 1445 4847 1451 4922
rect 1457 6859 1463 6933
rect 1485 6909 1488 6919
rect 1468 6889 1471 6892
rect 1457 6719 1463 6855
rect 1468 6881 1471 6885
rect 1484 6883 1487 6892
rect 1505 6877 1508 6890
rect 1521 6883 1524 6892
rect 1530 6881 1533 6886
rect 1468 6830 1471 6877
rect 1536 6866 1539 6919
rect 1548 6905 1549 6909
rect 1587 6907 1590 6919
rect 1542 6883 1545 6892
rect 1542 6873 1546 6877
rect 1483 6852 1486 6862
rect 1550 6852 1553 6905
rect 1563 6877 1566 6890
rect 1579 6883 1582 6892
rect 1600 6883 1603 6892
rect 1586 6852 1589 6862
rect 1600 6845 1603 6877
rect 1608 6838 1612 6933
rect 1617 6909 1620 6919
rect 1616 6883 1619 6892
rect 1637 6877 1640 6890
rect 1653 6883 1656 6892
rect 1662 6881 1665 6886
rect 1668 6866 1671 6919
rect 1680 6905 1681 6909
rect 1719 6907 1722 6919
rect 1674 6883 1677 6892
rect 1674 6873 1678 6877
rect 1615 6852 1618 6862
rect 1682 6852 1685 6905
rect 1695 6877 1698 6890
rect 1711 6883 1714 6892
rect 1718 6852 1721 6862
rect 1592 6834 1596 6838
rect 1608 6833 1612 6834
rect 1468 6790 1471 6818
rect 1592 6815 1596 6830
rect 1592 6808 1596 6811
rect 1592 6800 1596 6804
rect 1608 6804 1612 6818
rect 1624 6815 1628 6830
rect 1624 6808 1628 6811
rect 1468 6756 1471 6786
rect 1485 6769 1488 6779
rect 1468 6741 1471 6752
rect 1484 6743 1487 6752
rect 1505 6737 1508 6750
rect 1521 6743 1524 6752
rect 1530 6741 1533 6746
rect 1536 6726 1539 6779
rect 1548 6765 1549 6769
rect 1587 6767 1590 6779
rect 1542 6743 1545 6752
rect 1542 6733 1546 6737
rect 1457 6633 1463 6715
rect 1483 6712 1486 6722
rect 1550 6712 1553 6765
rect 1600 6756 1603 6793
rect 1563 6737 1566 6750
rect 1579 6743 1582 6752
rect 1600 6743 1603 6752
rect 1586 6712 1589 6722
rect 1457 6603 1463 6629
rect 1468 6670 1471 6700
rect 1485 6683 1488 6693
rect 1468 6655 1471 6666
rect 1484 6657 1487 6666
rect 1505 6651 1508 6664
rect 1521 6657 1524 6666
rect 1530 6655 1533 6660
rect 1468 6604 1471 6651
rect 1536 6640 1539 6693
rect 1548 6679 1549 6683
rect 1587 6681 1590 6693
rect 1542 6657 1545 6666
rect 1542 6647 1546 6651
rect 1483 6626 1486 6636
rect 1550 6626 1553 6679
rect 1563 6651 1566 6664
rect 1579 6657 1582 6666
rect 1600 6657 1603 6666
rect 1586 6626 1589 6636
rect 1600 6619 1603 6651
rect 1457 6561 1463 6599
rect 1457 6491 1463 6557
rect 1468 6562 1471 6592
rect 1468 6528 1471 6558
rect 1485 6541 1488 6551
rect 1468 6513 1471 6524
rect 1484 6515 1487 6524
rect 1505 6509 1508 6522
rect 1521 6515 1524 6524
rect 1530 6513 1533 6518
rect 1536 6498 1539 6551
rect 1548 6537 1549 6541
rect 1587 6539 1590 6551
rect 1542 6515 1545 6524
rect 1542 6505 1546 6509
rect 1457 6429 1463 6487
rect 1483 6484 1486 6494
rect 1550 6484 1553 6537
rect 1600 6528 1603 6565
rect 1563 6509 1566 6522
rect 1579 6515 1582 6524
rect 1600 6515 1603 6524
rect 1586 6484 1589 6494
rect 1457 6297 1463 6425
rect 1457 6165 1463 6293
rect 1457 6091 1463 6161
rect 1457 6033 1463 6087
rect 1584 6067 1588 6072
rect 1608 6067 1612 6800
rect 1617 6769 1620 6779
rect 1616 6743 1619 6752
rect 1637 6737 1640 6750
rect 1653 6743 1656 6752
rect 1662 6741 1665 6746
rect 1668 6726 1671 6779
rect 1680 6765 1681 6769
rect 1719 6767 1722 6779
rect 1674 6743 1677 6752
rect 1674 6733 1678 6737
rect 1615 6712 1618 6722
rect 1682 6712 1685 6765
rect 1695 6737 1698 6750
rect 1711 6743 1714 6752
rect 1718 6712 1721 6722
rect 1617 6683 1620 6693
rect 1616 6657 1619 6666
rect 1637 6651 1640 6664
rect 1653 6657 1656 6666
rect 1662 6655 1665 6660
rect 1668 6640 1671 6693
rect 1680 6679 1681 6683
rect 1719 6681 1722 6693
rect 1674 6657 1677 6666
rect 1674 6647 1678 6651
rect 1615 6626 1618 6636
rect 1682 6626 1685 6679
rect 1695 6651 1698 6664
rect 1711 6657 1714 6666
rect 1718 6626 1721 6636
rect 1725 6612 1729 6933
rect 1749 6909 1752 6919
rect 1732 6883 1735 6892
rect 1748 6883 1751 6892
rect 1769 6877 1772 6890
rect 1785 6883 1788 6892
rect 1794 6881 1797 6886
rect 1732 6845 1735 6877
rect 1800 6866 1803 6919
rect 1812 6905 1813 6909
rect 1851 6907 1854 6919
rect 1806 6883 1809 6892
rect 1806 6873 1810 6877
rect 1747 6852 1750 6862
rect 1814 6852 1817 6905
rect 1827 6877 1830 6890
rect 1843 6883 1846 6892
rect 1850 6852 1853 6862
rect 1732 6756 1735 6793
rect 1857 6790 1860 6882
rect 1749 6769 1752 6779
rect 1732 6743 1735 6752
rect 1748 6743 1751 6752
rect 1769 6737 1772 6750
rect 1785 6743 1788 6752
rect 1794 6741 1797 6746
rect 1800 6726 1803 6779
rect 1812 6765 1813 6769
rect 1851 6767 1854 6779
rect 1806 6743 1809 6752
rect 1806 6733 1810 6737
rect 1747 6712 1750 6722
rect 1814 6712 1817 6765
rect 1827 6737 1830 6750
rect 1843 6743 1846 6752
rect 1850 6712 1853 6722
rect 1857 6704 1860 6742
rect 1872 6729 1876 6811
rect 1911 6739 1914 6749
rect 1894 6716 1897 6717
rect 1749 6683 1752 6693
rect 1732 6657 1735 6666
rect 1748 6657 1751 6666
rect 1769 6651 1772 6664
rect 1785 6657 1788 6666
rect 1794 6655 1797 6660
rect 1732 6619 1735 6651
rect 1800 6640 1803 6693
rect 1812 6679 1813 6683
rect 1851 6681 1854 6693
rect 1806 6657 1809 6666
rect 1806 6647 1810 6651
rect 1747 6626 1750 6636
rect 1814 6626 1817 6679
rect 1827 6651 1830 6664
rect 1843 6657 1846 6666
rect 1850 6626 1853 6636
rect 1709 6608 1713 6612
rect 1725 6607 1729 6608
rect 1709 6589 1713 6604
rect 1709 6580 1713 6585
rect 1709 6572 1713 6576
rect 1725 6576 1729 6592
rect 1741 6589 1745 6604
rect 1741 6580 1745 6585
rect 1617 6541 1620 6551
rect 1616 6515 1619 6524
rect 1637 6509 1640 6522
rect 1653 6515 1656 6524
rect 1662 6513 1665 6518
rect 1668 6498 1671 6551
rect 1680 6537 1681 6541
rect 1719 6539 1722 6551
rect 1674 6515 1677 6524
rect 1674 6505 1678 6509
rect 1615 6484 1618 6494
rect 1682 6484 1685 6537
rect 1695 6509 1698 6522
rect 1711 6515 1714 6524
rect 1718 6484 1721 6494
rect 1615 6139 1618 6151
rect 1656 6137 1657 6141
rect 1623 6115 1626 6124
rect 1639 6109 1642 6122
rect 1616 6084 1619 6094
rect 1652 6084 1655 6137
rect 1660 6115 1663 6124
rect 1659 6105 1663 6109
rect 1666 6098 1669 6151
rect 1717 6141 1720 6151
rect 1672 6113 1675 6118
rect 1681 6115 1684 6124
rect 1697 6109 1700 6122
rect 1718 6115 1721 6124
rect 1719 6084 1722 6094
rect 1457 5989 1463 6029
rect 1600 6026 1603 6056
rect 1600 6019 1603 6022
rect 1599 6018 1603 6019
rect 1600 6013 1603 6014
rect 1457 5956 1463 5985
rect 1457 5877 1463 5952
rect 1485 5927 1488 5937
rect 1468 5907 1471 5910
rect 1457 5737 1463 5873
rect 1468 5899 1471 5903
rect 1484 5901 1487 5910
rect 1505 5895 1508 5908
rect 1521 5901 1524 5910
rect 1530 5899 1533 5904
rect 1468 5848 1471 5895
rect 1536 5884 1539 5937
rect 1548 5923 1549 5927
rect 1587 5925 1590 5937
rect 1542 5901 1545 5910
rect 1542 5891 1546 5895
rect 1483 5870 1486 5880
rect 1550 5870 1553 5923
rect 1563 5895 1566 5908
rect 1579 5901 1582 5910
rect 1600 5901 1603 5910
rect 1586 5870 1589 5880
rect 1600 5863 1603 5895
rect 1608 5856 1612 6063
rect 1725 6076 1729 6572
rect 1732 6528 1735 6565
rect 1857 6562 1860 6656
rect 1872 6567 1876 6709
rect 1894 6711 1897 6712
rect 1910 6713 1913 6722
rect 1931 6707 1934 6720
rect 1947 6713 1950 6722
rect 1956 6711 1959 6716
rect 1962 6696 1965 6749
rect 1974 6735 1975 6739
rect 2013 6737 2016 6749
rect 1968 6713 1971 6722
rect 1968 6703 1972 6707
rect 1909 6682 1912 6692
rect 1976 6682 1979 6735
rect 1989 6707 1992 6720
rect 2005 6713 2008 6722
rect 2012 6682 2015 6692
rect 2019 6675 2022 6712
rect 1894 6640 1897 6670
rect 1911 6653 1914 6663
rect 1894 6627 1897 6636
rect 1910 6627 1913 6636
rect 1931 6621 1934 6634
rect 1947 6627 1950 6636
rect 1956 6625 1959 6630
rect 1894 6575 1897 6621
rect 1962 6610 1965 6663
rect 1974 6649 1975 6653
rect 2013 6651 2016 6663
rect 1968 6627 1971 6636
rect 1968 6617 1972 6621
rect 1909 6596 1912 6606
rect 1976 6596 1979 6649
rect 1989 6621 1992 6634
rect 2005 6627 2008 6636
rect 2012 6596 2015 6606
rect 2026 6603 2030 6685
rect 2330 6582 2336 6933
rect 1894 6572 1895 6575
rect 1749 6541 1752 6551
rect 1732 6515 1735 6524
rect 1748 6515 1751 6524
rect 1769 6509 1772 6522
rect 1785 6515 1788 6524
rect 1794 6513 1797 6518
rect 1800 6498 1803 6551
rect 1812 6537 1813 6541
rect 1851 6539 1854 6551
rect 1806 6515 1809 6524
rect 1806 6505 1810 6509
rect 1747 6484 1750 6494
rect 1814 6484 1817 6537
rect 1827 6509 1830 6522
rect 1843 6515 1846 6524
rect 1850 6484 1853 6494
rect 1884 6327 1888 6563
rect 1901 6544 1904 6557
rect 1908 6547 1911 6550
rect 1929 6544 1932 6557
rect 1945 6544 1948 6557
rect 1902 6495 1905 6510
rect 1922 6502 1926 6505
rect 1930 6495 1933 6510
rect 1945 6495 1948 6510
rect 1954 6502 1957 6543
rect 1973 6510 1976 6550
rect 1979 6502 1982 6543
rect 1995 6509 1998 6550
rect 2002 6544 2005 6557
rect 2019 6544 2022 6557
rect 2026 6547 2029 6550
rect 2052 6544 2056 6557
rect 2001 6495 2004 6510
rect 2020 6495 2023 6510
rect 2038 6502 2041 6506
rect 2060 6502 2063 6571
rect 2070 6554 2073 6564
rect 2078 6544 2082 6557
rect 2090 6458 2094 6530
rect 2098 6436 2101 6514
rect 2109 6472 2112 6550
rect 2162 6544 2165 6557
rect 2169 6547 2172 6550
rect 2190 6544 2193 6557
rect 2206 6544 2209 6557
rect 2163 6495 2166 6510
rect 2183 6502 2187 6505
rect 2191 6495 2194 6510
rect 2206 6495 2209 6510
rect 2215 6502 2218 6543
rect 2234 6510 2237 6550
rect 2240 6502 2243 6543
rect 2256 6509 2259 6550
rect 2263 6544 2266 6557
rect 2280 6544 2283 6557
rect 2304 6554 2308 6564
rect 2287 6547 2290 6550
rect 2313 6544 2316 6557
rect 2262 6495 2265 6510
rect 2281 6495 2284 6510
rect 2299 6502 2302 6506
rect 2163 6476 2166 6491
rect 2183 6481 2187 6484
rect 2191 6476 2194 6491
rect 2206 6476 2209 6491
rect 2102 6433 2106 6436
rect 1919 6326 1923 6394
rect 1927 6304 1930 6378
rect 1938 6340 1941 6414
rect 1938 6317 1941 6336
rect 2009 6326 2013 6394
rect 1938 6314 1958 6317
rect 1973 6304 1976 6314
rect 1931 6301 1976 6304
rect 1734 6115 1737 6124
rect 1617 6039 1620 6049
rect 1616 6013 1619 6022
rect 1637 6007 1640 6020
rect 1653 6013 1656 6022
rect 1662 6011 1665 6016
rect 1668 5996 1671 6049
rect 1680 6035 1681 6039
rect 1719 6037 1722 6049
rect 1674 6013 1677 6022
rect 1674 6003 1678 6007
rect 1615 5982 1618 5992
rect 1682 5982 1685 6035
rect 1695 6007 1698 6020
rect 1711 6013 1714 6022
rect 1718 5982 1721 5992
rect 1617 5927 1620 5937
rect 1616 5901 1619 5910
rect 1637 5895 1640 5908
rect 1653 5901 1656 5910
rect 1662 5899 1665 5904
rect 1668 5884 1671 5937
rect 1680 5923 1681 5927
rect 1719 5925 1722 5937
rect 1674 5901 1677 5910
rect 1674 5891 1678 5895
rect 1615 5870 1618 5880
rect 1682 5870 1685 5923
rect 1695 5895 1698 5908
rect 1711 5901 1714 5910
rect 1718 5870 1721 5880
rect 1592 5852 1596 5856
rect 1608 5851 1612 5852
rect 1468 5808 1471 5836
rect 1592 5833 1596 5848
rect 1592 5826 1596 5829
rect 1592 5818 1596 5822
rect 1608 5822 1612 5836
rect 1624 5833 1628 5848
rect 1624 5826 1628 5829
rect 1468 5774 1471 5804
rect 1485 5787 1488 5797
rect 1468 5759 1471 5770
rect 1484 5761 1487 5770
rect 1505 5755 1508 5768
rect 1521 5761 1524 5770
rect 1530 5759 1533 5764
rect 1536 5744 1539 5797
rect 1548 5783 1549 5787
rect 1587 5785 1590 5797
rect 1542 5761 1545 5770
rect 1542 5751 1546 5755
rect 1457 5651 1463 5733
rect 1483 5730 1486 5740
rect 1550 5730 1553 5783
rect 1600 5774 1603 5811
rect 1563 5755 1566 5768
rect 1579 5761 1582 5770
rect 1600 5761 1603 5770
rect 1586 5730 1589 5740
rect 1457 5621 1463 5647
rect 1468 5688 1471 5718
rect 1485 5701 1488 5711
rect 1468 5673 1471 5684
rect 1484 5675 1487 5684
rect 1505 5669 1508 5682
rect 1521 5675 1524 5684
rect 1530 5673 1533 5678
rect 1468 5622 1471 5669
rect 1536 5658 1539 5711
rect 1548 5697 1549 5701
rect 1587 5699 1590 5711
rect 1542 5675 1545 5684
rect 1542 5665 1546 5669
rect 1483 5644 1486 5654
rect 1550 5644 1553 5697
rect 1563 5669 1566 5682
rect 1579 5675 1582 5684
rect 1600 5675 1603 5684
rect 1586 5644 1589 5654
rect 1600 5637 1603 5669
rect 1457 5579 1463 5617
rect 1457 5509 1463 5575
rect 1468 5580 1471 5610
rect 1468 5546 1471 5576
rect 1485 5559 1488 5569
rect 1468 5531 1471 5542
rect 1484 5533 1487 5542
rect 1505 5527 1508 5540
rect 1521 5533 1524 5542
rect 1530 5531 1533 5536
rect 1536 5516 1539 5569
rect 1548 5555 1549 5559
rect 1587 5557 1590 5569
rect 1542 5533 1545 5542
rect 1542 5523 1546 5527
rect 1457 5447 1463 5505
rect 1483 5502 1486 5512
rect 1550 5502 1553 5555
rect 1600 5546 1603 5583
rect 1563 5527 1566 5540
rect 1579 5533 1582 5542
rect 1600 5533 1603 5542
rect 1586 5502 1589 5512
rect 1608 5496 1612 5818
rect 1617 5787 1620 5797
rect 1616 5761 1619 5770
rect 1637 5755 1640 5768
rect 1653 5761 1656 5770
rect 1662 5759 1665 5764
rect 1668 5744 1671 5797
rect 1680 5783 1681 5787
rect 1719 5785 1722 5797
rect 1674 5761 1677 5770
rect 1674 5751 1678 5755
rect 1615 5730 1618 5740
rect 1682 5730 1685 5783
rect 1695 5755 1698 5768
rect 1711 5761 1714 5770
rect 1718 5730 1721 5740
rect 1617 5701 1620 5711
rect 1616 5675 1619 5684
rect 1637 5669 1640 5682
rect 1653 5675 1656 5684
rect 1662 5673 1665 5678
rect 1668 5658 1671 5711
rect 1680 5697 1681 5701
rect 1719 5699 1722 5711
rect 1674 5675 1677 5684
rect 1674 5665 1678 5669
rect 1615 5644 1618 5654
rect 1682 5644 1685 5697
rect 1695 5669 1698 5682
rect 1711 5675 1714 5684
rect 1718 5644 1721 5654
rect 1725 5630 1729 6072
rect 1734 6069 1737 6109
rect 1734 6016 1737 6065
rect 1797 6030 1865 6033
rect 1973 6033 1976 6301
rect 2017 6304 2020 6378
rect 2028 6340 2031 6414
rect 2028 6317 2031 6336
rect 2090 6326 2094 6394
rect 2098 6382 2101 6432
rect 2109 6418 2112 6468
rect 2162 6429 2165 6442
rect 2169 6436 2172 6439
rect 2190 6429 2193 6442
rect 2028 6314 2048 6317
rect 2063 6304 2066 6314
rect 2021 6301 2066 6304
rect 2098 6304 2101 6378
rect 2109 6340 2112 6414
rect 2162 6412 2165 6425
rect 2169 6415 2172 6418
rect 2190 6412 2193 6425
rect 2206 6429 2209 6442
rect 2215 6443 2218 6484
rect 2234 6436 2237 6476
rect 2240 6443 2243 6484
rect 2256 6436 2259 6477
rect 2262 6476 2265 6491
rect 2281 6476 2284 6491
rect 2289 6488 2293 6498
rect 2313 6495 2316 6510
rect 2299 6480 2302 6484
rect 2313 6476 2316 6491
rect 2263 6429 2266 6442
rect 2280 6429 2283 6442
rect 2287 6436 2290 6439
rect 2206 6412 2209 6425
rect 2163 6363 2166 6378
rect 2183 6370 2187 6373
rect 2191 6363 2194 6378
rect 2206 6363 2209 6378
rect 2215 6370 2218 6411
rect 2234 6378 2237 6418
rect 2240 6370 2243 6411
rect 2256 6377 2259 6418
rect 2263 6412 2266 6425
rect 2280 6412 2283 6425
rect 2313 6429 2316 6442
rect 2287 6415 2290 6418
rect 2313 6412 2316 6425
rect 2262 6363 2265 6378
rect 2281 6363 2284 6378
rect 2299 6370 2302 6374
rect 2313 6363 2316 6378
rect 2163 6344 2166 6359
rect 2183 6349 2187 6352
rect 2191 6344 2194 6359
rect 2206 6344 2209 6359
rect 1985 6194 1989 6259
rect 1993 6172 1996 6243
rect 2004 6208 2007 6279
rect 2004 6185 2007 6204
rect 2039 6186 2042 6187
rect 2004 6182 2024 6185
rect 2039 6172 2042 6182
rect 1997 6169 2042 6172
rect 2039 6165 2042 6169
rect 2001 6161 2042 6165
rect 1869 6030 1976 6033
rect 1797 6001 1800 6030
rect 2001 6027 2004 6161
rect 2009 6062 2013 6128
rect 2017 6040 2020 6112
rect 2028 6076 2031 6148
rect 2028 6053 2031 6072
rect 2028 6050 2048 6053
rect 2060 6050 2063 6301
rect 2102 6301 2106 6304
rect 2090 6194 2094 6259
rect 2098 6247 2101 6300
rect 2109 6283 2112 6336
rect 2162 6297 2165 6310
rect 2169 6304 2172 6307
rect 2190 6297 2193 6310
rect 2098 6172 2101 6243
rect 2109 6208 2112 6279
rect 2162 6280 2165 6293
rect 2169 6283 2172 6286
rect 2190 6280 2193 6293
rect 2206 6297 2209 6310
rect 2215 6311 2218 6352
rect 2234 6304 2237 6344
rect 2240 6311 2243 6352
rect 2256 6304 2259 6345
rect 2262 6344 2265 6359
rect 2281 6344 2284 6359
rect 2299 6348 2302 6352
rect 2313 6344 2316 6359
rect 2263 6297 2266 6310
rect 2280 6297 2283 6310
rect 2287 6304 2290 6307
rect 2206 6280 2209 6293
rect 2163 6231 2166 6246
rect 2183 6238 2187 6241
rect 2191 6231 2194 6246
rect 2206 6231 2209 6246
rect 2215 6238 2218 6279
rect 2234 6246 2237 6286
rect 2240 6238 2243 6279
rect 2256 6245 2259 6286
rect 2263 6280 2266 6293
rect 2280 6280 2283 6293
rect 2313 6297 2316 6310
rect 2287 6283 2290 6286
rect 2313 6280 2316 6293
rect 2262 6231 2265 6246
rect 2281 6231 2284 6246
rect 2299 6238 2302 6242
rect 2313 6231 2316 6246
rect 2163 6212 2166 6227
rect 2183 6217 2187 6220
rect 2191 6212 2194 6227
rect 2206 6212 2209 6227
rect 2109 6185 2112 6204
rect 2109 6182 2113 6185
rect 2102 6169 2106 6172
rect 2090 6062 2094 6128
rect 2098 6116 2101 6168
rect 2109 6152 2112 6182
rect 2162 6165 2165 6178
rect 2169 6172 2172 6175
rect 2190 6165 2193 6178
rect 2063 6040 2066 6050
rect 2021 6037 2066 6040
rect 2063 6034 2066 6037
rect 2098 6040 2101 6112
rect 2109 6076 2112 6148
rect 2162 6148 2165 6161
rect 2169 6151 2172 6154
rect 2190 6148 2193 6161
rect 2206 6165 2209 6178
rect 2215 6179 2218 6220
rect 2234 6172 2237 6212
rect 2240 6179 2243 6220
rect 2256 6172 2259 6213
rect 2262 6212 2265 6227
rect 2281 6212 2284 6227
rect 2299 6216 2302 6220
rect 2313 6212 2316 6227
rect 2263 6165 2266 6178
rect 2280 6165 2283 6178
rect 2287 6172 2290 6175
rect 2206 6148 2209 6161
rect 2163 6099 2166 6114
rect 2183 6106 2187 6109
rect 2191 6099 2194 6114
rect 2206 6099 2209 6114
rect 2215 6106 2218 6147
rect 2234 6114 2237 6154
rect 2240 6106 2243 6147
rect 2256 6113 2259 6154
rect 2263 6148 2266 6161
rect 2280 6148 2283 6161
rect 2302 6158 2306 6168
rect 2313 6165 2316 6178
rect 2287 6151 2290 6154
rect 2313 6148 2316 6161
rect 2262 6099 2265 6114
rect 2281 6099 2284 6114
rect 2299 6106 2302 6110
rect 2313 6099 2316 6114
rect 2163 6080 2166 6095
rect 2183 6085 2187 6088
rect 2191 6080 2194 6095
rect 2206 6080 2209 6095
rect 2109 6053 2112 6072
rect 2109 6050 2129 6053
rect 2144 6040 2147 6050
rect 2102 6037 2147 6040
rect 1929 6023 2004 6027
rect 2061 6029 2066 6034
rect 1814 6006 1817 6016
rect 1797 5993 1800 5997
rect 1797 5983 1800 5989
rect 1796 5980 1800 5983
rect 1797 5978 1800 5980
rect 1813 5980 1816 5989
rect 1834 5974 1837 5987
rect 1850 5980 1853 5989
rect 1859 5978 1862 5983
rect 1865 5963 1868 6016
rect 1877 6002 1878 6006
rect 1916 6004 1919 6016
rect 1871 5980 1874 5989
rect 1871 5970 1875 5974
rect 1812 5949 1815 5959
rect 1879 5949 1882 6002
rect 1929 6001 1932 6023
rect 1946 6006 1949 6016
rect 1892 5974 1895 5987
rect 1908 5980 1911 5989
rect 1929 5983 1932 5989
rect 1925 5980 1932 5983
rect 1929 5978 1932 5980
rect 1945 5980 1948 5989
rect 1966 5974 1969 5987
rect 1982 5980 1985 5989
rect 1991 5978 1994 5983
rect 1997 5963 2000 6016
rect 2009 6002 2010 6006
rect 2048 6004 2051 6016
rect 2003 5980 2006 5989
rect 2003 5970 2007 5974
rect 1915 5949 1918 5959
rect 1944 5949 1947 5959
rect 2011 5949 2014 6002
rect 2061 5993 2064 6029
rect 2144 6026 2147 6037
rect 2162 6033 2165 6046
rect 2169 6040 2172 6043
rect 2190 6033 2193 6046
rect 2206 6033 2209 6046
rect 2215 6047 2218 6088
rect 2234 6040 2237 6080
rect 2240 6047 2243 6088
rect 2256 6040 2259 6081
rect 2262 6080 2265 6095
rect 2281 6080 2284 6095
rect 2299 6084 2302 6088
rect 2313 6080 2316 6095
rect 2263 6033 2266 6046
rect 2280 6033 2283 6046
rect 2287 6040 2290 6043
rect 2313 6033 2316 6046
rect 2144 6023 2196 6026
rect 2078 6006 2081 6016
rect 2024 5974 2027 5987
rect 2040 5980 2043 5989
rect 2061 5983 2064 5989
rect 2057 5980 2064 5983
rect 2061 5978 2064 5980
rect 2077 5980 2080 5989
rect 2098 5974 2101 5987
rect 2114 5980 2117 5989
rect 2123 5978 2126 5983
rect 2129 5963 2132 6016
rect 2141 6002 2142 6006
rect 2180 6004 2183 6016
rect 2135 5980 2138 5989
rect 2135 5970 2139 5974
rect 2047 5949 2050 5959
rect 2076 5949 2079 5959
rect 2143 5949 2146 6002
rect 2193 5993 2196 6023
rect 2210 6006 2213 6016
rect 2156 5974 2159 5987
rect 2172 5980 2175 5989
rect 2193 5983 2196 5989
rect 2189 5980 2196 5983
rect 2193 5978 2196 5980
rect 2209 5980 2212 5989
rect 2230 5974 2233 5987
rect 2246 5980 2249 5989
rect 2255 5978 2258 5983
rect 2261 5963 2264 6016
rect 2273 6002 2274 6006
rect 2312 6004 2315 6016
rect 2267 5980 2270 5989
rect 2267 5970 2271 5974
rect 2179 5949 2182 5959
rect 2208 5949 2211 5959
rect 2275 5949 2278 6002
rect 2288 5974 2291 5987
rect 2304 5980 2307 5989
rect 2311 5949 2314 5959
rect 1749 5927 1752 5937
rect 1732 5901 1735 5910
rect 1748 5901 1751 5910
rect 1769 5895 1772 5908
rect 1785 5901 1788 5910
rect 1794 5899 1797 5904
rect 1732 5863 1735 5895
rect 1800 5884 1803 5937
rect 1812 5923 1813 5927
rect 1851 5925 1854 5937
rect 1806 5901 1809 5910
rect 1806 5891 1810 5895
rect 1747 5870 1750 5880
rect 1814 5870 1817 5923
rect 1827 5895 1830 5908
rect 1843 5901 1846 5910
rect 1850 5870 1853 5880
rect 1732 5774 1735 5811
rect 1857 5808 1860 5900
rect 1749 5787 1752 5797
rect 1732 5761 1735 5770
rect 1748 5761 1751 5770
rect 1769 5755 1772 5768
rect 1785 5761 1788 5770
rect 1794 5759 1797 5764
rect 1800 5744 1803 5797
rect 1812 5783 1813 5787
rect 1851 5785 1854 5797
rect 1806 5761 1809 5770
rect 1806 5751 1810 5755
rect 1747 5730 1750 5740
rect 1814 5730 1817 5783
rect 1827 5755 1830 5768
rect 1843 5761 1846 5770
rect 1850 5730 1853 5740
rect 1857 5722 1860 5760
rect 1872 5747 1876 5829
rect 1911 5757 1914 5767
rect 1894 5734 1897 5735
rect 1749 5701 1752 5711
rect 1732 5675 1735 5684
rect 1748 5675 1751 5684
rect 1769 5669 1772 5682
rect 1785 5675 1788 5684
rect 1794 5673 1797 5678
rect 1732 5637 1735 5669
rect 1800 5658 1803 5711
rect 1812 5697 1813 5701
rect 1851 5699 1854 5711
rect 1806 5675 1809 5684
rect 1806 5665 1810 5669
rect 1747 5644 1750 5654
rect 1814 5644 1817 5697
rect 1827 5669 1830 5682
rect 1843 5675 1846 5684
rect 1850 5644 1853 5654
rect 1709 5626 1713 5630
rect 1725 5625 1729 5626
rect 1709 5607 1713 5622
rect 1709 5599 1713 5603
rect 1709 5590 1713 5595
rect 1725 5594 1729 5610
rect 1741 5607 1745 5622
rect 1741 5599 1745 5603
rect 1617 5559 1620 5569
rect 1616 5533 1619 5542
rect 1637 5527 1640 5540
rect 1653 5533 1656 5542
rect 1662 5531 1665 5536
rect 1668 5516 1671 5569
rect 1680 5555 1681 5559
rect 1719 5557 1722 5569
rect 1674 5533 1677 5542
rect 1674 5523 1678 5527
rect 1615 5502 1618 5512
rect 1682 5502 1685 5555
rect 1695 5527 1698 5540
rect 1711 5533 1714 5542
rect 1718 5502 1721 5512
rect 1725 5495 1729 5590
rect 1732 5546 1735 5583
rect 1857 5580 1860 5674
rect 1872 5585 1876 5727
rect 1894 5729 1897 5730
rect 1910 5731 1913 5740
rect 1931 5725 1934 5738
rect 1947 5731 1950 5740
rect 1956 5729 1959 5734
rect 1962 5714 1965 5767
rect 1974 5753 1975 5757
rect 2013 5755 2016 5767
rect 1968 5731 1971 5740
rect 1968 5721 1972 5725
rect 1909 5700 1912 5710
rect 1976 5700 1979 5753
rect 1989 5725 1992 5738
rect 2005 5731 2008 5740
rect 2012 5700 2015 5710
rect 2019 5693 2022 5730
rect 1894 5658 1897 5688
rect 1911 5671 1914 5681
rect 1894 5645 1897 5654
rect 1910 5645 1913 5654
rect 1931 5639 1934 5652
rect 1947 5645 1950 5654
rect 1956 5643 1959 5648
rect 1894 5593 1897 5639
rect 1962 5628 1965 5681
rect 1974 5667 1975 5671
rect 2013 5669 2016 5681
rect 1968 5645 1971 5654
rect 1968 5635 1972 5639
rect 1909 5614 1912 5624
rect 1976 5614 1979 5667
rect 1989 5639 1992 5652
rect 2005 5645 2008 5654
rect 2012 5614 2015 5624
rect 2026 5621 2030 5703
rect 2330 5600 2336 6578
rect 1894 5590 1895 5593
rect 1749 5559 1752 5569
rect 1732 5533 1735 5542
rect 1748 5533 1751 5542
rect 1769 5527 1772 5540
rect 1785 5533 1788 5542
rect 1794 5531 1797 5536
rect 1800 5516 1803 5569
rect 1812 5555 1813 5559
rect 1851 5557 1854 5569
rect 1806 5533 1809 5542
rect 1806 5523 1810 5527
rect 1747 5502 1750 5512
rect 1814 5502 1817 5555
rect 1827 5527 1830 5540
rect 1843 5533 1846 5542
rect 1850 5502 1853 5512
rect 1608 5490 1612 5491
rect 1725 5489 1729 5490
rect 1457 5315 1463 5443
rect 1457 5281 1463 5311
rect 1457 5183 1463 5277
rect 1492 5297 1496 5481
rect 1492 5249 1496 5293
rect 1500 5472 1504 5481
rect 1500 5342 1504 5468
rect 1500 5281 1504 5338
rect 1500 5212 1504 5277
rect 1507 5422 1512 5481
rect 1507 5292 1512 5418
rect 1680 5391 1684 5428
rect 1754 5371 1758 5441
rect 1762 5349 1765 5425
rect 1773 5385 1776 5461
rect 1844 5440 1846 5444
rect 1773 5362 1776 5381
rect 1789 5368 1833 5371
rect 1830 5363 1833 5368
rect 1773 5359 1793 5362
rect 1808 5349 1811 5359
rect 1766 5346 1811 5349
rect 1507 5249 1512 5288
rect 1575 5261 1579 5302
rect 1754 5241 1758 5311
rect 1762 5219 1765 5295
rect 1773 5255 1776 5331
rect 1773 5232 1776 5251
rect 1789 5238 1811 5241
rect 1808 5233 1811 5238
rect 1830 5233 1833 5359
rect 1842 5314 1846 5440
rect 1884 5345 1888 5581
rect 1901 5562 1904 5575
rect 1908 5565 1911 5568
rect 1929 5562 1932 5575
rect 1945 5562 1948 5575
rect 1902 5513 1905 5528
rect 1922 5520 1926 5523
rect 1930 5513 1933 5528
rect 1945 5513 1948 5528
rect 1954 5520 1957 5561
rect 1973 5528 1976 5568
rect 1979 5520 1982 5561
rect 1995 5527 1998 5568
rect 2002 5562 2005 5575
rect 2019 5562 2022 5575
rect 2026 5565 2029 5568
rect 2052 5562 2056 5575
rect 2001 5513 2004 5528
rect 2020 5513 2023 5528
rect 2038 5520 2041 5524
rect 2060 5520 2063 5589
rect 2070 5572 2073 5582
rect 2078 5562 2082 5575
rect 2090 5476 2094 5548
rect 2098 5454 2101 5532
rect 2109 5490 2112 5568
rect 2162 5562 2165 5575
rect 2169 5565 2172 5568
rect 2190 5562 2193 5575
rect 2206 5562 2209 5575
rect 2163 5513 2166 5528
rect 2183 5520 2187 5523
rect 2191 5513 2194 5528
rect 2206 5513 2209 5528
rect 2215 5520 2218 5561
rect 2234 5528 2237 5568
rect 2240 5520 2243 5561
rect 2256 5527 2259 5568
rect 2263 5562 2266 5575
rect 2280 5562 2283 5575
rect 2304 5572 2308 5582
rect 2287 5565 2290 5568
rect 2313 5562 2316 5575
rect 2262 5513 2265 5528
rect 2281 5513 2284 5528
rect 2299 5520 2302 5524
rect 2163 5494 2166 5509
rect 2183 5499 2187 5502
rect 2191 5494 2194 5509
rect 2206 5494 2209 5509
rect 2102 5451 2106 5454
rect 1919 5344 1923 5412
rect 1927 5322 1930 5396
rect 1938 5358 1941 5432
rect 1938 5335 1941 5354
rect 2009 5344 2013 5412
rect 1938 5332 1958 5335
rect 1973 5322 1976 5332
rect 1931 5319 1976 5322
rect 1846 5310 1857 5314
rect 1842 5296 1857 5310
rect 1773 5229 1793 5232
rect 1812 5229 1833 5233
rect 1808 5219 1811 5229
rect 1766 5216 1811 5219
rect 1808 5194 1811 5216
rect 1457 5109 1463 5179
rect 1457 5051 1463 5105
rect 1584 5085 1588 5090
rect 1608 5085 1612 5173
rect 1615 5157 1618 5169
rect 1656 5155 1657 5159
rect 1623 5133 1626 5142
rect 1639 5127 1642 5140
rect 1616 5102 1619 5112
rect 1652 5102 1655 5155
rect 1660 5133 1663 5142
rect 1659 5123 1663 5127
rect 1666 5116 1669 5169
rect 1717 5159 1720 5169
rect 1672 5131 1675 5136
rect 1681 5133 1684 5142
rect 1697 5127 1700 5140
rect 1718 5133 1721 5142
rect 1719 5102 1722 5112
rect 1457 5007 1463 5047
rect 1600 5044 1603 5074
rect 1600 5037 1603 5040
rect 1600 5031 1603 5033
rect 1457 4974 1463 5003
rect 1608 4981 1612 5081
rect 1725 5094 1729 5174
rect 1734 5133 1737 5142
rect 1617 5057 1620 5067
rect 1616 5031 1619 5040
rect 1637 5025 1640 5038
rect 1653 5031 1656 5040
rect 1662 5029 1665 5034
rect 1668 5014 1671 5067
rect 1680 5053 1681 5057
rect 1719 5055 1722 5067
rect 1674 5031 1677 5040
rect 1674 5021 1678 5025
rect 1615 5000 1618 5010
rect 1682 5000 1685 5053
rect 1695 5025 1698 5038
rect 1711 5031 1714 5040
rect 1718 5000 1721 5010
rect 1725 4981 1729 5090
rect 1734 5087 1737 5127
rect 1734 5034 1737 5083
rect 1807 5073 1811 5190
rect 1457 4934 1463 4970
rect 1457 4854 1463 4930
rect 1745 4870 1749 5069
rect 1844 5064 1857 5296
rect 1756 4880 1761 5056
rect 1797 5048 1865 5051
rect 1973 5051 1976 5319
rect 2017 5322 2020 5396
rect 2028 5358 2031 5432
rect 2028 5335 2031 5354
rect 2090 5344 2094 5412
rect 2098 5400 2101 5450
rect 2109 5436 2112 5486
rect 2162 5447 2165 5460
rect 2169 5454 2172 5457
rect 2190 5447 2193 5460
rect 2028 5332 2048 5335
rect 2063 5322 2066 5332
rect 2021 5319 2066 5322
rect 2098 5322 2101 5396
rect 2109 5358 2112 5432
rect 2162 5430 2165 5443
rect 2169 5433 2172 5436
rect 2190 5430 2193 5443
rect 2206 5447 2209 5460
rect 2215 5461 2218 5502
rect 2234 5454 2237 5494
rect 2240 5461 2243 5502
rect 2256 5454 2259 5495
rect 2262 5494 2265 5509
rect 2281 5494 2284 5509
rect 2289 5506 2293 5516
rect 2313 5513 2316 5528
rect 2299 5498 2302 5502
rect 2313 5494 2316 5509
rect 2263 5447 2266 5460
rect 2280 5447 2283 5460
rect 2287 5454 2290 5457
rect 2206 5430 2209 5443
rect 2163 5381 2166 5396
rect 2183 5388 2187 5391
rect 2191 5381 2194 5396
rect 2206 5381 2209 5396
rect 2215 5388 2218 5429
rect 2234 5396 2237 5436
rect 2240 5388 2243 5429
rect 2256 5395 2259 5436
rect 2263 5430 2266 5443
rect 2280 5430 2283 5443
rect 2313 5447 2316 5460
rect 2287 5433 2290 5436
rect 2313 5430 2316 5443
rect 2262 5381 2265 5396
rect 2281 5381 2284 5396
rect 2299 5388 2302 5392
rect 2313 5381 2316 5396
rect 2163 5362 2166 5377
rect 2183 5367 2187 5370
rect 2191 5362 2194 5377
rect 2206 5362 2209 5377
rect 1985 5212 1989 5277
rect 1993 5190 1996 5261
rect 2004 5226 2007 5297
rect 2004 5203 2007 5222
rect 2039 5204 2042 5205
rect 2004 5200 2024 5203
rect 2039 5190 2042 5200
rect 1997 5187 2042 5190
rect 2039 5183 2042 5187
rect 2001 5179 2042 5183
rect 1869 5048 1976 5051
rect 1797 5019 1800 5048
rect 2001 5045 2004 5179
rect 2009 5080 2013 5146
rect 2017 5058 2020 5130
rect 2028 5094 2031 5166
rect 2028 5071 2031 5090
rect 2028 5068 2048 5071
rect 2060 5068 2063 5319
rect 2102 5319 2106 5322
rect 2090 5212 2094 5277
rect 2098 5265 2101 5318
rect 2109 5301 2112 5354
rect 2162 5315 2165 5328
rect 2169 5322 2172 5325
rect 2190 5315 2193 5328
rect 2098 5190 2101 5261
rect 2109 5226 2112 5297
rect 2162 5298 2165 5311
rect 2169 5301 2172 5304
rect 2190 5298 2193 5311
rect 2206 5315 2209 5328
rect 2215 5329 2218 5370
rect 2234 5322 2237 5362
rect 2240 5329 2243 5370
rect 2256 5322 2259 5363
rect 2262 5362 2265 5377
rect 2281 5362 2284 5377
rect 2299 5366 2302 5370
rect 2313 5362 2316 5377
rect 2263 5315 2266 5328
rect 2280 5315 2283 5328
rect 2287 5322 2290 5325
rect 2206 5298 2209 5311
rect 2163 5249 2166 5264
rect 2183 5256 2187 5259
rect 2191 5249 2194 5264
rect 2206 5249 2209 5264
rect 2215 5256 2218 5297
rect 2234 5264 2237 5304
rect 2240 5256 2243 5297
rect 2256 5263 2259 5304
rect 2263 5298 2266 5311
rect 2280 5298 2283 5311
rect 2313 5315 2316 5328
rect 2287 5301 2290 5304
rect 2313 5298 2316 5311
rect 2262 5249 2265 5264
rect 2281 5249 2284 5264
rect 2299 5256 2302 5260
rect 2313 5249 2316 5264
rect 2163 5230 2166 5245
rect 2183 5235 2187 5238
rect 2191 5230 2194 5245
rect 2206 5230 2209 5245
rect 2109 5203 2112 5222
rect 2109 5200 2113 5203
rect 2102 5187 2106 5190
rect 2090 5080 2094 5146
rect 2098 5134 2101 5186
rect 2109 5170 2112 5200
rect 2162 5183 2165 5196
rect 2169 5190 2172 5193
rect 2190 5183 2193 5196
rect 2063 5058 2066 5068
rect 2021 5055 2066 5058
rect 2063 5052 2066 5055
rect 2098 5058 2101 5130
rect 2109 5094 2112 5166
rect 2162 5166 2165 5179
rect 2169 5169 2172 5172
rect 2190 5166 2193 5179
rect 2206 5183 2209 5196
rect 2215 5197 2218 5238
rect 2234 5190 2237 5230
rect 2240 5197 2243 5238
rect 2256 5190 2259 5231
rect 2262 5230 2265 5245
rect 2281 5230 2284 5245
rect 2299 5234 2302 5238
rect 2313 5230 2316 5245
rect 2263 5183 2266 5196
rect 2280 5183 2283 5196
rect 2287 5190 2290 5193
rect 2206 5166 2209 5179
rect 2163 5117 2166 5132
rect 2183 5124 2187 5127
rect 2191 5117 2194 5132
rect 2206 5117 2209 5132
rect 2215 5124 2218 5165
rect 2234 5132 2237 5172
rect 2240 5124 2243 5165
rect 2256 5131 2259 5172
rect 2263 5166 2266 5179
rect 2280 5166 2283 5179
rect 2302 5176 2306 5186
rect 2313 5183 2316 5196
rect 2287 5169 2290 5172
rect 2313 5166 2316 5179
rect 2262 5117 2265 5132
rect 2281 5117 2284 5132
rect 2299 5124 2302 5128
rect 2313 5117 2316 5132
rect 2163 5098 2166 5113
rect 2183 5103 2187 5106
rect 2191 5098 2194 5113
rect 2206 5098 2209 5113
rect 2109 5071 2112 5090
rect 2109 5068 2129 5071
rect 2144 5058 2147 5068
rect 2102 5055 2147 5058
rect 1929 5041 2004 5045
rect 2061 5047 2066 5052
rect 1814 5024 1817 5034
rect 1797 5011 1800 5015
rect 1797 5001 1800 5007
rect 1796 4998 1800 5001
rect 1797 4996 1800 4998
rect 1813 4998 1816 5007
rect 1834 4992 1837 5005
rect 1850 4998 1853 5007
rect 1859 4996 1862 5001
rect 1865 4981 1868 5034
rect 1877 5020 1878 5024
rect 1916 5022 1919 5034
rect 1871 4998 1874 5007
rect 1871 4988 1875 4992
rect 1812 4967 1815 4977
rect 1879 4967 1882 5020
rect 1929 5019 1932 5041
rect 1946 5024 1949 5034
rect 1892 4992 1895 5005
rect 1908 4998 1911 5007
rect 1929 5001 1932 5007
rect 1925 4998 1932 5001
rect 1929 4996 1932 4998
rect 1945 4998 1948 5007
rect 1966 4992 1969 5005
rect 1982 4998 1985 5007
rect 1991 4996 1994 5001
rect 1997 4981 2000 5034
rect 2009 5020 2010 5024
rect 2048 5022 2051 5034
rect 2003 4998 2006 5007
rect 2003 4988 2007 4992
rect 1915 4967 1918 4977
rect 1944 4967 1947 4977
rect 2011 4967 2014 5020
rect 2061 5011 2064 5047
rect 2144 5044 2147 5055
rect 2162 5051 2165 5064
rect 2169 5058 2172 5061
rect 2190 5051 2193 5064
rect 2206 5051 2209 5064
rect 2215 5065 2218 5106
rect 2234 5058 2237 5098
rect 2240 5065 2243 5106
rect 2256 5058 2259 5099
rect 2262 5098 2265 5113
rect 2281 5098 2284 5113
rect 2299 5102 2302 5106
rect 2313 5098 2316 5113
rect 2263 5051 2266 5064
rect 2280 5051 2283 5064
rect 2287 5058 2290 5061
rect 2313 5051 2316 5064
rect 2144 5041 2196 5044
rect 2078 5024 2081 5034
rect 2024 4992 2027 5005
rect 2040 4998 2043 5007
rect 2061 5001 2064 5007
rect 2057 4998 2064 5001
rect 2061 4996 2064 4998
rect 2077 4998 2080 5007
rect 2098 4992 2101 5005
rect 2114 4998 2117 5007
rect 2123 4996 2126 5001
rect 2129 4981 2132 5034
rect 2141 5020 2142 5024
rect 2180 5022 2183 5034
rect 2135 4998 2138 5007
rect 2135 4988 2139 4992
rect 2047 4967 2050 4977
rect 2076 4967 2079 4977
rect 2143 4967 2146 5020
rect 2193 5011 2196 5041
rect 2210 5024 2213 5034
rect 2156 4992 2159 5005
rect 2172 4998 2175 5007
rect 2193 5001 2196 5007
rect 2189 4998 2196 5001
rect 2193 4996 2196 4998
rect 2209 4998 2212 5007
rect 2230 4992 2233 5005
rect 2246 4998 2249 5007
rect 2255 4996 2258 5001
rect 2261 4981 2264 5034
rect 2273 5020 2274 5024
rect 2312 5022 2315 5034
rect 2267 4998 2270 5007
rect 2267 4988 2271 4992
rect 2179 4967 2182 4977
rect 2208 4967 2211 4977
rect 2275 4967 2278 5020
rect 2288 4992 2291 5005
rect 2304 4998 2307 5007
rect 2321 4996 2325 4997
rect 2311 4967 2314 4977
rect 1482 4845 1537 4851
rect 1790 4847 1845 4848
rect 617 4810 618 4814
rect 622 4810 623 4814
rect 627 4810 628 4814
rect 632 4810 633 4814
rect 637 4810 638 4814
rect 642 4810 643 4814
rect 613 4809 647 4810
rect 617 4805 618 4809
rect 622 4805 623 4809
rect 627 4805 628 4809
rect 632 4805 633 4809
rect 637 4805 638 4809
rect 642 4805 643 4809
rect 613 4804 647 4805
rect 617 4800 618 4804
rect 622 4800 623 4804
rect 627 4800 628 4804
rect 632 4800 633 4804
rect 637 4800 638 4804
rect 642 4800 643 4804
rect 613 4799 647 4800
rect 617 4795 618 4799
rect 622 4795 623 4799
rect 627 4795 628 4799
rect 632 4795 633 4799
rect 637 4795 638 4799
rect 642 4795 643 4799
rect 663 4810 664 4814
rect 668 4810 669 4814
rect 673 4810 674 4814
rect 678 4810 679 4814
rect 683 4810 684 4814
rect 688 4810 689 4814
rect 659 4809 693 4810
rect 663 4805 664 4809
rect 668 4805 669 4809
rect 673 4805 674 4809
rect 678 4805 679 4809
rect 683 4805 684 4809
rect 688 4805 689 4809
rect 659 4804 693 4805
rect 663 4800 664 4804
rect 668 4800 669 4804
rect 673 4800 674 4804
rect 678 4800 679 4804
rect 683 4800 684 4804
rect 688 4800 689 4804
rect 659 4799 693 4800
rect 663 4795 664 4799
rect 668 4795 669 4799
rect 673 4795 674 4799
rect 678 4795 679 4799
rect 683 4795 684 4799
rect 688 4795 689 4799
rect 617 4781 618 4785
rect 622 4781 623 4785
rect 627 4781 628 4785
rect 632 4781 633 4785
rect 637 4781 638 4785
rect 642 4781 643 4785
rect 613 4780 647 4781
rect 617 4776 618 4780
rect 622 4776 623 4780
rect 627 4776 628 4780
rect 632 4776 633 4780
rect 637 4776 638 4780
rect 642 4776 643 4780
rect 613 4775 647 4776
rect 617 4771 618 4775
rect 622 4771 623 4775
rect 627 4771 628 4775
rect 632 4771 633 4775
rect 637 4771 638 4775
rect 642 4771 643 4775
rect 613 4770 647 4771
rect 617 4766 618 4770
rect 622 4766 623 4770
rect 627 4766 628 4770
rect 632 4766 633 4770
rect 637 4766 638 4770
rect 642 4766 643 4770
rect 663 4781 664 4785
rect 668 4781 669 4785
rect 673 4781 674 4785
rect 678 4781 679 4785
rect 683 4781 684 4785
rect 688 4781 689 4785
rect 659 4780 693 4781
rect 663 4776 664 4780
rect 668 4776 669 4780
rect 673 4776 674 4780
rect 678 4776 679 4780
rect 683 4776 684 4780
rect 688 4776 689 4780
rect 659 4775 693 4776
rect 663 4771 664 4775
rect 668 4771 669 4775
rect 673 4771 674 4775
rect 678 4771 679 4775
rect 683 4771 684 4775
rect 688 4771 689 4775
rect 659 4770 693 4771
rect 663 4766 664 4770
rect 668 4766 669 4770
rect 673 4766 674 4770
rect 678 4766 679 4770
rect 683 4766 684 4770
rect 688 4766 689 4770
rect 617 4752 618 4756
rect 622 4752 623 4756
rect 627 4752 628 4756
rect 632 4752 633 4756
rect 637 4752 638 4756
rect 642 4752 643 4756
rect 613 4751 647 4752
rect 617 4747 618 4751
rect 622 4747 623 4751
rect 627 4747 628 4751
rect 632 4747 633 4751
rect 637 4747 638 4751
rect 642 4747 643 4751
rect 613 4746 647 4747
rect 617 4742 618 4746
rect 622 4742 623 4746
rect 627 4742 628 4746
rect 632 4742 633 4746
rect 637 4742 638 4746
rect 642 4742 643 4746
rect 613 4741 647 4742
rect 617 4737 618 4741
rect 622 4737 623 4741
rect 627 4737 628 4741
rect 632 4737 633 4741
rect 637 4737 638 4741
rect 642 4737 643 4741
rect 663 4752 664 4756
rect 668 4752 669 4756
rect 673 4752 674 4756
rect 678 4752 679 4756
rect 683 4752 684 4756
rect 688 4752 689 4756
rect 659 4751 693 4752
rect 663 4747 664 4751
rect 668 4747 669 4751
rect 673 4747 674 4751
rect 678 4747 679 4751
rect 683 4747 684 4751
rect 688 4747 689 4751
rect 659 4746 693 4747
rect 663 4742 664 4746
rect 668 4742 669 4746
rect 673 4742 674 4746
rect 678 4742 679 4746
rect 683 4742 684 4746
rect 688 4742 689 4746
rect 659 4741 693 4742
rect 663 4737 664 4741
rect 668 4737 669 4741
rect 673 4737 674 4741
rect 678 4737 679 4741
rect 683 4737 684 4741
rect 688 4737 689 4741
rect 1482 4710 1538 4845
rect 1790 4708 1845 4843
rect 1790 4706 1793 4708
rect 2119 4707 2132 4866
rect 2146 4709 2151 4876
rect 2330 4862 2336 5596
rect 2342 6852 2348 6933
rect 2342 6712 2348 6848
rect 2342 6682 2348 6708
rect 2342 6626 2348 6678
rect 2342 6596 2348 6622
rect 2342 6484 2348 6592
rect 2342 6084 2348 6480
rect 2342 5982 2348 6080
rect 2342 5949 2348 5978
rect 2342 5870 2348 5945
rect 2342 5730 2348 5866
rect 2342 5700 2348 5726
rect 2342 5644 2348 5696
rect 2342 5614 2348 5640
rect 2342 5502 2348 5610
rect 2342 5102 2348 5498
rect 2342 5000 2348 5098
rect 2342 4967 2348 4996
rect 2342 4817 2348 4963
rect 2354 6923 2360 6933
rect 2354 6783 2360 6919
rect 2354 6753 2360 6779
rect 2354 6697 2360 6749
rect 2354 6667 2360 6693
rect 2354 6554 2360 6663
rect 2354 6155 2360 6550
rect 2354 6053 2360 6151
rect 2354 6020 2360 6049
rect 2354 5941 2360 6016
rect 2354 5801 2360 5937
rect 2354 5771 2360 5797
rect 2354 5715 2360 5767
rect 2354 5685 2360 5711
rect 2354 5572 2360 5681
rect 2354 5173 2360 5568
rect 2354 5071 2360 5169
rect 2354 5038 2360 5067
rect 2354 4825 2360 5034
rect 2354 4813 2360 4821
rect 2366 6568 2372 6933
rect 2366 6436 2372 6564
rect 2366 6422 2372 6432
rect 2366 6304 2372 6418
rect 2366 6290 2372 6300
rect 2366 6172 2372 6286
rect 2366 6040 2372 6168
rect 2366 5586 2372 6036
rect 2366 5454 2372 5582
rect 2366 5440 2372 5450
rect 2366 5322 2372 5436
rect 2366 5308 2372 5318
rect 2366 5190 2372 5304
rect 2366 5058 2372 5186
rect 2366 4832 2372 5054
rect 2366 4813 2372 4828
rect 2378 6576 2384 6933
rect 2378 6502 2384 6572
rect 2378 6370 2384 6498
rect 2378 6356 2384 6366
rect 2378 6238 2384 6352
rect 2378 6224 2384 6234
rect 2378 6106 2384 6220
rect 2378 6092 2384 6102
rect 2378 5594 2384 6088
rect 2378 5520 2384 5590
rect 2378 5388 2384 5516
rect 2378 5374 2384 5384
rect 2378 5256 2384 5370
rect 2378 5242 2384 5252
rect 2378 5124 2384 5238
rect 2378 5110 2384 5120
rect 2378 4839 2384 5106
rect 2390 6916 2396 6933
rect 2390 6776 2396 6912
rect 2390 6746 2396 6772
rect 2390 6690 2396 6742
rect 2390 6660 2396 6686
rect 2390 6548 2396 6656
rect 2390 6495 2396 6544
rect 2390 6363 2396 6491
rect 2390 6231 2396 6359
rect 2390 6148 2396 6227
rect 2390 6099 2396 6144
rect 2390 6046 2396 6095
rect 2390 6013 2396 6042
rect 2390 5934 2396 6009
rect 2390 5794 2396 5930
rect 2390 5764 2396 5790
rect 2390 5708 2396 5760
rect 2390 5678 2396 5704
rect 2390 5566 2396 5674
rect 2390 5513 2396 5562
rect 2390 5381 2396 5509
rect 2390 5249 2396 5377
rect 2390 5166 2396 5245
rect 2390 5117 2396 5162
rect 2390 5064 2396 5113
rect 2390 5031 2396 5060
rect 2390 4848 2396 5027
rect 2402 6859 2408 6933
rect 2430 6909 2433 6919
rect 2413 6889 2416 6892
rect 2402 6719 2408 6855
rect 2413 6881 2416 6885
rect 2429 6883 2432 6892
rect 2450 6877 2453 6890
rect 2466 6883 2469 6892
rect 2475 6881 2478 6886
rect 2413 6830 2416 6877
rect 2481 6866 2484 6919
rect 2493 6905 2494 6909
rect 2532 6907 2535 6919
rect 2487 6883 2490 6892
rect 2487 6873 2491 6877
rect 2428 6852 2431 6862
rect 2495 6852 2498 6905
rect 2508 6877 2511 6890
rect 2524 6883 2527 6892
rect 2545 6883 2548 6892
rect 2531 6852 2534 6862
rect 2545 6845 2548 6877
rect 2553 6838 2557 6933
rect 2562 6909 2565 6919
rect 2561 6883 2564 6892
rect 2582 6877 2585 6890
rect 2598 6883 2601 6892
rect 2607 6881 2610 6886
rect 2613 6866 2616 6919
rect 2625 6905 2626 6909
rect 2664 6907 2667 6919
rect 2619 6883 2622 6892
rect 2619 6873 2623 6877
rect 2560 6852 2563 6862
rect 2627 6852 2630 6905
rect 2640 6877 2643 6890
rect 2656 6883 2659 6892
rect 2663 6852 2666 6862
rect 2537 6834 2541 6838
rect 2553 6833 2557 6834
rect 2413 6790 2416 6818
rect 2537 6815 2541 6830
rect 2537 6808 2541 6811
rect 2537 6800 2541 6804
rect 2553 6804 2557 6818
rect 2569 6815 2573 6830
rect 2569 6808 2573 6811
rect 2413 6756 2416 6786
rect 2430 6769 2433 6779
rect 2413 6741 2416 6752
rect 2429 6743 2432 6752
rect 2450 6737 2453 6750
rect 2466 6743 2469 6752
rect 2475 6741 2478 6746
rect 2481 6726 2484 6779
rect 2493 6765 2494 6769
rect 2532 6767 2535 6779
rect 2487 6743 2490 6752
rect 2487 6733 2491 6737
rect 2402 6633 2408 6715
rect 2428 6712 2431 6722
rect 2495 6712 2498 6765
rect 2545 6756 2548 6793
rect 2508 6737 2511 6750
rect 2524 6743 2527 6752
rect 2545 6743 2548 6752
rect 2531 6712 2534 6722
rect 2402 6603 2408 6629
rect 2413 6670 2416 6700
rect 2430 6683 2433 6693
rect 2413 6655 2416 6666
rect 2429 6657 2432 6666
rect 2450 6651 2453 6664
rect 2466 6657 2469 6666
rect 2475 6655 2478 6660
rect 2413 6604 2416 6651
rect 2481 6640 2484 6693
rect 2493 6679 2494 6683
rect 2532 6681 2535 6693
rect 2487 6657 2490 6666
rect 2487 6647 2491 6651
rect 2428 6626 2431 6636
rect 2495 6626 2498 6679
rect 2508 6651 2511 6664
rect 2524 6657 2527 6666
rect 2545 6657 2548 6666
rect 2531 6626 2534 6636
rect 2545 6619 2548 6651
rect 2402 6561 2408 6599
rect 2402 6491 2408 6557
rect 2413 6562 2416 6592
rect 2413 6528 2416 6558
rect 2430 6541 2433 6551
rect 2413 6513 2416 6524
rect 2429 6515 2432 6524
rect 2450 6509 2453 6522
rect 2466 6515 2469 6524
rect 2475 6513 2478 6518
rect 2481 6498 2484 6551
rect 2493 6537 2494 6541
rect 2532 6539 2535 6551
rect 2487 6515 2490 6524
rect 2487 6505 2491 6509
rect 2402 6429 2408 6487
rect 2428 6484 2431 6494
rect 2495 6484 2498 6537
rect 2545 6528 2548 6565
rect 2508 6509 2511 6522
rect 2524 6515 2527 6524
rect 2545 6515 2548 6524
rect 2531 6484 2534 6494
rect 2402 6297 2408 6425
rect 2402 6165 2408 6293
rect 2402 6091 2408 6161
rect 2402 6033 2408 6087
rect 2529 6067 2533 6072
rect 2553 6067 2557 6800
rect 2562 6769 2565 6779
rect 2561 6743 2564 6752
rect 2582 6737 2585 6750
rect 2598 6743 2601 6752
rect 2607 6741 2610 6746
rect 2613 6726 2616 6779
rect 2625 6765 2626 6769
rect 2664 6767 2667 6779
rect 2619 6743 2622 6752
rect 2619 6733 2623 6737
rect 2560 6712 2563 6722
rect 2627 6712 2630 6765
rect 2640 6737 2643 6750
rect 2656 6743 2659 6752
rect 2663 6712 2666 6722
rect 2562 6683 2565 6693
rect 2561 6657 2564 6666
rect 2582 6651 2585 6664
rect 2598 6657 2601 6666
rect 2607 6655 2610 6660
rect 2613 6640 2616 6693
rect 2625 6679 2626 6683
rect 2664 6681 2667 6693
rect 2619 6657 2622 6666
rect 2619 6647 2623 6651
rect 2560 6626 2563 6636
rect 2627 6626 2630 6679
rect 2640 6651 2643 6664
rect 2656 6657 2659 6666
rect 2663 6626 2666 6636
rect 2670 6612 2674 6933
rect 2694 6909 2697 6919
rect 2677 6883 2680 6892
rect 2693 6883 2696 6892
rect 2714 6877 2717 6890
rect 2730 6883 2733 6892
rect 2739 6881 2742 6886
rect 2677 6845 2680 6877
rect 2745 6866 2748 6919
rect 2757 6905 2758 6909
rect 2796 6907 2799 6919
rect 2751 6883 2754 6892
rect 2751 6873 2755 6877
rect 2692 6852 2695 6862
rect 2759 6852 2762 6905
rect 2772 6877 2775 6890
rect 2788 6883 2791 6892
rect 2795 6852 2798 6862
rect 2677 6756 2680 6793
rect 2802 6790 2805 6882
rect 2694 6769 2697 6779
rect 2677 6743 2680 6752
rect 2693 6743 2696 6752
rect 2714 6737 2717 6750
rect 2730 6743 2733 6752
rect 2739 6741 2742 6746
rect 2745 6726 2748 6779
rect 2757 6765 2758 6769
rect 2796 6767 2799 6779
rect 2751 6743 2754 6752
rect 2751 6733 2755 6737
rect 2692 6712 2695 6722
rect 2759 6712 2762 6765
rect 2772 6737 2775 6750
rect 2788 6743 2791 6752
rect 2795 6712 2798 6722
rect 2802 6704 2805 6742
rect 2694 6683 2697 6693
rect 2677 6657 2680 6666
rect 2693 6657 2696 6666
rect 2714 6651 2717 6664
rect 2730 6657 2733 6666
rect 2739 6655 2742 6660
rect 2677 6619 2680 6651
rect 2745 6640 2748 6693
rect 2757 6679 2758 6683
rect 2796 6681 2799 6693
rect 2751 6657 2754 6666
rect 2751 6647 2755 6651
rect 2692 6626 2695 6636
rect 2759 6626 2762 6679
rect 2772 6651 2775 6664
rect 2788 6657 2791 6666
rect 2795 6626 2798 6636
rect 2654 6608 2658 6612
rect 2670 6607 2674 6608
rect 2654 6589 2658 6604
rect 2654 6580 2658 6585
rect 2654 6572 2658 6576
rect 2670 6576 2674 6592
rect 2686 6589 2690 6604
rect 2686 6580 2690 6585
rect 2562 6541 2565 6551
rect 2561 6515 2564 6524
rect 2582 6509 2585 6522
rect 2598 6515 2601 6524
rect 2607 6513 2610 6518
rect 2613 6498 2616 6551
rect 2625 6537 2626 6541
rect 2664 6539 2667 6551
rect 2619 6515 2622 6524
rect 2619 6505 2623 6509
rect 2560 6484 2563 6494
rect 2627 6484 2630 6537
rect 2640 6509 2643 6522
rect 2656 6515 2659 6524
rect 2663 6484 2666 6494
rect 2560 6139 2563 6151
rect 2601 6137 2602 6141
rect 2568 6115 2571 6124
rect 2584 6109 2587 6122
rect 2561 6084 2564 6094
rect 2597 6084 2600 6137
rect 2605 6115 2608 6124
rect 2604 6105 2608 6109
rect 2611 6098 2614 6151
rect 2662 6141 2665 6151
rect 2617 6113 2620 6118
rect 2626 6115 2629 6124
rect 2642 6109 2645 6122
rect 2663 6115 2666 6124
rect 2664 6084 2667 6094
rect 2402 5989 2408 6029
rect 2545 6026 2548 6056
rect 2545 6019 2548 6022
rect 2545 6013 2548 6015
rect 2402 5956 2408 5985
rect 2402 5877 2408 5952
rect 2430 5927 2433 5937
rect 2413 5907 2416 5910
rect 2402 5737 2408 5873
rect 2413 5899 2416 5903
rect 2429 5901 2432 5910
rect 2450 5895 2453 5908
rect 2466 5901 2469 5910
rect 2475 5899 2478 5904
rect 2413 5848 2416 5895
rect 2481 5884 2484 5937
rect 2493 5923 2494 5927
rect 2532 5925 2535 5937
rect 2487 5901 2490 5910
rect 2487 5891 2491 5895
rect 2428 5870 2431 5880
rect 2495 5870 2498 5923
rect 2508 5895 2511 5908
rect 2524 5901 2527 5910
rect 2545 5901 2548 5910
rect 2531 5870 2534 5880
rect 2545 5863 2548 5895
rect 2553 5856 2557 6063
rect 2670 6076 2674 6572
rect 2677 6528 2680 6565
rect 2802 6562 2805 6656
rect 2694 6541 2697 6551
rect 2677 6515 2680 6524
rect 2693 6515 2696 6524
rect 2714 6509 2717 6522
rect 2730 6515 2733 6524
rect 2739 6513 2742 6518
rect 2745 6498 2748 6551
rect 2757 6537 2758 6541
rect 2796 6539 2799 6551
rect 2751 6515 2754 6524
rect 2751 6505 2755 6509
rect 2692 6484 2695 6494
rect 2759 6484 2762 6537
rect 2772 6509 2775 6522
rect 2788 6515 2791 6524
rect 2795 6484 2798 6494
rect 2679 6115 2682 6124
rect 2562 6039 2565 6049
rect 2561 6013 2564 6022
rect 2582 6007 2585 6020
rect 2598 6013 2601 6022
rect 2607 6011 2610 6016
rect 2613 5996 2616 6049
rect 2625 6035 2626 6039
rect 2664 6037 2667 6049
rect 2619 6013 2622 6022
rect 2619 6003 2623 6007
rect 2560 5982 2563 5992
rect 2627 5982 2630 6035
rect 2640 6007 2643 6020
rect 2656 6013 2659 6022
rect 2663 5982 2666 5992
rect 2562 5927 2565 5937
rect 2561 5901 2564 5910
rect 2582 5895 2585 5908
rect 2598 5901 2601 5910
rect 2607 5899 2610 5904
rect 2613 5884 2616 5937
rect 2625 5923 2626 5927
rect 2664 5925 2667 5937
rect 2619 5901 2622 5910
rect 2619 5891 2623 5895
rect 2560 5870 2563 5880
rect 2627 5870 2630 5923
rect 2640 5895 2643 5908
rect 2656 5901 2659 5910
rect 2663 5870 2666 5880
rect 2537 5852 2541 5856
rect 2553 5851 2557 5852
rect 2413 5808 2416 5836
rect 2537 5833 2541 5848
rect 2537 5826 2541 5829
rect 2537 5818 2541 5822
rect 2553 5822 2557 5836
rect 2569 5833 2573 5848
rect 2569 5826 2573 5829
rect 2413 5774 2416 5804
rect 2430 5787 2433 5797
rect 2413 5759 2416 5770
rect 2429 5761 2432 5770
rect 2450 5755 2453 5768
rect 2466 5761 2469 5770
rect 2475 5759 2478 5764
rect 2481 5744 2484 5797
rect 2493 5783 2494 5787
rect 2532 5785 2535 5797
rect 2487 5761 2490 5770
rect 2487 5751 2491 5755
rect 2402 5651 2408 5733
rect 2428 5730 2431 5740
rect 2495 5730 2498 5783
rect 2545 5774 2548 5811
rect 2508 5755 2511 5768
rect 2524 5761 2527 5770
rect 2545 5761 2548 5770
rect 2531 5730 2534 5740
rect 2402 5621 2408 5647
rect 2413 5688 2416 5718
rect 2430 5701 2433 5711
rect 2413 5673 2416 5684
rect 2429 5675 2432 5684
rect 2450 5669 2453 5682
rect 2466 5675 2469 5684
rect 2475 5673 2478 5678
rect 2413 5622 2416 5669
rect 2481 5658 2484 5711
rect 2493 5697 2494 5701
rect 2532 5699 2535 5711
rect 2487 5675 2490 5684
rect 2487 5665 2491 5669
rect 2428 5644 2431 5654
rect 2495 5644 2498 5697
rect 2508 5669 2511 5682
rect 2524 5675 2527 5684
rect 2545 5675 2548 5684
rect 2531 5644 2534 5654
rect 2545 5637 2548 5669
rect 2402 5579 2408 5617
rect 2402 5509 2408 5575
rect 2413 5580 2416 5610
rect 2413 5546 2416 5576
rect 2430 5559 2433 5569
rect 2413 5531 2416 5542
rect 2429 5533 2432 5542
rect 2450 5527 2453 5540
rect 2466 5533 2469 5542
rect 2475 5531 2478 5536
rect 2481 5516 2484 5569
rect 2493 5555 2494 5559
rect 2532 5557 2535 5569
rect 2487 5533 2490 5542
rect 2487 5523 2491 5527
rect 2402 5447 2408 5505
rect 2428 5502 2431 5512
rect 2495 5502 2498 5555
rect 2545 5546 2548 5583
rect 2508 5527 2511 5540
rect 2524 5533 2527 5542
rect 2545 5533 2548 5542
rect 2531 5502 2534 5512
rect 2402 5315 2408 5443
rect 2402 5183 2408 5311
rect 2402 5109 2408 5179
rect 2402 5051 2408 5105
rect 2529 5085 2533 5090
rect 2553 5085 2557 5818
rect 2562 5787 2565 5797
rect 2561 5761 2564 5770
rect 2582 5755 2585 5768
rect 2598 5761 2601 5770
rect 2607 5759 2610 5764
rect 2613 5744 2616 5797
rect 2625 5783 2626 5787
rect 2664 5785 2667 5797
rect 2619 5761 2622 5770
rect 2619 5751 2623 5755
rect 2560 5730 2563 5740
rect 2627 5730 2630 5783
rect 2640 5755 2643 5768
rect 2656 5761 2659 5770
rect 2663 5730 2666 5740
rect 2562 5701 2565 5711
rect 2561 5675 2564 5684
rect 2582 5669 2585 5682
rect 2598 5675 2601 5684
rect 2607 5673 2610 5678
rect 2613 5658 2616 5711
rect 2625 5697 2626 5701
rect 2664 5699 2667 5711
rect 2619 5675 2622 5684
rect 2619 5665 2623 5669
rect 2560 5644 2563 5654
rect 2627 5644 2630 5697
rect 2640 5669 2643 5682
rect 2656 5675 2659 5684
rect 2663 5644 2666 5654
rect 2670 5630 2674 6072
rect 2679 6069 2682 6109
rect 2679 6016 2682 6065
rect 2694 5927 2697 5937
rect 2677 5901 2680 5910
rect 2693 5901 2696 5910
rect 2714 5895 2717 5908
rect 2730 5901 2733 5910
rect 2739 5899 2742 5904
rect 2677 5863 2680 5895
rect 2745 5884 2748 5937
rect 2757 5923 2758 5927
rect 2796 5925 2799 5937
rect 2751 5901 2754 5910
rect 2751 5891 2755 5895
rect 2692 5870 2695 5880
rect 2759 5870 2762 5923
rect 2772 5895 2775 5908
rect 2788 5901 2791 5910
rect 2795 5870 2798 5880
rect 2677 5774 2680 5811
rect 2802 5808 2805 5900
rect 2694 5787 2697 5797
rect 2677 5761 2680 5770
rect 2693 5761 2696 5770
rect 2714 5755 2717 5768
rect 2730 5761 2733 5770
rect 2739 5759 2742 5764
rect 2745 5744 2748 5797
rect 2757 5783 2758 5787
rect 2796 5785 2799 5797
rect 2751 5761 2754 5770
rect 2751 5751 2755 5755
rect 2692 5730 2695 5740
rect 2759 5730 2762 5783
rect 2772 5755 2775 5768
rect 2788 5761 2791 5770
rect 2795 5730 2798 5740
rect 2802 5722 2805 5760
rect 2694 5701 2697 5711
rect 2677 5675 2680 5684
rect 2693 5675 2696 5684
rect 2714 5669 2717 5682
rect 2730 5675 2733 5684
rect 2739 5673 2742 5678
rect 2677 5637 2680 5669
rect 2745 5658 2748 5711
rect 2757 5697 2758 5701
rect 2796 5699 2799 5711
rect 2751 5675 2754 5684
rect 2751 5665 2755 5669
rect 2692 5644 2695 5654
rect 2759 5644 2762 5697
rect 2772 5669 2775 5682
rect 2788 5675 2791 5684
rect 2795 5644 2798 5654
rect 2654 5626 2658 5630
rect 2670 5625 2674 5626
rect 2654 5607 2658 5622
rect 2654 5599 2658 5603
rect 2654 5590 2658 5595
rect 2670 5594 2674 5610
rect 2686 5607 2690 5622
rect 2686 5599 2690 5603
rect 2562 5559 2565 5569
rect 2561 5533 2564 5542
rect 2582 5527 2585 5540
rect 2598 5533 2601 5542
rect 2607 5531 2610 5536
rect 2613 5516 2616 5569
rect 2625 5555 2626 5559
rect 2664 5557 2667 5569
rect 2619 5533 2622 5542
rect 2619 5523 2623 5527
rect 2560 5502 2563 5512
rect 2627 5502 2630 5555
rect 2640 5527 2643 5540
rect 2656 5533 2659 5542
rect 2663 5502 2666 5512
rect 2560 5157 2563 5169
rect 2601 5155 2602 5159
rect 2568 5133 2571 5142
rect 2584 5127 2587 5140
rect 2561 5102 2564 5112
rect 2597 5102 2600 5155
rect 2605 5133 2608 5142
rect 2604 5123 2608 5127
rect 2611 5116 2614 5169
rect 2662 5159 2665 5169
rect 2617 5131 2620 5136
rect 2626 5133 2629 5142
rect 2642 5127 2645 5140
rect 2663 5133 2666 5142
rect 2664 5102 2667 5112
rect 2402 5007 2408 5047
rect 2545 5044 2548 5074
rect 2545 5037 2548 5040
rect 2545 5031 2548 5033
rect 2402 4974 2408 5003
rect 2402 4855 2408 4970
rect 2553 4947 2557 5081
rect 2670 5094 2674 5590
rect 2677 5546 2680 5583
rect 2802 5580 2805 5674
rect 2694 5559 2697 5569
rect 2677 5533 2680 5542
rect 2693 5533 2696 5542
rect 2714 5527 2717 5540
rect 2730 5533 2733 5542
rect 2739 5531 2742 5536
rect 2745 5516 2748 5569
rect 2757 5555 2758 5559
rect 2796 5557 2799 5569
rect 2751 5533 2754 5542
rect 2751 5523 2755 5527
rect 2692 5502 2695 5512
rect 2759 5502 2762 5555
rect 2772 5527 2775 5540
rect 2788 5533 2791 5542
rect 2795 5502 2798 5512
rect 2679 5133 2682 5142
rect 2562 5057 2565 5067
rect 2561 5031 2564 5040
rect 2582 5025 2585 5038
rect 2598 5031 2601 5040
rect 2607 5029 2610 5034
rect 2613 5014 2616 5067
rect 2625 5053 2626 5057
rect 2664 5055 2667 5067
rect 2619 5031 2622 5040
rect 2619 5021 2623 5025
rect 2560 5000 2563 5010
rect 2627 5000 2630 5053
rect 2640 5025 2643 5038
rect 2656 5031 2659 5040
rect 2663 5000 2666 5010
rect 2670 4936 2674 5090
rect 2679 5087 2682 5127
rect 2679 5034 2682 5083
rect 3836 4936 3844 7464
rect 3918 7366 3922 7472
rect 4493 7475 4641 7477
rect 4493 7471 4496 7475
rect 4500 7471 4501 7475
rect 4505 7473 4641 7475
rect 4505 7471 4645 7473
rect 4493 7470 4645 7471
rect 4493 7466 4496 7470
rect 4500 7466 4501 7470
rect 4505 7466 4641 7470
rect 4493 7465 4645 7466
rect 4493 7461 4496 7465
rect 4500 7461 4501 7465
rect 4505 7461 4641 7465
rect 4493 7460 4645 7461
rect 4493 7456 4496 7460
rect 4500 7456 4501 7460
rect 4505 7456 4641 7460
rect 4493 7455 4645 7456
rect 4493 7451 4496 7455
rect 4500 7451 4501 7455
rect 4505 7451 4641 7455
rect 4493 7450 4645 7451
rect 4493 7446 4496 7450
rect 4500 7446 4501 7450
rect 4505 7446 4641 7450
rect 4493 7445 4645 7446
rect 4493 7441 4496 7445
rect 4500 7441 4501 7445
rect 4505 7441 4641 7445
rect 4493 7440 4645 7441
rect 4493 7436 4496 7440
rect 4500 7436 4501 7440
rect 4505 7436 4641 7440
rect 4493 7435 4645 7436
rect 4493 7431 4496 7435
rect 4500 7431 4501 7435
rect 4505 7431 4641 7435
rect 4493 7430 4645 7431
rect 4493 7426 4496 7430
rect 4500 7426 4501 7430
rect 4505 7426 4641 7430
rect 4493 7425 4645 7426
rect 4493 7421 4496 7425
rect 4500 7421 4501 7425
rect 4505 7421 4641 7425
rect 4493 7420 4645 7421
rect 4493 7416 4496 7420
rect 4500 7416 4501 7420
rect 4505 7416 4641 7420
rect 4493 7415 4645 7416
rect 4493 7411 4496 7415
rect 4500 7411 4501 7415
rect 4505 7413 4645 7415
rect 4505 7411 4641 7413
rect 4493 7409 4641 7411
rect 4657 7461 4662 7465
rect 4666 7461 4672 7465
rect 4676 7461 4682 7465
rect 4686 7461 4692 7465
rect 4696 7461 4702 7465
rect 4706 7461 4712 7465
rect 4716 7461 4722 7465
rect 4726 7461 4732 7465
rect 4736 7461 4742 7465
rect 4657 7460 4746 7461
rect 4661 7456 4667 7460
rect 4671 7456 4677 7460
rect 4681 7456 4687 7460
rect 4691 7456 4697 7460
rect 4701 7456 4707 7460
rect 4711 7456 4717 7460
rect 4721 7456 4727 7460
rect 4731 7456 4737 7460
rect 4741 7456 4746 7460
rect 4657 7455 4746 7456
rect 4657 7451 4662 7455
rect 4666 7451 4672 7455
rect 4676 7451 4682 7455
rect 4686 7451 4692 7455
rect 4696 7451 4702 7455
rect 4706 7451 4712 7455
rect 4716 7451 4722 7455
rect 4726 7451 4732 7455
rect 4736 7451 4742 7455
rect 4657 7450 4746 7451
rect 4661 7446 4667 7450
rect 4671 7446 4677 7450
rect 4681 7446 4687 7450
rect 4691 7446 4697 7450
rect 4701 7446 4707 7450
rect 4711 7446 4717 7450
rect 4721 7446 4727 7450
rect 4731 7446 4737 7450
rect 4741 7446 4746 7450
rect 4657 7445 4746 7446
rect 4657 7441 4662 7445
rect 4666 7441 4672 7445
rect 4676 7441 4682 7445
rect 4686 7441 4692 7445
rect 4696 7441 4702 7445
rect 4706 7441 4712 7445
rect 4716 7441 4722 7445
rect 4726 7441 4732 7445
rect 4736 7441 4742 7445
rect 4657 7440 4746 7441
rect 4661 7436 4667 7440
rect 4671 7436 4677 7440
rect 4681 7436 4687 7440
rect 4691 7436 4697 7440
rect 4701 7436 4707 7440
rect 4711 7436 4717 7440
rect 4721 7436 4727 7440
rect 4731 7436 4737 7440
rect 4741 7436 4746 7440
rect 4657 7435 4746 7436
rect 4657 7431 4662 7435
rect 4666 7431 4672 7435
rect 4676 7431 4682 7435
rect 4686 7431 4692 7435
rect 4696 7431 4702 7435
rect 4706 7431 4712 7435
rect 4716 7431 4722 7435
rect 4726 7431 4732 7435
rect 4736 7431 4742 7435
rect 4657 7430 4746 7431
rect 4661 7426 4667 7430
rect 4671 7426 4677 7430
rect 4681 7426 4687 7430
rect 4691 7426 4697 7430
rect 4701 7426 4707 7430
rect 4711 7426 4717 7430
rect 4721 7426 4727 7430
rect 4731 7426 4737 7430
rect 4741 7426 4746 7430
rect 4657 7425 4746 7426
rect 4657 7421 4662 7425
rect 4666 7421 4672 7425
rect 4676 7421 4682 7425
rect 4686 7421 4692 7425
rect 4696 7421 4702 7425
rect 4706 7421 4712 7425
rect 4716 7421 4722 7425
rect 4726 7421 4732 7425
rect 4736 7421 4742 7425
rect 4657 7411 4746 7421
rect 4786 7411 4795 7421
rect 4657 7408 4795 7411
rect 4657 7404 4775 7408
rect 4779 7404 4780 7408
rect 4784 7404 4785 7408
rect 4789 7404 4790 7408
rect 4794 7404 4795 7408
rect 4657 7401 4795 7404
rect 4657 7397 4775 7401
rect 4779 7397 4780 7401
rect 4784 7397 4785 7401
rect 4789 7397 4790 7401
rect 4794 7397 4795 7401
rect 4657 7394 4795 7397
rect 4576 7389 4588 7393
rect 4592 7389 4604 7393
rect 4608 7389 4620 7393
rect 4657 7390 4775 7394
rect 4779 7390 4780 7394
rect 4784 7390 4785 7394
rect 4789 7390 4790 7394
rect 4794 7390 4795 7394
rect 4657 7387 4795 7390
rect 4657 7383 4775 7387
rect 4779 7383 4780 7387
rect 4784 7383 4785 7387
rect 4789 7383 4790 7387
rect 4794 7383 4795 7387
rect 4657 7380 4795 7383
rect 4657 7376 4775 7380
rect 4779 7376 4780 7380
rect 4784 7376 4785 7380
rect 4789 7376 4790 7380
rect 4794 7376 4795 7380
rect 4657 7373 4795 7376
rect 4657 7369 4775 7373
rect 4779 7369 4780 7373
rect 4784 7369 4785 7373
rect 4789 7369 4790 7373
rect 4794 7369 4795 7373
rect 4657 7366 4795 7369
rect 4657 7362 4775 7366
rect 4779 7362 4780 7366
rect 4784 7362 4785 7366
rect 4789 7362 4790 7366
rect 4794 7362 4795 7366
rect 4657 7359 4795 7362
rect 4657 7355 4775 7359
rect 4779 7355 4780 7359
rect 4784 7355 4785 7359
rect 4789 7355 4790 7359
rect 4794 7355 4795 7359
rect 4657 7352 4795 7355
rect 4657 7348 4775 7352
rect 4779 7348 4780 7352
rect 4784 7348 4785 7352
rect 4789 7348 4790 7352
rect 4794 7348 4795 7352
rect 4657 7345 4795 7348
rect 4657 7341 4775 7345
rect 4779 7341 4780 7345
rect 4784 7341 4785 7345
rect 4789 7341 4790 7345
rect 4794 7341 4795 7345
rect 4657 7338 4795 7341
rect 4576 7331 4588 7335
rect 4592 7331 4604 7335
rect 4608 7331 4620 7335
rect 4657 7334 4775 7338
rect 4779 7334 4780 7338
rect 4784 7334 4785 7338
rect 4789 7334 4790 7338
rect 4794 7334 4795 7338
rect 4657 7331 4795 7334
rect 4657 7327 4775 7331
rect 4779 7327 4780 7331
rect 4784 7327 4785 7331
rect 4789 7327 4790 7331
rect 4794 7327 4795 7331
rect 4657 7324 4795 7327
rect 4657 7320 4775 7324
rect 4779 7320 4780 7324
rect 4784 7320 4785 7324
rect 4789 7320 4790 7324
rect 4794 7320 4795 7324
rect 4550 7315 4641 7317
rect 4550 7311 4553 7315
rect 4557 7311 4558 7315
rect 4562 7313 4641 7315
rect 4562 7311 4645 7313
rect 4550 7310 4645 7311
rect 4550 7306 4553 7310
rect 4557 7306 4558 7310
rect 4562 7306 4641 7310
rect 4550 7305 4645 7306
rect 4550 7301 4553 7305
rect 4557 7301 4558 7305
rect 4562 7301 4641 7305
rect 4550 7300 4645 7301
rect 4550 7296 4553 7300
rect 4557 7296 4558 7300
rect 4562 7296 4641 7300
rect 4550 7295 4645 7296
rect 4494 7289 4496 7293
rect 4500 7289 4501 7293
rect 4505 7289 4506 7293
rect 4510 7289 4511 7293
rect 4494 7288 4515 7289
rect 4494 7284 4496 7288
rect 4500 7284 4501 7288
rect 4505 7284 4506 7288
rect 4510 7284 4511 7288
rect 4494 7283 4515 7284
rect 4494 7279 4496 7283
rect 4500 7279 4501 7283
rect 4505 7279 4506 7283
rect 4510 7279 4511 7283
rect 4494 7278 4515 7279
rect 4494 7274 4496 7278
rect 4500 7274 4501 7278
rect 4505 7274 4506 7278
rect 4510 7274 4511 7278
rect 4494 7273 4515 7274
rect 4494 7269 4496 7273
rect 4500 7269 4501 7273
rect 4505 7269 4506 7273
rect 4510 7269 4511 7273
rect 4494 7268 4515 7269
rect 4494 7264 4496 7268
rect 4500 7264 4501 7268
rect 4505 7264 4506 7268
rect 4510 7264 4511 7268
rect 4494 7263 4515 7264
rect 4494 7259 4496 7263
rect 4500 7259 4501 7263
rect 4505 7259 4506 7263
rect 4510 7259 4511 7263
rect 4494 7258 4515 7259
rect 4494 7254 4496 7258
rect 4500 7254 4501 7258
rect 4505 7254 4506 7258
rect 4510 7254 4511 7258
rect 4494 7253 4515 7254
rect 4494 7249 4496 7253
rect 4500 7249 4501 7253
rect 4505 7249 4506 7253
rect 4510 7249 4511 7253
rect 4550 7291 4553 7295
rect 4557 7291 4558 7295
rect 4562 7291 4641 7295
rect 4550 7290 4645 7291
rect 4550 7286 4553 7290
rect 4557 7286 4558 7290
rect 4562 7286 4641 7290
rect 4550 7285 4645 7286
rect 4550 7281 4553 7285
rect 4557 7281 4558 7285
rect 4562 7281 4641 7285
rect 4550 7280 4645 7281
rect 4550 7276 4553 7280
rect 4557 7276 4558 7280
rect 4562 7276 4641 7280
rect 4550 7275 4645 7276
rect 4550 7271 4553 7275
rect 4557 7271 4558 7275
rect 4562 7271 4641 7275
rect 4550 7270 4645 7271
rect 4550 7266 4553 7270
rect 4557 7266 4558 7270
rect 4562 7266 4641 7270
rect 4550 7265 4645 7266
rect 4550 7261 4553 7265
rect 4557 7261 4558 7265
rect 4562 7261 4641 7265
rect 4657 7315 4795 7320
rect 4657 7305 4746 7315
rect 4786 7305 4795 7315
rect 4657 7301 4662 7305
rect 4666 7301 4672 7305
rect 4676 7301 4682 7305
rect 4686 7301 4692 7305
rect 4696 7301 4702 7305
rect 4706 7301 4712 7305
rect 4716 7301 4722 7305
rect 4726 7301 4732 7305
rect 4736 7301 4742 7305
rect 4657 7300 4746 7301
rect 4661 7296 4667 7300
rect 4671 7296 4677 7300
rect 4681 7296 4687 7300
rect 4691 7296 4697 7300
rect 4701 7296 4707 7300
rect 4711 7296 4717 7300
rect 4721 7296 4727 7300
rect 4731 7296 4737 7300
rect 4741 7296 4746 7300
rect 4657 7295 4746 7296
rect 4657 7291 4662 7295
rect 4666 7291 4672 7295
rect 4676 7291 4682 7295
rect 4686 7291 4692 7295
rect 4696 7291 4702 7295
rect 4706 7291 4712 7295
rect 4716 7291 4722 7295
rect 4726 7291 4732 7295
rect 4736 7291 4742 7295
rect 4657 7290 4746 7291
rect 4661 7286 4667 7290
rect 4671 7286 4677 7290
rect 4681 7286 4687 7290
rect 4691 7286 4697 7290
rect 4701 7286 4707 7290
rect 4711 7286 4717 7290
rect 4721 7286 4727 7290
rect 4731 7286 4737 7290
rect 4741 7286 4746 7290
rect 4657 7285 4746 7286
rect 4657 7281 4662 7285
rect 4666 7281 4672 7285
rect 4676 7281 4682 7285
rect 4686 7281 4692 7285
rect 4696 7281 4702 7285
rect 4706 7281 4712 7285
rect 4716 7281 4722 7285
rect 4726 7281 4732 7285
rect 4736 7281 4742 7285
rect 4657 7280 4746 7281
rect 4661 7276 4667 7280
rect 4671 7276 4677 7280
rect 4681 7276 4687 7280
rect 4691 7276 4697 7280
rect 4701 7276 4707 7280
rect 4711 7276 4717 7280
rect 4721 7276 4727 7280
rect 4731 7276 4737 7280
rect 4741 7276 4746 7280
rect 4657 7275 4746 7276
rect 4657 7271 4662 7275
rect 4666 7271 4672 7275
rect 4676 7271 4682 7275
rect 4686 7271 4692 7275
rect 4696 7271 4702 7275
rect 4706 7271 4712 7275
rect 4716 7271 4722 7275
rect 4726 7271 4732 7275
rect 4736 7271 4742 7275
rect 4657 7270 4746 7271
rect 4661 7266 4667 7270
rect 4671 7266 4677 7270
rect 4681 7266 4687 7270
rect 4691 7266 4697 7270
rect 4701 7266 4707 7270
rect 4711 7266 4717 7270
rect 4721 7266 4727 7270
rect 4731 7266 4737 7270
rect 4741 7266 4746 7270
rect 4657 7265 4746 7266
rect 4657 7261 4662 7265
rect 4666 7261 4672 7265
rect 4676 7261 4682 7265
rect 4686 7261 4692 7265
rect 4696 7261 4702 7265
rect 4706 7261 4712 7265
rect 4716 7261 4722 7265
rect 4726 7261 4732 7265
rect 4736 7261 4742 7265
rect 4550 7260 4645 7261
rect 4550 7256 4553 7260
rect 4557 7256 4558 7260
rect 4562 7256 4641 7260
rect 4550 7255 4645 7256
rect 4550 7251 4553 7255
rect 4557 7251 4558 7255
rect 4562 7253 4645 7255
rect 4562 7251 4641 7253
rect 4550 7249 4641 7251
rect 4494 7248 4515 7249
rect 4494 7244 4496 7248
rect 4500 7244 4501 7248
rect 4505 7244 4506 7248
rect 4510 7244 4511 7248
rect 4494 7243 4515 7244
rect 4494 7239 4496 7243
rect 4500 7239 4501 7243
rect 4505 7239 4506 7243
rect 4510 7239 4511 7243
rect 4494 7237 4515 7239
rect 4826 7236 4829 7490
rect 5083 7236 5086 7490
rect 4483 7230 4484 7234
rect 4488 7230 4489 7234
rect 4493 7230 4494 7234
rect 4498 7230 4499 7234
rect 4503 7230 4504 7234
rect 4508 7230 4509 7234
rect 4479 7229 4513 7230
rect 4483 7225 4484 7229
rect 4488 7225 4489 7229
rect 4493 7225 4494 7229
rect 4498 7225 4499 7229
rect 4503 7225 4504 7229
rect 4508 7225 4509 7229
rect 4479 7224 4513 7225
rect 4483 7220 4484 7224
rect 4488 7220 4489 7224
rect 4493 7220 4494 7224
rect 4498 7220 4499 7224
rect 4503 7220 4504 7224
rect 4508 7220 4509 7224
rect 4479 7219 4513 7220
rect 4483 7215 4484 7219
rect 4488 7215 4489 7219
rect 4493 7215 4494 7219
rect 4498 7215 4499 7219
rect 4503 7215 4504 7219
rect 4508 7215 4509 7219
rect 4529 7230 4530 7234
rect 4534 7230 4535 7234
rect 4539 7230 4540 7234
rect 4544 7230 4545 7234
rect 4549 7230 4550 7234
rect 4554 7230 4555 7234
rect 4826 7233 5086 7236
rect 4525 7229 4559 7230
rect 4529 7225 4530 7229
rect 4534 7225 4535 7229
rect 4539 7225 4540 7229
rect 4544 7225 4545 7229
rect 4549 7225 4550 7229
rect 4554 7225 4555 7229
rect 4525 7224 4559 7225
rect 4529 7220 4530 7224
rect 4534 7220 4535 7224
rect 4539 7220 4540 7224
rect 4544 7220 4545 7224
rect 4549 7220 4550 7224
rect 4554 7220 4555 7224
rect 4525 7219 4559 7220
rect 4529 7215 4530 7219
rect 4534 7215 4535 7219
rect 4539 7215 4540 7219
rect 4544 7215 4545 7219
rect 4549 7215 4550 7219
rect 4554 7215 4555 7219
rect 4483 7202 4484 7206
rect 4488 7202 4489 7206
rect 4493 7202 4494 7206
rect 4498 7202 4499 7206
rect 4503 7202 4504 7206
rect 4508 7202 4509 7206
rect 4479 7201 4513 7202
rect 4483 7197 4484 7201
rect 4488 7197 4489 7201
rect 4493 7197 4494 7201
rect 4498 7197 4499 7201
rect 4503 7197 4504 7201
rect 4508 7197 4509 7201
rect 4479 7196 4513 7197
rect 4483 7192 4484 7196
rect 4488 7192 4489 7196
rect 4493 7192 4494 7196
rect 4498 7192 4499 7196
rect 4503 7192 4504 7196
rect 4508 7192 4509 7196
rect 4479 7191 4513 7192
rect 4483 7187 4484 7191
rect 4488 7187 4489 7191
rect 4493 7187 4494 7191
rect 4498 7187 4499 7191
rect 4503 7187 4504 7191
rect 4508 7187 4509 7191
rect 4529 7202 4530 7206
rect 4534 7202 4535 7206
rect 4539 7202 4540 7206
rect 4544 7202 4545 7206
rect 4549 7202 4550 7206
rect 4554 7202 4555 7206
rect 4525 7201 4559 7202
rect 4529 7197 4530 7201
rect 4534 7197 4535 7201
rect 4539 7197 4540 7201
rect 4544 7197 4545 7201
rect 4549 7197 4550 7201
rect 4554 7197 4555 7201
rect 4525 7196 4559 7197
rect 4529 7192 4530 7196
rect 4534 7192 4535 7196
rect 4539 7192 4540 7196
rect 4544 7192 4545 7196
rect 4549 7192 4550 7196
rect 4554 7192 4555 7196
rect 4525 7191 4559 7192
rect 4529 7187 4530 7191
rect 4534 7187 4535 7191
rect 4539 7187 4540 7191
rect 4544 7187 4545 7191
rect 4549 7187 4550 7191
rect 4554 7187 4555 7191
rect 4479 7156 4513 7157
rect 4483 7152 4484 7156
rect 4488 7152 4489 7156
rect 4493 7152 4494 7156
rect 4498 7152 4499 7156
rect 4503 7152 4504 7156
rect 4508 7152 4509 7156
rect 4525 7156 4559 7157
rect 4529 7152 4530 7156
rect 4534 7152 4535 7156
rect 4539 7152 4540 7156
rect 4544 7152 4545 7156
rect 4549 7152 4550 7156
rect 4554 7152 4555 7156
rect 4826 7118 5086 7121
rect 4826 6864 4829 7118
rect 5083 6864 5086 7118
rect 4483 6858 4484 6862
rect 4488 6858 4489 6862
rect 4493 6858 4494 6862
rect 4498 6858 4499 6862
rect 4503 6858 4504 6862
rect 4508 6858 4509 6862
rect 4479 6857 4513 6858
rect 4483 6853 4484 6857
rect 4488 6853 4489 6857
rect 4493 6853 4494 6857
rect 4498 6853 4499 6857
rect 4503 6853 4504 6857
rect 4508 6853 4509 6857
rect 4479 6852 4513 6853
rect 4483 6848 4484 6852
rect 4488 6848 4489 6852
rect 4493 6848 4494 6852
rect 4498 6848 4499 6852
rect 4503 6848 4504 6852
rect 4508 6848 4509 6852
rect 4479 6847 4513 6848
rect 4483 6843 4484 6847
rect 4488 6843 4489 6847
rect 4493 6843 4494 6847
rect 4498 6843 4499 6847
rect 4503 6843 4504 6847
rect 4508 6843 4509 6847
rect 4529 6858 4530 6862
rect 4534 6858 4535 6862
rect 4539 6858 4540 6862
rect 4544 6858 4545 6862
rect 4549 6858 4550 6862
rect 4554 6858 4555 6862
rect 4826 6861 5086 6864
rect 4525 6857 4559 6858
rect 4529 6853 4530 6857
rect 4534 6853 4535 6857
rect 4539 6853 4540 6857
rect 4544 6853 4545 6857
rect 4549 6853 4550 6857
rect 4554 6853 4555 6857
rect 4525 6852 4559 6853
rect 4529 6848 4530 6852
rect 4534 6848 4535 6852
rect 4539 6848 4540 6852
rect 4544 6848 4545 6852
rect 4549 6848 4550 6852
rect 4554 6848 4555 6852
rect 4525 6847 4559 6848
rect 4529 6843 4530 6847
rect 4534 6843 4535 6847
rect 4539 6843 4540 6847
rect 4544 6843 4545 6847
rect 4549 6843 4550 6847
rect 4554 6843 4555 6847
rect 4826 6809 5086 6812
rect 4826 6555 4829 6809
rect 5083 6555 5086 6809
rect 4483 6549 4484 6553
rect 4488 6549 4489 6553
rect 4493 6549 4494 6553
rect 4498 6549 4499 6553
rect 4503 6549 4504 6553
rect 4508 6549 4509 6553
rect 4479 6548 4513 6549
rect 4483 6544 4484 6548
rect 4488 6544 4489 6548
rect 4493 6544 4494 6548
rect 4498 6544 4499 6548
rect 4503 6544 4504 6548
rect 4508 6544 4509 6548
rect 4479 6543 4513 6544
rect 4483 6539 4484 6543
rect 4488 6539 4489 6543
rect 4493 6539 4494 6543
rect 4498 6539 4499 6543
rect 4503 6539 4504 6543
rect 4508 6539 4509 6543
rect 4479 6538 4513 6539
rect 4483 6534 4484 6538
rect 4488 6534 4489 6538
rect 4493 6534 4494 6538
rect 4498 6534 4499 6538
rect 4503 6534 4504 6538
rect 4508 6534 4509 6538
rect 4529 6549 4530 6553
rect 4534 6549 4535 6553
rect 4539 6549 4540 6553
rect 4544 6549 4545 6553
rect 4549 6549 4550 6553
rect 4554 6549 4555 6553
rect 4826 6552 5086 6555
rect 4525 6548 4559 6549
rect 4529 6544 4530 6548
rect 4534 6544 4535 6548
rect 4539 6544 4540 6548
rect 4544 6544 4545 6548
rect 4549 6544 4550 6548
rect 4554 6544 4555 6548
rect 4525 6543 4559 6544
rect 4529 6539 4530 6543
rect 4534 6539 4535 6543
rect 4539 6539 4540 6543
rect 4544 6539 4545 6543
rect 4549 6539 4550 6543
rect 4554 6539 4555 6543
rect 4525 6538 4559 6539
rect 4529 6534 4530 6538
rect 4534 6534 4535 6538
rect 4539 6534 4540 6538
rect 4544 6534 4545 6538
rect 4549 6534 4550 6538
rect 4554 6534 4555 6538
rect 4826 6500 5086 6503
rect 4826 6246 4829 6500
rect 5083 6246 5086 6500
rect 4483 6240 4484 6244
rect 4488 6240 4489 6244
rect 4493 6240 4494 6244
rect 4498 6240 4499 6244
rect 4503 6240 4504 6244
rect 4508 6240 4509 6244
rect 4479 6239 4513 6240
rect 4483 6235 4484 6239
rect 4488 6235 4489 6239
rect 4493 6235 4494 6239
rect 4498 6235 4499 6239
rect 4503 6235 4504 6239
rect 4508 6235 4509 6239
rect 4479 6234 4513 6235
rect 4483 6230 4484 6234
rect 4488 6230 4489 6234
rect 4493 6230 4494 6234
rect 4498 6230 4499 6234
rect 4503 6230 4504 6234
rect 4508 6230 4509 6234
rect 4479 6229 4513 6230
rect 4483 6225 4484 6229
rect 4488 6225 4489 6229
rect 4493 6225 4494 6229
rect 4498 6225 4499 6229
rect 4503 6225 4504 6229
rect 4508 6225 4509 6229
rect 4529 6240 4530 6244
rect 4534 6240 4535 6244
rect 4539 6240 4540 6244
rect 4544 6240 4545 6244
rect 4549 6240 4550 6244
rect 4554 6240 4555 6244
rect 4826 6243 5086 6246
rect 4525 6239 4559 6240
rect 4529 6235 4530 6239
rect 4534 6235 4535 6239
rect 4539 6235 4540 6239
rect 4544 6235 4545 6239
rect 4549 6235 4550 6239
rect 4554 6235 4555 6239
rect 4525 6234 4559 6235
rect 4529 6230 4530 6234
rect 4534 6230 4535 6234
rect 4539 6230 4540 6234
rect 4544 6230 4545 6234
rect 4549 6230 4550 6234
rect 4554 6230 4555 6234
rect 4525 6229 4559 6230
rect 4529 6225 4530 6229
rect 4534 6225 4535 6229
rect 4539 6225 4540 6229
rect 4544 6225 4545 6229
rect 4549 6225 4550 6229
rect 4554 6225 4555 6229
rect 4826 6191 5086 6194
rect 4826 5937 4829 6191
rect 5083 5937 5086 6191
rect 4483 5931 4484 5935
rect 4488 5931 4489 5935
rect 4493 5931 4494 5935
rect 4498 5931 4499 5935
rect 4503 5931 4504 5935
rect 4508 5931 4509 5935
rect 4479 5930 4513 5931
rect 4483 5926 4484 5930
rect 4488 5926 4489 5930
rect 4493 5926 4494 5930
rect 4498 5926 4499 5930
rect 4503 5926 4504 5930
rect 4508 5926 4509 5930
rect 4479 5925 4513 5926
rect 4483 5921 4484 5925
rect 4488 5921 4489 5925
rect 4493 5921 4494 5925
rect 4498 5921 4499 5925
rect 4503 5921 4504 5925
rect 4508 5921 4509 5925
rect 4479 5920 4513 5921
rect 4483 5916 4484 5920
rect 4488 5916 4489 5920
rect 4493 5916 4494 5920
rect 4498 5916 4499 5920
rect 4503 5916 4504 5920
rect 4508 5916 4509 5920
rect 4529 5931 4530 5935
rect 4534 5931 4535 5935
rect 4539 5931 4540 5935
rect 4544 5931 4545 5935
rect 4549 5931 4550 5935
rect 4554 5931 4555 5935
rect 4826 5934 5086 5937
rect 4525 5930 4559 5931
rect 4529 5926 4530 5930
rect 4534 5926 4535 5930
rect 4539 5926 4540 5930
rect 4544 5926 4545 5930
rect 4549 5926 4550 5930
rect 4554 5926 4555 5930
rect 4525 5925 4559 5926
rect 4529 5921 4530 5925
rect 4534 5921 4535 5925
rect 4539 5921 4540 5925
rect 4544 5921 4545 5925
rect 4549 5921 4550 5925
rect 4554 5921 4555 5925
rect 4525 5920 4559 5921
rect 4529 5916 4530 5920
rect 4534 5916 4535 5920
rect 4539 5916 4540 5920
rect 4544 5916 4545 5920
rect 4549 5916 4550 5920
rect 4554 5916 4555 5920
rect 4826 5882 5086 5885
rect 4826 5628 4829 5882
rect 5083 5628 5086 5882
rect 4483 5622 4484 5626
rect 4488 5622 4489 5626
rect 4493 5622 4494 5626
rect 4498 5622 4499 5626
rect 4503 5622 4504 5626
rect 4508 5622 4509 5626
rect 4479 5621 4513 5622
rect 4483 5617 4484 5621
rect 4488 5617 4489 5621
rect 4493 5617 4494 5621
rect 4498 5617 4499 5621
rect 4503 5617 4504 5621
rect 4508 5617 4509 5621
rect 4479 5616 4513 5617
rect 4483 5612 4484 5616
rect 4488 5612 4489 5616
rect 4493 5612 4494 5616
rect 4498 5612 4499 5616
rect 4503 5612 4504 5616
rect 4508 5612 4509 5616
rect 4479 5611 4513 5612
rect 4483 5607 4484 5611
rect 4488 5607 4489 5611
rect 4493 5607 4494 5611
rect 4498 5607 4499 5611
rect 4503 5607 4504 5611
rect 4508 5607 4509 5611
rect 4529 5622 4530 5626
rect 4534 5622 4535 5626
rect 4539 5622 4540 5626
rect 4544 5622 4545 5626
rect 4549 5622 4550 5626
rect 4554 5622 4555 5626
rect 4826 5625 5086 5628
rect 4525 5621 4559 5622
rect 4529 5617 4530 5621
rect 4534 5617 4535 5621
rect 4539 5617 4540 5621
rect 4544 5617 4545 5621
rect 4549 5617 4550 5621
rect 4554 5617 4555 5621
rect 4525 5616 4559 5617
rect 4529 5612 4530 5616
rect 4534 5612 4535 5616
rect 4539 5612 4540 5616
rect 4544 5612 4545 5616
rect 4549 5612 4550 5616
rect 4554 5612 4555 5616
rect 4525 5611 4559 5612
rect 4529 5607 4530 5611
rect 4534 5607 4535 5611
rect 4539 5607 4540 5611
rect 4544 5607 4545 5611
rect 4549 5607 4550 5611
rect 4554 5607 4555 5611
rect 4826 5573 5086 5576
rect 4826 5319 4829 5573
rect 5083 5319 5086 5573
rect 4483 5313 4484 5317
rect 4488 5313 4489 5317
rect 4493 5313 4494 5317
rect 4498 5313 4499 5317
rect 4503 5313 4504 5317
rect 4508 5313 4509 5317
rect 4479 5312 4513 5313
rect 4483 5308 4484 5312
rect 4488 5308 4489 5312
rect 4493 5308 4494 5312
rect 4498 5308 4499 5312
rect 4503 5308 4504 5312
rect 4508 5308 4509 5312
rect 4479 5307 4513 5308
rect 4483 5303 4484 5307
rect 4488 5303 4489 5307
rect 4493 5303 4494 5307
rect 4498 5303 4499 5307
rect 4503 5303 4504 5307
rect 4508 5303 4509 5307
rect 4479 5302 4513 5303
rect 4483 5298 4484 5302
rect 4488 5298 4489 5302
rect 4493 5298 4494 5302
rect 4498 5298 4499 5302
rect 4503 5298 4504 5302
rect 4508 5298 4509 5302
rect 4529 5313 4530 5317
rect 4534 5313 4535 5317
rect 4539 5313 4540 5317
rect 4544 5313 4545 5317
rect 4549 5313 4550 5317
rect 4554 5313 4555 5317
rect 4826 5316 5086 5319
rect 4525 5312 4559 5313
rect 4529 5308 4530 5312
rect 4534 5308 4535 5312
rect 4539 5308 4540 5312
rect 4544 5308 4545 5312
rect 4549 5308 4550 5312
rect 4554 5308 4555 5312
rect 4525 5307 4559 5308
rect 4529 5303 4530 5307
rect 4534 5303 4535 5307
rect 4539 5303 4540 5307
rect 4544 5303 4545 5307
rect 4549 5303 4550 5307
rect 4554 5303 4555 5307
rect 4525 5302 4559 5303
rect 4529 5298 4530 5302
rect 4534 5298 4535 5302
rect 4539 5298 4540 5302
rect 4544 5298 4545 5302
rect 4549 5298 4550 5302
rect 4554 5298 4555 5302
rect 4826 5264 5086 5267
rect 4826 5010 4829 5264
rect 5083 5010 5086 5264
rect 4483 5004 4484 5008
rect 4488 5004 4489 5008
rect 4493 5004 4494 5008
rect 4498 5004 4499 5008
rect 4503 5004 4504 5008
rect 4508 5004 4509 5008
rect 4479 5003 4513 5004
rect 4483 4999 4484 5003
rect 4488 4999 4489 5003
rect 4493 4999 4494 5003
rect 4498 4999 4499 5003
rect 4503 4999 4504 5003
rect 4508 4999 4509 5003
rect 4479 4998 4513 4999
rect 4483 4994 4484 4998
rect 4488 4994 4489 4998
rect 4493 4994 4494 4998
rect 4498 4994 4499 4998
rect 4503 4994 4504 4998
rect 4508 4994 4509 4998
rect 4479 4993 4513 4994
rect 4483 4989 4484 4993
rect 4488 4989 4489 4993
rect 4493 4989 4494 4993
rect 4498 4989 4499 4993
rect 4503 4989 4504 4993
rect 4508 4989 4509 4993
rect 4529 5004 4530 5008
rect 4534 5004 4535 5008
rect 4539 5004 4540 5008
rect 4544 5004 4545 5008
rect 4549 5004 4550 5008
rect 4554 5004 4555 5008
rect 4826 5007 5086 5010
rect 4525 5003 4559 5004
rect 4529 4999 4530 5003
rect 4534 4999 4535 5003
rect 4539 4999 4540 5003
rect 4544 4999 4545 5003
rect 4549 4999 4550 5003
rect 4554 4999 4555 5003
rect 4525 4998 4559 4999
rect 4529 4994 4530 4998
rect 4534 4994 4535 4998
rect 4539 4994 4540 4998
rect 4544 4994 4545 4998
rect 4549 4994 4550 4998
rect 4554 4994 4555 4998
rect 4525 4993 4559 4994
rect 4529 4989 4530 4993
rect 4534 4989 4535 4993
rect 4539 4989 4540 4993
rect 4544 4989 4545 4993
rect 4549 4989 4550 4993
rect 4554 4989 4555 4993
rect 2670 4928 2674 4932
rect 2378 4813 2384 4835
rect 2670 4739 2675 4928
rect 4483 4811 4484 4815
rect 4488 4811 4489 4815
rect 4493 4811 4494 4815
rect 4498 4811 4499 4815
rect 4503 4811 4504 4815
rect 4508 4811 4509 4815
rect 4479 4810 4513 4811
rect 4483 4806 4484 4810
rect 4488 4806 4489 4810
rect 4493 4806 4494 4810
rect 4498 4806 4499 4810
rect 4503 4806 4504 4810
rect 4508 4806 4509 4810
rect 4479 4805 4513 4806
rect 4483 4801 4484 4805
rect 4488 4801 4489 4805
rect 4493 4801 4494 4805
rect 4498 4801 4499 4805
rect 4503 4801 4504 4805
rect 4508 4801 4509 4805
rect 4479 4800 4513 4801
rect 4483 4796 4484 4800
rect 4488 4796 4489 4800
rect 4493 4796 4494 4800
rect 4498 4796 4499 4800
rect 4503 4796 4504 4800
rect 4508 4796 4509 4800
rect 4529 4811 4530 4815
rect 4534 4811 4535 4815
rect 4539 4811 4540 4815
rect 4544 4811 4545 4815
rect 4549 4811 4550 4815
rect 4554 4811 4555 4815
rect 4525 4810 4559 4811
rect 4529 4806 4530 4810
rect 4534 4806 4535 4810
rect 4539 4806 4540 4810
rect 4544 4806 4545 4810
rect 4549 4806 4550 4810
rect 4554 4806 4555 4810
rect 4525 4805 4559 4806
rect 4529 4801 4530 4805
rect 4534 4801 4535 4805
rect 4539 4801 4540 4805
rect 4544 4801 4545 4805
rect 4549 4801 4550 4805
rect 4554 4801 4555 4805
rect 4525 4800 4559 4801
rect 4529 4796 4530 4800
rect 4534 4796 4535 4800
rect 4539 4796 4540 4800
rect 4544 4796 4545 4800
rect 4549 4796 4550 4800
rect 4554 4796 4555 4800
rect 4483 4785 4484 4789
rect 4488 4785 4489 4789
rect 4493 4785 4494 4789
rect 4498 4785 4499 4789
rect 4503 4785 4504 4789
rect 4508 4785 4509 4789
rect 4479 4784 4513 4785
rect 4483 4780 4484 4784
rect 4488 4780 4489 4784
rect 4493 4780 4494 4784
rect 4498 4780 4499 4784
rect 4503 4780 4504 4784
rect 4508 4780 4509 4784
rect 4479 4779 4513 4780
rect 4483 4775 4484 4779
rect 4488 4775 4489 4779
rect 4493 4775 4494 4779
rect 4498 4775 4499 4779
rect 4503 4775 4504 4779
rect 4508 4775 4509 4779
rect 4479 4774 4513 4775
rect 4483 4770 4484 4774
rect 4488 4770 4489 4774
rect 4493 4770 4494 4774
rect 4498 4770 4499 4774
rect 4503 4770 4504 4774
rect 4508 4770 4509 4774
rect 4529 4785 4530 4789
rect 4534 4785 4535 4789
rect 4539 4785 4540 4789
rect 4544 4785 4545 4789
rect 4549 4785 4550 4789
rect 4554 4785 4555 4789
rect 4525 4784 4559 4785
rect 4529 4780 4530 4784
rect 4534 4780 4535 4784
rect 4539 4780 4540 4784
rect 4544 4780 4545 4784
rect 4549 4780 4550 4784
rect 4554 4780 4555 4784
rect 4525 4779 4559 4780
rect 4529 4775 4530 4779
rect 4534 4775 4535 4779
rect 4539 4775 4540 4779
rect 4544 4775 4545 4779
rect 4549 4775 4550 4779
rect 4554 4775 4555 4779
rect 4525 4774 4559 4775
rect 4529 4770 4530 4774
rect 4534 4770 4535 4774
rect 4539 4770 4540 4774
rect 4544 4770 4545 4774
rect 4549 4770 4550 4774
rect 4554 4770 4555 4774
rect 4483 4759 4484 4763
rect 4488 4759 4489 4763
rect 4493 4759 4494 4763
rect 4498 4759 4499 4763
rect 4503 4759 4504 4763
rect 4508 4759 4509 4763
rect 4479 4758 4513 4759
rect 4483 4754 4484 4758
rect 4488 4754 4489 4758
rect 4493 4754 4494 4758
rect 4498 4754 4499 4758
rect 4503 4754 4504 4758
rect 4508 4754 4509 4758
rect 4479 4753 4513 4754
rect 4483 4749 4484 4753
rect 4488 4749 4489 4753
rect 4493 4749 4494 4753
rect 4498 4749 4499 4753
rect 4503 4749 4504 4753
rect 4508 4749 4509 4753
rect 4479 4748 4513 4749
rect 4483 4744 4484 4748
rect 4488 4744 4489 4748
rect 4493 4744 4494 4748
rect 4498 4744 4499 4748
rect 4503 4744 4504 4748
rect 4508 4744 4509 4748
rect 4529 4759 4530 4763
rect 4534 4759 4535 4763
rect 4539 4759 4540 4763
rect 4544 4759 4545 4763
rect 4549 4759 4550 4763
rect 4554 4759 4555 4763
rect 4525 4758 4559 4759
rect 4529 4754 4530 4758
rect 4534 4754 4535 4758
rect 4539 4754 4540 4758
rect 4544 4754 4545 4758
rect 4549 4754 4550 4758
rect 4554 4754 4555 4758
rect 4525 4753 4559 4754
rect 4529 4749 4530 4753
rect 4534 4749 4535 4753
rect 4539 4749 4540 4753
rect 4544 4749 4545 4753
rect 4549 4749 4550 4753
rect 4554 4749 4555 4753
rect 4525 4748 4559 4749
rect 4529 4744 4530 4748
rect 4534 4744 4535 4748
rect 4539 4744 4540 4748
rect 4544 4744 4545 4748
rect 4549 4744 4550 4748
rect 4554 4744 4555 4748
rect 4483 4733 4484 4737
rect 4488 4733 4489 4737
rect 4493 4733 4494 4737
rect 4498 4733 4499 4737
rect 4503 4733 4504 4737
rect 4508 4733 4509 4737
rect 4479 4732 4513 4733
rect 4483 4728 4484 4732
rect 4488 4728 4489 4732
rect 4493 4728 4494 4732
rect 4498 4728 4499 4732
rect 4503 4728 4504 4732
rect 4508 4728 4509 4732
rect 4479 4727 4513 4728
rect 4483 4723 4484 4727
rect 4488 4723 4489 4727
rect 4493 4723 4494 4727
rect 4498 4723 4499 4727
rect 4503 4723 4504 4727
rect 4508 4723 4509 4727
rect 4479 4722 4513 4723
rect 2911 4695 2915 4721
rect 2914 4691 2915 4695
rect 2993 4698 2999 4721
rect 4483 4718 4484 4722
rect 4488 4718 4489 4722
rect 4493 4718 4494 4722
rect 4498 4718 4499 4722
rect 4503 4718 4504 4722
rect 4508 4718 4509 4722
rect 4529 4733 4530 4737
rect 4534 4733 4535 4737
rect 4539 4733 4540 4737
rect 4544 4733 4545 4737
rect 4549 4733 4550 4737
rect 4554 4733 4555 4737
rect 4525 4732 4559 4733
rect 4529 4728 4530 4732
rect 4534 4728 4535 4732
rect 4539 4728 4540 4732
rect 4544 4728 4545 4732
rect 4549 4728 4550 4732
rect 4554 4728 4555 4732
rect 4525 4727 4559 4728
rect 4529 4723 4530 4727
rect 4534 4723 4535 4727
rect 4539 4723 4540 4727
rect 4544 4723 4545 4727
rect 4549 4723 4550 4727
rect 4554 4723 4555 4727
rect 4525 4722 4559 4723
rect 4529 4718 4530 4722
rect 4534 4718 4535 4722
rect 4539 4718 4540 4722
rect 4544 4718 4545 4722
rect 4549 4718 4550 4722
rect 4554 4718 4555 4722
rect 4483 4707 4484 4711
rect 4488 4707 4489 4711
rect 4493 4707 4494 4711
rect 4498 4707 4499 4711
rect 4503 4707 4504 4711
rect 4508 4707 4509 4711
rect 4479 4706 4513 4707
rect 4483 4702 4484 4706
rect 4488 4702 4489 4706
rect 4493 4702 4494 4706
rect 4498 4702 4499 4706
rect 4503 4702 4504 4706
rect 4508 4702 4509 4706
rect 4479 4701 4513 4702
rect 2993 4691 3006 4698
rect 4483 4697 4484 4701
rect 4488 4697 4489 4701
rect 4493 4697 4494 4701
rect 4498 4697 4499 4701
rect 4503 4697 4504 4701
rect 4508 4697 4509 4701
rect 4479 4696 4513 4697
rect 4483 4692 4484 4696
rect 4488 4692 4489 4696
rect 4493 4692 4494 4696
rect 4498 4692 4499 4696
rect 4503 4692 4504 4696
rect 4508 4692 4509 4696
rect 4529 4707 4530 4711
rect 4534 4707 4535 4711
rect 4539 4707 4540 4711
rect 4544 4707 4545 4711
rect 4549 4707 4550 4711
rect 4554 4707 4555 4711
rect 4525 4706 4559 4707
rect 4529 4702 4530 4706
rect 4534 4702 4535 4706
rect 4539 4702 4540 4706
rect 4544 4702 4545 4706
rect 4549 4702 4550 4706
rect 4554 4702 4555 4706
rect 4525 4701 4559 4702
rect 4529 4697 4530 4701
rect 4534 4697 4535 4701
rect 4539 4697 4540 4701
rect 4544 4697 4545 4701
rect 4549 4697 4550 4701
rect 4554 4697 4555 4701
rect 4525 4696 4559 4697
rect 4529 4692 4530 4696
rect 4534 4692 4535 4696
rect 4539 4692 4540 4696
rect 4544 4692 4545 4696
rect 4549 4692 4550 4696
rect 4554 4692 4555 4696
rect 1810 4653 1830 4655
rect 1814 4649 1815 4653
rect 1819 4649 1820 4653
rect 1824 4649 1825 4653
rect 1829 4649 1830 4653
rect 1810 4648 1830 4649
rect 1814 4644 1815 4648
rect 1819 4644 1820 4648
rect 1824 4644 1825 4648
rect 1829 4644 1830 4648
rect 1810 4643 1830 4644
rect 1814 4639 1815 4643
rect 1819 4639 1820 4643
rect 1824 4639 1825 4643
rect 1829 4639 1830 4643
rect 1810 4638 1830 4639
rect 1814 4634 1815 4638
rect 1819 4634 1820 4638
rect 1824 4634 1825 4638
rect 1829 4634 1830 4638
rect 1810 4633 1830 4634
rect 1814 4629 1815 4633
rect 1819 4629 1820 4633
rect 1824 4629 1825 4633
rect 1829 4629 1830 4633
rect 1810 4628 1830 4629
rect 761 4624 762 4628
rect 766 4624 767 4628
rect 771 4624 772 4628
rect 757 4623 776 4624
rect 761 4619 762 4623
rect 766 4619 767 4623
rect 771 4619 772 4623
rect 757 4618 776 4619
rect 761 4614 762 4618
rect 766 4614 767 4618
rect 771 4614 772 4618
rect 757 4613 776 4614
rect 761 4609 762 4613
rect 766 4609 767 4613
rect 771 4609 772 4613
rect 757 4608 776 4609
rect 761 4604 762 4608
rect 766 4604 767 4608
rect 771 4604 772 4608
rect 757 4603 776 4604
rect 761 4599 762 4603
rect 766 4599 767 4603
rect 771 4599 772 4603
rect 757 4598 776 4599
rect 761 4594 762 4598
rect 766 4594 767 4598
rect 771 4594 772 4598
rect 787 4624 788 4628
rect 792 4624 793 4628
rect 797 4624 798 4628
rect 783 4623 802 4624
rect 787 4619 788 4623
rect 792 4619 793 4623
rect 797 4619 798 4623
rect 783 4618 802 4619
rect 787 4614 788 4618
rect 792 4614 793 4618
rect 797 4614 798 4618
rect 783 4613 802 4614
rect 787 4609 788 4613
rect 792 4609 793 4613
rect 797 4609 798 4613
rect 783 4608 802 4609
rect 787 4604 788 4608
rect 792 4604 793 4608
rect 797 4604 798 4608
rect 783 4603 802 4604
rect 787 4599 788 4603
rect 792 4599 793 4603
rect 797 4599 798 4603
rect 783 4598 802 4599
rect 787 4594 788 4598
rect 792 4594 793 4598
rect 797 4594 798 4598
rect 813 4624 814 4628
rect 818 4624 819 4628
rect 823 4624 824 4628
rect 809 4623 828 4624
rect 813 4619 814 4623
rect 818 4619 819 4623
rect 823 4619 824 4623
rect 809 4618 828 4619
rect 813 4614 814 4618
rect 818 4614 819 4618
rect 823 4614 824 4618
rect 809 4613 828 4614
rect 813 4609 814 4613
rect 818 4609 819 4613
rect 823 4609 824 4613
rect 809 4608 828 4609
rect 813 4604 814 4608
rect 818 4604 819 4608
rect 823 4604 824 4608
rect 809 4603 828 4604
rect 813 4599 814 4603
rect 818 4599 819 4603
rect 823 4599 824 4603
rect 809 4598 828 4599
rect 813 4594 814 4598
rect 818 4594 819 4598
rect 823 4594 824 4598
rect 839 4624 840 4628
rect 844 4624 845 4628
rect 849 4624 850 4628
rect 835 4623 854 4624
rect 839 4619 840 4623
rect 844 4619 845 4623
rect 849 4619 850 4623
rect 835 4618 854 4619
rect 839 4614 840 4618
rect 844 4614 845 4618
rect 849 4614 850 4618
rect 835 4613 854 4614
rect 839 4609 840 4613
rect 844 4609 845 4613
rect 849 4609 850 4613
rect 835 4608 854 4609
rect 839 4604 840 4608
rect 844 4604 845 4608
rect 849 4604 850 4608
rect 835 4603 854 4604
rect 839 4599 840 4603
rect 844 4599 845 4603
rect 849 4599 850 4603
rect 835 4598 854 4599
rect 839 4594 840 4598
rect 844 4594 845 4598
rect 849 4594 850 4598
rect 865 4624 866 4628
rect 870 4624 871 4628
rect 875 4624 876 4628
rect 861 4623 880 4624
rect 865 4619 866 4623
rect 870 4619 871 4623
rect 875 4619 876 4623
rect 861 4618 880 4619
rect 865 4614 866 4618
rect 870 4614 871 4618
rect 875 4614 876 4618
rect 861 4613 880 4614
rect 865 4609 866 4613
rect 870 4609 871 4613
rect 875 4609 876 4613
rect 861 4608 880 4609
rect 865 4604 866 4608
rect 870 4604 871 4608
rect 875 4604 876 4608
rect 861 4603 880 4604
rect 865 4599 866 4603
rect 870 4599 871 4603
rect 875 4599 876 4603
rect 861 4598 880 4599
rect 865 4594 866 4598
rect 870 4594 871 4598
rect 875 4594 876 4598
rect 1057 4624 1058 4628
rect 1062 4624 1063 4628
rect 1067 4624 1068 4628
rect 1053 4623 1072 4624
rect 1057 4619 1058 4623
rect 1062 4619 1063 4623
rect 1067 4619 1068 4623
rect 1053 4618 1072 4619
rect 1057 4614 1058 4618
rect 1062 4614 1063 4618
rect 1067 4614 1068 4618
rect 1366 4624 1367 4628
rect 1371 4624 1372 4628
rect 1376 4624 1377 4628
rect 1362 4623 1381 4624
rect 1366 4619 1367 4623
rect 1371 4619 1372 4623
rect 1376 4619 1377 4623
rect 1362 4618 1381 4619
rect 1366 4614 1367 4618
rect 1371 4614 1372 4618
rect 1376 4614 1377 4618
rect 1675 4624 1676 4628
rect 1680 4624 1681 4628
rect 1685 4624 1686 4628
rect 1671 4623 1690 4624
rect 1675 4619 1676 4623
rect 1680 4619 1681 4623
rect 1685 4619 1686 4623
rect 1671 4618 1690 4619
rect 1675 4614 1676 4618
rect 1680 4614 1681 4618
rect 1685 4614 1686 4618
rect 1053 4613 1072 4614
rect 1057 4609 1058 4613
rect 1062 4609 1063 4613
rect 1067 4609 1068 4613
rect 1053 4608 1072 4609
rect 1057 4604 1058 4608
rect 1062 4604 1063 4608
rect 1067 4604 1068 4608
rect 1053 4603 1072 4604
rect 1057 4599 1058 4603
rect 1062 4599 1063 4603
rect 1067 4599 1068 4603
rect 1053 4598 1072 4599
rect 1057 4594 1058 4598
rect 1062 4594 1063 4598
rect 1067 4594 1068 4598
rect 1075 4611 1131 4613
rect 1075 4607 1077 4611
rect 1081 4607 1082 4611
rect 1086 4607 1087 4611
rect 1091 4607 1092 4611
rect 1096 4607 1097 4611
rect 1101 4607 1102 4611
rect 1106 4607 1107 4611
rect 1111 4607 1112 4611
rect 1116 4607 1117 4611
rect 1121 4607 1122 4611
rect 1126 4607 1127 4611
rect 1075 4606 1131 4607
rect 1075 4602 1077 4606
rect 1081 4602 1082 4606
rect 1086 4602 1087 4606
rect 1091 4602 1092 4606
rect 1096 4602 1097 4606
rect 1101 4602 1102 4606
rect 1106 4602 1107 4606
rect 1111 4602 1112 4606
rect 1116 4602 1117 4606
rect 1121 4602 1122 4606
rect 1126 4602 1127 4606
rect 1075 4601 1131 4602
rect 1075 4597 1077 4601
rect 1081 4597 1082 4601
rect 1086 4597 1087 4601
rect 1091 4597 1092 4601
rect 1096 4597 1097 4601
rect 1101 4597 1102 4601
rect 1106 4597 1107 4601
rect 1111 4597 1112 4601
rect 1116 4597 1117 4601
rect 1121 4597 1122 4601
rect 1126 4597 1127 4601
rect 1075 4596 1131 4597
rect 1075 4592 1077 4596
rect 1081 4592 1082 4596
rect 1086 4592 1087 4596
rect 1091 4592 1092 4596
rect 1096 4592 1097 4596
rect 1101 4592 1102 4596
rect 1106 4592 1107 4596
rect 1111 4592 1112 4596
rect 1116 4592 1117 4596
rect 1121 4592 1122 4596
rect 1126 4592 1127 4596
rect 1247 4611 1315 4614
rect 1247 4607 1249 4611
rect 1253 4607 1254 4611
rect 1258 4607 1259 4611
rect 1263 4607 1264 4611
rect 1268 4607 1269 4611
rect 1273 4607 1274 4611
rect 1278 4607 1279 4611
rect 1283 4607 1284 4611
rect 1288 4607 1289 4611
rect 1293 4607 1294 4611
rect 1298 4607 1299 4611
rect 1303 4607 1304 4611
rect 1308 4607 1309 4611
rect 1313 4607 1315 4611
rect 1247 4606 1315 4607
rect 1247 4602 1249 4606
rect 1253 4602 1254 4606
rect 1258 4602 1259 4606
rect 1263 4602 1264 4606
rect 1268 4602 1269 4606
rect 1273 4602 1274 4606
rect 1278 4602 1279 4606
rect 1283 4602 1284 4606
rect 1288 4602 1289 4606
rect 1293 4602 1294 4606
rect 1298 4602 1299 4606
rect 1303 4602 1304 4606
rect 1308 4602 1309 4606
rect 1313 4602 1315 4606
rect 761 4578 762 4582
rect 766 4578 767 4582
rect 771 4578 772 4582
rect 757 4577 776 4578
rect 761 4573 762 4577
rect 766 4573 767 4577
rect 771 4573 772 4577
rect 757 4572 776 4573
rect 761 4568 762 4572
rect 766 4568 767 4572
rect 771 4568 772 4572
rect 757 4567 776 4568
rect 761 4563 762 4567
rect 766 4563 767 4567
rect 771 4563 772 4567
rect 757 4562 776 4563
rect 761 4558 762 4562
rect 766 4558 767 4562
rect 771 4558 772 4562
rect 757 4557 776 4558
rect 761 4553 762 4557
rect 766 4553 767 4557
rect 771 4553 772 4557
rect 757 4552 776 4553
rect 761 4548 762 4552
rect 766 4548 767 4552
rect 771 4548 772 4552
rect 787 4578 788 4582
rect 792 4578 793 4582
rect 797 4578 798 4582
rect 783 4577 802 4578
rect 787 4573 788 4577
rect 792 4573 793 4577
rect 797 4573 798 4577
rect 783 4572 802 4573
rect 787 4568 788 4572
rect 792 4568 793 4572
rect 797 4568 798 4572
rect 783 4567 802 4568
rect 787 4563 788 4567
rect 792 4563 793 4567
rect 797 4563 798 4567
rect 783 4562 802 4563
rect 787 4558 788 4562
rect 792 4558 793 4562
rect 797 4558 798 4562
rect 783 4557 802 4558
rect 787 4553 788 4557
rect 792 4553 793 4557
rect 797 4553 798 4557
rect 783 4552 802 4553
rect 787 4548 788 4552
rect 792 4548 793 4552
rect 797 4548 798 4552
rect 813 4578 814 4582
rect 818 4578 819 4582
rect 823 4578 824 4582
rect 809 4577 828 4578
rect 813 4573 814 4577
rect 818 4573 819 4577
rect 823 4573 824 4577
rect 809 4572 828 4573
rect 813 4568 814 4572
rect 818 4568 819 4572
rect 823 4568 824 4572
rect 809 4567 828 4568
rect 813 4563 814 4567
rect 818 4563 819 4567
rect 823 4563 824 4567
rect 809 4562 828 4563
rect 813 4558 814 4562
rect 818 4558 819 4562
rect 823 4558 824 4562
rect 809 4557 828 4558
rect 813 4553 814 4557
rect 818 4553 819 4557
rect 823 4553 824 4557
rect 809 4552 828 4553
rect 813 4548 814 4552
rect 818 4548 819 4552
rect 823 4548 824 4552
rect 839 4578 840 4582
rect 844 4578 845 4582
rect 849 4578 850 4582
rect 835 4577 854 4578
rect 839 4573 840 4577
rect 844 4573 845 4577
rect 849 4573 850 4577
rect 835 4572 854 4573
rect 839 4568 840 4572
rect 844 4568 845 4572
rect 849 4568 850 4572
rect 835 4567 854 4568
rect 839 4563 840 4567
rect 844 4563 845 4567
rect 849 4563 850 4567
rect 835 4562 854 4563
rect 839 4558 840 4562
rect 844 4558 845 4562
rect 849 4558 850 4562
rect 835 4557 854 4558
rect 839 4553 840 4557
rect 844 4553 845 4557
rect 849 4553 850 4557
rect 835 4552 854 4553
rect 839 4548 840 4552
rect 844 4548 845 4552
rect 849 4548 850 4552
rect 865 4578 866 4582
rect 870 4578 871 4582
rect 875 4578 876 4582
rect 861 4577 880 4578
rect 865 4573 866 4577
rect 870 4573 871 4577
rect 875 4573 876 4577
rect 861 4572 880 4573
rect 865 4568 866 4572
rect 870 4568 871 4572
rect 875 4568 876 4572
rect 861 4567 880 4568
rect 865 4563 866 4567
rect 870 4563 871 4567
rect 875 4563 876 4567
rect 861 4562 880 4563
rect 865 4558 866 4562
rect 870 4558 871 4562
rect 875 4558 876 4562
rect 861 4557 880 4558
rect 865 4553 866 4557
rect 870 4553 871 4557
rect 875 4553 876 4557
rect 861 4552 880 4553
rect 865 4548 866 4552
rect 870 4548 871 4552
rect 875 4548 876 4552
rect 1057 4578 1058 4582
rect 1062 4578 1063 4582
rect 1067 4578 1068 4582
rect 1053 4577 1072 4578
rect 1057 4573 1058 4577
rect 1062 4573 1063 4577
rect 1067 4573 1068 4577
rect 1053 4572 1072 4573
rect 1057 4568 1058 4572
rect 1062 4568 1063 4572
rect 1067 4568 1068 4572
rect 1053 4567 1072 4568
rect 1057 4563 1058 4567
rect 1062 4563 1063 4567
rect 1067 4563 1068 4567
rect 1053 4562 1072 4563
rect 1057 4558 1058 4562
rect 1062 4558 1063 4562
rect 1067 4558 1068 4562
rect 1053 4557 1072 4558
rect 1057 4553 1058 4557
rect 1062 4553 1063 4557
rect 1067 4553 1068 4557
rect 1053 4552 1072 4553
rect 1057 4548 1058 4552
rect 1062 4548 1063 4552
rect 1067 4548 1068 4552
rect 1087 4554 1155 4557
rect 1087 4550 1089 4554
rect 1093 4550 1094 4554
rect 1098 4550 1099 4554
rect 1103 4550 1104 4554
rect 1108 4550 1109 4554
rect 1113 4550 1114 4554
rect 1118 4550 1119 4554
rect 1123 4550 1124 4554
rect 1128 4550 1129 4554
rect 1133 4550 1134 4554
rect 1138 4550 1139 4554
rect 1143 4550 1144 4554
rect 1148 4550 1149 4554
rect 1153 4550 1155 4554
rect 1087 4549 1155 4550
rect 1087 4545 1089 4549
rect 1093 4545 1094 4549
rect 1098 4545 1099 4549
rect 1103 4545 1104 4549
rect 1108 4545 1109 4549
rect 1113 4545 1114 4549
rect 1118 4545 1119 4549
rect 1123 4545 1124 4549
rect 1128 4545 1129 4549
rect 1133 4545 1134 4549
rect 1138 4545 1139 4549
rect 1143 4545 1144 4549
rect 1148 4545 1149 4549
rect 1153 4545 1155 4549
rect 99 4053 1031 4528
rect 1087 4466 1155 4545
rect 1169 4519 1173 4531
rect 1169 4503 1173 4515
rect 1169 4487 1173 4499
rect 1227 4519 1231 4531
rect 1227 4503 1231 4515
rect 1227 4487 1231 4499
rect 1091 4462 1094 4466
rect 1098 4462 1099 4466
rect 1103 4462 1104 4466
rect 1108 4462 1109 4466
rect 1113 4462 1114 4466
rect 1118 4462 1119 4466
rect 1123 4462 1124 4466
rect 1128 4462 1129 4466
rect 1133 4462 1134 4466
rect 1138 4462 1139 4466
rect 1143 4462 1144 4466
rect 1148 4462 1151 4466
rect 1247 4466 1315 4602
rect 1362 4613 1381 4614
rect 1366 4609 1367 4613
rect 1371 4609 1372 4613
rect 1376 4609 1377 4613
rect 1362 4608 1381 4609
rect 1366 4604 1367 4608
rect 1371 4604 1372 4608
rect 1376 4604 1377 4608
rect 1362 4603 1381 4604
rect 1366 4599 1367 4603
rect 1371 4599 1372 4603
rect 1376 4599 1377 4603
rect 1362 4598 1381 4599
rect 1366 4594 1367 4598
rect 1371 4594 1372 4598
rect 1376 4594 1377 4598
rect 1384 4611 1440 4613
rect 1384 4607 1386 4611
rect 1390 4607 1391 4611
rect 1395 4607 1396 4611
rect 1400 4607 1401 4611
rect 1405 4607 1406 4611
rect 1410 4607 1411 4611
rect 1415 4607 1416 4611
rect 1420 4607 1421 4611
rect 1425 4607 1426 4611
rect 1430 4607 1431 4611
rect 1435 4607 1436 4611
rect 1384 4606 1440 4607
rect 1384 4602 1386 4606
rect 1390 4602 1391 4606
rect 1395 4602 1396 4606
rect 1400 4602 1401 4606
rect 1405 4602 1406 4606
rect 1410 4602 1411 4606
rect 1415 4602 1416 4606
rect 1420 4602 1421 4606
rect 1425 4602 1426 4606
rect 1430 4602 1431 4606
rect 1435 4602 1436 4606
rect 1384 4601 1440 4602
rect 1384 4597 1386 4601
rect 1390 4597 1391 4601
rect 1395 4597 1396 4601
rect 1400 4597 1401 4601
rect 1405 4597 1406 4601
rect 1410 4597 1411 4601
rect 1415 4597 1416 4601
rect 1420 4597 1421 4601
rect 1425 4597 1426 4601
rect 1430 4597 1431 4601
rect 1435 4597 1436 4601
rect 1384 4596 1440 4597
rect 1384 4592 1386 4596
rect 1390 4592 1391 4596
rect 1395 4592 1396 4596
rect 1400 4592 1401 4596
rect 1405 4592 1406 4596
rect 1410 4592 1411 4596
rect 1415 4592 1416 4596
rect 1420 4592 1421 4596
rect 1425 4592 1426 4596
rect 1430 4592 1431 4596
rect 1435 4592 1436 4596
rect 1556 4611 1624 4614
rect 1556 4607 1558 4611
rect 1562 4607 1563 4611
rect 1567 4607 1568 4611
rect 1572 4607 1573 4611
rect 1577 4607 1578 4611
rect 1582 4607 1583 4611
rect 1587 4607 1588 4611
rect 1592 4607 1593 4611
rect 1597 4607 1598 4611
rect 1602 4607 1603 4611
rect 1607 4607 1608 4611
rect 1612 4607 1613 4611
rect 1617 4607 1618 4611
rect 1622 4607 1624 4611
rect 1556 4606 1624 4607
rect 1556 4602 1558 4606
rect 1562 4602 1563 4606
rect 1567 4602 1568 4606
rect 1572 4602 1573 4606
rect 1577 4602 1578 4606
rect 1582 4602 1583 4606
rect 1587 4602 1588 4606
rect 1592 4602 1593 4606
rect 1597 4602 1598 4606
rect 1602 4602 1603 4606
rect 1607 4602 1608 4606
rect 1612 4602 1613 4606
rect 1617 4602 1618 4606
rect 1622 4602 1624 4606
rect 1327 4578 1348 4580
rect 1331 4574 1332 4578
rect 1336 4574 1337 4578
rect 1341 4574 1342 4578
rect 1346 4574 1348 4578
rect 1327 4573 1348 4574
rect 1331 4569 1332 4573
rect 1336 4569 1337 4573
rect 1341 4569 1342 4573
rect 1346 4569 1348 4573
rect 1327 4568 1348 4569
rect 1331 4564 1332 4568
rect 1336 4564 1337 4568
rect 1341 4564 1342 4568
rect 1346 4564 1348 4568
rect 1327 4563 1348 4564
rect 1331 4559 1332 4563
rect 1336 4559 1337 4563
rect 1341 4559 1342 4563
rect 1346 4559 1348 4563
rect 1327 4558 1348 4559
rect 1331 4554 1332 4558
rect 1336 4554 1337 4558
rect 1341 4554 1342 4558
rect 1346 4554 1348 4558
rect 1327 4553 1348 4554
rect 1331 4549 1332 4553
rect 1336 4549 1337 4553
rect 1341 4549 1342 4553
rect 1346 4549 1348 4553
rect 1327 4548 1348 4549
rect 1366 4578 1367 4582
rect 1371 4578 1372 4582
rect 1376 4578 1377 4582
rect 1362 4577 1381 4578
rect 1366 4573 1367 4577
rect 1371 4573 1372 4577
rect 1376 4573 1377 4577
rect 1362 4572 1381 4573
rect 1366 4568 1367 4572
rect 1371 4568 1372 4572
rect 1376 4568 1377 4572
rect 1362 4567 1381 4568
rect 1366 4563 1367 4567
rect 1371 4563 1372 4567
rect 1376 4563 1377 4567
rect 1362 4562 1381 4563
rect 1366 4558 1367 4562
rect 1371 4558 1372 4562
rect 1376 4558 1377 4562
rect 1362 4557 1381 4558
rect 1501 4573 1521 4575
rect 1505 4569 1506 4573
rect 1510 4569 1511 4573
rect 1515 4569 1516 4573
rect 1520 4569 1521 4573
rect 1501 4568 1521 4569
rect 1505 4564 1506 4568
rect 1510 4564 1511 4568
rect 1515 4564 1516 4568
rect 1520 4564 1521 4568
rect 1501 4563 1521 4564
rect 1505 4559 1506 4563
rect 1510 4559 1511 4563
rect 1515 4559 1516 4563
rect 1520 4559 1521 4563
rect 1501 4558 1521 4559
rect 1366 4553 1367 4557
rect 1371 4553 1372 4557
rect 1376 4553 1377 4557
rect 1362 4552 1381 4553
rect 1366 4548 1367 4552
rect 1371 4548 1372 4552
rect 1376 4548 1377 4552
rect 1396 4554 1464 4557
rect 1396 4550 1398 4554
rect 1402 4550 1403 4554
rect 1407 4550 1408 4554
rect 1412 4550 1413 4554
rect 1417 4550 1418 4554
rect 1422 4550 1423 4554
rect 1427 4550 1428 4554
rect 1432 4550 1433 4554
rect 1437 4550 1438 4554
rect 1442 4550 1443 4554
rect 1447 4550 1448 4554
rect 1452 4550 1453 4554
rect 1457 4550 1458 4554
rect 1462 4550 1464 4554
rect 1396 4549 1464 4550
rect 1331 4544 1332 4548
rect 1336 4544 1337 4548
rect 1341 4544 1342 4548
rect 1346 4544 1348 4548
rect 1327 4543 1348 4544
rect 1331 4539 1332 4543
rect 1336 4539 1337 4543
rect 1341 4539 1342 4543
rect 1346 4539 1348 4543
rect 1327 4538 1348 4539
rect 1331 4534 1332 4538
rect 1336 4534 1337 4538
rect 1341 4534 1342 4538
rect 1346 4534 1348 4538
rect 1327 4533 1348 4534
rect 1331 4529 1332 4533
rect 1336 4529 1337 4533
rect 1341 4529 1342 4533
rect 1346 4529 1348 4533
rect 1327 4528 1348 4529
rect 1331 4524 1332 4528
rect 1336 4524 1337 4528
rect 1341 4524 1342 4528
rect 1346 4524 1348 4528
rect 1327 4523 1348 4524
rect 1331 4519 1332 4523
rect 1336 4519 1337 4523
rect 1341 4519 1342 4523
rect 1346 4519 1348 4523
rect 1327 4518 1348 4519
rect 1331 4514 1332 4518
rect 1336 4514 1337 4518
rect 1341 4514 1342 4518
rect 1346 4514 1348 4518
rect 1327 4512 1348 4514
rect 1396 4545 1398 4549
rect 1402 4545 1403 4549
rect 1407 4545 1408 4549
rect 1412 4545 1413 4549
rect 1417 4545 1418 4549
rect 1422 4545 1423 4549
rect 1427 4545 1428 4549
rect 1432 4545 1433 4549
rect 1437 4545 1438 4549
rect 1442 4545 1443 4549
rect 1447 4545 1448 4549
rect 1452 4545 1453 4549
rect 1457 4545 1458 4549
rect 1462 4545 1464 4549
rect 1251 4462 1254 4466
rect 1258 4462 1259 4466
rect 1263 4462 1264 4466
rect 1268 4462 1269 4466
rect 1273 4462 1274 4466
rect 1278 4462 1279 4466
rect 1283 4462 1284 4466
rect 1288 4462 1289 4466
rect 1293 4462 1294 4466
rect 1298 4462 1299 4466
rect 1303 4462 1304 4466
rect 1308 4462 1311 4466
rect 1396 4466 1464 4545
rect 1505 4554 1506 4558
rect 1510 4554 1511 4558
rect 1515 4554 1516 4558
rect 1520 4554 1521 4558
rect 1501 4553 1521 4554
rect 1505 4549 1506 4553
rect 1510 4549 1511 4553
rect 1515 4549 1516 4553
rect 1520 4549 1521 4553
rect 1501 4548 1521 4549
rect 1505 4544 1506 4548
rect 1510 4544 1511 4548
rect 1515 4544 1516 4548
rect 1520 4544 1521 4548
rect 1501 4543 1521 4544
rect 1505 4539 1506 4543
rect 1510 4539 1511 4543
rect 1515 4539 1516 4543
rect 1520 4539 1521 4543
rect 1501 4538 1521 4539
rect 1505 4534 1506 4538
rect 1510 4534 1511 4538
rect 1515 4534 1516 4538
rect 1520 4534 1521 4538
rect 1501 4533 1521 4534
rect 1505 4529 1506 4533
rect 1510 4529 1511 4533
rect 1515 4529 1516 4533
rect 1520 4529 1521 4533
rect 1501 4528 1521 4529
rect 1505 4524 1506 4528
rect 1510 4524 1511 4528
rect 1515 4524 1516 4528
rect 1520 4524 1521 4528
rect 1501 4523 1521 4524
rect 1505 4519 1506 4523
rect 1510 4519 1511 4523
rect 1515 4519 1516 4523
rect 1520 4519 1521 4523
rect 1400 4462 1403 4466
rect 1407 4462 1408 4466
rect 1412 4462 1413 4466
rect 1417 4462 1418 4466
rect 1422 4462 1423 4466
rect 1427 4462 1428 4466
rect 1432 4462 1433 4466
rect 1437 4462 1438 4466
rect 1442 4462 1443 4466
rect 1447 4462 1448 4466
rect 1452 4462 1453 4466
rect 1457 4462 1460 4466
rect 1556 4466 1624 4602
rect 1671 4613 1690 4614
rect 1814 4624 1815 4628
rect 1819 4624 1820 4628
rect 1824 4624 1825 4628
rect 1829 4624 1830 4628
rect 1810 4623 1830 4624
rect 1814 4619 1815 4623
rect 1819 4619 1820 4623
rect 1824 4619 1825 4623
rect 1829 4619 1830 4623
rect 1810 4618 1830 4619
rect 1814 4614 1815 4618
rect 1819 4614 1820 4618
rect 1824 4614 1825 4618
rect 1829 4614 1830 4618
rect 1984 4624 1985 4628
rect 1989 4624 1990 4628
rect 1994 4624 1995 4628
rect 1980 4623 1999 4624
rect 1984 4619 1985 4623
rect 1989 4619 1990 4623
rect 1994 4619 1995 4623
rect 1980 4618 1999 4619
rect 1984 4614 1985 4618
rect 1989 4614 1990 4618
rect 1994 4614 1995 4618
rect 2293 4624 2294 4628
rect 2298 4624 2299 4628
rect 2303 4624 2304 4628
rect 2289 4623 2308 4624
rect 2293 4619 2294 4623
rect 2298 4619 2299 4623
rect 2303 4619 2304 4623
rect 2289 4618 2308 4619
rect 2293 4614 2294 4618
rect 2298 4614 2299 4618
rect 2303 4614 2304 4618
rect 2602 4624 2603 4628
rect 2607 4624 2608 4628
rect 2612 4624 2613 4628
rect 2598 4623 2617 4624
rect 2602 4619 2603 4623
rect 2607 4619 2608 4623
rect 2612 4619 2613 4623
rect 2598 4618 2617 4619
rect 2602 4614 2603 4618
rect 2607 4614 2608 4618
rect 2612 4614 2613 4618
rect 2911 4624 2912 4628
rect 2916 4624 2917 4628
rect 2921 4624 2922 4628
rect 2907 4623 2926 4624
rect 2911 4619 2912 4623
rect 2916 4619 2917 4623
rect 2921 4619 2922 4623
rect 2907 4618 2926 4619
rect 2911 4614 2912 4618
rect 2916 4614 2917 4618
rect 2921 4614 2922 4618
rect 1810 4613 1830 4614
rect 1675 4609 1676 4613
rect 1680 4609 1681 4613
rect 1685 4609 1686 4613
rect 1671 4608 1690 4609
rect 1675 4604 1676 4608
rect 1680 4604 1681 4608
rect 1685 4604 1686 4608
rect 1671 4603 1690 4604
rect 1675 4599 1676 4603
rect 1680 4599 1681 4603
rect 1685 4599 1686 4603
rect 1671 4598 1690 4599
rect 1675 4594 1676 4598
rect 1680 4594 1681 4598
rect 1685 4594 1686 4598
rect 1693 4611 1749 4613
rect 1693 4607 1695 4611
rect 1699 4607 1700 4611
rect 1704 4607 1705 4611
rect 1709 4607 1710 4611
rect 1714 4607 1715 4611
rect 1719 4607 1720 4611
rect 1724 4607 1725 4611
rect 1729 4607 1730 4611
rect 1734 4607 1735 4611
rect 1739 4607 1740 4611
rect 1744 4607 1745 4611
rect 1693 4606 1749 4607
rect 1693 4602 1695 4606
rect 1699 4602 1700 4606
rect 1704 4602 1705 4606
rect 1709 4602 1710 4606
rect 1714 4602 1715 4606
rect 1719 4602 1720 4606
rect 1724 4602 1725 4606
rect 1729 4602 1730 4606
rect 1734 4602 1735 4606
rect 1739 4602 1740 4606
rect 1744 4602 1745 4606
rect 1693 4601 1749 4602
rect 1693 4597 1695 4601
rect 1699 4597 1700 4601
rect 1704 4597 1705 4601
rect 1709 4597 1710 4601
rect 1714 4597 1715 4601
rect 1719 4597 1720 4601
rect 1724 4597 1725 4601
rect 1729 4597 1730 4601
rect 1734 4597 1735 4601
rect 1739 4597 1740 4601
rect 1744 4597 1745 4601
rect 1814 4609 1815 4613
rect 1819 4609 1820 4613
rect 1824 4609 1825 4613
rect 1829 4609 1830 4613
rect 1810 4608 1830 4609
rect 1814 4604 1815 4608
rect 1819 4604 1820 4608
rect 1824 4604 1825 4608
rect 1829 4604 1830 4608
rect 1810 4603 1830 4604
rect 1814 4599 1815 4603
rect 1819 4599 1820 4603
rect 1824 4599 1825 4603
rect 1829 4599 1830 4603
rect 1865 4611 1933 4614
rect 1865 4607 1867 4611
rect 1871 4607 1872 4611
rect 1876 4607 1877 4611
rect 1881 4607 1882 4611
rect 1886 4607 1887 4611
rect 1891 4607 1892 4611
rect 1896 4607 1897 4611
rect 1901 4607 1902 4611
rect 1906 4607 1907 4611
rect 1911 4607 1912 4611
rect 1916 4607 1917 4611
rect 1921 4607 1922 4611
rect 1926 4607 1927 4611
rect 1931 4607 1933 4611
rect 1865 4606 1933 4607
rect 1865 4602 1867 4606
rect 1871 4602 1872 4606
rect 1876 4602 1877 4606
rect 1881 4602 1882 4606
rect 1886 4602 1887 4606
rect 1891 4602 1892 4606
rect 1896 4602 1897 4606
rect 1901 4602 1902 4606
rect 1906 4602 1907 4606
rect 1911 4602 1912 4606
rect 1916 4602 1917 4606
rect 1921 4602 1922 4606
rect 1926 4602 1927 4606
rect 1931 4602 1933 4606
rect 1693 4596 1749 4597
rect 1693 4592 1695 4596
rect 1699 4592 1700 4596
rect 1704 4592 1705 4596
rect 1709 4592 1710 4596
rect 1714 4592 1715 4596
rect 1719 4592 1720 4596
rect 1724 4592 1725 4596
rect 1729 4592 1730 4596
rect 1734 4592 1735 4596
rect 1739 4592 1740 4596
rect 1744 4592 1745 4596
rect 1636 4578 1657 4580
rect 1640 4574 1641 4578
rect 1645 4574 1646 4578
rect 1650 4574 1651 4578
rect 1655 4574 1657 4578
rect 1636 4573 1657 4574
rect 1640 4569 1641 4573
rect 1645 4569 1646 4573
rect 1650 4569 1651 4573
rect 1655 4569 1657 4573
rect 1636 4568 1657 4569
rect 1640 4564 1641 4568
rect 1645 4564 1646 4568
rect 1650 4564 1651 4568
rect 1655 4564 1657 4568
rect 1636 4563 1657 4564
rect 1640 4559 1641 4563
rect 1645 4559 1646 4563
rect 1650 4559 1651 4563
rect 1655 4559 1657 4563
rect 1636 4558 1657 4559
rect 1640 4554 1641 4558
rect 1645 4554 1646 4558
rect 1650 4554 1651 4558
rect 1655 4554 1657 4558
rect 1636 4553 1657 4554
rect 1640 4549 1641 4553
rect 1645 4549 1646 4553
rect 1650 4549 1651 4553
rect 1655 4549 1657 4553
rect 1636 4548 1657 4549
rect 1675 4578 1676 4582
rect 1680 4578 1681 4582
rect 1685 4578 1686 4582
rect 1671 4577 1690 4578
rect 1675 4573 1676 4577
rect 1680 4573 1681 4577
rect 1685 4573 1686 4577
rect 1671 4572 1690 4573
rect 1675 4568 1676 4572
rect 1680 4568 1681 4572
rect 1685 4568 1686 4572
rect 1671 4567 1690 4568
rect 1675 4563 1676 4567
rect 1680 4563 1681 4567
rect 1685 4563 1686 4567
rect 1671 4562 1690 4563
rect 1675 4558 1676 4562
rect 1680 4558 1681 4562
rect 1685 4558 1686 4562
rect 1671 4557 1690 4558
rect 1675 4553 1676 4557
rect 1680 4553 1681 4557
rect 1685 4553 1686 4557
rect 1671 4552 1690 4553
rect 1675 4548 1676 4552
rect 1680 4548 1681 4552
rect 1685 4548 1686 4552
rect 1705 4554 1773 4557
rect 1705 4550 1707 4554
rect 1711 4550 1712 4554
rect 1716 4550 1717 4554
rect 1721 4550 1722 4554
rect 1726 4550 1727 4554
rect 1731 4550 1732 4554
rect 1736 4550 1737 4554
rect 1741 4550 1742 4554
rect 1746 4550 1747 4554
rect 1751 4550 1752 4554
rect 1756 4550 1757 4554
rect 1761 4550 1762 4554
rect 1766 4550 1767 4554
rect 1771 4550 1773 4554
rect 1705 4549 1773 4550
rect 1640 4544 1641 4548
rect 1645 4544 1646 4548
rect 1650 4544 1651 4548
rect 1655 4544 1657 4548
rect 1636 4543 1657 4544
rect 1640 4539 1641 4543
rect 1645 4539 1646 4543
rect 1650 4539 1651 4543
rect 1655 4539 1657 4543
rect 1636 4538 1657 4539
rect 1640 4534 1641 4538
rect 1645 4534 1646 4538
rect 1650 4534 1651 4538
rect 1655 4534 1657 4538
rect 1636 4533 1657 4534
rect 1640 4529 1641 4533
rect 1645 4529 1646 4533
rect 1650 4529 1651 4533
rect 1655 4529 1657 4533
rect 1636 4528 1657 4529
rect 1640 4524 1641 4528
rect 1645 4524 1646 4528
rect 1650 4524 1651 4528
rect 1655 4524 1657 4528
rect 1636 4523 1657 4524
rect 1640 4519 1641 4523
rect 1645 4519 1646 4523
rect 1650 4519 1651 4523
rect 1655 4519 1657 4523
rect 1636 4518 1657 4519
rect 1640 4514 1641 4518
rect 1645 4514 1646 4518
rect 1650 4514 1651 4518
rect 1655 4514 1657 4518
rect 1636 4512 1657 4514
rect 1705 4545 1707 4549
rect 1711 4545 1712 4549
rect 1716 4545 1717 4549
rect 1721 4545 1722 4549
rect 1726 4545 1727 4549
rect 1731 4545 1732 4549
rect 1736 4545 1737 4549
rect 1741 4545 1742 4549
rect 1746 4545 1747 4549
rect 1751 4545 1752 4549
rect 1756 4545 1757 4549
rect 1761 4545 1762 4549
rect 1766 4545 1767 4549
rect 1771 4545 1773 4549
rect 1560 4462 1563 4466
rect 1567 4462 1568 4466
rect 1572 4462 1573 4466
rect 1577 4462 1578 4466
rect 1582 4462 1583 4466
rect 1587 4462 1588 4466
rect 1592 4462 1593 4466
rect 1597 4462 1598 4466
rect 1602 4462 1603 4466
rect 1607 4462 1608 4466
rect 1612 4462 1613 4466
rect 1617 4462 1620 4466
rect 1705 4466 1773 4545
rect 1709 4462 1712 4466
rect 1716 4462 1717 4466
rect 1721 4462 1722 4466
rect 1726 4462 1727 4466
rect 1731 4462 1732 4466
rect 1736 4462 1737 4466
rect 1741 4462 1742 4466
rect 1746 4462 1747 4466
rect 1751 4462 1752 4466
rect 1756 4462 1757 4466
rect 1761 4462 1762 4466
rect 1766 4462 1769 4466
rect 1865 4466 1933 4602
rect 1980 4613 1999 4614
rect 1984 4609 1985 4613
rect 1989 4609 1990 4613
rect 1994 4609 1995 4613
rect 1980 4608 1999 4609
rect 1984 4604 1985 4608
rect 1989 4604 1990 4608
rect 1994 4604 1995 4608
rect 1980 4603 1999 4604
rect 1984 4599 1985 4603
rect 1989 4599 1990 4603
rect 1994 4599 1995 4603
rect 1980 4598 1999 4599
rect 1984 4594 1985 4598
rect 1989 4594 1990 4598
rect 1994 4594 1995 4598
rect 2002 4611 2058 4613
rect 2002 4607 2004 4611
rect 2008 4607 2009 4611
rect 2013 4607 2014 4611
rect 2018 4607 2019 4611
rect 2023 4607 2024 4611
rect 2028 4607 2029 4611
rect 2033 4607 2034 4611
rect 2038 4607 2039 4611
rect 2043 4607 2044 4611
rect 2048 4607 2049 4611
rect 2053 4607 2054 4611
rect 2002 4606 2058 4607
rect 2002 4602 2004 4606
rect 2008 4602 2009 4606
rect 2013 4602 2014 4606
rect 2018 4602 2019 4606
rect 2023 4602 2024 4606
rect 2028 4602 2029 4606
rect 2033 4602 2034 4606
rect 2038 4602 2039 4606
rect 2043 4602 2044 4606
rect 2048 4602 2049 4606
rect 2053 4602 2054 4606
rect 2002 4601 2058 4602
rect 2002 4597 2004 4601
rect 2008 4597 2009 4601
rect 2013 4597 2014 4601
rect 2018 4597 2019 4601
rect 2023 4597 2024 4601
rect 2028 4597 2029 4601
rect 2033 4597 2034 4601
rect 2038 4597 2039 4601
rect 2043 4597 2044 4601
rect 2048 4597 2049 4601
rect 2053 4597 2054 4601
rect 2002 4596 2058 4597
rect 2002 4592 2004 4596
rect 2008 4592 2009 4596
rect 2013 4592 2014 4596
rect 2018 4592 2019 4596
rect 2023 4592 2024 4596
rect 2028 4592 2029 4596
rect 2033 4592 2034 4596
rect 2038 4592 2039 4596
rect 2043 4592 2044 4596
rect 2048 4592 2049 4596
rect 2053 4592 2054 4596
rect 2174 4611 2242 4614
rect 2174 4607 2176 4611
rect 2180 4607 2181 4611
rect 2185 4607 2186 4611
rect 2190 4607 2191 4611
rect 2195 4607 2196 4611
rect 2200 4607 2201 4611
rect 2205 4607 2206 4611
rect 2210 4607 2211 4611
rect 2215 4607 2216 4611
rect 2220 4607 2221 4611
rect 2225 4607 2226 4611
rect 2230 4607 2231 4611
rect 2235 4607 2236 4611
rect 2240 4607 2242 4611
rect 2174 4606 2242 4607
rect 2174 4602 2176 4606
rect 2180 4602 2181 4606
rect 2185 4602 2186 4606
rect 2190 4602 2191 4606
rect 2195 4602 2196 4606
rect 2200 4602 2201 4606
rect 2205 4602 2206 4606
rect 2210 4602 2211 4606
rect 2215 4602 2216 4606
rect 2220 4602 2221 4606
rect 2225 4602 2226 4606
rect 2230 4602 2231 4606
rect 2235 4602 2236 4606
rect 2240 4602 2242 4606
rect 1945 4578 1966 4580
rect 1949 4574 1950 4578
rect 1954 4574 1955 4578
rect 1959 4574 1960 4578
rect 1964 4574 1966 4578
rect 1945 4573 1966 4574
rect 1949 4569 1950 4573
rect 1954 4569 1955 4573
rect 1959 4569 1960 4573
rect 1964 4569 1966 4573
rect 1945 4568 1966 4569
rect 1949 4564 1950 4568
rect 1954 4564 1955 4568
rect 1959 4564 1960 4568
rect 1964 4564 1966 4568
rect 1945 4563 1966 4564
rect 1949 4559 1950 4563
rect 1954 4559 1955 4563
rect 1959 4559 1960 4563
rect 1964 4559 1966 4563
rect 1945 4558 1966 4559
rect 1949 4554 1950 4558
rect 1954 4554 1955 4558
rect 1959 4554 1960 4558
rect 1964 4554 1966 4558
rect 1945 4553 1966 4554
rect 1949 4549 1950 4553
rect 1954 4549 1955 4553
rect 1959 4549 1960 4553
rect 1964 4549 1966 4553
rect 1945 4548 1966 4549
rect 1984 4578 1985 4582
rect 1989 4578 1990 4582
rect 1994 4578 1995 4582
rect 1980 4577 1999 4578
rect 1984 4573 1985 4577
rect 1989 4573 1990 4577
rect 1994 4573 1995 4577
rect 1980 4572 1999 4573
rect 1984 4568 1985 4572
rect 1989 4568 1990 4572
rect 1994 4568 1995 4572
rect 1980 4567 1999 4568
rect 1984 4563 1985 4567
rect 1989 4563 1990 4567
rect 1994 4563 1995 4567
rect 1980 4562 1999 4563
rect 1984 4558 1985 4562
rect 1989 4558 1990 4562
rect 1994 4558 1995 4562
rect 1980 4557 1999 4558
rect 1984 4553 1985 4557
rect 1989 4553 1990 4557
rect 1994 4553 1995 4557
rect 1980 4552 1999 4553
rect 1984 4548 1985 4552
rect 1989 4548 1990 4552
rect 1994 4548 1995 4552
rect 2014 4554 2082 4557
rect 2014 4550 2016 4554
rect 2020 4550 2021 4554
rect 2025 4550 2026 4554
rect 2030 4550 2031 4554
rect 2035 4550 2036 4554
rect 2040 4550 2041 4554
rect 2045 4550 2046 4554
rect 2050 4550 2051 4554
rect 2055 4550 2056 4554
rect 2060 4550 2061 4554
rect 2065 4550 2066 4554
rect 2070 4550 2071 4554
rect 2075 4550 2076 4554
rect 2080 4550 2082 4554
rect 2014 4549 2082 4550
rect 1949 4544 1950 4548
rect 1954 4544 1955 4548
rect 1959 4544 1960 4548
rect 1964 4544 1966 4548
rect 1945 4543 1966 4544
rect 1949 4539 1950 4543
rect 1954 4539 1955 4543
rect 1959 4539 1960 4543
rect 1964 4539 1966 4543
rect 1945 4538 1966 4539
rect 1949 4534 1950 4538
rect 1954 4534 1955 4538
rect 1959 4534 1960 4538
rect 1964 4534 1966 4538
rect 1945 4533 1966 4534
rect 1949 4529 1950 4533
rect 1954 4529 1955 4533
rect 1959 4529 1960 4533
rect 1964 4529 1966 4533
rect 1945 4528 1966 4529
rect 1949 4524 1950 4528
rect 1954 4524 1955 4528
rect 1959 4524 1960 4528
rect 1964 4524 1966 4528
rect 1945 4523 1966 4524
rect 1949 4519 1950 4523
rect 1954 4519 1955 4523
rect 1959 4519 1960 4523
rect 1964 4519 1966 4523
rect 1945 4518 1966 4519
rect 1949 4514 1950 4518
rect 1954 4514 1955 4518
rect 1959 4514 1960 4518
rect 1964 4514 1966 4518
rect 1945 4512 1966 4514
rect 2014 4545 2016 4549
rect 2020 4545 2021 4549
rect 2025 4545 2026 4549
rect 2030 4545 2031 4549
rect 2035 4545 2036 4549
rect 2040 4545 2041 4549
rect 2045 4545 2046 4549
rect 2050 4545 2051 4549
rect 2055 4545 2056 4549
rect 2060 4545 2061 4549
rect 2065 4545 2066 4549
rect 2070 4545 2071 4549
rect 2075 4545 2076 4549
rect 2080 4545 2082 4549
rect 1869 4462 1872 4466
rect 1876 4462 1877 4466
rect 1881 4462 1882 4466
rect 1886 4462 1887 4466
rect 1891 4462 1892 4466
rect 1896 4462 1897 4466
rect 1901 4462 1902 4466
rect 1906 4462 1907 4466
rect 1911 4462 1912 4466
rect 1916 4462 1917 4466
rect 1921 4462 1922 4466
rect 1926 4462 1929 4466
rect 2014 4466 2082 4545
rect 2096 4519 2100 4531
rect 2096 4503 2100 4515
rect 2096 4487 2100 4499
rect 2154 4519 2158 4531
rect 2154 4503 2158 4515
rect 2154 4487 2158 4499
rect 2018 4462 2021 4466
rect 2025 4462 2026 4466
rect 2030 4462 2031 4466
rect 2035 4462 2036 4466
rect 2040 4462 2041 4466
rect 2045 4462 2046 4466
rect 2050 4462 2051 4466
rect 2055 4462 2056 4466
rect 2060 4462 2061 4466
rect 2065 4462 2066 4466
rect 2070 4462 2071 4466
rect 2075 4462 2078 4466
rect 2174 4466 2242 4602
rect 2289 4613 2308 4614
rect 2293 4609 2294 4613
rect 2298 4609 2299 4613
rect 2303 4609 2304 4613
rect 2289 4608 2308 4609
rect 2293 4604 2294 4608
rect 2298 4604 2299 4608
rect 2303 4604 2304 4608
rect 2289 4603 2308 4604
rect 2293 4599 2294 4603
rect 2298 4599 2299 4603
rect 2303 4599 2304 4603
rect 2289 4598 2308 4599
rect 2293 4594 2294 4598
rect 2298 4594 2299 4598
rect 2303 4594 2304 4598
rect 2311 4611 2367 4613
rect 2311 4607 2313 4611
rect 2317 4607 2318 4611
rect 2322 4607 2323 4611
rect 2327 4607 2328 4611
rect 2332 4607 2333 4611
rect 2337 4607 2338 4611
rect 2342 4607 2343 4611
rect 2347 4607 2348 4611
rect 2352 4607 2353 4611
rect 2357 4607 2358 4611
rect 2362 4607 2363 4611
rect 2311 4606 2367 4607
rect 2311 4602 2313 4606
rect 2317 4602 2318 4606
rect 2322 4602 2323 4606
rect 2327 4602 2328 4606
rect 2332 4602 2333 4606
rect 2337 4602 2338 4606
rect 2342 4602 2343 4606
rect 2347 4602 2348 4606
rect 2352 4602 2353 4606
rect 2357 4602 2358 4606
rect 2362 4602 2363 4606
rect 2311 4601 2367 4602
rect 2311 4597 2313 4601
rect 2317 4597 2318 4601
rect 2322 4597 2323 4601
rect 2327 4597 2328 4601
rect 2332 4597 2333 4601
rect 2337 4597 2338 4601
rect 2342 4597 2343 4601
rect 2347 4597 2348 4601
rect 2352 4597 2353 4601
rect 2357 4597 2358 4601
rect 2362 4597 2363 4601
rect 2311 4596 2367 4597
rect 2311 4592 2313 4596
rect 2317 4592 2318 4596
rect 2322 4592 2323 4596
rect 2327 4592 2328 4596
rect 2332 4592 2333 4596
rect 2337 4592 2338 4596
rect 2342 4592 2343 4596
rect 2347 4592 2348 4596
rect 2352 4592 2353 4596
rect 2357 4592 2358 4596
rect 2362 4592 2363 4596
rect 2483 4611 2551 4614
rect 2483 4607 2485 4611
rect 2489 4607 2490 4611
rect 2494 4607 2495 4611
rect 2499 4607 2500 4611
rect 2504 4607 2505 4611
rect 2509 4607 2510 4611
rect 2514 4607 2515 4611
rect 2519 4607 2520 4611
rect 2524 4607 2525 4611
rect 2529 4607 2530 4611
rect 2534 4607 2535 4611
rect 2539 4607 2540 4611
rect 2544 4607 2545 4611
rect 2549 4607 2551 4611
rect 2483 4606 2551 4607
rect 2483 4602 2485 4606
rect 2489 4602 2490 4606
rect 2494 4602 2495 4606
rect 2499 4602 2500 4606
rect 2504 4602 2505 4606
rect 2509 4602 2510 4606
rect 2514 4602 2515 4606
rect 2519 4602 2520 4606
rect 2524 4602 2525 4606
rect 2529 4602 2530 4606
rect 2534 4602 2535 4606
rect 2539 4602 2540 4606
rect 2544 4602 2545 4606
rect 2549 4602 2551 4606
rect 2254 4578 2275 4580
rect 2258 4574 2259 4578
rect 2263 4574 2264 4578
rect 2268 4574 2269 4578
rect 2273 4574 2275 4578
rect 2254 4573 2275 4574
rect 2258 4569 2259 4573
rect 2263 4569 2264 4573
rect 2268 4569 2269 4573
rect 2273 4569 2275 4573
rect 2254 4568 2275 4569
rect 2258 4564 2259 4568
rect 2263 4564 2264 4568
rect 2268 4564 2269 4568
rect 2273 4564 2275 4568
rect 2254 4563 2275 4564
rect 2258 4559 2259 4563
rect 2263 4559 2264 4563
rect 2268 4559 2269 4563
rect 2273 4559 2275 4563
rect 2254 4558 2275 4559
rect 2258 4554 2259 4558
rect 2263 4554 2264 4558
rect 2268 4554 2269 4558
rect 2273 4554 2275 4558
rect 2254 4553 2275 4554
rect 2258 4549 2259 4553
rect 2263 4549 2264 4553
rect 2268 4549 2269 4553
rect 2273 4549 2275 4553
rect 2254 4548 2275 4549
rect 2293 4578 2294 4582
rect 2298 4578 2299 4582
rect 2303 4578 2304 4582
rect 2289 4577 2308 4578
rect 2293 4573 2294 4577
rect 2298 4573 2299 4577
rect 2303 4573 2304 4577
rect 2289 4572 2308 4573
rect 2293 4568 2294 4572
rect 2298 4568 2299 4572
rect 2303 4568 2304 4572
rect 2289 4567 2308 4568
rect 2293 4563 2294 4567
rect 2298 4563 2299 4567
rect 2303 4563 2304 4567
rect 2289 4562 2308 4563
rect 2293 4558 2294 4562
rect 2298 4558 2299 4562
rect 2303 4558 2304 4562
rect 2289 4557 2308 4558
rect 2293 4553 2294 4557
rect 2298 4553 2299 4557
rect 2303 4553 2304 4557
rect 2289 4552 2308 4553
rect 2293 4548 2294 4552
rect 2298 4548 2299 4552
rect 2303 4548 2304 4552
rect 2323 4554 2391 4557
rect 2323 4550 2325 4554
rect 2329 4550 2330 4554
rect 2334 4550 2335 4554
rect 2339 4550 2340 4554
rect 2344 4550 2345 4554
rect 2349 4550 2350 4554
rect 2354 4550 2355 4554
rect 2359 4550 2360 4554
rect 2364 4550 2365 4554
rect 2369 4550 2370 4554
rect 2374 4550 2375 4554
rect 2379 4550 2380 4554
rect 2384 4550 2385 4554
rect 2389 4550 2391 4554
rect 2323 4549 2391 4550
rect 2258 4544 2259 4548
rect 2263 4544 2264 4548
rect 2268 4544 2269 4548
rect 2273 4544 2275 4548
rect 2254 4543 2275 4544
rect 2258 4539 2259 4543
rect 2263 4539 2264 4543
rect 2268 4539 2269 4543
rect 2273 4539 2275 4543
rect 2254 4538 2275 4539
rect 2258 4534 2259 4538
rect 2263 4534 2264 4538
rect 2268 4534 2269 4538
rect 2273 4534 2275 4538
rect 2254 4533 2275 4534
rect 2258 4529 2259 4533
rect 2263 4529 2264 4533
rect 2268 4529 2269 4533
rect 2273 4529 2275 4533
rect 2254 4528 2275 4529
rect 2258 4524 2259 4528
rect 2263 4524 2264 4528
rect 2268 4524 2269 4528
rect 2273 4524 2275 4528
rect 2254 4523 2275 4524
rect 2258 4519 2259 4523
rect 2263 4519 2264 4523
rect 2268 4519 2269 4523
rect 2273 4519 2275 4523
rect 2254 4518 2275 4519
rect 2258 4514 2259 4518
rect 2263 4514 2264 4518
rect 2268 4514 2269 4518
rect 2273 4514 2275 4518
rect 2254 4512 2275 4514
rect 2323 4545 2325 4549
rect 2329 4545 2330 4549
rect 2334 4545 2335 4549
rect 2339 4545 2340 4549
rect 2344 4545 2345 4549
rect 2349 4545 2350 4549
rect 2354 4545 2355 4549
rect 2359 4545 2360 4549
rect 2364 4545 2365 4549
rect 2369 4545 2370 4549
rect 2374 4545 2375 4549
rect 2379 4545 2380 4549
rect 2384 4545 2385 4549
rect 2389 4545 2391 4549
rect 2178 4462 2181 4466
rect 2185 4462 2186 4466
rect 2190 4462 2191 4466
rect 2195 4462 2196 4466
rect 2200 4462 2201 4466
rect 2205 4462 2206 4466
rect 2210 4462 2211 4466
rect 2215 4462 2216 4466
rect 2220 4462 2221 4466
rect 2225 4462 2226 4466
rect 2230 4462 2231 4466
rect 2235 4462 2238 4466
rect 2323 4466 2391 4545
rect 2405 4519 2409 4531
rect 2405 4503 2409 4515
rect 2405 4487 2409 4499
rect 2463 4519 2467 4531
rect 2463 4503 2467 4515
rect 2463 4487 2467 4499
rect 2327 4462 2330 4466
rect 2334 4462 2335 4466
rect 2339 4462 2340 4466
rect 2344 4462 2345 4466
rect 2349 4462 2350 4466
rect 2354 4462 2355 4466
rect 2359 4462 2360 4466
rect 2364 4462 2365 4466
rect 2369 4462 2370 4466
rect 2374 4462 2375 4466
rect 2379 4462 2380 4466
rect 2384 4462 2387 4466
rect 2483 4466 2551 4602
rect 2598 4613 2617 4614
rect 2602 4609 2603 4613
rect 2607 4609 2608 4613
rect 2612 4609 2613 4613
rect 2598 4608 2617 4609
rect 2602 4604 2603 4608
rect 2607 4604 2608 4608
rect 2612 4604 2613 4608
rect 2598 4603 2617 4604
rect 2602 4599 2603 4603
rect 2607 4599 2608 4603
rect 2612 4599 2613 4603
rect 2598 4598 2617 4599
rect 2602 4594 2603 4598
rect 2607 4594 2608 4598
rect 2612 4594 2613 4598
rect 2620 4611 2676 4613
rect 2620 4607 2622 4611
rect 2626 4607 2627 4611
rect 2631 4607 2632 4611
rect 2636 4607 2637 4611
rect 2641 4607 2642 4611
rect 2646 4607 2647 4611
rect 2651 4607 2652 4611
rect 2656 4607 2657 4611
rect 2661 4607 2662 4611
rect 2666 4607 2667 4611
rect 2671 4607 2672 4611
rect 2620 4606 2676 4607
rect 2620 4602 2622 4606
rect 2626 4602 2627 4606
rect 2631 4602 2632 4606
rect 2636 4602 2637 4606
rect 2641 4602 2642 4606
rect 2646 4602 2647 4606
rect 2651 4602 2652 4606
rect 2656 4602 2657 4606
rect 2661 4602 2662 4606
rect 2666 4602 2667 4606
rect 2671 4602 2672 4606
rect 2620 4601 2676 4602
rect 2620 4597 2622 4601
rect 2626 4597 2627 4601
rect 2631 4597 2632 4601
rect 2636 4597 2637 4601
rect 2641 4597 2642 4601
rect 2646 4597 2647 4601
rect 2651 4597 2652 4601
rect 2656 4597 2657 4601
rect 2661 4597 2662 4601
rect 2666 4597 2667 4601
rect 2671 4597 2672 4601
rect 2620 4596 2676 4597
rect 2620 4592 2622 4596
rect 2626 4592 2627 4596
rect 2631 4592 2632 4596
rect 2636 4592 2637 4596
rect 2641 4592 2642 4596
rect 2646 4592 2647 4596
rect 2651 4592 2652 4596
rect 2656 4592 2657 4596
rect 2661 4592 2662 4596
rect 2666 4592 2667 4596
rect 2671 4592 2672 4596
rect 2792 4611 2860 4614
rect 2792 4607 2794 4611
rect 2798 4607 2799 4611
rect 2803 4607 2804 4611
rect 2808 4607 2809 4611
rect 2813 4607 2814 4611
rect 2818 4607 2819 4611
rect 2823 4607 2824 4611
rect 2828 4607 2829 4611
rect 2833 4607 2834 4611
rect 2838 4607 2839 4611
rect 2843 4607 2844 4611
rect 2848 4607 2849 4611
rect 2853 4607 2854 4611
rect 2858 4607 2860 4611
rect 2792 4606 2860 4607
rect 2792 4602 2794 4606
rect 2798 4602 2799 4606
rect 2803 4602 2804 4606
rect 2808 4602 2809 4606
rect 2813 4602 2814 4606
rect 2818 4602 2819 4606
rect 2823 4602 2824 4606
rect 2828 4602 2829 4606
rect 2833 4602 2834 4606
rect 2838 4602 2839 4606
rect 2843 4602 2844 4606
rect 2848 4602 2849 4606
rect 2853 4602 2854 4606
rect 2858 4602 2860 4606
rect 2563 4578 2584 4580
rect 2567 4574 2568 4578
rect 2572 4574 2573 4578
rect 2577 4574 2578 4578
rect 2582 4574 2584 4578
rect 2563 4573 2584 4574
rect 2567 4569 2568 4573
rect 2572 4569 2573 4573
rect 2577 4569 2578 4573
rect 2582 4569 2584 4573
rect 2563 4568 2584 4569
rect 2567 4564 2568 4568
rect 2572 4564 2573 4568
rect 2577 4564 2578 4568
rect 2582 4564 2584 4568
rect 2563 4563 2584 4564
rect 2567 4559 2568 4563
rect 2572 4559 2573 4563
rect 2577 4559 2578 4563
rect 2582 4559 2584 4563
rect 2563 4558 2584 4559
rect 2567 4554 2568 4558
rect 2572 4554 2573 4558
rect 2577 4554 2578 4558
rect 2582 4554 2584 4558
rect 2563 4553 2584 4554
rect 2567 4549 2568 4553
rect 2572 4549 2573 4553
rect 2577 4549 2578 4553
rect 2582 4549 2584 4553
rect 2563 4548 2584 4549
rect 2602 4578 2603 4582
rect 2607 4578 2608 4582
rect 2612 4578 2613 4582
rect 2598 4577 2617 4578
rect 2602 4573 2603 4577
rect 2607 4573 2608 4577
rect 2612 4573 2613 4577
rect 2598 4572 2617 4573
rect 2602 4568 2603 4572
rect 2607 4568 2608 4572
rect 2612 4568 2613 4572
rect 2598 4567 2617 4568
rect 2602 4563 2603 4567
rect 2607 4563 2608 4567
rect 2612 4563 2613 4567
rect 2598 4562 2617 4563
rect 2602 4558 2603 4562
rect 2607 4558 2608 4562
rect 2612 4558 2613 4562
rect 2598 4557 2617 4558
rect 2602 4553 2603 4557
rect 2607 4553 2608 4557
rect 2612 4553 2613 4557
rect 2598 4552 2617 4553
rect 2602 4548 2603 4552
rect 2607 4548 2608 4552
rect 2612 4548 2613 4552
rect 2632 4554 2700 4557
rect 2632 4550 2634 4554
rect 2638 4550 2639 4554
rect 2643 4550 2644 4554
rect 2648 4550 2649 4554
rect 2653 4550 2654 4554
rect 2658 4550 2659 4554
rect 2663 4550 2664 4554
rect 2668 4550 2669 4554
rect 2673 4550 2674 4554
rect 2678 4550 2679 4554
rect 2683 4550 2684 4554
rect 2688 4550 2689 4554
rect 2693 4550 2694 4554
rect 2698 4550 2700 4554
rect 2632 4549 2700 4550
rect 2567 4544 2568 4548
rect 2572 4544 2573 4548
rect 2577 4544 2578 4548
rect 2582 4544 2584 4548
rect 2563 4543 2584 4544
rect 2567 4539 2568 4543
rect 2572 4539 2573 4543
rect 2577 4539 2578 4543
rect 2582 4539 2584 4543
rect 2563 4538 2584 4539
rect 2567 4534 2568 4538
rect 2572 4534 2573 4538
rect 2577 4534 2578 4538
rect 2582 4534 2584 4538
rect 2563 4533 2584 4534
rect 2567 4529 2568 4533
rect 2572 4529 2573 4533
rect 2577 4529 2578 4533
rect 2582 4529 2584 4533
rect 2563 4528 2584 4529
rect 2567 4524 2568 4528
rect 2572 4524 2573 4528
rect 2577 4524 2578 4528
rect 2582 4524 2584 4528
rect 2563 4523 2584 4524
rect 2567 4519 2568 4523
rect 2572 4519 2573 4523
rect 2577 4519 2578 4523
rect 2582 4519 2584 4523
rect 2563 4518 2584 4519
rect 2567 4514 2568 4518
rect 2572 4514 2573 4518
rect 2577 4514 2578 4518
rect 2582 4514 2584 4518
rect 2563 4512 2584 4514
rect 2632 4545 2634 4549
rect 2638 4545 2639 4549
rect 2643 4545 2644 4549
rect 2648 4545 2649 4549
rect 2653 4545 2654 4549
rect 2658 4545 2659 4549
rect 2663 4545 2664 4549
rect 2668 4545 2669 4549
rect 2673 4545 2674 4549
rect 2678 4545 2679 4549
rect 2683 4545 2684 4549
rect 2688 4545 2689 4549
rect 2693 4545 2694 4549
rect 2698 4545 2700 4549
rect 2487 4462 2490 4466
rect 2494 4462 2495 4466
rect 2499 4462 2500 4466
rect 2504 4462 2505 4466
rect 2509 4462 2510 4466
rect 2514 4462 2515 4466
rect 2519 4462 2520 4466
rect 2524 4462 2525 4466
rect 2529 4462 2530 4466
rect 2534 4462 2535 4466
rect 2539 4462 2540 4466
rect 2544 4462 2547 4466
rect 2632 4466 2700 4545
rect 2714 4519 2718 4531
rect 2714 4503 2718 4515
rect 2714 4487 2718 4499
rect 2772 4519 2776 4531
rect 2772 4503 2776 4515
rect 2772 4487 2776 4499
rect 2636 4462 2639 4466
rect 2643 4462 2644 4466
rect 2648 4462 2649 4466
rect 2653 4462 2654 4466
rect 2658 4462 2659 4466
rect 2663 4462 2664 4466
rect 2668 4462 2669 4466
rect 2673 4462 2674 4466
rect 2678 4462 2679 4466
rect 2683 4462 2684 4466
rect 2688 4462 2689 4466
rect 2693 4462 2696 4466
rect 2792 4466 2860 4602
rect 2907 4613 2926 4614
rect 2911 4609 2912 4613
rect 2916 4609 2917 4613
rect 2921 4609 2922 4613
rect 2907 4608 2926 4609
rect 2911 4604 2912 4608
rect 2916 4604 2917 4608
rect 2921 4604 2922 4608
rect 2907 4603 2926 4604
rect 2911 4599 2912 4603
rect 2916 4599 2917 4603
rect 2921 4599 2922 4603
rect 2907 4598 2926 4599
rect 2911 4594 2912 4598
rect 2916 4594 2917 4598
rect 2921 4594 2922 4598
rect 2929 4611 2985 4613
rect 2929 4607 2931 4611
rect 2935 4607 2936 4611
rect 2940 4607 2941 4611
rect 2945 4607 2946 4611
rect 2950 4607 2951 4611
rect 2955 4607 2956 4611
rect 2960 4607 2961 4611
rect 2965 4607 2966 4611
rect 2970 4607 2971 4611
rect 2975 4607 2976 4611
rect 2980 4607 2981 4611
rect 2929 4606 2985 4607
rect 2929 4602 2931 4606
rect 2935 4602 2936 4606
rect 2940 4602 2941 4606
rect 2945 4602 2946 4606
rect 2950 4602 2951 4606
rect 2955 4602 2956 4606
rect 2960 4602 2961 4606
rect 2965 4602 2966 4606
rect 2970 4602 2971 4606
rect 2975 4602 2976 4606
rect 2980 4602 2981 4606
rect 2929 4601 2985 4602
rect 2929 4597 2931 4601
rect 2935 4597 2936 4601
rect 2940 4597 2941 4601
rect 2945 4597 2946 4601
rect 2950 4597 2951 4601
rect 2955 4597 2956 4601
rect 2960 4597 2961 4601
rect 2965 4597 2966 4601
rect 2970 4597 2971 4601
rect 2975 4597 2976 4601
rect 2980 4597 2981 4601
rect 2929 4596 2985 4597
rect 2929 4592 2931 4596
rect 2935 4592 2936 4596
rect 2940 4592 2941 4596
rect 2945 4592 2946 4596
rect 2950 4592 2951 4596
rect 2955 4592 2956 4596
rect 2960 4592 2961 4596
rect 2965 4592 2966 4596
rect 2970 4592 2971 4596
rect 2975 4592 2976 4596
rect 2980 4592 2981 4596
rect 2872 4578 2893 4580
rect 2876 4574 2877 4578
rect 2881 4574 2882 4578
rect 2886 4574 2887 4578
rect 2891 4574 2893 4578
rect 2872 4573 2893 4574
rect 2876 4569 2877 4573
rect 2881 4569 2882 4573
rect 2886 4569 2887 4573
rect 2891 4569 2893 4573
rect 2872 4568 2893 4569
rect 2876 4564 2877 4568
rect 2881 4564 2882 4568
rect 2886 4564 2887 4568
rect 2891 4564 2893 4568
rect 2872 4563 2893 4564
rect 2876 4559 2877 4563
rect 2881 4559 2882 4563
rect 2886 4559 2887 4563
rect 2891 4559 2893 4563
rect 2872 4558 2893 4559
rect 2876 4554 2877 4558
rect 2881 4554 2882 4558
rect 2886 4554 2887 4558
rect 2891 4554 2893 4558
rect 2872 4553 2893 4554
rect 2876 4549 2877 4553
rect 2881 4549 2882 4553
rect 2886 4549 2887 4553
rect 2891 4549 2893 4553
rect 2872 4548 2893 4549
rect 2911 4578 2912 4582
rect 2916 4578 2917 4582
rect 2921 4578 2922 4582
rect 2907 4577 2926 4578
rect 2911 4573 2912 4577
rect 2916 4573 2917 4577
rect 2921 4573 2922 4577
rect 2907 4572 2926 4573
rect 2911 4568 2912 4572
rect 2916 4568 2917 4572
rect 2921 4568 2922 4572
rect 2998 4578 3006 4691
rect 3664 4653 3684 4655
rect 3668 4649 3669 4653
rect 3673 4649 3674 4653
rect 3678 4649 3679 4653
rect 3683 4649 3684 4653
rect 3664 4648 3684 4649
rect 3668 4644 3669 4648
rect 3673 4644 3674 4648
rect 3678 4644 3679 4648
rect 3683 4644 3684 4648
rect 3664 4643 3684 4644
rect 3668 4639 3669 4643
rect 3673 4639 3674 4643
rect 3678 4639 3679 4643
rect 3683 4639 3684 4643
rect 3664 4638 3684 4639
rect 3668 4634 3669 4638
rect 3673 4634 3674 4638
rect 3678 4634 3679 4638
rect 3683 4634 3684 4638
rect 3664 4633 3684 4634
rect 3668 4629 3669 4633
rect 3673 4629 3674 4633
rect 3678 4629 3679 4633
rect 3683 4629 3684 4633
rect 3664 4628 3684 4629
rect 3220 4624 3221 4628
rect 3225 4624 3226 4628
rect 3230 4624 3231 4628
rect 3216 4623 3235 4624
rect 3220 4619 3221 4623
rect 3225 4619 3226 4623
rect 3230 4619 3231 4623
rect 3216 4618 3235 4619
rect 3220 4614 3221 4618
rect 3225 4614 3226 4618
rect 3230 4614 3231 4618
rect 3529 4624 3530 4628
rect 3534 4624 3535 4628
rect 3539 4624 3540 4628
rect 3525 4623 3544 4624
rect 3529 4619 3530 4623
rect 3534 4619 3535 4623
rect 3539 4619 3540 4623
rect 3525 4618 3544 4619
rect 3529 4614 3530 4618
rect 3534 4614 3535 4618
rect 3539 4614 3540 4618
rect 2998 4573 3000 4578
rect 3005 4573 3006 4578
rect 2998 4571 3006 4573
rect 3101 4611 3169 4614
rect 3101 4607 3103 4611
rect 3107 4607 3108 4611
rect 3112 4607 3113 4611
rect 3117 4607 3118 4611
rect 3122 4607 3123 4611
rect 3127 4607 3128 4611
rect 3132 4607 3133 4611
rect 3137 4607 3138 4611
rect 3142 4607 3143 4611
rect 3147 4607 3148 4611
rect 3152 4607 3153 4611
rect 3157 4607 3158 4611
rect 3162 4607 3163 4611
rect 3167 4607 3169 4611
rect 3101 4606 3169 4607
rect 3101 4602 3103 4606
rect 3107 4602 3108 4606
rect 3112 4602 3113 4606
rect 3117 4602 3118 4606
rect 3122 4602 3123 4606
rect 3127 4602 3128 4606
rect 3132 4602 3133 4606
rect 3137 4602 3138 4606
rect 3142 4602 3143 4606
rect 3147 4602 3148 4606
rect 3152 4602 3153 4606
rect 3157 4602 3158 4606
rect 3162 4602 3163 4606
rect 3167 4602 3169 4606
rect 2907 4567 2926 4568
rect 2911 4563 2912 4567
rect 2916 4563 2917 4567
rect 2921 4563 2922 4567
rect 2907 4562 2926 4563
rect 2911 4558 2912 4562
rect 2916 4558 2917 4562
rect 2921 4558 2922 4562
rect 2907 4557 2926 4558
rect 2911 4553 2912 4557
rect 2916 4553 2917 4557
rect 2921 4553 2922 4557
rect 2907 4552 2926 4553
rect 2911 4548 2912 4552
rect 2916 4548 2917 4552
rect 2921 4548 2922 4552
rect 2941 4554 3009 4557
rect 2941 4550 2943 4554
rect 2947 4550 2948 4554
rect 2952 4550 2953 4554
rect 2957 4550 2958 4554
rect 2962 4550 2963 4554
rect 2967 4550 2968 4554
rect 2972 4550 2973 4554
rect 2977 4550 2978 4554
rect 2982 4550 2983 4554
rect 2987 4550 2988 4554
rect 2992 4550 2993 4554
rect 2997 4550 2998 4554
rect 3002 4550 3003 4554
rect 3007 4550 3009 4554
rect 2941 4549 3009 4550
rect 2876 4544 2877 4548
rect 2881 4544 2882 4548
rect 2886 4544 2887 4548
rect 2891 4544 2893 4548
rect 2872 4543 2893 4544
rect 2876 4539 2877 4543
rect 2881 4539 2882 4543
rect 2886 4539 2887 4543
rect 2891 4539 2893 4543
rect 2872 4538 2893 4539
rect 2876 4534 2877 4538
rect 2881 4534 2882 4538
rect 2886 4534 2887 4538
rect 2891 4534 2893 4538
rect 2872 4533 2893 4534
rect 2876 4529 2877 4533
rect 2881 4529 2882 4533
rect 2886 4529 2887 4533
rect 2891 4529 2893 4533
rect 2872 4528 2893 4529
rect 2876 4524 2877 4528
rect 2881 4524 2882 4528
rect 2886 4524 2887 4528
rect 2891 4524 2893 4528
rect 2872 4523 2893 4524
rect 2876 4519 2877 4523
rect 2881 4519 2882 4523
rect 2886 4519 2887 4523
rect 2891 4519 2893 4523
rect 2872 4518 2893 4519
rect 2876 4514 2877 4518
rect 2881 4514 2882 4518
rect 2886 4514 2887 4518
rect 2891 4514 2893 4518
rect 2872 4512 2893 4514
rect 2941 4545 2943 4549
rect 2947 4545 2948 4549
rect 2952 4545 2953 4549
rect 2957 4545 2958 4549
rect 2962 4545 2963 4549
rect 2967 4545 2968 4549
rect 2972 4545 2973 4549
rect 2977 4545 2978 4549
rect 2982 4545 2983 4549
rect 2987 4545 2988 4549
rect 2992 4545 2993 4549
rect 2997 4545 2998 4549
rect 3002 4545 3003 4549
rect 3007 4545 3009 4549
rect 2796 4462 2799 4466
rect 2803 4462 2804 4466
rect 2808 4462 2809 4466
rect 2813 4462 2814 4466
rect 2818 4462 2819 4466
rect 2823 4462 2824 4466
rect 2828 4462 2829 4466
rect 2833 4462 2834 4466
rect 2838 4462 2839 4466
rect 2843 4462 2844 4466
rect 2848 4462 2849 4466
rect 2853 4462 2856 4466
rect 2941 4466 3009 4545
rect 3023 4519 3027 4531
rect 3023 4503 3027 4515
rect 3023 4487 3027 4499
rect 3081 4519 3085 4531
rect 3081 4503 3085 4515
rect 3081 4487 3085 4499
rect 2945 4462 2948 4466
rect 2952 4462 2953 4466
rect 2957 4462 2958 4466
rect 2962 4462 2963 4466
rect 2967 4462 2968 4466
rect 2972 4462 2973 4466
rect 2977 4462 2978 4466
rect 2982 4462 2983 4466
rect 2987 4462 2988 4466
rect 2992 4462 2993 4466
rect 2997 4462 2998 4466
rect 3002 4462 3005 4466
rect 3101 4466 3169 4602
rect 3216 4613 3235 4614
rect 3220 4609 3221 4613
rect 3225 4609 3226 4613
rect 3230 4609 3231 4613
rect 3216 4608 3235 4609
rect 3220 4604 3221 4608
rect 3225 4604 3226 4608
rect 3230 4604 3231 4608
rect 3216 4603 3235 4604
rect 3220 4599 3221 4603
rect 3225 4599 3226 4603
rect 3230 4599 3231 4603
rect 3216 4598 3235 4599
rect 3220 4594 3221 4598
rect 3225 4594 3226 4598
rect 3230 4594 3231 4598
rect 3238 4611 3294 4613
rect 3238 4607 3240 4611
rect 3244 4607 3245 4611
rect 3249 4607 3250 4611
rect 3254 4607 3255 4611
rect 3259 4607 3260 4611
rect 3264 4607 3265 4611
rect 3269 4607 3270 4611
rect 3274 4607 3275 4611
rect 3279 4607 3280 4611
rect 3284 4607 3285 4611
rect 3289 4607 3290 4611
rect 3238 4606 3294 4607
rect 3238 4602 3240 4606
rect 3244 4602 3245 4606
rect 3249 4602 3250 4606
rect 3254 4602 3255 4606
rect 3259 4602 3260 4606
rect 3264 4602 3265 4606
rect 3269 4602 3270 4606
rect 3274 4602 3275 4606
rect 3279 4602 3280 4606
rect 3284 4602 3285 4606
rect 3289 4602 3290 4606
rect 3238 4601 3294 4602
rect 3238 4597 3240 4601
rect 3244 4597 3245 4601
rect 3249 4597 3250 4601
rect 3254 4597 3255 4601
rect 3259 4597 3260 4601
rect 3264 4597 3265 4601
rect 3269 4597 3270 4601
rect 3274 4597 3275 4601
rect 3279 4597 3280 4601
rect 3284 4597 3285 4601
rect 3289 4597 3290 4601
rect 3238 4596 3294 4597
rect 3238 4592 3240 4596
rect 3244 4592 3245 4596
rect 3249 4592 3250 4596
rect 3254 4592 3255 4596
rect 3259 4592 3260 4596
rect 3264 4592 3265 4596
rect 3269 4592 3270 4596
rect 3274 4592 3275 4596
rect 3279 4592 3280 4596
rect 3284 4592 3285 4596
rect 3289 4592 3290 4596
rect 3410 4611 3478 4614
rect 3410 4607 3412 4611
rect 3416 4607 3417 4611
rect 3421 4607 3422 4611
rect 3426 4607 3427 4611
rect 3431 4607 3432 4611
rect 3436 4607 3437 4611
rect 3441 4607 3442 4611
rect 3446 4607 3447 4611
rect 3451 4607 3452 4611
rect 3456 4607 3457 4611
rect 3461 4607 3462 4611
rect 3466 4607 3467 4611
rect 3471 4607 3472 4611
rect 3476 4607 3478 4611
rect 3410 4606 3478 4607
rect 3410 4602 3412 4606
rect 3416 4602 3417 4606
rect 3421 4602 3422 4606
rect 3426 4602 3427 4606
rect 3431 4602 3432 4606
rect 3436 4602 3437 4606
rect 3441 4602 3442 4606
rect 3446 4602 3447 4606
rect 3451 4602 3452 4606
rect 3456 4602 3457 4606
rect 3461 4602 3462 4606
rect 3466 4602 3467 4606
rect 3471 4602 3472 4606
rect 3476 4602 3478 4606
rect 3181 4578 3202 4580
rect 3185 4574 3186 4578
rect 3190 4574 3191 4578
rect 3195 4574 3196 4578
rect 3200 4574 3202 4578
rect 3181 4573 3202 4574
rect 3185 4569 3186 4573
rect 3190 4569 3191 4573
rect 3195 4569 3196 4573
rect 3200 4569 3202 4573
rect 3181 4568 3202 4569
rect 3185 4564 3186 4568
rect 3190 4564 3191 4568
rect 3195 4564 3196 4568
rect 3200 4564 3202 4568
rect 3181 4563 3202 4564
rect 3185 4559 3186 4563
rect 3190 4559 3191 4563
rect 3195 4559 3196 4563
rect 3200 4559 3202 4563
rect 3181 4558 3202 4559
rect 3185 4554 3186 4558
rect 3190 4554 3191 4558
rect 3195 4554 3196 4558
rect 3200 4554 3202 4558
rect 3181 4553 3202 4554
rect 3185 4549 3186 4553
rect 3190 4549 3191 4553
rect 3195 4549 3196 4553
rect 3200 4549 3202 4553
rect 3181 4548 3202 4549
rect 3220 4578 3221 4582
rect 3225 4578 3226 4582
rect 3230 4578 3231 4582
rect 3216 4577 3235 4578
rect 3220 4573 3221 4577
rect 3225 4573 3226 4577
rect 3230 4573 3231 4577
rect 3216 4572 3235 4573
rect 3220 4568 3221 4572
rect 3225 4568 3226 4572
rect 3230 4568 3231 4572
rect 3216 4567 3235 4568
rect 3220 4563 3221 4567
rect 3225 4563 3226 4567
rect 3230 4563 3231 4567
rect 3216 4562 3235 4563
rect 3220 4558 3221 4562
rect 3225 4558 3226 4562
rect 3230 4558 3231 4562
rect 3216 4557 3235 4558
rect 3220 4553 3221 4557
rect 3225 4553 3226 4557
rect 3230 4553 3231 4557
rect 3216 4552 3235 4553
rect 3220 4548 3221 4552
rect 3225 4548 3226 4552
rect 3230 4548 3231 4552
rect 3250 4554 3318 4557
rect 3250 4550 3252 4554
rect 3256 4550 3257 4554
rect 3261 4550 3262 4554
rect 3266 4550 3267 4554
rect 3271 4550 3272 4554
rect 3276 4550 3277 4554
rect 3281 4550 3282 4554
rect 3286 4550 3287 4554
rect 3291 4550 3292 4554
rect 3296 4550 3297 4554
rect 3301 4550 3302 4554
rect 3306 4550 3307 4554
rect 3311 4550 3312 4554
rect 3316 4550 3318 4554
rect 3250 4549 3318 4550
rect 3185 4544 3186 4548
rect 3190 4544 3191 4548
rect 3195 4544 3196 4548
rect 3200 4544 3202 4548
rect 3181 4543 3202 4544
rect 3185 4539 3186 4543
rect 3190 4539 3191 4543
rect 3195 4539 3196 4543
rect 3200 4539 3202 4543
rect 3181 4538 3202 4539
rect 3185 4534 3186 4538
rect 3190 4534 3191 4538
rect 3195 4534 3196 4538
rect 3200 4534 3202 4538
rect 3181 4533 3202 4534
rect 3185 4529 3186 4533
rect 3190 4529 3191 4533
rect 3195 4529 3196 4533
rect 3200 4529 3202 4533
rect 3181 4528 3202 4529
rect 3185 4524 3186 4528
rect 3190 4524 3191 4528
rect 3195 4524 3196 4528
rect 3200 4524 3202 4528
rect 3181 4523 3202 4524
rect 3185 4519 3186 4523
rect 3190 4519 3191 4523
rect 3195 4519 3196 4523
rect 3200 4519 3202 4523
rect 3181 4518 3202 4519
rect 3185 4514 3186 4518
rect 3190 4514 3191 4518
rect 3195 4514 3196 4518
rect 3200 4514 3202 4518
rect 3181 4512 3202 4514
rect 3250 4545 3252 4549
rect 3256 4545 3257 4549
rect 3261 4545 3262 4549
rect 3266 4545 3267 4549
rect 3271 4545 3272 4549
rect 3276 4545 3277 4549
rect 3281 4545 3282 4549
rect 3286 4545 3287 4549
rect 3291 4545 3292 4549
rect 3296 4545 3297 4549
rect 3301 4545 3302 4549
rect 3306 4545 3307 4549
rect 3311 4545 3312 4549
rect 3316 4545 3318 4549
rect 3105 4462 3108 4466
rect 3112 4462 3113 4466
rect 3117 4462 3118 4466
rect 3122 4462 3123 4466
rect 3127 4462 3128 4466
rect 3132 4462 3133 4466
rect 3137 4462 3138 4466
rect 3142 4462 3143 4466
rect 3147 4462 3148 4466
rect 3152 4462 3153 4466
rect 3157 4462 3158 4466
rect 3162 4462 3165 4466
rect 3250 4466 3318 4545
rect 3332 4519 3336 4531
rect 3332 4503 3336 4515
rect 3332 4487 3336 4499
rect 3390 4519 3394 4531
rect 3390 4503 3394 4515
rect 3390 4487 3394 4499
rect 3254 4462 3257 4466
rect 3261 4462 3262 4466
rect 3266 4462 3267 4466
rect 3271 4462 3272 4466
rect 3276 4462 3277 4466
rect 3281 4462 3282 4466
rect 3286 4462 3287 4466
rect 3291 4462 3292 4466
rect 3296 4462 3297 4466
rect 3301 4462 3302 4466
rect 3306 4462 3307 4466
rect 3311 4462 3314 4466
rect 3410 4466 3478 4602
rect 3525 4613 3544 4614
rect 3668 4624 3669 4628
rect 3673 4624 3674 4628
rect 3678 4624 3679 4628
rect 3683 4624 3684 4628
rect 3664 4623 3684 4624
rect 3668 4619 3669 4623
rect 3673 4619 3674 4623
rect 3678 4619 3679 4623
rect 3683 4619 3684 4623
rect 3664 4618 3684 4619
rect 3668 4614 3669 4618
rect 3673 4614 3674 4618
rect 3678 4614 3679 4618
rect 3683 4614 3684 4618
rect 3838 4624 3839 4628
rect 3843 4624 3844 4628
rect 3848 4624 3849 4628
rect 3834 4623 3853 4624
rect 3838 4619 3839 4623
rect 3843 4619 3844 4623
rect 3848 4619 3849 4623
rect 3834 4618 3853 4619
rect 3838 4614 3839 4618
rect 3843 4614 3844 4618
rect 3848 4614 3849 4618
rect 3664 4613 3684 4614
rect 3529 4609 3530 4613
rect 3534 4609 3535 4613
rect 3539 4609 3540 4613
rect 3525 4608 3544 4609
rect 3529 4604 3530 4608
rect 3534 4604 3535 4608
rect 3539 4604 3540 4608
rect 3525 4603 3544 4604
rect 3529 4599 3530 4603
rect 3534 4599 3535 4603
rect 3539 4599 3540 4603
rect 3525 4598 3544 4599
rect 3529 4594 3530 4598
rect 3534 4594 3535 4598
rect 3539 4594 3540 4598
rect 3547 4611 3603 4613
rect 3547 4607 3549 4611
rect 3553 4607 3554 4611
rect 3558 4607 3559 4611
rect 3563 4607 3564 4611
rect 3568 4607 3569 4611
rect 3573 4607 3574 4611
rect 3578 4607 3579 4611
rect 3583 4607 3584 4611
rect 3588 4607 3589 4611
rect 3593 4607 3594 4611
rect 3598 4607 3599 4611
rect 3547 4606 3603 4607
rect 3547 4602 3549 4606
rect 3553 4602 3554 4606
rect 3558 4602 3559 4606
rect 3563 4602 3564 4606
rect 3568 4602 3569 4606
rect 3573 4602 3574 4606
rect 3578 4602 3579 4606
rect 3583 4602 3584 4606
rect 3588 4602 3589 4606
rect 3593 4602 3594 4606
rect 3598 4602 3599 4606
rect 3547 4601 3603 4602
rect 3547 4597 3549 4601
rect 3553 4597 3554 4601
rect 3558 4597 3559 4601
rect 3563 4597 3564 4601
rect 3568 4597 3569 4601
rect 3573 4597 3574 4601
rect 3578 4597 3579 4601
rect 3583 4597 3584 4601
rect 3588 4597 3589 4601
rect 3593 4597 3594 4601
rect 3598 4597 3599 4601
rect 3668 4609 3669 4613
rect 3673 4609 3674 4613
rect 3678 4609 3679 4613
rect 3683 4609 3684 4613
rect 3664 4608 3684 4609
rect 3668 4604 3669 4608
rect 3673 4604 3674 4608
rect 3678 4604 3679 4608
rect 3683 4604 3684 4608
rect 3664 4603 3684 4604
rect 3668 4599 3669 4603
rect 3673 4599 3674 4603
rect 3678 4599 3679 4603
rect 3683 4599 3684 4603
rect 3719 4611 3787 4614
rect 3719 4607 3721 4611
rect 3725 4607 3726 4611
rect 3730 4607 3731 4611
rect 3735 4607 3736 4611
rect 3740 4607 3741 4611
rect 3745 4607 3746 4611
rect 3750 4607 3751 4611
rect 3755 4607 3756 4611
rect 3760 4607 3761 4611
rect 3765 4607 3766 4611
rect 3770 4607 3771 4611
rect 3775 4607 3776 4611
rect 3780 4607 3781 4611
rect 3785 4607 3787 4611
rect 3719 4606 3787 4607
rect 3719 4602 3721 4606
rect 3725 4602 3726 4606
rect 3730 4602 3731 4606
rect 3735 4602 3736 4606
rect 3740 4602 3741 4606
rect 3745 4602 3746 4606
rect 3750 4602 3751 4606
rect 3755 4602 3756 4606
rect 3760 4602 3761 4606
rect 3765 4602 3766 4606
rect 3770 4602 3771 4606
rect 3775 4602 3776 4606
rect 3780 4602 3781 4606
rect 3785 4602 3787 4606
rect 3547 4596 3603 4597
rect 3547 4592 3549 4596
rect 3553 4592 3554 4596
rect 3558 4592 3559 4596
rect 3563 4592 3564 4596
rect 3568 4592 3569 4596
rect 3573 4592 3574 4596
rect 3578 4592 3579 4596
rect 3583 4592 3584 4596
rect 3588 4592 3589 4596
rect 3593 4592 3594 4596
rect 3598 4592 3599 4596
rect 3490 4578 3511 4580
rect 3494 4574 3495 4578
rect 3499 4574 3500 4578
rect 3504 4574 3505 4578
rect 3509 4574 3511 4578
rect 3490 4573 3511 4574
rect 3494 4569 3495 4573
rect 3499 4569 3500 4573
rect 3504 4569 3505 4573
rect 3509 4569 3511 4573
rect 3490 4568 3511 4569
rect 3494 4564 3495 4568
rect 3499 4564 3500 4568
rect 3504 4564 3505 4568
rect 3509 4564 3511 4568
rect 3490 4563 3511 4564
rect 3494 4559 3495 4563
rect 3499 4559 3500 4563
rect 3504 4559 3505 4563
rect 3509 4559 3511 4563
rect 3490 4558 3511 4559
rect 3494 4554 3495 4558
rect 3499 4554 3500 4558
rect 3504 4554 3505 4558
rect 3509 4554 3511 4558
rect 3490 4553 3511 4554
rect 3494 4549 3495 4553
rect 3499 4549 3500 4553
rect 3504 4549 3505 4553
rect 3509 4549 3511 4553
rect 3490 4548 3511 4549
rect 3529 4578 3530 4582
rect 3534 4578 3535 4582
rect 3539 4578 3540 4582
rect 3525 4577 3544 4578
rect 3529 4573 3530 4577
rect 3534 4573 3535 4577
rect 3539 4573 3540 4577
rect 3525 4572 3544 4573
rect 3529 4568 3530 4572
rect 3534 4568 3535 4572
rect 3539 4568 3540 4572
rect 3525 4567 3544 4568
rect 3529 4563 3530 4567
rect 3534 4563 3535 4567
rect 3539 4563 3540 4567
rect 3525 4562 3544 4563
rect 3529 4558 3530 4562
rect 3534 4558 3535 4562
rect 3539 4558 3540 4562
rect 3525 4557 3544 4558
rect 3529 4553 3530 4557
rect 3534 4553 3535 4557
rect 3539 4553 3540 4557
rect 3525 4552 3544 4553
rect 3529 4548 3530 4552
rect 3534 4548 3535 4552
rect 3539 4548 3540 4552
rect 3559 4554 3627 4557
rect 3559 4550 3561 4554
rect 3565 4550 3566 4554
rect 3570 4550 3571 4554
rect 3575 4550 3576 4554
rect 3580 4550 3581 4554
rect 3585 4550 3586 4554
rect 3590 4550 3591 4554
rect 3595 4550 3596 4554
rect 3600 4550 3601 4554
rect 3605 4550 3606 4554
rect 3610 4550 3611 4554
rect 3615 4550 3616 4554
rect 3620 4550 3621 4554
rect 3625 4550 3627 4554
rect 3559 4549 3627 4550
rect 3494 4544 3495 4548
rect 3499 4544 3500 4548
rect 3504 4544 3505 4548
rect 3509 4544 3511 4548
rect 3490 4543 3511 4544
rect 3494 4539 3495 4543
rect 3499 4539 3500 4543
rect 3504 4539 3505 4543
rect 3509 4539 3511 4543
rect 3490 4538 3511 4539
rect 3494 4534 3495 4538
rect 3499 4534 3500 4538
rect 3504 4534 3505 4538
rect 3509 4534 3511 4538
rect 3490 4533 3511 4534
rect 3494 4529 3495 4533
rect 3499 4529 3500 4533
rect 3504 4529 3505 4533
rect 3509 4529 3511 4533
rect 3490 4528 3511 4529
rect 3494 4524 3495 4528
rect 3499 4524 3500 4528
rect 3504 4524 3505 4528
rect 3509 4524 3511 4528
rect 3490 4523 3511 4524
rect 3494 4519 3495 4523
rect 3499 4519 3500 4523
rect 3504 4519 3505 4523
rect 3509 4519 3511 4523
rect 3490 4518 3511 4519
rect 3494 4514 3495 4518
rect 3499 4514 3500 4518
rect 3504 4514 3505 4518
rect 3509 4514 3511 4518
rect 3490 4512 3511 4514
rect 3559 4545 3561 4549
rect 3565 4545 3566 4549
rect 3570 4545 3571 4549
rect 3575 4545 3576 4549
rect 3580 4545 3581 4549
rect 3585 4545 3586 4549
rect 3590 4545 3591 4549
rect 3595 4545 3596 4549
rect 3600 4545 3601 4549
rect 3605 4545 3606 4549
rect 3610 4545 3611 4549
rect 3615 4545 3616 4549
rect 3620 4545 3621 4549
rect 3625 4545 3627 4549
rect 3414 4462 3417 4466
rect 3421 4462 3422 4466
rect 3426 4462 3427 4466
rect 3431 4462 3432 4466
rect 3436 4462 3437 4466
rect 3441 4462 3442 4466
rect 3446 4462 3447 4466
rect 3451 4462 3452 4466
rect 3456 4462 3457 4466
rect 3461 4462 3462 4466
rect 3466 4462 3467 4466
rect 3471 4462 3474 4466
rect 3559 4466 3627 4545
rect 3563 4462 3566 4466
rect 3570 4462 3571 4466
rect 3575 4462 3576 4466
rect 3580 4462 3581 4466
rect 3585 4462 3586 4466
rect 3590 4462 3591 4466
rect 3595 4462 3596 4466
rect 3600 4462 3601 4466
rect 3605 4462 3606 4466
rect 3610 4462 3611 4466
rect 3615 4462 3616 4466
rect 3620 4462 3623 4466
rect 3719 4466 3787 4602
rect 3834 4613 3853 4614
rect 3838 4609 3839 4613
rect 3843 4609 3844 4613
rect 3848 4609 3849 4613
rect 3834 4608 3853 4609
rect 3838 4604 3839 4608
rect 3843 4604 3844 4608
rect 3848 4604 3849 4608
rect 3834 4603 3853 4604
rect 3838 4599 3839 4603
rect 3843 4599 3844 4603
rect 3848 4599 3849 4603
rect 3834 4598 3853 4599
rect 3838 4594 3839 4598
rect 3843 4594 3844 4598
rect 3848 4594 3849 4598
rect 4239 4624 4240 4628
rect 4244 4624 4245 4628
rect 4249 4624 4250 4628
rect 4235 4623 4254 4624
rect 4239 4619 4240 4623
rect 4244 4619 4245 4623
rect 4249 4619 4250 4623
rect 4235 4618 4254 4619
rect 4239 4614 4240 4618
rect 4244 4614 4245 4618
rect 4249 4614 4250 4618
rect 4235 4613 4254 4614
rect 4239 4609 4240 4613
rect 4244 4609 4245 4613
rect 4249 4609 4250 4613
rect 4235 4608 4254 4609
rect 4239 4604 4240 4608
rect 4244 4604 4245 4608
rect 4249 4604 4250 4608
rect 4235 4603 4254 4604
rect 4239 4599 4240 4603
rect 4244 4599 4245 4603
rect 4249 4599 4250 4603
rect 4235 4598 4254 4599
rect 4239 4594 4240 4598
rect 4244 4594 4245 4598
rect 4249 4594 4250 4598
rect 4268 4624 4269 4628
rect 4273 4624 4274 4628
rect 4278 4624 4279 4628
rect 4264 4623 4283 4624
rect 4268 4619 4269 4623
rect 4273 4619 4274 4623
rect 4278 4619 4279 4623
rect 4264 4618 4283 4619
rect 4268 4614 4269 4618
rect 4273 4614 4274 4618
rect 4278 4614 4279 4618
rect 4264 4613 4283 4614
rect 4268 4609 4269 4613
rect 4273 4609 4274 4613
rect 4278 4609 4279 4613
rect 4264 4608 4283 4609
rect 4268 4604 4269 4608
rect 4273 4604 4274 4608
rect 4278 4604 4279 4608
rect 4264 4603 4283 4604
rect 4268 4599 4269 4603
rect 4273 4599 4274 4603
rect 4278 4599 4279 4603
rect 4264 4598 4283 4599
rect 4268 4594 4269 4598
rect 4273 4594 4274 4598
rect 4278 4594 4279 4598
rect 4297 4624 4298 4628
rect 4302 4624 4303 4628
rect 4307 4624 4308 4628
rect 4293 4623 4312 4624
rect 4297 4619 4298 4623
rect 4302 4619 4303 4623
rect 4307 4619 4308 4623
rect 4293 4618 4312 4619
rect 4297 4614 4298 4618
rect 4302 4614 4303 4618
rect 4307 4614 4308 4618
rect 4293 4613 4312 4614
rect 4297 4609 4298 4613
rect 4302 4609 4303 4613
rect 4307 4609 4308 4613
rect 4293 4608 4312 4609
rect 4297 4604 4298 4608
rect 4302 4604 4303 4608
rect 4307 4604 4308 4608
rect 4293 4603 4312 4604
rect 4297 4599 4298 4603
rect 4302 4599 4303 4603
rect 4307 4599 4308 4603
rect 4293 4598 4312 4599
rect 4297 4594 4298 4598
rect 4302 4594 4303 4598
rect 4307 4594 4308 4598
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4336 4624 4337 4628
rect 4322 4623 4341 4624
rect 4326 4619 4327 4623
rect 4331 4619 4332 4623
rect 4336 4619 4337 4623
rect 4322 4618 4341 4619
rect 4326 4614 4327 4618
rect 4331 4614 4332 4618
rect 4336 4614 4337 4618
rect 4322 4613 4341 4614
rect 4326 4609 4327 4613
rect 4331 4609 4332 4613
rect 4336 4609 4337 4613
rect 4322 4608 4341 4609
rect 4326 4604 4327 4608
rect 4331 4604 4332 4608
rect 4336 4604 4337 4608
rect 4322 4603 4341 4604
rect 4326 4599 4327 4603
rect 4331 4599 4332 4603
rect 4336 4599 4337 4603
rect 4322 4598 4341 4599
rect 4326 4594 4327 4598
rect 4331 4594 4332 4598
rect 4336 4594 4337 4598
rect 4355 4624 4356 4628
rect 4360 4624 4361 4628
rect 4365 4624 4366 4628
rect 4351 4623 4370 4624
rect 4355 4619 4356 4623
rect 4360 4619 4361 4623
rect 4365 4619 4366 4623
rect 4351 4618 4370 4619
rect 4355 4614 4356 4618
rect 4360 4614 4361 4618
rect 4365 4614 4366 4618
rect 4351 4613 4370 4614
rect 4355 4609 4356 4613
rect 4360 4609 4361 4613
rect 4365 4609 4366 4613
rect 4351 4608 4370 4609
rect 4355 4604 4356 4608
rect 4360 4604 4361 4608
rect 4365 4604 4366 4608
rect 4351 4603 4370 4604
rect 4355 4599 4356 4603
rect 4360 4599 4361 4603
rect 4365 4599 4366 4603
rect 4351 4598 4370 4599
rect 4355 4594 4356 4598
rect 4360 4594 4361 4598
rect 4365 4594 4366 4598
rect 3799 4578 3820 4580
rect 3803 4574 3804 4578
rect 3808 4574 3809 4578
rect 3813 4574 3814 4578
rect 3818 4574 3820 4578
rect 3799 4573 3820 4574
rect 3803 4569 3804 4573
rect 3808 4569 3809 4573
rect 3813 4569 3814 4573
rect 3818 4569 3820 4573
rect 3799 4568 3820 4569
rect 3803 4564 3804 4568
rect 3808 4564 3809 4568
rect 3813 4564 3814 4568
rect 3818 4564 3820 4568
rect 3799 4563 3820 4564
rect 3803 4559 3804 4563
rect 3808 4559 3809 4563
rect 3813 4559 3814 4563
rect 3818 4559 3820 4563
rect 3799 4558 3820 4559
rect 3803 4554 3804 4558
rect 3808 4554 3809 4558
rect 3813 4554 3814 4558
rect 3818 4554 3820 4558
rect 3799 4553 3820 4554
rect 3803 4549 3804 4553
rect 3808 4549 3809 4553
rect 3813 4549 3814 4553
rect 3818 4549 3820 4553
rect 3799 4548 3820 4549
rect 3838 4578 3839 4582
rect 3843 4578 3844 4582
rect 3848 4578 3849 4582
rect 3834 4577 3853 4578
rect 3838 4573 3839 4577
rect 3843 4573 3844 4577
rect 3848 4573 3849 4577
rect 3834 4572 3853 4573
rect 3838 4568 3839 4572
rect 3843 4568 3844 4572
rect 3848 4568 3849 4572
rect 3834 4567 3853 4568
rect 3838 4563 3839 4567
rect 3843 4563 3844 4567
rect 3848 4563 3849 4567
rect 3834 4562 3853 4563
rect 3838 4558 3839 4562
rect 3843 4558 3844 4562
rect 3848 4558 3849 4562
rect 3834 4557 3853 4558
rect 3838 4553 3839 4557
rect 3843 4553 3844 4557
rect 3848 4553 3849 4557
rect 3834 4552 3853 4553
rect 3838 4548 3839 4552
rect 3843 4548 3844 4552
rect 3848 4548 3849 4552
rect 4239 4578 4240 4582
rect 4244 4578 4245 4582
rect 4249 4578 4250 4582
rect 4235 4577 4254 4578
rect 4239 4573 4240 4577
rect 4244 4573 4245 4577
rect 4249 4573 4250 4577
rect 4235 4572 4254 4573
rect 4239 4568 4240 4572
rect 4244 4568 4245 4572
rect 4249 4568 4250 4572
rect 4235 4567 4254 4568
rect 4239 4563 4240 4567
rect 4244 4563 4245 4567
rect 4249 4563 4250 4567
rect 4235 4562 4254 4563
rect 4239 4558 4240 4562
rect 4244 4558 4245 4562
rect 4249 4558 4250 4562
rect 4235 4557 4254 4558
rect 4239 4553 4240 4557
rect 4244 4553 4245 4557
rect 4249 4553 4250 4557
rect 4235 4552 4254 4553
rect 4239 4548 4240 4552
rect 4244 4548 4245 4552
rect 4249 4548 4250 4552
rect 4268 4578 4269 4582
rect 4273 4578 4274 4582
rect 4278 4578 4279 4582
rect 4264 4577 4283 4578
rect 4268 4573 4269 4577
rect 4273 4573 4274 4577
rect 4278 4573 4279 4577
rect 4264 4572 4283 4573
rect 4268 4568 4269 4572
rect 4273 4568 4274 4572
rect 4278 4568 4279 4572
rect 4264 4567 4283 4568
rect 4268 4563 4269 4567
rect 4273 4563 4274 4567
rect 4278 4563 4279 4567
rect 4264 4562 4283 4563
rect 4268 4558 4269 4562
rect 4273 4558 4274 4562
rect 4278 4558 4279 4562
rect 4264 4557 4283 4558
rect 4268 4553 4269 4557
rect 4273 4553 4274 4557
rect 4278 4553 4279 4557
rect 4264 4552 4283 4553
rect 4268 4548 4269 4552
rect 4273 4548 4274 4552
rect 4278 4548 4279 4552
rect 4297 4578 4298 4582
rect 4302 4578 4303 4582
rect 4307 4578 4308 4582
rect 4293 4577 4312 4578
rect 4297 4573 4298 4577
rect 4302 4573 4303 4577
rect 4307 4573 4308 4577
rect 4293 4572 4312 4573
rect 4297 4568 4298 4572
rect 4302 4568 4303 4572
rect 4307 4568 4308 4572
rect 4293 4567 4312 4568
rect 4297 4563 4298 4567
rect 4302 4563 4303 4567
rect 4307 4563 4308 4567
rect 4293 4562 4312 4563
rect 4297 4558 4298 4562
rect 4302 4558 4303 4562
rect 4307 4558 4308 4562
rect 4293 4557 4312 4558
rect 4297 4553 4298 4557
rect 4302 4553 4303 4557
rect 4307 4553 4308 4557
rect 4293 4552 4312 4553
rect 4297 4548 4298 4552
rect 4302 4548 4303 4552
rect 4307 4548 4308 4552
rect 4326 4578 4327 4582
rect 4331 4578 4332 4582
rect 4336 4578 4337 4582
rect 4322 4577 4341 4578
rect 4326 4573 4327 4577
rect 4331 4573 4332 4577
rect 4336 4573 4337 4577
rect 4322 4572 4341 4573
rect 4326 4568 4327 4572
rect 4331 4568 4332 4572
rect 4336 4568 4337 4572
rect 4322 4567 4341 4568
rect 4326 4563 4327 4567
rect 4331 4563 4332 4567
rect 4336 4563 4337 4567
rect 4322 4562 4341 4563
rect 4326 4558 4327 4562
rect 4331 4558 4332 4562
rect 4336 4558 4337 4562
rect 4322 4557 4341 4558
rect 4326 4553 4327 4557
rect 4331 4553 4332 4557
rect 4336 4553 4337 4557
rect 4322 4552 4341 4553
rect 4326 4548 4327 4552
rect 4331 4548 4332 4552
rect 4336 4548 4337 4552
rect 4355 4578 4356 4582
rect 4360 4578 4361 4582
rect 4365 4578 4366 4582
rect 4351 4577 4370 4578
rect 4355 4573 4356 4577
rect 4360 4573 4361 4577
rect 4365 4573 4366 4577
rect 4351 4572 4370 4573
rect 4355 4568 4356 4572
rect 4360 4568 4361 4572
rect 4365 4568 4366 4572
rect 4351 4567 4370 4568
rect 4355 4563 4356 4567
rect 4360 4563 4361 4567
rect 4365 4563 4366 4567
rect 4351 4562 4370 4563
rect 4355 4558 4356 4562
rect 4360 4558 4361 4562
rect 4365 4558 4366 4562
rect 4351 4557 4370 4558
rect 4355 4553 4356 4557
rect 4360 4553 4361 4557
rect 4365 4553 4366 4557
rect 4351 4552 4370 4553
rect 4355 4548 4356 4552
rect 4360 4548 4361 4552
rect 4365 4548 4366 4552
rect 3803 4544 3804 4548
rect 3808 4544 3809 4548
rect 3813 4544 3814 4548
rect 3818 4544 3820 4548
rect 3799 4543 3820 4544
rect 3803 4539 3804 4543
rect 3808 4539 3809 4543
rect 3813 4539 3814 4543
rect 3818 4539 3820 4543
rect 3799 4538 3820 4539
rect 3803 4534 3804 4538
rect 3808 4534 3809 4538
rect 3813 4534 3814 4538
rect 3818 4534 3820 4538
rect 3799 4533 3820 4534
rect 3803 4529 3804 4533
rect 3808 4529 3809 4533
rect 3813 4529 3814 4533
rect 3818 4529 3820 4533
rect 3799 4528 3820 4529
rect 4579 4528 5054 4966
rect 3803 4524 3804 4528
rect 3808 4524 3809 4528
rect 3813 4524 3814 4528
rect 3818 4524 3820 4528
rect 3799 4523 3820 4524
rect 3803 4519 3804 4523
rect 3808 4519 3809 4523
rect 3813 4519 3814 4523
rect 3818 4519 3820 4523
rect 3799 4518 3820 4519
rect 3803 4514 3804 4518
rect 3808 4514 3809 4518
rect 3813 4514 3814 4518
rect 3818 4514 3820 4518
rect 3799 4512 3820 4514
rect 3723 4462 3726 4466
rect 3730 4462 3731 4466
rect 3735 4462 3736 4466
rect 3740 4462 3741 4466
rect 3745 4462 3746 4466
rect 3750 4462 3751 4466
rect 3755 4462 3756 4466
rect 3760 4462 3761 4466
rect 3765 4462 3766 4466
rect 3770 4462 3771 4466
rect 3775 4462 3776 4466
rect 3780 4462 3783 4466
rect 1099 4446 1104 4450
rect 1108 4446 1114 4450
rect 1118 4446 1124 4450
rect 1128 4446 1134 4450
rect 1138 4446 1264 4450
rect 1268 4446 1274 4450
rect 1278 4446 1284 4450
rect 1288 4446 1294 4450
rect 1298 4446 1303 4450
rect 1099 4445 1303 4446
rect 1103 4441 1109 4445
rect 1113 4441 1119 4445
rect 1123 4441 1129 4445
rect 1133 4441 1139 4445
rect 1143 4441 1259 4445
rect 1263 4441 1269 4445
rect 1273 4441 1279 4445
rect 1283 4441 1289 4445
rect 1293 4441 1299 4445
rect 1099 4440 1303 4441
rect 1099 4436 1104 4440
rect 1108 4436 1114 4440
rect 1118 4436 1124 4440
rect 1128 4436 1134 4440
rect 1138 4436 1264 4440
rect 1268 4436 1274 4440
rect 1278 4436 1284 4440
rect 1288 4436 1294 4440
rect 1298 4436 1303 4440
rect 1099 4435 1303 4436
rect 1103 4431 1109 4435
rect 1113 4431 1119 4435
rect 1123 4431 1129 4435
rect 1133 4431 1139 4435
rect 1143 4431 1259 4435
rect 1263 4431 1269 4435
rect 1273 4431 1279 4435
rect 1283 4431 1289 4435
rect 1293 4431 1299 4435
rect 1099 4430 1303 4431
rect 1099 4426 1104 4430
rect 1108 4426 1114 4430
rect 1118 4426 1124 4430
rect 1128 4426 1134 4430
rect 1138 4426 1264 4430
rect 1268 4426 1274 4430
rect 1278 4426 1284 4430
rect 1288 4426 1294 4430
rect 1298 4426 1303 4430
rect 1099 4425 1303 4426
rect 1103 4421 1109 4425
rect 1113 4421 1119 4425
rect 1123 4421 1129 4425
rect 1133 4421 1139 4425
rect 1143 4421 1259 4425
rect 1263 4421 1269 4425
rect 1273 4421 1279 4425
rect 1283 4421 1289 4425
rect 1293 4421 1299 4425
rect 1099 4420 1303 4421
rect 1099 4416 1104 4420
rect 1108 4416 1114 4420
rect 1118 4416 1124 4420
rect 1128 4416 1134 4420
rect 1138 4416 1264 4420
rect 1268 4416 1274 4420
rect 1278 4416 1284 4420
rect 1288 4416 1294 4420
rect 1298 4416 1303 4420
rect 1099 4415 1303 4416
rect 1103 4411 1109 4415
rect 1113 4411 1119 4415
rect 1123 4411 1129 4415
rect 1133 4411 1139 4415
rect 1143 4411 1259 4415
rect 1263 4411 1269 4415
rect 1273 4411 1279 4415
rect 1283 4411 1289 4415
rect 1293 4411 1299 4415
rect 1099 4410 1303 4411
rect 1099 4406 1104 4410
rect 1108 4406 1114 4410
rect 1118 4406 1124 4410
rect 1128 4406 1134 4410
rect 1138 4406 1264 4410
rect 1268 4406 1274 4410
rect 1278 4406 1284 4410
rect 1288 4406 1294 4410
rect 1298 4406 1303 4410
rect 1099 4405 1303 4406
rect 1103 4401 1109 4405
rect 1113 4401 1119 4405
rect 1123 4401 1129 4405
rect 1133 4401 1139 4405
rect 1143 4401 1259 4405
rect 1263 4401 1269 4405
rect 1273 4401 1279 4405
rect 1283 4401 1289 4405
rect 1293 4401 1299 4405
rect 1099 4400 1303 4401
rect 1099 4396 1104 4400
rect 1108 4396 1114 4400
rect 1118 4396 1124 4400
rect 1128 4396 1134 4400
rect 1138 4396 1264 4400
rect 1268 4396 1274 4400
rect 1278 4396 1284 4400
rect 1288 4396 1294 4400
rect 1298 4396 1303 4400
rect 1099 4395 1303 4396
rect 1103 4391 1109 4395
rect 1113 4391 1119 4395
rect 1123 4391 1129 4395
rect 1133 4391 1139 4395
rect 1143 4391 1259 4395
rect 1263 4391 1269 4395
rect 1273 4391 1279 4395
rect 1283 4391 1289 4395
rect 1293 4391 1299 4395
rect 1099 4390 1303 4391
rect 1099 4386 1104 4390
rect 1108 4386 1114 4390
rect 1118 4386 1124 4390
rect 1128 4386 1134 4390
rect 1138 4386 1264 4390
rect 1268 4386 1274 4390
rect 1278 4386 1284 4390
rect 1288 4386 1294 4390
rect 1298 4386 1303 4390
rect 1099 4385 1303 4386
rect 1103 4381 1109 4385
rect 1113 4381 1119 4385
rect 1123 4381 1129 4385
rect 1133 4381 1139 4385
rect 1143 4381 1259 4385
rect 1263 4381 1269 4385
rect 1273 4381 1279 4385
rect 1283 4381 1289 4385
rect 1293 4381 1299 4385
rect 1099 4380 1303 4381
rect 1099 4376 1104 4380
rect 1108 4376 1114 4380
rect 1118 4376 1124 4380
rect 1128 4376 1134 4380
rect 1138 4376 1264 4380
rect 1268 4376 1274 4380
rect 1278 4376 1284 4380
rect 1288 4376 1294 4380
rect 1298 4376 1303 4380
rect 1099 4375 1303 4376
rect 1103 4371 1109 4375
rect 1113 4371 1119 4375
rect 1123 4371 1129 4375
rect 1133 4371 1139 4375
rect 1143 4371 1259 4375
rect 1263 4371 1269 4375
rect 1273 4371 1279 4375
rect 1283 4371 1289 4375
rect 1293 4371 1299 4375
rect 1099 4370 1303 4371
rect 1099 4366 1104 4370
rect 1108 4366 1114 4370
rect 1118 4366 1124 4370
rect 1128 4366 1134 4370
rect 1138 4366 1264 4370
rect 1268 4366 1274 4370
rect 1278 4366 1284 4370
rect 1288 4366 1294 4370
rect 1298 4366 1303 4370
rect 1099 4365 1303 4366
rect 1103 4361 1109 4365
rect 1113 4361 1119 4365
rect 1123 4361 1129 4365
rect 1133 4361 1139 4365
rect 1143 4361 1259 4365
rect 1263 4361 1269 4365
rect 1273 4361 1279 4365
rect 1283 4361 1289 4365
rect 1293 4361 1299 4365
rect 1408 4446 1413 4450
rect 1417 4446 1423 4450
rect 1427 4446 1433 4450
rect 1437 4446 1443 4450
rect 1447 4446 1573 4450
rect 1577 4446 1583 4450
rect 1587 4446 1593 4450
rect 1597 4446 1603 4450
rect 1607 4446 1612 4450
rect 1408 4445 1612 4446
rect 1412 4441 1418 4445
rect 1422 4441 1428 4445
rect 1432 4441 1438 4445
rect 1442 4441 1448 4445
rect 1452 4441 1568 4445
rect 1572 4441 1578 4445
rect 1582 4441 1588 4445
rect 1592 4441 1598 4445
rect 1602 4441 1608 4445
rect 1408 4440 1612 4441
rect 1408 4436 1413 4440
rect 1417 4436 1423 4440
rect 1427 4436 1433 4440
rect 1437 4436 1443 4440
rect 1447 4436 1573 4440
rect 1577 4436 1583 4440
rect 1587 4436 1593 4440
rect 1597 4436 1603 4440
rect 1607 4436 1612 4440
rect 1408 4435 1612 4436
rect 1412 4431 1418 4435
rect 1422 4431 1428 4435
rect 1432 4431 1438 4435
rect 1442 4431 1448 4435
rect 1452 4431 1568 4435
rect 1572 4431 1578 4435
rect 1582 4431 1588 4435
rect 1592 4431 1598 4435
rect 1602 4431 1608 4435
rect 1408 4430 1612 4431
rect 1408 4426 1413 4430
rect 1417 4426 1423 4430
rect 1427 4426 1433 4430
rect 1437 4426 1443 4430
rect 1447 4426 1573 4430
rect 1577 4426 1583 4430
rect 1587 4426 1593 4430
rect 1597 4426 1603 4430
rect 1607 4426 1612 4430
rect 1408 4425 1612 4426
rect 1412 4421 1418 4425
rect 1422 4421 1428 4425
rect 1432 4421 1438 4425
rect 1442 4421 1448 4425
rect 1452 4421 1568 4425
rect 1572 4421 1578 4425
rect 1582 4421 1588 4425
rect 1592 4421 1598 4425
rect 1602 4421 1608 4425
rect 1408 4420 1612 4421
rect 1408 4416 1413 4420
rect 1417 4416 1423 4420
rect 1427 4416 1433 4420
rect 1437 4416 1443 4420
rect 1447 4416 1573 4420
rect 1577 4416 1583 4420
rect 1587 4416 1593 4420
rect 1597 4416 1603 4420
rect 1607 4416 1612 4420
rect 1408 4415 1612 4416
rect 1412 4411 1418 4415
rect 1422 4411 1428 4415
rect 1432 4411 1438 4415
rect 1442 4411 1448 4415
rect 1452 4411 1568 4415
rect 1572 4411 1578 4415
rect 1582 4411 1588 4415
rect 1592 4411 1598 4415
rect 1602 4411 1608 4415
rect 1408 4410 1612 4411
rect 1408 4406 1413 4410
rect 1417 4406 1423 4410
rect 1427 4406 1433 4410
rect 1437 4406 1443 4410
rect 1447 4406 1573 4410
rect 1577 4406 1583 4410
rect 1587 4406 1593 4410
rect 1597 4406 1603 4410
rect 1607 4406 1612 4410
rect 1408 4405 1612 4406
rect 1412 4401 1418 4405
rect 1422 4401 1428 4405
rect 1432 4401 1438 4405
rect 1442 4401 1448 4405
rect 1452 4401 1568 4405
rect 1572 4401 1578 4405
rect 1582 4401 1588 4405
rect 1592 4401 1598 4405
rect 1602 4401 1608 4405
rect 1408 4400 1612 4401
rect 1408 4396 1413 4400
rect 1417 4396 1423 4400
rect 1427 4396 1433 4400
rect 1437 4396 1443 4400
rect 1447 4396 1573 4400
rect 1577 4396 1583 4400
rect 1587 4396 1593 4400
rect 1597 4396 1603 4400
rect 1607 4396 1612 4400
rect 1408 4395 1612 4396
rect 1412 4391 1418 4395
rect 1422 4391 1428 4395
rect 1432 4391 1438 4395
rect 1442 4391 1448 4395
rect 1452 4391 1568 4395
rect 1572 4391 1578 4395
rect 1582 4391 1588 4395
rect 1592 4391 1598 4395
rect 1602 4391 1608 4395
rect 1408 4390 1612 4391
rect 1408 4386 1413 4390
rect 1417 4386 1423 4390
rect 1427 4386 1433 4390
rect 1437 4386 1443 4390
rect 1447 4386 1573 4390
rect 1577 4386 1583 4390
rect 1587 4386 1593 4390
rect 1597 4386 1603 4390
rect 1607 4386 1612 4390
rect 1408 4385 1612 4386
rect 1412 4381 1418 4385
rect 1422 4381 1428 4385
rect 1432 4381 1438 4385
rect 1442 4381 1448 4385
rect 1452 4381 1568 4385
rect 1572 4381 1578 4385
rect 1582 4381 1588 4385
rect 1592 4381 1598 4385
rect 1602 4381 1608 4385
rect 1408 4380 1612 4381
rect 1408 4376 1413 4380
rect 1417 4376 1423 4380
rect 1427 4376 1433 4380
rect 1437 4376 1443 4380
rect 1447 4376 1573 4380
rect 1577 4376 1583 4380
rect 1587 4376 1593 4380
rect 1597 4376 1603 4380
rect 1607 4376 1612 4380
rect 1408 4375 1612 4376
rect 1412 4371 1418 4375
rect 1422 4371 1428 4375
rect 1432 4371 1438 4375
rect 1442 4371 1448 4375
rect 1452 4371 1568 4375
rect 1572 4371 1578 4375
rect 1582 4371 1588 4375
rect 1592 4371 1598 4375
rect 1602 4371 1608 4375
rect 1408 4370 1612 4371
rect 1408 4366 1413 4370
rect 1417 4366 1423 4370
rect 1427 4366 1433 4370
rect 1437 4366 1443 4370
rect 1447 4366 1573 4370
rect 1577 4366 1583 4370
rect 1587 4366 1593 4370
rect 1597 4366 1603 4370
rect 1607 4366 1612 4370
rect 1408 4365 1612 4366
rect 1412 4361 1418 4365
rect 1422 4361 1428 4365
rect 1432 4361 1438 4365
rect 1442 4361 1448 4365
rect 1452 4361 1568 4365
rect 1572 4361 1578 4365
rect 1582 4361 1588 4365
rect 1592 4361 1598 4365
rect 1602 4361 1608 4365
rect 1717 4446 1722 4450
rect 1726 4446 1732 4450
rect 1736 4446 1742 4450
rect 1746 4446 1752 4450
rect 1756 4446 1882 4450
rect 1886 4446 1892 4450
rect 1896 4446 1902 4450
rect 1906 4446 1912 4450
rect 1916 4446 1921 4450
rect 1717 4445 1921 4446
rect 1721 4441 1727 4445
rect 1731 4441 1737 4445
rect 1741 4441 1747 4445
rect 1751 4441 1757 4445
rect 1761 4441 1877 4445
rect 1881 4441 1887 4445
rect 1891 4441 1897 4445
rect 1901 4441 1907 4445
rect 1911 4441 1917 4445
rect 1717 4440 1921 4441
rect 1717 4436 1722 4440
rect 1726 4436 1732 4440
rect 1736 4436 1742 4440
rect 1746 4436 1752 4440
rect 1756 4436 1882 4440
rect 1886 4436 1892 4440
rect 1896 4436 1902 4440
rect 1906 4436 1912 4440
rect 1916 4436 1921 4440
rect 1717 4435 1921 4436
rect 1721 4431 1727 4435
rect 1731 4431 1737 4435
rect 1741 4431 1747 4435
rect 1751 4431 1757 4435
rect 1761 4431 1877 4435
rect 1881 4431 1887 4435
rect 1891 4431 1897 4435
rect 1901 4431 1907 4435
rect 1911 4431 1917 4435
rect 1717 4430 1921 4431
rect 1717 4426 1722 4430
rect 1726 4426 1732 4430
rect 1736 4426 1742 4430
rect 1746 4426 1752 4430
rect 1756 4426 1882 4430
rect 1886 4426 1892 4430
rect 1896 4426 1902 4430
rect 1906 4426 1912 4430
rect 1916 4426 1921 4430
rect 1717 4425 1921 4426
rect 1721 4421 1727 4425
rect 1731 4421 1737 4425
rect 1741 4421 1747 4425
rect 1751 4421 1757 4425
rect 1761 4421 1877 4425
rect 1881 4421 1887 4425
rect 1891 4421 1897 4425
rect 1901 4421 1907 4425
rect 1911 4421 1917 4425
rect 1717 4420 1921 4421
rect 1717 4416 1722 4420
rect 1726 4416 1732 4420
rect 1736 4416 1742 4420
rect 1746 4416 1752 4420
rect 1756 4416 1882 4420
rect 1886 4416 1892 4420
rect 1896 4416 1902 4420
rect 1906 4416 1912 4420
rect 1916 4416 1921 4420
rect 1717 4415 1921 4416
rect 1721 4411 1727 4415
rect 1731 4411 1737 4415
rect 1741 4411 1747 4415
rect 1751 4411 1757 4415
rect 1761 4411 1877 4415
rect 1881 4411 1887 4415
rect 1891 4411 1897 4415
rect 1901 4411 1907 4415
rect 1911 4411 1917 4415
rect 1717 4410 1921 4411
rect 1717 4406 1722 4410
rect 1726 4406 1732 4410
rect 1736 4406 1742 4410
rect 1746 4406 1752 4410
rect 1756 4406 1882 4410
rect 1886 4406 1892 4410
rect 1896 4406 1902 4410
rect 1906 4406 1912 4410
rect 1916 4406 1921 4410
rect 1717 4405 1921 4406
rect 1721 4401 1727 4405
rect 1731 4401 1737 4405
rect 1741 4401 1747 4405
rect 1751 4401 1757 4405
rect 1761 4401 1877 4405
rect 1881 4401 1887 4405
rect 1891 4401 1897 4405
rect 1901 4401 1907 4405
rect 1911 4401 1917 4405
rect 1717 4400 1921 4401
rect 1717 4396 1722 4400
rect 1726 4396 1732 4400
rect 1736 4396 1742 4400
rect 1746 4396 1752 4400
rect 1756 4396 1882 4400
rect 1886 4396 1892 4400
rect 1896 4396 1902 4400
rect 1906 4396 1912 4400
rect 1916 4396 1921 4400
rect 1717 4395 1921 4396
rect 1721 4391 1727 4395
rect 1731 4391 1737 4395
rect 1741 4391 1747 4395
rect 1751 4391 1757 4395
rect 1761 4391 1877 4395
rect 1881 4391 1887 4395
rect 1891 4391 1897 4395
rect 1901 4391 1907 4395
rect 1911 4391 1917 4395
rect 1717 4390 1921 4391
rect 1717 4386 1722 4390
rect 1726 4386 1732 4390
rect 1736 4386 1742 4390
rect 1746 4386 1752 4390
rect 1756 4386 1882 4390
rect 1886 4386 1892 4390
rect 1896 4386 1902 4390
rect 1906 4386 1912 4390
rect 1916 4386 1921 4390
rect 1717 4385 1921 4386
rect 1721 4381 1727 4385
rect 1731 4381 1737 4385
rect 1741 4381 1747 4385
rect 1751 4381 1757 4385
rect 1761 4381 1877 4385
rect 1881 4381 1887 4385
rect 1891 4381 1897 4385
rect 1901 4381 1907 4385
rect 1911 4381 1917 4385
rect 1717 4380 1921 4381
rect 1717 4376 1722 4380
rect 1726 4376 1732 4380
rect 1736 4376 1742 4380
rect 1746 4376 1752 4380
rect 1756 4376 1882 4380
rect 1886 4376 1892 4380
rect 1896 4376 1902 4380
rect 1906 4376 1912 4380
rect 1916 4376 1921 4380
rect 1717 4375 1921 4376
rect 1721 4371 1727 4375
rect 1731 4371 1737 4375
rect 1741 4371 1747 4375
rect 1751 4371 1757 4375
rect 1761 4371 1877 4375
rect 1881 4371 1887 4375
rect 1891 4371 1897 4375
rect 1901 4371 1907 4375
rect 1911 4371 1917 4375
rect 1717 4370 1921 4371
rect 1717 4366 1722 4370
rect 1726 4366 1732 4370
rect 1736 4366 1742 4370
rect 1746 4366 1752 4370
rect 1756 4366 1882 4370
rect 1886 4366 1892 4370
rect 1896 4366 1902 4370
rect 1906 4366 1912 4370
rect 1916 4366 1921 4370
rect 1717 4365 1921 4366
rect 1721 4361 1727 4365
rect 1731 4361 1737 4365
rect 1741 4361 1747 4365
rect 1751 4361 1757 4365
rect 1761 4361 1877 4365
rect 1881 4361 1887 4365
rect 1891 4361 1897 4365
rect 1901 4361 1907 4365
rect 1911 4361 1917 4365
rect 2026 4446 2031 4450
rect 2035 4446 2041 4450
rect 2045 4446 2051 4450
rect 2055 4446 2061 4450
rect 2065 4446 2191 4450
rect 2195 4446 2201 4450
rect 2205 4446 2211 4450
rect 2215 4446 2221 4450
rect 2225 4446 2230 4450
rect 2026 4445 2230 4446
rect 2030 4441 2036 4445
rect 2040 4441 2046 4445
rect 2050 4441 2056 4445
rect 2060 4441 2066 4445
rect 2070 4441 2186 4445
rect 2190 4441 2196 4445
rect 2200 4441 2206 4445
rect 2210 4441 2216 4445
rect 2220 4441 2226 4445
rect 2026 4440 2230 4441
rect 2026 4436 2031 4440
rect 2035 4436 2041 4440
rect 2045 4436 2051 4440
rect 2055 4436 2061 4440
rect 2065 4436 2191 4440
rect 2195 4436 2201 4440
rect 2205 4436 2211 4440
rect 2215 4436 2221 4440
rect 2225 4436 2230 4440
rect 2026 4435 2230 4436
rect 2030 4431 2036 4435
rect 2040 4431 2046 4435
rect 2050 4431 2056 4435
rect 2060 4431 2066 4435
rect 2070 4431 2186 4435
rect 2190 4431 2196 4435
rect 2200 4431 2206 4435
rect 2210 4431 2216 4435
rect 2220 4431 2226 4435
rect 2026 4430 2230 4431
rect 2026 4426 2031 4430
rect 2035 4426 2041 4430
rect 2045 4426 2051 4430
rect 2055 4426 2061 4430
rect 2065 4426 2191 4430
rect 2195 4426 2201 4430
rect 2205 4426 2211 4430
rect 2215 4426 2221 4430
rect 2225 4426 2230 4430
rect 2026 4425 2230 4426
rect 2030 4421 2036 4425
rect 2040 4421 2046 4425
rect 2050 4421 2056 4425
rect 2060 4421 2066 4425
rect 2070 4421 2186 4425
rect 2190 4421 2196 4425
rect 2200 4421 2206 4425
rect 2210 4421 2216 4425
rect 2220 4421 2226 4425
rect 2026 4420 2230 4421
rect 2026 4416 2031 4420
rect 2035 4416 2041 4420
rect 2045 4416 2051 4420
rect 2055 4416 2061 4420
rect 2065 4416 2191 4420
rect 2195 4416 2201 4420
rect 2205 4416 2211 4420
rect 2215 4416 2221 4420
rect 2225 4416 2230 4420
rect 2026 4415 2230 4416
rect 2030 4411 2036 4415
rect 2040 4411 2046 4415
rect 2050 4411 2056 4415
rect 2060 4411 2066 4415
rect 2070 4411 2186 4415
rect 2190 4411 2196 4415
rect 2200 4411 2206 4415
rect 2210 4411 2216 4415
rect 2220 4411 2226 4415
rect 2026 4410 2230 4411
rect 2026 4406 2031 4410
rect 2035 4406 2041 4410
rect 2045 4406 2051 4410
rect 2055 4406 2061 4410
rect 2065 4406 2191 4410
rect 2195 4406 2201 4410
rect 2205 4406 2211 4410
rect 2215 4406 2221 4410
rect 2225 4406 2230 4410
rect 2026 4405 2230 4406
rect 2030 4401 2036 4405
rect 2040 4401 2046 4405
rect 2050 4401 2056 4405
rect 2060 4401 2066 4405
rect 2070 4401 2186 4405
rect 2190 4401 2196 4405
rect 2200 4401 2206 4405
rect 2210 4401 2216 4405
rect 2220 4401 2226 4405
rect 2026 4400 2230 4401
rect 2026 4396 2031 4400
rect 2035 4396 2041 4400
rect 2045 4396 2051 4400
rect 2055 4396 2061 4400
rect 2065 4396 2191 4400
rect 2195 4396 2201 4400
rect 2205 4396 2211 4400
rect 2215 4396 2221 4400
rect 2225 4396 2230 4400
rect 2026 4395 2230 4396
rect 2030 4391 2036 4395
rect 2040 4391 2046 4395
rect 2050 4391 2056 4395
rect 2060 4391 2066 4395
rect 2070 4391 2186 4395
rect 2190 4391 2196 4395
rect 2200 4391 2206 4395
rect 2210 4391 2216 4395
rect 2220 4391 2226 4395
rect 2026 4390 2230 4391
rect 2026 4386 2031 4390
rect 2035 4386 2041 4390
rect 2045 4386 2051 4390
rect 2055 4386 2061 4390
rect 2065 4386 2191 4390
rect 2195 4386 2201 4390
rect 2205 4386 2211 4390
rect 2215 4386 2221 4390
rect 2225 4386 2230 4390
rect 2026 4385 2230 4386
rect 2030 4381 2036 4385
rect 2040 4381 2046 4385
rect 2050 4381 2056 4385
rect 2060 4381 2066 4385
rect 2070 4381 2186 4385
rect 2190 4381 2196 4385
rect 2200 4381 2206 4385
rect 2210 4381 2216 4385
rect 2220 4381 2226 4385
rect 2026 4380 2230 4381
rect 2026 4376 2031 4380
rect 2035 4376 2041 4380
rect 2045 4376 2051 4380
rect 2055 4376 2061 4380
rect 2065 4376 2191 4380
rect 2195 4376 2201 4380
rect 2205 4376 2211 4380
rect 2215 4376 2221 4380
rect 2225 4376 2230 4380
rect 2026 4375 2230 4376
rect 2030 4371 2036 4375
rect 2040 4371 2046 4375
rect 2050 4371 2056 4375
rect 2060 4371 2066 4375
rect 2070 4371 2186 4375
rect 2190 4371 2196 4375
rect 2200 4371 2206 4375
rect 2210 4371 2216 4375
rect 2220 4371 2226 4375
rect 2026 4370 2230 4371
rect 2026 4366 2031 4370
rect 2035 4366 2041 4370
rect 2045 4366 2051 4370
rect 2055 4366 2061 4370
rect 2065 4366 2191 4370
rect 2195 4366 2201 4370
rect 2205 4366 2211 4370
rect 2215 4366 2221 4370
rect 2225 4366 2230 4370
rect 2026 4365 2230 4366
rect 2030 4361 2036 4365
rect 2040 4361 2046 4365
rect 2050 4361 2056 4365
rect 2060 4361 2066 4365
rect 2070 4361 2186 4365
rect 2190 4361 2196 4365
rect 2200 4361 2206 4365
rect 2210 4361 2216 4365
rect 2220 4361 2226 4365
rect 2335 4446 2340 4450
rect 2344 4446 2350 4450
rect 2354 4446 2360 4450
rect 2364 4446 2370 4450
rect 2374 4446 2500 4450
rect 2504 4446 2510 4450
rect 2514 4446 2520 4450
rect 2524 4446 2530 4450
rect 2534 4446 2539 4450
rect 2335 4445 2539 4446
rect 2339 4441 2345 4445
rect 2349 4441 2355 4445
rect 2359 4441 2365 4445
rect 2369 4441 2375 4445
rect 2379 4441 2495 4445
rect 2499 4441 2505 4445
rect 2509 4441 2515 4445
rect 2519 4441 2525 4445
rect 2529 4441 2535 4445
rect 2335 4440 2539 4441
rect 2335 4436 2340 4440
rect 2344 4436 2350 4440
rect 2354 4436 2360 4440
rect 2364 4436 2370 4440
rect 2374 4436 2500 4440
rect 2504 4436 2510 4440
rect 2514 4436 2520 4440
rect 2524 4436 2530 4440
rect 2534 4436 2539 4440
rect 2335 4435 2539 4436
rect 2339 4431 2345 4435
rect 2349 4431 2355 4435
rect 2359 4431 2365 4435
rect 2369 4431 2375 4435
rect 2379 4431 2495 4435
rect 2499 4431 2505 4435
rect 2509 4431 2515 4435
rect 2519 4431 2525 4435
rect 2529 4431 2535 4435
rect 2335 4430 2539 4431
rect 2335 4426 2340 4430
rect 2344 4426 2350 4430
rect 2354 4426 2360 4430
rect 2364 4426 2370 4430
rect 2374 4426 2500 4430
rect 2504 4426 2510 4430
rect 2514 4426 2520 4430
rect 2524 4426 2530 4430
rect 2534 4426 2539 4430
rect 2335 4425 2539 4426
rect 2339 4421 2345 4425
rect 2349 4421 2355 4425
rect 2359 4421 2365 4425
rect 2369 4421 2375 4425
rect 2379 4421 2495 4425
rect 2499 4421 2505 4425
rect 2509 4421 2515 4425
rect 2519 4421 2525 4425
rect 2529 4421 2535 4425
rect 2335 4420 2539 4421
rect 2335 4416 2340 4420
rect 2344 4416 2350 4420
rect 2354 4416 2360 4420
rect 2364 4416 2370 4420
rect 2374 4416 2500 4420
rect 2504 4416 2510 4420
rect 2514 4416 2520 4420
rect 2524 4416 2530 4420
rect 2534 4416 2539 4420
rect 2335 4415 2539 4416
rect 2339 4411 2345 4415
rect 2349 4411 2355 4415
rect 2359 4411 2365 4415
rect 2369 4411 2375 4415
rect 2379 4411 2495 4415
rect 2499 4411 2505 4415
rect 2509 4411 2515 4415
rect 2519 4411 2525 4415
rect 2529 4411 2535 4415
rect 2335 4410 2539 4411
rect 2335 4406 2340 4410
rect 2344 4406 2350 4410
rect 2354 4406 2360 4410
rect 2364 4406 2370 4410
rect 2374 4406 2500 4410
rect 2504 4406 2510 4410
rect 2514 4406 2520 4410
rect 2524 4406 2530 4410
rect 2534 4406 2539 4410
rect 2335 4405 2539 4406
rect 2339 4401 2345 4405
rect 2349 4401 2355 4405
rect 2359 4401 2365 4405
rect 2369 4401 2375 4405
rect 2379 4401 2495 4405
rect 2499 4401 2505 4405
rect 2509 4401 2515 4405
rect 2519 4401 2525 4405
rect 2529 4401 2535 4405
rect 2335 4400 2539 4401
rect 2335 4396 2340 4400
rect 2344 4396 2350 4400
rect 2354 4396 2360 4400
rect 2364 4396 2370 4400
rect 2374 4396 2500 4400
rect 2504 4396 2510 4400
rect 2514 4396 2520 4400
rect 2524 4396 2530 4400
rect 2534 4396 2539 4400
rect 2335 4395 2539 4396
rect 2339 4391 2345 4395
rect 2349 4391 2355 4395
rect 2359 4391 2365 4395
rect 2369 4391 2375 4395
rect 2379 4391 2495 4395
rect 2499 4391 2505 4395
rect 2509 4391 2515 4395
rect 2519 4391 2525 4395
rect 2529 4391 2535 4395
rect 2335 4390 2539 4391
rect 2335 4386 2340 4390
rect 2344 4386 2350 4390
rect 2354 4386 2360 4390
rect 2364 4386 2370 4390
rect 2374 4386 2500 4390
rect 2504 4386 2510 4390
rect 2514 4386 2520 4390
rect 2524 4386 2530 4390
rect 2534 4386 2539 4390
rect 2335 4385 2539 4386
rect 2339 4381 2345 4385
rect 2349 4381 2355 4385
rect 2359 4381 2365 4385
rect 2369 4381 2375 4385
rect 2379 4381 2495 4385
rect 2499 4381 2505 4385
rect 2509 4381 2515 4385
rect 2519 4381 2525 4385
rect 2529 4381 2535 4385
rect 2335 4380 2539 4381
rect 2335 4376 2340 4380
rect 2344 4376 2350 4380
rect 2354 4376 2360 4380
rect 2364 4376 2370 4380
rect 2374 4376 2500 4380
rect 2504 4376 2510 4380
rect 2514 4376 2520 4380
rect 2524 4376 2530 4380
rect 2534 4376 2539 4380
rect 2335 4375 2539 4376
rect 2339 4371 2345 4375
rect 2349 4371 2355 4375
rect 2359 4371 2365 4375
rect 2369 4371 2375 4375
rect 2379 4371 2495 4375
rect 2499 4371 2505 4375
rect 2509 4371 2515 4375
rect 2519 4371 2525 4375
rect 2529 4371 2535 4375
rect 2335 4370 2539 4371
rect 2335 4366 2340 4370
rect 2344 4366 2350 4370
rect 2354 4366 2360 4370
rect 2364 4366 2370 4370
rect 2374 4366 2500 4370
rect 2504 4366 2510 4370
rect 2514 4366 2520 4370
rect 2524 4366 2530 4370
rect 2534 4366 2539 4370
rect 2335 4365 2539 4366
rect 2339 4361 2345 4365
rect 2349 4361 2355 4365
rect 2359 4361 2365 4365
rect 2369 4361 2375 4365
rect 2379 4361 2495 4365
rect 2499 4361 2505 4365
rect 2509 4361 2515 4365
rect 2519 4361 2525 4365
rect 2529 4361 2535 4365
rect 2644 4446 2649 4450
rect 2653 4446 2659 4450
rect 2663 4446 2669 4450
rect 2673 4446 2679 4450
rect 2683 4446 2809 4450
rect 2813 4446 2819 4450
rect 2823 4446 2829 4450
rect 2833 4446 2839 4450
rect 2843 4446 2848 4450
rect 2644 4445 2848 4446
rect 2648 4441 2654 4445
rect 2658 4441 2664 4445
rect 2668 4441 2674 4445
rect 2678 4441 2684 4445
rect 2688 4441 2804 4445
rect 2808 4441 2814 4445
rect 2818 4441 2824 4445
rect 2828 4441 2834 4445
rect 2838 4441 2844 4445
rect 2644 4440 2848 4441
rect 2644 4436 2649 4440
rect 2653 4436 2659 4440
rect 2663 4436 2669 4440
rect 2673 4436 2679 4440
rect 2683 4436 2809 4440
rect 2813 4436 2819 4440
rect 2823 4436 2829 4440
rect 2833 4436 2839 4440
rect 2843 4436 2848 4440
rect 2644 4435 2848 4436
rect 2648 4431 2654 4435
rect 2658 4431 2664 4435
rect 2668 4431 2674 4435
rect 2678 4431 2684 4435
rect 2688 4431 2804 4435
rect 2808 4431 2814 4435
rect 2818 4431 2824 4435
rect 2828 4431 2834 4435
rect 2838 4431 2844 4435
rect 2644 4430 2848 4431
rect 2644 4426 2649 4430
rect 2653 4426 2659 4430
rect 2663 4426 2669 4430
rect 2673 4426 2679 4430
rect 2683 4426 2809 4430
rect 2813 4426 2819 4430
rect 2823 4426 2829 4430
rect 2833 4426 2839 4430
rect 2843 4426 2848 4430
rect 2644 4425 2848 4426
rect 2648 4421 2654 4425
rect 2658 4421 2664 4425
rect 2668 4421 2674 4425
rect 2678 4421 2684 4425
rect 2688 4421 2804 4425
rect 2808 4421 2814 4425
rect 2818 4421 2824 4425
rect 2828 4421 2834 4425
rect 2838 4421 2844 4425
rect 2644 4420 2848 4421
rect 2644 4416 2649 4420
rect 2653 4416 2659 4420
rect 2663 4416 2669 4420
rect 2673 4416 2679 4420
rect 2683 4416 2809 4420
rect 2813 4416 2819 4420
rect 2823 4416 2829 4420
rect 2833 4416 2839 4420
rect 2843 4416 2848 4420
rect 2644 4415 2848 4416
rect 2648 4411 2654 4415
rect 2658 4411 2664 4415
rect 2668 4411 2674 4415
rect 2678 4411 2684 4415
rect 2688 4411 2804 4415
rect 2808 4411 2814 4415
rect 2818 4411 2824 4415
rect 2828 4411 2834 4415
rect 2838 4411 2844 4415
rect 2644 4410 2848 4411
rect 2644 4406 2649 4410
rect 2653 4406 2659 4410
rect 2663 4406 2669 4410
rect 2673 4406 2679 4410
rect 2683 4406 2809 4410
rect 2813 4406 2819 4410
rect 2823 4406 2829 4410
rect 2833 4406 2839 4410
rect 2843 4406 2848 4410
rect 2644 4405 2848 4406
rect 2648 4401 2654 4405
rect 2658 4401 2664 4405
rect 2668 4401 2674 4405
rect 2678 4401 2684 4405
rect 2688 4401 2804 4405
rect 2808 4401 2814 4405
rect 2818 4401 2824 4405
rect 2828 4401 2834 4405
rect 2838 4401 2844 4405
rect 2644 4400 2848 4401
rect 2644 4396 2649 4400
rect 2653 4396 2659 4400
rect 2663 4396 2669 4400
rect 2673 4396 2679 4400
rect 2683 4396 2809 4400
rect 2813 4396 2819 4400
rect 2823 4396 2829 4400
rect 2833 4396 2839 4400
rect 2843 4396 2848 4400
rect 2644 4395 2848 4396
rect 2648 4391 2654 4395
rect 2658 4391 2664 4395
rect 2668 4391 2674 4395
rect 2678 4391 2684 4395
rect 2688 4391 2804 4395
rect 2808 4391 2814 4395
rect 2818 4391 2824 4395
rect 2828 4391 2834 4395
rect 2838 4391 2844 4395
rect 2644 4390 2848 4391
rect 2644 4386 2649 4390
rect 2653 4386 2659 4390
rect 2663 4386 2669 4390
rect 2673 4386 2679 4390
rect 2683 4386 2809 4390
rect 2813 4386 2819 4390
rect 2823 4386 2829 4390
rect 2833 4386 2839 4390
rect 2843 4386 2848 4390
rect 2644 4385 2848 4386
rect 2648 4381 2654 4385
rect 2658 4381 2664 4385
rect 2668 4381 2674 4385
rect 2678 4381 2684 4385
rect 2688 4381 2804 4385
rect 2808 4381 2814 4385
rect 2818 4381 2824 4385
rect 2828 4381 2834 4385
rect 2838 4381 2844 4385
rect 2644 4380 2848 4381
rect 2644 4376 2649 4380
rect 2653 4376 2659 4380
rect 2663 4376 2669 4380
rect 2673 4376 2679 4380
rect 2683 4376 2809 4380
rect 2813 4376 2819 4380
rect 2823 4376 2829 4380
rect 2833 4376 2839 4380
rect 2843 4376 2848 4380
rect 2644 4375 2848 4376
rect 2648 4371 2654 4375
rect 2658 4371 2664 4375
rect 2668 4371 2674 4375
rect 2678 4371 2684 4375
rect 2688 4371 2804 4375
rect 2808 4371 2814 4375
rect 2818 4371 2824 4375
rect 2828 4371 2834 4375
rect 2838 4371 2844 4375
rect 2644 4370 2848 4371
rect 2644 4366 2649 4370
rect 2653 4366 2659 4370
rect 2663 4366 2669 4370
rect 2673 4366 2679 4370
rect 2683 4366 2809 4370
rect 2813 4366 2819 4370
rect 2823 4366 2829 4370
rect 2833 4366 2839 4370
rect 2843 4366 2848 4370
rect 2644 4365 2848 4366
rect 2648 4361 2654 4365
rect 2658 4361 2664 4365
rect 2668 4361 2674 4365
rect 2678 4361 2684 4365
rect 2688 4361 2804 4365
rect 2808 4361 2814 4365
rect 2818 4361 2824 4365
rect 2828 4361 2834 4365
rect 2838 4361 2844 4365
rect 2953 4446 2958 4450
rect 2962 4446 2968 4450
rect 2972 4446 2978 4450
rect 2982 4446 2988 4450
rect 2992 4446 3118 4450
rect 3122 4446 3128 4450
rect 3132 4446 3138 4450
rect 3142 4446 3148 4450
rect 3152 4446 3157 4450
rect 2953 4445 3157 4446
rect 2957 4441 2963 4445
rect 2967 4441 2973 4445
rect 2977 4441 2983 4445
rect 2987 4441 2993 4445
rect 2997 4441 3113 4445
rect 3117 4441 3123 4445
rect 3127 4441 3133 4445
rect 3137 4441 3143 4445
rect 3147 4441 3153 4445
rect 2953 4440 3157 4441
rect 2953 4436 2958 4440
rect 2962 4436 2968 4440
rect 2972 4436 2978 4440
rect 2982 4436 2988 4440
rect 2992 4436 3118 4440
rect 3122 4436 3128 4440
rect 3132 4436 3138 4440
rect 3142 4436 3148 4440
rect 3152 4436 3157 4440
rect 2953 4435 3157 4436
rect 2957 4431 2963 4435
rect 2967 4431 2973 4435
rect 2977 4431 2983 4435
rect 2987 4431 2993 4435
rect 2997 4431 3113 4435
rect 3117 4431 3123 4435
rect 3127 4431 3133 4435
rect 3137 4431 3143 4435
rect 3147 4431 3153 4435
rect 2953 4430 3157 4431
rect 2953 4426 2958 4430
rect 2962 4426 2968 4430
rect 2972 4426 2978 4430
rect 2982 4426 2988 4430
rect 2992 4426 3118 4430
rect 3122 4426 3128 4430
rect 3132 4426 3138 4430
rect 3142 4426 3148 4430
rect 3152 4426 3157 4430
rect 2953 4425 3157 4426
rect 2957 4421 2963 4425
rect 2967 4421 2973 4425
rect 2977 4421 2983 4425
rect 2987 4421 2993 4425
rect 2997 4421 3113 4425
rect 3117 4421 3123 4425
rect 3127 4421 3133 4425
rect 3137 4421 3143 4425
rect 3147 4421 3153 4425
rect 2953 4420 3157 4421
rect 2953 4416 2958 4420
rect 2962 4416 2968 4420
rect 2972 4416 2978 4420
rect 2982 4416 2988 4420
rect 2992 4416 3118 4420
rect 3122 4416 3128 4420
rect 3132 4416 3138 4420
rect 3142 4416 3148 4420
rect 3152 4416 3157 4420
rect 2953 4415 3157 4416
rect 2957 4411 2963 4415
rect 2967 4411 2973 4415
rect 2977 4411 2983 4415
rect 2987 4411 2993 4415
rect 2997 4411 3113 4415
rect 3117 4411 3123 4415
rect 3127 4411 3133 4415
rect 3137 4411 3143 4415
rect 3147 4411 3153 4415
rect 2953 4410 3157 4411
rect 2953 4406 2958 4410
rect 2962 4406 2968 4410
rect 2972 4406 2978 4410
rect 2982 4406 2988 4410
rect 2992 4406 3118 4410
rect 3122 4406 3128 4410
rect 3132 4406 3138 4410
rect 3142 4406 3148 4410
rect 3152 4406 3157 4410
rect 2953 4405 3157 4406
rect 2957 4401 2963 4405
rect 2967 4401 2973 4405
rect 2977 4401 2983 4405
rect 2987 4401 2993 4405
rect 2997 4401 3113 4405
rect 3117 4401 3123 4405
rect 3127 4401 3133 4405
rect 3137 4401 3143 4405
rect 3147 4401 3153 4405
rect 2953 4400 3157 4401
rect 2953 4396 2958 4400
rect 2962 4396 2968 4400
rect 2972 4396 2978 4400
rect 2982 4396 2988 4400
rect 2992 4396 3118 4400
rect 3122 4396 3128 4400
rect 3132 4396 3138 4400
rect 3142 4396 3148 4400
rect 3152 4396 3157 4400
rect 2953 4395 3157 4396
rect 2957 4391 2963 4395
rect 2967 4391 2973 4395
rect 2977 4391 2983 4395
rect 2987 4391 2993 4395
rect 2997 4391 3113 4395
rect 3117 4391 3123 4395
rect 3127 4391 3133 4395
rect 3137 4391 3143 4395
rect 3147 4391 3153 4395
rect 2953 4390 3157 4391
rect 2953 4386 2958 4390
rect 2962 4386 2968 4390
rect 2972 4386 2978 4390
rect 2982 4386 2988 4390
rect 2992 4386 3118 4390
rect 3122 4386 3128 4390
rect 3132 4386 3138 4390
rect 3142 4386 3148 4390
rect 3152 4386 3157 4390
rect 2953 4385 3157 4386
rect 2957 4381 2963 4385
rect 2967 4381 2973 4385
rect 2977 4381 2983 4385
rect 2987 4381 2993 4385
rect 2997 4381 3113 4385
rect 3117 4381 3123 4385
rect 3127 4381 3133 4385
rect 3137 4381 3143 4385
rect 3147 4381 3153 4385
rect 2953 4380 3157 4381
rect 2953 4376 2958 4380
rect 2962 4376 2968 4380
rect 2972 4376 2978 4380
rect 2982 4376 2988 4380
rect 2992 4376 3118 4380
rect 3122 4376 3128 4380
rect 3132 4376 3138 4380
rect 3142 4376 3148 4380
rect 3152 4376 3157 4380
rect 2953 4375 3157 4376
rect 2957 4371 2963 4375
rect 2967 4371 2973 4375
rect 2977 4371 2983 4375
rect 2987 4371 2993 4375
rect 2997 4371 3113 4375
rect 3117 4371 3123 4375
rect 3127 4371 3133 4375
rect 3137 4371 3143 4375
rect 3147 4371 3153 4375
rect 2953 4370 3157 4371
rect 2953 4366 2958 4370
rect 2962 4366 2968 4370
rect 2972 4366 2978 4370
rect 2982 4366 2988 4370
rect 2992 4366 3118 4370
rect 3122 4366 3128 4370
rect 3132 4366 3138 4370
rect 3142 4366 3148 4370
rect 3152 4366 3157 4370
rect 2953 4365 3157 4366
rect 2957 4361 2963 4365
rect 2967 4361 2973 4365
rect 2977 4361 2983 4365
rect 2987 4361 2993 4365
rect 2997 4361 3113 4365
rect 3117 4361 3123 4365
rect 3127 4361 3133 4365
rect 3137 4361 3143 4365
rect 3147 4361 3153 4365
rect 3262 4446 3267 4450
rect 3271 4446 3277 4450
rect 3281 4446 3287 4450
rect 3291 4446 3297 4450
rect 3301 4446 3427 4450
rect 3431 4446 3437 4450
rect 3441 4446 3447 4450
rect 3451 4446 3457 4450
rect 3461 4446 3466 4450
rect 3262 4445 3466 4446
rect 3266 4441 3272 4445
rect 3276 4441 3282 4445
rect 3286 4441 3292 4445
rect 3296 4441 3302 4445
rect 3306 4441 3422 4445
rect 3426 4441 3432 4445
rect 3436 4441 3442 4445
rect 3446 4441 3452 4445
rect 3456 4441 3462 4445
rect 3262 4440 3466 4441
rect 3262 4436 3267 4440
rect 3271 4436 3277 4440
rect 3281 4436 3287 4440
rect 3291 4436 3297 4440
rect 3301 4436 3427 4440
rect 3431 4436 3437 4440
rect 3441 4436 3447 4440
rect 3451 4436 3457 4440
rect 3461 4436 3466 4440
rect 3262 4435 3466 4436
rect 3266 4431 3272 4435
rect 3276 4431 3282 4435
rect 3286 4431 3292 4435
rect 3296 4431 3302 4435
rect 3306 4431 3422 4435
rect 3426 4431 3432 4435
rect 3436 4431 3442 4435
rect 3446 4431 3452 4435
rect 3456 4431 3462 4435
rect 3262 4430 3466 4431
rect 3262 4426 3267 4430
rect 3271 4426 3277 4430
rect 3281 4426 3287 4430
rect 3291 4426 3297 4430
rect 3301 4426 3427 4430
rect 3431 4426 3437 4430
rect 3441 4426 3447 4430
rect 3451 4426 3457 4430
rect 3461 4426 3466 4430
rect 3262 4425 3466 4426
rect 3266 4421 3272 4425
rect 3276 4421 3282 4425
rect 3286 4421 3292 4425
rect 3296 4421 3302 4425
rect 3306 4421 3422 4425
rect 3426 4421 3432 4425
rect 3436 4421 3442 4425
rect 3446 4421 3452 4425
rect 3456 4421 3462 4425
rect 3262 4420 3466 4421
rect 3262 4416 3267 4420
rect 3271 4416 3277 4420
rect 3281 4416 3287 4420
rect 3291 4416 3297 4420
rect 3301 4416 3427 4420
rect 3431 4416 3437 4420
rect 3441 4416 3447 4420
rect 3451 4416 3457 4420
rect 3461 4416 3466 4420
rect 3262 4415 3466 4416
rect 3266 4411 3272 4415
rect 3276 4411 3282 4415
rect 3286 4411 3292 4415
rect 3296 4411 3302 4415
rect 3306 4411 3422 4415
rect 3426 4411 3432 4415
rect 3436 4411 3442 4415
rect 3446 4411 3452 4415
rect 3456 4411 3462 4415
rect 3262 4410 3466 4411
rect 3262 4406 3267 4410
rect 3271 4406 3277 4410
rect 3281 4406 3287 4410
rect 3291 4406 3297 4410
rect 3301 4406 3427 4410
rect 3431 4406 3437 4410
rect 3441 4406 3447 4410
rect 3451 4406 3457 4410
rect 3461 4406 3466 4410
rect 3262 4405 3466 4406
rect 3266 4401 3272 4405
rect 3276 4401 3282 4405
rect 3286 4401 3292 4405
rect 3296 4401 3302 4405
rect 3306 4401 3422 4405
rect 3426 4401 3432 4405
rect 3436 4401 3442 4405
rect 3446 4401 3452 4405
rect 3456 4401 3462 4405
rect 3262 4400 3466 4401
rect 3262 4396 3267 4400
rect 3271 4396 3277 4400
rect 3281 4396 3287 4400
rect 3291 4396 3297 4400
rect 3301 4396 3427 4400
rect 3431 4396 3437 4400
rect 3441 4396 3447 4400
rect 3451 4396 3457 4400
rect 3461 4396 3466 4400
rect 3262 4395 3466 4396
rect 3266 4391 3272 4395
rect 3276 4391 3282 4395
rect 3286 4391 3292 4395
rect 3296 4391 3302 4395
rect 3306 4391 3422 4395
rect 3426 4391 3432 4395
rect 3436 4391 3442 4395
rect 3446 4391 3452 4395
rect 3456 4391 3462 4395
rect 3262 4390 3466 4391
rect 3262 4386 3267 4390
rect 3271 4386 3277 4390
rect 3281 4386 3287 4390
rect 3291 4386 3297 4390
rect 3301 4386 3427 4390
rect 3431 4386 3437 4390
rect 3441 4386 3447 4390
rect 3451 4386 3457 4390
rect 3461 4386 3466 4390
rect 3262 4385 3466 4386
rect 3266 4381 3272 4385
rect 3276 4381 3282 4385
rect 3286 4381 3292 4385
rect 3296 4381 3302 4385
rect 3306 4381 3422 4385
rect 3426 4381 3432 4385
rect 3436 4381 3442 4385
rect 3446 4381 3452 4385
rect 3456 4381 3462 4385
rect 3262 4380 3466 4381
rect 3262 4376 3267 4380
rect 3271 4376 3277 4380
rect 3281 4376 3287 4380
rect 3291 4376 3297 4380
rect 3301 4376 3427 4380
rect 3431 4376 3437 4380
rect 3441 4376 3447 4380
rect 3451 4376 3457 4380
rect 3461 4376 3466 4380
rect 3262 4375 3466 4376
rect 3266 4371 3272 4375
rect 3276 4371 3282 4375
rect 3286 4371 3292 4375
rect 3296 4371 3302 4375
rect 3306 4371 3422 4375
rect 3426 4371 3432 4375
rect 3436 4371 3442 4375
rect 3446 4371 3452 4375
rect 3456 4371 3462 4375
rect 3262 4370 3466 4371
rect 3262 4366 3267 4370
rect 3271 4366 3277 4370
rect 3281 4366 3287 4370
rect 3291 4366 3297 4370
rect 3301 4366 3427 4370
rect 3431 4366 3437 4370
rect 3441 4366 3447 4370
rect 3451 4366 3457 4370
rect 3461 4366 3466 4370
rect 3262 4365 3466 4366
rect 3266 4361 3272 4365
rect 3276 4361 3282 4365
rect 3286 4361 3292 4365
rect 3296 4361 3302 4365
rect 3306 4361 3422 4365
rect 3426 4361 3432 4365
rect 3436 4361 3442 4365
rect 3446 4361 3452 4365
rect 3456 4361 3462 4365
rect 3571 4446 3576 4450
rect 3580 4446 3586 4450
rect 3590 4446 3596 4450
rect 3600 4446 3606 4450
rect 3610 4446 3736 4450
rect 3740 4446 3746 4450
rect 3750 4446 3756 4450
rect 3760 4446 3766 4450
rect 3770 4446 3775 4450
rect 3571 4445 3775 4446
rect 3575 4441 3581 4445
rect 3585 4441 3591 4445
rect 3595 4441 3601 4445
rect 3605 4441 3611 4445
rect 3615 4441 3731 4445
rect 3735 4441 3741 4445
rect 3745 4441 3751 4445
rect 3755 4441 3761 4445
rect 3765 4441 3771 4445
rect 3571 4440 3775 4441
rect 3571 4436 3576 4440
rect 3580 4436 3586 4440
rect 3590 4436 3596 4440
rect 3600 4436 3606 4440
rect 3610 4436 3736 4440
rect 3740 4436 3746 4440
rect 3750 4436 3756 4440
rect 3760 4436 3766 4440
rect 3770 4436 3775 4440
rect 3571 4435 3775 4436
rect 3575 4431 3581 4435
rect 3585 4431 3591 4435
rect 3595 4431 3601 4435
rect 3605 4431 3611 4435
rect 3615 4431 3731 4435
rect 3735 4431 3741 4435
rect 3745 4431 3751 4435
rect 3755 4431 3761 4435
rect 3765 4431 3771 4435
rect 3571 4430 3775 4431
rect 3571 4426 3576 4430
rect 3580 4426 3586 4430
rect 3590 4426 3596 4430
rect 3600 4426 3606 4430
rect 3610 4426 3736 4430
rect 3740 4426 3746 4430
rect 3750 4426 3756 4430
rect 3760 4426 3766 4430
rect 3770 4426 3775 4430
rect 3571 4425 3775 4426
rect 3575 4421 3581 4425
rect 3585 4421 3591 4425
rect 3595 4421 3601 4425
rect 3605 4421 3611 4425
rect 3615 4421 3731 4425
rect 3735 4421 3741 4425
rect 3745 4421 3751 4425
rect 3755 4421 3761 4425
rect 3765 4421 3771 4425
rect 3571 4420 3775 4421
rect 3571 4416 3576 4420
rect 3580 4416 3586 4420
rect 3590 4416 3596 4420
rect 3600 4416 3606 4420
rect 3610 4416 3736 4420
rect 3740 4416 3746 4420
rect 3750 4416 3756 4420
rect 3760 4416 3766 4420
rect 3770 4416 3775 4420
rect 3571 4415 3775 4416
rect 3575 4411 3581 4415
rect 3585 4411 3591 4415
rect 3595 4411 3601 4415
rect 3605 4411 3611 4415
rect 3615 4411 3731 4415
rect 3735 4411 3741 4415
rect 3745 4411 3751 4415
rect 3755 4411 3761 4415
rect 3765 4411 3771 4415
rect 3571 4410 3775 4411
rect 3571 4406 3576 4410
rect 3580 4406 3586 4410
rect 3590 4406 3596 4410
rect 3600 4406 3606 4410
rect 3610 4406 3736 4410
rect 3740 4406 3746 4410
rect 3750 4406 3756 4410
rect 3760 4406 3766 4410
rect 3770 4406 3775 4410
rect 3571 4405 3775 4406
rect 3575 4401 3581 4405
rect 3585 4401 3591 4405
rect 3595 4401 3601 4405
rect 3605 4401 3611 4405
rect 3615 4401 3731 4405
rect 3735 4401 3741 4405
rect 3745 4401 3751 4405
rect 3755 4401 3761 4405
rect 3765 4401 3771 4405
rect 3571 4400 3775 4401
rect 3571 4396 3576 4400
rect 3580 4396 3586 4400
rect 3590 4396 3596 4400
rect 3600 4396 3606 4400
rect 3610 4396 3736 4400
rect 3740 4396 3746 4400
rect 3750 4396 3756 4400
rect 3760 4396 3766 4400
rect 3770 4396 3775 4400
rect 3571 4395 3775 4396
rect 3575 4391 3581 4395
rect 3585 4391 3591 4395
rect 3595 4391 3601 4395
rect 3605 4391 3611 4395
rect 3615 4391 3731 4395
rect 3735 4391 3741 4395
rect 3745 4391 3751 4395
rect 3755 4391 3761 4395
rect 3765 4391 3771 4395
rect 3571 4390 3775 4391
rect 3571 4386 3576 4390
rect 3580 4386 3586 4390
rect 3590 4386 3596 4390
rect 3600 4386 3606 4390
rect 3610 4386 3736 4390
rect 3740 4386 3746 4390
rect 3750 4386 3756 4390
rect 3760 4386 3766 4390
rect 3770 4386 3775 4390
rect 3571 4385 3775 4386
rect 3575 4381 3581 4385
rect 3585 4381 3591 4385
rect 3595 4381 3601 4385
rect 3605 4381 3611 4385
rect 3615 4381 3731 4385
rect 3735 4381 3741 4385
rect 3745 4381 3751 4385
rect 3755 4381 3761 4385
rect 3765 4381 3771 4385
rect 3571 4380 3775 4381
rect 3571 4376 3576 4380
rect 3580 4376 3586 4380
rect 3590 4376 3596 4380
rect 3600 4376 3606 4380
rect 3610 4376 3736 4380
rect 3740 4376 3746 4380
rect 3750 4376 3756 4380
rect 3760 4376 3766 4380
rect 3770 4376 3775 4380
rect 3571 4375 3775 4376
rect 3575 4371 3581 4375
rect 3585 4371 3591 4375
rect 3595 4371 3601 4375
rect 3605 4371 3611 4375
rect 3615 4371 3731 4375
rect 3735 4371 3741 4375
rect 3745 4371 3751 4375
rect 3755 4371 3761 4375
rect 3765 4371 3771 4375
rect 3571 4370 3775 4371
rect 3571 4366 3576 4370
rect 3580 4366 3586 4370
rect 3590 4366 3596 4370
rect 3600 4366 3606 4370
rect 3610 4366 3736 4370
rect 3740 4366 3746 4370
rect 3750 4366 3756 4370
rect 3760 4366 3766 4370
rect 3770 4366 3775 4370
rect 3571 4365 3775 4366
rect 3575 4361 3581 4365
rect 3585 4361 3591 4365
rect 3595 4361 3601 4365
rect 3605 4361 3611 4365
rect 3615 4361 3731 4365
rect 3735 4361 3741 4365
rect 3745 4361 3751 4365
rect 3755 4361 3761 4365
rect 3765 4361 3771 4365
rect 1153 4332 1249 4361
rect 1153 4328 1158 4332
rect 1162 4328 1165 4332
rect 1169 4328 1172 4332
rect 1176 4328 1179 4332
rect 1183 4328 1186 4332
rect 1190 4328 1193 4332
rect 1197 4328 1200 4332
rect 1204 4328 1207 4332
rect 1211 4328 1214 4332
rect 1218 4328 1221 4332
rect 1225 4328 1228 4332
rect 1232 4328 1235 4332
rect 1239 4328 1242 4332
rect 1246 4328 1249 4332
rect 1153 4327 1249 4328
rect 1153 4323 1158 4327
rect 1162 4323 1165 4327
rect 1169 4323 1172 4327
rect 1176 4323 1179 4327
rect 1183 4323 1186 4327
rect 1190 4323 1193 4327
rect 1197 4323 1200 4327
rect 1204 4323 1207 4327
rect 1211 4323 1214 4327
rect 1218 4323 1221 4327
rect 1225 4323 1228 4327
rect 1232 4323 1235 4327
rect 1239 4323 1242 4327
rect 1246 4323 1249 4327
rect 1153 4322 1249 4323
rect 1153 4321 1158 4322
rect 1143 4318 1158 4321
rect 1162 4318 1165 4322
rect 1169 4318 1172 4322
rect 1176 4318 1179 4322
rect 1183 4318 1186 4322
rect 1190 4318 1193 4322
rect 1197 4318 1200 4322
rect 1204 4318 1207 4322
rect 1211 4318 1214 4322
rect 1218 4318 1221 4322
rect 1225 4318 1228 4322
rect 1232 4318 1235 4322
rect 1239 4318 1242 4322
rect 1246 4321 1249 4322
rect 1462 4332 1558 4361
rect 1462 4328 1467 4332
rect 1471 4328 1474 4332
rect 1478 4328 1481 4332
rect 1485 4328 1488 4332
rect 1492 4328 1495 4332
rect 1499 4328 1502 4332
rect 1506 4328 1509 4332
rect 1513 4328 1516 4332
rect 1520 4328 1523 4332
rect 1527 4328 1530 4332
rect 1534 4328 1537 4332
rect 1541 4328 1544 4332
rect 1548 4328 1551 4332
rect 1555 4328 1558 4332
rect 1462 4327 1558 4328
rect 1462 4323 1467 4327
rect 1471 4323 1474 4327
rect 1478 4323 1481 4327
rect 1485 4323 1488 4327
rect 1492 4323 1495 4327
rect 1499 4323 1502 4327
rect 1506 4323 1509 4327
rect 1513 4323 1516 4327
rect 1520 4323 1523 4327
rect 1527 4323 1530 4327
rect 1534 4323 1537 4327
rect 1541 4323 1544 4327
rect 1548 4323 1551 4327
rect 1555 4323 1558 4327
rect 1462 4322 1558 4323
rect 1462 4321 1467 4322
rect 1246 4318 1259 4321
rect 1143 4317 1259 4318
rect 1143 4313 1158 4317
rect 1162 4313 1165 4317
rect 1169 4313 1172 4317
rect 1176 4313 1179 4317
rect 1183 4313 1186 4317
rect 1190 4313 1193 4317
rect 1197 4313 1200 4317
rect 1204 4313 1207 4317
rect 1211 4313 1214 4317
rect 1218 4313 1221 4317
rect 1225 4313 1228 4317
rect 1232 4313 1235 4317
rect 1239 4313 1242 4317
rect 1246 4313 1259 4317
rect 1143 4312 1259 4313
rect 1452 4318 1467 4321
rect 1471 4318 1474 4322
rect 1478 4318 1481 4322
rect 1485 4318 1488 4322
rect 1492 4318 1495 4322
rect 1499 4318 1502 4322
rect 1506 4318 1509 4322
rect 1513 4318 1516 4322
rect 1520 4318 1523 4322
rect 1527 4318 1530 4322
rect 1534 4318 1537 4322
rect 1541 4318 1544 4322
rect 1548 4318 1551 4322
rect 1555 4321 1558 4322
rect 1771 4332 1867 4361
rect 1771 4328 1776 4332
rect 1780 4328 1783 4332
rect 1787 4328 1790 4332
rect 1794 4328 1797 4332
rect 1801 4328 1804 4332
rect 1808 4328 1811 4332
rect 1815 4328 1818 4332
rect 1822 4328 1825 4332
rect 1829 4328 1832 4332
rect 1836 4328 1839 4332
rect 1843 4328 1846 4332
rect 1850 4328 1853 4332
rect 1857 4328 1860 4332
rect 1864 4328 1867 4332
rect 1771 4327 1867 4328
rect 1771 4323 1776 4327
rect 1780 4323 1783 4327
rect 1787 4323 1790 4327
rect 1794 4323 1797 4327
rect 1801 4323 1804 4327
rect 1808 4323 1811 4327
rect 1815 4323 1818 4327
rect 1822 4323 1825 4327
rect 1829 4323 1832 4327
rect 1836 4323 1839 4327
rect 1843 4323 1846 4327
rect 1850 4323 1853 4327
rect 1857 4323 1860 4327
rect 1864 4323 1867 4327
rect 1771 4322 1867 4323
rect 1771 4321 1776 4322
rect 1555 4318 1568 4321
rect 1452 4317 1568 4318
rect 1452 4313 1467 4317
rect 1471 4313 1474 4317
rect 1478 4313 1481 4317
rect 1485 4313 1488 4317
rect 1492 4313 1495 4317
rect 1499 4313 1502 4317
rect 1506 4313 1509 4317
rect 1513 4313 1516 4317
rect 1520 4313 1523 4317
rect 1527 4313 1530 4317
rect 1534 4313 1537 4317
rect 1541 4313 1544 4317
rect 1548 4313 1551 4317
rect 1555 4313 1568 4317
rect 1452 4312 1568 4313
rect 1761 4318 1776 4321
rect 1780 4318 1783 4322
rect 1787 4318 1790 4322
rect 1794 4318 1797 4322
rect 1801 4318 1804 4322
rect 1808 4318 1811 4322
rect 1815 4318 1818 4322
rect 1822 4318 1825 4322
rect 1829 4318 1832 4322
rect 1836 4318 1839 4322
rect 1843 4318 1846 4322
rect 1850 4318 1853 4322
rect 1857 4318 1860 4322
rect 1864 4321 1867 4322
rect 2080 4332 2176 4361
rect 2080 4328 2085 4332
rect 2089 4328 2092 4332
rect 2096 4328 2099 4332
rect 2103 4328 2106 4332
rect 2110 4328 2113 4332
rect 2117 4328 2120 4332
rect 2124 4328 2127 4332
rect 2131 4328 2134 4332
rect 2138 4328 2141 4332
rect 2145 4328 2148 4332
rect 2152 4328 2155 4332
rect 2159 4328 2162 4332
rect 2166 4328 2169 4332
rect 2173 4328 2176 4332
rect 2080 4327 2176 4328
rect 2080 4323 2085 4327
rect 2089 4323 2092 4327
rect 2096 4323 2099 4327
rect 2103 4323 2106 4327
rect 2110 4323 2113 4327
rect 2117 4323 2120 4327
rect 2124 4323 2127 4327
rect 2131 4323 2134 4327
rect 2138 4323 2141 4327
rect 2145 4323 2148 4327
rect 2152 4323 2155 4327
rect 2159 4323 2162 4327
rect 2166 4323 2169 4327
rect 2173 4323 2176 4327
rect 2080 4322 2176 4323
rect 2080 4321 2085 4322
rect 1864 4318 1877 4321
rect 1761 4317 1877 4318
rect 1761 4313 1776 4317
rect 1780 4313 1783 4317
rect 1787 4313 1790 4317
rect 1794 4313 1797 4317
rect 1801 4313 1804 4317
rect 1808 4313 1811 4317
rect 1815 4313 1818 4317
rect 1822 4313 1825 4317
rect 1829 4313 1832 4317
rect 1836 4313 1839 4317
rect 1843 4313 1846 4317
rect 1850 4313 1853 4317
rect 1857 4313 1860 4317
rect 1864 4313 1877 4317
rect 1761 4312 1877 4313
rect 2070 4318 2085 4321
rect 2089 4318 2092 4322
rect 2096 4318 2099 4322
rect 2103 4318 2106 4322
rect 2110 4318 2113 4322
rect 2117 4318 2120 4322
rect 2124 4318 2127 4322
rect 2131 4318 2134 4322
rect 2138 4318 2141 4322
rect 2145 4318 2148 4322
rect 2152 4318 2155 4322
rect 2159 4318 2162 4322
rect 2166 4318 2169 4322
rect 2173 4321 2176 4322
rect 2389 4332 2485 4361
rect 2389 4328 2394 4332
rect 2398 4328 2401 4332
rect 2405 4328 2408 4332
rect 2412 4328 2415 4332
rect 2419 4328 2422 4332
rect 2426 4328 2429 4332
rect 2433 4328 2436 4332
rect 2440 4328 2443 4332
rect 2447 4328 2450 4332
rect 2454 4328 2457 4332
rect 2461 4328 2464 4332
rect 2468 4328 2471 4332
rect 2475 4328 2478 4332
rect 2482 4328 2485 4332
rect 2389 4327 2485 4328
rect 2389 4323 2394 4327
rect 2398 4323 2401 4327
rect 2405 4323 2408 4327
rect 2412 4323 2415 4327
rect 2419 4323 2422 4327
rect 2426 4323 2429 4327
rect 2433 4323 2436 4327
rect 2440 4323 2443 4327
rect 2447 4323 2450 4327
rect 2454 4323 2457 4327
rect 2461 4323 2464 4327
rect 2468 4323 2471 4327
rect 2475 4323 2478 4327
rect 2482 4323 2485 4327
rect 2389 4322 2485 4323
rect 2389 4321 2394 4322
rect 2173 4318 2186 4321
rect 2070 4317 2186 4318
rect 2070 4313 2085 4317
rect 2089 4313 2092 4317
rect 2096 4313 2099 4317
rect 2103 4313 2106 4317
rect 2110 4313 2113 4317
rect 2117 4313 2120 4317
rect 2124 4313 2127 4317
rect 2131 4313 2134 4317
rect 2138 4313 2141 4317
rect 2145 4313 2148 4317
rect 2152 4313 2155 4317
rect 2159 4313 2162 4317
rect 2166 4313 2169 4317
rect 2173 4313 2186 4317
rect 2070 4312 2186 4313
rect 2379 4318 2394 4321
rect 2398 4318 2401 4322
rect 2405 4318 2408 4322
rect 2412 4318 2415 4322
rect 2419 4318 2422 4322
rect 2426 4318 2429 4322
rect 2433 4318 2436 4322
rect 2440 4318 2443 4322
rect 2447 4318 2450 4322
rect 2454 4318 2457 4322
rect 2461 4318 2464 4322
rect 2468 4318 2471 4322
rect 2475 4318 2478 4322
rect 2482 4321 2485 4322
rect 2698 4332 2794 4361
rect 2698 4328 2703 4332
rect 2707 4328 2710 4332
rect 2714 4328 2717 4332
rect 2721 4328 2724 4332
rect 2728 4328 2731 4332
rect 2735 4328 2738 4332
rect 2742 4328 2745 4332
rect 2749 4328 2752 4332
rect 2756 4328 2759 4332
rect 2763 4328 2766 4332
rect 2770 4328 2773 4332
rect 2777 4328 2780 4332
rect 2784 4328 2787 4332
rect 2791 4328 2794 4332
rect 2698 4327 2794 4328
rect 2698 4323 2703 4327
rect 2707 4323 2710 4327
rect 2714 4323 2717 4327
rect 2721 4323 2724 4327
rect 2728 4323 2731 4327
rect 2735 4323 2738 4327
rect 2742 4323 2745 4327
rect 2749 4323 2752 4327
rect 2756 4323 2759 4327
rect 2763 4323 2766 4327
rect 2770 4323 2773 4327
rect 2777 4323 2780 4327
rect 2784 4323 2787 4327
rect 2791 4323 2794 4327
rect 2698 4322 2794 4323
rect 2698 4321 2703 4322
rect 2482 4318 2495 4321
rect 2379 4317 2495 4318
rect 2379 4313 2394 4317
rect 2398 4313 2401 4317
rect 2405 4313 2408 4317
rect 2412 4313 2415 4317
rect 2419 4313 2422 4317
rect 2426 4313 2429 4317
rect 2433 4313 2436 4317
rect 2440 4313 2443 4317
rect 2447 4313 2450 4317
rect 2454 4313 2457 4317
rect 2461 4313 2464 4317
rect 2468 4313 2471 4317
rect 2475 4313 2478 4317
rect 2482 4313 2495 4317
rect 2379 4312 2495 4313
rect 2688 4318 2703 4321
rect 2707 4318 2710 4322
rect 2714 4318 2717 4322
rect 2721 4318 2724 4322
rect 2728 4318 2731 4322
rect 2735 4318 2738 4322
rect 2742 4318 2745 4322
rect 2749 4318 2752 4322
rect 2756 4318 2759 4322
rect 2763 4318 2766 4322
rect 2770 4318 2773 4322
rect 2777 4318 2780 4322
rect 2784 4318 2787 4322
rect 2791 4321 2794 4322
rect 3007 4332 3103 4361
rect 3007 4328 3012 4332
rect 3016 4328 3019 4332
rect 3023 4328 3026 4332
rect 3030 4328 3033 4332
rect 3037 4328 3040 4332
rect 3044 4328 3047 4332
rect 3051 4328 3054 4332
rect 3058 4328 3061 4332
rect 3065 4328 3068 4332
rect 3072 4328 3075 4332
rect 3079 4328 3082 4332
rect 3086 4328 3089 4332
rect 3093 4328 3096 4332
rect 3100 4328 3103 4332
rect 3007 4327 3103 4328
rect 3007 4323 3012 4327
rect 3016 4323 3019 4327
rect 3023 4323 3026 4327
rect 3030 4323 3033 4327
rect 3037 4323 3040 4327
rect 3044 4323 3047 4327
rect 3051 4323 3054 4327
rect 3058 4323 3061 4327
rect 3065 4323 3068 4327
rect 3072 4323 3075 4327
rect 3079 4323 3082 4327
rect 3086 4323 3089 4327
rect 3093 4323 3096 4327
rect 3100 4323 3103 4327
rect 3007 4322 3103 4323
rect 3007 4321 3012 4322
rect 2791 4318 2804 4321
rect 2688 4317 2804 4318
rect 2688 4313 2703 4317
rect 2707 4313 2710 4317
rect 2714 4313 2717 4317
rect 2721 4313 2724 4317
rect 2728 4313 2731 4317
rect 2735 4313 2738 4317
rect 2742 4313 2745 4317
rect 2749 4313 2752 4317
rect 2756 4313 2759 4317
rect 2763 4313 2766 4317
rect 2770 4313 2773 4317
rect 2777 4313 2780 4317
rect 2784 4313 2787 4317
rect 2791 4313 2804 4317
rect 2688 4312 2804 4313
rect 2997 4318 3012 4321
rect 3016 4318 3019 4322
rect 3023 4318 3026 4322
rect 3030 4318 3033 4322
rect 3037 4318 3040 4322
rect 3044 4318 3047 4322
rect 3051 4318 3054 4322
rect 3058 4318 3061 4322
rect 3065 4318 3068 4322
rect 3072 4318 3075 4322
rect 3079 4318 3082 4322
rect 3086 4318 3089 4322
rect 3093 4318 3096 4322
rect 3100 4321 3103 4322
rect 3316 4332 3412 4361
rect 3316 4328 3321 4332
rect 3325 4328 3328 4332
rect 3332 4328 3335 4332
rect 3339 4328 3342 4332
rect 3346 4328 3349 4332
rect 3353 4328 3356 4332
rect 3360 4328 3363 4332
rect 3367 4328 3370 4332
rect 3374 4328 3377 4332
rect 3381 4328 3384 4332
rect 3388 4328 3391 4332
rect 3395 4328 3398 4332
rect 3402 4328 3405 4332
rect 3409 4328 3412 4332
rect 3316 4327 3412 4328
rect 3316 4323 3321 4327
rect 3325 4323 3328 4327
rect 3332 4323 3335 4327
rect 3339 4323 3342 4327
rect 3346 4323 3349 4327
rect 3353 4323 3356 4327
rect 3360 4323 3363 4327
rect 3367 4323 3370 4327
rect 3374 4323 3377 4327
rect 3381 4323 3384 4327
rect 3388 4323 3391 4327
rect 3395 4323 3398 4327
rect 3402 4323 3405 4327
rect 3409 4323 3412 4327
rect 3316 4322 3412 4323
rect 3316 4321 3321 4322
rect 3100 4318 3113 4321
rect 2997 4317 3113 4318
rect 2997 4313 3012 4317
rect 3016 4313 3019 4317
rect 3023 4313 3026 4317
rect 3030 4313 3033 4317
rect 3037 4313 3040 4317
rect 3044 4313 3047 4317
rect 3051 4313 3054 4317
rect 3058 4313 3061 4317
rect 3065 4313 3068 4317
rect 3072 4313 3075 4317
rect 3079 4313 3082 4317
rect 3086 4313 3089 4317
rect 3093 4313 3096 4317
rect 3100 4313 3113 4317
rect 2997 4312 3113 4313
rect 3306 4318 3321 4321
rect 3325 4318 3328 4322
rect 3332 4318 3335 4322
rect 3339 4318 3342 4322
rect 3346 4318 3349 4322
rect 3353 4318 3356 4322
rect 3360 4318 3363 4322
rect 3367 4318 3370 4322
rect 3374 4318 3377 4322
rect 3381 4318 3384 4322
rect 3388 4318 3391 4322
rect 3395 4318 3398 4322
rect 3402 4318 3405 4322
rect 3409 4321 3412 4322
rect 3625 4332 3721 4361
rect 3625 4328 3630 4332
rect 3634 4328 3637 4332
rect 3641 4328 3644 4332
rect 3648 4328 3651 4332
rect 3655 4328 3658 4332
rect 3662 4328 3665 4332
rect 3669 4328 3672 4332
rect 3676 4328 3679 4332
rect 3683 4328 3686 4332
rect 3690 4328 3693 4332
rect 3697 4328 3700 4332
rect 3704 4328 3707 4332
rect 3711 4328 3714 4332
rect 3718 4328 3721 4332
rect 3625 4327 3721 4328
rect 3625 4323 3630 4327
rect 3634 4323 3637 4327
rect 3641 4323 3644 4327
rect 3648 4323 3651 4327
rect 3655 4323 3658 4327
rect 3662 4323 3665 4327
rect 3669 4323 3672 4327
rect 3676 4323 3679 4327
rect 3683 4323 3686 4327
rect 3690 4323 3693 4327
rect 3697 4323 3700 4327
rect 3704 4323 3707 4327
rect 3711 4323 3714 4327
rect 3718 4323 3721 4327
rect 3625 4322 3721 4323
rect 3625 4321 3630 4322
rect 3409 4318 3422 4321
rect 3306 4317 3422 4318
rect 3306 4313 3321 4317
rect 3325 4313 3328 4317
rect 3332 4313 3335 4317
rect 3339 4313 3342 4317
rect 3346 4313 3349 4317
rect 3353 4313 3356 4317
rect 3360 4313 3363 4317
rect 3367 4313 3370 4317
rect 3374 4313 3377 4317
rect 3381 4313 3384 4317
rect 3388 4313 3391 4317
rect 3395 4313 3398 4317
rect 3402 4313 3405 4317
rect 3409 4313 3422 4317
rect 3306 4312 3422 4313
rect 3615 4318 3630 4321
rect 3634 4318 3637 4322
rect 3641 4318 3644 4322
rect 3648 4318 3651 4322
rect 3655 4318 3658 4322
rect 3662 4318 3665 4322
rect 3669 4318 3672 4322
rect 3676 4318 3679 4322
rect 3683 4318 3686 4322
rect 3690 4318 3693 4322
rect 3697 4318 3700 4322
rect 3704 4318 3707 4322
rect 3711 4318 3714 4322
rect 3718 4321 3721 4322
rect 3718 4318 3731 4321
rect 3615 4317 3731 4318
rect 3615 4313 3630 4317
rect 3634 4313 3637 4317
rect 3641 4313 3644 4317
rect 3648 4313 3651 4317
rect 3655 4313 3658 4317
rect 3662 4313 3665 4317
rect 3669 4313 3672 4317
rect 3676 4313 3679 4317
rect 3683 4313 3686 4317
rect 3690 4313 3693 4317
rect 3697 4313 3700 4317
rect 3704 4313 3707 4317
rect 3711 4313 3714 4317
rect 3718 4313 3731 4317
rect 3615 4312 3731 4313
rect 1071 4278 1331 4281
rect 1071 4024 1074 4278
rect 1328 4024 1331 4278
rect 1071 4021 1331 4024
rect 1380 4278 1640 4281
rect 1380 4024 1383 4278
rect 1637 4024 1640 4278
rect 1380 4021 1640 4024
rect 1689 4278 1949 4281
rect 1689 4024 1692 4278
rect 1946 4024 1949 4278
rect 1689 4021 1949 4024
rect 1998 4278 2258 4281
rect 1998 4024 2001 4278
rect 2255 4024 2258 4278
rect 1998 4021 2258 4024
rect 2307 4278 2567 4281
rect 2307 4024 2310 4278
rect 2564 4024 2567 4278
rect 2307 4021 2567 4024
rect 2616 4278 2876 4281
rect 2616 4024 2619 4278
rect 2873 4024 2876 4278
rect 2616 4021 2876 4024
rect 2925 4278 3185 4281
rect 2925 4024 2928 4278
rect 3182 4024 3185 4278
rect 2925 4021 3185 4024
rect 3234 4278 3494 4281
rect 3234 4024 3237 4278
rect 3491 4024 3494 4278
rect 3234 4021 3494 4024
rect 3543 4278 3803 4281
rect 3543 4024 3546 4278
rect 3800 4024 3803 4278
rect 3543 4021 3803 4024
rect 3852 4278 4112 4281
rect 3852 4024 3855 4278
rect 4109 4024 4112 4278
rect 4148 4034 5054 4528
rect 3852 4021 4112 4024
<< m3contact >>
rect 1354 9796 1358 9800
rect 1359 9796 1363 9800
rect 1354 9791 1358 9795
rect 1359 9791 1363 9795
rect 1354 9786 1358 9790
rect 1359 9786 1363 9790
rect 1354 9781 1358 9785
rect 1359 9781 1363 9785
rect 1354 9776 1358 9780
rect 1359 9776 1363 9780
rect 1354 9771 1358 9775
rect 1359 9771 1363 9775
rect 1354 9766 1358 9770
rect 1359 9766 1363 9770
rect 802 9762 806 9766
rect 807 9762 811 9766
rect 812 9762 816 9766
rect 817 9762 821 9766
rect 802 9752 806 9756
rect 807 9752 811 9756
rect 812 9752 816 9756
rect 817 9752 821 9756
rect 802 9742 806 9746
rect 807 9742 811 9746
rect 812 9742 816 9746
rect 817 9742 821 9746
rect 802 9732 806 9736
rect 807 9732 811 9736
rect 812 9732 816 9736
rect 817 9732 821 9736
rect 831 9762 835 9766
rect 836 9762 840 9766
rect 841 9762 845 9766
rect 846 9762 850 9766
rect 831 9752 835 9756
rect 836 9752 840 9756
rect 841 9752 845 9756
rect 846 9752 850 9756
rect 831 9742 835 9746
rect 836 9742 840 9746
rect 841 9742 845 9746
rect 846 9742 850 9746
rect 831 9732 835 9736
rect 836 9732 840 9736
rect 841 9732 845 9736
rect 846 9732 850 9736
rect 860 9762 864 9766
rect 865 9762 869 9766
rect 870 9762 874 9766
rect 875 9762 879 9766
rect 860 9752 864 9756
rect 865 9752 869 9756
rect 870 9752 874 9756
rect 875 9752 879 9756
rect 860 9742 864 9746
rect 865 9742 869 9746
rect 870 9742 874 9746
rect 875 9742 879 9746
rect 860 9732 864 9736
rect 865 9732 869 9736
rect 870 9732 874 9736
rect 875 9732 879 9736
rect 889 9762 893 9766
rect 894 9762 898 9766
rect 899 9762 903 9766
rect 904 9762 908 9766
rect 889 9752 893 9756
rect 894 9752 898 9756
rect 899 9752 903 9756
rect 904 9752 908 9756
rect 889 9742 893 9746
rect 894 9742 898 9746
rect 899 9742 903 9746
rect 904 9742 908 9746
rect 889 9732 893 9736
rect 894 9732 898 9736
rect 899 9732 903 9736
rect 904 9732 908 9736
rect 918 9762 922 9766
rect 923 9762 927 9766
rect 928 9762 932 9766
rect 933 9762 937 9766
rect 918 9752 922 9756
rect 923 9752 927 9756
rect 928 9752 932 9756
rect 933 9752 937 9756
rect 918 9742 922 9746
rect 923 9742 927 9746
rect 928 9742 932 9746
rect 933 9742 937 9746
rect 918 9732 922 9736
rect 923 9732 927 9736
rect 928 9732 932 9736
rect 933 9732 937 9736
rect 1319 9762 1323 9766
rect 1324 9762 1328 9766
rect 1329 9762 1333 9766
rect 1334 9762 1338 9766
rect 1319 9752 1323 9756
rect 1324 9752 1328 9756
rect 1329 9752 1333 9756
rect 1334 9752 1338 9756
rect 1319 9742 1323 9746
rect 1324 9742 1328 9746
rect 1329 9742 1333 9746
rect 1334 9742 1338 9746
rect 1319 9732 1323 9736
rect 1324 9732 1328 9736
rect 1329 9732 1333 9736
rect 1334 9732 1338 9736
rect 1354 9761 1358 9765
rect 1359 9761 1363 9765
rect 1354 9756 1358 9760
rect 1359 9756 1363 9760
rect 1354 9751 1358 9755
rect 1359 9751 1363 9755
rect 1354 9746 1358 9750
rect 1359 9746 1363 9750
rect 1354 9741 1358 9745
rect 1359 9741 1363 9745
rect 1354 9736 1358 9740
rect 1359 9736 1363 9740
rect 802 9716 806 9720
rect 807 9716 811 9720
rect 812 9716 816 9720
rect 817 9716 821 9720
rect 802 9706 806 9710
rect 807 9706 811 9710
rect 812 9706 816 9710
rect 817 9706 821 9710
rect 802 9696 806 9700
rect 807 9696 811 9700
rect 812 9696 816 9700
rect 817 9696 821 9700
rect 802 9686 806 9690
rect 807 9686 811 9690
rect 812 9686 816 9690
rect 817 9686 821 9690
rect 831 9716 835 9720
rect 836 9716 840 9720
rect 841 9716 845 9720
rect 846 9716 850 9720
rect 831 9706 835 9710
rect 836 9706 840 9710
rect 841 9706 845 9710
rect 846 9706 850 9710
rect 831 9696 835 9700
rect 836 9696 840 9700
rect 841 9696 845 9700
rect 846 9696 850 9700
rect 831 9686 835 9690
rect 836 9686 840 9690
rect 841 9686 845 9690
rect 846 9686 850 9690
rect 860 9716 864 9720
rect 865 9716 869 9720
rect 870 9716 874 9720
rect 875 9716 879 9720
rect 860 9706 864 9710
rect 865 9706 869 9710
rect 870 9706 874 9710
rect 875 9706 879 9710
rect 860 9696 864 9700
rect 865 9696 869 9700
rect 870 9696 874 9700
rect 875 9696 879 9700
rect 860 9686 864 9690
rect 865 9686 869 9690
rect 870 9686 874 9690
rect 875 9686 879 9690
rect 889 9716 893 9720
rect 894 9716 898 9720
rect 899 9716 903 9720
rect 904 9716 908 9720
rect 889 9706 893 9710
rect 894 9706 898 9710
rect 899 9706 903 9710
rect 904 9706 908 9710
rect 889 9696 893 9700
rect 894 9696 898 9700
rect 899 9696 903 9700
rect 904 9696 908 9700
rect 889 9686 893 9690
rect 894 9686 898 9690
rect 899 9686 903 9690
rect 904 9686 908 9690
rect 918 9716 922 9720
rect 923 9716 927 9720
rect 928 9716 932 9720
rect 933 9716 937 9720
rect 918 9706 922 9710
rect 923 9706 927 9710
rect 928 9706 932 9710
rect 933 9706 937 9710
rect 918 9696 922 9700
rect 923 9696 927 9700
rect 928 9696 932 9700
rect 933 9696 937 9700
rect 918 9686 922 9690
rect 923 9686 927 9690
rect 928 9686 932 9690
rect 933 9686 937 9690
rect 1319 9716 1323 9720
rect 1324 9716 1328 9720
rect 1329 9716 1333 9720
rect 1334 9716 1338 9720
rect 1319 9706 1323 9710
rect 1324 9706 1328 9710
rect 1329 9706 1333 9710
rect 1334 9706 1338 9710
rect 1547 9765 1551 9769
rect 1552 9765 1556 9769
rect 1557 9765 1561 9769
rect 1562 9765 1566 9769
rect 1567 9765 1571 9769
rect 1572 9765 1576 9769
rect 1577 9765 1581 9769
rect 1582 9765 1586 9769
rect 1587 9765 1591 9769
rect 1592 9765 1596 9769
rect 1597 9765 1601 9769
rect 1602 9765 1606 9769
rect 1607 9765 1611 9769
rect 1663 9796 1667 9800
rect 1668 9796 1672 9800
rect 1663 9791 1667 9795
rect 1668 9791 1672 9795
rect 1663 9786 1667 9790
rect 1668 9786 1672 9790
rect 1663 9781 1667 9785
rect 1668 9781 1672 9785
rect 1663 9776 1667 9780
rect 1668 9776 1672 9780
rect 1663 9771 1667 9775
rect 1668 9771 1672 9775
rect 1663 9766 1667 9770
rect 1668 9766 1672 9770
rect 1547 9760 1551 9764
rect 1552 9760 1556 9764
rect 1557 9760 1561 9764
rect 1562 9760 1566 9764
rect 1567 9760 1571 9764
rect 1572 9760 1576 9764
rect 1577 9760 1581 9764
rect 1582 9760 1586 9764
rect 1587 9760 1591 9764
rect 1592 9760 1596 9764
rect 1597 9760 1601 9764
rect 1602 9760 1606 9764
rect 1607 9760 1611 9764
rect 1628 9762 1632 9766
rect 1633 9762 1637 9766
rect 1638 9762 1642 9766
rect 1643 9762 1647 9766
rect 1628 9752 1632 9756
rect 1633 9752 1637 9756
rect 1638 9752 1642 9756
rect 1643 9752 1647 9756
rect 1628 9742 1632 9746
rect 1633 9742 1637 9746
rect 1638 9742 1642 9746
rect 1643 9742 1647 9746
rect 1628 9732 1632 9736
rect 1633 9732 1637 9736
rect 1638 9732 1642 9736
rect 1643 9732 1647 9736
rect 1663 9761 1667 9765
rect 1668 9761 1672 9765
rect 1663 9756 1667 9760
rect 1668 9756 1672 9760
rect 1663 9751 1667 9755
rect 1668 9751 1672 9755
rect 1663 9746 1667 9750
rect 1668 9746 1672 9750
rect 1663 9741 1667 9745
rect 1668 9741 1672 9745
rect 1663 9736 1667 9740
rect 1668 9736 1672 9740
rect 1387 9708 1391 9712
rect 1392 9708 1396 9712
rect 1397 9708 1401 9712
rect 1402 9708 1406 9712
rect 1407 9708 1411 9712
rect 1412 9708 1416 9712
rect 1417 9708 1421 9712
rect 1422 9708 1426 9712
rect 1427 9708 1431 9712
rect 1432 9708 1436 9712
rect 1437 9708 1441 9712
rect 1442 9708 1446 9712
rect 1447 9708 1451 9712
rect 1387 9703 1391 9707
rect 1392 9703 1396 9707
rect 1397 9703 1401 9707
rect 1402 9703 1406 9707
rect 1407 9703 1411 9707
rect 1412 9703 1416 9707
rect 1417 9703 1421 9707
rect 1422 9703 1426 9707
rect 1427 9703 1431 9707
rect 1432 9703 1436 9707
rect 1437 9703 1441 9707
rect 1442 9703 1446 9707
rect 1447 9703 1451 9707
rect 1489 9711 1493 9715
rect 1494 9711 1498 9715
rect 1489 9706 1493 9710
rect 1494 9706 1498 9710
rect 1489 9701 1493 9705
rect 1494 9701 1498 9705
rect 1569 9708 1573 9712
rect 1574 9708 1578 9712
rect 1579 9708 1583 9712
rect 1584 9708 1588 9712
rect 1589 9708 1593 9712
rect 1594 9708 1598 9712
rect 1599 9708 1603 9712
rect 1604 9708 1608 9712
rect 1609 9708 1613 9712
rect 1614 9708 1618 9712
rect 1619 9708 1623 9712
rect 1569 9703 1573 9707
rect 1574 9703 1578 9707
rect 1579 9703 1583 9707
rect 1584 9703 1588 9707
rect 1589 9703 1593 9707
rect 1594 9703 1598 9707
rect 1599 9703 1603 9707
rect 1604 9703 1608 9707
rect 1609 9703 1613 9707
rect 1614 9703 1618 9707
rect 1619 9703 1623 9707
rect 1628 9716 1632 9720
rect 1633 9716 1637 9720
rect 1638 9716 1642 9720
rect 1643 9716 1647 9720
rect 1628 9706 1632 9710
rect 1633 9706 1637 9710
rect 1638 9706 1642 9710
rect 1643 9706 1647 9710
rect 1319 9696 1323 9700
rect 1324 9696 1328 9700
rect 1329 9696 1333 9700
rect 1334 9696 1338 9700
rect 1319 9686 1323 9690
rect 1324 9686 1328 9690
rect 1329 9686 1333 9690
rect 1334 9686 1338 9690
rect 1489 9696 1493 9700
rect 1494 9696 1498 9700
rect 1489 9691 1493 9695
rect 1494 9691 1498 9695
rect 1489 9686 1493 9690
rect 1494 9686 1498 9690
rect 1856 9765 1860 9769
rect 1861 9765 1865 9769
rect 1866 9765 1870 9769
rect 1871 9765 1875 9769
rect 1876 9765 1880 9769
rect 1881 9765 1885 9769
rect 1886 9765 1890 9769
rect 1891 9765 1895 9769
rect 1896 9765 1900 9769
rect 1901 9765 1905 9769
rect 1906 9765 1910 9769
rect 1911 9765 1915 9769
rect 1916 9765 1920 9769
rect 1972 9796 1976 9800
rect 1977 9796 1981 9800
rect 1972 9791 1976 9795
rect 1977 9791 1981 9795
rect 1972 9786 1976 9790
rect 1977 9786 1981 9790
rect 1972 9781 1976 9785
rect 1977 9781 1981 9785
rect 1972 9776 1976 9780
rect 1977 9776 1981 9780
rect 1972 9771 1976 9775
rect 1977 9771 1981 9775
rect 1972 9766 1976 9770
rect 1977 9766 1981 9770
rect 1856 9760 1860 9764
rect 1861 9760 1865 9764
rect 1866 9760 1870 9764
rect 1871 9760 1875 9764
rect 1876 9760 1880 9764
rect 1881 9760 1885 9764
rect 1886 9760 1890 9764
rect 1891 9760 1895 9764
rect 1896 9760 1900 9764
rect 1901 9760 1905 9764
rect 1906 9760 1910 9764
rect 1911 9760 1915 9764
rect 1916 9760 1920 9764
rect 1937 9762 1941 9766
rect 1942 9762 1946 9766
rect 1947 9762 1951 9766
rect 1952 9762 1956 9766
rect 1937 9752 1941 9756
rect 1942 9752 1946 9756
rect 1947 9752 1951 9756
rect 1952 9752 1956 9756
rect 1937 9742 1941 9746
rect 1942 9742 1946 9746
rect 1947 9742 1951 9746
rect 1952 9742 1956 9746
rect 1937 9732 1941 9736
rect 1942 9732 1946 9736
rect 1947 9732 1951 9736
rect 1952 9732 1956 9736
rect 1972 9761 1976 9765
rect 1977 9761 1981 9765
rect 1972 9756 1976 9760
rect 1977 9756 1981 9760
rect 1972 9751 1976 9755
rect 1977 9751 1981 9755
rect 1972 9746 1976 9750
rect 1977 9746 1981 9750
rect 1972 9741 1976 9745
rect 1977 9741 1981 9745
rect 1972 9736 1976 9740
rect 1977 9736 1981 9740
rect 1696 9708 1700 9712
rect 1701 9708 1705 9712
rect 1706 9708 1710 9712
rect 1711 9708 1715 9712
rect 1716 9708 1720 9712
rect 1721 9708 1725 9712
rect 1726 9708 1730 9712
rect 1731 9708 1735 9712
rect 1736 9708 1740 9712
rect 1741 9708 1745 9712
rect 1746 9708 1750 9712
rect 1751 9708 1755 9712
rect 1756 9708 1760 9712
rect 1696 9703 1700 9707
rect 1701 9703 1705 9707
rect 1706 9703 1710 9707
rect 1711 9703 1715 9707
rect 1716 9703 1720 9707
rect 1721 9703 1725 9707
rect 1726 9703 1730 9707
rect 1731 9703 1735 9707
rect 1736 9703 1740 9707
rect 1741 9703 1745 9707
rect 1746 9703 1750 9707
rect 1751 9703 1755 9707
rect 1756 9703 1760 9707
rect 1878 9708 1882 9712
rect 1883 9708 1887 9712
rect 1888 9708 1892 9712
rect 1893 9708 1897 9712
rect 1898 9708 1902 9712
rect 1903 9708 1907 9712
rect 1908 9708 1912 9712
rect 1913 9708 1917 9712
rect 1918 9708 1922 9712
rect 1923 9708 1927 9712
rect 1928 9708 1932 9712
rect 1878 9703 1882 9707
rect 1883 9703 1887 9707
rect 1888 9703 1892 9707
rect 1893 9703 1897 9707
rect 1898 9703 1902 9707
rect 1903 9703 1907 9707
rect 1908 9703 1912 9707
rect 1913 9703 1917 9707
rect 1918 9703 1922 9707
rect 1923 9703 1927 9707
rect 1928 9703 1932 9707
rect 1937 9716 1941 9720
rect 1942 9716 1946 9720
rect 1947 9716 1951 9720
rect 1952 9716 1956 9720
rect 1937 9706 1941 9710
rect 1942 9706 1946 9710
rect 1947 9706 1951 9710
rect 1952 9706 1956 9710
rect 2165 9765 2169 9769
rect 2170 9765 2174 9769
rect 2175 9765 2179 9769
rect 2180 9765 2184 9769
rect 2185 9765 2189 9769
rect 2190 9765 2194 9769
rect 2195 9765 2199 9769
rect 2200 9765 2204 9769
rect 2205 9765 2209 9769
rect 2210 9765 2214 9769
rect 2215 9765 2219 9769
rect 2220 9765 2224 9769
rect 2225 9765 2229 9769
rect 2281 9796 2285 9800
rect 2286 9796 2290 9800
rect 2281 9791 2285 9795
rect 2286 9791 2290 9795
rect 2281 9786 2285 9790
rect 2286 9786 2290 9790
rect 2281 9781 2285 9785
rect 2286 9781 2290 9785
rect 2281 9776 2285 9780
rect 2286 9776 2290 9780
rect 2281 9771 2285 9775
rect 2286 9771 2290 9775
rect 2281 9766 2285 9770
rect 2286 9766 2290 9770
rect 2165 9760 2169 9764
rect 2170 9760 2174 9764
rect 2175 9760 2179 9764
rect 2180 9760 2184 9764
rect 2185 9760 2189 9764
rect 2190 9760 2194 9764
rect 2195 9760 2199 9764
rect 2200 9760 2204 9764
rect 2205 9760 2209 9764
rect 2210 9760 2214 9764
rect 2215 9760 2219 9764
rect 2220 9760 2224 9764
rect 2225 9760 2229 9764
rect 2246 9762 2250 9766
rect 2251 9762 2255 9766
rect 2256 9762 2260 9766
rect 2261 9762 2265 9766
rect 2246 9752 2250 9756
rect 2251 9752 2255 9756
rect 2256 9752 2260 9756
rect 2261 9752 2265 9756
rect 2005 9708 2009 9712
rect 2010 9708 2014 9712
rect 2015 9708 2019 9712
rect 2020 9708 2024 9712
rect 2025 9708 2029 9712
rect 2030 9708 2034 9712
rect 2035 9708 2039 9712
rect 2040 9708 2044 9712
rect 2045 9708 2049 9712
rect 2050 9708 2054 9712
rect 2055 9708 2059 9712
rect 2060 9708 2064 9712
rect 2065 9708 2069 9712
rect 2005 9703 2009 9707
rect 2010 9703 2014 9707
rect 2015 9703 2019 9707
rect 2020 9703 2024 9707
rect 2025 9703 2029 9707
rect 2030 9703 2034 9707
rect 2035 9703 2039 9707
rect 2040 9703 2044 9707
rect 2045 9703 2049 9707
rect 2050 9703 2054 9707
rect 2055 9703 2059 9707
rect 2060 9703 2064 9707
rect 2065 9703 2069 9707
rect 2167 9736 2172 9741
rect 1628 9696 1632 9700
rect 1633 9696 1637 9700
rect 1638 9696 1642 9700
rect 1643 9696 1647 9700
rect 1628 9686 1632 9690
rect 1633 9686 1637 9690
rect 1638 9686 1642 9690
rect 1643 9686 1647 9690
rect 1937 9696 1941 9700
rect 1942 9696 1946 9700
rect 1947 9696 1951 9700
rect 1952 9696 1956 9700
rect 1937 9686 1941 9690
rect 1942 9686 1946 9690
rect 1947 9686 1951 9690
rect 1952 9686 1956 9690
rect 1489 9681 1493 9685
rect 1494 9681 1498 9685
rect 1489 9676 1493 9680
rect 1494 9676 1498 9680
rect 1489 9671 1493 9675
rect 1494 9671 1498 9675
rect 1489 9666 1493 9670
rect 1494 9666 1498 9670
rect 1489 9661 1493 9665
rect 1494 9661 1498 9665
rect 2246 9742 2250 9746
rect 2251 9742 2255 9746
rect 2256 9742 2260 9746
rect 2261 9742 2265 9746
rect 2246 9732 2250 9736
rect 2251 9732 2255 9736
rect 2256 9732 2260 9736
rect 2261 9732 2265 9736
rect 2281 9761 2285 9765
rect 2286 9761 2290 9765
rect 2281 9756 2285 9760
rect 2286 9756 2290 9760
rect 2281 9751 2285 9755
rect 2286 9751 2290 9755
rect 2281 9746 2285 9750
rect 2286 9746 2290 9750
rect 2281 9741 2285 9745
rect 2286 9741 2290 9745
rect 2281 9736 2285 9740
rect 2286 9736 2290 9740
rect 2187 9708 2191 9712
rect 2192 9708 2196 9712
rect 2197 9708 2201 9712
rect 2202 9708 2206 9712
rect 2207 9708 2211 9712
rect 2212 9708 2216 9712
rect 2217 9708 2221 9712
rect 2222 9708 2226 9712
rect 2227 9708 2231 9712
rect 2232 9708 2236 9712
rect 2237 9708 2241 9712
rect 2187 9703 2191 9707
rect 2192 9703 2196 9707
rect 2197 9703 2201 9707
rect 2202 9703 2206 9707
rect 2207 9703 2211 9707
rect 2212 9703 2216 9707
rect 2217 9703 2221 9707
rect 2222 9703 2226 9707
rect 2227 9703 2231 9707
rect 2232 9703 2236 9707
rect 2237 9703 2241 9707
rect 2246 9716 2250 9720
rect 2251 9716 2255 9720
rect 2256 9716 2260 9720
rect 2261 9716 2265 9720
rect 2246 9706 2250 9710
rect 2251 9706 2255 9710
rect 2256 9706 2260 9710
rect 2261 9706 2265 9710
rect 2474 9765 2478 9769
rect 2479 9765 2483 9769
rect 2484 9765 2488 9769
rect 2489 9765 2493 9769
rect 2494 9765 2498 9769
rect 2499 9765 2503 9769
rect 2504 9765 2508 9769
rect 2509 9765 2513 9769
rect 2514 9765 2518 9769
rect 2519 9765 2523 9769
rect 2524 9765 2528 9769
rect 2529 9765 2533 9769
rect 2534 9765 2538 9769
rect 2590 9796 2594 9800
rect 2595 9796 2599 9800
rect 2590 9791 2594 9795
rect 2595 9791 2599 9795
rect 2590 9786 2594 9790
rect 2595 9786 2599 9790
rect 2590 9781 2594 9785
rect 2595 9781 2599 9785
rect 2590 9776 2594 9780
rect 2595 9776 2599 9780
rect 2590 9771 2594 9775
rect 2595 9771 2599 9775
rect 2590 9766 2594 9770
rect 2595 9766 2599 9770
rect 2474 9760 2478 9764
rect 2479 9760 2483 9764
rect 2484 9760 2488 9764
rect 2489 9760 2493 9764
rect 2494 9760 2498 9764
rect 2499 9760 2503 9764
rect 2504 9760 2508 9764
rect 2509 9760 2513 9764
rect 2514 9760 2518 9764
rect 2519 9760 2523 9764
rect 2524 9760 2528 9764
rect 2529 9760 2533 9764
rect 2534 9760 2538 9764
rect 2555 9762 2559 9766
rect 2560 9762 2564 9766
rect 2565 9762 2569 9766
rect 2570 9762 2574 9766
rect 2555 9752 2559 9756
rect 2560 9752 2564 9756
rect 2565 9752 2569 9756
rect 2570 9752 2574 9756
rect 2555 9742 2559 9746
rect 2560 9742 2564 9746
rect 2565 9742 2569 9746
rect 2570 9742 2574 9746
rect 2555 9732 2559 9736
rect 2560 9732 2564 9736
rect 2565 9732 2569 9736
rect 2570 9732 2574 9736
rect 2590 9761 2594 9765
rect 2595 9761 2599 9765
rect 2590 9756 2594 9760
rect 2595 9756 2599 9760
rect 2590 9751 2594 9755
rect 2595 9751 2599 9755
rect 2590 9746 2594 9750
rect 2595 9746 2599 9750
rect 2590 9741 2594 9745
rect 2595 9741 2599 9745
rect 2590 9736 2594 9740
rect 2595 9736 2599 9740
rect 2314 9708 2318 9712
rect 2319 9708 2323 9712
rect 2324 9708 2328 9712
rect 2329 9708 2333 9712
rect 2334 9708 2338 9712
rect 2339 9708 2343 9712
rect 2344 9708 2348 9712
rect 2349 9708 2353 9712
rect 2354 9708 2358 9712
rect 2359 9708 2363 9712
rect 2364 9708 2368 9712
rect 2369 9708 2373 9712
rect 2374 9708 2378 9712
rect 2314 9703 2318 9707
rect 2319 9703 2323 9707
rect 2324 9703 2328 9707
rect 2329 9703 2333 9707
rect 2334 9703 2338 9707
rect 2339 9703 2343 9707
rect 2344 9703 2348 9707
rect 2349 9703 2353 9707
rect 2354 9703 2358 9707
rect 2359 9703 2363 9707
rect 2364 9703 2368 9707
rect 2369 9703 2373 9707
rect 2374 9703 2378 9707
rect 2496 9708 2500 9712
rect 2501 9708 2505 9712
rect 2506 9708 2510 9712
rect 2511 9708 2515 9712
rect 2516 9708 2520 9712
rect 2521 9708 2525 9712
rect 2526 9708 2530 9712
rect 2531 9708 2535 9712
rect 2536 9708 2540 9712
rect 2541 9708 2545 9712
rect 2546 9708 2550 9712
rect 2496 9703 2500 9707
rect 2501 9703 2505 9707
rect 2506 9703 2510 9707
rect 2511 9703 2515 9707
rect 2516 9703 2520 9707
rect 2521 9703 2525 9707
rect 2526 9703 2530 9707
rect 2531 9703 2535 9707
rect 2536 9703 2540 9707
rect 2541 9703 2545 9707
rect 2546 9703 2550 9707
rect 2555 9716 2559 9720
rect 2560 9716 2564 9720
rect 2565 9716 2569 9720
rect 2570 9716 2574 9720
rect 2555 9706 2559 9710
rect 2560 9706 2564 9710
rect 2565 9706 2569 9710
rect 2570 9706 2574 9710
rect 2783 9765 2787 9769
rect 2788 9765 2792 9769
rect 2793 9765 2797 9769
rect 2798 9765 2802 9769
rect 2803 9765 2807 9769
rect 2808 9765 2812 9769
rect 2813 9765 2817 9769
rect 2818 9765 2822 9769
rect 2823 9765 2827 9769
rect 2828 9765 2832 9769
rect 2833 9765 2837 9769
rect 2838 9765 2842 9769
rect 2843 9765 2847 9769
rect 2899 9796 2903 9800
rect 2904 9796 2908 9800
rect 2899 9791 2903 9795
rect 2904 9791 2908 9795
rect 2899 9786 2903 9790
rect 2904 9786 2908 9790
rect 2899 9781 2903 9785
rect 2904 9781 2908 9785
rect 2899 9776 2903 9780
rect 2904 9776 2908 9780
rect 2899 9771 2903 9775
rect 2904 9771 2908 9775
rect 2899 9766 2903 9770
rect 2904 9766 2908 9770
rect 2783 9760 2787 9764
rect 2788 9760 2792 9764
rect 2793 9760 2797 9764
rect 2798 9760 2802 9764
rect 2803 9760 2807 9764
rect 2808 9760 2812 9764
rect 2813 9760 2817 9764
rect 2818 9760 2822 9764
rect 2823 9760 2827 9764
rect 2828 9760 2832 9764
rect 2833 9760 2837 9764
rect 2838 9760 2842 9764
rect 2843 9760 2847 9764
rect 2864 9762 2868 9766
rect 2869 9762 2873 9766
rect 2874 9762 2878 9766
rect 2879 9762 2883 9766
rect 2864 9752 2868 9756
rect 2869 9752 2873 9756
rect 2874 9752 2878 9756
rect 2879 9752 2883 9756
rect 2864 9742 2868 9746
rect 2869 9742 2873 9746
rect 2874 9742 2878 9746
rect 2879 9742 2883 9746
rect 2864 9732 2868 9736
rect 2869 9732 2873 9736
rect 2874 9732 2878 9736
rect 2879 9732 2883 9736
rect 2899 9761 2903 9765
rect 2904 9761 2908 9765
rect 2899 9756 2903 9760
rect 2904 9756 2908 9760
rect 2899 9751 2903 9755
rect 2904 9751 2908 9755
rect 2899 9746 2903 9750
rect 2904 9746 2908 9750
rect 2899 9741 2903 9745
rect 2904 9741 2908 9745
rect 2899 9736 2903 9740
rect 2904 9736 2908 9740
rect 2623 9708 2627 9712
rect 2628 9708 2632 9712
rect 2633 9708 2637 9712
rect 2638 9708 2642 9712
rect 2643 9708 2647 9712
rect 2648 9708 2652 9712
rect 2653 9708 2657 9712
rect 2658 9708 2662 9712
rect 2663 9708 2667 9712
rect 2668 9708 2672 9712
rect 2673 9708 2677 9712
rect 2678 9708 2682 9712
rect 2683 9708 2687 9712
rect 2623 9703 2627 9707
rect 2628 9703 2632 9707
rect 2633 9703 2637 9707
rect 2638 9703 2642 9707
rect 2643 9703 2647 9707
rect 2648 9703 2652 9707
rect 2653 9703 2657 9707
rect 2658 9703 2662 9707
rect 2663 9703 2667 9707
rect 2668 9703 2672 9707
rect 2673 9703 2677 9707
rect 2678 9703 2682 9707
rect 2683 9703 2687 9707
rect 2805 9708 2809 9712
rect 2810 9708 2814 9712
rect 2815 9708 2819 9712
rect 2820 9708 2824 9712
rect 2825 9708 2829 9712
rect 2830 9708 2834 9712
rect 2835 9708 2839 9712
rect 2840 9708 2844 9712
rect 2845 9708 2849 9712
rect 2850 9708 2854 9712
rect 2855 9708 2859 9712
rect 2805 9703 2809 9707
rect 2810 9703 2814 9707
rect 2815 9703 2819 9707
rect 2820 9703 2824 9707
rect 2825 9703 2829 9707
rect 2830 9703 2834 9707
rect 2835 9703 2839 9707
rect 2840 9703 2844 9707
rect 2845 9703 2849 9707
rect 2850 9703 2854 9707
rect 2855 9703 2859 9707
rect 2864 9716 2868 9720
rect 2869 9716 2873 9720
rect 2874 9716 2878 9720
rect 2879 9716 2883 9720
rect 2864 9706 2868 9710
rect 2869 9706 2873 9710
rect 2874 9706 2878 9710
rect 2879 9706 2883 9710
rect 3092 9765 3096 9769
rect 3097 9765 3101 9769
rect 3102 9765 3106 9769
rect 3107 9765 3111 9769
rect 3112 9765 3116 9769
rect 3117 9765 3121 9769
rect 3122 9765 3126 9769
rect 3127 9765 3131 9769
rect 3132 9765 3136 9769
rect 3137 9765 3141 9769
rect 3142 9765 3146 9769
rect 3147 9765 3151 9769
rect 3152 9765 3156 9769
rect 3208 9796 3212 9800
rect 3213 9796 3217 9800
rect 3208 9791 3212 9795
rect 3213 9791 3217 9795
rect 3208 9786 3212 9790
rect 3213 9786 3217 9790
rect 3208 9781 3212 9785
rect 3213 9781 3217 9785
rect 3208 9776 3212 9780
rect 3213 9776 3217 9780
rect 3208 9771 3212 9775
rect 3213 9771 3217 9775
rect 3208 9766 3212 9770
rect 3213 9766 3217 9770
rect 3092 9760 3096 9764
rect 3097 9760 3101 9764
rect 3102 9760 3106 9764
rect 3107 9760 3111 9764
rect 3112 9760 3116 9764
rect 3117 9760 3121 9764
rect 3122 9760 3126 9764
rect 3127 9760 3131 9764
rect 3132 9760 3136 9764
rect 3137 9760 3141 9764
rect 3142 9760 3146 9764
rect 3147 9760 3151 9764
rect 3152 9760 3156 9764
rect 3173 9762 3177 9766
rect 3178 9762 3182 9766
rect 3183 9762 3187 9766
rect 3188 9762 3192 9766
rect 3173 9752 3177 9756
rect 3178 9752 3182 9756
rect 3183 9752 3187 9756
rect 3188 9752 3192 9756
rect 3173 9742 3177 9746
rect 3178 9742 3182 9746
rect 3183 9742 3187 9746
rect 3188 9742 3192 9746
rect 3173 9732 3177 9736
rect 3178 9732 3182 9736
rect 3183 9732 3187 9736
rect 3188 9732 3192 9736
rect 3208 9761 3212 9765
rect 3213 9761 3217 9765
rect 3208 9756 3212 9760
rect 3213 9756 3217 9760
rect 3208 9751 3212 9755
rect 3213 9751 3217 9755
rect 3208 9746 3212 9750
rect 3213 9746 3217 9750
rect 3208 9741 3212 9745
rect 3213 9741 3217 9745
rect 3208 9736 3212 9740
rect 3213 9736 3217 9740
rect 2932 9708 2936 9712
rect 2937 9708 2941 9712
rect 2942 9708 2946 9712
rect 2947 9708 2951 9712
rect 2952 9708 2956 9712
rect 2957 9708 2961 9712
rect 2962 9708 2966 9712
rect 2967 9708 2971 9712
rect 2972 9708 2976 9712
rect 2977 9708 2981 9712
rect 2982 9708 2986 9712
rect 2987 9708 2991 9712
rect 2992 9708 2996 9712
rect 2932 9703 2936 9707
rect 2937 9703 2941 9707
rect 2942 9703 2946 9707
rect 2947 9703 2951 9707
rect 2952 9703 2956 9707
rect 2957 9703 2961 9707
rect 2962 9703 2966 9707
rect 2967 9703 2971 9707
rect 2972 9703 2976 9707
rect 2977 9703 2981 9707
rect 2982 9703 2986 9707
rect 2987 9703 2991 9707
rect 2992 9703 2996 9707
rect 3114 9708 3118 9712
rect 3119 9708 3123 9712
rect 3124 9708 3128 9712
rect 3129 9708 3133 9712
rect 3134 9708 3138 9712
rect 3139 9708 3143 9712
rect 3144 9708 3148 9712
rect 3149 9708 3153 9712
rect 3154 9708 3158 9712
rect 3159 9708 3163 9712
rect 3164 9708 3168 9712
rect 3114 9703 3118 9707
rect 3119 9703 3123 9707
rect 3124 9703 3128 9707
rect 3129 9703 3133 9707
rect 3134 9703 3138 9707
rect 3139 9703 3143 9707
rect 3144 9703 3148 9707
rect 3149 9703 3153 9707
rect 3154 9703 3158 9707
rect 3159 9703 3163 9707
rect 3164 9703 3168 9707
rect 3173 9716 3177 9720
rect 3178 9716 3182 9720
rect 3183 9716 3187 9720
rect 3188 9716 3192 9720
rect 3173 9706 3177 9710
rect 3178 9706 3182 9710
rect 3183 9706 3187 9710
rect 3188 9706 3192 9710
rect 3401 9765 3405 9769
rect 3406 9765 3410 9769
rect 3411 9765 3415 9769
rect 3416 9765 3420 9769
rect 3421 9765 3425 9769
rect 3426 9765 3430 9769
rect 3431 9765 3435 9769
rect 3436 9765 3440 9769
rect 3441 9765 3445 9769
rect 3446 9765 3450 9769
rect 3451 9765 3455 9769
rect 3456 9765 3460 9769
rect 3461 9765 3465 9769
rect 3517 9796 3521 9800
rect 3522 9796 3526 9800
rect 3517 9791 3521 9795
rect 3522 9791 3526 9795
rect 3517 9786 3521 9790
rect 3522 9786 3526 9790
rect 3517 9781 3521 9785
rect 3522 9781 3526 9785
rect 3517 9776 3521 9780
rect 3522 9776 3526 9780
rect 3517 9771 3521 9775
rect 3522 9771 3526 9775
rect 3517 9766 3521 9770
rect 3522 9766 3526 9770
rect 3401 9760 3405 9764
rect 3406 9760 3410 9764
rect 3411 9760 3415 9764
rect 3416 9760 3420 9764
rect 3421 9760 3425 9764
rect 3426 9760 3430 9764
rect 3431 9760 3435 9764
rect 3436 9760 3440 9764
rect 3441 9760 3445 9764
rect 3446 9760 3450 9764
rect 3451 9760 3455 9764
rect 3456 9760 3460 9764
rect 3461 9760 3465 9764
rect 3482 9762 3486 9766
rect 3487 9762 3491 9766
rect 3492 9762 3496 9766
rect 3497 9762 3501 9766
rect 3482 9752 3486 9756
rect 3487 9752 3491 9756
rect 3492 9752 3496 9756
rect 3497 9752 3501 9756
rect 3482 9742 3486 9746
rect 3487 9742 3491 9746
rect 3492 9742 3496 9746
rect 3497 9742 3501 9746
rect 3482 9732 3486 9736
rect 3487 9732 3491 9736
rect 3492 9732 3496 9736
rect 3497 9732 3501 9736
rect 3517 9761 3521 9765
rect 3522 9761 3526 9765
rect 3517 9756 3521 9760
rect 3522 9756 3526 9760
rect 3517 9751 3521 9755
rect 3522 9751 3526 9755
rect 3517 9746 3521 9750
rect 3522 9746 3526 9750
rect 3517 9741 3521 9745
rect 3522 9741 3526 9745
rect 3517 9736 3521 9740
rect 3522 9736 3526 9740
rect 3241 9708 3245 9712
rect 3246 9708 3250 9712
rect 3251 9708 3255 9712
rect 3256 9708 3260 9712
rect 3261 9708 3265 9712
rect 3266 9708 3270 9712
rect 3271 9708 3275 9712
rect 3276 9708 3280 9712
rect 3281 9708 3285 9712
rect 3286 9708 3290 9712
rect 3291 9708 3295 9712
rect 3296 9708 3300 9712
rect 3301 9708 3305 9712
rect 3241 9703 3245 9707
rect 3246 9703 3250 9707
rect 3251 9703 3255 9707
rect 3256 9703 3260 9707
rect 3261 9703 3265 9707
rect 3266 9703 3270 9707
rect 3271 9703 3275 9707
rect 3276 9703 3280 9707
rect 3281 9703 3285 9707
rect 3286 9703 3290 9707
rect 3291 9703 3295 9707
rect 3296 9703 3300 9707
rect 3301 9703 3305 9707
rect 3343 9711 3347 9715
rect 3348 9711 3352 9715
rect 3343 9706 3347 9710
rect 3348 9706 3352 9710
rect 3343 9701 3347 9705
rect 3348 9701 3352 9705
rect 3423 9708 3427 9712
rect 3428 9708 3432 9712
rect 3433 9708 3437 9712
rect 3438 9708 3442 9712
rect 3443 9708 3447 9712
rect 3448 9708 3452 9712
rect 3453 9708 3457 9712
rect 3458 9708 3462 9712
rect 3463 9708 3467 9712
rect 3468 9708 3472 9712
rect 3473 9708 3477 9712
rect 3423 9703 3427 9707
rect 3428 9703 3432 9707
rect 3433 9703 3437 9707
rect 3438 9703 3442 9707
rect 3443 9703 3447 9707
rect 3448 9703 3452 9707
rect 3453 9703 3457 9707
rect 3458 9703 3462 9707
rect 3463 9703 3467 9707
rect 3468 9703 3472 9707
rect 3473 9703 3477 9707
rect 3482 9716 3486 9720
rect 3487 9716 3491 9720
rect 3492 9716 3496 9720
rect 3497 9716 3501 9720
rect 3482 9706 3486 9710
rect 3487 9706 3491 9710
rect 3492 9706 3496 9710
rect 3497 9706 3501 9710
rect 2246 9696 2250 9700
rect 2251 9696 2255 9700
rect 2256 9696 2260 9700
rect 2261 9696 2265 9700
rect 2246 9686 2250 9690
rect 2251 9686 2255 9690
rect 2256 9686 2260 9690
rect 2261 9686 2265 9690
rect 2555 9696 2559 9700
rect 2560 9696 2564 9700
rect 2565 9696 2569 9700
rect 2570 9696 2574 9700
rect 2555 9686 2559 9690
rect 2560 9686 2564 9690
rect 2565 9686 2569 9690
rect 2570 9686 2574 9690
rect 2864 9696 2868 9700
rect 2869 9696 2873 9700
rect 2874 9696 2878 9700
rect 2879 9696 2883 9700
rect 2864 9686 2868 9690
rect 2869 9686 2873 9690
rect 2874 9686 2878 9690
rect 2879 9686 2883 9690
rect 3173 9696 3177 9700
rect 3178 9696 3182 9700
rect 3183 9696 3187 9700
rect 3188 9696 3192 9700
rect 3173 9686 3177 9690
rect 3178 9686 3182 9690
rect 3183 9686 3187 9690
rect 3188 9686 3192 9690
rect 3343 9696 3347 9700
rect 3348 9696 3352 9700
rect 3343 9691 3347 9695
rect 3348 9691 3352 9695
rect 3343 9686 3347 9690
rect 3348 9686 3352 9690
rect 3652 9791 3656 9795
rect 3657 9791 3661 9795
rect 3652 9786 3656 9790
rect 3657 9786 3661 9790
rect 3652 9781 3656 9785
rect 3657 9781 3661 9785
rect 3652 9776 3656 9780
rect 3657 9776 3661 9780
rect 3652 9771 3656 9775
rect 3657 9771 3661 9775
rect 3652 9766 3656 9770
rect 3657 9766 3661 9770
rect 3652 9761 3656 9765
rect 3657 9761 3661 9765
rect 3652 9756 3656 9760
rect 3657 9756 3661 9760
rect 3710 9765 3714 9769
rect 3715 9765 3719 9769
rect 3720 9765 3724 9769
rect 3725 9765 3729 9769
rect 3730 9765 3734 9769
rect 3735 9765 3739 9769
rect 3740 9765 3744 9769
rect 3745 9765 3749 9769
rect 3750 9765 3754 9769
rect 3755 9765 3759 9769
rect 3760 9765 3764 9769
rect 3765 9765 3769 9769
rect 3770 9765 3774 9769
rect 3826 9796 3830 9800
rect 3831 9796 3835 9800
rect 3826 9791 3830 9795
rect 3831 9791 3835 9795
rect 3826 9786 3830 9790
rect 3831 9786 3835 9790
rect 3826 9781 3830 9785
rect 3831 9781 3835 9785
rect 3826 9776 3830 9780
rect 3831 9776 3835 9780
rect 3826 9771 3830 9775
rect 3831 9771 3835 9775
rect 3826 9766 3830 9770
rect 3831 9766 3835 9770
rect 3710 9760 3714 9764
rect 3715 9760 3719 9764
rect 3720 9760 3724 9764
rect 3725 9760 3729 9764
rect 3730 9760 3734 9764
rect 3735 9760 3739 9764
rect 3740 9760 3744 9764
rect 3745 9760 3749 9764
rect 3750 9760 3754 9764
rect 3755 9760 3759 9764
rect 3760 9760 3764 9764
rect 3765 9760 3769 9764
rect 3770 9760 3774 9764
rect 3791 9762 3795 9766
rect 3796 9762 3800 9766
rect 3801 9762 3805 9766
rect 3806 9762 3810 9766
rect 3652 9751 3656 9755
rect 3657 9751 3661 9755
rect 3652 9746 3656 9750
rect 3657 9746 3661 9750
rect 3652 9741 3656 9745
rect 3657 9741 3661 9745
rect 3791 9752 3795 9756
rect 3796 9752 3800 9756
rect 3801 9752 3805 9756
rect 3806 9752 3810 9756
rect 3791 9742 3795 9746
rect 3796 9742 3800 9746
rect 3801 9742 3805 9746
rect 3806 9742 3810 9746
rect 3791 9732 3795 9736
rect 3796 9732 3800 9736
rect 3801 9732 3805 9736
rect 3806 9732 3810 9736
rect 3826 9761 3830 9765
rect 3831 9761 3835 9765
rect 3826 9756 3830 9760
rect 3831 9756 3835 9760
rect 3826 9751 3830 9755
rect 3831 9751 3835 9755
rect 3826 9746 3830 9750
rect 3831 9746 3835 9750
rect 3826 9741 3830 9745
rect 3831 9741 3835 9745
rect 3826 9736 3830 9740
rect 3831 9736 3835 9740
rect 3550 9708 3554 9712
rect 3555 9708 3559 9712
rect 3560 9708 3564 9712
rect 3565 9708 3569 9712
rect 3570 9708 3574 9712
rect 3575 9708 3579 9712
rect 3580 9708 3584 9712
rect 3585 9708 3589 9712
rect 3590 9708 3594 9712
rect 3595 9708 3599 9712
rect 3600 9708 3604 9712
rect 3605 9708 3609 9712
rect 3610 9708 3614 9712
rect 3550 9703 3554 9707
rect 3555 9703 3559 9707
rect 3560 9703 3564 9707
rect 3565 9703 3569 9707
rect 3570 9703 3574 9707
rect 3575 9703 3579 9707
rect 3580 9703 3584 9707
rect 3585 9703 3589 9707
rect 3590 9703 3594 9707
rect 3595 9703 3599 9707
rect 3600 9703 3604 9707
rect 3605 9703 3609 9707
rect 3610 9703 3614 9707
rect 3732 9708 3736 9712
rect 3737 9708 3741 9712
rect 3742 9708 3746 9712
rect 3747 9708 3751 9712
rect 3752 9708 3756 9712
rect 3757 9708 3761 9712
rect 3762 9708 3766 9712
rect 3767 9708 3771 9712
rect 3772 9708 3776 9712
rect 3777 9708 3781 9712
rect 3782 9708 3786 9712
rect 3732 9703 3736 9707
rect 3737 9703 3741 9707
rect 3742 9703 3746 9707
rect 3747 9703 3751 9707
rect 3752 9703 3756 9707
rect 3757 9703 3761 9707
rect 3762 9703 3766 9707
rect 3767 9703 3771 9707
rect 3772 9703 3776 9707
rect 3777 9703 3781 9707
rect 3782 9703 3786 9707
rect 3791 9716 3795 9720
rect 3796 9716 3800 9720
rect 3801 9716 3805 9720
rect 3806 9716 3810 9720
rect 3791 9706 3795 9710
rect 3796 9706 3800 9710
rect 3801 9706 3805 9710
rect 3806 9706 3810 9710
rect 4019 9765 4023 9769
rect 4024 9765 4028 9769
rect 4029 9765 4033 9769
rect 4034 9765 4038 9769
rect 4039 9765 4043 9769
rect 4044 9765 4048 9769
rect 4049 9765 4053 9769
rect 4054 9765 4058 9769
rect 4059 9765 4063 9769
rect 4064 9765 4068 9769
rect 4069 9765 4073 9769
rect 4074 9765 4078 9769
rect 4079 9765 4083 9769
rect 4019 9760 4023 9764
rect 4024 9760 4028 9764
rect 4029 9760 4033 9764
rect 4034 9760 4038 9764
rect 4039 9760 4043 9764
rect 4044 9760 4048 9764
rect 4049 9760 4053 9764
rect 4054 9760 4058 9764
rect 4059 9760 4063 9764
rect 4064 9760 4068 9764
rect 4069 9760 4073 9764
rect 4074 9760 4078 9764
rect 4079 9760 4083 9764
rect 4100 9762 4104 9766
rect 4105 9762 4109 9766
rect 4110 9762 4114 9766
rect 4115 9762 4119 9766
rect 4100 9752 4104 9756
rect 4105 9752 4109 9756
rect 4110 9752 4114 9756
rect 4115 9752 4119 9756
rect 4100 9742 4104 9746
rect 4105 9742 4109 9746
rect 4110 9742 4114 9746
rect 4115 9742 4119 9746
rect 4100 9732 4104 9736
rect 4105 9732 4109 9736
rect 4110 9732 4114 9736
rect 4115 9732 4119 9736
rect 4292 9762 4296 9766
rect 4297 9762 4301 9766
rect 4302 9762 4306 9766
rect 4307 9762 4311 9766
rect 4292 9752 4296 9756
rect 4297 9752 4301 9756
rect 4302 9752 4306 9756
rect 4307 9752 4311 9756
rect 4292 9742 4296 9746
rect 4297 9742 4301 9746
rect 4302 9742 4306 9746
rect 4307 9742 4311 9746
rect 4292 9732 4296 9736
rect 4297 9732 4301 9736
rect 4302 9732 4306 9736
rect 4307 9732 4311 9736
rect 4318 9762 4322 9766
rect 4323 9762 4327 9766
rect 4328 9762 4332 9766
rect 4333 9762 4337 9766
rect 4318 9752 4322 9756
rect 4323 9752 4327 9756
rect 4328 9752 4332 9756
rect 4333 9752 4337 9756
rect 4318 9742 4322 9746
rect 4323 9742 4327 9746
rect 4328 9742 4332 9746
rect 4333 9742 4337 9746
rect 4318 9732 4322 9736
rect 4323 9732 4327 9736
rect 4328 9732 4332 9736
rect 4333 9732 4337 9736
rect 4344 9762 4348 9766
rect 4349 9762 4353 9766
rect 4354 9762 4358 9766
rect 4359 9762 4363 9766
rect 4344 9752 4348 9756
rect 4349 9752 4353 9756
rect 4354 9752 4358 9756
rect 4359 9752 4363 9756
rect 4344 9742 4348 9746
rect 4349 9742 4353 9746
rect 4354 9742 4358 9746
rect 4359 9742 4363 9746
rect 4344 9732 4348 9736
rect 4349 9732 4353 9736
rect 4354 9732 4358 9736
rect 4359 9732 4363 9736
rect 4370 9762 4374 9766
rect 4375 9762 4379 9766
rect 4380 9762 4384 9766
rect 4385 9762 4389 9766
rect 4370 9752 4374 9756
rect 4375 9752 4379 9756
rect 4380 9752 4384 9756
rect 4385 9752 4389 9756
rect 4370 9742 4374 9746
rect 4375 9742 4379 9746
rect 4380 9742 4384 9746
rect 4385 9742 4389 9746
rect 4370 9732 4374 9736
rect 4375 9732 4379 9736
rect 4380 9732 4384 9736
rect 4385 9732 4389 9736
rect 4396 9762 4400 9766
rect 4401 9762 4405 9766
rect 4406 9762 4410 9766
rect 4411 9762 4415 9766
rect 4396 9752 4400 9756
rect 4401 9752 4405 9756
rect 4406 9752 4410 9756
rect 4411 9752 4415 9756
rect 4396 9742 4400 9746
rect 4401 9742 4405 9746
rect 4406 9742 4410 9746
rect 4411 9742 4415 9746
rect 4396 9732 4400 9736
rect 4401 9732 4405 9736
rect 4406 9732 4410 9736
rect 4411 9732 4415 9736
rect 3859 9708 3863 9712
rect 3864 9708 3868 9712
rect 3869 9708 3873 9712
rect 3874 9708 3878 9712
rect 3879 9708 3883 9712
rect 3884 9708 3888 9712
rect 3889 9708 3893 9712
rect 3894 9708 3898 9712
rect 3899 9708 3903 9712
rect 3904 9708 3908 9712
rect 3909 9708 3913 9712
rect 3914 9708 3918 9712
rect 3919 9708 3923 9712
rect 3859 9703 3863 9707
rect 3864 9703 3868 9707
rect 3869 9703 3873 9707
rect 3874 9703 3878 9707
rect 3879 9703 3883 9707
rect 3884 9703 3888 9707
rect 3889 9703 3893 9707
rect 3894 9703 3898 9707
rect 3899 9703 3903 9707
rect 3904 9703 3908 9707
rect 3909 9703 3913 9707
rect 3914 9703 3918 9707
rect 3919 9703 3923 9707
rect 4041 9708 4045 9712
rect 4046 9708 4050 9712
rect 4051 9708 4055 9712
rect 4056 9708 4060 9712
rect 4061 9708 4065 9712
rect 4066 9708 4070 9712
rect 4071 9708 4075 9712
rect 4076 9708 4080 9712
rect 4081 9708 4085 9712
rect 4086 9708 4090 9712
rect 4091 9708 4095 9712
rect 4041 9703 4045 9707
rect 4046 9703 4050 9707
rect 4051 9703 4055 9707
rect 4056 9703 4060 9707
rect 4061 9703 4065 9707
rect 4066 9703 4070 9707
rect 4071 9703 4075 9707
rect 4076 9703 4080 9707
rect 4081 9703 4085 9707
rect 4086 9703 4090 9707
rect 4091 9703 4095 9707
rect 4100 9716 4104 9720
rect 4105 9716 4109 9720
rect 4110 9716 4114 9720
rect 4115 9716 4119 9720
rect 4100 9706 4104 9710
rect 4105 9706 4109 9710
rect 4110 9706 4114 9710
rect 4115 9706 4119 9710
rect 3482 9696 3486 9700
rect 3487 9696 3491 9700
rect 3492 9696 3496 9700
rect 3497 9696 3501 9700
rect 3482 9686 3486 9690
rect 3487 9686 3491 9690
rect 3492 9686 3496 9690
rect 3497 9686 3501 9690
rect 3791 9696 3795 9700
rect 3796 9696 3800 9700
rect 3801 9696 3805 9700
rect 3806 9696 3810 9700
rect 3791 9686 3795 9690
rect 3796 9686 3800 9690
rect 3801 9686 3805 9690
rect 3806 9686 3810 9690
rect 4100 9696 4104 9700
rect 4105 9696 4109 9700
rect 4110 9696 4114 9700
rect 4115 9696 4119 9700
rect 4100 9686 4104 9690
rect 4105 9686 4109 9690
rect 4110 9686 4114 9690
rect 4115 9686 4119 9690
rect 4292 9716 4296 9720
rect 4297 9716 4301 9720
rect 4302 9716 4306 9720
rect 4307 9716 4311 9720
rect 4292 9706 4296 9710
rect 4297 9706 4301 9710
rect 4302 9706 4306 9710
rect 4307 9706 4311 9710
rect 4292 9696 4296 9700
rect 4297 9696 4301 9700
rect 4302 9696 4306 9700
rect 4307 9696 4311 9700
rect 4292 9686 4296 9690
rect 4297 9686 4301 9690
rect 4302 9686 4306 9690
rect 4307 9686 4311 9690
rect 4318 9716 4322 9720
rect 4323 9716 4327 9720
rect 4328 9716 4332 9720
rect 4333 9716 4337 9720
rect 4318 9706 4322 9710
rect 4323 9706 4327 9710
rect 4328 9706 4332 9710
rect 4333 9706 4337 9710
rect 4318 9696 4322 9700
rect 4323 9696 4327 9700
rect 4328 9696 4332 9700
rect 4333 9696 4337 9700
rect 4318 9686 4322 9690
rect 4323 9686 4327 9690
rect 4328 9686 4332 9690
rect 4333 9686 4337 9690
rect 4344 9716 4348 9720
rect 4349 9716 4353 9720
rect 4354 9716 4358 9720
rect 4359 9716 4363 9720
rect 4344 9706 4348 9710
rect 4349 9706 4353 9710
rect 4354 9706 4358 9710
rect 4359 9706 4363 9710
rect 4344 9696 4348 9700
rect 4349 9696 4353 9700
rect 4354 9696 4358 9700
rect 4359 9696 4363 9700
rect 4344 9686 4348 9690
rect 4349 9686 4353 9690
rect 4354 9686 4358 9690
rect 4359 9686 4363 9690
rect 4370 9716 4374 9720
rect 4375 9716 4379 9720
rect 4380 9716 4384 9720
rect 4385 9716 4389 9720
rect 4370 9706 4374 9710
rect 4375 9706 4379 9710
rect 4380 9706 4384 9710
rect 4385 9706 4389 9710
rect 4370 9696 4374 9700
rect 4375 9696 4379 9700
rect 4380 9696 4384 9700
rect 4385 9696 4389 9700
rect 4370 9686 4374 9690
rect 4375 9686 4379 9690
rect 4380 9686 4384 9690
rect 4385 9686 4389 9690
rect 4396 9716 4400 9720
rect 4401 9716 4405 9720
rect 4406 9716 4410 9720
rect 4411 9716 4415 9720
rect 4396 9706 4400 9710
rect 4401 9706 4405 9710
rect 4406 9706 4410 9710
rect 4411 9706 4415 9710
rect 4396 9696 4400 9700
rect 4401 9696 4405 9700
rect 4406 9696 4410 9700
rect 4411 9696 4415 9700
rect 4396 9686 4400 9690
rect 4401 9686 4405 9690
rect 4406 9686 4410 9690
rect 4411 9686 4415 9690
rect 3343 9681 3347 9685
rect 3348 9681 3352 9685
rect 3343 9676 3347 9680
rect 3348 9676 3352 9680
rect 3343 9671 3347 9675
rect 3348 9671 3352 9675
rect 3343 9666 3347 9670
rect 3348 9666 3352 9670
rect 3343 9661 3347 9665
rect 3348 9661 3352 9665
rect 613 9618 617 9622
rect 623 9618 627 9622
rect 633 9618 637 9622
rect 643 9618 647 9622
rect 613 9613 617 9617
rect 623 9613 627 9617
rect 633 9613 637 9617
rect 643 9613 647 9617
rect 613 9608 617 9612
rect 623 9608 627 9612
rect 633 9608 637 9612
rect 643 9608 647 9612
rect 613 9603 617 9607
rect 623 9603 627 9607
rect 633 9603 637 9607
rect 643 9603 647 9607
rect 659 9618 663 9622
rect 669 9618 673 9622
rect 679 9618 683 9622
rect 689 9618 693 9622
rect 659 9613 663 9617
rect 669 9613 673 9617
rect 679 9613 683 9617
rect 689 9613 693 9617
rect 659 9608 663 9612
rect 669 9608 673 9612
rect 679 9608 683 9612
rect 689 9608 693 9612
rect 659 9603 663 9607
rect 669 9603 673 9607
rect 679 9603 683 9607
rect 689 9603 693 9607
rect 613 9592 617 9596
rect 623 9592 627 9596
rect 633 9592 637 9596
rect 643 9592 647 9596
rect 613 9587 617 9591
rect 623 9587 627 9591
rect 633 9587 637 9591
rect 643 9587 647 9591
rect 613 9582 617 9586
rect 623 9582 627 9586
rect 633 9582 637 9586
rect 643 9582 647 9586
rect 613 9577 617 9581
rect 623 9577 627 9581
rect 633 9577 637 9581
rect 643 9577 647 9581
rect 659 9592 663 9596
rect 669 9592 673 9596
rect 679 9592 683 9596
rect 689 9592 693 9596
rect 659 9587 663 9591
rect 669 9587 673 9591
rect 679 9587 683 9591
rect 689 9587 693 9591
rect 659 9582 663 9586
rect 669 9582 673 9586
rect 679 9582 683 9586
rect 689 9582 693 9586
rect 659 9577 663 9581
rect 669 9577 673 9581
rect 679 9577 683 9581
rect 689 9577 693 9581
rect 2258 9619 2262 9623
rect 613 9566 617 9570
rect 623 9566 627 9570
rect 633 9566 637 9570
rect 643 9566 647 9570
rect 613 9561 617 9565
rect 623 9561 627 9565
rect 633 9561 637 9565
rect 643 9561 647 9565
rect 613 9556 617 9560
rect 623 9556 627 9560
rect 633 9556 637 9560
rect 643 9556 647 9560
rect 613 9551 617 9555
rect 623 9551 627 9555
rect 633 9551 637 9555
rect 643 9551 647 9555
rect 659 9566 663 9570
rect 669 9566 673 9570
rect 679 9566 683 9570
rect 689 9566 693 9570
rect 659 9561 663 9565
rect 669 9561 673 9565
rect 679 9561 683 9565
rect 689 9561 693 9565
rect 659 9556 663 9560
rect 669 9556 673 9560
rect 679 9556 683 9560
rect 689 9556 693 9560
rect 659 9551 663 9555
rect 669 9551 673 9555
rect 679 9551 683 9555
rect 689 9551 693 9555
rect 613 9540 617 9544
rect 623 9540 627 9544
rect 633 9540 637 9544
rect 643 9540 647 9544
rect 613 9535 617 9539
rect 623 9535 627 9539
rect 633 9535 637 9539
rect 643 9535 647 9539
rect 613 9530 617 9534
rect 623 9530 627 9534
rect 633 9530 637 9534
rect 643 9530 647 9534
rect 613 9525 617 9529
rect 623 9525 627 9529
rect 633 9525 637 9529
rect 643 9525 647 9529
rect 659 9540 663 9544
rect 669 9540 673 9544
rect 679 9540 683 9544
rect 689 9540 693 9544
rect 659 9535 663 9539
rect 669 9535 673 9539
rect 679 9535 683 9539
rect 689 9535 693 9539
rect 659 9530 663 9534
rect 669 9530 673 9534
rect 679 9530 683 9534
rect 689 9530 693 9534
rect 659 9525 663 9529
rect 669 9525 673 9529
rect 679 9525 683 9529
rect 689 9525 693 9529
rect 613 9514 617 9518
rect 623 9514 627 9518
rect 633 9514 637 9518
rect 643 9514 647 9518
rect 613 9509 617 9513
rect 623 9509 627 9513
rect 633 9509 637 9513
rect 643 9509 647 9513
rect 613 9504 617 9508
rect 623 9504 627 9508
rect 633 9504 637 9508
rect 643 9504 647 9508
rect 613 9499 617 9503
rect 623 9499 627 9503
rect 633 9499 637 9503
rect 643 9499 647 9503
rect 659 9514 663 9518
rect 669 9514 673 9518
rect 679 9514 683 9518
rect 689 9514 693 9518
rect 659 9509 663 9513
rect 669 9509 673 9513
rect 679 9509 683 9513
rect 689 9509 693 9513
rect 659 9504 663 9508
rect 669 9504 673 9508
rect 679 9504 683 9508
rect 689 9504 693 9508
rect 659 9499 663 9503
rect 669 9499 673 9503
rect 679 9499 683 9503
rect 689 9499 693 9503
rect 613 9321 617 9325
rect 623 9321 627 9325
rect 633 9321 637 9325
rect 643 9321 647 9325
rect 613 9316 617 9320
rect 623 9316 627 9320
rect 633 9316 637 9320
rect 643 9316 647 9320
rect 613 9311 617 9315
rect 623 9311 627 9315
rect 633 9311 637 9315
rect 643 9311 647 9315
rect 613 9306 617 9310
rect 623 9306 627 9310
rect 633 9306 637 9310
rect 643 9306 647 9310
rect 659 9321 663 9325
rect 669 9321 673 9325
rect 679 9321 683 9325
rect 689 9321 693 9325
rect 659 9316 663 9320
rect 669 9316 673 9320
rect 679 9316 683 9320
rect 689 9316 693 9320
rect 659 9311 663 9315
rect 669 9311 673 9315
rect 679 9311 683 9315
rect 689 9311 693 9315
rect 659 9306 663 9310
rect 669 9306 673 9310
rect 679 9306 683 9310
rect 689 9306 693 9310
rect 613 9012 617 9016
rect 623 9012 627 9016
rect 633 9012 637 9016
rect 643 9012 647 9016
rect 613 9007 617 9011
rect 623 9007 627 9011
rect 633 9007 637 9011
rect 643 9007 647 9011
rect 613 9002 617 9006
rect 623 9002 627 9006
rect 633 9002 637 9006
rect 643 9002 647 9006
rect 613 8997 617 9001
rect 623 8997 627 9001
rect 633 8997 637 9001
rect 643 8997 647 9001
rect 659 9012 663 9016
rect 669 9012 673 9016
rect 679 9012 683 9016
rect 689 9012 693 9016
rect 659 9007 663 9011
rect 669 9007 673 9011
rect 679 9007 683 9011
rect 689 9007 693 9011
rect 659 9002 663 9006
rect 669 9002 673 9006
rect 679 9002 683 9006
rect 689 9002 693 9006
rect 659 8997 663 9001
rect 669 8997 673 9001
rect 679 8997 683 9001
rect 689 8997 693 9001
rect 613 8703 617 8707
rect 623 8703 627 8707
rect 633 8703 637 8707
rect 643 8703 647 8707
rect 613 8698 617 8702
rect 623 8698 627 8702
rect 633 8698 637 8702
rect 643 8698 647 8702
rect 613 8693 617 8697
rect 623 8693 627 8697
rect 633 8693 637 8697
rect 643 8693 647 8697
rect 613 8688 617 8692
rect 623 8688 627 8692
rect 633 8688 637 8692
rect 643 8688 647 8692
rect 659 8703 663 8707
rect 669 8703 673 8707
rect 679 8703 683 8707
rect 689 8703 693 8707
rect 659 8698 663 8702
rect 669 8698 673 8702
rect 679 8698 683 8702
rect 689 8698 693 8702
rect 659 8693 663 8697
rect 669 8693 673 8697
rect 679 8693 683 8697
rect 689 8693 693 8697
rect 659 8688 663 8692
rect 669 8688 673 8692
rect 679 8688 683 8692
rect 689 8688 693 8692
rect 2624 9277 2628 9281
rect 613 8394 617 8398
rect 623 8394 627 8398
rect 633 8394 637 8398
rect 643 8394 647 8398
rect 613 8389 617 8393
rect 623 8389 627 8393
rect 633 8389 637 8393
rect 643 8389 647 8393
rect 613 8384 617 8388
rect 623 8384 627 8388
rect 633 8384 637 8388
rect 643 8384 647 8388
rect 613 8379 617 8383
rect 623 8379 627 8383
rect 633 8379 637 8383
rect 643 8379 647 8383
rect 659 8394 663 8398
rect 669 8394 673 8398
rect 679 8394 683 8398
rect 689 8394 693 8398
rect 659 8389 663 8393
rect 669 8389 673 8393
rect 679 8389 683 8393
rect 689 8389 693 8393
rect 659 8384 663 8388
rect 669 8384 673 8388
rect 679 8384 683 8388
rect 689 8384 693 8388
rect 659 8379 663 8383
rect 669 8379 673 8383
rect 679 8379 683 8383
rect 689 8379 693 8383
rect 2623 9174 2627 9178
rect 613 8085 617 8089
rect 623 8085 627 8089
rect 633 8085 637 8089
rect 643 8085 647 8089
rect 613 8080 617 8084
rect 623 8080 627 8084
rect 633 8080 637 8084
rect 643 8080 647 8084
rect 613 8075 617 8079
rect 623 8075 627 8079
rect 633 8075 637 8079
rect 643 8075 647 8079
rect 613 8070 617 8074
rect 623 8070 627 8074
rect 633 8070 637 8074
rect 643 8070 647 8074
rect 659 8085 663 8089
rect 669 8085 673 8089
rect 679 8085 683 8089
rect 689 8085 693 8089
rect 659 8080 663 8084
rect 669 8080 673 8084
rect 679 8080 683 8084
rect 689 8080 693 8084
rect 659 8075 663 8079
rect 669 8075 673 8079
rect 679 8075 683 8079
rect 689 8075 693 8079
rect 659 8070 663 8074
rect 669 8070 673 8074
rect 679 8070 683 8074
rect 689 8070 693 8074
rect 2367 7792 2371 7796
rect 613 7776 617 7780
rect 623 7776 627 7780
rect 633 7776 637 7780
rect 643 7776 647 7780
rect 613 7771 617 7775
rect 623 7771 627 7775
rect 633 7771 637 7775
rect 643 7771 647 7775
rect 613 7766 617 7770
rect 623 7766 627 7770
rect 633 7766 637 7770
rect 643 7766 647 7770
rect 613 7761 617 7765
rect 623 7761 627 7765
rect 633 7761 637 7765
rect 643 7761 647 7765
rect 659 7776 663 7780
rect 669 7776 673 7780
rect 679 7776 683 7780
rect 689 7776 693 7780
rect 659 7771 663 7775
rect 669 7771 673 7775
rect 679 7771 683 7775
rect 689 7771 693 7775
rect 659 7766 663 7770
rect 669 7766 673 7770
rect 679 7766 683 7770
rect 689 7766 693 7770
rect 659 7761 663 7765
rect 669 7761 673 7765
rect 679 7761 683 7765
rect 689 7761 693 7765
rect 2756 8407 2760 8411
rect 2624 8295 2628 8299
rect 613 7467 617 7471
rect 623 7467 627 7471
rect 633 7467 637 7471
rect 643 7467 647 7471
rect 613 7462 617 7466
rect 623 7462 627 7466
rect 633 7462 637 7466
rect 643 7462 647 7466
rect 613 7457 617 7461
rect 623 7457 627 7461
rect 633 7457 637 7461
rect 643 7457 647 7461
rect 613 7452 617 7456
rect 623 7452 627 7456
rect 633 7452 637 7456
rect 643 7452 647 7456
rect 659 7467 663 7471
rect 669 7467 673 7471
rect 679 7467 683 7471
rect 689 7467 693 7471
rect 659 7462 663 7466
rect 669 7462 673 7466
rect 679 7462 683 7466
rect 689 7462 693 7466
rect 659 7457 663 7461
rect 669 7457 673 7461
rect 679 7457 683 7461
rect 689 7457 693 7461
rect 659 7452 663 7456
rect 669 7452 673 7456
rect 679 7452 683 7456
rect 689 7452 693 7456
rect 2623 8192 2627 8196
rect 2756 7425 2760 7429
rect 4479 9573 4483 9577
rect 4489 9573 4493 9577
rect 4499 9573 4503 9577
rect 4509 9573 4513 9577
rect 4479 9568 4483 9572
rect 4489 9568 4493 9572
rect 4499 9568 4503 9572
rect 4509 9568 4513 9572
rect 4479 9563 4483 9567
rect 4489 9563 4493 9567
rect 4499 9563 4503 9567
rect 4509 9563 4513 9567
rect 4479 9558 4483 9562
rect 4489 9558 4493 9562
rect 4499 9558 4503 9562
rect 4509 9558 4513 9562
rect 4525 9573 4529 9577
rect 4535 9573 4539 9577
rect 4545 9573 4549 9577
rect 4555 9573 4559 9577
rect 4525 9568 4529 9572
rect 4535 9568 4539 9572
rect 4545 9568 4549 9572
rect 4555 9568 4559 9572
rect 4525 9563 4529 9567
rect 4535 9563 4539 9567
rect 4545 9563 4549 9567
rect 4555 9563 4559 9567
rect 4525 9558 4529 9562
rect 4535 9558 4539 9562
rect 4545 9558 4549 9562
rect 4555 9558 4559 9562
rect 4479 9544 4483 9548
rect 4489 9544 4493 9548
rect 4499 9544 4503 9548
rect 4509 9544 4513 9548
rect 4479 9539 4483 9543
rect 4489 9539 4493 9543
rect 4499 9539 4503 9543
rect 4509 9539 4513 9543
rect 4479 9534 4483 9538
rect 4489 9534 4493 9538
rect 4499 9534 4503 9538
rect 4509 9534 4513 9538
rect 4479 9529 4483 9533
rect 4489 9529 4493 9533
rect 4499 9529 4503 9533
rect 4509 9529 4513 9533
rect 4525 9544 4529 9548
rect 4535 9544 4539 9548
rect 4545 9544 4549 9548
rect 4555 9544 4559 9548
rect 4525 9539 4529 9543
rect 4535 9539 4539 9543
rect 4545 9539 4549 9543
rect 4555 9539 4559 9543
rect 4525 9534 4529 9538
rect 4535 9534 4539 9538
rect 4545 9534 4549 9538
rect 4555 9534 4559 9538
rect 4525 9529 4529 9533
rect 4535 9529 4539 9533
rect 4545 9529 4549 9533
rect 4555 9529 4559 9533
rect 4479 9515 4483 9519
rect 4489 9515 4493 9519
rect 4499 9515 4503 9519
rect 4509 9515 4513 9519
rect 4479 9510 4483 9514
rect 4489 9510 4493 9514
rect 4499 9510 4503 9514
rect 4509 9510 4513 9514
rect 4479 9505 4483 9509
rect 4489 9505 4493 9509
rect 4499 9505 4503 9509
rect 4509 9505 4513 9509
rect 4479 9500 4483 9504
rect 4489 9500 4493 9504
rect 4499 9500 4503 9504
rect 4509 9500 4513 9504
rect 4525 9515 4529 9519
rect 4535 9515 4539 9519
rect 4545 9515 4549 9519
rect 4555 9515 4559 9519
rect 4525 9510 4529 9514
rect 4535 9510 4539 9514
rect 4545 9510 4549 9514
rect 4555 9510 4559 9514
rect 4525 9505 4529 9509
rect 4535 9505 4539 9509
rect 4545 9505 4549 9509
rect 4555 9505 4559 9509
rect 4525 9500 4529 9504
rect 4535 9500 4539 9504
rect 4545 9500 4549 9504
rect 4555 9500 4559 9504
rect 2847 9313 2851 9317
rect 2887 9230 2892 9235
rect 2898 9226 2903 9231
rect 2921 9235 2926 9240
rect 2945 9230 2950 9235
rect 2960 9234 2965 9240
rect 2990 9230 2995 9235
rect 3019 9229 3024 9234
rect 2974 9224 2979 9229
rect 3003 9224 3007 9229
rect 3045 9223 3050 9228
rect 2851 9170 2856 9175
rect 2887 9163 2892 9168
rect 2898 9167 2903 9172
rect 2921 9158 2926 9163
rect 2945 9163 2950 9168
rect 2974 9169 2979 9174
rect 3003 9169 3007 9174
rect 2960 9158 2965 9164
rect 2990 9163 2995 9168
rect 3019 9164 3024 9169
rect 3045 9164 3050 9169
rect 2850 9101 2855 9106
rect 2887 9098 2892 9103
rect 2898 9094 2903 9099
rect 2921 9103 2926 9108
rect 2945 9098 2950 9103
rect 3101 9229 3106 9234
rect 2960 9102 2965 9108
rect 2990 9098 2995 9103
rect 3019 9097 3024 9102
rect 2974 9092 2979 9097
rect 3003 9092 3007 9097
rect 3045 9091 3050 9096
rect 2851 9038 2856 9043
rect 2887 9031 2892 9036
rect 2898 9035 2903 9040
rect 2921 9026 2926 9031
rect 2945 9031 2950 9036
rect 2974 9037 2979 9042
rect 3003 9037 3007 9042
rect 2960 9026 2965 9032
rect 2990 9031 2995 9036
rect 3019 9032 3024 9037
rect 3044 9033 3049 9038
rect 2850 8969 2855 8974
rect 2887 8966 2892 8971
rect 2898 8962 2903 8967
rect 2921 8971 2926 8976
rect 2945 8966 2950 8971
rect 2960 8970 2965 8976
rect 2990 8966 2995 8971
rect 3019 8965 3024 8970
rect 2974 8960 2979 8965
rect 3003 8960 3007 8965
rect 3045 8959 3050 8964
rect 3101 9105 3106 9110
rect 3126 9223 3131 9228
rect 3125 9164 3130 9169
rect 3186 9229 3191 9234
rect 3150 9091 3155 9096
rect 3150 9033 3155 9038
rect 2851 8906 2856 8911
rect 2887 8899 2892 8904
rect 2898 8903 2903 8908
rect 2921 8894 2926 8899
rect 2945 8899 2950 8904
rect 2974 8905 2979 8910
rect 3003 8905 3007 8910
rect 2960 8894 2965 8900
rect 2990 8899 2995 8904
rect 3019 8900 3024 8905
rect 3045 8898 3050 8903
rect 2850 8837 2855 8842
rect 2887 8834 2892 8839
rect 2898 8830 2903 8835
rect 2921 8839 2926 8844
rect 2945 8834 2950 8839
rect 2960 8838 2965 8844
rect 2990 8834 2995 8839
rect 3019 8833 3024 8838
rect 2974 8828 2979 8833
rect 3003 8828 3007 8833
rect 3045 8827 3050 8832
rect 3101 8965 3106 8970
rect 3126 8959 3131 8964
rect 3125 8898 3130 8903
rect 3303 9262 3307 9266
rect 3208 9102 3213 9107
rect 3569 9277 3573 9281
rect 3568 9174 3572 9178
rect 3443 9135 3448 9140
rect 3560 9136 3565 9141
rect 3183 8974 3188 8979
rect 3217 8967 3222 8972
rect 3214 8894 3219 8899
rect 2851 8774 2856 8779
rect 2887 8767 2892 8772
rect 2898 8771 2903 8776
rect 2921 8762 2926 8767
rect 2945 8767 2950 8772
rect 2974 8773 2979 8778
rect 3003 8773 3007 8778
rect 2960 8762 2965 8768
rect 2990 8767 2995 8772
rect 3019 8768 3024 8773
rect 3044 8762 3049 8767
rect 3101 8841 3106 8846
rect 3089 8773 3094 8778
rect 3148 8767 3153 8772
rect 3159 8771 3164 8776
rect 3182 8762 3187 8767
rect 3206 8767 3211 8772
rect 3235 8773 3240 8778
rect 3264 8773 3268 8778
rect 3221 8762 3226 8768
rect 3251 8767 3256 8772
rect 3276 8773 3281 8778
rect 3443 8819 3448 8824
rect 3312 8774 3316 8778
rect 3150 8662 3154 8666
rect 3560 8818 3565 8823
rect 3275 8580 3279 8584
rect 2847 8331 2851 8335
rect 2887 8248 2892 8253
rect 2898 8244 2903 8249
rect 2921 8253 2926 8258
rect 2945 8248 2950 8253
rect 2960 8252 2965 8258
rect 2990 8248 2995 8253
rect 3019 8247 3024 8252
rect 2974 8242 2979 8247
rect 3003 8242 3007 8247
rect 3045 8241 3050 8246
rect 2851 8188 2856 8193
rect 2887 8181 2892 8186
rect 2898 8185 2903 8190
rect 2921 8176 2926 8181
rect 2945 8181 2950 8186
rect 2974 8187 2979 8192
rect 3003 8187 3007 8192
rect 2960 8176 2965 8182
rect 2990 8181 2995 8186
rect 3019 8182 3024 8187
rect 3045 8182 3050 8187
rect 2850 8119 2855 8124
rect 2887 8116 2892 8121
rect 2898 8112 2903 8117
rect 2921 8121 2926 8126
rect 2945 8116 2950 8121
rect 3101 8247 3106 8252
rect 2960 8120 2965 8126
rect 2990 8116 2995 8121
rect 3019 8115 3024 8120
rect 2974 8110 2979 8115
rect 3003 8110 3007 8115
rect 3045 8109 3050 8114
rect 2851 8056 2856 8061
rect 2887 8049 2892 8054
rect 2898 8053 2903 8058
rect 2921 8044 2926 8049
rect 2945 8049 2950 8054
rect 2974 8055 2979 8060
rect 3003 8055 3007 8060
rect 2960 8044 2965 8050
rect 2990 8049 2995 8054
rect 3019 8050 3024 8055
rect 3044 8051 3049 8056
rect 2850 7987 2855 7992
rect 2887 7984 2892 7989
rect 2898 7980 2903 7985
rect 2921 7989 2926 7994
rect 2945 7984 2950 7989
rect 2960 7988 2965 7994
rect 2990 7984 2995 7989
rect 3019 7983 3024 7988
rect 2974 7978 2979 7983
rect 3003 7978 3007 7983
rect 3045 7977 3050 7982
rect 3101 8123 3106 8128
rect 3126 8241 3131 8246
rect 3125 8182 3130 8187
rect 3186 8247 3191 8252
rect 3150 8109 3155 8114
rect 3150 8051 3155 8056
rect 2851 7924 2856 7929
rect 2887 7917 2892 7922
rect 2898 7921 2903 7926
rect 2921 7912 2926 7917
rect 2945 7917 2950 7922
rect 2974 7923 2979 7928
rect 3003 7923 3007 7928
rect 2960 7912 2965 7918
rect 2990 7917 2995 7922
rect 3019 7918 3024 7923
rect 3045 7916 3050 7921
rect 2850 7855 2855 7860
rect 2887 7852 2892 7857
rect 2898 7848 2903 7853
rect 2921 7857 2926 7862
rect 2945 7852 2950 7857
rect 2960 7856 2965 7862
rect 2990 7852 2995 7857
rect 3019 7851 3024 7856
rect 2974 7846 2979 7851
rect 3003 7846 3007 7851
rect 3045 7845 3050 7850
rect 3101 7983 3106 7988
rect 3126 7977 3131 7982
rect 3125 7916 3130 7921
rect 3303 8280 3307 8284
rect 3208 8120 3213 8125
rect 3183 7992 3188 7997
rect 3217 7985 3222 7990
rect 3214 7912 3219 7917
rect 2851 7792 2856 7797
rect 2887 7785 2892 7790
rect 2898 7789 2903 7794
rect 2921 7780 2926 7785
rect 2945 7785 2950 7790
rect 2974 7791 2979 7796
rect 3003 7791 3007 7796
rect 2960 7780 2965 7786
rect 2990 7785 2995 7790
rect 3019 7786 3024 7791
rect 3044 7780 3049 7785
rect 3101 7859 3106 7864
rect 3089 7791 3094 7796
rect 3148 7785 3153 7790
rect 3159 7789 3164 7794
rect 3182 7780 3187 7785
rect 3206 7785 3211 7790
rect 3235 7791 3240 7796
rect 3264 7791 3268 7796
rect 3221 7780 3226 7786
rect 3251 7785 3256 7790
rect 3276 7791 3281 7796
rect 3312 7792 3316 7796
rect 3150 7680 3154 7684
rect 3701 8407 3705 8411
rect 3569 8296 3573 8300
rect 3275 7598 3279 7602
rect 3568 8192 3572 8196
rect 3701 7425 3705 7429
rect 4479 9486 4483 9490
rect 4489 9486 4493 9490
rect 4499 9486 4503 9490
rect 4509 9486 4513 9490
rect 4479 9481 4483 9485
rect 4489 9481 4493 9485
rect 4499 9481 4503 9485
rect 4509 9481 4513 9485
rect 4479 9476 4483 9480
rect 4489 9476 4493 9480
rect 4499 9476 4503 9480
rect 4509 9476 4513 9480
rect 4479 9471 4483 9475
rect 4489 9471 4493 9475
rect 4499 9471 4503 9475
rect 4509 9471 4513 9475
rect 4525 9486 4529 9490
rect 4535 9486 4539 9490
rect 4545 9486 4549 9490
rect 4555 9486 4559 9490
rect 4525 9481 4529 9485
rect 4535 9481 4539 9485
rect 4545 9481 4549 9485
rect 4555 9481 4559 9485
rect 4525 9476 4529 9480
rect 4535 9476 4539 9480
rect 4545 9476 4549 9480
rect 4555 9476 4559 9480
rect 4525 9471 4529 9475
rect 4535 9471 4539 9475
rect 4545 9471 4549 9475
rect 4555 9471 4559 9475
rect 4479 9457 4483 9461
rect 4489 9457 4493 9461
rect 4499 9457 4503 9461
rect 4509 9457 4513 9461
rect 4479 9452 4483 9456
rect 4489 9452 4493 9456
rect 4499 9452 4503 9456
rect 4509 9452 4513 9456
rect 4479 9447 4483 9451
rect 4489 9447 4493 9451
rect 4499 9447 4503 9451
rect 4509 9447 4513 9451
rect 4479 9442 4483 9446
rect 4489 9442 4493 9446
rect 4499 9442 4503 9446
rect 4509 9442 4513 9446
rect 4525 9457 4529 9461
rect 4535 9457 4539 9461
rect 4545 9457 4549 9461
rect 4555 9457 4559 9461
rect 4525 9452 4529 9456
rect 4535 9452 4539 9456
rect 4545 9452 4549 9456
rect 4555 9452 4559 9456
rect 4525 9447 4529 9451
rect 4535 9447 4539 9451
rect 4545 9447 4549 9451
rect 4555 9447 4559 9451
rect 4525 9442 4529 9446
rect 4535 9442 4539 9446
rect 4545 9442 4549 9446
rect 4555 9442 4559 9446
rect 3792 9313 3796 9317
rect 3832 9230 3837 9235
rect 3843 9226 3848 9231
rect 3866 9235 3871 9240
rect 3890 9230 3895 9235
rect 3905 9234 3910 9240
rect 3935 9230 3940 9235
rect 3964 9229 3969 9234
rect 3919 9224 3924 9229
rect 3948 9224 3952 9229
rect 3990 9223 3995 9228
rect 3796 9170 3801 9175
rect 3832 9163 3837 9168
rect 3843 9167 3848 9172
rect 3866 9158 3871 9163
rect 3890 9163 3895 9168
rect 3919 9169 3924 9174
rect 3948 9169 3952 9174
rect 3905 9158 3910 9164
rect 3935 9163 3940 9168
rect 3964 9164 3969 9169
rect 3990 9164 3995 9169
rect 3795 9101 3800 9106
rect 3832 9098 3837 9103
rect 3843 9094 3848 9099
rect 3866 9103 3871 9108
rect 3890 9098 3895 9103
rect 4046 9229 4051 9234
rect 3905 9102 3910 9108
rect 3935 9098 3940 9103
rect 3964 9097 3969 9102
rect 3919 9092 3924 9097
rect 3948 9092 3952 9097
rect 3990 9091 3995 9096
rect 3796 9038 3801 9043
rect 3832 9031 3837 9036
rect 3843 9035 3848 9040
rect 3866 9026 3871 9031
rect 3890 9031 3895 9036
rect 3919 9037 3924 9042
rect 3948 9037 3952 9042
rect 3905 9026 3910 9032
rect 3935 9031 3940 9036
rect 3964 9032 3969 9037
rect 3989 9033 3994 9038
rect 3795 8969 3800 8974
rect 3832 8966 3837 8971
rect 3843 8962 3848 8967
rect 3866 8971 3871 8976
rect 3890 8966 3895 8971
rect 3905 8970 3910 8976
rect 3935 8966 3940 8971
rect 3964 8965 3969 8970
rect 3919 8960 3924 8965
rect 3948 8960 3952 8965
rect 3990 8959 3995 8964
rect 4046 9105 4051 9110
rect 4071 9223 4076 9228
rect 4070 9164 4075 9169
rect 4131 9229 4136 9234
rect 4095 9091 4100 9096
rect 4095 9033 4100 9038
rect 3796 8906 3801 8911
rect 3832 8899 3837 8904
rect 3843 8903 3848 8908
rect 3866 8894 3871 8899
rect 3890 8899 3895 8904
rect 3919 8905 3924 8910
rect 3948 8905 3952 8910
rect 3905 8894 3910 8900
rect 3935 8899 3940 8904
rect 3964 8900 3969 8905
rect 3990 8898 3995 8903
rect 3795 8837 3800 8842
rect 3832 8834 3837 8839
rect 3843 8830 3848 8835
rect 3866 8839 3871 8844
rect 3890 8834 3895 8839
rect 3905 8838 3910 8844
rect 3935 8834 3940 8839
rect 3964 8833 3969 8838
rect 3919 8828 3924 8833
rect 3948 8828 3952 8833
rect 3990 8827 3995 8832
rect 4046 8965 4051 8970
rect 4071 8959 4076 8964
rect 4070 8898 4075 8903
rect 4248 9262 4252 9266
rect 4153 9102 4158 9107
rect 4479 9056 4483 9060
rect 4489 9056 4493 9060
rect 4499 9056 4503 9060
rect 4509 9056 4513 9060
rect 4479 9051 4483 9055
rect 4489 9051 4493 9055
rect 4499 9051 4503 9055
rect 4509 9051 4513 9055
rect 4479 9046 4483 9050
rect 4489 9046 4493 9050
rect 4499 9046 4503 9050
rect 4509 9046 4513 9050
rect 4479 9041 4483 9045
rect 4489 9041 4493 9045
rect 4499 9041 4503 9045
rect 4509 9041 4513 9045
rect 4525 9056 4529 9060
rect 4535 9056 4539 9060
rect 4545 9056 4549 9060
rect 4555 9056 4559 9060
rect 4525 9051 4529 9055
rect 4535 9051 4539 9055
rect 4545 9051 4549 9055
rect 4555 9051 4559 9055
rect 4525 9046 4529 9050
rect 4535 9046 4539 9050
rect 4545 9046 4549 9050
rect 4555 9046 4559 9050
rect 4525 9041 4529 9045
rect 4535 9041 4539 9045
rect 4545 9041 4549 9045
rect 4555 9041 4559 9045
rect 4128 8974 4133 8979
rect 4162 8967 4167 8972
rect 4159 8894 4164 8899
rect 3796 8774 3801 8779
rect 3832 8767 3837 8772
rect 3843 8771 3848 8776
rect 3866 8762 3871 8767
rect 3890 8767 3895 8772
rect 3919 8773 3924 8778
rect 3948 8773 3952 8778
rect 3905 8762 3910 8768
rect 3935 8767 3940 8772
rect 3964 8768 3969 8773
rect 3989 8762 3994 8767
rect 4046 8841 4051 8846
rect 4034 8773 4039 8778
rect 4093 8767 4098 8772
rect 4104 8771 4109 8776
rect 4127 8762 4132 8767
rect 4151 8767 4156 8772
rect 4180 8773 4185 8778
rect 4209 8773 4213 8778
rect 4166 8762 4171 8768
rect 4196 8767 4201 8772
rect 4221 8773 4226 8778
rect 4479 8747 4483 8751
rect 4489 8747 4493 8751
rect 4499 8747 4503 8751
rect 4509 8747 4513 8751
rect 4479 8742 4483 8746
rect 4489 8742 4493 8746
rect 4499 8742 4503 8746
rect 4509 8742 4513 8746
rect 4479 8737 4483 8741
rect 4489 8737 4493 8741
rect 4499 8737 4503 8741
rect 4509 8737 4513 8741
rect 4479 8732 4483 8736
rect 4489 8732 4493 8736
rect 4499 8732 4503 8736
rect 4509 8732 4513 8736
rect 4525 8747 4529 8751
rect 4535 8747 4539 8751
rect 4545 8747 4549 8751
rect 4555 8747 4559 8751
rect 4525 8742 4529 8746
rect 4535 8742 4539 8746
rect 4545 8742 4549 8746
rect 4555 8742 4559 8746
rect 4525 8737 4529 8741
rect 4535 8737 4539 8741
rect 4545 8737 4549 8741
rect 4555 8737 4559 8741
rect 4525 8732 4529 8736
rect 4535 8732 4539 8736
rect 4545 8732 4549 8736
rect 4555 8732 4559 8736
rect 4095 8662 4099 8666
rect 4220 8580 4224 8584
rect 4479 8438 4483 8442
rect 4489 8438 4493 8442
rect 4499 8438 4503 8442
rect 4509 8438 4513 8442
rect 4479 8433 4483 8437
rect 4489 8433 4493 8437
rect 4499 8433 4503 8437
rect 4509 8433 4513 8437
rect 4479 8428 4483 8432
rect 4489 8428 4493 8432
rect 4499 8428 4503 8432
rect 4509 8428 4513 8432
rect 4479 8423 4483 8427
rect 4489 8423 4493 8427
rect 4499 8423 4503 8427
rect 4509 8423 4513 8427
rect 4525 8438 4529 8442
rect 4535 8438 4539 8442
rect 4545 8438 4549 8442
rect 4555 8438 4559 8442
rect 4525 8433 4529 8437
rect 4535 8433 4539 8437
rect 4545 8433 4549 8437
rect 4555 8433 4559 8437
rect 4525 8428 4529 8432
rect 4535 8428 4539 8432
rect 4545 8428 4549 8432
rect 4555 8428 4559 8432
rect 4525 8423 4529 8427
rect 4535 8423 4539 8427
rect 4545 8423 4549 8427
rect 4555 8423 4559 8427
rect 3792 8331 3796 8335
rect 3832 8248 3837 8253
rect 3843 8244 3848 8249
rect 3866 8253 3871 8258
rect 3890 8248 3895 8253
rect 3905 8252 3910 8258
rect 3935 8248 3940 8253
rect 3964 8247 3969 8252
rect 3919 8242 3924 8247
rect 3948 8242 3952 8247
rect 3990 8241 3995 8246
rect 3796 8188 3801 8193
rect 3832 8181 3837 8186
rect 3843 8185 3848 8190
rect 3866 8176 3871 8181
rect 3890 8181 3895 8186
rect 3919 8187 3924 8192
rect 3948 8187 3952 8192
rect 3905 8176 3910 8182
rect 3935 8181 3940 8186
rect 3964 8182 3969 8187
rect 3990 8182 3995 8187
rect 3795 8119 3800 8124
rect 3832 8116 3837 8121
rect 3843 8112 3848 8117
rect 3866 8121 3871 8126
rect 3890 8116 3895 8121
rect 4046 8247 4051 8252
rect 3905 8120 3910 8126
rect 3935 8116 3940 8121
rect 3964 8115 3969 8120
rect 3919 8110 3924 8115
rect 3948 8110 3952 8115
rect 3990 8109 3995 8114
rect 3796 8056 3801 8061
rect 3832 8049 3837 8054
rect 3843 8053 3848 8058
rect 3866 8044 3871 8049
rect 3890 8049 3895 8054
rect 3919 8055 3924 8060
rect 3948 8055 3952 8060
rect 3905 8044 3910 8050
rect 3935 8049 3940 8054
rect 3964 8050 3969 8055
rect 3989 8051 3994 8056
rect 3795 7987 3800 7992
rect 3832 7984 3837 7989
rect 3843 7980 3848 7985
rect 3866 7989 3871 7994
rect 3890 7984 3895 7989
rect 3905 7988 3910 7994
rect 3935 7984 3940 7989
rect 3964 7983 3969 7988
rect 3919 7978 3924 7983
rect 3948 7978 3952 7983
rect 3990 7977 3995 7982
rect 4046 8123 4051 8128
rect 4071 8241 4076 8246
rect 4070 8182 4075 8187
rect 4131 8247 4136 8252
rect 4095 8109 4100 8114
rect 4095 8051 4100 8056
rect 3796 7924 3801 7929
rect 3832 7917 3837 7922
rect 3843 7921 3848 7926
rect 3866 7912 3871 7917
rect 3890 7917 3895 7922
rect 3919 7923 3924 7928
rect 3948 7923 3952 7928
rect 3905 7912 3910 7918
rect 3935 7917 3940 7922
rect 3964 7918 3969 7923
rect 3990 7916 3995 7921
rect 3795 7855 3800 7860
rect 3832 7852 3837 7857
rect 3843 7848 3848 7853
rect 3866 7857 3871 7862
rect 3890 7852 3895 7857
rect 3905 7856 3910 7862
rect 3935 7852 3940 7857
rect 3964 7851 3969 7856
rect 3919 7846 3924 7851
rect 3948 7846 3952 7851
rect 3990 7845 3995 7850
rect 4046 7983 4051 7988
rect 4071 7977 4076 7982
rect 4070 7916 4075 7921
rect 4248 8280 4252 8284
rect 4479 8129 4483 8133
rect 4489 8129 4493 8133
rect 4499 8129 4503 8133
rect 4509 8129 4513 8133
rect 4153 8120 4158 8125
rect 4479 8124 4483 8128
rect 4489 8124 4493 8128
rect 4499 8124 4503 8128
rect 4509 8124 4513 8128
rect 4479 8119 4483 8123
rect 4489 8119 4493 8123
rect 4499 8119 4503 8123
rect 4509 8119 4513 8123
rect 4479 8114 4483 8118
rect 4489 8114 4493 8118
rect 4499 8114 4503 8118
rect 4509 8114 4513 8118
rect 4525 8129 4529 8133
rect 4535 8129 4539 8133
rect 4545 8129 4549 8133
rect 4555 8129 4559 8133
rect 4525 8124 4529 8128
rect 4535 8124 4539 8128
rect 4545 8124 4549 8128
rect 4555 8124 4559 8128
rect 4525 8119 4529 8123
rect 4535 8119 4539 8123
rect 4545 8119 4549 8123
rect 4555 8119 4559 8123
rect 4525 8114 4529 8118
rect 4535 8114 4539 8118
rect 4545 8114 4549 8118
rect 4555 8114 4559 8118
rect 4479 8098 4483 8102
rect 4489 8098 4493 8102
rect 4499 8098 4503 8102
rect 4509 8098 4513 8102
rect 4479 8093 4483 8097
rect 4489 8093 4493 8097
rect 4499 8093 4503 8097
rect 4509 8093 4513 8097
rect 4479 8088 4483 8092
rect 4489 8088 4493 8092
rect 4499 8088 4503 8092
rect 4509 8088 4513 8092
rect 4479 8083 4483 8087
rect 4489 8083 4493 8087
rect 4499 8083 4503 8087
rect 4509 8083 4513 8087
rect 4525 8098 4529 8102
rect 4535 8098 4539 8102
rect 4545 8098 4549 8102
rect 4555 8098 4559 8102
rect 4525 8093 4529 8097
rect 4535 8093 4539 8097
rect 4545 8093 4549 8097
rect 4555 8093 4559 8097
rect 4525 8088 4529 8092
rect 4535 8088 4539 8092
rect 4545 8088 4549 8092
rect 4555 8088 4559 8092
rect 4525 8083 4529 8087
rect 4535 8083 4539 8087
rect 4545 8083 4549 8087
rect 4555 8083 4559 8087
rect 4496 8074 4500 8078
rect 4501 8074 4505 8078
rect 4496 8069 4500 8073
rect 4501 8069 4505 8073
rect 4496 8064 4500 8068
rect 4501 8064 4505 8068
rect 4496 8059 4500 8063
rect 4501 8059 4505 8063
rect 4496 8054 4500 8058
rect 4501 8054 4505 8058
rect 4496 8049 4500 8053
rect 4501 8049 4505 8053
rect 4496 8044 4500 8048
rect 4501 8044 4505 8048
rect 4496 8039 4500 8043
rect 4501 8039 4505 8043
rect 4496 8034 4500 8038
rect 4501 8034 4505 8038
rect 4496 8029 4500 8033
rect 4501 8029 4505 8033
rect 4496 8024 4500 8028
rect 4501 8024 4505 8028
rect 4128 7992 4133 7997
rect 4162 7985 4167 7990
rect 4159 7912 4164 7917
rect 3796 7792 3801 7797
rect 3832 7785 3837 7790
rect 3843 7789 3848 7794
rect 3866 7780 3871 7785
rect 3890 7785 3895 7790
rect 3919 7791 3924 7796
rect 3948 7791 3952 7796
rect 3905 7780 3910 7786
rect 3935 7785 3940 7790
rect 3964 7786 3969 7791
rect 3989 7780 3994 7785
rect 4046 7859 4051 7864
rect 4034 7791 4039 7796
rect 4093 7785 4098 7790
rect 4104 7789 4109 7794
rect 4127 7780 4132 7785
rect 4151 7785 4156 7790
rect 4180 7791 4185 7796
rect 4209 7791 4213 7796
rect 4166 7780 4171 7786
rect 4196 7785 4201 7790
rect 4221 7791 4226 7796
rect 4095 7680 4099 7684
rect 4220 7598 4224 7602
rect 4529 7814 4533 7818
rect 4534 7814 4538 7818
rect 4539 7814 4543 7818
rect 4544 7814 4548 7818
rect 4549 7814 4553 7818
rect 4554 7814 4558 7818
rect 4559 7814 4563 7818
rect 4564 7814 4568 7818
rect 4569 7814 4573 7818
rect 4574 7814 4578 7818
rect 4579 7814 4583 7818
rect 4584 7814 4588 7818
rect 4589 7814 4593 7818
rect 4529 7809 4533 7813
rect 4534 7809 4538 7813
rect 4539 7809 4543 7813
rect 4544 7809 4548 7813
rect 4549 7809 4553 7813
rect 4554 7809 4558 7813
rect 4559 7809 4563 7813
rect 4564 7809 4568 7813
rect 4569 7809 4573 7813
rect 4574 7809 4578 7813
rect 4579 7809 4583 7813
rect 4584 7809 4588 7813
rect 4589 7809 4593 7813
rect 4479 7789 4483 7793
rect 4489 7789 4493 7793
rect 4499 7789 4503 7793
rect 4509 7789 4513 7793
rect 4479 7784 4483 7788
rect 4489 7784 4493 7788
rect 4499 7784 4503 7788
rect 4509 7784 4513 7788
rect 4479 7779 4483 7783
rect 4489 7779 4493 7783
rect 4499 7779 4503 7783
rect 4509 7779 4513 7783
rect 4479 7774 4483 7778
rect 4489 7774 4493 7778
rect 4499 7774 4503 7778
rect 4509 7774 4513 7778
rect 4525 7789 4529 7793
rect 4535 7789 4539 7793
rect 4545 7789 4549 7793
rect 4555 7789 4559 7793
rect 4525 7784 4529 7788
rect 4535 7784 4539 7788
rect 4545 7784 4549 7788
rect 4555 7784 4559 7788
rect 4525 7779 4529 7783
rect 4535 7779 4539 7783
rect 4545 7779 4549 7783
rect 4555 7779 4559 7783
rect 4525 7774 4529 7778
rect 4535 7774 4539 7778
rect 4545 7774 4549 7778
rect 4555 7774 4559 7778
rect 4529 7499 4533 7503
rect 4534 7499 4538 7503
rect 4539 7499 4543 7503
rect 4544 7499 4548 7503
rect 4549 7499 4553 7503
rect 4554 7499 4558 7503
rect 4559 7499 4563 7503
rect 4564 7499 4568 7503
rect 4569 7499 4573 7503
rect 4574 7499 4578 7503
rect 4579 7499 4583 7503
rect 4584 7499 4588 7503
rect 4589 7499 4593 7503
rect 613 7158 617 7162
rect 623 7158 627 7162
rect 633 7158 637 7162
rect 643 7158 647 7162
rect 659 7158 663 7162
rect 669 7158 673 7162
rect 679 7158 683 7162
rect 689 7158 693 7162
rect 613 7123 617 7127
rect 623 7123 627 7127
rect 633 7123 637 7127
rect 643 7123 647 7127
rect 613 7118 617 7122
rect 623 7118 627 7122
rect 633 7118 637 7122
rect 643 7118 647 7122
rect 613 7113 617 7117
rect 623 7113 627 7117
rect 633 7113 637 7117
rect 643 7113 647 7117
rect 613 7108 617 7112
rect 623 7108 627 7112
rect 633 7108 637 7112
rect 643 7108 647 7112
rect 659 7123 663 7127
rect 669 7123 673 7127
rect 679 7123 683 7127
rect 689 7123 693 7127
rect 659 7118 663 7122
rect 669 7118 673 7122
rect 679 7118 683 7122
rect 689 7118 693 7122
rect 659 7113 663 7117
rect 669 7113 673 7117
rect 679 7113 683 7117
rect 689 7113 693 7117
rect 659 7108 663 7112
rect 669 7108 673 7112
rect 679 7108 683 7112
rect 689 7108 693 7112
rect 613 6536 617 6540
rect 623 6536 627 6540
rect 633 6536 637 6540
rect 643 6536 647 6540
rect 613 6531 617 6535
rect 623 6531 627 6535
rect 633 6531 637 6535
rect 643 6531 647 6535
rect 613 6526 617 6530
rect 623 6526 627 6530
rect 633 6526 637 6530
rect 643 6526 647 6530
rect 613 6521 617 6525
rect 623 6521 627 6525
rect 633 6521 637 6525
rect 643 6521 647 6525
rect 659 6536 663 6540
rect 669 6536 673 6540
rect 679 6536 683 6540
rect 689 6536 693 6540
rect 659 6531 663 6535
rect 669 6531 673 6535
rect 679 6531 683 6535
rect 689 6531 693 6535
rect 659 6526 663 6530
rect 669 6526 673 6530
rect 679 6526 683 6530
rect 689 6526 693 6530
rect 659 6521 663 6525
rect 669 6521 673 6525
rect 679 6521 683 6525
rect 689 6521 693 6525
rect 579 6501 583 6505
rect 584 6501 588 6505
rect 589 6501 593 6505
rect 594 6501 598 6505
rect 599 6501 603 6505
rect 604 6501 608 6505
rect 609 6501 613 6505
rect 614 6501 618 6505
rect 619 6501 623 6505
rect 624 6501 628 6505
rect 629 6501 633 6505
rect 634 6501 638 6505
rect 639 6501 643 6505
rect 579 6496 583 6500
rect 584 6496 588 6500
rect 589 6496 593 6500
rect 594 6496 598 6500
rect 599 6496 603 6500
rect 604 6496 608 6500
rect 609 6496 613 6500
rect 614 6496 618 6500
rect 619 6496 623 6500
rect 624 6496 628 6500
rect 629 6496 633 6500
rect 634 6496 638 6500
rect 639 6496 643 6500
rect 948 6712 952 6716
rect 1073 6630 1077 6634
rect 946 6518 951 6523
rect 971 6524 976 6529
rect 1001 6528 1006 6534
rect 959 6518 963 6523
rect 987 6518 992 6523
rect 1016 6524 1021 6529
rect 1040 6529 1045 6534
rect 1063 6520 1068 6525
rect 1074 6524 1079 6529
rect 1133 6518 1138 6523
rect 1121 6450 1126 6455
rect 1178 6529 1183 6534
rect 1203 6523 1208 6528
rect 1232 6524 1237 6529
rect 1262 6528 1267 6534
rect 1220 6518 1224 6523
rect 1248 6518 1253 6523
rect 1277 6524 1282 6529
rect 1301 6529 1306 6534
rect 1324 6520 1329 6525
rect 1335 6524 1340 6529
rect 1371 6517 1376 6522
rect 1008 6397 1013 6402
rect 1005 6324 1010 6329
rect 1039 6317 1044 6322
rect 667 6286 671 6290
rect 672 6286 676 6290
rect 667 6281 671 6285
rect 672 6281 676 6285
rect 667 6276 671 6280
rect 672 6276 676 6280
rect 667 6271 671 6275
rect 672 6271 676 6275
rect 667 6266 671 6270
rect 672 6266 676 6270
rect 667 6261 671 6265
rect 672 6261 676 6265
rect 667 6256 671 6260
rect 672 6256 676 6260
rect 667 6251 671 6255
rect 672 6251 676 6255
rect 667 6246 671 6250
rect 672 6246 676 6250
rect 667 6241 671 6245
rect 672 6241 676 6245
rect 667 6236 671 6240
rect 672 6236 676 6240
rect 613 6227 617 6231
rect 623 6227 627 6231
rect 633 6227 637 6231
rect 643 6227 647 6231
rect 613 6222 617 6226
rect 623 6222 627 6226
rect 633 6222 637 6226
rect 643 6222 647 6226
rect 613 6217 617 6221
rect 623 6217 627 6221
rect 633 6217 637 6221
rect 643 6217 647 6221
rect 613 6212 617 6216
rect 623 6212 627 6216
rect 633 6212 637 6216
rect 643 6212 647 6216
rect 659 6227 663 6231
rect 669 6227 673 6231
rect 679 6227 683 6231
rect 689 6227 693 6231
rect 659 6222 663 6226
rect 669 6222 673 6226
rect 679 6222 683 6226
rect 689 6222 693 6226
rect 659 6217 663 6221
rect 669 6217 673 6221
rect 679 6217 683 6221
rect 689 6217 693 6221
rect 659 6212 663 6216
rect 669 6212 673 6216
rect 679 6212 683 6216
rect 689 6212 693 6216
rect 613 6196 617 6200
rect 623 6196 627 6200
rect 633 6196 637 6200
rect 643 6196 647 6200
rect 613 6191 617 6195
rect 623 6191 627 6195
rect 633 6191 637 6195
rect 643 6191 647 6195
rect 613 6186 617 6190
rect 623 6186 627 6190
rect 633 6186 637 6190
rect 643 6186 647 6190
rect 613 6181 617 6185
rect 623 6181 627 6185
rect 633 6181 637 6185
rect 643 6181 647 6185
rect 659 6196 663 6200
rect 669 6196 673 6200
rect 679 6196 683 6200
rect 689 6196 693 6200
rect 659 6191 663 6195
rect 669 6191 673 6195
rect 679 6191 683 6195
rect 689 6191 693 6195
rect 659 6186 663 6190
rect 669 6186 673 6190
rect 679 6186 683 6190
rect 689 6186 693 6190
rect 1014 6189 1019 6194
rect 659 6181 663 6185
rect 669 6181 673 6185
rect 679 6181 683 6185
rect 689 6181 693 6185
rect 920 6030 924 6034
rect 1097 6393 1102 6398
rect 1096 6332 1101 6337
rect 1121 6326 1126 6331
rect 1177 6464 1182 6469
rect 1220 6463 1224 6468
rect 1248 6463 1253 6468
rect 1203 6458 1208 6463
rect 1232 6457 1237 6462
rect 1262 6452 1267 6458
rect 1277 6457 1282 6462
rect 1301 6452 1306 6457
rect 1324 6461 1329 6466
rect 1335 6457 1340 6462
rect 1372 6454 1377 6459
rect 1177 6393 1182 6398
rect 1203 6391 1208 6396
rect 1232 6392 1237 6397
rect 1262 6396 1267 6402
rect 1220 6386 1224 6391
rect 1248 6386 1253 6391
rect 1277 6392 1282 6397
rect 1301 6397 1306 6402
rect 1324 6388 1329 6393
rect 1335 6392 1340 6397
rect 1371 6385 1376 6390
rect 1072 6258 1077 6263
rect 1072 6200 1077 6205
rect 1036 6062 1041 6067
rect 1097 6127 1102 6132
rect 1096 6068 1101 6073
rect 1121 6186 1126 6191
rect 1177 6332 1182 6337
rect 1220 6331 1224 6336
rect 1248 6331 1253 6336
rect 1203 6326 1208 6331
rect 1232 6325 1237 6330
rect 1262 6320 1267 6326
rect 1277 6325 1282 6330
rect 1301 6320 1306 6325
rect 1324 6329 1329 6334
rect 1335 6325 1340 6330
rect 1372 6322 1377 6327
rect 1178 6258 1183 6263
rect 1203 6259 1208 6264
rect 1232 6260 1237 6265
rect 1262 6264 1267 6270
rect 1220 6254 1224 6259
rect 1248 6254 1253 6259
rect 1277 6260 1282 6265
rect 1301 6265 1306 6270
rect 1324 6256 1329 6261
rect 1335 6260 1340 6265
rect 1371 6253 1376 6258
rect 1177 6200 1182 6205
rect 1220 6199 1224 6204
rect 1248 6199 1253 6204
rect 1203 6194 1208 6199
rect 1232 6193 1237 6198
rect 1262 6188 1267 6194
rect 1121 6062 1126 6067
rect 1277 6193 1282 6198
rect 1301 6188 1306 6193
rect 1324 6197 1329 6202
rect 1335 6193 1340 6198
rect 1372 6190 1377 6195
rect 1177 6127 1182 6132
rect 1203 6127 1208 6132
rect 1232 6128 1237 6133
rect 1262 6132 1267 6138
rect 1220 6122 1224 6127
rect 1248 6122 1253 6127
rect 1277 6128 1282 6133
rect 1301 6133 1306 6138
rect 1324 6124 1329 6129
rect 1335 6128 1340 6133
rect 1371 6121 1376 6126
rect 1177 6068 1182 6073
rect 1220 6067 1224 6072
rect 1248 6067 1253 6072
rect 1203 6062 1208 6067
rect 1232 6061 1237 6066
rect 1262 6056 1267 6062
rect 1277 6061 1282 6066
rect 1301 6056 1306 6061
rect 1324 6065 1329 6070
rect 1335 6061 1340 6066
rect 1376 5979 1380 5983
rect 613 5887 617 5891
rect 623 5887 627 5891
rect 633 5887 637 5891
rect 643 5887 647 5891
rect 613 5882 617 5886
rect 623 5882 627 5886
rect 633 5882 637 5886
rect 643 5882 647 5886
rect 613 5877 617 5881
rect 623 5877 627 5881
rect 633 5877 637 5881
rect 643 5877 647 5881
rect 613 5872 617 5876
rect 623 5872 627 5876
rect 633 5872 637 5876
rect 643 5872 647 5876
rect 659 5887 663 5891
rect 669 5887 673 5891
rect 679 5887 683 5891
rect 689 5887 693 5891
rect 659 5882 663 5886
rect 669 5882 673 5886
rect 679 5882 683 5886
rect 689 5882 693 5886
rect 659 5877 663 5881
rect 669 5877 673 5881
rect 679 5877 683 5881
rect 689 5877 693 5881
rect 659 5872 663 5876
rect 669 5872 673 5876
rect 679 5872 683 5876
rect 689 5872 693 5876
rect 948 5730 952 5734
rect 1073 5648 1077 5652
rect 613 5578 617 5582
rect 623 5578 627 5582
rect 633 5578 637 5582
rect 643 5578 647 5582
rect 613 5573 617 5577
rect 623 5573 627 5577
rect 633 5573 637 5577
rect 643 5573 647 5577
rect 613 5568 617 5572
rect 623 5568 627 5572
rect 633 5568 637 5572
rect 643 5568 647 5572
rect 613 5563 617 5567
rect 623 5563 627 5567
rect 633 5563 637 5567
rect 643 5563 647 5567
rect 659 5578 663 5582
rect 669 5578 673 5582
rect 679 5578 683 5582
rect 689 5578 693 5582
rect 659 5573 663 5577
rect 669 5573 673 5577
rect 679 5573 683 5577
rect 689 5573 693 5577
rect 659 5568 663 5572
rect 669 5568 673 5572
rect 679 5568 683 5572
rect 689 5568 693 5572
rect 659 5563 663 5567
rect 669 5563 673 5567
rect 679 5563 683 5567
rect 689 5563 693 5567
rect 946 5536 951 5541
rect 971 5542 976 5547
rect 1001 5546 1006 5552
rect 959 5536 963 5541
rect 987 5536 992 5541
rect 1016 5542 1021 5547
rect 1040 5547 1045 5552
rect 1063 5538 1068 5543
rect 1074 5542 1079 5547
rect 1133 5536 1138 5541
rect 1121 5468 1126 5473
rect 1178 5547 1183 5552
rect 1203 5541 1208 5546
rect 1232 5542 1237 5547
rect 1262 5546 1267 5552
rect 1220 5536 1224 5541
rect 1248 5536 1253 5541
rect 1277 5542 1282 5547
rect 1301 5547 1306 5552
rect 1324 5538 1329 5543
rect 1335 5542 1340 5547
rect 1371 5535 1376 5540
rect 1008 5415 1013 5420
rect 1005 5342 1010 5347
rect 1039 5335 1044 5340
rect 613 5269 617 5273
rect 623 5269 627 5273
rect 633 5269 637 5273
rect 643 5269 647 5273
rect 613 5264 617 5268
rect 623 5264 627 5268
rect 633 5264 637 5268
rect 643 5264 647 5268
rect 613 5259 617 5263
rect 623 5259 627 5263
rect 633 5259 637 5263
rect 643 5259 647 5263
rect 613 5254 617 5258
rect 623 5254 627 5258
rect 633 5254 637 5258
rect 643 5254 647 5258
rect 659 5269 663 5273
rect 669 5269 673 5273
rect 679 5269 683 5273
rect 689 5269 693 5273
rect 659 5264 663 5268
rect 669 5264 673 5268
rect 679 5264 683 5268
rect 689 5264 693 5268
rect 659 5259 663 5263
rect 669 5259 673 5263
rect 679 5259 683 5263
rect 689 5259 693 5263
rect 659 5254 663 5258
rect 669 5254 673 5258
rect 679 5254 683 5258
rect 689 5254 693 5258
rect 1014 5207 1019 5212
rect 920 5048 924 5052
rect 1097 5411 1102 5416
rect 1096 5350 1101 5355
rect 1121 5344 1126 5349
rect 1177 5482 1182 5487
rect 1220 5481 1224 5486
rect 1248 5481 1253 5486
rect 1203 5476 1208 5481
rect 1232 5475 1237 5480
rect 1262 5470 1267 5476
rect 1277 5475 1282 5480
rect 1301 5470 1306 5475
rect 1324 5479 1329 5484
rect 1335 5475 1340 5480
rect 1372 5472 1377 5477
rect 1177 5411 1182 5416
rect 1203 5409 1208 5414
rect 1232 5410 1237 5415
rect 1262 5414 1267 5420
rect 1220 5404 1224 5409
rect 1248 5404 1253 5409
rect 1277 5410 1282 5415
rect 1301 5415 1306 5420
rect 1324 5406 1329 5411
rect 1335 5410 1340 5415
rect 1371 5403 1376 5408
rect 1072 5276 1077 5281
rect 1072 5218 1077 5223
rect 1036 5080 1041 5085
rect 1097 5145 1102 5150
rect 1096 5086 1101 5091
rect 1121 5204 1126 5209
rect 1177 5350 1182 5355
rect 1220 5349 1224 5354
rect 1248 5349 1253 5354
rect 1203 5344 1208 5349
rect 1232 5343 1237 5348
rect 1262 5338 1267 5344
rect 1277 5343 1282 5348
rect 1301 5338 1306 5343
rect 1324 5347 1329 5352
rect 1335 5343 1340 5348
rect 1372 5340 1377 5345
rect 1178 5276 1183 5281
rect 1203 5277 1208 5282
rect 1232 5278 1237 5283
rect 1262 5282 1267 5288
rect 1220 5272 1224 5277
rect 1248 5272 1253 5277
rect 1277 5278 1282 5283
rect 1301 5283 1306 5288
rect 1324 5274 1329 5279
rect 1335 5278 1340 5283
rect 1371 5271 1376 5276
rect 1177 5218 1182 5223
rect 1220 5217 1224 5222
rect 1248 5217 1253 5222
rect 1203 5212 1208 5217
rect 1232 5211 1237 5216
rect 1262 5206 1267 5212
rect 1121 5080 1126 5085
rect 1277 5211 1282 5216
rect 1301 5206 1306 5211
rect 1324 5215 1329 5220
rect 1335 5211 1340 5216
rect 1372 5208 1377 5213
rect 1177 5145 1182 5150
rect 1203 5145 1208 5150
rect 1232 5146 1237 5151
rect 1262 5150 1267 5156
rect 1220 5140 1224 5145
rect 1248 5140 1253 5145
rect 1277 5146 1282 5151
rect 1301 5151 1306 5156
rect 1324 5142 1329 5147
rect 1335 5146 1340 5151
rect 1371 5139 1376 5144
rect 1177 5086 1182 5091
rect 1220 5085 1224 5090
rect 1248 5085 1253 5090
rect 1203 5080 1208 5085
rect 1232 5079 1237 5084
rect 1262 5074 1267 5080
rect 1277 5079 1282 5084
rect 1301 5074 1306 5079
rect 1324 5083 1329 5088
rect 1335 5079 1340 5084
rect 1376 4997 1380 5001
rect 613 4868 617 4872
rect 623 4868 627 4872
rect 633 4868 637 4872
rect 643 4868 647 4872
rect 613 4863 617 4867
rect 623 4863 627 4867
rect 633 4863 637 4867
rect 643 4863 647 4867
rect 613 4858 617 4862
rect 623 4858 627 4862
rect 633 4858 637 4862
rect 643 4858 647 4862
rect 613 4853 617 4857
rect 623 4853 627 4857
rect 633 4853 637 4857
rect 643 4853 647 4857
rect 659 4868 663 4872
rect 669 4868 673 4872
rect 679 4868 683 4872
rect 689 4868 693 4872
rect 659 4863 663 4867
rect 669 4863 673 4867
rect 679 4863 683 4867
rect 689 4863 693 4867
rect 659 4858 663 4862
rect 669 4858 673 4862
rect 679 4858 683 4862
rect 689 4858 693 4862
rect 659 4853 663 4857
rect 669 4853 673 4857
rect 679 4853 683 4857
rect 689 4853 693 4857
rect 613 4839 617 4843
rect 623 4839 627 4843
rect 633 4839 637 4843
rect 643 4839 647 4843
rect 613 4834 617 4838
rect 623 4834 627 4838
rect 633 4834 637 4838
rect 643 4834 647 4838
rect 613 4829 617 4833
rect 623 4829 627 4833
rect 633 4829 637 4833
rect 643 4829 647 4833
rect 613 4824 617 4828
rect 623 4824 627 4828
rect 633 4824 637 4828
rect 643 4824 647 4828
rect 659 4839 663 4843
rect 669 4839 673 4843
rect 679 4839 683 4843
rect 689 4839 693 4843
rect 659 4834 663 4838
rect 669 4834 673 4838
rect 679 4834 683 4838
rect 689 4834 693 4838
rect 659 4829 663 4833
rect 669 4829 673 4833
rect 679 4829 683 4833
rect 689 4829 693 4833
rect 659 4824 663 4828
rect 669 4824 673 4828
rect 679 4824 683 4828
rect 689 4824 693 4828
rect 1467 6885 1471 6889
rect 1600 6118 1604 6122
rect 1893 6712 1897 6716
rect 1599 6014 1603 6018
rect 1467 5903 1471 5907
rect 2018 6630 2022 6634
rect 1856 6518 1860 6522
rect 1891 6518 1896 6523
rect 1916 6524 1921 6529
rect 1946 6528 1951 6534
rect 1904 6518 1908 6523
rect 1932 6518 1937 6523
rect 1961 6524 1966 6529
rect 1985 6529 1990 6534
rect 2008 6520 2013 6525
rect 2019 6524 2024 6529
rect 2078 6518 2083 6523
rect 2066 6450 2071 6455
rect 2123 6529 2128 6534
rect 2148 6523 2153 6528
rect 2177 6524 2182 6529
rect 2207 6528 2212 6534
rect 2165 6518 2169 6523
rect 2193 6518 2198 6523
rect 2222 6524 2227 6529
rect 2246 6529 2251 6534
rect 2269 6520 2274 6525
rect 2280 6524 2285 6529
rect 2316 6517 2321 6522
rect 1953 6397 1958 6402
rect 1950 6324 1955 6329
rect 1984 6317 1989 6322
rect 1959 6189 1964 6194
rect 1865 6030 1869 6034
rect 2042 6393 2047 6398
rect 2041 6332 2046 6337
rect 2066 6326 2071 6331
rect 2122 6464 2127 6469
rect 2165 6463 2169 6468
rect 2193 6463 2198 6468
rect 2148 6458 2153 6463
rect 2177 6457 2182 6462
rect 2207 6452 2212 6458
rect 2222 6457 2227 6462
rect 2246 6452 2251 6457
rect 2269 6461 2274 6466
rect 2280 6457 2285 6462
rect 2317 6454 2322 6459
rect 2122 6393 2127 6398
rect 2148 6391 2153 6396
rect 2177 6392 2182 6397
rect 2207 6396 2212 6402
rect 2165 6386 2169 6391
rect 2193 6386 2198 6391
rect 2222 6392 2227 6397
rect 2246 6397 2251 6402
rect 2269 6388 2274 6393
rect 2280 6392 2285 6397
rect 2316 6385 2321 6390
rect 2017 6258 2022 6263
rect 2017 6200 2022 6205
rect 1981 6062 1986 6067
rect 2042 6127 2047 6132
rect 2041 6068 2046 6073
rect 2066 6186 2071 6191
rect 2122 6332 2127 6337
rect 2165 6331 2169 6336
rect 2193 6331 2198 6336
rect 2148 6326 2153 6331
rect 2177 6325 2182 6330
rect 2207 6320 2212 6326
rect 2222 6325 2227 6330
rect 2246 6320 2251 6325
rect 2269 6329 2274 6334
rect 2280 6325 2285 6330
rect 2317 6322 2322 6327
rect 2123 6258 2128 6263
rect 2148 6259 2153 6264
rect 2177 6260 2182 6265
rect 2207 6264 2212 6270
rect 2165 6254 2169 6259
rect 2193 6254 2198 6259
rect 2222 6260 2227 6265
rect 2246 6265 2251 6270
rect 2269 6256 2274 6261
rect 2280 6260 2285 6265
rect 2316 6253 2321 6258
rect 2122 6200 2127 6205
rect 2165 6199 2169 6204
rect 2193 6199 2198 6204
rect 2148 6194 2153 6199
rect 2177 6193 2182 6198
rect 2207 6188 2212 6194
rect 2066 6062 2071 6067
rect 2222 6193 2227 6198
rect 2246 6188 2251 6193
rect 2269 6197 2274 6202
rect 2280 6193 2285 6198
rect 2317 6190 2322 6195
rect 2122 6127 2127 6132
rect 2148 6127 2153 6132
rect 2177 6128 2182 6133
rect 2207 6132 2212 6138
rect 2165 6122 2169 6127
rect 2193 6122 2198 6127
rect 2222 6128 2227 6133
rect 2246 6133 2251 6138
rect 2269 6124 2274 6129
rect 2280 6128 2285 6133
rect 2316 6121 2321 6126
rect 2122 6068 2127 6073
rect 2165 6067 2169 6072
rect 2193 6067 2198 6072
rect 2148 6062 2153 6067
rect 2177 6061 2182 6066
rect 2207 6056 2212 6062
rect 2222 6061 2227 6066
rect 2246 6056 2251 6061
rect 2269 6065 2274 6070
rect 2280 6061 2285 6066
rect 2321 5979 2325 5983
rect 1893 5730 1897 5734
rect 1607 5491 1612 5496
rect 2018 5648 2022 5652
rect 1856 5536 1860 5540
rect 1724 5490 1729 5495
rect 1891 5536 1896 5541
rect 1916 5542 1921 5547
rect 1946 5546 1951 5552
rect 1904 5536 1908 5541
rect 1932 5536 1937 5541
rect 1961 5542 1966 5547
rect 1985 5547 1990 5552
rect 2008 5538 2013 5543
rect 2019 5542 2024 5547
rect 2078 5536 2083 5541
rect 2066 5468 2071 5473
rect 2123 5547 2128 5552
rect 2148 5541 2153 5546
rect 2177 5542 2182 5547
rect 2207 5546 2212 5552
rect 2165 5536 2169 5541
rect 2193 5536 2198 5541
rect 2222 5542 2227 5547
rect 2246 5547 2251 5552
rect 2269 5538 2274 5543
rect 2280 5542 2285 5547
rect 2316 5535 2321 5540
rect 1953 5415 1958 5420
rect 1950 5342 1955 5347
rect 1984 5335 1989 5340
rect 1607 5173 1612 5178
rect 1724 5174 1729 5179
rect 1600 5136 1604 5140
rect 1599 5033 1603 5037
rect 1959 5207 1964 5212
rect 1865 5048 1869 5052
rect 2042 5411 2047 5416
rect 2041 5350 2046 5355
rect 2066 5344 2071 5349
rect 2122 5482 2127 5487
rect 2165 5481 2169 5486
rect 2193 5481 2198 5486
rect 2148 5476 2153 5481
rect 2177 5475 2182 5480
rect 2207 5470 2212 5476
rect 2222 5475 2227 5480
rect 2246 5470 2251 5475
rect 2269 5479 2274 5484
rect 2280 5475 2285 5480
rect 2317 5472 2322 5477
rect 2122 5411 2127 5416
rect 2148 5409 2153 5414
rect 2177 5410 2182 5415
rect 2207 5414 2212 5420
rect 2165 5404 2169 5409
rect 2193 5404 2198 5409
rect 2222 5410 2227 5415
rect 2246 5415 2251 5420
rect 2269 5406 2274 5411
rect 2280 5410 2285 5415
rect 2316 5403 2321 5408
rect 2017 5276 2022 5281
rect 2017 5218 2022 5223
rect 1981 5080 1986 5085
rect 2042 5145 2047 5150
rect 2041 5086 2046 5091
rect 2066 5204 2071 5209
rect 2122 5350 2127 5355
rect 2165 5349 2169 5354
rect 2193 5349 2198 5354
rect 2148 5344 2153 5349
rect 2177 5343 2182 5348
rect 2207 5338 2212 5344
rect 2222 5343 2227 5348
rect 2246 5338 2251 5343
rect 2269 5347 2274 5352
rect 2280 5343 2285 5348
rect 2317 5340 2322 5345
rect 2123 5276 2128 5281
rect 2148 5277 2153 5282
rect 2177 5278 2182 5283
rect 2207 5282 2212 5288
rect 2165 5272 2169 5277
rect 2193 5272 2198 5277
rect 2222 5278 2227 5283
rect 2246 5283 2251 5288
rect 2269 5274 2274 5279
rect 2280 5278 2285 5283
rect 2316 5271 2321 5276
rect 2122 5218 2127 5223
rect 2165 5217 2169 5222
rect 2193 5217 2198 5222
rect 2148 5212 2153 5217
rect 2177 5211 2182 5216
rect 2207 5206 2212 5212
rect 2066 5080 2071 5085
rect 2222 5211 2227 5216
rect 2246 5206 2251 5211
rect 2269 5215 2274 5220
rect 2280 5211 2285 5216
rect 2317 5208 2322 5213
rect 2122 5145 2127 5150
rect 2148 5145 2153 5150
rect 2177 5146 2182 5151
rect 2207 5150 2212 5156
rect 2165 5140 2169 5145
rect 2193 5140 2198 5145
rect 2222 5146 2227 5151
rect 2246 5151 2251 5156
rect 2269 5142 2274 5147
rect 2280 5146 2285 5151
rect 2316 5139 2321 5144
rect 2122 5086 2127 5091
rect 2165 5085 2169 5090
rect 2193 5085 2198 5090
rect 2148 5080 2153 5085
rect 2177 5079 2182 5084
rect 2207 5074 2212 5080
rect 2222 5079 2227 5084
rect 2246 5074 2251 5079
rect 2269 5083 2274 5088
rect 2280 5079 2285 5084
rect 2321 4997 2325 5001
rect 613 4810 617 4814
rect 623 4810 627 4814
rect 633 4810 637 4814
rect 643 4810 647 4814
rect 613 4805 617 4809
rect 623 4805 627 4809
rect 633 4805 637 4809
rect 643 4805 647 4809
rect 613 4800 617 4804
rect 623 4800 627 4804
rect 633 4800 637 4804
rect 643 4800 647 4804
rect 613 4795 617 4799
rect 623 4795 627 4799
rect 633 4795 637 4799
rect 643 4795 647 4799
rect 659 4810 663 4814
rect 669 4810 673 4814
rect 679 4810 683 4814
rect 689 4810 693 4814
rect 659 4805 663 4809
rect 669 4805 673 4809
rect 679 4805 683 4809
rect 689 4805 693 4809
rect 659 4800 663 4804
rect 669 4800 673 4804
rect 679 4800 683 4804
rect 689 4800 693 4804
rect 659 4795 663 4799
rect 669 4795 673 4799
rect 679 4795 683 4799
rect 689 4795 693 4799
rect 613 4781 617 4785
rect 623 4781 627 4785
rect 633 4781 637 4785
rect 643 4781 647 4785
rect 613 4776 617 4780
rect 623 4776 627 4780
rect 633 4776 637 4780
rect 643 4776 647 4780
rect 613 4771 617 4775
rect 623 4771 627 4775
rect 633 4771 637 4775
rect 643 4771 647 4775
rect 613 4766 617 4770
rect 623 4766 627 4770
rect 633 4766 637 4770
rect 643 4766 647 4770
rect 659 4781 663 4785
rect 669 4781 673 4785
rect 679 4781 683 4785
rect 689 4781 693 4785
rect 659 4776 663 4780
rect 669 4776 673 4780
rect 679 4776 683 4780
rect 689 4776 693 4780
rect 659 4771 663 4775
rect 669 4771 673 4775
rect 679 4771 683 4775
rect 689 4771 693 4775
rect 659 4766 663 4770
rect 669 4766 673 4770
rect 679 4766 683 4770
rect 689 4766 693 4770
rect 613 4752 617 4756
rect 623 4752 627 4756
rect 633 4752 637 4756
rect 643 4752 647 4756
rect 613 4747 617 4751
rect 623 4747 627 4751
rect 633 4747 637 4751
rect 643 4747 647 4751
rect 613 4742 617 4746
rect 623 4742 627 4746
rect 633 4742 637 4746
rect 643 4742 647 4746
rect 613 4737 617 4741
rect 623 4737 627 4741
rect 633 4737 637 4741
rect 643 4737 647 4741
rect 659 4752 663 4756
rect 669 4752 673 4756
rect 679 4752 683 4756
rect 689 4752 693 4756
rect 659 4747 663 4751
rect 669 4747 673 4751
rect 679 4747 683 4751
rect 689 4747 693 4751
rect 659 4742 663 4746
rect 669 4742 673 4746
rect 679 4742 683 4746
rect 689 4742 693 4746
rect 659 4737 663 4741
rect 669 4737 673 4741
rect 679 4737 683 4741
rect 689 4737 693 4741
rect 2412 6885 2416 6889
rect 2545 6118 2549 6122
rect 2544 6015 2548 6019
rect 2412 5903 2416 5907
rect 2801 6518 2805 6522
rect 2545 5136 2549 5140
rect 2544 5033 2548 5037
rect 4496 7471 4500 7475
rect 4501 7471 4505 7475
rect 4496 7466 4500 7470
rect 4501 7466 4505 7470
rect 4496 7461 4500 7465
rect 4501 7461 4505 7465
rect 4496 7456 4500 7460
rect 4501 7456 4505 7460
rect 4496 7451 4500 7455
rect 4501 7451 4505 7455
rect 4496 7446 4500 7450
rect 4501 7446 4505 7450
rect 4496 7441 4500 7445
rect 4501 7441 4505 7445
rect 4496 7436 4500 7440
rect 4501 7436 4505 7440
rect 4496 7431 4500 7435
rect 4501 7431 4505 7435
rect 4496 7426 4500 7430
rect 4501 7426 4505 7430
rect 4496 7421 4500 7425
rect 4501 7421 4505 7425
rect 4496 7416 4500 7420
rect 4501 7416 4505 7420
rect 4496 7411 4500 7415
rect 4501 7411 4505 7415
rect 4553 7311 4557 7315
rect 4558 7311 4562 7315
rect 4553 7306 4557 7310
rect 4558 7306 4562 7310
rect 4553 7301 4557 7305
rect 4558 7301 4562 7305
rect 4553 7296 4557 7300
rect 4558 7296 4562 7300
rect 4496 7289 4500 7293
rect 4501 7289 4505 7293
rect 4496 7284 4500 7288
rect 4501 7284 4505 7288
rect 4496 7279 4500 7283
rect 4501 7279 4505 7283
rect 4496 7274 4500 7278
rect 4501 7274 4505 7278
rect 4496 7269 4500 7273
rect 4501 7269 4505 7273
rect 4496 7264 4500 7268
rect 4501 7264 4505 7268
rect 4496 7259 4500 7263
rect 4501 7259 4505 7263
rect 4496 7254 4500 7258
rect 4501 7254 4505 7258
rect 4496 7249 4500 7253
rect 4501 7249 4505 7253
rect 4553 7291 4557 7295
rect 4558 7291 4562 7295
rect 4553 7286 4557 7290
rect 4558 7286 4562 7290
rect 4553 7281 4557 7285
rect 4558 7281 4562 7285
rect 4553 7276 4557 7280
rect 4558 7276 4562 7280
rect 4553 7271 4557 7275
rect 4558 7271 4562 7275
rect 4553 7266 4557 7270
rect 4558 7266 4562 7270
rect 4553 7261 4557 7265
rect 4558 7261 4562 7265
rect 4553 7256 4557 7260
rect 4558 7256 4562 7260
rect 4553 7251 4557 7255
rect 4558 7251 4562 7255
rect 4496 7244 4500 7248
rect 4501 7244 4505 7248
rect 4496 7239 4500 7243
rect 4501 7239 4505 7243
rect 4479 7230 4483 7234
rect 4489 7230 4493 7234
rect 4499 7230 4503 7234
rect 4509 7230 4513 7234
rect 4479 7225 4483 7229
rect 4489 7225 4493 7229
rect 4499 7225 4503 7229
rect 4509 7225 4513 7229
rect 4479 7220 4483 7224
rect 4489 7220 4493 7224
rect 4499 7220 4503 7224
rect 4509 7220 4513 7224
rect 4479 7215 4483 7219
rect 4489 7215 4493 7219
rect 4499 7215 4503 7219
rect 4509 7215 4513 7219
rect 4525 7230 4529 7234
rect 4535 7230 4539 7234
rect 4545 7230 4549 7234
rect 4555 7230 4559 7234
rect 4525 7225 4529 7229
rect 4535 7225 4539 7229
rect 4545 7225 4549 7229
rect 4555 7225 4559 7229
rect 4525 7220 4529 7224
rect 4535 7220 4539 7224
rect 4545 7220 4549 7224
rect 4555 7220 4559 7224
rect 4525 7215 4529 7219
rect 4535 7215 4539 7219
rect 4545 7215 4549 7219
rect 4555 7215 4559 7219
rect 4479 7202 4483 7206
rect 4489 7202 4493 7206
rect 4499 7202 4503 7206
rect 4509 7202 4513 7206
rect 4479 7197 4483 7201
rect 4489 7197 4493 7201
rect 4499 7197 4503 7201
rect 4509 7197 4513 7201
rect 4479 7192 4483 7196
rect 4489 7192 4493 7196
rect 4499 7192 4503 7196
rect 4509 7192 4513 7196
rect 4479 7187 4483 7191
rect 4489 7187 4493 7191
rect 4499 7187 4503 7191
rect 4509 7187 4513 7191
rect 4525 7202 4529 7206
rect 4535 7202 4539 7206
rect 4545 7202 4549 7206
rect 4555 7202 4559 7206
rect 4525 7197 4529 7201
rect 4535 7197 4539 7201
rect 4545 7197 4549 7201
rect 4555 7197 4559 7201
rect 4525 7192 4529 7196
rect 4535 7192 4539 7196
rect 4545 7192 4549 7196
rect 4555 7192 4559 7196
rect 4525 7187 4529 7191
rect 4535 7187 4539 7191
rect 4545 7187 4549 7191
rect 4555 7187 4559 7191
rect 4479 7152 4483 7156
rect 4489 7152 4493 7156
rect 4499 7152 4503 7156
rect 4509 7152 4513 7156
rect 4525 7152 4529 7156
rect 4535 7152 4539 7156
rect 4545 7152 4549 7156
rect 4555 7152 4559 7156
rect 4479 6858 4483 6862
rect 4489 6858 4493 6862
rect 4499 6858 4503 6862
rect 4509 6858 4513 6862
rect 4479 6853 4483 6857
rect 4489 6853 4493 6857
rect 4499 6853 4503 6857
rect 4509 6853 4513 6857
rect 4479 6848 4483 6852
rect 4489 6848 4493 6852
rect 4499 6848 4503 6852
rect 4509 6848 4513 6852
rect 4479 6843 4483 6847
rect 4489 6843 4493 6847
rect 4499 6843 4503 6847
rect 4509 6843 4513 6847
rect 4525 6858 4529 6862
rect 4535 6858 4539 6862
rect 4545 6858 4549 6862
rect 4555 6858 4559 6862
rect 4525 6853 4529 6857
rect 4535 6853 4539 6857
rect 4545 6853 4549 6857
rect 4555 6853 4559 6857
rect 4525 6848 4529 6852
rect 4535 6848 4539 6852
rect 4545 6848 4549 6852
rect 4555 6848 4559 6852
rect 4525 6843 4529 6847
rect 4535 6843 4539 6847
rect 4545 6843 4549 6847
rect 4555 6843 4559 6847
rect 4479 6549 4483 6553
rect 4489 6549 4493 6553
rect 4499 6549 4503 6553
rect 4509 6549 4513 6553
rect 4479 6544 4483 6548
rect 4489 6544 4493 6548
rect 4499 6544 4503 6548
rect 4509 6544 4513 6548
rect 4479 6539 4483 6543
rect 4489 6539 4493 6543
rect 4499 6539 4503 6543
rect 4509 6539 4513 6543
rect 4479 6534 4483 6538
rect 4489 6534 4493 6538
rect 4499 6534 4503 6538
rect 4509 6534 4513 6538
rect 4525 6549 4529 6553
rect 4535 6549 4539 6553
rect 4545 6549 4549 6553
rect 4555 6549 4559 6553
rect 4525 6544 4529 6548
rect 4535 6544 4539 6548
rect 4545 6544 4549 6548
rect 4555 6544 4559 6548
rect 4525 6539 4529 6543
rect 4535 6539 4539 6543
rect 4545 6539 4549 6543
rect 4555 6539 4559 6543
rect 4525 6534 4529 6538
rect 4535 6534 4539 6538
rect 4545 6534 4549 6538
rect 4555 6534 4559 6538
rect 4479 6240 4483 6244
rect 4489 6240 4493 6244
rect 4499 6240 4503 6244
rect 4509 6240 4513 6244
rect 4479 6235 4483 6239
rect 4489 6235 4493 6239
rect 4499 6235 4503 6239
rect 4509 6235 4513 6239
rect 4479 6230 4483 6234
rect 4489 6230 4493 6234
rect 4499 6230 4503 6234
rect 4509 6230 4513 6234
rect 4479 6225 4483 6229
rect 4489 6225 4493 6229
rect 4499 6225 4503 6229
rect 4509 6225 4513 6229
rect 4525 6240 4529 6244
rect 4535 6240 4539 6244
rect 4545 6240 4549 6244
rect 4555 6240 4559 6244
rect 4525 6235 4529 6239
rect 4535 6235 4539 6239
rect 4545 6235 4549 6239
rect 4555 6235 4559 6239
rect 4525 6230 4529 6234
rect 4535 6230 4539 6234
rect 4545 6230 4549 6234
rect 4555 6230 4559 6234
rect 4525 6225 4529 6229
rect 4535 6225 4539 6229
rect 4545 6225 4549 6229
rect 4555 6225 4559 6229
rect 4479 5931 4483 5935
rect 4489 5931 4493 5935
rect 4499 5931 4503 5935
rect 4509 5931 4513 5935
rect 4479 5926 4483 5930
rect 4489 5926 4493 5930
rect 4499 5926 4503 5930
rect 4509 5926 4513 5930
rect 4479 5921 4483 5925
rect 4489 5921 4493 5925
rect 4499 5921 4503 5925
rect 4509 5921 4513 5925
rect 4479 5916 4483 5920
rect 4489 5916 4493 5920
rect 4499 5916 4503 5920
rect 4509 5916 4513 5920
rect 4525 5931 4529 5935
rect 4535 5931 4539 5935
rect 4545 5931 4549 5935
rect 4555 5931 4559 5935
rect 4525 5926 4529 5930
rect 4535 5926 4539 5930
rect 4545 5926 4549 5930
rect 4555 5926 4559 5930
rect 4525 5921 4529 5925
rect 4535 5921 4539 5925
rect 4545 5921 4549 5925
rect 4555 5921 4559 5925
rect 4525 5916 4529 5920
rect 4535 5916 4539 5920
rect 4545 5916 4549 5920
rect 4555 5916 4559 5920
rect 4479 5622 4483 5626
rect 4489 5622 4493 5626
rect 4499 5622 4503 5626
rect 4509 5622 4513 5626
rect 4479 5617 4483 5621
rect 4489 5617 4493 5621
rect 4499 5617 4503 5621
rect 4509 5617 4513 5621
rect 4479 5612 4483 5616
rect 4489 5612 4493 5616
rect 4499 5612 4503 5616
rect 4509 5612 4513 5616
rect 4479 5607 4483 5611
rect 4489 5607 4493 5611
rect 4499 5607 4503 5611
rect 4509 5607 4513 5611
rect 4525 5622 4529 5626
rect 4535 5622 4539 5626
rect 4545 5622 4549 5626
rect 4555 5622 4559 5626
rect 4525 5617 4529 5621
rect 4535 5617 4539 5621
rect 4545 5617 4549 5621
rect 4555 5617 4559 5621
rect 4525 5612 4529 5616
rect 4535 5612 4539 5616
rect 4545 5612 4549 5616
rect 4555 5612 4559 5616
rect 4525 5607 4529 5611
rect 4535 5607 4539 5611
rect 4545 5607 4549 5611
rect 4555 5607 4559 5611
rect 4251 5532 4255 5536
rect 4479 5313 4483 5317
rect 4489 5313 4493 5317
rect 4499 5313 4503 5317
rect 4509 5313 4513 5317
rect 4479 5308 4483 5312
rect 4489 5308 4493 5312
rect 4499 5308 4503 5312
rect 4509 5308 4513 5312
rect 4479 5303 4483 5307
rect 4489 5303 4493 5307
rect 4499 5303 4503 5307
rect 4509 5303 4513 5307
rect 4479 5298 4483 5302
rect 4489 5298 4493 5302
rect 4499 5298 4503 5302
rect 4509 5298 4513 5302
rect 4525 5313 4529 5317
rect 4535 5313 4539 5317
rect 4545 5313 4549 5317
rect 4555 5313 4559 5317
rect 4525 5308 4529 5312
rect 4535 5308 4539 5312
rect 4545 5308 4549 5312
rect 4555 5308 4559 5312
rect 4525 5303 4529 5307
rect 4535 5303 4539 5307
rect 4545 5303 4549 5307
rect 4555 5303 4559 5307
rect 4525 5298 4529 5302
rect 4535 5298 4539 5302
rect 4545 5298 4549 5302
rect 4555 5298 4559 5302
rect 4479 5004 4483 5008
rect 4489 5004 4493 5008
rect 4499 5004 4503 5008
rect 4509 5004 4513 5008
rect 4479 4999 4483 5003
rect 4489 4999 4493 5003
rect 4499 4999 4503 5003
rect 4509 4999 4513 5003
rect 4479 4994 4483 4998
rect 4489 4994 4493 4998
rect 4499 4994 4503 4998
rect 4509 4994 4513 4998
rect 4479 4989 4483 4993
rect 4489 4989 4493 4993
rect 4499 4989 4503 4993
rect 4509 4989 4513 4993
rect 4525 5004 4529 5008
rect 4535 5004 4539 5008
rect 4545 5004 4549 5008
rect 4555 5004 4559 5008
rect 4525 4999 4529 5003
rect 4535 4999 4539 5003
rect 4545 4999 4549 5003
rect 4555 4999 4559 5003
rect 4525 4994 4529 4998
rect 4535 4994 4539 4998
rect 4545 4994 4549 4998
rect 4555 4994 4559 4998
rect 4525 4989 4529 4993
rect 4535 4989 4539 4993
rect 4545 4989 4549 4993
rect 4555 4989 4559 4993
rect 4479 4811 4483 4815
rect 4489 4811 4493 4815
rect 4499 4811 4503 4815
rect 4509 4811 4513 4815
rect 4479 4806 4483 4810
rect 4489 4806 4493 4810
rect 4499 4806 4503 4810
rect 4509 4806 4513 4810
rect 4479 4801 4483 4805
rect 4489 4801 4493 4805
rect 4499 4801 4503 4805
rect 4509 4801 4513 4805
rect 4479 4796 4483 4800
rect 4489 4796 4493 4800
rect 4499 4796 4503 4800
rect 4509 4796 4513 4800
rect 4525 4811 4529 4815
rect 4535 4811 4539 4815
rect 4545 4811 4549 4815
rect 4555 4811 4559 4815
rect 4525 4806 4529 4810
rect 4535 4806 4539 4810
rect 4545 4806 4549 4810
rect 4555 4806 4559 4810
rect 4525 4801 4529 4805
rect 4535 4801 4539 4805
rect 4545 4801 4549 4805
rect 4555 4801 4559 4805
rect 4525 4796 4529 4800
rect 4535 4796 4539 4800
rect 4545 4796 4549 4800
rect 4555 4796 4559 4800
rect 4479 4785 4483 4789
rect 4489 4785 4493 4789
rect 4499 4785 4503 4789
rect 4509 4785 4513 4789
rect 4479 4780 4483 4784
rect 4489 4780 4493 4784
rect 4499 4780 4503 4784
rect 4509 4780 4513 4784
rect 4479 4775 4483 4779
rect 4489 4775 4493 4779
rect 4499 4775 4503 4779
rect 4509 4775 4513 4779
rect 4479 4770 4483 4774
rect 4489 4770 4493 4774
rect 4499 4770 4503 4774
rect 4509 4770 4513 4774
rect 4525 4785 4529 4789
rect 4535 4785 4539 4789
rect 4545 4785 4549 4789
rect 4555 4785 4559 4789
rect 4525 4780 4529 4784
rect 4535 4780 4539 4784
rect 4545 4780 4549 4784
rect 4555 4780 4559 4784
rect 4525 4775 4529 4779
rect 4535 4775 4539 4779
rect 4545 4775 4549 4779
rect 4555 4775 4559 4779
rect 4525 4770 4529 4774
rect 4535 4770 4539 4774
rect 4545 4770 4549 4774
rect 4555 4770 4559 4774
rect 4479 4759 4483 4763
rect 4489 4759 4493 4763
rect 4499 4759 4503 4763
rect 4509 4759 4513 4763
rect 4479 4754 4483 4758
rect 4489 4754 4493 4758
rect 4499 4754 4503 4758
rect 4509 4754 4513 4758
rect 4479 4749 4483 4753
rect 4489 4749 4493 4753
rect 4499 4749 4503 4753
rect 4509 4749 4513 4753
rect 4479 4744 4483 4748
rect 4489 4744 4493 4748
rect 4499 4744 4503 4748
rect 4509 4744 4513 4748
rect 4525 4759 4529 4763
rect 4535 4759 4539 4763
rect 4545 4759 4549 4763
rect 4555 4759 4559 4763
rect 4525 4754 4529 4758
rect 4535 4754 4539 4758
rect 4545 4754 4549 4758
rect 4555 4754 4559 4758
rect 4525 4749 4529 4753
rect 4535 4749 4539 4753
rect 4545 4749 4549 4753
rect 4555 4749 4559 4753
rect 4525 4744 4529 4748
rect 4535 4744 4539 4748
rect 4545 4744 4549 4748
rect 4555 4744 4559 4748
rect 4479 4733 4483 4737
rect 4489 4733 4493 4737
rect 4499 4733 4503 4737
rect 4509 4733 4513 4737
rect 4479 4728 4483 4732
rect 4489 4728 4493 4732
rect 4499 4728 4503 4732
rect 4509 4728 4513 4732
rect 4479 4723 4483 4727
rect 4489 4723 4493 4727
rect 4499 4723 4503 4727
rect 4509 4723 4513 4727
rect 2910 4691 2914 4695
rect 4479 4718 4483 4722
rect 4489 4718 4493 4722
rect 4499 4718 4503 4722
rect 4509 4718 4513 4722
rect 4525 4733 4529 4737
rect 4535 4733 4539 4737
rect 4545 4733 4549 4737
rect 4555 4733 4559 4737
rect 4525 4728 4529 4732
rect 4535 4728 4539 4732
rect 4545 4728 4549 4732
rect 4555 4728 4559 4732
rect 4525 4723 4529 4727
rect 4535 4723 4539 4727
rect 4545 4723 4549 4727
rect 4555 4723 4559 4727
rect 4525 4718 4529 4722
rect 4535 4718 4539 4722
rect 4545 4718 4549 4722
rect 4555 4718 4559 4722
rect 4479 4707 4483 4711
rect 4489 4707 4493 4711
rect 4499 4707 4503 4711
rect 4509 4707 4513 4711
rect 4479 4702 4483 4706
rect 4489 4702 4493 4706
rect 4499 4702 4503 4706
rect 4509 4702 4513 4706
rect 4479 4697 4483 4701
rect 4489 4697 4493 4701
rect 4499 4697 4503 4701
rect 4509 4697 4513 4701
rect 4479 4692 4483 4696
rect 4489 4692 4493 4696
rect 4499 4692 4503 4696
rect 4509 4692 4513 4696
rect 4525 4707 4529 4711
rect 4535 4707 4539 4711
rect 4545 4707 4549 4711
rect 4555 4707 4559 4711
rect 4525 4702 4529 4706
rect 4535 4702 4539 4706
rect 4545 4702 4549 4706
rect 4555 4702 4559 4706
rect 4525 4697 4529 4701
rect 4535 4697 4539 4701
rect 4545 4697 4549 4701
rect 4555 4697 4559 4701
rect 4525 4692 4529 4696
rect 4535 4692 4539 4696
rect 4545 4692 4549 4696
rect 4555 4692 4559 4696
rect 1820 4649 1824 4653
rect 1825 4649 1829 4653
rect 1820 4644 1824 4648
rect 1825 4644 1829 4648
rect 1820 4639 1824 4643
rect 1825 4639 1829 4643
rect 1820 4634 1824 4638
rect 1825 4634 1829 4638
rect 1820 4629 1824 4633
rect 1825 4629 1829 4633
rect 757 4624 761 4628
rect 762 4624 766 4628
rect 767 4624 771 4628
rect 772 4624 776 4628
rect 757 4614 761 4618
rect 762 4614 766 4618
rect 767 4614 771 4618
rect 772 4614 776 4618
rect 757 4604 761 4608
rect 762 4604 766 4608
rect 767 4604 771 4608
rect 772 4604 776 4608
rect 757 4594 761 4598
rect 762 4594 766 4598
rect 767 4594 771 4598
rect 772 4594 776 4598
rect 783 4624 787 4628
rect 788 4624 792 4628
rect 793 4624 797 4628
rect 798 4624 802 4628
rect 783 4614 787 4618
rect 788 4614 792 4618
rect 793 4614 797 4618
rect 798 4614 802 4618
rect 783 4604 787 4608
rect 788 4604 792 4608
rect 793 4604 797 4608
rect 798 4604 802 4608
rect 783 4594 787 4598
rect 788 4594 792 4598
rect 793 4594 797 4598
rect 798 4594 802 4598
rect 809 4624 813 4628
rect 814 4624 818 4628
rect 819 4624 823 4628
rect 824 4624 828 4628
rect 809 4614 813 4618
rect 814 4614 818 4618
rect 819 4614 823 4618
rect 824 4614 828 4618
rect 809 4604 813 4608
rect 814 4604 818 4608
rect 819 4604 823 4608
rect 824 4604 828 4608
rect 809 4594 813 4598
rect 814 4594 818 4598
rect 819 4594 823 4598
rect 824 4594 828 4598
rect 835 4624 839 4628
rect 840 4624 844 4628
rect 845 4624 849 4628
rect 850 4624 854 4628
rect 835 4614 839 4618
rect 840 4614 844 4618
rect 845 4614 849 4618
rect 850 4614 854 4618
rect 835 4604 839 4608
rect 840 4604 844 4608
rect 845 4604 849 4608
rect 850 4604 854 4608
rect 835 4594 839 4598
rect 840 4594 844 4598
rect 845 4594 849 4598
rect 850 4594 854 4598
rect 861 4624 865 4628
rect 866 4624 870 4628
rect 871 4624 875 4628
rect 876 4624 880 4628
rect 861 4614 865 4618
rect 866 4614 870 4618
rect 871 4614 875 4618
rect 876 4614 880 4618
rect 861 4604 865 4608
rect 866 4604 870 4608
rect 871 4604 875 4608
rect 876 4604 880 4608
rect 861 4594 865 4598
rect 866 4594 870 4598
rect 871 4594 875 4598
rect 876 4594 880 4598
rect 1053 4624 1057 4628
rect 1058 4624 1062 4628
rect 1063 4624 1067 4628
rect 1068 4624 1072 4628
rect 1053 4614 1057 4618
rect 1058 4614 1062 4618
rect 1063 4614 1067 4618
rect 1068 4614 1072 4618
rect 1362 4624 1366 4628
rect 1367 4624 1371 4628
rect 1372 4624 1376 4628
rect 1377 4624 1381 4628
rect 1362 4614 1366 4618
rect 1367 4614 1371 4618
rect 1372 4614 1376 4618
rect 1377 4614 1381 4618
rect 1671 4624 1675 4628
rect 1676 4624 1680 4628
rect 1681 4624 1685 4628
rect 1686 4624 1690 4628
rect 1671 4614 1675 4618
rect 1676 4614 1680 4618
rect 1681 4614 1685 4618
rect 1686 4614 1690 4618
rect 1053 4604 1057 4608
rect 1058 4604 1062 4608
rect 1063 4604 1067 4608
rect 1068 4604 1072 4608
rect 1053 4594 1057 4598
rect 1058 4594 1062 4598
rect 1063 4594 1067 4598
rect 1068 4594 1072 4598
rect 1077 4607 1081 4611
rect 1082 4607 1086 4611
rect 1087 4607 1091 4611
rect 1092 4607 1096 4611
rect 1097 4607 1101 4611
rect 1102 4607 1106 4611
rect 1107 4607 1111 4611
rect 1112 4607 1116 4611
rect 1117 4607 1121 4611
rect 1122 4607 1126 4611
rect 1127 4607 1131 4611
rect 1077 4602 1081 4606
rect 1082 4602 1086 4606
rect 1087 4602 1091 4606
rect 1092 4602 1096 4606
rect 1097 4602 1101 4606
rect 1102 4602 1106 4606
rect 1107 4602 1111 4606
rect 1112 4602 1116 4606
rect 1117 4602 1121 4606
rect 1122 4602 1126 4606
rect 1127 4602 1131 4606
rect 1249 4607 1253 4611
rect 1254 4607 1258 4611
rect 1259 4607 1263 4611
rect 1264 4607 1268 4611
rect 1269 4607 1273 4611
rect 1274 4607 1278 4611
rect 1279 4607 1283 4611
rect 1284 4607 1288 4611
rect 1289 4607 1293 4611
rect 1294 4607 1298 4611
rect 1299 4607 1303 4611
rect 1304 4607 1308 4611
rect 1309 4607 1313 4611
rect 1249 4602 1253 4606
rect 1254 4602 1258 4606
rect 1259 4602 1263 4606
rect 1264 4602 1268 4606
rect 1269 4602 1273 4606
rect 1274 4602 1278 4606
rect 1279 4602 1283 4606
rect 1284 4602 1288 4606
rect 1289 4602 1293 4606
rect 1294 4602 1298 4606
rect 1299 4602 1303 4606
rect 1304 4602 1308 4606
rect 1309 4602 1313 4606
rect 757 4578 761 4582
rect 762 4578 766 4582
rect 767 4578 771 4582
rect 772 4578 776 4582
rect 757 4568 761 4572
rect 762 4568 766 4572
rect 767 4568 771 4572
rect 772 4568 776 4572
rect 757 4558 761 4562
rect 762 4558 766 4562
rect 767 4558 771 4562
rect 772 4558 776 4562
rect 757 4548 761 4552
rect 762 4548 766 4552
rect 767 4548 771 4552
rect 772 4548 776 4552
rect 783 4578 787 4582
rect 788 4578 792 4582
rect 793 4578 797 4582
rect 798 4578 802 4582
rect 783 4568 787 4572
rect 788 4568 792 4572
rect 793 4568 797 4572
rect 798 4568 802 4572
rect 783 4558 787 4562
rect 788 4558 792 4562
rect 793 4558 797 4562
rect 798 4558 802 4562
rect 783 4548 787 4552
rect 788 4548 792 4552
rect 793 4548 797 4552
rect 798 4548 802 4552
rect 809 4578 813 4582
rect 814 4578 818 4582
rect 819 4578 823 4582
rect 824 4578 828 4582
rect 809 4568 813 4572
rect 814 4568 818 4572
rect 819 4568 823 4572
rect 824 4568 828 4572
rect 809 4558 813 4562
rect 814 4558 818 4562
rect 819 4558 823 4562
rect 824 4558 828 4562
rect 809 4548 813 4552
rect 814 4548 818 4552
rect 819 4548 823 4552
rect 824 4548 828 4552
rect 835 4578 839 4582
rect 840 4578 844 4582
rect 845 4578 849 4582
rect 850 4578 854 4582
rect 835 4568 839 4572
rect 840 4568 844 4572
rect 845 4568 849 4572
rect 850 4568 854 4572
rect 835 4558 839 4562
rect 840 4558 844 4562
rect 845 4558 849 4562
rect 850 4558 854 4562
rect 835 4548 839 4552
rect 840 4548 844 4552
rect 845 4548 849 4552
rect 850 4548 854 4552
rect 861 4578 865 4582
rect 866 4578 870 4582
rect 871 4578 875 4582
rect 876 4578 880 4582
rect 861 4568 865 4572
rect 866 4568 870 4572
rect 871 4568 875 4572
rect 876 4568 880 4572
rect 861 4558 865 4562
rect 866 4558 870 4562
rect 871 4558 875 4562
rect 876 4558 880 4562
rect 861 4548 865 4552
rect 866 4548 870 4552
rect 871 4548 875 4552
rect 876 4548 880 4552
rect 1053 4578 1057 4582
rect 1058 4578 1062 4582
rect 1063 4578 1067 4582
rect 1068 4578 1072 4582
rect 1053 4568 1057 4572
rect 1058 4568 1062 4572
rect 1063 4568 1067 4572
rect 1068 4568 1072 4572
rect 1053 4558 1057 4562
rect 1058 4558 1062 4562
rect 1063 4558 1067 4562
rect 1068 4558 1072 4562
rect 1053 4548 1057 4552
rect 1058 4548 1062 4552
rect 1063 4548 1067 4552
rect 1068 4548 1072 4552
rect 1089 4550 1093 4554
rect 1094 4550 1098 4554
rect 1099 4550 1103 4554
rect 1104 4550 1108 4554
rect 1109 4550 1113 4554
rect 1114 4550 1118 4554
rect 1119 4550 1123 4554
rect 1124 4550 1128 4554
rect 1129 4550 1133 4554
rect 1134 4550 1138 4554
rect 1139 4550 1143 4554
rect 1144 4550 1148 4554
rect 1149 4550 1153 4554
rect 1089 4545 1093 4549
rect 1094 4545 1098 4549
rect 1099 4545 1103 4549
rect 1104 4545 1108 4549
rect 1109 4545 1113 4549
rect 1114 4545 1118 4549
rect 1119 4545 1123 4549
rect 1124 4545 1128 4549
rect 1129 4545 1133 4549
rect 1134 4545 1138 4549
rect 1139 4545 1143 4549
rect 1144 4545 1148 4549
rect 1149 4545 1153 4549
rect 1362 4604 1366 4608
rect 1367 4604 1371 4608
rect 1372 4604 1376 4608
rect 1377 4604 1381 4608
rect 1362 4594 1366 4598
rect 1367 4594 1371 4598
rect 1372 4594 1376 4598
rect 1377 4594 1381 4598
rect 1386 4607 1390 4611
rect 1391 4607 1395 4611
rect 1396 4607 1400 4611
rect 1401 4607 1405 4611
rect 1406 4607 1410 4611
rect 1411 4607 1415 4611
rect 1416 4607 1420 4611
rect 1421 4607 1425 4611
rect 1426 4607 1430 4611
rect 1431 4607 1435 4611
rect 1436 4607 1440 4611
rect 1386 4602 1390 4606
rect 1391 4602 1395 4606
rect 1396 4602 1400 4606
rect 1401 4602 1405 4606
rect 1406 4602 1410 4606
rect 1411 4602 1415 4606
rect 1416 4602 1420 4606
rect 1421 4602 1425 4606
rect 1426 4602 1430 4606
rect 1431 4602 1435 4606
rect 1436 4602 1440 4606
rect 1558 4607 1562 4611
rect 1563 4607 1567 4611
rect 1568 4607 1572 4611
rect 1573 4607 1577 4611
rect 1578 4607 1582 4611
rect 1583 4607 1587 4611
rect 1588 4607 1592 4611
rect 1593 4607 1597 4611
rect 1598 4607 1602 4611
rect 1603 4607 1607 4611
rect 1608 4607 1612 4611
rect 1613 4607 1617 4611
rect 1618 4607 1622 4611
rect 1558 4602 1562 4606
rect 1563 4602 1567 4606
rect 1568 4602 1572 4606
rect 1573 4602 1577 4606
rect 1578 4602 1582 4606
rect 1583 4602 1587 4606
rect 1588 4602 1592 4606
rect 1593 4602 1597 4606
rect 1598 4602 1602 4606
rect 1603 4602 1607 4606
rect 1608 4602 1612 4606
rect 1613 4602 1617 4606
rect 1618 4602 1622 4606
rect 1337 4574 1341 4578
rect 1342 4574 1346 4578
rect 1337 4569 1341 4573
rect 1342 4569 1346 4573
rect 1337 4564 1341 4568
rect 1342 4564 1346 4568
rect 1337 4559 1341 4563
rect 1342 4559 1346 4563
rect 1337 4554 1341 4558
rect 1342 4554 1346 4558
rect 1337 4549 1341 4553
rect 1342 4549 1346 4553
rect 1362 4578 1366 4582
rect 1367 4578 1371 4582
rect 1372 4578 1376 4582
rect 1377 4578 1381 4582
rect 1362 4568 1366 4572
rect 1367 4568 1371 4572
rect 1372 4568 1376 4572
rect 1377 4568 1381 4572
rect 1362 4558 1366 4562
rect 1367 4558 1371 4562
rect 1372 4558 1376 4562
rect 1377 4558 1381 4562
rect 1511 4569 1515 4573
rect 1516 4569 1520 4573
rect 1511 4564 1515 4568
rect 1516 4564 1520 4568
rect 1511 4559 1515 4563
rect 1516 4559 1520 4563
rect 1362 4548 1366 4552
rect 1367 4548 1371 4552
rect 1372 4548 1376 4552
rect 1377 4548 1381 4552
rect 1398 4550 1402 4554
rect 1403 4550 1407 4554
rect 1408 4550 1412 4554
rect 1413 4550 1417 4554
rect 1418 4550 1422 4554
rect 1423 4550 1427 4554
rect 1428 4550 1432 4554
rect 1433 4550 1437 4554
rect 1438 4550 1442 4554
rect 1443 4550 1447 4554
rect 1448 4550 1452 4554
rect 1453 4550 1457 4554
rect 1458 4550 1462 4554
rect 1337 4544 1341 4548
rect 1342 4544 1346 4548
rect 1337 4539 1341 4543
rect 1342 4539 1346 4543
rect 1337 4534 1341 4538
rect 1342 4534 1346 4538
rect 1337 4529 1341 4533
rect 1342 4529 1346 4533
rect 1337 4524 1341 4528
rect 1342 4524 1346 4528
rect 1337 4519 1341 4523
rect 1342 4519 1346 4523
rect 1337 4514 1341 4518
rect 1342 4514 1346 4518
rect 1398 4545 1402 4549
rect 1403 4545 1407 4549
rect 1408 4545 1412 4549
rect 1413 4545 1417 4549
rect 1418 4545 1422 4549
rect 1423 4545 1427 4549
rect 1428 4545 1432 4549
rect 1433 4545 1437 4549
rect 1438 4545 1442 4549
rect 1443 4545 1447 4549
rect 1448 4545 1452 4549
rect 1453 4545 1457 4549
rect 1458 4545 1462 4549
rect 1511 4554 1515 4558
rect 1516 4554 1520 4558
rect 1511 4549 1515 4553
rect 1516 4549 1520 4553
rect 1511 4544 1515 4548
rect 1516 4544 1520 4548
rect 1511 4539 1515 4543
rect 1516 4539 1520 4543
rect 1511 4534 1515 4538
rect 1516 4534 1520 4538
rect 1511 4529 1515 4533
rect 1516 4529 1520 4533
rect 1511 4524 1515 4528
rect 1516 4524 1520 4528
rect 1511 4519 1515 4523
rect 1516 4519 1520 4523
rect 1820 4624 1824 4628
rect 1825 4624 1829 4628
rect 1820 4619 1824 4623
rect 1825 4619 1829 4623
rect 1820 4614 1824 4618
rect 1825 4614 1829 4618
rect 1980 4624 1984 4628
rect 1985 4624 1989 4628
rect 1990 4624 1994 4628
rect 1995 4624 1999 4628
rect 1980 4614 1984 4618
rect 1985 4614 1989 4618
rect 1990 4614 1994 4618
rect 1995 4614 1999 4618
rect 2289 4624 2293 4628
rect 2294 4624 2298 4628
rect 2299 4624 2303 4628
rect 2304 4624 2308 4628
rect 2289 4614 2293 4618
rect 2294 4614 2298 4618
rect 2299 4614 2303 4618
rect 2304 4614 2308 4618
rect 2598 4624 2602 4628
rect 2603 4624 2607 4628
rect 2608 4624 2612 4628
rect 2613 4624 2617 4628
rect 2598 4614 2602 4618
rect 2603 4614 2607 4618
rect 2608 4614 2612 4618
rect 2613 4614 2617 4618
rect 2907 4624 2911 4628
rect 2912 4624 2916 4628
rect 2917 4624 2921 4628
rect 2922 4624 2926 4628
rect 2907 4614 2911 4618
rect 2912 4614 2916 4618
rect 2917 4614 2921 4618
rect 2922 4614 2926 4618
rect 1671 4604 1675 4608
rect 1676 4604 1680 4608
rect 1681 4604 1685 4608
rect 1686 4604 1690 4608
rect 1671 4594 1675 4598
rect 1676 4594 1680 4598
rect 1681 4594 1685 4598
rect 1686 4594 1690 4598
rect 1695 4607 1699 4611
rect 1700 4607 1704 4611
rect 1705 4607 1709 4611
rect 1710 4607 1714 4611
rect 1715 4607 1719 4611
rect 1720 4607 1724 4611
rect 1725 4607 1729 4611
rect 1730 4607 1734 4611
rect 1735 4607 1739 4611
rect 1740 4607 1744 4611
rect 1745 4607 1749 4611
rect 1695 4602 1699 4606
rect 1700 4602 1704 4606
rect 1705 4602 1709 4606
rect 1710 4602 1714 4606
rect 1715 4602 1719 4606
rect 1720 4602 1724 4606
rect 1725 4602 1729 4606
rect 1730 4602 1734 4606
rect 1735 4602 1739 4606
rect 1740 4602 1744 4606
rect 1745 4602 1749 4606
rect 1820 4609 1824 4613
rect 1825 4609 1829 4613
rect 1820 4604 1824 4608
rect 1825 4604 1829 4608
rect 1820 4599 1824 4603
rect 1825 4599 1829 4603
rect 1867 4607 1871 4611
rect 1872 4607 1876 4611
rect 1877 4607 1881 4611
rect 1882 4607 1886 4611
rect 1887 4607 1891 4611
rect 1892 4607 1896 4611
rect 1897 4607 1901 4611
rect 1902 4607 1906 4611
rect 1907 4607 1911 4611
rect 1912 4607 1916 4611
rect 1917 4607 1921 4611
rect 1922 4607 1926 4611
rect 1927 4607 1931 4611
rect 1867 4602 1871 4606
rect 1872 4602 1876 4606
rect 1877 4602 1881 4606
rect 1882 4602 1886 4606
rect 1887 4602 1891 4606
rect 1892 4602 1896 4606
rect 1897 4602 1901 4606
rect 1902 4602 1906 4606
rect 1907 4602 1911 4606
rect 1912 4602 1916 4606
rect 1917 4602 1921 4606
rect 1922 4602 1926 4606
rect 1927 4602 1931 4606
rect 1646 4574 1650 4578
rect 1651 4574 1655 4578
rect 1646 4569 1650 4573
rect 1651 4569 1655 4573
rect 1646 4564 1650 4568
rect 1651 4564 1655 4568
rect 1646 4559 1650 4563
rect 1651 4559 1655 4563
rect 1646 4554 1650 4558
rect 1651 4554 1655 4558
rect 1646 4549 1650 4553
rect 1651 4549 1655 4553
rect 1671 4578 1675 4582
rect 1676 4578 1680 4582
rect 1681 4578 1685 4582
rect 1686 4578 1690 4582
rect 1671 4568 1675 4572
rect 1676 4568 1680 4572
rect 1681 4568 1685 4572
rect 1686 4568 1690 4572
rect 1671 4558 1675 4562
rect 1676 4558 1680 4562
rect 1681 4558 1685 4562
rect 1686 4558 1690 4562
rect 1671 4548 1675 4552
rect 1676 4548 1680 4552
rect 1681 4548 1685 4552
rect 1686 4548 1690 4552
rect 1707 4550 1711 4554
rect 1712 4550 1716 4554
rect 1717 4550 1721 4554
rect 1722 4550 1726 4554
rect 1727 4550 1731 4554
rect 1732 4550 1736 4554
rect 1737 4550 1741 4554
rect 1742 4550 1746 4554
rect 1747 4550 1751 4554
rect 1752 4550 1756 4554
rect 1757 4550 1761 4554
rect 1762 4550 1766 4554
rect 1767 4550 1771 4554
rect 1646 4544 1650 4548
rect 1651 4544 1655 4548
rect 1646 4539 1650 4543
rect 1651 4539 1655 4543
rect 1646 4534 1650 4538
rect 1651 4534 1655 4538
rect 1646 4529 1650 4533
rect 1651 4529 1655 4533
rect 1646 4524 1650 4528
rect 1651 4524 1655 4528
rect 1646 4519 1650 4523
rect 1651 4519 1655 4523
rect 1646 4514 1650 4518
rect 1651 4514 1655 4518
rect 1707 4545 1711 4549
rect 1712 4545 1716 4549
rect 1717 4545 1721 4549
rect 1722 4545 1726 4549
rect 1727 4545 1731 4549
rect 1732 4545 1736 4549
rect 1737 4545 1741 4549
rect 1742 4545 1746 4549
rect 1747 4545 1751 4549
rect 1752 4545 1756 4549
rect 1757 4545 1761 4549
rect 1762 4545 1766 4549
rect 1767 4545 1771 4549
rect 1980 4604 1984 4608
rect 1985 4604 1989 4608
rect 1990 4604 1994 4608
rect 1995 4604 1999 4608
rect 1980 4594 1984 4598
rect 1985 4594 1989 4598
rect 1990 4594 1994 4598
rect 1995 4594 1999 4598
rect 2004 4607 2008 4611
rect 2009 4607 2013 4611
rect 2014 4607 2018 4611
rect 2019 4607 2023 4611
rect 2024 4607 2028 4611
rect 2029 4607 2033 4611
rect 2034 4607 2038 4611
rect 2039 4607 2043 4611
rect 2044 4607 2048 4611
rect 2049 4607 2053 4611
rect 2054 4607 2058 4611
rect 2004 4602 2008 4606
rect 2009 4602 2013 4606
rect 2014 4602 2018 4606
rect 2019 4602 2023 4606
rect 2024 4602 2028 4606
rect 2029 4602 2033 4606
rect 2034 4602 2038 4606
rect 2039 4602 2043 4606
rect 2044 4602 2048 4606
rect 2049 4602 2053 4606
rect 2054 4602 2058 4606
rect 2176 4607 2180 4611
rect 2181 4607 2185 4611
rect 2186 4607 2190 4611
rect 2191 4607 2195 4611
rect 2196 4607 2200 4611
rect 2201 4607 2205 4611
rect 2206 4607 2210 4611
rect 2211 4607 2215 4611
rect 2216 4607 2220 4611
rect 2221 4607 2225 4611
rect 2226 4607 2230 4611
rect 2231 4607 2235 4611
rect 2236 4607 2240 4611
rect 2176 4602 2180 4606
rect 2181 4602 2185 4606
rect 2186 4602 2190 4606
rect 2191 4602 2195 4606
rect 2196 4602 2200 4606
rect 2201 4602 2205 4606
rect 2206 4602 2210 4606
rect 2211 4602 2215 4606
rect 2216 4602 2220 4606
rect 2221 4602 2225 4606
rect 2226 4602 2230 4606
rect 2231 4602 2235 4606
rect 2236 4602 2240 4606
rect 1955 4574 1959 4578
rect 1960 4574 1964 4578
rect 1955 4569 1959 4573
rect 1960 4569 1964 4573
rect 1955 4564 1959 4568
rect 1960 4564 1964 4568
rect 1955 4559 1959 4563
rect 1960 4559 1964 4563
rect 1955 4554 1959 4558
rect 1960 4554 1964 4558
rect 1955 4549 1959 4553
rect 1960 4549 1964 4553
rect 1980 4578 1984 4582
rect 1985 4578 1989 4582
rect 1990 4578 1994 4582
rect 1995 4578 1999 4582
rect 1980 4568 1984 4572
rect 1985 4568 1989 4572
rect 1990 4568 1994 4572
rect 1995 4568 1999 4572
rect 1980 4558 1984 4562
rect 1985 4558 1989 4562
rect 1990 4558 1994 4562
rect 1995 4558 1999 4562
rect 1980 4548 1984 4552
rect 1985 4548 1989 4552
rect 1990 4548 1994 4552
rect 1995 4548 1999 4552
rect 2016 4550 2020 4554
rect 2021 4550 2025 4554
rect 2026 4550 2030 4554
rect 2031 4550 2035 4554
rect 2036 4550 2040 4554
rect 2041 4550 2045 4554
rect 2046 4550 2050 4554
rect 2051 4550 2055 4554
rect 2056 4550 2060 4554
rect 2061 4550 2065 4554
rect 2066 4550 2070 4554
rect 2071 4550 2075 4554
rect 2076 4550 2080 4554
rect 1955 4544 1959 4548
rect 1960 4544 1964 4548
rect 1955 4539 1959 4543
rect 1960 4539 1964 4543
rect 1955 4534 1959 4538
rect 1960 4534 1964 4538
rect 1955 4529 1959 4533
rect 1960 4529 1964 4533
rect 1955 4524 1959 4528
rect 1960 4524 1964 4528
rect 1955 4519 1959 4523
rect 1960 4519 1964 4523
rect 1955 4514 1959 4518
rect 1960 4514 1964 4518
rect 2016 4545 2020 4549
rect 2021 4545 2025 4549
rect 2026 4545 2030 4549
rect 2031 4545 2035 4549
rect 2036 4545 2040 4549
rect 2041 4545 2045 4549
rect 2046 4545 2050 4549
rect 2051 4545 2055 4549
rect 2056 4545 2060 4549
rect 2061 4545 2065 4549
rect 2066 4545 2070 4549
rect 2071 4545 2075 4549
rect 2076 4545 2080 4549
rect 2289 4604 2293 4608
rect 2294 4604 2298 4608
rect 2299 4604 2303 4608
rect 2304 4604 2308 4608
rect 2289 4594 2293 4598
rect 2294 4594 2298 4598
rect 2299 4594 2303 4598
rect 2304 4594 2308 4598
rect 2313 4607 2317 4611
rect 2318 4607 2322 4611
rect 2323 4607 2327 4611
rect 2328 4607 2332 4611
rect 2333 4607 2337 4611
rect 2338 4607 2342 4611
rect 2343 4607 2347 4611
rect 2348 4607 2352 4611
rect 2353 4607 2357 4611
rect 2358 4607 2362 4611
rect 2363 4607 2367 4611
rect 2313 4602 2317 4606
rect 2318 4602 2322 4606
rect 2323 4602 2327 4606
rect 2328 4602 2332 4606
rect 2333 4602 2337 4606
rect 2338 4602 2342 4606
rect 2343 4602 2347 4606
rect 2348 4602 2352 4606
rect 2353 4602 2357 4606
rect 2358 4602 2362 4606
rect 2363 4602 2367 4606
rect 2485 4607 2489 4611
rect 2490 4607 2494 4611
rect 2495 4607 2499 4611
rect 2500 4607 2504 4611
rect 2505 4607 2509 4611
rect 2510 4607 2514 4611
rect 2515 4607 2519 4611
rect 2520 4607 2524 4611
rect 2525 4607 2529 4611
rect 2530 4607 2534 4611
rect 2535 4607 2539 4611
rect 2540 4607 2544 4611
rect 2545 4607 2549 4611
rect 2485 4602 2489 4606
rect 2490 4602 2494 4606
rect 2495 4602 2499 4606
rect 2500 4602 2504 4606
rect 2505 4602 2509 4606
rect 2510 4602 2514 4606
rect 2515 4602 2519 4606
rect 2520 4602 2524 4606
rect 2525 4602 2529 4606
rect 2530 4602 2534 4606
rect 2535 4602 2539 4606
rect 2540 4602 2544 4606
rect 2545 4602 2549 4606
rect 2264 4574 2268 4578
rect 2269 4574 2273 4578
rect 2264 4569 2268 4573
rect 2269 4569 2273 4573
rect 2264 4564 2268 4568
rect 2269 4564 2273 4568
rect 2264 4559 2268 4563
rect 2269 4559 2273 4563
rect 2264 4554 2268 4558
rect 2269 4554 2273 4558
rect 2264 4549 2268 4553
rect 2269 4549 2273 4553
rect 2289 4578 2293 4582
rect 2294 4578 2298 4582
rect 2299 4578 2303 4582
rect 2304 4578 2308 4582
rect 2289 4568 2293 4572
rect 2294 4568 2298 4572
rect 2299 4568 2303 4572
rect 2304 4568 2308 4572
rect 2289 4558 2293 4562
rect 2294 4558 2298 4562
rect 2299 4558 2303 4562
rect 2304 4558 2308 4562
rect 2289 4548 2293 4552
rect 2294 4548 2298 4552
rect 2299 4548 2303 4552
rect 2304 4548 2308 4552
rect 2325 4550 2329 4554
rect 2330 4550 2334 4554
rect 2335 4550 2339 4554
rect 2340 4550 2344 4554
rect 2345 4550 2349 4554
rect 2350 4550 2354 4554
rect 2355 4550 2359 4554
rect 2360 4550 2364 4554
rect 2365 4550 2369 4554
rect 2370 4550 2374 4554
rect 2375 4550 2379 4554
rect 2380 4550 2384 4554
rect 2385 4550 2389 4554
rect 2264 4544 2268 4548
rect 2269 4544 2273 4548
rect 2264 4539 2268 4543
rect 2269 4539 2273 4543
rect 2264 4534 2268 4538
rect 2269 4534 2273 4538
rect 2264 4529 2268 4533
rect 2269 4529 2273 4533
rect 2264 4524 2268 4528
rect 2269 4524 2273 4528
rect 2264 4519 2268 4523
rect 2269 4519 2273 4523
rect 2264 4514 2268 4518
rect 2269 4514 2273 4518
rect 2325 4545 2329 4549
rect 2330 4545 2334 4549
rect 2335 4545 2339 4549
rect 2340 4545 2344 4549
rect 2345 4545 2349 4549
rect 2350 4545 2354 4549
rect 2355 4545 2359 4549
rect 2360 4545 2364 4549
rect 2365 4545 2369 4549
rect 2370 4545 2374 4549
rect 2375 4545 2379 4549
rect 2380 4545 2384 4549
rect 2385 4545 2389 4549
rect 2598 4604 2602 4608
rect 2603 4604 2607 4608
rect 2608 4604 2612 4608
rect 2613 4604 2617 4608
rect 2598 4594 2602 4598
rect 2603 4594 2607 4598
rect 2608 4594 2612 4598
rect 2613 4594 2617 4598
rect 2622 4607 2626 4611
rect 2627 4607 2631 4611
rect 2632 4607 2636 4611
rect 2637 4607 2641 4611
rect 2642 4607 2646 4611
rect 2647 4607 2651 4611
rect 2652 4607 2656 4611
rect 2657 4607 2661 4611
rect 2662 4607 2666 4611
rect 2667 4607 2671 4611
rect 2672 4607 2676 4611
rect 2622 4602 2626 4606
rect 2627 4602 2631 4606
rect 2632 4602 2636 4606
rect 2637 4602 2641 4606
rect 2642 4602 2646 4606
rect 2647 4602 2651 4606
rect 2652 4602 2656 4606
rect 2657 4602 2661 4606
rect 2662 4602 2666 4606
rect 2667 4602 2671 4606
rect 2672 4602 2676 4606
rect 2794 4607 2798 4611
rect 2799 4607 2803 4611
rect 2804 4607 2808 4611
rect 2809 4607 2813 4611
rect 2814 4607 2818 4611
rect 2819 4607 2823 4611
rect 2824 4607 2828 4611
rect 2829 4607 2833 4611
rect 2834 4607 2838 4611
rect 2839 4607 2843 4611
rect 2844 4607 2848 4611
rect 2849 4607 2853 4611
rect 2854 4607 2858 4611
rect 2794 4602 2798 4606
rect 2799 4602 2803 4606
rect 2804 4602 2808 4606
rect 2809 4602 2813 4606
rect 2814 4602 2818 4606
rect 2819 4602 2823 4606
rect 2824 4602 2828 4606
rect 2829 4602 2833 4606
rect 2834 4602 2838 4606
rect 2839 4602 2843 4606
rect 2844 4602 2848 4606
rect 2849 4602 2853 4606
rect 2854 4602 2858 4606
rect 2573 4574 2577 4578
rect 2578 4574 2582 4578
rect 2573 4569 2577 4573
rect 2578 4569 2582 4573
rect 2573 4564 2577 4568
rect 2578 4564 2582 4568
rect 2573 4559 2577 4563
rect 2578 4559 2582 4563
rect 2573 4554 2577 4558
rect 2578 4554 2582 4558
rect 2573 4549 2577 4553
rect 2578 4549 2582 4553
rect 2598 4578 2602 4582
rect 2603 4578 2607 4582
rect 2608 4578 2612 4582
rect 2613 4578 2617 4582
rect 2598 4568 2602 4572
rect 2603 4568 2607 4572
rect 2608 4568 2612 4572
rect 2613 4568 2617 4572
rect 2598 4558 2602 4562
rect 2603 4558 2607 4562
rect 2608 4558 2612 4562
rect 2613 4558 2617 4562
rect 2598 4548 2602 4552
rect 2603 4548 2607 4552
rect 2608 4548 2612 4552
rect 2613 4548 2617 4552
rect 2634 4550 2638 4554
rect 2639 4550 2643 4554
rect 2644 4550 2648 4554
rect 2649 4550 2653 4554
rect 2654 4550 2658 4554
rect 2659 4550 2663 4554
rect 2664 4550 2668 4554
rect 2669 4550 2673 4554
rect 2674 4550 2678 4554
rect 2679 4550 2683 4554
rect 2684 4550 2688 4554
rect 2689 4550 2693 4554
rect 2694 4550 2698 4554
rect 2573 4544 2577 4548
rect 2578 4544 2582 4548
rect 2573 4539 2577 4543
rect 2578 4539 2582 4543
rect 2573 4534 2577 4538
rect 2578 4534 2582 4538
rect 2573 4529 2577 4533
rect 2578 4529 2582 4533
rect 2573 4524 2577 4528
rect 2578 4524 2582 4528
rect 2573 4519 2577 4523
rect 2578 4519 2582 4523
rect 2573 4514 2577 4518
rect 2578 4514 2582 4518
rect 2634 4545 2638 4549
rect 2639 4545 2643 4549
rect 2644 4545 2648 4549
rect 2649 4545 2653 4549
rect 2654 4545 2658 4549
rect 2659 4545 2663 4549
rect 2664 4545 2668 4549
rect 2669 4545 2673 4549
rect 2674 4545 2678 4549
rect 2679 4545 2683 4549
rect 2684 4545 2688 4549
rect 2689 4545 2693 4549
rect 2694 4545 2698 4549
rect 2907 4604 2911 4608
rect 2912 4604 2916 4608
rect 2917 4604 2921 4608
rect 2922 4604 2926 4608
rect 2907 4594 2911 4598
rect 2912 4594 2916 4598
rect 2917 4594 2921 4598
rect 2922 4594 2926 4598
rect 2931 4607 2935 4611
rect 2936 4607 2940 4611
rect 2941 4607 2945 4611
rect 2946 4607 2950 4611
rect 2951 4607 2955 4611
rect 2956 4607 2960 4611
rect 2961 4607 2965 4611
rect 2966 4607 2970 4611
rect 2971 4607 2975 4611
rect 2976 4607 2980 4611
rect 2981 4607 2985 4611
rect 2931 4602 2935 4606
rect 2936 4602 2940 4606
rect 2941 4602 2945 4606
rect 2946 4602 2950 4606
rect 2951 4602 2955 4606
rect 2956 4602 2960 4606
rect 2961 4602 2965 4606
rect 2966 4602 2970 4606
rect 2971 4602 2975 4606
rect 2976 4602 2980 4606
rect 2981 4602 2985 4606
rect 2882 4574 2886 4578
rect 2887 4574 2891 4578
rect 2882 4569 2886 4573
rect 2887 4569 2891 4573
rect 2882 4564 2886 4568
rect 2887 4564 2891 4568
rect 2882 4559 2886 4563
rect 2887 4559 2891 4563
rect 2882 4554 2886 4558
rect 2887 4554 2891 4558
rect 2882 4549 2886 4553
rect 2887 4549 2891 4553
rect 2907 4578 2911 4582
rect 2912 4578 2916 4582
rect 2917 4578 2921 4582
rect 2922 4578 2926 4582
rect 2907 4568 2911 4572
rect 2912 4568 2916 4572
rect 2917 4568 2921 4572
rect 2922 4568 2926 4572
rect 3674 4649 3678 4653
rect 3679 4649 3683 4653
rect 3674 4644 3678 4648
rect 3679 4644 3683 4648
rect 3674 4639 3678 4643
rect 3679 4639 3683 4643
rect 3674 4634 3678 4638
rect 3679 4634 3683 4638
rect 3674 4629 3678 4633
rect 3679 4629 3683 4633
rect 3216 4624 3220 4628
rect 3221 4624 3225 4628
rect 3226 4624 3230 4628
rect 3231 4624 3235 4628
rect 3216 4614 3220 4618
rect 3221 4614 3225 4618
rect 3226 4614 3230 4618
rect 3231 4614 3235 4618
rect 3525 4624 3529 4628
rect 3530 4624 3534 4628
rect 3535 4624 3539 4628
rect 3540 4624 3544 4628
rect 3525 4614 3529 4618
rect 3530 4614 3534 4618
rect 3535 4614 3539 4618
rect 3540 4614 3544 4618
rect 3000 4573 3005 4578
rect 3103 4607 3107 4611
rect 3108 4607 3112 4611
rect 3113 4607 3117 4611
rect 3118 4607 3122 4611
rect 3123 4607 3127 4611
rect 3128 4607 3132 4611
rect 3133 4607 3137 4611
rect 3138 4607 3142 4611
rect 3143 4607 3147 4611
rect 3148 4607 3152 4611
rect 3153 4607 3157 4611
rect 3158 4607 3162 4611
rect 3163 4607 3167 4611
rect 3103 4602 3107 4606
rect 3108 4602 3112 4606
rect 3113 4602 3117 4606
rect 3118 4602 3122 4606
rect 3123 4602 3127 4606
rect 3128 4602 3132 4606
rect 3133 4602 3137 4606
rect 3138 4602 3142 4606
rect 3143 4602 3147 4606
rect 3148 4602 3152 4606
rect 3153 4602 3157 4606
rect 3158 4602 3162 4606
rect 3163 4602 3167 4606
rect 2907 4558 2911 4562
rect 2912 4558 2916 4562
rect 2917 4558 2921 4562
rect 2922 4558 2926 4562
rect 2907 4548 2911 4552
rect 2912 4548 2916 4552
rect 2917 4548 2921 4552
rect 2922 4548 2926 4552
rect 2943 4550 2947 4554
rect 2948 4550 2952 4554
rect 2953 4550 2957 4554
rect 2958 4550 2962 4554
rect 2963 4550 2967 4554
rect 2968 4550 2972 4554
rect 2973 4550 2977 4554
rect 2978 4550 2982 4554
rect 2983 4550 2987 4554
rect 2988 4550 2992 4554
rect 2993 4550 2997 4554
rect 2998 4550 3002 4554
rect 3003 4550 3007 4554
rect 2882 4544 2886 4548
rect 2887 4544 2891 4548
rect 2882 4539 2886 4543
rect 2887 4539 2891 4543
rect 2882 4534 2886 4538
rect 2887 4534 2891 4538
rect 2882 4529 2886 4533
rect 2887 4529 2891 4533
rect 2882 4524 2886 4528
rect 2887 4524 2891 4528
rect 2882 4519 2886 4523
rect 2887 4519 2891 4523
rect 2882 4514 2886 4518
rect 2887 4514 2891 4518
rect 2943 4545 2947 4549
rect 2948 4545 2952 4549
rect 2953 4545 2957 4549
rect 2958 4545 2962 4549
rect 2963 4545 2967 4549
rect 2968 4545 2972 4549
rect 2973 4545 2977 4549
rect 2978 4545 2982 4549
rect 2983 4545 2987 4549
rect 2988 4545 2992 4549
rect 2993 4545 2997 4549
rect 2998 4545 3002 4549
rect 3003 4545 3007 4549
rect 3216 4604 3220 4608
rect 3221 4604 3225 4608
rect 3226 4604 3230 4608
rect 3231 4604 3235 4608
rect 3216 4594 3220 4598
rect 3221 4594 3225 4598
rect 3226 4594 3230 4598
rect 3231 4594 3235 4598
rect 3240 4607 3244 4611
rect 3245 4607 3249 4611
rect 3250 4607 3254 4611
rect 3255 4607 3259 4611
rect 3260 4607 3264 4611
rect 3265 4607 3269 4611
rect 3270 4607 3274 4611
rect 3275 4607 3279 4611
rect 3280 4607 3284 4611
rect 3285 4607 3289 4611
rect 3290 4607 3294 4611
rect 3240 4602 3244 4606
rect 3245 4602 3249 4606
rect 3250 4602 3254 4606
rect 3255 4602 3259 4606
rect 3260 4602 3264 4606
rect 3265 4602 3269 4606
rect 3270 4602 3274 4606
rect 3275 4602 3279 4606
rect 3280 4602 3284 4606
rect 3285 4602 3289 4606
rect 3290 4602 3294 4606
rect 3412 4607 3416 4611
rect 3417 4607 3421 4611
rect 3422 4607 3426 4611
rect 3427 4607 3431 4611
rect 3432 4607 3436 4611
rect 3437 4607 3441 4611
rect 3442 4607 3446 4611
rect 3447 4607 3451 4611
rect 3452 4607 3456 4611
rect 3457 4607 3461 4611
rect 3462 4607 3466 4611
rect 3467 4607 3471 4611
rect 3472 4607 3476 4611
rect 3412 4602 3416 4606
rect 3417 4602 3421 4606
rect 3422 4602 3426 4606
rect 3427 4602 3431 4606
rect 3432 4602 3436 4606
rect 3437 4602 3441 4606
rect 3442 4602 3446 4606
rect 3447 4602 3451 4606
rect 3452 4602 3456 4606
rect 3457 4602 3461 4606
rect 3462 4602 3466 4606
rect 3467 4602 3471 4606
rect 3472 4602 3476 4606
rect 3191 4574 3195 4578
rect 3196 4574 3200 4578
rect 3191 4569 3195 4573
rect 3196 4569 3200 4573
rect 3191 4564 3195 4568
rect 3196 4564 3200 4568
rect 3191 4559 3195 4563
rect 3196 4559 3200 4563
rect 3191 4554 3195 4558
rect 3196 4554 3200 4558
rect 3191 4549 3195 4553
rect 3196 4549 3200 4553
rect 3216 4578 3220 4582
rect 3221 4578 3225 4582
rect 3226 4578 3230 4582
rect 3231 4578 3235 4582
rect 3216 4568 3220 4572
rect 3221 4568 3225 4572
rect 3226 4568 3230 4572
rect 3231 4568 3235 4572
rect 3216 4558 3220 4562
rect 3221 4558 3225 4562
rect 3226 4558 3230 4562
rect 3231 4558 3235 4562
rect 3216 4548 3220 4552
rect 3221 4548 3225 4552
rect 3226 4548 3230 4552
rect 3231 4548 3235 4552
rect 3252 4550 3256 4554
rect 3257 4550 3261 4554
rect 3262 4550 3266 4554
rect 3267 4550 3271 4554
rect 3272 4550 3276 4554
rect 3277 4550 3281 4554
rect 3282 4550 3286 4554
rect 3287 4550 3291 4554
rect 3292 4550 3296 4554
rect 3297 4550 3301 4554
rect 3302 4550 3306 4554
rect 3307 4550 3311 4554
rect 3312 4550 3316 4554
rect 3191 4544 3195 4548
rect 3196 4544 3200 4548
rect 3191 4539 3195 4543
rect 3196 4539 3200 4543
rect 3191 4534 3195 4538
rect 3196 4534 3200 4538
rect 3191 4529 3195 4533
rect 3196 4529 3200 4533
rect 3191 4524 3195 4528
rect 3196 4524 3200 4528
rect 3191 4519 3195 4523
rect 3196 4519 3200 4523
rect 3191 4514 3195 4518
rect 3196 4514 3200 4518
rect 3252 4545 3256 4549
rect 3257 4545 3261 4549
rect 3262 4545 3266 4549
rect 3267 4545 3271 4549
rect 3272 4545 3276 4549
rect 3277 4545 3281 4549
rect 3282 4545 3286 4549
rect 3287 4545 3291 4549
rect 3292 4545 3296 4549
rect 3297 4545 3301 4549
rect 3302 4545 3306 4549
rect 3307 4545 3311 4549
rect 3312 4545 3316 4549
rect 3674 4624 3678 4628
rect 3679 4624 3683 4628
rect 3674 4619 3678 4623
rect 3679 4619 3683 4623
rect 3674 4614 3678 4618
rect 3679 4614 3683 4618
rect 3834 4624 3838 4628
rect 3839 4624 3843 4628
rect 3844 4624 3848 4628
rect 3849 4624 3853 4628
rect 3834 4614 3838 4618
rect 3839 4614 3843 4618
rect 3844 4614 3848 4618
rect 3849 4614 3853 4618
rect 3525 4604 3529 4608
rect 3530 4604 3534 4608
rect 3535 4604 3539 4608
rect 3540 4604 3544 4608
rect 3525 4594 3529 4598
rect 3530 4594 3534 4598
rect 3535 4594 3539 4598
rect 3540 4594 3544 4598
rect 3549 4607 3553 4611
rect 3554 4607 3558 4611
rect 3559 4607 3563 4611
rect 3564 4607 3568 4611
rect 3569 4607 3573 4611
rect 3574 4607 3578 4611
rect 3579 4607 3583 4611
rect 3584 4607 3588 4611
rect 3589 4607 3593 4611
rect 3594 4607 3598 4611
rect 3599 4607 3603 4611
rect 3549 4602 3553 4606
rect 3554 4602 3558 4606
rect 3559 4602 3563 4606
rect 3564 4602 3568 4606
rect 3569 4602 3573 4606
rect 3574 4602 3578 4606
rect 3579 4602 3583 4606
rect 3584 4602 3588 4606
rect 3589 4602 3593 4606
rect 3594 4602 3598 4606
rect 3599 4602 3603 4606
rect 3674 4609 3678 4613
rect 3679 4609 3683 4613
rect 3674 4604 3678 4608
rect 3679 4604 3683 4608
rect 3674 4599 3678 4603
rect 3679 4599 3683 4603
rect 3721 4607 3725 4611
rect 3726 4607 3730 4611
rect 3731 4607 3735 4611
rect 3736 4607 3740 4611
rect 3741 4607 3745 4611
rect 3746 4607 3750 4611
rect 3751 4607 3755 4611
rect 3756 4607 3760 4611
rect 3761 4607 3765 4611
rect 3766 4607 3770 4611
rect 3771 4607 3775 4611
rect 3776 4607 3780 4611
rect 3781 4607 3785 4611
rect 3721 4602 3725 4606
rect 3726 4602 3730 4606
rect 3731 4602 3735 4606
rect 3736 4602 3740 4606
rect 3741 4602 3745 4606
rect 3746 4602 3750 4606
rect 3751 4602 3755 4606
rect 3756 4602 3760 4606
rect 3761 4602 3765 4606
rect 3766 4602 3770 4606
rect 3771 4602 3775 4606
rect 3776 4602 3780 4606
rect 3781 4602 3785 4606
rect 3500 4574 3504 4578
rect 3505 4574 3509 4578
rect 3500 4569 3504 4573
rect 3505 4569 3509 4573
rect 3500 4564 3504 4568
rect 3505 4564 3509 4568
rect 3500 4559 3504 4563
rect 3505 4559 3509 4563
rect 3500 4554 3504 4558
rect 3505 4554 3509 4558
rect 3500 4549 3504 4553
rect 3505 4549 3509 4553
rect 3525 4578 3529 4582
rect 3530 4578 3534 4582
rect 3535 4578 3539 4582
rect 3540 4578 3544 4582
rect 3525 4568 3529 4572
rect 3530 4568 3534 4572
rect 3535 4568 3539 4572
rect 3540 4568 3544 4572
rect 3525 4558 3529 4562
rect 3530 4558 3534 4562
rect 3535 4558 3539 4562
rect 3540 4558 3544 4562
rect 3525 4548 3529 4552
rect 3530 4548 3534 4552
rect 3535 4548 3539 4552
rect 3540 4548 3544 4552
rect 3561 4550 3565 4554
rect 3566 4550 3570 4554
rect 3571 4550 3575 4554
rect 3576 4550 3580 4554
rect 3581 4550 3585 4554
rect 3586 4550 3590 4554
rect 3591 4550 3595 4554
rect 3596 4550 3600 4554
rect 3601 4550 3605 4554
rect 3606 4550 3610 4554
rect 3611 4550 3615 4554
rect 3616 4550 3620 4554
rect 3621 4550 3625 4554
rect 3500 4544 3504 4548
rect 3505 4544 3509 4548
rect 3500 4539 3504 4543
rect 3505 4539 3509 4543
rect 3500 4534 3504 4538
rect 3505 4534 3509 4538
rect 3500 4529 3504 4533
rect 3505 4529 3509 4533
rect 3500 4524 3504 4528
rect 3505 4524 3509 4528
rect 3500 4519 3504 4523
rect 3505 4519 3509 4523
rect 3500 4514 3504 4518
rect 3505 4514 3509 4518
rect 3561 4545 3565 4549
rect 3566 4545 3570 4549
rect 3571 4545 3575 4549
rect 3576 4545 3580 4549
rect 3581 4545 3585 4549
rect 3586 4545 3590 4549
rect 3591 4545 3595 4549
rect 3596 4545 3600 4549
rect 3601 4545 3605 4549
rect 3606 4545 3610 4549
rect 3611 4545 3615 4549
rect 3616 4545 3620 4549
rect 3621 4545 3625 4549
rect 3834 4604 3838 4608
rect 3839 4604 3843 4608
rect 3844 4604 3848 4608
rect 3849 4604 3853 4608
rect 3834 4594 3838 4598
rect 3839 4594 3843 4598
rect 3844 4594 3848 4598
rect 3849 4594 3853 4598
rect 4235 4624 4239 4628
rect 4240 4624 4244 4628
rect 4245 4624 4249 4628
rect 4250 4624 4254 4628
rect 4235 4614 4239 4618
rect 4240 4614 4244 4618
rect 4245 4614 4249 4618
rect 4250 4614 4254 4618
rect 4235 4604 4239 4608
rect 4240 4604 4244 4608
rect 4245 4604 4249 4608
rect 4250 4604 4254 4608
rect 4235 4594 4239 4598
rect 4240 4594 4244 4598
rect 4245 4594 4249 4598
rect 4250 4594 4254 4598
rect 4264 4624 4268 4628
rect 4269 4624 4273 4628
rect 4274 4624 4278 4628
rect 4279 4624 4283 4628
rect 4264 4614 4268 4618
rect 4269 4614 4273 4618
rect 4274 4614 4278 4618
rect 4279 4614 4283 4618
rect 4264 4604 4268 4608
rect 4269 4604 4273 4608
rect 4274 4604 4278 4608
rect 4279 4604 4283 4608
rect 4264 4594 4268 4598
rect 4269 4594 4273 4598
rect 4274 4594 4278 4598
rect 4279 4594 4283 4598
rect 4293 4624 4297 4628
rect 4298 4624 4302 4628
rect 4303 4624 4307 4628
rect 4308 4624 4312 4628
rect 4293 4614 4297 4618
rect 4298 4614 4302 4618
rect 4303 4614 4307 4618
rect 4308 4614 4312 4618
rect 4293 4604 4297 4608
rect 4298 4604 4302 4608
rect 4303 4604 4307 4608
rect 4308 4604 4312 4608
rect 4293 4594 4297 4598
rect 4298 4594 4302 4598
rect 4303 4594 4307 4598
rect 4308 4594 4312 4598
rect 4322 4624 4326 4628
rect 4327 4624 4331 4628
rect 4332 4624 4336 4628
rect 4337 4624 4341 4628
rect 4322 4614 4326 4618
rect 4327 4614 4331 4618
rect 4332 4614 4336 4618
rect 4337 4614 4341 4618
rect 4322 4604 4326 4608
rect 4327 4604 4331 4608
rect 4332 4604 4336 4608
rect 4337 4604 4341 4608
rect 4322 4594 4326 4598
rect 4327 4594 4331 4598
rect 4332 4594 4336 4598
rect 4337 4594 4341 4598
rect 4351 4624 4355 4628
rect 4356 4624 4360 4628
rect 4361 4624 4365 4628
rect 4366 4624 4370 4628
rect 4351 4614 4355 4618
rect 4356 4614 4360 4618
rect 4361 4614 4365 4618
rect 4366 4614 4370 4618
rect 4351 4604 4355 4608
rect 4356 4604 4360 4608
rect 4361 4604 4365 4608
rect 4366 4604 4370 4608
rect 4351 4594 4355 4598
rect 4356 4594 4360 4598
rect 4361 4594 4365 4598
rect 4366 4594 4370 4598
rect 3809 4574 3813 4578
rect 3814 4574 3818 4578
rect 3809 4569 3813 4573
rect 3814 4569 3818 4573
rect 3809 4564 3813 4568
rect 3814 4564 3818 4568
rect 3809 4559 3813 4563
rect 3814 4559 3818 4563
rect 3809 4554 3813 4558
rect 3814 4554 3818 4558
rect 3809 4549 3813 4553
rect 3814 4549 3818 4553
rect 3834 4578 3838 4582
rect 3839 4578 3843 4582
rect 3844 4578 3848 4582
rect 3849 4578 3853 4582
rect 3834 4568 3838 4572
rect 3839 4568 3843 4572
rect 3844 4568 3848 4572
rect 3849 4568 3853 4572
rect 3834 4558 3838 4562
rect 3839 4558 3843 4562
rect 3844 4558 3848 4562
rect 3849 4558 3853 4562
rect 3834 4548 3838 4552
rect 3839 4548 3843 4552
rect 3844 4548 3848 4552
rect 3849 4548 3853 4552
rect 4235 4578 4239 4582
rect 4240 4578 4244 4582
rect 4245 4578 4249 4582
rect 4250 4578 4254 4582
rect 4235 4568 4239 4572
rect 4240 4568 4244 4572
rect 4245 4568 4249 4572
rect 4250 4568 4254 4572
rect 4235 4558 4239 4562
rect 4240 4558 4244 4562
rect 4245 4558 4249 4562
rect 4250 4558 4254 4562
rect 4235 4548 4239 4552
rect 4240 4548 4244 4552
rect 4245 4548 4249 4552
rect 4250 4548 4254 4552
rect 4264 4578 4268 4582
rect 4269 4578 4273 4582
rect 4274 4578 4278 4582
rect 4279 4578 4283 4582
rect 4264 4568 4268 4572
rect 4269 4568 4273 4572
rect 4274 4568 4278 4572
rect 4279 4568 4283 4572
rect 4264 4558 4268 4562
rect 4269 4558 4273 4562
rect 4274 4558 4278 4562
rect 4279 4558 4283 4562
rect 4264 4548 4268 4552
rect 4269 4548 4273 4552
rect 4274 4548 4278 4552
rect 4279 4548 4283 4552
rect 4293 4578 4297 4582
rect 4298 4578 4302 4582
rect 4303 4578 4307 4582
rect 4308 4578 4312 4582
rect 4293 4568 4297 4572
rect 4298 4568 4302 4572
rect 4303 4568 4307 4572
rect 4308 4568 4312 4572
rect 4293 4558 4297 4562
rect 4298 4558 4302 4562
rect 4303 4558 4307 4562
rect 4308 4558 4312 4562
rect 4293 4548 4297 4552
rect 4298 4548 4302 4552
rect 4303 4548 4307 4552
rect 4308 4548 4312 4552
rect 4322 4578 4326 4582
rect 4327 4578 4331 4582
rect 4332 4578 4336 4582
rect 4337 4578 4341 4582
rect 4322 4568 4326 4572
rect 4327 4568 4331 4572
rect 4332 4568 4336 4572
rect 4337 4568 4341 4572
rect 4322 4558 4326 4562
rect 4327 4558 4331 4562
rect 4332 4558 4336 4562
rect 4337 4558 4341 4562
rect 4322 4548 4326 4552
rect 4327 4548 4331 4552
rect 4332 4548 4336 4552
rect 4337 4548 4341 4552
rect 4351 4578 4355 4582
rect 4356 4578 4360 4582
rect 4361 4578 4365 4582
rect 4366 4578 4370 4582
rect 4351 4568 4355 4572
rect 4356 4568 4360 4572
rect 4361 4568 4365 4572
rect 4366 4568 4370 4572
rect 4351 4558 4355 4562
rect 4356 4558 4360 4562
rect 4361 4558 4365 4562
rect 4366 4558 4370 4562
rect 4351 4548 4355 4552
rect 4356 4548 4360 4552
rect 4361 4548 4365 4552
rect 4366 4548 4370 4552
rect 3809 4544 3813 4548
rect 3814 4544 3818 4548
rect 3809 4539 3813 4543
rect 3814 4539 3818 4543
rect 3809 4534 3813 4538
rect 3814 4534 3818 4538
rect 3809 4529 3813 4533
rect 3814 4529 3818 4533
rect 3809 4524 3813 4528
rect 3814 4524 3818 4528
rect 3809 4519 3813 4523
rect 3814 4519 3818 4523
rect 3809 4514 3813 4518
rect 3814 4514 3818 4518
<< metal3 >>
rect 570 9800 4602 9809
rect 570 9796 1354 9800
rect 1358 9796 1359 9800
rect 1363 9796 1663 9800
rect 1667 9796 1668 9800
rect 1672 9796 1972 9800
rect 1976 9796 1977 9800
rect 1981 9796 2281 9800
rect 2285 9796 2286 9800
rect 2290 9796 2590 9800
rect 2594 9796 2595 9800
rect 2599 9796 2899 9800
rect 2903 9796 2904 9800
rect 2908 9796 3208 9800
rect 3212 9796 3213 9800
rect 3217 9796 3517 9800
rect 3521 9796 3522 9800
rect 3526 9796 3826 9800
rect 3830 9796 3831 9800
rect 3835 9796 4602 9800
rect 570 9795 4602 9796
rect 570 9791 1354 9795
rect 1358 9791 1359 9795
rect 1363 9791 1663 9795
rect 1667 9791 1668 9795
rect 1672 9791 1972 9795
rect 1976 9791 1977 9795
rect 1981 9791 2281 9795
rect 2285 9791 2286 9795
rect 2290 9791 2590 9795
rect 2594 9791 2595 9795
rect 2599 9791 2899 9795
rect 2903 9791 2904 9795
rect 2908 9791 3208 9795
rect 3212 9791 3213 9795
rect 3217 9791 3517 9795
rect 3521 9791 3522 9795
rect 3526 9791 3652 9795
rect 3656 9791 3657 9795
rect 3661 9791 3826 9795
rect 3830 9791 3831 9795
rect 3835 9791 4602 9795
rect 570 9790 4602 9791
rect 570 9786 1354 9790
rect 1358 9786 1359 9790
rect 1363 9786 1663 9790
rect 1667 9786 1668 9790
rect 1672 9786 1972 9790
rect 1976 9786 1977 9790
rect 1981 9786 2281 9790
rect 2285 9786 2286 9790
rect 2290 9786 2590 9790
rect 2594 9786 2595 9790
rect 2599 9786 2899 9790
rect 2903 9786 2904 9790
rect 2908 9786 3208 9790
rect 3212 9786 3213 9790
rect 3217 9786 3517 9790
rect 3521 9786 3522 9790
rect 3526 9786 3652 9790
rect 3656 9786 3657 9790
rect 3661 9786 3826 9790
rect 3830 9786 3831 9790
rect 3835 9786 4602 9790
rect 570 9785 4602 9786
rect 570 9781 1354 9785
rect 1358 9781 1359 9785
rect 1363 9781 1663 9785
rect 1667 9781 1668 9785
rect 1672 9781 1972 9785
rect 1976 9781 1977 9785
rect 1981 9781 2281 9785
rect 2285 9781 2286 9785
rect 2290 9781 2590 9785
rect 2594 9781 2595 9785
rect 2599 9781 2899 9785
rect 2903 9781 2904 9785
rect 2908 9781 3208 9785
rect 3212 9781 3213 9785
rect 3217 9781 3517 9785
rect 3521 9781 3522 9785
rect 3526 9781 3652 9785
rect 3656 9781 3657 9785
rect 3661 9781 3826 9785
rect 3830 9781 3831 9785
rect 3835 9781 4602 9785
rect 570 9780 4602 9781
rect 570 9776 1354 9780
rect 1358 9776 1359 9780
rect 1363 9776 1663 9780
rect 1667 9776 1668 9780
rect 1672 9776 1972 9780
rect 1976 9776 1977 9780
rect 1981 9776 2281 9780
rect 2285 9776 2286 9780
rect 2290 9776 2590 9780
rect 2594 9776 2595 9780
rect 2599 9776 2899 9780
rect 2903 9776 2904 9780
rect 2908 9776 3208 9780
rect 3212 9776 3213 9780
rect 3217 9776 3517 9780
rect 3521 9776 3522 9780
rect 3526 9776 3652 9780
rect 3656 9776 3657 9780
rect 3661 9776 3826 9780
rect 3830 9776 3831 9780
rect 3835 9776 4602 9780
rect 570 9775 4602 9776
rect 570 9771 1354 9775
rect 1358 9771 1359 9775
rect 1363 9771 1663 9775
rect 1667 9771 1668 9775
rect 1672 9771 1972 9775
rect 1976 9771 1977 9775
rect 1981 9771 2281 9775
rect 2285 9771 2286 9775
rect 2290 9771 2590 9775
rect 2594 9771 2595 9775
rect 2599 9771 2899 9775
rect 2903 9771 2904 9775
rect 2908 9771 3208 9775
rect 3212 9771 3213 9775
rect 3217 9771 3517 9775
rect 3521 9771 3522 9775
rect 3526 9771 3652 9775
rect 3656 9771 3657 9775
rect 3661 9771 3826 9775
rect 3830 9771 3831 9775
rect 3835 9771 4602 9775
rect 570 9770 4602 9771
rect 570 9766 1354 9770
rect 1358 9766 1359 9770
rect 1363 9769 1663 9770
rect 1363 9766 1547 9769
rect 570 9762 802 9766
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 821 9762 831 9766
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 850 9762 860 9766
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 879 9762 889 9766
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 908 9762 918 9766
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 937 9762 1319 9766
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1338 9765 1547 9766
rect 1551 9765 1552 9769
rect 1556 9765 1557 9769
rect 1561 9765 1562 9769
rect 1566 9765 1567 9769
rect 1571 9765 1572 9769
rect 1576 9765 1577 9769
rect 1581 9765 1582 9769
rect 1586 9765 1587 9769
rect 1591 9765 1592 9769
rect 1596 9765 1597 9769
rect 1601 9765 1602 9769
rect 1606 9765 1607 9769
rect 1611 9766 1663 9769
rect 1667 9766 1668 9770
rect 1672 9769 1972 9770
rect 1672 9766 1856 9769
rect 1611 9765 1628 9766
rect 1338 9762 1354 9765
rect 570 9761 1354 9762
rect 1358 9761 1359 9765
rect 1363 9764 1628 9765
rect 1363 9761 1547 9764
rect 570 9760 1547 9761
rect 1551 9760 1552 9764
rect 1556 9760 1557 9764
rect 1561 9760 1562 9764
rect 1566 9760 1567 9764
rect 1571 9760 1572 9764
rect 1576 9760 1577 9764
rect 1581 9760 1582 9764
rect 1586 9760 1587 9764
rect 1591 9760 1592 9764
rect 1596 9760 1597 9764
rect 1601 9760 1602 9764
rect 1606 9760 1607 9764
rect 1611 9762 1628 9764
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1647 9765 1856 9766
rect 1860 9765 1861 9769
rect 1865 9765 1866 9769
rect 1870 9765 1871 9769
rect 1875 9765 1876 9769
rect 1880 9765 1881 9769
rect 1885 9765 1886 9769
rect 1890 9765 1891 9769
rect 1895 9765 1896 9769
rect 1900 9765 1901 9769
rect 1905 9765 1906 9769
rect 1910 9765 1911 9769
rect 1915 9765 1916 9769
rect 1920 9766 1972 9769
rect 1976 9766 1977 9770
rect 1981 9769 2281 9770
rect 1981 9766 2165 9769
rect 1920 9765 1937 9766
rect 1647 9762 1663 9765
rect 1611 9761 1663 9762
rect 1667 9761 1668 9765
rect 1672 9764 1937 9765
rect 1672 9761 1856 9764
rect 1611 9760 1856 9761
rect 1860 9760 1861 9764
rect 1865 9760 1866 9764
rect 1870 9760 1871 9764
rect 1875 9760 1876 9764
rect 1880 9760 1881 9764
rect 1885 9760 1886 9764
rect 1890 9760 1891 9764
rect 1895 9760 1896 9764
rect 1900 9760 1901 9764
rect 1905 9760 1906 9764
rect 1910 9760 1911 9764
rect 1915 9760 1916 9764
rect 1920 9762 1937 9764
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1956 9765 2165 9766
rect 2169 9765 2170 9769
rect 2174 9765 2175 9769
rect 2179 9765 2180 9769
rect 2184 9765 2185 9769
rect 2189 9765 2190 9769
rect 2194 9765 2195 9769
rect 2199 9765 2200 9769
rect 2204 9765 2205 9769
rect 2209 9765 2210 9769
rect 2214 9765 2215 9769
rect 2219 9765 2220 9769
rect 2224 9765 2225 9769
rect 2229 9766 2281 9769
rect 2285 9766 2286 9770
rect 2290 9769 2590 9770
rect 2290 9766 2474 9769
rect 2229 9765 2246 9766
rect 1956 9762 1972 9765
rect 1920 9761 1972 9762
rect 1976 9761 1977 9765
rect 1981 9764 2246 9765
rect 1981 9761 2165 9764
rect 1920 9760 2165 9761
rect 2169 9760 2170 9764
rect 2174 9760 2175 9764
rect 2179 9760 2180 9764
rect 2184 9760 2185 9764
rect 2189 9760 2190 9764
rect 2194 9760 2195 9764
rect 2199 9760 2200 9764
rect 2204 9760 2205 9764
rect 2209 9760 2210 9764
rect 2214 9760 2215 9764
rect 2219 9760 2220 9764
rect 2224 9760 2225 9764
rect 2229 9762 2246 9764
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2265 9765 2474 9766
rect 2478 9765 2479 9769
rect 2483 9765 2484 9769
rect 2488 9765 2489 9769
rect 2493 9765 2494 9769
rect 2498 9765 2499 9769
rect 2503 9765 2504 9769
rect 2508 9765 2509 9769
rect 2513 9765 2514 9769
rect 2518 9765 2519 9769
rect 2523 9765 2524 9769
rect 2528 9765 2529 9769
rect 2533 9765 2534 9769
rect 2538 9766 2590 9769
rect 2594 9766 2595 9770
rect 2599 9769 2899 9770
rect 2599 9766 2783 9769
rect 2538 9765 2555 9766
rect 2265 9762 2281 9765
rect 2229 9761 2281 9762
rect 2285 9761 2286 9765
rect 2290 9764 2555 9765
rect 2290 9761 2474 9764
rect 2229 9760 2474 9761
rect 2478 9760 2479 9764
rect 2483 9760 2484 9764
rect 2488 9760 2489 9764
rect 2493 9760 2494 9764
rect 2498 9760 2499 9764
rect 2503 9760 2504 9764
rect 2508 9760 2509 9764
rect 2513 9760 2514 9764
rect 2518 9760 2519 9764
rect 2523 9760 2524 9764
rect 2528 9760 2529 9764
rect 2533 9760 2534 9764
rect 2538 9762 2555 9764
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2574 9765 2783 9766
rect 2787 9765 2788 9769
rect 2792 9765 2793 9769
rect 2797 9765 2798 9769
rect 2802 9765 2803 9769
rect 2807 9765 2808 9769
rect 2812 9765 2813 9769
rect 2817 9765 2818 9769
rect 2822 9765 2823 9769
rect 2827 9765 2828 9769
rect 2832 9765 2833 9769
rect 2837 9765 2838 9769
rect 2842 9765 2843 9769
rect 2847 9766 2899 9769
rect 2903 9766 2904 9770
rect 2908 9769 3208 9770
rect 2908 9766 3092 9769
rect 2847 9765 2864 9766
rect 2574 9762 2590 9765
rect 2538 9761 2590 9762
rect 2594 9761 2595 9765
rect 2599 9764 2864 9765
rect 2599 9761 2783 9764
rect 2538 9760 2783 9761
rect 2787 9760 2788 9764
rect 2792 9760 2793 9764
rect 2797 9760 2798 9764
rect 2802 9760 2803 9764
rect 2807 9760 2808 9764
rect 2812 9760 2813 9764
rect 2817 9760 2818 9764
rect 2822 9760 2823 9764
rect 2827 9760 2828 9764
rect 2832 9760 2833 9764
rect 2837 9760 2838 9764
rect 2842 9760 2843 9764
rect 2847 9762 2864 9764
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2883 9765 3092 9766
rect 3096 9765 3097 9769
rect 3101 9765 3102 9769
rect 3106 9765 3107 9769
rect 3111 9765 3112 9769
rect 3116 9765 3117 9769
rect 3121 9765 3122 9769
rect 3126 9765 3127 9769
rect 3131 9765 3132 9769
rect 3136 9765 3137 9769
rect 3141 9765 3142 9769
rect 3146 9765 3147 9769
rect 3151 9765 3152 9769
rect 3156 9766 3208 9769
rect 3212 9766 3213 9770
rect 3217 9769 3517 9770
rect 3217 9766 3401 9769
rect 3156 9765 3173 9766
rect 2883 9762 2899 9765
rect 2847 9761 2899 9762
rect 2903 9761 2904 9765
rect 2908 9764 3173 9765
rect 2908 9761 3092 9764
rect 2847 9760 3092 9761
rect 3096 9760 3097 9764
rect 3101 9760 3102 9764
rect 3106 9760 3107 9764
rect 3111 9760 3112 9764
rect 3116 9760 3117 9764
rect 3121 9760 3122 9764
rect 3126 9760 3127 9764
rect 3131 9760 3132 9764
rect 3136 9760 3137 9764
rect 3141 9760 3142 9764
rect 3146 9760 3147 9764
rect 3151 9760 3152 9764
rect 3156 9762 3173 9764
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3192 9765 3401 9766
rect 3405 9765 3406 9769
rect 3410 9765 3411 9769
rect 3415 9765 3416 9769
rect 3420 9765 3421 9769
rect 3425 9765 3426 9769
rect 3430 9765 3431 9769
rect 3435 9765 3436 9769
rect 3440 9765 3441 9769
rect 3445 9765 3446 9769
rect 3450 9765 3451 9769
rect 3455 9765 3456 9769
rect 3460 9765 3461 9769
rect 3465 9766 3517 9769
rect 3521 9766 3522 9770
rect 3526 9766 3652 9770
rect 3656 9766 3657 9770
rect 3661 9769 3826 9770
rect 3661 9766 3710 9769
rect 3465 9765 3482 9766
rect 3192 9762 3208 9765
rect 3156 9761 3208 9762
rect 3212 9761 3213 9765
rect 3217 9764 3482 9765
rect 3217 9761 3401 9764
rect 3156 9760 3401 9761
rect 3405 9760 3406 9764
rect 3410 9760 3411 9764
rect 3415 9760 3416 9764
rect 3420 9760 3421 9764
rect 3425 9760 3426 9764
rect 3430 9760 3431 9764
rect 3435 9760 3436 9764
rect 3440 9760 3441 9764
rect 3445 9760 3446 9764
rect 3450 9760 3451 9764
rect 3455 9760 3456 9764
rect 3460 9760 3461 9764
rect 3465 9762 3482 9764
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3501 9765 3710 9766
rect 3714 9765 3715 9769
rect 3719 9765 3720 9769
rect 3724 9765 3725 9769
rect 3729 9765 3730 9769
rect 3734 9765 3735 9769
rect 3739 9765 3740 9769
rect 3744 9765 3745 9769
rect 3749 9765 3750 9769
rect 3754 9765 3755 9769
rect 3759 9765 3760 9769
rect 3764 9765 3765 9769
rect 3769 9765 3770 9769
rect 3774 9766 3826 9769
rect 3830 9766 3831 9770
rect 3835 9769 4602 9770
rect 3835 9766 4019 9769
rect 3774 9765 3791 9766
rect 3501 9762 3517 9765
rect 3465 9761 3517 9762
rect 3521 9761 3522 9765
rect 3526 9761 3652 9765
rect 3656 9761 3657 9765
rect 3661 9764 3791 9765
rect 3661 9761 3710 9764
rect 3465 9760 3710 9761
rect 3714 9760 3715 9764
rect 3719 9760 3720 9764
rect 3724 9760 3725 9764
rect 3729 9760 3730 9764
rect 3734 9760 3735 9764
rect 3739 9760 3740 9764
rect 3744 9760 3745 9764
rect 3749 9760 3750 9764
rect 3754 9760 3755 9764
rect 3759 9760 3760 9764
rect 3764 9760 3765 9764
rect 3769 9760 3770 9764
rect 3774 9762 3791 9764
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3810 9765 4019 9766
rect 4023 9765 4024 9769
rect 4028 9765 4029 9769
rect 4033 9765 4034 9769
rect 4038 9765 4039 9769
rect 4043 9765 4044 9769
rect 4048 9765 4049 9769
rect 4053 9765 4054 9769
rect 4058 9765 4059 9769
rect 4063 9765 4064 9769
rect 4068 9765 4069 9769
rect 4073 9765 4074 9769
rect 4078 9765 4079 9769
rect 4083 9766 4602 9769
rect 4083 9765 4100 9766
rect 3810 9762 3826 9765
rect 3774 9761 3826 9762
rect 3830 9761 3831 9765
rect 3835 9764 4100 9765
rect 3835 9761 4019 9764
rect 3774 9760 4019 9761
rect 4023 9760 4024 9764
rect 4028 9760 4029 9764
rect 4033 9760 4034 9764
rect 4038 9760 4039 9764
rect 4043 9760 4044 9764
rect 4048 9760 4049 9764
rect 4053 9760 4054 9764
rect 4058 9760 4059 9764
rect 4063 9760 4064 9764
rect 4068 9760 4069 9764
rect 4073 9760 4074 9764
rect 4078 9760 4079 9764
rect 4083 9762 4100 9764
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4119 9762 4292 9766
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4311 9762 4318 9766
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4337 9762 4344 9766
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4363 9762 4370 9766
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4389 9762 4396 9766
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4415 9762 4602 9766
rect 4083 9760 4602 9762
rect 570 9756 1354 9760
rect 1358 9756 1359 9760
rect 1363 9756 1663 9760
rect 1667 9756 1668 9760
rect 1672 9756 1972 9760
rect 1976 9756 1977 9760
rect 1981 9756 2281 9760
rect 2285 9756 2286 9760
rect 2290 9756 2590 9760
rect 2594 9756 2595 9760
rect 2599 9756 2899 9760
rect 2903 9756 2904 9760
rect 2908 9756 3208 9760
rect 3212 9756 3213 9760
rect 3217 9756 3517 9760
rect 3521 9756 3522 9760
rect 3526 9756 3652 9760
rect 3656 9756 3657 9760
rect 3661 9756 3826 9760
rect 3830 9756 3831 9760
rect 3835 9756 4602 9760
rect 570 9752 802 9756
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 821 9752 831 9756
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 850 9752 860 9756
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 879 9752 889 9756
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 908 9752 918 9756
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 937 9752 1319 9756
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1338 9755 1628 9756
rect 1338 9752 1354 9755
rect 570 9751 1354 9752
rect 1358 9751 1359 9755
rect 1363 9752 1628 9755
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1647 9755 1937 9756
rect 1647 9752 1663 9755
rect 1363 9751 1663 9752
rect 1667 9751 1668 9755
rect 1672 9752 1937 9755
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1956 9755 2246 9756
rect 1956 9752 1972 9755
rect 1672 9751 1972 9752
rect 1976 9751 1977 9755
rect 1981 9752 2246 9755
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2265 9755 2555 9756
rect 2265 9752 2281 9755
rect 1981 9751 2281 9752
rect 2285 9751 2286 9755
rect 2290 9752 2555 9755
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2574 9755 2864 9756
rect 2574 9752 2590 9755
rect 2290 9751 2590 9752
rect 2594 9751 2595 9755
rect 2599 9752 2864 9755
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2883 9755 3173 9756
rect 2883 9752 2899 9755
rect 2599 9751 2899 9752
rect 2903 9751 2904 9755
rect 2908 9752 3173 9755
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3192 9755 3482 9756
rect 3192 9752 3208 9755
rect 2908 9751 3208 9752
rect 3212 9751 3213 9755
rect 3217 9752 3482 9755
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3501 9755 3791 9756
rect 3501 9752 3517 9755
rect 3217 9751 3517 9752
rect 3521 9751 3522 9755
rect 3526 9751 3652 9755
rect 3656 9751 3657 9755
rect 3661 9752 3791 9755
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3810 9755 4100 9756
rect 3810 9752 3826 9755
rect 3661 9751 3826 9752
rect 3830 9751 3831 9755
rect 3835 9752 4100 9755
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4119 9752 4292 9756
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4311 9752 4318 9756
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4337 9752 4344 9756
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4363 9752 4370 9756
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4389 9752 4396 9756
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4415 9752 4602 9756
rect 3835 9751 4602 9752
rect 570 9750 4602 9751
rect 570 9746 1354 9750
rect 1358 9746 1359 9750
rect 1363 9746 1663 9750
rect 1667 9746 1668 9750
rect 1672 9746 1972 9750
rect 1976 9746 1977 9750
rect 1981 9746 2281 9750
rect 2285 9746 2286 9750
rect 2290 9746 2590 9750
rect 2594 9746 2595 9750
rect 2599 9746 2899 9750
rect 2903 9746 2904 9750
rect 2908 9746 3208 9750
rect 3212 9746 3213 9750
rect 3217 9746 3517 9750
rect 3521 9746 3522 9750
rect 3526 9746 3652 9750
rect 3656 9746 3657 9750
rect 3661 9746 3826 9750
rect 3830 9746 3831 9750
rect 3835 9746 4602 9750
rect 570 9742 802 9746
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 821 9742 831 9746
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 850 9742 860 9746
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 879 9742 889 9746
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 908 9742 918 9746
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 937 9742 1319 9746
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1338 9745 1628 9746
rect 1338 9742 1354 9745
rect 570 9741 1354 9742
rect 1358 9741 1359 9745
rect 1363 9742 1628 9745
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1647 9745 1937 9746
rect 1647 9742 1663 9745
rect 1363 9741 1663 9742
rect 1667 9741 1668 9745
rect 1672 9742 1937 9745
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1956 9745 2246 9746
rect 1956 9742 1972 9745
rect 1672 9741 1972 9742
rect 1976 9741 1977 9745
rect 1981 9742 2246 9745
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2265 9745 2555 9746
rect 2265 9742 2281 9745
rect 1981 9741 2281 9742
rect 2285 9741 2286 9745
rect 2290 9742 2555 9745
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2574 9745 2864 9746
rect 2574 9742 2590 9745
rect 2290 9741 2590 9742
rect 2594 9741 2595 9745
rect 2599 9742 2864 9745
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2883 9745 3173 9746
rect 2883 9742 2899 9745
rect 2599 9741 2899 9742
rect 2903 9741 2904 9745
rect 2908 9742 3173 9745
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3192 9745 3482 9746
rect 3192 9742 3208 9745
rect 2908 9741 3208 9742
rect 3212 9741 3213 9745
rect 3217 9742 3482 9745
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3501 9745 3791 9746
rect 3501 9742 3517 9745
rect 3217 9741 3517 9742
rect 3521 9741 3522 9745
rect 3526 9741 3652 9745
rect 3656 9741 3657 9745
rect 3661 9742 3791 9745
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3810 9745 4100 9746
rect 3810 9742 3826 9745
rect 3661 9741 3826 9742
rect 3830 9741 3831 9745
rect 3835 9742 4100 9745
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4119 9742 4292 9746
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4311 9742 4318 9746
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4337 9742 4344 9746
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4363 9742 4370 9746
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4389 9742 4396 9746
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4415 9742 4602 9746
rect 3835 9741 4602 9742
rect 570 9740 2167 9741
rect 570 9736 1354 9740
rect 1358 9736 1359 9740
rect 1363 9736 1663 9740
rect 1667 9736 1668 9740
rect 1672 9736 1972 9740
rect 1976 9736 1977 9740
rect 1981 9736 2167 9740
rect 2172 9740 4602 9741
rect 2172 9736 2281 9740
rect 2285 9736 2286 9740
rect 2290 9736 2590 9740
rect 2594 9736 2595 9740
rect 2599 9736 2899 9740
rect 2903 9736 2904 9740
rect 2908 9736 3208 9740
rect 3212 9736 3213 9740
rect 3217 9736 3517 9740
rect 3521 9736 3522 9740
rect 3526 9736 3826 9740
rect 3830 9736 3831 9740
rect 3835 9736 4602 9740
rect 570 9732 802 9736
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 821 9732 831 9736
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 850 9732 860 9736
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 879 9732 889 9736
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 908 9732 918 9736
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 937 9732 1319 9736
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1338 9732 1628 9736
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1647 9732 1937 9736
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1956 9732 2246 9736
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2265 9732 2555 9736
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2574 9732 2864 9736
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2883 9732 3173 9736
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3192 9732 3482 9736
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3501 9732 3791 9736
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3810 9732 4100 9736
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4119 9732 4292 9736
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4311 9732 4318 9736
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4337 9732 4344 9736
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4363 9732 4370 9736
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4389 9732 4396 9736
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 4415 9732 4602 9736
rect 570 9729 4602 9732
rect 570 9622 650 9729
rect 570 9618 613 9622
rect 617 9618 623 9622
rect 627 9618 633 9622
rect 637 9618 643 9622
rect 647 9618 650 9622
rect 570 9617 650 9618
rect 570 9613 613 9617
rect 617 9613 623 9617
rect 627 9613 633 9617
rect 637 9613 643 9617
rect 647 9613 650 9617
rect 570 9612 650 9613
rect 570 9608 613 9612
rect 617 9608 623 9612
rect 627 9608 633 9612
rect 637 9608 643 9612
rect 647 9608 650 9612
rect 570 9607 650 9608
rect 570 9603 613 9607
rect 617 9603 623 9607
rect 627 9603 633 9607
rect 637 9603 643 9607
rect 647 9603 650 9607
rect 570 9596 650 9603
rect 570 9592 613 9596
rect 617 9592 623 9596
rect 627 9592 633 9596
rect 637 9592 643 9596
rect 647 9592 650 9596
rect 570 9591 650 9592
rect 570 9587 613 9591
rect 617 9587 623 9591
rect 627 9587 633 9591
rect 637 9587 643 9591
rect 647 9587 650 9591
rect 570 9586 650 9587
rect 570 9582 613 9586
rect 617 9582 623 9586
rect 627 9582 633 9586
rect 637 9582 643 9586
rect 647 9582 650 9586
rect 570 9581 650 9582
rect 570 9577 613 9581
rect 617 9577 623 9581
rect 627 9577 633 9581
rect 637 9577 643 9581
rect 647 9577 650 9581
rect 570 9570 650 9577
rect 570 9566 613 9570
rect 617 9566 623 9570
rect 627 9566 633 9570
rect 637 9566 643 9570
rect 647 9566 650 9570
rect 570 9565 650 9566
rect 570 9561 613 9565
rect 617 9561 623 9565
rect 627 9561 633 9565
rect 637 9561 643 9565
rect 647 9561 650 9565
rect 570 9560 650 9561
rect 570 9556 613 9560
rect 617 9556 623 9560
rect 627 9556 633 9560
rect 637 9556 643 9560
rect 647 9556 650 9560
rect 570 9555 650 9556
rect 570 9551 613 9555
rect 617 9551 623 9555
rect 627 9551 633 9555
rect 637 9551 643 9555
rect 647 9551 650 9555
rect 570 9544 650 9551
rect 570 9540 613 9544
rect 617 9540 623 9544
rect 627 9540 633 9544
rect 637 9540 643 9544
rect 647 9540 650 9544
rect 570 9539 650 9540
rect 570 9535 613 9539
rect 617 9535 623 9539
rect 627 9535 633 9539
rect 637 9535 643 9539
rect 647 9535 650 9539
rect 570 9534 650 9535
rect 570 9530 613 9534
rect 617 9530 623 9534
rect 627 9530 633 9534
rect 637 9530 643 9534
rect 647 9530 650 9534
rect 570 9529 650 9530
rect 570 9525 613 9529
rect 617 9525 623 9529
rect 627 9525 633 9529
rect 637 9525 643 9529
rect 647 9525 650 9529
rect 570 9518 650 9525
rect 570 9514 613 9518
rect 617 9514 623 9518
rect 627 9514 633 9518
rect 637 9514 643 9518
rect 647 9514 650 9518
rect 570 9513 650 9514
rect 570 9509 613 9513
rect 617 9509 623 9513
rect 627 9509 633 9513
rect 637 9509 643 9513
rect 647 9509 650 9513
rect 570 9508 650 9509
rect 570 9504 613 9508
rect 617 9504 623 9508
rect 627 9504 633 9508
rect 637 9504 643 9508
rect 647 9504 650 9508
rect 570 9503 650 9504
rect 570 9499 613 9503
rect 617 9499 623 9503
rect 627 9499 633 9503
rect 637 9499 643 9503
rect 647 9499 650 9503
rect 570 9325 650 9499
rect 570 9321 613 9325
rect 617 9321 623 9325
rect 627 9321 633 9325
rect 637 9321 643 9325
rect 647 9321 650 9325
rect 570 9320 650 9321
rect 570 9316 613 9320
rect 617 9316 623 9320
rect 627 9316 633 9320
rect 637 9316 643 9320
rect 647 9316 650 9320
rect 570 9315 650 9316
rect 570 9311 613 9315
rect 617 9311 623 9315
rect 627 9311 633 9315
rect 637 9311 643 9315
rect 647 9311 650 9315
rect 570 9310 650 9311
rect 570 9306 613 9310
rect 617 9306 623 9310
rect 627 9306 633 9310
rect 637 9306 643 9310
rect 647 9306 650 9310
rect 570 9016 650 9306
rect 570 9012 613 9016
rect 617 9012 623 9016
rect 627 9012 633 9016
rect 637 9012 643 9016
rect 647 9012 650 9016
rect 570 9011 650 9012
rect 570 9007 613 9011
rect 617 9007 623 9011
rect 627 9007 633 9011
rect 637 9007 643 9011
rect 647 9007 650 9011
rect 570 9006 650 9007
rect 570 9002 613 9006
rect 617 9002 623 9006
rect 627 9002 633 9006
rect 637 9002 643 9006
rect 647 9002 650 9006
rect 570 9001 650 9002
rect 570 8997 613 9001
rect 617 8997 623 9001
rect 627 8997 633 9001
rect 637 8997 643 9001
rect 647 8997 650 9001
rect 570 8707 650 8997
rect 570 8703 613 8707
rect 617 8703 623 8707
rect 627 8703 633 8707
rect 637 8703 643 8707
rect 647 8703 650 8707
rect 570 8702 650 8703
rect 570 8698 613 8702
rect 617 8698 623 8702
rect 627 8698 633 8702
rect 637 8698 643 8702
rect 647 8698 650 8702
rect 570 8697 650 8698
rect 570 8693 613 8697
rect 617 8693 623 8697
rect 627 8693 633 8697
rect 637 8693 643 8697
rect 647 8693 650 8697
rect 570 8692 650 8693
rect 570 8688 613 8692
rect 617 8688 623 8692
rect 627 8688 633 8692
rect 637 8688 643 8692
rect 647 8688 650 8692
rect 570 8398 650 8688
rect 570 8394 613 8398
rect 617 8394 623 8398
rect 627 8394 633 8398
rect 637 8394 643 8398
rect 647 8394 650 8398
rect 570 8393 650 8394
rect 570 8389 613 8393
rect 617 8389 623 8393
rect 627 8389 633 8393
rect 637 8389 643 8393
rect 647 8389 650 8393
rect 570 8388 650 8389
rect 570 8384 613 8388
rect 617 8384 623 8388
rect 627 8384 633 8388
rect 637 8384 643 8388
rect 647 8384 650 8388
rect 570 8383 650 8384
rect 570 8379 613 8383
rect 617 8379 623 8383
rect 627 8379 633 8383
rect 637 8379 643 8383
rect 647 8379 650 8383
rect 570 8089 650 8379
rect 570 8085 613 8089
rect 617 8085 623 8089
rect 627 8085 633 8089
rect 637 8085 643 8089
rect 647 8085 650 8089
rect 570 8084 650 8085
rect 570 8080 613 8084
rect 617 8080 623 8084
rect 627 8080 633 8084
rect 637 8080 643 8084
rect 647 8080 650 8084
rect 570 8079 650 8080
rect 570 8075 613 8079
rect 617 8075 623 8079
rect 627 8075 633 8079
rect 637 8075 643 8079
rect 647 8075 650 8079
rect 570 8074 650 8075
rect 570 8070 613 8074
rect 617 8070 623 8074
rect 627 8070 633 8074
rect 637 8070 643 8074
rect 647 8070 650 8074
rect 570 7780 650 8070
rect 570 7776 613 7780
rect 617 7776 623 7780
rect 627 7776 633 7780
rect 637 7776 643 7780
rect 647 7776 650 7780
rect 570 7775 650 7776
rect 570 7771 613 7775
rect 617 7771 623 7775
rect 627 7771 633 7775
rect 637 7771 643 7775
rect 647 7771 650 7775
rect 570 7770 650 7771
rect 570 7766 613 7770
rect 617 7766 623 7770
rect 627 7766 633 7770
rect 637 7766 643 7770
rect 647 7766 650 7770
rect 570 7765 650 7766
rect 570 7761 613 7765
rect 617 7761 623 7765
rect 627 7761 633 7765
rect 637 7761 643 7765
rect 647 7761 650 7765
rect 570 7471 650 7761
rect 570 7467 613 7471
rect 617 7467 623 7471
rect 627 7467 633 7471
rect 637 7467 643 7471
rect 647 7467 650 7471
rect 570 7466 650 7467
rect 570 7462 613 7466
rect 617 7462 623 7466
rect 627 7462 633 7466
rect 637 7462 643 7466
rect 647 7462 650 7466
rect 570 7461 650 7462
rect 570 7457 613 7461
rect 617 7457 623 7461
rect 627 7457 633 7461
rect 637 7457 643 7461
rect 647 7457 650 7461
rect 570 7456 650 7457
rect 570 7452 613 7456
rect 617 7452 623 7456
rect 627 7452 633 7456
rect 637 7452 643 7456
rect 647 7452 650 7456
rect 570 7162 650 7452
rect 570 7158 613 7162
rect 617 7158 623 7162
rect 627 7158 633 7162
rect 637 7158 643 7162
rect 647 7158 650 7162
rect 570 7127 650 7158
rect 570 7123 613 7127
rect 617 7123 623 7127
rect 627 7123 633 7127
rect 637 7123 643 7127
rect 647 7123 650 7127
rect 570 7122 650 7123
rect 570 7118 613 7122
rect 617 7118 623 7122
rect 627 7118 633 7122
rect 637 7118 643 7122
rect 647 7118 650 7122
rect 570 7117 650 7118
rect 570 7113 613 7117
rect 617 7113 623 7117
rect 627 7113 633 7117
rect 637 7113 643 7117
rect 647 7113 650 7117
rect 570 7112 650 7113
rect 570 7108 613 7112
rect 617 7108 623 7112
rect 627 7108 633 7112
rect 637 7108 643 7112
rect 647 7108 650 7112
rect 570 6540 650 7108
rect 570 6536 613 6540
rect 617 6536 623 6540
rect 627 6536 633 6540
rect 637 6536 643 6540
rect 647 6536 650 6540
rect 570 6535 650 6536
rect 570 6531 613 6535
rect 617 6531 623 6535
rect 627 6531 633 6535
rect 637 6531 643 6535
rect 647 6531 650 6535
rect 570 6530 650 6531
rect 570 6526 613 6530
rect 617 6526 623 6530
rect 627 6526 633 6530
rect 637 6526 643 6530
rect 647 6526 650 6530
rect 570 6525 650 6526
rect 570 6521 613 6525
rect 617 6521 623 6525
rect 627 6521 633 6525
rect 637 6521 643 6525
rect 647 6521 650 6525
rect 570 6505 650 6521
rect 570 6501 579 6505
rect 583 6501 584 6505
rect 588 6501 589 6505
rect 593 6501 594 6505
rect 598 6501 599 6505
rect 603 6501 604 6505
rect 608 6501 609 6505
rect 613 6501 614 6505
rect 618 6501 619 6505
rect 623 6501 624 6505
rect 628 6501 629 6505
rect 633 6501 634 6505
rect 638 6501 639 6505
rect 643 6501 650 6505
rect 570 6500 650 6501
rect 570 6496 579 6500
rect 583 6496 584 6500
rect 588 6496 589 6500
rect 593 6496 594 6500
rect 598 6496 599 6500
rect 603 6496 604 6500
rect 608 6496 609 6500
rect 613 6496 614 6500
rect 618 6496 619 6500
rect 623 6496 624 6500
rect 628 6496 629 6500
rect 633 6496 634 6500
rect 638 6496 639 6500
rect 643 6496 650 6500
rect 570 6231 650 6496
rect 570 6227 613 6231
rect 617 6227 623 6231
rect 627 6227 633 6231
rect 637 6227 643 6231
rect 647 6227 650 6231
rect 570 6226 650 6227
rect 570 6222 613 6226
rect 617 6222 623 6226
rect 627 6222 633 6226
rect 637 6222 643 6226
rect 647 6222 650 6226
rect 570 6221 650 6222
rect 570 6217 613 6221
rect 617 6217 623 6221
rect 627 6217 633 6221
rect 637 6217 643 6221
rect 647 6217 650 6221
rect 570 6216 650 6217
rect 570 6212 613 6216
rect 617 6212 623 6216
rect 627 6212 633 6216
rect 637 6212 643 6216
rect 647 6212 650 6216
rect 570 6200 650 6212
rect 570 6196 613 6200
rect 617 6196 623 6200
rect 627 6196 633 6200
rect 637 6196 643 6200
rect 647 6196 650 6200
rect 570 6195 650 6196
rect 570 6191 613 6195
rect 617 6191 623 6195
rect 627 6191 633 6195
rect 637 6191 643 6195
rect 647 6191 650 6195
rect 570 6190 650 6191
rect 570 6186 613 6190
rect 617 6186 623 6190
rect 627 6186 633 6190
rect 637 6186 643 6190
rect 647 6186 650 6190
rect 570 6185 650 6186
rect 570 6181 613 6185
rect 617 6181 623 6185
rect 627 6181 633 6185
rect 637 6181 643 6185
rect 647 6181 650 6185
rect 570 5891 650 6181
rect 570 5887 613 5891
rect 617 5887 623 5891
rect 627 5887 633 5891
rect 637 5887 643 5891
rect 647 5887 650 5891
rect 570 5886 650 5887
rect 570 5882 613 5886
rect 617 5882 623 5886
rect 627 5882 633 5886
rect 637 5882 643 5886
rect 647 5882 650 5886
rect 570 5881 650 5882
rect 570 5877 613 5881
rect 617 5877 623 5881
rect 627 5877 633 5881
rect 637 5877 643 5881
rect 647 5877 650 5881
rect 570 5876 650 5877
rect 570 5872 613 5876
rect 617 5872 623 5876
rect 627 5872 633 5876
rect 637 5872 643 5876
rect 647 5872 650 5876
rect 570 5582 650 5872
rect 570 5578 613 5582
rect 617 5578 623 5582
rect 627 5578 633 5582
rect 637 5578 643 5582
rect 647 5578 650 5582
rect 570 5577 650 5578
rect 570 5573 613 5577
rect 617 5573 623 5577
rect 627 5573 633 5577
rect 637 5573 643 5577
rect 647 5573 650 5577
rect 570 5572 650 5573
rect 570 5568 613 5572
rect 617 5568 623 5572
rect 627 5568 633 5572
rect 637 5568 643 5572
rect 647 5568 650 5572
rect 570 5567 650 5568
rect 570 5563 613 5567
rect 617 5563 623 5567
rect 627 5563 633 5567
rect 637 5563 643 5567
rect 647 5563 650 5567
rect 570 5273 650 5563
rect 570 5269 613 5273
rect 617 5269 623 5273
rect 627 5269 633 5273
rect 637 5269 643 5273
rect 647 5269 650 5273
rect 570 5268 650 5269
rect 570 5264 613 5268
rect 617 5264 623 5268
rect 627 5264 633 5268
rect 637 5264 643 5268
rect 647 5264 650 5268
rect 570 5263 650 5264
rect 570 5259 613 5263
rect 617 5259 623 5263
rect 627 5259 633 5263
rect 637 5259 643 5263
rect 647 5259 650 5263
rect 570 5258 650 5259
rect 570 5254 613 5258
rect 617 5254 623 5258
rect 627 5254 633 5258
rect 637 5254 643 5258
rect 647 5254 650 5258
rect 570 4872 650 5254
rect 570 4868 613 4872
rect 617 4868 623 4872
rect 627 4868 633 4872
rect 637 4868 643 4872
rect 647 4868 650 4872
rect 570 4867 650 4868
rect 570 4863 613 4867
rect 617 4863 623 4867
rect 627 4863 633 4867
rect 637 4863 643 4867
rect 647 4863 650 4867
rect 570 4862 650 4863
rect 570 4858 613 4862
rect 617 4858 623 4862
rect 627 4858 633 4862
rect 637 4858 643 4862
rect 647 4858 650 4862
rect 570 4857 650 4858
rect 570 4853 613 4857
rect 617 4853 623 4857
rect 627 4853 633 4857
rect 637 4853 643 4857
rect 647 4853 650 4857
rect 570 4843 650 4853
rect 570 4839 613 4843
rect 617 4839 623 4843
rect 627 4839 633 4843
rect 637 4839 643 4843
rect 647 4839 650 4843
rect 570 4838 650 4839
rect 570 4834 613 4838
rect 617 4834 623 4838
rect 627 4834 633 4838
rect 637 4834 643 4838
rect 647 4834 650 4838
rect 570 4833 650 4834
rect 570 4829 613 4833
rect 617 4829 623 4833
rect 627 4829 633 4833
rect 637 4829 643 4833
rect 647 4829 650 4833
rect 570 4828 650 4829
rect 570 4824 613 4828
rect 617 4824 623 4828
rect 627 4824 633 4828
rect 637 4824 643 4828
rect 647 4824 650 4828
rect 570 4814 650 4824
rect 570 4810 613 4814
rect 617 4810 623 4814
rect 627 4810 633 4814
rect 637 4810 643 4814
rect 647 4810 650 4814
rect 570 4809 650 4810
rect 570 4805 613 4809
rect 617 4805 623 4809
rect 627 4805 633 4809
rect 637 4805 643 4809
rect 647 4805 650 4809
rect 570 4804 650 4805
rect 570 4800 613 4804
rect 617 4800 623 4804
rect 627 4800 633 4804
rect 637 4800 643 4804
rect 647 4800 650 4804
rect 570 4799 650 4800
rect 570 4795 613 4799
rect 617 4795 623 4799
rect 627 4795 633 4799
rect 637 4795 643 4799
rect 647 4795 650 4799
rect 570 4785 650 4795
rect 570 4781 613 4785
rect 617 4781 623 4785
rect 627 4781 633 4785
rect 637 4781 643 4785
rect 647 4781 650 4785
rect 570 4780 650 4781
rect 570 4776 613 4780
rect 617 4776 623 4780
rect 627 4776 633 4780
rect 637 4776 643 4780
rect 647 4776 650 4780
rect 570 4775 650 4776
rect 570 4771 613 4775
rect 617 4771 623 4775
rect 627 4771 633 4775
rect 637 4771 643 4775
rect 647 4771 650 4775
rect 570 4770 650 4771
rect 570 4766 613 4770
rect 617 4766 623 4770
rect 627 4766 633 4770
rect 637 4766 643 4770
rect 647 4766 650 4770
rect 570 4756 650 4766
rect 570 4752 613 4756
rect 617 4752 623 4756
rect 627 4752 633 4756
rect 637 4752 643 4756
rect 647 4752 650 4756
rect 570 4751 650 4752
rect 570 4747 613 4751
rect 617 4747 623 4751
rect 627 4747 633 4751
rect 637 4747 643 4751
rect 647 4747 650 4751
rect 570 4746 650 4747
rect 570 4742 613 4746
rect 617 4742 623 4746
rect 627 4742 633 4746
rect 637 4742 643 4746
rect 647 4742 650 4746
rect 570 4741 650 4742
rect 570 4737 613 4741
rect 617 4737 623 4741
rect 627 4737 633 4741
rect 637 4737 643 4741
rect 647 4737 650 4741
rect 570 4585 650 4737
rect 654 9720 4518 9725
rect 654 9716 802 9720
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 821 9716 831 9720
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 850 9716 860 9720
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 879 9716 889 9720
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 908 9716 918 9720
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 937 9716 1319 9720
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1338 9716 1628 9720
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1647 9716 1937 9720
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1956 9716 2246 9720
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2265 9716 2555 9720
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2574 9716 2864 9720
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2883 9716 3173 9720
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3192 9716 3482 9720
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3501 9716 3791 9720
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3810 9716 4100 9720
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4119 9716 4292 9720
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4311 9716 4318 9720
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4337 9716 4344 9720
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4363 9716 4370 9720
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4389 9716 4396 9720
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4415 9716 4518 9720
rect 654 9715 4518 9716
rect 654 9712 1489 9715
rect 654 9710 1387 9712
rect 654 9706 802 9710
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 821 9706 831 9710
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 850 9706 860 9710
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 879 9706 889 9710
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 908 9706 918 9710
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 937 9706 1319 9710
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1338 9708 1387 9710
rect 1391 9708 1392 9712
rect 1396 9708 1397 9712
rect 1401 9708 1402 9712
rect 1406 9708 1407 9712
rect 1411 9708 1412 9712
rect 1416 9708 1417 9712
rect 1421 9708 1422 9712
rect 1426 9708 1427 9712
rect 1431 9708 1432 9712
rect 1436 9708 1437 9712
rect 1441 9708 1442 9712
rect 1446 9708 1447 9712
rect 1451 9711 1489 9712
rect 1493 9711 1494 9715
rect 1498 9712 3343 9715
rect 1498 9711 1569 9712
rect 1451 9710 1569 9711
rect 1451 9708 1489 9710
rect 1338 9707 1489 9708
rect 1338 9706 1387 9707
rect 654 9703 1387 9706
rect 1391 9703 1392 9707
rect 1396 9703 1397 9707
rect 1401 9703 1402 9707
rect 1406 9703 1407 9707
rect 1411 9703 1412 9707
rect 1416 9703 1417 9707
rect 1421 9703 1422 9707
rect 1426 9703 1427 9707
rect 1431 9703 1432 9707
rect 1436 9703 1437 9707
rect 1441 9703 1442 9707
rect 1446 9703 1447 9707
rect 1451 9706 1489 9707
rect 1493 9706 1494 9710
rect 1498 9708 1569 9710
rect 1573 9708 1574 9712
rect 1578 9708 1579 9712
rect 1583 9708 1584 9712
rect 1588 9708 1589 9712
rect 1593 9708 1594 9712
rect 1598 9708 1599 9712
rect 1603 9708 1604 9712
rect 1608 9708 1609 9712
rect 1613 9708 1614 9712
rect 1618 9708 1619 9712
rect 1623 9710 1696 9712
rect 1623 9708 1628 9710
rect 1498 9707 1628 9708
rect 1498 9706 1569 9707
rect 1451 9705 1569 9706
rect 1451 9703 1489 9705
rect 654 9701 1489 9703
rect 1493 9701 1494 9705
rect 1498 9703 1569 9705
rect 1573 9703 1574 9707
rect 1578 9703 1579 9707
rect 1583 9703 1584 9707
rect 1588 9703 1589 9707
rect 1593 9703 1594 9707
rect 1598 9703 1599 9707
rect 1603 9703 1604 9707
rect 1608 9703 1609 9707
rect 1613 9703 1614 9707
rect 1618 9703 1619 9707
rect 1623 9706 1628 9707
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1647 9708 1696 9710
rect 1700 9708 1701 9712
rect 1705 9708 1706 9712
rect 1710 9708 1711 9712
rect 1715 9708 1716 9712
rect 1720 9708 1721 9712
rect 1725 9708 1726 9712
rect 1730 9708 1731 9712
rect 1735 9708 1736 9712
rect 1740 9708 1741 9712
rect 1745 9708 1746 9712
rect 1750 9708 1751 9712
rect 1755 9708 1756 9712
rect 1760 9708 1878 9712
rect 1882 9708 1883 9712
rect 1887 9708 1888 9712
rect 1892 9708 1893 9712
rect 1897 9708 1898 9712
rect 1902 9708 1903 9712
rect 1907 9708 1908 9712
rect 1912 9708 1913 9712
rect 1917 9708 1918 9712
rect 1922 9708 1923 9712
rect 1927 9708 1928 9712
rect 1932 9710 2005 9712
rect 1932 9708 1937 9710
rect 1647 9707 1937 9708
rect 1647 9706 1696 9707
rect 1623 9703 1696 9706
rect 1700 9703 1701 9707
rect 1705 9703 1706 9707
rect 1710 9703 1711 9707
rect 1715 9703 1716 9707
rect 1720 9703 1721 9707
rect 1725 9703 1726 9707
rect 1730 9703 1731 9707
rect 1735 9703 1736 9707
rect 1740 9703 1741 9707
rect 1745 9703 1746 9707
rect 1750 9703 1751 9707
rect 1755 9703 1756 9707
rect 1760 9703 1878 9707
rect 1882 9703 1883 9707
rect 1887 9703 1888 9707
rect 1892 9703 1893 9707
rect 1897 9703 1898 9707
rect 1902 9703 1903 9707
rect 1907 9703 1908 9707
rect 1912 9703 1913 9707
rect 1917 9703 1918 9707
rect 1922 9703 1923 9707
rect 1927 9703 1928 9707
rect 1932 9706 1937 9707
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1956 9708 2005 9710
rect 2009 9708 2010 9712
rect 2014 9708 2015 9712
rect 2019 9708 2020 9712
rect 2024 9708 2025 9712
rect 2029 9708 2030 9712
rect 2034 9708 2035 9712
rect 2039 9708 2040 9712
rect 2044 9708 2045 9712
rect 2049 9708 2050 9712
rect 2054 9708 2055 9712
rect 2059 9708 2060 9712
rect 2064 9708 2065 9712
rect 2069 9708 2187 9712
rect 2191 9708 2192 9712
rect 2196 9708 2197 9712
rect 2201 9708 2202 9712
rect 2206 9708 2207 9712
rect 2211 9708 2212 9712
rect 2216 9708 2217 9712
rect 2221 9708 2222 9712
rect 2226 9708 2227 9712
rect 2231 9708 2232 9712
rect 2236 9708 2237 9712
rect 2241 9710 2314 9712
rect 2241 9708 2246 9710
rect 1956 9707 2246 9708
rect 1956 9706 2005 9707
rect 1932 9703 2005 9706
rect 2009 9703 2010 9707
rect 2014 9703 2015 9707
rect 2019 9703 2020 9707
rect 2024 9703 2025 9707
rect 2029 9703 2030 9707
rect 2034 9703 2035 9707
rect 2039 9703 2040 9707
rect 2044 9703 2045 9707
rect 2049 9703 2050 9707
rect 2054 9703 2055 9707
rect 2059 9703 2060 9707
rect 2064 9703 2065 9707
rect 2069 9703 2187 9707
rect 2191 9703 2192 9707
rect 2196 9703 2197 9707
rect 2201 9703 2202 9707
rect 2206 9703 2207 9707
rect 2211 9703 2212 9707
rect 2216 9703 2217 9707
rect 2221 9703 2222 9707
rect 2226 9703 2227 9707
rect 2231 9703 2232 9707
rect 2236 9703 2237 9707
rect 2241 9706 2246 9707
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2265 9708 2314 9710
rect 2318 9708 2319 9712
rect 2323 9708 2324 9712
rect 2328 9708 2329 9712
rect 2333 9708 2334 9712
rect 2338 9708 2339 9712
rect 2343 9708 2344 9712
rect 2348 9708 2349 9712
rect 2353 9708 2354 9712
rect 2358 9708 2359 9712
rect 2363 9708 2364 9712
rect 2368 9708 2369 9712
rect 2373 9708 2374 9712
rect 2378 9708 2496 9712
rect 2500 9708 2501 9712
rect 2505 9708 2506 9712
rect 2510 9708 2511 9712
rect 2515 9708 2516 9712
rect 2520 9708 2521 9712
rect 2525 9708 2526 9712
rect 2530 9708 2531 9712
rect 2535 9708 2536 9712
rect 2540 9708 2541 9712
rect 2545 9708 2546 9712
rect 2550 9710 2623 9712
rect 2550 9708 2555 9710
rect 2265 9707 2555 9708
rect 2265 9706 2314 9707
rect 2241 9703 2314 9706
rect 2318 9703 2319 9707
rect 2323 9703 2324 9707
rect 2328 9703 2329 9707
rect 2333 9703 2334 9707
rect 2338 9703 2339 9707
rect 2343 9703 2344 9707
rect 2348 9703 2349 9707
rect 2353 9703 2354 9707
rect 2358 9703 2359 9707
rect 2363 9703 2364 9707
rect 2368 9703 2369 9707
rect 2373 9703 2374 9707
rect 2378 9703 2496 9707
rect 2500 9703 2501 9707
rect 2505 9703 2506 9707
rect 2510 9703 2511 9707
rect 2515 9703 2516 9707
rect 2520 9703 2521 9707
rect 2525 9703 2526 9707
rect 2530 9703 2531 9707
rect 2535 9703 2536 9707
rect 2540 9703 2541 9707
rect 2545 9703 2546 9707
rect 2550 9706 2555 9707
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2574 9708 2623 9710
rect 2627 9708 2628 9712
rect 2632 9708 2633 9712
rect 2637 9708 2638 9712
rect 2642 9708 2643 9712
rect 2647 9708 2648 9712
rect 2652 9708 2653 9712
rect 2657 9708 2658 9712
rect 2662 9708 2663 9712
rect 2667 9708 2668 9712
rect 2672 9708 2673 9712
rect 2677 9708 2678 9712
rect 2682 9708 2683 9712
rect 2687 9708 2805 9712
rect 2809 9708 2810 9712
rect 2814 9708 2815 9712
rect 2819 9708 2820 9712
rect 2824 9708 2825 9712
rect 2829 9708 2830 9712
rect 2834 9708 2835 9712
rect 2839 9708 2840 9712
rect 2844 9708 2845 9712
rect 2849 9708 2850 9712
rect 2854 9708 2855 9712
rect 2859 9710 2932 9712
rect 2859 9708 2864 9710
rect 2574 9707 2864 9708
rect 2574 9706 2623 9707
rect 2550 9703 2623 9706
rect 2627 9703 2628 9707
rect 2632 9703 2633 9707
rect 2637 9703 2638 9707
rect 2642 9703 2643 9707
rect 2647 9703 2648 9707
rect 2652 9703 2653 9707
rect 2657 9703 2658 9707
rect 2662 9703 2663 9707
rect 2667 9703 2668 9707
rect 2672 9703 2673 9707
rect 2677 9703 2678 9707
rect 2682 9703 2683 9707
rect 2687 9703 2805 9707
rect 2809 9703 2810 9707
rect 2814 9703 2815 9707
rect 2819 9703 2820 9707
rect 2824 9703 2825 9707
rect 2829 9703 2830 9707
rect 2834 9703 2835 9707
rect 2839 9703 2840 9707
rect 2844 9703 2845 9707
rect 2849 9703 2850 9707
rect 2854 9703 2855 9707
rect 2859 9706 2864 9707
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2883 9708 2932 9710
rect 2936 9708 2937 9712
rect 2941 9708 2942 9712
rect 2946 9708 2947 9712
rect 2951 9708 2952 9712
rect 2956 9708 2957 9712
rect 2961 9708 2962 9712
rect 2966 9708 2967 9712
rect 2971 9708 2972 9712
rect 2976 9708 2977 9712
rect 2981 9708 2982 9712
rect 2986 9708 2987 9712
rect 2991 9708 2992 9712
rect 2996 9708 3114 9712
rect 3118 9708 3119 9712
rect 3123 9708 3124 9712
rect 3128 9708 3129 9712
rect 3133 9708 3134 9712
rect 3138 9708 3139 9712
rect 3143 9708 3144 9712
rect 3148 9708 3149 9712
rect 3153 9708 3154 9712
rect 3158 9708 3159 9712
rect 3163 9708 3164 9712
rect 3168 9710 3241 9712
rect 3168 9708 3173 9710
rect 2883 9707 3173 9708
rect 2883 9706 2932 9707
rect 2859 9703 2932 9706
rect 2936 9703 2937 9707
rect 2941 9703 2942 9707
rect 2946 9703 2947 9707
rect 2951 9703 2952 9707
rect 2956 9703 2957 9707
rect 2961 9703 2962 9707
rect 2966 9703 2967 9707
rect 2971 9703 2972 9707
rect 2976 9703 2977 9707
rect 2981 9703 2982 9707
rect 2986 9703 2987 9707
rect 2991 9703 2992 9707
rect 2996 9703 3114 9707
rect 3118 9703 3119 9707
rect 3123 9703 3124 9707
rect 3128 9703 3129 9707
rect 3133 9703 3134 9707
rect 3138 9703 3139 9707
rect 3143 9703 3144 9707
rect 3148 9703 3149 9707
rect 3153 9703 3154 9707
rect 3158 9703 3159 9707
rect 3163 9703 3164 9707
rect 3168 9706 3173 9707
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3192 9708 3241 9710
rect 3245 9708 3246 9712
rect 3250 9708 3251 9712
rect 3255 9708 3256 9712
rect 3260 9708 3261 9712
rect 3265 9708 3266 9712
rect 3270 9708 3271 9712
rect 3275 9708 3276 9712
rect 3280 9708 3281 9712
rect 3285 9708 3286 9712
rect 3290 9708 3291 9712
rect 3295 9708 3296 9712
rect 3300 9708 3301 9712
rect 3305 9711 3343 9712
rect 3347 9711 3348 9715
rect 3352 9712 4518 9715
rect 3352 9711 3423 9712
rect 3305 9710 3423 9711
rect 3305 9708 3343 9710
rect 3192 9707 3343 9708
rect 3192 9706 3241 9707
rect 3168 9703 3241 9706
rect 3245 9703 3246 9707
rect 3250 9703 3251 9707
rect 3255 9703 3256 9707
rect 3260 9703 3261 9707
rect 3265 9703 3266 9707
rect 3270 9703 3271 9707
rect 3275 9703 3276 9707
rect 3280 9703 3281 9707
rect 3285 9703 3286 9707
rect 3290 9703 3291 9707
rect 3295 9703 3296 9707
rect 3300 9703 3301 9707
rect 3305 9706 3343 9707
rect 3347 9706 3348 9710
rect 3352 9708 3423 9710
rect 3427 9708 3428 9712
rect 3432 9708 3433 9712
rect 3437 9708 3438 9712
rect 3442 9708 3443 9712
rect 3447 9708 3448 9712
rect 3452 9708 3453 9712
rect 3457 9708 3458 9712
rect 3462 9708 3463 9712
rect 3467 9708 3468 9712
rect 3472 9708 3473 9712
rect 3477 9710 3550 9712
rect 3477 9708 3482 9710
rect 3352 9707 3482 9708
rect 3352 9706 3423 9707
rect 3305 9705 3423 9706
rect 3305 9703 3343 9705
rect 1498 9701 3343 9703
rect 3347 9701 3348 9705
rect 3352 9703 3423 9705
rect 3427 9703 3428 9707
rect 3432 9703 3433 9707
rect 3437 9703 3438 9707
rect 3442 9703 3443 9707
rect 3447 9703 3448 9707
rect 3452 9703 3453 9707
rect 3457 9703 3458 9707
rect 3462 9703 3463 9707
rect 3467 9703 3468 9707
rect 3472 9703 3473 9707
rect 3477 9706 3482 9707
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3501 9708 3550 9710
rect 3554 9708 3555 9712
rect 3559 9708 3560 9712
rect 3564 9708 3565 9712
rect 3569 9708 3570 9712
rect 3574 9708 3575 9712
rect 3579 9708 3580 9712
rect 3584 9708 3585 9712
rect 3589 9708 3590 9712
rect 3594 9708 3595 9712
rect 3599 9708 3600 9712
rect 3604 9708 3605 9712
rect 3609 9708 3610 9712
rect 3614 9708 3732 9712
rect 3736 9708 3737 9712
rect 3741 9708 3742 9712
rect 3746 9708 3747 9712
rect 3751 9708 3752 9712
rect 3756 9708 3757 9712
rect 3761 9708 3762 9712
rect 3766 9708 3767 9712
rect 3771 9708 3772 9712
rect 3776 9708 3777 9712
rect 3781 9708 3782 9712
rect 3786 9710 3859 9712
rect 3786 9708 3791 9710
rect 3501 9707 3791 9708
rect 3501 9706 3550 9707
rect 3477 9703 3550 9706
rect 3554 9703 3555 9707
rect 3559 9703 3560 9707
rect 3564 9703 3565 9707
rect 3569 9703 3570 9707
rect 3574 9703 3575 9707
rect 3579 9703 3580 9707
rect 3584 9703 3585 9707
rect 3589 9703 3590 9707
rect 3594 9703 3595 9707
rect 3599 9703 3600 9707
rect 3604 9703 3605 9707
rect 3609 9703 3610 9707
rect 3614 9703 3732 9707
rect 3736 9703 3737 9707
rect 3741 9703 3742 9707
rect 3746 9703 3747 9707
rect 3751 9703 3752 9707
rect 3756 9703 3757 9707
rect 3761 9703 3762 9707
rect 3766 9703 3767 9707
rect 3771 9703 3772 9707
rect 3776 9703 3777 9707
rect 3781 9703 3782 9707
rect 3786 9706 3791 9707
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3810 9708 3859 9710
rect 3863 9708 3864 9712
rect 3868 9708 3869 9712
rect 3873 9708 3874 9712
rect 3878 9708 3879 9712
rect 3883 9708 3884 9712
rect 3888 9708 3889 9712
rect 3893 9708 3894 9712
rect 3898 9708 3899 9712
rect 3903 9708 3904 9712
rect 3908 9708 3909 9712
rect 3913 9708 3914 9712
rect 3918 9708 3919 9712
rect 3923 9708 4041 9712
rect 4045 9708 4046 9712
rect 4050 9708 4051 9712
rect 4055 9708 4056 9712
rect 4060 9708 4061 9712
rect 4065 9708 4066 9712
rect 4070 9708 4071 9712
rect 4075 9708 4076 9712
rect 4080 9708 4081 9712
rect 4085 9708 4086 9712
rect 4090 9708 4091 9712
rect 4095 9710 4518 9712
rect 4095 9708 4100 9710
rect 3810 9707 4100 9708
rect 3810 9706 3859 9707
rect 3786 9703 3859 9706
rect 3863 9703 3864 9707
rect 3868 9703 3869 9707
rect 3873 9703 3874 9707
rect 3878 9703 3879 9707
rect 3883 9703 3884 9707
rect 3888 9703 3889 9707
rect 3893 9703 3894 9707
rect 3898 9703 3899 9707
rect 3903 9703 3904 9707
rect 3908 9703 3909 9707
rect 3913 9703 3914 9707
rect 3918 9703 3919 9707
rect 3923 9703 4041 9707
rect 4045 9703 4046 9707
rect 4050 9703 4051 9707
rect 4055 9703 4056 9707
rect 4060 9703 4061 9707
rect 4065 9703 4066 9707
rect 4070 9703 4071 9707
rect 4075 9703 4076 9707
rect 4080 9703 4081 9707
rect 4085 9703 4086 9707
rect 4090 9703 4091 9707
rect 4095 9706 4100 9707
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4119 9706 4292 9710
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4311 9706 4318 9710
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4337 9706 4344 9710
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4363 9706 4370 9710
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4389 9706 4396 9710
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4415 9706 4518 9710
rect 4095 9703 4518 9706
rect 3352 9701 4518 9703
rect 654 9700 4518 9701
rect 654 9696 802 9700
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 821 9696 831 9700
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 850 9696 860 9700
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 879 9696 889 9700
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 908 9696 918 9700
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 937 9696 1319 9700
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1338 9696 1489 9700
rect 1493 9696 1494 9700
rect 1498 9696 1628 9700
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1647 9696 1937 9700
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1956 9696 2246 9700
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2265 9696 2555 9700
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2574 9696 2864 9700
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2883 9696 3173 9700
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3192 9696 3343 9700
rect 3347 9696 3348 9700
rect 3352 9696 3482 9700
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3501 9696 3791 9700
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3810 9696 4100 9700
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4119 9696 4292 9700
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4311 9696 4318 9700
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4337 9696 4344 9700
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4363 9696 4370 9700
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4389 9696 4396 9700
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4415 9696 4518 9700
rect 654 9695 4518 9696
rect 654 9691 1489 9695
rect 1493 9691 1494 9695
rect 1498 9691 3343 9695
rect 3347 9691 3348 9695
rect 3352 9691 4518 9695
rect 654 9690 4518 9691
rect 654 9686 802 9690
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 821 9686 831 9690
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 850 9686 860 9690
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 879 9686 889 9690
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 908 9686 918 9690
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 937 9686 1319 9690
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1338 9686 1489 9690
rect 1493 9686 1494 9690
rect 1498 9686 1628 9690
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1647 9686 1937 9690
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 1956 9686 2246 9690
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2265 9686 2555 9690
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2574 9686 2864 9690
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 2883 9686 3173 9690
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3192 9686 3343 9690
rect 3347 9686 3348 9690
rect 3352 9686 3482 9690
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 3501 9686 3791 9690
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 3810 9686 4100 9690
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4119 9686 4292 9690
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4311 9686 4318 9690
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4337 9686 4344 9690
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4363 9686 4370 9690
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4389 9686 4396 9690
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 4415 9686 4518 9690
rect 654 9685 4518 9686
rect 654 9681 1489 9685
rect 1493 9681 1494 9685
rect 1498 9681 3343 9685
rect 3347 9681 3348 9685
rect 3352 9681 4518 9685
rect 654 9680 4518 9681
rect 654 9676 1489 9680
rect 1493 9676 1494 9680
rect 1498 9676 3343 9680
rect 3347 9676 3348 9680
rect 3352 9676 4518 9680
rect 654 9675 4518 9676
rect 654 9671 1489 9675
rect 1493 9671 1494 9675
rect 1498 9671 3343 9675
rect 3347 9671 3348 9675
rect 3352 9671 4518 9675
rect 654 9670 4518 9671
rect 654 9666 1489 9670
rect 1493 9666 1494 9670
rect 1498 9666 3343 9670
rect 3347 9666 3348 9670
rect 3352 9666 4518 9670
rect 654 9665 4518 9666
rect 654 9661 1489 9665
rect 1493 9661 1494 9665
rect 1498 9661 3343 9665
rect 3347 9661 3348 9665
rect 3352 9661 4518 9665
rect 654 9623 4518 9661
rect 654 9622 2258 9623
rect 654 9618 659 9622
rect 663 9618 669 9622
rect 673 9618 679 9622
rect 683 9618 689 9622
rect 693 9619 2258 9622
rect 2262 9619 4518 9623
rect 693 9618 4518 9619
rect 654 9617 4518 9618
rect 654 9613 659 9617
rect 663 9613 669 9617
rect 673 9613 679 9617
rect 683 9613 689 9617
rect 693 9613 4518 9617
rect 654 9612 4518 9613
rect 654 9608 659 9612
rect 663 9608 669 9612
rect 673 9608 679 9612
rect 683 9608 689 9612
rect 693 9610 4518 9612
rect 693 9608 769 9610
rect 654 9607 769 9608
rect 654 9603 659 9607
rect 663 9603 669 9607
rect 673 9603 679 9607
rect 683 9603 689 9607
rect 693 9603 769 9607
rect 654 9596 769 9603
rect 654 9592 659 9596
rect 663 9592 669 9596
rect 673 9592 679 9596
rect 683 9592 689 9596
rect 693 9592 769 9596
rect 654 9591 769 9592
rect 654 9587 659 9591
rect 663 9587 669 9591
rect 673 9587 679 9591
rect 683 9587 689 9591
rect 693 9587 769 9591
rect 654 9586 769 9587
rect 654 9582 659 9586
rect 663 9582 669 9586
rect 673 9582 679 9586
rect 683 9582 689 9586
rect 693 9582 769 9586
rect 654 9581 769 9582
rect 654 9577 659 9581
rect 663 9577 669 9581
rect 673 9577 679 9581
rect 683 9577 689 9581
rect 693 9577 769 9581
rect 654 9570 769 9577
rect 654 9566 659 9570
rect 663 9566 669 9570
rect 673 9566 679 9570
rect 683 9566 689 9570
rect 693 9566 769 9570
rect 654 9565 769 9566
rect 654 9561 659 9565
rect 663 9561 669 9565
rect 673 9561 679 9565
rect 683 9561 689 9565
rect 693 9561 769 9565
rect 654 9560 769 9561
rect 654 9556 659 9560
rect 663 9556 669 9560
rect 673 9556 679 9560
rect 683 9556 689 9560
rect 693 9556 769 9560
rect 654 9555 769 9556
rect 654 9551 659 9555
rect 663 9551 669 9555
rect 673 9551 679 9555
rect 683 9551 689 9555
rect 693 9551 769 9555
rect 654 9544 769 9551
rect 654 9540 659 9544
rect 663 9540 669 9544
rect 673 9540 679 9544
rect 683 9540 689 9544
rect 693 9540 769 9544
rect 654 9539 769 9540
rect 654 9535 659 9539
rect 663 9535 669 9539
rect 673 9535 679 9539
rect 683 9535 689 9539
rect 693 9535 769 9539
rect 654 9534 769 9535
rect 654 9530 659 9534
rect 663 9530 669 9534
rect 673 9530 679 9534
rect 683 9530 689 9534
rect 693 9530 769 9534
rect 654 9529 769 9530
rect 654 9525 659 9529
rect 663 9525 669 9529
rect 673 9525 679 9529
rect 683 9525 689 9529
rect 693 9525 769 9529
rect 654 9518 769 9525
rect 654 9514 659 9518
rect 663 9514 669 9518
rect 673 9514 679 9518
rect 683 9514 689 9518
rect 693 9514 769 9518
rect 654 9513 769 9514
rect 654 9509 659 9513
rect 663 9509 669 9513
rect 673 9509 679 9513
rect 683 9509 689 9513
rect 693 9509 769 9513
rect 654 9508 769 9509
rect 654 9504 659 9508
rect 663 9504 669 9508
rect 673 9504 679 9508
rect 683 9504 689 9508
rect 693 9504 769 9508
rect 654 9503 769 9504
rect 654 9499 659 9503
rect 663 9499 669 9503
rect 673 9499 679 9503
rect 683 9499 689 9503
rect 693 9499 769 9503
rect 654 9325 769 9499
rect 654 9321 659 9325
rect 663 9321 669 9325
rect 673 9321 679 9325
rect 683 9321 689 9325
rect 693 9321 769 9325
rect 654 9320 769 9321
rect 654 9316 659 9320
rect 663 9316 669 9320
rect 673 9316 679 9320
rect 683 9316 689 9320
rect 693 9316 769 9320
rect 4403 9577 4518 9610
rect 4403 9573 4479 9577
rect 4483 9573 4489 9577
rect 4493 9573 4499 9577
rect 4503 9573 4509 9577
rect 4513 9573 4518 9577
rect 4403 9572 4518 9573
rect 4403 9568 4479 9572
rect 4483 9568 4489 9572
rect 4493 9568 4499 9572
rect 4503 9568 4509 9572
rect 4513 9568 4518 9572
rect 4403 9567 4518 9568
rect 4403 9563 4479 9567
rect 4483 9563 4489 9567
rect 4493 9563 4499 9567
rect 4503 9563 4509 9567
rect 4513 9563 4518 9567
rect 4403 9562 4518 9563
rect 4403 9558 4479 9562
rect 4483 9558 4489 9562
rect 4493 9558 4499 9562
rect 4503 9558 4509 9562
rect 4513 9558 4518 9562
rect 4403 9548 4518 9558
rect 4403 9544 4479 9548
rect 4483 9544 4489 9548
rect 4493 9544 4499 9548
rect 4503 9544 4509 9548
rect 4513 9544 4518 9548
rect 4403 9543 4518 9544
rect 4403 9539 4479 9543
rect 4483 9539 4489 9543
rect 4493 9539 4499 9543
rect 4503 9539 4509 9543
rect 4513 9539 4518 9543
rect 4403 9538 4518 9539
rect 4403 9534 4479 9538
rect 4483 9534 4489 9538
rect 4493 9534 4499 9538
rect 4503 9534 4509 9538
rect 4513 9534 4518 9538
rect 4403 9533 4518 9534
rect 4403 9529 4479 9533
rect 4483 9529 4489 9533
rect 4493 9529 4499 9533
rect 4503 9529 4509 9533
rect 4513 9529 4518 9533
rect 4403 9519 4518 9529
rect 4403 9515 4479 9519
rect 4483 9515 4489 9519
rect 4493 9515 4499 9519
rect 4503 9515 4509 9519
rect 4513 9515 4518 9519
rect 4403 9514 4518 9515
rect 4403 9510 4479 9514
rect 4483 9510 4489 9514
rect 4493 9510 4499 9514
rect 4503 9510 4509 9514
rect 4513 9510 4518 9514
rect 4403 9509 4518 9510
rect 4403 9505 4479 9509
rect 4483 9505 4489 9509
rect 4493 9505 4499 9509
rect 4503 9505 4509 9509
rect 4513 9505 4518 9509
rect 4403 9504 4518 9505
rect 4403 9500 4479 9504
rect 4483 9500 4489 9504
rect 4493 9500 4499 9504
rect 4503 9500 4509 9504
rect 4513 9500 4518 9504
rect 4403 9490 4518 9500
rect 4403 9486 4479 9490
rect 4483 9486 4489 9490
rect 4493 9486 4499 9490
rect 4503 9486 4509 9490
rect 4513 9486 4518 9490
rect 4403 9485 4518 9486
rect 4403 9481 4479 9485
rect 4483 9481 4489 9485
rect 4493 9481 4499 9485
rect 4503 9481 4509 9485
rect 4513 9481 4518 9485
rect 4403 9480 4518 9481
rect 4403 9476 4479 9480
rect 4483 9476 4489 9480
rect 4493 9476 4499 9480
rect 4503 9476 4509 9480
rect 4513 9476 4518 9480
rect 4403 9475 4518 9476
rect 4403 9471 4479 9475
rect 4483 9471 4489 9475
rect 4493 9471 4499 9475
rect 4503 9471 4509 9475
rect 4513 9471 4518 9475
rect 4403 9461 4518 9471
rect 4403 9457 4479 9461
rect 4483 9457 4489 9461
rect 4493 9457 4499 9461
rect 4503 9457 4509 9461
rect 4513 9457 4518 9461
rect 4403 9456 4518 9457
rect 4403 9452 4479 9456
rect 4483 9452 4489 9456
rect 4493 9452 4499 9456
rect 4503 9452 4509 9456
rect 4513 9452 4518 9456
rect 4403 9451 4518 9452
rect 4403 9447 4479 9451
rect 4483 9447 4489 9451
rect 4493 9447 4499 9451
rect 4503 9447 4509 9451
rect 4513 9447 4518 9451
rect 4403 9446 4518 9447
rect 4403 9442 4479 9446
rect 4483 9442 4489 9446
rect 4493 9442 4499 9446
rect 4503 9442 4509 9446
rect 4513 9442 4518 9446
rect 654 9315 769 9316
rect 654 9311 659 9315
rect 663 9311 669 9315
rect 673 9311 679 9315
rect 683 9311 689 9315
rect 693 9311 769 9315
rect 654 9310 769 9311
rect 654 9306 659 9310
rect 663 9306 669 9310
rect 673 9306 679 9310
rect 683 9306 689 9310
rect 693 9306 769 9310
rect 654 9016 769 9306
rect 2846 9317 2852 9318
rect 2846 9313 2847 9317
rect 2851 9313 2852 9317
rect 2846 9312 2852 9313
rect 3791 9317 3797 9318
rect 3791 9313 3792 9317
rect 3796 9313 3797 9317
rect 3791 9312 3797 9313
rect 2846 9282 2851 9312
rect 3791 9282 3796 9312
rect 2623 9281 2851 9282
rect 2623 9277 2624 9281
rect 2628 9277 2851 9281
rect 3568 9281 3796 9282
rect 3568 9277 3569 9281
rect 3573 9277 3796 9281
rect 2623 9276 2629 9277
rect 3568 9276 3574 9277
rect 3302 9266 3308 9267
rect 3302 9262 3303 9266
rect 3307 9262 3308 9266
rect 3302 9261 3308 9262
rect 4247 9266 4253 9267
rect 4247 9262 4248 9266
rect 4252 9262 4253 9266
rect 4247 9261 4253 9262
rect 2887 9240 2927 9241
rect 2887 9236 2921 9240
rect 2886 9235 2893 9236
rect 2886 9230 2887 9235
rect 2892 9230 2893 9235
rect 2920 9235 2921 9236
rect 2926 9235 2927 9240
rect 2959 9240 2995 9245
rect 2920 9234 2927 9235
rect 2944 9235 2951 9236
rect 2886 9229 2893 9230
rect 2897 9231 2904 9232
rect 2897 9226 2898 9231
rect 2903 9226 2904 9231
rect 2944 9230 2945 9235
rect 2950 9230 2951 9235
rect 2959 9234 2960 9240
rect 2965 9239 2995 9240
rect 2965 9234 2966 9239
rect 2990 9236 2995 9239
rect 2959 9233 2966 9234
rect 2989 9235 2996 9236
rect 2989 9230 2990 9235
rect 2995 9230 2996 9235
rect 3018 9234 3025 9235
rect 2944 9229 2951 9230
rect 2973 9229 2980 9230
rect 2989 9229 2996 9230
rect 3002 9229 3008 9230
rect 2945 9226 2950 9229
rect 2897 9221 2950 9226
rect 2973 9224 2974 9229
rect 2979 9224 2980 9229
rect 3002 9224 3003 9229
rect 3007 9224 3008 9229
rect 2973 9223 3008 9224
rect 2974 9219 3008 9223
rect 3018 9229 3019 9234
rect 3024 9229 3025 9234
rect 3100 9234 3107 9235
rect 3100 9229 3101 9234
rect 3106 9229 3107 9234
rect 3185 9234 3192 9235
rect 3185 9229 3186 9234
rect 3191 9229 3192 9234
rect 3018 9228 3025 9229
rect 3044 9228 3051 9229
rect 3100 9228 3107 9229
rect 3125 9228 3132 9229
rect 3185 9228 3192 9229
rect 3018 9223 3045 9228
rect 3050 9223 3051 9228
rect 3101 9223 3126 9228
rect 3131 9223 3132 9228
rect 3018 9202 3023 9223
rect 3044 9222 3051 9223
rect 3125 9222 3132 9223
rect 3182 9223 3191 9228
rect 2851 9196 3023 9202
rect 2622 9178 2628 9179
rect 2622 9174 2623 9178
rect 2627 9174 2760 9178
rect 2851 9176 2856 9196
rect 2622 9173 2760 9174
rect 654 9012 659 9016
rect 663 9012 669 9016
rect 673 9012 679 9016
rect 683 9012 689 9016
rect 693 9012 769 9016
rect 654 9011 769 9012
rect 654 9007 659 9011
rect 663 9007 669 9011
rect 673 9007 679 9011
rect 683 9007 689 9011
rect 693 9007 769 9011
rect 654 9006 769 9007
rect 654 9002 659 9006
rect 663 9002 669 9006
rect 673 9002 679 9006
rect 683 9002 689 9006
rect 693 9002 769 9006
rect 654 9001 769 9002
rect 654 8997 659 9001
rect 663 8997 669 9001
rect 673 8997 679 9001
rect 683 8997 689 9001
rect 693 8997 769 9001
rect 654 8707 769 8997
rect 654 8703 659 8707
rect 663 8703 669 8707
rect 673 8703 679 8707
rect 683 8703 689 8707
rect 693 8703 769 8707
rect 654 8702 769 8703
rect 654 8698 659 8702
rect 663 8698 669 8702
rect 673 8698 679 8702
rect 683 8698 689 8702
rect 693 8698 769 8702
rect 654 8697 769 8698
rect 654 8693 659 8697
rect 663 8693 669 8697
rect 673 8693 679 8697
rect 683 8693 689 8697
rect 693 8693 769 8697
rect 654 8692 769 8693
rect 654 8688 659 8692
rect 663 8688 669 8692
rect 673 8688 679 8692
rect 683 8688 689 8692
rect 693 8688 769 8692
rect 654 8398 769 8688
rect 2755 8412 2760 9173
rect 2850 9175 2857 9176
rect 2850 9170 2851 9175
rect 2856 9170 2857 9175
rect 2850 9169 2857 9170
rect 2897 9172 2950 9177
rect 2974 9175 3008 9179
rect 2886 9168 2893 9169
rect 2886 9163 2887 9168
rect 2892 9163 2893 9168
rect 2897 9167 2898 9172
rect 2903 9167 2904 9172
rect 2945 9169 2950 9172
rect 2973 9174 3008 9175
rect 2973 9169 2974 9174
rect 2979 9169 2980 9174
rect 3002 9169 3003 9174
rect 3007 9169 3008 9174
rect 2897 9166 2904 9167
rect 2944 9168 2951 9169
rect 2973 9168 2980 9169
rect 2989 9168 2996 9169
rect 3002 9168 3008 9169
rect 3018 9169 3025 9170
rect 3044 9169 3051 9170
rect 3124 9169 3131 9170
rect 2886 9162 2893 9163
rect 2920 9163 2927 9164
rect 2920 9162 2921 9163
rect 2887 9158 2921 9162
rect 2926 9158 2927 9163
rect 2944 9163 2945 9168
rect 2950 9163 2951 9168
rect 2944 9162 2951 9163
rect 2959 9164 2966 9165
rect 2887 9157 2927 9158
rect 2959 9158 2960 9164
rect 2965 9159 2966 9164
rect 2989 9163 2990 9168
rect 2995 9163 2996 9168
rect 3018 9164 3019 9169
rect 3024 9164 3045 9169
rect 3050 9164 3051 9169
rect 3018 9163 3025 9164
rect 3044 9163 3051 9164
rect 3101 9164 3125 9169
rect 3130 9164 3131 9169
rect 2989 9162 2996 9163
rect 2990 9159 2995 9162
rect 2965 9158 2995 9159
rect 2959 9153 2995 9158
rect 3019 9136 3024 9163
rect 2850 9130 3024 9136
rect 2850 9107 2855 9130
rect 2887 9108 2927 9109
rect 2849 9106 2856 9107
rect 2849 9101 2850 9106
rect 2855 9101 2856 9106
rect 2887 9104 2921 9108
rect 2849 9100 2856 9101
rect 2886 9103 2893 9104
rect 2886 9098 2887 9103
rect 2892 9098 2893 9103
rect 2920 9103 2921 9104
rect 2926 9103 2927 9108
rect 2959 9108 2995 9113
rect 3101 9111 3106 9164
rect 3124 9163 3131 9164
rect 3182 9135 3187 9223
rect 3144 9130 3187 9135
rect 2920 9102 2927 9103
rect 2944 9103 2951 9104
rect 2886 9097 2893 9098
rect 2897 9099 2904 9100
rect 2897 9094 2898 9099
rect 2903 9094 2904 9099
rect 2944 9098 2945 9103
rect 2950 9098 2951 9103
rect 2959 9102 2960 9108
rect 2965 9107 2995 9108
rect 2965 9102 2966 9107
rect 2990 9104 2995 9107
rect 3100 9110 3107 9111
rect 3100 9105 3101 9110
rect 3106 9105 3107 9110
rect 3100 9104 3107 9105
rect 2959 9101 2966 9102
rect 2989 9103 2996 9104
rect 2989 9098 2990 9103
rect 2995 9098 2996 9103
rect 3018 9102 3025 9103
rect 2944 9097 2951 9098
rect 2973 9097 2980 9098
rect 2989 9097 2996 9098
rect 3002 9097 3008 9098
rect 2945 9094 2950 9097
rect 2897 9089 2950 9094
rect 2973 9092 2974 9097
rect 2979 9092 2980 9097
rect 3002 9092 3003 9097
rect 3007 9092 3008 9097
rect 2973 9091 3008 9092
rect 2974 9087 3008 9091
rect 3018 9097 3019 9102
rect 3024 9097 3025 9102
rect 3144 9097 3149 9130
rect 3207 9107 3214 9108
rect 3207 9102 3208 9107
rect 3213 9102 3214 9107
rect 3207 9101 3214 9102
rect 3018 9096 3025 9097
rect 3044 9096 3051 9097
rect 3018 9091 3045 9096
rect 3050 9091 3051 9096
rect 3144 9096 3156 9097
rect 3144 9091 3150 9096
rect 3155 9091 3156 9096
rect 3018 9070 3023 9091
rect 3044 9090 3051 9091
rect 3149 9090 3156 9091
rect 2851 9064 3023 9070
rect 2851 9044 2856 9064
rect 2850 9043 2857 9044
rect 2850 9038 2851 9043
rect 2856 9038 2857 9043
rect 2850 9037 2857 9038
rect 2897 9040 2950 9045
rect 2974 9043 3008 9047
rect 2886 9036 2893 9037
rect 2886 9031 2887 9036
rect 2892 9031 2893 9036
rect 2897 9035 2898 9040
rect 2903 9035 2904 9040
rect 2945 9037 2950 9040
rect 2973 9042 3008 9043
rect 2973 9037 2974 9042
rect 2979 9037 2980 9042
rect 3002 9037 3003 9042
rect 3007 9037 3008 9042
rect 3043 9038 3050 9039
rect 3149 9038 3156 9039
rect 2897 9034 2904 9035
rect 2944 9036 2951 9037
rect 2973 9036 2980 9037
rect 2989 9036 2996 9037
rect 3002 9036 3008 9037
rect 3018 9037 3044 9038
rect 2886 9030 2893 9031
rect 2920 9031 2927 9032
rect 2920 9030 2921 9031
rect 2887 9026 2921 9030
rect 2926 9026 2927 9031
rect 2944 9031 2945 9036
rect 2950 9031 2951 9036
rect 2944 9030 2951 9031
rect 2959 9032 2966 9033
rect 2887 9025 2927 9026
rect 2959 9026 2960 9032
rect 2965 9027 2966 9032
rect 2989 9031 2990 9036
rect 2995 9031 2996 9036
rect 2989 9030 2996 9031
rect 3018 9032 3019 9037
rect 3024 9033 3044 9037
rect 3049 9033 3050 9038
rect 3024 9032 3025 9033
rect 3043 9032 3050 9033
rect 3145 9033 3150 9038
rect 3155 9033 3156 9038
rect 3145 9032 3156 9033
rect 3018 9031 3025 9032
rect 2990 9027 2995 9030
rect 2965 9026 2995 9027
rect 2959 9021 2995 9026
rect 3018 9004 3023 9031
rect 2850 8998 3023 9004
rect 3145 9004 3150 9032
rect 3145 8999 3188 9004
rect 2850 8975 2855 8998
rect 2887 8976 2927 8977
rect 2849 8974 2856 8975
rect 2849 8969 2850 8974
rect 2855 8969 2856 8974
rect 2887 8972 2921 8976
rect 2849 8968 2856 8969
rect 2886 8971 2893 8972
rect 2886 8966 2887 8971
rect 2892 8966 2893 8971
rect 2920 8971 2921 8972
rect 2926 8971 2927 8976
rect 2959 8976 2995 8981
rect 3183 8980 3188 8999
rect 2920 8970 2927 8971
rect 2944 8971 2951 8972
rect 2886 8965 2893 8966
rect 2897 8967 2904 8968
rect 2897 8962 2898 8967
rect 2903 8962 2904 8967
rect 2944 8966 2945 8971
rect 2950 8966 2951 8971
rect 2959 8970 2960 8976
rect 2965 8975 2995 8976
rect 2965 8970 2966 8975
rect 2990 8972 2995 8975
rect 3182 8979 3189 8980
rect 3182 8974 3183 8979
rect 3188 8974 3189 8979
rect 3182 8973 3189 8974
rect 3208 8972 3213 9101
rect 3216 8972 3223 8973
rect 2959 8969 2966 8970
rect 2989 8971 2996 8972
rect 2989 8966 2990 8971
rect 2995 8966 2996 8971
rect 3018 8970 3025 8971
rect 2944 8965 2951 8966
rect 2973 8965 2980 8966
rect 2989 8965 2996 8966
rect 3002 8965 3008 8966
rect 2945 8962 2950 8965
rect 2897 8957 2950 8962
rect 2973 8960 2974 8965
rect 2979 8960 2980 8965
rect 3002 8960 3003 8965
rect 3007 8960 3008 8965
rect 2973 8959 3008 8960
rect 2974 8955 3008 8959
rect 3018 8965 3019 8970
rect 3024 8965 3025 8970
rect 3100 8970 3107 8971
rect 3100 8965 3101 8970
rect 3106 8965 3107 8970
rect 3196 8967 3217 8972
rect 3222 8967 3223 8972
rect 3196 8966 3208 8967
rect 3216 8966 3223 8967
rect 3018 8964 3025 8965
rect 3044 8964 3051 8965
rect 3100 8964 3107 8965
rect 3125 8964 3132 8965
rect 3018 8959 3045 8964
rect 3050 8959 3051 8964
rect 3101 8959 3126 8964
rect 3131 8959 3132 8964
rect 3018 8938 3023 8959
rect 3044 8958 3051 8959
rect 3125 8958 3132 8959
rect 3196 8958 3201 8966
rect 2851 8932 3023 8938
rect 3163 8937 3201 8958
rect 2851 8912 2856 8932
rect 2850 8911 2857 8912
rect 2850 8906 2851 8911
rect 2856 8906 2857 8911
rect 2850 8905 2857 8906
rect 2897 8908 2950 8913
rect 2974 8911 3008 8915
rect 2886 8904 2893 8905
rect 2886 8899 2887 8904
rect 2892 8899 2893 8904
rect 2897 8903 2898 8908
rect 2903 8903 2904 8908
rect 2945 8905 2950 8908
rect 2973 8910 3008 8911
rect 2973 8905 2974 8910
rect 2979 8905 2980 8910
rect 3002 8905 3003 8910
rect 3007 8905 3008 8910
rect 2897 8902 2904 8903
rect 2944 8904 2951 8905
rect 2973 8904 2980 8905
rect 2989 8904 2996 8905
rect 3002 8904 3008 8905
rect 3018 8905 3025 8906
rect 2886 8898 2893 8899
rect 2920 8899 2927 8900
rect 2920 8898 2921 8899
rect 2887 8894 2921 8898
rect 2926 8894 2927 8899
rect 2944 8899 2945 8904
rect 2950 8899 2951 8904
rect 2944 8898 2951 8899
rect 2959 8900 2966 8901
rect 2887 8893 2927 8894
rect 2959 8894 2960 8900
rect 2965 8895 2966 8900
rect 2989 8899 2990 8904
rect 2995 8899 2996 8904
rect 3018 8900 3019 8905
rect 3024 8903 3025 8905
rect 3044 8903 3051 8904
rect 3124 8903 3131 8904
rect 3024 8900 3045 8903
rect 3018 8899 3045 8900
rect 2989 8898 2996 8899
rect 3019 8898 3045 8899
rect 3050 8898 3051 8903
rect 2990 8895 2995 8898
rect 2965 8894 2995 8895
rect 2959 8889 2995 8894
rect 3019 8872 3024 8898
rect 3044 8897 3051 8898
rect 3101 8898 3125 8903
rect 3130 8898 3131 8903
rect 2850 8866 3024 8872
rect 2850 8843 2855 8866
rect 2887 8844 2927 8845
rect 2849 8842 2856 8843
rect 2849 8837 2850 8842
rect 2855 8837 2856 8842
rect 2887 8840 2921 8844
rect 2849 8836 2856 8837
rect 2886 8839 2893 8840
rect 2886 8834 2887 8839
rect 2892 8834 2893 8839
rect 2920 8839 2921 8840
rect 2926 8839 2927 8844
rect 2959 8844 2995 8849
rect 3101 8847 3106 8898
rect 3124 8897 3131 8898
rect 2920 8838 2927 8839
rect 2944 8839 2951 8840
rect 2886 8833 2893 8834
rect 2897 8835 2904 8836
rect 2897 8830 2898 8835
rect 2903 8830 2904 8835
rect 2944 8834 2945 8839
rect 2950 8834 2951 8839
rect 2959 8838 2960 8844
rect 2965 8843 2995 8844
rect 2965 8838 2966 8843
rect 2990 8840 2995 8843
rect 3100 8846 3107 8847
rect 3100 8841 3101 8846
rect 3106 8841 3107 8846
rect 3100 8840 3107 8841
rect 2959 8837 2966 8838
rect 2989 8839 2996 8840
rect 2989 8834 2990 8839
rect 2995 8834 2996 8839
rect 3018 8838 3025 8839
rect 2944 8833 2951 8834
rect 2973 8833 2980 8834
rect 2989 8833 2996 8834
rect 3002 8833 3008 8834
rect 2945 8830 2950 8833
rect 2897 8825 2950 8830
rect 2973 8828 2974 8833
rect 2979 8828 2980 8833
rect 3002 8828 3003 8833
rect 3007 8828 3008 8833
rect 2973 8827 3008 8828
rect 2974 8823 3008 8827
rect 3018 8833 3019 8838
rect 3024 8833 3025 8838
rect 3018 8832 3025 8833
rect 3044 8832 3051 8833
rect 3018 8827 3045 8832
rect 3050 8827 3051 8832
rect 3163 8828 3168 8937
rect 3213 8899 3220 8900
rect 3213 8894 3214 8899
rect 3219 8894 3220 8899
rect 3213 8893 3220 8894
rect 3120 8827 3168 8828
rect 3018 8806 3023 8827
rect 3044 8826 3051 8827
rect 2851 8800 3023 8806
rect 3089 8822 3168 8827
rect 3214 8831 3219 8893
rect 3214 8825 3281 8831
rect 2851 8780 2856 8800
rect 2850 8779 2857 8780
rect 2850 8774 2851 8779
rect 2856 8774 2857 8779
rect 2850 8773 2857 8774
rect 2897 8776 2950 8781
rect 2974 8779 3008 8783
rect 3089 8779 3094 8822
rect 2886 8772 2893 8773
rect 2886 8767 2887 8772
rect 2892 8767 2893 8772
rect 2897 8771 2898 8776
rect 2903 8771 2904 8776
rect 2945 8773 2950 8776
rect 2973 8778 3008 8779
rect 2973 8773 2974 8778
rect 2979 8773 2980 8778
rect 3002 8773 3003 8778
rect 3007 8773 3008 8778
rect 3088 8778 3095 8779
rect 2897 8770 2904 8771
rect 2944 8772 2951 8773
rect 2973 8772 2980 8773
rect 2989 8772 2996 8773
rect 3002 8772 3008 8773
rect 3018 8773 3025 8774
rect 2886 8766 2893 8767
rect 2920 8767 2927 8768
rect 2920 8766 2921 8767
rect 2887 8762 2921 8766
rect 2926 8762 2927 8767
rect 2944 8767 2945 8772
rect 2950 8767 2951 8772
rect 2944 8766 2951 8767
rect 2959 8768 2966 8769
rect 2887 8761 2927 8762
rect 2959 8762 2960 8768
rect 2965 8763 2966 8768
rect 2989 8767 2990 8772
rect 2995 8767 2996 8772
rect 3018 8768 3019 8773
rect 3024 8768 3025 8773
rect 3088 8773 3089 8778
rect 3094 8773 3095 8778
rect 3158 8776 3211 8781
rect 3235 8779 3269 8783
rect 3276 8779 3281 8825
rect 3088 8772 3095 8773
rect 3147 8772 3154 8773
rect 3018 8767 3025 8768
rect 3043 8767 3050 8768
rect 2989 8766 2996 8767
rect 2990 8763 2995 8766
rect 2965 8762 2995 8763
rect 2959 8757 2995 8762
rect 3020 8762 3044 8767
rect 3049 8762 3050 8767
rect 3147 8767 3148 8772
rect 3153 8767 3154 8772
rect 3158 8771 3159 8776
rect 3164 8771 3165 8776
rect 3206 8773 3211 8776
rect 3234 8778 3269 8779
rect 3234 8773 3235 8778
rect 3240 8773 3241 8778
rect 3263 8773 3264 8778
rect 3268 8773 3269 8778
rect 3158 8770 3165 8771
rect 3205 8772 3212 8773
rect 3234 8772 3241 8773
rect 3250 8772 3257 8773
rect 3263 8772 3269 8773
rect 3275 8778 3282 8779
rect 3275 8773 3276 8778
rect 3281 8773 3282 8778
rect 3275 8772 3282 8773
rect 3147 8766 3154 8767
rect 3181 8767 3188 8768
rect 3181 8766 3182 8767
rect 2755 8411 2761 8412
rect 2755 8407 2756 8411
rect 2760 8407 2761 8411
rect 2755 8406 2761 8407
rect 654 8394 659 8398
rect 663 8394 669 8398
rect 673 8394 679 8398
rect 683 8394 689 8398
rect 693 8394 769 8398
rect 654 8393 769 8394
rect 654 8389 659 8393
rect 663 8389 669 8393
rect 673 8389 679 8393
rect 683 8389 689 8393
rect 693 8389 769 8393
rect 654 8388 769 8389
rect 3020 8394 3025 8762
rect 3043 8761 3050 8762
rect 3148 8762 3182 8766
rect 3187 8762 3188 8767
rect 3205 8767 3206 8772
rect 3211 8767 3212 8772
rect 3205 8766 3212 8767
rect 3220 8768 3227 8769
rect 3148 8761 3188 8762
rect 3220 8762 3221 8768
rect 3226 8763 3227 8768
rect 3250 8767 3251 8772
rect 3256 8767 3257 8772
rect 3250 8766 3257 8767
rect 3251 8763 3256 8766
rect 3226 8762 3256 8763
rect 3220 8757 3256 8762
rect 3303 8734 3308 9261
rect 3832 9240 3872 9241
rect 3792 9238 3799 9239
rect 3770 9233 3799 9238
rect 3832 9236 3866 9240
rect 3567 9178 3573 9179
rect 3567 9174 3568 9178
rect 3572 9174 3705 9178
rect 3567 9173 3705 9174
rect 3559 9141 3566 9142
rect 3442 9140 3449 9141
rect 3442 9135 3443 9140
rect 3448 9135 3449 9140
rect 3559 9136 3560 9141
rect 3565 9136 3566 9141
rect 3559 9135 3566 9136
rect 3442 9134 3449 9135
rect 3443 8825 3448 9134
rect 3442 8824 3449 8825
rect 3560 8824 3565 9135
rect 3442 8819 3443 8824
rect 3448 8819 3449 8824
rect 3442 8818 3449 8819
rect 3559 8823 3566 8824
rect 3559 8818 3560 8823
rect 3565 8818 3566 8823
rect 3559 8817 3566 8818
rect 3311 8778 3317 8779
rect 3311 8774 3312 8778
rect 3316 8774 3317 8778
rect 3311 8773 3317 8774
rect 3150 8729 3308 8734
rect 3150 8667 3155 8729
rect 3149 8666 3155 8667
rect 3149 8662 3150 8666
rect 3154 8662 3155 8666
rect 3149 8661 3155 8662
rect 3312 8604 3317 8773
rect 3275 8599 3317 8604
rect 3275 8585 3280 8599
rect 3274 8584 3280 8585
rect 3274 8580 3275 8584
rect 3279 8580 3280 8584
rect 3274 8579 3280 8580
rect 3700 8412 3705 9173
rect 3700 8411 3706 8412
rect 3700 8407 3701 8411
rect 3705 8407 3706 8411
rect 3700 8406 3706 8407
rect 3770 8394 3775 9233
rect 3792 9232 3799 9233
rect 3831 9235 3838 9236
rect 3831 9230 3832 9235
rect 3837 9230 3838 9235
rect 3865 9235 3866 9236
rect 3871 9235 3872 9240
rect 3904 9240 3940 9245
rect 3865 9234 3872 9235
rect 3889 9235 3896 9236
rect 3831 9229 3838 9230
rect 3842 9231 3849 9232
rect 3842 9226 3843 9231
rect 3848 9226 3849 9231
rect 3889 9230 3890 9235
rect 3895 9230 3896 9235
rect 3904 9234 3905 9240
rect 3910 9239 3940 9240
rect 3910 9234 3911 9239
rect 3935 9236 3940 9239
rect 3904 9233 3911 9234
rect 3934 9235 3941 9236
rect 3934 9230 3935 9235
rect 3940 9230 3941 9235
rect 3963 9234 3970 9235
rect 3889 9229 3896 9230
rect 3918 9229 3925 9230
rect 3934 9229 3941 9230
rect 3947 9229 3953 9230
rect 3890 9226 3895 9229
rect 3842 9221 3895 9226
rect 3918 9224 3919 9229
rect 3924 9224 3925 9229
rect 3947 9224 3948 9229
rect 3952 9224 3953 9229
rect 3918 9223 3953 9224
rect 3919 9219 3953 9223
rect 3963 9229 3964 9234
rect 3969 9229 3970 9234
rect 4045 9234 4052 9235
rect 4045 9229 4046 9234
rect 4051 9229 4052 9234
rect 4130 9234 4137 9235
rect 4130 9229 4131 9234
rect 4136 9229 4137 9234
rect 3963 9228 3970 9229
rect 3989 9228 3996 9229
rect 4045 9228 4052 9229
rect 4070 9228 4077 9229
rect 4130 9228 4137 9229
rect 3963 9223 3990 9228
rect 3995 9223 3996 9228
rect 4046 9223 4071 9228
rect 4076 9223 4077 9228
rect 3963 9202 3968 9223
rect 3989 9222 3996 9223
rect 4070 9222 4077 9223
rect 4127 9223 4136 9228
rect 3796 9196 3968 9202
rect 3796 9176 3801 9196
rect 3795 9175 3802 9176
rect 3795 9170 3796 9175
rect 3801 9170 3802 9175
rect 3795 9169 3802 9170
rect 3842 9172 3895 9177
rect 3919 9175 3953 9179
rect 3831 9168 3838 9169
rect 3831 9163 3832 9168
rect 3837 9163 3838 9168
rect 3842 9167 3843 9172
rect 3848 9167 3849 9172
rect 3890 9169 3895 9172
rect 3918 9174 3953 9175
rect 3918 9169 3919 9174
rect 3924 9169 3925 9174
rect 3947 9169 3948 9174
rect 3952 9169 3953 9174
rect 3842 9166 3849 9167
rect 3889 9168 3896 9169
rect 3918 9168 3925 9169
rect 3934 9168 3941 9169
rect 3947 9168 3953 9169
rect 3963 9169 3970 9170
rect 3989 9169 3996 9170
rect 4069 9169 4076 9170
rect 3831 9162 3838 9163
rect 3865 9163 3872 9164
rect 3865 9162 3866 9163
rect 3832 9158 3866 9162
rect 3871 9158 3872 9163
rect 3889 9163 3890 9168
rect 3895 9163 3896 9168
rect 3889 9162 3896 9163
rect 3904 9164 3911 9165
rect 3832 9157 3872 9158
rect 3904 9158 3905 9164
rect 3910 9159 3911 9164
rect 3934 9163 3935 9168
rect 3940 9163 3941 9168
rect 3963 9164 3964 9169
rect 3969 9164 3990 9169
rect 3995 9164 3996 9169
rect 3963 9163 3970 9164
rect 3989 9163 3996 9164
rect 4046 9164 4070 9169
rect 4075 9164 4076 9169
rect 3934 9162 3941 9163
rect 3935 9159 3940 9162
rect 3910 9158 3940 9159
rect 3904 9153 3940 9158
rect 3964 9136 3969 9163
rect 3795 9130 3969 9136
rect 3795 9107 3800 9130
rect 3832 9108 3872 9109
rect 3794 9106 3801 9107
rect 3794 9101 3795 9106
rect 3800 9101 3801 9106
rect 3832 9104 3866 9108
rect 3794 9100 3801 9101
rect 3831 9103 3838 9104
rect 3831 9098 3832 9103
rect 3837 9098 3838 9103
rect 3865 9103 3866 9104
rect 3871 9103 3872 9108
rect 3904 9108 3940 9113
rect 4046 9111 4051 9164
rect 4069 9163 4076 9164
rect 4127 9135 4132 9223
rect 4089 9130 4132 9135
rect 3865 9102 3872 9103
rect 3889 9103 3896 9104
rect 3831 9097 3838 9098
rect 3842 9099 3849 9100
rect 3842 9094 3843 9099
rect 3848 9094 3849 9099
rect 3889 9098 3890 9103
rect 3895 9098 3896 9103
rect 3904 9102 3905 9108
rect 3910 9107 3940 9108
rect 3910 9102 3911 9107
rect 3935 9104 3940 9107
rect 4045 9110 4052 9111
rect 4045 9105 4046 9110
rect 4051 9105 4052 9110
rect 4045 9104 4052 9105
rect 3904 9101 3911 9102
rect 3934 9103 3941 9104
rect 3934 9098 3935 9103
rect 3940 9098 3941 9103
rect 3963 9102 3970 9103
rect 3889 9097 3896 9098
rect 3918 9097 3925 9098
rect 3934 9097 3941 9098
rect 3947 9097 3953 9098
rect 3890 9094 3895 9097
rect 3842 9089 3895 9094
rect 3918 9092 3919 9097
rect 3924 9092 3925 9097
rect 3947 9092 3948 9097
rect 3952 9092 3953 9097
rect 3918 9091 3953 9092
rect 3919 9087 3953 9091
rect 3963 9097 3964 9102
rect 3969 9097 3970 9102
rect 4089 9097 4094 9130
rect 4152 9107 4159 9108
rect 4152 9102 4153 9107
rect 4158 9102 4159 9107
rect 4152 9101 4159 9102
rect 3963 9096 3970 9097
rect 3989 9096 3996 9097
rect 3963 9091 3990 9096
rect 3995 9091 3996 9096
rect 4089 9096 4101 9097
rect 4089 9091 4095 9096
rect 4100 9091 4101 9096
rect 3963 9070 3968 9091
rect 3989 9090 3996 9091
rect 4094 9090 4101 9091
rect 3796 9064 3968 9070
rect 3796 9044 3801 9064
rect 3795 9043 3802 9044
rect 3795 9038 3796 9043
rect 3801 9038 3802 9043
rect 3795 9037 3802 9038
rect 3842 9040 3895 9045
rect 3919 9043 3953 9047
rect 3831 9036 3838 9037
rect 3831 9031 3832 9036
rect 3837 9031 3838 9036
rect 3842 9035 3843 9040
rect 3848 9035 3849 9040
rect 3890 9037 3895 9040
rect 3918 9042 3953 9043
rect 3918 9037 3919 9042
rect 3924 9037 3925 9042
rect 3947 9037 3948 9042
rect 3952 9037 3953 9042
rect 3988 9038 3995 9039
rect 4094 9038 4101 9039
rect 3842 9034 3849 9035
rect 3889 9036 3896 9037
rect 3918 9036 3925 9037
rect 3934 9036 3941 9037
rect 3947 9036 3953 9037
rect 3963 9037 3989 9038
rect 3831 9030 3838 9031
rect 3865 9031 3872 9032
rect 3865 9030 3866 9031
rect 3832 9026 3866 9030
rect 3871 9026 3872 9031
rect 3889 9031 3890 9036
rect 3895 9031 3896 9036
rect 3889 9030 3896 9031
rect 3904 9032 3911 9033
rect 3832 9025 3872 9026
rect 3904 9026 3905 9032
rect 3910 9027 3911 9032
rect 3934 9031 3935 9036
rect 3940 9031 3941 9036
rect 3934 9030 3941 9031
rect 3963 9032 3964 9037
rect 3969 9033 3989 9037
rect 3994 9033 3995 9038
rect 3969 9032 3970 9033
rect 3988 9032 3995 9033
rect 4090 9033 4095 9038
rect 4100 9033 4101 9038
rect 4090 9032 4101 9033
rect 3963 9031 3970 9032
rect 3935 9027 3940 9030
rect 3910 9026 3940 9027
rect 3904 9021 3940 9026
rect 3963 9004 3968 9031
rect 3795 8998 3968 9004
rect 4090 9004 4095 9032
rect 4090 8999 4133 9004
rect 3795 8975 3800 8998
rect 3832 8976 3872 8977
rect 3794 8974 3801 8975
rect 3794 8969 3795 8974
rect 3800 8969 3801 8974
rect 3832 8972 3866 8976
rect 3794 8968 3801 8969
rect 3831 8971 3838 8972
rect 3831 8966 3832 8971
rect 3837 8966 3838 8971
rect 3865 8971 3866 8972
rect 3871 8971 3872 8976
rect 3904 8976 3940 8981
rect 4128 8980 4133 8999
rect 3865 8970 3872 8971
rect 3889 8971 3896 8972
rect 3831 8965 3838 8966
rect 3842 8967 3849 8968
rect 3842 8962 3843 8967
rect 3848 8962 3849 8967
rect 3889 8966 3890 8971
rect 3895 8966 3896 8971
rect 3904 8970 3905 8976
rect 3910 8975 3940 8976
rect 3910 8970 3911 8975
rect 3935 8972 3940 8975
rect 4127 8979 4134 8980
rect 4127 8974 4128 8979
rect 4133 8974 4134 8979
rect 4127 8973 4134 8974
rect 4153 8972 4158 9101
rect 4161 8972 4168 8973
rect 3904 8969 3911 8970
rect 3934 8971 3941 8972
rect 3934 8966 3935 8971
rect 3940 8966 3941 8971
rect 3963 8970 3970 8971
rect 3889 8965 3896 8966
rect 3918 8965 3925 8966
rect 3934 8965 3941 8966
rect 3947 8965 3953 8966
rect 3890 8962 3895 8965
rect 3842 8957 3895 8962
rect 3918 8960 3919 8965
rect 3924 8960 3925 8965
rect 3947 8960 3948 8965
rect 3952 8960 3953 8965
rect 3918 8959 3953 8960
rect 3919 8955 3953 8959
rect 3963 8965 3964 8970
rect 3969 8965 3970 8970
rect 4045 8970 4052 8971
rect 4045 8965 4046 8970
rect 4051 8965 4052 8970
rect 4141 8967 4162 8972
rect 4167 8967 4168 8972
rect 4141 8966 4153 8967
rect 4161 8966 4168 8967
rect 3963 8964 3970 8965
rect 3989 8964 3996 8965
rect 4045 8964 4052 8965
rect 4070 8964 4077 8965
rect 3963 8959 3990 8964
rect 3995 8959 3996 8964
rect 4046 8959 4071 8964
rect 4076 8959 4077 8964
rect 3963 8938 3968 8959
rect 3989 8958 3996 8959
rect 4070 8958 4077 8959
rect 4141 8958 4146 8966
rect 3796 8932 3968 8938
rect 4108 8937 4146 8958
rect 3796 8912 3801 8932
rect 3795 8911 3802 8912
rect 3795 8906 3796 8911
rect 3801 8906 3802 8911
rect 3795 8905 3802 8906
rect 3842 8908 3895 8913
rect 3919 8911 3953 8915
rect 3831 8904 3838 8905
rect 3831 8899 3832 8904
rect 3837 8899 3838 8904
rect 3842 8903 3843 8908
rect 3848 8903 3849 8908
rect 3890 8905 3895 8908
rect 3918 8910 3953 8911
rect 3918 8905 3919 8910
rect 3924 8905 3925 8910
rect 3947 8905 3948 8910
rect 3952 8905 3953 8910
rect 3842 8902 3849 8903
rect 3889 8904 3896 8905
rect 3918 8904 3925 8905
rect 3934 8904 3941 8905
rect 3947 8904 3953 8905
rect 3963 8905 3970 8906
rect 3831 8898 3838 8899
rect 3865 8899 3872 8900
rect 3865 8898 3866 8899
rect 3832 8894 3866 8898
rect 3871 8894 3872 8899
rect 3889 8899 3890 8904
rect 3895 8899 3896 8904
rect 3889 8898 3896 8899
rect 3904 8900 3911 8901
rect 3832 8893 3872 8894
rect 3904 8894 3905 8900
rect 3910 8895 3911 8900
rect 3934 8899 3935 8904
rect 3940 8899 3941 8904
rect 3963 8900 3964 8905
rect 3969 8903 3970 8905
rect 3989 8903 3996 8904
rect 4069 8903 4076 8904
rect 3969 8900 3990 8903
rect 3963 8899 3990 8900
rect 3934 8898 3941 8899
rect 3964 8898 3990 8899
rect 3995 8898 3996 8903
rect 3935 8895 3940 8898
rect 3910 8894 3940 8895
rect 3904 8889 3940 8894
rect 3964 8872 3969 8898
rect 3989 8897 3996 8898
rect 4046 8898 4070 8903
rect 4075 8898 4076 8903
rect 3795 8866 3969 8872
rect 3795 8843 3800 8866
rect 3832 8844 3872 8845
rect 3794 8842 3801 8843
rect 3794 8837 3795 8842
rect 3800 8837 3801 8842
rect 3832 8840 3866 8844
rect 3794 8836 3801 8837
rect 3831 8839 3838 8840
rect 3831 8834 3832 8839
rect 3837 8834 3838 8839
rect 3865 8839 3866 8840
rect 3871 8839 3872 8844
rect 3904 8844 3940 8849
rect 4046 8847 4051 8898
rect 4069 8897 4076 8898
rect 3865 8838 3872 8839
rect 3889 8839 3896 8840
rect 3831 8833 3838 8834
rect 3842 8835 3849 8836
rect 3842 8830 3843 8835
rect 3848 8830 3849 8835
rect 3889 8834 3890 8839
rect 3895 8834 3896 8839
rect 3904 8838 3905 8844
rect 3910 8843 3940 8844
rect 3910 8838 3911 8843
rect 3935 8840 3940 8843
rect 4045 8846 4052 8847
rect 4045 8841 4046 8846
rect 4051 8841 4052 8846
rect 4045 8840 4052 8841
rect 3904 8837 3911 8838
rect 3934 8839 3941 8840
rect 3934 8834 3935 8839
rect 3940 8834 3941 8839
rect 3963 8838 3970 8839
rect 3889 8833 3896 8834
rect 3918 8833 3925 8834
rect 3934 8833 3941 8834
rect 3947 8833 3953 8834
rect 3890 8830 3895 8833
rect 3842 8825 3895 8830
rect 3918 8828 3919 8833
rect 3924 8828 3925 8833
rect 3947 8828 3948 8833
rect 3952 8828 3953 8833
rect 3918 8827 3953 8828
rect 3919 8823 3953 8827
rect 3963 8833 3964 8838
rect 3969 8833 3970 8838
rect 3963 8832 3970 8833
rect 3989 8832 3996 8833
rect 3963 8827 3990 8832
rect 3995 8827 3996 8832
rect 4108 8828 4113 8937
rect 4158 8899 4165 8900
rect 4158 8894 4159 8899
rect 4164 8894 4165 8899
rect 4158 8893 4165 8894
rect 4065 8827 4113 8828
rect 3963 8806 3968 8827
rect 3989 8826 3996 8827
rect 3796 8800 3968 8806
rect 4034 8822 4113 8827
rect 4159 8831 4164 8893
rect 4159 8825 4226 8831
rect 3796 8780 3801 8800
rect 3795 8779 3802 8780
rect 3795 8774 3796 8779
rect 3801 8774 3802 8779
rect 3795 8773 3802 8774
rect 3842 8776 3895 8781
rect 3919 8779 3953 8783
rect 4034 8779 4039 8822
rect 3831 8772 3838 8773
rect 3831 8767 3832 8772
rect 3837 8767 3838 8772
rect 3842 8771 3843 8776
rect 3848 8771 3849 8776
rect 3890 8773 3895 8776
rect 3918 8778 3953 8779
rect 3918 8773 3919 8778
rect 3924 8773 3925 8778
rect 3947 8773 3948 8778
rect 3952 8773 3953 8778
rect 4033 8778 4040 8779
rect 3842 8770 3849 8771
rect 3889 8772 3896 8773
rect 3918 8772 3925 8773
rect 3934 8772 3941 8773
rect 3947 8772 3953 8773
rect 3963 8773 3970 8774
rect 3831 8766 3838 8767
rect 3865 8767 3872 8768
rect 3865 8766 3866 8767
rect 3832 8762 3866 8766
rect 3871 8762 3872 8767
rect 3889 8767 3890 8772
rect 3895 8767 3896 8772
rect 3889 8766 3896 8767
rect 3904 8768 3911 8769
rect 3832 8761 3872 8762
rect 3904 8762 3905 8768
rect 3910 8763 3911 8768
rect 3934 8767 3935 8772
rect 3940 8767 3941 8772
rect 3963 8768 3964 8773
rect 3969 8768 3970 8773
rect 4033 8773 4034 8778
rect 4039 8773 4040 8778
rect 4103 8776 4156 8781
rect 4180 8779 4214 8783
rect 4221 8779 4226 8825
rect 4033 8772 4040 8773
rect 4092 8772 4099 8773
rect 3963 8767 3970 8768
rect 3988 8767 3995 8768
rect 3934 8766 3941 8767
rect 3935 8763 3940 8766
rect 3910 8762 3940 8763
rect 3904 8757 3940 8762
rect 3965 8762 3989 8767
rect 3994 8762 3995 8767
rect 4092 8767 4093 8772
rect 4098 8767 4099 8772
rect 4103 8771 4104 8776
rect 4109 8771 4110 8776
rect 4151 8773 4156 8776
rect 4179 8778 4214 8779
rect 4179 8773 4180 8778
rect 4185 8773 4186 8778
rect 4208 8773 4209 8778
rect 4213 8773 4214 8778
rect 4103 8770 4110 8771
rect 4150 8772 4157 8773
rect 4179 8772 4186 8773
rect 4195 8772 4202 8773
rect 4208 8772 4214 8773
rect 4220 8778 4227 8779
rect 4220 8773 4221 8778
rect 4226 8773 4227 8778
rect 4220 8772 4227 8773
rect 4092 8766 4099 8767
rect 4126 8767 4133 8768
rect 4126 8766 4127 8767
rect 3965 8631 3970 8762
rect 3988 8761 3995 8762
rect 4093 8762 4127 8766
rect 4132 8762 4133 8767
rect 4150 8767 4151 8772
rect 4156 8767 4157 8772
rect 4150 8766 4157 8767
rect 4165 8768 4172 8769
rect 4093 8761 4133 8762
rect 4165 8762 4166 8768
rect 4171 8763 4172 8768
rect 4195 8767 4196 8772
rect 4201 8767 4202 8772
rect 4195 8766 4202 8767
rect 4196 8763 4201 8766
rect 4171 8762 4201 8763
rect 4165 8757 4201 8762
rect 4248 8734 4253 9261
rect 4095 8729 4253 8734
rect 4403 9060 4518 9442
rect 4403 9056 4479 9060
rect 4483 9056 4489 9060
rect 4493 9056 4499 9060
rect 4503 9056 4509 9060
rect 4513 9056 4518 9060
rect 4403 9055 4518 9056
rect 4403 9051 4479 9055
rect 4483 9051 4489 9055
rect 4493 9051 4499 9055
rect 4503 9051 4509 9055
rect 4513 9051 4518 9055
rect 4403 9050 4518 9051
rect 4403 9046 4479 9050
rect 4483 9046 4489 9050
rect 4493 9046 4499 9050
rect 4503 9046 4509 9050
rect 4513 9046 4518 9050
rect 4403 9045 4518 9046
rect 4403 9041 4479 9045
rect 4483 9041 4489 9045
rect 4493 9041 4499 9045
rect 4503 9041 4509 9045
rect 4513 9041 4518 9045
rect 4403 8751 4518 9041
rect 4403 8747 4479 8751
rect 4483 8747 4489 8751
rect 4493 8747 4499 8751
rect 4503 8747 4509 8751
rect 4513 8747 4518 8751
rect 4403 8746 4518 8747
rect 4403 8742 4479 8746
rect 4483 8742 4489 8746
rect 4493 8742 4499 8746
rect 4503 8742 4509 8746
rect 4513 8742 4518 8746
rect 4403 8741 4518 8742
rect 4403 8737 4479 8741
rect 4483 8737 4489 8741
rect 4493 8737 4499 8741
rect 4503 8737 4509 8741
rect 4513 8737 4518 8741
rect 4403 8736 4518 8737
rect 4403 8732 4479 8736
rect 4483 8732 4489 8736
rect 4493 8732 4499 8736
rect 4503 8732 4509 8736
rect 4513 8732 4518 8736
rect 4095 8667 4100 8729
rect 4094 8666 4100 8667
rect 4094 8662 4095 8666
rect 4099 8662 4100 8666
rect 4094 8661 4100 8662
rect 3965 8625 4276 8631
rect 4219 8584 4225 8585
rect 4219 8580 4220 8584
rect 4224 8580 4225 8584
rect 4219 8579 4225 8580
rect 3020 8388 3775 8394
rect 654 8384 659 8388
rect 663 8384 669 8388
rect 673 8384 679 8388
rect 683 8384 689 8388
rect 693 8384 769 8388
rect 654 8383 769 8384
rect 654 8379 659 8383
rect 663 8379 669 8383
rect 673 8379 679 8383
rect 683 8379 689 8383
rect 693 8379 769 8383
rect 654 8089 769 8379
rect 4220 8375 4225 8579
rect 654 8085 659 8089
rect 663 8085 669 8089
rect 673 8085 679 8089
rect 683 8085 689 8089
rect 693 8085 769 8089
rect 654 8084 769 8085
rect 654 8080 659 8084
rect 663 8080 669 8084
rect 673 8080 679 8084
rect 683 8080 689 8084
rect 693 8080 769 8084
rect 654 8079 769 8080
rect 654 8075 659 8079
rect 663 8075 669 8079
rect 673 8075 679 8079
rect 683 8075 689 8079
rect 693 8075 769 8079
rect 654 8074 769 8075
rect 654 8070 659 8074
rect 663 8070 669 8074
rect 673 8070 679 8074
rect 683 8070 689 8074
rect 693 8070 769 8074
rect 654 7780 769 8070
rect 2367 8370 4225 8375
rect 2367 7797 2372 8370
rect 2761 8335 2852 8336
rect 2761 8331 2847 8335
rect 2851 8331 2852 8335
rect 2762 8300 2767 8331
rect 2846 8330 2852 8331
rect 3791 8335 3797 8336
rect 3791 8331 3792 8335
rect 3796 8331 3797 8335
rect 3791 8330 3797 8331
rect 2623 8299 2767 8300
rect 2623 8295 2624 8299
rect 2628 8295 2767 8299
rect 3568 8300 3574 8301
rect 3791 8300 3796 8330
rect 2623 8294 2629 8295
rect 2849 8292 3329 8297
rect 3568 8296 3569 8300
rect 3573 8296 3796 8300
rect 4271 8297 4276 8625
rect 3568 8295 3796 8296
rect 3934 8292 4276 8297
rect 4403 8442 4518 8732
rect 4403 8438 4479 8442
rect 4483 8438 4489 8442
rect 4493 8438 4499 8442
rect 4503 8438 4509 8442
rect 4513 8438 4518 8442
rect 4403 8437 4518 8438
rect 4403 8433 4479 8437
rect 4483 8433 4489 8437
rect 4493 8433 4499 8437
rect 4503 8433 4509 8437
rect 4513 8433 4518 8437
rect 4403 8432 4518 8433
rect 4403 8428 4479 8432
rect 4483 8428 4489 8432
rect 4493 8428 4499 8432
rect 4503 8428 4509 8432
rect 4513 8428 4518 8432
rect 4403 8427 4518 8428
rect 4403 8423 4479 8427
rect 4483 8423 4489 8427
rect 4493 8423 4499 8427
rect 4503 8423 4509 8427
rect 4513 8423 4518 8427
rect 2849 8257 2854 8292
rect 3324 8287 3962 8292
rect 3302 8284 3308 8285
rect 3302 8280 3303 8284
rect 3307 8280 3308 8284
rect 3302 8279 3308 8280
rect 4247 8284 4253 8285
rect 4247 8280 4248 8284
rect 4252 8280 4253 8284
rect 4247 8279 4253 8280
rect 2887 8258 2927 8259
rect 2848 8250 2855 8257
rect 2887 8254 2921 8258
rect 2886 8253 2893 8254
rect 2886 8248 2887 8253
rect 2892 8248 2893 8253
rect 2920 8253 2921 8254
rect 2926 8253 2927 8258
rect 2959 8258 2995 8263
rect 2920 8252 2927 8253
rect 2944 8253 2951 8254
rect 2886 8247 2893 8248
rect 2897 8249 2904 8250
rect 2897 8244 2898 8249
rect 2903 8244 2904 8249
rect 2944 8248 2945 8253
rect 2950 8248 2951 8253
rect 2959 8252 2960 8258
rect 2965 8257 2995 8258
rect 2965 8252 2966 8257
rect 2990 8254 2995 8257
rect 2959 8251 2966 8252
rect 2989 8253 2996 8254
rect 2989 8248 2990 8253
rect 2995 8248 2996 8253
rect 3018 8252 3025 8253
rect 2944 8247 2951 8248
rect 2973 8247 2980 8248
rect 2989 8247 2996 8248
rect 3002 8247 3008 8248
rect 2945 8244 2950 8247
rect 2897 8239 2950 8244
rect 2973 8242 2974 8247
rect 2979 8242 2980 8247
rect 3002 8242 3003 8247
rect 3007 8242 3008 8247
rect 2973 8241 3008 8242
rect 2974 8237 3008 8241
rect 3018 8247 3019 8252
rect 3024 8247 3025 8252
rect 3100 8252 3107 8253
rect 3100 8247 3101 8252
rect 3106 8247 3107 8252
rect 3185 8252 3192 8253
rect 3185 8247 3186 8252
rect 3191 8247 3192 8252
rect 3018 8246 3025 8247
rect 3044 8246 3051 8247
rect 3100 8246 3107 8247
rect 3125 8246 3132 8247
rect 3185 8246 3192 8247
rect 3018 8241 3045 8246
rect 3050 8241 3051 8246
rect 3101 8241 3126 8246
rect 3131 8241 3132 8246
rect 3018 8220 3023 8241
rect 3044 8240 3051 8241
rect 3125 8240 3132 8241
rect 3182 8241 3191 8246
rect 2851 8214 3023 8220
rect 2622 8196 2628 8197
rect 2622 8192 2623 8196
rect 2627 8192 2760 8196
rect 2851 8194 2856 8214
rect 2622 8191 2760 8192
rect 2366 7796 2372 7797
rect 2366 7792 2367 7796
rect 2371 7792 2372 7796
rect 2366 7791 2372 7792
rect 654 7776 659 7780
rect 663 7776 669 7780
rect 673 7776 679 7780
rect 683 7776 689 7780
rect 693 7776 769 7780
rect 654 7775 769 7776
rect 654 7771 659 7775
rect 663 7771 669 7775
rect 673 7771 679 7775
rect 683 7771 689 7775
rect 693 7771 769 7775
rect 654 7770 769 7771
rect 654 7766 659 7770
rect 663 7766 669 7770
rect 673 7766 679 7770
rect 683 7766 689 7770
rect 693 7766 769 7770
rect 654 7765 769 7766
rect 654 7761 659 7765
rect 663 7761 669 7765
rect 673 7761 679 7765
rect 683 7761 689 7765
rect 693 7761 769 7765
rect 654 7471 769 7761
rect 654 7467 659 7471
rect 663 7467 669 7471
rect 673 7467 679 7471
rect 683 7467 689 7471
rect 693 7467 769 7471
rect 654 7466 769 7467
rect 654 7462 659 7466
rect 663 7462 669 7466
rect 673 7462 679 7466
rect 683 7462 689 7466
rect 693 7462 769 7466
rect 654 7461 769 7462
rect 654 7457 659 7461
rect 663 7457 669 7461
rect 673 7457 679 7461
rect 683 7457 689 7461
rect 693 7457 769 7461
rect 654 7456 769 7457
rect 654 7452 659 7456
rect 663 7452 669 7456
rect 673 7452 679 7456
rect 683 7452 689 7456
rect 693 7452 769 7456
rect 654 7162 769 7452
rect 2755 7430 2760 8191
rect 2850 8193 2857 8194
rect 2850 8188 2851 8193
rect 2856 8188 2857 8193
rect 2850 8187 2857 8188
rect 2897 8190 2950 8195
rect 2974 8193 3008 8197
rect 2886 8186 2893 8187
rect 2886 8181 2887 8186
rect 2892 8181 2893 8186
rect 2897 8185 2898 8190
rect 2903 8185 2904 8190
rect 2945 8187 2950 8190
rect 2973 8192 3008 8193
rect 2973 8187 2974 8192
rect 2979 8187 2980 8192
rect 3002 8187 3003 8192
rect 3007 8187 3008 8192
rect 2897 8184 2904 8185
rect 2944 8186 2951 8187
rect 2973 8186 2980 8187
rect 2989 8186 2996 8187
rect 3002 8186 3008 8187
rect 3018 8187 3025 8188
rect 3044 8187 3051 8188
rect 3124 8187 3131 8188
rect 2886 8180 2893 8181
rect 2920 8181 2927 8182
rect 2920 8180 2921 8181
rect 2887 8176 2921 8180
rect 2926 8176 2927 8181
rect 2944 8181 2945 8186
rect 2950 8181 2951 8186
rect 2944 8180 2951 8181
rect 2959 8182 2966 8183
rect 2887 8175 2927 8176
rect 2959 8176 2960 8182
rect 2965 8177 2966 8182
rect 2989 8181 2990 8186
rect 2995 8181 2996 8186
rect 3018 8182 3019 8187
rect 3024 8182 3045 8187
rect 3050 8182 3051 8187
rect 3018 8181 3025 8182
rect 3044 8181 3051 8182
rect 3101 8182 3125 8187
rect 3130 8182 3131 8187
rect 2989 8180 2996 8181
rect 2990 8177 2995 8180
rect 2965 8176 2995 8177
rect 2959 8171 2995 8176
rect 3019 8154 3024 8181
rect 2850 8148 3024 8154
rect 2850 8125 2855 8148
rect 2887 8126 2927 8127
rect 2849 8124 2856 8125
rect 2849 8119 2850 8124
rect 2855 8119 2856 8124
rect 2887 8122 2921 8126
rect 2849 8118 2856 8119
rect 2886 8121 2893 8122
rect 2886 8116 2887 8121
rect 2892 8116 2893 8121
rect 2920 8121 2921 8122
rect 2926 8121 2927 8126
rect 2959 8126 2995 8131
rect 3101 8129 3106 8182
rect 3124 8181 3131 8182
rect 3182 8153 3187 8241
rect 3144 8148 3187 8153
rect 2920 8120 2927 8121
rect 2944 8121 2951 8122
rect 2886 8115 2893 8116
rect 2897 8117 2904 8118
rect 2897 8112 2898 8117
rect 2903 8112 2904 8117
rect 2944 8116 2945 8121
rect 2950 8116 2951 8121
rect 2959 8120 2960 8126
rect 2965 8125 2995 8126
rect 2965 8120 2966 8125
rect 2990 8122 2995 8125
rect 3100 8128 3107 8129
rect 3100 8123 3101 8128
rect 3106 8123 3107 8128
rect 3100 8122 3107 8123
rect 2959 8119 2966 8120
rect 2989 8121 2996 8122
rect 2989 8116 2990 8121
rect 2995 8116 2996 8121
rect 3018 8120 3025 8121
rect 2944 8115 2951 8116
rect 2973 8115 2980 8116
rect 2989 8115 2996 8116
rect 3002 8115 3008 8116
rect 2945 8112 2950 8115
rect 2897 8107 2950 8112
rect 2973 8110 2974 8115
rect 2979 8110 2980 8115
rect 3002 8110 3003 8115
rect 3007 8110 3008 8115
rect 2973 8109 3008 8110
rect 2974 8105 3008 8109
rect 3018 8115 3019 8120
rect 3024 8115 3025 8120
rect 3144 8115 3149 8148
rect 3207 8125 3214 8126
rect 3207 8120 3208 8125
rect 3213 8120 3214 8125
rect 3207 8119 3214 8120
rect 3018 8114 3025 8115
rect 3044 8114 3051 8115
rect 3018 8109 3045 8114
rect 3050 8109 3051 8114
rect 3144 8114 3156 8115
rect 3144 8109 3150 8114
rect 3155 8109 3156 8114
rect 3018 8088 3023 8109
rect 3044 8108 3051 8109
rect 3149 8108 3156 8109
rect 2851 8082 3023 8088
rect 2851 8062 2856 8082
rect 2850 8061 2857 8062
rect 2850 8056 2851 8061
rect 2856 8056 2857 8061
rect 2850 8055 2857 8056
rect 2897 8058 2950 8063
rect 2974 8061 3008 8065
rect 2886 8054 2893 8055
rect 2886 8049 2887 8054
rect 2892 8049 2893 8054
rect 2897 8053 2898 8058
rect 2903 8053 2904 8058
rect 2945 8055 2950 8058
rect 2973 8060 3008 8061
rect 2973 8055 2974 8060
rect 2979 8055 2980 8060
rect 3002 8055 3003 8060
rect 3007 8055 3008 8060
rect 3043 8056 3050 8057
rect 3149 8056 3156 8057
rect 2897 8052 2904 8053
rect 2944 8054 2951 8055
rect 2973 8054 2980 8055
rect 2989 8054 2996 8055
rect 3002 8054 3008 8055
rect 3018 8055 3044 8056
rect 2886 8048 2893 8049
rect 2920 8049 2927 8050
rect 2920 8048 2921 8049
rect 2887 8044 2921 8048
rect 2926 8044 2927 8049
rect 2944 8049 2945 8054
rect 2950 8049 2951 8054
rect 2944 8048 2951 8049
rect 2959 8050 2966 8051
rect 2887 8043 2927 8044
rect 2959 8044 2960 8050
rect 2965 8045 2966 8050
rect 2989 8049 2990 8054
rect 2995 8049 2996 8054
rect 2989 8048 2996 8049
rect 3018 8050 3019 8055
rect 3024 8051 3044 8055
rect 3049 8051 3050 8056
rect 3024 8050 3025 8051
rect 3043 8050 3050 8051
rect 3145 8051 3150 8056
rect 3155 8051 3156 8056
rect 3145 8050 3156 8051
rect 3018 8049 3025 8050
rect 2990 8045 2995 8048
rect 2965 8044 2995 8045
rect 2959 8039 2995 8044
rect 3018 8022 3023 8049
rect 2850 8016 3023 8022
rect 3145 8022 3150 8050
rect 3145 8017 3188 8022
rect 2850 7993 2855 8016
rect 2887 7994 2927 7995
rect 2849 7992 2856 7993
rect 2849 7987 2850 7992
rect 2855 7987 2856 7992
rect 2887 7990 2921 7994
rect 2849 7986 2856 7987
rect 2886 7989 2893 7990
rect 2886 7984 2887 7989
rect 2892 7984 2893 7989
rect 2920 7989 2921 7990
rect 2926 7989 2927 7994
rect 2959 7994 2995 7999
rect 3183 7998 3188 8017
rect 2920 7988 2927 7989
rect 2944 7989 2951 7990
rect 2886 7983 2893 7984
rect 2897 7985 2904 7986
rect 2897 7980 2898 7985
rect 2903 7980 2904 7985
rect 2944 7984 2945 7989
rect 2950 7984 2951 7989
rect 2959 7988 2960 7994
rect 2965 7993 2995 7994
rect 2965 7988 2966 7993
rect 2990 7990 2995 7993
rect 3182 7997 3189 7998
rect 3182 7992 3183 7997
rect 3188 7992 3189 7997
rect 3182 7991 3189 7992
rect 3208 7990 3213 8119
rect 3216 7990 3223 7991
rect 2959 7987 2966 7988
rect 2989 7989 2996 7990
rect 2989 7984 2990 7989
rect 2995 7984 2996 7989
rect 3018 7988 3025 7989
rect 2944 7983 2951 7984
rect 2973 7983 2980 7984
rect 2989 7983 2996 7984
rect 3002 7983 3008 7984
rect 2945 7980 2950 7983
rect 2897 7975 2950 7980
rect 2973 7978 2974 7983
rect 2979 7978 2980 7983
rect 3002 7978 3003 7983
rect 3007 7978 3008 7983
rect 2973 7977 3008 7978
rect 2974 7973 3008 7977
rect 3018 7983 3019 7988
rect 3024 7983 3025 7988
rect 3100 7988 3107 7989
rect 3100 7983 3101 7988
rect 3106 7983 3107 7988
rect 3196 7985 3217 7990
rect 3222 7985 3223 7990
rect 3196 7984 3208 7985
rect 3216 7984 3223 7985
rect 3018 7982 3025 7983
rect 3044 7982 3051 7983
rect 3100 7982 3107 7983
rect 3125 7982 3132 7983
rect 3018 7977 3045 7982
rect 3050 7977 3051 7982
rect 3101 7977 3126 7982
rect 3131 7977 3132 7982
rect 3018 7956 3023 7977
rect 3044 7976 3051 7977
rect 3125 7976 3132 7977
rect 3196 7976 3201 7984
rect 2851 7950 3023 7956
rect 3163 7955 3201 7976
rect 2851 7930 2856 7950
rect 2850 7929 2857 7930
rect 2850 7924 2851 7929
rect 2856 7924 2857 7929
rect 2850 7923 2857 7924
rect 2897 7926 2950 7931
rect 2974 7929 3008 7933
rect 2886 7922 2893 7923
rect 2886 7917 2887 7922
rect 2892 7917 2893 7922
rect 2897 7921 2898 7926
rect 2903 7921 2904 7926
rect 2945 7923 2950 7926
rect 2973 7928 3008 7929
rect 2973 7923 2974 7928
rect 2979 7923 2980 7928
rect 3002 7923 3003 7928
rect 3007 7923 3008 7928
rect 2897 7920 2904 7921
rect 2944 7922 2951 7923
rect 2973 7922 2980 7923
rect 2989 7922 2996 7923
rect 3002 7922 3008 7923
rect 3018 7923 3025 7924
rect 2886 7916 2893 7917
rect 2920 7917 2927 7918
rect 2920 7916 2921 7917
rect 2887 7912 2921 7916
rect 2926 7912 2927 7917
rect 2944 7917 2945 7922
rect 2950 7917 2951 7922
rect 2944 7916 2951 7917
rect 2959 7918 2966 7919
rect 2887 7911 2927 7912
rect 2959 7912 2960 7918
rect 2965 7913 2966 7918
rect 2989 7917 2990 7922
rect 2995 7917 2996 7922
rect 3018 7918 3019 7923
rect 3024 7921 3025 7923
rect 3044 7921 3051 7922
rect 3124 7921 3131 7922
rect 3024 7918 3045 7921
rect 3018 7917 3045 7918
rect 2989 7916 2996 7917
rect 3019 7916 3045 7917
rect 3050 7916 3051 7921
rect 2990 7913 2995 7916
rect 2965 7912 2995 7913
rect 2959 7907 2995 7912
rect 3019 7890 3024 7916
rect 3044 7915 3051 7916
rect 3101 7916 3125 7921
rect 3130 7916 3131 7921
rect 2850 7884 3024 7890
rect 2850 7861 2855 7884
rect 2887 7862 2927 7863
rect 2849 7860 2856 7861
rect 2849 7855 2850 7860
rect 2855 7855 2856 7860
rect 2887 7858 2921 7862
rect 2849 7854 2856 7855
rect 2886 7857 2893 7858
rect 2886 7852 2887 7857
rect 2892 7852 2893 7857
rect 2920 7857 2921 7858
rect 2926 7857 2927 7862
rect 2959 7862 2995 7867
rect 3101 7865 3106 7916
rect 3124 7915 3131 7916
rect 2920 7856 2927 7857
rect 2944 7857 2951 7858
rect 2886 7851 2893 7852
rect 2897 7853 2904 7854
rect 2897 7848 2898 7853
rect 2903 7848 2904 7853
rect 2944 7852 2945 7857
rect 2950 7852 2951 7857
rect 2959 7856 2960 7862
rect 2965 7861 2995 7862
rect 2965 7856 2966 7861
rect 2990 7858 2995 7861
rect 3100 7864 3107 7865
rect 3100 7859 3101 7864
rect 3106 7859 3107 7864
rect 3100 7858 3107 7859
rect 2959 7855 2966 7856
rect 2989 7857 2996 7858
rect 2989 7852 2990 7857
rect 2995 7852 2996 7857
rect 3018 7856 3025 7857
rect 2944 7851 2951 7852
rect 2973 7851 2980 7852
rect 2989 7851 2996 7852
rect 3002 7851 3008 7852
rect 2945 7848 2950 7851
rect 2897 7843 2950 7848
rect 2973 7846 2974 7851
rect 2979 7846 2980 7851
rect 3002 7846 3003 7851
rect 3007 7846 3008 7851
rect 2973 7845 3008 7846
rect 2974 7841 3008 7845
rect 3018 7851 3019 7856
rect 3024 7851 3025 7856
rect 3018 7850 3025 7851
rect 3044 7850 3051 7851
rect 3018 7845 3045 7850
rect 3050 7845 3051 7850
rect 3163 7846 3168 7955
rect 3213 7917 3220 7918
rect 3213 7912 3214 7917
rect 3219 7912 3220 7917
rect 3213 7911 3220 7912
rect 3120 7845 3168 7846
rect 3018 7824 3023 7845
rect 3044 7844 3051 7845
rect 2851 7818 3023 7824
rect 3089 7840 3168 7845
rect 3214 7849 3219 7911
rect 3214 7843 3281 7849
rect 2851 7798 2856 7818
rect 2850 7797 2857 7798
rect 2850 7792 2851 7797
rect 2856 7792 2857 7797
rect 2850 7791 2857 7792
rect 2897 7794 2950 7799
rect 2974 7797 3008 7801
rect 3089 7797 3094 7840
rect 2886 7790 2893 7791
rect 2886 7785 2887 7790
rect 2892 7785 2893 7790
rect 2897 7789 2898 7794
rect 2903 7789 2904 7794
rect 2945 7791 2950 7794
rect 2973 7796 3008 7797
rect 2973 7791 2974 7796
rect 2979 7791 2980 7796
rect 3002 7791 3003 7796
rect 3007 7791 3008 7796
rect 3088 7796 3095 7797
rect 2897 7788 2904 7789
rect 2944 7790 2951 7791
rect 2973 7790 2980 7791
rect 2989 7790 2996 7791
rect 3002 7790 3008 7791
rect 3018 7791 3025 7792
rect 2886 7784 2893 7785
rect 2920 7785 2927 7786
rect 2920 7784 2921 7785
rect 2887 7780 2921 7784
rect 2926 7780 2927 7785
rect 2944 7785 2945 7790
rect 2950 7785 2951 7790
rect 2944 7784 2951 7785
rect 2959 7786 2966 7787
rect 2887 7779 2927 7780
rect 2959 7780 2960 7786
rect 2965 7781 2966 7786
rect 2989 7785 2990 7790
rect 2995 7785 2996 7790
rect 3018 7786 3019 7791
rect 3024 7786 3025 7791
rect 3088 7791 3089 7796
rect 3094 7791 3095 7796
rect 3158 7794 3211 7799
rect 3235 7797 3269 7801
rect 3276 7797 3281 7843
rect 3088 7790 3095 7791
rect 3147 7790 3154 7791
rect 3018 7785 3025 7786
rect 3043 7785 3050 7786
rect 2989 7784 2996 7785
rect 2990 7781 2995 7784
rect 2965 7780 2995 7781
rect 2959 7775 2995 7780
rect 3020 7780 3044 7785
rect 3049 7780 3050 7785
rect 3147 7785 3148 7790
rect 3153 7785 3154 7790
rect 3158 7789 3159 7794
rect 3164 7789 3165 7794
rect 3206 7791 3211 7794
rect 3234 7796 3269 7797
rect 3234 7791 3235 7796
rect 3240 7791 3241 7796
rect 3263 7791 3264 7796
rect 3268 7791 3269 7796
rect 3158 7788 3165 7789
rect 3205 7790 3212 7791
rect 3234 7790 3241 7791
rect 3250 7790 3257 7791
rect 3263 7790 3269 7791
rect 3275 7796 3282 7797
rect 3275 7791 3276 7796
rect 3281 7791 3282 7796
rect 3275 7790 3282 7791
rect 3147 7784 3154 7785
rect 3181 7785 3188 7786
rect 3181 7784 3182 7785
rect 2755 7429 2761 7430
rect 2755 7425 2756 7429
rect 2760 7425 2761 7429
rect 2755 7424 2761 7425
rect 3020 7427 3025 7780
rect 3043 7779 3050 7780
rect 3148 7780 3182 7784
rect 3187 7780 3188 7785
rect 3205 7785 3206 7790
rect 3211 7785 3212 7790
rect 3205 7784 3212 7785
rect 3220 7786 3227 7787
rect 3148 7779 3188 7780
rect 3220 7780 3221 7786
rect 3226 7781 3227 7786
rect 3250 7785 3251 7790
rect 3256 7785 3257 7790
rect 3250 7784 3257 7785
rect 3251 7781 3256 7784
rect 3226 7780 3256 7781
rect 3220 7775 3256 7780
rect 3303 7752 3308 8279
rect 3832 8258 3872 8259
rect 3793 8256 3800 8257
rect 3770 8251 3800 8256
rect 3832 8254 3866 8258
rect 3567 8196 3573 8197
rect 3567 8192 3568 8196
rect 3572 8192 3705 8196
rect 3567 8191 3705 8192
rect 3311 7796 3317 7797
rect 3311 7792 3312 7796
rect 3316 7792 3317 7796
rect 3311 7791 3317 7792
rect 3150 7747 3308 7752
rect 3150 7685 3155 7747
rect 3149 7684 3155 7685
rect 3149 7680 3150 7684
rect 3154 7680 3155 7684
rect 3149 7679 3155 7680
rect 3312 7622 3317 7791
rect 3275 7617 3317 7622
rect 3275 7603 3280 7617
rect 3274 7602 3280 7603
rect 3274 7598 3275 7602
rect 3279 7598 3280 7602
rect 3274 7597 3280 7598
rect 3700 7430 3705 8191
rect 3700 7429 3706 7430
rect 3020 7422 3059 7427
rect 3700 7425 3701 7429
rect 3705 7425 3706 7429
rect 3700 7424 3706 7425
rect 3770 7418 3775 8251
rect 3793 8250 3800 8251
rect 3831 8253 3838 8254
rect 3831 8248 3832 8253
rect 3837 8248 3838 8253
rect 3865 8253 3866 8254
rect 3871 8253 3872 8258
rect 3904 8258 3940 8263
rect 3865 8252 3872 8253
rect 3889 8253 3896 8254
rect 3831 8247 3838 8248
rect 3842 8249 3849 8250
rect 3842 8244 3843 8249
rect 3848 8244 3849 8249
rect 3889 8248 3890 8253
rect 3895 8248 3896 8253
rect 3904 8252 3905 8258
rect 3910 8257 3940 8258
rect 3910 8252 3911 8257
rect 3935 8254 3940 8257
rect 3904 8251 3911 8252
rect 3934 8253 3941 8254
rect 3934 8248 3935 8253
rect 3940 8248 3941 8253
rect 3963 8252 3970 8253
rect 3889 8247 3896 8248
rect 3918 8247 3925 8248
rect 3934 8247 3941 8248
rect 3947 8247 3953 8248
rect 3890 8244 3895 8247
rect 3842 8239 3895 8244
rect 3918 8242 3919 8247
rect 3924 8242 3925 8247
rect 3947 8242 3948 8247
rect 3952 8242 3953 8247
rect 3918 8241 3953 8242
rect 3919 8237 3953 8241
rect 3963 8247 3964 8252
rect 3969 8247 3970 8252
rect 4045 8252 4052 8253
rect 4045 8247 4046 8252
rect 4051 8247 4052 8252
rect 4130 8252 4137 8253
rect 4130 8247 4131 8252
rect 4136 8247 4137 8252
rect 3963 8246 3970 8247
rect 3989 8246 3996 8247
rect 4045 8246 4052 8247
rect 4070 8246 4077 8247
rect 4130 8246 4137 8247
rect 3963 8241 3990 8246
rect 3995 8241 3996 8246
rect 4046 8241 4071 8246
rect 4076 8241 4077 8246
rect 3963 8220 3968 8241
rect 3989 8240 3996 8241
rect 4070 8240 4077 8241
rect 4127 8241 4136 8246
rect 3796 8214 3968 8220
rect 3796 8194 3801 8214
rect 3795 8193 3802 8194
rect 3795 8188 3796 8193
rect 3801 8188 3802 8193
rect 3795 8187 3802 8188
rect 3842 8190 3895 8195
rect 3919 8193 3953 8197
rect 3831 8186 3838 8187
rect 3831 8181 3832 8186
rect 3837 8181 3838 8186
rect 3842 8185 3843 8190
rect 3848 8185 3849 8190
rect 3890 8187 3895 8190
rect 3918 8192 3953 8193
rect 3918 8187 3919 8192
rect 3924 8187 3925 8192
rect 3947 8187 3948 8192
rect 3952 8187 3953 8192
rect 3842 8184 3849 8185
rect 3889 8186 3896 8187
rect 3918 8186 3925 8187
rect 3934 8186 3941 8187
rect 3947 8186 3953 8187
rect 3963 8187 3970 8188
rect 3989 8187 3996 8188
rect 4069 8187 4076 8188
rect 3831 8180 3838 8181
rect 3865 8181 3872 8182
rect 3865 8180 3866 8181
rect 3832 8176 3866 8180
rect 3871 8176 3872 8181
rect 3889 8181 3890 8186
rect 3895 8181 3896 8186
rect 3889 8180 3896 8181
rect 3904 8182 3911 8183
rect 3832 8175 3872 8176
rect 3904 8176 3905 8182
rect 3910 8177 3911 8182
rect 3934 8181 3935 8186
rect 3940 8181 3941 8186
rect 3963 8182 3964 8187
rect 3969 8182 3990 8187
rect 3995 8182 3996 8187
rect 3963 8181 3970 8182
rect 3989 8181 3996 8182
rect 4046 8182 4070 8187
rect 4075 8182 4076 8187
rect 3934 8180 3941 8181
rect 3935 8177 3940 8180
rect 3910 8176 3940 8177
rect 3904 8171 3940 8176
rect 3964 8154 3969 8181
rect 3795 8148 3969 8154
rect 3795 8125 3800 8148
rect 3832 8126 3872 8127
rect 3794 8124 3801 8125
rect 3794 8119 3795 8124
rect 3800 8119 3801 8124
rect 3832 8122 3866 8126
rect 3794 8118 3801 8119
rect 3831 8121 3838 8122
rect 3831 8116 3832 8121
rect 3837 8116 3838 8121
rect 3865 8121 3866 8122
rect 3871 8121 3872 8126
rect 3904 8126 3940 8131
rect 4046 8129 4051 8182
rect 4069 8181 4076 8182
rect 4127 8153 4132 8241
rect 4089 8148 4132 8153
rect 3865 8120 3872 8121
rect 3889 8121 3896 8122
rect 3831 8115 3838 8116
rect 3842 8117 3849 8118
rect 3842 8112 3843 8117
rect 3848 8112 3849 8117
rect 3889 8116 3890 8121
rect 3895 8116 3896 8121
rect 3904 8120 3905 8126
rect 3910 8125 3940 8126
rect 3910 8120 3911 8125
rect 3935 8122 3940 8125
rect 4045 8128 4052 8129
rect 4045 8123 4046 8128
rect 4051 8123 4052 8128
rect 4045 8122 4052 8123
rect 3904 8119 3911 8120
rect 3934 8121 3941 8122
rect 3934 8116 3935 8121
rect 3940 8116 3941 8121
rect 3963 8120 3970 8121
rect 3889 8115 3896 8116
rect 3918 8115 3925 8116
rect 3934 8115 3941 8116
rect 3947 8115 3953 8116
rect 3890 8112 3895 8115
rect 3842 8107 3895 8112
rect 3918 8110 3919 8115
rect 3924 8110 3925 8115
rect 3947 8110 3948 8115
rect 3952 8110 3953 8115
rect 3918 8109 3953 8110
rect 3919 8105 3953 8109
rect 3963 8115 3964 8120
rect 3969 8115 3970 8120
rect 4089 8115 4094 8148
rect 4152 8125 4159 8126
rect 4152 8120 4153 8125
rect 4158 8120 4159 8125
rect 4152 8119 4159 8120
rect 3963 8114 3970 8115
rect 3989 8114 3996 8115
rect 3963 8109 3990 8114
rect 3995 8109 3996 8114
rect 4089 8114 4101 8115
rect 4089 8109 4095 8114
rect 4100 8109 4101 8114
rect 3963 8088 3968 8109
rect 3989 8108 3996 8109
rect 4094 8108 4101 8109
rect 3796 8082 3968 8088
rect 3796 8062 3801 8082
rect 3795 8061 3802 8062
rect 3795 8056 3796 8061
rect 3801 8056 3802 8061
rect 3795 8055 3802 8056
rect 3842 8058 3895 8063
rect 3919 8061 3953 8065
rect 3831 8054 3838 8055
rect 3831 8049 3832 8054
rect 3837 8049 3838 8054
rect 3842 8053 3843 8058
rect 3848 8053 3849 8058
rect 3890 8055 3895 8058
rect 3918 8060 3953 8061
rect 3918 8055 3919 8060
rect 3924 8055 3925 8060
rect 3947 8055 3948 8060
rect 3952 8055 3953 8060
rect 3988 8056 3995 8057
rect 4094 8056 4101 8057
rect 3842 8052 3849 8053
rect 3889 8054 3896 8055
rect 3918 8054 3925 8055
rect 3934 8054 3941 8055
rect 3947 8054 3953 8055
rect 3963 8055 3989 8056
rect 3831 8048 3838 8049
rect 3865 8049 3872 8050
rect 3865 8048 3866 8049
rect 3832 8044 3866 8048
rect 3871 8044 3872 8049
rect 3889 8049 3890 8054
rect 3895 8049 3896 8054
rect 3889 8048 3896 8049
rect 3904 8050 3911 8051
rect 3832 8043 3872 8044
rect 3904 8044 3905 8050
rect 3910 8045 3911 8050
rect 3934 8049 3935 8054
rect 3940 8049 3941 8054
rect 3934 8048 3941 8049
rect 3963 8050 3964 8055
rect 3969 8051 3989 8055
rect 3994 8051 3995 8056
rect 3969 8050 3970 8051
rect 3988 8050 3995 8051
rect 4090 8051 4095 8056
rect 4100 8051 4101 8056
rect 4090 8050 4101 8051
rect 3963 8049 3970 8050
rect 3935 8045 3940 8048
rect 3910 8044 3940 8045
rect 3904 8039 3940 8044
rect 3963 8022 3968 8049
rect 3795 8016 3968 8022
rect 4090 8022 4095 8050
rect 4090 8017 4133 8022
rect 3795 7993 3800 8016
rect 3832 7994 3872 7995
rect 3794 7992 3801 7993
rect 3794 7987 3795 7992
rect 3800 7987 3801 7992
rect 3832 7990 3866 7994
rect 3794 7986 3801 7987
rect 3831 7989 3838 7990
rect 3831 7984 3832 7989
rect 3837 7984 3838 7989
rect 3865 7989 3866 7990
rect 3871 7989 3872 7994
rect 3904 7994 3940 7999
rect 4128 7998 4133 8017
rect 3865 7988 3872 7989
rect 3889 7989 3896 7990
rect 3831 7983 3838 7984
rect 3842 7985 3849 7986
rect 3842 7980 3843 7985
rect 3848 7980 3849 7985
rect 3889 7984 3890 7989
rect 3895 7984 3896 7989
rect 3904 7988 3905 7994
rect 3910 7993 3940 7994
rect 3910 7988 3911 7993
rect 3935 7990 3940 7993
rect 4127 7997 4134 7998
rect 4127 7992 4128 7997
rect 4133 7992 4134 7997
rect 4127 7991 4134 7992
rect 4153 7990 4158 8119
rect 4161 7990 4168 7991
rect 3904 7987 3911 7988
rect 3934 7989 3941 7990
rect 3934 7984 3935 7989
rect 3940 7984 3941 7989
rect 3963 7988 3970 7989
rect 3889 7983 3896 7984
rect 3918 7983 3925 7984
rect 3934 7983 3941 7984
rect 3947 7983 3953 7984
rect 3890 7980 3895 7983
rect 3842 7975 3895 7980
rect 3918 7978 3919 7983
rect 3924 7978 3925 7983
rect 3947 7978 3948 7983
rect 3952 7978 3953 7983
rect 3918 7977 3953 7978
rect 3919 7973 3953 7977
rect 3963 7983 3964 7988
rect 3969 7983 3970 7988
rect 4045 7988 4052 7989
rect 4045 7983 4046 7988
rect 4051 7983 4052 7988
rect 4141 7985 4162 7990
rect 4167 7985 4168 7990
rect 4141 7984 4153 7985
rect 4161 7984 4168 7985
rect 3963 7982 3970 7983
rect 3989 7982 3996 7983
rect 4045 7982 4052 7983
rect 4070 7982 4077 7983
rect 3963 7977 3990 7982
rect 3995 7977 3996 7982
rect 4046 7977 4071 7982
rect 4076 7977 4077 7982
rect 3963 7956 3968 7977
rect 3989 7976 3996 7977
rect 4070 7976 4077 7977
rect 4141 7976 4146 7984
rect 3796 7950 3968 7956
rect 4108 7955 4146 7976
rect 3796 7930 3801 7950
rect 3795 7929 3802 7930
rect 3795 7924 3796 7929
rect 3801 7924 3802 7929
rect 3795 7923 3802 7924
rect 3842 7926 3895 7931
rect 3919 7929 3953 7933
rect 3831 7922 3838 7923
rect 3831 7917 3832 7922
rect 3837 7917 3838 7922
rect 3842 7921 3843 7926
rect 3848 7921 3849 7926
rect 3890 7923 3895 7926
rect 3918 7928 3953 7929
rect 3918 7923 3919 7928
rect 3924 7923 3925 7928
rect 3947 7923 3948 7928
rect 3952 7923 3953 7928
rect 3842 7920 3849 7921
rect 3889 7922 3896 7923
rect 3918 7922 3925 7923
rect 3934 7922 3941 7923
rect 3947 7922 3953 7923
rect 3963 7923 3970 7924
rect 3831 7916 3838 7917
rect 3865 7917 3872 7918
rect 3865 7916 3866 7917
rect 3832 7912 3866 7916
rect 3871 7912 3872 7917
rect 3889 7917 3890 7922
rect 3895 7917 3896 7922
rect 3889 7916 3896 7917
rect 3904 7918 3911 7919
rect 3832 7911 3872 7912
rect 3904 7912 3905 7918
rect 3910 7913 3911 7918
rect 3934 7917 3935 7922
rect 3940 7917 3941 7922
rect 3963 7918 3964 7923
rect 3969 7921 3970 7923
rect 3989 7921 3996 7922
rect 4069 7921 4076 7922
rect 3969 7918 3990 7921
rect 3963 7917 3990 7918
rect 3934 7916 3941 7917
rect 3964 7916 3990 7917
rect 3995 7916 3996 7921
rect 3935 7913 3940 7916
rect 3910 7912 3940 7913
rect 3904 7907 3940 7912
rect 3964 7890 3969 7916
rect 3989 7915 3996 7916
rect 4046 7916 4070 7921
rect 4075 7916 4076 7921
rect 3795 7884 3969 7890
rect 3795 7861 3800 7884
rect 3832 7862 3872 7863
rect 3794 7860 3801 7861
rect 3794 7855 3795 7860
rect 3800 7855 3801 7860
rect 3832 7858 3866 7862
rect 3794 7854 3801 7855
rect 3831 7857 3838 7858
rect 3831 7852 3832 7857
rect 3837 7852 3838 7857
rect 3865 7857 3866 7858
rect 3871 7857 3872 7862
rect 3904 7862 3940 7867
rect 4046 7865 4051 7916
rect 4069 7915 4076 7916
rect 3865 7856 3872 7857
rect 3889 7857 3896 7858
rect 3831 7851 3838 7852
rect 3842 7853 3849 7854
rect 3842 7848 3843 7853
rect 3848 7848 3849 7853
rect 3889 7852 3890 7857
rect 3895 7852 3896 7857
rect 3904 7856 3905 7862
rect 3910 7861 3940 7862
rect 3910 7856 3911 7861
rect 3935 7858 3940 7861
rect 4045 7864 4052 7865
rect 4045 7859 4046 7864
rect 4051 7859 4052 7864
rect 4045 7858 4052 7859
rect 3904 7855 3911 7856
rect 3934 7857 3941 7858
rect 3934 7852 3935 7857
rect 3940 7852 3941 7857
rect 3963 7856 3970 7857
rect 3889 7851 3896 7852
rect 3918 7851 3925 7852
rect 3934 7851 3941 7852
rect 3947 7851 3953 7852
rect 3890 7848 3895 7851
rect 3842 7843 3895 7848
rect 3918 7846 3919 7851
rect 3924 7846 3925 7851
rect 3947 7846 3948 7851
rect 3952 7846 3953 7851
rect 3918 7845 3953 7846
rect 3919 7841 3953 7845
rect 3963 7851 3964 7856
rect 3969 7851 3970 7856
rect 3963 7850 3970 7851
rect 3989 7850 3996 7851
rect 3963 7845 3990 7850
rect 3995 7845 3996 7850
rect 4108 7846 4113 7955
rect 4158 7917 4165 7918
rect 4158 7912 4159 7917
rect 4164 7912 4165 7917
rect 4158 7911 4165 7912
rect 4065 7845 4113 7846
rect 3963 7824 3968 7845
rect 3989 7844 3996 7845
rect 3796 7818 3968 7824
rect 4034 7840 4113 7845
rect 4159 7849 4164 7911
rect 4159 7843 4226 7849
rect 3796 7798 3801 7818
rect 3795 7797 3802 7798
rect 3795 7792 3796 7797
rect 3801 7792 3802 7797
rect 3795 7791 3802 7792
rect 3842 7794 3895 7799
rect 3919 7797 3953 7801
rect 4034 7797 4039 7840
rect 3831 7790 3838 7791
rect 3831 7785 3832 7790
rect 3837 7785 3838 7790
rect 3842 7789 3843 7794
rect 3848 7789 3849 7794
rect 3890 7791 3895 7794
rect 3918 7796 3953 7797
rect 3918 7791 3919 7796
rect 3924 7791 3925 7796
rect 3947 7791 3948 7796
rect 3952 7791 3953 7796
rect 4033 7796 4040 7797
rect 3842 7788 3849 7789
rect 3889 7790 3896 7791
rect 3918 7790 3925 7791
rect 3934 7790 3941 7791
rect 3947 7790 3953 7791
rect 3963 7791 3970 7792
rect 3831 7784 3838 7785
rect 3865 7785 3872 7786
rect 3865 7784 3866 7785
rect 3832 7780 3866 7784
rect 3871 7780 3872 7785
rect 3889 7785 3890 7790
rect 3895 7785 3896 7790
rect 3889 7784 3896 7785
rect 3904 7786 3911 7787
rect 3832 7779 3872 7780
rect 3904 7780 3905 7786
rect 3910 7781 3911 7786
rect 3934 7785 3935 7790
rect 3940 7785 3941 7790
rect 3963 7786 3964 7791
rect 3969 7786 3970 7791
rect 4033 7791 4034 7796
rect 4039 7791 4040 7796
rect 4103 7794 4156 7799
rect 4180 7797 4214 7801
rect 4221 7797 4226 7843
rect 4033 7790 4040 7791
rect 4092 7790 4099 7791
rect 3963 7785 3970 7786
rect 3988 7785 3995 7786
rect 3934 7784 3941 7785
rect 3935 7781 3940 7784
rect 3910 7780 3940 7781
rect 3965 7780 3989 7785
rect 3994 7780 3995 7785
rect 4092 7785 4093 7790
rect 4098 7785 4099 7790
rect 4103 7789 4104 7794
rect 4109 7789 4110 7794
rect 4151 7791 4156 7794
rect 4179 7796 4214 7797
rect 4179 7791 4180 7796
rect 4185 7791 4186 7796
rect 4208 7791 4209 7796
rect 4213 7791 4214 7796
rect 4103 7788 4110 7789
rect 4150 7790 4157 7791
rect 4179 7790 4186 7791
rect 4195 7790 4202 7791
rect 4208 7790 4214 7791
rect 4220 7796 4227 7797
rect 4220 7791 4221 7796
rect 4226 7791 4227 7796
rect 4220 7790 4227 7791
rect 4092 7784 4099 7785
rect 4126 7785 4133 7786
rect 4126 7784 4127 7785
rect 3904 7775 3940 7780
rect 3988 7779 3995 7780
rect 4093 7780 4127 7784
rect 4132 7780 4133 7785
rect 4150 7785 4151 7790
rect 4156 7785 4157 7790
rect 4150 7784 4157 7785
rect 4165 7786 4172 7787
rect 4093 7779 4133 7780
rect 4165 7780 4166 7786
rect 4171 7781 4172 7786
rect 4195 7785 4196 7790
rect 4201 7785 4202 7790
rect 4195 7784 4202 7785
rect 4196 7781 4201 7784
rect 4171 7780 4201 7781
rect 4165 7775 4201 7780
rect 4248 7752 4253 8279
rect 4095 7747 4253 7752
rect 4403 8133 4518 8423
rect 4403 8129 4479 8133
rect 4483 8129 4489 8133
rect 4493 8129 4499 8133
rect 4503 8129 4509 8133
rect 4513 8129 4518 8133
rect 4403 8128 4518 8129
rect 4403 8124 4479 8128
rect 4483 8124 4489 8128
rect 4493 8124 4499 8128
rect 4503 8124 4509 8128
rect 4513 8124 4518 8128
rect 4403 8123 4518 8124
rect 4403 8119 4479 8123
rect 4483 8119 4489 8123
rect 4493 8119 4499 8123
rect 4503 8119 4509 8123
rect 4513 8119 4518 8123
rect 4403 8118 4518 8119
rect 4403 8114 4479 8118
rect 4483 8114 4489 8118
rect 4493 8114 4499 8118
rect 4503 8114 4509 8118
rect 4513 8114 4518 8118
rect 4403 8102 4518 8114
rect 4403 8098 4479 8102
rect 4483 8098 4489 8102
rect 4493 8098 4499 8102
rect 4503 8098 4509 8102
rect 4513 8098 4518 8102
rect 4403 8097 4518 8098
rect 4403 8093 4479 8097
rect 4483 8093 4489 8097
rect 4493 8093 4499 8097
rect 4503 8093 4509 8097
rect 4513 8093 4518 8097
rect 4403 8092 4518 8093
rect 4403 8088 4479 8092
rect 4483 8088 4489 8092
rect 4493 8088 4499 8092
rect 4503 8088 4509 8092
rect 4513 8088 4518 8092
rect 4403 8087 4518 8088
rect 4403 8083 4479 8087
rect 4483 8083 4489 8087
rect 4493 8083 4499 8087
rect 4503 8083 4509 8087
rect 4513 8083 4518 8087
rect 4403 8078 4518 8083
rect 4403 8074 4496 8078
rect 4500 8074 4501 8078
rect 4505 8074 4518 8078
rect 4403 8073 4518 8074
rect 4403 8069 4496 8073
rect 4500 8069 4501 8073
rect 4505 8069 4518 8073
rect 4403 8068 4518 8069
rect 4403 8064 4496 8068
rect 4500 8064 4501 8068
rect 4505 8064 4518 8068
rect 4403 8063 4518 8064
rect 4403 8059 4496 8063
rect 4500 8059 4501 8063
rect 4505 8059 4518 8063
rect 4403 8058 4518 8059
rect 4403 8054 4496 8058
rect 4500 8054 4501 8058
rect 4505 8054 4518 8058
rect 4403 8053 4518 8054
rect 4403 8049 4496 8053
rect 4500 8049 4501 8053
rect 4505 8049 4518 8053
rect 4403 8048 4518 8049
rect 4403 8044 4496 8048
rect 4500 8044 4501 8048
rect 4505 8044 4518 8048
rect 4403 8043 4518 8044
rect 4403 8039 4496 8043
rect 4500 8039 4501 8043
rect 4505 8039 4518 8043
rect 4403 8038 4518 8039
rect 4403 8034 4496 8038
rect 4500 8034 4501 8038
rect 4505 8034 4518 8038
rect 4403 8033 4518 8034
rect 4403 8029 4496 8033
rect 4500 8029 4501 8033
rect 4505 8029 4518 8033
rect 4403 8028 4518 8029
rect 4403 8024 4496 8028
rect 4500 8024 4501 8028
rect 4505 8024 4518 8028
rect 4403 7793 4518 8024
rect 4403 7789 4479 7793
rect 4483 7789 4489 7793
rect 4493 7789 4499 7793
rect 4503 7789 4509 7793
rect 4513 7789 4518 7793
rect 4403 7788 4518 7789
rect 4403 7784 4479 7788
rect 4483 7784 4489 7788
rect 4493 7784 4499 7788
rect 4503 7784 4509 7788
rect 4513 7784 4518 7788
rect 4403 7783 4518 7784
rect 4403 7779 4479 7783
rect 4483 7779 4489 7783
rect 4493 7779 4499 7783
rect 4503 7779 4509 7783
rect 4513 7779 4518 7783
rect 4403 7778 4518 7779
rect 4403 7774 4479 7778
rect 4483 7774 4489 7778
rect 4493 7774 4499 7778
rect 4503 7774 4509 7778
rect 4513 7774 4518 7778
rect 4095 7685 4100 7747
rect 4094 7684 4100 7685
rect 4094 7680 4095 7684
rect 4099 7680 4100 7684
rect 4094 7679 4100 7680
rect 4220 7617 4255 7622
rect 4220 7603 4225 7617
rect 4219 7602 4225 7603
rect 4219 7598 4220 7602
rect 4224 7598 4225 7602
rect 4219 7597 4225 7598
rect 3020 7413 3775 7418
rect 654 7158 659 7162
rect 663 7158 669 7162
rect 673 7158 679 7162
rect 683 7158 689 7162
rect 693 7158 769 7162
rect 654 7127 769 7158
rect 654 7123 659 7127
rect 663 7123 669 7127
rect 673 7123 679 7127
rect 683 7123 689 7127
rect 693 7123 769 7127
rect 654 7122 769 7123
rect 654 7118 659 7122
rect 663 7118 669 7122
rect 673 7118 679 7122
rect 683 7118 689 7122
rect 693 7118 769 7122
rect 654 7117 769 7118
rect 654 7113 659 7117
rect 663 7113 669 7117
rect 673 7113 679 7117
rect 683 7113 689 7117
rect 693 7113 769 7117
rect 654 7112 769 7113
rect 654 7108 659 7112
rect 663 7108 669 7112
rect 673 7108 679 7112
rect 683 7108 689 7112
rect 693 7108 769 7112
rect 654 6540 769 7108
rect 1397 6896 2152 6901
rect 947 6716 953 6717
rect 947 6712 948 6716
rect 952 6712 953 6716
rect 947 6711 953 6712
rect 947 6697 952 6711
rect 917 6692 952 6697
rect 1072 6634 1078 6635
rect 1072 6630 1073 6634
rect 1077 6630 1078 6634
rect 1072 6629 1078 6630
rect 1072 6567 1077 6629
rect 654 6536 659 6540
rect 663 6536 669 6540
rect 673 6536 679 6540
rect 683 6536 689 6540
rect 693 6536 769 6540
rect 654 6535 769 6536
rect 654 6531 659 6535
rect 663 6531 669 6535
rect 673 6531 679 6535
rect 683 6531 689 6535
rect 693 6531 769 6535
rect 654 6530 769 6531
rect 654 6526 659 6530
rect 663 6526 669 6530
rect 673 6526 679 6530
rect 683 6526 689 6530
rect 693 6526 769 6530
rect 654 6525 769 6526
rect 654 6521 659 6525
rect 663 6521 669 6525
rect 673 6521 679 6525
rect 683 6521 689 6525
rect 693 6521 769 6525
rect 654 6290 769 6521
rect 654 6286 667 6290
rect 671 6286 672 6290
rect 676 6286 769 6290
rect 654 6285 769 6286
rect 654 6281 667 6285
rect 671 6281 672 6285
rect 676 6281 769 6285
rect 654 6280 769 6281
rect 654 6276 667 6280
rect 671 6276 672 6280
rect 676 6276 769 6280
rect 654 6275 769 6276
rect 654 6271 667 6275
rect 671 6271 672 6275
rect 676 6271 769 6275
rect 654 6270 769 6271
rect 654 6266 667 6270
rect 671 6266 672 6270
rect 676 6266 769 6270
rect 654 6265 769 6266
rect 654 6261 667 6265
rect 671 6261 672 6265
rect 676 6261 769 6265
rect 654 6260 769 6261
rect 654 6256 667 6260
rect 671 6256 672 6260
rect 676 6256 769 6260
rect 654 6255 769 6256
rect 654 6251 667 6255
rect 671 6251 672 6255
rect 676 6251 769 6255
rect 654 6250 769 6251
rect 654 6246 667 6250
rect 671 6246 672 6250
rect 676 6246 769 6250
rect 654 6245 769 6246
rect 654 6241 667 6245
rect 671 6241 672 6245
rect 676 6241 769 6245
rect 654 6240 769 6241
rect 654 6236 667 6240
rect 671 6236 672 6240
rect 676 6236 769 6240
rect 654 6231 769 6236
rect 654 6227 659 6231
rect 663 6227 669 6231
rect 673 6227 679 6231
rect 683 6227 689 6231
rect 693 6227 769 6231
rect 654 6226 769 6227
rect 654 6222 659 6226
rect 663 6222 669 6226
rect 673 6222 679 6226
rect 683 6222 689 6226
rect 693 6222 769 6226
rect 654 6221 769 6222
rect 654 6217 659 6221
rect 663 6217 669 6221
rect 673 6217 679 6221
rect 683 6217 689 6221
rect 693 6217 769 6221
rect 654 6216 769 6217
rect 654 6212 659 6216
rect 663 6212 669 6216
rect 673 6212 679 6216
rect 683 6212 689 6216
rect 693 6212 769 6216
rect 654 6200 769 6212
rect 654 6196 659 6200
rect 663 6196 669 6200
rect 673 6196 679 6200
rect 683 6196 689 6200
rect 693 6196 769 6200
rect 654 6195 769 6196
rect 654 6191 659 6195
rect 663 6191 669 6195
rect 673 6191 679 6195
rect 683 6191 689 6195
rect 693 6191 769 6195
rect 654 6190 769 6191
rect 654 6186 659 6190
rect 663 6186 669 6190
rect 673 6186 679 6190
rect 683 6186 689 6190
rect 693 6186 769 6190
rect 654 6185 769 6186
rect 654 6181 659 6185
rect 663 6181 669 6185
rect 673 6181 679 6185
rect 683 6181 689 6185
rect 693 6181 769 6185
rect 654 5891 769 6181
rect 919 6562 1077 6567
rect 919 6035 924 6562
rect 971 6534 1007 6539
rect 971 6533 1001 6534
rect 971 6530 976 6533
rect 970 6529 977 6530
rect 970 6524 971 6529
rect 976 6524 977 6529
rect 1000 6528 1001 6533
rect 1006 6528 1007 6534
rect 1039 6534 1079 6535
rect 1000 6527 1007 6528
rect 1015 6529 1022 6530
rect 1015 6524 1016 6529
rect 1021 6524 1022 6529
rect 1039 6529 1040 6534
rect 1045 6530 1079 6534
rect 1177 6534 1184 6535
rect 1232 6534 1268 6539
rect 1045 6529 1046 6530
rect 1039 6528 1046 6529
rect 1073 6529 1080 6530
rect 945 6523 952 6524
rect 945 6518 946 6523
rect 951 6518 952 6523
rect 945 6517 952 6518
rect 958 6523 964 6524
rect 970 6523 977 6524
rect 986 6523 993 6524
rect 1015 6523 1022 6524
rect 1062 6525 1069 6526
rect 958 6518 959 6523
rect 963 6518 964 6523
rect 986 6518 987 6523
rect 992 6518 993 6523
rect 958 6517 993 6518
rect 1016 6520 1021 6523
rect 1062 6520 1063 6525
rect 1068 6520 1069 6525
rect 1073 6524 1074 6529
rect 1079 6524 1080 6529
rect 1177 6529 1178 6534
rect 1183 6529 1207 6534
rect 1232 6533 1262 6534
rect 1232 6530 1237 6533
rect 1231 6529 1238 6530
rect 1177 6528 1184 6529
rect 1202 6528 1209 6529
rect 1073 6523 1080 6524
rect 1132 6523 1139 6524
rect 946 6471 951 6517
rect 958 6513 992 6517
rect 1016 6515 1069 6520
rect 1132 6518 1133 6523
rect 1138 6518 1139 6523
rect 1202 6523 1203 6528
rect 1208 6523 1209 6528
rect 1231 6524 1232 6529
rect 1237 6524 1238 6529
rect 1261 6528 1262 6533
rect 1267 6528 1268 6534
rect 1300 6534 1340 6535
rect 1261 6527 1268 6528
rect 1276 6529 1283 6530
rect 1276 6524 1277 6529
rect 1282 6524 1283 6529
rect 1300 6529 1301 6534
rect 1306 6530 1340 6534
rect 1306 6529 1307 6530
rect 1300 6528 1307 6529
rect 1334 6529 1341 6530
rect 1202 6522 1209 6523
rect 1219 6523 1225 6524
rect 1231 6523 1238 6524
rect 1247 6523 1254 6524
rect 1276 6523 1283 6524
rect 1323 6525 1330 6526
rect 1132 6517 1139 6518
rect 1219 6518 1220 6523
rect 1224 6518 1225 6523
rect 1247 6518 1248 6523
rect 1253 6518 1254 6523
rect 1219 6517 1254 6518
rect 1277 6520 1282 6523
rect 1323 6520 1324 6525
rect 1329 6520 1330 6525
rect 1334 6524 1335 6529
rect 1340 6524 1341 6529
rect 1334 6523 1341 6524
rect 1133 6474 1138 6517
rect 1219 6513 1253 6517
rect 1277 6515 1330 6520
rect 1370 6522 1377 6523
rect 1370 6517 1371 6522
rect 1376 6517 1377 6522
rect 1370 6516 1377 6517
rect 1371 6496 1376 6516
rect 946 6465 1013 6471
rect 1008 6403 1013 6465
rect 1059 6469 1138 6474
rect 1204 6490 1376 6496
rect 1176 6469 1183 6470
rect 1204 6469 1209 6490
rect 1059 6468 1107 6469
rect 1007 6402 1014 6403
rect 1007 6397 1008 6402
rect 1013 6397 1014 6402
rect 1007 6396 1014 6397
rect 1059 6359 1064 6468
rect 1176 6464 1177 6469
rect 1182 6464 1209 6469
rect 1176 6463 1183 6464
rect 1202 6463 1209 6464
rect 1202 6458 1203 6463
rect 1208 6458 1209 6463
rect 1219 6469 1253 6473
rect 1219 6468 1254 6469
rect 1219 6463 1220 6468
rect 1224 6463 1225 6468
rect 1247 6463 1248 6468
rect 1253 6463 1254 6468
rect 1277 6466 1330 6471
rect 1277 6463 1282 6466
rect 1219 6462 1225 6463
rect 1231 6462 1238 6463
rect 1247 6462 1254 6463
rect 1276 6462 1283 6463
rect 1202 6457 1209 6458
rect 1231 6457 1232 6462
rect 1237 6457 1238 6462
rect 1231 6456 1238 6457
rect 1261 6458 1268 6459
rect 1120 6455 1127 6456
rect 1120 6450 1121 6455
rect 1126 6450 1127 6455
rect 1120 6449 1127 6450
rect 1232 6453 1237 6456
rect 1261 6453 1262 6458
rect 1232 6452 1262 6453
rect 1267 6452 1268 6458
rect 1276 6457 1277 6462
rect 1282 6457 1283 6462
rect 1323 6461 1324 6466
rect 1329 6461 1330 6466
rect 1323 6460 1330 6461
rect 1334 6462 1341 6463
rect 1276 6456 1283 6457
rect 1300 6457 1307 6458
rect 1096 6398 1103 6399
rect 1121 6398 1126 6449
rect 1232 6447 1268 6452
rect 1300 6452 1301 6457
rect 1306 6456 1307 6457
rect 1334 6457 1335 6462
rect 1340 6457 1341 6462
rect 1334 6456 1341 6457
rect 1371 6459 1378 6460
rect 1306 6452 1340 6456
rect 1371 6454 1372 6459
rect 1377 6454 1378 6459
rect 1371 6453 1378 6454
rect 1300 6451 1340 6452
rect 1372 6430 1377 6453
rect 1203 6424 1377 6430
rect 1096 6393 1097 6398
rect 1102 6393 1126 6398
rect 1176 6398 1183 6399
rect 1203 6398 1208 6424
rect 1232 6402 1268 6407
rect 1232 6401 1262 6402
rect 1232 6398 1237 6401
rect 1176 6393 1177 6398
rect 1182 6397 1208 6398
rect 1231 6397 1238 6398
rect 1182 6396 1209 6397
rect 1182 6393 1203 6396
rect 1096 6392 1103 6393
rect 1176 6392 1183 6393
rect 1202 6391 1203 6393
rect 1208 6391 1209 6396
rect 1231 6392 1232 6397
rect 1237 6392 1238 6397
rect 1261 6396 1262 6401
rect 1267 6396 1268 6402
rect 1300 6402 1340 6403
rect 1261 6395 1268 6396
rect 1276 6397 1283 6398
rect 1276 6392 1277 6397
rect 1282 6392 1283 6397
rect 1300 6397 1301 6402
rect 1306 6398 1340 6402
rect 1306 6397 1307 6398
rect 1300 6396 1307 6397
rect 1334 6397 1341 6398
rect 1202 6390 1209 6391
rect 1219 6391 1225 6392
rect 1231 6391 1238 6392
rect 1247 6391 1254 6392
rect 1276 6391 1283 6392
rect 1323 6393 1330 6394
rect 1219 6386 1220 6391
rect 1224 6386 1225 6391
rect 1247 6386 1248 6391
rect 1253 6386 1254 6391
rect 1219 6385 1254 6386
rect 1277 6388 1282 6391
rect 1323 6388 1324 6393
rect 1329 6388 1330 6393
rect 1334 6392 1335 6397
rect 1340 6392 1341 6397
rect 1334 6391 1341 6392
rect 1219 6381 1253 6385
rect 1277 6383 1330 6388
rect 1370 6390 1377 6391
rect 1370 6385 1371 6390
rect 1376 6385 1377 6390
rect 1370 6384 1377 6385
rect 1371 6364 1376 6384
rect 1026 6338 1064 6359
rect 1204 6358 1376 6364
rect 1026 6330 1031 6338
rect 1095 6337 1102 6338
rect 1176 6337 1183 6338
rect 1204 6337 1209 6358
rect 1095 6332 1096 6337
rect 1101 6332 1126 6337
rect 1176 6332 1177 6337
rect 1182 6332 1209 6337
rect 1095 6331 1102 6332
rect 1120 6331 1127 6332
rect 1176 6331 1183 6332
rect 1202 6331 1209 6332
rect 1004 6329 1011 6330
rect 1019 6329 1031 6330
rect 1004 6324 1005 6329
rect 1010 6324 1031 6329
rect 1120 6326 1121 6331
rect 1126 6326 1127 6331
rect 1120 6325 1127 6326
rect 1202 6326 1203 6331
rect 1208 6326 1209 6331
rect 1219 6337 1253 6341
rect 1219 6336 1254 6337
rect 1219 6331 1220 6336
rect 1224 6331 1225 6336
rect 1247 6331 1248 6336
rect 1253 6331 1254 6336
rect 1277 6334 1330 6339
rect 1277 6331 1282 6334
rect 1219 6330 1225 6331
rect 1231 6330 1238 6331
rect 1247 6330 1254 6331
rect 1276 6330 1283 6331
rect 1202 6325 1209 6326
rect 1231 6325 1232 6330
rect 1237 6325 1238 6330
rect 1231 6324 1238 6325
rect 1261 6326 1268 6327
rect 1004 6323 1011 6324
rect 1014 6195 1019 6324
rect 1038 6322 1045 6323
rect 1038 6317 1039 6322
rect 1044 6317 1045 6322
rect 1038 6316 1045 6317
rect 1232 6321 1237 6324
rect 1261 6321 1262 6326
rect 1232 6320 1262 6321
rect 1267 6320 1268 6326
rect 1276 6325 1277 6330
rect 1282 6325 1283 6330
rect 1323 6329 1324 6334
rect 1329 6329 1330 6334
rect 1323 6328 1330 6329
rect 1334 6330 1341 6331
rect 1276 6324 1283 6325
rect 1300 6325 1307 6326
rect 1039 6297 1044 6316
rect 1232 6315 1268 6320
rect 1300 6320 1301 6325
rect 1306 6324 1307 6325
rect 1334 6325 1335 6330
rect 1340 6325 1341 6330
rect 1334 6324 1341 6325
rect 1371 6327 1378 6328
rect 1306 6320 1340 6324
rect 1371 6322 1372 6327
rect 1377 6322 1378 6327
rect 1371 6321 1378 6322
rect 1300 6319 1340 6320
rect 1372 6298 1377 6321
rect 1039 6292 1082 6297
rect 1077 6264 1082 6292
rect 1204 6292 1377 6298
rect 1204 6265 1209 6292
rect 1232 6270 1268 6275
rect 1232 6269 1262 6270
rect 1232 6266 1237 6269
rect 1202 6264 1209 6265
rect 1071 6263 1082 6264
rect 1071 6258 1072 6263
rect 1077 6258 1082 6263
rect 1177 6263 1184 6264
rect 1202 6263 1203 6264
rect 1177 6258 1178 6263
rect 1183 6259 1203 6263
rect 1208 6259 1209 6264
rect 1231 6265 1238 6266
rect 1231 6260 1232 6265
rect 1237 6260 1238 6265
rect 1261 6264 1262 6269
rect 1267 6264 1268 6270
rect 1300 6270 1340 6271
rect 1261 6263 1268 6264
rect 1276 6265 1283 6266
rect 1276 6260 1277 6265
rect 1282 6260 1283 6265
rect 1300 6265 1301 6270
rect 1306 6266 1340 6270
rect 1306 6265 1307 6266
rect 1300 6264 1307 6265
rect 1334 6265 1341 6266
rect 1183 6258 1209 6259
rect 1219 6259 1225 6260
rect 1231 6259 1238 6260
rect 1247 6259 1254 6260
rect 1276 6259 1283 6260
rect 1323 6261 1330 6262
rect 1071 6257 1078 6258
rect 1177 6257 1184 6258
rect 1219 6254 1220 6259
rect 1224 6254 1225 6259
rect 1247 6254 1248 6259
rect 1253 6254 1254 6259
rect 1219 6253 1254 6254
rect 1277 6256 1282 6259
rect 1323 6256 1324 6261
rect 1329 6256 1330 6261
rect 1334 6260 1335 6265
rect 1340 6260 1341 6265
rect 1334 6259 1341 6260
rect 1219 6249 1253 6253
rect 1277 6251 1330 6256
rect 1370 6258 1377 6259
rect 1370 6253 1371 6258
rect 1376 6253 1377 6258
rect 1370 6252 1377 6253
rect 1371 6232 1376 6252
rect 1204 6226 1376 6232
rect 1071 6205 1078 6206
rect 1176 6205 1183 6206
rect 1204 6205 1209 6226
rect 1071 6200 1072 6205
rect 1077 6200 1083 6205
rect 1071 6199 1083 6200
rect 1176 6200 1177 6205
rect 1182 6200 1209 6205
rect 1176 6199 1183 6200
rect 1202 6199 1209 6200
rect 1013 6194 1020 6195
rect 1013 6189 1014 6194
rect 1019 6189 1020 6194
rect 1013 6188 1020 6189
rect 1078 6166 1083 6199
rect 1202 6194 1203 6199
rect 1208 6194 1209 6199
rect 1219 6205 1253 6209
rect 1219 6204 1254 6205
rect 1219 6199 1220 6204
rect 1224 6199 1225 6204
rect 1247 6199 1248 6204
rect 1253 6199 1254 6204
rect 1277 6202 1330 6207
rect 1277 6199 1282 6202
rect 1219 6198 1225 6199
rect 1231 6198 1238 6199
rect 1247 6198 1254 6199
rect 1276 6198 1283 6199
rect 1202 6193 1209 6194
rect 1231 6193 1232 6198
rect 1237 6193 1238 6198
rect 1231 6192 1238 6193
rect 1261 6194 1268 6195
rect 1120 6191 1127 6192
rect 1120 6186 1121 6191
rect 1126 6186 1127 6191
rect 1120 6185 1127 6186
rect 1232 6189 1237 6192
rect 1261 6189 1262 6194
rect 1232 6188 1262 6189
rect 1267 6188 1268 6194
rect 1276 6193 1277 6198
rect 1282 6193 1283 6198
rect 1323 6197 1324 6202
rect 1329 6197 1330 6202
rect 1323 6196 1330 6197
rect 1334 6198 1341 6199
rect 1276 6192 1283 6193
rect 1300 6193 1307 6194
rect 1040 6161 1083 6166
rect 1040 6073 1045 6161
rect 1096 6132 1103 6133
rect 1121 6132 1126 6185
rect 1232 6183 1268 6188
rect 1300 6188 1301 6193
rect 1306 6192 1307 6193
rect 1334 6193 1335 6198
rect 1340 6193 1341 6198
rect 1334 6192 1341 6193
rect 1371 6195 1378 6196
rect 1306 6188 1340 6192
rect 1371 6190 1372 6195
rect 1377 6190 1378 6195
rect 1371 6189 1378 6190
rect 1300 6187 1340 6188
rect 1372 6166 1377 6189
rect 1203 6160 1377 6166
rect 1203 6133 1208 6160
rect 1232 6138 1268 6143
rect 1232 6137 1262 6138
rect 1232 6134 1237 6137
rect 1231 6133 1238 6134
rect 1096 6127 1097 6132
rect 1102 6127 1126 6132
rect 1176 6132 1183 6133
rect 1202 6132 1209 6133
rect 1176 6127 1177 6132
rect 1182 6127 1203 6132
rect 1208 6127 1209 6132
rect 1231 6128 1232 6133
rect 1237 6128 1238 6133
rect 1261 6132 1262 6137
rect 1267 6132 1268 6138
rect 1300 6138 1340 6139
rect 1261 6131 1268 6132
rect 1276 6133 1283 6134
rect 1276 6128 1277 6133
rect 1282 6128 1283 6133
rect 1300 6133 1301 6138
rect 1306 6134 1340 6138
rect 1306 6133 1307 6134
rect 1300 6132 1307 6133
rect 1334 6133 1341 6134
rect 1096 6126 1103 6127
rect 1176 6126 1183 6127
rect 1202 6126 1209 6127
rect 1219 6127 1225 6128
rect 1231 6127 1238 6128
rect 1247 6127 1254 6128
rect 1276 6127 1283 6128
rect 1323 6129 1330 6130
rect 1219 6122 1220 6127
rect 1224 6122 1225 6127
rect 1247 6122 1248 6127
rect 1253 6122 1254 6127
rect 1219 6121 1254 6122
rect 1277 6124 1282 6127
rect 1323 6124 1324 6129
rect 1329 6124 1330 6129
rect 1334 6128 1335 6133
rect 1340 6128 1341 6133
rect 1334 6127 1341 6128
rect 1219 6117 1253 6121
rect 1277 6119 1330 6124
rect 1370 6126 1377 6127
rect 1370 6121 1371 6126
rect 1376 6121 1377 6126
rect 1370 6120 1377 6121
rect 1371 6100 1376 6120
rect 1204 6094 1376 6100
rect 1036 6068 1045 6073
rect 1095 6073 1102 6074
rect 1176 6073 1183 6074
rect 1204 6073 1209 6094
rect 1095 6068 1096 6073
rect 1101 6068 1126 6073
rect 1176 6068 1177 6073
rect 1182 6068 1209 6073
rect 1035 6067 1042 6068
rect 1095 6067 1102 6068
rect 1120 6067 1127 6068
rect 1176 6067 1183 6068
rect 1202 6067 1209 6068
rect 1035 6062 1036 6067
rect 1041 6062 1042 6067
rect 1035 6061 1042 6062
rect 1120 6062 1121 6067
rect 1126 6062 1127 6067
rect 1120 6061 1127 6062
rect 1202 6062 1203 6067
rect 1208 6062 1209 6067
rect 1219 6073 1253 6077
rect 1219 6072 1254 6073
rect 1219 6067 1220 6072
rect 1224 6067 1225 6072
rect 1247 6067 1248 6072
rect 1253 6067 1254 6072
rect 1277 6070 1330 6075
rect 1277 6067 1282 6070
rect 1219 6066 1225 6067
rect 1231 6066 1238 6067
rect 1247 6066 1254 6067
rect 1276 6066 1283 6067
rect 1202 6061 1209 6062
rect 1231 6061 1232 6066
rect 1237 6061 1238 6066
rect 1231 6060 1238 6061
rect 1261 6062 1268 6063
rect 1232 6057 1237 6060
rect 1261 6057 1262 6062
rect 1232 6056 1262 6057
rect 1267 6056 1268 6062
rect 1276 6061 1277 6066
rect 1282 6061 1283 6066
rect 1323 6065 1324 6070
rect 1329 6065 1330 6070
rect 1323 6064 1330 6065
rect 1334 6066 1341 6067
rect 1276 6060 1283 6061
rect 1300 6061 1307 6062
rect 1232 6051 1268 6056
rect 1300 6056 1301 6061
rect 1306 6060 1307 6061
rect 1334 6061 1335 6066
rect 1340 6061 1341 6066
rect 1334 6060 1341 6061
rect 1372 6063 1379 6064
rect 1397 6063 1402 6896
rect 1466 6889 1472 6890
rect 1466 6885 1467 6889
rect 1471 6885 1472 6889
rect 2113 6887 2152 6892
rect 1466 6884 1472 6885
rect 1467 6123 1472 6884
rect 1892 6716 1898 6717
rect 1892 6712 1893 6716
rect 1897 6712 1898 6716
rect 1892 6711 1898 6712
rect 1892 6697 1897 6711
rect 1855 6692 1897 6697
rect 1855 6523 1860 6692
rect 2017 6634 2023 6635
rect 2017 6630 2018 6634
rect 2022 6630 2023 6634
rect 2017 6629 2023 6630
rect 2017 6567 2022 6629
rect 1864 6562 2022 6567
rect 1855 6522 1861 6523
rect 1855 6518 1856 6522
rect 1860 6518 1861 6522
rect 1855 6517 1861 6518
rect 1467 6122 1605 6123
rect 1467 6118 1600 6122
rect 1604 6118 1605 6122
rect 1599 6117 1605 6118
rect 1306 6056 1340 6060
rect 1372 6058 1402 6063
rect 1372 6057 1379 6058
rect 1300 6055 1340 6056
rect 1864 6035 1869 6562
rect 1916 6534 1952 6539
rect 1916 6533 1946 6534
rect 1916 6530 1921 6533
rect 1915 6529 1922 6530
rect 1915 6524 1916 6529
rect 1921 6524 1922 6529
rect 1945 6528 1946 6533
rect 1951 6528 1952 6534
rect 1984 6534 2024 6535
rect 1945 6527 1952 6528
rect 1960 6529 1967 6530
rect 1960 6524 1961 6529
rect 1966 6524 1967 6529
rect 1984 6529 1985 6534
rect 1990 6530 2024 6534
rect 2122 6534 2129 6535
rect 2147 6534 2152 6887
rect 2411 6889 2417 6890
rect 2411 6885 2412 6889
rect 2416 6885 2417 6889
rect 2411 6884 2417 6885
rect 1990 6529 1991 6530
rect 1984 6528 1991 6529
rect 2018 6529 2025 6530
rect 1890 6523 1897 6524
rect 1890 6518 1891 6523
rect 1896 6518 1897 6523
rect 1890 6517 1897 6518
rect 1903 6523 1909 6524
rect 1915 6523 1922 6524
rect 1931 6523 1938 6524
rect 1960 6523 1967 6524
rect 2007 6525 2014 6526
rect 1903 6518 1904 6523
rect 1908 6518 1909 6523
rect 1931 6518 1932 6523
rect 1937 6518 1938 6523
rect 1903 6517 1938 6518
rect 1961 6520 1966 6523
rect 2007 6520 2008 6525
rect 2013 6520 2014 6525
rect 2018 6524 2019 6529
rect 2024 6524 2025 6529
rect 2122 6529 2123 6534
rect 2128 6529 2152 6534
rect 2177 6534 2213 6539
rect 2177 6533 2207 6534
rect 2177 6530 2182 6533
rect 2176 6529 2183 6530
rect 2122 6528 2129 6529
rect 2147 6528 2154 6529
rect 2018 6523 2025 6524
rect 2077 6523 2084 6524
rect 1891 6471 1896 6517
rect 1903 6513 1937 6517
rect 1961 6515 2014 6520
rect 2077 6518 2078 6523
rect 2083 6518 2084 6523
rect 2147 6523 2148 6528
rect 2153 6523 2154 6528
rect 2176 6524 2177 6529
rect 2182 6524 2183 6529
rect 2206 6528 2207 6533
rect 2212 6528 2213 6534
rect 2245 6534 2285 6535
rect 2206 6527 2213 6528
rect 2221 6529 2228 6530
rect 2221 6524 2222 6529
rect 2227 6524 2228 6529
rect 2245 6529 2246 6534
rect 2251 6530 2285 6534
rect 2251 6529 2252 6530
rect 2245 6528 2252 6529
rect 2279 6529 2286 6530
rect 2147 6522 2154 6523
rect 2164 6523 2170 6524
rect 2176 6523 2183 6524
rect 2192 6523 2199 6524
rect 2221 6523 2228 6524
rect 2268 6525 2275 6526
rect 2077 6517 2084 6518
rect 2164 6518 2165 6523
rect 2169 6518 2170 6523
rect 2192 6518 2193 6523
rect 2198 6518 2199 6523
rect 2164 6517 2199 6518
rect 2222 6520 2227 6523
rect 2268 6520 2269 6525
rect 2274 6520 2275 6525
rect 2279 6524 2280 6529
rect 2285 6524 2286 6529
rect 2279 6523 2286 6524
rect 2078 6474 2083 6517
rect 2164 6513 2198 6517
rect 2222 6515 2275 6520
rect 2315 6522 2322 6523
rect 2315 6517 2316 6522
rect 2321 6517 2322 6522
rect 2315 6516 2322 6517
rect 2316 6496 2321 6516
rect 1891 6465 1958 6471
rect 1953 6403 1958 6465
rect 2004 6469 2083 6474
rect 2149 6490 2321 6496
rect 2121 6469 2128 6470
rect 2149 6469 2154 6490
rect 2004 6468 2052 6469
rect 1952 6402 1959 6403
rect 1952 6397 1953 6402
rect 1958 6397 1959 6402
rect 1952 6396 1959 6397
rect 2004 6359 2009 6468
rect 2121 6464 2122 6469
rect 2127 6464 2154 6469
rect 2121 6463 2128 6464
rect 2147 6463 2154 6464
rect 2147 6458 2148 6463
rect 2153 6458 2154 6463
rect 2164 6469 2198 6473
rect 2164 6468 2199 6469
rect 2164 6463 2165 6468
rect 2169 6463 2170 6468
rect 2192 6463 2193 6468
rect 2198 6463 2199 6468
rect 2222 6466 2275 6471
rect 2222 6463 2227 6466
rect 2164 6462 2170 6463
rect 2176 6462 2183 6463
rect 2192 6462 2199 6463
rect 2221 6462 2228 6463
rect 2147 6457 2154 6458
rect 2176 6457 2177 6462
rect 2182 6457 2183 6462
rect 2176 6456 2183 6457
rect 2206 6458 2213 6459
rect 2065 6455 2072 6456
rect 2065 6450 2066 6455
rect 2071 6450 2072 6455
rect 2065 6449 2072 6450
rect 2177 6453 2182 6456
rect 2206 6453 2207 6458
rect 2177 6452 2207 6453
rect 2212 6452 2213 6458
rect 2221 6457 2222 6462
rect 2227 6457 2228 6462
rect 2268 6461 2269 6466
rect 2274 6461 2275 6466
rect 2268 6460 2275 6461
rect 2279 6462 2286 6463
rect 2221 6456 2228 6457
rect 2245 6457 2252 6458
rect 2041 6398 2048 6399
rect 2066 6398 2071 6449
rect 2177 6447 2213 6452
rect 2245 6452 2246 6457
rect 2251 6456 2252 6457
rect 2279 6457 2280 6462
rect 2285 6457 2286 6462
rect 2279 6456 2286 6457
rect 2316 6459 2323 6460
rect 2251 6452 2285 6456
rect 2316 6454 2317 6459
rect 2322 6454 2323 6459
rect 2316 6453 2323 6454
rect 2245 6451 2285 6452
rect 2317 6430 2322 6453
rect 2148 6424 2322 6430
rect 2041 6393 2042 6398
rect 2047 6393 2071 6398
rect 2121 6398 2128 6399
rect 2148 6398 2153 6424
rect 2177 6402 2213 6407
rect 2177 6401 2207 6402
rect 2177 6398 2182 6401
rect 2121 6393 2122 6398
rect 2127 6397 2153 6398
rect 2176 6397 2183 6398
rect 2127 6396 2154 6397
rect 2127 6393 2148 6396
rect 2041 6392 2048 6393
rect 2121 6392 2128 6393
rect 2147 6391 2148 6393
rect 2153 6391 2154 6396
rect 2176 6392 2177 6397
rect 2182 6392 2183 6397
rect 2206 6396 2207 6401
rect 2212 6396 2213 6402
rect 2245 6402 2285 6403
rect 2206 6395 2213 6396
rect 2221 6397 2228 6398
rect 2221 6392 2222 6397
rect 2227 6392 2228 6397
rect 2245 6397 2246 6402
rect 2251 6398 2285 6402
rect 2251 6397 2252 6398
rect 2245 6396 2252 6397
rect 2279 6397 2286 6398
rect 2147 6390 2154 6391
rect 2164 6391 2170 6392
rect 2176 6391 2183 6392
rect 2192 6391 2199 6392
rect 2221 6391 2228 6392
rect 2268 6393 2275 6394
rect 2164 6386 2165 6391
rect 2169 6386 2170 6391
rect 2192 6386 2193 6391
rect 2198 6386 2199 6391
rect 2164 6385 2199 6386
rect 2222 6388 2227 6391
rect 2268 6388 2269 6393
rect 2274 6388 2275 6393
rect 2279 6392 2280 6397
rect 2285 6392 2286 6397
rect 2279 6391 2286 6392
rect 2164 6381 2198 6385
rect 2222 6383 2275 6388
rect 2315 6390 2322 6391
rect 2315 6385 2316 6390
rect 2321 6385 2322 6390
rect 2315 6384 2322 6385
rect 2316 6364 2321 6384
rect 1971 6338 2009 6359
rect 2149 6358 2321 6364
rect 1971 6330 1976 6338
rect 2040 6337 2047 6338
rect 2121 6337 2128 6338
rect 2149 6337 2154 6358
rect 2040 6332 2041 6337
rect 2046 6332 2071 6337
rect 2121 6332 2122 6337
rect 2127 6332 2154 6337
rect 2040 6331 2047 6332
rect 2065 6331 2072 6332
rect 2121 6331 2128 6332
rect 2147 6331 2154 6332
rect 1949 6329 1956 6330
rect 1964 6329 1976 6330
rect 1949 6324 1950 6329
rect 1955 6324 1976 6329
rect 2065 6326 2066 6331
rect 2071 6326 2072 6331
rect 2065 6325 2072 6326
rect 2147 6326 2148 6331
rect 2153 6326 2154 6331
rect 2164 6337 2198 6341
rect 2164 6336 2199 6337
rect 2164 6331 2165 6336
rect 2169 6331 2170 6336
rect 2192 6331 2193 6336
rect 2198 6331 2199 6336
rect 2222 6334 2275 6339
rect 2222 6331 2227 6334
rect 2164 6330 2170 6331
rect 2176 6330 2183 6331
rect 2192 6330 2199 6331
rect 2221 6330 2228 6331
rect 2147 6325 2154 6326
rect 2176 6325 2177 6330
rect 2182 6325 2183 6330
rect 2176 6324 2183 6325
rect 2206 6326 2213 6327
rect 1949 6323 1956 6324
rect 1959 6195 1964 6324
rect 1983 6322 1990 6323
rect 1983 6317 1984 6322
rect 1989 6317 1990 6322
rect 1983 6316 1990 6317
rect 2177 6321 2182 6324
rect 2206 6321 2207 6326
rect 2177 6320 2207 6321
rect 2212 6320 2213 6326
rect 2221 6325 2222 6330
rect 2227 6325 2228 6330
rect 2268 6329 2269 6334
rect 2274 6329 2275 6334
rect 2268 6328 2275 6329
rect 2279 6330 2286 6331
rect 2221 6324 2228 6325
rect 2245 6325 2252 6326
rect 1984 6297 1989 6316
rect 2177 6315 2213 6320
rect 2245 6320 2246 6325
rect 2251 6324 2252 6325
rect 2279 6325 2280 6330
rect 2285 6325 2286 6330
rect 2279 6324 2286 6325
rect 2316 6327 2323 6328
rect 2251 6320 2285 6324
rect 2316 6322 2317 6327
rect 2322 6322 2323 6327
rect 2316 6321 2323 6322
rect 2245 6319 2285 6320
rect 2317 6298 2322 6321
rect 1984 6292 2027 6297
rect 2022 6264 2027 6292
rect 2149 6292 2322 6298
rect 2149 6265 2154 6292
rect 2177 6270 2213 6275
rect 2177 6269 2207 6270
rect 2177 6266 2182 6269
rect 2147 6264 2154 6265
rect 2016 6263 2027 6264
rect 2016 6258 2017 6263
rect 2022 6258 2027 6263
rect 2122 6263 2129 6264
rect 2147 6263 2148 6264
rect 2122 6258 2123 6263
rect 2128 6259 2148 6263
rect 2153 6259 2154 6264
rect 2176 6265 2183 6266
rect 2176 6260 2177 6265
rect 2182 6260 2183 6265
rect 2206 6264 2207 6269
rect 2212 6264 2213 6270
rect 2245 6270 2285 6271
rect 2206 6263 2213 6264
rect 2221 6265 2228 6266
rect 2221 6260 2222 6265
rect 2227 6260 2228 6265
rect 2245 6265 2246 6270
rect 2251 6266 2285 6270
rect 2251 6265 2252 6266
rect 2245 6264 2252 6265
rect 2279 6265 2286 6266
rect 2128 6258 2154 6259
rect 2164 6259 2170 6260
rect 2176 6259 2183 6260
rect 2192 6259 2199 6260
rect 2221 6259 2228 6260
rect 2268 6261 2275 6262
rect 2016 6257 2023 6258
rect 2122 6257 2129 6258
rect 2164 6254 2165 6259
rect 2169 6254 2170 6259
rect 2192 6254 2193 6259
rect 2198 6254 2199 6259
rect 2164 6253 2199 6254
rect 2222 6256 2227 6259
rect 2268 6256 2269 6261
rect 2274 6256 2275 6261
rect 2279 6260 2280 6265
rect 2285 6260 2286 6265
rect 2279 6259 2286 6260
rect 2164 6249 2198 6253
rect 2222 6251 2275 6256
rect 2315 6258 2322 6259
rect 2315 6253 2316 6258
rect 2321 6253 2322 6258
rect 2315 6252 2322 6253
rect 2316 6232 2321 6252
rect 2149 6226 2321 6232
rect 2016 6205 2023 6206
rect 2121 6205 2128 6206
rect 2149 6205 2154 6226
rect 2016 6200 2017 6205
rect 2022 6200 2028 6205
rect 2016 6199 2028 6200
rect 2121 6200 2122 6205
rect 2127 6200 2154 6205
rect 2121 6199 2128 6200
rect 2147 6199 2154 6200
rect 1958 6194 1965 6195
rect 1958 6189 1959 6194
rect 1964 6189 1965 6194
rect 1958 6188 1965 6189
rect 2023 6166 2028 6199
rect 2147 6194 2148 6199
rect 2153 6194 2154 6199
rect 2164 6205 2198 6209
rect 2164 6204 2199 6205
rect 2164 6199 2165 6204
rect 2169 6199 2170 6204
rect 2192 6199 2193 6204
rect 2198 6199 2199 6204
rect 2222 6202 2275 6207
rect 2222 6199 2227 6202
rect 2164 6198 2170 6199
rect 2176 6198 2183 6199
rect 2192 6198 2199 6199
rect 2221 6198 2228 6199
rect 2147 6193 2154 6194
rect 2176 6193 2177 6198
rect 2182 6193 2183 6198
rect 2176 6192 2183 6193
rect 2206 6194 2213 6195
rect 2065 6191 2072 6192
rect 2065 6186 2066 6191
rect 2071 6186 2072 6191
rect 2065 6185 2072 6186
rect 2177 6189 2182 6192
rect 2206 6189 2207 6194
rect 2177 6188 2207 6189
rect 2212 6188 2213 6194
rect 2221 6193 2222 6198
rect 2227 6193 2228 6198
rect 2268 6197 2269 6202
rect 2274 6197 2275 6202
rect 2268 6196 2275 6197
rect 2279 6198 2286 6199
rect 2221 6192 2228 6193
rect 2245 6193 2252 6194
rect 1985 6161 2028 6166
rect 1985 6073 1990 6161
rect 2041 6132 2048 6133
rect 2066 6132 2071 6185
rect 2177 6183 2213 6188
rect 2245 6188 2246 6193
rect 2251 6192 2252 6193
rect 2279 6193 2280 6198
rect 2285 6193 2286 6198
rect 2279 6192 2286 6193
rect 2316 6195 2323 6196
rect 2251 6188 2285 6192
rect 2316 6190 2317 6195
rect 2322 6190 2323 6195
rect 2316 6189 2323 6190
rect 2245 6187 2285 6188
rect 2317 6166 2322 6189
rect 2148 6160 2322 6166
rect 2148 6133 2153 6160
rect 2177 6138 2213 6143
rect 2177 6137 2207 6138
rect 2177 6134 2182 6137
rect 2176 6133 2183 6134
rect 2041 6127 2042 6132
rect 2047 6127 2071 6132
rect 2121 6132 2128 6133
rect 2147 6132 2154 6133
rect 2121 6127 2122 6132
rect 2127 6127 2148 6132
rect 2153 6127 2154 6132
rect 2176 6128 2177 6133
rect 2182 6128 2183 6133
rect 2206 6132 2207 6137
rect 2212 6132 2213 6138
rect 2245 6138 2285 6139
rect 2206 6131 2213 6132
rect 2221 6133 2228 6134
rect 2221 6128 2222 6133
rect 2227 6128 2228 6133
rect 2245 6133 2246 6138
rect 2251 6134 2285 6138
rect 2251 6133 2252 6134
rect 2245 6132 2252 6133
rect 2279 6133 2286 6134
rect 2041 6126 2048 6127
rect 2121 6126 2128 6127
rect 2147 6126 2154 6127
rect 2164 6127 2170 6128
rect 2176 6127 2183 6128
rect 2192 6127 2199 6128
rect 2221 6127 2228 6128
rect 2268 6129 2275 6130
rect 2164 6122 2165 6127
rect 2169 6122 2170 6127
rect 2192 6122 2193 6127
rect 2198 6122 2199 6127
rect 2164 6121 2199 6122
rect 2222 6124 2227 6127
rect 2268 6124 2269 6129
rect 2274 6124 2275 6129
rect 2279 6128 2280 6133
rect 2285 6128 2286 6133
rect 2279 6127 2286 6128
rect 2164 6117 2198 6121
rect 2222 6119 2275 6124
rect 2315 6126 2322 6127
rect 2315 6121 2316 6126
rect 2321 6121 2322 6126
rect 2315 6120 2322 6121
rect 2412 6123 2417 6884
rect 2800 6522 2806 6523
rect 2800 6518 2801 6522
rect 2805 6518 2806 6522
rect 2800 6517 2806 6518
rect 2412 6122 2550 6123
rect 2316 6100 2321 6120
rect 2412 6118 2545 6122
rect 2549 6118 2550 6122
rect 2544 6117 2550 6118
rect 2149 6094 2321 6100
rect 1981 6068 1990 6073
rect 2040 6073 2047 6074
rect 2121 6073 2128 6074
rect 2149 6073 2154 6094
rect 2040 6068 2041 6073
rect 2046 6068 2071 6073
rect 2121 6068 2122 6073
rect 2127 6068 2154 6073
rect 1980 6067 1987 6068
rect 2040 6067 2047 6068
rect 2065 6067 2072 6068
rect 2121 6067 2128 6068
rect 2147 6067 2154 6068
rect 1980 6062 1981 6067
rect 1986 6062 1987 6067
rect 1980 6061 1987 6062
rect 2065 6062 2066 6067
rect 2071 6062 2072 6067
rect 2065 6061 2072 6062
rect 2147 6062 2148 6067
rect 2153 6062 2154 6067
rect 2164 6073 2198 6077
rect 2164 6072 2199 6073
rect 2164 6067 2165 6072
rect 2169 6067 2170 6072
rect 2192 6067 2193 6072
rect 2198 6067 2199 6072
rect 2222 6070 2275 6075
rect 2222 6067 2227 6070
rect 2164 6066 2170 6067
rect 2176 6066 2183 6067
rect 2192 6066 2199 6067
rect 2221 6066 2228 6067
rect 2147 6061 2154 6062
rect 2176 6061 2177 6066
rect 2182 6061 2183 6066
rect 2176 6060 2183 6061
rect 2206 6062 2213 6063
rect 2177 6057 2182 6060
rect 2206 6057 2207 6062
rect 2177 6056 2207 6057
rect 2212 6056 2213 6062
rect 2221 6061 2222 6066
rect 2227 6061 2228 6066
rect 2268 6065 2269 6070
rect 2274 6065 2275 6070
rect 2268 6064 2275 6065
rect 2279 6066 2286 6067
rect 2221 6060 2228 6061
rect 2245 6061 2252 6062
rect 2177 6051 2213 6056
rect 2245 6056 2246 6061
rect 2251 6060 2252 6061
rect 2279 6061 2280 6066
rect 2285 6061 2286 6066
rect 2279 6060 2286 6061
rect 2251 6056 2285 6060
rect 2317 6057 2324 6064
rect 2245 6055 2285 6056
rect 919 6034 925 6035
rect 919 6030 920 6034
rect 924 6030 925 6034
rect 919 6029 925 6030
rect 1864 6034 1870 6035
rect 1864 6030 1865 6034
rect 1869 6030 1870 6034
rect 1864 6029 1870 6030
rect 1210 6022 1848 6027
rect 2318 6022 2323 6057
rect 654 5887 659 5891
rect 663 5887 669 5891
rect 673 5887 679 5891
rect 683 5887 689 5891
rect 693 5887 769 5891
rect 654 5886 769 5887
rect 654 5882 659 5886
rect 663 5882 669 5886
rect 673 5882 679 5886
rect 683 5882 689 5886
rect 693 5882 769 5886
rect 654 5881 769 5882
rect 654 5877 659 5881
rect 663 5877 669 5881
rect 673 5877 679 5881
rect 683 5877 689 5881
rect 693 5877 769 5881
rect 654 5876 769 5877
rect 654 5872 659 5876
rect 663 5872 669 5876
rect 673 5872 679 5876
rect 683 5872 689 5876
rect 693 5872 769 5876
rect 654 5582 769 5872
rect 896 6017 1238 6022
rect 1376 6018 1604 6019
rect 896 5689 901 6017
rect 1376 6014 1599 6018
rect 1603 6014 1604 6018
rect 1843 6017 2323 6022
rect 2543 6019 2549 6020
rect 1376 5984 1381 6014
rect 1598 6013 1604 6014
rect 2405 6015 2544 6019
rect 2548 6015 2549 6019
rect 2405 6014 2549 6015
rect 1375 5983 1381 5984
rect 1375 5979 1376 5983
rect 1380 5979 1381 5983
rect 1375 5978 1381 5979
rect 2320 5983 2326 5984
rect 2405 5983 2410 6014
rect 2320 5979 2321 5983
rect 2325 5979 2411 5983
rect 2320 5978 2411 5979
rect 2800 5944 2805 6517
rect 947 5939 2805 5944
rect 947 5735 952 5939
rect 1397 5920 2152 5926
rect 947 5734 953 5735
rect 947 5730 948 5734
rect 952 5730 953 5734
rect 947 5729 953 5730
rect 896 5683 1207 5689
rect 1072 5652 1078 5653
rect 1072 5648 1073 5652
rect 1077 5648 1078 5652
rect 1072 5647 1078 5648
rect 1072 5585 1077 5647
rect 654 5578 659 5582
rect 663 5578 669 5582
rect 673 5578 679 5582
rect 683 5578 689 5582
rect 693 5578 769 5582
rect 654 5577 769 5578
rect 654 5573 659 5577
rect 663 5573 669 5577
rect 673 5573 679 5577
rect 683 5573 689 5577
rect 693 5573 769 5577
rect 654 5572 769 5573
rect 654 5568 659 5572
rect 663 5568 669 5572
rect 673 5568 679 5572
rect 683 5568 689 5572
rect 693 5568 769 5572
rect 654 5567 769 5568
rect 654 5563 659 5567
rect 663 5563 669 5567
rect 673 5563 679 5567
rect 683 5563 689 5567
rect 693 5563 769 5567
rect 654 5273 769 5563
rect 654 5269 659 5273
rect 663 5269 669 5273
rect 673 5269 679 5273
rect 683 5269 689 5273
rect 693 5269 769 5273
rect 654 5268 769 5269
rect 654 5264 659 5268
rect 663 5264 669 5268
rect 673 5264 679 5268
rect 683 5264 689 5268
rect 693 5264 769 5268
rect 654 5263 769 5264
rect 654 5259 659 5263
rect 663 5259 669 5263
rect 673 5259 679 5263
rect 683 5259 689 5263
rect 693 5259 769 5263
rect 654 5258 769 5259
rect 654 5254 659 5258
rect 663 5254 669 5258
rect 673 5254 679 5258
rect 683 5254 689 5258
rect 693 5254 769 5258
rect 654 4872 769 5254
rect 919 5580 1077 5585
rect 919 5053 924 5580
rect 971 5552 1007 5557
rect 971 5551 1001 5552
rect 971 5548 976 5551
rect 970 5547 977 5548
rect 970 5542 971 5547
rect 976 5542 977 5547
rect 1000 5546 1001 5551
rect 1006 5546 1007 5552
rect 1039 5552 1079 5553
rect 1000 5545 1007 5546
rect 1015 5547 1022 5548
rect 1015 5542 1016 5547
rect 1021 5542 1022 5547
rect 1039 5547 1040 5552
rect 1045 5548 1079 5552
rect 1177 5552 1184 5553
rect 1202 5552 1207 5683
rect 1045 5547 1046 5548
rect 1039 5546 1046 5547
rect 1073 5547 1080 5548
rect 945 5541 952 5542
rect 945 5536 946 5541
rect 951 5536 952 5541
rect 945 5535 952 5536
rect 958 5541 964 5542
rect 970 5541 977 5542
rect 986 5541 993 5542
rect 1015 5541 1022 5542
rect 1062 5543 1069 5544
rect 958 5536 959 5541
rect 963 5536 964 5541
rect 986 5536 987 5541
rect 992 5536 993 5541
rect 958 5535 993 5536
rect 1016 5538 1021 5541
rect 1062 5538 1063 5543
rect 1068 5538 1069 5543
rect 1073 5542 1074 5547
rect 1079 5542 1080 5547
rect 1177 5547 1178 5552
rect 1183 5547 1207 5552
rect 1232 5552 1268 5557
rect 1232 5551 1262 5552
rect 1232 5548 1237 5551
rect 1231 5547 1238 5548
rect 1177 5546 1184 5547
rect 1202 5546 1209 5547
rect 1073 5541 1080 5542
rect 1132 5541 1139 5542
rect 946 5489 951 5535
rect 958 5531 992 5535
rect 1016 5533 1069 5538
rect 1132 5536 1133 5541
rect 1138 5536 1139 5541
rect 1202 5541 1203 5546
rect 1208 5541 1209 5546
rect 1231 5542 1232 5547
rect 1237 5542 1238 5547
rect 1261 5546 1262 5551
rect 1267 5546 1268 5552
rect 1300 5552 1340 5553
rect 1261 5545 1268 5546
rect 1276 5547 1283 5548
rect 1276 5542 1277 5547
rect 1282 5542 1283 5547
rect 1300 5547 1301 5552
rect 1306 5548 1340 5552
rect 1306 5547 1307 5548
rect 1300 5546 1307 5547
rect 1334 5547 1341 5548
rect 1202 5540 1209 5541
rect 1219 5541 1225 5542
rect 1231 5541 1238 5542
rect 1247 5541 1254 5542
rect 1276 5541 1283 5542
rect 1323 5543 1330 5544
rect 1132 5535 1139 5536
rect 1219 5536 1220 5541
rect 1224 5536 1225 5541
rect 1247 5536 1248 5541
rect 1253 5536 1254 5541
rect 1219 5535 1254 5536
rect 1277 5538 1282 5541
rect 1323 5538 1324 5543
rect 1329 5538 1330 5543
rect 1334 5542 1335 5547
rect 1340 5542 1341 5547
rect 1334 5541 1341 5542
rect 1133 5492 1138 5535
rect 1219 5531 1253 5535
rect 1277 5533 1330 5538
rect 1370 5540 1377 5541
rect 1370 5535 1371 5540
rect 1376 5535 1377 5540
rect 1370 5534 1377 5535
rect 1371 5514 1376 5534
rect 946 5483 1013 5489
rect 1008 5421 1013 5483
rect 1059 5487 1138 5492
rect 1204 5508 1376 5514
rect 1176 5487 1183 5488
rect 1204 5487 1209 5508
rect 1059 5486 1107 5487
rect 1007 5420 1014 5421
rect 1007 5415 1008 5420
rect 1013 5415 1014 5420
rect 1007 5414 1014 5415
rect 1059 5377 1064 5486
rect 1176 5482 1177 5487
rect 1182 5482 1209 5487
rect 1176 5481 1183 5482
rect 1202 5481 1209 5482
rect 1202 5476 1203 5481
rect 1208 5476 1209 5481
rect 1219 5487 1253 5491
rect 1219 5486 1254 5487
rect 1219 5481 1220 5486
rect 1224 5481 1225 5486
rect 1247 5481 1248 5486
rect 1253 5481 1254 5486
rect 1277 5484 1330 5489
rect 1277 5481 1282 5484
rect 1219 5480 1225 5481
rect 1231 5480 1238 5481
rect 1247 5480 1254 5481
rect 1276 5480 1283 5481
rect 1202 5475 1209 5476
rect 1231 5475 1232 5480
rect 1237 5475 1238 5480
rect 1231 5474 1238 5475
rect 1261 5476 1268 5477
rect 1120 5473 1127 5474
rect 1120 5468 1121 5473
rect 1126 5468 1127 5473
rect 1120 5467 1127 5468
rect 1232 5471 1237 5474
rect 1261 5471 1262 5476
rect 1232 5470 1262 5471
rect 1267 5470 1268 5476
rect 1276 5475 1277 5480
rect 1282 5475 1283 5480
rect 1323 5479 1324 5484
rect 1329 5479 1330 5484
rect 1323 5478 1330 5479
rect 1334 5480 1341 5481
rect 1276 5474 1283 5475
rect 1300 5475 1307 5476
rect 1096 5416 1103 5417
rect 1121 5416 1126 5467
rect 1232 5465 1268 5470
rect 1300 5470 1301 5475
rect 1306 5474 1307 5475
rect 1334 5475 1335 5480
rect 1340 5475 1341 5480
rect 1334 5474 1341 5475
rect 1371 5477 1378 5478
rect 1306 5470 1340 5474
rect 1371 5472 1372 5477
rect 1377 5472 1378 5477
rect 1371 5471 1378 5472
rect 1300 5469 1340 5470
rect 1372 5448 1377 5471
rect 1203 5442 1377 5448
rect 1096 5411 1097 5416
rect 1102 5411 1126 5416
rect 1176 5416 1183 5417
rect 1203 5416 1208 5442
rect 1232 5420 1268 5425
rect 1232 5419 1262 5420
rect 1232 5416 1237 5419
rect 1176 5411 1177 5416
rect 1182 5415 1208 5416
rect 1231 5415 1238 5416
rect 1182 5414 1209 5415
rect 1182 5411 1203 5414
rect 1096 5410 1103 5411
rect 1176 5410 1183 5411
rect 1202 5409 1203 5411
rect 1208 5409 1209 5414
rect 1231 5410 1232 5415
rect 1237 5410 1238 5415
rect 1261 5414 1262 5419
rect 1267 5414 1268 5420
rect 1300 5420 1340 5421
rect 1261 5413 1268 5414
rect 1276 5415 1283 5416
rect 1276 5410 1277 5415
rect 1282 5410 1283 5415
rect 1300 5415 1301 5420
rect 1306 5416 1340 5420
rect 1306 5415 1307 5416
rect 1300 5414 1307 5415
rect 1334 5415 1341 5416
rect 1202 5408 1209 5409
rect 1219 5409 1225 5410
rect 1231 5409 1238 5410
rect 1247 5409 1254 5410
rect 1276 5409 1283 5410
rect 1323 5411 1330 5412
rect 1219 5404 1220 5409
rect 1224 5404 1225 5409
rect 1247 5404 1248 5409
rect 1253 5404 1254 5409
rect 1219 5403 1254 5404
rect 1277 5406 1282 5409
rect 1323 5406 1324 5411
rect 1329 5406 1330 5411
rect 1334 5410 1335 5415
rect 1340 5410 1341 5415
rect 1334 5409 1341 5410
rect 1219 5399 1253 5403
rect 1277 5401 1330 5406
rect 1370 5408 1377 5409
rect 1370 5403 1371 5408
rect 1376 5403 1377 5408
rect 1370 5402 1377 5403
rect 1371 5382 1376 5402
rect 1026 5356 1064 5377
rect 1204 5376 1376 5382
rect 1026 5348 1031 5356
rect 1095 5355 1102 5356
rect 1176 5355 1183 5356
rect 1204 5355 1209 5376
rect 1095 5350 1096 5355
rect 1101 5350 1126 5355
rect 1176 5350 1177 5355
rect 1182 5350 1209 5355
rect 1095 5349 1102 5350
rect 1120 5349 1127 5350
rect 1176 5349 1183 5350
rect 1202 5349 1209 5350
rect 1004 5347 1011 5348
rect 1019 5347 1031 5348
rect 1004 5342 1005 5347
rect 1010 5342 1031 5347
rect 1120 5344 1121 5349
rect 1126 5344 1127 5349
rect 1120 5343 1127 5344
rect 1202 5344 1203 5349
rect 1208 5344 1209 5349
rect 1219 5355 1253 5359
rect 1219 5354 1254 5355
rect 1219 5349 1220 5354
rect 1224 5349 1225 5354
rect 1247 5349 1248 5354
rect 1253 5349 1254 5354
rect 1277 5352 1330 5357
rect 1277 5349 1282 5352
rect 1219 5348 1225 5349
rect 1231 5348 1238 5349
rect 1247 5348 1254 5349
rect 1276 5348 1283 5349
rect 1202 5343 1209 5344
rect 1231 5343 1232 5348
rect 1237 5343 1238 5348
rect 1231 5342 1238 5343
rect 1261 5344 1268 5345
rect 1004 5341 1011 5342
rect 1014 5213 1019 5342
rect 1038 5340 1045 5341
rect 1038 5335 1039 5340
rect 1044 5335 1045 5340
rect 1038 5334 1045 5335
rect 1232 5339 1237 5342
rect 1261 5339 1262 5344
rect 1232 5338 1262 5339
rect 1267 5338 1268 5344
rect 1276 5343 1277 5348
rect 1282 5343 1283 5348
rect 1323 5347 1324 5352
rect 1329 5347 1330 5352
rect 1323 5346 1330 5347
rect 1334 5348 1341 5349
rect 1276 5342 1283 5343
rect 1300 5343 1307 5344
rect 1039 5315 1044 5334
rect 1232 5333 1268 5338
rect 1300 5338 1301 5343
rect 1306 5342 1307 5343
rect 1334 5343 1335 5348
rect 1340 5343 1341 5348
rect 1334 5342 1341 5343
rect 1371 5345 1378 5346
rect 1306 5338 1340 5342
rect 1371 5340 1372 5345
rect 1377 5340 1378 5345
rect 1371 5339 1378 5340
rect 1300 5337 1340 5338
rect 1372 5316 1377 5339
rect 1039 5310 1082 5315
rect 1077 5282 1082 5310
rect 1204 5310 1377 5316
rect 1204 5283 1209 5310
rect 1232 5288 1268 5293
rect 1232 5287 1262 5288
rect 1232 5284 1237 5287
rect 1202 5282 1209 5283
rect 1071 5281 1082 5282
rect 1071 5276 1072 5281
rect 1077 5276 1082 5281
rect 1177 5281 1184 5282
rect 1202 5281 1203 5282
rect 1177 5276 1178 5281
rect 1183 5277 1203 5281
rect 1208 5277 1209 5282
rect 1231 5283 1238 5284
rect 1231 5278 1232 5283
rect 1237 5278 1238 5283
rect 1261 5282 1262 5287
rect 1267 5282 1268 5288
rect 1300 5288 1340 5289
rect 1261 5281 1268 5282
rect 1276 5283 1283 5284
rect 1276 5278 1277 5283
rect 1282 5278 1283 5283
rect 1300 5283 1301 5288
rect 1306 5284 1340 5288
rect 1306 5283 1307 5284
rect 1300 5282 1307 5283
rect 1334 5283 1341 5284
rect 1183 5276 1209 5277
rect 1219 5277 1225 5278
rect 1231 5277 1238 5278
rect 1247 5277 1254 5278
rect 1276 5277 1283 5278
rect 1323 5279 1330 5280
rect 1071 5275 1078 5276
rect 1177 5275 1184 5276
rect 1219 5272 1220 5277
rect 1224 5272 1225 5277
rect 1247 5272 1248 5277
rect 1253 5272 1254 5277
rect 1219 5271 1254 5272
rect 1277 5274 1282 5277
rect 1323 5274 1324 5279
rect 1329 5274 1330 5279
rect 1334 5278 1335 5283
rect 1340 5278 1341 5283
rect 1334 5277 1341 5278
rect 1219 5267 1253 5271
rect 1277 5269 1330 5274
rect 1370 5276 1377 5277
rect 1370 5271 1371 5276
rect 1376 5271 1377 5276
rect 1370 5270 1377 5271
rect 1371 5250 1376 5270
rect 1204 5244 1376 5250
rect 1071 5223 1078 5224
rect 1176 5223 1183 5224
rect 1204 5223 1209 5244
rect 1071 5218 1072 5223
rect 1077 5218 1083 5223
rect 1071 5217 1083 5218
rect 1176 5218 1177 5223
rect 1182 5218 1209 5223
rect 1176 5217 1183 5218
rect 1202 5217 1209 5218
rect 1013 5212 1020 5213
rect 1013 5207 1014 5212
rect 1019 5207 1020 5212
rect 1013 5206 1020 5207
rect 1078 5184 1083 5217
rect 1202 5212 1203 5217
rect 1208 5212 1209 5217
rect 1219 5223 1253 5227
rect 1219 5222 1254 5223
rect 1219 5217 1220 5222
rect 1224 5217 1225 5222
rect 1247 5217 1248 5222
rect 1253 5217 1254 5222
rect 1277 5220 1330 5225
rect 1277 5217 1282 5220
rect 1219 5216 1225 5217
rect 1231 5216 1238 5217
rect 1247 5216 1254 5217
rect 1276 5216 1283 5217
rect 1202 5211 1209 5212
rect 1231 5211 1232 5216
rect 1237 5211 1238 5216
rect 1231 5210 1238 5211
rect 1261 5212 1268 5213
rect 1120 5209 1127 5210
rect 1120 5204 1121 5209
rect 1126 5204 1127 5209
rect 1120 5203 1127 5204
rect 1232 5207 1237 5210
rect 1261 5207 1262 5212
rect 1232 5206 1262 5207
rect 1267 5206 1268 5212
rect 1276 5211 1277 5216
rect 1282 5211 1283 5216
rect 1323 5215 1324 5220
rect 1329 5215 1330 5220
rect 1323 5214 1330 5215
rect 1334 5216 1341 5217
rect 1276 5210 1283 5211
rect 1300 5211 1307 5212
rect 1040 5179 1083 5184
rect 1040 5091 1045 5179
rect 1096 5150 1103 5151
rect 1121 5150 1126 5203
rect 1232 5201 1268 5206
rect 1300 5206 1301 5211
rect 1306 5210 1307 5211
rect 1334 5211 1335 5216
rect 1340 5211 1341 5216
rect 1334 5210 1341 5211
rect 1371 5213 1378 5214
rect 1306 5206 1340 5210
rect 1371 5208 1372 5213
rect 1377 5208 1378 5213
rect 1371 5207 1378 5208
rect 1300 5205 1340 5206
rect 1372 5184 1377 5207
rect 1203 5178 1377 5184
rect 1203 5151 1208 5178
rect 1232 5156 1268 5161
rect 1232 5155 1262 5156
rect 1232 5152 1237 5155
rect 1231 5151 1238 5152
rect 1096 5145 1097 5150
rect 1102 5145 1126 5150
rect 1176 5150 1183 5151
rect 1202 5150 1209 5151
rect 1176 5145 1177 5150
rect 1182 5145 1203 5150
rect 1208 5145 1209 5150
rect 1231 5146 1232 5151
rect 1237 5146 1238 5151
rect 1261 5150 1262 5155
rect 1267 5150 1268 5156
rect 1300 5156 1340 5157
rect 1261 5149 1268 5150
rect 1276 5151 1283 5152
rect 1276 5146 1277 5151
rect 1282 5146 1283 5151
rect 1300 5151 1301 5156
rect 1306 5152 1340 5156
rect 1306 5151 1307 5152
rect 1300 5150 1307 5151
rect 1334 5151 1341 5152
rect 1096 5144 1103 5145
rect 1176 5144 1183 5145
rect 1202 5144 1209 5145
rect 1219 5145 1225 5146
rect 1231 5145 1238 5146
rect 1247 5145 1254 5146
rect 1276 5145 1283 5146
rect 1323 5147 1330 5148
rect 1219 5140 1220 5145
rect 1224 5140 1225 5145
rect 1247 5140 1248 5145
rect 1253 5140 1254 5145
rect 1219 5139 1254 5140
rect 1277 5142 1282 5145
rect 1323 5142 1324 5147
rect 1329 5142 1330 5147
rect 1334 5146 1335 5151
rect 1340 5146 1341 5151
rect 1334 5145 1341 5146
rect 1219 5135 1253 5139
rect 1277 5137 1330 5142
rect 1370 5144 1377 5145
rect 1370 5139 1371 5144
rect 1376 5139 1377 5144
rect 1370 5138 1377 5139
rect 1371 5118 1376 5138
rect 1204 5112 1376 5118
rect 1036 5086 1045 5091
rect 1095 5091 1102 5092
rect 1176 5091 1183 5092
rect 1204 5091 1209 5112
rect 1095 5086 1096 5091
rect 1101 5086 1126 5091
rect 1176 5086 1177 5091
rect 1182 5086 1209 5091
rect 1035 5085 1042 5086
rect 1095 5085 1102 5086
rect 1120 5085 1127 5086
rect 1176 5085 1183 5086
rect 1202 5085 1209 5086
rect 1035 5080 1036 5085
rect 1041 5080 1042 5085
rect 1035 5079 1042 5080
rect 1120 5080 1121 5085
rect 1126 5080 1127 5085
rect 1120 5079 1127 5080
rect 1202 5080 1203 5085
rect 1208 5080 1209 5085
rect 1219 5091 1253 5095
rect 1219 5090 1254 5091
rect 1219 5085 1220 5090
rect 1224 5085 1225 5090
rect 1247 5085 1248 5090
rect 1253 5085 1254 5090
rect 1277 5088 1330 5093
rect 1277 5085 1282 5088
rect 1219 5084 1225 5085
rect 1231 5084 1238 5085
rect 1247 5084 1254 5085
rect 1276 5084 1283 5085
rect 1202 5079 1209 5080
rect 1231 5079 1232 5084
rect 1237 5079 1238 5084
rect 1231 5078 1238 5079
rect 1261 5080 1268 5081
rect 1232 5075 1237 5078
rect 1261 5075 1262 5080
rect 1232 5074 1262 5075
rect 1267 5074 1268 5080
rect 1276 5079 1277 5084
rect 1282 5079 1283 5084
rect 1323 5083 1324 5088
rect 1329 5083 1330 5088
rect 1323 5082 1330 5083
rect 1334 5084 1341 5085
rect 1276 5078 1283 5079
rect 1300 5079 1307 5080
rect 1232 5069 1268 5074
rect 1300 5074 1301 5079
rect 1306 5078 1307 5079
rect 1334 5079 1335 5084
rect 1340 5079 1341 5084
rect 1334 5078 1341 5079
rect 1373 5081 1380 5082
rect 1397 5081 1402 5920
rect 1466 5907 1472 5908
rect 1466 5903 1467 5907
rect 1471 5903 1472 5907
rect 1466 5902 1472 5903
rect 1467 5141 1472 5902
rect 1892 5734 1898 5735
rect 1892 5730 1893 5734
rect 1897 5730 1898 5734
rect 1892 5729 1898 5730
rect 1892 5715 1897 5729
rect 1855 5710 1897 5715
rect 1855 5541 1860 5710
rect 2017 5652 2023 5653
rect 2017 5648 2018 5652
rect 2022 5648 2023 5652
rect 2017 5647 2023 5648
rect 2017 5585 2022 5647
rect 1864 5580 2022 5585
rect 1855 5540 1861 5541
rect 1855 5536 1856 5540
rect 1860 5536 1861 5540
rect 1855 5535 1861 5536
rect 1606 5496 1613 5497
rect 1606 5491 1607 5496
rect 1612 5491 1613 5496
rect 1606 5490 1613 5491
rect 1723 5495 1730 5496
rect 1723 5490 1724 5495
rect 1729 5490 1730 5495
rect 1607 5179 1612 5490
rect 1723 5489 1730 5490
rect 1724 5180 1729 5489
rect 1723 5179 1730 5180
rect 1606 5178 1613 5179
rect 1606 5173 1607 5178
rect 1612 5173 1613 5178
rect 1723 5174 1724 5179
rect 1729 5174 1730 5179
rect 1723 5173 1730 5174
rect 1606 5172 1613 5173
rect 1467 5140 1605 5141
rect 1467 5136 1600 5140
rect 1604 5136 1605 5140
rect 1599 5135 1605 5136
rect 1306 5074 1340 5078
rect 1373 5076 1402 5081
rect 1373 5075 1380 5076
rect 1300 5073 1340 5074
rect 1864 5053 1869 5580
rect 1916 5552 1952 5557
rect 1916 5551 1946 5552
rect 1916 5548 1921 5551
rect 1915 5547 1922 5548
rect 1915 5542 1916 5547
rect 1921 5542 1922 5547
rect 1945 5546 1946 5551
rect 1951 5546 1952 5552
rect 1984 5552 2024 5553
rect 1945 5545 1952 5546
rect 1960 5547 1967 5548
rect 1960 5542 1961 5547
rect 1966 5542 1967 5547
rect 1984 5547 1985 5552
rect 1990 5548 2024 5552
rect 2122 5552 2129 5553
rect 2147 5552 2152 5920
rect 2411 5907 2417 5908
rect 2411 5903 2412 5907
rect 2416 5903 2417 5907
rect 2411 5902 2417 5903
rect 1990 5547 1991 5548
rect 1984 5546 1991 5547
rect 2018 5547 2025 5548
rect 1890 5541 1897 5542
rect 1890 5536 1891 5541
rect 1896 5536 1897 5541
rect 1890 5535 1897 5536
rect 1903 5541 1909 5542
rect 1915 5541 1922 5542
rect 1931 5541 1938 5542
rect 1960 5541 1967 5542
rect 2007 5543 2014 5544
rect 1903 5536 1904 5541
rect 1908 5536 1909 5541
rect 1931 5536 1932 5541
rect 1937 5536 1938 5541
rect 1903 5535 1938 5536
rect 1961 5538 1966 5541
rect 2007 5538 2008 5543
rect 2013 5538 2014 5543
rect 2018 5542 2019 5547
rect 2024 5542 2025 5547
rect 2122 5547 2123 5552
rect 2128 5547 2152 5552
rect 2177 5552 2213 5557
rect 2177 5551 2207 5552
rect 2177 5548 2182 5551
rect 2176 5547 2183 5548
rect 2122 5546 2129 5547
rect 2147 5546 2154 5547
rect 2018 5541 2025 5542
rect 2077 5541 2084 5542
rect 1891 5489 1896 5535
rect 1903 5531 1937 5535
rect 1961 5533 2014 5538
rect 2077 5536 2078 5541
rect 2083 5536 2084 5541
rect 2147 5541 2148 5546
rect 2153 5541 2154 5546
rect 2176 5542 2177 5547
rect 2182 5542 2183 5547
rect 2206 5546 2207 5551
rect 2212 5546 2213 5552
rect 2245 5552 2285 5553
rect 2206 5545 2213 5546
rect 2221 5547 2228 5548
rect 2221 5542 2222 5547
rect 2227 5542 2228 5547
rect 2245 5547 2246 5552
rect 2251 5548 2285 5552
rect 2251 5547 2252 5548
rect 2245 5546 2252 5547
rect 2279 5547 2286 5548
rect 2147 5540 2154 5541
rect 2164 5541 2170 5542
rect 2176 5541 2183 5542
rect 2192 5541 2199 5542
rect 2221 5541 2228 5542
rect 2268 5543 2275 5544
rect 2077 5535 2084 5536
rect 2164 5536 2165 5541
rect 2169 5536 2170 5541
rect 2192 5536 2193 5541
rect 2198 5536 2199 5541
rect 2164 5535 2199 5536
rect 2222 5538 2227 5541
rect 2268 5538 2269 5543
rect 2274 5538 2275 5543
rect 2279 5542 2280 5547
rect 2285 5542 2286 5547
rect 2279 5541 2286 5542
rect 2078 5492 2083 5535
rect 2164 5531 2198 5535
rect 2222 5533 2275 5538
rect 2315 5540 2322 5541
rect 2315 5535 2316 5540
rect 2321 5535 2322 5540
rect 2315 5534 2322 5535
rect 2316 5514 2321 5534
rect 1891 5483 1958 5489
rect 1953 5421 1958 5483
rect 2004 5487 2083 5492
rect 2149 5508 2321 5514
rect 2121 5487 2128 5488
rect 2149 5487 2154 5508
rect 2004 5486 2052 5487
rect 1952 5420 1959 5421
rect 1952 5415 1953 5420
rect 1958 5415 1959 5420
rect 1952 5414 1959 5415
rect 2004 5377 2009 5486
rect 2121 5482 2122 5487
rect 2127 5482 2154 5487
rect 2121 5481 2128 5482
rect 2147 5481 2154 5482
rect 2147 5476 2148 5481
rect 2153 5476 2154 5481
rect 2164 5487 2198 5491
rect 2164 5486 2199 5487
rect 2164 5481 2165 5486
rect 2169 5481 2170 5486
rect 2192 5481 2193 5486
rect 2198 5481 2199 5486
rect 2222 5484 2275 5489
rect 2222 5481 2227 5484
rect 2164 5480 2170 5481
rect 2176 5480 2183 5481
rect 2192 5480 2199 5481
rect 2221 5480 2228 5481
rect 2147 5475 2154 5476
rect 2176 5475 2177 5480
rect 2182 5475 2183 5480
rect 2176 5474 2183 5475
rect 2206 5476 2213 5477
rect 2065 5473 2072 5474
rect 2065 5468 2066 5473
rect 2071 5468 2072 5473
rect 2065 5467 2072 5468
rect 2177 5471 2182 5474
rect 2206 5471 2207 5476
rect 2177 5470 2207 5471
rect 2212 5470 2213 5476
rect 2221 5475 2222 5480
rect 2227 5475 2228 5480
rect 2268 5479 2269 5484
rect 2274 5479 2275 5484
rect 2268 5478 2275 5479
rect 2279 5480 2286 5481
rect 2221 5474 2228 5475
rect 2245 5475 2252 5476
rect 2041 5416 2048 5417
rect 2066 5416 2071 5467
rect 2177 5465 2213 5470
rect 2245 5470 2246 5475
rect 2251 5474 2252 5475
rect 2279 5475 2280 5480
rect 2285 5475 2286 5480
rect 2279 5474 2286 5475
rect 2316 5477 2323 5478
rect 2251 5470 2285 5474
rect 2316 5472 2317 5477
rect 2322 5472 2323 5477
rect 2316 5471 2323 5472
rect 2245 5469 2285 5470
rect 2317 5448 2322 5471
rect 2148 5442 2322 5448
rect 2041 5411 2042 5416
rect 2047 5411 2071 5416
rect 2121 5416 2128 5417
rect 2148 5416 2153 5442
rect 2177 5420 2213 5425
rect 2177 5419 2207 5420
rect 2177 5416 2182 5419
rect 2121 5411 2122 5416
rect 2127 5415 2153 5416
rect 2176 5415 2183 5416
rect 2127 5414 2154 5415
rect 2127 5411 2148 5414
rect 2041 5410 2048 5411
rect 2121 5410 2128 5411
rect 2147 5409 2148 5411
rect 2153 5409 2154 5414
rect 2176 5410 2177 5415
rect 2182 5410 2183 5415
rect 2206 5414 2207 5419
rect 2212 5414 2213 5420
rect 2245 5420 2285 5421
rect 2206 5413 2213 5414
rect 2221 5415 2228 5416
rect 2221 5410 2222 5415
rect 2227 5410 2228 5415
rect 2245 5415 2246 5420
rect 2251 5416 2285 5420
rect 2251 5415 2252 5416
rect 2245 5414 2252 5415
rect 2279 5415 2286 5416
rect 2147 5408 2154 5409
rect 2164 5409 2170 5410
rect 2176 5409 2183 5410
rect 2192 5409 2199 5410
rect 2221 5409 2228 5410
rect 2268 5411 2275 5412
rect 2164 5404 2165 5409
rect 2169 5404 2170 5409
rect 2192 5404 2193 5409
rect 2198 5404 2199 5409
rect 2164 5403 2199 5404
rect 2222 5406 2227 5409
rect 2268 5406 2269 5411
rect 2274 5406 2275 5411
rect 2279 5410 2280 5415
rect 2285 5410 2286 5415
rect 2279 5409 2286 5410
rect 2164 5399 2198 5403
rect 2222 5401 2275 5406
rect 2315 5408 2322 5409
rect 2315 5403 2316 5408
rect 2321 5403 2322 5408
rect 2315 5402 2322 5403
rect 2316 5382 2321 5402
rect 1971 5356 2009 5377
rect 2149 5376 2321 5382
rect 1971 5348 1976 5356
rect 2040 5355 2047 5356
rect 2121 5355 2128 5356
rect 2149 5355 2154 5376
rect 2040 5350 2041 5355
rect 2046 5350 2071 5355
rect 2121 5350 2122 5355
rect 2127 5350 2154 5355
rect 2040 5349 2047 5350
rect 2065 5349 2072 5350
rect 2121 5349 2128 5350
rect 2147 5349 2154 5350
rect 1949 5347 1956 5348
rect 1964 5347 1976 5348
rect 1949 5342 1950 5347
rect 1955 5342 1976 5347
rect 2065 5344 2066 5349
rect 2071 5344 2072 5349
rect 2065 5343 2072 5344
rect 2147 5344 2148 5349
rect 2153 5344 2154 5349
rect 2164 5355 2198 5359
rect 2164 5354 2199 5355
rect 2164 5349 2165 5354
rect 2169 5349 2170 5354
rect 2192 5349 2193 5354
rect 2198 5349 2199 5354
rect 2222 5352 2275 5357
rect 2222 5349 2227 5352
rect 2164 5348 2170 5349
rect 2176 5348 2183 5349
rect 2192 5348 2199 5349
rect 2221 5348 2228 5349
rect 2147 5343 2154 5344
rect 2176 5343 2177 5348
rect 2182 5343 2183 5348
rect 2176 5342 2183 5343
rect 2206 5344 2213 5345
rect 1949 5341 1956 5342
rect 1959 5213 1964 5342
rect 1983 5340 1990 5341
rect 1983 5335 1984 5340
rect 1989 5335 1990 5340
rect 1983 5334 1990 5335
rect 2177 5339 2182 5342
rect 2206 5339 2207 5344
rect 2177 5338 2207 5339
rect 2212 5338 2213 5344
rect 2221 5343 2222 5348
rect 2227 5343 2228 5348
rect 2268 5347 2269 5352
rect 2274 5347 2275 5352
rect 2268 5346 2275 5347
rect 2279 5348 2286 5349
rect 2221 5342 2228 5343
rect 2245 5343 2252 5344
rect 1984 5315 1989 5334
rect 2177 5333 2213 5338
rect 2245 5338 2246 5343
rect 2251 5342 2252 5343
rect 2279 5343 2280 5348
rect 2285 5343 2286 5348
rect 2279 5342 2286 5343
rect 2316 5345 2323 5346
rect 2251 5338 2285 5342
rect 2316 5340 2317 5345
rect 2322 5340 2323 5345
rect 2316 5339 2323 5340
rect 2245 5337 2285 5338
rect 2317 5316 2322 5339
rect 1984 5310 2027 5315
rect 2022 5282 2027 5310
rect 2149 5310 2322 5316
rect 2149 5283 2154 5310
rect 2177 5288 2213 5293
rect 2177 5287 2207 5288
rect 2177 5284 2182 5287
rect 2147 5282 2154 5283
rect 2016 5281 2027 5282
rect 2016 5276 2017 5281
rect 2022 5276 2027 5281
rect 2122 5281 2129 5282
rect 2147 5281 2148 5282
rect 2122 5276 2123 5281
rect 2128 5277 2148 5281
rect 2153 5277 2154 5282
rect 2176 5283 2183 5284
rect 2176 5278 2177 5283
rect 2182 5278 2183 5283
rect 2206 5282 2207 5287
rect 2212 5282 2213 5288
rect 2245 5288 2285 5289
rect 2206 5281 2213 5282
rect 2221 5283 2228 5284
rect 2221 5278 2222 5283
rect 2227 5278 2228 5283
rect 2245 5283 2246 5288
rect 2251 5284 2285 5288
rect 2251 5283 2252 5284
rect 2245 5282 2252 5283
rect 2279 5283 2286 5284
rect 2128 5276 2154 5277
rect 2164 5277 2170 5278
rect 2176 5277 2183 5278
rect 2192 5277 2199 5278
rect 2221 5277 2228 5278
rect 2268 5279 2275 5280
rect 2016 5275 2023 5276
rect 2122 5275 2129 5276
rect 2164 5272 2165 5277
rect 2169 5272 2170 5277
rect 2192 5272 2193 5277
rect 2198 5272 2199 5277
rect 2164 5271 2199 5272
rect 2222 5274 2227 5277
rect 2268 5274 2269 5279
rect 2274 5274 2275 5279
rect 2279 5278 2280 5283
rect 2285 5278 2286 5283
rect 2279 5277 2286 5278
rect 2164 5267 2198 5271
rect 2222 5269 2275 5274
rect 2315 5276 2322 5277
rect 2315 5271 2316 5276
rect 2321 5271 2322 5276
rect 2315 5270 2322 5271
rect 2316 5250 2321 5270
rect 2149 5244 2321 5250
rect 2016 5223 2023 5224
rect 2121 5223 2128 5224
rect 2149 5223 2154 5244
rect 2016 5218 2017 5223
rect 2022 5218 2028 5223
rect 2016 5217 2028 5218
rect 2121 5218 2122 5223
rect 2127 5218 2154 5223
rect 2121 5217 2128 5218
rect 2147 5217 2154 5218
rect 1958 5212 1965 5213
rect 1958 5207 1959 5212
rect 1964 5207 1965 5212
rect 1958 5206 1965 5207
rect 2023 5184 2028 5217
rect 2147 5212 2148 5217
rect 2153 5212 2154 5217
rect 2164 5223 2198 5227
rect 2164 5222 2199 5223
rect 2164 5217 2165 5222
rect 2169 5217 2170 5222
rect 2192 5217 2193 5222
rect 2198 5217 2199 5222
rect 2222 5220 2275 5225
rect 2222 5217 2227 5220
rect 2164 5216 2170 5217
rect 2176 5216 2183 5217
rect 2192 5216 2199 5217
rect 2221 5216 2228 5217
rect 2147 5211 2154 5212
rect 2176 5211 2177 5216
rect 2182 5211 2183 5216
rect 2176 5210 2183 5211
rect 2206 5212 2213 5213
rect 2065 5209 2072 5210
rect 2065 5204 2066 5209
rect 2071 5204 2072 5209
rect 2065 5203 2072 5204
rect 2177 5207 2182 5210
rect 2206 5207 2207 5212
rect 2177 5206 2207 5207
rect 2212 5206 2213 5212
rect 2221 5211 2222 5216
rect 2227 5211 2228 5216
rect 2268 5215 2269 5220
rect 2274 5215 2275 5220
rect 2268 5214 2275 5215
rect 2279 5216 2286 5217
rect 2221 5210 2228 5211
rect 2245 5211 2252 5212
rect 1985 5179 2028 5184
rect 1985 5091 1990 5179
rect 2041 5150 2048 5151
rect 2066 5150 2071 5203
rect 2177 5201 2213 5206
rect 2245 5206 2246 5211
rect 2251 5210 2252 5211
rect 2279 5211 2280 5216
rect 2285 5211 2286 5216
rect 2279 5210 2286 5211
rect 2316 5213 2323 5214
rect 2251 5206 2285 5210
rect 2316 5208 2317 5213
rect 2322 5208 2323 5213
rect 2316 5207 2323 5208
rect 2245 5205 2285 5206
rect 2317 5184 2322 5207
rect 2148 5178 2322 5184
rect 2148 5151 2153 5178
rect 2177 5156 2213 5161
rect 2177 5155 2207 5156
rect 2177 5152 2182 5155
rect 2176 5151 2183 5152
rect 2041 5145 2042 5150
rect 2047 5145 2071 5150
rect 2121 5150 2128 5151
rect 2147 5150 2154 5151
rect 2121 5145 2122 5150
rect 2127 5145 2148 5150
rect 2153 5145 2154 5150
rect 2176 5146 2177 5151
rect 2182 5146 2183 5151
rect 2206 5150 2207 5155
rect 2212 5150 2213 5156
rect 2245 5156 2285 5157
rect 2206 5149 2213 5150
rect 2221 5151 2228 5152
rect 2221 5146 2222 5151
rect 2227 5146 2228 5151
rect 2245 5151 2246 5156
rect 2251 5152 2285 5156
rect 2251 5151 2252 5152
rect 2245 5150 2252 5151
rect 2279 5151 2286 5152
rect 2041 5144 2048 5145
rect 2121 5144 2128 5145
rect 2147 5144 2154 5145
rect 2164 5145 2170 5146
rect 2176 5145 2183 5146
rect 2192 5145 2199 5146
rect 2221 5145 2228 5146
rect 2268 5147 2275 5148
rect 2164 5140 2165 5145
rect 2169 5140 2170 5145
rect 2192 5140 2193 5145
rect 2198 5140 2199 5145
rect 2164 5139 2199 5140
rect 2222 5142 2227 5145
rect 2268 5142 2269 5147
rect 2274 5142 2275 5147
rect 2279 5146 2280 5151
rect 2285 5146 2286 5151
rect 2279 5145 2286 5146
rect 2164 5135 2198 5139
rect 2222 5137 2275 5142
rect 2315 5144 2322 5145
rect 2315 5139 2316 5144
rect 2321 5139 2322 5144
rect 2315 5138 2322 5139
rect 2412 5141 2417 5902
rect 4250 5537 4255 7617
rect 4403 7504 4518 7774
rect 4406 7475 4518 7504
rect 4406 7471 4496 7475
rect 4500 7471 4501 7475
rect 4505 7471 4518 7475
rect 4406 7470 4518 7471
rect 4406 7466 4496 7470
rect 4500 7466 4501 7470
rect 4505 7466 4518 7470
rect 4406 7465 4518 7466
rect 4406 7461 4496 7465
rect 4500 7461 4501 7465
rect 4505 7461 4518 7465
rect 4406 7460 4518 7461
rect 4406 7456 4496 7460
rect 4500 7456 4501 7460
rect 4505 7456 4518 7460
rect 4406 7455 4518 7456
rect 4406 7451 4496 7455
rect 4500 7451 4501 7455
rect 4505 7451 4518 7455
rect 4406 7450 4518 7451
rect 4406 7446 4496 7450
rect 4500 7446 4501 7450
rect 4505 7446 4518 7450
rect 4406 7445 4518 7446
rect 4406 7441 4496 7445
rect 4500 7441 4501 7445
rect 4505 7441 4518 7445
rect 4406 7440 4518 7441
rect 4406 7436 4496 7440
rect 4500 7436 4501 7440
rect 4505 7436 4518 7440
rect 4406 7435 4518 7436
rect 4406 7431 4496 7435
rect 4500 7431 4501 7435
rect 4505 7431 4518 7435
rect 4406 7430 4518 7431
rect 4406 7426 4496 7430
rect 4500 7426 4501 7430
rect 4505 7426 4518 7430
rect 4406 7425 4518 7426
rect 4406 7421 4496 7425
rect 4500 7421 4501 7425
rect 4505 7421 4518 7425
rect 4406 7420 4518 7421
rect 4406 7416 4496 7420
rect 4500 7416 4501 7420
rect 4505 7416 4518 7420
rect 4406 7415 4518 7416
rect 4406 7411 4496 7415
rect 4500 7411 4501 7415
rect 4505 7411 4518 7415
rect 4406 7293 4518 7411
rect 4406 7289 4496 7293
rect 4500 7289 4501 7293
rect 4505 7289 4518 7293
rect 4406 7288 4518 7289
rect 4406 7284 4496 7288
rect 4500 7284 4501 7288
rect 4505 7284 4518 7288
rect 4406 7283 4518 7284
rect 4406 7279 4496 7283
rect 4500 7279 4501 7283
rect 4505 7279 4518 7283
rect 4406 7278 4518 7279
rect 4406 7274 4496 7278
rect 4500 7274 4501 7278
rect 4505 7274 4518 7278
rect 4406 7273 4518 7274
rect 4406 7269 4496 7273
rect 4500 7269 4501 7273
rect 4505 7269 4518 7273
rect 4406 7268 4518 7269
rect 4406 7264 4496 7268
rect 4500 7264 4501 7268
rect 4505 7264 4518 7268
rect 4406 7263 4518 7264
rect 4406 7259 4496 7263
rect 4500 7259 4501 7263
rect 4505 7259 4518 7263
rect 4406 7258 4518 7259
rect 4406 7254 4496 7258
rect 4500 7254 4501 7258
rect 4505 7254 4518 7258
rect 4406 7253 4518 7254
rect 4406 7249 4496 7253
rect 4500 7249 4501 7253
rect 4505 7249 4518 7253
rect 4406 7248 4518 7249
rect 4406 7244 4496 7248
rect 4500 7244 4501 7248
rect 4505 7244 4518 7248
rect 4406 7243 4518 7244
rect 4406 7239 4496 7243
rect 4500 7239 4501 7243
rect 4505 7239 4518 7243
rect 4406 7234 4518 7239
rect 4406 7230 4479 7234
rect 4483 7230 4489 7234
rect 4493 7230 4499 7234
rect 4503 7230 4509 7234
rect 4513 7230 4518 7234
rect 4406 7229 4518 7230
rect 4406 7225 4479 7229
rect 4483 7225 4489 7229
rect 4493 7225 4499 7229
rect 4503 7225 4509 7229
rect 4513 7225 4518 7229
rect 4406 7224 4518 7225
rect 4406 7220 4479 7224
rect 4483 7220 4489 7224
rect 4493 7220 4499 7224
rect 4503 7220 4509 7224
rect 4513 7220 4518 7224
rect 4406 7219 4518 7220
rect 4406 7215 4479 7219
rect 4483 7215 4489 7219
rect 4493 7215 4499 7219
rect 4503 7215 4509 7219
rect 4513 7215 4518 7219
rect 4406 7208 4518 7215
rect 4403 7206 4518 7208
rect 4403 7202 4479 7206
rect 4483 7202 4489 7206
rect 4493 7202 4499 7206
rect 4503 7202 4509 7206
rect 4513 7202 4518 7206
rect 4403 7201 4518 7202
rect 4403 7197 4479 7201
rect 4483 7197 4489 7201
rect 4493 7197 4499 7201
rect 4503 7197 4509 7201
rect 4513 7197 4518 7201
rect 4403 7196 4518 7197
rect 4403 7192 4479 7196
rect 4483 7192 4489 7196
rect 4493 7192 4499 7196
rect 4503 7192 4509 7196
rect 4513 7192 4518 7196
rect 4403 7191 4518 7192
rect 4403 7187 4479 7191
rect 4483 7187 4489 7191
rect 4493 7187 4499 7191
rect 4503 7187 4509 7191
rect 4513 7187 4518 7191
rect 4403 7156 4518 7187
rect 4403 7152 4479 7156
rect 4483 7152 4489 7156
rect 4493 7152 4499 7156
rect 4503 7152 4509 7156
rect 4513 7152 4518 7156
rect 4403 6862 4518 7152
rect 4403 6858 4479 6862
rect 4483 6858 4489 6862
rect 4493 6858 4499 6862
rect 4503 6858 4509 6862
rect 4513 6858 4518 6862
rect 4403 6857 4518 6858
rect 4403 6853 4479 6857
rect 4483 6853 4489 6857
rect 4493 6853 4499 6857
rect 4503 6853 4509 6857
rect 4513 6853 4518 6857
rect 4403 6852 4518 6853
rect 4403 6848 4479 6852
rect 4483 6848 4489 6852
rect 4493 6848 4499 6852
rect 4503 6848 4509 6852
rect 4513 6848 4518 6852
rect 4403 6847 4518 6848
rect 4403 6843 4479 6847
rect 4483 6843 4489 6847
rect 4493 6843 4499 6847
rect 4503 6843 4509 6847
rect 4513 6843 4518 6847
rect 4403 6553 4518 6843
rect 4403 6549 4479 6553
rect 4483 6549 4489 6553
rect 4493 6549 4499 6553
rect 4503 6549 4509 6553
rect 4513 6549 4518 6553
rect 4403 6548 4518 6549
rect 4403 6544 4479 6548
rect 4483 6544 4489 6548
rect 4493 6544 4499 6548
rect 4503 6544 4509 6548
rect 4513 6544 4518 6548
rect 4403 6543 4518 6544
rect 4403 6539 4479 6543
rect 4483 6539 4489 6543
rect 4493 6539 4499 6543
rect 4503 6539 4509 6543
rect 4513 6539 4518 6543
rect 4403 6538 4518 6539
rect 4403 6534 4479 6538
rect 4483 6534 4489 6538
rect 4493 6534 4499 6538
rect 4503 6534 4509 6538
rect 4513 6534 4518 6538
rect 4403 6244 4518 6534
rect 4403 6240 4479 6244
rect 4483 6240 4489 6244
rect 4493 6240 4499 6244
rect 4503 6240 4509 6244
rect 4513 6240 4518 6244
rect 4403 6239 4518 6240
rect 4403 6235 4479 6239
rect 4483 6235 4489 6239
rect 4493 6235 4499 6239
rect 4503 6235 4509 6239
rect 4513 6235 4518 6239
rect 4403 6234 4518 6235
rect 4403 6230 4479 6234
rect 4483 6230 4489 6234
rect 4493 6230 4499 6234
rect 4503 6230 4509 6234
rect 4513 6230 4518 6234
rect 4403 6229 4518 6230
rect 4403 6225 4479 6229
rect 4483 6225 4489 6229
rect 4493 6225 4499 6229
rect 4503 6225 4509 6229
rect 4513 6225 4518 6229
rect 4403 5935 4518 6225
rect 4403 5931 4479 5935
rect 4483 5931 4489 5935
rect 4493 5931 4499 5935
rect 4503 5931 4509 5935
rect 4513 5931 4518 5935
rect 4403 5930 4518 5931
rect 4403 5926 4479 5930
rect 4483 5926 4489 5930
rect 4493 5926 4499 5930
rect 4503 5926 4509 5930
rect 4513 5926 4518 5930
rect 4403 5925 4518 5926
rect 4403 5921 4479 5925
rect 4483 5921 4489 5925
rect 4493 5921 4499 5925
rect 4503 5921 4509 5925
rect 4513 5921 4518 5925
rect 4403 5920 4518 5921
rect 4403 5916 4479 5920
rect 4483 5916 4489 5920
rect 4493 5916 4499 5920
rect 4503 5916 4509 5920
rect 4513 5916 4518 5920
rect 4403 5626 4518 5916
rect 4403 5622 4479 5626
rect 4483 5622 4489 5626
rect 4493 5622 4499 5626
rect 4503 5622 4509 5626
rect 4513 5622 4518 5626
rect 4403 5621 4518 5622
rect 4403 5617 4479 5621
rect 4483 5617 4489 5621
rect 4493 5617 4499 5621
rect 4503 5617 4509 5621
rect 4513 5617 4518 5621
rect 4403 5616 4518 5617
rect 4403 5612 4479 5616
rect 4483 5612 4489 5616
rect 4493 5612 4499 5616
rect 4503 5612 4509 5616
rect 4513 5612 4518 5616
rect 4403 5611 4518 5612
rect 4403 5607 4479 5611
rect 4483 5607 4489 5611
rect 4493 5607 4499 5611
rect 4503 5607 4509 5611
rect 4513 5607 4518 5611
rect 4249 5536 4256 5537
rect 4249 5532 4251 5536
rect 4255 5532 4256 5536
rect 4249 5531 4256 5532
rect 4250 5530 4255 5531
rect 4403 5317 4518 5607
rect 4403 5313 4479 5317
rect 4483 5313 4489 5317
rect 4493 5313 4499 5317
rect 4503 5313 4509 5317
rect 4513 5313 4518 5317
rect 4403 5312 4518 5313
rect 4403 5308 4479 5312
rect 4483 5308 4489 5312
rect 4493 5308 4499 5312
rect 4503 5308 4509 5312
rect 4513 5308 4518 5312
rect 4403 5307 4518 5308
rect 4403 5303 4479 5307
rect 4483 5303 4489 5307
rect 4493 5303 4499 5307
rect 4503 5303 4509 5307
rect 4513 5303 4518 5307
rect 4403 5302 4518 5303
rect 4403 5298 4479 5302
rect 4483 5298 4489 5302
rect 4493 5298 4499 5302
rect 4503 5298 4509 5302
rect 4513 5298 4518 5302
rect 2412 5140 2550 5141
rect 2316 5118 2321 5138
rect 2412 5136 2545 5140
rect 2549 5136 2550 5140
rect 2544 5135 2550 5136
rect 2149 5112 2321 5118
rect 1981 5086 1990 5091
rect 2040 5091 2047 5092
rect 2121 5091 2128 5092
rect 2149 5091 2154 5112
rect 2040 5086 2041 5091
rect 2046 5086 2071 5091
rect 2121 5086 2122 5091
rect 2127 5086 2154 5091
rect 1980 5085 1987 5086
rect 2040 5085 2047 5086
rect 2065 5085 2072 5086
rect 2121 5085 2128 5086
rect 2147 5085 2154 5086
rect 1980 5080 1981 5085
rect 1986 5080 1987 5085
rect 1980 5079 1987 5080
rect 2065 5080 2066 5085
rect 2071 5080 2072 5085
rect 2065 5079 2072 5080
rect 2147 5080 2148 5085
rect 2153 5080 2154 5085
rect 2164 5091 2198 5095
rect 2164 5090 2199 5091
rect 2164 5085 2165 5090
rect 2169 5085 2170 5090
rect 2192 5085 2193 5090
rect 2198 5085 2199 5090
rect 2222 5088 2275 5093
rect 2222 5085 2227 5088
rect 2164 5084 2170 5085
rect 2176 5084 2183 5085
rect 2192 5084 2199 5085
rect 2221 5084 2228 5085
rect 2147 5079 2154 5080
rect 2176 5079 2177 5084
rect 2182 5079 2183 5084
rect 2176 5078 2183 5079
rect 2206 5080 2213 5081
rect 2177 5075 2182 5078
rect 2206 5075 2207 5080
rect 2177 5074 2207 5075
rect 2212 5074 2213 5080
rect 2221 5079 2222 5084
rect 2227 5079 2228 5084
rect 2268 5083 2269 5088
rect 2274 5083 2275 5088
rect 2268 5082 2275 5083
rect 2279 5084 2286 5085
rect 2221 5078 2228 5079
rect 2245 5079 2252 5080
rect 2177 5069 2213 5074
rect 2245 5074 2246 5079
rect 2251 5078 2252 5079
rect 2279 5079 2280 5084
rect 2285 5079 2286 5084
rect 2279 5078 2286 5079
rect 2251 5074 2285 5078
rect 2245 5073 2285 5074
rect 919 5052 925 5053
rect 919 5048 920 5052
rect 924 5048 925 5052
rect 919 5047 925 5048
rect 1864 5052 1870 5053
rect 1864 5048 1865 5052
rect 1869 5048 1870 5052
rect 1864 5047 1870 5048
rect 1598 5037 1604 5038
rect 2543 5037 2549 5038
rect 1376 5033 1599 5037
rect 1603 5033 1604 5037
rect 1376 5032 1604 5033
rect 2321 5033 2544 5037
rect 2548 5033 2549 5037
rect 2321 5032 2549 5033
rect 1376 5002 1381 5032
rect 2321 5002 2326 5032
rect 1375 5001 1381 5002
rect 1375 4997 1376 5001
rect 1380 4997 1381 5001
rect 1375 4996 1381 4997
rect 2320 5001 2326 5002
rect 2320 4997 2321 5001
rect 2325 4997 2326 5001
rect 2320 4996 2326 4997
rect 4403 5008 4518 5298
rect 4403 5004 4479 5008
rect 4483 5004 4489 5008
rect 4493 5004 4499 5008
rect 4503 5004 4509 5008
rect 4513 5004 4518 5008
rect 4403 5003 4518 5004
rect 4403 4999 4479 5003
rect 4483 4999 4489 5003
rect 4493 4999 4499 5003
rect 4503 4999 4509 5003
rect 4513 4999 4518 5003
rect 4403 4998 4518 4999
rect 654 4868 659 4872
rect 663 4868 669 4872
rect 673 4868 679 4872
rect 683 4868 689 4872
rect 693 4868 769 4872
rect 654 4867 769 4868
rect 654 4863 659 4867
rect 663 4863 669 4867
rect 673 4863 679 4867
rect 683 4863 689 4867
rect 693 4863 769 4867
rect 654 4862 769 4863
rect 654 4858 659 4862
rect 663 4858 669 4862
rect 673 4858 679 4862
rect 683 4858 689 4862
rect 693 4858 769 4862
rect 654 4857 769 4858
rect 654 4853 659 4857
rect 663 4853 669 4857
rect 673 4853 679 4857
rect 683 4853 689 4857
rect 693 4853 769 4857
rect 654 4843 769 4853
rect 654 4839 659 4843
rect 663 4839 669 4843
rect 673 4839 679 4843
rect 683 4839 689 4843
rect 693 4839 769 4843
rect 654 4838 769 4839
rect 654 4834 659 4838
rect 663 4834 669 4838
rect 673 4834 679 4838
rect 683 4834 689 4838
rect 693 4834 769 4838
rect 654 4833 769 4834
rect 654 4829 659 4833
rect 663 4829 669 4833
rect 673 4829 679 4833
rect 683 4829 689 4833
rect 693 4829 769 4833
rect 654 4828 769 4829
rect 654 4824 659 4828
rect 663 4824 669 4828
rect 673 4824 679 4828
rect 683 4824 689 4828
rect 693 4824 769 4828
rect 654 4814 769 4824
rect 654 4810 659 4814
rect 663 4810 669 4814
rect 673 4810 679 4814
rect 683 4810 689 4814
rect 693 4810 769 4814
rect 654 4809 769 4810
rect 654 4805 659 4809
rect 663 4805 669 4809
rect 673 4805 679 4809
rect 683 4805 689 4809
rect 693 4805 769 4809
rect 654 4804 769 4805
rect 654 4800 659 4804
rect 663 4800 669 4804
rect 673 4800 679 4804
rect 683 4800 689 4804
rect 693 4800 769 4804
rect 654 4799 769 4800
rect 654 4795 659 4799
rect 663 4795 669 4799
rect 673 4795 679 4799
rect 683 4795 689 4799
rect 693 4795 769 4799
rect 654 4785 769 4795
rect 654 4781 659 4785
rect 663 4781 669 4785
rect 673 4781 679 4785
rect 683 4781 689 4785
rect 693 4781 769 4785
rect 654 4780 769 4781
rect 654 4776 659 4780
rect 663 4776 669 4780
rect 673 4776 679 4780
rect 683 4776 689 4780
rect 693 4776 769 4780
rect 654 4775 769 4776
rect 654 4771 659 4775
rect 663 4771 669 4775
rect 673 4771 679 4775
rect 683 4771 689 4775
rect 693 4771 769 4775
rect 654 4770 769 4771
rect 654 4766 659 4770
rect 663 4766 669 4770
rect 673 4766 679 4770
rect 683 4766 689 4770
rect 693 4766 769 4770
rect 654 4756 769 4766
rect 654 4752 659 4756
rect 663 4752 669 4756
rect 673 4752 679 4756
rect 683 4752 689 4756
rect 693 4752 769 4756
rect 654 4751 769 4752
rect 654 4747 659 4751
rect 663 4747 669 4751
rect 673 4747 679 4751
rect 683 4747 689 4751
rect 693 4747 769 4751
rect 654 4746 769 4747
rect 654 4742 659 4746
rect 663 4742 669 4746
rect 673 4742 679 4746
rect 683 4742 689 4746
rect 693 4742 769 4746
rect 654 4741 769 4742
rect 654 4737 659 4741
rect 663 4737 669 4741
rect 673 4737 679 4741
rect 683 4737 689 4741
rect 693 4737 769 4741
rect 654 4704 769 4737
rect 4403 4994 4479 4998
rect 4483 4994 4489 4998
rect 4493 4994 4499 4998
rect 4503 4994 4509 4998
rect 4513 4994 4518 4998
rect 4403 4993 4518 4994
rect 4403 4989 4479 4993
rect 4483 4989 4489 4993
rect 4493 4989 4499 4993
rect 4503 4989 4509 4993
rect 4513 4989 4518 4993
rect 4403 4815 4518 4989
rect 4403 4811 4479 4815
rect 4483 4811 4489 4815
rect 4493 4811 4499 4815
rect 4503 4811 4509 4815
rect 4513 4811 4518 4815
rect 4403 4810 4518 4811
rect 4403 4806 4479 4810
rect 4483 4806 4489 4810
rect 4493 4806 4499 4810
rect 4503 4806 4509 4810
rect 4513 4806 4518 4810
rect 4403 4805 4518 4806
rect 4403 4801 4479 4805
rect 4483 4801 4489 4805
rect 4493 4801 4499 4805
rect 4503 4801 4509 4805
rect 4513 4801 4518 4805
rect 4403 4800 4518 4801
rect 4403 4796 4479 4800
rect 4483 4796 4489 4800
rect 4493 4796 4499 4800
rect 4503 4796 4509 4800
rect 4513 4796 4518 4800
rect 4403 4789 4518 4796
rect 4403 4785 4479 4789
rect 4483 4785 4489 4789
rect 4493 4785 4499 4789
rect 4503 4785 4509 4789
rect 4513 4785 4518 4789
rect 4403 4784 4518 4785
rect 4403 4780 4479 4784
rect 4483 4780 4489 4784
rect 4493 4780 4499 4784
rect 4503 4780 4509 4784
rect 4513 4780 4518 4784
rect 4403 4779 4518 4780
rect 4403 4775 4479 4779
rect 4483 4775 4489 4779
rect 4493 4775 4499 4779
rect 4503 4775 4509 4779
rect 4513 4775 4518 4779
rect 4403 4774 4518 4775
rect 4403 4770 4479 4774
rect 4483 4770 4489 4774
rect 4493 4770 4499 4774
rect 4503 4770 4509 4774
rect 4513 4770 4518 4774
rect 4403 4763 4518 4770
rect 4403 4759 4479 4763
rect 4483 4759 4489 4763
rect 4493 4759 4499 4763
rect 4503 4759 4509 4763
rect 4513 4759 4518 4763
rect 4403 4758 4518 4759
rect 4403 4754 4479 4758
rect 4483 4754 4489 4758
rect 4493 4754 4499 4758
rect 4503 4754 4509 4758
rect 4513 4754 4518 4758
rect 4403 4753 4518 4754
rect 4403 4749 4479 4753
rect 4483 4749 4489 4753
rect 4493 4749 4499 4753
rect 4503 4749 4509 4753
rect 4513 4749 4518 4753
rect 4403 4748 4518 4749
rect 4403 4744 4479 4748
rect 4483 4744 4489 4748
rect 4493 4744 4499 4748
rect 4503 4744 4509 4748
rect 4513 4744 4518 4748
rect 4403 4737 4518 4744
rect 4403 4733 4479 4737
rect 4483 4733 4489 4737
rect 4493 4733 4499 4737
rect 4503 4733 4509 4737
rect 4513 4733 4518 4737
rect 4403 4732 4518 4733
rect 4403 4728 4479 4732
rect 4483 4728 4489 4732
rect 4493 4728 4499 4732
rect 4503 4728 4509 4732
rect 4513 4728 4518 4732
rect 4403 4727 4518 4728
rect 4403 4723 4479 4727
rect 4483 4723 4489 4727
rect 4493 4723 4499 4727
rect 4503 4723 4509 4727
rect 4513 4723 4518 4727
rect 4403 4722 4518 4723
rect 4403 4718 4479 4722
rect 4483 4718 4489 4722
rect 4493 4718 4499 4722
rect 4503 4718 4509 4722
rect 4513 4718 4518 4722
rect 4403 4711 4518 4718
rect 4403 4707 4479 4711
rect 4483 4707 4489 4711
rect 4493 4707 4499 4711
rect 4503 4707 4509 4711
rect 4513 4707 4518 4711
rect 4403 4706 4518 4707
rect 4403 4704 4479 4706
rect 654 4702 4479 4704
rect 4483 4702 4489 4706
rect 4493 4702 4499 4706
rect 4503 4702 4509 4706
rect 4513 4702 4518 4706
rect 654 4701 4518 4702
rect 654 4697 4479 4701
rect 4483 4697 4489 4701
rect 4493 4697 4499 4701
rect 4503 4697 4509 4701
rect 4513 4697 4518 4701
rect 654 4696 4518 4697
rect 654 4695 4479 4696
rect 654 4691 2910 4695
rect 2914 4692 4479 4695
rect 4483 4692 4489 4696
rect 4493 4692 4499 4696
rect 4503 4692 4509 4696
rect 4513 4692 4518 4696
rect 2914 4691 4518 4692
rect 654 4653 4518 4691
rect 654 4649 1820 4653
rect 1824 4649 1825 4653
rect 1829 4649 3674 4653
rect 3678 4649 3679 4653
rect 3683 4649 4518 4653
rect 654 4648 4518 4649
rect 654 4644 1820 4648
rect 1824 4644 1825 4648
rect 1829 4644 3674 4648
rect 3678 4644 3679 4648
rect 3683 4644 4518 4648
rect 654 4643 4518 4644
rect 654 4639 1820 4643
rect 1824 4639 1825 4643
rect 1829 4639 3674 4643
rect 3678 4639 3679 4643
rect 3683 4639 4518 4643
rect 654 4638 4518 4639
rect 654 4634 1820 4638
rect 1824 4634 1825 4638
rect 1829 4634 3674 4638
rect 3678 4634 3679 4638
rect 3683 4634 4518 4638
rect 654 4633 4518 4634
rect 654 4629 1820 4633
rect 1824 4629 1825 4633
rect 1829 4629 3674 4633
rect 3678 4629 3679 4633
rect 3683 4629 4518 4633
rect 654 4628 4518 4629
rect 654 4624 757 4628
rect 761 4624 762 4628
rect 766 4624 767 4628
rect 771 4624 772 4628
rect 776 4624 783 4628
rect 787 4624 788 4628
rect 792 4624 793 4628
rect 797 4624 798 4628
rect 802 4624 809 4628
rect 813 4624 814 4628
rect 818 4624 819 4628
rect 823 4624 824 4628
rect 828 4624 835 4628
rect 839 4624 840 4628
rect 844 4624 845 4628
rect 849 4624 850 4628
rect 854 4624 861 4628
rect 865 4624 866 4628
rect 870 4624 871 4628
rect 875 4624 876 4628
rect 880 4624 1053 4628
rect 1057 4624 1058 4628
rect 1062 4624 1063 4628
rect 1067 4624 1068 4628
rect 1072 4624 1362 4628
rect 1366 4624 1367 4628
rect 1371 4624 1372 4628
rect 1376 4624 1377 4628
rect 1381 4624 1671 4628
rect 1675 4624 1676 4628
rect 1680 4624 1681 4628
rect 1685 4624 1686 4628
rect 1690 4624 1820 4628
rect 1824 4624 1825 4628
rect 1829 4624 1980 4628
rect 1984 4624 1985 4628
rect 1989 4624 1990 4628
rect 1994 4624 1995 4628
rect 1999 4624 2289 4628
rect 2293 4624 2294 4628
rect 2298 4624 2299 4628
rect 2303 4624 2304 4628
rect 2308 4624 2598 4628
rect 2602 4624 2603 4628
rect 2607 4624 2608 4628
rect 2612 4624 2613 4628
rect 2617 4624 2907 4628
rect 2911 4624 2912 4628
rect 2916 4624 2917 4628
rect 2921 4624 2922 4628
rect 2926 4624 3216 4628
rect 3220 4624 3221 4628
rect 3225 4624 3226 4628
rect 3230 4624 3231 4628
rect 3235 4624 3525 4628
rect 3529 4624 3530 4628
rect 3534 4624 3535 4628
rect 3539 4624 3540 4628
rect 3544 4624 3674 4628
rect 3678 4624 3679 4628
rect 3683 4624 3834 4628
rect 3838 4624 3839 4628
rect 3843 4624 3844 4628
rect 3848 4624 3849 4628
rect 3853 4624 4235 4628
rect 4239 4624 4240 4628
rect 4244 4624 4245 4628
rect 4249 4624 4250 4628
rect 4254 4624 4264 4628
rect 4268 4624 4269 4628
rect 4273 4624 4274 4628
rect 4278 4624 4279 4628
rect 4283 4624 4293 4628
rect 4297 4624 4298 4628
rect 4302 4624 4303 4628
rect 4307 4624 4308 4628
rect 4312 4624 4322 4628
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4336 4624 4337 4628
rect 4341 4624 4351 4628
rect 4355 4624 4356 4628
rect 4360 4624 4361 4628
rect 4365 4624 4366 4628
rect 4370 4624 4518 4628
rect 654 4623 4518 4624
rect 654 4619 1820 4623
rect 1824 4619 1825 4623
rect 1829 4619 3674 4623
rect 3678 4619 3679 4623
rect 3683 4619 4518 4623
rect 654 4618 4518 4619
rect 654 4614 757 4618
rect 761 4614 762 4618
rect 766 4614 767 4618
rect 771 4614 772 4618
rect 776 4614 783 4618
rect 787 4614 788 4618
rect 792 4614 793 4618
rect 797 4614 798 4618
rect 802 4614 809 4618
rect 813 4614 814 4618
rect 818 4614 819 4618
rect 823 4614 824 4618
rect 828 4614 835 4618
rect 839 4614 840 4618
rect 844 4614 845 4618
rect 849 4614 850 4618
rect 854 4614 861 4618
rect 865 4614 866 4618
rect 870 4614 871 4618
rect 875 4614 876 4618
rect 880 4614 1053 4618
rect 1057 4614 1058 4618
rect 1062 4614 1063 4618
rect 1067 4614 1068 4618
rect 1072 4614 1362 4618
rect 1366 4614 1367 4618
rect 1371 4614 1372 4618
rect 1376 4614 1377 4618
rect 1381 4614 1671 4618
rect 1675 4614 1676 4618
rect 1680 4614 1681 4618
rect 1685 4614 1686 4618
rect 1690 4614 1820 4618
rect 1824 4614 1825 4618
rect 1829 4614 1980 4618
rect 1984 4614 1985 4618
rect 1989 4614 1990 4618
rect 1994 4614 1995 4618
rect 1999 4614 2289 4618
rect 2293 4614 2294 4618
rect 2298 4614 2299 4618
rect 2303 4614 2304 4618
rect 2308 4614 2598 4618
rect 2602 4614 2603 4618
rect 2607 4614 2608 4618
rect 2612 4614 2613 4618
rect 2617 4614 2907 4618
rect 2911 4614 2912 4618
rect 2916 4614 2917 4618
rect 2921 4614 2922 4618
rect 2926 4614 3216 4618
rect 3220 4614 3221 4618
rect 3225 4614 3226 4618
rect 3230 4614 3231 4618
rect 3235 4614 3525 4618
rect 3529 4614 3530 4618
rect 3534 4614 3535 4618
rect 3539 4614 3540 4618
rect 3544 4614 3674 4618
rect 3678 4614 3679 4618
rect 3683 4614 3834 4618
rect 3838 4614 3839 4618
rect 3843 4614 3844 4618
rect 3848 4614 3849 4618
rect 3853 4614 4235 4618
rect 4239 4614 4240 4618
rect 4244 4614 4245 4618
rect 4249 4614 4250 4618
rect 4254 4614 4264 4618
rect 4268 4614 4269 4618
rect 4273 4614 4274 4618
rect 4278 4614 4279 4618
rect 4283 4614 4293 4618
rect 4297 4614 4298 4618
rect 4302 4614 4303 4618
rect 4307 4614 4308 4618
rect 4312 4614 4322 4618
rect 4326 4614 4327 4618
rect 4331 4614 4332 4618
rect 4336 4614 4337 4618
rect 4341 4614 4351 4618
rect 4355 4614 4356 4618
rect 4360 4614 4361 4618
rect 4365 4614 4366 4618
rect 4370 4614 4518 4618
rect 654 4613 4518 4614
rect 654 4611 1820 4613
rect 654 4608 1077 4611
rect 654 4604 757 4608
rect 761 4604 762 4608
rect 766 4604 767 4608
rect 771 4604 772 4608
rect 776 4604 783 4608
rect 787 4604 788 4608
rect 792 4604 793 4608
rect 797 4604 798 4608
rect 802 4604 809 4608
rect 813 4604 814 4608
rect 818 4604 819 4608
rect 823 4604 824 4608
rect 828 4604 835 4608
rect 839 4604 840 4608
rect 844 4604 845 4608
rect 849 4604 850 4608
rect 854 4604 861 4608
rect 865 4604 866 4608
rect 870 4604 871 4608
rect 875 4604 876 4608
rect 880 4604 1053 4608
rect 1057 4604 1058 4608
rect 1062 4604 1063 4608
rect 1067 4604 1068 4608
rect 1072 4607 1077 4608
rect 1081 4607 1082 4611
rect 1086 4607 1087 4611
rect 1091 4607 1092 4611
rect 1096 4607 1097 4611
rect 1101 4607 1102 4611
rect 1106 4607 1107 4611
rect 1111 4607 1112 4611
rect 1116 4607 1117 4611
rect 1121 4607 1122 4611
rect 1126 4607 1127 4611
rect 1131 4607 1249 4611
rect 1253 4607 1254 4611
rect 1258 4607 1259 4611
rect 1263 4607 1264 4611
rect 1268 4607 1269 4611
rect 1273 4607 1274 4611
rect 1278 4607 1279 4611
rect 1283 4607 1284 4611
rect 1288 4607 1289 4611
rect 1293 4607 1294 4611
rect 1298 4607 1299 4611
rect 1303 4607 1304 4611
rect 1308 4607 1309 4611
rect 1313 4608 1386 4611
rect 1313 4607 1362 4608
rect 1072 4606 1362 4607
rect 1072 4604 1077 4606
rect 654 4602 1077 4604
rect 1081 4602 1082 4606
rect 1086 4602 1087 4606
rect 1091 4602 1092 4606
rect 1096 4602 1097 4606
rect 1101 4602 1102 4606
rect 1106 4602 1107 4606
rect 1111 4602 1112 4606
rect 1116 4602 1117 4606
rect 1121 4602 1122 4606
rect 1126 4602 1127 4606
rect 1131 4602 1249 4606
rect 1253 4602 1254 4606
rect 1258 4602 1259 4606
rect 1263 4602 1264 4606
rect 1268 4602 1269 4606
rect 1273 4602 1274 4606
rect 1278 4602 1279 4606
rect 1283 4602 1284 4606
rect 1288 4602 1289 4606
rect 1293 4602 1294 4606
rect 1298 4602 1299 4606
rect 1303 4602 1304 4606
rect 1308 4602 1309 4606
rect 1313 4604 1362 4606
rect 1366 4604 1367 4608
rect 1371 4604 1372 4608
rect 1376 4604 1377 4608
rect 1381 4607 1386 4608
rect 1390 4607 1391 4611
rect 1395 4607 1396 4611
rect 1400 4607 1401 4611
rect 1405 4607 1406 4611
rect 1410 4607 1411 4611
rect 1415 4607 1416 4611
rect 1420 4607 1421 4611
rect 1425 4607 1426 4611
rect 1430 4607 1431 4611
rect 1435 4607 1436 4611
rect 1440 4607 1558 4611
rect 1562 4607 1563 4611
rect 1567 4607 1568 4611
rect 1572 4607 1573 4611
rect 1577 4607 1578 4611
rect 1582 4607 1583 4611
rect 1587 4607 1588 4611
rect 1592 4607 1593 4611
rect 1597 4607 1598 4611
rect 1602 4607 1603 4611
rect 1607 4607 1608 4611
rect 1612 4607 1613 4611
rect 1617 4607 1618 4611
rect 1622 4608 1695 4611
rect 1622 4607 1671 4608
rect 1381 4606 1671 4607
rect 1381 4604 1386 4606
rect 1313 4602 1386 4604
rect 1390 4602 1391 4606
rect 1395 4602 1396 4606
rect 1400 4602 1401 4606
rect 1405 4602 1406 4606
rect 1410 4602 1411 4606
rect 1415 4602 1416 4606
rect 1420 4602 1421 4606
rect 1425 4602 1426 4606
rect 1430 4602 1431 4606
rect 1435 4602 1436 4606
rect 1440 4602 1558 4606
rect 1562 4602 1563 4606
rect 1567 4602 1568 4606
rect 1572 4602 1573 4606
rect 1577 4602 1578 4606
rect 1582 4602 1583 4606
rect 1587 4602 1588 4606
rect 1592 4602 1593 4606
rect 1597 4602 1598 4606
rect 1602 4602 1603 4606
rect 1607 4602 1608 4606
rect 1612 4602 1613 4606
rect 1617 4602 1618 4606
rect 1622 4604 1671 4606
rect 1675 4604 1676 4608
rect 1680 4604 1681 4608
rect 1685 4604 1686 4608
rect 1690 4607 1695 4608
rect 1699 4607 1700 4611
rect 1704 4607 1705 4611
rect 1709 4607 1710 4611
rect 1714 4607 1715 4611
rect 1719 4607 1720 4611
rect 1724 4607 1725 4611
rect 1729 4607 1730 4611
rect 1734 4607 1735 4611
rect 1739 4607 1740 4611
rect 1744 4607 1745 4611
rect 1749 4609 1820 4611
rect 1824 4609 1825 4613
rect 1829 4611 3674 4613
rect 1829 4609 1867 4611
rect 1749 4608 1867 4609
rect 1749 4607 1820 4608
rect 1690 4606 1820 4607
rect 1690 4604 1695 4606
rect 1622 4602 1695 4604
rect 1699 4602 1700 4606
rect 1704 4602 1705 4606
rect 1709 4602 1710 4606
rect 1714 4602 1715 4606
rect 1719 4602 1720 4606
rect 1724 4602 1725 4606
rect 1729 4602 1730 4606
rect 1734 4602 1735 4606
rect 1739 4602 1740 4606
rect 1744 4602 1745 4606
rect 1749 4604 1820 4606
rect 1824 4604 1825 4608
rect 1829 4607 1867 4608
rect 1871 4607 1872 4611
rect 1876 4607 1877 4611
rect 1881 4607 1882 4611
rect 1886 4607 1887 4611
rect 1891 4607 1892 4611
rect 1896 4607 1897 4611
rect 1901 4607 1902 4611
rect 1906 4607 1907 4611
rect 1911 4607 1912 4611
rect 1916 4607 1917 4611
rect 1921 4607 1922 4611
rect 1926 4607 1927 4611
rect 1931 4608 2004 4611
rect 1931 4607 1980 4608
rect 1829 4606 1980 4607
rect 1829 4604 1867 4606
rect 1749 4603 1867 4604
rect 1749 4602 1820 4603
rect 654 4599 1820 4602
rect 1824 4599 1825 4603
rect 1829 4602 1867 4603
rect 1871 4602 1872 4606
rect 1876 4602 1877 4606
rect 1881 4602 1882 4606
rect 1886 4602 1887 4606
rect 1891 4602 1892 4606
rect 1896 4602 1897 4606
rect 1901 4602 1902 4606
rect 1906 4602 1907 4606
rect 1911 4602 1912 4606
rect 1916 4602 1917 4606
rect 1921 4602 1922 4606
rect 1926 4602 1927 4606
rect 1931 4604 1980 4606
rect 1984 4604 1985 4608
rect 1989 4604 1990 4608
rect 1994 4604 1995 4608
rect 1999 4607 2004 4608
rect 2008 4607 2009 4611
rect 2013 4607 2014 4611
rect 2018 4607 2019 4611
rect 2023 4607 2024 4611
rect 2028 4607 2029 4611
rect 2033 4607 2034 4611
rect 2038 4607 2039 4611
rect 2043 4607 2044 4611
rect 2048 4607 2049 4611
rect 2053 4607 2054 4611
rect 2058 4607 2176 4611
rect 2180 4607 2181 4611
rect 2185 4607 2186 4611
rect 2190 4607 2191 4611
rect 2195 4607 2196 4611
rect 2200 4607 2201 4611
rect 2205 4607 2206 4611
rect 2210 4607 2211 4611
rect 2215 4607 2216 4611
rect 2220 4607 2221 4611
rect 2225 4607 2226 4611
rect 2230 4607 2231 4611
rect 2235 4607 2236 4611
rect 2240 4608 2313 4611
rect 2240 4607 2289 4608
rect 1999 4606 2289 4607
rect 1999 4604 2004 4606
rect 1931 4602 2004 4604
rect 2008 4602 2009 4606
rect 2013 4602 2014 4606
rect 2018 4602 2019 4606
rect 2023 4602 2024 4606
rect 2028 4602 2029 4606
rect 2033 4602 2034 4606
rect 2038 4602 2039 4606
rect 2043 4602 2044 4606
rect 2048 4602 2049 4606
rect 2053 4602 2054 4606
rect 2058 4602 2176 4606
rect 2180 4602 2181 4606
rect 2185 4602 2186 4606
rect 2190 4602 2191 4606
rect 2195 4602 2196 4606
rect 2200 4602 2201 4606
rect 2205 4602 2206 4606
rect 2210 4602 2211 4606
rect 2215 4602 2216 4606
rect 2220 4602 2221 4606
rect 2225 4602 2226 4606
rect 2230 4602 2231 4606
rect 2235 4602 2236 4606
rect 2240 4604 2289 4606
rect 2293 4604 2294 4608
rect 2298 4604 2299 4608
rect 2303 4604 2304 4608
rect 2308 4607 2313 4608
rect 2317 4607 2318 4611
rect 2322 4607 2323 4611
rect 2327 4607 2328 4611
rect 2332 4607 2333 4611
rect 2337 4607 2338 4611
rect 2342 4607 2343 4611
rect 2347 4607 2348 4611
rect 2352 4607 2353 4611
rect 2357 4607 2358 4611
rect 2362 4607 2363 4611
rect 2367 4607 2485 4611
rect 2489 4607 2490 4611
rect 2494 4607 2495 4611
rect 2499 4607 2500 4611
rect 2504 4607 2505 4611
rect 2509 4607 2510 4611
rect 2514 4607 2515 4611
rect 2519 4607 2520 4611
rect 2524 4607 2525 4611
rect 2529 4607 2530 4611
rect 2534 4607 2535 4611
rect 2539 4607 2540 4611
rect 2544 4607 2545 4611
rect 2549 4608 2622 4611
rect 2549 4607 2598 4608
rect 2308 4606 2598 4607
rect 2308 4604 2313 4606
rect 2240 4602 2313 4604
rect 2317 4602 2318 4606
rect 2322 4602 2323 4606
rect 2327 4602 2328 4606
rect 2332 4602 2333 4606
rect 2337 4602 2338 4606
rect 2342 4602 2343 4606
rect 2347 4602 2348 4606
rect 2352 4602 2353 4606
rect 2357 4602 2358 4606
rect 2362 4602 2363 4606
rect 2367 4602 2485 4606
rect 2489 4602 2490 4606
rect 2494 4602 2495 4606
rect 2499 4602 2500 4606
rect 2504 4602 2505 4606
rect 2509 4602 2510 4606
rect 2514 4602 2515 4606
rect 2519 4602 2520 4606
rect 2524 4602 2525 4606
rect 2529 4602 2530 4606
rect 2534 4602 2535 4606
rect 2539 4602 2540 4606
rect 2544 4602 2545 4606
rect 2549 4604 2598 4606
rect 2602 4604 2603 4608
rect 2607 4604 2608 4608
rect 2612 4604 2613 4608
rect 2617 4607 2622 4608
rect 2626 4607 2627 4611
rect 2631 4607 2632 4611
rect 2636 4607 2637 4611
rect 2641 4607 2642 4611
rect 2646 4607 2647 4611
rect 2651 4607 2652 4611
rect 2656 4607 2657 4611
rect 2661 4607 2662 4611
rect 2666 4607 2667 4611
rect 2671 4607 2672 4611
rect 2676 4607 2794 4611
rect 2798 4607 2799 4611
rect 2803 4607 2804 4611
rect 2808 4607 2809 4611
rect 2813 4607 2814 4611
rect 2818 4607 2819 4611
rect 2823 4607 2824 4611
rect 2828 4607 2829 4611
rect 2833 4607 2834 4611
rect 2838 4607 2839 4611
rect 2843 4607 2844 4611
rect 2848 4607 2849 4611
rect 2853 4607 2854 4611
rect 2858 4608 2931 4611
rect 2858 4607 2907 4608
rect 2617 4606 2907 4607
rect 2617 4604 2622 4606
rect 2549 4602 2622 4604
rect 2626 4602 2627 4606
rect 2631 4602 2632 4606
rect 2636 4602 2637 4606
rect 2641 4602 2642 4606
rect 2646 4602 2647 4606
rect 2651 4602 2652 4606
rect 2656 4602 2657 4606
rect 2661 4602 2662 4606
rect 2666 4602 2667 4606
rect 2671 4602 2672 4606
rect 2676 4602 2794 4606
rect 2798 4602 2799 4606
rect 2803 4602 2804 4606
rect 2808 4602 2809 4606
rect 2813 4602 2814 4606
rect 2818 4602 2819 4606
rect 2823 4602 2824 4606
rect 2828 4602 2829 4606
rect 2833 4602 2834 4606
rect 2838 4602 2839 4606
rect 2843 4602 2844 4606
rect 2848 4602 2849 4606
rect 2853 4602 2854 4606
rect 2858 4604 2907 4606
rect 2911 4604 2912 4608
rect 2916 4604 2917 4608
rect 2921 4604 2922 4608
rect 2926 4607 2931 4608
rect 2935 4607 2936 4611
rect 2940 4607 2941 4611
rect 2945 4607 2946 4611
rect 2950 4607 2951 4611
rect 2955 4607 2956 4611
rect 2960 4607 2961 4611
rect 2965 4607 2966 4611
rect 2970 4607 2971 4611
rect 2975 4607 2976 4611
rect 2980 4607 2981 4611
rect 2985 4607 3103 4611
rect 3107 4607 3108 4611
rect 3112 4607 3113 4611
rect 3117 4607 3118 4611
rect 3122 4607 3123 4611
rect 3127 4607 3128 4611
rect 3132 4607 3133 4611
rect 3137 4607 3138 4611
rect 3142 4607 3143 4611
rect 3147 4607 3148 4611
rect 3152 4607 3153 4611
rect 3157 4607 3158 4611
rect 3162 4607 3163 4611
rect 3167 4608 3240 4611
rect 3167 4607 3216 4608
rect 2926 4606 3216 4607
rect 2926 4604 2931 4606
rect 2858 4602 2931 4604
rect 2935 4602 2936 4606
rect 2940 4602 2941 4606
rect 2945 4602 2946 4606
rect 2950 4602 2951 4606
rect 2955 4602 2956 4606
rect 2960 4602 2961 4606
rect 2965 4602 2966 4606
rect 2970 4602 2971 4606
rect 2975 4602 2976 4606
rect 2980 4602 2981 4606
rect 2985 4602 3103 4606
rect 3107 4602 3108 4606
rect 3112 4602 3113 4606
rect 3117 4602 3118 4606
rect 3122 4602 3123 4606
rect 3127 4602 3128 4606
rect 3132 4602 3133 4606
rect 3137 4602 3138 4606
rect 3142 4602 3143 4606
rect 3147 4602 3148 4606
rect 3152 4602 3153 4606
rect 3157 4602 3158 4606
rect 3162 4602 3163 4606
rect 3167 4604 3216 4606
rect 3220 4604 3221 4608
rect 3225 4604 3226 4608
rect 3230 4604 3231 4608
rect 3235 4607 3240 4608
rect 3244 4607 3245 4611
rect 3249 4607 3250 4611
rect 3254 4607 3255 4611
rect 3259 4607 3260 4611
rect 3264 4607 3265 4611
rect 3269 4607 3270 4611
rect 3274 4607 3275 4611
rect 3279 4607 3280 4611
rect 3284 4607 3285 4611
rect 3289 4607 3290 4611
rect 3294 4607 3412 4611
rect 3416 4607 3417 4611
rect 3421 4607 3422 4611
rect 3426 4607 3427 4611
rect 3431 4607 3432 4611
rect 3436 4607 3437 4611
rect 3441 4607 3442 4611
rect 3446 4607 3447 4611
rect 3451 4607 3452 4611
rect 3456 4607 3457 4611
rect 3461 4607 3462 4611
rect 3466 4607 3467 4611
rect 3471 4607 3472 4611
rect 3476 4608 3549 4611
rect 3476 4607 3525 4608
rect 3235 4606 3525 4607
rect 3235 4604 3240 4606
rect 3167 4602 3240 4604
rect 3244 4602 3245 4606
rect 3249 4602 3250 4606
rect 3254 4602 3255 4606
rect 3259 4602 3260 4606
rect 3264 4602 3265 4606
rect 3269 4602 3270 4606
rect 3274 4602 3275 4606
rect 3279 4602 3280 4606
rect 3284 4602 3285 4606
rect 3289 4602 3290 4606
rect 3294 4602 3412 4606
rect 3416 4602 3417 4606
rect 3421 4602 3422 4606
rect 3426 4602 3427 4606
rect 3431 4602 3432 4606
rect 3436 4602 3437 4606
rect 3441 4602 3442 4606
rect 3446 4602 3447 4606
rect 3451 4602 3452 4606
rect 3456 4602 3457 4606
rect 3461 4602 3462 4606
rect 3466 4602 3467 4606
rect 3471 4602 3472 4606
rect 3476 4604 3525 4606
rect 3529 4604 3530 4608
rect 3534 4604 3535 4608
rect 3539 4604 3540 4608
rect 3544 4607 3549 4608
rect 3553 4607 3554 4611
rect 3558 4607 3559 4611
rect 3563 4607 3564 4611
rect 3568 4607 3569 4611
rect 3573 4607 3574 4611
rect 3578 4607 3579 4611
rect 3583 4607 3584 4611
rect 3588 4607 3589 4611
rect 3593 4607 3594 4611
rect 3598 4607 3599 4611
rect 3603 4609 3674 4611
rect 3678 4609 3679 4613
rect 3683 4611 4518 4613
rect 3683 4609 3721 4611
rect 3603 4608 3721 4609
rect 3603 4607 3674 4608
rect 3544 4606 3674 4607
rect 3544 4604 3549 4606
rect 3476 4602 3549 4604
rect 3553 4602 3554 4606
rect 3558 4602 3559 4606
rect 3563 4602 3564 4606
rect 3568 4602 3569 4606
rect 3573 4602 3574 4606
rect 3578 4602 3579 4606
rect 3583 4602 3584 4606
rect 3588 4602 3589 4606
rect 3593 4602 3594 4606
rect 3598 4602 3599 4606
rect 3603 4604 3674 4606
rect 3678 4604 3679 4608
rect 3683 4607 3721 4608
rect 3725 4607 3726 4611
rect 3730 4607 3731 4611
rect 3735 4607 3736 4611
rect 3740 4607 3741 4611
rect 3745 4607 3746 4611
rect 3750 4607 3751 4611
rect 3755 4607 3756 4611
rect 3760 4607 3761 4611
rect 3765 4607 3766 4611
rect 3770 4607 3771 4611
rect 3775 4607 3776 4611
rect 3780 4607 3781 4611
rect 3785 4608 4518 4611
rect 3785 4607 3834 4608
rect 3683 4606 3834 4607
rect 3683 4604 3721 4606
rect 3603 4603 3721 4604
rect 3603 4602 3674 4603
rect 1829 4599 3674 4602
rect 3678 4599 3679 4603
rect 3683 4602 3721 4603
rect 3725 4602 3726 4606
rect 3730 4602 3731 4606
rect 3735 4602 3736 4606
rect 3740 4602 3741 4606
rect 3745 4602 3746 4606
rect 3750 4602 3751 4606
rect 3755 4602 3756 4606
rect 3760 4602 3761 4606
rect 3765 4602 3766 4606
rect 3770 4602 3771 4606
rect 3775 4602 3776 4606
rect 3780 4602 3781 4606
rect 3785 4604 3834 4606
rect 3838 4604 3839 4608
rect 3843 4604 3844 4608
rect 3848 4604 3849 4608
rect 3853 4604 4235 4608
rect 4239 4604 4240 4608
rect 4244 4604 4245 4608
rect 4249 4604 4250 4608
rect 4254 4604 4264 4608
rect 4268 4604 4269 4608
rect 4273 4604 4274 4608
rect 4278 4604 4279 4608
rect 4283 4604 4293 4608
rect 4297 4604 4298 4608
rect 4302 4604 4303 4608
rect 4307 4604 4308 4608
rect 4312 4604 4322 4608
rect 4326 4604 4327 4608
rect 4331 4604 4332 4608
rect 4336 4604 4337 4608
rect 4341 4604 4351 4608
rect 4355 4604 4356 4608
rect 4360 4604 4361 4608
rect 4365 4604 4366 4608
rect 4370 4604 4518 4608
rect 3785 4602 4518 4604
rect 3683 4599 4518 4602
rect 654 4598 4518 4599
rect 654 4594 757 4598
rect 761 4594 762 4598
rect 766 4594 767 4598
rect 771 4594 772 4598
rect 776 4594 783 4598
rect 787 4594 788 4598
rect 792 4594 793 4598
rect 797 4594 798 4598
rect 802 4594 809 4598
rect 813 4594 814 4598
rect 818 4594 819 4598
rect 823 4594 824 4598
rect 828 4594 835 4598
rect 839 4594 840 4598
rect 844 4594 845 4598
rect 849 4594 850 4598
rect 854 4594 861 4598
rect 865 4594 866 4598
rect 870 4594 871 4598
rect 875 4594 876 4598
rect 880 4594 1053 4598
rect 1057 4594 1058 4598
rect 1062 4594 1063 4598
rect 1067 4594 1068 4598
rect 1072 4594 1362 4598
rect 1366 4594 1367 4598
rect 1371 4594 1372 4598
rect 1376 4594 1377 4598
rect 1381 4594 1671 4598
rect 1675 4594 1676 4598
rect 1680 4594 1681 4598
rect 1685 4594 1686 4598
rect 1690 4594 1980 4598
rect 1984 4594 1985 4598
rect 1989 4594 1990 4598
rect 1994 4594 1995 4598
rect 1999 4594 2289 4598
rect 2293 4594 2294 4598
rect 2298 4594 2299 4598
rect 2303 4594 2304 4598
rect 2308 4594 2598 4598
rect 2602 4594 2603 4598
rect 2607 4594 2608 4598
rect 2612 4594 2613 4598
rect 2617 4594 2907 4598
rect 2911 4594 2912 4598
rect 2916 4594 2917 4598
rect 2921 4594 2922 4598
rect 2926 4594 3216 4598
rect 3220 4594 3221 4598
rect 3225 4594 3226 4598
rect 3230 4594 3231 4598
rect 3235 4594 3525 4598
rect 3529 4594 3530 4598
rect 3534 4594 3535 4598
rect 3539 4594 3540 4598
rect 3544 4594 3834 4598
rect 3838 4594 3839 4598
rect 3843 4594 3844 4598
rect 3848 4594 3849 4598
rect 3853 4594 4235 4598
rect 4239 4594 4240 4598
rect 4244 4594 4245 4598
rect 4249 4594 4250 4598
rect 4254 4594 4264 4598
rect 4268 4594 4269 4598
rect 4273 4594 4274 4598
rect 4278 4594 4279 4598
rect 4283 4594 4293 4598
rect 4297 4594 4298 4598
rect 4302 4594 4303 4598
rect 4307 4594 4308 4598
rect 4312 4594 4322 4598
rect 4326 4594 4327 4598
rect 4331 4594 4332 4598
rect 4336 4594 4337 4598
rect 4341 4594 4351 4598
rect 4355 4594 4356 4598
rect 4360 4594 4361 4598
rect 4365 4594 4366 4598
rect 4370 4594 4518 4598
rect 654 4589 4518 4594
rect 4522 9577 4602 9729
rect 4522 9573 4525 9577
rect 4529 9573 4535 9577
rect 4539 9573 4545 9577
rect 4549 9573 4555 9577
rect 4559 9573 4602 9577
rect 4522 9572 4602 9573
rect 4522 9568 4525 9572
rect 4529 9568 4535 9572
rect 4539 9568 4545 9572
rect 4549 9568 4555 9572
rect 4559 9568 4602 9572
rect 4522 9567 4602 9568
rect 4522 9563 4525 9567
rect 4529 9563 4535 9567
rect 4539 9563 4545 9567
rect 4549 9563 4555 9567
rect 4559 9563 4602 9567
rect 4522 9562 4602 9563
rect 4522 9558 4525 9562
rect 4529 9558 4535 9562
rect 4539 9558 4545 9562
rect 4549 9558 4555 9562
rect 4559 9558 4602 9562
rect 4522 9548 4602 9558
rect 4522 9544 4525 9548
rect 4529 9544 4535 9548
rect 4539 9544 4545 9548
rect 4549 9544 4555 9548
rect 4559 9544 4602 9548
rect 4522 9543 4602 9544
rect 4522 9539 4525 9543
rect 4529 9539 4535 9543
rect 4539 9539 4545 9543
rect 4549 9539 4555 9543
rect 4559 9539 4602 9543
rect 4522 9538 4602 9539
rect 4522 9534 4525 9538
rect 4529 9534 4535 9538
rect 4539 9534 4545 9538
rect 4549 9534 4555 9538
rect 4559 9534 4602 9538
rect 4522 9533 4602 9534
rect 4522 9529 4525 9533
rect 4529 9529 4535 9533
rect 4539 9529 4545 9533
rect 4549 9529 4555 9533
rect 4559 9529 4602 9533
rect 4522 9519 4602 9529
rect 4522 9515 4525 9519
rect 4529 9515 4535 9519
rect 4539 9515 4545 9519
rect 4549 9515 4555 9519
rect 4559 9515 4602 9519
rect 4522 9514 4602 9515
rect 4522 9510 4525 9514
rect 4529 9510 4535 9514
rect 4539 9510 4545 9514
rect 4549 9510 4555 9514
rect 4559 9510 4602 9514
rect 4522 9509 4602 9510
rect 4522 9505 4525 9509
rect 4529 9505 4535 9509
rect 4539 9505 4545 9509
rect 4549 9505 4555 9509
rect 4559 9505 4602 9509
rect 4522 9504 4602 9505
rect 4522 9500 4525 9504
rect 4529 9500 4535 9504
rect 4539 9500 4545 9504
rect 4549 9500 4555 9504
rect 4559 9500 4602 9504
rect 4522 9490 4602 9500
rect 4522 9486 4525 9490
rect 4529 9486 4535 9490
rect 4539 9486 4545 9490
rect 4549 9486 4555 9490
rect 4559 9486 4602 9490
rect 4522 9485 4602 9486
rect 4522 9481 4525 9485
rect 4529 9481 4535 9485
rect 4539 9481 4545 9485
rect 4549 9481 4555 9485
rect 4559 9481 4602 9485
rect 4522 9480 4602 9481
rect 4522 9476 4525 9480
rect 4529 9476 4535 9480
rect 4539 9476 4545 9480
rect 4549 9476 4555 9480
rect 4559 9476 4602 9480
rect 4522 9475 4602 9476
rect 4522 9471 4525 9475
rect 4529 9471 4535 9475
rect 4539 9471 4545 9475
rect 4549 9471 4555 9475
rect 4559 9471 4602 9475
rect 4522 9461 4602 9471
rect 4522 9457 4525 9461
rect 4529 9457 4535 9461
rect 4539 9457 4545 9461
rect 4549 9457 4555 9461
rect 4559 9457 4602 9461
rect 4522 9456 4602 9457
rect 4522 9452 4525 9456
rect 4529 9452 4535 9456
rect 4539 9452 4545 9456
rect 4549 9452 4555 9456
rect 4559 9452 4602 9456
rect 4522 9451 4602 9452
rect 4522 9447 4525 9451
rect 4529 9447 4535 9451
rect 4539 9447 4545 9451
rect 4549 9447 4555 9451
rect 4559 9447 4602 9451
rect 4522 9446 4602 9447
rect 4522 9442 4525 9446
rect 4529 9442 4535 9446
rect 4539 9442 4545 9446
rect 4549 9442 4555 9446
rect 4559 9442 4602 9446
rect 4522 9060 4602 9442
rect 4522 9056 4525 9060
rect 4529 9056 4535 9060
rect 4539 9056 4545 9060
rect 4549 9056 4555 9060
rect 4559 9056 4602 9060
rect 4522 9055 4602 9056
rect 4522 9051 4525 9055
rect 4529 9051 4535 9055
rect 4539 9051 4545 9055
rect 4549 9051 4555 9055
rect 4559 9051 4602 9055
rect 4522 9050 4602 9051
rect 4522 9046 4525 9050
rect 4529 9046 4535 9050
rect 4539 9046 4545 9050
rect 4549 9046 4555 9050
rect 4559 9046 4602 9050
rect 4522 9045 4602 9046
rect 4522 9041 4525 9045
rect 4529 9041 4535 9045
rect 4539 9041 4545 9045
rect 4549 9041 4555 9045
rect 4559 9041 4602 9045
rect 4522 8751 4602 9041
rect 4522 8747 4525 8751
rect 4529 8747 4535 8751
rect 4539 8747 4545 8751
rect 4549 8747 4555 8751
rect 4559 8747 4602 8751
rect 4522 8746 4602 8747
rect 4522 8742 4525 8746
rect 4529 8742 4535 8746
rect 4539 8742 4545 8746
rect 4549 8742 4555 8746
rect 4559 8742 4602 8746
rect 4522 8741 4602 8742
rect 4522 8737 4525 8741
rect 4529 8737 4535 8741
rect 4539 8737 4545 8741
rect 4549 8737 4555 8741
rect 4559 8737 4602 8741
rect 4522 8736 4602 8737
rect 4522 8732 4525 8736
rect 4529 8732 4535 8736
rect 4539 8732 4545 8736
rect 4549 8732 4555 8736
rect 4559 8732 4602 8736
rect 4522 8442 4602 8732
rect 4522 8438 4525 8442
rect 4529 8438 4535 8442
rect 4539 8438 4545 8442
rect 4549 8438 4555 8442
rect 4559 8438 4602 8442
rect 4522 8437 4602 8438
rect 4522 8433 4525 8437
rect 4529 8433 4535 8437
rect 4539 8433 4545 8437
rect 4549 8433 4555 8437
rect 4559 8433 4602 8437
rect 4522 8432 4602 8433
rect 4522 8428 4525 8432
rect 4529 8428 4535 8432
rect 4539 8428 4545 8432
rect 4549 8428 4555 8432
rect 4559 8428 4602 8432
rect 4522 8427 4602 8428
rect 4522 8423 4525 8427
rect 4529 8423 4535 8427
rect 4539 8423 4545 8427
rect 4549 8423 4555 8427
rect 4559 8423 4602 8427
rect 4522 8133 4602 8423
rect 4522 8129 4525 8133
rect 4529 8129 4535 8133
rect 4539 8129 4545 8133
rect 4549 8129 4555 8133
rect 4559 8129 4602 8133
rect 4522 8128 4602 8129
rect 4522 8124 4525 8128
rect 4529 8124 4535 8128
rect 4539 8124 4545 8128
rect 4549 8124 4555 8128
rect 4559 8124 4602 8128
rect 4522 8123 4602 8124
rect 4522 8119 4525 8123
rect 4529 8119 4535 8123
rect 4539 8119 4545 8123
rect 4549 8119 4555 8123
rect 4559 8119 4602 8123
rect 4522 8118 4602 8119
rect 4522 8114 4525 8118
rect 4529 8114 4535 8118
rect 4539 8114 4545 8118
rect 4549 8114 4555 8118
rect 4559 8114 4602 8118
rect 4522 8102 4602 8114
rect 4522 8098 4525 8102
rect 4529 8098 4535 8102
rect 4539 8098 4545 8102
rect 4549 8098 4555 8102
rect 4559 8098 4602 8102
rect 4522 8097 4602 8098
rect 4522 8093 4525 8097
rect 4529 8093 4535 8097
rect 4539 8093 4545 8097
rect 4549 8093 4555 8097
rect 4559 8093 4602 8097
rect 4522 8092 4602 8093
rect 4522 8088 4525 8092
rect 4529 8088 4535 8092
rect 4539 8088 4545 8092
rect 4549 8088 4555 8092
rect 4559 8088 4602 8092
rect 4522 8087 4602 8088
rect 4522 8083 4525 8087
rect 4529 8083 4535 8087
rect 4539 8083 4545 8087
rect 4549 8083 4555 8087
rect 4559 8083 4602 8087
rect 4522 7818 4602 8083
rect 4522 7814 4529 7818
rect 4533 7814 4534 7818
rect 4538 7814 4539 7818
rect 4543 7814 4544 7818
rect 4548 7814 4549 7818
rect 4553 7814 4554 7818
rect 4558 7814 4559 7818
rect 4563 7814 4564 7818
rect 4568 7814 4569 7818
rect 4573 7814 4574 7818
rect 4578 7814 4579 7818
rect 4583 7814 4584 7818
rect 4588 7814 4589 7818
rect 4593 7814 4602 7818
rect 4522 7813 4602 7814
rect 4522 7809 4529 7813
rect 4533 7809 4534 7813
rect 4538 7809 4539 7813
rect 4543 7809 4544 7813
rect 4548 7809 4549 7813
rect 4553 7809 4554 7813
rect 4558 7809 4559 7813
rect 4563 7809 4564 7813
rect 4568 7809 4569 7813
rect 4573 7809 4574 7813
rect 4578 7809 4579 7813
rect 4583 7809 4584 7813
rect 4588 7809 4589 7813
rect 4593 7809 4602 7813
rect 4522 7793 4602 7809
rect 4522 7789 4525 7793
rect 4529 7789 4535 7793
rect 4539 7789 4545 7793
rect 4549 7789 4555 7793
rect 4559 7789 4602 7793
rect 4522 7788 4602 7789
rect 4522 7784 4525 7788
rect 4529 7784 4535 7788
rect 4539 7784 4545 7788
rect 4549 7784 4555 7788
rect 4559 7784 4602 7788
rect 4522 7783 4602 7784
rect 4522 7779 4525 7783
rect 4529 7779 4535 7783
rect 4539 7779 4545 7783
rect 4549 7779 4555 7783
rect 4559 7779 4602 7783
rect 4522 7778 4602 7779
rect 4522 7774 4525 7778
rect 4529 7774 4535 7778
rect 4539 7774 4545 7778
rect 4549 7774 4555 7778
rect 4559 7774 4602 7778
rect 4522 7503 4602 7774
rect 4522 7499 4529 7503
rect 4533 7499 4534 7503
rect 4538 7499 4539 7503
rect 4543 7499 4544 7503
rect 4548 7499 4549 7503
rect 4553 7499 4554 7503
rect 4558 7499 4559 7503
rect 4563 7499 4564 7503
rect 4568 7499 4569 7503
rect 4573 7499 4574 7503
rect 4578 7499 4579 7503
rect 4583 7499 4584 7503
rect 4588 7499 4589 7503
rect 4593 7499 4602 7503
rect 4522 7315 4602 7499
rect 4522 7311 4553 7315
rect 4557 7311 4558 7315
rect 4562 7311 4602 7315
rect 4522 7310 4602 7311
rect 4522 7306 4553 7310
rect 4557 7306 4558 7310
rect 4562 7306 4602 7310
rect 4522 7305 4602 7306
rect 4522 7301 4553 7305
rect 4557 7301 4558 7305
rect 4562 7301 4602 7305
rect 4522 7300 4602 7301
rect 4522 7296 4553 7300
rect 4557 7296 4558 7300
rect 4562 7296 4602 7300
rect 4522 7295 4602 7296
rect 4522 7291 4553 7295
rect 4557 7291 4558 7295
rect 4562 7291 4602 7295
rect 4522 7290 4602 7291
rect 4522 7286 4553 7290
rect 4557 7286 4558 7290
rect 4562 7286 4602 7290
rect 4522 7285 4602 7286
rect 4522 7281 4553 7285
rect 4557 7281 4558 7285
rect 4562 7281 4602 7285
rect 4522 7280 4602 7281
rect 4522 7276 4553 7280
rect 4557 7276 4558 7280
rect 4562 7276 4602 7280
rect 4522 7275 4602 7276
rect 4522 7271 4553 7275
rect 4557 7271 4558 7275
rect 4562 7271 4602 7275
rect 4522 7270 4602 7271
rect 4522 7266 4553 7270
rect 4557 7266 4558 7270
rect 4562 7266 4602 7270
rect 4522 7265 4602 7266
rect 4522 7261 4553 7265
rect 4557 7261 4558 7265
rect 4562 7261 4602 7265
rect 4522 7260 4602 7261
rect 4522 7256 4553 7260
rect 4557 7256 4558 7260
rect 4562 7256 4602 7260
rect 4522 7255 4602 7256
rect 4522 7251 4553 7255
rect 4557 7251 4558 7255
rect 4562 7251 4602 7255
rect 4522 7234 4602 7251
rect 4522 7230 4525 7234
rect 4529 7230 4535 7234
rect 4539 7230 4545 7234
rect 4549 7230 4555 7234
rect 4559 7230 4602 7234
rect 4522 7229 4602 7230
rect 4522 7225 4525 7229
rect 4529 7225 4535 7229
rect 4539 7225 4545 7229
rect 4549 7225 4555 7229
rect 4559 7225 4602 7229
rect 4522 7224 4602 7225
rect 4522 7220 4525 7224
rect 4529 7220 4535 7224
rect 4539 7220 4545 7224
rect 4549 7220 4555 7224
rect 4559 7220 4602 7224
rect 4522 7219 4602 7220
rect 4522 7215 4525 7219
rect 4529 7215 4535 7219
rect 4539 7215 4545 7219
rect 4549 7215 4555 7219
rect 4559 7215 4602 7219
rect 4522 7206 4602 7215
rect 4522 7202 4525 7206
rect 4529 7202 4535 7206
rect 4539 7202 4545 7206
rect 4549 7202 4555 7206
rect 4559 7202 4602 7206
rect 4522 7201 4602 7202
rect 4522 7197 4525 7201
rect 4529 7197 4535 7201
rect 4539 7197 4545 7201
rect 4549 7197 4555 7201
rect 4559 7197 4602 7201
rect 4522 7196 4602 7197
rect 4522 7192 4525 7196
rect 4529 7192 4535 7196
rect 4539 7192 4545 7196
rect 4549 7192 4555 7196
rect 4559 7192 4602 7196
rect 4522 7191 4602 7192
rect 4522 7187 4525 7191
rect 4529 7187 4535 7191
rect 4539 7187 4545 7191
rect 4549 7187 4555 7191
rect 4559 7187 4602 7191
rect 4522 7156 4602 7187
rect 4522 7152 4525 7156
rect 4529 7152 4535 7156
rect 4539 7152 4545 7156
rect 4549 7152 4555 7156
rect 4559 7152 4602 7156
rect 4522 6862 4602 7152
rect 4522 6858 4525 6862
rect 4529 6858 4535 6862
rect 4539 6858 4545 6862
rect 4549 6858 4555 6862
rect 4559 6858 4602 6862
rect 4522 6857 4602 6858
rect 4522 6853 4525 6857
rect 4529 6853 4535 6857
rect 4539 6853 4545 6857
rect 4549 6853 4555 6857
rect 4559 6853 4602 6857
rect 4522 6852 4602 6853
rect 4522 6848 4525 6852
rect 4529 6848 4535 6852
rect 4539 6848 4545 6852
rect 4549 6848 4555 6852
rect 4559 6848 4602 6852
rect 4522 6847 4602 6848
rect 4522 6843 4525 6847
rect 4529 6843 4535 6847
rect 4539 6843 4545 6847
rect 4549 6843 4555 6847
rect 4559 6843 4602 6847
rect 4522 6553 4602 6843
rect 4522 6549 4525 6553
rect 4529 6549 4535 6553
rect 4539 6549 4545 6553
rect 4549 6549 4555 6553
rect 4559 6549 4602 6553
rect 4522 6548 4602 6549
rect 4522 6544 4525 6548
rect 4529 6544 4535 6548
rect 4539 6544 4545 6548
rect 4549 6544 4555 6548
rect 4559 6544 4602 6548
rect 4522 6543 4602 6544
rect 4522 6539 4525 6543
rect 4529 6539 4535 6543
rect 4539 6539 4545 6543
rect 4549 6539 4555 6543
rect 4559 6539 4602 6543
rect 4522 6538 4602 6539
rect 4522 6534 4525 6538
rect 4529 6534 4535 6538
rect 4539 6534 4545 6538
rect 4549 6534 4555 6538
rect 4559 6534 4602 6538
rect 4522 6244 4602 6534
rect 4522 6240 4525 6244
rect 4529 6240 4535 6244
rect 4539 6240 4545 6244
rect 4549 6240 4555 6244
rect 4559 6240 4602 6244
rect 4522 6239 4602 6240
rect 4522 6235 4525 6239
rect 4529 6235 4535 6239
rect 4539 6235 4545 6239
rect 4549 6235 4555 6239
rect 4559 6235 4602 6239
rect 4522 6234 4602 6235
rect 4522 6230 4525 6234
rect 4529 6230 4535 6234
rect 4539 6230 4545 6234
rect 4549 6230 4555 6234
rect 4559 6230 4602 6234
rect 4522 6229 4602 6230
rect 4522 6225 4525 6229
rect 4529 6225 4535 6229
rect 4539 6225 4545 6229
rect 4549 6225 4555 6229
rect 4559 6225 4602 6229
rect 4522 5935 4602 6225
rect 4522 5931 4525 5935
rect 4529 5931 4535 5935
rect 4539 5931 4545 5935
rect 4549 5931 4555 5935
rect 4559 5931 4602 5935
rect 4522 5930 4602 5931
rect 4522 5926 4525 5930
rect 4529 5926 4535 5930
rect 4539 5926 4545 5930
rect 4549 5926 4555 5930
rect 4559 5926 4602 5930
rect 4522 5925 4602 5926
rect 4522 5921 4525 5925
rect 4529 5921 4535 5925
rect 4539 5921 4545 5925
rect 4549 5921 4555 5925
rect 4559 5921 4602 5925
rect 4522 5920 4602 5921
rect 4522 5916 4525 5920
rect 4529 5916 4535 5920
rect 4539 5916 4545 5920
rect 4549 5916 4555 5920
rect 4559 5916 4602 5920
rect 4522 5626 4602 5916
rect 4522 5622 4525 5626
rect 4529 5622 4535 5626
rect 4539 5622 4545 5626
rect 4549 5622 4555 5626
rect 4559 5622 4602 5626
rect 4522 5621 4602 5622
rect 4522 5617 4525 5621
rect 4529 5617 4535 5621
rect 4539 5617 4545 5621
rect 4549 5617 4555 5621
rect 4559 5617 4602 5621
rect 4522 5616 4602 5617
rect 4522 5612 4525 5616
rect 4529 5612 4535 5616
rect 4539 5612 4545 5616
rect 4549 5612 4555 5616
rect 4559 5612 4602 5616
rect 4522 5611 4602 5612
rect 4522 5607 4525 5611
rect 4529 5607 4535 5611
rect 4539 5607 4545 5611
rect 4549 5607 4555 5611
rect 4559 5607 4602 5611
rect 4522 5317 4602 5607
rect 4522 5313 4525 5317
rect 4529 5313 4535 5317
rect 4539 5313 4545 5317
rect 4549 5313 4555 5317
rect 4559 5313 4602 5317
rect 4522 5312 4602 5313
rect 4522 5308 4525 5312
rect 4529 5308 4535 5312
rect 4539 5308 4545 5312
rect 4549 5308 4555 5312
rect 4559 5308 4602 5312
rect 4522 5307 4602 5308
rect 4522 5303 4525 5307
rect 4529 5303 4535 5307
rect 4539 5303 4545 5307
rect 4549 5303 4555 5307
rect 4559 5303 4602 5307
rect 4522 5302 4602 5303
rect 4522 5298 4525 5302
rect 4529 5298 4535 5302
rect 4539 5298 4545 5302
rect 4549 5298 4555 5302
rect 4559 5298 4602 5302
rect 4522 5008 4602 5298
rect 4522 5004 4525 5008
rect 4529 5004 4535 5008
rect 4539 5004 4545 5008
rect 4549 5004 4555 5008
rect 4559 5004 4602 5008
rect 4522 5003 4602 5004
rect 4522 4999 4525 5003
rect 4529 4999 4535 5003
rect 4539 4999 4545 5003
rect 4549 4999 4555 5003
rect 4559 4999 4602 5003
rect 4522 4998 4602 4999
rect 4522 4994 4525 4998
rect 4529 4994 4535 4998
rect 4539 4994 4545 4998
rect 4549 4994 4555 4998
rect 4559 4994 4602 4998
rect 4522 4993 4602 4994
rect 4522 4989 4525 4993
rect 4529 4989 4535 4993
rect 4539 4989 4545 4993
rect 4549 4989 4555 4993
rect 4559 4989 4602 4993
rect 4522 4815 4602 4989
rect 4522 4811 4525 4815
rect 4529 4811 4535 4815
rect 4539 4811 4545 4815
rect 4549 4811 4555 4815
rect 4559 4811 4602 4815
rect 4522 4810 4602 4811
rect 4522 4806 4525 4810
rect 4529 4806 4535 4810
rect 4539 4806 4545 4810
rect 4549 4806 4555 4810
rect 4559 4806 4602 4810
rect 4522 4805 4602 4806
rect 4522 4801 4525 4805
rect 4529 4801 4535 4805
rect 4539 4801 4545 4805
rect 4549 4801 4555 4805
rect 4559 4801 4602 4805
rect 4522 4800 4602 4801
rect 4522 4796 4525 4800
rect 4529 4796 4535 4800
rect 4539 4796 4545 4800
rect 4549 4796 4555 4800
rect 4559 4796 4602 4800
rect 4522 4789 4602 4796
rect 4522 4785 4525 4789
rect 4529 4785 4535 4789
rect 4539 4785 4545 4789
rect 4549 4785 4555 4789
rect 4559 4785 4602 4789
rect 4522 4784 4602 4785
rect 4522 4780 4525 4784
rect 4529 4780 4535 4784
rect 4539 4780 4545 4784
rect 4549 4780 4555 4784
rect 4559 4780 4602 4784
rect 4522 4779 4602 4780
rect 4522 4775 4525 4779
rect 4529 4775 4535 4779
rect 4539 4775 4545 4779
rect 4549 4775 4555 4779
rect 4559 4775 4602 4779
rect 4522 4774 4602 4775
rect 4522 4770 4525 4774
rect 4529 4770 4535 4774
rect 4539 4770 4545 4774
rect 4549 4770 4555 4774
rect 4559 4770 4602 4774
rect 4522 4763 4602 4770
rect 4522 4759 4525 4763
rect 4529 4759 4535 4763
rect 4539 4759 4545 4763
rect 4549 4759 4555 4763
rect 4559 4759 4602 4763
rect 4522 4758 4602 4759
rect 4522 4754 4525 4758
rect 4529 4754 4535 4758
rect 4539 4754 4545 4758
rect 4549 4754 4555 4758
rect 4559 4754 4602 4758
rect 4522 4753 4602 4754
rect 4522 4749 4525 4753
rect 4529 4749 4535 4753
rect 4539 4749 4545 4753
rect 4549 4749 4555 4753
rect 4559 4749 4602 4753
rect 4522 4748 4602 4749
rect 4522 4744 4525 4748
rect 4529 4744 4535 4748
rect 4539 4744 4545 4748
rect 4549 4744 4555 4748
rect 4559 4744 4602 4748
rect 4522 4737 4602 4744
rect 4522 4733 4525 4737
rect 4529 4733 4535 4737
rect 4539 4733 4545 4737
rect 4549 4733 4555 4737
rect 4559 4733 4602 4737
rect 4522 4732 4602 4733
rect 4522 4728 4525 4732
rect 4529 4728 4535 4732
rect 4539 4728 4545 4732
rect 4549 4728 4555 4732
rect 4559 4728 4602 4732
rect 4522 4727 4602 4728
rect 4522 4723 4525 4727
rect 4529 4723 4535 4727
rect 4539 4723 4545 4727
rect 4549 4723 4555 4727
rect 4559 4723 4602 4727
rect 4522 4722 4602 4723
rect 4522 4718 4525 4722
rect 4529 4718 4535 4722
rect 4539 4718 4545 4722
rect 4549 4718 4555 4722
rect 4559 4718 4602 4722
rect 4522 4711 4602 4718
rect 4522 4707 4525 4711
rect 4529 4707 4535 4711
rect 4539 4707 4545 4711
rect 4549 4707 4555 4711
rect 4559 4707 4602 4711
rect 4522 4706 4602 4707
rect 4522 4702 4525 4706
rect 4529 4702 4535 4706
rect 4539 4702 4545 4706
rect 4549 4702 4555 4706
rect 4559 4702 4602 4706
rect 4522 4701 4602 4702
rect 4522 4697 4525 4701
rect 4529 4697 4535 4701
rect 4539 4697 4545 4701
rect 4549 4697 4555 4701
rect 4559 4697 4602 4701
rect 4522 4696 4602 4697
rect 4522 4692 4525 4696
rect 4529 4692 4535 4696
rect 4539 4692 4545 4696
rect 4549 4692 4555 4696
rect 4559 4692 4602 4696
rect 4522 4585 4602 4692
rect 570 4582 4602 4585
rect 570 4578 757 4582
rect 761 4578 762 4582
rect 766 4578 767 4582
rect 771 4578 772 4582
rect 776 4578 783 4582
rect 787 4578 788 4582
rect 792 4578 793 4582
rect 797 4578 798 4582
rect 802 4578 809 4582
rect 813 4578 814 4582
rect 818 4578 819 4582
rect 823 4578 824 4582
rect 828 4578 835 4582
rect 839 4578 840 4582
rect 844 4578 845 4582
rect 849 4578 850 4582
rect 854 4578 861 4582
rect 865 4578 866 4582
rect 870 4578 871 4582
rect 875 4578 876 4582
rect 880 4578 1053 4582
rect 1057 4578 1058 4582
rect 1062 4578 1063 4582
rect 1067 4578 1068 4582
rect 1072 4578 1362 4582
rect 1366 4578 1367 4582
rect 1371 4578 1372 4582
rect 1376 4578 1377 4582
rect 1381 4578 1671 4582
rect 1675 4578 1676 4582
rect 1680 4578 1681 4582
rect 1685 4578 1686 4582
rect 1690 4578 1980 4582
rect 1984 4578 1985 4582
rect 1989 4578 1990 4582
rect 1994 4578 1995 4582
rect 1999 4578 2289 4582
rect 2293 4578 2294 4582
rect 2298 4578 2299 4582
rect 2303 4578 2304 4582
rect 2308 4578 2598 4582
rect 2602 4578 2603 4582
rect 2607 4578 2608 4582
rect 2612 4578 2613 4582
rect 2617 4578 2907 4582
rect 2911 4578 2912 4582
rect 2916 4578 2917 4582
rect 2921 4578 2922 4582
rect 2926 4578 3216 4582
rect 3220 4578 3221 4582
rect 3225 4578 3226 4582
rect 3230 4578 3231 4582
rect 3235 4578 3525 4582
rect 3529 4578 3530 4582
rect 3534 4578 3535 4582
rect 3539 4578 3540 4582
rect 3544 4578 3834 4582
rect 3838 4578 3839 4582
rect 3843 4578 3844 4582
rect 3848 4578 3849 4582
rect 3853 4578 4235 4582
rect 4239 4578 4240 4582
rect 4244 4578 4245 4582
rect 4249 4578 4250 4582
rect 4254 4578 4264 4582
rect 4268 4578 4269 4582
rect 4273 4578 4274 4582
rect 4278 4578 4279 4582
rect 4283 4578 4293 4582
rect 4297 4578 4298 4582
rect 4302 4578 4303 4582
rect 4307 4578 4308 4582
rect 4312 4578 4322 4582
rect 4326 4578 4327 4582
rect 4331 4578 4332 4582
rect 4336 4578 4337 4582
rect 4341 4578 4351 4582
rect 4355 4578 4356 4582
rect 4360 4578 4361 4582
rect 4365 4578 4366 4582
rect 4370 4578 4602 4582
rect 570 4574 1337 4578
rect 1341 4574 1342 4578
rect 1346 4574 1646 4578
rect 1650 4574 1651 4578
rect 1655 4574 1955 4578
rect 1959 4574 1960 4578
rect 1964 4574 2264 4578
rect 2268 4574 2269 4578
rect 2273 4574 2573 4578
rect 2577 4574 2578 4578
rect 2582 4574 2882 4578
rect 2886 4574 2887 4578
rect 2891 4574 3000 4578
rect 570 4573 3000 4574
rect 3005 4574 3191 4578
rect 3195 4574 3196 4578
rect 3200 4574 3500 4578
rect 3504 4574 3505 4578
rect 3509 4574 3809 4578
rect 3813 4574 3814 4578
rect 3818 4574 4602 4578
rect 3005 4573 4602 4574
rect 570 4572 1337 4573
rect 570 4568 757 4572
rect 761 4568 762 4572
rect 766 4568 767 4572
rect 771 4568 772 4572
rect 776 4568 783 4572
rect 787 4568 788 4572
rect 792 4568 793 4572
rect 797 4568 798 4572
rect 802 4568 809 4572
rect 813 4568 814 4572
rect 818 4568 819 4572
rect 823 4568 824 4572
rect 828 4568 835 4572
rect 839 4568 840 4572
rect 844 4568 845 4572
rect 849 4568 850 4572
rect 854 4568 861 4572
rect 865 4568 866 4572
rect 870 4568 871 4572
rect 875 4568 876 4572
rect 880 4568 1053 4572
rect 1057 4568 1058 4572
rect 1062 4568 1063 4572
rect 1067 4568 1068 4572
rect 1072 4569 1337 4572
rect 1341 4569 1342 4573
rect 1346 4572 1511 4573
rect 1346 4569 1362 4572
rect 1072 4568 1362 4569
rect 1366 4568 1367 4572
rect 1371 4568 1372 4572
rect 1376 4568 1377 4572
rect 1381 4569 1511 4572
rect 1515 4569 1516 4573
rect 1520 4569 1646 4573
rect 1650 4569 1651 4573
rect 1655 4572 1955 4573
rect 1655 4569 1671 4572
rect 1381 4568 1671 4569
rect 1675 4568 1676 4572
rect 1680 4568 1681 4572
rect 1685 4568 1686 4572
rect 1690 4569 1955 4572
rect 1959 4569 1960 4573
rect 1964 4572 2264 4573
rect 1964 4569 1980 4572
rect 1690 4568 1980 4569
rect 1984 4568 1985 4572
rect 1989 4568 1990 4572
rect 1994 4568 1995 4572
rect 1999 4569 2264 4572
rect 2268 4569 2269 4573
rect 2273 4572 2573 4573
rect 2273 4569 2289 4572
rect 1999 4568 2289 4569
rect 2293 4568 2294 4572
rect 2298 4568 2299 4572
rect 2303 4568 2304 4572
rect 2308 4569 2573 4572
rect 2577 4569 2578 4573
rect 2582 4572 2882 4573
rect 2582 4569 2598 4572
rect 2308 4568 2598 4569
rect 2602 4568 2603 4572
rect 2607 4568 2608 4572
rect 2612 4568 2613 4572
rect 2617 4569 2882 4572
rect 2886 4569 2887 4573
rect 2891 4572 3191 4573
rect 2891 4569 2907 4572
rect 2617 4568 2907 4569
rect 2911 4568 2912 4572
rect 2916 4568 2917 4572
rect 2921 4568 2922 4572
rect 2926 4569 3191 4572
rect 3195 4569 3196 4573
rect 3200 4572 3500 4573
rect 3200 4569 3216 4572
rect 2926 4568 3216 4569
rect 3220 4568 3221 4572
rect 3225 4568 3226 4572
rect 3230 4568 3231 4572
rect 3235 4569 3500 4572
rect 3504 4569 3505 4573
rect 3509 4572 3809 4573
rect 3509 4569 3525 4572
rect 3235 4568 3525 4569
rect 3529 4568 3530 4572
rect 3534 4568 3535 4572
rect 3539 4568 3540 4572
rect 3544 4569 3809 4572
rect 3813 4569 3814 4573
rect 3818 4572 4602 4573
rect 3818 4569 3834 4572
rect 3544 4568 3834 4569
rect 3838 4568 3839 4572
rect 3843 4568 3844 4572
rect 3848 4568 3849 4572
rect 3853 4568 4235 4572
rect 4239 4568 4240 4572
rect 4244 4568 4245 4572
rect 4249 4568 4250 4572
rect 4254 4568 4264 4572
rect 4268 4568 4269 4572
rect 4273 4568 4274 4572
rect 4278 4568 4279 4572
rect 4283 4568 4293 4572
rect 4297 4568 4298 4572
rect 4302 4568 4303 4572
rect 4307 4568 4308 4572
rect 4312 4568 4322 4572
rect 4326 4568 4327 4572
rect 4331 4568 4332 4572
rect 4336 4568 4337 4572
rect 4341 4568 4351 4572
rect 4355 4568 4356 4572
rect 4360 4568 4361 4572
rect 4365 4568 4366 4572
rect 4370 4568 4602 4572
rect 570 4564 1337 4568
rect 1341 4564 1342 4568
rect 1346 4564 1511 4568
rect 1515 4564 1516 4568
rect 1520 4564 1646 4568
rect 1650 4564 1651 4568
rect 1655 4564 1955 4568
rect 1959 4564 1960 4568
rect 1964 4564 2264 4568
rect 2268 4564 2269 4568
rect 2273 4564 2573 4568
rect 2577 4564 2578 4568
rect 2582 4564 2882 4568
rect 2886 4564 2887 4568
rect 2891 4564 3191 4568
rect 3195 4564 3196 4568
rect 3200 4564 3500 4568
rect 3504 4564 3505 4568
rect 3509 4564 3809 4568
rect 3813 4564 3814 4568
rect 3818 4564 4602 4568
rect 570 4563 4602 4564
rect 570 4562 1337 4563
rect 570 4558 757 4562
rect 761 4558 762 4562
rect 766 4558 767 4562
rect 771 4558 772 4562
rect 776 4558 783 4562
rect 787 4558 788 4562
rect 792 4558 793 4562
rect 797 4558 798 4562
rect 802 4558 809 4562
rect 813 4558 814 4562
rect 818 4558 819 4562
rect 823 4558 824 4562
rect 828 4558 835 4562
rect 839 4558 840 4562
rect 844 4558 845 4562
rect 849 4558 850 4562
rect 854 4558 861 4562
rect 865 4558 866 4562
rect 870 4558 871 4562
rect 875 4558 876 4562
rect 880 4558 1053 4562
rect 1057 4558 1058 4562
rect 1062 4558 1063 4562
rect 1067 4558 1068 4562
rect 1072 4559 1337 4562
rect 1341 4559 1342 4563
rect 1346 4562 1511 4563
rect 1346 4559 1362 4562
rect 1072 4558 1362 4559
rect 1366 4558 1367 4562
rect 1371 4558 1372 4562
rect 1376 4558 1377 4562
rect 1381 4559 1511 4562
rect 1515 4559 1516 4563
rect 1520 4559 1646 4563
rect 1650 4559 1651 4563
rect 1655 4562 1955 4563
rect 1655 4559 1671 4562
rect 1381 4558 1671 4559
rect 1675 4558 1676 4562
rect 1680 4558 1681 4562
rect 1685 4558 1686 4562
rect 1690 4559 1955 4562
rect 1959 4559 1960 4563
rect 1964 4562 2264 4563
rect 1964 4559 1980 4562
rect 1690 4558 1980 4559
rect 1984 4558 1985 4562
rect 1989 4558 1990 4562
rect 1994 4558 1995 4562
rect 1999 4559 2264 4562
rect 2268 4559 2269 4563
rect 2273 4562 2573 4563
rect 2273 4559 2289 4562
rect 1999 4558 2289 4559
rect 2293 4558 2294 4562
rect 2298 4558 2299 4562
rect 2303 4558 2304 4562
rect 2308 4559 2573 4562
rect 2577 4559 2578 4563
rect 2582 4562 2882 4563
rect 2582 4559 2598 4562
rect 2308 4558 2598 4559
rect 2602 4558 2603 4562
rect 2607 4558 2608 4562
rect 2612 4558 2613 4562
rect 2617 4559 2882 4562
rect 2886 4559 2887 4563
rect 2891 4562 3191 4563
rect 2891 4559 2907 4562
rect 2617 4558 2907 4559
rect 2911 4558 2912 4562
rect 2916 4558 2917 4562
rect 2921 4558 2922 4562
rect 2926 4559 3191 4562
rect 3195 4559 3196 4563
rect 3200 4562 3500 4563
rect 3200 4559 3216 4562
rect 2926 4558 3216 4559
rect 3220 4558 3221 4562
rect 3225 4558 3226 4562
rect 3230 4558 3231 4562
rect 3235 4559 3500 4562
rect 3504 4559 3505 4563
rect 3509 4562 3809 4563
rect 3509 4559 3525 4562
rect 3235 4558 3525 4559
rect 3529 4558 3530 4562
rect 3534 4558 3535 4562
rect 3539 4558 3540 4562
rect 3544 4559 3809 4562
rect 3813 4559 3814 4563
rect 3818 4562 4602 4563
rect 3818 4559 3834 4562
rect 3544 4558 3834 4559
rect 3838 4558 3839 4562
rect 3843 4558 3844 4562
rect 3848 4558 3849 4562
rect 3853 4558 4235 4562
rect 4239 4558 4240 4562
rect 4244 4558 4245 4562
rect 4249 4558 4250 4562
rect 4254 4558 4264 4562
rect 4268 4558 4269 4562
rect 4273 4558 4274 4562
rect 4278 4558 4279 4562
rect 4283 4558 4293 4562
rect 4297 4558 4298 4562
rect 4302 4558 4303 4562
rect 4307 4558 4308 4562
rect 4312 4558 4322 4562
rect 4326 4558 4327 4562
rect 4331 4558 4332 4562
rect 4336 4558 4337 4562
rect 4341 4558 4351 4562
rect 4355 4558 4356 4562
rect 4360 4558 4361 4562
rect 4365 4558 4366 4562
rect 4370 4558 4602 4562
rect 570 4554 1337 4558
rect 1341 4554 1342 4558
rect 1346 4554 1511 4558
rect 1515 4554 1516 4558
rect 1520 4554 1646 4558
rect 1650 4554 1651 4558
rect 1655 4554 1955 4558
rect 1959 4554 1960 4558
rect 1964 4554 2264 4558
rect 2268 4554 2269 4558
rect 2273 4554 2573 4558
rect 2577 4554 2578 4558
rect 2582 4554 2882 4558
rect 2886 4554 2887 4558
rect 2891 4554 3191 4558
rect 3195 4554 3196 4558
rect 3200 4554 3500 4558
rect 3504 4554 3505 4558
rect 3509 4554 3809 4558
rect 3813 4554 3814 4558
rect 3818 4554 4602 4558
rect 570 4552 1089 4554
rect 570 4548 757 4552
rect 761 4548 762 4552
rect 766 4548 767 4552
rect 771 4548 772 4552
rect 776 4548 783 4552
rect 787 4548 788 4552
rect 792 4548 793 4552
rect 797 4548 798 4552
rect 802 4548 809 4552
rect 813 4548 814 4552
rect 818 4548 819 4552
rect 823 4548 824 4552
rect 828 4548 835 4552
rect 839 4548 840 4552
rect 844 4548 845 4552
rect 849 4548 850 4552
rect 854 4548 861 4552
rect 865 4548 866 4552
rect 870 4548 871 4552
rect 875 4548 876 4552
rect 880 4548 1053 4552
rect 1057 4548 1058 4552
rect 1062 4548 1063 4552
rect 1067 4548 1068 4552
rect 1072 4550 1089 4552
rect 1093 4550 1094 4554
rect 1098 4550 1099 4554
rect 1103 4550 1104 4554
rect 1108 4550 1109 4554
rect 1113 4550 1114 4554
rect 1118 4550 1119 4554
rect 1123 4550 1124 4554
rect 1128 4550 1129 4554
rect 1133 4550 1134 4554
rect 1138 4550 1139 4554
rect 1143 4550 1144 4554
rect 1148 4550 1149 4554
rect 1153 4553 1398 4554
rect 1153 4550 1337 4553
rect 1072 4549 1337 4550
rect 1341 4549 1342 4553
rect 1346 4552 1398 4553
rect 1346 4549 1362 4552
rect 1072 4548 1089 4549
rect 570 4545 1089 4548
rect 1093 4545 1094 4549
rect 1098 4545 1099 4549
rect 1103 4545 1104 4549
rect 1108 4545 1109 4549
rect 1113 4545 1114 4549
rect 1118 4545 1119 4549
rect 1123 4545 1124 4549
rect 1128 4545 1129 4549
rect 1133 4545 1134 4549
rect 1138 4545 1139 4549
rect 1143 4545 1144 4549
rect 1148 4545 1149 4549
rect 1153 4548 1362 4549
rect 1366 4548 1367 4552
rect 1371 4548 1372 4552
rect 1376 4548 1377 4552
rect 1381 4550 1398 4552
rect 1402 4550 1403 4554
rect 1407 4550 1408 4554
rect 1412 4550 1413 4554
rect 1417 4550 1418 4554
rect 1422 4550 1423 4554
rect 1427 4550 1428 4554
rect 1432 4550 1433 4554
rect 1437 4550 1438 4554
rect 1442 4550 1443 4554
rect 1447 4550 1448 4554
rect 1452 4550 1453 4554
rect 1457 4550 1458 4554
rect 1462 4553 1707 4554
rect 1462 4550 1511 4553
rect 1381 4549 1511 4550
rect 1515 4549 1516 4553
rect 1520 4549 1646 4553
rect 1650 4549 1651 4553
rect 1655 4552 1707 4553
rect 1655 4549 1671 4552
rect 1381 4548 1398 4549
rect 1153 4545 1337 4548
rect 570 4544 1337 4545
rect 1341 4544 1342 4548
rect 1346 4545 1398 4548
rect 1402 4545 1403 4549
rect 1407 4545 1408 4549
rect 1412 4545 1413 4549
rect 1417 4545 1418 4549
rect 1422 4545 1423 4549
rect 1427 4545 1428 4549
rect 1432 4545 1433 4549
rect 1437 4545 1438 4549
rect 1442 4545 1443 4549
rect 1447 4545 1448 4549
rect 1452 4545 1453 4549
rect 1457 4545 1458 4549
rect 1462 4548 1671 4549
rect 1675 4548 1676 4552
rect 1680 4548 1681 4552
rect 1685 4548 1686 4552
rect 1690 4550 1707 4552
rect 1711 4550 1712 4554
rect 1716 4550 1717 4554
rect 1721 4550 1722 4554
rect 1726 4550 1727 4554
rect 1731 4550 1732 4554
rect 1736 4550 1737 4554
rect 1741 4550 1742 4554
rect 1746 4550 1747 4554
rect 1751 4550 1752 4554
rect 1756 4550 1757 4554
rect 1761 4550 1762 4554
rect 1766 4550 1767 4554
rect 1771 4553 2016 4554
rect 1771 4550 1955 4553
rect 1690 4549 1955 4550
rect 1959 4549 1960 4553
rect 1964 4552 2016 4553
rect 1964 4549 1980 4552
rect 1690 4548 1707 4549
rect 1462 4545 1511 4548
rect 1346 4544 1511 4545
rect 1515 4544 1516 4548
rect 1520 4544 1646 4548
rect 1650 4544 1651 4548
rect 1655 4545 1707 4548
rect 1711 4545 1712 4549
rect 1716 4545 1717 4549
rect 1721 4545 1722 4549
rect 1726 4545 1727 4549
rect 1731 4545 1732 4549
rect 1736 4545 1737 4549
rect 1741 4545 1742 4549
rect 1746 4545 1747 4549
rect 1751 4545 1752 4549
rect 1756 4545 1757 4549
rect 1761 4545 1762 4549
rect 1766 4545 1767 4549
rect 1771 4548 1980 4549
rect 1984 4548 1985 4552
rect 1989 4548 1990 4552
rect 1994 4548 1995 4552
rect 1999 4550 2016 4552
rect 2020 4550 2021 4554
rect 2025 4550 2026 4554
rect 2030 4550 2031 4554
rect 2035 4550 2036 4554
rect 2040 4550 2041 4554
rect 2045 4550 2046 4554
rect 2050 4550 2051 4554
rect 2055 4550 2056 4554
rect 2060 4550 2061 4554
rect 2065 4550 2066 4554
rect 2070 4550 2071 4554
rect 2075 4550 2076 4554
rect 2080 4553 2325 4554
rect 2080 4550 2264 4553
rect 1999 4549 2264 4550
rect 2268 4549 2269 4553
rect 2273 4552 2325 4553
rect 2273 4549 2289 4552
rect 1999 4548 2016 4549
rect 1771 4545 1955 4548
rect 1655 4544 1955 4545
rect 1959 4544 1960 4548
rect 1964 4545 2016 4548
rect 2020 4545 2021 4549
rect 2025 4545 2026 4549
rect 2030 4545 2031 4549
rect 2035 4545 2036 4549
rect 2040 4545 2041 4549
rect 2045 4545 2046 4549
rect 2050 4545 2051 4549
rect 2055 4545 2056 4549
rect 2060 4545 2061 4549
rect 2065 4545 2066 4549
rect 2070 4545 2071 4549
rect 2075 4545 2076 4549
rect 2080 4548 2289 4549
rect 2293 4548 2294 4552
rect 2298 4548 2299 4552
rect 2303 4548 2304 4552
rect 2308 4550 2325 4552
rect 2329 4550 2330 4554
rect 2334 4550 2335 4554
rect 2339 4550 2340 4554
rect 2344 4550 2345 4554
rect 2349 4550 2350 4554
rect 2354 4550 2355 4554
rect 2359 4550 2360 4554
rect 2364 4550 2365 4554
rect 2369 4550 2370 4554
rect 2374 4550 2375 4554
rect 2379 4550 2380 4554
rect 2384 4550 2385 4554
rect 2389 4553 2634 4554
rect 2389 4550 2573 4553
rect 2308 4549 2573 4550
rect 2577 4549 2578 4553
rect 2582 4552 2634 4553
rect 2582 4549 2598 4552
rect 2308 4548 2325 4549
rect 2080 4545 2264 4548
rect 1964 4544 2264 4545
rect 2268 4544 2269 4548
rect 2273 4545 2325 4548
rect 2329 4545 2330 4549
rect 2334 4545 2335 4549
rect 2339 4545 2340 4549
rect 2344 4545 2345 4549
rect 2349 4545 2350 4549
rect 2354 4545 2355 4549
rect 2359 4545 2360 4549
rect 2364 4545 2365 4549
rect 2369 4545 2370 4549
rect 2374 4545 2375 4549
rect 2379 4545 2380 4549
rect 2384 4545 2385 4549
rect 2389 4548 2598 4549
rect 2602 4548 2603 4552
rect 2607 4548 2608 4552
rect 2612 4548 2613 4552
rect 2617 4550 2634 4552
rect 2638 4550 2639 4554
rect 2643 4550 2644 4554
rect 2648 4550 2649 4554
rect 2653 4550 2654 4554
rect 2658 4550 2659 4554
rect 2663 4550 2664 4554
rect 2668 4550 2669 4554
rect 2673 4550 2674 4554
rect 2678 4550 2679 4554
rect 2683 4550 2684 4554
rect 2688 4550 2689 4554
rect 2693 4550 2694 4554
rect 2698 4553 2943 4554
rect 2698 4550 2882 4553
rect 2617 4549 2882 4550
rect 2886 4549 2887 4553
rect 2891 4552 2943 4553
rect 2891 4549 2907 4552
rect 2617 4548 2634 4549
rect 2389 4545 2573 4548
rect 2273 4544 2573 4545
rect 2577 4544 2578 4548
rect 2582 4545 2634 4548
rect 2638 4545 2639 4549
rect 2643 4545 2644 4549
rect 2648 4545 2649 4549
rect 2653 4545 2654 4549
rect 2658 4545 2659 4549
rect 2663 4545 2664 4549
rect 2668 4545 2669 4549
rect 2673 4545 2674 4549
rect 2678 4545 2679 4549
rect 2683 4545 2684 4549
rect 2688 4545 2689 4549
rect 2693 4545 2694 4549
rect 2698 4548 2907 4549
rect 2911 4548 2912 4552
rect 2916 4548 2917 4552
rect 2921 4548 2922 4552
rect 2926 4550 2943 4552
rect 2947 4550 2948 4554
rect 2952 4550 2953 4554
rect 2957 4550 2958 4554
rect 2962 4550 2963 4554
rect 2967 4550 2968 4554
rect 2972 4550 2973 4554
rect 2977 4550 2978 4554
rect 2982 4550 2983 4554
rect 2987 4550 2988 4554
rect 2992 4550 2993 4554
rect 2997 4550 2998 4554
rect 3002 4550 3003 4554
rect 3007 4553 3252 4554
rect 3007 4550 3191 4553
rect 2926 4549 3191 4550
rect 3195 4549 3196 4553
rect 3200 4552 3252 4553
rect 3200 4549 3216 4552
rect 2926 4548 2943 4549
rect 2698 4545 2882 4548
rect 2582 4544 2882 4545
rect 2886 4544 2887 4548
rect 2891 4545 2943 4548
rect 2947 4545 2948 4549
rect 2952 4545 2953 4549
rect 2957 4545 2958 4549
rect 2962 4545 2963 4549
rect 2967 4545 2968 4549
rect 2972 4545 2973 4549
rect 2977 4545 2978 4549
rect 2982 4545 2983 4549
rect 2987 4545 2988 4549
rect 2992 4545 2993 4549
rect 2997 4545 2998 4549
rect 3002 4545 3003 4549
rect 3007 4548 3216 4549
rect 3220 4548 3221 4552
rect 3225 4548 3226 4552
rect 3230 4548 3231 4552
rect 3235 4550 3252 4552
rect 3256 4550 3257 4554
rect 3261 4550 3262 4554
rect 3266 4550 3267 4554
rect 3271 4550 3272 4554
rect 3276 4550 3277 4554
rect 3281 4550 3282 4554
rect 3286 4550 3287 4554
rect 3291 4550 3292 4554
rect 3296 4550 3297 4554
rect 3301 4550 3302 4554
rect 3306 4550 3307 4554
rect 3311 4550 3312 4554
rect 3316 4553 3561 4554
rect 3316 4550 3500 4553
rect 3235 4549 3500 4550
rect 3504 4549 3505 4553
rect 3509 4552 3561 4553
rect 3509 4549 3525 4552
rect 3235 4548 3252 4549
rect 3007 4545 3191 4548
rect 2891 4544 3191 4545
rect 3195 4544 3196 4548
rect 3200 4545 3252 4548
rect 3256 4545 3257 4549
rect 3261 4545 3262 4549
rect 3266 4545 3267 4549
rect 3271 4545 3272 4549
rect 3276 4545 3277 4549
rect 3281 4545 3282 4549
rect 3286 4545 3287 4549
rect 3291 4545 3292 4549
rect 3296 4545 3297 4549
rect 3301 4545 3302 4549
rect 3306 4545 3307 4549
rect 3311 4545 3312 4549
rect 3316 4548 3525 4549
rect 3529 4548 3530 4552
rect 3534 4548 3535 4552
rect 3539 4548 3540 4552
rect 3544 4550 3561 4552
rect 3565 4550 3566 4554
rect 3570 4550 3571 4554
rect 3575 4550 3576 4554
rect 3580 4550 3581 4554
rect 3585 4550 3586 4554
rect 3590 4550 3591 4554
rect 3595 4550 3596 4554
rect 3600 4550 3601 4554
rect 3605 4550 3606 4554
rect 3610 4550 3611 4554
rect 3615 4550 3616 4554
rect 3620 4550 3621 4554
rect 3625 4553 4602 4554
rect 3625 4550 3809 4553
rect 3544 4549 3809 4550
rect 3813 4549 3814 4553
rect 3818 4552 4602 4553
rect 3818 4549 3834 4552
rect 3544 4548 3561 4549
rect 3316 4545 3500 4548
rect 3200 4544 3500 4545
rect 3504 4544 3505 4548
rect 3509 4545 3561 4548
rect 3565 4545 3566 4549
rect 3570 4545 3571 4549
rect 3575 4545 3576 4549
rect 3580 4545 3581 4549
rect 3585 4545 3586 4549
rect 3590 4545 3591 4549
rect 3595 4545 3596 4549
rect 3600 4545 3601 4549
rect 3605 4545 3606 4549
rect 3610 4545 3611 4549
rect 3615 4545 3616 4549
rect 3620 4545 3621 4549
rect 3625 4548 3834 4549
rect 3838 4548 3839 4552
rect 3843 4548 3844 4552
rect 3848 4548 3849 4552
rect 3853 4548 4235 4552
rect 4239 4548 4240 4552
rect 4244 4548 4245 4552
rect 4249 4548 4250 4552
rect 4254 4548 4264 4552
rect 4268 4548 4269 4552
rect 4273 4548 4274 4552
rect 4278 4548 4279 4552
rect 4283 4548 4293 4552
rect 4297 4548 4298 4552
rect 4302 4548 4303 4552
rect 4307 4548 4308 4552
rect 4312 4548 4322 4552
rect 4326 4548 4327 4552
rect 4331 4548 4332 4552
rect 4336 4548 4337 4552
rect 4341 4548 4351 4552
rect 4355 4548 4356 4552
rect 4360 4548 4361 4552
rect 4365 4548 4366 4552
rect 4370 4548 4602 4552
rect 3625 4545 3809 4548
rect 3509 4544 3809 4545
rect 3813 4544 3814 4548
rect 3818 4544 4602 4548
rect 570 4543 4602 4544
rect 570 4539 1337 4543
rect 1341 4539 1342 4543
rect 1346 4539 1511 4543
rect 1515 4539 1516 4543
rect 1520 4539 1646 4543
rect 1650 4539 1651 4543
rect 1655 4539 1955 4543
rect 1959 4539 1960 4543
rect 1964 4539 2264 4543
rect 2268 4539 2269 4543
rect 2273 4539 2573 4543
rect 2577 4539 2578 4543
rect 2582 4539 2882 4543
rect 2886 4539 2887 4543
rect 2891 4539 3191 4543
rect 3195 4539 3196 4543
rect 3200 4539 3500 4543
rect 3504 4539 3505 4543
rect 3509 4539 3809 4543
rect 3813 4539 3814 4543
rect 3818 4539 4602 4543
rect 570 4538 4602 4539
rect 570 4534 1337 4538
rect 1341 4534 1342 4538
rect 1346 4534 1511 4538
rect 1515 4534 1516 4538
rect 1520 4534 1646 4538
rect 1650 4534 1651 4538
rect 1655 4534 1955 4538
rect 1959 4534 1960 4538
rect 1964 4534 2264 4538
rect 2268 4534 2269 4538
rect 2273 4534 2573 4538
rect 2577 4534 2578 4538
rect 2582 4534 2882 4538
rect 2886 4534 2887 4538
rect 2891 4534 3191 4538
rect 3195 4534 3196 4538
rect 3200 4534 3500 4538
rect 3504 4534 3505 4538
rect 3509 4534 3809 4538
rect 3813 4534 3814 4538
rect 3818 4534 4602 4538
rect 570 4533 4602 4534
rect 570 4529 1337 4533
rect 1341 4529 1342 4533
rect 1346 4529 1511 4533
rect 1515 4529 1516 4533
rect 1520 4529 1646 4533
rect 1650 4529 1651 4533
rect 1655 4529 1955 4533
rect 1959 4529 1960 4533
rect 1964 4529 2264 4533
rect 2268 4529 2269 4533
rect 2273 4529 2573 4533
rect 2577 4529 2578 4533
rect 2582 4529 2882 4533
rect 2886 4529 2887 4533
rect 2891 4529 3191 4533
rect 3195 4529 3196 4533
rect 3200 4529 3500 4533
rect 3504 4529 3505 4533
rect 3509 4529 3809 4533
rect 3813 4529 3814 4533
rect 3818 4529 4602 4533
rect 570 4528 4602 4529
rect 570 4524 1337 4528
rect 1341 4524 1342 4528
rect 1346 4524 1511 4528
rect 1515 4524 1516 4528
rect 1520 4524 1646 4528
rect 1650 4524 1651 4528
rect 1655 4524 1955 4528
rect 1959 4524 1960 4528
rect 1964 4524 2264 4528
rect 2268 4524 2269 4528
rect 2273 4524 2573 4528
rect 2577 4524 2578 4528
rect 2582 4524 2882 4528
rect 2886 4524 2887 4528
rect 2891 4524 3191 4528
rect 3195 4524 3196 4528
rect 3200 4524 3500 4528
rect 3504 4524 3505 4528
rect 3509 4524 3809 4528
rect 3813 4524 3814 4528
rect 3818 4524 4602 4528
rect 570 4523 4602 4524
rect 570 4519 1337 4523
rect 1341 4519 1342 4523
rect 1346 4519 1511 4523
rect 1515 4519 1516 4523
rect 1520 4519 1646 4523
rect 1650 4519 1651 4523
rect 1655 4519 1955 4523
rect 1959 4519 1960 4523
rect 1964 4519 2264 4523
rect 2268 4519 2269 4523
rect 2273 4519 2573 4523
rect 2577 4519 2578 4523
rect 2582 4519 2882 4523
rect 2886 4519 2887 4523
rect 2891 4519 3191 4523
rect 3195 4519 3196 4523
rect 3200 4519 3500 4523
rect 3504 4519 3505 4523
rect 3509 4519 3809 4523
rect 3813 4519 3814 4523
rect 3818 4519 4602 4523
rect 570 4518 4602 4519
rect 570 4514 1337 4518
rect 1341 4514 1342 4518
rect 1346 4514 1646 4518
rect 1650 4514 1651 4518
rect 1655 4514 1955 4518
rect 1959 4514 1960 4518
rect 1964 4514 2264 4518
rect 2268 4514 2269 4518
rect 2273 4514 2573 4518
rect 2577 4514 2578 4518
rect 2582 4514 2882 4518
rect 2886 4514 2887 4518
rect 2891 4514 3191 4518
rect 3195 4514 3196 4518
rect 3200 4514 3500 4518
rect 3504 4514 3505 4518
rect 3509 4514 3809 4518
rect 3813 4514 3814 4518
rect 3818 4514 4602 4518
rect 570 4505 4602 4514
<< pad >>
rect 1063 10036 1317 10290
rect 1372 10036 1626 10290
rect 1681 10036 1935 10290
rect 1990 10036 2244 10290
rect 2299 10036 2553 10290
rect 2608 10036 2862 10290
rect 2917 10036 3171 10290
rect 3226 10036 3480 10290
rect 3535 10036 3789 10290
rect 3844 10036 4098 10290
rect 89 9050 343 9304
rect 89 8741 343 8995
rect 89 8432 343 8686
rect 89 8123 343 8377
rect 89 7814 343 8068
rect 89 7505 343 7759
rect 89 7196 343 7450
rect 89 6852 343 7106
rect 89 6542 343 6796
rect 89 6233 343 6487
rect 89 5925 343 6179
rect 89 5616 343 5870
rect 89 5307 343 5561
rect 89 4998 343 5252
rect 4829 9062 5083 9316
rect 4829 8753 5083 9007
rect 4829 8444 5083 8698
rect 4829 8135 5083 8389
rect 4829 7827 5083 8081
rect 4829 7518 5083 7772
rect 4829 7236 5083 7490
rect 4829 6864 5083 7118
rect 4829 6555 5083 6809
rect 4829 6246 5083 6500
rect 4829 5937 5083 6191
rect 4829 5628 5083 5882
rect 4829 5319 5083 5573
rect 4829 5010 5083 5264
rect 1074 4024 1328 4278
rect 1383 4024 1637 4278
rect 1692 4024 1946 4278
rect 2001 4024 2255 4278
rect 2310 4024 2564 4278
rect 2619 4024 2873 4278
rect 2928 4024 3182 4278
rect 3237 4024 3491 4278
rect 3546 4024 3800 4278
rect 3855 4024 4109 4278
<< labels >>
rlabel pad 3886 10068 4035 10201 1 rst_b
rlabel metal1 3645 9817 3676 9851 1 Vdd!
rlabel metal1 3341 9819 3372 9853 1 GND!
rlabel pad 3037 10120 3068 10154 1 mode
rlabel pad 2739 10147 2770 10181 1 clk
rlabel pad 2404 10136 2435 10170 1 data
rlabel pad 2100 10131 2131 10165 1 program
rlabel pad 4906 7918 4937 7952 1 out
rlabel pad 1189 4108 1290 4244 1 rst_b1
rlabel pad 2386 4086 2487 4222 1 clk
rlabel pad 2070 4086 2206 4244 1 mode
rlabel pad 2692 4074 2828 4232 1 data1
rlabel pad 170 6251 306 6409 1 out1
rlabel pad 4846 7292 5003 7471 1 s_or_p
<< end >>
