magic
tech scmos
timestamp 1608330800
<< nwell >>
rect 1060 10033 1320 10293
rect 1369 10033 1629 10293
rect 1678 10033 1938 10293
rect 1987 10033 2247 10293
rect 2296 10033 2556 10293
rect 2605 10033 2865 10293
rect 2914 10033 3174 10293
rect 3223 10033 3483 10293
rect 3532 10033 3792 10293
rect 3841 10033 4101 10293
rect 86 9047 346 9307
rect 4826 9059 5086 9319
rect 86 8738 346 8998
rect 4826 8750 5086 9010
rect 86 8429 346 8689
rect 4826 8441 5086 8701
rect 86 8120 346 8380
rect 4826 8132 5086 8392
rect 86 7811 346 8071
rect 4826 7824 5086 8084
rect 86 7502 346 7762
rect 4826 7515 5086 7775
rect 86 7193 346 7453
rect 4826 7205 5086 7465
rect 86 6884 346 7144
rect 4826 6896 5086 7156
rect 86 6575 346 6835
rect 4826 6587 5086 6847
rect 86 6266 346 6526
rect 4826 6278 5086 6538
rect 1072 5293 1332 5553
rect 1381 5293 1641 5553
rect 1690 5293 1950 5553
rect 1999 5293 2259 5553
rect 2308 5293 2568 5553
rect 2617 5293 2877 5553
rect 2926 5293 3186 5553
rect 3235 5293 3495 5553
rect 3544 5293 3804 5553
rect 3853 5293 4113 5553
<< ntransistor >>
rect 1829 9824 1869 9826
rect 2138 9824 2178 9826
rect 2447 9824 2487 9826
rect 2756 9824 2796 9826
rect 3065 9824 3105 9826
rect 3992 9824 4032 9826
rect 1829 9816 1869 9818
rect 2138 9816 2178 9818
rect 2447 9816 2487 9818
rect 2756 9816 2796 9818
rect 3065 9816 3105 9818
rect 3992 9816 4032 9818
rect 1829 9808 1869 9810
rect 1829 9800 1869 9802
rect 1829 9792 1869 9794
rect 1829 9784 1869 9786
rect 2138 9808 2178 9810
rect 2138 9800 2178 9802
rect 2138 9792 2178 9794
rect 2138 9784 2178 9786
rect 2447 9808 2487 9810
rect 2447 9800 2487 9802
rect 2447 9792 2487 9794
rect 2447 9784 2487 9786
rect 2756 9808 2796 9810
rect 2756 9800 2796 9802
rect 2756 9792 2796 9794
rect 2756 9784 2796 9786
rect 3065 9808 3105 9810
rect 3065 9800 3105 9802
rect 3065 9792 3105 9794
rect 3065 9784 3105 9786
rect 3992 9808 4032 9810
rect 3992 9800 4032 9802
rect 3992 9792 4032 9794
rect 3992 9784 4032 9786
rect 2856 9299 2858 9303
rect 2861 9299 2863 9303
rect 2877 9299 2879 9303
rect 2893 9299 2895 9303
rect 2898 9299 2900 9303
rect 2919 9299 2921 9303
rect 2935 9299 2937 9303
rect 2951 9299 2953 9303
rect 2956 9299 2958 9303
rect 2972 9299 2974 9303
rect 2988 9299 2990 9303
rect 2993 9299 2995 9303
rect 3009 9299 3011 9303
rect 3025 9299 3027 9303
rect 3030 9299 3032 9303
rect 3051 9299 3053 9303
rect 3067 9299 3069 9303
rect 3083 9299 3085 9303
rect 3088 9299 3090 9303
rect 3104 9299 3106 9303
rect 3120 9299 3122 9303
rect 3125 9299 3127 9303
rect 3141 9299 3143 9303
rect 3157 9299 3159 9303
rect 3162 9299 3164 9303
rect 3183 9299 3185 9303
rect 3199 9299 3201 9303
rect 3215 9299 3217 9303
rect 3220 9299 3222 9303
rect 3236 9299 3238 9303
rect 3252 9299 3254 9303
rect 3257 9299 3259 9303
rect 3273 9299 3275 9303
rect 3289 9299 3291 9303
rect 3294 9299 3296 9303
rect 3315 9299 3317 9303
rect 3331 9299 3333 9303
rect 3347 9299 3349 9303
rect 3352 9299 3354 9303
rect 3368 9299 3370 9303
rect 3801 9299 3803 9303
rect 3806 9299 3808 9303
rect 3822 9299 3824 9303
rect 3838 9299 3840 9303
rect 3843 9299 3845 9303
rect 3864 9299 3866 9303
rect 3880 9299 3882 9303
rect 3896 9299 3898 9303
rect 3901 9299 3903 9303
rect 3917 9299 3919 9303
rect 3933 9299 3935 9303
rect 3938 9299 3940 9303
rect 3954 9299 3956 9303
rect 3970 9299 3972 9303
rect 3975 9299 3977 9303
rect 3996 9299 3998 9303
rect 4012 9299 4014 9303
rect 4028 9299 4030 9303
rect 4033 9299 4035 9303
rect 4049 9299 4051 9303
rect 4065 9299 4067 9303
rect 4070 9299 4072 9303
rect 4086 9299 4088 9303
rect 4102 9299 4104 9303
rect 4107 9299 4109 9303
rect 4128 9299 4130 9303
rect 4144 9299 4146 9303
rect 4160 9299 4162 9303
rect 4165 9299 4167 9303
rect 4181 9299 4183 9303
rect 4197 9299 4199 9303
rect 4202 9299 4204 9303
rect 4218 9299 4220 9303
rect 4234 9299 4236 9303
rect 4239 9299 4241 9303
rect 4260 9299 4262 9303
rect 4276 9299 4278 9303
rect 4292 9299 4294 9303
rect 4297 9299 4299 9303
rect 4313 9299 4315 9303
rect 2504 9266 2506 9270
rect 2509 9266 2511 9270
rect 2525 9266 2527 9270
rect 2541 9266 2543 9270
rect 2546 9266 2548 9270
rect 2567 9266 2569 9270
rect 2583 9266 2585 9270
rect 2599 9266 2601 9270
rect 2604 9266 2606 9270
rect 2620 9266 2622 9270
rect 3449 9266 3451 9270
rect 3454 9266 3456 9270
rect 3470 9266 3472 9270
rect 3486 9266 3488 9270
rect 3491 9266 3493 9270
rect 3512 9266 3514 9270
rect 3528 9266 3530 9270
rect 3544 9266 3546 9270
rect 3549 9266 3551 9270
rect 3565 9266 3567 9270
rect 2628 9229 2630 9233
rect 3035 9233 3037 9237
rect 3061 9229 3063 9233
rect 3066 9229 3068 9233
rect 3116 9233 3118 9237
rect 3142 9229 3144 9233
rect 3147 9229 3149 9233
rect 3089 9225 3091 9229
rect 2511 9220 2513 9224
rect 2861 9220 2863 9224
rect 2877 9220 2879 9224
rect 2893 9220 2895 9224
rect 2916 9220 2918 9224
rect 2921 9220 2923 9224
rect 2947 9220 2949 9224
rect 2968 9220 2970 9224
rect 2988 9220 2990 9224
rect 2993 9220 2995 9224
rect 3011 9220 3013 9224
rect 3170 9225 3172 9229
rect 3573 9229 3575 9233
rect 3980 9233 3982 9237
rect 4006 9229 4008 9233
rect 4011 9229 4013 9233
rect 4061 9233 4063 9237
rect 4087 9229 4089 9233
rect 4092 9229 4094 9233
rect 4034 9225 4036 9229
rect 3456 9220 3458 9224
rect 3806 9220 3808 9224
rect 3822 9220 3824 9224
rect 3838 9220 3840 9224
rect 3861 9220 3863 9224
rect 3866 9220 3868 9224
rect 3892 9220 3894 9224
rect 3913 9220 3915 9224
rect 3933 9220 3935 9224
rect 3938 9220 3940 9224
rect 3956 9220 3958 9224
rect 4115 9225 4117 9229
rect 2861 9174 2863 9178
rect 2877 9174 2879 9178
rect 2893 9174 2895 9178
rect 2916 9174 2918 9178
rect 2921 9174 2923 9178
rect 2947 9174 2949 9178
rect 2968 9174 2970 9178
rect 2988 9174 2990 9178
rect 2993 9174 2995 9178
rect 3011 9174 3013 9178
rect 2495 9164 2497 9168
rect 2511 9164 2513 9168
rect 2516 9164 2518 9168
rect 2532 9164 2534 9168
rect 2548 9164 2550 9168
rect 2569 9164 2571 9168
rect 2574 9164 2576 9168
rect 2590 9164 2592 9168
rect 2606 9164 2608 9168
rect 2611 9164 2613 9168
rect 3061 9173 3063 9177
rect 3066 9173 3068 9177
rect 3142 9173 3144 9177
rect 3147 9173 3149 9177
rect 3806 9174 3808 9178
rect 3822 9174 3824 9178
rect 3838 9174 3840 9178
rect 3861 9174 3863 9178
rect 3866 9174 3868 9178
rect 3892 9174 3894 9178
rect 3913 9174 3915 9178
rect 3933 9174 3935 9178
rect 3938 9174 3940 9178
rect 3956 9174 3958 9178
rect 3440 9164 3442 9168
rect 3456 9164 3458 9168
rect 3461 9164 3463 9168
rect 3477 9164 3479 9168
rect 3493 9164 3495 9168
rect 3514 9164 3516 9168
rect 3519 9164 3521 9168
rect 3535 9164 3537 9168
rect 3551 9164 3553 9168
rect 3556 9164 3558 9168
rect 4006 9173 4008 9177
rect 4011 9173 4013 9177
rect 4087 9173 4089 9177
rect 4092 9173 4094 9177
rect 3061 9097 3063 9101
rect 3066 9097 3068 9101
rect 3140 9101 3142 9105
rect 3166 9097 3168 9101
rect 3171 9097 3173 9101
rect 3089 9093 3091 9097
rect 2861 9088 2863 9092
rect 2877 9088 2879 9092
rect 2893 9088 2895 9092
rect 2916 9088 2918 9092
rect 2921 9088 2923 9092
rect 2947 9088 2949 9092
rect 2968 9088 2970 9092
rect 2988 9088 2990 9092
rect 2993 9088 2995 9092
rect 3011 9088 3013 9092
rect 3194 9093 3196 9097
rect 3371 9072 3373 9076
rect 3397 9068 3399 9072
rect 3402 9068 3404 9072
rect 3425 9064 3427 9068
rect 4006 9097 4008 9101
rect 4011 9097 4013 9101
rect 4085 9101 4087 9105
rect 4111 9097 4113 9101
rect 4116 9097 4118 9101
rect 4034 9093 4036 9097
rect 3806 9088 3808 9092
rect 3822 9088 3824 9092
rect 3838 9088 3840 9092
rect 3861 9088 3863 9092
rect 3866 9088 3868 9092
rect 3892 9088 3894 9092
rect 3913 9088 3915 9092
rect 3933 9088 3935 9092
rect 3938 9088 3940 9092
rect 3956 9088 3958 9092
rect 4139 9093 4141 9097
rect 2861 9042 2863 9046
rect 2877 9042 2879 9046
rect 2893 9042 2895 9046
rect 2916 9042 2918 9046
rect 2921 9042 2923 9046
rect 2947 9042 2949 9046
rect 2968 9042 2970 9046
rect 2988 9042 2990 9046
rect 2993 9042 2995 9046
rect 3011 9042 3013 9046
rect 3061 9042 3063 9046
rect 3066 9042 3068 9046
rect 3166 9042 3168 9046
rect 3171 9042 3173 9046
rect 3557 9033 3559 9045
rect 3610 9033 3612 9045
rect 3806 9042 3808 9046
rect 3822 9042 3824 9046
rect 3838 9042 3840 9046
rect 3861 9042 3863 9046
rect 3866 9042 3868 9046
rect 3892 9042 3894 9046
rect 3913 9042 3915 9046
rect 3933 9042 3935 9046
rect 3938 9042 3940 9046
rect 3956 9042 3958 9046
rect 4006 9042 4008 9046
rect 4011 9042 4013 9046
rect 4111 9042 4113 9046
rect 4116 9042 4118 9046
rect 3397 9008 3399 9012
rect 3402 9008 3404 9012
rect 3061 8965 3063 8969
rect 3066 8965 3068 8969
rect 3116 8969 3118 8973
rect 3142 8965 3144 8969
rect 3147 8965 3149 8969
rect 3206 8969 3208 8973
rect 3232 8965 3234 8969
rect 3237 8965 3239 8969
rect 3089 8961 3091 8965
rect 2861 8956 2863 8960
rect 2877 8956 2879 8960
rect 2893 8956 2895 8960
rect 2916 8956 2918 8960
rect 2921 8956 2923 8960
rect 2947 8956 2949 8960
rect 2968 8956 2970 8960
rect 2988 8956 2990 8960
rect 2993 8956 2995 8960
rect 3011 8956 3013 8960
rect 3170 8961 3172 8965
rect 3260 8961 3262 8965
rect 3349 8942 3351 8946
rect 3371 8942 3373 8946
rect 3397 8938 3399 8942
rect 3402 8938 3404 8942
rect 3425 8934 3427 8938
rect 4006 8965 4008 8969
rect 4011 8965 4013 8969
rect 4061 8969 4063 8973
rect 4087 8965 4089 8969
rect 4092 8965 4094 8969
rect 4151 8969 4153 8973
rect 4177 8965 4179 8969
rect 4182 8965 4184 8969
rect 4034 8961 4036 8965
rect 3806 8956 3808 8960
rect 3822 8956 3824 8960
rect 3838 8956 3840 8960
rect 3861 8956 3863 8960
rect 3866 8956 3868 8960
rect 3892 8956 3894 8960
rect 3913 8956 3915 8960
rect 3933 8956 3935 8960
rect 3938 8956 3940 8960
rect 3956 8956 3958 8960
rect 4115 8961 4117 8965
rect 4205 8961 4207 8965
rect 2861 8910 2863 8914
rect 2877 8910 2879 8914
rect 2893 8910 2895 8914
rect 2916 8910 2918 8914
rect 2921 8910 2923 8914
rect 2947 8910 2949 8914
rect 2968 8910 2970 8914
rect 2988 8910 2990 8914
rect 2993 8910 2995 8914
rect 3011 8910 3013 8914
rect 3061 8907 3063 8911
rect 3066 8907 3068 8911
rect 3142 8907 3144 8911
rect 3147 8907 3149 8911
rect 3232 8907 3234 8911
rect 3237 8907 3239 8911
rect 3463 8903 3465 8915
rect 3516 8903 3518 8915
rect 3806 8910 3808 8914
rect 3822 8910 3824 8914
rect 3838 8910 3840 8914
rect 3861 8910 3863 8914
rect 3866 8910 3868 8914
rect 3892 8910 3894 8914
rect 3913 8910 3915 8914
rect 3933 8910 3935 8914
rect 3938 8910 3940 8914
rect 3956 8910 3958 8914
rect 4006 8907 4008 8911
rect 4011 8907 4013 8911
rect 4087 8907 4089 8911
rect 4092 8907 4094 8911
rect 4177 8907 4179 8911
rect 4182 8907 4184 8911
rect 3397 8878 3399 8882
rect 3402 8878 3404 8882
rect 3061 8833 3063 8837
rect 3066 8833 3068 8837
rect 3089 8829 3091 8833
rect 2861 8824 2863 8828
rect 2877 8824 2879 8828
rect 2893 8824 2895 8828
rect 2916 8824 2918 8828
rect 2921 8824 2923 8828
rect 2947 8824 2949 8828
rect 2968 8824 2970 8828
rect 2988 8824 2990 8828
rect 2993 8824 2995 8828
rect 3011 8824 3013 8828
rect 4006 8833 4008 8837
rect 4011 8833 4013 8837
rect 4034 8829 4036 8833
rect 3806 8824 3808 8828
rect 3822 8824 3824 8828
rect 3838 8824 3840 8828
rect 3861 8824 3863 8828
rect 3866 8824 3868 8828
rect 3892 8824 3894 8828
rect 3913 8824 3915 8828
rect 3933 8824 3935 8828
rect 3938 8824 3940 8828
rect 3956 8824 3958 8828
rect 2861 8778 2863 8782
rect 2877 8778 2879 8782
rect 2893 8778 2895 8782
rect 2916 8778 2918 8782
rect 2921 8778 2923 8782
rect 2947 8778 2949 8782
rect 2968 8778 2970 8782
rect 2988 8778 2990 8782
rect 2993 8778 2995 8782
rect 3011 8778 3013 8782
rect 3095 8778 3097 8782
rect 3113 8778 3115 8782
rect 3138 8778 3140 8782
rect 3154 8778 3156 8782
rect 3177 8778 3179 8782
rect 3182 8778 3184 8782
rect 3208 8778 3210 8782
rect 3229 8778 3231 8782
rect 3249 8778 3251 8782
rect 3254 8778 3256 8782
rect 3272 8778 3274 8782
rect 2372 8764 2374 8768
rect 2377 8764 2379 8768
rect 2393 8764 2395 8768
rect 2409 8764 2411 8768
rect 2414 8764 2416 8768
rect 2435 8764 2437 8768
rect 2451 8764 2453 8768
rect 2467 8764 2469 8768
rect 2472 8764 2474 8768
rect 2488 8764 2490 8768
rect 2504 8764 2506 8768
rect 2509 8764 2511 8768
rect 2525 8764 2527 8768
rect 2541 8764 2543 8768
rect 2546 8764 2548 8768
rect 2567 8764 2569 8768
rect 2583 8764 2585 8768
rect 2599 8764 2601 8768
rect 2604 8764 2606 8768
rect 2620 8764 2622 8768
rect 2636 8764 2638 8768
rect 2641 8764 2643 8768
rect 2657 8764 2659 8768
rect 2673 8764 2675 8768
rect 2678 8764 2680 8768
rect 2699 8764 2701 8768
rect 2715 8764 2717 8768
rect 2731 8764 2733 8768
rect 2736 8764 2738 8768
rect 2752 8764 2754 8768
rect 3061 8771 3063 8775
rect 3066 8771 3068 8775
rect 3806 8778 3808 8782
rect 3822 8778 3824 8782
rect 3838 8778 3840 8782
rect 3861 8778 3863 8782
rect 3866 8778 3868 8782
rect 3892 8778 3894 8782
rect 3913 8778 3915 8782
rect 3933 8778 3935 8782
rect 3938 8778 3940 8782
rect 3956 8778 3958 8782
rect 4040 8778 4042 8782
rect 4058 8778 4060 8782
rect 4083 8778 4085 8782
rect 4099 8778 4101 8782
rect 4122 8778 4124 8782
rect 4127 8778 4129 8782
rect 4153 8778 4155 8782
rect 4174 8778 4176 8782
rect 4194 8778 4196 8782
rect 4199 8778 4201 8782
rect 4217 8778 4219 8782
rect 3317 8764 3319 8768
rect 3322 8764 3324 8768
rect 3338 8764 3340 8768
rect 3354 8764 3356 8768
rect 3359 8764 3361 8768
rect 3380 8764 3382 8768
rect 3396 8764 3398 8768
rect 3412 8764 3414 8768
rect 3417 8764 3419 8768
rect 3433 8764 3435 8768
rect 3449 8764 3451 8768
rect 3454 8764 3456 8768
rect 3470 8764 3472 8768
rect 3486 8764 3488 8768
rect 3491 8764 3493 8768
rect 3512 8764 3514 8768
rect 3528 8764 3530 8768
rect 3544 8764 3546 8768
rect 3549 8764 3551 8768
rect 3565 8764 3567 8768
rect 3581 8764 3583 8768
rect 3586 8764 3588 8768
rect 3602 8764 3604 8768
rect 3618 8764 3620 8768
rect 3623 8764 3625 8768
rect 3644 8764 3646 8768
rect 3660 8764 3662 8768
rect 3676 8764 3678 8768
rect 3681 8764 3683 8768
rect 3697 8764 3699 8768
rect 4006 8771 4008 8775
rect 4011 8771 4013 8775
rect 2487 8720 2489 8724
rect 2511 8720 2513 8724
rect 3284 8722 3288 8724
rect 3432 8720 3434 8724
rect 3456 8720 3458 8724
rect 4229 8722 4233 8724
rect 2507 8707 2509 8711
rect 3452 8707 3454 8711
rect 2498 8693 2502 8695
rect 3443 8693 3447 8695
rect 2487 8684 2489 8688
rect 2511 8684 2513 8688
rect 3432 8684 3434 8688
rect 3456 8684 3458 8688
rect 3155 8652 3157 8656
rect 3160 8652 3162 8656
rect 3176 8652 3178 8656
rect 3192 8652 3194 8656
rect 3197 8652 3199 8656
rect 3218 8652 3220 8656
rect 3234 8652 3236 8656
rect 3250 8652 3252 8656
rect 3255 8652 3257 8656
rect 3271 8652 3273 8656
rect 4100 8652 4102 8656
rect 4105 8652 4107 8656
rect 4121 8652 4123 8656
rect 4137 8652 4139 8656
rect 4142 8652 4144 8656
rect 4163 8652 4165 8656
rect 4179 8652 4181 8656
rect 4195 8652 4197 8656
rect 4200 8652 4202 8656
rect 4216 8652 4218 8656
rect 2372 8622 2374 8626
rect 2377 8622 2379 8626
rect 2393 8622 2395 8626
rect 2409 8622 2411 8626
rect 2414 8622 2416 8626
rect 2435 8622 2437 8626
rect 2451 8622 2453 8626
rect 2467 8622 2469 8626
rect 2472 8622 2474 8626
rect 2488 8622 2490 8626
rect 2504 8622 2506 8626
rect 2509 8622 2511 8626
rect 2525 8622 2527 8626
rect 2541 8622 2543 8626
rect 2546 8622 2548 8626
rect 2567 8622 2569 8626
rect 2583 8622 2585 8626
rect 2599 8622 2601 8626
rect 2604 8622 2606 8626
rect 2620 8622 2622 8626
rect 2636 8622 2638 8626
rect 2641 8622 2643 8626
rect 2657 8622 2659 8626
rect 2673 8622 2675 8626
rect 2678 8622 2680 8626
rect 2699 8622 2701 8626
rect 2715 8622 2717 8626
rect 2731 8622 2733 8626
rect 2736 8622 2738 8626
rect 2752 8622 2754 8626
rect 3317 8622 3319 8626
rect 3322 8622 3324 8626
rect 3338 8622 3340 8626
rect 3354 8622 3356 8626
rect 3359 8622 3361 8626
rect 3380 8622 3382 8626
rect 3396 8622 3398 8626
rect 3412 8622 3414 8626
rect 3417 8622 3419 8626
rect 3433 8622 3435 8626
rect 3449 8622 3451 8626
rect 3454 8622 3456 8626
rect 3470 8622 3472 8626
rect 3486 8622 3488 8626
rect 3491 8622 3493 8626
rect 3512 8622 3514 8626
rect 3528 8622 3530 8626
rect 3544 8622 3546 8626
rect 3549 8622 3551 8626
rect 3565 8622 3567 8626
rect 3581 8622 3583 8626
rect 3586 8622 3588 8626
rect 3602 8622 3604 8626
rect 3618 8622 3620 8626
rect 3623 8622 3625 8626
rect 3644 8622 3646 8626
rect 3660 8622 3662 8626
rect 3676 8622 3678 8626
rect 3681 8622 3683 8626
rect 3697 8622 3699 8626
rect 3296 8576 3300 8578
rect 4241 8576 4245 8578
rect 3155 8566 3157 8570
rect 3160 8566 3162 8570
rect 3176 8566 3178 8570
rect 3192 8566 3194 8570
rect 3197 8566 3199 8570
rect 3218 8566 3220 8570
rect 3234 8566 3236 8570
rect 3250 8566 3252 8570
rect 3255 8566 3257 8570
rect 3271 8566 3273 8570
rect 4100 8566 4102 8570
rect 4105 8566 4107 8570
rect 4121 8566 4123 8570
rect 4137 8566 4139 8570
rect 4142 8566 4144 8570
rect 4163 8566 4165 8570
rect 4179 8566 4181 8570
rect 4195 8566 4197 8570
rect 4200 8566 4202 8570
rect 4216 8566 4218 8570
rect 2372 8536 2374 8540
rect 2377 8536 2379 8540
rect 2393 8536 2395 8540
rect 2409 8536 2411 8540
rect 2414 8536 2416 8540
rect 2435 8536 2437 8540
rect 2451 8536 2453 8540
rect 2467 8536 2469 8540
rect 2472 8536 2474 8540
rect 2488 8536 2490 8540
rect 2504 8536 2506 8540
rect 2509 8536 2511 8540
rect 2525 8536 2527 8540
rect 2541 8536 2543 8540
rect 2546 8536 2548 8540
rect 2567 8536 2569 8540
rect 2583 8536 2585 8540
rect 2599 8536 2601 8540
rect 2604 8536 2606 8540
rect 2620 8536 2622 8540
rect 2636 8536 2638 8540
rect 2641 8536 2643 8540
rect 2657 8536 2659 8540
rect 2673 8536 2675 8540
rect 2678 8536 2680 8540
rect 2699 8536 2701 8540
rect 2715 8536 2717 8540
rect 2731 8536 2733 8540
rect 2736 8536 2738 8540
rect 2752 8536 2754 8540
rect 3317 8536 3319 8540
rect 3322 8536 3324 8540
rect 3338 8536 3340 8540
rect 3354 8536 3356 8540
rect 3359 8536 3361 8540
rect 3380 8536 3382 8540
rect 3396 8536 3398 8540
rect 3412 8536 3414 8540
rect 3417 8536 3419 8540
rect 3433 8536 3435 8540
rect 3449 8536 3451 8540
rect 3454 8536 3456 8540
rect 3470 8536 3472 8540
rect 3486 8536 3488 8540
rect 3491 8536 3493 8540
rect 3512 8536 3514 8540
rect 3528 8536 3530 8540
rect 3544 8536 3546 8540
rect 3549 8536 3551 8540
rect 3565 8536 3567 8540
rect 3581 8536 3583 8540
rect 3586 8536 3588 8540
rect 3602 8536 3604 8540
rect 3618 8536 3620 8540
rect 3623 8536 3625 8540
rect 3644 8536 3646 8540
rect 3660 8536 3662 8540
rect 3676 8536 3678 8540
rect 3681 8536 3683 8540
rect 3697 8536 3699 8540
rect 2604 8492 2606 8496
rect 2628 8492 2630 8496
rect 3549 8492 3551 8496
rect 3573 8492 3575 8496
rect 2624 8481 2626 8485
rect 3569 8481 3571 8485
rect 2615 8467 2619 8469
rect 3560 8467 3564 8469
rect 2604 8458 2606 8462
rect 2628 8458 2630 8462
rect 3549 8458 3551 8462
rect 3573 8458 3575 8462
rect 2372 8396 2374 8400
rect 2377 8396 2379 8400
rect 2393 8396 2395 8400
rect 2409 8396 2411 8400
rect 2414 8396 2416 8400
rect 2435 8396 2437 8400
rect 2451 8396 2453 8400
rect 2467 8396 2469 8400
rect 2472 8396 2474 8400
rect 2488 8396 2490 8400
rect 2504 8396 2506 8400
rect 2509 8396 2511 8400
rect 2525 8396 2527 8400
rect 2541 8396 2543 8400
rect 2546 8396 2548 8400
rect 2567 8396 2569 8400
rect 2583 8396 2585 8400
rect 2599 8396 2601 8400
rect 2604 8396 2606 8400
rect 2620 8396 2622 8400
rect 2636 8396 2638 8400
rect 2641 8396 2643 8400
rect 2657 8396 2659 8400
rect 2673 8396 2675 8400
rect 2678 8396 2680 8400
rect 2699 8396 2701 8400
rect 2715 8396 2717 8400
rect 2731 8396 2733 8400
rect 2736 8396 2738 8400
rect 2752 8396 2754 8400
rect 3317 8396 3319 8400
rect 3322 8396 3324 8400
rect 3338 8396 3340 8400
rect 3354 8396 3356 8400
rect 3359 8396 3361 8400
rect 3380 8396 3382 8400
rect 3396 8396 3398 8400
rect 3412 8396 3414 8400
rect 3417 8396 3419 8400
rect 3433 8396 3435 8400
rect 3449 8396 3451 8400
rect 3454 8396 3456 8400
rect 3470 8396 3472 8400
rect 3486 8396 3488 8400
rect 3491 8396 3493 8400
rect 3512 8396 3514 8400
rect 3528 8396 3530 8400
rect 3544 8396 3546 8400
rect 3549 8396 3551 8400
rect 3565 8396 3567 8400
rect 3581 8396 3583 8400
rect 3586 8396 3588 8400
rect 3602 8396 3604 8400
rect 3618 8396 3620 8400
rect 3623 8396 3625 8400
rect 3644 8396 3646 8400
rect 3660 8396 3662 8400
rect 3676 8396 3678 8400
rect 3681 8396 3683 8400
rect 3697 8396 3699 8400
rect 2856 8317 2858 8321
rect 2861 8317 2863 8321
rect 2877 8317 2879 8321
rect 2893 8317 2895 8321
rect 2898 8317 2900 8321
rect 2919 8317 2921 8321
rect 2935 8317 2937 8321
rect 2951 8317 2953 8321
rect 2956 8317 2958 8321
rect 2972 8317 2974 8321
rect 2988 8317 2990 8321
rect 2993 8317 2995 8321
rect 3009 8317 3011 8321
rect 3025 8317 3027 8321
rect 3030 8317 3032 8321
rect 3051 8317 3053 8321
rect 3067 8317 3069 8321
rect 3083 8317 3085 8321
rect 3088 8317 3090 8321
rect 3104 8317 3106 8321
rect 3120 8317 3122 8321
rect 3125 8317 3127 8321
rect 3141 8317 3143 8321
rect 3157 8317 3159 8321
rect 3162 8317 3164 8321
rect 3183 8317 3185 8321
rect 3199 8317 3201 8321
rect 3215 8317 3217 8321
rect 3220 8317 3222 8321
rect 3236 8317 3238 8321
rect 3252 8317 3254 8321
rect 3257 8317 3259 8321
rect 3273 8317 3275 8321
rect 3289 8317 3291 8321
rect 3294 8317 3296 8321
rect 3315 8317 3317 8321
rect 3331 8317 3333 8321
rect 3347 8317 3349 8321
rect 3352 8317 3354 8321
rect 3368 8317 3370 8321
rect 3801 8317 3803 8321
rect 3806 8317 3808 8321
rect 3822 8317 3824 8321
rect 3838 8317 3840 8321
rect 3843 8317 3845 8321
rect 3864 8317 3866 8321
rect 3880 8317 3882 8321
rect 3896 8317 3898 8321
rect 3901 8317 3903 8321
rect 3917 8317 3919 8321
rect 3933 8317 3935 8321
rect 3938 8317 3940 8321
rect 3954 8317 3956 8321
rect 3970 8317 3972 8321
rect 3975 8317 3977 8321
rect 3996 8317 3998 8321
rect 4012 8317 4014 8321
rect 4028 8317 4030 8321
rect 4033 8317 4035 8321
rect 4049 8317 4051 8321
rect 4065 8317 4067 8321
rect 4070 8317 4072 8321
rect 4086 8317 4088 8321
rect 4102 8317 4104 8321
rect 4107 8317 4109 8321
rect 4128 8317 4130 8321
rect 4144 8317 4146 8321
rect 4160 8317 4162 8321
rect 4165 8317 4167 8321
rect 4181 8317 4183 8321
rect 4197 8317 4199 8321
rect 4202 8317 4204 8321
rect 4218 8317 4220 8321
rect 4234 8317 4236 8321
rect 4239 8317 4241 8321
rect 4260 8317 4262 8321
rect 4276 8317 4278 8321
rect 4292 8317 4294 8321
rect 4297 8317 4299 8321
rect 4313 8317 4315 8321
rect 2504 8284 2506 8288
rect 2509 8284 2511 8288
rect 2525 8284 2527 8288
rect 2541 8284 2543 8288
rect 2546 8284 2548 8288
rect 2567 8284 2569 8288
rect 2583 8284 2585 8288
rect 2599 8284 2601 8288
rect 2604 8284 2606 8288
rect 2620 8284 2622 8288
rect 3449 8284 3451 8288
rect 3454 8284 3456 8288
rect 3470 8284 3472 8288
rect 3486 8284 3488 8288
rect 3491 8284 3493 8288
rect 3512 8284 3514 8288
rect 3528 8284 3530 8288
rect 3544 8284 3546 8288
rect 3549 8284 3551 8288
rect 3565 8284 3567 8288
rect 2628 8247 2630 8251
rect 3035 8251 3037 8255
rect 3061 8247 3063 8251
rect 3066 8247 3068 8251
rect 3116 8251 3118 8255
rect 3142 8247 3144 8251
rect 3147 8247 3149 8251
rect 3089 8243 3091 8247
rect 2511 8238 2513 8242
rect 2861 8238 2863 8242
rect 2877 8238 2879 8242
rect 2893 8238 2895 8242
rect 2916 8238 2918 8242
rect 2921 8238 2923 8242
rect 2947 8238 2949 8242
rect 2968 8238 2970 8242
rect 2988 8238 2990 8242
rect 2993 8238 2995 8242
rect 3011 8238 3013 8242
rect 3170 8243 3172 8247
rect 3573 8247 3575 8251
rect 3980 8251 3982 8255
rect 4006 8247 4008 8251
rect 4011 8247 4013 8251
rect 4061 8251 4063 8255
rect 4087 8247 4089 8251
rect 4092 8247 4094 8251
rect 4034 8243 4036 8247
rect 3456 8238 3458 8242
rect 3806 8238 3808 8242
rect 3822 8238 3824 8242
rect 3838 8238 3840 8242
rect 3861 8238 3863 8242
rect 3866 8238 3868 8242
rect 3892 8238 3894 8242
rect 3913 8238 3915 8242
rect 3933 8238 3935 8242
rect 3938 8238 3940 8242
rect 3956 8238 3958 8242
rect 4115 8243 4117 8247
rect 2861 8192 2863 8196
rect 2877 8192 2879 8196
rect 2893 8192 2895 8196
rect 2916 8192 2918 8196
rect 2921 8192 2923 8196
rect 2947 8192 2949 8196
rect 2968 8192 2970 8196
rect 2988 8192 2990 8196
rect 2993 8192 2995 8196
rect 3011 8192 3013 8196
rect 2495 8182 2497 8186
rect 2511 8182 2513 8186
rect 2516 8182 2518 8186
rect 2532 8182 2534 8186
rect 2548 8182 2550 8186
rect 2569 8182 2571 8186
rect 2574 8182 2576 8186
rect 2590 8182 2592 8186
rect 2606 8182 2608 8186
rect 2611 8182 2613 8186
rect 3061 8191 3063 8195
rect 3066 8191 3068 8195
rect 3142 8191 3144 8195
rect 3147 8191 3149 8195
rect 3806 8192 3808 8196
rect 3822 8192 3824 8196
rect 3838 8192 3840 8196
rect 3861 8192 3863 8196
rect 3866 8192 3868 8196
rect 3892 8192 3894 8196
rect 3913 8192 3915 8196
rect 3933 8192 3935 8196
rect 3938 8192 3940 8196
rect 3956 8192 3958 8196
rect 3440 8182 3442 8186
rect 3456 8182 3458 8186
rect 3461 8182 3463 8186
rect 3477 8182 3479 8186
rect 3493 8182 3495 8186
rect 3514 8182 3516 8186
rect 3519 8182 3521 8186
rect 3535 8182 3537 8186
rect 3551 8182 3553 8186
rect 3556 8182 3558 8186
rect 4006 8191 4008 8195
rect 4011 8191 4013 8195
rect 4087 8191 4089 8195
rect 4092 8191 4094 8195
rect 3061 8115 3063 8119
rect 3066 8115 3068 8119
rect 3140 8119 3142 8123
rect 3166 8115 3168 8119
rect 3171 8115 3173 8119
rect 3089 8111 3091 8115
rect 2861 8106 2863 8110
rect 2877 8106 2879 8110
rect 2893 8106 2895 8110
rect 2916 8106 2918 8110
rect 2921 8106 2923 8110
rect 2947 8106 2949 8110
rect 2968 8106 2970 8110
rect 2988 8106 2990 8110
rect 2993 8106 2995 8110
rect 3011 8106 3013 8110
rect 3194 8111 3196 8115
rect 4006 8115 4008 8119
rect 4011 8115 4013 8119
rect 4085 8119 4087 8123
rect 4111 8115 4113 8119
rect 4116 8115 4118 8119
rect 4034 8111 4036 8115
rect 3806 8106 3808 8110
rect 3822 8106 3824 8110
rect 3838 8106 3840 8110
rect 3861 8106 3863 8110
rect 3866 8106 3868 8110
rect 3892 8106 3894 8110
rect 3913 8106 3915 8110
rect 3933 8106 3935 8110
rect 3938 8106 3940 8110
rect 3956 8106 3958 8110
rect 4139 8111 4141 8115
rect 2861 8060 2863 8064
rect 2877 8060 2879 8064
rect 2893 8060 2895 8064
rect 2916 8060 2918 8064
rect 2921 8060 2923 8064
rect 2947 8060 2949 8064
rect 2968 8060 2970 8064
rect 2988 8060 2990 8064
rect 2993 8060 2995 8064
rect 3011 8060 3013 8064
rect 3061 8060 3063 8064
rect 3066 8060 3068 8064
rect 3166 8060 3168 8064
rect 3171 8060 3173 8064
rect 3806 8060 3808 8064
rect 3822 8060 3824 8064
rect 3838 8060 3840 8064
rect 3861 8060 3863 8064
rect 3866 8060 3868 8064
rect 3892 8060 3894 8064
rect 3913 8060 3915 8064
rect 3933 8060 3935 8064
rect 3938 8060 3940 8064
rect 3956 8060 3958 8064
rect 4006 8060 4008 8064
rect 4011 8060 4013 8064
rect 4111 8060 4113 8064
rect 4116 8060 4118 8064
rect 3061 7983 3063 7987
rect 3066 7983 3068 7987
rect 3116 7987 3118 7991
rect 3142 7983 3144 7987
rect 3147 7983 3149 7987
rect 3206 7987 3208 7991
rect 3232 7983 3234 7987
rect 3237 7983 3239 7987
rect 3089 7979 3091 7983
rect 2861 7974 2863 7978
rect 2877 7974 2879 7978
rect 2893 7974 2895 7978
rect 2916 7974 2918 7978
rect 2921 7974 2923 7978
rect 2947 7974 2949 7978
rect 2968 7974 2970 7978
rect 2988 7974 2990 7978
rect 2993 7974 2995 7978
rect 3011 7974 3013 7978
rect 3170 7979 3172 7983
rect 3260 7979 3262 7983
rect 4006 7983 4008 7987
rect 4011 7983 4013 7987
rect 4061 7987 4063 7991
rect 4087 7983 4089 7987
rect 4092 7983 4094 7987
rect 4151 7987 4153 7991
rect 4177 7983 4179 7987
rect 4182 7983 4184 7987
rect 4034 7979 4036 7983
rect 3806 7974 3808 7978
rect 3822 7974 3824 7978
rect 3838 7974 3840 7978
rect 3861 7974 3863 7978
rect 3866 7974 3868 7978
rect 3892 7974 3894 7978
rect 3913 7974 3915 7978
rect 3933 7974 3935 7978
rect 3938 7974 3940 7978
rect 3956 7974 3958 7978
rect 4115 7979 4117 7983
rect 4205 7979 4207 7983
rect 2861 7928 2863 7932
rect 2877 7928 2879 7932
rect 2893 7928 2895 7932
rect 2916 7928 2918 7932
rect 2921 7928 2923 7932
rect 2947 7928 2949 7932
rect 2968 7928 2970 7932
rect 2988 7928 2990 7932
rect 2993 7928 2995 7932
rect 3011 7928 3013 7932
rect 3061 7925 3063 7929
rect 3066 7925 3068 7929
rect 3142 7925 3144 7929
rect 3147 7925 3149 7929
rect 3232 7925 3234 7929
rect 3237 7925 3239 7929
rect 3806 7928 3808 7932
rect 3822 7928 3824 7932
rect 3838 7928 3840 7932
rect 3861 7928 3863 7932
rect 3866 7928 3868 7932
rect 3892 7928 3894 7932
rect 3913 7928 3915 7932
rect 3933 7928 3935 7932
rect 3938 7928 3940 7932
rect 3956 7928 3958 7932
rect 4006 7925 4008 7929
rect 4011 7925 4013 7929
rect 4087 7925 4089 7929
rect 4092 7925 4094 7929
rect 4177 7925 4179 7929
rect 4182 7925 4184 7929
rect 3061 7851 3063 7855
rect 3066 7851 3068 7855
rect 3089 7847 3091 7851
rect 2861 7842 2863 7846
rect 2877 7842 2879 7846
rect 2893 7842 2895 7846
rect 2916 7842 2918 7846
rect 2921 7842 2923 7846
rect 2947 7842 2949 7846
rect 2968 7842 2970 7846
rect 2988 7842 2990 7846
rect 2993 7842 2995 7846
rect 3011 7842 3013 7846
rect 4006 7851 4008 7855
rect 4011 7851 4013 7855
rect 4034 7847 4036 7851
rect 3806 7842 3808 7846
rect 3822 7842 3824 7846
rect 3838 7842 3840 7846
rect 3861 7842 3863 7846
rect 3866 7842 3868 7846
rect 3892 7842 3894 7846
rect 3913 7842 3915 7846
rect 3933 7842 3935 7846
rect 3938 7842 3940 7846
rect 3956 7842 3958 7846
rect 2861 7796 2863 7800
rect 2877 7796 2879 7800
rect 2893 7796 2895 7800
rect 2916 7796 2918 7800
rect 2921 7796 2923 7800
rect 2947 7796 2949 7800
rect 2968 7796 2970 7800
rect 2988 7796 2990 7800
rect 2993 7796 2995 7800
rect 3011 7796 3013 7800
rect 3095 7796 3097 7800
rect 3113 7796 3115 7800
rect 3138 7796 3140 7800
rect 3154 7796 3156 7800
rect 3177 7796 3179 7800
rect 3182 7796 3184 7800
rect 3208 7796 3210 7800
rect 3229 7796 3231 7800
rect 3249 7796 3251 7800
rect 3254 7796 3256 7800
rect 3272 7796 3274 7800
rect 2372 7782 2374 7786
rect 2377 7782 2379 7786
rect 2393 7782 2395 7786
rect 2409 7782 2411 7786
rect 2414 7782 2416 7786
rect 2435 7782 2437 7786
rect 2451 7782 2453 7786
rect 2467 7782 2469 7786
rect 2472 7782 2474 7786
rect 2488 7782 2490 7786
rect 2504 7782 2506 7786
rect 2509 7782 2511 7786
rect 2525 7782 2527 7786
rect 2541 7782 2543 7786
rect 2546 7782 2548 7786
rect 2567 7782 2569 7786
rect 2583 7782 2585 7786
rect 2599 7782 2601 7786
rect 2604 7782 2606 7786
rect 2620 7782 2622 7786
rect 2636 7782 2638 7786
rect 2641 7782 2643 7786
rect 2657 7782 2659 7786
rect 2673 7782 2675 7786
rect 2678 7782 2680 7786
rect 2699 7782 2701 7786
rect 2715 7782 2717 7786
rect 2731 7782 2733 7786
rect 2736 7782 2738 7786
rect 2752 7782 2754 7786
rect 3061 7789 3063 7793
rect 3066 7789 3068 7793
rect 3806 7796 3808 7800
rect 3822 7796 3824 7800
rect 3838 7796 3840 7800
rect 3861 7796 3863 7800
rect 3866 7796 3868 7800
rect 3892 7796 3894 7800
rect 3913 7796 3915 7800
rect 3933 7796 3935 7800
rect 3938 7796 3940 7800
rect 3956 7796 3958 7800
rect 4040 7796 4042 7800
rect 4058 7796 4060 7800
rect 4083 7796 4085 7800
rect 4099 7796 4101 7800
rect 4122 7796 4124 7800
rect 4127 7796 4129 7800
rect 4153 7796 4155 7800
rect 4174 7796 4176 7800
rect 4194 7796 4196 7800
rect 4199 7796 4201 7800
rect 4217 7796 4219 7800
rect 3317 7782 3319 7786
rect 3322 7782 3324 7786
rect 3338 7782 3340 7786
rect 3354 7782 3356 7786
rect 3359 7782 3361 7786
rect 3380 7782 3382 7786
rect 3396 7782 3398 7786
rect 3412 7782 3414 7786
rect 3417 7782 3419 7786
rect 3433 7782 3435 7786
rect 3449 7782 3451 7786
rect 3454 7782 3456 7786
rect 3470 7782 3472 7786
rect 3486 7782 3488 7786
rect 3491 7782 3493 7786
rect 3512 7782 3514 7786
rect 3528 7782 3530 7786
rect 3544 7782 3546 7786
rect 3549 7782 3551 7786
rect 3565 7782 3567 7786
rect 3581 7782 3583 7786
rect 3586 7782 3588 7786
rect 3602 7782 3604 7786
rect 3618 7782 3620 7786
rect 3623 7782 3625 7786
rect 3644 7782 3646 7786
rect 3660 7782 3662 7786
rect 3676 7782 3678 7786
rect 3681 7782 3683 7786
rect 3697 7782 3699 7786
rect 4006 7789 4008 7793
rect 4011 7789 4013 7793
rect 2487 7738 2489 7742
rect 2511 7738 2513 7742
rect 3284 7740 3288 7742
rect 3432 7738 3434 7742
rect 3456 7738 3458 7742
rect 4229 7740 4233 7742
rect 2507 7725 2509 7729
rect 3452 7725 3454 7729
rect 2498 7711 2502 7713
rect 3443 7711 3447 7713
rect 2487 7702 2489 7706
rect 2511 7702 2513 7706
rect 3432 7702 3434 7706
rect 3456 7702 3458 7706
rect 3155 7670 3157 7674
rect 3160 7670 3162 7674
rect 3176 7670 3178 7674
rect 3192 7670 3194 7674
rect 3197 7670 3199 7674
rect 3218 7670 3220 7674
rect 3234 7670 3236 7674
rect 3250 7670 3252 7674
rect 3255 7670 3257 7674
rect 3271 7670 3273 7674
rect 4100 7670 4102 7674
rect 4105 7670 4107 7674
rect 4121 7670 4123 7674
rect 4137 7670 4139 7674
rect 4142 7670 4144 7674
rect 4163 7670 4165 7674
rect 4179 7670 4181 7674
rect 4195 7670 4197 7674
rect 4200 7670 4202 7674
rect 4216 7670 4218 7674
rect 2372 7640 2374 7644
rect 2377 7640 2379 7644
rect 2393 7640 2395 7644
rect 2409 7640 2411 7644
rect 2414 7640 2416 7644
rect 2435 7640 2437 7644
rect 2451 7640 2453 7644
rect 2467 7640 2469 7644
rect 2472 7640 2474 7644
rect 2488 7640 2490 7644
rect 2504 7640 2506 7644
rect 2509 7640 2511 7644
rect 2525 7640 2527 7644
rect 2541 7640 2543 7644
rect 2546 7640 2548 7644
rect 2567 7640 2569 7644
rect 2583 7640 2585 7644
rect 2599 7640 2601 7644
rect 2604 7640 2606 7644
rect 2620 7640 2622 7644
rect 2636 7640 2638 7644
rect 2641 7640 2643 7644
rect 2657 7640 2659 7644
rect 2673 7640 2675 7644
rect 2678 7640 2680 7644
rect 2699 7640 2701 7644
rect 2715 7640 2717 7644
rect 2731 7640 2733 7644
rect 2736 7640 2738 7644
rect 2752 7640 2754 7644
rect 3317 7640 3319 7644
rect 3322 7640 3324 7644
rect 3338 7640 3340 7644
rect 3354 7640 3356 7644
rect 3359 7640 3361 7644
rect 3380 7640 3382 7644
rect 3396 7640 3398 7644
rect 3412 7640 3414 7644
rect 3417 7640 3419 7644
rect 3433 7640 3435 7644
rect 3449 7640 3451 7644
rect 3454 7640 3456 7644
rect 3470 7640 3472 7644
rect 3486 7640 3488 7644
rect 3491 7640 3493 7644
rect 3512 7640 3514 7644
rect 3528 7640 3530 7644
rect 3544 7640 3546 7644
rect 3549 7640 3551 7644
rect 3565 7640 3567 7644
rect 3581 7640 3583 7644
rect 3586 7640 3588 7644
rect 3602 7640 3604 7644
rect 3618 7640 3620 7644
rect 3623 7640 3625 7644
rect 3644 7640 3646 7644
rect 3660 7640 3662 7644
rect 3676 7640 3678 7644
rect 3681 7640 3683 7644
rect 3697 7640 3699 7644
rect 3296 7594 3300 7596
rect 4241 7594 4245 7596
rect 3155 7584 3157 7588
rect 3160 7584 3162 7588
rect 3176 7584 3178 7588
rect 3192 7584 3194 7588
rect 3197 7584 3199 7588
rect 3218 7584 3220 7588
rect 3234 7584 3236 7588
rect 3250 7584 3252 7588
rect 3255 7584 3257 7588
rect 3271 7584 3273 7588
rect 4100 7584 4102 7588
rect 4105 7584 4107 7588
rect 4121 7584 4123 7588
rect 4137 7584 4139 7588
rect 4142 7584 4144 7588
rect 4163 7584 4165 7588
rect 4179 7584 4181 7588
rect 4195 7584 4197 7588
rect 4200 7584 4202 7588
rect 4216 7584 4218 7588
rect 2372 7554 2374 7558
rect 2377 7554 2379 7558
rect 2393 7554 2395 7558
rect 2409 7554 2411 7558
rect 2414 7554 2416 7558
rect 2435 7554 2437 7558
rect 2451 7554 2453 7558
rect 2467 7554 2469 7558
rect 2472 7554 2474 7558
rect 2488 7554 2490 7558
rect 2504 7554 2506 7558
rect 2509 7554 2511 7558
rect 2525 7554 2527 7558
rect 2541 7554 2543 7558
rect 2546 7554 2548 7558
rect 2567 7554 2569 7558
rect 2583 7554 2585 7558
rect 2599 7554 2601 7558
rect 2604 7554 2606 7558
rect 2620 7554 2622 7558
rect 2636 7554 2638 7558
rect 2641 7554 2643 7558
rect 2657 7554 2659 7558
rect 2673 7554 2675 7558
rect 2678 7554 2680 7558
rect 2699 7554 2701 7558
rect 2715 7554 2717 7558
rect 2731 7554 2733 7558
rect 2736 7554 2738 7558
rect 2752 7554 2754 7558
rect 3317 7554 3319 7558
rect 3322 7554 3324 7558
rect 3338 7554 3340 7558
rect 3354 7554 3356 7558
rect 3359 7554 3361 7558
rect 3380 7554 3382 7558
rect 3396 7554 3398 7558
rect 3412 7554 3414 7558
rect 3417 7554 3419 7558
rect 3433 7554 3435 7558
rect 3449 7554 3451 7558
rect 3454 7554 3456 7558
rect 3470 7554 3472 7558
rect 3486 7554 3488 7558
rect 3491 7554 3493 7558
rect 3512 7554 3514 7558
rect 3528 7554 3530 7558
rect 3544 7554 3546 7558
rect 3549 7554 3551 7558
rect 3565 7554 3567 7558
rect 3581 7554 3583 7558
rect 3586 7554 3588 7558
rect 3602 7554 3604 7558
rect 3618 7554 3620 7558
rect 3623 7554 3625 7558
rect 3644 7554 3646 7558
rect 3660 7554 3662 7558
rect 3676 7554 3678 7558
rect 3681 7554 3683 7558
rect 3697 7554 3699 7558
rect 2604 7510 2606 7514
rect 2628 7510 2630 7514
rect 3549 7510 3551 7514
rect 3573 7510 3575 7514
rect 2624 7499 2626 7503
rect 3569 7499 3571 7503
rect 2615 7485 2619 7487
rect 3560 7485 3564 7487
rect 2604 7476 2606 7480
rect 2628 7476 2630 7480
rect 3549 7476 3551 7480
rect 3573 7476 3575 7480
rect 2372 7414 2374 7418
rect 2377 7414 2379 7418
rect 2393 7414 2395 7418
rect 2409 7414 2411 7418
rect 2414 7414 2416 7418
rect 2435 7414 2437 7418
rect 2451 7414 2453 7418
rect 2467 7414 2469 7418
rect 2472 7414 2474 7418
rect 2488 7414 2490 7418
rect 2504 7414 2506 7418
rect 2509 7414 2511 7418
rect 2525 7414 2527 7418
rect 2541 7414 2543 7418
rect 2546 7414 2548 7418
rect 2567 7414 2569 7418
rect 2583 7414 2585 7418
rect 2599 7414 2601 7418
rect 2604 7414 2606 7418
rect 2620 7414 2622 7418
rect 2636 7414 2638 7418
rect 2641 7414 2643 7418
rect 2657 7414 2659 7418
rect 2673 7414 2675 7418
rect 2678 7414 2680 7418
rect 2699 7414 2701 7418
rect 2715 7414 2717 7418
rect 2731 7414 2733 7418
rect 2736 7414 2738 7418
rect 2752 7414 2754 7418
rect 3317 7414 3319 7418
rect 3322 7414 3324 7418
rect 3338 7414 3340 7418
rect 3354 7414 3356 7418
rect 3359 7414 3361 7418
rect 3380 7414 3382 7418
rect 3396 7414 3398 7418
rect 3412 7414 3414 7418
rect 3417 7414 3419 7418
rect 3433 7414 3435 7418
rect 3449 7414 3451 7418
rect 3454 7414 3456 7418
rect 3470 7414 3472 7418
rect 3486 7414 3488 7418
rect 3491 7414 3493 7418
rect 3512 7414 3514 7418
rect 3528 7414 3530 7418
rect 3544 7414 3546 7418
rect 3549 7414 3551 7418
rect 3565 7414 3567 7418
rect 3581 7414 3583 7418
rect 3586 7414 3588 7418
rect 3602 7414 3604 7418
rect 3618 7414 3620 7418
rect 3623 7414 3625 7418
rect 3644 7414 3646 7418
rect 3660 7414 3662 7418
rect 3676 7414 3678 7418
rect 3681 7414 3683 7418
rect 3697 7414 3699 7418
rect 4579 7975 4581 8015
rect 4587 7975 4589 8015
rect 4595 7975 4597 8015
rect 4603 7975 4605 8015
rect 4611 7975 4613 8015
rect 4619 7975 4621 8015
rect 4634 7975 4636 8034
rect 4642 7975 4644 8034
rect 4650 7975 4652 8034
rect 4658 7975 4660 8034
rect 4677 7975 4679 8034
rect 4685 7975 4687 8034
rect 4693 7975 4695 8034
rect 4701 7975 4703 8034
rect 4718 7975 4720 8034
rect 4726 7975 4728 8034
rect 4734 7975 4736 8034
rect 4742 7975 4744 8034
<< ptransistor >>
rect 1743 9824 1799 9826
rect 2052 9824 2108 9826
rect 2361 9824 2417 9826
rect 2670 9824 2726 9826
rect 2979 9824 3035 9826
rect 3906 9824 3962 9826
rect 1743 9816 1799 9818
rect 2052 9816 2108 9818
rect 2361 9816 2417 9818
rect 2670 9816 2726 9818
rect 2979 9816 3035 9818
rect 3906 9816 3962 9818
rect 1743 9808 1799 9810
rect 1743 9800 1799 9802
rect 1743 9792 1799 9794
rect 1743 9784 1799 9786
rect 2052 9808 2108 9810
rect 2052 9800 2108 9802
rect 2052 9792 2108 9794
rect 2052 9784 2108 9786
rect 2361 9808 2417 9810
rect 2361 9800 2417 9802
rect 2361 9792 2417 9794
rect 2361 9784 2417 9786
rect 2670 9808 2726 9810
rect 2670 9800 2726 9802
rect 2670 9792 2726 9794
rect 2670 9784 2726 9786
rect 2979 9808 3035 9810
rect 2979 9800 3035 9802
rect 2979 9792 3035 9794
rect 2979 9784 3035 9786
rect 3906 9808 3962 9810
rect 3906 9800 3962 9802
rect 3906 9792 3962 9794
rect 3906 9784 3962 9786
rect 2856 9322 2858 9330
rect 2861 9322 2863 9330
rect 2877 9322 2879 9330
rect 2893 9322 2895 9330
rect 2898 9322 2900 9330
rect 2919 9322 2921 9330
rect 2935 9322 2937 9330
rect 2951 9322 2953 9330
rect 2956 9322 2958 9330
rect 2972 9322 2974 9330
rect 2988 9322 2990 9330
rect 2993 9322 2995 9330
rect 3009 9322 3011 9330
rect 3025 9322 3027 9330
rect 3030 9322 3032 9330
rect 3051 9322 3053 9330
rect 3067 9322 3069 9330
rect 3083 9322 3085 9330
rect 3088 9322 3090 9330
rect 3104 9322 3106 9330
rect 3120 9322 3122 9330
rect 3125 9322 3127 9330
rect 3141 9322 3143 9330
rect 3157 9322 3159 9330
rect 3162 9322 3164 9330
rect 3183 9322 3185 9330
rect 3199 9322 3201 9330
rect 3215 9322 3217 9330
rect 3220 9322 3222 9330
rect 3236 9322 3238 9330
rect 3252 9322 3254 9330
rect 3257 9322 3259 9330
rect 3273 9322 3275 9330
rect 3289 9322 3291 9330
rect 3294 9322 3296 9330
rect 3315 9322 3317 9330
rect 3331 9322 3333 9330
rect 3347 9322 3349 9330
rect 3352 9322 3354 9330
rect 3368 9322 3370 9330
rect 3801 9322 3803 9330
rect 3806 9322 3808 9330
rect 3822 9322 3824 9330
rect 3838 9322 3840 9330
rect 3843 9322 3845 9330
rect 3864 9322 3866 9330
rect 3880 9322 3882 9330
rect 3896 9322 3898 9330
rect 3901 9322 3903 9330
rect 3917 9322 3919 9330
rect 3933 9322 3935 9330
rect 3938 9322 3940 9330
rect 3954 9322 3956 9330
rect 3970 9322 3972 9330
rect 3975 9322 3977 9330
rect 3996 9322 3998 9330
rect 4012 9322 4014 9330
rect 4028 9322 4030 9330
rect 4033 9322 4035 9330
rect 4049 9322 4051 9330
rect 4065 9322 4067 9330
rect 4070 9322 4072 9330
rect 4086 9322 4088 9330
rect 4102 9322 4104 9330
rect 4107 9322 4109 9330
rect 4128 9322 4130 9330
rect 4144 9322 4146 9330
rect 4160 9322 4162 9330
rect 4165 9322 4167 9330
rect 4181 9322 4183 9330
rect 4197 9322 4199 9330
rect 4202 9322 4204 9330
rect 4218 9322 4220 9330
rect 4234 9322 4236 9330
rect 4239 9322 4241 9330
rect 4260 9322 4262 9330
rect 4276 9322 4278 9330
rect 4292 9322 4294 9330
rect 4297 9322 4299 9330
rect 4313 9322 4315 9330
rect 2504 9289 2506 9297
rect 2509 9289 2511 9297
rect 2525 9289 2527 9297
rect 2541 9289 2543 9297
rect 2546 9289 2548 9297
rect 2567 9289 2569 9297
rect 2583 9289 2585 9297
rect 2599 9289 2601 9297
rect 2604 9289 2606 9297
rect 2620 9289 2622 9297
rect 3449 9289 3451 9297
rect 3454 9289 3456 9297
rect 3470 9289 3472 9297
rect 3486 9289 3488 9297
rect 3491 9289 3493 9297
rect 3512 9289 3514 9297
rect 3528 9289 3530 9297
rect 3544 9289 3546 9297
rect 3549 9289 3551 9297
rect 3565 9289 3567 9297
rect 3035 9251 3037 9259
rect 2861 9238 2863 9246
rect 2877 9238 2879 9246
rect 2893 9238 2895 9246
rect 2916 9238 2918 9246
rect 2921 9238 2923 9246
rect 2947 9238 2949 9246
rect 2968 9238 2970 9246
rect 2988 9238 2990 9246
rect 2993 9238 2995 9246
rect 3011 9238 3013 9246
rect 3061 9245 3063 9253
rect 3066 9245 3068 9253
rect 3089 9251 3091 9259
rect 3116 9251 3118 9259
rect 3142 9245 3144 9253
rect 3147 9245 3149 9253
rect 3170 9251 3172 9259
rect 3980 9251 3982 9259
rect 3806 9238 3808 9246
rect 3822 9238 3824 9246
rect 3838 9238 3840 9246
rect 3861 9238 3863 9246
rect 3866 9238 3868 9246
rect 3892 9238 3894 9246
rect 3913 9238 3915 9246
rect 3933 9238 3935 9246
rect 3938 9238 3940 9246
rect 3956 9238 3958 9246
rect 4006 9245 4008 9253
rect 4011 9245 4013 9253
rect 4034 9251 4036 9259
rect 4061 9251 4063 9259
rect 4087 9245 4089 9253
rect 4092 9245 4094 9253
rect 4115 9251 4117 9259
rect 2495 9187 2497 9195
rect 2511 9187 2513 9195
rect 2516 9187 2518 9195
rect 2532 9187 2534 9195
rect 2548 9187 2550 9195
rect 2569 9187 2571 9195
rect 2574 9187 2576 9195
rect 2590 9187 2592 9195
rect 2606 9187 2608 9195
rect 2611 9187 2613 9195
rect 3440 9187 3442 9195
rect 3456 9187 3458 9195
rect 3461 9187 3463 9195
rect 3477 9187 3479 9195
rect 3493 9187 3495 9195
rect 3514 9187 3516 9195
rect 3519 9187 3521 9195
rect 3535 9187 3537 9195
rect 3551 9187 3553 9195
rect 3556 9187 3558 9195
rect 2861 9152 2863 9160
rect 2877 9152 2879 9160
rect 2893 9152 2895 9160
rect 2916 9152 2918 9160
rect 2921 9152 2923 9160
rect 2947 9152 2949 9160
rect 2968 9152 2970 9160
rect 2988 9152 2990 9160
rect 2993 9152 2995 9160
rect 3011 9152 3013 9160
rect 3061 9153 3063 9161
rect 3066 9153 3068 9161
rect 3142 9153 3144 9161
rect 3147 9153 3149 9161
rect 3806 9152 3808 9160
rect 3822 9152 3824 9160
rect 3838 9152 3840 9160
rect 3861 9152 3863 9160
rect 3866 9152 3868 9160
rect 3892 9152 3894 9160
rect 3913 9152 3915 9160
rect 3933 9152 3935 9160
rect 3938 9152 3940 9160
rect 3956 9152 3958 9160
rect 4006 9153 4008 9161
rect 4011 9153 4013 9161
rect 4087 9153 4089 9161
rect 4092 9153 4094 9161
rect 2861 9106 2863 9114
rect 2877 9106 2879 9114
rect 2893 9106 2895 9114
rect 2916 9106 2918 9114
rect 2921 9106 2923 9114
rect 2947 9106 2949 9114
rect 2968 9106 2970 9114
rect 2988 9106 2990 9114
rect 2993 9106 2995 9114
rect 3011 9106 3013 9114
rect 3061 9113 3063 9121
rect 3066 9113 3068 9121
rect 3089 9119 3091 9127
rect 3140 9119 3142 9127
rect 3166 9113 3168 9121
rect 3171 9113 3173 9121
rect 3194 9119 3196 9127
rect 3806 9106 3808 9114
rect 3822 9106 3824 9114
rect 3838 9106 3840 9114
rect 3861 9106 3863 9114
rect 3866 9106 3868 9114
rect 3892 9106 3894 9114
rect 3913 9106 3915 9114
rect 3933 9106 3935 9114
rect 3938 9106 3940 9114
rect 3956 9106 3958 9114
rect 4006 9113 4008 9121
rect 4011 9113 4013 9121
rect 4034 9119 4036 9127
rect 4085 9119 4087 9127
rect 3371 9090 3373 9098
rect 3397 9084 3399 9092
rect 3402 9084 3404 9092
rect 3425 9090 3427 9098
rect 3557 9065 3559 9095
rect 3610 9065 3612 9095
rect 4111 9113 4113 9121
rect 4116 9113 4118 9121
rect 4139 9119 4141 9127
rect 2861 9020 2863 9028
rect 2877 9020 2879 9028
rect 2893 9020 2895 9028
rect 2916 9020 2918 9028
rect 2921 9020 2923 9028
rect 2947 9020 2949 9028
rect 2968 9020 2970 9028
rect 2988 9020 2990 9028
rect 2993 9020 2995 9028
rect 3011 9020 3013 9028
rect 3061 9022 3063 9030
rect 3066 9022 3068 9030
rect 3166 9022 3168 9030
rect 3171 9022 3173 9030
rect 3806 9020 3808 9028
rect 3822 9020 3824 9028
rect 3838 9020 3840 9028
rect 3861 9020 3863 9028
rect 3866 9020 3868 9028
rect 3892 9020 3894 9028
rect 3913 9020 3915 9028
rect 3933 9020 3935 9028
rect 3938 9020 3940 9028
rect 3956 9020 3958 9028
rect 4006 9022 4008 9030
rect 4011 9022 4013 9030
rect 4111 9022 4113 9030
rect 4116 9022 4118 9030
rect 2861 8974 2863 8982
rect 2877 8974 2879 8982
rect 2893 8974 2895 8982
rect 2916 8974 2918 8982
rect 2921 8974 2923 8982
rect 2947 8974 2949 8982
rect 2968 8974 2970 8982
rect 2988 8974 2990 8982
rect 2993 8974 2995 8982
rect 3011 8974 3013 8982
rect 3061 8981 3063 8989
rect 3066 8981 3068 8989
rect 3089 8987 3091 8995
rect 3116 8987 3118 8995
rect 3142 8981 3144 8989
rect 3147 8981 3149 8989
rect 3170 8987 3172 8995
rect 3206 8987 3208 8995
rect 3232 8981 3234 8989
rect 3237 8981 3239 8989
rect 3260 8987 3262 8995
rect 3397 8988 3399 8996
rect 3402 8988 3404 8996
rect 3806 8974 3808 8982
rect 3822 8974 3824 8982
rect 3838 8974 3840 8982
rect 3861 8974 3863 8982
rect 3866 8974 3868 8982
rect 3892 8974 3894 8982
rect 3913 8974 3915 8982
rect 3933 8974 3935 8982
rect 3938 8974 3940 8982
rect 3956 8974 3958 8982
rect 4006 8981 4008 8989
rect 4011 8981 4013 8989
rect 4034 8987 4036 8995
rect 4061 8987 4063 8995
rect 3349 8960 3351 8968
rect 3371 8960 3373 8968
rect 3397 8954 3399 8962
rect 3402 8954 3404 8962
rect 3425 8960 3427 8968
rect 3463 8935 3465 8965
rect 3516 8935 3518 8965
rect 4087 8981 4089 8989
rect 4092 8981 4094 8989
rect 4115 8987 4117 8995
rect 4151 8987 4153 8995
rect 4177 8981 4179 8989
rect 4182 8981 4184 8989
rect 4205 8987 4207 8995
rect 2861 8888 2863 8896
rect 2877 8888 2879 8896
rect 2893 8888 2895 8896
rect 2916 8888 2918 8896
rect 2921 8888 2923 8896
rect 2947 8888 2949 8896
rect 2968 8888 2970 8896
rect 2988 8888 2990 8896
rect 2993 8888 2995 8896
rect 3011 8888 3013 8896
rect 3061 8887 3063 8895
rect 3066 8887 3068 8895
rect 3142 8887 3144 8895
rect 3147 8887 3149 8895
rect 3232 8887 3234 8895
rect 3237 8887 3239 8895
rect 3806 8888 3808 8896
rect 3822 8888 3824 8896
rect 3838 8888 3840 8896
rect 3861 8888 3863 8896
rect 3866 8888 3868 8896
rect 3892 8888 3894 8896
rect 3913 8888 3915 8896
rect 3933 8888 3935 8896
rect 3938 8888 3940 8896
rect 3956 8888 3958 8896
rect 4006 8887 4008 8895
rect 4011 8887 4013 8895
rect 4087 8887 4089 8895
rect 4092 8887 4094 8895
rect 4177 8887 4179 8895
rect 4182 8887 4184 8895
rect 2861 8842 2863 8850
rect 2877 8842 2879 8850
rect 2893 8842 2895 8850
rect 2916 8842 2918 8850
rect 2921 8842 2923 8850
rect 2947 8842 2949 8850
rect 2968 8842 2970 8850
rect 2988 8842 2990 8850
rect 2993 8842 2995 8850
rect 3011 8842 3013 8850
rect 3061 8849 3063 8857
rect 3066 8849 3068 8857
rect 3089 8855 3091 8863
rect 3397 8858 3399 8866
rect 3402 8858 3404 8866
rect 3806 8842 3808 8850
rect 3822 8842 3824 8850
rect 3838 8842 3840 8850
rect 3861 8842 3863 8850
rect 3866 8842 3868 8850
rect 3892 8842 3894 8850
rect 3913 8842 3915 8850
rect 3933 8842 3935 8850
rect 3938 8842 3940 8850
rect 3956 8842 3958 8850
rect 4006 8849 4008 8857
rect 4011 8849 4013 8857
rect 4034 8855 4036 8863
rect 2372 8787 2374 8795
rect 2377 8787 2379 8795
rect 2393 8787 2395 8795
rect 2409 8787 2411 8795
rect 2414 8787 2416 8795
rect 2435 8787 2437 8795
rect 2451 8787 2453 8795
rect 2467 8787 2469 8795
rect 2472 8787 2474 8795
rect 2488 8787 2490 8795
rect 2504 8787 2506 8795
rect 2509 8787 2511 8795
rect 2525 8787 2527 8795
rect 2541 8787 2543 8795
rect 2546 8787 2548 8795
rect 2567 8787 2569 8795
rect 2583 8787 2585 8795
rect 2599 8787 2601 8795
rect 2604 8787 2606 8795
rect 2620 8787 2622 8795
rect 2636 8787 2638 8795
rect 2641 8787 2643 8795
rect 2657 8787 2659 8795
rect 2673 8787 2675 8795
rect 2678 8787 2680 8795
rect 2699 8787 2701 8795
rect 2715 8787 2717 8795
rect 2731 8787 2733 8795
rect 2736 8787 2738 8795
rect 2752 8787 2754 8795
rect 3317 8787 3319 8795
rect 3322 8787 3324 8795
rect 3338 8787 3340 8795
rect 3354 8787 3356 8795
rect 3359 8787 3361 8795
rect 3380 8787 3382 8795
rect 3396 8787 3398 8795
rect 3412 8787 3414 8795
rect 3417 8787 3419 8795
rect 3433 8787 3435 8795
rect 3449 8787 3451 8795
rect 3454 8787 3456 8795
rect 3470 8787 3472 8795
rect 3486 8787 3488 8795
rect 3491 8787 3493 8795
rect 3512 8787 3514 8795
rect 3528 8787 3530 8795
rect 3544 8787 3546 8795
rect 3549 8787 3551 8795
rect 3565 8787 3567 8795
rect 3581 8787 3583 8795
rect 3586 8787 3588 8795
rect 3602 8787 3604 8795
rect 3618 8787 3620 8795
rect 3623 8787 3625 8795
rect 3644 8787 3646 8795
rect 3660 8787 3662 8795
rect 3676 8787 3678 8795
rect 3681 8787 3683 8795
rect 3697 8787 3699 8795
rect 2861 8756 2863 8764
rect 2877 8756 2879 8764
rect 2893 8756 2895 8764
rect 2916 8756 2918 8764
rect 2921 8756 2923 8764
rect 2947 8756 2949 8764
rect 2968 8756 2970 8764
rect 2988 8756 2990 8764
rect 2993 8756 2995 8764
rect 3011 8756 3013 8764
rect 3061 8751 3063 8759
rect 3066 8751 3068 8759
rect 3095 8756 3097 8764
rect 3113 8756 3115 8764
rect 3138 8756 3140 8764
rect 3154 8756 3156 8764
rect 3177 8756 3179 8764
rect 3182 8756 3184 8764
rect 3208 8756 3210 8764
rect 3229 8756 3231 8764
rect 3249 8756 3251 8764
rect 3254 8756 3256 8764
rect 3272 8756 3274 8764
rect 3806 8756 3808 8764
rect 3822 8756 3824 8764
rect 3838 8756 3840 8764
rect 3861 8756 3863 8764
rect 3866 8756 3868 8764
rect 3892 8756 3894 8764
rect 3913 8756 3915 8764
rect 3933 8756 3935 8764
rect 3938 8756 3940 8764
rect 3956 8756 3958 8764
rect 4006 8751 4008 8759
rect 4011 8751 4013 8759
rect 4040 8756 4042 8764
rect 4058 8756 4060 8764
rect 4083 8756 4085 8764
rect 4099 8756 4101 8764
rect 4122 8756 4124 8764
rect 4127 8756 4129 8764
rect 4153 8756 4155 8764
rect 4174 8756 4176 8764
rect 4194 8756 4196 8764
rect 4199 8756 4201 8764
rect 4217 8756 4219 8764
rect 3155 8675 3157 8683
rect 3160 8675 3162 8683
rect 3176 8675 3178 8683
rect 3192 8675 3194 8683
rect 3197 8675 3199 8683
rect 3218 8675 3220 8683
rect 3234 8675 3236 8683
rect 3250 8675 3252 8683
rect 3255 8675 3257 8683
rect 3271 8675 3273 8683
rect 4100 8675 4102 8683
rect 4105 8675 4107 8683
rect 4121 8675 4123 8683
rect 4137 8675 4139 8683
rect 4142 8675 4144 8683
rect 4163 8675 4165 8683
rect 4179 8675 4181 8683
rect 4195 8675 4197 8683
rect 4200 8675 4202 8683
rect 4216 8675 4218 8683
rect 2372 8645 2374 8653
rect 2377 8645 2379 8653
rect 2393 8645 2395 8653
rect 2409 8645 2411 8653
rect 2414 8645 2416 8653
rect 2435 8645 2437 8653
rect 2451 8645 2453 8653
rect 2467 8645 2469 8653
rect 2472 8645 2474 8653
rect 2488 8645 2490 8653
rect 2504 8645 2506 8653
rect 2509 8645 2511 8653
rect 2525 8645 2527 8653
rect 2541 8645 2543 8653
rect 2546 8645 2548 8653
rect 2567 8645 2569 8653
rect 2583 8645 2585 8653
rect 2599 8645 2601 8653
rect 2604 8645 2606 8653
rect 2620 8645 2622 8653
rect 2636 8645 2638 8653
rect 2641 8645 2643 8653
rect 2657 8645 2659 8653
rect 2673 8645 2675 8653
rect 2678 8645 2680 8653
rect 2699 8645 2701 8653
rect 2715 8645 2717 8653
rect 2731 8645 2733 8653
rect 2736 8645 2738 8653
rect 2752 8645 2754 8653
rect 3317 8645 3319 8653
rect 3322 8645 3324 8653
rect 3338 8645 3340 8653
rect 3354 8645 3356 8653
rect 3359 8645 3361 8653
rect 3380 8645 3382 8653
rect 3396 8645 3398 8653
rect 3412 8645 3414 8653
rect 3417 8645 3419 8653
rect 3433 8645 3435 8653
rect 3449 8645 3451 8653
rect 3454 8645 3456 8653
rect 3470 8645 3472 8653
rect 3486 8645 3488 8653
rect 3491 8645 3493 8653
rect 3512 8645 3514 8653
rect 3528 8645 3530 8653
rect 3544 8645 3546 8653
rect 3549 8645 3551 8653
rect 3565 8645 3567 8653
rect 3581 8645 3583 8653
rect 3586 8645 3588 8653
rect 3602 8645 3604 8653
rect 3618 8645 3620 8653
rect 3623 8645 3625 8653
rect 3644 8645 3646 8653
rect 3660 8645 3662 8653
rect 3676 8645 3678 8653
rect 3681 8645 3683 8653
rect 3697 8645 3699 8653
rect 3155 8589 3157 8597
rect 3160 8589 3162 8597
rect 3176 8589 3178 8597
rect 3192 8589 3194 8597
rect 3197 8589 3199 8597
rect 3218 8589 3220 8597
rect 3234 8589 3236 8597
rect 3250 8589 3252 8597
rect 3255 8589 3257 8597
rect 3271 8589 3273 8597
rect 4100 8589 4102 8597
rect 4105 8589 4107 8597
rect 4121 8589 4123 8597
rect 4137 8589 4139 8597
rect 4142 8589 4144 8597
rect 4163 8589 4165 8597
rect 4179 8589 4181 8597
rect 4195 8589 4197 8597
rect 4200 8589 4202 8597
rect 4216 8589 4218 8597
rect 2372 8559 2374 8567
rect 2377 8559 2379 8567
rect 2393 8559 2395 8567
rect 2409 8559 2411 8567
rect 2414 8559 2416 8567
rect 2435 8559 2437 8567
rect 2451 8559 2453 8567
rect 2467 8559 2469 8567
rect 2472 8559 2474 8567
rect 2488 8559 2490 8567
rect 2504 8559 2506 8567
rect 2509 8559 2511 8567
rect 2525 8559 2527 8567
rect 2541 8559 2543 8567
rect 2546 8559 2548 8567
rect 2567 8559 2569 8567
rect 2583 8559 2585 8567
rect 2599 8559 2601 8567
rect 2604 8559 2606 8567
rect 2620 8559 2622 8567
rect 2636 8559 2638 8567
rect 2641 8559 2643 8567
rect 2657 8559 2659 8567
rect 2673 8559 2675 8567
rect 2678 8559 2680 8567
rect 2699 8559 2701 8567
rect 2715 8559 2717 8567
rect 2731 8559 2733 8567
rect 2736 8559 2738 8567
rect 2752 8559 2754 8567
rect 3317 8559 3319 8567
rect 3322 8559 3324 8567
rect 3338 8559 3340 8567
rect 3354 8559 3356 8567
rect 3359 8559 3361 8567
rect 3380 8559 3382 8567
rect 3396 8559 3398 8567
rect 3412 8559 3414 8567
rect 3417 8559 3419 8567
rect 3433 8559 3435 8567
rect 3449 8559 3451 8567
rect 3454 8559 3456 8567
rect 3470 8559 3472 8567
rect 3486 8559 3488 8567
rect 3491 8559 3493 8567
rect 3512 8559 3514 8567
rect 3528 8559 3530 8567
rect 3544 8559 3546 8567
rect 3549 8559 3551 8567
rect 3565 8559 3567 8567
rect 3581 8559 3583 8567
rect 3586 8559 3588 8567
rect 3602 8559 3604 8567
rect 3618 8559 3620 8567
rect 3623 8559 3625 8567
rect 3644 8559 3646 8567
rect 3660 8559 3662 8567
rect 3676 8559 3678 8567
rect 3681 8559 3683 8567
rect 3697 8559 3699 8567
rect 2372 8419 2374 8427
rect 2377 8419 2379 8427
rect 2393 8419 2395 8427
rect 2409 8419 2411 8427
rect 2414 8419 2416 8427
rect 2435 8419 2437 8427
rect 2451 8419 2453 8427
rect 2467 8419 2469 8427
rect 2472 8419 2474 8427
rect 2488 8419 2490 8427
rect 2504 8419 2506 8427
rect 2509 8419 2511 8427
rect 2525 8419 2527 8427
rect 2541 8419 2543 8427
rect 2546 8419 2548 8427
rect 2567 8419 2569 8427
rect 2583 8419 2585 8427
rect 2599 8419 2601 8427
rect 2604 8419 2606 8427
rect 2620 8419 2622 8427
rect 2636 8419 2638 8427
rect 2641 8419 2643 8427
rect 2657 8419 2659 8427
rect 2673 8419 2675 8427
rect 2678 8419 2680 8427
rect 2699 8419 2701 8427
rect 2715 8419 2717 8427
rect 2731 8419 2733 8427
rect 2736 8419 2738 8427
rect 2752 8419 2754 8427
rect 3317 8419 3319 8427
rect 3322 8419 3324 8427
rect 3338 8419 3340 8427
rect 3354 8419 3356 8427
rect 3359 8419 3361 8427
rect 3380 8419 3382 8427
rect 3396 8419 3398 8427
rect 3412 8419 3414 8427
rect 3417 8419 3419 8427
rect 3433 8419 3435 8427
rect 3449 8419 3451 8427
rect 3454 8419 3456 8427
rect 3470 8419 3472 8427
rect 3486 8419 3488 8427
rect 3491 8419 3493 8427
rect 3512 8419 3514 8427
rect 3528 8419 3530 8427
rect 3544 8419 3546 8427
rect 3549 8419 3551 8427
rect 3565 8419 3567 8427
rect 3581 8419 3583 8427
rect 3586 8419 3588 8427
rect 3602 8419 3604 8427
rect 3618 8419 3620 8427
rect 3623 8419 3625 8427
rect 3644 8419 3646 8427
rect 3660 8419 3662 8427
rect 3676 8419 3678 8427
rect 3681 8419 3683 8427
rect 3697 8419 3699 8427
rect 2856 8340 2858 8348
rect 2861 8340 2863 8348
rect 2877 8340 2879 8348
rect 2893 8340 2895 8348
rect 2898 8340 2900 8348
rect 2919 8340 2921 8348
rect 2935 8340 2937 8348
rect 2951 8340 2953 8348
rect 2956 8340 2958 8348
rect 2972 8340 2974 8348
rect 2988 8340 2990 8348
rect 2993 8340 2995 8348
rect 3009 8340 3011 8348
rect 3025 8340 3027 8348
rect 3030 8340 3032 8348
rect 3051 8340 3053 8348
rect 3067 8340 3069 8348
rect 3083 8340 3085 8348
rect 3088 8340 3090 8348
rect 3104 8340 3106 8348
rect 3120 8340 3122 8348
rect 3125 8340 3127 8348
rect 3141 8340 3143 8348
rect 3157 8340 3159 8348
rect 3162 8340 3164 8348
rect 3183 8340 3185 8348
rect 3199 8340 3201 8348
rect 3215 8340 3217 8348
rect 3220 8340 3222 8348
rect 3236 8340 3238 8348
rect 3252 8340 3254 8348
rect 3257 8340 3259 8348
rect 3273 8340 3275 8348
rect 3289 8340 3291 8348
rect 3294 8340 3296 8348
rect 3315 8340 3317 8348
rect 3331 8340 3333 8348
rect 3347 8340 3349 8348
rect 3352 8340 3354 8348
rect 3368 8340 3370 8348
rect 3801 8340 3803 8348
rect 3806 8340 3808 8348
rect 3822 8340 3824 8348
rect 3838 8340 3840 8348
rect 3843 8340 3845 8348
rect 3864 8340 3866 8348
rect 3880 8340 3882 8348
rect 3896 8340 3898 8348
rect 3901 8340 3903 8348
rect 3917 8340 3919 8348
rect 3933 8340 3935 8348
rect 3938 8340 3940 8348
rect 3954 8340 3956 8348
rect 3970 8340 3972 8348
rect 3975 8340 3977 8348
rect 3996 8340 3998 8348
rect 4012 8340 4014 8348
rect 4028 8340 4030 8348
rect 4033 8340 4035 8348
rect 4049 8340 4051 8348
rect 4065 8340 4067 8348
rect 4070 8340 4072 8348
rect 4086 8340 4088 8348
rect 4102 8340 4104 8348
rect 4107 8340 4109 8348
rect 4128 8340 4130 8348
rect 4144 8340 4146 8348
rect 4160 8340 4162 8348
rect 4165 8340 4167 8348
rect 4181 8340 4183 8348
rect 4197 8340 4199 8348
rect 4202 8340 4204 8348
rect 4218 8340 4220 8348
rect 4234 8340 4236 8348
rect 4239 8340 4241 8348
rect 4260 8340 4262 8348
rect 4276 8340 4278 8348
rect 4292 8340 4294 8348
rect 4297 8340 4299 8348
rect 4313 8340 4315 8348
rect 2504 8307 2506 8315
rect 2509 8307 2511 8315
rect 2525 8307 2527 8315
rect 2541 8307 2543 8315
rect 2546 8307 2548 8315
rect 2567 8307 2569 8315
rect 2583 8307 2585 8315
rect 2599 8307 2601 8315
rect 2604 8307 2606 8315
rect 2620 8307 2622 8315
rect 3449 8307 3451 8315
rect 3454 8307 3456 8315
rect 3470 8307 3472 8315
rect 3486 8307 3488 8315
rect 3491 8307 3493 8315
rect 3512 8307 3514 8315
rect 3528 8307 3530 8315
rect 3544 8307 3546 8315
rect 3549 8307 3551 8315
rect 3565 8307 3567 8315
rect 3035 8269 3037 8277
rect 2861 8256 2863 8264
rect 2877 8256 2879 8264
rect 2893 8256 2895 8264
rect 2916 8256 2918 8264
rect 2921 8256 2923 8264
rect 2947 8256 2949 8264
rect 2968 8256 2970 8264
rect 2988 8256 2990 8264
rect 2993 8256 2995 8264
rect 3011 8256 3013 8264
rect 3061 8263 3063 8271
rect 3066 8263 3068 8271
rect 3089 8269 3091 8277
rect 3116 8269 3118 8277
rect 3142 8263 3144 8271
rect 3147 8263 3149 8271
rect 3170 8269 3172 8277
rect 3980 8269 3982 8277
rect 3806 8256 3808 8264
rect 3822 8256 3824 8264
rect 3838 8256 3840 8264
rect 3861 8256 3863 8264
rect 3866 8256 3868 8264
rect 3892 8256 3894 8264
rect 3913 8256 3915 8264
rect 3933 8256 3935 8264
rect 3938 8256 3940 8264
rect 3956 8256 3958 8264
rect 4006 8263 4008 8271
rect 4011 8263 4013 8271
rect 4034 8269 4036 8277
rect 4061 8269 4063 8277
rect 4087 8263 4089 8271
rect 4092 8263 4094 8271
rect 4115 8269 4117 8277
rect 2495 8205 2497 8213
rect 2511 8205 2513 8213
rect 2516 8205 2518 8213
rect 2532 8205 2534 8213
rect 2548 8205 2550 8213
rect 2569 8205 2571 8213
rect 2574 8205 2576 8213
rect 2590 8205 2592 8213
rect 2606 8205 2608 8213
rect 2611 8205 2613 8213
rect 3440 8205 3442 8213
rect 3456 8205 3458 8213
rect 3461 8205 3463 8213
rect 3477 8205 3479 8213
rect 3493 8205 3495 8213
rect 3514 8205 3516 8213
rect 3519 8205 3521 8213
rect 3535 8205 3537 8213
rect 3551 8205 3553 8213
rect 3556 8205 3558 8213
rect 2861 8170 2863 8178
rect 2877 8170 2879 8178
rect 2893 8170 2895 8178
rect 2916 8170 2918 8178
rect 2921 8170 2923 8178
rect 2947 8170 2949 8178
rect 2968 8170 2970 8178
rect 2988 8170 2990 8178
rect 2993 8170 2995 8178
rect 3011 8170 3013 8178
rect 3061 8171 3063 8179
rect 3066 8171 3068 8179
rect 3142 8171 3144 8179
rect 3147 8171 3149 8179
rect 3806 8170 3808 8178
rect 3822 8170 3824 8178
rect 3838 8170 3840 8178
rect 3861 8170 3863 8178
rect 3866 8170 3868 8178
rect 3892 8170 3894 8178
rect 3913 8170 3915 8178
rect 3933 8170 3935 8178
rect 3938 8170 3940 8178
rect 3956 8170 3958 8178
rect 4006 8171 4008 8179
rect 4011 8171 4013 8179
rect 4087 8171 4089 8179
rect 4092 8171 4094 8179
rect 2861 8124 2863 8132
rect 2877 8124 2879 8132
rect 2893 8124 2895 8132
rect 2916 8124 2918 8132
rect 2921 8124 2923 8132
rect 2947 8124 2949 8132
rect 2968 8124 2970 8132
rect 2988 8124 2990 8132
rect 2993 8124 2995 8132
rect 3011 8124 3013 8132
rect 3061 8131 3063 8139
rect 3066 8131 3068 8139
rect 3089 8137 3091 8145
rect 3140 8137 3142 8145
rect 3166 8131 3168 8139
rect 3171 8131 3173 8139
rect 3194 8137 3196 8145
rect 3806 8124 3808 8132
rect 3822 8124 3824 8132
rect 3838 8124 3840 8132
rect 3861 8124 3863 8132
rect 3866 8124 3868 8132
rect 3892 8124 3894 8132
rect 3913 8124 3915 8132
rect 3933 8124 3935 8132
rect 3938 8124 3940 8132
rect 3956 8124 3958 8132
rect 4006 8131 4008 8139
rect 4011 8131 4013 8139
rect 4034 8137 4036 8145
rect 4085 8137 4087 8145
rect 4111 8131 4113 8139
rect 4116 8131 4118 8139
rect 4139 8137 4141 8145
rect 2861 8038 2863 8046
rect 2877 8038 2879 8046
rect 2893 8038 2895 8046
rect 2916 8038 2918 8046
rect 2921 8038 2923 8046
rect 2947 8038 2949 8046
rect 2968 8038 2970 8046
rect 2988 8038 2990 8046
rect 2993 8038 2995 8046
rect 3011 8038 3013 8046
rect 3061 8040 3063 8048
rect 3066 8040 3068 8048
rect 3166 8040 3168 8048
rect 3171 8040 3173 8048
rect 3806 8038 3808 8046
rect 3822 8038 3824 8046
rect 3838 8038 3840 8046
rect 3861 8038 3863 8046
rect 3866 8038 3868 8046
rect 3892 8038 3894 8046
rect 3913 8038 3915 8046
rect 3933 8038 3935 8046
rect 3938 8038 3940 8046
rect 3956 8038 3958 8046
rect 4006 8040 4008 8048
rect 4011 8040 4013 8048
rect 4111 8040 4113 8048
rect 4116 8040 4118 8048
rect 2861 7992 2863 8000
rect 2877 7992 2879 8000
rect 2893 7992 2895 8000
rect 2916 7992 2918 8000
rect 2921 7992 2923 8000
rect 2947 7992 2949 8000
rect 2968 7992 2970 8000
rect 2988 7992 2990 8000
rect 2993 7992 2995 8000
rect 3011 7992 3013 8000
rect 3061 7999 3063 8007
rect 3066 7999 3068 8007
rect 3089 8005 3091 8013
rect 3116 8005 3118 8013
rect 3142 7999 3144 8007
rect 3147 7999 3149 8007
rect 3170 8005 3172 8013
rect 3206 8005 3208 8013
rect 3232 7999 3234 8007
rect 3237 7999 3239 8007
rect 3260 8005 3262 8013
rect 3806 7992 3808 8000
rect 3822 7992 3824 8000
rect 3838 7992 3840 8000
rect 3861 7992 3863 8000
rect 3866 7992 3868 8000
rect 3892 7992 3894 8000
rect 3913 7992 3915 8000
rect 3933 7992 3935 8000
rect 3938 7992 3940 8000
rect 3956 7992 3958 8000
rect 4006 7999 4008 8007
rect 4011 7999 4013 8007
rect 4034 8005 4036 8013
rect 4061 8005 4063 8013
rect 4087 7999 4089 8007
rect 4092 7999 4094 8007
rect 4115 8005 4117 8013
rect 4151 8005 4153 8013
rect 4177 7999 4179 8007
rect 4182 7999 4184 8007
rect 4205 8005 4207 8013
rect 2861 7906 2863 7914
rect 2877 7906 2879 7914
rect 2893 7906 2895 7914
rect 2916 7906 2918 7914
rect 2921 7906 2923 7914
rect 2947 7906 2949 7914
rect 2968 7906 2970 7914
rect 2988 7906 2990 7914
rect 2993 7906 2995 7914
rect 3011 7906 3013 7914
rect 3061 7905 3063 7913
rect 3066 7905 3068 7913
rect 3142 7905 3144 7913
rect 3147 7905 3149 7913
rect 3232 7905 3234 7913
rect 3237 7905 3239 7913
rect 3806 7906 3808 7914
rect 3822 7906 3824 7914
rect 3838 7906 3840 7914
rect 3861 7906 3863 7914
rect 3866 7906 3868 7914
rect 3892 7906 3894 7914
rect 3913 7906 3915 7914
rect 3933 7906 3935 7914
rect 3938 7906 3940 7914
rect 3956 7906 3958 7914
rect 4006 7905 4008 7913
rect 4011 7905 4013 7913
rect 4087 7905 4089 7913
rect 4092 7905 4094 7913
rect 4177 7905 4179 7913
rect 4182 7905 4184 7913
rect 2861 7860 2863 7868
rect 2877 7860 2879 7868
rect 2893 7860 2895 7868
rect 2916 7860 2918 7868
rect 2921 7860 2923 7868
rect 2947 7860 2949 7868
rect 2968 7860 2970 7868
rect 2988 7860 2990 7868
rect 2993 7860 2995 7868
rect 3011 7860 3013 7868
rect 3061 7867 3063 7875
rect 3066 7867 3068 7875
rect 3089 7873 3091 7881
rect 3806 7860 3808 7868
rect 3822 7860 3824 7868
rect 3838 7860 3840 7868
rect 3861 7860 3863 7868
rect 3866 7860 3868 7868
rect 3892 7860 3894 7868
rect 3913 7860 3915 7868
rect 3933 7860 3935 7868
rect 3938 7860 3940 7868
rect 3956 7860 3958 7868
rect 4006 7867 4008 7875
rect 4011 7867 4013 7875
rect 4034 7873 4036 7881
rect 2372 7805 2374 7813
rect 2377 7805 2379 7813
rect 2393 7805 2395 7813
rect 2409 7805 2411 7813
rect 2414 7805 2416 7813
rect 2435 7805 2437 7813
rect 2451 7805 2453 7813
rect 2467 7805 2469 7813
rect 2472 7805 2474 7813
rect 2488 7805 2490 7813
rect 2504 7805 2506 7813
rect 2509 7805 2511 7813
rect 2525 7805 2527 7813
rect 2541 7805 2543 7813
rect 2546 7805 2548 7813
rect 2567 7805 2569 7813
rect 2583 7805 2585 7813
rect 2599 7805 2601 7813
rect 2604 7805 2606 7813
rect 2620 7805 2622 7813
rect 2636 7805 2638 7813
rect 2641 7805 2643 7813
rect 2657 7805 2659 7813
rect 2673 7805 2675 7813
rect 2678 7805 2680 7813
rect 2699 7805 2701 7813
rect 2715 7805 2717 7813
rect 2731 7805 2733 7813
rect 2736 7805 2738 7813
rect 2752 7805 2754 7813
rect 3317 7805 3319 7813
rect 3322 7805 3324 7813
rect 3338 7805 3340 7813
rect 3354 7805 3356 7813
rect 3359 7805 3361 7813
rect 3380 7805 3382 7813
rect 3396 7805 3398 7813
rect 3412 7805 3414 7813
rect 3417 7805 3419 7813
rect 3433 7805 3435 7813
rect 3449 7805 3451 7813
rect 3454 7805 3456 7813
rect 3470 7805 3472 7813
rect 3486 7805 3488 7813
rect 3491 7805 3493 7813
rect 3512 7805 3514 7813
rect 3528 7805 3530 7813
rect 3544 7805 3546 7813
rect 3549 7805 3551 7813
rect 3565 7805 3567 7813
rect 3581 7805 3583 7813
rect 3586 7805 3588 7813
rect 3602 7805 3604 7813
rect 3618 7805 3620 7813
rect 3623 7805 3625 7813
rect 3644 7805 3646 7813
rect 3660 7805 3662 7813
rect 3676 7805 3678 7813
rect 3681 7805 3683 7813
rect 3697 7805 3699 7813
rect 2861 7774 2863 7782
rect 2877 7774 2879 7782
rect 2893 7774 2895 7782
rect 2916 7774 2918 7782
rect 2921 7774 2923 7782
rect 2947 7774 2949 7782
rect 2968 7774 2970 7782
rect 2988 7774 2990 7782
rect 2993 7774 2995 7782
rect 3011 7774 3013 7782
rect 3061 7769 3063 7777
rect 3066 7769 3068 7777
rect 3095 7774 3097 7782
rect 3113 7774 3115 7782
rect 3138 7774 3140 7782
rect 3154 7774 3156 7782
rect 3177 7774 3179 7782
rect 3182 7774 3184 7782
rect 3208 7774 3210 7782
rect 3229 7774 3231 7782
rect 3249 7774 3251 7782
rect 3254 7774 3256 7782
rect 3272 7774 3274 7782
rect 3806 7774 3808 7782
rect 3822 7774 3824 7782
rect 3838 7774 3840 7782
rect 3861 7774 3863 7782
rect 3866 7774 3868 7782
rect 3892 7774 3894 7782
rect 3913 7774 3915 7782
rect 3933 7774 3935 7782
rect 3938 7774 3940 7782
rect 3956 7774 3958 7782
rect 4006 7769 4008 7777
rect 4011 7769 4013 7777
rect 4040 7774 4042 7782
rect 4058 7774 4060 7782
rect 4083 7774 4085 7782
rect 4099 7774 4101 7782
rect 4122 7774 4124 7782
rect 4127 7774 4129 7782
rect 4153 7774 4155 7782
rect 4174 7774 4176 7782
rect 4194 7774 4196 7782
rect 4199 7774 4201 7782
rect 4217 7774 4219 7782
rect 3155 7693 3157 7701
rect 3160 7693 3162 7701
rect 3176 7693 3178 7701
rect 3192 7693 3194 7701
rect 3197 7693 3199 7701
rect 3218 7693 3220 7701
rect 3234 7693 3236 7701
rect 3250 7693 3252 7701
rect 3255 7693 3257 7701
rect 3271 7693 3273 7701
rect 4100 7693 4102 7701
rect 4105 7693 4107 7701
rect 4121 7693 4123 7701
rect 4137 7693 4139 7701
rect 4142 7693 4144 7701
rect 4163 7693 4165 7701
rect 4179 7693 4181 7701
rect 4195 7693 4197 7701
rect 4200 7693 4202 7701
rect 4216 7693 4218 7701
rect 2372 7663 2374 7671
rect 2377 7663 2379 7671
rect 2393 7663 2395 7671
rect 2409 7663 2411 7671
rect 2414 7663 2416 7671
rect 2435 7663 2437 7671
rect 2451 7663 2453 7671
rect 2467 7663 2469 7671
rect 2472 7663 2474 7671
rect 2488 7663 2490 7671
rect 2504 7663 2506 7671
rect 2509 7663 2511 7671
rect 2525 7663 2527 7671
rect 2541 7663 2543 7671
rect 2546 7663 2548 7671
rect 2567 7663 2569 7671
rect 2583 7663 2585 7671
rect 2599 7663 2601 7671
rect 2604 7663 2606 7671
rect 2620 7663 2622 7671
rect 2636 7663 2638 7671
rect 2641 7663 2643 7671
rect 2657 7663 2659 7671
rect 2673 7663 2675 7671
rect 2678 7663 2680 7671
rect 2699 7663 2701 7671
rect 2715 7663 2717 7671
rect 2731 7663 2733 7671
rect 2736 7663 2738 7671
rect 2752 7663 2754 7671
rect 3317 7663 3319 7671
rect 3322 7663 3324 7671
rect 3338 7663 3340 7671
rect 3354 7663 3356 7671
rect 3359 7663 3361 7671
rect 3380 7663 3382 7671
rect 3396 7663 3398 7671
rect 3412 7663 3414 7671
rect 3417 7663 3419 7671
rect 3433 7663 3435 7671
rect 3449 7663 3451 7671
rect 3454 7663 3456 7671
rect 3470 7663 3472 7671
rect 3486 7663 3488 7671
rect 3491 7663 3493 7671
rect 3512 7663 3514 7671
rect 3528 7663 3530 7671
rect 3544 7663 3546 7671
rect 3549 7663 3551 7671
rect 3565 7663 3567 7671
rect 3581 7663 3583 7671
rect 3586 7663 3588 7671
rect 3602 7663 3604 7671
rect 3618 7663 3620 7671
rect 3623 7663 3625 7671
rect 3644 7663 3646 7671
rect 3660 7663 3662 7671
rect 3676 7663 3678 7671
rect 3681 7663 3683 7671
rect 3697 7663 3699 7671
rect 3155 7607 3157 7615
rect 3160 7607 3162 7615
rect 3176 7607 3178 7615
rect 3192 7607 3194 7615
rect 3197 7607 3199 7615
rect 3218 7607 3220 7615
rect 3234 7607 3236 7615
rect 3250 7607 3252 7615
rect 3255 7607 3257 7615
rect 3271 7607 3273 7615
rect 4100 7607 4102 7615
rect 4105 7607 4107 7615
rect 4121 7607 4123 7615
rect 4137 7607 4139 7615
rect 4142 7607 4144 7615
rect 4163 7607 4165 7615
rect 4179 7607 4181 7615
rect 4195 7607 4197 7615
rect 4200 7607 4202 7615
rect 4216 7607 4218 7615
rect 2372 7577 2374 7585
rect 2377 7577 2379 7585
rect 2393 7577 2395 7585
rect 2409 7577 2411 7585
rect 2414 7577 2416 7585
rect 2435 7577 2437 7585
rect 2451 7577 2453 7585
rect 2467 7577 2469 7585
rect 2472 7577 2474 7585
rect 2488 7577 2490 7585
rect 2504 7577 2506 7585
rect 2509 7577 2511 7585
rect 2525 7577 2527 7585
rect 2541 7577 2543 7585
rect 2546 7577 2548 7585
rect 2567 7577 2569 7585
rect 2583 7577 2585 7585
rect 2599 7577 2601 7585
rect 2604 7577 2606 7585
rect 2620 7577 2622 7585
rect 2636 7577 2638 7585
rect 2641 7577 2643 7585
rect 2657 7577 2659 7585
rect 2673 7577 2675 7585
rect 2678 7577 2680 7585
rect 2699 7577 2701 7585
rect 2715 7577 2717 7585
rect 2731 7577 2733 7585
rect 2736 7577 2738 7585
rect 2752 7577 2754 7585
rect 3317 7577 3319 7585
rect 3322 7577 3324 7585
rect 3338 7577 3340 7585
rect 3354 7577 3356 7585
rect 3359 7577 3361 7585
rect 3380 7577 3382 7585
rect 3396 7577 3398 7585
rect 3412 7577 3414 7585
rect 3417 7577 3419 7585
rect 3433 7577 3435 7585
rect 3449 7577 3451 7585
rect 3454 7577 3456 7585
rect 3470 7577 3472 7585
rect 3486 7577 3488 7585
rect 3491 7577 3493 7585
rect 3512 7577 3514 7585
rect 3528 7577 3530 7585
rect 3544 7577 3546 7585
rect 3549 7577 3551 7585
rect 3565 7577 3567 7585
rect 3581 7577 3583 7585
rect 3586 7577 3588 7585
rect 3602 7577 3604 7585
rect 3618 7577 3620 7585
rect 3623 7577 3625 7585
rect 3644 7577 3646 7585
rect 3660 7577 3662 7585
rect 3676 7577 3678 7585
rect 3681 7577 3683 7585
rect 3697 7577 3699 7585
rect 2372 7437 2374 7445
rect 2377 7437 2379 7445
rect 2393 7437 2395 7445
rect 2409 7437 2411 7445
rect 2414 7437 2416 7445
rect 2435 7437 2437 7445
rect 2451 7437 2453 7445
rect 2467 7437 2469 7445
rect 2472 7437 2474 7445
rect 2488 7437 2490 7445
rect 2504 7437 2506 7445
rect 2509 7437 2511 7445
rect 2525 7437 2527 7445
rect 2541 7437 2543 7445
rect 2546 7437 2548 7445
rect 2567 7437 2569 7445
rect 2583 7437 2585 7445
rect 2599 7437 2601 7445
rect 2604 7437 2606 7445
rect 2620 7437 2622 7445
rect 2636 7437 2638 7445
rect 2641 7437 2643 7445
rect 2657 7437 2659 7445
rect 2673 7437 2675 7445
rect 2678 7437 2680 7445
rect 2699 7437 2701 7445
rect 2715 7437 2717 7445
rect 2731 7437 2733 7445
rect 2736 7437 2738 7445
rect 2752 7437 2754 7445
rect 3317 7437 3319 7445
rect 3322 7437 3324 7445
rect 3338 7437 3340 7445
rect 3354 7437 3356 7445
rect 3359 7437 3361 7445
rect 3380 7437 3382 7445
rect 3396 7437 3398 7445
rect 3412 7437 3414 7445
rect 3417 7437 3419 7445
rect 3433 7437 3435 7445
rect 3449 7437 3451 7445
rect 3454 7437 3456 7445
rect 3470 7437 3472 7445
rect 3486 7437 3488 7445
rect 3491 7437 3493 7445
rect 3512 7437 3514 7445
rect 3528 7437 3530 7445
rect 3544 7437 3546 7445
rect 3549 7437 3551 7445
rect 3565 7437 3567 7445
rect 3581 7437 3583 7445
rect 3586 7437 3588 7445
rect 3602 7437 3604 7445
rect 3618 7437 3620 7445
rect 3623 7437 3625 7445
rect 3644 7437 3646 7445
rect 3660 7437 3662 7445
rect 3676 7437 3678 7445
rect 3681 7437 3683 7445
rect 3697 7437 3699 7445
rect 4579 7889 4581 7945
rect 4587 7889 4589 7945
rect 4595 7889 4597 7945
rect 4603 7889 4605 7945
rect 4611 7889 4613 7945
rect 4619 7889 4621 7945
rect 4634 7857 4636 7945
rect 4642 7857 4644 7945
rect 4650 7857 4652 7945
rect 4658 7857 4660 7945
rect 4677 7857 4679 7945
rect 4685 7857 4687 7945
rect 4693 7857 4695 7945
rect 4701 7857 4703 7945
rect 4718 7857 4720 7945
rect 4726 7857 4728 7945
rect 4734 7857 4736 7945
rect 4742 7857 4744 7945
<< ndiffusion >>
rect 1397 9949 1402 9953
rect 1406 9949 1412 9953
rect 1416 9949 1422 9953
rect 1426 9949 1432 9953
rect 1436 9949 1441 9953
rect 1397 9948 1441 9949
rect 1401 9944 1407 9948
rect 1411 9944 1417 9948
rect 1421 9944 1427 9948
rect 1431 9944 1437 9948
rect 1397 9943 1441 9944
rect 1397 9939 1402 9943
rect 1406 9939 1412 9943
rect 1416 9939 1422 9943
rect 1426 9939 1432 9943
rect 1436 9939 1441 9943
rect 1397 9938 1441 9939
rect 1401 9934 1407 9938
rect 1411 9934 1417 9938
rect 1421 9934 1427 9938
rect 1431 9934 1437 9938
rect 1397 9933 1441 9934
rect 1397 9929 1402 9933
rect 1406 9929 1412 9933
rect 1416 9929 1422 9933
rect 1426 9929 1432 9933
rect 1436 9929 1441 9933
rect 1397 9928 1441 9929
rect 1401 9924 1407 9928
rect 1411 9924 1417 9928
rect 1421 9924 1427 9928
rect 1431 9924 1437 9928
rect 1397 9923 1441 9924
rect 1397 9919 1402 9923
rect 1406 9919 1412 9923
rect 1416 9919 1422 9923
rect 1426 9919 1432 9923
rect 1436 9919 1441 9923
rect 1397 9918 1441 9919
rect 1401 9914 1407 9918
rect 1411 9914 1417 9918
rect 1421 9914 1427 9918
rect 1431 9914 1437 9918
rect 1397 9913 1441 9914
rect 1397 9909 1402 9913
rect 1406 9909 1412 9913
rect 1416 9909 1422 9913
rect 1426 9909 1432 9913
rect 1436 9909 1441 9913
rect 1397 9908 1441 9909
rect 1401 9904 1407 9908
rect 1411 9904 1417 9908
rect 1421 9904 1427 9908
rect 1431 9904 1437 9908
rect 1397 9903 1441 9904
rect 1397 9899 1402 9903
rect 1406 9899 1412 9903
rect 1416 9899 1422 9903
rect 1426 9899 1432 9903
rect 1436 9899 1441 9903
rect 1397 9898 1441 9899
rect 1401 9894 1407 9898
rect 1411 9894 1417 9898
rect 1421 9894 1427 9898
rect 1431 9894 1437 9898
rect 1397 9893 1441 9894
rect 1397 9889 1402 9893
rect 1406 9889 1412 9893
rect 1416 9889 1422 9893
rect 1426 9889 1432 9893
rect 1436 9889 1441 9893
rect 1397 9888 1441 9889
rect 1401 9884 1407 9888
rect 1411 9884 1417 9888
rect 1421 9884 1427 9888
rect 1431 9884 1437 9888
rect 1397 9883 1441 9884
rect 1397 9879 1402 9883
rect 1406 9879 1412 9883
rect 1416 9879 1422 9883
rect 1426 9879 1432 9883
rect 1436 9879 1441 9883
rect 1397 9878 1441 9879
rect 1401 9874 1407 9878
rect 1411 9874 1417 9878
rect 1421 9874 1427 9878
rect 1431 9874 1437 9878
rect 1397 9873 1441 9874
rect 1397 9869 1402 9873
rect 1406 9869 1412 9873
rect 1416 9869 1422 9873
rect 1426 9869 1432 9873
rect 1436 9869 1441 9873
rect 1397 9868 1441 9869
rect 1401 9864 1407 9868
rect 1411 9864 1417 9868
rect 1421 9864 1427 9868
rect 1431 9864 1437 9868
rect 1706 9949 1711 9953
rect 1715 9949 1721 9953
rect 1725 9949 1731 9953
rect 1735 9949 1741 9953
rect 1745 9949 1750 9953
rect 1706 9948 1750 9949
rect 1710 9944 1716 9948
rect 1720 9944 1726 9948
rect 1730 9944 1736 9948
rect 1740 9944 1746 9948
rect 1706 9943 1750 9944
rect 1706 9939 1711 9943
rect 1715 9939 1721 9943
rect 1725 9939 1731 9943
rect 1735 9939 1741 9943
rect 1745 9939 1750 9943
rect 1706 9938 1750 9939
rect 1710 9934 1716 9938
rect 1720 9934 1726 9938
rect 1730 9934 1736 9938
rect 1740 9934 1746 9938
rect 1706 9933 1750 9934
rect 1706 9929 1711 9933
rect 1715 9929 1721 9933
rect 1725 9929 1731 9933
rect 1735 9929 1741 9933
rect 1745 9929 1750 9933
rect 1706 9928 1750 9929
rect 1710 9924 1716 9928
rect 1720 9924 1726 9928
rect 1730 9924 1736 9928
rect 1740 9924 1746 9928
rect 1706 9923 1750 9924
rect 1706 9919 1711 9923
rect 1715 9919 1721 9923
rect 1725 9919 1731 9923
rect 1735 9919 1741 9923
rect 1745 9919 1750 9923
rect 1706 9918 1750 9919
rect 1710 9914 1716 9918
rect 1720 9914 1726 9918
rect 1730 9914 1736 9918
rect 1740 9914 1746 9918
rect 1706 9913 1750 9914
rect 1706 9909 1711 9913
rect 1715 9909 1721 9913
rect 1725 9909 1731 9913
rect 1735 9909 1741 9913
rect 1745 9909 1750 9913
rect 1706 9908 1750 9909
rect 1710 9904 1716 9908
rect 1720 9904 1726 9908
rect 1730 9904 1736 9908
rect 1740 9904 1746 9908
rect 1706 9903 1750 9904
rect 1706 9899 1711 9903
rect 1715 9899 1721 9903
rect 1725 9899 1731 9903
rect 1735 9899 1741 9903
rect 1745 9899 1750 9903
rect 1706 9898 1750 9899
rect 1710 9894 1716 9898
rect 1720 9894 1726 9898
rect 1730 9894 1736 9898
rect 1740 9894 1746 9898
rect 1706 9893 1750 9894
rect 1706 9889 1711 9893
rect 1715 9889 1721 9893
rect 1725 9889 1731 9893
rect 1735 9889 1741 9893
rect 1745 9889 1750 9893
rect 1706 9888 1750 9889
rect 1710 9884 1716 9888
rect 1720 9884 1726 9888
rect 1730 9884 1736 9888
rect 1740 9884 1746 9888
rect 1706 9883 1750 9884
rect 1706 9879 1711 9883
rect 1715 9879 1721 9883
rect 1725 9879 1731 9883
rect 1735 9879 1741 9883
rect 1745 9879 1750 9883
rect 1706 9878 1750 9879
rect 1710 9874 1716 9878
rect 1720 9874 1726 9878
rect 1730 9874 1736 9878
rect 1740 9874 1746 9878
rect 1706 9873 1750 9874
rect 1706 9869 1711 9873
rect 1715 9869 1721 9873
rect 1725 9869 1731 9873
rect 1735 9869 1741 9873
rect 1745 9869 1750 9873
rect 1706 9868 1750 9869
rect 1710 9864 1716 9868
rect 1720 9864 1726 9868
rect 1730 9864 1736 9868
rect 1740 9864 1746 9868
rect 2015 9949 2020 9953
rect 2024 9949 2030 9953
rect 2034 9949 2040 9953
rect 2044 9949 2050 9953
rect 2054 9949 2059 9953
rect 2015 9948 2059 9949
rect 2019 9944 2025 9948
rect 2029 9944 2035 9948
rect 2039 9944 2045 9948
rect 2049 9944 2055 9948
rect 2015 9943 2059 9944
rect 2015 9939 2020 9943
rect 2024 9939 2030 9943
rect 2034 9939 2040 9943
rect 2044 9939 2050 9943
rect 2054 9939 2059 9943
rect 2015 9938 2059 9939
rect 2019 9934 2025 9938
rect 2029 9934 2035 9938
rect 2039 9934 2045 9938
rect 2049 9934 2055 9938
rect 2015 9933 2059 9934
rect 2015 9929 2020 9933
rect 2024 9929 2030 9933
rect 2034 9929 2040 9933
rect 2044 9929 2050 9933
rect 2054 9929 2059 9933
rect 2015 9928 2059 9929
rect 2019 9924 2025 9928
rect 2029 9924 2035 9928
rect 2039 9924 2045 9928
rect 2049 9924 2055 9928
rect 2015 9923 2059 9924
rect 2015 9919 2020 9923
rect 2024 9919 2030 9923
rect 2034 9919 2040 9923
rect 2044 9919 2050 9923
rect 2054 9919 2059 9923
rect 2015 9918 2059 9919
rect 2019 9914 2025 9918
rect 2029 9914 2035 9918
rect 2039 9914 2045 9918
rect 2049 9914 2055 9918
rect 2015 9913 2059 9914
rect 2015 9909 2020 9913
rect 2024 9909 2030 9913
rect 2034 9909 2040 9913
rect 2044 9909 2050 9913
rect 2054 9909 2059 9913
rect 2015 9908 2059 9909
rect 2019 9904 2025 9908
rect 2029 9904 2035 9908
rect 2039 9904 2045 9908
rect 2049 9904 2055 9908
rect 2015 9903 2059 9904
rect 2015 9899 2020 9903
rect 2024 9899 2030 9903
rect 2034 9899 2040 9903
rect 2044 9899 2050 9903
rect 2054 9899 2059 9903
rect 2015 9898 2059 9899
rect 2019 9894 2025 9898
rect 2029 9894 2035 9898
rect 2039 9894 2045 9898
rect 2049 9894 2055 9898
rect 2015 9893 2059 9894
rect 2015 9889 2020 9893
rect 2024 9889 2030 9893
rect 2034 9889 2040 9893
rect 2044 9889 2050 9893
rect 2054 9889 2059 9893
rect 2015 9888 2059 9889
rect 2019 9884 2025 9888
rect 2029 9884 2035 9888
rect 2039 9884 2045 9888
rect 2049 9884 2055 9888
rect 2015 9883 2059 9884
rect 2015 9879 2020 9883
rect 2024 9879 2030 9883
rect 2034 9879 2040 9883
rect 2044 9879 2050 9883
rect 2054 9879 2059 9883
rect 2015 9878 2059 9879
rect 2019 9874 2025 9878
rect 2029 9874 2035 9878
rect 2039 9874 2045 9878
rect 2049 9874 2055 9878
rect 2015 9873 2059 9874
rect 2015 9869 2020 9873
rect 2024 9869 2030 9873
rect 2034 9869 2040 9873
rect 2044 9869 2050 9873
rect 2054 9869 2059 9873
rect 2015 9868 2059 9869
rect 2019 9864 2025 9868
rect 2029 9864 2035 9868
rect 2039 9864 2045 9868
rect 2049 9864 2055 9868
rect 2324 9949 2329 9953
rect 2333 9949 2339 9953
rect 2343 9949 2349 9953
rect 2353 9949 2359 9953
rect 2363 9949 2368 9953
rect 2324 9948 2368 9949
rect 2328 9944 2334 9948
rect 2338 9944 2344 9948
rect 2348 9944 2354 9948
rect 2358 9944 2364 9948
rect 2324 9943 2368 9944
rect 2324 9939 2329 9943
rect 2333 9939 2339 9943
rect 2343 9939 2349 9943
rect 2353 9939 2359 9943
rect 2363 9939 2368 9943
rect 2324 9938 2368 9939
rect 2328 9934 2334 9938
rect 2338 9934 2344 9938
rect 2348 9934 2354 9938
rect 2358 9934 2364 9938
rect 2324 9933 2368 9934
rect 2324 9929 2329 9933
rect 2333 9929 2339 9933
rect 2343 9929 2349 9933
rect 2353 9929 2359 9933
rect 2363 9929 2368 9933
rect 2324 9928 2368 9929
rect 2328 9924 2334 9928
rect 2338 9924 2344 9928
rect 2348 9924 2354 9928
rect 2358 9924 2364 9928
rect 2324 9923 2368 9924
rect 2324 9919 2329 9923
rect 2333 9919 2339 9923
rect 2343 9919 2349 9923
rect 2353 9919 2359 9923
rect 2363 9919 2368 9923
rect 2324 9918 2368 9919
rect 2328 9914 2334 9918
rect 2338 9914 2344 9918
rect 2348 9914 2354 9918
rect 2358 9914 2364 9918
rect 2324 9913 2368 9914
rect 2324 9909 2329 9913
rect 2333 9909 2339 9913
rect 2343 9909 2349 9913
rect 2353 9909 2359 9913
rect 2363 9909 2368 9913
rect 2324 9908 2368 9909
rect 2328 9904 2334 9908
rect 2338 9904 2344 9908
rect 2348 9904 2354 9908
rect 2358 9904 2364 9908
rect 2324 9903 2368 9904
rect 2324 9899 2329 9903
rect 2333 9899 2339 9903
rect 2343 9899 2349 9903
rect 2353 9899 2359 9903
rect 2363 9899 2368 9903
rect 2324 9898 2368 9899
rect 2328 9894 2334 9898
rect 2338 9894 2344 9898
rect 2348 9894 2354 9898
rect 2358 9894 2364 9898
rect 2324 9893 2368 9894
rect 2324 9889 2329 9893
rect 2333 9889 2339 9893
rect 2343 9889 2349 9893
rect 2353 9889 2359 9893
rect 2363 9889 2368 9893
rect 2324 9888 2368 9889
rect 2328 9884 2334 9888
rect 2338 9884 2344 9888
rect 2348 9884 2354 9888
rect 2358 9884 2364 9888
rect 2324 9883 2368 9884
rect 2324 9879 2329 9883
rect 2333 9879 2339 9883
rect 2343 9879 2349 9883
rect 2353 9879 2359 9883
rect 2363 9879 2368 9883
rect 2324 9878 2368 9879
rect 2328 9874 2334 9878
rect 2338 9874 2344 9878
rect 2348 9874 2354 9878
rect 2358 9874 2364 9878
rect 2324 9873 2368 9874
rect 2324 9869 2329 9873
rect 2333 9869 2339 9873
rect 2343 9869 2349 9873
rect 2353 9869 2359 9873
rect 2363 9869 2368 9873
rect 2324 9868 2368 9869
rect 2328 9864 2334 9868
rect 2338 9864 2344 9868
rect 2348 9864 2354 9868
rect 2358 9864 2364 9868
rect 2633 9949 2638 9953
rect 2642 9949 2648 9953
rect 2652 9949 2658 9953
rect 2662 9949 2668 9953
rect 2672 9949 2677 9953
rect 2633 9948 2677 9949
rect 2637 9944 2643 9948
rect 2647 9944 2653 9948
rect 2657 9944 2663 9948
rect 2667 9944 2673 9948
rect 2633 9943 2677 9944
rect 2633 9939 2638 9943
rect 2642 9939 2648 9943
rect 2652 9939 2658 9943
rect 2662 9939 2668 9943
rect 2672 9939 2677 9943
rect 2633 9938 2677 9939
rect 2637 9934 2643 9938
rect 2647 9934 2653 9938
rect 2657 9934 2663 9938
rect 2667 9934 2673 9938
rect 2633 9933 2677 9934
rect 2633 9929 2638 9933
rect 2642 9929 2648 9933
rect 2652 9929 2658 9933
rect 2662 9929 2668 9933
rect 2672 9929 2677 9933
rect 2633 9928 2677 9929
rect 2637 9924 2643 9928
rect 2647 9924 2653 9928
rect 2657 9924 2663 9928
rect 2667 9924 2673 9928
rect 2633 9923 2677 9924
rect 2633 9919 2638 9923
rect 2642 9919 2648 9923
rect 2652 9919 2658 9923
rect 2662 9919 2668 9923
rect 2672 9919 2677 9923
rect 2633 9918 2677 9919
rect 2637 9914 2643 9918
rect 2647 9914 2653 9918
rect 2657 9914 2663 9918
rect 2667 9914 2673 9918
rect 2633 9913 2677 9914
rect 2633 9909 2638 9913
rect 2642 9909 2648 9913
rect 2652 9909 2658 9913
rect 2662 9909 2668 9913
rect 2672 9909 2677 9913
rect 2633 9908 2677 9909
rect 2637 9904 2643 9908
rect 2647 9904 2653 9908
rect 2657 9904 2663 9908
rect 2667 9904 2673 9908
rect 2633 9903 2677 9904
rect 2633 9899 2638 9903
rect 2642 9899 2648 9903
rect 2652 9899 2658 9903
rect 2662 9899 2668 9903
rect 2672 9899 2677 9903
rect 2633 9898 2677 9899
rect 2637 9894 2643 9898
rect 2647 9894 2653 9898
rect 2657 9894 2663 9898
rect 2667 9894 2673 9898
rect 2633 9893 2677 9894
rect 2633 9889 2638 9893
rect 2642 9889 2648 9893
rect 2652 9889 2658 9893
rect 2662 9889 2668 9893
rect 2672 9889 2677 9893
rect 2633 9888 2677 9889
rect 2637 9884 2643 9888
rect 2647 9884 2653 9888
rect 2657 9884 2663 9888
rect 2667 9884 2673 9888
rect 2633 9883 2677 9884
rect 2633 9879 2638 9883
rect 2642 9879 2648 9883
rect 2652 9879 2658 9883
rect 2662 9879 2668 9883
rect 2672 9879 2677 9883
rect 2633 9878 2677 9879
rect 2637 9874 2643 9878
rect 2647 9874 2653 9878
rect 2657 9874 2663 9878
rect 2667 9874 2673 9878
rect 2633 9873 2677 9874
rect 2633 9869 2638 9873
rect 2642 9869 2648 9873
rect 2652 9869 2658 9873
rect 2662 9869 2668 9873
rect 2672 9869 2677 9873
rect 2633 9868 2677 9869
rect 2637 9864 2643 9868
rect 2647 9864 2653 9868
rect 2657 9864 2663 9868
rect 2667 9864 2673 9868
rect 2942 9949 2947 9953
rect 2951 9949 2957 9953
rect 2961 9949 2967 9953
rect 2971 9949 2977 9953
rect 2981 9949 2986 9953
rect 2942 9948 2986 9949
rect 2946 9944 2952 9948
rect 2956 9944 2962 9948
rect 2966 9944 2972 9948
rect 2976 9944 2982 9948
rect 2942 9943 2986 9944
rect 2942 9939 2947 9943
rect 2951 9939 2957 9943
rect 2961 9939 2967 9943
rect 2971 9939 2977 9943
rect 2981 9939 2986 9943
rect 2942 9938 2986 9939
rect 2946 9934 2952 9938
rect 2956 9934 2962 9938
rect 2966 9934 2972 9938
rect 2976 9934 2982 9938
rect 2942 9933 2986 9934
rect 2942 9929 2947 9933
rect 2951 9929 2957 9933
rect 2961 9929 2967 9933
rect 2971 9929 2977 9933
rect 2981 9929 2986 9933
rect 2942 9928 2986 9929
rect 2946 9924 2952 9928
rect 2956 9924 2962 9928
rect 2966 9924 2972 9928
rect 2976 9924 2982 9928
rect 2942 9923 2986 9924
rect 2942 9919 2947 9923
rect 2951 9919 2957 9923
rect 2961 9919 2967 9923
rect 2971 9919 2977 9923
rect 2981 9919 2986 9923
rect 2942 9918 2986 9919
rect 2946 9914 2952 9918
rect 2956 9914 2962 9918
rect 2966 9914 2972 9918
rect 2976 9914 2982 9918
rect 2942 9913 2986 9914
rect 2942 9909 2947 9913
rect 2951 9909 2957 9913
rect 2961 9909 2967 9913
rect 2971 9909 2977 9913
rect 2981 9909 2986 9913
rect 2942 9908 2986 9909
rect 2946 9904 2952 9908
rect 2956 9904 2962 9908
rect 2966 9904 2972 9908
rect 2976 9904 2982 9908
rect 2942 9903 2986 9904
rect 2942 9899 2947 9903
rect 2951 9899 2957 9903
rect 2961 9899 2967 9903
rect 2971 9899 2977 9903
rect 2981 9899 2986 9903
rect 2942 9898 2986 9899
rect 2946 9894 2952 9898
rect 2956 9894 2962 9898
rect 2966 9894 2972 9898
rect 2976 9894 2982 9898
rect 2942 9893 2986 9894
rect 2942 9889 2947 9893
rect 2951 9889 2957 9893
rect 2961 9889 2967 9893
rect 2971 9889 2977 9893
rect 2981 9889 2986 9893
rect 2942 9888 2986 9889
rect 2946 9884 2952 9888
rect 2956 9884 2962 9888
rect 2966 9884 2972 9888
rect 2976 9884 2982 9888
rect 2942 9883 2986 9884
rect 2942 9879 2947 9883
rect 2951 9879 2957 9883
rect 2961 9879 2967 9883
rect 2971 9879 2977 9883
rect 2981 9879 2986 9883
rect 2942 9878 2986 9879
rect 2946 9874 2952 9878
rect 2956 9874 2962 9878
rect 2966 9874 2972 9878
rect 2976 9874 2982 9878
rect 2942 9873 2986 9874
rect 2942 9869 2947 9873
rect 2951 9869 2957 9873
rect 2961 9869 2967 9873
rect 2971 9869 2977 9873
rect 2981 9869 2986 9873
rect 2942 9868 2986 9869
rect 2946 9864 2952 9868
rect 2956 9864 2962 9868
rect 2966 9864 2972 9868
rect 2976 9864 2982 9868
rect 3251 9949 3256 9953
rect 3260 9949 3266 9953
rect 3270 9949 3276 9953
rect 3280 9949 3286 9953
rect 3290 9949 3295 9953
rect 3251 9948 3295 9949
rect 3255 9944 3261 9948
rect 3265 9944 3271 9948
rect 3275 9944 3281 9948
rect 3285 9944 3291 9948
rect 3251 9943 3295 9944
rect 3251 9939 3256 9943
rect 3260 9939 3266 9943
rect 3270 9939 3276 9943
rect 3280 9939 3286 9943
rect 3290 9939 3295 9943
rect 3251 9938 3295 9939
rect 3255 9934 3261 9938
rect 3265 9934 3271 9938
rect 3275 9934 3281 9938
rect 3285 9934 3291 9938
rect 3251 9933 3295 9934
rect 3251 9929 3256 9933
rect 3260 9929 3266 9933
rect 3270 9929 3276 9933
rect 3280 9929 3286 9933
rect 3290 9929 3295 9933
rect 3251 9928 3295 9929
rect 3255 9924 3261 9928
rect 3265 9924 3271 9928
rect 3275 9924 3281 9928
rect 3285 9924 3291 9928
rect 3251 9923 3295 9924
rect 3251 9919 3256 9923
rect 3260 9919 3266 9923
rect 3270 9919 3276 9923
rect 3280 9919 3286 9923
rect 3290 9919 3295 9923
rect 3251 9918 3295 9919
rect 3255 9914 3261 9918
rect 3265 9914 3271 9918
rect 3275 9914 3281 9918
rect 3285 9914 3291 9918
rect 3251 9913 3295 9914
rect 3251 9909 3256 9913
rect 3260 9909 3266 9913
rect 3270 9909 3276 9913
rect 3280 9909 3286 9913
rect 3290 9909 3295 9913
rect 3251 9908 3295 9909
rect 3255 9904 3261 9908
rect 3265 9904 3271 9908
rect 3275 9904 3281 9908
rect 3285 9904 3291 9908
rect 3251 9903 3295 9904
rect 3251 9899 3256 9903
rect 3260 9899 3266 9903
rect 3270 9899 3276 9903
rect 3280 9899 3286 9903
rect 3290 9899 3295 9903
rect 3251 9898 3295 9899
rect 3255 9894 3261 9898
rect 3265 9894 3271 9898
rect 3275 9894 3281 9898
rect 3285 9894 3291 9898
rect 3251 9893 3295 9894
rect 3251 9889 3256 9893
rect 3260 9889 3266 9893
rect 3270 9889 3276 9893
rect 3280 9889 3286 9893
rect 3290 9889 3295 9893
rect 3251 9888 3295 9889
rect 3255 9884 3261 9888
rect 3265 9884 3271 9888
rect 3275 9884 3281 9888
rect 3285 9884 3291 9888
rect 3251 9883 3295 9884
rect 3251 9879 3256 9883
rect 3260 9879 3266 9883
rect 3270 9879 3276 9883
rect 3280 9879 3286 9883
rect 3290 9879 3295 9883
rect 3251 9878 3295 9879
rect 3255 9874 3261 9878
rect 3265 9874 3271 9878
rect 3275 9874 3281 9878
rect 3285 9874 3291 9878
rect 3251 9873 3295 9874
rect 3251 9869 3256 9873
rect 3260 9869 3266 9873
rect 3270 9869 3276 9873
rect 3280 9869 3286 9873
rect 3290 9869 3295 9873
rect 3251 9868 3295 9869
rect 3255 9864 3261 9868
rect 3265 9864 3271 9868
rect 3275 9864 3281 9868
rect 3285 9864 3291 9868
rect 3560 9949 3565 9953
rect 3569 9949 3575 9953
rect 3579 9949 3585 9953
rect 3589 9949 3595 9953
rect 3599 9949 3604 9953
rect 3560 9948 3604 9949
rect 3564 9944 3570 9948
rect 3574 9944 3580 9948
rect 3584 9944 3590 9948
rect 3594 9944 3600 9948
rect 3560 9943 3604 9944
rect 3560 9939 3565 9943
rect 3569 9939 3575 9943
rect 3579 9939 3585 9943
rect 3589 9939 3595 9943
rect 3599 9939 3604 9943
rect 3560 9938 3604 9939
rect 3564 9934 3570 9938
rect 3574 9934 3580 9938
rect 3584 9934 3590 9938
rect 3594 9934 3600 9938
rect 3560 9933 3604 9934
rect 3560 9929 3565 9933
rect 3569 9929 3575 9933
rect 3579 9929 3585 9933
rect 3589 9929 3595 9933
rect 3599 9929 3604 9933
rect 3560 9928 3604 9929
rect 3564 9924 3570 9928
rect 3574 9924 3580 9928
rect 3584 9924 3590 9928
rect 3594 9924 3600 9928
rect 3560 9923 3604 9924
rect 3560 9919 3565 9923
rect 3569 9919 3575 9923
rect 3579 9919 3585 9923
rect 3589 9919 3595 9923
rect 3599 9919 3604 9923
rect 3560 9918 3604 9919
rect 3564 9914 3570 9918
rect 3574 9914 3580 9918
rect 3584 9914 3590 9918
rect 3594 9914 3600 9918
rect 3560 9913 3604 9914
rect 3560 9909 3565 9913
rect 3569 9909 3575 9913
rect 3579 9909 3585 9913
rect 3589 9909 3595 9913
rect 3599 9909 3604 9913
rect 3560 9908 3604 9909
rect 3564 9904 3570 9908
rect 3574 9904 3580 9908
rect 3584 9904 3590 9908
rect 3594 9904 3600 9908
rect 3560 9903 3604 9904
rect 3560 9899 3565 9903
rect 3569 9899 3575 9903
rect 3579 9899 3585 9903
rect 3589 9899 3595 9903
rect 3599 9899 3604 9903
rect 3560 9898 3604 9899
rect 3564 9894 3570 9898
rect 3574 9894 3580 9898
rect 3584 9894 3590 9898
rect 3594 9894 3600 9898
rect 3560 9893 3604 9894
rect 3560 9889 3565 9893
rect 3569 9889 3575 9893
rect 3579 9889 3585 9893
rect 3589 9889 3595 9893
rect 3599 9889 3604 9893
rect 3560 9888 3604 9889
rect 3564 9884 3570 9888
rect 3574 9884 3580 9888
rect 3584 9884 3590 9888
rect 3594 9884 3600 9888
rect 3560 9883 3604 9884
rect 3560 9879 3565 9883
rect 3569 9879 3575 9883
rect 3579 9879 3585 9883
rect 3589 9879 3595 9883
rect 3599 9879 3604 9883
rect 3560 9878 3604 9879
rect 3564 9874 3570 9878
rect 3574 9874 3580 9878
rect 3584 9874 3590 9878
rect 3594 9874 3600 9878
rect 3560 9873 3604 9874
rect 3560 9869 3565 9873
rect 3569 9869 3575 9873
rect 3579 9869 3585 9873
rect 3589 9869 3595 9873
rect 3599 9869 3604 9873
rect 3560 9868 3604 9869
rect 3564 9864 3570 9868
rect 3574 9864 3580 9868
rect 3584 9864 3590 9868
rect 3594 9864 3600 9868
rect 3869 9949 3874 9953
rect 3878 9949 3884 9953
rect 3888 9949 3894 9953
rect 3898 9949 3904 9953
rect 3908 9949 3913 9953
rect 3869 9948 3913 9949
rect 3873 9944 3879 9948
rect 3883 9944 3889 9948
rect 3893 9944 3899 9948
rect 3903 9944 3909 9948
rect 3869 9943 3913 9944
rect 3869 9939 3874 9943
rect 3878 9939 3884 9943
rect 3888 9939 3894 9943
rect 3898 9939 3904 9943
rect 3908 9939 3913 9943
rect 3869 9938 3913 9939
rect 3873 9934 3879 9938
rect 3883 9934 3889 9938
rect 3893 9934 3899 9938
rect 3903 9934 3909 9938
rect 3869 9933 3913 9934
rect 3869 9929 3874 9933
rect 3878 9929 3884 9933
rect 3888 9929 3894 9933
rect 3898 9929 3904 9933
rect 3908 9929 3913 9933
rect 3869 9928 3913 9929
rect 3873 9924 3879 9928
rect 3883 9924 3889 9928
rect 3893 9924 3899 9928
rect 3903 9924 3909 9928
rect 3869 9923 3913 9924
rect 3869 9919 3874 9923
rect 3878 9919 3884 9923
rect 3888 9919 3894 9923
rect 3898 9919 3904 9923
rect 3908 9919 3913 9923
rect 3869 9918 3913 9919
rect 3873 9914 3879 9918
rect 3883 9914 3889 9918
rect 3893 9914 3899 9918
rect 3903 9914 3909 9918
rect 3869 9913 3913 9914
rect 3869 9909 3874 9913
rect 3878 9909 3884 9913
rect 3888 9909 3894 9913
rect 3898 9909 3904 9913
rect 3908 9909 3913 9913
rect 3869 9908 3913 9909
rect 3873 9904 3879 9908
rect 3883 9904 3889 9908
rect 3893 9904 3899 9908
rect 3903 9904 3909 9908
rect 3869 9903 3913 9904
rect 3869 9899 3874 9903
rect 3878 9899 3884 9903
rect 3888 9899 3894 9903
rect 3898 9899 3904 9903
rect 3908 9899 3913 9903
rect 3869 9898 3913 9899
rect 3873 9894 3879 9898
rect 3883 9894 3889 9898
rect 3893 9894 3899 9898
rect 3903 9894 3909 9898
rect 3869 9893 3913 9894
rect 3869 9889 3874 9893
rect 3878 9889 3884 9893
rect 3888 9889 3894 9893
rect 3898 9889 3904 9893
rect 3908 9889 3913 9893
rect 3869 9888 3913 9889
rect 3873 9884 3879 9888
rect 3883 9884 3889 9888
rect 3893 9884 3899 9888
rect 3903 9884 3909 9888
rect 3869 9883 3913 9884
rect 3869 9879 3874 9883
rect 3878 9879 3884 9883
rect 3888 9879 3894 9883
rect 3898 9879 3904 9883
rect 3908 9879 3913 9883
rect 3869 9878 3913 9879
rect 3873 9874 3879 9878
rect 3883 9874 3889 9878
rect 3893 9874 3899 9878
rect 3903 9874 3909 9878
rect 3869 9873 3913 9874
rect 3869 9869 3874 9873
rect 3878 9869 3884 9873
rect 3888 9869 3894 9873
rect 3898 9869 3904 9873
rect 3908 9869 3913 9873
rect 3869 9868 3913 9869
rect 3873 9864 3879 9868
rect 3883 9864 3889 9868
rect 3893 9864 3899 9868
rect 3903 9864 3909 9868
rect 1836 9827 1840 9831
rect 1829 9826 1869 9827
rect 2145 9827 2149 9831
rect 2138 9826 2178 9827
rect 2454 9827 2458 9831
rect 2447 9826 2487 9827
rect 2763 9827 2767 9831
rect 2756 9826 2796 9827
rect 3072 9827 3076 9831
rect 3065 9826 3105 9827
rect 3999 9827 4003 9831
rect 3992 9826 4032 9827
rect 1829 9823 1869 9824
rect 1829 9818 1869 9819
rect 2138 9823 2178 9824
rect 2138 9818 2178 9819
rect 2447 9823 2487 9824
rect 2447 9818 2487 9819
rect 2756 9823 2796 9824
rect 2756 9818 2796 9819
rect 3065 9823 3105 9824
rect 3065 9818 3105 9819
rect 3992 9823 4032 9824
rect 3992 9818 4032 9819
rect 1829 9815 1869 9816
rect 1836 9811 1840 9815
rect 1829 9810 1869 9811
rect 2138 9815 2178 9816
rect 1829 9807 1869 9808
rect 1829 9802 1869 9803
rect 1829 9799 1869 9800
rect 1836 9795 1840 9799
rect 1829 9794 1869 9795
rect 1829 9791 1869 9792
rect 1829 9786 1869 9787
rect 2145 9811 2149 9815
rect 2138 9810 2178 9811
rect 2447 9815 2487 9816
rect 2138 9807 2178 9808
rect 2138 9802 2178 9803
rect 2138 9799 2178 9800
rect 2145 9795 2149 9799
rect 2138 9794 2178 9795
rect 2138 9791 2178 9792
rect 2138 9786 2178 9787
rect 2454 9811 2458 9815
rect 2447 9810 2487 9811
rect 2756 9815 2796 9816
rect 2447 9807 2487 9808
rect 2447 9802 2487 9803
rect 2447 9799 2487 9800
rect 2454 9795 2458 9799
rect 2447 9794 2487 9795
rect 2447 9791 2487 9792
rect 2447 9786 2487 9787
rect 2763 9811 2767 9815
rect 2756 9810 2796 9811
rect 3065 9815 3105 9816
rect 2756 9807 2796 9808
rect 2756 9802 2796 9803
rect 2756 9799 2796 9800
rect 2763 9795 2767 9799
rect 2756 9794 2796 9795
rect 2756 9791 2796 9792
rect 2756 9786 2796 9787
rect 3072 9811 3076 9815
rect 3065 9810 3105 9811
rect 3992 9815 4032 9816
rect 3065 9807 3105 9808
rect 3065 9802 3105 9803
rect 3065 9799 3105 9800
rect 3072 9795 3076 9799
rect 3065 9794 3105 9795
rect 3065 9791 3105 9792
rect 3065 9786 3105 9787
rect 3999 9811 4003 9815
rect 3992 9810 4032 9811
rect 3992 9807 4032 9808
rect 3992 9802 4032 9803
rect 3992 9799 4032 9800
rect 3999 9795 4003 9799
rect 3992 9794 4032 9795
rect 3992 9791 4032 9792
rect 3992 9786 4032 9787
rect 1829 9783 1869 9784
rect 1836 9779 1840 9783
rect 2138 9783 2178 9784
rect 2145 9779 2149 9783
rect 2447 9783 2487 9784
rect 2454 9779 2458 9783
rect 2756 9783 2796 9784
rect 2763 9779 2767 9783
rect 3065 9783 3105 9784
rect 3072 9779 3076 9783
rect 3992 9783 4032 9784
rect 3999 9779 4003 9783
rect 2855 9299 2856 9303
rect 2858 9299 2861 9303
rect 2863 9299 2864 9303
rect 2876 9299 2877 9303
rect 2879 9299 2880 9303
rect 2892 9299 2893 9303
rect 2895 9299 2898 9303
rect 2900 9299 2901 9303
rect 2918 9299 2919 9303
rect 2921 9299 2922 9303
rect 2934 9299 2935 9303
rect 2937 9299 2938 9303
rect 2950 9299 2951 9303
rect 2953 9299 2956 9303
rect 2958 9299 2959 9303
rect 2971 9299 2972 9303
rect 2974 9299 2975 9303
rect 2987 9299 2988 9303
rect 2990 9299 2993 9303
rect 2995 9299 2996 9303
rect 3008 9299 3009 9303
rect 3011 9299 3012 9303
rect 3024 9299 3025 9303
rect 3027 9299 3030 9303
rect 3032 9299 3033 9303
rect 3050 9299 3051 9303
rect 3053 9299 3054 9303
rect 3066 9299 3067 9303
rect 3069 9299 3070 9303
rect 3082 9299 3083 9303
rect 3085 9299 3088 9303
rect 3090 9299 3091 9303
rect 3103 9299 3104 9303
rect 3106 9299 3107 9303
rect 3119 9299 3120 9303
rect 3122 9299 3125 9303
rect 3127 9299 3128 9303
rect 3140 9299 3141 9303
rect 3143 9299 3144 9303
rect 3156 9299 3157 9303
rect 3159 9299 3162 9303
rect 3164 9299 3165 9303
rect 3182 9299 3183 9303
rect 3185 9299 3186 9303
rect 3198 9299 3199 9303
rect 3201 9299 3202 9303
rect 3214 9299 3215 9303
rect 3217 9299 3220 9303
rect 3222 9299 3223 9303
rect 3235 9299 3236 9303
rect 3238 9299 3239 9303
rect 3251 9299 3252 9303
rect 3254 9299 3257 9303
rect 3259 9299 3260 9303
rect 3272 9299 3273 9303
rect 3275 9299 3276 9303
rect 3288 9299 3289 9303
rect 3291 9299 3294 9303
rect 3296 9299 3297 9303
rect 3314 9299 3315 9303
rect 3317 9299 3318 9303
rect 3330 9299 3331 9303
rect 3333 9299 3334 9303
rect 3346 9299 3347 9303
rect 3349 9299 3352 9303
rect 3354 9299 3355 9303
rect 3367 9299 3368 9303
rect 3370 9299 3371 9303
rect 3800 9299 3801 9303
rect 3803 9299 3806 9303
rect 3808 9299 3809 9303
rect 3821 9299 3822 9303
rect 3824 9299 3825 9303
rect 3837 9299 3838 9303
rect 3840 9299 3843 9303
rect 3845 9299 3846 9303
rect 3863 9299 3864 9303
rect 3866 9299 3867 9303
rect 3879 9299 3880 9303
rect 3882 9299 3883 9303
rect 3895 9299 3896 9303
rect 3898 9299 3901 9303
rect 3903 9299 3904 9303
rect 3916 9299 3917 9303
rect 3919 9299 3920 9303
rect 3932 9299 3933 9303
rect 3935 9299 3938 9303
rect 3940 9299 3941 9303
rect 3953 9299 3954 9303
rect 3956 9299 3957 9303
rect 3969 9299 3970 9303
rect 3972 9299 3975 9303
rect 3977 9299 3978 9303
rect 3995 9299 3996 9303
rect 3998 9299 3999 9303
rect 4011 9299 4012 9303
rect 4014 9299 4015 9303
rect 4027 9299 4028 9303
rect 4030 9299 4033 9303
rect 4035 9299 4036 9303
rect 4048 9299 4049 9303
rect 4051 9299 4052 9303
rect 4064 9299 4065 9303
rect 4067 9299 4070 9303
rect 4072 9299 4073 9303
rect 4085 9299 4086 9303
rect 4088 9299 4089 9303
rect 4101 9299 4102 9303
rect 4104 9299 4107 9303
rect 4109 9299 4110 9303
rect 4127 9299 4128 9303
rect 4130 9299 4131 9303
rect 4143 9299 4144 9303
rect 4146 9299 4147 9303
rect 4159 9299 4160 9303
rect 4162 9299 4165 9303
rect 4167 9299 4168 9303
rect 4180 9299 4181 9303
rect 4183 9299 4184 9303
rect 4196 9299 4197 9303
rect 4199 9299 4202 9303
rect 4204 9299 4205 9303
rect 4217 9299 4218 9303
rect 4220 9299 4221 9303
rect 4233 9299 4234 9303
rect 4236 9299 4239 9303
rect 4241 9299 4242 9303
rect 4259 9299 4260 9303
rect 4262 9299 4263 9303
rect 4275 9299 4276 9303
rect 4278 9299 4279 9303
rect 4291 9299 4292 9303
rect 4294 9299 4297 9303
rect 4299 9299 4300 9303
rect 4312 9299 4313 9303
rect 4315 9299 4316 9303
rect 2503 9266 2504 9270
rect 2506 9266 2509 9270
rect 2511 9266 2512 9270
rect 2524 9266 2525 9270
rect 2527 9266 2528 9270
rect 2540 9266 2541 9270
rect 2543 9266 2546 9270
rect 2548 9266 2549 9270
rect 2566 9266 2567 9270
rect 2569 9266 2570 9270
rect 2582 9266 2583 9270
rect 2585 9266 2586 9270
rect 2598 9266 2599 9270
rect 2601 9266 2604 9270
rect 2606 9266 2607 9270
rect 2619 9266 2620 9270
rect 2622 9266 2623 9270
rect 3448 9266 3449 9270
rect 3451 9266 3454 9270
rect 3456 9266 3457 9270
rect 3469 9266 3470 9270
rect 3472 9266 3473 9270
rect 3485 9266 3486 9270
rect 3488 9266 3491 9270
rect 3493 9266 3494 9270
rect 3511 9266 3512 9270
rect 3514 9266 3515 9270
rect 3527 9266 3528 9270
rect 3530 9266 3531 9270
rect 3543 9266 3544 9270
rect 3546 9266 3549 9270
rect 3551 9266 3552 9270
rect 3564 9266 3565 9270
rect 3567 9266 3568 9270
rect 2627 9229 2628 9233
rect 2630 9229 2631 9233
rect 3034 9233 3035 9237
rect 3037 9233 3038 9237
rect 3058 9229 3061 9233
rect 3063 9229 3066 9233
rect 3068 9229 3069 9233
rect 3115 9233 3116 9237
rect 3118 9233 3119 9237
rect 3139 9229 3142 9233
rect 3144 9229 3147 9233
rect 3149 9229 3150 9233
rect 3088 9225 3089 9229
rect 3091 9225 3092 9229
rect 2510 9220 2511 9224
rect 2513 9220 2514 9224
rect 2860 9220 2861 9224
rect 2863 9220 2864 9224
rect 2876 9220 2877 9224
rect 2879 9220 2880 9224
rect 2892 9220 2893 9224
rect 2895 9220 2896 9224
rect 2911 9220 2916 9224
rect 2918 9220 2921 9224
rect 2923 9220 2924 9224
rect 2945 9220 2947 9224
rect 2949 9220 2950 9224
rect 2967 9220 2968 9224
rect 2970 9220 2971 9224
rect 2983 9220 2988 9224
rect 2990 9220 2993 9224
rect 2995 9220 2996 9224
rect 3010 9220 3011 9224
rect 3013 9220 3014 9224
rect 3169 9225 3170 9229
rect 3172 9225 3173 9229
rect 3572 9229 3573 9233
rect 3575 9229 3576 9233
rect 3979 9233 3980 9237
rect 3982 9233 3983 9237
rect 4003 9229 4006 9233
rect 4008 9229 4011 9233
rect 4013 9229 4014 9233
rect 4060 9233 4061 9237
rect 4063 9233 4064 9237
rect 4084 9229 4087 9233
rect 4089 9229 4092 9233
rect 4094 9229 4095 9233
rect 4033 9225 4034 9229
rect 4036 9225 4037 9229
rect 3455 9220 3456 9224
rect 3458 9220 3459 9224
rect 3805 9220 3806 9224
rect 3808 9220 3809 9224
rect 3821 9220 3822 9224
rect 3824 9220 3825 9224
rect 3837 9220 3838 9224
rect 3840 9220 3841 9224
rect 3856 9220 3861 9224
rect 3863 9220 3866 9224
rect 3868 9220 3869 9224
rect 3890 9220 3892 9224
rect 3894 9220 3895 9224
rect 3912 9220 3913 9224
rect 3915 9220 3916 9224
rect 3928 9220 3933 9224
rect 3935 9220 3938 9224
rect 3940 9220 3941 9224
rect 3955 9220 3956 9224
rect 3958 9220 3959 9224
rect 4114 9225 4115 9229
rect 4117 9225 4118 9229
rect 2860 9174 2861 9178
rect 2863 9174 2864 9178
rect 2876 9174 2877 9178
rect 2879 9174 2880 9178
rect 2892 9174 2893 9178
rect 2895 9174 2896 9178
rect 2911 9174 2916 9178
rect 2918 9174 2921 9178
rect 2923 9174 2924 9178
rect 2945 9174 2947 9178
rect 2949 9174 2950 9178
rect 2967 9174 2968 9178
rect 2970 9174 2971 9178
rect 2983 9174 2988 9178
rect 2990 9174 2993 9178
rect 2995 9174 2996 9178
rect 3010 9174 3011 9178
rect 3013 9174 3014 9178
rect 2494 9164 2495 9168
rect 2497 9164 2498 9168
rect 2510 9164 2511 9168
rect 2513 9164 2516 9168
rect 2518 9164 2519 9168
rect 2531 9164 2532 9168
rect 2534 9164 2535 9168
rect 2547 9164 2548 9168
rect 2550 9164 2551 9168
rect 2568 9164 2569 9168
rect 2571 9164 2574 9168
rect 2576 9164 2577 9168
rect 2589 9164 2590 9168
rect 2592 9164 2593 9168
rect 2605 9164 2606 9168
rect 2608 9164 2611 9168
rect 2613 9164 2614 9168
rect 3058 9173 3061 9177
rect 3063 9173 3066 9177
rect 3068 9173 3069 9177
rect 3139 9173 3142 9177
rect 3144 9173 3147 9177
rect 3149 9173 3150 9177
rect 3805 9174 3806 9178
rect 3808 9174 3809 9178
rect 3821 9174 3822 9178
rect 3824 9174 3825 9178
rect 3837 9174 3838 9178
rect 3840 9174 3841 9178
rect 3856 9174 3861 9178
rect 3863 9174 3866 9178
rect 3868 9174 3869 9178
rect 3890 9174 3892 9178
rect 3894 9174 3895 9178
rect 3912 9174 3913 9178
rect 3915 9174 3916 9178
rect 3928 9174 3933 9178
rect 3935 9174 3938 9178
rect 3940 9174 3941 9178
rect 3955 9174 3956 9178
rect 3958 9174 3959 9178
rect 3439 9164 3440 9168
rect 3442 9164 3443 9168
rect 3455 9164 3456 9168
rect 3458 9164 3461 9168
rect 3463 9164 3464 9168
rect 3476 9164 3477 9168
rect 3479 9164 3480 9168
rect 3492 9164 3493 9168
rect 3495 9164 3496 9168
rect 3513 9164 3514 9168
rect 3516 9164 3519 9168
rect 3521 9164 3522 9168
rect 3534 9164 3535 9168
rect 3537 9164 3538 9168
rect 3550 9164 3551 9168
rect 3553 9164 3556 9168
rect 3558 9164 3559 9168
rect 4003 9173 4006 9177
rect 4008 9173 4011 9177
rect 4013 9173 4014 9177
rect 4084 9173 4087 9177
rect 4089 9173 4092 9177
rect 4094 9173 4095 9177
rect 3058 9097 3061 9101
rect 3063 9097 3066 9101
rect 3068 9097 3069 9101
rect 3139 9101 3140 9105
rect 3142 9101 3143 9105
rect 3163 9097 3166 9101
rect 3168 9097 3171 9101
rect 3173 9097 3174 9101
rect 3088 9093 3089 9097
rect 3091 9093 3092 9097
rect 2860 9088 2861 9092
rect 2863 9088 2864 9092
rect 2876 9088 2877 9092
rect 2879 9088 2880 9092
rect 2892 9088 2893 9092
rect 2895 9088 2896 9092
rect 2911 9088 2916 9092
rect 2918 9088 2921 9092
rect 2923 9088 2924 9092
rect 2945 9088 2947 9092
rect 2949 9088 2950 9092
rect 2967 9088 2968 9092
rect 2970 9088 2971 9092
rect 2983 9088 2988 9092
rect 2990 9088 2993 9092
rect 2995 9088 2996 9092
rect 3010 9088 3011 9092
rect 3013 9088 3014 9092
rect 3193 9093 3194 9097
rect 3196 9093 3197 9097
rect 3370 9072 3371 9076
rect 3373 9072 3374 9076
rect 3394 9068 3397 9072
rect 3399 9068 3402 9072
rect 3404 9068 3405 9072
rect 3424 9064 3425 9068
rect 3427 9064 3428 9068
rect 4003 9097 4006 9101
rect 4008 9097 4011 9101
rect 4013 9097 4014 9101
rect 4084 9101 4085 9105
rect 4087 9101 4088 9105
rect 4108 9097 4111 9101
rect 4113 9097 4116 9101
rect 4118 9097 4119 9101
rect 4033 9093 4034 9097
rect 4036 9093 4037 9097
rect 3805 9088 3806 9092
rect 3808 9088 3809 9092
rect 3821 9088 3822 9092
rect 3824 9088 3825 9092
rect 3837 9088 3838 9092
rect 3840 9088 3841 9092
rect 3856 9088 3861 9092
rect 3863 9088 3866 9092
rect 3868 9088 3869 9092
rect 3890 9088 3892 9092
rect 3894 9088 3895 9092
rect 3912 9088 3913 9092
rect 3915 9088 3916 9092
rect 3928 9088 3933 9092
rect 3935 9088 3938 9092
rect 3940 9088 3941 9092
rect 3955 9088 3956 9092
rect 3958 9088 3959 9092
rect 4138 9093 4139 9097
rect 4141 9093 4142 9097
rect 2860 9042 2861 9046
rect 2863 9042 2864 9046
rect 2876 9042 2877 9046
rect 2879 9042 2880 9046
rect 2892 9042 2893 9046
rect 2895 9042 2896 9046
rect 2911 9042 2916 9046
rect 2918 9042 2921 9046
rect 2923 9042 2924 9046
rect 2945 9042 2947 9046
rect 2949 9042 2950 9046
rect 2967 9042 2968 9046
rect 2970 9042 2971 9046
rect 2983 9042 2988 9046
rect 2990 9042 2993 9046
rect 2995 9042 2996 9046
rect 3010 9042 3011 9046
rect 3013 9042 3014 9046
rect 3058 9042 3061 9046
rect 3063 9042 3066 9046
rect 3068 9042 3069 9046
rect 3163 9042 3166 9046
rect 3168 9042 3171 9046
rect 3173 9042 3174 9046
rect 3556 9033 3557 9045
rect 3559 9033 3560 9045
rect 3609 9033 3610 9045
rect 3612 9033 3613 9045
rect 3805 9042 3806 9046
rect 3808 9042 3809 9046
rect 3821 9042 3822 9046
rect 3824 9042 3825 9046
rect 3837 9042 3838 9046
rect 3840 9042 3841 9046
rect 3856 9042 3861 9046
rect 3863 9042 3866 9046
rect 3868 9042 3869 9046
rect 3890 9042 3892 9046
rect 3894 9042 3895 9046
rect 3912 9042 3913 9046
rect 3915 9042 3916 9046
rect 3928 9042 3933 9046
rect 3935 9042 3938 9046
rect 3940 9042 3941 9046
rect 3955 9042 3956 9046
rect 3958 9042 3959 9046
rect 4003 9042 4006 9046
rect 4008 9042 4011 9046
rect 4013 9042 4014 9046
rect 4108 9042 4111 9046
rect 4113 9042 4116 9046
rect 4118 9042 4119 9046
rect 3394 9008 3397 9012
rect 3399 9008 3402 9012
rect 3404 9008 3405 9012
rect 3058 8965 3061 8969
rect 3063 8965 3066 8969
rect 3068 8965 3069 8969
rect 3115 8969 3116 8973
rect 3118 8969 3119 8973
rect 3139 8965 3142 8969
rect 3144 8965 3147 8969
rect 3149 8965 3150 8969
rect 3205 8969 3206 8973
rect 3208 8969 3209 8973
rect 3229 8965 3232 8969
rect 3234 8965 3237 8969
rect 3239 8965 3240 8969
rect 3088 8961 3089 8965
rect 3091 8961 3092 8965
rect 2860 8956 2861 8960
rect 2863 8956 2864 8960
rect 2876 8956 2877 8960
rect 2879 8956 2880 8960
rect 2892 8956 2893 8960
rect 2895 8956 2896 8960
rect 2911 8956 2916 8960
rect 2918 8956 2921 8960
rect 2923 8956 2924 8960
rect 2945 8956 2947 8960
rect 2949 8956 2950 8960
rect 2967 8956 2968 8960
rect 2970 8956 2971 8960
rect 2983 8956 2988 8960
rect 2990 8956 2993 8960
rect 2995 8956 2996 8960
rect 3010 8956 3011 8960
rect 3013 8956 3014 8960
rect 3169 8961 3170 8965
rect 3172 8961 3173 8965
rect 3259 8961 3260 8965
rect 3262 8961 3263 8965
rect 3348 8942 3349 8946
rect 3351 8942 3352 8946
rect 3370 8942 3371 8946
rect 3373 8942 3374 8946
rect 3394 8938 3397 8942
rect 3399 8938 3402 8942
rect 3404 8938 3405 8942
rect 3424 8934 3425 8938
rect 3427 8934 3428 8938
rect 4003 8965 4006 8969
rect 4008 8965 4011 8969
rect 4013 8965 4014 8969
rect 4060 8969 4061 8973
rect 4063 8969 4064 8973
rect 4084 8965 4087 8969
rect 4089 8965 4092 8969
rect 4094 8965 4095 8969
rect 4150 8969 4151 8973
rect 4153 8969 4154 8973
rect 4174 8965 4177 8969
rect 4179 8965 4182 8969
rect 4184 8965 4185 8969
rect 4033 8961 4034 8965
rect 4036 8961 4037 8965
rect 3805 8956 3806 8960
rect 3808 8956 3809 8960
rect 3821 8956 3822 8960
rect 3824 8956 3825 8960
rect 3837 8956 3838 8960
rect 3840 8956 3841 8960
rect 3856 8956 3861 8960
rect 3863 8956 3866 8960
rect 3868 8956 3869 8960
rect 3890 8956 3892 8960
rect 3894 8956 3895 8960
rect 3912 8956 3913 8960
rect 3915 8956 3916 8960
rect 3928 8956 3933 8960
rect 3935 8956 3938 8960
rect 3940 8956 3941 8960
rect 3955 8956 3956 8960
rect 3958 8956 3959 8960
rect 4114 8961 4115 8965
rect 4117 8961 4118 8965
rect 4204 8961 4205 8965
rect 4207 8961 4208 8965
rect 2860 8910 2861 8914
rect 2863 8910 2864 8914
rect 2876 8910 2877 8914
rect 2879 8910 2880 8914
rect 2892 8910 2893 8914
rect 2895 8910 2896 8914
rect 2911 8910 2916 8914
rect 2918 8910 2921 8914
rect 2923 8910 2924 8914
rect 2945 8910 2947 8914
rect 2949 8910 2950 8914
rect 2967 8910 2968 8914
rect 2970 8910 2971 8914
rect 2983 8910 2988 8914
rect 2990 8910 2993 8914
rect 2995 8910 2996 8914
rect 3010 8910 3011 8914
rect 3013 8910 3014 8914
rect 3058 8907 3061 8911
rect 3063 8907 3066 8911
rect 3068 8907 3069 8911
rect 3139 8907 3142 8911
rect 3144 8907 3147 8911
rect 3149 8907 3150 8911
rect 3229 8907 3232 8911
rect 3234 8907 3237 8911
rect 3239 8907 3240 8911
rect 3462 8903 3463 8915
rect 3465 8903 3466 8915
rect 3515 8903 3516 8915
rect 3518 8903 3519 8915
rect 3805 8910 3806 8914
rect 3808 8910 3809 8914
rect 3821 8910 3822 8914
rect 3824 8910 3825 8914
rect 3837 8910 3838 8914
rect 3840 8910 3841 8914
rect 3856 8910 3861 8914
rect 3863 8910 3866 8914
rect 3868 8910 3869 8914
rect 3890 8910 3892 8914
rect 3894 8910 3895 8914
rect 3912 8910 3913 8914
rect 3915 8910 3916 8914
rect 3928 8910 3933 8914
rect 3935 8910 3938 8914
rect 3940 8910 3941 8914
rect 3955 8910 3956 8914
rect 3958 8910 3959 8914
rect 4003 8907 4006 8911
rect 4008 8907 4011 8911
rect 4013 8907 4014 8911
rect 4084 8907 4087 8911
rect 4089 8907 4092 8911
rect 4094 8907 4095 8911
rect 4174 8907 4177 8911
rect 4179 8907 4182 8911
rect 4184 8907 4185 8911
rect 3394 8878 3397 8882
rect 3399 8878 3402 8882
rect 3404 8878 3405 8882
rect 3058 8833 3061 8837
rect 3063 8833 3066 8837
rect 3068 8833 3069 8837
rect 3088 8829 3089 8833
rect 3091 8829 3092 8833
rect 2860 8824 2861 8828
rect 2863 8824 2864 8828
rect 2876 8824 2877 8828
rect 2879 8824 2880 8828
rect 2892 8824 2893 8828
rect 2895 8824 2896 8828
rect 2911 8824 2916 8828
rect 2918 8824 2921 8828
rect 2923 8824 2924 8828
rect 2945 8824 2947 8828
rect 2949 8824 2950 8828
rect 2967 8824 2968 8828
rect 2970 8824 2971 8828
rect 2983 8824 2988 8828
rect 2990 8824 2993 8828
rect 2995 8824 2996 8828
rect 3010 8824 3011 8828
rect 3013 8824 3014 8828
rect 4003 8833 4006 8837
rect 4008 8833 4011 8837
rect 4013 8833 4014 8837
rect 4033 8829 4034 8833
rect 4036 8829 4037 8833
rect 3805 8824 3806 8828
rect 3808 8824 3809 8828
rect 3821 8824 3822 8828
rect 3824 8824 3825 8828
rect 3837 8824 3838 8828
rect 3840 8824 3841 8828
rect 3856 8824 3861 8828
rect 3863 8824 3866 8828
rect 3868 8824 3869 8828
rect 3890 8824 3892 8828
rect 3894 8824 3895 8828
rect 3912 8824 3913 8828
rect 3915 8824 3916 8828
rect 3928 8824 3933 8828
rect 3935 8824 3938 8828
rect 3940 8824 3941 8828
rect 3955 8824 3956 8828
rect 3958 8824 3959 8828
rect 2860 8778 2861 8782
rect 2863 8778 2864 8782
rect 2876 8778 2877 8782
rect 2879 8778 2880 8782
rect 2892 8778 2893 8782
rect 2895 8778 2896 8782
rect 2911 8778 2916 8782
rect 2918 8778 2921 8782
rect 2923 8778 2924 8782
rect 2945 8778 2947 8782
rect 2949 8778 2950 8782
rect 2967 8778 2968 8782
rect 2970 8778 2971 8782
rect 2983 8778 2988 8782
rect 2990 8778 2993 8782
rect 2995 8778 2996 8782
rect 3010 8778 3011 8782
rect 3013 8778 3014 8782
rect 3094 8778 3095 8782
rect 3097 8778 3098 8782
rect 3102 8778 3108 8782
rect 3112 8778 3113 8782
rect 3115 8778 3116 8782
rect 3137 8778 3138 8782
rect 3140 8778 3141 8782
rect 3153 8778 3154 8782
rect 3156 8778 3157 8782
rect 3172 8778 3177 8782
rect 3179 8778 3182 8782
rect 3184 8778 3185 8782
rect 3206 8778 3208 8782
rect 3210 8778 3211 8782
rect 3228 8778 3229 8782
rect 3231 8778 3232 8782
rect 3244 8778 3249 8782
rect 3251 8778 3254 8782
rect 3256 8778 3257 8782
rect 3271 8778 3272 8782
rect 3274 8778 3275 8782
rect 2371 8764 2372 8768
rect 2374 8764 2377 8768
rect 2379 8764 2380 8768
rect 2392 8764 2393 8768
rect 2395 8764 2396 8768
rect 2408 8764 2409 8768
rect 2411 8764 2414 8768
rect 2416 8764 2417 8768
rect 2434 8764 2435 8768
rect 2437 8764 2438 8768
rect 2450 8764 2451 8768
rect 2453 8764 2454 8768
rect 2466 8764 2467 8768
rect 2469 8764 2472 8768
rect 2474 8764 2475 8768
rect 2487 8764 2488 8768
rect 2490 8764 2491 8768
rect 2503 8764 2504 8768
rect 2506 8764 2509 8768
rect 2511 8764 2512 8768
rect 2524 8764 2525 8768
rect 2527 8764 2528 8768
rect 2540 8764 2541 8768
rect 2543 8764 2546 8768
rect 2548 8764 2549 8768
rect 2566 8764 2567 8768
rect 2569 8764 2570 8768
rect 2582 8764 2583 8768
rect 2585 8764 2586 8768
rect 2598 8764 2599 8768
rect 2601 8764 2604 8768
rect 2606 8764 2607 8768
rect 2619 8764 2620 8768
rect 2622 8764 2623 8768
rect 2635 8764 2636 8768
rect 2638 8764 2641 8768
rect 2643 8764 2644 8768
rect 2656 8764 2657 8768
rect 2659 8764 2660 8768
rect 2672 8764 2673 8768
rect 2675 8764 2678 8768
rect 2680 8764 2681 8768
rect 2698 8764 2699 8768
rect 2701 8764 2702 8768
rect 2714 8764 2715 8768
rect 2717 8764 2718 8768
rect 2730 8764 2731 8768
rect 2733 8764 2736 8768
rect 2738 8764 2739 8768
rect 2751 8764 2752 8768
rect 2754 8764 2755 8768
rect 3058 8771 3061 8775
rect 3063 8771 3066 8775
rect 3068 8771 3069 8775
rect 3805 8778 3806 8782
rect 3808 8778 3809 8782
rect 3821 8778 3822 8782
rect 3824 8778 3825 8782
rect 3837 8778 3838 8782
rect 3840 8778 3841 8782
rect 3856 8778 3861 8782
rect 3863 8778 3866 8782
rect 3868 8778 3869 8782
rect 3890 8778 3892 8782
rect 3894 8778 3895 8782
rect 3912 8778 3913 8782
rect 3915 8778 3916 8782
rect 3928 8778 3933 8782
rect 3935 8778 3938 8782
rect 3940 8778 3941 8782
rect 3955 8778 3956 8782
rect 3958 8778 3959 8782
rect 4039 8778 4040 8782
rect 4042 8778 4043 8782
rect 4047 8778 4053 8782
rect 4057 8778 4058 8782
rect 4060 8778 4061 8782
rect 4082 8778 4083 8782
rect 4085 8778 4086 8782
rect 4098 8778 4099 8782
rect 4101 8778 4102 8782
rect 4117 8778 4122 8782
rect 4124 8778 4127 8782
rect 4129 8778 4130 8782
rect 4151 8778 4153 8782
rect 4155 8778 4156 8782
rect 4173 8778 4174 8782
rect 4176 8778 4177 8782
rect 4189 8778 4194 8782
rect 4196 8778 4199 8782
rect 4201 8778 4202 8782
rect 4216 8778 4217 8782
rect 4219 8778 4220 8782
rect 3316 8764 3317 8768
rect 3319 8764 3322 8768
rect 3324 8764 3325 8768
rect 3337 8764 3338 8768
rect 3340 8764 3341 8768
rect 3353 8764 3354 8768
rect 3356 8764 3359 8768
rect 3361 8764 3362 8768
rect 3379 8764 3380 8768
rect 3382 8764 3383 8768
rect 3395 8764 3396 8768
rect 3398 8764 3399 8768
rect 3411 8764 3412 8768
rect 3414 8764 3417 8768
rect 3419 8764 3420 8768
rect 3432 8764 3433 8768
rect 3435 8764 3436 8768
rect 3448 8764 3449 8768
rect 3451 8764 3454 8768
rect 3456 8764 3457 8768
rect 3469 8764 3470 8768
rect 3472 8764 3473 8768
rect 3485 8764 3486 8768
rect 3488 8764 3491 8768
rect 3493 8764 3494 8768
rect 3511 8764 3512 8768
rect 3514 8764 3515 8768
rect 3527 8764 3528 8768
rect 3530 8764 3531 8768
rect 3543 8764 3544 8768
rect 3546 8764 3549 8768
rect 3551 8764 3552 8768
rect 3564 8764 3565 8768
rect 3567 8764 3568 8768
rect 3580 8764 3581 8768
rect 3583 8764 3586 8768
rect 3588 8764 3589 8768
rect 3601 8764 3602 8768
rect 3604 8764 3605 8768
rect 3617 8764 3618 8768
rect 3620 8764 3623 8768
rect 3625 8764 3626 8768
rect 3643 8764 3644 8768
rect 3646 8764 3647 8768
rect 3659 8764 3660 8768
rect 3662 8764 3663 8768
rect 3675 8764 3676 8768
rect 3678 8764 3681 8768
rect 3683 8764 3684 8768
rect 3696 8764 3697 8768
rect 3699 8764 3700 8768
rect 4003 8771 4006 8775
rect 4008 8771 4011 8775
rect 4013 8771 4014 8775
rect 2486 8720 2487 8724
rect 2489 8720 2490 8724
rect 2510 8720 2511 8724
rect 2513 8720 2514 8724
rect 3284 8724 3288 8725
rect 3284 8721 3288 8722
rect 3431 8720 3432 8724
rect 3434 8720 3435 8724
rect 3455 8720 3456 8724
rect 3458 8720 3459 8724
rect 4229 8724 4233 8725
rect 4229 8721 4233 8722
rect 2506 8707 2507 8711
rect 2509 8707 2510 8711
rect 3451 8707 3452 8711
rect 3454 8707 3455 8711
rect 2498 8695 2502 8696
rect 2498 8692 2502 8693
rect 3443 8695 3447 8696
rect 3443 8692 3447 8693
rect 2486 8684 2487 8688
rect 2489 8684 2490 8688
rect 2510 8684 2511 8688
rect 2513 8684 2514 8688
rect 3431 8684 3432 8688
rect 3434 8684 3435 8688
rect 3455 8684 3456 8688
rect 3458 8684 3459 8688
rect 3154 8652 3155 8656
rect 3157 8652 3160 8656
rect 3162 8652 3163 8656
rect 3175 8652 3176 8656
rect 3178 8652 3179 8656
rect 3191 8652 3192 8656
rect 3194 8652 3197 8656
rect 3199 8652 3200 8656
rect 3217 8652 3218 8656
rect 3220 8652 3221 8656
rect 3233 8652 3234 8656
rect 3236 8652 3237 8656
rect 3249 8652 3250 8656
rect 3252 8652 3255 8656
rect 3257 8652 3258 8656
rect 3270 8652 3271 8656
rect 3273 8652 3274 8656
rect 4099 8652 4100 8656
rect 4102 8652 4105 8656
rect 4107 8652 4108 8656
rect 4120 8652 4121 8656
rect 4123 8652 4124 8656
rect 4136 8652 4137 8656
rect 4139 8652 4142 8656
rect 4144 8652 4145 8656
rect 4162 8652 4163 8656
rect 4165 8652 4166 8656
rect 4178 8652 4179 8656
rect 4181 8652 4182 8656
rect 4194 8652 4195 8656
rect 4197 8652 4200 8656
rect 4202 8652 4203 8656
rect 4215 8652 4216 8656
rect 4218 8652 4219 8656
rect 2371 8622 2372 8626
rect 2374 8622 2377 8626
rect 2379 8622 2380 8626
rect 2392 8622 2393 8626
rect 2395 8622 2396 8626
rect 2408 8622 2409 8626
rect 2411 8622 2414 8626
rect 2416 8622 2417 8626
rect 2434 8622 2435 8626
rect 2437 8622 2438 8626
rect 2450 8622 2451 8626
rect 2453 8622 2454 8626
rect 2466 8622 2467 8626
rect 2469 8622 2472 8626
rect 2474 8622 2475 8626
rect 2487 8622 2488 8626
rect 2490 8622 2491 8626
rect 2503 8622 2504 8626
rect 2506 8622 2509 8626
rect 2511 8622 2512 8626
rect 2524 8622 2525 8626
rect 2527 8622 2528 8626
rect 2540 8622 2541 8626
rect 2543 8622 2546 8626
rect 2548 8622 2549 8626
rect 2566 8622 2567 8626
rect 2569 8622 2570 8626
rect 2582 8622 2583 8626
rect 2585 8622 2586 8626
rect 2598 8622 2599 8626
rect 2601 8622 2604 8626
rect 2606 8622 2607 8626
rect 2619 8622 2620 8626
rect 2622 8622 2623 8626
rect 2635 8622 2636 8626
rect 2638 8622 2641 8626
rect 2643 8622 2644 8626
rect 2656 8622 2657 8626
rect 2659 8622 2660 8626
rect 2672 8622 2673 8626
rect 2675 8622 2678 8626
rect 2680 8622 2681 8626
rect 2698 8622 2699 8626
rect 2701 8622 2702 8626
rect 2714 8622 2715 8626
rect 2717 8622 2718 8626
rect 2730 8622 2731 8626
rect 2733 8622 2736 8626
rect 2738 8622 2739 8626
rect 2751 8622 2752 8626
rect 2754 8622 2755 8626
rect 3316 8622 3317 8626
rect 3319 8622 3322 8626
rect 3324 8622 3325 8626
rect 3337 8622 3338 8626
rect 3340 8622 3341 8626
rect 3353 8622 3354 8626
rect 3356 8622 3359 8626
rect 3361 8622 3362 8626
rect 3379 8622 3380 8626
rect 3382 8622 3383 8626
rect 3395 8622 3396 8626
rect 3398 8622 3399 8626
rect 3411 8622 3412 8626
rect 3414 8622 3417 8626
rect 3419 8622 3420 8626
rect 3432 8622 3433 8626
rect 3435 8622 3436 8626
rect 3448 8622 3449 8626
rect 3451 8622 3454 8626
rect 3456 8622 3457 8626
rect 3469 8622 3470 8626
rect 3472 8622 3473 8626
rect 3485 8622 3486 8626
rect 3488 8622 3491 8626
rect 3493 8622 3494 8626
rect 3511 8622 3512 8626
rect 3514 8622 3515 8626
rect 3527 8622 3528 8626
rect 3530 8622 3531 8626
rect 3543 8622 3544 8626
rect 3546 8622 3549 8626
rect 3551 8622 3552 8626
rect 3564 8622 3565 8626
rect 3567 8622 3568 8626
rect 3580 8622 3581 8626
rect 3583 8622 3586 8626
rect 3588 8622 3589 8626
rect 3601 8622 3602 8626
rect 3604 8622 3605 8626
rect 3617 8622 3618 8626
rect 3620 8622 3623 8626
rect 3625 8622 3626 8626
rect 3643 8622 3644 8626
rect 3646 8622 3647 8626
rect 3659 8622 3660 8626
rect 3662 8622 3663 8626
rect 3675 8622 3676 8626
rect 3678 8622 3681 8626
rect 3683 8622 3684 8626
rect 3696 8622 3697 8626
rect 3699 8622 3700 8626
rect 3296 8578 3300 8579
rect 3296 8575 3300 8576
rect 4241 8578 4245 8579
rect 4241 8575 4245 8576
rect 3154 8566 3155 8570
rect 3157 8566 3160 8570
rect 3162 8566 3163 8570
rect 3175 8566 3176 8570
rect 3178 8566 3179 8570
rect 3191 8566 3192 8570
rect 3194 8566 3197 8570
rect 3199 8566 3200 8570
rect 3217 8566 3218 8570
rect 3220 8566 3221 8570
rect 3233 8566 3234 8570
rect 3236 8566 3237 8570
rect 3249 8566 3250 8570
rect 3252 8566 3255 8570
rect 3257 8566 3258 8570
rect 3270 8566 3271 8570
rect 3273 8566 3274 8570
rect 4099 8566 4100 8570
rect 4102 8566 4105 8570
rect 4107 8566 4108 8570
rect 4120 8566 4121 8570
rect 4123 8566 4124 8570
rect 4136 8566 4137 8570
rect 4139 8566 4142 8570
rect 4144 8566 4145 8570
rect 4162 8566 4163 8570
rect 4165 8566 4166 8570
rect 4178 8566 4179 8570
rect 4181 8566 4182 8570
rect 4194 8566 4195 8570
rect 4197 8566 4200 8570
rect 4202 8566 4203 8570
rect 4215 8566 4216 8570
rect 4218 8566 4219 8570
rect 2371 8536 2372 8540
rect 2374 8536 2377 8540
rect 2379 8536 2380 8540
rect 2392 8536 2393 8540
rect 2395 8536 2396 8540
rect 2408 8536 2409 8540
rect 2411 8536 2414 8540
rect 2416 8536 2417 8540
rect 2434 8536 2435 8540
rect 2437 8536 2438 8540
rect 2450 8536 2451 8540
rect 2453 8536 2454 8540
rect 2466 8536 2467 8540
rect 2469 8536 2472 8540
rect 2474 8536 2475 8540
rect 2487 8536 2488 8540
rect 2490 8536 2491 8540
rect 2503 8536 2504 8540
rect 2506 8536 2509 8540
rect 2511 8536 2512 8540
rect 2524 8536 2525 8540
rect 2527 8536 2528 8540
rect 2540 8536 2541 8540
rect 2543 8536 2546 8540
rect 2548 8536 2549 8540
rect 2566 8536 2567 8540
rect 2569 8536 2570 8540
rect 2582 8536 2583 8540
rect 2585 8536 2586 8540
rect 2598 8536 2599 8540
rect 2601 8536 2604 8540
rect 2606 8536 2607 8540
rect 2619 8536 2620 8540
rect 2622 8536 2623 8540
rect 2635 8536 2636 8540
rect 2638 8536 2641 8540
rect 2643 8536 2644 8540
rect 2656 8536 2657 8540
rect 2659 8536 2660 8540
rect 2672 8536 2673 8540
rect 2675 8536 2678 8540
rect 2680 8536 2681 8540
rect 2698 8536 2699 8540
rect 2701 8536 2702 8540
rect 2714 8536 2715 8540
rect 2717 8536 2718 8540
rect 2730 8536 2731 8540
rect 2733 8536 2736 8540
rect 2738 8536 2739 8540
rect 2751 8536 2752 8540
rect 2754 8536 2755 8540
rect 3316 8536 3317 8540
rect 3319 8536 3322 8540
rect 3324 8536 3325 8540
rect 3337 8536 3338 8540
rect 3340 8536 3341 8540
rect 3353 8536 3354 8540
rect 3356 8536 3359 8540
rect 3361 8536 3362 8540
rect 3379 8536 3380 8540
rect 3382 8536 3383 8540
rect 3395 8536 3396 8540
rect 3398 8536 3399 8540
rect 3411 8536 3412 8540
rect 3414 8536 3417 8540
rect 3419 8536 3420 8540
rect 3432 8536 3433 8540
rect 3435 8536 3436 8540
rect 3448 8536 3449 8540
rect 3451 8536 3454 8540
rect 3456 8536 3457 8540
rect 3469 8536 3470 8540
rect 3472 8536 3473 8540
rect 3485 8536 3486 8540
rect 3488 8536 3491 8540
rect 3493 8536 3494 8540
rect 3511 8536 3512 8540
rect 3514 8536 3515 8540
rect 3527 8536 3528 8540
rect 3530 8536 3531 8540
rect 3543 8536 3544 8540
rect 3546 8536 3549 8540
rect 3551 8536 3552 8540
rect 3564 8536 3565 8540
rect 3567 8536 3568 8540
rect 3580 8536 3581 8540
rect 3583 8536 3586 8540
rect 3588 8536 3589 8540
rect 3601 8536 3602 8540
rect 3604 8536 3605 8540
rect 3617 8536 3618 8540
rect 3620 8536 3623 8540
rect 3625 8536 3626 8540
rect 3643 8536 3644 8540
rect 3646 8536 3647 8540
rect 3659 8536 3660 8540
rect 3662 8536 3663 8540
rect 3675 8536 3676 8540
rect 3678 8536 3681 8540
rect 3683 8536 3684 8540
rect 3696 8536 3697 8540
rect 3699 8536 3700 8540
rect 2603 8492 2604 8496
rect 2606 8492 2607 8496
rect 2627 8492 2628 8496
rect 2630 8492 2631 8496
rect 3548 8492 3549 8496
rect 3551 8492 3552 8496
rect 3572 8492 3573 8496
rect 3575 8492 3576 8496
rect 2623 8481 2624 8485
rect 2626 8481 2627 8485
rect 3568 8481 3569 8485
rect 3571 8481 3572 8485
rect 2615 8469 2619 8470
rect 2615 8466 2619 8467
rect 3560 8469 3564 8470
rect 3560 8466 3564 8467
rect 2603 8458 2604 8462
rect 2606 8458 2607 8462
rect 2627 8458 2628 8462
rect 2630 8458 2631 8462
rect 3548 8458 3549 8462
rect 3551 8458 3552 8462
rect 3572 8458 3573 8462
rect 3575 8458 3576 8462
rect 2371 8396 2372 8400
rect 2374 8396 2377 8400
rect 2379 8396 2380 8400
rect 2392 8396 2393 8400
rect 2395 8396 2396 8400
rect 2408 8396 2409 8400
rect 2411 8396 2414 8400
rect 2416 8396 2417 8400
rect 2434 8396 2435 8400
rect 2437 8396 2438 8400
rect 2450 8396 2451 8400
rect 2453 8396 2454 8400
rect 2466 8396 2467 8400
rect 2469 8396 2472 8400
rect 2474 8396 2475 8400
rect 2487 8396 2488 8400
rect 2490 8396 2491 8400
rect 2503 8396 2504 8400
rect 2506 8396 2509 8400
rect 2511 8396 2512 8400
rect 2524 8396 2525 8400
rect 2527 8396 2528 8400
rect 2540 8396 2541 8400
rect 2543 8396 2546 8400
rect 2548 8396 2549 8400
rect 2566 8396 2567 8400
rect 2569 8396 2570 8400
rect 2582 8396 2583 8400
rect 2585 8396 2586 8400
rect 2598 8396 2599 8400
rect 2601 8396 2604 8400
rect 2606 8396 2607 8400
rect 2619 8396 2620 8400
rect 2622 8396 2623 8400
rect 2635 8396 2636 8400
rect 2638 8396 2641 8400
rect 2643 8396 2644 8400
rect 2656 8396 2657 8400
rect 2659 8396 2660 8400
rect 2672 8396 2673 8400
rect 2675 8396 2678 8400
rect 2680 8396 2681 8400
rect 2698 8396 2699 8400
rect 2701 8396 2702 8400
rect 2714 8396 2715 8400
rect 2717 8396 2718 8400
rect 2730 8396 2731 8400
rect 2733 8396 2736 8400
rect 2738 8396 2739 8400
rect 2751 8396 2752 8400
rect 2754 8396 2755 8400
rect 3316 8396 3317 8400
rect 3319 8396 3322 8400
rect 3324 8396 3325 8400
rect 3337 8396 3338 8400
rect 3340 8396 3341 8400
rect 3353 8396 3354 8400
rect 3356 8396 3359 8400
rect 3361 8396 3362 8400
rect 3379 8396 3380 8400
rect 3382 8396 3383 8400
rect 3395 8396 3396 8400
rect 3398 8396 3399 8400
rect 3411 8396 3412 8400
rect 3414 8396 3417 8400
rect 3419 8396 3420 8400
rect 3432 8396 3433 8400
rect 3435 8396 3436 8400
rect 3448 8396 3449 8400
rect 3451 8396 3454 8400
rect 3456 8396 3457 8400
rect 3469 8396 3470 8400
rect 3472 8396 3473 8400
rect 3485 8396 3486 8400
rect 3488 8396 3491 8400
rect 3493 8396 3494 8400
rect 3511 8396 3512 8400
rect 3514 8396 3515 8400
rect 3527 8396 3528 8400
rect 3530 8396 3531 8400
rect 3543 8396 3544 8400
rect 3546 8396 3549 8400
rect 3551 8396 3552 8400
rect 3564 8396 3565 8400
rect 3567 8396 3568 8400
rect 3580 8396 3581 8400
rect 3583 8396 3586 8400
rect 3588 8396 3589 8400
rect 3601 8396 3602 8400
rect 3604 8396 3605 8400
rect 3617 8396 3618 8400
rect 3620 8396 3623 8400
rect 3625 8396 3626 8400
rect 3643 8396 3644 8400
rect 3646 8396 3647 8400
rect 3659 8396 3660 8400
rect 3662 8396 3663 8400
rect 3675 8396 3676 8400
rect 3678 8396 3681 8400
rect 3683 8396 3684 8400
rect 3696 8396 3697 8400
rect 3699 8396 3700 8400
rect 2855 8317 2856 8321
rect 2858 8317 2861 8321
rect 2863 8317 2864 8321
rect 2876 8317 2877 8321
rect 2879 8317 2880 8321
rect 2892 8317 2893 8321
rect 2895 8317 2898 8321
rect 2900 8317 2901 8321
rect 2918 8317 2919 8321
rect 2921 8317 2922 8321
rect 2934 8317 2935 8321
rect 2937 8317 2938 8321
rect 2950 8317 2951 8321
rect 2953 8317 2956 8321
rect 2958 8317 2959 8321
rect 2971 8317 2972 8321
rect 2974 8317 2975 8321
rect 2987 8317 2988 8321
rect 2990 8317 2993 8321
rect 2995 8317 2996 8321
rect 3008 8317 3009 8321
rect 3011 8317 3012 8321
rect 3024 8317 3025 8321
rect 3027 8317 3030 8321
rect 3032 8317 3033 8321
rect 3050 8317 3051 8321
rect 3053 8317 3054 8321
rect 3066 8317 3067 8321
rect 3069 8317 3070 8321
rect 3082 8317 3083 8321
rect 3085 8317 3088 8321
rect 3090 8317 3091 8321
rect 3103 8317 3104 8321
rect 3106 8317 3107 8321
rect 3119 8317 3120 8321
rect 3122 8317 3125 8321
rect 3127 8317 3128 8321
rect 3140 8317 3141 8321
rect 3143 8317 3144 8321
rect 3156 8317 3157 8321
rect 3159 8317 3162 8321
rect 3164 8317 3165 8321
rect 3182 8317 3183 8321
rect 3185 8317 3186 8321
rect 3198 8317 3199 8321
rect 3201 8317 3202 8321
rect 3214 8317 3215 8321
rect 3217 8317 3220 8321
rect 3222 8317 3223 8321
rect 3235 8317 3236 8321
rect 3238 8317 3239 8321
rect 3251 8317 3252 8321
rect 3254 8317 3257 8321
rect 3259 8317 3260 8321
rect 3272 8317 3273 8321
rect 3275 8317 3276 8321
rect 3288 8317 3289 8321
rect 3291 8317 3294 8321
rect 3296 8317 3297 8321
rect 3314 8317 3315 8321
rect 3317 8317 3318 8321
rect 3330 8317 3331 8321
rect 3333 8317 3334 8321
rect 3346 8317 3347 8321
rect 3349 8317 3352 8321
rect 3354 8317 3355 8321
rect 3367 8317 3368 8321
rect 3370 8317 3371 8321
rect 3800 8317 3801 8321
rect 3803 8317 3806 8321
rect 3808 8317 3809 8321
rect 3821 8317 3822 8321
rect 3824 8317 3825 8321
rect 3837 8317 3838 8321
rect 3840 8317 3843 8321
rect 3845 8317 3846 8321
rect 3863 8317 3864 8321
rect 3866 8317 3867 8321
rect 3879 8317 3880 8321
rect 3882 8317 3883 8321
rect 3895 8317 3896 8321
rect 3898 8317 3901 8321
rect 3903 8317 3904 8321
rect 3916 8317 3917 8321
rect 3919 8317 3920 8321
rect 3932 8317 3933 8321
rect 3935 8317 3938 8321
rect 3940 8317 3941 8321
rect 3953 8317 3954 8321
rect 3956 8317 3957 8321
rect 3969 8317 3970 8321
rect 3972 8317 3975 8321
rect 3977 8317 3978 8321
rect 3995 8317 3996 8321
rect 3998 8317 3999 8321
rect 4011 8317 4012 8321
rect 4014 8317 4015 8321
rect 4027 8317 4028 8321
rect 4030 8317 4033 8321
rect 4035 8317 4036 8321
rect 4048 8317 4049 8321
rect 4051 8317 4052 8321
rect 4064 8317 4065 8321
rect 4067 8317 4070 8321
rect 4072 8317 4073 8321
rect 4085 8317 4086 8321
rect 4088 8317 4089 8321
rect 4101 8317 4102 8321
rect 4104 8317 4107 8321
rect 4109 8317 4110 8321
rect 4127 8317 4128 8321
rect 4130 8317 4131 8321
rect 4143 8317 4144 8321
rect 4146 8317 4147 8321
rect 4159 8317 4160 8321
rect 4162 8317 4165 8321
rect 4167 8317 4168 8321
rect 4180 8317 4181 8321
rect 4183 8317 4184 8321
rect 4196 8317 4197 8321
rect 4199 8317 4202 8321
rect 4204 8317 4205 8321
rect 4217 8317 4218 8321
rect 4220 8317 4221 8321
rect 4233 8317 4234 8321
rect 4236 8317 4239 8321
rect 4241 8317 4242 8321
rect 4259 8317 4260 8321
rect 4262 8317 4263 8321
rect 4275 8317 4276 8321
rect 4278 8317 4279 8321
rect 4291 8317 4292 8321
rect 4294 8317 4297 8321
rect 4299 8317 4300 8321
rect 4312 8317 4313 8321
rect 4315 8317 4316 8321
rect 2503 8284 2504 8288
rect 2506 8284 2509 8288
rect 2511 8284 2512 8288
rect 2524 8284 2525 8288
rect 2527 8284 2528 8288
rect 2540 8284 2541 8288
rect 2543 8284 2546 8288
rect 2548 8284 2549 8288
rect 2566 8284 2567 8288
rect 2569 8284 2570 8288
rect 2582 8284 2583 8288
rect 2585 8284 2586 8288
rect 2598 8284 2599 8288
rect 2601 8284 2604 8288
rect 2606 8284 2607 8288
rect 2619 8284 2620 8288
rect 2622 8284 2623 8288
rect 3448 8284 3449 8288
rect 3451 8284 3454 8288
rect 3456 8284 3457 8288
rect 3469 8284 3470 8288
rect 3472 8284 3473 8288
rect 3485 8284 3486 8288
rect 3488 8284 3491 8288
rect 3493 8284 3494 8288
rect 3511 8284 3512 8288
rect 3514 8284 3515 8288
rect 3527 8284 3528 8288
rect 3530 8284 3531 8288
rect 3543 8284 3544 8288
rect 3546 8284 3549 8288
rect 3551 8284 3552 8288
rect 3564 8284 3565 8288
rect 3567 8284 3568 8288
rect 2627 8247 2628 8251
rect 2630 8247 2631 8251
rect 3034 8251 3035 8255
rect 3037 8251 3038 8255
rect 3058 8247 3061 8251
rect 3063 8247 3066 8251
rect 3068 8247 3069 8251
rect 3115 8251 3116 8255
rect 3118 8251 3119 8255
rect 3139 8247 3142 8251
rect 3144 8247 3147 8251
rect 3149 8247 3150 8251
rect 3088 8243 3089 8247
rect 3091 8243 3092 8247
rect 2510 8238 2511 8242
rect 2513 8238 2514 8242
rect 2860 8238 2861 8242
rect 2863 8238 2864 8242
rect 2876 8238 2877 8242
rect 2879 8238 2880 8242
rect 2892 8238 2893 8242
rect 2895 8238 2896 8242
rect 2911 8238 2916 8242
rect 2918 8238 2921 8242
rect 2923 8238 2924 8242
rect 2945 8238 2947 8242
rect 2949 8238 2950 8242
rect 2967 8238 2968 8242
rect 2970 8238 2971 8242
rect 2983 8238 2988 8242
rect 2990 8238 2993 8242
rect 2995 8238 2996 8242
rect 3010 8238 3011 8242
rect 3013 8238 3014 8242
rect 3169 8243 3170 8247
rect 3172 8243 3173 8247
rect 3572 8247 3573 8251
rect 3575 8247 3576 8251
rect 3979 8251 3980 8255
rect 3982 8251 3983 8255
rect 4003 8247 4006 8251
rect 4008 8247 4011 8251
rect 4013 8247 4014 8251
rect 4060 8251 4061 8255
rect 4063 8251 4064 8255
rect 4084 8247 4087 8251
rect 4089 8247 4092 8251
rect 4094 8247 4095 8251
rect 4033 8243 4034 8247
rect 4036 8243 4037 8247
rect 3455 8238 3456 8242
rect 3458 8238 3459 8242
rect 3805 8238 3806 8242
rect 3808 8238 3809 8242
rect 3821 8238 3822 8242
rect 3824 8238 3825 8242
rect 3837 8238 3838 8242
rect 3840 8238 3841 8242
rect 3856 8238 3861 8242
rect 3863 8238 3866 8242
rect 3868 8238 3869 8242
rect 3890 8238 3892 8242
rect 3894 8238 3895 8242
rect 3912 8238 3913 8242
rect 3915 8238 3916 8242
rect 3928 8238 3933 8242
rect 3935 8238 3938 8242
rect 3940 8238 3941 8242
rect 3955 8238 3956 8242
rect 3958 8238 3959 8242
rect 4114 8243 4115 8247
rect 4117 8243 4118 8247
rect 2860 8192 2861 8196
rect 2863 8192 2864 8196
rect 2876 8192 2877 8196
rect 2879 8192 2880 8196
rect 2892 8192 2893 8196
rect 2895 8192 2896 8196
rect 2911 8192 2916 8196
rect 2918 8192 2921 8196
rect 2923 8192 2924 8196
rect 2945 8192 2947 8196
rect 2949 8192 2950 8196
rect 2967 8192 2968 8196
rect 2970 8192 2971 8196
rect 2983 8192 2988 8196
rect 2990 8192 2993 8196
rect 2995 8192 2996 8196
rect 3010 8192 3011 8196
rect 3013 8192 3014 8196
rect 2494 8182 2495 8186
rect 2497 8182 2498 8186
rect 2510 8182 2511 8186
rect 2513 8182 2516 8186
rect 2518 8182 2519 8186
rect 2531 8182 2532 8186
rect 2534 8182 2535 8186
rect 2547 8182 2548 8186
rect 2550 8182 2551 8186
rect 2568 8182 2569 8186
rect 2571 8182 2574 8186
rect 2576 8182 2577 8186
rect 2589 8182 2590 8186
rect 2592 8182 2593 8186
rect 2605 8182 2606 8186
rect 2608 8182 2611 8186
rect 2613 8182 2614 8186
rect 3058 8191 3061 8195
rect 3063 8191 3066 8195
rect 3068 8191 3069 8195
rect 3139 8191 3142 8195
rect 3144 8191 3147 8195
rect 3149 8191 3150 8195
rect 3805 8192 3806 8196
rect 3808 8192 3809 8196
rect 3821 8192 3822 8196
rect 3824 8192 3825 8196
rect 3837 8192 3838 8196
rect 3840 8192 3841 8196
rect 3856 8192 3861 8196
rect 3863 8192 3866 8196
rect 3868 8192 3869 8196
rect 3890 8192 3892 8196
rect 3894 8192 3895 8196
rect 3912 8192 3913 8196
rect 3915 8192 3916 8196
rect 3928 8192 3933 8196
rect 3935 8192 3938 8196
rect 3940 8192 3941 8196
rect 3955 8192 3956 8196
rect 3958 8192 3959 8196
rect 3439 8182 3440 8186
rect 3442 8182 3443 8186
rect 3455 8182 3456 8186
rect 3458 8182 3461 8186
rect 3463 8182 3464 8186
rect 3476 8182 3477 8186
rect 3479 8182 3480 8186
rect 3492 8182 3493 8186
rect 3495 8182 3496 8186
rect 3513 8182 3514 8186
rect 3516 8182 3519 8186
rect 3521 8182 3522 8186
rect 3534 8182 3535 8186
rect 3537 8182 3538 8186
rect 3550 8182 3551 8186
rect 3553 8182 3556 8186
rect 3558 8182 3559 8186
rect 4003 8191 4006 8195
rect 4008 8191 4011 8195
rect 4013 8191 4014 8195
rect 4084 8191 4087 8195
rect 4089 8191 4092 8195
rect 4094 8191 4095 8195
rect 3058 8115 3061 8119
rect 3063 8115 3066 8119
rect 3068 8115 3069 8119
rect 3139 8119 3140 8123
rect 3142 8119 3143 8123
rect 3163 8115 3166 8119
rect 3168 8115 3171 8119
rect 3173 8115 3174 8119
rect 3088 8111 3089 8115
rect 3091 8111 3092 8115
rect 2860 8106 2861 8110
rect 2863 8106 2864 8110
rect 2876 8106 2877 8110
rect 2879 8106 2880 8110
rect 2892 8106 2893 8110
rect 2895 8106 2896 8110
rect 2911 8106 2916 8110
rect 2918 8106 2921 8110
rect 2923 8106 2924 8110
rect 2945 8106 2947 8110
rect 2949 8106 2950 8110
rect 2967 8106 2968 8110
rect 2970 8106 2971 8110
rect 2983 8106 2988 8110
rect 2990 8106 2993 8110
rect 2995 8106 2996 8110
rect 3010 8106 3011 8110
rect 3013 8106 3014 8110
rect 3193 8111 3194 8115
rect 3196 8111 3197 8115
rect 4003 8115 4006 8119
rect 4008 8115 4011 8119
rect 4013 8115 4014 8119
rect 4084 8119 4085 8123
rect 4087 8119 4088 8123
rect 4108 8115 4111 8119
rect 4113 8115 4116 8119
rect 4118 8115 4119 8119
rect 4033 8111 4034 8115
rect 4036 8111 4037 8115
rect 3805 8106 3806 8110
rect 3808 8106 3809 8110
rect 3821 8106 3822 8110
rect 3824 8106 3825 8110
rect 3837 8106 3838 8110
rect 3840 8106 3841 8110
rect 3856 8106 3861 8110
rect 3863 8106 3866 8110
rect 3868 8106 3869 8110
rect 3890 8106 3892 8110
rect 3894 8106 3895 8110
rect 3912 8106 3913 8110
rect 3915 8106 3916 8110
rect 3928 8106 3933 8110
rect 3935 8106 3938 8110
rect 3940 8106 3941 8110
rect 3955 8106 3956 8110
rect 3958 8106 3959 8110
rect 4138 8111 4139 8115
rect 4141 8111 4142 8115
rect 2860 8060 2861 8064
rect 2863 8060 2864 8064
rect 2876 8060 2877 8064
rect 2879 8060 2880 8064
rect 2892 8060 2893 8064
rect 2895 8060 2896 8064
rect 2911 8060 2916 8064
rect 2918 8060 2921 8064
rect 2923 8060 2924 8064
rect 2945 8060 2947 8064
rect 2949 8060 2950 8064
rect 2967 8060 2968 8064
rect 2970 8060 2971 8064
rect 2983 8060 2988 8064
rect 2990 8060 2993 8064
rect 2995 8060 2996 8064
rect 3010 8060 3011 8064
rect 3013 8060 3014 8064
rect 3058 8060 3061 8064
rect 3063 8060 3066 8064
rect 3068 8060 3069 8064
rect 3163 8060 3166 8064
rect 3168 8060 3171 8064
rect 3173 8060 3174 8064
rect 3805 8060 3806 8064
rect 3808 8060 3809 8064
rect 3821 8060 3822 8064
rect 3824 8060 3825 8064
rect 3837 8060 3838 8064
rect 3840 8060 3841 8064
rect 3856 8060 3861 8064
rect 3863 8060 3866 8064
rect 3868 8060 3869 8064
rect 3890 8060 3892 8064
rect 3894 8060 3895 8064
rect 3912 8060 3913 8064
rect 3915 8060 3916 8064
rect 3928 8060 3933 8064
rect 3935 8060 3938 8064
rect 3940 8060 3941 8064
rect 3955 8060 3956 8064
rect 3958 8060 3959 8064
rect 4003 8060 4006 8064
rect 4008 8060 4011 8064
rect 4013 8060 4014 8064
rect 4108 8060 4111 8064
rect 4113 8060 4116 8064
rect 4118 8060 4119 8064
rect 3058 7983 3061 7987
rect 3063 7983 3066 7987
rect 3068 7983 3069 7987
rect 3115 7987 3116 7991
rect 3118 7987 3119 7991
rect 3139 7983 3142 7987
rect 3144 7983 3147 7987
rect 3149 7983 3150 7987
rect 3205 7987 3206 7991
rect 3208 7987 3209 7991
rect 3229 7983 3232 7987
rect 3234 7983 3237 7987
rect 3239 7983 3240 7987
rect 3088 7979 3089 7983
rect 3091 7979 3092 7983
rect 2860 7974 2861 7978
rect 2863 7974 2864 7978
rect 2876 7974 2877 7978
rect 2879 7974 2880 7978
rect 2892 7974 2893 7978
rect 2895 7974 2896 7978
rect 2911 7974 2916 7978
rect 2918 7974 2921 7978
rect 2923 7974 2924 7978
rect 2945 7974 2947 7978
rect 2949 7974 2950 7978
rect 2967 7974 2968 7978
rect 2970 7974 2971 7978
rect 2983 7974 2988 7978
rect 2990 7974 2993 7978
rect 2995 7974 2996 7978
rect 3010 7974 3011 7978
rect 3013 7974 3014 7978
rect 3169 7979 3170 7983
rect 3172 7979 3173 7983
rect 3259 7979 3260 7983
rect 3262 7979 3263 7983
rect 4003 7983 4006 7987
rect 4008 7983 4011 7987
rect 4013 7983 4014 7987
rect 4060 7987 4061 7991
rect 4063 7987 4064 7991
rect 4084 7983 4087 7987
rect 4089 7983 4092 7987
rect 4094 7983 4095 7987
rect 4150 7987 4151 7991
rect 4153 7987 4154 7991
rect 4174 7983 4177 7987
rect 4179 7983 4182 7987
rect 4184 7983 4185 7987
rect 4033 7979 4034 7983
rect 4036 7979 4037 7983
rect 3805 7974 3806 7978
rect 3808 7974 3809 7978
rect 3821 7974 3822 7978
rect 3824 7974 3825 7978
rect 3837 7974 3838 7978
rect 3840 7974 3841 7978
rect 3856 7974 3861 7978
rect 3863 7974 3866 7978
rect 3868 7974 3869 7978
rect 3890 7974 3892 7978
rect 3894 7974 3895 7978
rect 3912 7974 3913 7978
rect 3915 7974 3916 7978
rect 3928 7974 3933 7978
rect 3935 7974 3938 7978
rect 3940 7974 3941 7978
rect 3955 7974 3956 7978
rect 3958 7974 3959 7978
rect 4114 7979 4115 7983
rect 4117 7979 4118 7983
rect 4204 7979 4205 7983
rect 4207 7979 4208 7983
rect 2860 7928 2861 7932
rect 2863 7928 2864 7932
rect 2876 7928 2877 7932
rect 2879 7928 2880 7932
rect 2892 7928 2893 7932
rect 2895 7928 2896 7932
rect 2911 7928 2916 7932
rect 2918 7928 2921 7932
rect 2923 7928 2924 7932
rect 2945 7928 2947 7932
rect 2949 7928 2950 7932
rect 2967 7928 2968 7932
rect 2970 7928 2971 7932
rect 2983 7928 2988 7932
rect 2990 7928 2993 7932
rect 2995 7928 2996 7932
rect 3010 7928 3011 7932
rect 3013 7928 3014 7932
rect 3058 7925 3061 7929
rect 3063 7925 3066 7929
rect 3068 7925 3069 7929
rect 3139 7925 3142 7929
rect 3144 7925 3147 7929
rect 3149 7925 3150 7929
rect 3229 7925 3232 7929
rect 3234 7925 3237 7929
rect 3239 7925 3240 7929
rect 3805 7928 3806 7932
rect 3808 7928 3809 7932
rect 3821 7928 3822 7932
rect 3824 7928 3825 7932
rect 3837 7928 3838 7932
rect 3840 7928 3841 7932
rect 3856 7928 3861 7932
rect 3863 7928 3866 7932
rect 3868 7928 3869 7932
rect 3890 7928 3892 7932
rect 3894 7928 3895 7932
rect 3912 7928 3913 7932
rect 3915 7928 3916 7932
rect 3928 7928 3933 7932
rect 3935 7928 3938 7932
rect 3940 7928 3941 7932
rect 3955 7928 3956 7932
rect 3958 7928 3959 7932
rect 4003 7925 4006 7929
rect 4008 7925 4011 7929
rect 4013 7925 4014 7929
rect 4084 7925 4087 7929
rect 4089 7925 4092 7929
rect 4094 7925 4095 7929
rect 4174 7925 4177 7929
rect 4179 7925 4182 7929
rect 4184 7925 4185 7929
rect 3058 7851 3061 7855
rect 3063 7851 3066 7855
rect 3068 7851 3069 7855
rect 3088 7847 3089 7851
rect 3091 7847 3092 7851
rect 2860 7842 2861 7846
rect 2863 7842 2864 7846
rect 2876 7842 2877 7846
rect 2879 7842 2880 7846
rect 2892 7842 2893 7846
rect 2895 7842 2896 7846
rect 2911 7842 2916 7846
rect 2918 7842 2921 7846
rect 2923 7842 2924 7846
rect 2945 7842 2947 7846
rect 2949 7842 2950 7846
rect 2967 7842 2968 7846
rect 2970 7842 2971 7846
rect 2983 7842 2988 7846
rect 2990 7842 2993 7846
rect 2995 7842 2996 7846
rect 3010 7842 3011 7846
rect 3013 7842 3014 7846
rect 4003 7851 4006 7855
rect 4008 7851 4011 7855
rect 4013 7851 4014 7855
rect 4033 7847 4034 7851
rect 4036 7847 4037 7851
rect 3805 7842 3806 7846
rect 3808 7842 3809 7846
rect 3821 7842 3822 7846
rect 3824 7842 3825 7846
rect 3837 7842 3838 7846
rect 3840 7842 3841 7846
rect 3856 7842 3861 7846
rect 3863 7842 3866 7846
rect 3868 7842 3869 7846
rect 3890 7842 3892 7846
rect 3894 7842 3895 7846
rect 3912 7842 3913 7846
rect 3915 7842 3916 7846
rect 3928 7842 3933 7846
rect 3935 7842 3938 7846
rect 3940 7842 3941 7846
rect 3955 7842 3956 7846
rect 3958 7842 3959 7846
rect 2860 7796 2861 7800
rect 2863 7796 2864 7800
rect 2876 7796 2877 7800
rect 2879 7796 2880 7800
rect 2892 7796 2893 7800
rect 2895 7796 2896 7800
rect 2911 7796 2916 7800
rect 2918 7796 2921 7800
rect 2923 7796 2924 7800
rect 2945 7796 2947 7800
rect 2949 7796 2950 7800
rect 2967 7796 2968 7800
rect 2970 7796 2971 7800
rect 2983 7796 2988 7800
rect 2990 7796 2993 7800
rect 2995 7796 2996 7800
rect 3010 7796 3011 7800
rect 3013 7796 3014 7800
rect 3094 7796 3095 7800
rect 3097 7796 3098 7800
rect 3102 7796 3108 7800
rect 3112 7796 3113 7800
rect 3115 7796 3116 7800
rect 3137 7796 3138 7800
rect 3140 7796 3141 7800
rect 3153 7796 3154 7800
rect 3156 7796 3157 7800
rect 3172 7796 3177 7800
rect 3179 7796 3182 7800
rect 3184 7796 3185 7800
rect 3206 7796 3208 7800
rect 3210 7796 3211 7800
rect 3228 7796 3229 7800
rect 3231 7796 3232 7800
rect 3244 7796 3249 7800
rect 3251 7796 3254 7800
rect 3256 7796 3257 7800
rect 3271 7796 3272 7800
rect 3274 7796 3275 7800
rect 2371 7782 2372 7786
rect 2374 7782 2377 7786
rect 2379 7782 2380 7786
rect 2392 7782 2393 7786
rect 2395 7782 2396 7786
rect 2408 7782 2409 7786
rect 2411 7782 2414 7786
rect 2416 7782 2417 7786
rect 2434 7782 2435 7786
rect 2437 7782 2438 7786
rect 2450 7782 2451 7786
rect 2453 7782 2454 7786
rect 2466 7782 2467 7786
rect 2469 7782 2472 7786
rect 2474 7782 2475 7786
rect 2487 7782 2488 7786
rect 2490 7782 2491 7786
rect 2503 7782 2504 7786
rect 2506 7782 2509 7786
rect 2511 7782 2512 7786
rect 2524 7782 2525 7786
rect 2527 7782 2528 7786
rect 2540 7782 2541 7786
rect 2543 7782 2546 7786
rect 2548 7782 2549 7786
rect 2566 7782 2567 7786
rect 2569 7782 2570 7786
rect 2582 7782 2583 7786
rect 2585 7782 2586 7786
rect 2598 7782 2599 7786
rect 2601 7782 2604 7786
rect 2606 7782 2607 7786
rect 2619 7782 2620 7786
rect 2622 7782 2623 7786
rect 2635 7782 2636 7786
rect 2638 7782 2641 7786
rect 2643 7782 2644 7786
rect 2656 7782 2657 7786
rect 2659 7782 2660 7786
rect 2672 7782 2673 7786
rect 2675 7782 2678 7786
rect 2680 7782 2681 7786
rect 2698 7782 2699 7786
rect 2701 7782 2702 7786
rect 2714 7782 2715 7786
rect 2717 7782 2718 7786
rect 2730 7782 2731 7786
rect 2733 7782 2736 7786
rect 2738 7782 2739 7786
rect 2751 7782 2752 7786
rect 2754 7782 2755 7786
rect 3058 7789 3061 7793
rect 3063 7789 3066 7793
rect 3068 7789 3069 7793
rect 3805 7796 3806 7800
rect 3808 7796 3809 7800
rect 3821 7796 3822 7800
rect 3824 7796 3825 7800
rect 3837 7796 3838 7800
rect 3840 7796 3841 7800
rect 3856 7796 3861 7800
rect 3863 7796 3866 7800
rect 3868 7796 3869 7800
rect 3890 7796 3892 7800
rect 3894 7796 3895 7800
rect 3912 7796 3913 7800
rect 3915 7796 3916 7800
rect 3928 7796 3933 7800
rect 3935 7796 3938 7800
rect 3940 7796 3941 7800
rect 3955 7796 3956 7800
rect 3958 7796 3959 7800
rect 4039 7796 4040 7800
rect 4042 7796 4043 7800
rect 4047 7796 4053 7800
rect 4057 7796 4058 7800
rect 4060 7796 4061 7800
rect 4082 7796 4083 7800
rect 4085 7796 4086 7800
rect 4098 7796 4099 7800
rect 4101 7796 4102 7800
rect 4117 7796 4122 7800
rect 4124 7796 4127 7800
rect 4129 7796 4130 7800
rect 4151 7796 4153 7800
rect 4155 7796 4156 7800
rect 4173 7796 4174 7800
rect 4176 7796 4177 7800
rect 4189 7796 4194 7800
rect 4196 7796 4199 7800
rect 4201 7796 4202 7800
rect 4216 7796 4217 7800
rect 4219 7796 4220 7800
rect 3316 7782 3317 7786
rect 3319 7782 3322 7786
rect 3324 7782 3325 7786
rect 3337 7782 3338 7786
rect 3340 7782 3341 7786
rect 3353 7782 3354 7786
rect 3356 7782 3359 7786
rect 3361 7782 3362 7786
rect 3379 7782 3380 7786
rect 3382 7782 3383 7786
rect 3395 7782 3396 7786
rect 3398 7782 3399 7786
rect 3411 7782 3412 7786
rect 3414 7782 3417 7786
rect 3419 7782 3420 7786
rect 3432 7782 3433 7786
rect 3435 7782 3436 7786
rect 3448 7782 3449 7786
rect 3451 7782 3454 7786
rect 3456 7782 3457 7786
rect 3469 7782 3470 7786
rect 3472 7782 3473 7786
rect 3485 7782 3486 7786
rect 3488 7782 3491 7786
rect 3493 7782 3494 7786
rect 3511 7782 3512 7786
rect 3514 7782 3515 7786
rect 3527 7782 3528 7786
rect 3530 7782 3531 7786
rect 3543 7782 3544 7786
rect 3546 7782 3549 7786
rect 3551 7782 3552 7786
rect 3564 7782 3565 7786
rect 3567 7782 3568 7786
rect 3580 7782 3581 7786
rect 3583 7782 3586 7786
rect 3588 7782 3589 7786
rect 3601 7782 3602 7786
rect 3604 7782 3605 7786
rect 3617 7782 3618 7786
rect 3620 7782 3623 7786
rect 3625 7782 3626 7786
rect 3643 7782 3644 7786
rect 3646 7782 3647 7786
rect 3659 7782 3660 7786
rect 3662 7782 3663 7786
rect 3675 7782 3676 7786
rect 3678 7782 3681 7786
rect 3683 7782 3684 7786
rect 3696 7782 3697 7786
rect 3699 7782 3700 7786
rect 4003 7789 4006 7793
rect 4008 7789 4011 7793
rect 4013 7789 4014 7793
rect 2486 7738 2487 7742
rect 2489 7738 2490 7742
rect 2510 7738 2511 7742
rect 2513 7738 2514 7742
rect 3284 7742 3288 7743
rect 3284 7739 3288 7740
rect 3431 7738 3432 7742
rect 3434 7738 3435 7742
rect 3455 7738 3456 7742
rect 3458 7738 3459 7742
rect 4229 7742 4233 7743
rect 4229 7739 4233 7740
rect 2506 7725 2507 7729
rect 2509 7725 2510 7729
rect 3451 7725 3452 7729
rect 3454 7725 3455 7729
rect 2498 7713 2502 7714
rect 2498 7710 2502 7711
rect 3443 7713 3447 7714
rect 3443 7710 3447 7711
rect 2486 7702 2487 7706
rect 2489 7702 2490 7706
rect 2510 7702 2511 7706
rect 2513 7702 2514 7706
rect 3431 7702 3432 7706
rect 3434 7702 3435 7706
rect 3455 7702 3456 7706
rect 3458 7702 3459 7706
rect 3154 7670 3155 7674
rect 3157 7670 3160 7674
rect 3162 7670 3163 7674
rect 3175 7670 3176 7674
rect 3178 7670 3179 7674
rect 3191 7670 3192 7674
rect 3194 7670 3197 7674
rect 3199 7670 3200 7674
rect 3217 7670 3218 7674
rect 3220 7670 3221 7674
rect 3233 7670 3234 7674
rect 3236 7670 3237 7674
rect 3249 7670 3250 7674
rect 3252 7670 3255 7674
rect 3257 7670 3258 7674
rect 3270 7670 3271 7674
rect 3273 7670 3274 7674
rect 4099 7670 4100 7674
rect 4102 7670 4105 7674
rect 4107 7670 4108 7674
rect 4120 7670 4121 7674
rect 4123 7670 4124 7674
rect 4136 7670 4137 7674
rect 4139 7670 4142 7674
rect 4144 7670 4145 7674
rect 4162 7670 4163 7674
rect 4165 7670 4166 7674
rect 4178 7670 4179 7674
rect 4181 7670 4182 7674
rect 4194 7670 4195 7674
rect 4197 7670 4200 7674
rect 4202 7670 4203 7674
rect 4215 7670 4216 7674
rect 4218 7670 4219 7674
rect 2371 7640 2372 7644
rect 2374 7640 2377 7644
rect 2379 7640 2380 7644
rect 2392 7640 2393 7644
rect 2395 7640 2396 7644
rect 2408 7640 2409 7644
rect 2411 7640 2414 7644
rect 2416 7640 2417 7644
rect 2434 7640 2435 7644
rect 2437 7640 2438 7644
rect 2450 7640 2451 7644
rect 2453 7640 2454 7644
rect 2466 7640 2467 7644
rect 2469 7640 2472 7644
rect 2474 7640 2475 7644
rect 2487 7640 2488 7644
rect 2490 7640 2491 7644
rect 2503 7640 2504 7644
rect 2506 7640 2509 7644
rect 2511 7640 2512 7644
rect 2524 7640 2525 7644
rect 2527 7640 2528 7644
rect 2540 7640 2541 7644
rect 2543 7640 2546 7644
rect 2548 7640 2549 7644
rect 2566 7640 2567 7644
rect 2569 7640 2570 7644
rect 2582 7640 2583 7644
rect 2585 7640 2586 7644
rect 2598 7640 2599 7644
rect 2601 7640 2604 7644
rect 2606 7640 2607 7644
rect 2619 7640 2620 7644
rect 2622 7640 2623 7644
rect 2635 7640 2636 7644
rect 2638 7640 2641 7644
rect 2643 7640 2644 7644
rect 2656 7640 2657 7644
rect 2659 7640 2660 7644
rect 2672 7640 2673 7644
rect 2675 7640 2678 7644
rect 2680 7640 2681 7644
rect 2698 7640 2699 7644
rect 2701 7640 2702 7644
rect 2714 7640 2715 7644
rect 2717 7640 2718 7644
rect 2730 7640 2731 7644
rect 2733 7640 2736 7644
rect 2738 7640 2739 7644
rect 2751 7640 2752 7644
rect 2754 7640 2755 7644
rect 3316 7640 3317 7644
rect 3319 7640 3322 7644
rect 3324 7640 3325 7644
rect 3337 7640 3338 7644
rect 3340 7640 3341 7644
rect 3353 7640 3354 7644
rect 3356 7640 3359 7644
rect 3361 7640 3362 7644
rect 3379 7640 3380 7644
rect 3382 7640 3383 7644
rect 3395 7640 3396 7644
rect 3398 7640 3399 7644
rect 3411 7640 3412 7644
rect 3414 7640 3417 7644
rect 3419 7640 3420 7644
rect 3432 7640 3433 7644
rect 3435 7640 3436 7644
rect 3448 7640 3449 7644
rect 3451 7640 3454 7644
rect 3456 7640 3457 7644
rect 3469 7640 3470 7644
rect 3472 7640 3473 7644
rect 3485 7640 3486 7644
rect 3488 7640 3491 7644
rect 3493 7640 3494 7644
rect 3511 7640 3512 7644
rect 3514 7640 3515 7644
rect 3527 7640 3528 7644
rect 3530 7640 3531 7644
rect 3543 7640 3544 7644
rect 3546 7640 3549 7644
rect 3551 7640 3552 7644
rect 3564 7640 3565 7644
rect 3567 7640 3568 7644
rect 3580 7640 3581 7644
rect 3583 7640 3586 7644
rect 3588 7640 3589 7644
rect 3601 7640 3602 7644
rect 3604 7640 3605 7644
rect 3617 7640 3618 7644
rect 3620 7640 3623 7644
rect 3625 7640 3626 7644
rect 3643 7640 3644 7644
rect 3646 7640 3647 7644
rect 3659 7640 3660 7644
rect 3662 7640 3663 7644
rect 3675 7640 3676 7644
rect 3678 7640 3681 7644
rect 3683 7640 3684 7644
rect 3696 7640 3697 7644
rect 3699 7640 3700 7644
rect 3296 7596 3300 7597
rect 3296 7593 3300 7594
rect 4241 7596 4245 7597
rect 4241 7593 4245 7594
rect 3154 7584 3155 7588
rect 3157 7584 3160 7588
rect 3162 7584 3163 7588
rect 3175 7584 3176 7588
rect 3178 7584 3179 7588
rect 3191 7584 3192 7588
rect 3194 7584 3197 7588
rect 3199 7584 3200 7588
rect 3217 7584 3218 7588
rect 3220 7584 3221 7588
rect 3233 7584 3234 7588
rect 3236 7584 3237 7588
rect 3249 7584 3250 7588
rect 3252 7584 3255 7588
rect 3257 7584 3258 7588
rect 3270 7584 3271 7588
rect 3273 7584 3274 7588
rect 4099 7584 4100 7588
rect 4102 7584 4105 7588
rect 4107 7584 4108 7588
rect 4120 7584 4121 7588
rect 4123 7584 4124 7588
rect 4136 7584 4137 7588
rect 4139 7584 4142 7588
rect 4144 7584 4145 7588
rect 4162 7584 4163 7588
rect 4165 7584 4166 7588
rect 4178 7584 4179 7588
rect 4181 7584 4182 7588
rect 4194 7584 4195 7588
rect 4197 7584 4200 7588
rect 4202 7584 4203 7588
rect 4215 7584 4216 7588
rect 4218 7584 4219 7588
rect 2371 7554 2372 7558
rect 2374 7554 2377 7558
rect 2379 7554 2380 7558
rect 2392 7554 2393 7558
rect 2395 7554 2396 7558
rect 2408 7554 2409 7558
rect 2411 7554 2414 7558
rect 2416 7554 2417 7558
rect 2434 7554 2435 7558
rect 2437 7554 2438 7558
rect 2450 7554 2451 7558
rect 2453 7554 2454 7558
rect 2466 7554 2467 7558
rect 2469 7554 2472 7558
rect 2474 7554 2475 7558
rect 2487 7554 2488 7558
rect 2490 7554 2491 7558
rect 2503 7554 2504 7558
rect 2506 7554 2509 7558
rect 2511 7554 2512 7558
rect 2524 7554 2525 7558
rect 2527 7554 2528 7558
rect 2540 7554 2541 7558
rect 2543 7554 2546 7558
rect 2548 7554 2549 7558
rect 2566 7554 2567 7558
rect 2569 7554 2570 7558
rect 2582 7554 2583 7558
rect 2585 7554 2586 7558
rect 2598 7554 2599 7558
rect 2601 7554 2604 7558
rect 2606 7554 2607 7558
rect 2619 7554 2620 7558
rect 2622 7554 2623 7558
rect 2635 7554 2636 7558
rect 2638 7554 2641 7558
rect 2643 7554 2644 7558
rect 2656 7554 2657 7558
rect 2659 7554 2660 7558
rect 2672 7554 2673 7558
rect 2675 7554 2678 7558
rect 2680 7554 2681 7558
rect 2698 7554 2699 7558
rect 2701 7554 2702 7558
rect 2714 7554 2715 7558
rect 2717 7554 2718 7558
rect 2730 7554 2731 7558
rect 2733 7554 2736 7558
rect 2738 7554 2739 7558
rect 2751 7554 2752 7558
rect 2754 7554 2755 7558
rect 3316 7554 3317 7558
rect 3319 7554 3322 7558
rect 3324 7554 3325 7558
rect 3337 7554 3338 7558
rect 3340 7554 3341 7558
rect 3353 7554 3354 7558
rect 3356 7554 3359 7558
rect 3361 7554 3362 7558
rect 3379 7554 3380 7558
rect 3382 7554 3383 7558
rect 3395 7554 3396 7558
rect 3398 7554 3399 7558
rect 3411 7554 3412 7558
rect 3414 7554 3417 7558
rect 3419 7554 3420 7558
rect 3432 7554 3433 7558
rect 3435 7554 3436 7558
rect 3448 7554 3449 7558
rect 3451 7554 3454 7558
rect 3456 7554 3457 7558
rect 3469 7554 3470 7558
rect 3472 7554 3473 7558
rect 3485 7554 3486 7558
rect 3488 7554 3491 7558
rect 3493 7554 3494 7558
rect 3511 7554 3512 7558
rect 3514 7554 3515 7558
rect 3527 7554 3528 7558
rect 3530 7554 3531 7558
rect 3543 7554 3544 7558
rect 3546 7554 3549 7558
rect 3551 7554 3552 7558
rect 3564 7554 3565 7558
rect 3567 7554 3568 7558
rect 3580 7554 3581 7558
rect 3583 7554 3586 7558
rect 3588 7554 3589 7558
rect 3601 7554 3602 7558
rect 3604 7554 3605 7558
rect 3617 7554 3618 7558
rect 3620 7554 3623 7558
rect 3625 7554 3626 7558
rect 3643 7554 3644 7558
rect 3646 7554 3647 7558
rect 3659 7554 3660 7558
rect 3662 7554 3663 7558
rect 3675 7554 3676 7558
rect 3678 7554 3681 7558
rect 3683 7554 3684 7558
rect 3696 7554 3697 7558
rect 3699 7554 3700 7558
rect 2603 7510 2604 7514
rect 2606 7510 2607 7514
rect 2627 7510 2628 7514
rect 2630 7510 2631 7514
rect 3548 7510 3549 7514
rect 3551 7510 3552 7514
rect 3572 7510 3573 7514
rect 3575 7510 3576 7514
rect 2623 7499 2624 7503
rect 2626 7499 2627 7503
rect 3568 7499 3569 7503
rect 3571 7499 3572 7503
rect 2615 7487 2619 7488
rect 2615 7484 2619 7485
rect 3560 7487 3564 7488
rect 3560 7484 3564 7485
rect 2603 7476 2604 7480
rect 2606 7476 2607 7480
rect 2627 7476 2628 7480
rect 2630 7476 2631 7480
rect 3548 7476 3549 7480
rect 3551 7476 3552 7480
rect 3572 7476 3573 7480
rect 3575 7476 3576 7480
rect 2371 7414 2372 7418
rect 2374 7414 2377 7418
rect 2379 7414 2380 7418
rect 2392 7414 2393 7418
rect 2395 7414 2396 7418
rect 2408 7414 2409 7418
rect 2411 7414 2414 7418
rect 2416 7414 2417 7418
rect 2434 7414 2435 7418
rect 2437 7414 2438 7418
rect 2450 7414 2451 7418
rect 2453 7414 2454 7418
rect 2466 7414 2467 7418
rect 2469 7414 2472 7418
rect 2474 7414 2475 7418
rect 2487 7414 2488 7418
rect 2490 7414 2491 7418
rect 2503 7414 2504 7418
rect 2506 7414 2509 7418
rect 2511 7414 2512 7418
rect 2524 7414 2525 7418
rect 2527 7414 2528 7418
rect 2540 7414 2541 7418
rect 2543 7414 2546 7418
rect 2548 7414 2549 7418
rect 2566 7414 2567 7418
rect 2569 7414 2570 7418
rect 2582 7414 2583 7418
rect 2585 7414 2586 7418
rect 2598 7414 2599 7418
rect 2601 7414 2604 7418
rect 2606 7414 2607 7418
rect 2619 7414 2620 7418
rect 2622 7414 2623 7418
rect 2635 7414 2636 7418
rect 2638 7414 2641 7418
rect 2643 7414 2644 7418
rect 2656 7414 2657 7418
rect 2659 7414 2660 7418
rect 2672 7414 2673 7418
rect 2675 7414 2678 7418
rect 2680 7414 2681 7418
rect 2698 7414 2699 7418
rect 2701 7414 2702 7418
rect 2714 7414 2715 7418
rect 2717 7414 2718 7418
rect 2730 7414 2731 7418
rect 2733 7414 2736 7418
rect 2738 7414 2739 7418
rect 2751 7414 2752 7418
rect 2754 7414 2755 7418
rect 3316 7414 3317 7418
rect 3319 7414 3322 7418
rect 3324 7414 3325 7418
rect 3337 7414 3338 7418
rect 3340 7414 3341 7418
rect 3353 7414 3354 7418
rect 3356 7414 3359 7418
rect 3361 7414 3362 7418
rect 3379 7414 3380 7418
rect 3382 7414 3383 7418
rect 3395 7414 3396 7418
rect 3398 7414 3399 7418
rect 3411 7414 3412 7418
rect 3414 7414 3417 7418
rect 3419 7414 3420 7418
rect 3432 7414 3433 7418
rect 3435 7414 3436 7418
rect 3448 7414 3449 7418
rect 3451 7414 3454 7418
rect 3456 7414 3457 7418
rect 3469 7414 3470 7418
rect 3472 7414 3473 7418
rect 3485 7414 3486 7418
rect 3488 7414 3491 7418
rect 3493 7414 3494 7418
rect 3511 7414 3512 7418
rect 3514 7414 3515 7418
rect 3527 7414 3528 7418
rect 3530 7414 3531 7418
rect 3543 7414 3544 7418
rect 3546 7414 3549 7418
rect 3551 7414 3552 7418
rect 3564 7414 3565 7418
rect 3567 7414 3568 7418
rect 3580 7414 3581 7418
rect 3583 7414 3586 7418
rect 3588 7414 3589 7418
rect 3601 7414 3602 7418
rect 3604 7414 3605 7418
rect 3617 7414 3618 7418
rect 3620 7414 3623 7418
rect 3625 7414 3626 7418
rect 3643 7414 3644 7418
rect 3646 7414 3647 7418
rect 3659 7414 3660 7418
rect 3662 7414 3663 7418
rect 3675 7414 3676 7418
rect 3678 7414 3681 7418
rect 3683 7414 3684 7418
rect 3696 7414 3697 7418
rect 3699 7414 3700 7418
rect 4578 7986 4579 8015
rect 4574 7982 4579 7986
rect 4578 7975 4579 7982
rect 4581 7975 4582 8015
rect 4586 7975 4587 8015
rect 4589 7986 4590 8015
rect 4594 7986 4595 8015
rect 4589 7982 4595 7986
rect 4589 7975 4590 7982
rect 4594 7975 4595 7982
rect 4597 7975 4598 8015
rect 4602 7975 4603 8015
rect 4605 7986 4606 8015
rect 4610 7986 4611 8015
rect 4605 7982 4611 7986
rect 4605 7975 4606 7982
rect 4610 7975 4611 7982
rect 4613 7975 4614 8015
rect 4618 7975 4619 8015
rect 4621 7986 4622 8015
rect 4626 7986 4627 8015
rect 4621 7982 4627 7986
rect 4621 7975 4622 7982
rect 4626 7975 4627 7982
rect 4631 7975 4634 8034
rect 4636 7975 4637 8034
rect 4641 7975 4642 8034
rect 4644 7986 4645 8034
rect 4649 7986 4650 8034
rect 4644 7982 4650 7986
rect 4644 7975 4645 7982
rect 4649 7975 4650 7982
rect 4652 7975 4653 8034
rect 4657 7975 4658 8034
rect 4660 7986 4661 8034
rect 4665 7986 4666 8034
rect 4660 7982 4666 7986
rect 4660 7975 4661 7982
rect 4665 7975 4666 7982
rect 4670 7975 4677 8034
rect 4679 7975 4680 8034
rect 4684 7975 4685 8034
rect 4687 7986 4688 8034
rect 4692 7986 4693 8034
rect 4687 7975 4693 7986
rect 4695 7975 4696 8034
rect 4700 7975 4701 8034
rect 4703 7986 4704 8034
rect 4708 7986 4709 8034
rect 4703 7982 4709 7986
rect 4703 7975 4704 7982
rect 4708 7975 4709 7982
rect 4713 7975 4718 8034
rect 4720 7975 4721 8034
rect 4725 7975 4726 8034
rect 4728 7986 4729 8034
rect 4733 7986 4734 8034
rect 4728 7975 4734 7986
rect 4736 7975 4737 8034
rect 4741 7975 4742 8034
rect 4744 7986 4745 8034
rect 4749 7986 4750 8034
rect 4744 7982 4750 7986
rect 4744 7975 4745 7982
rect 4749 7975 4750 7982
<< pdiffusion >>
rect 1556 9949 1562 9953
rect 1566 9949 1572 9953
rect 1576 9949 1582 9953
rect 1586 9949 1592 9953
rect 1596 9949 1601 9953
rect 1556 9948 1601 9949
rect 1556 9944 1557 9948
rect 1561 9944 1567 9948
rect 1571 9944 1577 9948
rect 1581 9944 1587 9948
rect 1591 9944 1597 9948
rect 1556 9943 1601 9944
rect 1556 9939 1562 9943
rect 1566 9939 1572 9943
rect 1576 9939 1582 9943
rect 1586 9939 1592 9943
rect 1596 9939 1601 9943
rect 1556 9938 1601 9939
rect 1556 9934 1557 9938
rect 1561 9934 1567 9938
rect 1571 9934 1577 9938
rect 1581 9934 1587 9938
rect 1591 9934 1597 9938
rect 1556 9933 1601 9934
rect 1556 9929 1562 9933
rect 1566 9929 1572 9933
rect 1576 9929 1582 9933
rect 1586 9929 1592 9933
rect 1596 9929 1601 9933
rect 1556 9928 1601 9929
rect 1556 9924 1557 9928
rect 1561 9924 1567 9928
rect 1571 9924 1577 9928
rect 1581 9924 1587 9928
rect 1591 9924 1597 9928
rect 1556 9923 1601 9924
rect 1556 9919 1562 9923
rect 1566 9919 1572 9923
rect 1576 9919 1582 9923
rect 1586 9919 1592 9923
rect 1596 9919 1601 9923
rect 1556 9918 1601 9919
rect 1556 9914 1557 9918
rect 1561 9914 1567 9918
rect 1571 9914 1577 9918
rect 1581 9914 1587 9918
rect 1591 9914 1597 9918
rect 1556 9913 1601 9914
rect 1556 9909 1562 9913
rect 1566 9909 1572 9913
rect 1576 9909 1582 9913
rect 1586 9909 1592 9913
rect 1596 9909 1601 9913
rect 1556 9908 1601 9909
rect 1556 9904 1557 9908
rect 1561 9904 1567 9908
rect 1571 9904 1577 9908
rect 1581 9904 1587 9908
rect 1591 9904 1597 9908
rect 1556 9903 1601 9904
rect 1556 9899 1562 9903
rect 1566 9899 1572 9903
rect 1576 9899 1582 9903
rect 1586 9899 1592 9903
rect 1596 9899 1601 9903
rect 1556 9898 1601 9899
rect 1556 9894 1557 9898
rect 1561 9894 1567 9898
rect 1571 9894 1577 9898
rect 1581 9894 1587 9898
rect 1591 9894 1597 9898
rect 1556 9893 1601 9894
rect 1556 9889 1562 9893
rect 1566 9889 1572 9893
rect 1576 9889 1582 9893
rect 1586 9889 1592 9893
rect 1596 9889 1601 9893
rect 1556 9888 1601 9889
rect 1556 9884 1557 9888
rect 1561 9884 1567 9888
rect 1571 9884 1577 9888
rect 1581 9884 1587 9888
rect 1591 9884 1597 9888
rect 1556 9883 1601 9884
rect 1556 9879 1562 9883
rect 1566 9879 1572 9883
rect 1576 9879 1582 9883
rect 1586 9879 1592 9883
rect 1596 9879 1601 9883
rect 1556 9878 1601 9879
rect 1556 9874 1557 9878
rect 1561 9874 1567 9878
rect 1571 9874 1577 9878
rect 1581 9874 1587 9878
rect 1591 9874 1597 9878
rect 1556 9873 1601 9874
rect 1556 9869 1562 9873
rect 1566 9869 1572 9873
rect 1576 9869 1582 9873
rect 1586 9869 1592 9873
rect 1596 9869 1601 9873
rect 1556 9868 1601 9869
rect 1556 9864 1557 9868
rect 1561 9864 1567 9868
rect 1571 9864 1577 9868
rect 1581 9864 1587 9868
rect 1591 9864 1597 9868
rect 1865 9949 1871 9953
rect 1875 9949 1881 9953
rect 1885 9949 1891 9953
rect 1895 9949 1901 9953
rect 1905 9949 1910 9953
rect 1865 9948 1910 9949
rect 1865 9944 1866 9948
rect 1870 9944 1876 9948
rect 1880 9944 1886 9948
rect 1890 9944 1896 9948
rect 1900 9944 1906 9948
rect 1865 9943 1910 9944
rect 1865 9939 1871 9943
rect 1875 9939 1881 9943
rect 1885 9939 1891 9943
rect 1895 9939 1901 9943
rect 1905 9939 1910 9943
rect 1865 9938 1910 9939
rect 1865 9934 1866 9938
rect 1870 9934 1876 9938
rect 1880 9934 1886 9938
rect 1890 9934 1896 9938
rect 1900 9934 1906 9938
rect 1865 9933 1910 9934
rect 1865 9929 1871 9933
rect 1875 9929 1881 9933
rect 1885 9929 1891 9933
rect 1895 9929 1901 9933
rect 1905 9929 1910 9933
rect 1865 9928 1910 9929
rect 1865 9924 1866 9928
rect 1870 9924 1876 9928
rect 1880 9924 1886 9928
rect 1890 9924 1896 9928
rect 1900 9924 1906 9928
rect 1865 9923 1910 9924
rect 1865 9919 1871 9923
rect 1875 9919 1881 9923
rect 1885 9919 1891 9923
rect 1895 9919 1901 9923
rect 1905 9919 1910 9923
rect 1865 9918 1910 9919
rect 1865 9914 1866 9918
rect 1870 9914 1876 9918
rect 1880 9914 1886 9918
rect 1890 9914 1896 9918
rect 1900 9914 1906 9918
rect 1865 9913 1910 9914
rect 1865 9909 1871 9913
rect 1875 9909 1881 9913
rect 1885 9909 1891 9913
rect 1895 9909 1901 9913
rect 1905 9909 1910 9913
rect 1865 9908 1910 9909
rect 1865 9904 1866 9908
rect 1870 9904 1876 9908
rect 1880 9904 1886 9908
rect 1890 9904 1896 9908
rect 1900 9904 1906 9908
rect 1865 9903 1910 9904
rect 1865 9899 1871 9903
rect 1875 9899 1881 9903
rect 1885 9899 1891 9903
rect 1895 9899 1901 9903
rect 1905 9899 1910 9903
rect 1865 9898 1910 9899
rect 1865 9894 1866 9898
rect 1870 9894 1876 9898
rect 1880 9894 1886 9898
rect 1890 9894 1896 9898
rect 1900 9894 1906 9898
rect 1865 9893 1910 9894
rect 1865 9889 1871 9893
rect 1875 9889 1881 9893
rect 1885 9889 1891 9893
rect 1895 9889 1901 9893
rect 1905 9889 1910 9893
rect 1865 9888 1910 9889
rect 1865 9884 1866 9888
rect 1870 9884 1876 9888
rect 1880 9884 1886 9888
rect 1890 9884 1896 9888
rect 1900 9884 1906 9888
rect 1865 9883 1910 9884
rect 1865 9879 1871 9883
rect 1875 9879 1881 9883
rect 1885 9879 1891 9883
rect 1895 9879 1901 9883
rect 1905 9879 1910 9883
rect 1865 9878 1910 9879
rect 1865 9874 1866 9878
rect 1870 9874 1876 9878
rect 1880 9874 1886 9878
rect 1890 9874 1896 9878
rect 1900 9874 1906 9878
rect 1865 9873 1910 9874
rect 1865 9869 1871 9873
rect 1875 9869 1881 9873
rect 1885 9869 1891 9873
rect 1895 9869 1901 9873
rect 1905 9869 1910 9873
rect 1865 9868 1910 9869
rect 1865 9864 1866 9868
rect 1870 9864 1876 9868
rect 1880 9864 1886 9868
rect 1890 9864 1896 9868
rect 1900 9864 1906 9868
rect 2174 9949 2180 9953
rect 2184 9949 2190 9953
rect 2194 9949 2200 9953
rect 2204 9949 2210 9953
rect 2214 9949 2219 9953
rect 2174 9948 2219 9949
rect 2174 9944 2175 9948
rect 2179 9944 2185 9948
rect 2189 9944 2195 9948
rect 2199 9944 2205 9948
rect 2209 9944 2215 9948
rect 2174 9943 2219 9944
rect 2174 9939 2180 9943
rect 2184 9939 2190 9943
rect 2194 9939 2200 9943
rect 2204 9939 2210 9943
rect 2214 9939 2219 9943
rect 2174 9938 2219 9939
rect 2174 9934 2175 9938
rect 2179 9934 2185 9938
rect 2189 9934 2195 9938
rect 2199 9934 2205 9938
rect 2209 9934 2215 9938
rect 2174 9933 2219 9934
rect 2174 9929 2180 9933
rect 2184 9929 2190 9933
rect 2194 9929 2200 9933
rect 2204 9929 2210 9933
rect 2214 9929 2219 9933
rect 2174 9928 2219 9929
rect 2174 9924 2175 9928
rect 2179 9924 2185 9928
rect 2189 9924 2195 9928
rect 2199 9924 2205 9928
rect 2209 9924 2215 9928
rect 2174 9923 2219 9924
rect 2174 9919 2180 9923
rect 2184 9919 2190 9923
rect 2194 9919 2200 9923
rect 2204 9919 2210 9923
rect 2214 9919 2219 9923
rect 2174 9918 2219 9919
rect 2174 9914 2175 9918
rect 2179 9914 2185 9918
rect 2189 9914 2195 9918
rect 2199 9914 2205 9918
rect 2209 9914 2215 9918
rect 2174 9913 2219 9914
rect 2174 9909 2180 9913
rect 2184 9909 2190 9913
rect 2194 9909 2200 9913
rect 2204 9909 2210 9913
rect 2214 9909 2219 9913
rect 2174 9908 2219 9909
rect 2174 9904 2175 9908
rect 2179 9904 2185 9908
rect 2189 9904 2195 9908
rect 2199 9904 2205 9908
rect 2209 9904 2215 9908
rect 2174 9903 2219 9904
rect 2174 9899 2180 9903
rect 2184 9899 2190 9903
rect 2194 9899 2200 9903
rect 2204 9899 2210 9903
rect 2214 9899 2219 9903
rect 2174 9898 2219 9899
rect 2174 9894 2175 9898
rect 2179 9894 2185 9898
rect 2189 9894 2195 9898
rect 2199 9894 2205 9898
rect 2209 9894 2215 9898
rect 2174 9893 2219 9894
rect 2174 9889 2180 9893
rect 2184 9889 2190 9893
rect 2194 9889 2200 9893
rect 2204 9889 2210 9893
rect 2214 9889 2219 9893
rect 2174 9888 2219 9889
rect 2174 9884 2175 9888
rect 2179 9884 2185 9888
rect 2189 9884 2195 9888
rect 2199 9884 2205 9888
rect 2209 9884 2215 9888
rect 2174 9883 2219 9884
rect 2174 9879 2180 9883
rect 2184 9879 2190 9883
rect 2194 9879 2200 9883
rect 2204 9879 2210 9883
rect 2214 9879 2219 9883
rect 2174 9878 2219 9879
rect 2174 9874 2175 9878
rect 2179 9874 2185 9878
rect 2189 9874 2195 9878
rect 2199 9874 2205 9878
rect 2209 9874 2215 9878
rect 2174 9873 2219 9874
rect 2174 9869 2180 9873
rect 2184 9869 2190 9873
rect 2194 9869 2200 9873
rect 2204 9869 2210 9873
rect 2214 9869 2219 9873
rect 2174 9868 2219 9869
rect 2174 9864 2175 9868
rect 2179 9864 2185 9868
rect 2189 9864 2195 9868
rect 2199 9864 2205 9868
rect 2209 9864 2215 9868
rect 2483 9949 2489 9953
rect 2493 9949 2499 9953
rect 2503 9949 2509 9953
rect 2513 9949 2519 9953
rect 2523 9949 2528 9953
rect 2483 9948 2528 9949
rect 2483 9944 2484 9948
rect 2488 9944 2494 9948
rect 2498 9944 2504 9948
rect 2508 9944 2514 9948
rect 2518 9944 2524 9948
rect 2483 9943 2528 9944
rect 2483 9939 2489 9943
rect 2493 9939 2499 9943
rect 2503 9939 2509 9943
rect 2513 9939 2519 9943
rect 2523 9939 2528 9943
rect 2483 9938 2528 9939
rect 2483 9934 2484 9938
rect 2488 9934 2494 9938
rect 2498 9934 2504 9938
rect 2508 9934 2514 9938
rect 2518 9934 2524 9938
rect 2483 9933 2528 9934
rect 2483 9929 2489 9933
rect 2493 9929 2499 9933
rect 2503 9929 2509 9933
rect 2513 9929 2519 9933
rect 2523 9929 2528 9933
rect 2483 9928 2528 9929
rect 2483 9924 2484 9928
rect 2488 9924 2494 9928
rect 2498 9924 2504 9928
rect 2508 9924 2514 9928
rect 2518 9924 2524 9928
rect 2483 9923 2528 9924
rect 2483 9919 2489 9923
rect 2493 9919 2499 9923
rect 2503 9919 2509 9923
rect 2513 9919 2519 9923
rect 2523 9919 2528 9923
rect 2483 9918 2528 9919
rect 2483 9914 2484 9918
rect 2488 9914 2494 9918
rect 2498 9914 2504 9918
rect 2508 9914 2514 9918
rect 2518 9914 2524 9918
rect 2483 9913 2528 9914
rect 2483 9909 2489 9913
rect 2493 9909 2499 9913
rect 2503 9909 2509 9913
rect 2513 9909 2519 9913
rect 2523 9909 2528 9913
rect 2483 9908 2528 9909
rect 2483 9904 2484 9908
rect 2488 9904 2494 9908
rect 2498 9904 2504 9908
rect 2508 9904 2514 9908
rect 2518 9904 2524 9908
rect 2483 9903 2528 9904
rect 2483 9899 2489 9903
rect 2493 9899 2499 9903
rect 2503 9899 2509 9903
rect 2513 9899 2519 9903
rect 2523 9899 2528 9903
rect 2483 9898 2528 9899
rect 2483 9894 2484 9898
rect 2488 9894 2494 9898
rect 2498 9894 2504 9898
rect 2508 9894 2514 9898
rect 2518 9894 2524 9898
rect 2483 9893 2528 9894
rect 2483 9889 2489 9893
rect 2493 9889 2499 9893
rect 2503 9889 2509 9893
rect 2513 9889 2519 9893
rect 2523 9889 2528 9893
rect 2483 9888 2528 9889
rect 2483 9884 2484 9888
rect 2488 9884 2494 9888
rect 2498 9884 2504 9888
rect 2508 9884 2514 9888
rect 2518 9884 2524 9888
rect 2483 9883 2528 9884
rect 2483 9879 2489 9883
rect 2493 9879 2499 9883
rect 2503 9879 2509 9883
rect 2513 9879 2519 9883
rect 2523 9879 2528 9883
rect 2483 9878 2528 9879
rect 2483 9874 2484 9878
rect 2488 9874 2494 9878
rect 2498 9874 2504 9878
rect 2508 9874 2514 9878
rect 2518 9874 2524 9878
rect 2483 9873 2528 9874
rect 2483 9869 2489 9873
rect 2493 9869 2499 9873
rect 2503 9869 2509 9873
rect 2513 9869 2519 9873
rect 2523 9869 2528 9873
rect 2483 9868 2528 9869
rect 2483 9864 2484 9868
rect 2488 9864 2494 9868
rect 2498 9864 2504 9868
rect 2508 9864 2514 9868
rect 2518 9864 2524 9868
rect 2792 9949 2798 9953
rect 2802 9949 2808 9953
rect 2812 9949 2818 9953
rect 2822 9949 2828 9953
rect 2832 9949 2837 9953
rect 2792 9948 2837 9949
rect 2792 9944 2793 9948
rect 2797 9944 2803 9948
rect 2807 9944 2813 9948
rect 2817 9944 2823 9948
rect 2827 9944 2833 9948
rect 2792 9943 2837 9944
rect 2792 9939 2798 9943
rect 2802 9939 2808 9943
rect 2812 9939 2818 9943
rect 2822 9939 2828 9943
rect 2832 9939 2837 9943
rect 2792 9938 2837 9939
rect 2792 9934 2793 9938
rect 2797 9934 2803 9938
rect 2807 9934 2813 9938
rect 2817 9934 2823 9938
rect 2827 9934 2833 9938
rect 2792 9933 2837 9934
rect 2792 9929 2798 9933
rect 2802 9929 2808 9933
rect 2812 9929 2818 9933
rect 2822 9929 2828 9933
rect 2832 9929 2837 9933
rect 2792 9928 2837 9929
rect 2792 9924 2793 9928
rect 2797 9924 2803 9928
rect 2807 9924 2813 9928
rect 2817 9924 2823 9928
rect 2827 9924 2833 9928
rect 2792 9923 2837 9924
rect 2792 9919 2798 9923
rect 2802 9919 2808 9923
rect 2812 9919 2818 9923
rect 2822 9919 2828 9923
rect 2832 9919 2837 9923
rect 2792 9918 2837 9919
rect 2792 9914 2793 9918
rect 2797 9914 2803 9918
rect 2807 9914 2813 9918
rect 2817 9914 2823 9918
rect 2827 9914 2833 9918
rect 2792 9913 2837 9914
rect 2792 9909 2798 9913
rect 2802 9909 2808 9913
rect 2812 9909 2818 9913
rect 2822 9909 2828 9913
rect 2832 9909 2837 9913
rect 2792 9908 2837 9909
rect 2792 9904 2793 9908
rect 2797 9904 2803 9908
rect 2807 9904 2813 9908
rect 2817 9904 2823 9908
rect 2827 9904 2833 9908
rect 2792 9903 2837 9904
rect 2792 9899 2798 9903
rect 2802 9899 2808 9903
rect 2812 9899 2818 9903
rect 2822 9899 2828 9903
rect 2832 9899 2837 9903
rect 2792 9898 2837 9899
rect 2792 9894 2793 9898
rect 2797 9894 2803 9898
rect 2807 9894 2813 9898
rect 2817 9894 2823 9898
rect 2827 9894 2833 9898
rect 2792 9893 2837 9894
rect 2792 9889 2798 9893
rect 2802 9889 2808 9893
rect 2812 9889 2818 9893
rect 2822 9889 2828 9893
rect 2832 9889 2837 9893
rect 2792 9888 2837 9889
rect 2792 9884 2793 9888
rect 2797 9884 2803 9888
rect 2807 9884 2813 9888
rect 2817 9884 2823 9888
rect 2827 9884 2833 9888
rect 2792 9883 2837 9884
rect 2792 9879 2798 9883
rect 2802 9879 2808 9883
rect 2812 9879 2818 9883
rect 2822 9879 2828 9883
rect 2832 9879 2837 9883
rect 2792 9878 2837 9879
rect 2792 9874 2793 9878
rect 2797 9874 2803 9878
rect 2807 9874 2813 9878
rect 2817 9874 2823 9878
rect 2827 9874 2833 9878
rect 2792 9873 2837 9874
rect 2792 9869 2798 9873
rect 2802 9869 2808 9873
rect 2812 9869 2818 9873
rect 2822 9869 2828 9873
rect 2832 9869 2837 9873
rect 2792 9868 2837 9869
rect 2792 9864 2793 9868
rect 2797 9864 2803 9868
rect 2807 9864 2813 9868
rect 2817 9864 2823 9868
rect 2827 9864 2833 9868
rect 3101 9949 3107 9953
rect 3111 9949 3117 9953
rect 3121 9949 3127 9953
rect 3131 9949 3137 9953
rect 3141 9949 3146 9953
rect 3101 9948 3146 9949
rect 3101 9944 3102 9948
rect 3106 9944 3112 9948
rect 3116 9944 3122 9948
rect 3126 9944 3132 9948
rect 3136 9944 3142 9948
rect 3101 9943 3146 9944
rect 3101 9939 3107 9943
rect 3111 9939 3117 9943
rect 3121 9939 3127 9943
rect 3131 9939 3137 9943
rect 3141 9939 3146 9943
rect 3101 9938 3146 9939
rect 3101 9934 3102 9938
rect 3106 9934 3112 9938
rect 3116 9934 3122 9938
rect 3126 9934 3132 9938
rect 3136 9934 3142 9938
rect 3101 9933 3146 9934
rect 3101 9929 3107 9933
rect 3111 9929 3117 9933
rect 3121 9929 3127 9933
rect 3131 9929 3137 9933
rect 3141 9929 3146 9933
rect 3101 9928 3146 9929
rect 3101 9924 3102 9928
rect 3106 9924 3112 9928
rect 3116 9924 3122 9928
rect 3126 9924 3132 9928
rect 3136 9924 3142 9928
rect 3101 9923 3146 9924
rect 3101 9919 3107 9923
rect 3111 9919 3117 9923
rect 3121 9919 3127 9923
rect 3131 9919 3137 9923
rect 3141 9919 3146 9923
rect 3101 9918 3146 9919
rect 3101 9914 3102 9918
rect 3106 9914 3112 9918
rect 3116 9914 3122 9918
rect 3126 9914 3132 9918
rect 3136 9914 3142 9918
rect 3101 9913 3146 9914
rect 3101 9909 3107 9913
rect 3111 9909 3117 9913
rect 3121 9909 3127 9913
rect 3131 9909 3137 9913
rect 3141 9909 3146 9913
rect 3101 9908 3146 9909
rect 3101 9904 3102 9908
rect 3106 9904 3112 9908
rect 3116 9904 3122 9908
rect 3126 9904 3132 9908
rect 3136 9904 3142 9908
rect 3101 9903 3146 9904
rect 3101 9899 3107 9903
rect 3111 9899 3117 9903
rect 3121 9899 3127 9903
rect 3131 9899 3137 9903
rect 3141 9899 3146 9903
rect 3101 9898 3146 9899
rect 3101 9894 3102 9898
rect 3106 9894 3112 9898
rect 3116 9894 3122 9898
rect 3126 9894 3132 9898
rect 3136 9894 3142 9898
rect 3101 9893 3146 9894
rect 3101 9889 3107 9893
rect 3111 9889 3117 9893
rect 3121 9889 3127 9893
rect 3131 9889 3137 9893
rect 3141 9889 3146 9893
rect 3101 9888 3146 9889
rect 3101 9884 3102 9888
rect 3106 9884 3112 9888
rect 3116 9884 3122 9888
rect 3126 9884 3132 9888
rect 3136 9884 3142 9888
rect 3101 9883 3146 9884
rect 3101 9879 3107 9883
rect 3111 9879 3117 9883
rect 3121 9879 3127 9883
rect 3131 9879 3137 9883
rect 3141 9879 3146 9883
rect 3101 9878 3146 9879
rect 3101 9874 3102 9878
rect 3106 9874 3112 9878
rect 3116 9874 3122 9878
rect 3126 9874 3132 9878
rect 3136 9874 3142 9878
rect 3101 9873 3146 9874
rect 3101 9869 3107 9873
rect 3111 9869 3117 9873
rect 3121 9869 3127 9873
rect 3131 9869 3137 9873
rect 3141 9869 3146 9873
rect 3101 9868 3146 9869
rect 3101 9864 3102 9868
rect 3106 9864 3112 9868
rect 3116 9864 3122 9868
rect 3126 9864 3132 9868
rect 3136 9864 3142 9868
rect 3410 9949 3416 9953
rect 3420 9949 3426 9953
rect 3430 9949 3436 9953
rect 3440 9949 3446 9953
rect 3450 9949 3455 9953
rect 3410 9948 3455 9949
rect 3410 9944 3411 9948
rect 3415 9944 3421 9948
rect 3425 9944 3431 9948
rect 3435 9944 3441 9948
rect 3445 9944 3451 9948
rect 3410 9943 3455 9944
rect 3410 9939 3416 9943
rect 3420 9939 3426 9943
rect 3430 9939 3436 9943
rect 3440 9939 3446 9943
rect 3450 9939 3455 9943
rect 3410 9938 3455 9939
rect 3410 9934 3411 9938
rect 3415 9934 3421 9938
rect 3425 9934 3431 9938
rect 3435 9934 3441 9938
rect 3445 9934 3451 9938
rect 3410 9933 3455 9934
rect 3410 9929 3416 9933
rect 3420 9929 3426 9933
rect 3430 9929 3436 9933
rect 3440 9929 3446 9933
rect 3450 9929 3455 9933
rect 3410 9928 3455 9929
rect 3410 9924 3411 9928
rect 3415 9924 3421 9928
rect 3425 9924 3431 9928
rect 3435 9924 3441 9928
rect 3445 9924 3451 9928
rect 3410 9923 3455 9924
rect 3410 9919 3416 9923
rect 3420 9919 3426 9923
rect 3430 9919 3436 9923
rect 3440 9919 3446 9923
rect 3450 9919 3455 9923
rect 3410 9918 3455 9919
rect 3410 9914 3411 9918
rect 3415 9914 3421 9918
rect 3425 9914 3431 9918
rect 3435 9914 3441 9918
rect 3445 9914 3451 9918
rect 3410 9913 3455 9914
rect 3410 9909 3416 9913
rect 3420 9909 3426 9913
rect 3430 9909 3436 9913
rect 3440 9909 3446 9913
rect 3450 9909 3455 9913
rect 3410 9908 3455 9909
rect 3410 9904 3411 9908
rect 3415 9904 3421 9908
rect 3425 9904 3431 9908
rect 3435 9904 3441 9908
rect 3445 9904 3451 9908
rect 3410 9903 3455 9904
rect 3410 9899 3416 9903
rect 3420 9899 3426 9903
rect 3430 9899 3436 9903
rect 3440 9899 3446 9903
rect 3450 9899 3455 9903
rect 3410 9898 3455 9899
rect 3410 9894 3411 9898
rect 3415 9894 3421 9898
rect 3425 9894 3431 9898
rect 3435 9894 3441 9898
rect 3445 9894 3451 9898
rect 3410 9893 3455 9894
rect 3410 9889 3416 9893
rect 3420 9889 3426 9893
rect 3430 9889 3436 9893
rect 3440 9889 3446 9893
rect 3450 9889 3455 9893
rect 3410 9888 3455 9889
rect 3410 9884 3411 9888
rect 3415 9884 3421 9888
rect 3425 9884 3431 9888
rect 3435 9884 3441 9888
rect 3445 9884 3451 9888
rect 3410 9883 3455 9884
rect 3410 9879 3416 9883
rect 3420 9879 3426 9883
rect 3430 9879 3436 9883
rect 3440 9879 3446 9883
rect 3450 9879 3455 9883
rect 3410 9878 3455 9879
rect 3410 9874 3411 9878
rect 3415 9874 3421 9878
rect 3425 9874 3431 9878
rect 3435 9874 3441 9878
rect 3445 9874 3451 9878
rect 3410 9873 3455 9874
rect 3410 9869 3416 9873
rect 3420 9869 3426 9873
rect 3430 9869 3436 9873
rect 3440 9869 3446 9873
rect 3450 9869 3455 9873
rect 3410 9868 3455 9869
rect 3410 9864 3411 9868
rect 3415 9864 3421 9868
rect 3425 9864 3431 9868
rect 3435 9864 3441 9868
rect 3445 9864 3451 9868
rect 3719 9949 3725 9953
rect 3729 9949 3735 9953
rect 3739 9949 3745 9953
rect 3749 9949 3755 9953
rect 3759 9949 3764 9953
rect 3719 9948 3764 9949
rect 3719 9944 3720 9948
rect 3724 9944 3730 9948
rect 3734 9944 3740 9948
rect 3744 9944 3750 9948
rect 3754 9944 3760 9948
rect 3719 9943 3764 9944
rect 3719 9939 3725 9943
rect 3729 9939 3735 9943
rect 3739 9939 3745 9943
rect 3749 9939 3755 9943
rect 3759 9939 3764 9943
rect 3719 9938 3764 9939
rect 3719 9934 3720 9938
rect 3724 9934 3730 9938
rect 3734 9934 3740 9938
rect 3744 9934 3750 9938
rect 3754 9934 3760 9938
rect 3719 9933 3764 9934
rect 3719 9929 3725 9933
rect 3729 9929 3735 9933
rect 3739 9929 3745 9933
rect 3749 9929 3755 9933
rect 3759 9929 3764 9933
rect 3719 9928 3764 9929
rect 3719 9924 3720 9928
rect 3724 9924 3730 9928
rect 3734 9924 3740 9928
rect 3744 9924 3750 9928
rect 3754 9924 3760 9928
rect 3719 9923 3764 9924
rect 3719 9919 3725 9923
rect 3729 9919 3735 9923
rect 3739 9919 3745 9923
rect 3749 9919 3755 9923
rect 3759 9919 3764 9923
rect 3719 9918 3764 9919
rect 3719 9914 3720 9918
rect 3724 9914 3730 9918
rect 3734 9914 3740 9918
rect 3744 9914 3750 9918
rect 3754 9914 3760 9918
rect 3719 9913 3764 9914
rect 3719 9909 3725 9913
rect 3729 9909 3735 9913
rect 3739 9909 3745 9913
rect 3749 9909 3755 9913
rect 3759 9909 3764 9913
rect 3719 9908 3764 9909
rect 3719 9904 3720 9908
rect 3724 9904 3730 9908
rect 3734 9904 3740 9908
rect 3744 9904 3750 9908
rect 3754 9904 3760 9908
rect 3719 9903 3764 9904
rect 3719 9899 3725 9903
rect 3729 9899 3735 9903
rect 3739 9899 3745 9903
rect 3749 9899 3755 9903
rect 3759 9899 3764 9903
rect 3719 9898 3764 9899
rect 3719 9894 3720 9898
rect 3724 9894 3730 9898
rect 3734 9894 3740 9898
rect 3744 9894 3750 9898
rect 3754 9894 3760 9898
rect 3719 9893 3764 9894
rect 3719 9889 3725 9893
rect 3729 9889 3735 9893
rect 3739 9889 3745 9893
rect 3749 9889 3755 9893
rect 3759 9889 3764 9893
rect 3719 9888 3764 9889
rect 3719 9884 3720 9888
rect 3724 9884 3730 9888
rect 3734 9884 3740 9888
rect 3744 9884 3750 9888
rect 3754 9884 3760 9888
rect 3719 9883 3764 9884
rect 3719 9879 3725 9883
rect 3729 9879 3735 9883
rect 3739 9879 3745 9883
rect 3749 9879 3755 9883
rect 3759 9879 3764 9883
rect 3719 9878 3764 9879
rect 3719 9874 3720 9878
rect 3724 9874 3730 9878
rect 3734 9874 3740 9878
rect 3744 9874 3750 9878
rect 3754 9874 3760 9878
rect 3719 9873 3764 9874
rect 3719 9869 3725 9873
rect 3729 9869 3735 9873
rect 3739 9869 3745 9873
rect 3749 9869 3755 9873
rect 3759 9869 3764 9873
rect 3719 9868 3764 9869
rect 3719 9864 3720 9868
rect 3724 9864 3730 9868
rect 3734 9864 3740 9868
rect 3744 9864 3750 9868
rect 3754 9864 3760 9868
rect 4028 9949 4034 9953
rect 4038 9949 4044 9953
rect 4048 9949 4054 9953
rect 4058 9949 4064 9953
rect 4068 9949 4073 9953
rect 4028 9948 4073 9949
rect 4028 9944 4029 9948
rect 4033 9944 4039 9948
rect 4043 9944 4049 9948
rect 4053 9944 4059 9948
rect 4063 9944 4069 9948
rect 4028 9943 4073 9944
rect 4028 9939 4034 9943
rect 4038 9939 4044 9943
rect 4048 9939 4054 9943
rect 4058 9939 4064 9943
rect 4068 9939 4073 9943
rect 4028 9938 4073 9939
rect 4028 9934 4029 9938
rect 4033 9934 4039 9938
rect 4043 9934 4049 9938
rect 4053 9934 4059 9938
rect 4063 9934 4069 9938
rect 4028 9933 4073 9934
rect 4028 9929 4034 9933
rect 4038 9929 4044 9933
rect 4048 9929 4054 9933
rect 4058 9929 4064 9933
rect 4068 9929 4073 9933
rect 4028 9928 4073 9929
rect 4028 9924 4029 9928
rect 4033 9924 4039 9928
rect 4043 9924 4049 9928
rect 4053 9924 4059 9928
rect 4063 9924 4069 9928
rect 4028 9923 4073 9924
rect 4028 9919 4034 9923
rect 4038 9919 4044 9923
rect 4048 9919 4054 9923
rect 4058 9919 4064 9923
rect 4068 9919 4073 9923
rect 4028 9918 4073 9919
rect 4028 9914 4029 9918
rect 4033 9914 4039 9918
rect 4043 9914 4049 9918
rect 4053 9914 4059 9918
rect 4063 9914 4069 9918
rect 4028 9913 4073 9914
rect 4028 9909 4034 9913
rect 4038 9909 4044 9913
rect 4048 9909 4054 9913
rect 4058 9909 4064 9913
rect 4068 9909 4073 9913
rect 4028 9908 4073 9909
rect 4028 9904 4029 9908
rect 4033 9904 4039 9908
rect 4043 9904 4049 9908
rect 4053 9904 4059 9908
rect 4063 9904 4069 9908
rect 4028 9903 4073 9904
rect 4028 9899 4034 9903
rect 4038 9899 4044 9903
rect 4048 9899 4054 9903
rect 4058 9899 4064 9903
rect 4068 9899 4073 9903
rect 4028 9898 4073 9899
rect 4028 9894 4029 9898
rect 4033 9894 4039 9898
rect 4043 9894 4049 9898
rect 4053 9894 4059 9898
rect 4063 9894 4069 9898
rect 4028 9893 4073 9894
rect 4028 9889 4034 9893
rect 4038 9889 4044 9893
rect 4048 9889 4054 9893
rect 4058 9889 4064 9893
rect 4068 9889 4073 9893
rect 4028 9888 4073 9889
rect 4028 9884 4029 9888
rect 4033 9884 4039 9888
rect 4043 9884 4049 9888
rect 4053 9884 4059 9888
rect 4063 9884 4069 9888
rect 4028 9883 4073 9884
rect 4028 9879 4034 9883
rect 4038 9879 4044 9883
rect 4048 9879 4054 9883
rect 4058 9879 4064 9883
rect 4068 9879 4073 9883
rect 4028 9878 4073 9879
rect 4028 9874 4029 9878
rect 4033 9874 4039 9878
rect 4043 9874 4049 9878
rect 4053 9874 4059 9878
rect 4063 9874 4069 9878
rect 4028 9873 4073 9874
rect 4028 9869 4034 9873
rect 4038 9869 4044 9873
rect 4048 9869 4054 9873
rect 4058 9869 4064 9873
rect 4068 9869 4073 9873
rect 4028 9868 4073 9869
rect 4028 9864 4029 9868
rect 4033 9864 4039 9868
rect 4043 9864 4049 9868
rect 4053 9864 4059 9868
rect 4063 9864 4069 9868
rect 1778 9827 1782 9831
rect 1743 9826 1799 9827
rect 2087 9827 2091 9831
rect 2052 9826 2108 9827
rect 2396 9827 2400 9831
rect 2361 9826 2417 9827
rect 2705 9827 2709 9831
rect 2670 9826 2726 9827
rect 3014 9827 3018 9831
rect 2979 9826 3035 9827
rect 3941 9827 3945 9831
rect 3906 9826 3962 9827
rect 1743 9823 1799 9824
rect 1743 9818 1799 9819
rect 2052 9823 2108 9824
rect 2052 9818 2108 9819
rect 2361 9823 2417 9824
rect 2361 9818 2417 9819
rect 2670 9823 2726 9824
rect 2670 9818 2726 9819
rect 2979 9823 3035 9824
rect 2979 9818 3035 9819
rect 3906 9823 3962 9824
rect 3906 9818 3962 9819
rect 1743 9815 1799 9816
rect 1778 9811 1782 9815
rect 1743 9810 1799 9811
rect 2052 9815 2108 9816
rect 2087 9811 2091 9815
rect 2052 9810 2108 9811
rect 1743 9807 1799 9808
rect 1743 9802 1799 9803
rect 1743 9799 1799 9800
rect 1778 9795 1782 9799
rect 1743 9794 1799 9795
rect 1743 9791 1799 9792
rect 1743 9786 1799 9787
rect 2361 9815 2417 9816
rect 2396 9811 2400 9815
rect 2361 9810 2417 9811
rect 2052 9807 2108 9808
rect 2052 9802 2108 9803
rect 2052 9799 2108 9800
rect 2087 9795 2091 9799
rect 2052 9794 2108 9795
rect 2052 9791 2108 9792
rect 2052 9786 2108 9787
rect 2670 9815 2726 9816
rect 2705 9811 2709 9815
rect 2670 9810 2726 9811
rect 2361 9807 2417 9808
rect 2361 9802 2417 9803
rect 2361 9799 2417 9800
rect 2396 9795 2400 9799
rect 2361 9794 2417 9795
rect 2361 9791 2417 9792
rect 2361 9786 2417 9787
rect 2979 9815 3035 9816
rect 3014 9811 3018 9815
rect 2979 9810 3035 9811
rect 2670 9807 2726 9808
rect 2670 9802 2726 9803
rect 2670 9799 2726 9800
rect 2705 9795 2709 9799
rect 2670 9794 2726 9795
rect 2670 9791 2726 9792
rect 2670 9786 2726 9787
rect 3906 9815 3962 9816
rect 3941 9811 3945 9815
rect 3906 9810 3962 9811
rect 2979 9807 3035 9808
rect 2979 9802 3035 9803
rect 2979 9799 3035 9800
rect 3014 9795 3018 9799
rect 2979 9794 3035 9795
rect 2979 9791 3035 9792
rect 2979 9786 3035 9787
rect 3906 9807 3962 9808
rect 3906 9802 3962 9803
rect 3906 9799 3962 9800
rect 3941 9795 3945 9799
rect 3906 9794 3962 9795
rect 3906 9791 3962 9792
rect 3906 9786 3962 9787
rect 1743 9783 1799 9784
rect 1778 9779 1782 9783
rect 2052 9783 2108 9784
rect 2087 9779 2091 9783
rect 2361 9783 2417 9784
rect 2396 9779 2400 9783
rect 2670 9783 2726 9784
rect 2705 9779 2709 9783
rect 2979 9783 3035 9784
rect 3014 9779 3018 9783
rect 3906 9783 3962 9784
rect 3941 9779 3945 9783
rect 2855 9322 2856 9330
rect 2858 9322 2861 9330
rect 2863 9322 2864 9330
rect 2876 9322 2877 9330
rect 2879 9326 2880 9330
rect 2879 9322 2884 9326
rect 2892 9322 2893 9330
rect 2895 9322 2898 9330
rect 2900 9322 2901 9330
rect 2918 9322 2919 9330
rect 2921 9322 2922 9330
rect 2934 9322 2935 9330
rect 2937 9326 2938 9330
rect 2937 9322 2942 9326
rect 2950 9322 2951 9330
rect 2953 9322 2956 9330
rect 2958 9322 2959 9330
rect 2971 9322 2972 9330
rect 2974 9322 2975 9330
rect 2987 9322 2988 9330
rect 2990 9322 2993 9330
rect 2995 9322 2996 9330
rect 3008 9322 3009 9330
rect 3011 9326 3012 9330
rect 3011 9322 3016 9326
rect 3024 9322 3025 9330
rect 3027 9322 3030 9330
rect 3032 9322 3033 9330
rect 3050 9322 3051 9330
rect 3053 9322 3054 9330
rect 3066 9322 3067 9330
rect 3069 9326 3070 9330
rect 3069 9322 3074 9326
rect 3082 9322 3083 9330
rect 3085 9322 3088 9330
rect 3090 9322 3091 9330
rect 3103 9322 3104 9330
rect 3106 9322 3107 9330
rect 3119 9322 3120 9330
rect 3122 9322 3125 9330
rect 3127 9322 3128 9330
rect 3140 9322 3141 9330
rect 3143 9326 3144 9330
rect 3143 9322 3148 9326
rect 3156 9322 3157 9330
rect 3159 9322 3162 9330
rect 3164 9322 3165 9330
rect 3182 9322 3183 9330
rect 3185 9322 3186 9330
rect 3198 9322 3199 9330
rect 3201 9326 3202 9330
rect 3201 9322 3206 9326
rect 3214 9322 3215 9330
rect 3217 9322 3220 9330
rect 3222 9322 3223 9330
rect 3235 9322 3236 9330
rect 3238 9322 3239 9330
rect 3251 9322 3252 9330
rect 3254 9322 3257 9330
rect 3259 9322 3260 9330
rect 3272 9322 3273 9330
rect 3275 9326 3276 9330
rect 3275 9322 3280 9326
rect 3288 9322 3289 9330
rect 3291 9322 3294 9330
rect 3296 9322 3297 9330
rect 3314 9322 3315 9330
rect 3317 9322 3318 9330
rect 3330 9322 3331 9330
rect 3333 9326 3334 9330
rect 3333 9322 3338 9326
rect 3346 9322 3347 9330
rect 3349 9322 3352 9330
rect 3354 9322 3355 9330
rect 3367 9322 3368 9330
rect 3370 9322 3371 9330
rect 3800 9322 3801 9330
rect 3803 9322 3806 9330
rect 3808 9322 3809 9330
rect 3821 9322 3822 9330
rect 3824 9326 3825 9330
rect 3824 9322 3829 9326
rect 3837 9322 3838 9330
rect 3840 9322 3843 9330
rect 3845 9322 3846 9330
rect 3863 9322 3864 9330
rect 3866 9322 3867 9330
rect 3879 9322 3880 9330
rect 3882 9326 3883 9330
rect 3882 9322 3887 9326
rect 3895 9322 3896 9330
rect 3898 9322 3901 9330
rect 3903 9322 3904 9330
rect 3916 9322 3917 9330
rect 3919 9322 3920 9330
rect 3932 9322 3933 9330
rect 3935 9322 3938 9330
rect 3940 9322 3941 9330
rect 3953 9322 3954 9330
rect 3956 9326 3957 9330
rect 3956 9322 3961 9326
rect 3969 9322 3970 9330
rect 3972 9322 3975 9330
rect 3977 9322 3978 9330
rect 3995 9322 3996 9330
rect 3998 9322 3999 9330
rect 4011 9322 4012 9330
rect 4014 9326 4015 9330
rect 4014 9322 4019 9326
rect 4027 9322 4028 9330
rect 4030 9322 4033 9330
rect 4035 9322 4036 9330
rect 4048 9322 4049 9330
rect 4051 9322 4052 9330
rect 4064 9322 4065 9330
rect 4067 9322 4070 9330
rect 4072 9322 4073 9330
rect 4085 9322 4086 9330
rect 4088 9326 4089 9330
rect 4088 9322 4093 9326
rect 4101 9322 4102 9330
rect 4104 9322 4107 9330
rect 4109 9322 4110 9330
rect 4127 9322 4128 9330
rect 4130 9322 4131 9330
rect 4143 9322 4144 9330
rect 4146 9326 4147 9330
rect 4146 9322 4151 9326
rect 4159 9322 4160 9330
rect 4162 9322 4165 9330
rect 4167 9322 4168 9330
rect 4180 9322 4181 9330
rect 4183 9322 4184 9330
rect 4196 9322 4197 9330
rect 4199 9322 4202 9330
rect 4204 9322 4205 9330
rect 4217 9322 4218 9330
rect 4220 9326 4221 9330
rect 4220 9322 4225 9326
rect 4233 9322 4234 9330
rect 4236 9322 4239 9330
rect 4241 9322 4242 9330
rect 4259 9322 4260 9330
rect 4262 9322 4263 9330
rect 4275 9322 4276 9330
rect 4278 9326 4279 9330
rect 4278 9322 4283 9326
rect 4291 9322 4292 9330
rect 4294 9322 4297 9330
rect 4299 9322 4300 9330
rect 4312 9322 4313 9330
rect 4315 9322 4316 9330
rect 2503 9289 2504 9297
rect 2506 9289 2509 9297
rect 2511 9289 2512 9297
rect 2524 9289 2525 9297
rect 2527 9293 2528 9297
rect 2527 9289 2532 9293
rect 2540 9289 2541 9297
rect 2543 9289 2546 9297
rect 2548 9289 2549 9297
rect 2566 9289 2567 9297
rect 2569 9289 2570 9297
rect 2582 9289 2583 9297
rect 2585 9293 2586 9297
rect 2585 9289 2590 9293
rect 2598 9289 2599 9297
rect 2601 9289 2604 9297
rect 2606 9289 2607 9297
rect 2619 9289 2620 9297
rect 2622 9289 2623 9297
rect 3448 9289 3449 9297
rect 3451 9289 3454 9297
rect 3456 9289 3457 9297
rect 3469 9289 3470 9297
rect 3472 9293 3473 9297
rect 3472 9289 3477 9293
rect 3485 9289 3486 9297
rect 3488 9289 3491 9297
rect 3493 9289 3494 9297
rect 3511 9289 3512 9297
rect 3514 9289 3515 9297
rect 3527 9289 3528 9297
rect 3530 9293 3531 9297
rect 3530 9289 3535 9293
rect 3543 9289 3544 9297
rect 3546 9289 3549 9297
rect 3551 9289 3552 9297
rect 3564 9289 3565 9297
rect 3567 9289 3568 9297
rect 3034 9251 3035 9259
rect 3037 9251 3038 9259
rect 2860 9238 2861 9246
rect 2863 9238 2864 9246
rect 2876 9238 2877 9246
rect 2879 9238 2880 9246
rect 2892 9238 2893 9246
rect 2895 9238 2896 9246
rect 2911 9238 2916 9246
rect 2918 9238 2921 9246
rect 2923 9238 2924 9246
rect 2945 9238 2947 9246
rect 2949 9238 2950 9246
rect 2967 9238 2968 9246
rect 2970 9238 2971 9246
rect 2983 9238 2988 9246
rect 2990 9238 2993 9246
rect 2995 9238 2996 9246
rect 3010 9238 3011 9246
rect 3013 9238 3014 9246
rect 3058 9245 3061 9253
rect 3063 9245 3066 9253
rect 3068 9245 3069 9253
rect 3088 9251 3089 9259
rect 3091 9251 3092 9259
rect 3115 9251 3116 9259
rect 3118 9251 3119 9259
rect 3139 9245 3142 9253
rect 3144 9245 3147 9253
rect 3149 9245 3150 9253
rect 3169 9251 3170 9259
rect 3172 9251 3173 9259
rect 3979 9251 3980 9259
rect 3982 9251 3983 9259
rect 3805 9238 3806 9246
rect 3808 9238 3809 9246
rect 3821 9238 3822 9246
rect 3824 9238 3825 9246
rect 3837 9238 3838 9246
rect 3840 9238 3841 9246
rect 3856 9238 3861 9246
rect 3863 9238 3866 9246
rect 3868 9238 3869 9246
rect 3890 9238 3892 9246
rect 3894 9238 3895 9246
rect 3912 9238 3913 9246
rect 3915 9238 3916 9246
rect 3928 9238 3933 9246
rect 3935 9238 3938 9246
rect 3940 9238 3941 9246
rect 3955 9238 3956 9246
rect 3958 9238 3959 9246
rect 4003 9245 4006 9253
rect 4008 9245 4011 9253
rect 4013 9245 4014 9253
rect 4033 9251 4034 9259
rect 4036 9251 4037 9259
rect 4060 9251 4061 9259
rect 4063 9251 4064 9259
rect 4084 9245 4087 9253
rect 4089 9245 4092 9253
rect 4094 9245 4095 9253
rect 4114 9251 4115 9259
rect 4117 9251 4118 9259
rect 2494 9187 2495 9195
rect 2497 9187 2498 9195
rect 2510 9187 2511 9195
rect 2513 9187 2516 9195
rect 2518 9187 2519 9195
rect 2531 9191 2532 9195
rect 2527 9187 2532 9191
rect 2534 9187 2535 9195
rect 2547 9187 2548 9195
rect 2550 9187 2551 9195
rect 2568 9187 2569 9195
rect 2571 9187 2574 9195
rect 2576 9187 2577 9195
rect 2589 9191 2590 9195
rect 2585 9187 2590 9191
rect 2592 9187 2593 9195
rect 2605 9187 2606 9195
rect 2608 9187 2611 9195
rect 2613 9187 2614 9195
rect 3439 9187 3440 9195
rect 3442 9187 3443 9195
rect 3455 9187 3456 9195
rect 3458 9187 3461 9195
rect 3463 9187 3464 9195
rect 3476 9191 3477 9195
rect 3472 9187 3477 9191
rect 3479 9187 3480 9195
rect 3492 9187 3493 9195
rect 3495 9187 3496 9195
rect 3513 9187 3514 9195
rect 3516 9187 3519 9195
rect 3521 9187 3522 9195
rect 3534 9191 3535 9195
rect 3530 9187 3535 9191
rect 3537 9187 3538 9195
rect 3550 9187 3551 9195
rect 3553 9187 3556 9195
rect 3558 9187 3559 9195
rect 2860 9152 2861 9160
rect 2863 9152 2864 9160
rect 2876 9152 2877 9160
rect 2879 9152 2880 9160
rect 2892 9152 2893 9160
rect 2895 9152 2896 9160
rect 2911 9152 2916 9160
rect 2918 9152 2921 9160
rect 2923 9152 2924 9160
rect 2945 9152 2947 9160
rect 2949 9152 2950 9160
rect 2967 9152 2968 9160
rect 2970 9152 2971 9160
rect 2983 9152 2988 9160
rect 2990 9152 2993 9160
rect 2995 9152 2996 9160
rect 3010 9152 3011 9160
rect 3013 9152 3014 9160
rect 3058 9153 3061 9161
rect 3063 9153 3066 9161
rect 3068 9153 3069 9161
rect 3139 9153 3142 9161
rect 3144 9153 3147 9161
rect 3149 9153 3150 9161
rect 3805 9152 3806 9160
rect 3808 9152 3809 9160
rect 3821 9152 3822 9160
rect 3824 9152 3825 9160
rect 3837 9152 3838 9160
rect 3840 9152 3841 9160
rect 3856 9152 3861 9160
rect 3863 9152 3866 9160
rect 3868 9152 3869 9160
rect 3890 9152 3892 9160
rect 3894 9152 3895 9160
rect 3912 9152 3913 9160
rect 3915 9152 3916 9160
rect 3928 9152 3933 9160
rect 3935 9152 3938 9160
rect 3940 9152 3941 9160
rect 3955 9152 3956 9160
rect 3958 9152 3959 9160
rect 4003 9153 4006 9161
rect 4008 9153 4011 9161
rect 4013 9153 4014 9161
rect 4084 9153 4087 9161
rect 4089 9153 4092 9161
rect 4094 9153 4095 9161
rect 2860 9106 2861 9114
rect 2863 9106 2864 9114
rect 2876 9106 2877 9114
rect 2879 9106 2880 9114
rect 2892 9106 2893 9114
rect 2895 9106 2896 9114
rect 2911 9106 2916 9114
rect 2918 9106 2921 9114
rect 2923 9106 2924 9114
rect 2945 9106 2947 9114
rect 2949 9106 2950 9114
rect 2967 9106 2968 9114
rect 2970 9106 2971 9114
rect 2983 9106 2988 9114
rect 2990 9106 2993 9114
rect 2995 9106 2996 9114
rect 3010 9106 3011 9114
rect 3013 9106 3014 9114
rect 3058 9113 3061 9121
rect 3063 9113 3066 9121
rect 3068 9113 3069 9121
rect 3088 9119 3089 9127
rect 3091 9119 3092 9127
rect 3139 9119 3140 9127
rect 3142 9119 3143 9127
rect 3163 9113 3166 9121
rect 3168 9113 3171 9121
rect 3173 9113 3174 9121
rect 3193 9119 3194 9127
rect 3196 9119 3197 9127
rect 3805 9106 3806 9114
rect 3808 9106 3809 9114
rect 3821 9106 3822 9114
rect 3824 9106 3825 9114
rect 3837 9106 3838 9114
rect 3840 9106 3841 9114
rect 3856 9106 3861 9114
rect 3863 9106 3866 9114
rect 3868 9106 3869 9114
rect 3890 9106 3892 9114
rect 3894 9106 3895 9114
rect 3912 9106 3913 9114
rect 3915 9106 3916 9114
rect 3928 9106 3933 9114
rect 3935 9106 3938 9114
rect 3940 9106 3941 9114
rect 3955 9106 3956 9114
rect 3958 9106 3959 9114
rect 4003 9113 4006 9121
rect 4008 9113 4011 9121
rect 4013 9113 4014 9121
rect 4033 9119 4034 9127
rect 4036 9119 4037 9127
rect 4084 9119 4085 9127
rect 4087 9119 4088 9127
rect 3370 9090 3371 9098
rect 3373 9090 3374 9098
rect 3394 9084 3397 9092
rect 3399 9084 3402 9092
rect 3404 9084 3405 9092
rect 3424 9090 3425 9098
rect 3427 9090 3428 9098
rect 3556 9065 3557 9095
rect 3559 9065 3560 9095
rect 3609 9065 3610 9095
rect 3612 9065 3613 9095
rect 4108 9113 4111 9121
rect 4113 9113 4116 9121
rect 4118 9113 4119 9121
rect 4138 9119 4139 9127
rect 4141 9119 4142 9127
rect 2860 9020 2861 9028
rect 2863 9020 2864 9028
rect 2876 9020 2877 9028
rect 2879 9020 2880 9028
rect 2892 9020 2893 9028
rect 2895 9020 2896 9028
rect 2911 9020 2916 9028
rect 2918 9020 2921 9028
rect 2923 9020 2924 9028
rect 2945 9020 2947 9028
rect 2949 9020 2950 9028
rect 2967 9020 2968 9028
rect 2970 9020 2971 9028
rect 2983 9020 2988 9028
rect 2990 9020 2993 9028
rect 2995 9020 2996 9028
rect 3010 9020 3011 9028
rect 3013 9020 3014 9028
rect 3058 9022 3061 9030
rect 3063 9022 3066 9030
rect 3068 9022 3069 9030
rect 3163 9022 3166 9030
rect 3168 9022 3171 9030
rect 3173 9022 3174 9030
rect 3805 9020 3806 9028
rect 3808 9020 3809 9028
rect 3821 9020 3822 9028
rect 3824 9020 3825 9028
rect 3837 9020 3838 9028
rect 3840 9020 3841 9028
rect 3856 9020 3861 9028
rect 3863 9020 3866 9028
rect 3868 9020 3869 9028
rect 3890 9020 3892 9028
rect 3894 9020 3895 9028
rect 3912 9020 3913 9028
rect 3915 9020 3916 9028
rect 3928 9020 3933 9028
rect 3935 9020 3938 9028
rect 3940 9020 3941 9028
rect 3955 9020 3956 9028
rect 3958 9020 3959 9028
rect 4003 9022 4006 9030
rect 4008 9022 4011 9030
rect 4013 9022 4014 9030
rect 4108 9022 4111 9030
rect 4113 9022 4116 9030
rect 4118 9022 4119 9030
rect 2860 8974 2861 8982
rect 2863 8974 2864 8982
rect 2876 8974 2877 8982
rect 2879 8974 2880 8982
rect 2892 8974 2893 8982
rect 2895 8974 2896 8982
rect 2911 8974 2916 8982
rect 2918 8974 2921 8982
rect 2923 8974 2924 8982
rect 2945 8974 2947 8982
rect 2949 8974 2950 8982
rect 2967 8974 2968 8982
rect 2970 8974 2971 8982
rect 2983 8974 2988 8982
rect 2990 8974 2993 8982
rect 2995 8974 2996 8982
rect 3010 8974 3011 8982
rect 3013 8974 3014 8982
rect 3058 8981 3061 8989
rect 3063 8981 3066 8989
rect 3068 8981 3069 8989
rect 3088 8987 3089 8995
rect 3091 8987 3092 8995
rect 3115 8987 3116 8995
rect 3118 8987 3119 8995
rect 3139 8981 3142 8989
rect 3144 8981 3147 8989
rect 3149 8981 3150 8989
rect 3169 8987 3170 8995
rect 3172 8987 3173 8995
rect 3205 8987 3206 8995
rect 3208 8987 3209 8995
rect 3229 8981 3232 8989
rect 3234 8981 3237 8989
rect 3239 8981 3240 8989
rect 3259 8987 3260 8995
rect 3262 8987 3263 8995
rect 3394 8988 3397 8996
rect 3399 8988 3402 8996
rect 3404 8988 3405 8996
rect 3805 8974 3806 8982
rect 3808 8974 3809 8982
rect 3821 8974 3822 8982
rect 3824 8974 3825 8982
rect 3837 8974 3838 8982
rect 3840 8974 3841 8982
rect 3856 8974 3861 8982
rect 3863 8974 3866 8982
rect 3868 8974 3869 8982
rect 3890 8974 3892 8982
rect 3894 8974 3895 8982
rect 3912 8974 3913 8982
rect 3915 8974 3916 8982
rect 3928 8974 3933 8982
rect 3935 8974 3938 8982
rect 3940 8974 3941 8982
rect 3955 8974 3956 8982
rect 3958 8974 3959 8982
rect 4003 8981 4006 8989
rect 4008 8981 4011 8989
rect 4013 8981 4014 8989
rect 4033 8987 4034 8995
rect 4036 8987 4037 8995
rect 4060 8987 4061 8995
rect 4063 8987 4064 8995
rect 3348 8960 3349 8968
rect 3351 8960 3352 8968
rect 3370 8960 3371 8968
rect 3373 8960 3374 8968
rect 3394 8954 3397 8962
rect 3399 8954 3402 8962
rect 3404 8954 3405 8962
rect 3424 8960 3425 8968
rect 3427 8960 3428 8968
rect 3462 8935 3463 8965
rect 3465 8935 3466 8965
rect 3515 8935 3516 8965
rect 3518 8935 3519 8965
rect 4084 8981 4087 8989
rect 4089 8981 4092 8989
rect 4094 8981 4095 8989
rect 4114 8987 4115 8995
rect 4117 8987 4118 8995
rect 4150 8987 4151 8995
rect 4153 8987 4154 8995
rect 4174 8981 4177 8989
rect 4179 8981 4182 8989
rect 4184 8981 4185 8989
rect 4204 8987 4205 8995
rect 4207 8987 4208 8995
rect 2860 8888 2861 8896
rect 2863 8888 2864 8896
rect 2876 8888 2877 8896
rect 2879 8888 2880 8896
rect 2892 8888 2893 8896
rect 2895 8888 2896 8896
rect 2911 8888 2916 8896
rect 2918 8888 2921 8896
rect 2923 8888 2924 8896
rect 2945 8888 2947 8896
rect 2949 8888 2950 8896
rect 2967 8888 2968 8896
rect 2970 8888 2971 8896
rect 2983 8888 2988 8896
rect 2990 8888 2993 8896
rect 2995 8888 2996 8896
rect 3010 8888 3011 8896
rect 3013 8888 3014 8896
rect 3058 8887 3061 8895
rect 3063 8887 3066 8895
rect 3068 8887 3069 8895
rect 3139 8887 3142 8895
rect 3144 8887 3147 8895
rect 3149 8887 3150 8895
rect 3229 8887 3232 8895
rect 3234 8887 3237 8895
rect 3239 8887 3240 8895
rect 3805 8888 3806 8896
rect 3808 8888 3809 8896
rect 3821 8888 3822 8896
rect 3824 8888 3825 8896
rect 3837 8888 3838 8896
rect 3840 8888 3841 8896
rect 3856 8888 3861 8896
rect 3863 8888 3866 8896
rect 3868 8888 3869 8896
rect 3890 8888 3892 8896
rect 3894 8888 3895 8896
rect 3912 8888 3913 8896
rect 3915 8888 3916 8896
rect 3928 8888 3933 8896
rect 3935 8888 3938 8896
rect 3940 8888 3941 8896
rect 3955 8888 3956 8896
rect 3958 8888 3959 8896
rect 4003 8887 4006 8895
rect 4008 8887 4011 8895
rect 4013 8887 4014 8895
rect 4084 8887 4087 8895
rect 4089 8887 4092 8895
rect 4094 8887 4095 8895
rect 4174 8887 4177 8895
rect 4179 8887 4182 8895
rect 4184 8887 4185 8895
rect 2860 8842 2861 8850
rect 2863 8842 2864 8850
rect 2876 8842 2877 8850
rect 2879 8842 2880 8850
rect 2892 8842 2893 8850
rect 2895 8842 2896 8850
rect 2911 8842 2916 8850
rect 2918 8842 2921 8850
rect 2923 8842 2924 8850
rect 2945 8842 2947 8850
rect 2949 8842 2950 8850
rect 2967 8842 2968 8850
rect 2970 8842 2971 8850
rect 2983 8842 2988 8850
rect 2990 8842 2993 8850
rect 2995 8842 2996 8850
rect 3010 8842 3011 8850
rect 3013 8842 3014 8850
rect 3058 8849 3061 8857
rect 3063 8849 3066 8857
rect 3068 8849 3069 8857
rect 3088 8855 3089 8863
rect 3091 8855 3092 8863
rect 3394 8858 3397 8866
rect 3399 8858 3402 8866
rect 3404 8858 3405 8866
rect 3805 8842 3806 8850
rect 3808 8842 3809 8850
rect 3821 8842 3822 8850
rect 3824 8842 3825 8850
rect 3837 8842 3838 8850
rect 3840 8842 3841 8850
rect 3856 8842 3861 8850
rect 3863 8842 3866 8850
rect 3868 8842 3869 8850
rect 3890 8842 3892 8850
rect 3894 8842 3895 8850
rect 3912 8842 3913 8850
rect 3915 8842 3916 8850
rect 3928 8842 3933 8850
rect 3935 8842 3938 8850
rect 3940 8842 3941 8850
rect 3955 8842 3956 8850
rect 3958 8842 3959 8850
rect 4003 8849 4006 8857
rect 4008 8849 4011 8857
rect 4013 8849 4014 8857
rect 4033 8855 4034 8863
rect 4036 8855 4037 8863
rect 2371 8787 2372 8795
rect 2374 8787 2377 8795
rect 2379 8787 2380 8795
rect 2392 8787 2393 8795
rect 2395 8791 2396 8795
rect 2395 8787 2400 8791
rect 2408 8787 2409 8795
rect 2411 8787 2414 8795
rect 2416 8787 2417 8795
rect 2434 8787 2435 8795
rect 2437 8787 2438 8795
rect 2450 8787 2451 8795
rect 2453 8791 2454 8795
rect 2453 8787 2458 8791
rect 2466 8787 2467 8795
rect 2469 8787 2472 8795
rect 2474 8787 2475 8795
rect 2487 8787 2488 8795
rect 2490 8787 2491 8795
rect 2503 8787 2504 8795
rect 2506 8787 2509 8795
rect 2511 8787 2512 8795
rect 2524 8787 2525 8795
rect 2527 8791 2528 8795
rect 2527 8787 2532 8791
rect 2540 8787 2541 8795
rect 2543 8787 2546 8795
rect 2548 8787 2549 8795
rect 2566 8787 2567 8795
rect 2569 8787 2570 8795
rect 2582 8787 2583 8795
rect 2585 8791 2586 8795
rect 2585 8787 2590 8791
rect 2598 8787 2599 8795
rect 2601 8787 2604 8795
rect 2606 8787 2607 8795
rect 2619 8787 2620 8795
rect 2622 8787 2623 8795
rect 2635 8787 2636 8795
rect 2638 8787 2641 8795
rect 2643 8787 2644 8795
rect 2656 8787 2657 8795
rect 2659 8791 2660 8795
rect 2659 8787 2664 8791
rect 2672 8787 2673 8795
rect 2675 8787 2678 8795
rect 2680 8787 2681 8795
rect 2698 8787 2699 8795
rect 2701 8787 2702 8795
rect 2714 8787 2715 8795
rect 2717 8791 2718 8795
rect 2717 8787 2722 8791
rect 2730 8787 2731 8795
rect 2733 8787 2736 8795
rect 2738 8787 2739 8795
rect 2751 8787 2752 8795
rect 2754 8787 2755 8795
rect 3316 8787 3317 8795
rect 3319 8787 3322 8795
rect 3324 8787 3325 8795
rect 3337 8787 3338 8795
rect 3340 8791 3341 8795
rect 3340 8787 3345 8791
rect 3353 8787 3354 8795
rect 3356 8787 3359 8795
rect 3361 8787 3362 8795
rect 3379 8787 3380 8795
rect 3382 8787 3383 8795
rect 3395 8787 3396 8795
rect 3398 8791 3399 8795
rect 3398 8787 3403 8791
rect 3411 8787 3412 8795
rect 3414 8787 3417 8795
rect 3419 8787 3420 8795
rect 3432 8787 3433 8795
rect 3435 8787 3436 8795
rect 3448 8787 3449 8795
rect 3451 8787 3454 8795
rect 3456 8787 3457 8795
rect 3469 8787 3470 8795
rect 3472 8791 3473 8795
rect 3472 8787 3477 8791
rect 3485 8787 3486 8795
rect 3488 8787 3491 8795
rect 3493 8787 3494 8795
rect 3511 8787 3512 8795
rect 3514 8787 3515 8795
rect 3527 8787 3528 8795
rect 3530 8791 3531 8795
rect 3530 8787 3535 8791
rect 3543 8787 3544 8795
rect 3546 8787 3549 8795
rect 3551 8787 3552 8795
rect 3564 8787 3565 8795
rect 3567 8787 3568 8795
rect 3580 8787 3581 8795
rect 3583 8787 3586 8795
rect 3588 8787 3589 8795
rect 3601 8787 3602 8795
rect 3604 8791 3605 8795
rect 3604 8787 3609 8791
rect 3617 8787 3618 8795
rect 3620 8787 3623 8795
rect 3625 8787 3626 8795
rect 3643 8787 3644 8795
rect 3646 8787 3647 8795
rect 3659 8787 3660 8795
rect 3662 8791 3663 8795
rect 3662 8787 3667 8791
rect 3675 8787 3676 8795
rect 3678 8787 3681 8795
rect 3683 8787 3684 8795
rect 3696 8787 3697 8795
rect 3699 8787 3700 8795
rect 2860 8756 2861 8764
rect 2863 8756 2864 8764
rect 2876 8756 2877 8764
rect 2879 8756 2880 8764
rect 2892 8756 2893 8764
rect 2895 8756 2896 8764
rect 2911 8756 2916 8764
rect 2918 8756 2921 8764
rect 2923 8756 2924 8764
rect 2945 8756 2947 8764
rect 2949 8756 2950 8764
rect 2967 8756 2968 8764
rect 2970 8756 2971 8764
rect 2983 8756 2988 8764
rect 2990 8756 2993 8764
rect 2995 8756 2996 8764
rect 3010 8756 3011 8764
rect 3013 8756 3014 8764
rect 3058 8751 3061 8759
rect 3063 8751 3066 8759
rect 3068 8751 3069 8759
rect 3094 8756 3095 8764
rect 3097 8756 3098 8764
rect 3102 8756 3108 8764
rect 3112 8756 3113 8764
rect 3115 8756 3116 8764
rect 3137 8756 3138 8764
rect 3140 8756 3141 8764
rect 3153 8756 3154 8764
rect 3156 8756 3157 8764
rect 3172 8756 3177 8764
rect 3179 8756 3182 8764
rect 3184 8756 3185 8764
rect 3206 8756 3208 8764
rect 3210 8756 3211 8764
rect 3228 8756 3229 8764
rect 3231 8756 3232 8764
rect 3244 8756 3249 8764
rect 3251 8756 3254 8764
rect 3256 8756 3257 8764
rect 3271 8756 3272 8764
rect 3274 8756 3275 8764
rect 3805 8756 3806 8764
rect 3808 8756 3809 8764
rect 3821 8756 3822 8764
rect 3824 8756 3825 8764
rect 3837 8756 3838 8764
rect 3840 8756 3841 8764
rect 3856 8756 3861 8764
rect 3863 8756 3866 8764
rect 3868 8756 3869 8764
rect 3890 8756 3892 8764
rect 3894 8756 3895 8764
rect 3912 8756 3913 8764
rect 3915 8756 3916 8764
rect 3928 8756 3933 8764
rect 3935 8756 3938 8764
rect 3940 8756 3941 8764
rect 3955 8756 3956 8764
rect 3958 8756 3959 8764
rect 4003 8751 4006 8759
rect 4008 8751 4011 8759
rect 4013 8751 4014 8759
rect 4039 8756 4040 8764
rect 4042 8756 4043 8764
rect 4047 8756 4053 8764
rect 4057 8756 4058 8764
rect 4060 8756 4061 8764
rect 4082 8756 4083 8764
rect 4085 8756 4086 8764
rect 4098 8756 4099 8764
rect 4101 8756 4102 8764
rect 4117 8756 4122 8764
rect 4124 8756 4127 8764
rect 4129 8756 4130 8764
rect 4151 8756 4153 8764
rect 4155 8756 4156 8764
rect 4173 8756 4174 8764
rect 4176 8756 4177 8764
rect 4189 8756 4194 8764
rect 4196 8756 4199 8764
rect 4201 8756 4202 8764
rect 4216 8756 4217 8764
rect 4219 8756 4220 8764
rect 3154 8675 3155 8683
rect 3157 8675 3160 8683
rect 3162 8675 3163 8683
rect 3175 8675 3176 8683
rect 3178 8679 3179 8683
rect 3178 8675 3183 8679
rect 3191 8675 3192 8683
rect 3194 8675 3197 8683
rect 3199 8675 3200 8683
rect 3217 8675 3218 8683
rect 3220 8675 3221 8683
rect 3233 8675 3234 8683
rect 3236 8679 3237 8683
rect 3236 8675 3241 8679
rect 3249 8675 3250 8683
rect 3252 8675 3255 8683
rect 3257 8675 3258 8683
rect 3270 8675 3271 8683
rect 3273 8675 3274 8683
rect 4099 8675 4100 8683
rect 4102 8675 4105 8683
rect 4107 8675 4108 8683
rect 4120 8675 4121 8683
rect 4123 8679 4124 8683
rect 4123 8675 4128 8679
rect 4136 8675 4137 8683
rect 4139 8675 4142 8683
rect 4144 8675 4145 8683
rect 4162 8675 4163 8683
rect 4165 8675 4166 8683
rect 4178 8675 4179 8683
rect 4181 8679 4182 8683
rect 4181 8675 4186 8679
rect 4194 8675 4195 8683
rect 4197 8675 4200 8683
rect 4202 8675 4203 8683
rect 4215 8675 4216 8683
rect 4218 8675 4219 8683
rect 2371 8645 2372 8653
rect 2374 8645 2377 8653
rect 2379 8645 2380 8653
rect 2392 8645 2393 8653
rect 2395 8649 2396 8653
rect 2395 8645 2400 8649
rect 2408 8645 2409 8653
rect 2411 8645 2414 8653
rect 2416 8645 2417 8653
rect 2434 8645 2435 8653
rect 2437 8645 2438 8653
rect 2450 8645 2451 8653
rect 2453 8649 2454 8653
rect 2453 8645 2458 8649
rect 2466 8645 2467 8653
rect 2469 8645 2472 8653
rect 2474 8645 2475 8653
rect 2487 8645 2488 8653
rect 2490 8645 2491 8653
rect 2503 8645 2504 8653
rect 2506 8645 2509 8653
rect 2511 8645 2512 8653
rect 2524 8645 2525 8653
rect 2527 8649 2528 8653
rect 2527 8645 2532 8649
rect 2540 8645 2541 8653
rect 2543 8645 2546 8653
rect 2548 8645 2549 8653
rect 2566 8645 2567 8653
rect 2569 8645 2570 8653
rect 2582 8645 2583 8653
rect 2585 8649 2586 8653
rect 2585 8645 2590 8649
rect 2598 8645 2599 8653
rect 2601 8645 2604 8653
rect 2606 8645 2607 8653
rect 2619 8645 2620 8653
rect 2622 8645 2623 8653
rect 2635 8645 2636 8653
rect 2638 8645 2641 8653
rect 2643 8645 2644 8653
rect 2656 8645 2657 8653
rect 2659 8649 2660 8653
rect 2659 8645 2664 8649
rect 2672 8645 2673 8653
rect 2675 8645 2678 8653
rect 2680 8645 2681 8653
rect 2698 8645 2699 8653
rect 2701 8645 2702 8653
rect 2714 8645 2715 8653
rect 2717 8649 2718 8653
rect 2717 8645 2722 8649
rect 2730 8645 2731 8653
rect 2733 8645 2736 8653
rect 2738 8645 2739 8653
rect 2751 8645 2752 8653
rect 2754 8645 2755 8653
rect 3316 8645 3317 8653
rect 3319 8645 3322 8653
rect 3324 8645 3325 8653
rect 3337 8645 3338 8653
rect 3340 8649 3341 8653
rect 3340 8645 3345 8649
rect 3353 8645 3354 8653
rect 3356 8645 3359 8653
rect 3361 8645 3362 8653
rect 3379 8645 3380 8653
rect 3382 8645 3383 8653
rect 3395 8645 3396 8653
rect 3398 8649 3399 8653
rect 3398 8645 3403 8649
rect 3411 8645 3412 8653
rect 3414 8645 3417 8653
rect 3419 8645 3420 8653
rect 3432 8645 3433 8653
rect 3435 8645 3436 8653
rect 3448 8645 3449 8653
rect 3451 8645 3454 8653
rect 3456 8645 3457 8653
rect 3469 8645 3470 8653
rect 3472 8649 3473 8653
rect 3472 8645 3477 8649
rect 3485 8645 3486 8653
rect 3488 8645 3491 8653
rect 3493 8645 3494 8653
rect 3511 8645 3512 8653
rect 3514 8645 3515 8653
rect 3527 8645 3528 8653
rect 3530 8649 3531 8653
rect 3530 8645 3535 8649
rect 3543 8645 3544 8653
rect 3546 8645 3549 8653
rect 3551 8645 3552 8653
rect 3564 8645 3565 8653
rect 3567 8645 3568 8653
rect 3580 8645 3581 8653
rect 3583 8645 3586 8653
rect 3588 8645 3589 8653
rect 3601 8645 3602 8653
rect 3604 8649 3605 8653
rect 3604 8645 3609 8649
rect 3617 8645 3618 8653
rect 3620 8645 3623 8653
rect 3625 8645 3626 8653
rect 3643 8645 3644 8653
rect 3646 8645 3647 8653
rect 3659 8645 3660 8653
rect 3662 8649 3663 8653
rect 3662 8645 3667 8649
rect 3675 8645 3676 8653
rect 3678 8645 3681 8653
rect 3683 8645 3684 8653
rect 3696 8645 3697 8653
rect 3699 8645 3700 8653
rect 3154 8589 3155 8597
rect 3157 8589 3160 8597
rect 3162 8589 3163 8597
rect 3175 8589 3176 8597
rect 3178 8593 3179 8597
rect 3178 8589 3183 8593
rect 3191 8589 3192 8597
rect 3194 8589 3197 8597
rect 3199 8589 3200 8597
rect 3217 8589 3218 8597
rect 3220 8589 3221 8597
rect 3233 8589 3234 8597
rect 3236 8593 3237 8597
rect 3236 8589 3241 8593
rect 3249 8589 3250 8597
rect 3252 8589 3255 8597
rect 3257 8589 3258 8597
rect 3270 8589 3271 8597
rect 3273 8589 3274 8597
rect 4099 8589 4100 8597
rect 4102 8589 4105 8597
rect 4107 8589 4108 8597
rect 4120 8589 4121 8597
rect 4123 8593 4124 8597
rect 4123 8589 4128 8593
rect 4136 8589 4137 8597
rect 4139 8589 4142 8597
rect 4144 8589 4145 8597
rect 4162 8589 4163 8597
rect 4165 8589 4166 8597
rect 4178 8589 4179 8597
rect 4181 8593 4182 8597
rect 4181 8589 4186 8593
rect 4194 8589 4195 8597
rect 4197 8589 4200 8597
rect 4202 8589 4203 8597
rect 4215 8589 4216 8597
rect 4218 8589 4219 8597
rect 2371 8559 2372 8567
rect 2374 8559 2377 8567
rect 2379 8559 2380 8567
rect 2392 8559 2393 8567
rect 2395 8563 2396 8567
rect 2395 8559 2400 8563
rect 2408 8559 2409 8567
rect 2411 8559 2414 8567
rect 2416 8559 2417 8567
rect 2434 8559 2435 8567
rect 2437 8559 2438 8567
rect 2450 8559 2451 8567
rect 2453 8563 2454 8567
rect 2453 8559 2458 8563
rect 2466 8559 2467 8567
rect 2469 8559 2472 8567
rect 2474 8559 2475 8567
rect 2487 8559 2488 8567
rect 2490 8559 2491 8567
rect 2503 8559 2504 8567
rect 2506 8559 2509 8567
rect 2511 8559 2512 8567
rect 2524 8559 2525 8567
rect 2527 8563 2528 8567
rect 2527 8559 2532 8563
rect 2540 8559 2541 8567
rect 2543 8559 2546 8567
rect 2548 8559 2549 8567
rect 2566 8559 2567 8567
rect 2569 8559 2570 8567
rect 2582 8559 2583 8567
rect 2585 8563 2586 8567
rect 2585 8559 2590 8563
rect 2598 8559 2599 8567
rect 2601 8559 2604 8567
rect 2606 8559 2607 8567
rect 2619 8559 2620 8567
rect 2622 8559 2623 8567
rect 2635 8559 2636 8567
rect 2638 8559 2641 8567
rect 2643 8559 2644 8567
rect 2656 8559 2657 8567
rect 2659 8563 2660 8567
rect 2659 8559 2664 8563
rect 2672 8559 2673 8567
rect 2675 8559 2678 8567
rect 2680 8559 2681 8567
rect 2698 8559 2699 8567
rect 2701 8559 2702 8567
rect 2714 8559 2715 8567
rect 2717 8563 2718 8567
rect 2717 8559 2722 8563
rect 2730 8559 2731 8567
rect 2733 8559 2736 8567
rect 2738 8559 2739 8567
rect 2751 8559 2752 8567
rect 2754 8559 2755 8567
rect 3316 8559 3317 8567
rect 3319 8559 3322 8567
rect 3324 8559 3325 8567
rect 3337 8559 3338 8567
rect 3340 8563 3341 8567
rect 3340 8559 3345 8563
rect 3353 8559 3354 8567
rect 3356 8559 3359 8567
rect 3361 8559 3362 8567
rect 3379 8559 3380 8567
rect 3382 8559 3383 8567
rect 3395 8559 3396 8567
rect 3398 8563 3399 8567
rect 3398 8559 3403 8563
rect 3411 8559 3412 8567
rect 3414 8559 3417 8567
rect 3419 8559 3420 8567
rect 3432 8559 3433 8567
rect 3435 8559 3436 8567
rect 3448 8559 3449 8567
rect 3451 8559 3454 8567
rect 3456 8559 3457 8567
rect 3469 8559 3470 8567
rect 3472 8563 3473 8567
rect 3472 8559 3477 8563
rect 3485 8559 3486 8567
rect 3488 8559 3491 8567
rect 3493 8559 3494 8567
rect 3511 8559 3512 8567
rect 3514 8559 3515 8567
rect 3527 8559 3528 8567
rect 3530 8563 3531 8567
rect 3530 8559 3535 8563
rect 3543 8559 3544 8567
rect 3546 8559 3549 8567
rect 3551 8559 3552 8567
rect 3564 8559 3565 8567
rect 3567 8559 3568 8567
rect 3580 8559 3581 8567
rect 3583 8559 3586 8567
rect 3588 8559 3589 8567
rect 3601 8559 3602 8567
rect 3604 8563 3605 8567
rect 3604 8559 3609 8563
rect 3617 8559 3618 8567
rect 3620 8559 3623 8567
rect 3625 8559 3626 8567
rect 3643 8559 3644 8567
rect 3646 8559 3647 8567
rect 3659 8559 3660 8567
rect 3662 8563 3663 8567
rect 3662 8559 3667 8563
rect 3675 8559 3676 8567
rect 3678 8559 3681 8567
rect 3683 8559 3684 8567
rect 3696 8559 3697 8567
rect 3699 8559 3700 8567
rect 2371 8419 2372 8427
rect 2374 8419 2377 8427
rect 2379 8419 2380 8427
rect 2392 8419 2393 8427
rect 2395 8423 2396 8427
rect 2395 8419 2400 8423
rect 2408 8419 2409 8427
rect 2411 8419 2414 8427
rect 2416 8419 2417 8427
rect 2434 8419 2435 8427
rect 2437 8419 2438 8427
rect 2450 8419 2451 8427
rect 2453 8423 2454 8427
rect 2453 8419 2458 8423
rect 2466 8419 2467 8427
rect 2469 8419 2472 8427
rect 2474 8419 2475 8427
rect 2487 8419 2488 8427
rect 2490 8419 2491 8427
rect 2503 8419 2504 8427
rect 2506 8419 2509 8427
rect 2511 8419 2512 8427
rect 2524 8419 2525 8427
rect 2527 8423 2528 8427
rect 2527 8419 2532 8423
rect 2540 8419 2541 8427
rect 2543 8419 2546 8427
rect 2548 8419 2549 8427
rect 2566 8419 2567 8427
rect 2569 8419 2570 8427
rect 2582 8419 2583 8427
rect 2585 8423 2586 8427
rect 2585 8419 2590 8423
rect 2598 8419 2599 8427
rect 2601 8419 2604 8427
rect 2606 8419 2607 8427
rect 2619 8419 2620 8427
rect 2622 8419 2623 8427
rect 2635 8419 2636 8427
rect 2638 8419 2641 8427
rect 2643 8419 2644 8427
rect 2656 8419 2657 8427
rect 2659 8423 2660 8427
rect 2659 8419 2664 8423
rect 2672 8419 2673 8427
rect 2675 8419 2678 8427
rect 2680 8419 2681 8427
rect 2698 8419 2699 8427
rect 2701 8419 2702 8427
rect 2714 8419 2715 8427
rect 2717 8423 2718 8427
rect 2717 8419 2722 8423
rect 2730 8419 2731 8427
rect 2733 8419 2736 8427
rect 2738 8419 2739 8427
rect 2751 8419 2752 8427
rect 2754 8419 2755 8427
rect 3316 8419 3317 8427
rect 3319 8419 3322 8427
rect 3324 8419 3325 8427
rect 3337 8419 3338 8427
rect 3340 8423 3341 8427
rect 3340 8419 3345 8423
rect 3353 8419 3354 8427
rect 3356 8419 3359 8427
rect 3361 8419 3362 8427
rect 3379 8419 3380 8427
rect 3382 8419 3383 8427
rect 3395 8419 3396 8427
rect 3398 8423 3399 8427
rect 3398 8419 3403 8423
rect 3411 8419 3412 8427
rect 3414 8419 3417 8427
rect 3419 8419 3420 8427
rect 3432 8419 3433 8427
rect 3435 8419 3436 8427
rect 3448 8419 3449 8427
rect 3451 8419 3454 8427
rect 3456 8419 3457 8427
rect 3469 8419 3470 8427
rect 3472 8423 3473 8427
rect 3472 8419 3477 8423
rect 3485 8419 3486 8427
rect 3488 8419 3491 8427
rect 3493 8419 3494 8427
rect 3511 8419 3512 8427
rect 3514 8419 3515 8427
rect 3527 8419 3528 8427
rect 3530 8423 3531 8427
rect 3530 8419 3535 8423
rect 3543 8419 3544 8427
rect 3546 8419 3549 8427
rect 3551 8419 3552 8427
rect 3564 8419 3565 8427
rect 3567 8419 3568 8427
rect 3580 8419 3581 8427
rect 3583 8419 3586 8427
rect 3588 8419 3589 8427
rect 3601 8419 3602 8427
rect 3604 8423 3605 8427
rect 3604 8419 3609 8423
rect 3617 8419 3618 8427
rect 3620 8419 3623 8427
rect 3625 8419 3626 8427
rect 3643 8419 3644 8427
rect 3646 8419 3647 8427
rect 3659 8419 3660 8427
rect 3662 8423 3663 8427
rect 3662 8419 3667 8423
rect 3675 8419 3676 8427
rect 3678 8419 3681 8427
rect 3683 8419 3684 8427
rect 3696 8419 3697 8427
rect 3699 8419 3700 8427
rect 2855 8340 2856 8348
rect 2858 8340 2861 8348
rect 2863 8340 2864 8348
rect 2876 8340 2877 8348
rect 2879 8344 2880 8348
rect 2879 8340 2884 8344
rect 2892 8340 2893 8348
rect 2895 8340 2898 8348
rect 2900 8340 2901 8348
rect 2918 8340 2919 8348
rect 2921 8340 2922 8348
rect 2934 8340 2935 8348
rect 2937 8344 2938 8348
rect 2937 8340 2942 8344
rect 2950 8340 2951 8348
rect 2953 8340 2956 8348
rect 2958 8340 2959 8348
rect 2971 8340 2972 8348
rect 2974 8340 2975 8348
rect 2987 8340 2988 8348
rect 2990 8340 2993 8348
rect 2995 8340 2996 8348
rect 3008 8340 3009 8348
rect 3011 8344 3012 8348
rect 3011 8340 3016 8344
rect 3024 8340 3025 8348
rect 3027 8340 3030 8348
rect 3032 8340 3033 8348
rect 3050 8340 3051 8348
rect 3053 8340 3054 8348
rect 3066 8340 3067 8348
rect 3069 8344 3070 8348
rect 3069 8340 3074 8344
rect 3082 8340 3083 8348
rect 3085 8340 3088 8348
rect 3090 8340 3091 8348
rect 3103 8340 3104 8348
rect 3106 8340 3107 8348
rect 3119 8340 3120 8348
rect 3122 8340 3125 8348
rect 3127 8340 3128 8348
rect 3140 8340 3141 8348
rect 3143 8344 3144 8348
rect 3143 8340 3148 8344
rect 3156 8340 3157 8348
rect 3159 8340 3162 8348
rect 3164 8340 3165 8348
rect 3182 8340 3183 8348
rect 3185 8340 3186 8348
rect 3198 8340 3199 8348
rect 3201 8344 3202 8348
rect 3201 8340 3206 8344
rect 3214 8340 3215 8348
rect 3217 8340 3220 8348
rect 3222 8340 3223 8348
rect 3235 8340 3236 8348
rect 3238 8340 3239 8348
rect 3251 8340 3252 8348
rect 3254 8340 3257 8348
rect 3259 8340 3260 8348
rect 3272 8340 3273 8348
rect 3275 8344 3276 8348
rect 3275 8340 3280 8344
rect 3288 8340 3289 8348
rect 3291 8340 3294 8348
rect 3296 8340 3297 8348
rect 3314 8340 3315 8348
rect 3317 8340 3318 8348
rect 3330 8340 3331 8348
rect 3333 8344 3334 8348
rect 3333 8340 3338 8344
rect 3346 8340 3347 8348
rect 3349 8340 3352 8348
rect 3354 8340 3355 8348
rect 3367 8340 3368 8348
rect 3370 8340 3371 8348
rect 3800 8340 3801 8348
rect 3803 8340 3806 8348
rect 3808 8340 3809 8348
rect 3821 8340 3822 8348
rect 3824 8344 3825 8348
rect 3824 8340 3829 8344
rect 3837 8340 3838 8348
rect 3840 8340 3843 8348
rect 3845 8340 3846 8348
rect 3863 8340 3864 8348
rect 3866 8340 3867 8348
rect 3879 8340 3880 8348
rect 3882 8344 3883 8348
rect 3882 8340 3887 8344
rect 3895 8340 3896 8348
rect 3898 8340 3901 8348
rect 3903 8340 3904 8348
rect 3916 8340 3917 8348
rect 3919 8340 3920 8348
rect 3932 8340 3933 8348
rect 3935 8340 3938 8348
rect 3940 8340 3941 8348
rect 3953 8340 3954 8348
rect 3956 8344 3957 8348
rect 3956 8340 3961 8344
rect 3969 8340 3970 8348
rect 3972 8340 3975 8348
rect 3977 8340 3978 8348
rect 3995 8340 3996 8348
rect 3998 8340 3999 8348
rect 4011 8340 4012 8348
rect 4014 8344 4015 8348
rect 4014 8340 4019 8344
rect 4027 8340 4028 8348
rect 4030 8340 4033 8348
rect 4035 8340 4036 8348
rect 4048 8340 4049 8348
rect 4051 8340 4052 8348
rect 4064 8340 4065 8348
rect 4067 8340 4070 8348
rect 4072 8340 4073 8348
rect 4085 8340 4086 8348
rect 4088 8344 4089 8348
rect 4088 8340 4093 8344
rect 4101 8340 4102 8348
rect 4104 8340 4107 8348
rect 4109 8340 4110 8348
rect 4127 8340 4128 8348
rect 4130 8340 4131 8348
rect 4143 8340 4144 8348
rect 4146 8344 4147 8348
rect 4146 8340 4151 8344
rect 4159 8340 4160 8348
rect 4162 8340 4165 8348
rect 4167 8340 4168 8348
rect 4180 8340 4181 8348
rect 4183 8340 4184 8348
rect 4196 8340 4197 8348
rect 4199 8340 4202 8348
rect 4204 8340 4205 8348
rect 4217 8340 4218 8348
rect 4220 8344 4221 8348
rect 4220 8340 4225 8344
rect 4233 8340 4234 8348
rect 4236 8340 4239 8348
rect 4241 8340 4242 8348
rect 4259 8340 4260 8348
rect 4262 8340 4263 8348
rect 4275 8340 4276 8348
rect 4278 8344 4279 8348
rect 4278 8340 4283 8344
rect 4291 8340 4292 8348
rect 4294 8340 4297 8348
rect 4299 8340 4300 8348
rect 4312 8340 4313 8348
rect 4315 8340 4316 8348
rect 2503 8307 2504 8315
rect 2506 8307 2509 8315
rect 2511 8307 2512 8315
rect 2524 8307 2525 8315
rect 2527 8311 2528 8315
rect 2527 8307 2532 8311
rect 2540 8307 2541 8315
rect 2543 8307 2546 8315
rect 2548 8307 2549 8315
rect 2566 8307 2567 8315
rect 2569 8307 2570 8315
rect 2582 8307 2583 8315
rect 2585 8311 2586 8315
rect 2585 8307 2590 8311
rect 2598 8307 2599 8315
rect 2601 8307 2604 8315
rect 2606 8307 2607 8315
rect 2619 8307 2620 8315
rect 2622 8307 2623 8315
rect 3448 8307 3449 8315
rect 3451 8307 3454 8315
rect 3456 8307 3457 8315
rect 3469 8307 3470 8315
rect 3472 8311 3473 8315
rect 3472 8307 3477 8311
rect 3485 8307 3486 8315
rect 3488 8307 3491 8315
rect 3493 8307 3494 8315
rect 3511 8307 3512 8315
rect 3514 8307 3515 8315
rect 3527 8307 3528 8315
rect 3530 8311 3531 8315
rect 3530 8307 3535 8311
rect 3543 8307 3544 8315
rect 3546 8307 3549 8315
rect 3551 8307 3552 8315
rect 3564 8307 3565 8315
rect 3567 8307 3568 8315
rect 3034 8269 3035 8277
rect 3037 8269 3038 8277
rect 2860 8256 2861 8264
rect 2863 8256 2864 8264
rect 2876 8256 2877 8264
rect 2879 8256 2880 8264
rect 2892 8256 2893 8264
rect 2895 8256 2896 8264
rect 2911 8256 2916 8264
rect 2918 8256 2921 8264
rect 2923 8256 2924 8264
rect 2945 8256 2947 8264
rect 2949 8256 2950 8264
rect 2967 8256 2968 8264
rect 2970 8256 2971 8264
rect 2983 8256 2988 8264
rect 2990 8256 2993 8264
rect 2995 8256 2996 8264
rect 3010 8256 3011 8264
rect 3013 8256 3014 8264
rect 3058 8263 3061 8271
rect 3063 8263 3066 8271
rect 3068 8263 3069 8271
rect 3088 8269 3089 8277
rect 3091 8269 3092 8277
rect 3115 8269 3116 8277
rect 3118 8269 3119 8277
rect 3139 8263 3142 8271
rect 3144 8263 3147 8271
rect 3149 8263 3150 8271
rect 3169 8269 3170 8277
rect 3172 8269 3173 8277
rect 3979 8269 3980 8277
rect 3982 8269 3983 8277
rect 3805 8256 3806 8264
rect 3808 8256 3809 8264
rect 3821 8256 3822 8264
rect 3824 8256 3825 8264
rect 3837 8256 3838 8264
rect 3840 8256 3841 8264
rect 3856 8256 3861 8264
rect 3863 8256 3866 8264
rect 3868 8256 3869 8264
rect 3890 8256 3892 8264
rect 3894 8256 3895 8264
rect 3912 8256 3913 8264
rect 3915 8256 3916 8264
rect 3928 8256 3933 8264
rect 3935 8256 3938 8264
rect 3940 8256 3941 8264
rect 3955 8256 3956 8264
rect 3958 8256 3959 8264
rect 4003 8263 4006 8271
rect 4008 8263 4011 8271
rect 4013 8263 4014 8271
rect 4033 8269 4034 8277
rect 4036 8269 4037 8277
rect 4060 8269 4061 8277
rect 4063 8269 4064 8277
rect 4084 8263 4087 8271
rect 4089 8263 4092 8271
rect 4094 8263 4095 8271
rect 4114 8269 4115 8277
rect 4117 8269 4118 8277
rect 2494 8205 2495 8213
rect 2497 8205 2498 8213
rect 2510 8205 2511 8213
rect 2513 8205 2516 8213
rect 2518 8205 2519 8213
rect 2531 8209 2532 8213
rect 2527 8205 2532 8209
rect 2534 8205 2535 8213
rect 2547 8205 2548 8213
rect 2550 8205 2551 8213
rect 2568 8205 2569 8213
rect 2571 8205 2574 8213
rect 2576 8205 2577 8213
rect 2589 8209 2590 8213
rect 2585 8205 2590 8209
rect 2592 8205 2593 8213
rect 2605 8205 2606 8213
rect 2608 8205 2611 8213
rect 2613 8205 2614 8213
rect 3439 8205 3440 8213
rect 3442 8205 3443 8213
rect 3455 8205 3456 8213
rect 3458 8205 3461 8213
rect 3463 8205 3464 8213
rect 3476 8209 3477 8213
rect 3472 8205 3477 8209
rect 3479 8205 3480 8213
rect 3492 8205 3493 8213
rect 3495 8205 3496 8213
rect 3513 8205 3514 8213
rect 3516 8205 3519 8213
rect 3521 8205 3522 8213
rect 3534 8209 3535 8213
rect 3530 8205 3535 8209
rect 3537 8205 3538 8213
rect 3550 8205 3551 8213
rect 3553 8205 3556 8213
rect 3558 8205 3559 8213
rect 2860 8170 2861 8178
rect 2863 8170 2864 8178
rect 2876 8170 2877 8178
rect 2879 8170 2880 8178
rect 2892 8170 2893 8178
rect 2895 8170 2896 8178
rect 2911 8170 2916 8178
rect 2918 8170 2921 8178
rect 2923 8170 2924 8178
rect 2945 8170 2947 8178
rect 2949 8170 2950 8178
rect 2967 8170 2968 8178
rect 2970 8170 2971 8178
rect 2983 8170 2988 8178
rect 2990 8170 2993 8178
rect 2995 8170 2996 8178
rect 3010 8170 3011 8178
rect 3013 8170 3014 8178
rect 3058 8171 3061 8179
rect 3063 8171 3066 8179
rect 3068 8171 3069 8179
rect 3139 8171 3142 8179
rect 3144 8171 3147 8179
rect 3149 8171 3150 8179
rect 3805 8170 3806 8178
rect 3808 8170 3809 8178
rect 3821 8170 3822 8178
rect 3824 8170 3825 8178
rect 3837 8170 3838 8178
rect 3840 8170 3841 8178
rect 3856 8170 3861 8178
rect 3863 8170 3866 8178
rect 3868 8170 3869 8178
rect 3890 8170 3892 8178
rect 3894 8170 3895 8178
rect 3912 8170 3913 8178
rect 3915 8170 3916 8178
rect 3928 8170 3933 8178
rect 3935 8170 3938 8178
rect 3940 8170 3941 8178
rect 3955 8170 3956 8178
rect 3958 8170 3959 8178
rect 4003 8171 4006 8179
rect 4008 8171 4011 8179
rect 4013 8171 4014 8179
rect 4084 8171 4087 8179
rect 4089 8171 4092 8179
rect 4094 8171 4095 8179
rect 2860 8124 2861 8132
rect 2863 8124 2864 8132
rect 2876 8124 2877 8132
rect 2879 8124 2880 8132
rect 2892 8124 2893 8132
rect 2895 8124 2896 8132
rect 2911 8124 2916 8132
rect 2918 8124 2921 8132
rect 2923 8124 2924 8132
rect 2945 8124 2947 8132
rect 2949 8124 2950 8132
rect 2967 8124 2968 8132
rect 2970 8124 2971 8132
rect 2983 8124 2988 8132
rect 2990 8124 2993 8132
rect 2995 8124 2996 8132
rect 3010 8124 3011 8132
rect 3013 8124 3014 8132
rect 3058 8131 3061 8139
rect 3063 8131 3066 8139
rect 3068 8131 3069 8139
rect 3088 8137 3089 8145
rect 3091 8137 3092 8145
rect 3139 8137 3140 8145
rect 3142 8137 3143 8145
rect 3163 8131 3166 8139
rect 3168 8131 3171 8139
rect 3173 8131 3174 8139
rect 3193 8137 3194 8145
rect 3196 8137 3197 8145
rect 3805 8124 3806 8132
rect 3808 8124 3809 8132
rect 3821 8124 3822 8132
rect 3824 8124 3825 8132
rect 3837 8124 3838 8132
rect 3840 8124 3841 8132
rect 3856 8124 3861 8132
rect 3863 8124 3866 8132
rect 3868 8124 3869 8132
rect 3890 8124 3892 8132
rect 3894 8124 3895 8132
rect 3912 8124 3913 8132
rect 3915 8124 3916 8132
rect 3928 8124 3933 8132
rect 3935 8124 3938 8132
rect 3940 8124 3941 8132
rect 3955 8124 3956 8132
rect 3958 8124 3959 8132
rect 4003 8131 4006 8139
rect 4008 8131 4011 8139
rect 4013 8131 4014 8139
rect 4033 8137 4034 8145
rect 4036 8137 4037 8145
rect 4084 8137 4085 8145
rect 4087 8137 4088 8145
rect 4108 8131 4111 8139
rect 4113 8131 4116 8139
rect 4118 8131 4119 8139
rect 4138 8137 4139 8145
rect 4141 8137 4142 8145
rect 2860 8038 2861 8046
rect 2863 8038 2864 8046
rect 2876 8038 2877 8046
rect 2879 8038 2880 8046
rect 2892 8038 2893 8046
rect 2895 8038 2896 8046
rect 2911 8038 2916 8046
rect 2918 8038 2921 8046
rect 2923 8038 2924 8046
rect 2945 8038 2947 8046
rect 2949 8038 2950 8046
rect 2967 8038 2968 8046
rect 2970 8038 2971 8046
rect 2983 8038 2988 8046
rect 2990 8038 2993 8046
rect 2995 8038 2996 8046
rect 3010 8038 3011 8046
rect 3013 8038 3014 8046
rect 3058 8040 3061 8048
rect 3063 8040 3066 8048
rect 3068 8040 3069 8048
rect 3163 8040 3166 8048
rect 3168 8040 3171 8048
rect 3173 8040 3174 8048
rect 3805 8038 3806 8046
rect 3808 8038 3809 8046
rect 3821 8038 3822 8046
rect 3824 8038 3825 8046
rect 3837 8038 3838 8046
rect 3840 8038 3841 8046
rect 3856 8038 3861 8046
rect 3863 8038 3866 8046
rect 3868 8038 3869 8046
rect 3890 8038 3892 8046
rect 3894 8038 3895 8046
rect 3912 8038 3913 8046
rect 3915 8038 3916 8046
rect 3928 8038 3933 8046
rect 3935 8038 3938 8046
rect 3940 8038 3941 8046
rect 3955 8038 3956 8046
rect 3958 8038 3959 8046
rect 4003 8040 4006 8048
rect 4008 8040 4011 8048
rect 4013 8040 4014 8048
rect 4108 8040 4111 8048
rect 4113 8040 4116 8048
rect 4118 8040 4119 8048
rect 2860 7992 2861 8000
rect 2863 7992 2864 8000
rect 2876 7992 2877 8000
rect 2879 7992 2880 8000
rect 2892 7992 2893 8000
rect 2895 7992 2896 8000
rect 2911 7992 2916 8000
rect 2918 7992 2921 8000
rect 2923 7992 2924 8000
rect 2945 7992 2947 8000
rect 2949 7992 2950 8000
rect 2967 7992 2968 8000
rect 2970 7992 2971 8000
rect 2983 7992 2988 8000
rect 2990 7992 2993 8000
rect 2995 7992 2996 8000
rect 3010 7992 3011 8000
rect 3013 7992 3014 8000
rect 3058 7999 3061 8007
rect 3063 7999 3066 8007
rect 3068 7999 3069 8007
rect 3088 8005 3089 8013
rect 3091 8005 3092 8013
rect 3115 8005 3116 8013
rect 3118 8005 3119 8013
rect 3139 7999 3142 8007
rect 3144 7999 3147 8007
rect 3149 7999 3150 8007
rect 3169 8005 3170 8013
rect 3172 8005 3173 8013
rect 3205 8005 3206 8013
rect 3208 8005 3209 8013
rect 3229 7999 3232 8007
rect 3234 7999 3237 8007
rect 3239 7999 3240 8007
rect 3259 8005 3260 8013
rect 3262 8005 3263 8013
rect 3805 7992 3806 8000
rect 3808 7992 3809 8000
rect 3821 7992 3822 8000
rect 3824 7992 3825 8000
rect 3837 7992 3838 8000
rect 3840 7992 3841 8000
rect 3856 7992 3861 8000
rect 3863 7992 3866 8000
rect 3868 7992 3869 8000
rect 3890 7992 3892 8000
rect 3894 7992 3895 8000
rect 3912 7992 3913 8000
rect 3915 7992 3916 8000
rect 3928 7992 3933 8000
rect 3935 7992 3938 8000
rect 3940 7992 3941 8000
rect 3955 7992 3956 8000
rect 3958 7992 3959 8000
rect 4003 7999 4006 8007
rect 4008 7999 4011 8007
rect 4013 7999 4014 8007
rect 4033 8005 4034 8013
rect 4036 8005 4037 8013
rect 4060 8005 4061 8013
rect 4063 8005 4064 8013
rect 4084 7999 4087 8007
rect 4089 7999 4092 8007
rect 4094 7999 4095 8007
rect 4114 8005 4115 8013
rect 4117 8005 4118 8013
rect 4150 8005 4151 8013
rect 4153 8005 4154 8013
rect 4174 7999 4177 8007
rect 4179 7999 4182 8007
rect 4184 7999 4185 8007
rect 4204 8005 4205 8013
rect 4207 8005 4208 8013
rect 2860 7906 2861 7914
rect 2863 7906 2864 7914
rect 2876 7906 2877 7914
rect 2879 7906 2880 7914
rect 2892 7906 2893 7914
rect 2895 7906 2896 7914
rect 2911 7906 2916 7914
rect 2918 7906 2921 7914
rect 2923 7906 2924 7914
rect 2945 7906 2947 7914
rect 2949 7906 2950 7914
rect 2967 7906 2968 7914
rect 2970 7906 2971 7914
rect 2983 7906 2988 7914
rect 2990 7906 2993 7914
rect 2995 7906 2996 7914
rect 3010 7906 3011 7914
rect 3013 7906 3014 7914
rect 3058 7905 3061 7913
rect 3063 7905 3066 7913
rect 3068 7905 3069 7913
rect 3139 7905 3142 7913
rect 3144 7905 3147 7913
rect 3149 7905 3150 7913
rect 3229 7905 3232 7913
rect 3234 7905 3237 7913
rect 3239 7905 3240 7913
rect 3805 7906 3806 7914
rect 3808 7906 3809 7914
rect 3821 7906 3822 7914
rect 3824 7906 3825 7914
rect 3837 7906 3838 7914
rect 3840 7906 3841 7914
rect 3856 7906 3861 7914
rect 3863 7906 3866 7914
rect 3868 7906 3869 7914
rect 3890 7906 3892 7914
rect 3894 7906 3895 7914
rect 3912 7906 3913 7914
rect 3915 7906 3916 7914
rect 3928 7906 3933 7914
rect 3935 7906 3938 7914
rect 3940 7906 3941 7914
rect 3955 7906 3956 7914
rect 3958 7906 3959 7914
rect 4003 7905 4006 7913
rect 4008 7905 4011 7913
rect 4013 7905 4014 7913
rect 4084 7905 4087 7913
rect 4089 7905 4092 7913
rect 4094 7905 4095 7913
rect 4174 7905 4177 7913
rect 4179 7905 4182 7913
rect 4184 7905 4185 7913
rect 2860 7860 2861 7868
rect 2863 7860 2864 7868
rect 2876 7860 2877 7868
rect 2879 7860 2880 7868
rect 2892 7860 2893 7868
rect 2895 7860 2896 7868
rect 2911 7860 2916 7868
rect 2918 7860 2921 7868
rect 2923 7860 2924 7868
rect 2945 7860 2947 7868
rect 2949 7860 2950 7868
rect 2967 7860 2968 7868
rect 2970 7860 2971 7868
rect 2983 7860 2988 7868
rect 2990 7860 2993 7868
rect 2995 7860 2996 7868
rect 3010 7860 3011 7868
rect 3013 7860 3014 7868
rect 3058 7867 3061 7875
rect 3063 7867 3066 7875
rect 3068 7867 3069 7875
rect 3088 7873 3089 7881
rect 3091 7873 3092 7881
rect 3805 7860 3806 7868
rect 3808 7860 3809 7868
rect 3821 7860 3822 7868
rect 3824 7860 3825 7868
rect 3837 7860 3838 7868
rect 3840 7860 3841 7868
rect 3856 7860 3861 7868
rect 3863 7860 3866 7868
rect 3868 7860 3869 7868
rect 3890 7860 3892 7868
rect 3894 7860 3895 7868
rect 3912 7860 3913 7868
rect 3915 7860 3916 7868
rect 3928 7860 3933 7868
rect 3935 7860 3938 7868
rect 3940 7860 3941 7868
rect 3955 7860 3956 7868
rect 3958 7860 3959 7868
rect 4003 7867 4006 7875
rect 4008 7867 4011 7875
rect 4013 7867 4014 7875
rect 4033 7873 4034 7881
rect 4036 7873 4037 7881
rect 2371 7805 2372 7813
rect 2374 7805 2377 7813
rect 2379 7805 2380 7813
rect 2392 7805 2393 7813
rect 2395 7809 2396 7813
rect 2395 7805 2400 7809
rect 2408 7805 2409 7813
rect 2411 7805 2414 7813
rect 2416 7805 2417 7813
rect 2434 7805 2435 7813
rect 2437 7805 2438 7813
rect 2450 7805 2451 7813
rect 2453 7809 2454 7813
rect 2453 7805 2458 7809
rect 2466 7805 2467 7813
rect 2469 7805 2472 7813
rect 2474 7805 2475 7813
rect 2487 7805 2488 7813
rect 2490 7805 2491 7813
rect 2503 7805 2504 7813
rect 2506 7805 2509 7813
rect 2511 7805 2512 7813
rect 2524 7805 2525 7813
rect 2527 7809 2528 7813
rect 2527 7805 2532 7809
rect 2540 7805 2541 7813
rect 2543 7805 2546 7813
rect 2548 7805 2549 7813
rect 2566 7805 2567 7813
rect 2569 7805 2570 7813
rect 2582 7805 2583 7813
rect 2585 7809 2586 7813
rect 2585 7805 2590 7809
rect 2598 7805 2599 7813
rect 2601 7805 2604 7813
rect 2606 7805 2607 7813
rect 2619 7805 2620 7813
rect 2622 7805 2623 7813
rect 2635 7805 2636 7813
rect 2638 7805 2641 7813
rect 2643 7805 2644 7813
rect 2656 7805 2657 7813
rect 2659 7809 2660 7813
rect 2659 7805 2664 7809
rect 2672 7805 2673 7813
rect 2675 7805 2678 7813
rect 2680 7805 2681 7813
rect 2698 7805 2699 7813
rect 2701 7805 2702 7813
rect 2714 7805 2715 7813
rect 2717 7809 2718 7813
rect 2717 7805 2722 7809
rect 2730 7805 2731 7813
rect 2733 7805 2736 7813
rect 2738 7805 2739 7813
rect 2751 7805 2752 7813
rect 2754 7805 2755 7813
rect 3316 7805 3317 7813
rect 3319 7805 3322 7813
rect 3324 7805 3325 7813
rect 3337 7805 3338 7813
rect 3340 7809 3341 7813
rect 3340 7805 3345 7809
rect 3353 7805 3354 7813
rect 3356 7805 3359 7813
rect 3361 7805 3362 7813
rect 3379 7805 3380 7813
rect 3382 7805 3383 7813
rect 3395 7805 3396 7813
rect 3398 7809 3399 7813
rect 3398 7805 3403 7809
rect 3411 7805 3412 7813
rect 3414 7805 3417 7813
rect 3419 7805 3420 7813
rect 3432 7805 3433 7813
rect 3435 7805 3436 7813
rect 3448 7805 3449 7813
rect 3451 7805 3454 7813
rect 3456 7805 3457 7813
rect 3469 7805 3470 7813
rect 3472 7809 3473 7813
rect 3472 7805 3477 7809
rect 3485 7805 3486 7813
rect 3488 7805 3491 7813
rect 3493 7805 3494 7813
rect 3511 7805 3512 7813
rect 3514 7805 3515 7813
rect 3527 7805 3528 7813
rect 3530 7809 3531 7813
rect 3530 7805 3535 7809
rect 3543 7805 3544 7813
rect 3546 7805 3549 7813
rect 3551 7805 3552 7813
rect 3564 7805 3565 7813
rect 3567 7805 3568 7813
rect 3580 7805 3581 7813
rect 3583 7805 3586 7813
rect 3588 7805 3589 7813
rect 3601 7805 3602 7813
rect 3604 7809 3605 7813
rect 3604 7805 3609 7809
rect 3617 7805 3618 7813
rect 3620 7805 3623 7813
rect 3625 7805 3626 7813
rect 3643 7805 3644 7813
rect 3646 7805 3647 7813
rect 3659 7805 3660 7813
rect 3662 7809 3663 7813
rect 3662 7805 3667 7809
rect 3675 7805 3676 7813
rect 3678 7805 3681 7813
rect 3683 7805 3684 7813
rect 3696 7805 3697 7813
rect 3699 7805 3700 7813
rect 2860 7774 2861 7782
rect 2863 7774 2864 7782
rect 2876 7774 2877 7782
rect 2879 7774 2880 7782
rect 2892 7774 2893 7782
rect 2895 7774 2896 7782
rect 2911 7774 2916 7782
rect 2918 7774 2921 7782
rect 2923 7774 2924 7782
rect 2945 7774 2947 7782
rect 2949 7774 2950 7782
rect 2967 7774 2968 7782
rect 2970 7774 2971 7782
rect 2983 7774 2988 7782
rect 2990 7774 2993 7782
rect 2995 7774 2996 7782
rect 3010 7774 3011 7782
rect 3013 7774 3014 7782
rect 3058 7769 3061 7777
rect 3063 7769 3066 7777
rect 3068 7769 3069 7777
rect 3094 7774 3095 7782
rect 3097 7774 3098 7782
rect 3102 7774 3108 7782
rect 3112 7774 3113 7782
rect 3115 7774 3116 7782
rect 3137 7774 3138 7782
rect 3140 7774 3141 7782
rect 3153 7774 3154 7782
rect 3156 7774 3157 7782
rect 3172 7774 3177 7782
rect 3179 7774 3182 7782
rect 3184 7774 3185 7782
rect 3206 7774 3208 7782
rect 3210 7774 3211 7782
rect 3228 7774 3229 7782
rect 3231 7774 3232 7782
rect 3244 7774 3249 7782
rect 3251 7774 3254 7782
rect 3256 7774 3257 7782
rect 3271 7774 3272 7782
rect 3274 7774 3275 7782
rect 3805 7774 3806 7782
rect 3808 7774 3809 7782
rect 3821 7774 3822 7782
rect 3824 7774 3825 7782
rect 3837 7774 3838 7782
rect 3840 7774 3841 7782
rect 3856 7774 3861 7782
rect 3863 7774 3866 7782
rect 3868 7774 3869 7782
rect 3890 7774 3892 7782
rect 3894 7774 3895 7782
rect 3912 7774 3913 7782
rect 3915 7774 3916 7782
rect 3928 7774 3933 7782
rect 3935 7774 3938 7782
rect 3940 7774 3941 7782
rect 3955 7774 3956 7782
rect 3958 7774 3959 7782
rect 4003 7769 4006 7777
rect 4008 7769 4011 7777
rect 4013 7769 4014 7777
rect 4039 7774 4040 7782
rect 4042 7774 4043 7782
rect 4047 7774 4053 7782
rect 4057 7774 4058 7782
rect 4060 7774 4061 7782
rect 4082 7774 4083 7782
rect 4085 7774 4086 7782
rect 4098 7774 4099 7782
rect 4101 7774 4102 7782
rect 4117 7774 4122 7782
rect 4124 7774 4127 7782
rect 4129 7774 4130 7782
rect 4151 7774 4153 7782
rect 4155 7774 4156 7782
rect 4173 7774 4174 7782
rect 4176 7774 4177 7782
rect 4189 7774 4194 7782
rect 4196 7774 4199 7782
rect 4201 7774 4202 7782
rect 4216 7774 4217 7782
rect 4219 7774 4220 7782
rect 3154 7693 3155 7701
rect 3157 7693 3160 7701
rect 3162 7693 3163 7701
rect 3175 7693 3176 7701
rect 3178 7697 3179 7701
rect 3178 7693 3183 7697
rect 3191 7693 3192 7701
rect 3194 7693 3197 7701
rect 3199 7693 3200 7701
rect 3217 7693 3218 7701
rect 3220 7693 3221 7701
rect 3233 7693 3234 7701
rect 3236 7697 3237 7701
rect 3236 7693 3241 7697
rect 3249 7693 3250 7701
rect 3252 7693 3255 7701
rect 3257 7693 3258 7701
rect 3270 7693 3271 7701
rect 3273 7693 3274 7701
rect 4099 7693 4100 7701
rect 4102 7693 4105 7701
rect 4107 7693 4108 7701
rect 4120 7693 4121 7701
rect 4123 7697 4124 7701
rect 4123 7693 4128 7697
rect 4136 7693 4137 7701
rect 4139 7693 4142 7701
rect 4144 7693 4145 7701
rect 4162 7693 4163 7701
rect 4165 7693 4166 7701
rect 4178 7693 4179 7701
rect 4181 7697 4182 7701
rect 4181 7693 4186 7697
rect 4194 7693 4195 7701
rect 4197 7693 4200 7701
rect 4202 7693 4203 7701
rect 4215 7693 4216 7701
rect 4218 7693 4219 7701
rect 2371 7663 2372 7671
rect 2374 7663 2377 7671
rect 2379 7663 2380 7671
rect 2392 7663 2393 7671
rect 2395 7667 2396 7671
rect 2395 7663 2400 7667
rect 2408 7663 2409 7671
rect 2411 7663 2414 7671
rect 2416 7663 2417 7671
rect 2434 7663 2435 7671
rect 2437 7663 2438 7671
rect 2450 7663 2451 7671
rect 2453 7667 2454 7671
rect 2453 7663 2458 7667
rect 2466 7663 2467 7671
rect 2469 7663 2472 7671
rect 2474 7663 2475 7671
rect 2487 7663 2488 7671
rect 2490 7663 2491 7671
rect 2503 7663 2504 7671
rect 2506 7663 2509 7671
rect 2511 7663 2512 7671
rect 2524 7663 2525 7671
rect 2527 7667 2528 7671
rect 2527 7663 2532 7667
rect 2540 7663 2541 7671
rect 2543 7663 2546 7671
rect 2548 7663 2549 7671
rect 2566 7663 2567 7671
rect 2569 7663 2570 7671
rect 2582 7663 2583 7671
rect 2585 7667 2586 7671
rect 2585 7663 2590 7667
rect 2598 7663 2599 7671
rect 2601 7663 2604 7671
rect 2606 7663 2607 7671
rect 2619 7663 2620 7671
rect 2622 7663 2623 7671
rect 2635 7663 2636 7671
rect 2638 7663 2641 7671
rect 2643 7663 2644 7671
rect 2656 7663 2657 7671
rect 2659 7667 2660 7671
rect 2659 7663 2664 7667
rect 2672 7663 2673 7671
rect 2675 7663 2678 7671
rect 2680 7663 2681 7671
rect 2698 7663 2699 7671
rect 2701 7663 2702 7671
rect 2714 7663 2715 7671
rect 2717 7667 2718 7671
rect 2717 7663 2722 7667
rect 2730 7663 2731 7671
rect 2733 7663 2736 7671
rect 2738 7663 2739 7671
rect 2751 7663 2752 7671
rect 2754 7663 2755 7671
rect 3316 7663 3317 7671
rect 3319 7663 3322 7671
rect 3324 7663 3325 7671
rect 3337 7663 3338 7671
rect 3340 7667 3341 7671
rect 3340 7663 3345 7667
rect 3353 7663 3354 7671
rect 3356 7663 3359 7671
rect 3361 7663 3362 7671
rect 3379 7663 3380 7671
rect 3382 7663 3383 7671
rect 3395 7663 3396 7671
rect 3398 7667 3399 7671
rect 3398 7663 3403 7667
rect 3411 7663 3412 7671
rect 3414 7663 3417 7671
rect 3419 7663 3420 7671
rect 3432 7663 3433 7671
rect 3435 7663 3436 7671
rect 3448 7663 3449 7671
rect 3451 7663 3454 7671
rect 3456 7663 3457 7671
rect 3469 7663 3470 7671
rect 3472 7667 3473 7671
rect 3472 7663 3477 7667
rect 3485 7663 3486 7671
rect 3488 7663 3491 7671
rect 3493 7663 3494 7671
rect 3511 7663 3512 7671
rect 3514 7663 3515 7671
rect 3527 7663 3528 7671
rect 3530 7667 3531 7671
rect 3530 7663 3535 7667
rect 3543 7663 3544 7671
rect 3546 7663 3549 7671
rect 3551 7663 3552 7671
rect 3564 7663 3565 7671
rect 3567 7663 3568 7671
rect 3580 7663 3581 7671
rect 3583 7663 3586 7671
rect 3588 7663 3589 7671
rect 3601 7663 3602 7671
rect 3604 7667 3605 7671
rect 3604 7663 3609 7667
rect 3617 7663 3618 7671
rect 3620 7663 3623 7671
rect 3625 7663 3626 7671
rect 3643 7663 3644 7671
rect 3646 7663 3647 7671
rect 3659 7663 3660 7671
rect 3662 7667 3663 7671
rect 3662 7663 3667 7667
rect 3675 7663 3676 7671
rect 3678 7663 3681 7671
rect 3683 7663 3684 7671
rect 3696 7663 3697 7671
rect 3699 7663 3700 7671
rect 3154 7607 3155 7615
rect 3157 7607 3160 7615
rect 3162 7607 3163 7615
rect 3175 7607 3176 7615
rect 3178 7611 3179 7615
rect 3178 7607 3183 7611
rect 3191 7607 3192 7615
rect 3194 7607 3197 7615
rect 3199 7607 3200 7615
rect 3217 7607 3218 7615
rect 3220 7607 3221 7615
rect 3233 7607 3234 7615
rect 3236 7611 3237 7615
rect 3236 7607 3241 7611
rect 3249 7607 3250 7615
rect 3252 7607 3255 7615
rect 3257 7607 3258 7615
rect 3270 7607 3271 7615
rect 3273 7607 3274 7615
rect 4099 7607 4100 7615
rect 4102 7607 4105 7615
rect 4107 7607 4108 7615
rect 4120 7607 4121 7615
rect 4123 7611 4124 7615
rect 4123 7607 4128 7611
rect 4136 7607 4137 7615
rect 4139 7607 4142 7615
rect 4144 7607 4145 7615
rect 4162 7607 4163 7615
rect 4165 7607 4166 7615
rect 4178 7607 4179 7615
rect 4181 7611 4182 7615
rect 4181 7607 4186 7611
rect 4194 7607 4195 7615
rect 4197 7607 4200 7615
rect 4202 7607 4203 7615
rect 4215 7607 4216 7615
rect 4218 7607 4219 7615
rect 2371 7577 2372 7585
rect 2374 7577 2377 7585
rect 2379 7577 2380 7585
rect 2392 7577 2393 7585
rect 2395 7581 2396 7585
rect 2395 7577 2400 7581
rect 2408 7577 2409 7585
rect 2411 7577 2414 7585
rect 2416 7577 2417 7585
rect 2434 7577 2435 7585
rect 2437 7577 2438 7585
rect 2450 7577 2451 7585
rect 2453 7581 2454 7585
rect 2453 7577 2458 7581
rect 2466 7577 2467 7585
rect 2469 7577 2472 7585
rect 2474 7577 2475 7585
rect 2487 7577 2488 7585
rect 2490 7577 2491 7585
rect 2503 7577 2504 7585
rect 2506 7577 2509 7585
rect 2511 7577 2512 7585
rect 2524 7577 2525 7585
rect 2527 7581 2528 7585
rect 2527 7577 2532 7581
rect 2540 7577 2541 7585
rect 2543 7577 2546 7585
rect 2548 7577 2549 7585
rect 2566 7577 2567 7585
rect 2569 7577 2570 7585
rect 2582 7577 2583 7585
rect 2585 7581 2586 7585
rect 2585 7577 2590 7581
rect 2598 7577 2599 7585
rect 2601 7577 2604 7585
rect 2606 7577 2607 7585
rect 2619 7577 2620 7585
rect 2622 7577 2623 7585
rect 2635 7577 2636 7585
rect 2638 7577 2641 7585
rect 2643 7577 2644 7585
rect 2656 7577 2657 7585
rect 2659 7581 2660 7585
rect 2659 7577 2664 7581
rect 2672 7577 2673 7585
rect 2675 7577 2678 7585
rect 2680 7577 2681 7585
rect 2698 7577 2699 7585
rect 2701 7577 2702 7585
rect 2714 7577 2715 7585
rect 2717 7581 2718 7585
rect 2717 7577 2722 7581
rect 2730 7577 2731 7585
rect 2733 7577 2736 7585
rect 2738 7577 2739 7585
rect 2751 7577 2752 7585
rect 2754 7577 2755 7585
rect 3316 7577 3317 7585
rect 3319 7577 3322 7585
rect 3324 7577 3325 7585
rect 3337 7577 3338 7585
rect 3340 7581 3341 7585
rect 3340 7577 3345 7581
rect 3353 7577 3354 7585
rect 3356 7577 3359 7585
rect 3361 7577 3362 7585
rect 3379 7577 3380 7585
rect 3382 7577 3383 7585
rect 3395 7577 3396 7585
rect 3398 7581 3399 7585
rect 3398 7577 3403 7581
rect 3411 7577 3412 7585
rect 3414 7577 3417 7585
rect 3419 7577 3420 7585
rect 3432 7577 3433 7585
rect 3435 7577 3436 7585
rect 3448 7577 3449 7585
rect 3451 7577 3454 7585
rect 3456 7577 3457 7585
rect 3469 7577 3470 7585
rect 3472 7581 3473 7585
rect 3472 7577 3477 7581
rect 3485 7577 3486 7585
rect 3488 7577 3491 7585
rect 3493 7577 3494 7585
rect 3511 7577 3512 7585
rect 3514 7577 3515 7585
rect 3527 7577 3528 7585
rect 3530 7581 3531 7585
rect 3530 7577 3535 7581
rect 3543 7577 3544 7585
rect 3546 7577 3549 7585
rect 3551 7577 3552 7585
rect 3564 7577 3565 7585
rect 3567 7577 3568 7585
rect 3580 7577 3581 7585
rect 3583 7577 3586 7585
rect 3588 7577 3589 7585
rect 3601 7577 3602 7585
rect 3604 7581 3605 7585
rect 3604 7577 3609 7581
rect 3617 7577 3618 7585
rect 3620 7577 3623 7585
rect 3625 7577 3626 7585
rect 3643 7577 3644 7585
rect 3646 7577 3647 7585
rect 3659 7577 3660 7585
rect 3662 7581 3663 7585
rect 3662 7577 3667 7581
rect 3675 7577 3676 7585
rect 3678 7577 3681 7585
rect 3683 7577 3684 7585
rect 3696 7577 3697 7585
rect 3699 7577 3700 7585
rect 2371 7437 2372 7445
rect 2374 7437 2377 7445
rect 2379 7437 2380 7445
rect 2392 7437 2393 7445
rect 2395 7441 2396 7445
rect 2395 7437 2400 7441
rect 2408 7437 2409 7445
rect 2411 7437 2414 7445
rect 2416 7437 2417 7445
rect 2434 7437 2435 7445
rect 2437 7437 2438 7445
rect 2450 7437 2451 7445
rect 2453 7441 2454 7445
rect 2453 7437 2458 7441
rect 2466 7437 2467 7445
rect 2469 7437 2472 7445
rect 2474 7437 2475 7445
rect 2487 7437 2488 7445
rect 2490 7437 2491 7445
rect 2503 7437 2504 7445
rect 2506 7437 2509 7445
rect 2511 7437 2512 7445
rect 2524 7437 2525 7445
rect 2527 7441 2528 7445
rect 2527 7437 2532 7441
rect 2540 7437 2541 7445
rect 2543 7437 2546 7445
rect 2548 7437 2549 7445
rect 2566 7437 2567 7445
rect 2569 7437 2570 7445
rect 2582 7437 2583 7445
rect 2585 7441 2586 7445
rect 2585 7437 2590 7441
rect 2598 7437 2599 7445
rect 2601 7437 2604 7445
rect 2606 7437 2607 7445
rect 2619 7437 2620 7445
rect 2622 7437 2623 7445
rect 2635 7437 2636 7445
rect 2638 7437 2641 7445
rect 2643 7437 2644 7445
rect 2656 7437 2657 7445
rect 2659 7441 2660 7445
rect 2659 7437 2664 7441
rect 2672 7437 2673 7445
rect 2675 7437 2678 7445
rect 2680 7437 2681 7445
rect 2698 7437 2699 7445
rect 2701 7437 2702 7445
rect 2714 7437 2715 7445
rect 2717 7441 2718 7445
rect 2717 7437 2722 7441
rect 2730 7437 2731 7445
rect 2733 7437 2736 7445
rect 2738 7437 2739 7445
rect 2751 7437 2752 7445
rect 2754 7437 2755 7445
rect 3316 7437 3317 7445
rect 3319 7437 3322 7445
rect 3324 7437 3325 7445
rect 3337 7437 3338 7445
rect 3340 7441 3341 7445
rect 3340 7437 3345 7441
rect 3353 7437 3354 7445
rect 3356 7437 3359 7445
rect 3361 7437 3362 7445
rect 3379 7437 3380 7445
rect 3382 7437 3383 7445
rect 3395 7437 3396 7445
rect 3398 7441 3399 7445
rect 3398 7437 3403 7441
rect 3411 7437 3412 7445
rect 3414 7437 3417 7445
rect 3419 7437 3420 7445
rect 3432 7437 3433 7445
rect 3435 7437 3436 7445
rect 3448 7437 3449 7445
rect 3451 7437 3454 7445
rect 3456 7437 3457 7445
rect 3469 7437 3470 7445
rect 3472 7441 3473 7445
rect 3472 7437 3477 7441
rect 3485 7437 3486 7445
rect 3488 7437 3491 7445
rect 3493 7437 3494 7445
rect 3511 7437 3512 7445
rect 3514 7437 3515 7445
rect 3527 7437 3528 7445
rect 3530 7441 3531 7445
rect 3530 7437 3535 7441
rect 3543 7437 3544 7445
rect 3546 7437 3549 7445
rect 3551 7437 3552 7445
rect 3564 7437 3565 7445
rect 3567 7437 3568 7445
rect 3580 7437 3581 7445
rect 3583 7437 3586 7445
rect 3588 7437 3589 7445
rect 3601 7437 3602 7445
rect 3604 7441 3605 7445
rect 3604 7437 3609 7441
rect 3617 7437 3618 7445
rect 3620 7437 3623 7445
rect 3625 7437 3626 7445
rect 3643 7437 3644 7445
rect 3646 7437 3647 7445
rect 3659 7437 3660 7445
rect 3662 7441 3663 7445
rect 3662 7437 3667 7441
rect 3675 7437 3676 7445
rect 3678 7437 3681 7445
rect 3683 7437 3684 7445
rect 3696 7437 3697 7445
rect 3699 7437 3700 7445
rect 4578 7928 4579 7945
rect 4574 7924 4579 7928
rect 4578 7889 4579 7924
rect 4581 7889 4582 7945
rect 4586 7889 4587 7945
rect 4589 7928 4590 7945
rect 4594 7928 4595 7945
rect 4589 7924 4595 7928
rect 4589 7889 4590 7924
rect 4594 7889 4595 7924
rect 4597 7889 4598 7945
rect 4602 7889 4603 7945
rect 4605 7928 4606 7945
rect 4610 7928 4611 7945
rect 4605 7924 4611 7928
rect 4605 7889 4606 7924
rect 4610 7889 4611 7924
rect 4613 7889 4614 7945
rect 4618 7889 4619 7945
rect 4621 7928 4622 7945
rect 4626 7928 4627 7945
rect 4621 7924 4627 7928
rect 4621 7889 4622 7924
rect 4626 7889 4627 7924
rect 4631 7857 4634 7945
rect 4636 7857 4637 7945
rect 4641 7857 4642 7945
rect 4644 7936 4650 7945
rect 4644 7928 4645 7936
rect 4649 7928 4650 7936
rect 4644 7924 4650 7928
rect 4644 7857 4645 7924
rect 4649 7857 4650 7924
rect 4652 7857 4653 7945
rect 4657 7857 4658 7945
rect 4660 7928 4661 7945
rect 4665 7928 4666 7945
rect 4660 7924 4666 7928
rect 4660 7857 4661 7924
rect 4665 7857 4666 7924
rect 4674 7857 4677 7945
rect 4679 7857 4680 7945
rect 4684 7857 4685 7945
rect 4687 7936 4693 7945
rect 4687 7928 4688 7936
rect 4692 7928 4693 7936
rect 4687 7924 4693 7928
rect 4687 7857 4688 7924
rect 4692 7857 4693 7924
rect 4695 7857 4696 7945
rect 4700 7857 4701 7945
rect 4703 7928 4704 7945
rect 4708 7928 4709 7945
rect 4703 7924 4709 7928
rect 4703 7857 4704 7924
rect 4708 7857 4709 7924
rect 4713 7857 4718 7945
rect 4720 7857 4721 7945
rect 4725 7857 4726 7945
rect 4728 7936 4734 7945
rect 4728 7928 4729 7936
rect 4733 7928 4734 7936
rect 4728 7924 4734 7928
rect 4728 7857 4729 7924
rect 4733 7857 4734 7924
rect 4736 7857 4737 7945
rect 4741 7857 4742 7945
rect 4744 7928 4745 7945
rect 4749 7928 4750 7945
rect 4744 7924 4750 7928
rect 4744 7857 4745 7924
rect 4749 7857 4750 7924
<< ndcontact >>
rect 1402 9949 1406 9953
rect 1412 9949 1416 9953
rect 1422 9949 1426 9953
rect 1432 9949 1436 9953
rect 1397 9944 1401 9948
rect 1407 9944 1411 9948
rect 1417 9944 1421 9948
rect 1427 9944 1431 9948
rect 1437 9944 1441 9948
rect 1402 9939 1406 9943
rect 1412 9939 1416 9943
rect 1422 9939 1426 9943
rect 1432 9939 1436 9943
rect 1397 9934 1401 9938
rect 1407 9934 1411 9938
rect 1417 9934 1421 9938
rect 1427 9934 1431 9938
rect 1437 9934 1441 9938
rect 1402 9929 1406 9933
rect 1412 9929 1416 9933
rect 1422 9929 1426 9933
rect 1432 9929 1436 9933
rect 1397 9924 1401 9928
rect 1407 9924 1411 9928
rect 1417 9924 1421 9928
rect 1427 9924 1431 9928
rect 1437 9924 1441 9928
rect 1402 9919 1406 9923
rect 1412 9919 1416 9923
rect 1422 9919 1426 9923
rect 1432 9919 1436 9923
rect 1397 9914 1401 9918
rect 1407 9914 1411 9918
rect 1417 9914 1421 9918
rect 1427 9914 1431 9918
rect 1437 9914 1441 9918
rect 1402 9909 1406 9913
rect 1412 9909 1416 9913
rect 1422 9909 1426 9913
rect 1432 9909 1436 9913
rect 1397 9904 1401 9908
rect 1407 9904 1411 9908
rect 1417 9904 1421 9908
rect 1427 9904 1431 9908
rect 1437 9904 1441 9908
rect 1402 9899 1406 9903
rect 1412 9899 1416 9903
rect 1422 9899 1426 9903
rect 1432 9899 1436 9903
rect 1397 9894 1401 9898
rect 1407 9894 1411 9898
rect 1417 9894 1421 9898
rect 1427 9894 1431 9898
rect 1437 9894 1441 9898
rect 1402 9889 1406 9893
rect 1412 9889 1416 9893
rect 1422 9889 1426 9893
rect 1432 9889 1436 9893
rect 1397 9884 1401 9888
rect 1407 9884 1411 9888
rect 1417 9884 1421 9888
rect 1427 9884 1431 9888
rect 1437 9884 1441 9888
rect 1402 9879 1406 9883
rect 1412 9879 1416 9883
rect 1422 9879 1426 9883
rect 1432 9879 1436 9883
rect 1397 9874 1401 9878
rect 1407 9874 1411 9878
rect 1417 9874 1421 9878
rect 1427 9874 1431 9878
rect 1437 9874 1441 9878
rect 1402 9869 1406 9873
rect 1412 9869 1416 9873
rect 1422 9869 1426 9873
rect 1432 9869 1436 9873
rect 1397 9864 1401 9868
rect 1407 9864 1411 9868
rect 1417 9864 1421 9868
rect 1427 9864 1431 9868
rect 1437 9864 1441 9868
rect 1711 9949 1715 9953
rect 1721 9949 1725 9953
rect 1731 9949 1735 9953
rect 1741 9949 1745 9953
rect 1706 9944 1710 9948
rect 1716 9944 1720 9948
rect 1726 9944 1730 9948
rect 1736 9944 1740 9948
rect 1746 9944 1750 9948
rect 1711 9939 1715 9943
rect 1721 9939 1725 9943
rect 1731 9939 1735 9943
rect 1741 9939 1745 9943
rect 1706 9934 1710 9938
rect 1716 9934 1720 9938
rect 1726 9934 1730 9938
rect 1736 9934 1740 9938
rect 1746 9934 1750 9938
rect 1711 9929 1715 9933
rect 1721 9929 1725 9933
rect 1731 9929 1735 9933
rect 1741 9929 1745 9933
rect 1706 9924 1710 9928
rect 1716 9924 1720 9928
rect 1726 9924 1730 9928
rect 1736 9924 1740 9928
rect 1746 9924 1750 9928
rect 1711 9919 1715 9923
rect 1721 9919 1725 9923
rect 1731 9919 1735 9923
rect 1741 9919 1745 9923
rect 1706 9914 1710 9918
rect 1716 9914 1720 9918
rect 1726 9914 1730 9918
rect 1736 9914 1740 9918
rect 1746 9914 1750 9918
rect 1711 9909 1715 9913
rect 1721 9909 1725 9913
rect 1731 9909 1735 9913
rect 1741 9909 1745 9913
rect 1706 9904 1710 9908
rect 1716 9904 1720 9908
rect 1726 9904 1730 9908
rect 1736 9904 1740 9908
rect 1746 9904 1750 9908
rect 1711 9899 1715 9903
rect 1721 9899 1725 9903
rect 1731 9899 1735 9903
rect 1741 9899 1745 9903
rect 1706 9894 1710 9898
rect 1716 9894 1720 9898
rect 1726 9894 1730 9898
rect 1736 9894 1740 9898
rect 1746 9894 1750 9898
rect 1711 9889 1715 9893
rect 1721 9889 1725 9893
rect 1731 9889 1735 9893
rect 1741 9889 1745 9893
rect 1706 9884 1710 9888
rect 1716 9884 1720 9888
rect 1726 9884 1730 9888
rect 1736 9884 1740 9888
rect 1746 9884 1750 9888
rect 1711 9879 1715 9883
rect 1721 9879 1725 9883
rect 1731 9879 1735 9883
rect 1741 9879 1745 9883
rect 1706 9874 1710 9878
rect 1716 9874 1720 9878
rect 1726 9874 1730 9878
rect 1736 9874 1740 9878
rect 1746 9874 1750 9878
rect 1711 9869 1715 9873
rect 1721 9869 1725 9873
rect 1731 9869 1735 9873
rect 1741 9869 1745 9873
rect 1706 9864 1710 9868
rect 1716 9864 1720 9868
rect 1726 9864 1730 9868
rect 1736 9864 1740 9868
rect 1746 9864 1750 9868
rect 2020 9949 2024 9953
rect 2030 9949 2034 9953
rect 2040 9949 2044 9953
rect 2050 9949 2054 9953
rect 2015 9944 2019 9948
rect 2025 9944 2029 9948
rect 2035 9944 2039 9948
rect 2045 9944 2049 9948
rect 2055 9944 2059 9948
rect 2020 9939 2024 9943
rect 2030 9939 2034 9943
rect 2040 9939 2044 9943
rect 2050 9939 2054 9943
rect 2015 9934 2019 9938
rect 2025 9934 2029 9938
rect 2035 9934 2039 9938
rect 2045 9934 2049 9938
rect 2055 9934 2059 9938
rect 2020 9929 2024 9933
rect 2030 9929 2034 9933
rect 2040 9929 2044 9933
rect 2050 9929 2054 9933
rect 2015 9924 2019 9928
rect 2025 9924 2029 9928
rect 2035 9924 2039 9928
rect 2045 9924 2049 9928
rect 2055 9924 2059 9928
rect 2020 9919 2024 9923
rect 2030 9919 2034 9923
rect 2040 9919 2044 9923
rect 2050 9919 2054 9923
rect 2015 9914 2019 9918
rect 2025 9914 2029 9918
rect 2035 9914 2039 9918
rect 2045 9914 2049 9918
rect 2055 9914 2059 9918
rect 2020 9909 2024 9913
rect 2030 9909 2034 9913
rect 2040 9909 2044 9913
rect 2050 9909 2054 9913
rect 2015 9904 2019 9908
rect 2025 9904 2029 9908
rect 2035 9904 2039 9908
rect 2045 9904 2049 9908
rect 2055 9904 2059 9908
rect 2020 9899 2024 9903
rect 2030 9899 2034 9903
rect 2040 9899 2044 9903
rect 2050 9899 2054 9903
rect 2015 9894 2019 9898
rect 2025 9894 2029 9898
rect 2035 9894 2039 9898
rect 2045 9894 2049 9898
rect 2055 9894 2059 9898
rect 2020 9889 2024 9893
rect 2030 9889 2034 9893
rect 2040 9889 2044 9893
rect 2050 9889 2054 9893
rect 2015 9884 2019 9888
rect 2025 9884 2029 9888
rect 2035 9884 2039 9888
rect 2045 9884 2049 9888
rect 2055 9884 2059 9888
rect 2020 9879 2024 9883
rect 2030 9879 2034 9883
rect 2040 9879 2044 9883
rect 2050 9879 2054 9883
rect 2015 9874 2019 9878
rect 2025 9874 2029 9878
rect 2035 9874 2039 9878
rect 2045 9874 2049 9878
rect 2055 9874 2059 9878
rect 2020 9869 2024 9873
rect 2030 9869 2034 9873
rect 2040 9869 2044 9873
rect 2050 9869 2054 9873
rect 2015 9864 2019 9868
rect 2025 9864 2029 9868
rect 2035 9864 2039 9868
rect 2045 9864 2049 9868
rect 2055 9864 2059 9868
rect 2329 9949 2333 9953
rect 2339 9949 2343 9953
rect 2349 9949 2353 9953
rect 2359 9949 2363 9953
rect 2324 9944 2328 9948
rect 2334 9944 2338 9948
rect 2344 9944 2348 9948
rect 2354 9944 2358 9948
rect 2364 9944 2368 9948
rect 2329 9939 2333 9943
rect 2339 9939 2343 9943
rect 2349 9939 2353 9943
rect 2359 9939 2363 9943
rect 2324 9934 2328 9938
rect 2334 9934 2338 9938
rect 2344 9934 2348 9938
rect 2354 9934 2358 9938
rect 2364 9934 2368 9938
rect 2329 9929 2333 9933
rect 2339 9929 2343 9933
rect 2349 9929 2353 9933
rect 2359 9929 2363 9933
rect 2324 9924 2328 9928
rect 2334 9924 2338 9928
rect 2344 9924 2348 9928
rect 2354 9924 2358 9928
rect 2364 9924 2368 9928
rect 2329 9919 2333 9923
rect 2339 9919 2343 9923
rect 2349 9919 2353 9923
rect 2359 9919 2363 9923
rect 2324 9914 2328 9918
rect 2334 9914 2338 9918
rect 2344 9914 2348 9918
rect 2354 9914 2358 9918
rect 2364 9914 2368 9918
rect 2329 9909 2333 9913
rect 2339 9909 2343 9913
rect 2349 9909 2353 9913
rect 2359 9909 2363 9913
rect 2324 9904 2328 9908
rect 2334 9904 2338 9908
rect 2344 9904 2348 9908
rect 2354 9904 2358 9908
rect 2364 9904 2368 9908
rect 2329 9899 2333 9903
rect 2339 9899 2343 9903
rect 2349 9899 2353 9903
rect 2359 9899 2363 9903
rect 2324 9894 2328 9898
rect 2334 9894 2338 9898
rect 2344 9894 2348 9898
rect 2354 9894 2358 9898
rect 2364 9894 2368 9898
rect 2329 9889 2333 9893
rect 2339 9889 2343 9893
rect 2349 9889 2353 9893
rect 2359 9889 2363 9893
rect 2324 9884 2328 9888
rect 2334 9884 2338 9888
rect 2344 9884 2348 9888
rect 2354 9884 2358 9888
rect 2364 9884 2368 9888
rect 2329 9879 2333 9883
rect 2339 9879 2343 9883
rect 2349 9879 2353 9883
rect 2359 9879 2363 9883
rect 2324 9874 2328 9878
rect 2334 9874 2338 9878
rect 2344 9874 2348 9878
rect 2354 9874 2358 9878
rect 2364 9874 2368 9878
rect 2329 9869 2333 9873
rect 2339 9869 2343 9873
rect 2349 9869 2353 9873
rect 2359 9869 2363 9873
rect 2324 9864 2328 9868
rect 2334 9864 2338 9868
rect 2344 9864 2348 9868
rect 2354 9864 2358 9868
rect 2364 9864 2368 9868
rect 2638 9949 2642 9953
rect 2648 9949 2652 9953
rect 2658 9949 2662 9953
rect 2668 9949 2672 9953
rect 2633 9944 2637 9948
rect 2643 9944 2647 9948
rect 2653 9944 2657 9948
rect 2663 9944 2667 9948
rect 2673 9944 2677 9948
rect 2638 9939 2642 9943
rect 2648 9939 2652 9943
rect 2658 9939 2662 9943
rect 2668 9939 2672 9943
rect 2633 9934 2637 9938
rect 2643 9934 2647 9938
rect 2653 9934 2657 9938
rect 2663 9934 2667 9938
rect 2673 9934 2677 9938
rect 2638 9929 2642 9933
rect 2648 9929 2652 9933
rect 2658 9929 2662 9933
rect 2668 9929 2672 9933
rect 2633 9924 2637 9928
rect 2643 9924 2647 9928
rect 2653 9924 2657 9928
rect 2663 9924 2667 9928
rect 2673 9924 2677 9928
rect 2638 9919 2642 9923
rect 2648 9919 2652 9923
rect 2658 9919 2662 9923
rect 2668 9919 2672 9923
rect 2633 9914 2637 9918
rect 2643 9914 2647 9918
rect 2653 9914 2657 9918
rect 2663 9914 2667 9918
rect 2673 9914 2677 9918
rect 2638 9909 2642 9913
rect 2648 9909 2652 9913
rect 2658 9909 2662 9913
rect 2668 9909 2672 9913
rect 2633 9904 2637 9908
rect 2643 9904 2647 9908
rect 2653 9904 2657 9908
rect 2663 9904 2667 9908
rect 2673 9904 2677 9908
rect 2638 9899 2642 9903
rect 2648 9899 2652 9903
rect 2658 9899 2662 9903
rect 2668 9899 2672 9903
rect 2633 9894 2637 9898
rect 2643 9894 2647 9898
rect 2653 9894 2657 9898
rect 2663 9894 2667 9898
rect 2673 9894 2677 9898
rect 2638 9889 2642 9893
rect 2648 9889 2652 9893
rect 2658 9889 2662 9893
rect 2668 9889 2672 9893
rect 2633 9884 2637 9888
rect 2643 9884 2647 9888
rect 2653 9884 2657 9888
rect 2663 9884 2667 9888
rect 2673 9884 2677 9888
rect 2638 9879 2642 9883
rect 2648 9879 2652 9883
rect 2658 9879 2662 9883
rect 2668 9879 2672 9883
rect 2633 9874 2637 9878
rect 2643 9874 2647 9878
rect 2653 9874 2657 9878
rect 2663 9874 2667 9878
rect 2673 9874 2677 9878
rect 2638 9869 2642 9873
rect 2648 9869 2652 9873
rect 2658 9869 2662 9873
rect 2668 9869 2672 9873
rect 2633 9864 2637 9868
rect 2643 9864 2647 9868
rect 2653 9864 2657 9868
rect 2663 9864 2667 9868
rect 2673 9864 2677 9868
rect 2947 9949 2951 9953
rect 2957 9949 2961 9953
rect 2967 9949 2971 9953
rect 2977 9949 2981 9953
rect 2942 9944 2946 9948
rect 2952 9944 2956 9948
rect 2962 9944 2966 9948
rect 2972 9944 2976 9948
rect 2982 9944 2986 9948
rect 2947 9939 2951 9943
rect 2957 9939 2961 9943
rect 2967 9939 2971 9943
rect 2977 9939 2981 9943
rect 2942 9934 2946 9938
rect 2952 9934 2956 9938
rect 2962 9934 2966 9938
rect 2972 9934 2976 9938
rect 2982 9934 2986 9938
rect 2947 9929 2951 9933
rect 2957 9929 2961 9933
rect 2967 9929 2971 9933
rect 2977 9929 2981 9933
rect 2942 9924 2946 9928
rect 2952 9924 2956 9928
rect 2962 9924 2966 9928
rect 2972 9924 2976 9928
rect 2982 9924 2986 9928
rect 2947 9919 2951 9923
rect 2957 9919 2961 9923
rect 2967 9919 2971 9923
rect 2977 9919 2981 9923
rect 2942 9914 2946 9918
rect 2952 9914 2956 9918
rect 2962 9914 2966 9918
rect 2972 9914 2976 9918
rect 2982 9914 2986 9918
rect 2947 9909 2951 9913
rect 2957 9909 2961 9913
rect 2967 9909 2971 9913
rect 2977 9909 2981 9913
rect 2942 9904 2946 9908
rect 2952 9904 2956 9908
rect 2962 9904 2966 9908
rect 2972 9904 2976 9908
rect 2982 9904 2986 9908
rect 2947 9899 2951 9903
rect 2957 9899 2961 9903
rect 2967 9899 2971 9903
rect 2977 9899 2981 9903
rect 2942 9894 2946 9898
rect 2952 9894 2956 9898
rect 2962 9894 2966 9898
rect 2972 9894 2976 9898
rect 2982 9894 2986 9898
rect 2947 9889 2951 9893
rect 2957 9889 2961 9893
rect 2967 9889 2971 9893
rect 2977 9889 2981 9893
rect 2942 9884 2946 9888
rect 2952 9884 2956 9888
rect 2962 9884 2966 9888
rect 2972 9884 2976 9888
rect 2982 9884 2986 9888
rect 2947 9879 2951 9883
rect 2957 9879 2961 9883
rect 2967 9879 2971 9883
rect 2977 9879 2981 9883
rect 2942 9874 2946 9878
rect 2952 9874 2956 9878
rect 2962 9874 2966 9878
rect 2972 9874 2976 9878
rect 2982 9874 2986 9878
rect 2947 9869 2951 9873
rect 2957 9869 2961 9873
rect 2967 9869 2971 9873
rect 2977 9869 2981 9873
rect 2942 9864 2946 9868
rect 2952 9864 2956 9868
rect 2962 9864 2966 9868
rect 2972 9864 2976 9868
rect 2982 9864 2986 9868
rect 3256 9949 3260 9953
rect 3266 9949 3270 9953
rect 3276 9949 3280 9953
rect 3286 9949 3290 9953
rect 3251 9944 3255 9948
rect 3261 9944 3265 9948
rect 3271 9944 3275 9948
rect 3281 9944 3285 9948
rect 3291 9944 3295 9948
rect 3256 9939 3260 9943
rect 3266 9939 3270 9943
rect 3276 9939 3280 9943
rect 3286 9939 3290 9943
rect 3251 9934 3255 9938
rect 3261 9934 3265 9938
rect 3271 9934 3275 9938
rect 3281 9934 3285 9938
rect 3291 9934 3295 9938
rect 3256 9929 3260 9933
rect 3266 9929 3270 9933
rect 3276 9929 3280 9933
rect 3286 9929 3290 9933
rect 3251 9924 3255 9928
rect 3261 9924 3265 9928
rect 3271 9924 3275 9928
rect 3281 9924 3285 9928
rect 3291 9924 3295 9928
rect 3256 9919 3260 9923
rect 3266 9919 3270 9923
rect 3276 9919 3280 9923
rect 3286 9919 3290 9923
rect 3251 9914 3255 9918
rect 3261 9914 3265 9918
rect 3271 9914 3275 9918
rect 3281 9914 3285 9918
rect 3291 9914 3295 9918
rect 3256 9909 3260 9913
rect 3266 9909 3270 9913
rect 3276 9909 3280 9913
rect 3286 9909 3290 9913
rect 3251 9904 3255 9908
rect 3261 9904 3265 9908
rect 3271 9904 3275 9908
rect 3281 9904 3285 9908
rect 3291 9904 3295 9908
rect 3256 9899 3260 9903
rect 3266 9899 3270 9903
rect 3276 9899 3280 9903
rect 3286 9899 3290 9903
rect 3251 9894 3255 9898
rect 3261 9894 3265 9898
rect 3271 9894 3275 9898
rect 3281 9894 3285 9898
rect 3291 9894 3295 9898
rect 3256 9889 3260 9893
rect 3266 9889 3270 9893
rect 3276 9889 3280 9893
rect 3286 9889 3290 9893
rect 3251 9884 3255 9888
rect 3261 9884 3265 9888
rect 3271 9884 3275 9888
rect 3281 9884 3285 9888
rect 3291 9884 3295 9888
rect 3256 9879 3260 9883
rect 3266 9879 3270 9883
rect 3276 9879 3280 9883
rect 3286 9879 3290 9883
rect 3251 9874 3255 9878
rect 3261 9874 3265 9878
rect 3271 9874 3275 9878
rect 3281 9874 3285 9878
rect 3291 9874 3295 9878
rect 3256 9869 3260 9873
rect 3266 9869 3270 9873
rect 3276 9869 3280 9873
rect 3286 9869 3290 9873
rect 3251 9864 3255 9868
rect 3261 9864 3265 9868
rect 3271 9864 3275 9868
rect 3281 9864 3285 9868
rect 3291 9864 3295 9868
rect 3565 9949 3569 9953
rect 3575 9949 3579 9953
rect 3585 9949 3589 9953
rect 3595 9949 3599 9953
rect 3560 9944 3564 9948
rect 3570 9944 3574 9948
rect 3580 9944 3584 9948
rect 3590 9944 3594 9948
rect 3600 9944 3604 9948
rect 3565 9939 3569 9943
rect 3575 9939 3579 9943
rect 3585 9939 3589 9943
rect 3595 9939 3599 9943
rect 3560 9934 3564 9938
rect 3570 9934 3574 9938
rect 3580 9934 3584 9938
rect 3590 9934 3594 9938
rect 3600 9934 3604 9938
rect 3565 9929 3569 9933
rect 3575 9929 3579 9933
rect 3585 9929 3589 9933
rect 3595 9929 3599 9933
rect 3560 9924 3564 9928
rect 3570 9924 3574 9928
rect 3580 9924 3584 9928
rect 3590 9924 3594 9928
rect 3600 9924 3604 9928
rect 3565 9919 3569 9923
rect 3575 9919 3579 9923
rect 3585 9919 3589 9923
rect 3595 9919 3599 9923
rect 3560 9914 3564 9918
rect 3570 9914 3574 9918
rect 3580 9914 3584 9918
rect 3590 9914 3594 9918
rect 3600 9914 3604 9918
rect 3565 9909 3569 9913
rect 3575 9909 3579 9913
rect 3585 9909 3589 9913
rect 3595 9909 3599 9913
rect 3560 9904 3564 9908
rect 3570 9904 3574 9908
rect 3580 9904 3584 9908
rect 3590 9904 3594 9908
rect 3600 9904 3604 9908
rect 3565 9899 3569 9903
rect 3575 9899 3579 9903
rect 3585 9899 3589 9903
rect 3595 9899 3599 9903
rect 3560 9894 3564 9898
rect 3570 9894 3574 9898
rect 3580 9894 3584 9898
rect 3590 9894 3594 9898
rect 3600 9894 3604 9898
rect 3565 9889 3569 9893
rect 3575 9889 3579 9893
rect 3585 9889 3589 9893
rect 3595 9889 3599 9893
rect 3560 9884 3564 9888
rect 3570 9884 3574 9888
rect 3580 9884 3584 9888
rect 3590 9884 3594 9888
rect 3600 9884 3604 9888
rect 3565 9879 3569 9883
rect 3575 9879 3579 9883
rect 3585 9879 3589 9883
rect 3595 9879 3599 9883
rect 3560 9874 3564 9878
rect 3570 9874 3574 9878
rect 3580 9874 3584 9878
rect 3590 9874 3594 9878
rect 3600 9874 3604 9878
rect 3565 9869 3569 9873
rect 3575 9869 3579 9873
rect 3585 9869 3589 9873
rect 3595 9869 3599 9873
rect 3560 9864 3564 9868
rect 3570 9864 3574 9868
rect 3580 9864 3584 9868
rect 3590 9864 3594 9868
rect 3600 9864 3604 9868
rect 3874 9949 3878 9953
rect 3884 9949 3888 9953
rect 3894 9949 3898 9953
rect 3904 9949 3908 9953
rect 3869 9944 3873 9948
rect 3879 9944 3883 9948
rect 3889 9944 3893 9948
rect 3899 9944 3903 9948
rect 3909 9944 3913 9948
rect 3874 9939 3878 9943
rect 3884 9939 3888 9943
rect 3894 9939 3898 9943
rect 3904 9939 3908 9943
rect 3869 9934 3873 9938
rect 3879 9934 3883 9938
rect 3889 9934 3893 9938
rect 3899 9934 3903 9938
rect 3909 9934 3913 9938
rect 3874 9929 3878 9933
rect 3884 9929 3888 9933
rect 3894 9929 3898 9933
rect 3904 9929 3908 9933
rect 3869 9924 3873 9928
rect 3879 9924 3883 9928
rect 3889 9924 3893 9928
rect 3899 9924 3903 9928
rect 3909 9924 3913 9928
rect 3874 9919 3878 9923
rect 3884 9919 3888 9923
rect 3894 9919 3898 9923
rect 3904 9919 3908 9923
rect 3869 9914 3873 9918
rect 3879 9914 3883 9918
rect 3889 9914 3893 9918
rect 3899 9914 3903 9918
rect 3909 9914 3913 9918
rect 3874 9909 3878 9913
rect 3884 9909 3888 9913
rect 3894 9909 3898 9913
rect 3904 9909 3908 9913
rect 3869 9904 3873 9908
rect 3879 9904 3883 9908
rect 3889 9904 3893 9908
rect 3899 9904 3903 9908
rect 3909 9904 3913 9908
rect 3874 9899 3878 9903
rect 3884 9899 3888 9903
rect 3894 9899 3898 9903
rect 3904 9899 3908 9903
rect 3869 9894 3873 9898
rect 3879 9894 3883 9898
rect 3889 9894 3893 9898
rect 3899 9894 3903 9898
rect 3909 9894 3913 9898
rect 3874 9889 3878 9893
rect 3884 9889 3888 9893
rect 3894 9889 3898 9893
rect 3904 9889 3908 9893
rect 3869 9884 3873 9888
rect 3879 9884 3883 9888
rect 3889 9884 3893 9888
rect 3899 9884 3903 9888
rect 3909 9884 3913 9888
rect 3874 9879 3878 9883
rect 3884 9879 3888 9883
rect 3894 9879 3898 9883
rect 3904 9879 3908 9883
rect 3869 9874 3873 9878
rect 3879 9874 3883 9878
rect 3889 9874 3893 9878
rect 3899 9874 3903 9878
rect 3909 9874 3913 9878
rect 3874 9869 3878 9873
rect 3884 9869 3888 9873
rect 3894 9869 3898 9873
rect 3904 9869 3908 9873
rect 3869 9864 3873 9868
rect 3879 9864 3883 9868
rect 3889 9864 3893 9868
rect 3899 9864 3903 9868
rect 3909 9864 3913 9868
rect 1829 9827 1836 9831
rect 1840 9827 1869 9831
rect 2138 9827 2145 9831
rect 2149 9827 2178 9831
rect 2447 9827 2454 9831
rect 2458 9827 2487 9831
rect 2756 9827 2763 9831
rect 2767 9827 2796 9831
rect 3065 9827 3072 9831
rect 3076 9827 3105 9831
rect 3992 9827 3999 9831
rect 4003 9827 4032 9831
rect 1829 9819 1869 9823
rect 2138 9819 2178 9823
rect 2447 9819 2487 9823
rect 2756 9819 2796 9823
rect 3065 9819 3105 9823
rect 3992 9819 4032 9823
rect 1829 9811 1836 9815
rect 1840 9811 1869 9815
rect 1829 9803 1869 9807
rect 1829 9795 1836 9799
rect 1840 9795 1869 9799
rect 1829 9787 1869 9791
rect 2138 9811 2145 9815
rect 2149 9811 2178 9815
rect 2138 9803 2178 9807
rect 2138 9795 2145 9799
rect 2149 9795 2178 9799
rect 2138 9787 2178 9791
rect 2447 9811 2454 9815
rect 2458 9811 2487 9815
rect 2447 9803 2487 9807
rect 2447 9795 2454 9799
rect 2458 9795 2487 9799
rect 2447 9787 2487 9791
rect 2756 9811 2763 9815
rect 2767 9811 2796 9815
rect 2756 9803 2796 9807
rect 2756 9795 2763 9799
rect 2767 9795 2796 9799
rect 2756 9787 2796 9791
rect 3065 9811 3072 9815
rect 3076 9811 3105 9815
rect 3065 9803 3105 9807
rect 3065 9795 3072 9799
rect 3076 9795 3105 9799
rect 3065 9787 3105 9791
rect 3992 9811 3999 9815
rect 4003 9811 4032 9815
rect 3992 9803 4032 9807
rect 3992 9795 3999 9799
rect 4003 9795 4032 9799
rect 3992 9787 4032 9791
rect 1829 9779 1836 9783
rect 1840 9779 1869 9783
rect 2138 9779 2145 9783
rect 2149 9779 2178 9783
rect 2447 9779 2454 9783
rect 2458 9779 2487 9783
rect 2756 9779 2763 9783
rect 2767 9779 2796 9783
rect 3065 9779 3072 9783
rect 3076 9779 3105 9783
rect 3992 9779 3999 9783
rect 4003 9779 4032 9783
rect 2851 9299 2855 9303
rect 2864 9299 2868 9303
rect 2872 9299 2876 9303
rect 2880 9299 2884 9303
rect 2888 9299 2892 9303
rect 2901 9299 2905 9303
rect 2914 9299 2918 9303
rect 2922 9299 2926 9303
rect 2930 9299 2934 9303
rect 2938 9299 2942 9303
rect 2946 9299 2950 9303
rect 2959 9299 2963 9303
rect 2967 9299 2971 9303
rect 2975 9299 2979 9303
rect 2983 9299 2987 9303
rect 2996 9299 3000 9303
rect 3004 9299 3008 9303
rect 3012 9299 3016 9303
rect 3020 9299 3024 9303
rect 3033 9299 3037 9303
rect 3046 9299 3050 9303
rect 3054 9299 3058 9303
rect 3062 9299 3066 9303
rect 3070 9299 3074 9303
rect 3078 9299 3082 9303
rect 3091 9299 3095 9303
rect 3099 9299 3103 9303
rect 3107 9299 3111 9303
rect 3115 9299 3119 9303
rect 3128 9299 3132 9303
rect 3136 9299 3140 9303
rect 3144 9299 3148 9303
rect 3152 9299 3156 9303
rect 3165 9299 3169 9303
rect 3178 9299 3182 9303
rect 3186 9299 3190 9303
rect 3194 9299 3198 9303
rect 3202 9299 3206 9303
rect 3210 9299 3214 9303
rect 3223 9299 3227 9303
rect 3231 9299 3235 9303
rect 3239 9299 3243 9303
rect 3247 9299 3251 9303
rect 3260 9299 3264 9303
rect 3268 9299 3272 9303
rect 3276 9299 3280 9303
rect 3284 9299 3288 9303
rect 3297 9299 3301 9303
rect 3310 9299 3314 9303
rect 3318 9299 3322 9303
rect 3326 9299 3330 9303
rect 3334 9299 3338 9303
rect 3342 9299 3346 9303
rect 3355 9299 3359 9303
rect 3363 9299 3367 9303
rect 3371 9299 3375 9303
rect 3796 9299 3800 9303
rect 3809 9299 3813 9303
rect 3817 9299 3821 9303
rect 3825 9299 3829 9303
rect 3833 9299 3837 9303
rect 3846 9299 3850 9303
rect 3859 9299 3863 9303
rect 3867 9299 3871 9303
rect 3875 9299 3879 9303
rect 3883 9299 3887 9303
rect 3891 9299 3895 9303
rect 3904 9299 3908 9303
rect 3912 9299 3916 9303
rect 3920 9299 3924 9303
rect 3928 9299 3932 9303
rect 3941 9299 3945 9303
rect 3949 9299 3953 9303
rect 3957 9299 3961 9303
rect 3965 9299 3969 9303
rect 3978 9299 3982 9303
rect 3991 9299 3995 9303
rect 3999 9299 4003 9303
rect 4007 9299 4011 9303
rect 4015 9299 4019 9303
rect 4023 9299 4027 9303
rect 4036 9299 4040 9303
rect 4044 9299 4048 9303
rect 4052 9299 4056 9303
rect 4060 9299 4064 9303
rect 4073 9299 4077 9303
rect 4081 9299 4085 9303
rect 4089 9299 4093 9303
rect 4097 9299 4101 9303
rect 4110 9299 4114 9303
rect 4123 9299 4127 9303
rect 4131 9299 4135 9303
rect 4139 9299 4143 9303
rect 4147 9299 4151 9303
rect 4155 9299 4159 9303
rect 4168 9299 4172 9303
rect 4176 9299 4180 9303
rect 4184 9299 4188 9303
rect 4192 9299 4196 9303
rect 4205 9299 4209 9303
rect 4213 9299 4217 9303
rect 4221 9299 4225 9303
rect 4229 9299 4233 9303
rect 4242 9299 4246 9303
rect 4255 9299 4259 9303
rect 4263 9299 4267 9303
rect 4271 9299 4275 9303
rect 4279 9299 4283 9303
rect 4287 9299 4291 9303
rect 4300 9299 4304 9303
rect 4308 9299 4312 9303
rect 4316 9299 4320 9303
rect 2499 9266 2503 9270
rect 2512 9266 2516 9270
rect 2520 9266 2524 9270
rect 2528 9266 2532 9270
rect 2536 9266 2540 9270
rect 2549 9266 2553 9270
rect 2562 9266 2566 9270
rect 2570 9266 2574 9270
rect 2578 9266 2582 9270
rect 2586 9266 2590 9270
rect 2594 9266 2598 9270
rect 2607 9266 2611 9270
rect 2615 9266 2619 9270
rect 2623 9266 2627 9270
rect 3444 9266 3448 9270
rect 3457 9266 3461 9270
rect 3465 9266 3469 9270
rect 3473 9266 3477 9270
rect 3481 9266 3485 9270
rect 3494 9266 3498 9270
rect 3507 9266 3511 9270
rect 3515 9266 3519 9270
rect 3523 9266 3527 9270
rect 3531 9266 3535 9270
rect 3539 9266 3543 9270
rect 3552 9266 3556 9270
rect 3560 9266 3564 9270
rect 3568 9266 3572 9270
rect 2623 9229 2627 9233
rect 2631 9229 2635 9233
rect 3030 9233 3034 9237
rect 3038 9233 3042 9237
rect 3054 9229 3058 9233
rect 3069 9229 3073 9233
rect 3111 9233 3115 9237
rect 3119 9233 3123 9237
rect 3135 9229 3139 9233
rect 3150 9229 3154 9233
rect 3084 9225 3088 9229
rect 3092 9225 3096 9229
rect 2506 9220 2510 9224
rect 2514 9220 2518 9224
rect 2856 9220 2860 9224
rect 2864 9220 2868 9224
rect 2872 9220 2876 9224
rect 2880 9220 2884 9224
rect 2888 9220 2892 9224
rect 2896 9220 2900 9224
rect 2907 9220 2911 9224
rect 2924 9220 2928 9224
rect 2941 9220 2945 9224
rect 2950 9220 2954 9224
rect 2963 9220 2967 9224
rect 2971 9220 2975 9224
rect 2979 9220 2983 9224
rect 2996 9220 3000 9224
rect 3006 9220 3010 9224
rect 3014 9220 3018 9224
rect 3165 9225 3169 9229
rect 3173 9225 3177 9229
rect 3568 9229 3572 9233
rect 3576 9229 3580 9233
rect 3975 9233 3979 9237
rect 3983 9233 3987 9237
rect 3999 9229 4003 9233
rect 4014 9229 4018 9233
rect 4056 9233 4060 9237
rect 4064 9233 4068 9237
rect 4080 9229 4084 9233
rect 4095 9229 4099 9233
rect 4029 9225 4033 9229
rect 4037 9225 4041 9229
rect 3451 9220 3455 9224
rect 3459 9220 3463 9224
rect 3801 9220 3805 9224
rect 3809 9220 3813 9224
rect 3817 9220 3821 9224
rect 3825 9220 3829 9224
rect 3833 9220 3837 9224
rect 3841 9220 3845 9224
rect 3852 9220 3856 9224
rect 3869 9220 3873 9224
rect 3886 9220 3890 9224
rect 3895 9220 3899 9224
rect 3908 9220 3912 9224
rect 3916 9220 3920 9224
rect 3924 9220 3928 9224
rect 3941 9220 3945 9224
rect 3951 9220 3955 9224
rect 3959 9220 3963 9224
rect 4110 9225 4114 9229
rect 4118 9225 4122 9229
rect 2856 9174 2860 9178
rect 2864 9174 2868 9178
rect 2872 9174 2876 9178
rect 2880 9174 2884 9178
rect 2888 9174 2892 9178
rect 2896 9174 2900 9178
rect 2907 9174 2911 9178
rect 2924 9174 2928 9178
rect 2941 9174 2945 9178
rect 2950 9174 2954 9178
rect 2963 9174 2967 9178
rect 2971 9174 2975 9178
rect 2979 9174 2983 9178
rect 2996 9174 3000 9178
rect 3006 9174 3010 9178
rect 3014 9174 3018 9178
rect 2490 9164 2494 9168
rect 2498 9164 2502 9168
rect 2506 9164 2510 9168
rect 2519 9164 2523 9168
rect 2527 9164 2531 9168
rect 2535 9164 2539 9168
rect 2543 9164 2547 9168
rect 2551 9164 2555 9168
rect 2564 9164 2568 9168
rect 2577 9164 2581 9168
rect 2585 9164 2589 9168
rect 2593 9164 2597 9168
rect 2601 9164 2605 9168
rect 2614 9164 2618 9168
rect 3054 9173 3058 9177
rect 3069 9173 3073 9177
rect 3135 9173 3139 9177
rect 3150 9173 3154 9177
rect 3801 9174 3805 9178
rect 3809 9174 3813 9178
rect 3817 9174 3821 9178
rect 3825 9174 3829 9178
rect 3833 9174 3837 9178
rect 3841 9174 3845 9178
rect 3852 9174 3856 9178
rect 3869 9174 3873 9178
rect 3886 9174 3890 9178
rect 3895 9174 3899 9178
rect 3908 9174 3912 9178
rect 3916 9174 3920 9178
rect 3924 9174 3928 9178
rect 3941 9174 3945 9178
rect 3951 9174 3955 9178
rect 3959 9174 3963 9178
rect 3435 9164 3439 9168
rect 3443 9164 3447 9168
rect 3451 9164 3455 9168
rect 3464 9164 3468 9168
rect 3472 9164 3476 9168
rect 3480 9164 3484 9168
rect 3488 9164 3492 9168
rect 3496 9164 3500 9168
rect 3509 9164 3513 9168
rect 3522 9164 3526 9168
rect 3530 9164 3534 9168
rect 3538 9164 3542 9168
rect 3546 9164 3550 9168
rect 3559 9164 3563 9168
rect 3999 9173 4003 9177
rect 4014 9173 4018 9177
rect 4080 9173 4084 9177
rect 4095 9173 4099 9177
rect 3054 9097 3058 9101
rect 3069 9097 3073 9101
rect 3135 9101 3139 9105
rect 3143 9101 3147 9105
rect 3159 9097 3163 9101
rect 3174 9097 3178 9101
rect 3084 9093 3088 9097
rect 3092 9093 3096 9097
rect 2856 9088 2860 9092
rect 2864 9088 2868 9092
rect 2872 9088 2876 9092
rect 2880 9088 2884 9092
rect 2888 9088 2892 9092
rect 2896 9088 2900 9092
rect 2907 9088 2911 9092
rect 2924 9088 2928 9092
rect 2941 9088 2945 9092
rect 2950 9088 2954 9092
rect 2963 9088 2967 9092
rect 2971 9088 2975 9092
rect 2979 9088 2983 9092
rect 2996 9088 3000 9092
rect 3006 9088 3010 9092
rect 3014 9088 3018 9092
rect 3189 9093 3193 9097
rect 3197 9093 3201 9097
rect 3366 9072 3370 9076
rect 3374 9072 3378 9076
rect 3390 9068 3394 9072
rect 3405 9068 3409 9072
rect 3420 9064 3424 9068
rect 3428 9064 3432 9068
rect 3999 9097 4003 9101
rect 4014 9097 4018 9101
rect 4080 9101 4084 9105
rect 4088 9101 4092 9105
rect 4104 9097 4108 9101
rect 4119 9097 4123 9101
rect 4029 9093 4033 9097
rect 4037 9093 4041 9097
rect 3801 9088 3805 9092
rect 3809 9088 3813 9092
rect 3817 9088 3821 9092
rect 3825 9088 3829 9092
rect 3833 9088 3837 9092
rect 3841 9088 3845 9092
rect 3852 9088 3856 9092
rect 3869 9088 3873 9092
rect 3886 9088 3890 9092
rect 3895 9088 3899 9092
rect 3908 9088 3912 9092
rect 3916 9088 3920 9092
rect 3924 9088 3928 9092
rect 3941 9088 3945 9092
rect 3951 9088 3955 9092
rect 3959 9088 3963 9092
rect 4134 9093 4138 9097
rect 4142 9093 4146 9097
rect 2856 9042 2860 9046
rect 2864 9042 2868 9046
rect 2872 9042 2876 9046
rect 2880 9042 2884 9046
rect 2888 9042 2892 9046
rect 2896 9042 2900 9046
rect 2907 9042 2911 9046
rect 2924 9042 2928 9046
rect 2941 9042 2945 9046
rect 2950 9042 2954 9046
rect 2963 9042 2967 9046
rect 2971 9042 2975 9046
rect 2979 9042 2983 9046
rect 2996 9042 3000 9046
rect 3006 9042 3010 9046
rect 3014 9042 3018 9046
rect 3054 9042 3058 9046
rect 3069 9042 3073 9046
rect 3159 9042 3163 9046
rect 3174 9042 3178 9046
rect 3540 9033 3556 9045
rect 3560 9033 3576 9045
rect 3593 9033 3609 9045
rect 3613 9033 3629 9045
rect 3801 9042 3805 9046
rect 3809 9042 3813 9046
rect 3817 9042 3821 9046
rect 3825 9042 3829 9046
rect 3833 9042 3837 9046
rect 3841 9042 3845 9046
rect 3852 9042 3856 9046
rect 3869 9042 3873 9046
rect 3886 9042 3890 9046
rect 3895 9042 3899 9046
rect 3908 9042 3912 9046
rect 3916 9042 3920 9046
rect 3924 9042 3928 9046
rect 3941 9042 3945 9046
rect 3951 9042 3955 9046
rect 3959 9042 3963 9046
rect 3999 9042 4003 9046
rect 4014 9042 4018 9046
rect 4104 9042 4108 9046
rect 4119 9042 4123 9046
rect 3390 9008 3394 9012
rect 3405 9008 3409 9012
rect 3054 8965 3058 8969
rect 3069 8965 3073 8969
rect 3111 8969 3115 8973
rect 3119 8969 3123 8973
rect 3135 8965 3139 8969
rect 3150 8965 3154 8969
rect 3201 8969 3205 8973
rect 3209 8969 3213 8973
rect 3225 8965 3229 8969
rect 3240 8965 3244 8969
rect 3084 8961 3088 8965
rect 3092 8961 3096 8965
rect 2856 8956 2860 8960
rect 2864 8956 2868 8960
rect 2872 8956 2876 8960
rect 2880 8956 2884 8960
rect 2888 8956 2892 8960
rect 2896 8956 2900 8960
rect 2907 8956 2911 8960
rect 2924 8956 2928 8960
rect 2941 8956 2945 8960
rect 2950 8956 2954 8960
rect 2963 8956 2967 8960
rect 2971 8956 2975 8960
rect 2979 8956 2983 8960
rect 2996 8956 3000 8960
rect 3006 8956 3010 8960
rect 3014 8956 3018 8960
rect 3165 8961 3169 8965
rect 3173 8961 3177 8965
rect 3255 8961 3259 8965
rect 3263 8961 3267 8965
rect 3344 8942 3348 8946
rect 3352 8942 3356 8946
rect 3366 8942 3370 8946
rect 3374 8942 3378 8946
rect 3390 8938 3394 8942
rect 3405 8938 3409 8942
rect 3420 8934 3424 8938
rect 3428 8934 3432 8938
rect 3999 8965 4003 8969
rect 4014 8965 4018 8969
rect 4056 8969 4060 8973
rect 4064 8969 4068 8973
rect 4080 8965 4084 8969
rect 4095 8965 4099 8969
rect 4146 8969 4150 8973
rect 4154 8969 4158 8973
rect 4170 8965 4174 8969
rect 4185 8965 4189 8969
rect 4029 8961 4033 8965
rect 4037 8961 4041 8965
rect 3801 8956 3805 8960
rect 3809 8956 3813 8960
rect 3817 8956 3821 8960
rect 3825 8956 3829 8960
rect 3833 8956 3837 8960
rect 3841 8956 3845 8960
rect 3852 8956 3856 8960
rect 3869 8956 3873 8960
rect 3886 8956 3890 8960
rect 3895 8956 3899 8960
rect 3908 8956 3912 8960
rect 3916 8956 3920 8960
rect 3924 8956 3928 8960
rect 3941 8956 3945 8960
rect 3951 8956 3955 8960
rect 3959 8956 3963 8960
rect 4110 8961 4114 8965
rect 4118 8961 4122 8965
rect 4200 8961 4204 8965
rect 4208 8961 4212 8965
rect 2856 8910 2860 8914
rect 2864 8910 2868 8914
rect 2872 8910 2876 8914
rect 2880 8910 2884 8914
rect 2888 8910 2892 8914
rect 2896 8910 2900 8914
rect 2907 8910 2911 8914
rect 2924 8910 2928 8914
rect 2941 8910 2945 8914
rect 2950 8910 2954 8914
rect 2963 8910 2967 8914
rect 2971 8910 2975 8914
rect 2979 8910 2983 8914
rect 2996 8910 3000 8914
rect 3006 8910 3010 8914
rect 3014 8910 3018 8914
rect 3054 8907 3058 8911
rect 3069 8907 3073 8911
rect 3135 8907 3139 8911
rect 3150 8907 3154 8911
rect 3225 8907 3229 8911
rect 3240 8907 3244 8911
rect 3446 8903 3462 8915
rect 3466 8903 3482 8915
rect 3499 8903 3515 8915
rect 3519 8903 3535 8915
rect 3801 8910 3805 8914
rect 3809 8910 3813 8914
rect 3817 8910 3821 8914
rect 3825 8910 3829 8914
rect 3833 8910 3837 8914
rect 3841 8910 3845 8914
rect 3852 8910 3856 8914
rect 3869 8910 3873 8914
rect 3886 8910 3890 8914
rect 3895 8910 3899 8914
rect 3908 8910 3912 8914
rect 3916 8910 3920 8914
rect 3924 8910 3928 8914
rect 3941 8910 3945 8914
rect 3951 8910 3955 8914
rect 3959 8910 3963 8914
rect 3999 8907 4003 8911
rect 4014 8907 4018 8911
rect 4080 8907 4084 8911
rect 4095 8907 4099 8911
rect 4170 8907 4174 8911
rect 4185 8907 4189 8911
rect 3390 8878 3394 8882
rect 3405 8878 3409 8882
rect 3054 8833 3058 8837
rect 3069 8833 3073 8837
rect 3084 8829 3088 8833
rect 3092 8829 3096 8833
rect 2856 8824 2860 8828
rect 2864 8824 2868 8828
rect 2872 8824 2876 8828
rect 2880 8824 2884 8828
rect 2888 8824 2892 8828
rect 2896 8824 2900 8828
rect 2907 8824 2911 8828
rect 2924 8824 2928 8828
rect 2941 8824 2945 8828
rect 2950 8824 2954 8828
rect 2963 8824 2967 8828
rect 2971 8824 2975 8828
rect 2979 8824 2983 8828
rect 2996 8824 3000 8828
rect 3006 8824 3010 8828
rect 3014 8824 3018 8828
rect 3999 8833 4003 8837
rect 4014 8833 4018 8837
rect 4029 8829 4033 8833
rect 4037 8829 4041 8833
rect 3801 8824 3805 8828
rect 3809 8824 3813 8828
rect 3817 8824 3821 8828
rect 3825 8824 3829 8828
rect 3833 8824 3837 8828
rect 3841 8824 3845 8828
rect 3852 8824 3856 8828
rect 3869 8824 3873 8828
rect 3886 8824 3890 8828
rect 3895 8824 3899 8828
rect 3908 8824 3912 8828
rect 3916 8824 3920 8828
rect 3924 8824 3928 8828
rect 3941 8824 3945 8828
rect 3951 8824 3955 8828
rect 3959 8824 3963 8828
rect 2856 8778 2860 8782
rect 2864 8778 2868 8782
rect 2872 8778 2876 8782
rect 2880 8778 2884 8782
rect 2888 8778 2892 8782
rect 2896 8778 2900 8782
rect 2907 8778 2911 8782
rect 2924 8778 2928 8782
rect 2941 8778 2945 8782
rect 2950 8778 2954 8782
rect 2963 8778 2967 8782
rect 2971 8778 2975 8782
rect 2979 8778 2983 8782
rect 2996 8778 3000 8782
rect 3006 8778 3010 8782
rect 3014 8778 3018 8782
rect 3090 8778 3094 8782
rect 3098 8778 3102 8782
rect 3108 8778 3112 8782
rect 3116 8778 3120 8782
rect 3125 8778 3129 8782
rect 3133 8778 3137 8782
rect 3141 8778 3145 8782
rect 3149 8778 3153 8782
rect 3157 8778 3161 8782
rect 3168 8778 3172 8782
rect 3185 8778 3189 8782
rect 3202 8778 3206 8782
rect 3211 8778 3215 8782
rect 3224 8778 3228 8782
rect 3232 8778 3236 8782
rect 3240 8778 3244 8782
rect 3257 8778 3261 8782
rect 3267 8778 3271 8782
rect 3275 8778 3279 8782
rect 2367 8764 2371 8768
rect 2380 8764 2384 8768
rect 2388 8764 2392 8768
rect 2396 8764 2400 8768
rect 2404 8764 2408 8768
rect 2417 8764 2421 8768
rect 2430 8764 2434 8768
rect 2438 8764 2442 8768
rect 2446 8764 2450 8768
rect 2454 8764 2458 8768
rect 2462 8764 2466 8768
rect 2475 8764 2479 8768
rect 2483 8764 2487 8768
rect 2491 8764 2495 8768
rect 2499 8764 2503 8768
rect 2512 8764 2516 8768
rect 2520 8764 2524 8768
rect 2528 8764 2532 8768
rect 2536 8764 2540 8768
rect 2549 8764 2553 8768
rect 2562 8764 2566 8768
rect 2570 8764 2574 8768
rect 2578 8764 2582 8768
rect 2586 8764 2590 8768
rect 2594 8764 2598 8768
rect 2607 8764 2611 8768
rect 2615 8764 2619 8768
rect 2623 8764 2627 8768
rect 2631 8764 2635 8768
rect 2644 8764 2648 8768
rect 2652 8764 2656 8768
rect 2660 8764 2664 8768
rect 2668 8764 2672 8768
rect 2681 8764 2685 8768
rect 2694 8764 2698 8768
rect 2702 8764 2706 8768
rect 2710 8764 2714 8768
rect 2718 8764 2722 8768
rect 2726 8764 2730 8768
rect 2739 8764 2743 8768
rect 2747 8764 2751 8768
rect 2755 8764 2759 8768
rect 3054 8771 3058 8775
rect 3069 8771 3073 8775
rect 3801 8778 3805 8782
rect 3809 8778 3813 8782
rect 3817 8778 3821 8782
rect 3825 8778 3829 8782
rect 3833 8778 3837 8782
rect 3841 8778 3845 8782
rect 3852 8778 3856 8782
rect 3869 8778 3873 8782
rect 3886 8778 3890 8782
rect 3895 8778 3899 8782
rect 3908 8778 3912 8782
rect 3916 8778 3920 8782
rect 3924 8778 3928 8782
rect 3941 8778 3945 8782
rect 3951 8778 3955 8782
rect 3959 8778 3963 8782
rect 4035 8778 4039 8782
rect 4043 8778 4047 8782
rect 4053 8778 4057 8782
rect 4061 8778 4065 8782
rect 4070 8778 4074 8782
rect 4078 8778 4082 8782
rect 4086 8778 4090 8782
rect 4094 8778 4098 8782
rect 4102 8778 4106 8782
rect 4113 8778 4117 8782
rect 4130 8778 4134 8782
rect 4147 8778 4151 8782
rect 4156 8778 4160 8782
rect 4169 8778 4173 8782
rect 4177 8778 4181 8782
rect 4185 8778 4189 8782
rect 4202 8778 4206 8782
rect 4212 8778 4216 8782
rect 4220 8778 4224 8782
rect 3312 8764 3316 8768
rect 3325 8764 3329 8768
rect 3333 8764 3337 8768
rect 3341 8764 3345 8768
rect 3349 8764 3353 8768
rect 3362 8764 3366 8768
rect 3375 8764 3379 8768
rect 3383 8764 3387 8768
rect 3391 8764 3395 8768
rect 3399 8764 3403 8768
rect 3407 8764 3411 8768
rect 3420 8764 3424 8768
rect 3428 8764 3432 8768
rect 3436 8764 3440 8768
rect 3444 8764 3448 8768
rect 3457 8764 3461 8768
rect 3465 8764 3469 8768
rect 3473 8764 3477 8768
rect 3481 8764 3485 8768
rect 3494 8764 3498 8768
rect 3507 8764 3511 8768
rect 3515 8764 3519 8768
rect 3523 8764 3527 8768
rect 3531 8764 3535 8768
rect 3539 8764 3543 8768
rect 3552 8764 3556 8768
rect 3560 8764 3564 8768
rect 3568 8764 3572 8768
rect 3576 8764 3580 8768
rect 3589 8764 3593 8768
rect 3597 8764 3601 8768
rect 3605 8764 3609 8768
rect 3613 8764 3617 8768
rect 3626 8764 3630 8768
rect 3639 8764 3643 8768
rect 3647 8764 3651 8768
rect 3655 8764 3659 8768
rect 3663 8764 3667 8768
rect 3671 8764 3675 8768
rect 3684 8764 3688 8768
rect 3692 8764 3696 8768
rect 3700 8764 3704 8768
rect 3999 8771 4003 8775
rect 4014 8771 4018 8775
rect 2482 8720 2486 8724
rect 2490 8720 2494 8724
rect 2506 8720 2510 8724
rect 2514 8720 2518 8724
rect 3284 8725 3288 8729
rect 3284 8716 3288 8721
rect 3427 8720 3431 8724
rect 3435 8720 3439 8724
rect 3451 8720 3455 8724
rect 3459 8720 3463 8724
rect 4229 8725 4233 8729
rect 4229 8716 4233 8721
rect 2502 8707 2506 8711
rect 2510 8707 2514 8711
rect 3447 8707 3451 8711
rect 3455 8707 3459 8711
rect 2498 8696 2502 8700
rect 3443 8696 3447 8700
rect 2498 8688 2502 8692
rect 2482 8684 2486 8688
rect 2490 8684 2494 8688
rect 2506 8684 2510 8688
rect 2514 8684 2518 8688
rect 3443 8688 3447 8692
rect 3427 8684 3431 8688
rect 3435 8684 3439 8688
rect 3451 8684 3455 8688
rect 3459 8684 3463 8688
rect 3150 8652 3154 8656
rect 3163 8652 3167 8656
rect 3171 8652 3175 8656
rect 3179 8652 3183 8656
rect 3187 8652 3191 8656
rect 3200 8652 3204 8656
rect 3213 8652 3217 8656
rect 3221 8652 3225 8656
rect 3229 8652 3233 8656
rect 3237 8652 3241 8656
rect 3245 8652 3249 8656
rect 3258 8652 3262 8656
rect 3266 8652 3270 8656
rect 3274 8652 3278 8656
rect 4095 8652 4099 8656
rect 4108 8652 4112 8656
rect 4116 8652 4120 8656
rect 4124 8652 4128 8656
rect 4132 8652 4136 8656
rect 4145 8652 4149 8656
rect 4158 8652 4162 8656
rect 4166 8652 4170 8656
rect 4174 8652 4178 8656
rect 4182 8652 4186 8656
rect 4190 8652 4194 8656
rect 4203 8652 4207 8656
rect 4211 8652 4215 8656
rect 4219 8652 4223 8656
rect 2367 8622 2371 8626
rect 2380 8622 2384 8626
rect 2388 8622 2392 8626
rect 2396 8622 2400 8626
rect 2404 8622 2408 8626
rect 2417 8622 2421 8626
rect 2430 8622 2434 8626
rect 2438 8622 2442 8626
rect 2446 8622 2450 8626
rect 2454 8622 2458 8626
rect 2462 8622 2466 8626
rect 2475 8622 2479 8626
rect 2483 8622 2487 8626
rect 2491 8622 2495 8626
rect 2499 8622 2503 8626
rect 2512 8622 2516 8626
rect 2520 8622 2524 8626
rect 2528 8622 2532 8626
rect 2536 8622 2540 8626
rect 2549 8622 2553 8626
rect 2562 8622 2566 8626
rect 2570 8622 2574 8626
rect 2578 8622 2582 8626
rect 2586 8622 2590 8626
rect 2594 8622 2598 8626
rect 2607 8622 2611 8626
rect 2615 8622 2619 8626
rect 2623 8622 2627 8626
rect 2631 8622 2635 8626
rect 2644 8622 2648 8626
rect 2652 8622 2656 8626
rect 2660 8622 2664 8626
rect 2668 8622 2672 8626
rect 2681 8622 2685 8626
rect 2694 8622 2698 8626
rect 2702 8622 2706 8626
rect 2710 8622 2714 8626
rect 2718 8622 2722 8626
rect 2726 8622 2730 8626
rect 2739 8622 2743 8626
rect 2747 8622 2751 8626
rect 2755 8622 2759 8626
rect 3312 8622 3316 8626
rect 3325 8622 3329 8626
rect 3333 8622 3337 8626
rect 3341 8622 3345 8626
rect 3349 8622 3353 8626
rect 3362 8622 3366 8626
rect 3375 8622 3379 8626
rect 3383 8622 3387 8626
rect 3391 8622 3395 8626
rect 3399 8622 3403 8626
rect 3407 8622 3411 8626
rect 3420 8622 3424 8626
rect 3428 8622 3432 8626
rect 3436 8622 3440 8626
rect 3444 8622 3448 8626
rect 3457 8622 3461 8626
rect 3465 8622 3469 8626
rect 3473 8622 3477 8626
rect 3481 8622 3485 8626
rect 3494 8622 3498 8626
rect 3507 8622 3511 8626
rect 3515 8622 3519 8626
rect 3523 8622 3527 8626
rect 3531 8622 3535 8626
rect 3539 8622 3543 8626
rect 3552 8622 3556 8626
rect 3560 8622 3564 8626
rect 3568 8622 3572 8626
rect 3576 8622 3580 8626
rect 3589 8622 3593 8626
rect 3597 8622 3601 8626
rect 3605 8622 3609 8626
rect 3613 8622 3617 8626
rect 3626 8622 3630 8626
rect 3639 8622 3643 8626
rect 3647 8622 3651 8626
rect 3655 8622 3659 8626
rect 3663 8622 3667 8626
rect 3671 8622 3675 8626
rect 3684 8622 3688 8626
rect 3692 8622 3696 8626
rect 3700 8622 3704 8626
rect 3296 8579 3300 8583
rect 3296 8571 3300 8575
rect 4241 8579 4245 8583
rect 4241 8571 4245 8575
rect 3150 8566 3154 8570
rect 3163 8566 3167 8570
rect 3171 8566 3175 8570
rect 3179 8566 3183 8570
rect 3187 8566 3191 8570
rect 3200 8566 3204 8570
rect 3213 8566 3217 8570
rect 3221 8566 3225 8570
rect 3229 8566 3233 8570
rect 3237 8566 3241 8570
rect 3245 8566 3249 8570
rect 3258 8566 3262 8570
rect 3266 8566 3270 8570
rect 3274 8566 3278 8570
rect 4095 8566 4099 8570
rect 4108 8566 4112 8570
rect 4116 8566 4120 8570
rect 4124 8566 4128 8570
rect 4132 8566 4136 8570
rect 4145 8566 4149 8570
rect 4158 8566 4162 8570
rect 4166 8566 4170 8570
rect 4174 8566 4178 8570
rect 4182 8566 4186 8570
rect 4190 8566 4194 8570
rect 4203 8566 4207 8570
rect 4211 8566 4215 8570
rect 4219 8566 4223 8570
rect 2367 8536 2371 8540
rect 2380 8536 2384 8540
rect 2388 8536 2392 8540
rect 2396 8536 2400 8540
rect 2404 8536 2408 8540
rect 2417 8536 2421 8540
rect 2430 8536 2434 8540
rect 2438 8536 2442 8540
rect 2446 8536 2450 8540
rect 2454 8536 2458 8540
rect 2462 8536 2466 8540
rect 2475 8536 2479 8540
rect 2483 8536 2487 8540
rect 2491 8536 2495 8540
rect 2499 8536 2503 8540
rect 2512 8536 2516 8540
rect 2520 8536 2524 8540
rect 2528 8536 2532 8540
rect 2536 8536 2540 8540
rect 2549 8536 2553 8540
rect 2562 8536 2566 8540
rect 2570 8536 2574 8540
rect 2578 8536 2582 8540
rect 2586 8536 2590 8540
rect 2594 8536 2598 8540
rect 2607 8536 2611 8540
rect 2615 8536 2619 8540
rect 2623 8536 2627 8540
rect 2631 8536 2635 8540
rect 2644 8536 2648 8540
rect 2652 8536 2656 8540
rect 2660 8536 2664 8540
rect 2668 8536 2672 8540
rect 2681 8536 2685 8540
rect 2694 8536 2698 8540
rect 2702 8536 2706 8540
rect 2710 8536 2714 8540
rect 2718 8536 2722 8540
rect 2726 8536 2730 8540
rect 2739 8536 2743 8540
rect 2747 8536 2751 8540
rect 2755 8536 2759 8540
rect 3312 8536 3316 8540
rect 3325 8536 3329 8540
rect 3333 8536 3337 8540
rect 3341 8536 3345 8540
rect 3349 8536 3353 8540
rect 3362 8536 3366 8540
rect 3375 8536 3379 8540
rect 3383 8536 3387 8540
rect 3391 8536 3395 8540
rect 3399 8536 3403 8540
rect 3407 8536 3411 8540
rect 3420 8536 3424 8540
rect 3428 8536 3432 8540
rect 3436 8536 3440 8540
rect 3444 8536 3448 8540
rect 3457 8536 3461 8540
rect 3465 8536 3469 8540
rect 3473 8536 3477 8540
rect 3481 8536 3485 8540
rect 3494 8536 3498 8540
rect 3507 8536 3511 8540
rect 3515 8536 3519 8540
rect 3523 8536 3527 8540
rect 3531 8536 3535 8540
rect 3539 8536 3543 8540
rect 3552 8536 3556 8540
rect 3560 8536 3564 8540
rect 3568 8536 3572 8540
rect 3576 8536 3580 8540
rect 3589 8536 3593 8540
rect 3597 8536 3601 8540
rect 3605 8536 3609 8540
rect 3613 8536 3617 8540
rect 3626 8536 3630 8540
rect 3639 8536 3643 8540
rect 3647 8536 3651 8540
rect 3655 8536 3659 8540
rect 3663 8536 3667 8540
rect 3671 8536 3675 8540
rect 3684 8536 3688 8540
rect 3692 8536 3696 8540
rect 3700 8536 3704 8540
rect 2599 8492 2603 8496
rect 2607 8492 2611 8496
rect 2623 8492 2627 8496
rect 2631 8492 2635 8496
rect 3544 8492 3548 8496
rect 3552 8492 3556 8496
rect 3568 8492 3572 8496
rect 3576 8492 3580 8496
rect 2619 8481 2623 8485
rect 2627 8481 2631 8485
rect 3564 8481 3568 8485
rect 3572 8481 3576 8485
rect 2615 8470 2619 8474
rect 3560 8470 3564 8474
rect 2615 8462 2619 8466
rect 3560 8462 3564 8466
rect 2599 8458 2603 8462
rect 2607 8458 2611 8462
rect 2623 8458 2627 8462
rect 2631 8458 2635 8462
rect 3544 8458 3548 8462
rect 3552 8458 3556 8462
rect 3568 8458 3572 8462
rect 3576 8458 3580 8462
rect 2367 8396 2371 8400
rect 2380 8396 2384 8400
rect 2388 8396 2392 8400
rect 2396 8396 2400 8400
rect 2404 8396 2408 8400
rect 2417 8396 2421 8400
rect 2430 8396 2434 8400
rect 2438 8396 2442 8400
rect 2446 8396 2450 8400
rect 2454 8396 2458 8400
rect 2462 8396 2466 8400
rect 2475 8396 2479 8400
rect 2483 8396 2487 8400
rect 2491 8396 2495 8400
rect 2499 8396 2503 8400
rect 2512 8396 2516 8400
rect 2520 8396 2524 8400
rect 2528 8396 2532 8400
rect 2536 8396 2540 8400
rect 2549 8396 2553 8400
rect 2562 8396 2566 8400
rect 2570 8396 2574 8400
rect 2578 8396 2582 8400
rect 2586 8396 2590 8400
rect 2594 8396 2598 8400
rect 2607 8396 2611 8400
rect 2615 8396 2619 8400
rect 2623 8396 2627 8400
rect 2631 8396 2635 8400
rect 2644 8396 2648 8400
rect 2652 8396 2656 8400
rect 2660 8396 2664 8400
rect 2668 8396 2672 8400
rect 2681 8396 2685 8400
rect 2694 8396 2698 8400
rect 2702 8396 2706 8400
rect 2710 8396 2714 8400
rect 2718 8396 2722 8400
rect 2726 8396 2730 8400
rect 2739 8396 2743 8400
rect 2747 8396 2751 8400
rect 2755 8396 2759 8400
rect 3312 8396 3316 8400
rect 3325 8396 3329 8400
rect 3333 8396 3337 8400
rect 3341 8396 3345 8400
rect 3349 8396 3353 8400
rect 3362 8396 3366 8400
rect 3375 8396 3379 8400
rect 3383 8396 3387 8400
rect 3391 8396 3395 8400
rect 3399 8396 3403 8400
rect 3407 8396 3411 8400
rect 3420 8396 3424 8400
rect 3428 8396 3432 8400
rect 3436 8396 3440 8400
rect 3444 8396 3448 8400
rect 3457 8396 3461 8400
rect 3465 8396 3469 8400
rect 3473 8396 3477 8400
rect 3481 8396 3485 8400
rect 3494 8396 3498 8400
rect 3507 8396 3511 8400
rect 3515 8396 3519 8400
rect 3523 8396 3527 8400
rect 3531 8396 3535 8400
rect 3539 8396 3543 8400
rect 3552 8396 3556 8400
rect 3560 8396 3564 8400
rect 3568 8396 3572 8400
rect 3576 8396 3580 8400
rect 3589 8396 3593 8400
rect 3597 8396 3601 8400
rect 3605 8396 3609 8400
rect 3613 8396 3617 8400
rect 3626 8396 3630 8400
rect 3639 8396 3643 8400
rect 3647 8396 3651 8400
rect 3655 8396 3659 8400
rect 3663 8396 3667 8400
rect 3671 8396 3675 8400
rect 3684 8396 3688 8400
rect 3692 8396 3696 8400
rect 3700 8396 3704 8400
rect 2851 8317 2855 8321
rect 2864 8317 2868 8321
rect 2872 8317 2876 8321
rect 2880 8317 2884 8321
rect 2888 8317 2892 8321
rect 2901 8317 2905 8321
rect 2914 8317 2918 8321
rect 2922 8317 2926 8321
rect 2930 8317 2934 8321
rect 2938 8317 2942 8321
rect 2946 8317 2950 8321
rect 2959 8317 2963 8321
rect 2967 8317 2971 8321
rect 2975 8317 2979 8321
rect 2983 8317 2987 8321
rect 2996 8317 3000 8321
rect 3004 8317 3008 8321
rect 3012 8317 3016 8321
rect 3020 8317 3024 8321
rect 3033 8317 3037 8321
rect 3046 8317 3050 8321
rect 3054 8317 3058 8321
rect 3062 8317 3066 8321
rect 3070 8317 3074 8321
rect 3078 8317 3082 8321
rect 3091 8317 3095 8321
rect 3099 8317 3103 8321
rect 3107 8317 3111 8321
rect 3115 8317 3119 8321
rect 3128 8317 3132 8321
rect 3136 8317 3140 8321
rect 3144 8317 3148 8321
rect 3152 8317 3156 8321
rect 3165 8317 3169 8321
rect 3178 8317 3182 8321
rect 3186 8317 3190 8321
rect 3194 8317 3198 8321
rect 3202 8317 3206 8321
rect 3210 8317 3214 8321
rect 3223 8317 3227 8321
rect 3231 8317 3235 8321
rect 3239 8317 3243 8321
rect 3247 8317 3251 8321
rect 3260 8317 3264 8321
rect 3268 8317 3272 8321
rect 3276 8317 3280 8321
rect 3284 8317 3288 8321
rect 3297 8317 3301 8321
rect 3310 8317 3314 8321
rect 3318 8317 3322 8321
rect 3326 8317 3330 8321
rect 3334 8317 3338 8321
rect 3342 8317 3346 8321
rect 3355 8317 3359 8321
rect 3363 8317 3367 8321
rect 3371 8317 3375 8321
rect 3796 8317 3800 8321
rect 3809 8317 3813 8321
rect 3817 8317 3821 8321
rect 3825 8317 3829 8321
rect 3833 8317 3837 8321
rect 3846 8317 3850 8321
rect 3859 8317 3863 8321
rect 3867 8317 3871 8321
rect 3875 8317 3879 8321
rect 3883 8317 3887 8321
rect 3891 8317 3895 8321
rect 3904 8317 3908 8321
rect 3912 8317 3916 8321
rect 3920 8317 3924 8321
rect 3928 8317 3932 8321
rect 3941 8317 3945 8321
rect 3949 8317 3953 8321
rect 3957 8317 3961 8321
rect 3965 8317 3969 8321
rect 3978 8317 3982 8321
rect 3991 8317 3995 8321
rect 3999 8317 4003 8321
rect 4007 8317 4011 8321
rect 4015 8317 4019 8321
rect 4023 8317 4027 8321
rect 4036 8317 4040 8321
rect 4044 8317 4048 8321
rect 4052 8317 4056 8321
rect 4060 8317 4064 8321
rect 4073 8317 4077 8321
rect 4081 8317 4085 8321
rect 4089 8317 4093 8321
rect 4097 8317 4101 8321
rect 4110 8317 4114 8321
rect 4123 8317 4127 8321
rect 4131 8317 4135 8321
rect 4139 8317 4143 8321
rect 4147 8317 4151 8321
rect 4155 8317 4159 8321
rect 4168 8317 4172 8321
rect 4176 8317 4180 8321
rect 4184 8317 4188 8321
rect 4192 8317 4196 8321
rect 4205 8317 4209 8321
rect 4213 8317 4217 8321
rect 4221 8317 4225 8321
rect 4229 8317 4233 8321
rect 4242 8317 4246 8321
rect 4255 8317 4259 8321
rect 4263 8317 4267 8321
rect 4271 8317 4275 8321
rect 4279 8317 4283 8321
rect 4287 8317 4291 8321
rect 4300 8317 4304 8321
rect 4308 8317 4312 8321
rect 4316 8317 4320 8321
rect 2499 8284 2503 8288
rect 2512 8284 2516 8288
rect 2520 8284 2524 8288
rect 2528 8284 2532 8288
rect 2536 8284 2540 8288
rect 2549 8284 2553 8288
rect 2562 8284 2566 8288
rect 2570 8284 2574 8288
rect 2578 8284 2582 8288
rect 2586 8284 2590 8288
rect 2594 8284 2598 8288
rect 2607 8284 2611 8288
rect 2615 8284 2619 8288
rect 2623 8284 2627 8288
rect 3444 8284 3448 8288
rect 3457 8284 3461 8288
rect 3465 8284 3469 8288
rect 3473 8284 3477 8288
rect 3481 8284 3485 8288
rect 3494 8284 3498 8288
rect 3507 8284 3511 8288
rect 3515 8284 3519 8288
rect 3523 8284 3527 8288
rect 3531 8284 3535 8288
rect 3539 8284 3543 8288
rect 3552 8284 3556 8288
rect 3560 8284 3564 8288
rect 3568 8284 3572 8288
rect 2623 8247 2627 8251
rect 2631 8247 2635 8251
rect 3030 8251 3034 8255
rect 3038 8251 3042 8255
rect 3054 8247 3058 8251
rect 3069 8247 3073 8251
rect 3111 8251 3115 8255
rect 3119 8251 3123 8255
rect 3135 8247 3139 8251
rect 3150 8247 3154 8251
rect 3084 8243 3088 8247
rect 3092 8243 3096 8247
rect 2506 8238 2510 8242
rect 2514 8238 2518 8242
rect 2856 8238 2860 8242
rect 2864 8238 2868 8242
rect 2872 8238 2876 8242
rect 2880 8238 2884 8242
rect 2888 8238 2892 8242
rect 2896 8238 2900 8242
rect 2907 8238 2911 8242
rect 2924 8238 2928 8242
rect 2941 8238 2945 8242
rect 2950 8238 2954 8242
rect 2963 8238 2967 8242
rect 2971 8238 2975 8242
rect 2979 8238 2983 8242
rect 2996 8238 3000 8242
rect 3006 8238 3010 8242
rect 3014 8238 3018 8242
rect 3165 8243 3169 8247
rect 3173 8243 3177 8247
rect 3568 8247 3572 8251
rect 3576 8247 3580 8251
rect 3975 8251 3979 8255
rect 3983 8251 3987 8255
rect 3999 8247 4003 8251
rect 4014 8247 4018 8251
rect 4056 8251 4060 8255
rect 4064 8251 4068 8255
rect 4080 8247 4084 8251
rect 4095 8247 4099 8251
rect 4029 8243 4033 8247
rect 4037 8243 4041 8247
rect 3451 8238 3455 8242
rect 3459 8238 3463 8242
rect 3801 8238 3805 8242
rect 3809 8238 3813 8242
rect 3817 8238 3821 8242
rect 3825 8238 3829 8242
rect 3833 8238 3837 8242
rect 3841 8238 3845 8242
rect 3852 8238 3856 8242
rect 3869 8238 3873 8242
rect 3886 8238 3890 8242
rect 3895 8238 3899 8242
rect 3908 8238 3912 8242
rect 3916 8238 3920 8242
rect 3924 8238 3928 8242
rect 3941 8238 3945 8242
rect 3951 8238 3955 8242
rect 3959 8238 3963 8242
rect 4110 8243 4114 8247
rect 4118 8243 4122 8247
rect 2856 8192 2860 8196
rect 2864 8192 2868 8196
rect 2872 8192 2876 8196
rect 2880 8192 2884 8196
rect 2888 8192 2892 8196
rect 2896 8192 2900 8196
rect 2907 8192 2911 8196
rect 2924 8192 2928 8196
rect 2941 8192 2945 8196
rect 2950 8192 2954 8196
rect 2963 8192 2967 8196
rect 2971 8192 2975 8196
rect 2979 8192 2983 8196
rect 2996 8192 3000 8196
rect 3006 8192 3010 8196
rect 3014 8192 3018 8196
rect 2490 8182 2494 8186
rect 2498 8182 2502 8186
rect 2506 8182 2510 8186
rect 2519 8182 2523 8186
rect 2527 8182 2531 8186
rect 2535 8182 2539 8186
rect 2543 8182 2547 8186
rect 2551 8182 2555 8186
rect 2564 8182 2568 8186
rect 2577 8182 2581 8186
rect 2585 8182 2589 8186
rect 2593 8182 2597 8186
rect 2601 8182 2605 8186
rect 2614 8182 2618 8186
rect 3054 8191 3058 8195
rect 3069 8191 3073 8195
rect 3135 8191 3139 8195
rect 3150 8191 3154 8195
rect 3801 8192 3805 8196
rect 3809 8192 3813 8196
rect 3817 8192 3821 8196
rect 3825 8192 3829 8196
rect 3833 8192 3837 8196
rect 3841 8192 3845 8196
rect 3852 8192 3856 8196
rect 3869 8192 3873 8196
rect 3886 8192 3890 8196
rect 3895 8192 3899 8196
rect 3908 8192 3912 8196
rect 3916 8192 3920 8196
rect 3924 8192 3928 8196
rect 3941 8192 3945 8196
rect 3951 8192 3955 8196
rect 3959 8192 3963 8196
rect 3435 8182 3439 8186
rect 3443 8182 3447 8186
rect 3451 8182 3455 8186
rect 3464 8182 3468 8186
rect 3472 8182 3476 8186
rect 3480 8182 3484 8186
rect 3488 8182 3492 8186
rect 3496 8182 3500 8186
rect 3509 8182 3513 8186
rect 3522 8182 3526 8186
rect 3530 8182 3534 8186
rect 3538 8182 3542 8186
rect 3546 8182 3550 8186
rect 3559 8182 3563 8186
rect 3999 8191 4003 8195
rect 4014 8191 4018 8195
rect 4080 8191 4084 8195
rect 4095 8191 4099 8195
rect 3054 8115 3058 8119
rect 3069 8115 3073 8119
rect 3135 8119 3139 8123
rect 3143 8119 3147 8123
rect 3159 8115 3163 8119
rect 3174 8115 3178 8119
rect 3084 8111 3088 8115
rect 3092 8111 3096 8115
rect 2856 8106 2860 8110
rect 2864 8106 2868 8110
rect 2872 8106 2876 8110
rect 2880 8106 2884 8110
rect 2888 8106 2892 8110
rect 2896 8106 2900 8110
rect 2907 8106 2911 8110
rect 2924 8106 2928 8110
rect 2941 8106 2945 8110
rect 2950 8106 2954 8110
rect 2963 8106 2967 8110
rect 2971 8106 2975 8110
rect 2979 8106 2983 8110
rect 2996 8106 3000 8110
rect 3006 8106 3010 8110
rect 3014 8106 3018 8110
rect 3189 8111 3193 8115
rect 3197 8111 3201 8115
rect 3999 8115 4003 8119
rect 4014 8115 4018 8119
rect 4080 8119 4084 8123
rect 4088 8119 4092 8123
rect 4104 8115 4108 8119
rect 4119 8115 4123 8119
rect 4029 8111 4033 8115
rect 4037 8111 4041 8115
rect 3801 8106 3805 8110
rect 3809 8106 3813 8110
rect 3817 8106 3821 8110
rect 3825 8106 3829 8110
rect 3833 8106 3837 8110
rect 3841 8106 3845 8110
rect 3852 8106 3856 8110
rect 3869 8106 3873 8110
rect 3886 8106 3890 8110
rect 3895 8106 3899 8110
rect 3908 8106 3912 8110
rect 3916 8106 3920 8110
rect 3924 8106 3928 8110
rect 3941 8106 3945 8110
rect 3951 8106 3955 8110
rect 3959 8106 3963 8110
rect 4134 8111 4138 8115
rect 4142 8111 4146 8115
rect 2856 8060 2860 8064
rect 2864 8060 2868 8064
rect 2872 8060 2876 8064
rect 2880 8060 2884 8064
rect 2888 8060 2892 8064
rect 2896 8060 2900 8064
rect 2907 8060 2911 8064
rect 2924 8060 2928 8064
rect 2941 8060 2945 8064
rect 2950 8060 2954 8064
rect 2963 8060 2967 8064
rect 2971 8060 2975 8064
rect 2979 8060 2983 8064
rect 2996 8060 3000 8064
rect 3006 8060 3010 8064
rect 3014 8060 3018 8064
rect 3054 8060 3058 8064
rect 3069 8060 3073 8064
rect 3159 8060 3163 8064
rect 3174 8060 3178 8064
rect 3801 8060 3805 8064
rect 3809 8060 3813 8064
rect 3817 8060 3821 8064
rect 3825 8060 3829 8064
rect 3833 8060 3837 8064
rect 3841 8060 3845 8064
rect 3852 8060 3856 8064
rect 3869 8060 3873 8064
rect 3886 8060 3890 8064
rect 3895 8060 3899 8064
rect 3908 8060 3912 8064
rect 3916 8060 3920 8064
rect 3924 8060 3928 8064
rect 3941 8060 3945 8064
rect 3951 8060 3955 8064
rect 3959 8060 3963 8064
rect 3999 8060 4003 8064
rect 4014 8060 4018 8064
rect 4104 8060 4108 8064
rect 4119 8060 4123 8064
rect 3054 7983 3058 7987
rect 3069 7983 3073 7987
rect 3111 7987 3115 7991
rect 3119 7987 3123 7991
rect 3135 7983 3139 7987
rect 3150 7983 3154 7987
rect 3201 7987 3205 7991
rect 3209 7987 3213 7991
rect 3225 7983 3229 7987
rect 3240 7983 3244 7987
rect 3084 7979 3088 7983
rect 3092 7979 3096 7983
rect 2856 7974 2860 7978
rect 2864 7974 2868 7978
rect 2872 7974 2876 7978
rect 2880 7974 2884 7978
rect 2888 7974 2892 7978
rect 2896 7974 2900 7978
rect 2907 7974 2911 7978
rect 2924 7974 2928 7978
rect 2941 7974 2945 7978
rect 2950 7974 2954 7978
rect 2963 7974 2967 7978
rect 2971 7974 2975 7978
rect 2979 7974 2983 7978
rect 2996 7974 3000 7978
rect 3006 7974 3010 7978
rect 3014 7974 3018 7978
rect 3165 7979 3169 7983
rect 3173 7979 3177 7983
rect 3255 7979 3259 7983
rect 3263 7979 3267 7983
rect 3999 7983 4003 7987
rect 4014 7983 4018 7987
rect 4056 7987 4060 7991
rect 4064 7987 4068 7991
rect 4080 7983 4084 7987
rect 4095 7983 4099 7987
rect 4146 7987 4150 7991
rect 4154 7987 4158 7991
rect 4170 7983 4174 7987
rect 4185 7983 4189 7987
rect 4029 7979 4033 7983
rect 4037 7979 4041 7983
rect 3801 7974 3805 7978
rect 3809 7974 3813 7978
rect 3817 7974 3821 7978
rect 3825 7974 3829 7978
rect 3833 7974 3837 7978
rect 3841 7974 3845 7978
rect 3852 7974 3856 7978
rect 3869 7974 3873 7978
rect 3886 7974 3890 7978
rect 3895 7974 3899 7978
rect 3908 7974 3912 7978
rect 3916 7974 3920 7978
rect 3924 7974 3928 7978
rect 3941 7974 3945 7978
rect 3951 7974 3955 7978
rect 3959 7974 3963 7978
rect 4110 7979 4114 7983
rect 4118 7979 4122 7983
rect 4200 7979 4204 7983
rect 4208 7979 4212 7983
rect 2856 7928 2860 7932
rect 2864 7928 2868 7932
rect 2872 7928 2876 7932
rect 2880 7928 2884 7932
rect 2888 7928 2892 7932
rect 2896 7928 2900 7932
rect 2907 7928 2911 7932
rect 2924 7928 2928 7932
rect 2941 7928 2945 7932
rect 2950 7928 2954 7932
rect 2963 7928 2967 7932
rect 2971 7928 2975 7932
rect 2979 7928 2983 7932
rect 2996 7928 3000 7932
rect 3006 7928 3010 7932
rect 3014 7928 3018 7932
rect 3054 7925 3058 7929
rect 3069 7925 3073 7929
rect 3135 7925 3139 7929
rect 3150 7925 3154 7929
rect 3225 7925 3229 7929
rect 3240 7925 3244 7929
rect 3801 7928 3805 7932
rect 3809 7928 3813 7932
rect 3817 7928 3821 7932
rect 3825 7928 3829 7932
rect 3833 7928 3837 7932
rect 3841 7928 3845 7932
rect 3852 7928 3856 7932
rect 3869 7928 3873 7932
rect 3886 7928 3890 7932
rect 3895 7928 3899 7932
rect 3908 7928 3912 7932
rect 3916 7928 3920 7932
rect 3924 7928 3928 7932
rect 3941 7928 3945 7932
rect 3951 7928 3955 7932
rect 3959 7928 3963 7932
rect 3999 7925 4003 7929
rect 4014 7925 4018 7929
rect 4080 7925 4084 7929
rect 4095 7925 4099 7929
rect 4170 7925 4174 7929
rect 4185 7925 4189 7929
rect 3054 7851 3058 7855
rect 3069 7851 3073 7855
rect 3084 7847 3088 7851
rect 3092 7847 3096 7851
rect 2856 7842 2860 7846
rect 2864 7842 2868 7846
rect 2872 7842 2876 7846
rect 2880 7842 2884 7846
rect 2888 7842 2892 7846
rect 2896 7842 2900 7846
rect 2907 7842 2911 7846
rect 2924 7842 2928 7846
rect 2941 7842 2945 7846
rect 2950 7842 2954 7846
rect 2963 7842 2967 7846
rect 2971 7842 2975 7846
rect 2979 7842 2983 7846
rect 2996 7842 3000 7846
rect 3006 7842 3010 7846
rect 3014 7842 3018 7846
rect 3999 7851 4003 7855
rect 4014 7851 4018 7855
rect 4029 7847 4033 7851
rect 4037 7847 4041 7851
rect 3801 7842 3805 7846
rect 3809 7842 3813 7846
rect 3817 7842 3821 7846
rect 3825 7842 3829 7846
rect 3833 7842 3837 7846
rect 3841 7842 3845 7846
rect 3852 7842 3856 7846
rect 3869 7842 3873 7846
rect 3886 7842 3890 7846
rect 3895 7842 3899 7846
rect 3908 7842 3912 7846
rect 3916 7842 3920 7846
rect 3924 7842 3928 7846
rect 3941 7842 3945 7846
rect 3951 7842 3955 7846
rect 3959 7842 3963 7846
rect 2856 7796 2860 7800
rect 2864 7796 2868 7800
rect 2872 7796 2876 7800
rect 2880 7796 2884 7800
rect 2888 7796 2892 7800
rect 2896 7796 2900 7800
rect 2907 7796 2911 7800
rect 2924 7796 2928 7800
rect 2941 7796 2945 7800
rect 2950 7796 2954 7800
rect 2963 7796 2967 7800
rect 2971 7796 2975 7800
rect 2979 7796 2983 7800
rect 2996 7796 3000 7800
rect 3006 7796 3010 7800
rect 3014 7796 3018 7800
rect 3090 7796 3094 7800
rect 3098 7796 3102 7800
rect 3108 7796 3112 7800
rect 3116 7796 3120 7800
rect 3125 7796 3129 7800
rect 3133 7796 3137 7800
rect 3141 7796 3145 7800
rect 3149 7796 3153 7800
rect 3157 7796 3161 7800
rect 3168 7796 3172 7800
rect 3185 7796 3189 7800
rect 3202 7796 3206 7800
rect 3211 7796 3215 7800
rect 3224 7796 3228 7800
rect 3232 7796 3236 7800
rect 3240 7796 3244 7800
rect 3257 7796 3261 7800
rect 3267 7796 3271 7800
rect 3275 7796 3279 7800
rect 2367 7782 2371 7786
rect 2380 7782 2384 7786
rect 2388 7782 2392 7786
rect 2396 7782 2400 7786
rect 2404 7782 2408 7786
rect 2417 7782 2421 7786
rect 2430 7782 2434 7786
rect 2438 7782 2442 7786
rect 2446 7782 2450 7786
rect 2454 7782 2458 7786
rect 2462 7782 2466 7786
rect 2475 7782 2479 7786
rect 2483 7782 2487 7786
rect 2491 7782 2495 7786
rect 2499 7782 2503 7786
rect 2512 7782 2516 7786
rect 2520 7782 2524 7786
rect 2528 7782 2532 7786
rect 2536 7782 2540 7786
rect 2549 7782 2553 7786
rect 2562 7782 2566 7786
rect 2570 7782 2574 7786
rect 2578 7782 2582 7786
rect 2586 7782 2590 7786
rect 2594 7782 2598 7786
rect 2607 7782 2611 7786
rect 2615 7782 2619 7786
rect 2623 7782 2627 7786
rect 2631 7782 2635 7786
rect 2644 7782 2648 7786
rect 2652 7782 2656 7786
rect 2660 7782 2664 7786
rect 2668 7782 2672 7786
rect 2681 7782 2685 7786
rect 2694 7782 2698 7786
rect 2702 7782 2706 7786
rect 2710 7782 2714 7786
rect 2718 7782 2722 7786
rect 2726 7782 2730 7786
rect 2739 7782 2743 7786
rect 2747 7782 2751 7786
rect 2755 7782 2759 7786
rect 3054 7789 3058 7793
rect 3069 7789 3073 7793
rect 3801 7796 3805 7800
rect 3809 7796 3813 7800
rect 3817 7796 3821 7800
rect 3825 7796 3829 7800
rect 3833 7796 3837 7800
rect 3841 7796 3845 7800
rect 3852 7796 3856 7800
rect 3869 7796 3873 7800
rect 3886 7796 3890 7800
rect 3895 7796 3899 7800
rect 3908 7796 3912 7800
rect 3916 7796 3920 7800
rect 3924 7796 3928 7800
rect 3941 7796 3945 7800
rect 3951 7796 3955 7800
rect 3959 7796 3963 7800
rect 4035 7796 4039 7800
rect 4043 7796 4047 7800
rect 4053 7796 4057 7800
rect 4061 7796 4065 7800
rect 4070 7796 4074 7800
rect 4078 7796 4082 7800
rect 4086 7796 4090 7800
rect 4094 7796 4098 7800
rect 4102 7796 4106 7800
rect 4113 7796 4117 7800
rect 4130 7796 4134 7800
rect 4147 7796 4151 7800
rect 4156 7796 4160 7800
rect 4169 7796 4173 7800
rect 4177 7796 4181 7800
rect 4185 7796 4189 7800
rect 4202 7796 4206 7800
rect 4212 7796 4216 7800
rect 4220 7796 4224 7800
rect 3312 7782 3316 7786
rect 3325 7782 3329 7786
rect 3333 7782 3337 7786
rect 3341 7782 3345 7786
rect 3349 7782 3353 7786
rect 3362 7782 3366 7786
rect 3375 7782 3379 7786
rect 3383 7782 3387 7786
rect 3391 7782 3395 7786
rect 3399 7782 3403 7786
rect 3407 7782 3411 7786
rect 3420 7782 3424 7786
rect 3428 7782 3432 7786
rect 3436 7782 3440 7786
rect 3444 7782 3448 7786
rect 3457 7782 3461 7786
rect 3465 7782 3469 7786
rect 3473 7782 3477 7786
rect 3481 7782 3485 7786
rect 3494 7782 3498 7786
rect 3507 7782 3511 7786
rect 3515 7782 3519 7786
rect 3523 7782 3527 7786
rect 3531 7782 3535 7786
rect 3539 7782 3543 7786
rect 3552 7782 3556 7786
rect 3560 7782 3564 7786
rect 3568 7782 3572 7786
rect 3576 7782 3580 7786
rect 3589 7782 3593 7786
rect 3597 7782 3601 7786
rect 3605 7782 3609 7786
rect 3613 7782 3617 7786
rect 3626 7782 3630 7786
rect 3639 7782 3643 7786
rect 3647 7782 3651 7786
rect 3655 7782 3659 7786
rect 3663 7782 3667 7786
rect 3671 7782 3675 7786
rect 3684 7782 3688 7786
rect 3692 7782 3696 7786
rect 3700 7782 3704 7786
rect 3999 7789 4003 7793
rect 4014 7789 4018 7793
rect 2482 7738 2486 7742
rect 2490 7738 2494 7742
rect 2506 7738 2510 7742
rect 2514 7738 2518 7742
rect 3284 7743 3288 7747
rect 3284 7735 3288 7739
rect 3427 7738 3431 7742
rect 3435 7738 3439 7742
rect 3451 7738 3455 7742
rect 3459 7738 3463 7742
rect 4229 7743 4233 7747
rect 4229 7735 4233 7739
rect 2502 7725 2506 7729
rect 2510 7725 2514 7729
rect 3447 7725 3451 7729
rect 3455 7725 3459 7729
rect 2498 7714 2502 7718
rect 3443 7714 3447 7718
rect 2498 7706 2502 7710
rect 2482 7702 2486 7706
rect 2490 7702 2494 7706
rect 2506 7702 2510 7706
rect 2514 7702 2518 7706
rect 3443 7706 3447 7710
rect 3427 7702 3431 7706
rect 3435 7702 3439 7706
rect 3451 7702 3455 7706
rect 3459 7702 3463 7706
rect 3150 7670 3154 7674
rect 3163 7670 3167 7674
rect 3171 7670 3175 7674
rect 3179 7670 3183 7674
rect 3187 7670 3191 7674
rect 3200 7670 3204 7674
rect 3213 7670 3217 7674
rect 3221 7670 3225 7674
rect 3229 7670 3233 7674
rect 3237 7670 3241 7674
rect 3245 7670 3249 7674
rect 3258 7670 3262 7674
rect 3266 7670 3270 7674
rect 3274 7670 3278 7674
rect 4095 7670 4099 7674
rect 4108 7670 4112 7674
rect 4116 7670 4120 7674
rect 4124 7670 4128 7674
rect 4132 7670 4136 7674
rect 4145 7670 4149 7674
rect 4158 7670 4162 7674
rect 4166 7670 4170 7674
rect 4174 7670 4178 7674
rect 4182 7670 4186 7674
rect 4190 7670 4194 7674
rect 4203 7670 4207 7674
rect 4211 7670 4215 7674
rect 4219 7670 4223 7674
rect 2367 7640 2371 7644
rect 2380 7640 2384 7644
rect 2388 7640 2392 7644
rect 2396 7640 2400 7644
rect 2404 7640 2408 7644
rect 2417 7640 2421 7644
rect 2430 7640 2434 7644
rect 2438 7640 2442 7644
rect 2446 7640 2450 7644
rect 2454 7640 2458 7644
rect 2462 7640 2466 7644
rect 2475 7640 2479 7644
rect 2483 7640 2487 7644
rect 2491 7640 2495 7644
rect 2499 7640 2503 7644
rect 2512 7640 2516 7644
rect 2520 7640 2524 7644
rect 2528 7640 2532 7644
rect 2536 7640 2540 7644
rect 2549 7640 2553 7644
rect 2562 7640 2566 7644
rect 2570 7640 2574 7644
rect 2578 7640 2582 7644
rect 2586 7640 2590 7644
rect 2594 7640 2598 7644
rect 2607 7640 2611 7644
rect 2615 7640 2619 7644
rect 2623 7640 2627 7644
rect 2631 7640 2635 7644
rect 2644 7640 2648 7644
rect 2652 7640 2656 7644
rect 2660 7640 2664 7644
rect 2668 7640 2672 7644
rect 2681 7640 2685 7644
rect 2694 7640 2698 7644
rect 2702 7640 2706 7644
rect 2710 7640 2714 7644
rect 2718 7640 2722 7644
rect 2726 7640 2730 7644
rect 2739 7640 2743 7644
rect 2747 7640 2751 7644
rect 2755 7640 2759 7644
rect 3312 7640 3316 7644
rect 3325 7640 3329 7644
rect 3333 7640 3337 7644
rect 3341 7640 3345 7644
rect 3349 7640 3353 7644
rect 3362 7640 3366 7644
rect 3375 7640 3379 7644
rect 3383 7640 3387 7644
rect 3391 7640 3395 7644
rect 3399 7640 3403 7644
rect 3407 7640 3411 7644
rect 3420 7640 3424 7644
rect 3428 7640 3432 7644
rect 3436 7640 3440 7644
rect 3444 7640 3448 7644
rect 3457 7640 3461 7644
rect 3465 7640 3469 7644
rect 3473 7640 3477 7644
rect 3481 7640 3485 7644
rect 3494 7640 3498 7644
rect 3507 7640 3511 7644
rect 3515 7640 3519 7644
rect 3523 7640 3527 7644
rect 3531 7640 3535 7644
rect 3539 7640 3543 7644
rect 3552 7640 3556 7644
rect 3560 7640 3564 7644
rect 3568 7640 3572 7644
rect 3576 7640 3580 7644
rect 3589 7640 3593 7644
rect 3597 7640 3601 7644
rect 3605 7640 3609 7644
rect 3613 7640 3617 7644
rect 3626 7640 3630 7644
rect 3639 7640 3643 7644
rect 3647 7640 3651 7644
rect 3655 7640 3659 7644
rect 3663 7640 3667 7644
rect 3671 7640 3675 7644
rect 3684 7640 3688 7644
rect 3692 7640 3696 7644
rect 3700 7640 3704 7644
rect 3296 7597 3300 7601
rect 3296 7589 3300 7593
rect 4241 7597 4245 7601
rect 4241 7589 4245 7593
rect 3150 7584 3154 7588
rect 3163 7584 3167 7588
rect 3171 7584 3175 7588
rect 3179 7584 3183 7588
rect 3187 7584 3191 7588
rect 3200 7584 3204 7588
rect 3213 7584 3217 7588
rect 3221 7584 3225 7588
rect 3229 7584 3233 7588
rect 3237 7584 3241 7588
rect 3245 7584 3249 7588
rect 3258 7584 3262 7588
rect 3266 7584 3270 7588
rect 3274 7584 3278 7588
rect 4095 7584 4099 7588
rect 4108 7584 4112 7588
rect 4116 7584 4120 7588
rect 4124 7584 4128 7588
rect 4132 7584 4136 7588
rect 4145 7584 4149 7588
rect 4158 7584 4162 7588
rect 4166 7584 4170 7588
rect 4174 7584 4178 7588
rect 4182 7584 4186 7588
rect 4190 7584 4194 7588
rect 4203 7584 4207 7588
rect 4211 7584 4215 7588
rect 4219 7584 4223 7588
rect 2367 7554 2371 7558
rect 2380 7554 2384 7558
rect 2388 7554 2392 7558
rect 2396 7554 2400 7558
rect 2404 7554 2408 7558
rect 2417 7554 2421 7558
rect 2430 7554 2434 7558
rect 2438 7554 2442 7558
rect 2446 7554 2450 7558
rect 2454 7554 2458 7558
rect 2462 7554 2466 7558
rect 2475 7554 2479 7558
rect 2483 7554 2487 7558
rect 2491 7554 2495 7558
rect 2499 7554 2503 7558
rect 2512 7554 2516 7558
rect 2520 7554 2524 7558
rect 2528 7554 2532 7558
rect 2536 7554 2540 7558
rect 2549 7554 2553 7558
rect 2562 7554 2566 7558
rect 2570 7554 2574 7558
rect 2578 7554 2582 7558
rect 2586 7554 2590 7558
rect 2594 7554 2598 7558
rect 2607 7554 2611 7558
rect 2615 7554 2619 7558
rect 2623 7554 2627 7558
rect 2631 7554 2635 7558
rect 2644 7554 2648 7558
rect 2652 7554 2656 7558
rect 2660 7554 2664 7558
rect 2668 7554 2672 7558
rect 2681 7554 2685 7558
rect 2694 7554 2698 7558
rect 2702 7554 2706 7558
rect 2710 7554 2714 7558
rect 2718 7554 2722 7558
rect 2726 7554 2730 7558
rect 2739 7554 2743 7558
rect 2747 7554 2751 7558
rect 2755 7554 2759 7558
rect 3312 7554 3316 7558
rect 3325 7554 3329 7558
rect 3333 7554 3337 7558
rect 3341 7554 3345 7558
rect 3349 7554 3353 7558
rect 3362 7554 3366 7558
rect 3375 7554 3379 7558
rect 3383 7554 3387 7558
rect 3391 7554 3395 7558
rect 3399 7554 3403 7558
rect 3407 7554 3411 7558
rect 3420 7554 3424 7558
rect 3428 7554 3432 7558
rect 3436 7554 3440 7558
rect 3444 7554 3448 7558
rect 3457 7554 3461 7558
rect 3465 7554 3469 7558
rect 3473 7554 3477 7558
rect 3481 7554 3485 7558
rect 3494 7554 3498 7558
rect 3507 7554 3511 7558
rect 3515 7554 3519 7558
rect 3523 7554 3527 7558
rect 3531 7554 3535 7558
rect 3539 7554 3543 7558
rect 3552 7554 3556 7558
rect 3560 7554 3564 7558
rect 3568 7554 3572 7558
rect 3576 7554 3580 7558
rect 3589 7554 3593 7558
rect 3597 7554 3601 7558
rect 3605 7554 3609 7558
rect 3613 7554 3617 7558
rect 3626 7554 3630 7558
rect 3639 7554 3643 7558
rect 3647 7554 3651 7558
rect 3655 7554 3659 7558
rect 3663 7554 3667 7558
rect 3671 7554 3675 7558
rect 3684 7554 3688 7558
rect 3692 7554 3696 7558
rect 3700 7554 3704 7558
rect 2599 7510 2603 7514
rect 2607 7510 2611 7514
rect 2623 7510 2627 7514
rect 2631 7510 2635 7514
rect 3544 7510 3548 7514
rect 3552 7510 3556 7514
rect 3568 7510 3572 7514
rect 3576 7510 3580 7514
rect 2619 7499 2623 7503
rect 2627 7499 2631 7503
rect 3564 7499 3568 7503
rect 3572 7499 3576 7503
rect 2615 7488 2619 7492
rect 3560 7488 3564 7492
rect 2615 7480 2619 7484
rect 3560 7480 3564 7484
rect 2599 7476 2603 7480
rect 2607 7476 2611 7480
rect 2623 7476 2627 7480
rect 2631 7476 2635 7480
rect 3544 7476 3548 7480
rect 3552 7476 3556 7480
rect 3568 7476 3572 7480
rect 3576 7476 3580 7480
rect 2367 7414 2371 7418
rect 2380 7414 2384 7418
rect 2388 7414 2392 7418
rect 2396 7414 2400 7418
rect 2404 7414 2408 7418
rect 2417 7414 2421 7418
rect 2430 7414 2434 7418
rect 2438 7414 2442 7418
rect 2446 7414 2450 7418
rect 2454 7414 2458 7418
rect 2462 7414 2466 7418
rect 2475 7414 2479 7418
rect 2483 7414 2487 7418
rect 2491 7414 2495 7418
rect 2499 7414 2503 7418
rect 2512 7414 2516 7418
rect 2520 7414 2524 7418
rect 2528 7414 2532 7418
rect 2536 7414 2540 7418
rect 2549 7414 2553 7418
rect 2562 7414 2566 7418
rect 2570 7414 2574 7418
rect 2578 7414 2582 7418
rect 2586 7414 2590 7418
rect 2594 7414 2598 7418
rect 2607 7414 2611 7418
rect 2615 7414 2619 7418
rect 2623 7414 2627 7418
rect 2631 7414 2635 7418
rect 2644 7414 2648 7418
rect 2652 7414 2656 7418
rect 2660 7414 2664 7418
rect 2668 7414 2672 7418
rect 2681 7414 2685 7418
rect 2694 7414 2698 7418
rect 2702 7414 2706 7418
rect 2710 7414 2714 7418
rect 2718 7414 2722 7418
rect 2726 7414 2730 7418
rect 2739 7414 2743 7418
rect 2747 7414 2751 7418
rect 2755 7414 2759 7418
rect 3312 7414 3316 7418
rect 3325 7414 3329 7418
rect 3333 7414 3337 7418
rect 3341 7414 3345 7418
rect 3349 7414 3353 7418
rect 3362 7414 3366 7418
rect 3375 7414 3379 7418
rect 3383 7414 3387 7418
rect 3391 7414 3395 7418
rect 3399 7414 3403 7418
rect 3407 7414 3411 7418
rect 3420 7414 3424 7418
rect 3428 7414 3432 7418
rect 3436 7414 3440 7418
rect 3444 7414 3448 7418
rect 3457 7414 3461 7418
rect 3465 7414 3469 7418
rect 3473 7414 3477 7418
rect 3481 7414 3485 7418
rect 3494 7414 3498 7418
rect 3507 7414 3511 7418
rect 3515 7414 3519 7418
rect 3523 7414 3527 7418
rect 3531 7414 3535 7418
rect 3539 7414 3543 7418
rect 3552 7414 3556 7418
rect 3560 7414 3564 7418
rect 3568 7414 3572 7418
rect 3576 7414 3580 7418
rect 3589 7414 3593 7418
rect 3597 7414 3601 7418
rect 3605 7414 3609 7418
rect 3613 7414 3617 7418
rect 3626 7414 3630 7418
rect 3639 7414 3643 7418
rect 3647 7414 3651 7418
rect 3655 7414 3659 7418
rect 3663 7414 3667 7418
rect 3671 7414 3675 7418
rect 3684 7414 3688 7418
rect 3692 7414 3696 7418
rect 3700 7414 3704 7418
rect 4574 7986 4578 8015
rect 4574 7975 4578 7982
rect 4582 7975 4586 8015
rect 4590 7986 4594 8015
rect 4590 7975 4594 7982
rect 4598 7975 4602 8015
rect 4606 7986 4610 8015
rect 4606 7975 4610 7982
rect 4614 7975 4618 8015
rect 4622 7986 4626 8015
rect 4622 7975 4626 7982
rect 4637 7975 4641 8034
rect 4645 7986 4649 8034
rect 4645 7975 4649 7982
rect 4653 7975 4657 8034
rect 4661 7986 4665 8034
rect 4661 7975 4665 7982
rect 4680 7975 4684 8034
rect 4688 7986 4692 8034
rect 4696 7975 4700 8034
rect 4704 7986 4708 8034
rect 4704 7975 4708 7982
rect 4721 7975 4725 8034
rect 4729 7986 4733 8034
rect 4737 7975 4741 8034
rect 4745 7986 4749 8034
rect 4745 7975 4749 7982
<< pdcontact >>
rect 1562 9949 1566 9953
rect 1572 9949 1576 9953
rect 1582 9949 1586 9953
rect 1592 9949 1596 9953
rect 1557 9944 1561 9948
rect 1567 9944 1571 9948
rect 1577 9944 1581 9948
rect 1587 9944 1591 9948
rect 1597 9944 1601 9948
rect 1562 9939 1566 9943
rect 1572 9939 1576 9943
rect 1582 9939 1586 9943
rect 1592 9939 1596 9943
rect 1557 9934 1561 9938
rect 1567 9934 1571 9938
rect 1577 9934 1581 9938
rect 1587 9934 1591 9938
rect 1597 9934 1601 9938
rect 1562 9929 1566 9933
rect 1572 9929 1576 9933
rect 1582 9929 1586 9933
rect 1592 9929 1596 9933
rect 1557 9924 1561 9928
rect 1567 9924 1571 9928
rect 1577 9924 1581 9928
rect 1587 9924 1591 9928
rect 1597 9924 1601 9928
rect 1562 9919 1566 9923
rect 1572 9919 1576 9923
rect 1582 9919 1586 9923
rect 1592 9919 1596 9923
rect 1557 9914 1561 9918
rect 1567 9914 1571 9918
rect 1577 9914 1581 9918
rect 1587 9914 1591 9918
rect 1597 9914 1601 9918
rect 1562 9909 1566 9913
rect 1572 9909 1576 9913
rect 1582 9909 1586 9913
rect 1592 9909 1596 9913
rect 1557 9904 1561 9908
rect 1567 9904 1571 9908
rect 1577 9904 1581 9908
rect 1587 9904 1591 9908
rect 1597 9904 1601 9908
rect 1562 9899 1566 9903
rect 1572 9899 1576 9903
rect 1582 9899 1586 9903
rect 1592 9899 1596 9903
rect 1557 9894 1561 9898
rect 1567 9894 1571 9898
rect 1577 9894 1581 9898
rect 1587 9894 1591 9898
rect 1597 9894 1601 9898
rect 1562 9889 1566 9893
rect 1572 9889 1576 9893
rect 1582 9889 1586 9893
rect 1592 9889 1596 9893
rect 1557 9884 1561 9888
rect 1567 9884 1571 9888
rect 1577 9884 1581 9888
rect 1587 9884 1591 9888
rect 1597 9884 1601 9888
rect 1562 9879 1566 9883
rect 1572 9879 1576 9883
rect 1582 9879 1586 9883
rect 1592 9879 1596 9883
rect 1557 9874 1561 9878
rect 1567 9874 1571 9878
rect 1577 9874 1581 9878
rect 1587 9874 1591 9878
rect 1597 9874 1601 9878
rect 1562 9869 1566 9873
rect 1572 9869 1576 9873
rect 1582 9869 1586 9873
rect 1592 9869 1596 9873
rect 1557 9864 1561 9868
rect 1567 9864 1571 9868
rect 1577 9864 1581 9868
rect 1587 9864 1591 9868
rect 1597 9864 1601 9868
rect 1871 9949 1875 9953
rect 1881 9949 1885 9953
rect 1891 9949 1895 9953
rect 1901 9949 1905 9953
rect 1866 9944 1870 9948
rect 1876 9944 1880 9948
rect 1886 9944 1890 9948
rect 1896 9944 1900 9948
rect 1906 9944 1910 9948
rect 1871 9939 1875 9943
rect 1881 9939 1885 9943
rect 1891 9939 1895 9943
rect 1901 9939 1905 9943
rect 1866 9934 1870 9938
rect 1876 9934 1880 9938
rect 1886 9934 1890 9938
rect 1896 9934 1900 9938
rect 1906 9934 1910 9938
rect 1871 9929 1875 9933
rect 1881 9929 1885 9933
rect 1891 9929 1895 9933
rect 1901 9929 1905 9933
rect 1866 9924 1870 9928
rect 1876 9924 1880 9928
rect 1886 9924 1890 9928
rect 1896 9924 1900 9928
rect 1906 9924 1910 9928
rect 1871 9919 1875 9923
rect 1881 9919 1885 9923
rect 1891 9919 1895 9923
rect 1901 9919 1905 9923
rect 1866 9914 1870 9918
rect 1876 9914 1880 9918
rect 1886 9914 1890 9918
rect 1896 9914 1900 9918
rect 1906 9914 1910 9918
rect 1871 9909 1875 9913
rect 1881 9909 1885 9913
rect 1891 9909 1895 9913
rect 1901 9909 1905 9913
rect 1866 9904 1870 9908
rect 1876 9904 1880 9908
rect 1886 9904 1890 9908
rect 1896 9904 1900 9908
rect 1906 9904 1910 9908
rect 1871 9899 1875 9903
rect 1881 9899 1885 9903
rect 1891 9899 1895 9903
rect 1901 9899 1905 9903
rect 1866 9894 1870 9898
rect 1876 9894 1880 9898
rect 1886 9894 1890 9898
rect 1896 9894 1900 9898
rect 1906 9894 1910 9898
rect 1871 9889 1875 9893
rect 1881 9889 1885 9893
rect 1891 9889 1895 9893
rect 1901 9889 1905 9893
rect 1866 9884 1870 9888
rect 1876 9884 1880 9888
rect 1886 9884 1890 9888
rect 1896 9884 1900 9888
rect 1906 9884 1910 9888
rect 1871 9879 1875 9883
rect 1881 9879 1885 9883
rect 1891 9879 1895 9883
rect 1901 9879 1905 9883
rect 1866 9874 1870 9878
rect 1876 9874 1880 9878
rect 1886 9874 1890 9878
rect 1896 9874 1900 9878
rect 1906 9874 1910 9878
rect 1871 9869 1875 9873
rect 1881 9869 1885 9873
rect 1891 9869 1895 9873
rect 1901 9869 1905 9873
rect 1866 9864 1870 9868
rect 1876 9864 1880 9868
rect 1886 9864 1890 9868
rect 1896 9864 1900 9868
rect 1906 9864 1910 9868
rect 2180 9949 2184 9953
rect 2190 9949 2194 9953
rect 2200 9949 2204 9953
rect 2210 9949 2214 9953
rect 2175 9944 2179 9948
rect 2185 9944 2189 9948
rect 2195 9944 2199 9948
rect 2205 9944 2209 9948
rect 2215 9944 2219 9948
rect 2180 9939 2184 9943
rect 2190 9939 2194 9943
rect 2200 9939 2204 9943
rect 2210 9939 2214 9943
rect 2175 9934 2179 9938
rect 2185 9934 2189 9938
rect 2195 9934 2199 9938
rect 2205 9934 2209 9938
rect 2215 9934 2219 9938
rect 2180 9929 2184 9933
rect 2190 9929 2194 9933
rect 2200 9929 2204 9933
rect 2210 9929 2214 9933
rect 2175 9924 2179 9928
rect 2185 9924 2189 9928
rect 2195 9924 2199 9928
rect 2205 9924 2209 9928
rect 2215 9924 2219 9928
rect 2180 9919 2184 9923
rect 2190 9919 2194 9923
rect 2200 9919 2204 9923
rect 2210 9919 2214 9923
rect 2175 9914 2179 9918
rect 2185 9914 2189 9918
rect 2195 9914 2199 9918
rect 2205 9914 2209 9918
rect 2215 9914 2219 9918
rect 2180 9909 2184 9913
rect 2190 9909 2194 9913
rect 2200 9909 2204 9913
rect 2210 9909 2214 9913
rect 2175 9904 2179 9908
rect 2185 9904 2189 9908
rect 2195 9904 2199 9908
rect 2205 9904 2209 9908
rect 2215 9904 2219 9908
rect 2180 9899 2184 9903
rect 2190 9899 2194 9903
rect 2200 9899 2204 9903
rect 2210 9899 2214 9903
rect 2175 9894 2179 9898
rect 2185 9894 2189 9898
rect 2195 9894 2199 9898
rect 2205 9894 2209 9898
rect 2215 9894 2219 9898
rect 2180 9889 2184 9893
rect 2190 9889 2194 9893
rect 2200 9889 2204 9893
rect 2210 9889 2214 9893
rect 2175 9884 2179 9888
rect 2185 9884 2189 9888
rect 2195 9884 2199 9888
rect 2205 9884 2209 9888
rect 2215 9884 2219 9888
rect 2180 9879 2184 9883
rect 2190 9879 2194 9883
rect 2200 9879 2204 9883
rect 2210 9879 2214 9883
rect 2175 9874 2179 9878
rect 2185 9874 2189 9878
rect 2195 9874 2199 9878
rect 2205 9874 2209 9878
rect 2215 9874 2219 9878
rect 2180 9869 2184 9873
rect 2190 9869 2194 9873
rect 2200 9869 2204 9873
rect 2210 9869 2214 9873
rect 2175 9864 2179 9868
rect 2185 9864 2189 9868
rect 2195 9864 2199 9868
rect 2205 9864 2209 9868
rect 2215 9864 2219 9868
rect 2489 9949 2493 9953
rect 2499 9949 2503 9953
rect 2509 9949 2513 9953
rect 2519 9949 2523 9953
rect 2484 9944 2488 9948
rect 2494 9944 2498 9948
rect 2504 9944 2508 9948
rect 2514 9944 2518 9948
rect 2524 9944 2528 9948
rect 2489 9939 2493 9943
rect 2499 9939 2503 9943
rect 2509 9939 2513 9943
rect 2519 9939 2523 9943
rect 2484 9934 2488 9938
rect 2494 9934 2498 9938
rect 2504 9934 2508 9938
rect 2514 9934 2518 9938
rect 2524 9934 2528 9938
rect 2489 9929 2493 9933
rect 2499 9929 2503 9933
rect 2509 9929 2513 9933
rect 2519 9929 2523 9933
rect 2484 9924 2488 9928
rect 2494 9924 2498 9928
rect 2504 9924 2508 9928
rect 2514 9924 2518 9928
rect 2524 9924 2528 9928
rect 2489 9919 2493 9923
rect 2499 9919 2503 9923
rect 2509 9919 2513 9923
rect 2519 9919 2523 9923
rect 2484 9914 2488 9918
rect 2494 9914 2498 9918
rect 2504 9914 2508 9918
rect 2514 9914 2518 9918
rect 2524 9914 2528 9918
rect 2489 9909 2493 9913
rect 2499 9909 2503 9913
rect 2509 9909 2513 9913
rect 2519 9909 2523 9913
rect 2484 9904 2488 9908
rect 2494 9904 2498 9908
rect 2504 9904 2508 9908
rect 2514 9904 2518 9908
rect 2524 9904 2528 9908
rect 2489 9899 2493 9903
rect 2499 9899 2503 9903
rect 2509 9899 2513 9903
rect 2519 9899 2523 9903
rect 2484 9894 2488 9898
rect 2494 9894 2498 9898
rect 2504 9894 2508 9898
rect 2514 9894 2518 9898
rect 2524 9894 2528 9898
rect 2489 9889 2493 9893
rect 2499 9889 2503 9893
rect 2509 9889 2513 9893
rect 2519 9889 2523 9893
rect 2484 9884 2488 9888
rect 2494 9884 2498 9888
rect 2504 9884 2508 9888
rect 2514 9884 2518 9888
rect 2524 9884 2528 9888
rect 2489 9879 2493 9883
rect 2499 9879 2503 9883
rect 2509 9879 2513 9883
rect 2519 9879 2523 9883
rect 2484 9874 2488 9878
rect 2494 9874 2498 9878
rect 2504 9874 2508 9878
rect 2514 9874 2518 9878
rect 2524 9874 2528 9878
rect 2489 9869 2493 9873
rect 2499 9869 2503 9873
rect 2509 9869 2513 9873
rect 2519 9869 2523 9873
rect 2484 9864 2488 9868
rect 2494 9864 2498 9868
rect 2504 9864 2508 9868
rect 2514 9864 2518 9868
rect 2524 9864 2528 9868
rect 2798 9949 2802 9953
rect 2808 9949 2812 9953
rect 2818 9949 2822 9953
rect 2828 9949 2832 9953
rect 2793 9944 2797 9948
rect 2803 9944 2807 9948
rect 2813 9944 2817 9948
rect 2823 9944 2827 9948
rect 2833 9944 2837 9948
rect 2798 9939 2802 9943
rect 2808 9939 2812 9943
rect 2818 9939 2822 9943
rect 2828 9939 2832 9943
rect 2793 9934 2797 9938
rect 2803 9934 2807 9938
rect 2813 9934 2817 9938
rect 2823 9934 2827 9938
rect 2833 9934 2837 9938
rect 2798 9929 2802 9933
rect 2808 9929 2812 9933
rect 2818 9929 2822 9933
rect 2828 9929 2832 9933
rect 2793 9924 2797 9928
rect 2803 9924 2807 9928
rect 2813 9924 2817 9928
rect 2823 9924 2827 9928
rect 2833 9924 2837 9928
rect 2798 9919 2802 9923
rect 2808 9919 2812 9923
rect 2818 9919 2822 9923
rect 2828 9919 2832 9923
rect 2793 9914 2797 9918
rect 2803 9914 2807 9918
rect 2813 9914 2817 9918
rect 2823 9914 2827 9918
rect 2833 9914 2837 9918
rect 2798 9909 2802 9913
rect 2808 9909 2812 9913
rect 2818 9909 2822 9913
rect 2828 9909 2832 9913
rect 2793 9904 2797 9908
rect 2803 9904 2807 9908
rect 2813 9904 2817 9908
rect 2823 9904 2827 9908
rect 2833 9904 2837 9908
rect 2798 9899 2802 9903
rect 2808 9899 2812 9903
rect 2818 9899 2822 9903
rect 2828 9899 2832 9903
rect 2793 9894 2797 9898
rect 2803 9894 2807 9898
rect 2813 9894 2817 9898
rect 2823 9894 2827 9898
rect 2833 9894 2837 9898
rect 2798 9889 2802 9893
rect 2808 9889 2812 9893
rect 2818 9889 2822 9893
rect 2828 9889 2832 9893
rect 2793 9884 2797 9888
rect 2803 9884 2807 9888
rect 2813 9884 2817 9888
rect 2823 9884 2827 9888
rect 2833 9884 2837 9888
rect 2798 9879 2802 9883
rect 2808 9879 2812 9883
rect 2818 9879 2822 9883
rect 2828 9879 2832 9883
rect 2793 9874 2797 9878
rect 2803 9874 2807 9878
rect 2813 9874 2817 9878
rect 2823 9874 2827 9878
rect 2833 9874 2837 9878
rect 2798 9869 2802 9873
rect 2808 9869 2812 9873
rect 2818 9869 2822 9873
rect 2828 9869 2832 9873
rect 2793 9864 2797 9868
rect 2803 9864 2807 9868
rect 2813 9864 2817 9868
rect 2823 9864 2827 9868
rect 2833 9864 2837 9868
rect 3107 9949 3111 9953
rect 3117 9949 3121 9953
rect 3127 9949 3131 9953
rect 3137 9949 3141 9953
rect 3102 9944 3106 9948
rect 3112 9944 3116 9948
rect 3122 9944 3126 9948
rect 3132 9944 3136 9948
rect 3142 9944 3146 9948
rect 3107 9939 3111 9943
rect 3117 9939 3121 9943
rect 3127 9939 3131 9943
rect 3137 9939 3141 9943
rect 3102 9934 3106 9938
rect 3112 9934 3116 9938
rect 3122 9934 3126 9938
rect 3132 9934 3136 9938
rect 3142 9934 3146 9938
rect 3107 9929 3111 9933
rect 3117 9929 3121 9933
rect 3127 9929 3131 9933
rect 3137 9929 3141 9933
rect 3102 9924 3106 9928
rect 3112 9924 3116 9928
rect 3122 9924 3126 9928
rect 3132 9924 3136 9928
rect 3142 9924 3146 9928
rect 3107 9919 3111 9923
rect 3117 9919 3121 9923
rect 3127 9919 3131 9923
rect 3137 9919 3141 9923
rect 3102 9914 3106 9918
rect 3112 9914 3116 9918
rect 3122 9914 3126 9918
rect 3132 9914 3136 9918
rect 3142 9914 3146 9918
rect 3107 9909 3111 9913
rect 3117 9909 3121 9913
rect 3127 9909 3131 9913
rect 3137 9909 3141 9913
rect 3102 9904 3106 9908
rect 3112 9904 3116 9908
rect 3122 9904 3126 9908
rect 3132 9904 3136 9908
rect 3142 9904 3146 9908
rect 3107 9899 3111 9903
rect 3117 9899 3121 9903
rect 3127 9899 3131 9903
rect 3137 9899 3141 9903
rect 3102 9894 3106 9898
rect 3112 9894 3116 9898
rect 3122 9894 3126 9898
rect 3132 9894 3136 9898
rect 3142 9894 3146 9898
rect 3107 9889 3111 9893
rect 3117 9889 3121 9893
rect 3127 9889 3131 9893
rect 3137 9889 3141 9893
rect 3102 9884 3106 9888
rect 3112 9884 3116 9888
rect 3122 9884 3126 9888
rect 3132 9884 3136 9888
rect 3142 9884 3146 9888
rect 3107 9879 3111 9883
rect 3117 9879 3121 9883
rect 3127 9879 3131 9883
rect 3137 9879 3141 9883
rect 3102 9874 3106 9878
rect 3112 9874 3116 9878
rect 3122 9874 3126 9878
rect 3132 9874 3136 9878
rect 3142 9874 3146 9878
rect 3107 9869 3111 9873
rect 3117 9869 3121 9873
rect 3127 9869 3131 9873
rect 3137 9869 3141 9873
rect 3102 9864 3106 9868
rect 3112 9864 3116 9868
rect 3122 9864 3126 9868
rect 3132 9864 3136 9868
rect 3142 9864 3146 9868
rect 3416 9949 3420 9953
rect 3426 9949 3430 9953
rect 3436 9949 3440 9953
rect 3446 9949 3450 9953
rect 3411 9944 3415 9948
rect 3421 9944 3425 9948
rect 3431 9944 3435 9948
rect 3441 9944 3445 9948
rect 3451 9944 3455 9948
rect 3416 9939 3420 9943
rect 3426 9939 3430 9943
rect 3436 9939 3440 9943
rect 3446 9939 3450 9943
rect 3411 9934 3415 9938
rect 3421 9934 3425 9938
rect 3431 9934 3435 9938
rect 3441 9934 3445 9938
rect 3451 9934 3455 9938
rect 3416 9929 3420 9933
rect 3426 9929 3430 9933
rect 3436 9929 3440 9933
rect 3446 9929 3450 9933
rect 3411 9924 3415 9928
rect 3421 9924 3425 9928
rect 3431 9924 3435 9928
rect 3441 9924 3445 9928
rect 3451 9924 3455 9928
rect 3416 9919 3420 9923
rect 3426 9919 3430 9923
rect 3436 9919 3440 9923
rect 3446 9919 3450 9923
rect 3411 9914 3415 9918
rect 3421 9914 3425 9918
rect 3431 9914 3435 9918
rect 3441 9914 3445 9918
rect 3451 9914 3455 9918
rect 3416 9909 3420 9913
rect 3426 9909 3430 9913
rect 3436 9909 3440 9913
rect 3446 9909 3450 9913
rect 3411 9904 3415 9908
rect 3421 9904 3425 9908
rect 3431 9904 3435 9908
rect 3441 9904 3445 9908
rect 3451 9904 3455 9908
rect 3416 9899 3420 9903
rect 3426 9899 3430 9903
rect 3436 9899 3440 9903
rect 3446 9899 3450 9903
rect 3411 9894 3415 9898
rect 3421 9894 3425 9898
rect 3431 9894 3435 9898
rect 3441 9894 3445 9898
rect 3451 9894 3455 9898
rect 3416 9889 3420 9893
rect 3426 9889 3430 9893
rect 3436 9889 3440 9893
rect 3446 9889 3450 9893
rect 3411 9884 3415 9888
rect 3421 9884 3425 9888
rect 3431 9884 3435 9888
rect 3441 9884 3445 9888
rect 3451 9884 3455 9888
rect 3416 9879 3420 9883
rect 3426 9879 3430 9883
rect 3436 9879 3440 9883
rect 3446 9879 3450 9883
rect 3411 9874 3415 9878
rect 3421 9874 3425 9878
rect 3431 9874 3435 9878
rect 3441 9874 3445 9878
rect 3451 9874 3455 9878
rect 3416 9869 3420 9873
rect 3426 9869 3430 9873
rect 3436 9869 3440 9873
rect 3446 9869 3450 9873
rect 3411 9864 3415 9868
rect 3421 9864 3425 9868
rect 3431 9864 3435 9868
rect 3441 9864 3445 9868
rect 3451 9864 3455 9868
rect 3725 9949 3729 9953
rect 3735 9949 3739 9953
rect 3745 9949 3749 9953
rect 3755 9949 3759 9953
rect 3720 9944 3724 9948
rect 3730 9944 3734 9948
rect 3740 9944 3744 9948
rect 3750 9944 3754 9948
rect 3760 9944 3764 9948
rect 3725 9939 3729 9943
rect 3735 9939 3739 9943
rect 3745 9939 3749 9943
rect 3755 9939 3759 9943
rect 3720 9934 3724 9938
rect 3730 9934 3734 9938
rect 3740 9934 3744 9938
rect 3750 9934 3754 9938
rect 3760 9934 3764 9938
rect 3725 9929 3729 9933
rect 3735 9929 3739 9933
rect 3745 9929 3749 9933
rect 3755 9929 3759 9933
rect 3720 9924 3724 9928
rect 3730 9924 3734 9928
rect 3740 9924 3744 9928
rect 3750 9924 3754 9928
rect 3760 9924 3764 9928
rect 3725 9919 3729 9923
rect 3735 9919 3739 9923
rect 3745 9919 3749 9923
rect 3755 9919 3759 9923
rect 3720 9914 3724 9918
rect 3730 9914 3734 9918
rect 3740 9914 3744 9918
rect 3750 9914 3754 9918
rect 3760 9914 3764 9918
rect 3725 9909 3729 9913
rect 3735 9909 3739 9913
rect 3745 9909 3749 9913
rect 3755 9909 3759 9913
rect 3720 9904 3724 9908
rect 3730 9904 3734 9908
rect 3740 9904 3744 9908
rect 3750 9904 3754 9908
rect 3760 9904 3764 9908
rect 3725 9899 3729 9903
rect 3735 9899 3739 9903
rect 3745 9899 3749 9903
rect 3755 9899 3759 9903
rect 3720 9894 3724 9898
rect 3730 9894 3734 9898
rect 3740 9894 3744 9898
rect 3750 9894 3754 9898
rect 3760 9894 3764 9898
rect 3725 9889 3729 9893
rect 3735 9889 3739 9893
rect 3745 9889 3749 9893
rect 3755 9889 3759 9893
rect 3720 9884 3724 9888
rect 3730 9884 3734 9888
rect 3740 9884 3744 9888
rect 3750 9884 3754 9888
rect 3760 9884 3764 9888
rect 3725 9879 3729 9883
rect 3735 9879 3739 9883
rect 3745 9879 3749 9883
rect 3755 9879 3759 9883
rect 3720 9874 3724 9878
rect 3730 9874 3734 9878
rect 3740 9874 3744 9878
rect 3750 9874 3754 9878
rect 3760 9874 3764 9878
rect 3725 9869 3729 9873
rect 3735 9869 3739 9873
rect 3745 9869 3749 9873
rect 3755 9869 3759 9873
rect 3720 9864 3724 9868
rect 3730 9864 3734 9868
rect 3740 9864 3744 9868
rect 3750 9864 3754 9868
rect 3760 9864 3764 9868
rect 4034 9949 4038 9953
rect 4044 9949 4048 9953
rect 4054 9949 4058 9953
rect 4064 9949 4068 9953
rect 4029 9944 4033 9948
rect 4039 9944 4043 9948
rect 4049 9944 4053 9948
rect 4059 9944 4063 9948
rect 4069 9944 4073 9948
rect 4034 9939 4038 9943
rect 4044 9939 4048 9943
rect 4054 9939 4058 9943
rect 4064 9939 4068 9943
rect 4029 9934 4033 9938
rect 4039 9934 4043 9938
rect 4049 9934 4053 9938
rect 4059 9934 4063 9938
rect 4069 9934 4073 9938
rect 4034 9929 4038 9933
rect 4044 9929 4048 9933
rect 4054 9929 4058 9933
rect 4064 9929 4068 9933
rect 4029 9924 4033 9928
rect 4039 9924 4043 9928
rect 4049 9924 4053 9928
rect 4059 9924 4063 9928
rect 4069 9924 4073 9928
rect 4034 9919 4038 9923
rect 4044 9919 4048 9923
rect 4054 9919 4058 9923
rect 4064 9919 4068 9923
rect 4029 9914 4033 9918
rect 4039 9914 4043 9918
rect 4049 9914 4053 9918
rect 4059 9914 4063 9918
rect 4069 9914 4073 9918
rect 4034 9909 4038 9913
rect 4044 9909 4048 9913
rect 4054 9909 4058 9913
rect 4064 9909 4068 9913
rect 4029 9904 4033 9908
rect 4039 9904 4043 9908
rect 4049 9904 4053 9908
rect 4059 9904 4063 9908
rect 4069 9904 4073 9908
rect 4034 9899 4038 9903
rect 4044 9899 4048 9903
rect 4054 9899 4058 9903
rect 4064 9899 4068 9903
rect 4029 9894 4033 9898
rect 4039 9894 4043 9898
rect 4049 9894 4053 9898
rect 4059 9894 4063 9898
rect 4069 9894 4073 9898
rect 4034 9889 4038 9893
rect 4044 9889 4048 9893
rect 4054 9889 4058 9893
rect 4064 9889 4068 9893
rect 4029 9884 4033 9888
rect 4039 9884 4043 9888
rect 4049 9884 4053 9888
rect 4059 9884 4063 9888
rect 4069 9884 4073 9888
rect 4034 9879 4038 9883
rect 4044 9879 4048 9883
rect 4054 9879 4058 9883
rect 4064 9879 4068 9883
rect 4029 9874 4033 9878
rect 4039 9874 4043 9878
rect 4049 9874 4053 9878
rect 4059 9874 4063 9878
rect 4069 9874 4073 9878
rect 4034 9869 4038 9873
rect 4044 9869 4048 9873
rect 4054 9869 4058 9873
rect 4064 9869 4068 9873
rect 4029 9864 4033 9868
rect 4039 9864 4043 9868
rect 4049 9864 4053 9868
rect 4059 9864 4063 9868
rect 4069 9864 4073 9868
rect 1743 9827 1778 9831
rect 1782 9827 1799 9831
rect 2052 9827 2087 9831
rect 2091 9827 2108 9831
rect 2361 9827 2396 9831
rect 2400 9827 2417 9831
rect 2670 9827 2705 9831
rect 2709 9827 2726 9831
rect 2979 9827 3014 9831
rect 3018 9827 3035 9831
rect 3906 9827 3941 9831
rect 3945 9827 3962 9831
rect 1743 9819 1799 9823
rect 2052 9819 2108 9823
rect 2361 9819 2417 9823
rect 2670 9819 2726 9823
rect 2979 9819 3035 9823
rect 3906 9819 3962 9823
rect 1743 9811 1778 9815
rect 1782 9811 1799 9815
rect 2052 9811 2087 9815
rect 2091 9811 2108 9815
rect 1743 9803 1799 9807
rect 1743 9795 1778 9799
rect 1782 9795 1799 9799
rect 1743 9787 1799 9791
rect 2361 9811 2396 9815
rect 2400 9811 2417 9815
rect 2052 9803 2108 9807
rect 2052 9795 2087 9799
rect 2091 9795 2108 9799
rect 2052 9787 2108 9791
rect 2670 9811 2705 9815
rect 2709 9811 2726 9815
rect 2361 9803 2417 9807
rect 2361 9795 2396 9799
rect 2400 9795 2417 9799
rect 2361 9787 2417 9791
rect 2979 9811 3014 9815
rect 3018 9811 3035 9815
rect 2670 9803 2726 9807
rect 2670 9795 2705 9799
rect 2709 9795 2726 9799
rect 2670 9787 2726 9791
rect 3906 9811 3941 9815
rect 3945 9811 3962 9815
rect 2979 9803 3035 9807
rect 2979 9795 3014 9799
rect 3018 9795 3035 9799
rect 2979 9787 3035 9791
rect 3906 9803 3962 9807
rect 3906 9795 3941 9799
rect 3945 9795 3962 9799
rect 3906 9787 3962 9791
rect 1743 9779 1778 9783
rect 1782 9779 1799 9783
rect 2052 9779 2087 9783
rect 2091 9779 2108 9783
rect 2361 9779 2396 9783
rect 2400 9779 2417 9783
rect 2670 9779 2705 9783
rect 2709 9779 2726 9783
rect 2979 9779 3014 9783
rect 3018 9779 3035 9783
rect 3906 9779 3941 9783
rect 3945 9779 3962 9783
rect 2851 9322 2855 9330
rect 2864 9322 2868 9330
rect 2872 9322 2876 9330
rect 2880 9326 2884 9330
rect 2888 9322 2892 9330
rect 2901 9322 2905 9330
rect 2914 9322 2918 9330
rect 2922 9322 2926 9330
rect 2930 9322 2934 9330
rect 2938 9326 2942 9330
rect 2946 9322 2950 9330
rect 2959 9322 2963 9330
rect 2967 9322 2971 9330
rect 2975 9322 2979 9330
rect 2983 9322 2987 9330
rect 2996 9322 3000 9330
rect 3004 9322 3008 9330
rect 3012 9326 3016 9330
rect 3020 9322 3024 9330
rect 3033 9322 3037 9330
rect 3046 9322 3050 9330
rect 3054 9322 3058 9330
rect 3062 9322 3066 9330
rect 3070 9326 3074 9330
rect 3078 9322 3082 9330
rect 3091 9322 3095 9330
rect 3099 9322 3103 9330
rect 3107 9322 3111 9330
rect 3115 9322 3119 9330
rect 3128 9322 3132 9330
rect 3136 9322 3140 9330
rect 3144 9326 3148 9330
rect 3152 9322 3156 9330
rect 3165 9322 3169 9330
rect 3178 9322 3182 9330
rect 3186 9322 3190 9330
rect 3194 9322 3198 9330
rect 3202 9326 3206 9330
rect 3210 9322 3214 9330
rect 3223 9322 3227 9330
rect 3231 9322 3235 9330
rect 3239 9322 3243 9330
rect 3247 9322 3251 9330
rect 3260 9322 3264 9330
rect 3268 9322 3272 9330
rect 3276 9326 3280 9330
rect 3284 9322 3288 9330
rect 3297 9322 3301 9330
rect 3310 9322 3314 9330
rect 3318 9322 3322 9330
rect 3326 9322 3330 9330
rect 3334 9326 3338 9330
rect 3342 9322 3346 9330
rect 3355 9322 3359 9330
rect 3363 9322 3367 9330
rect 3371 9322 3375 9330
rect 3796 9322 3800 9330
rect 3809 9322 3813 9330
rect 3817 9322 3821 9330
rect 3825 9326 3829 9330
rect 3833 9322 3837 9330
rect 3846 9322 3850 9330
rect 3859 9322 3863 9330
rect 3867 9322 3871 9330
rect 3875 9322 3879 9330
rect 3883 9326 3887 9330
rect 3891 9322 3895 9330
rect 3904 9322 3908 9330
rect 3912 9322 3916 9330
rect 3920 9322 3924 9330
rect 3928 9322 3932 9330
rect 3941 9322 3945 9330
rect 3949 9322 3953 9330
rect 3957 9326 3961 9330
rect 3965 9322 3969 9330
rect 3978 9322 3982 9330
rect 3991 9322 3995 9330
rect 3999 9322 4003 9330
rect 4007 9322 4011 9330
rect 4015 9326 4019 9330
rect 4023 9322 4027 9330
rect 4036 9322 4040 9330
rect 4044 9322 4048 9330
rect 4052 9322 4056 9330
rect 4060 9322 4064 9330
rect 4073 9322 4077 9330
rect 4081 9322 4085 9330
rect 4089 9326 4093 9330
rect 4097 9322 4101 9330
rect 4110 9322 4114 9330
rect 4123 9322 4127 9330
rect 4131 9322 4135 9330
rect 4139 9322 4143 9330
rect 4147 9326 4151 9330
rect 4155 9322 4159 9330
rect 4168 9322 4172 9330
rect 4176 9322 4180 9330
rect 4184 9322 4188 9330
rect 4192 9322 4196 9330
rect 4205 9322 4209 9330
rect 4213 9322 4217 9330
rect 4221 9326 4225 9330
rect 4229 9322 4233 9330
rect 4242 9322 4246 9330
rect 4255 9322 4259 9330
rect 4263 9322 4267 9330
rect 4271 9322 4275 9330
rect 4279 9326 4283 9330
rect 4287 9322 4291 9330
rect 4300 9322 4304 9330
rect 4308 9322 4312 9330
rect 4316 9322 4320 9330
rect 2499 9289 2503 9297
rect 2512 9289 2516 9297
rect 2520 9289 2524 9297
rect 2528 9293 2532 9297
rect 2536 9289 2540 9297
rect 2549 9289 2553 9297
rect 2562 9289 2566 9297
rect 2570 9289 2574 9297
rect 2578 9289 2582 9297
rect 2586 9293 2590 9297
rect 2594 9289 2598 9297
rect 2607 9289 2611 9297
rect 2615 9289 2619 9297
rect 2623 9289 2627 9297
rect 3444 9289 3448 9297
rect 3457 9289 3461 9297
rect 3465 9289 3469 9297
rect 3473 9293 3477 9297
rect 3481 9289 3485 9297
rect 3494 9289 3498 9297
rect 3507 9289 3511 9297
rect 3515 9289 3519 9297
rect 3523 9289 3527 9297
rect 3531 9293 3535 9297
rect 3539 9289 3543 9297
rect 3552 9289 3556 9297
rect 3560 9289 3564 9297
rect 3568 9289 3572 9297
rect 3030 9251 3034 9259
rect 3038 9251 3042 9259
rect 2856 9238 2860 9246
rect 2864 9238 2868 9246
rect 2872 9238 2876 9246
rect 2880 9238 2884 9246
rect 2888 9238 2892 9246
rect 2896 9238 2900 9246
rect 2907 9238 2911 9246
rect 2924 9238 2928 9246
rect 2941 9238 2945 9246
rect 2950 9238 2954 9246
rect 2963 9238 2967 9246
rect 2971 9238 2975 9246
rect 2979 9238 2983 9246
rect 2996 9238 3000 9246
rect 3006 9238 3010 9246
rect 3014 9238 3018 9246
rect 3054 9245 3058 9253
rect 3069 9245 3073 9253
rect 3084 9251 3088 9259
rect 3092 9251 3096 9259
rect 3111 9251 3115 9259
rect 3119 9251 3123 9259
rect 3135 9245 3139 9253
rect 3150 9245 3154 9253
rect 3165 9251 3169 9259
rect 3173 9251 3177 9259
rect 3975 9251 3979 9259
rect 3983 9251 3987 9259
rect 3801 9238 3805 9246
rect 3809 9238 3813 9246
rect 3817 9238 3821 9246
rect 3825 9238 3829 9246
rect 3833 9238 3837 9246
rect 3841 9238 3845 9246
rect 3852 9238 3856 9246
rect 3869 9238 3873 9246
rect 3886 9238 3890 9246
rect 3895 9238 3899 9246
rect 3908 9238 3912 9246
rect 3916 9238 3920 9246
rect 3924 9238 3928 9246
rect 3941 9238 3945 9246
rect 3951 9238 3955 9246
rect 3959 9238 3963 9246
rect 3999 9245 4003 9253
rect 4014 9245 4018 9253
rect 4029 9251 4033 9259
rect 4037 9251 4041 9259
rect 4056 9251 4060 9259
rect 4064 9251 4068 9259
rect 4080 9245 4084 9253
rect 4095 9245 4099 9253
rect 4110 9251 4114 9259
rect 4118 9251 4122 9259
rect 2490 9187 2494 9195
rect 2498 9187 2502 9195
rect 2506 9187 2510 9195
rect 2519 9187 2523 9195
rect 2527 9191 2531 9195
rect 2535 9187 2539 9195
rect 2543 9187 2547 9195
rect 2551 9187 2555 9195
rect 2564 9187 2568 9195
rect 2577 9187 2581 9195
rect 2585 9191 2589 9195
rect 2593 9187 2597 9195
rect 2601 9187 2605 9195
rect 2614 9187 2618 9195
rect 3435 9187 3439 9195
rect 3443 9187 3447 9195
rect 3451 9187 3455 9195
rect 3464 9187 3468 9195
rect 3472 9191 3476 9195
rect 3480 9187 3484 9195
rect 3488 9187 3492 9195
rect 3496 9187 3500 9195
rect 3509 9187 3513 9195
rect 3522 9187 3526 9195
rect 3530 9191 3534 9195
rect 3538 9187 3542 9195
rect 3546 9187 3550 9195
rect 3559 9187 3563 9195
rect 2856 9152 2860 9160
rect 2864 9152 2868 9160
rect 2872 9152 2876 9160
rect 2880 9152 2884 9160
rect 2888 9152 2892 9160
rect 2896 9152 2900 9160
rect 2907 9152 2911 9160
rect 2924 9152 2928 9160
rect 2941 9152 2945 9160
rect 2950 9152 2954 9160
rect 2963 9152 2967 9160
rect 2971 9152 2975 9160
rect 2979 9152 2983 9160
rect 2996 9152 3000 9160
rect 3006 9152 3010 9160
rect 3014 9152 3018 9160
rect 3054 9153 3058 9161
rect 3069 9153 3073 9161
rect 3135 9153 3139 9161
rect 3150 9153 3154 9161
rect 3801 9152 3805 9160
rect 3809 9152 3813 9160
rect 3817 9152 3821 9160
rect 3825 9152 3829 9160
rect 3833 9152 3837 9160
rect 3841 9152 3845 9160
rect 3852 9152 3856 9160
rect 3869 9152 3873 9160
rect 3886 9152 3890 9160
rect 3895 9152 3899 9160
rect 3908 9152 3912 9160
rect 3916 9152 3920 9160
rect 3924 9152 3928 9160
rect 3941 9152 3945 9160
rect 3951 9152 3955 9160
rect 3959 9152 3963 9160
rect 3999 9153 4003 9161
rect 4014 9153 4018 9161
rect 4080 9153 4084 9161
rect 4095 9153 4099 9161
rect 2856 9106 2860 9114
rect 2864 9106 2868 9114
rect 2872 9106 2876 9114
rect 2880 9106 2884 9114
rect 2888 9106 2892 9114
rect 2896 9106 2900 9114
rect 2907 9106 2911 9114
rect 2924 9106 2928 9114
rect 2941 9106 2945 9114
rect 2950 9106 2954 9114
rect 2963 9106 2967 9114
rect 2971 9106 2975 9114
rect 2979 9106 2983 9114
rect 2996 9106 3000 9114
rect 3006 9106 3010 9114
rect 3014 9106 3018 9114
rect 3054 9113 3058 9121
rect 3069 9113 3073 9121
rect 3084 9119 3088 9127
rect 3092 9119 3096 9127
rect 3135 9119 3139 9127
rect 3143 9119 3147 9127
rect 3159 9113 3163 9121
rect 3174 9113 3178 9121
rect 3189 9119 3193 9127
rect 3197 9119 3201 9127
rect 3801 9106 3805 9114
rect 3809 9106 3813 9114
rect 3817 9106 3821 9114
rect 3825 9106 3829 9114
rect 3833 9106 3837 9114
rect 3841 9106 3845 9114
rect 3852 9106 3856 9114
rect 3869 9106 3873 9114
rect 3886 9106 3890 9114
rect 3895 9106 3899 9114
rect 3908 9106 3912 9114
rect 3916 9106 3920 9114
rect 3924 9106 3928 9114
rect 3941 9106 3945 9114
rect 3951 9106 3955 9114
rect 3959 9106 3963 9114
rect 3999 9113 4003 9121
rect 4014 9113 4018 9121
rect 4029 9119 4033 9127
rect 4037 9119 4041 9127
rect 4080 9119 4084 9127
rect 4088 9119 4092 9127
rect 3366 9090 3370 9098
rect 3374 9090 3378 9098
rect 3390 9084 3394 9092
rect 3405 9084 3409 9092
rect 3420 9090 3424 9098
rect 3428 9090 3432 9098
rect 3540 9065 3556 9095
rect 3560 9065 3576 9095
rect 3593 9065 3609 9095
rect 3613 9065 3629 9095
rect 4104 9113 4108 9121
rect 4119 9113 4123 9121
rect 4134 9119 4138 9127
rect 4142 9119 4146 9127
rect 2856 9020 2860 9028
rect 2864 9020 2868 9028
rect 2872 9020 2876 9028
rect 2880 9020 2884 9028
rect 2888 9020 2892 9028
rect 2896 9020 2900 9028
rect 2907 9020 2911 9028
rect 2924 9020 2928 9028
rect 2941 9020 2945 9028
rect 2950 9020 2954 9028
rect 2963 9020 2967 9028
rect 2971 9020 2975 9028
rect 2979 9020 2983 9028
rect 2996 9020 3000 9028
rect 3006 9020 3010 9028
rect 3014 9020 3018 9028
rect 3054 9022 3058 9030
rect 3069 9022 3073 9030
rect 3159 9022 3163 9030
rect 3174 9022 3178 9030
rect 3801 9020 3805 9028
rect 3809 9020 3813 9028
rect 3817 9020 3821 9028
rect 3825 9020 3829 9028
rect 3833 9020 3837 9028
rect 3841 9020 3845 9028
rect 3852 9020 3856 9028
rect 3869 9020 3873 9028
rect 3886 9020 3890 9028
rect 3895 9020 3899 9028
rect 3908 9020 3912 9028
rect 3916 9020 3920 9028
rect 3924 9020 3928 9028
rect 3941 9020 3945 9028
rect 3951 9020 3955 9028
rect 3959 9020 3963 9028
rect 3999 9022 4003 9030
rect 4014 9022 4018 9030
rect 4104 9022 4108 9030
rect 4119 9022 4123 9030
rect 2856 8974 2860 8982
rect 2864 8974 2868 8982
rect 2872 8974 2876 8982
rect 2880 8974 2884 8982
rect 2888 8974 2892 8982
rect 2896 8974 2900 8982
rect 2907 8974 2911 8982
rect 2924 8974 2928 8982
rect 2941 8974 2945 8982
rect 2950 8974 2954 8982
rect 2963 8974 2967 8982
rect 2971 8974 2975 8982
rect 2979 8974 2983 8982
rect 2996 8974 3000 8982
rect 3006 8974 3010 8982
rect 3014 8974 3018 8982
rect 3054 8981 3058 8989
rect 3069 8981 3073 8989
rect 3084 8987 3088 8995
rect 3092 8987 3096 8995
rect 3111 8987 3115 8995
rect 3119 8987 3123 8995
rect 3135 8981 3139 8989
rect 3150 8981 3154 8989
rect 3165 8987 3169 8995
rect 3173 8987 3177 8995
rect 3201 8987 3205 8995
rect 3209 8987 3213 8995
rect 3225 8981 3229 8989
rect 3240 8981 3244 8989
rect 3255 8987 3259 8995
rect 3263 8987 3267 8995
rect 3390 8988 3394 8996
rect 3405 8988 3409 8996
rect 3801 8974 3805 8982
rect 3809 8974 3813 8982
rect 3817 8974 3821 8982
rect 3825 8974 3829 8982
rect 3833 8974 3837 8982
rect 3841 8974 3845 8982
rect 3852 8974 3856 8982
rect 3869 8974 3873 8982
rect 3886 8974 3890 8982
rect 3895 8974 3899 8982
rect 3908 8974 3912 8982
rect 3916 8974 3920 8982
rect 3924 8974 3928 8982
rect 3941 8974 3945 8982
rect 3951 8974 3955 8982
rect 3959 8974 3963 8982
rect 3999 8981 4003 8989
rect 4014 8981 4018 8989
rect 4029 8987 4033 8995
rect 4037 8987 4041 8995
rect 4056 8987 4060 8995
rect 4064 8987 4068 8995
rect 3344 8960 3348 8968
rect 3352 8960 3356 8968
rect 3366 8960 3370 8968
rect 3374 8960 3378 8968
rect 3390 8954 3394 8962
rect 3405 8954 3409 8962
rect 3420 8960 3424 8968
rect 3428 8960 3432 8968
rect 3446 8935 3462 8965
rect 3466 8935 3482 8965
rect 3499 8935 3515 8965
rect 3519 8935 3535 8965
rect 4080 8981 4084 8989
rect 4095 8981 4099 8989
rect 4110 8987 4114 8995
rect 4118 8987 4122 8995
rect 4146 8987 4150 8995
rect 4154 8987 4158 8995
rect 4170 8981 4174 8989
rect 4185 8981 4189 8989
rect 4200 8987 4204 8995
rect 4208 8987 4212 8995
rect 2856 8888 2860 8896
rect 2864 8888 2868 8896
rect 2872 8888 2876 8896
rect 2880 8888 2884 8896
rect 2888 8888 2892 8896
rect 2896 8888 2900 8896
rect 2907 8888 2911 8896
rect 2924 8888 2928 8896
rect 2941 8888 2945 8896
rect 2950 8888 2954 8896
rect 2963 8888 2967 8896
rect 2971 8888 2975 8896
rect 2979 8888 2983 8896
rect 2996 8888 3000 8896
rect 3006 8888 3010 8896
rect 3014 8888 3018 8896
rect 3054 8887 3058 8895
rect 3069 8887 3073 8895
rect 3135 8887 3139 8895
rect 3150 8887 3154 8895
rect 3225 8887 3229 8895
rect 3240 8887 3244 8895
rect 3801 8888 3805 8896
rect 3809 8888 3813 8896
rect 3817 8888 3821 8896
rect 3825 8888 3829 8896
rect 3833 8888 3837 8896
rect 3841 8888 3845 8896
rect 3852 8888 3856 8896
rect 3869 8888 3873 8896
rect 3886 8888 3890 8896
rect 3895 8888 3899 8896
rect 3908 8888 3912 8896
rect 3916 8888 3920 8896
rect 3924 8888 3928 8896
rect 3941 8888 3945 8896
rect 3951 8888 3955 8896
rect 3959 8888 3963 8896
rect 3999 8887 4003 8895
rect 4014 8887 4018 8895
rect 4080 8887 4084 8895
rect 4095 8887 4099 8895
rect 4170 8887 4174 8895
rect 4185 8887 4189 8895
rect 2856 8842 2860 8850
rect 2864 8842 2868 8850
rect 2872 8842 2876 8850
rect 2880 8842 2884 8850
rect 2888 8842 2892 8850
rect 2896 8842 2900 8850
rect 2907 8842 2911 8850
rect 2924 8842 2928 8850
rect 2941 8842 2945 8850
rect 2950 8842 2954 8850
rect 2963 8842 2967 8850
rect 2971 8842 2975 8850
rect 2979 8842 2983 8850
rect 2996 8842 3000 8850
rect 3006 8842 3010 8850
rect 3014 8842 3018 8850
rect 3054 8849 3058 8857
rect 3069 8849 3073 8857
rect 3084 8855 3088 8863
rect 3092 8855 3096 8863
rect 3390 8858 3394 8866
rect 3405 8858 3409 8866
rect 3801 8842 3805 8850
rect 3809 8842 3813 8850
rect 3817 8842 3821 8850
rect 3825 8842 3829 8850
rect 3833 8842 3837 8850
rect 3841 8842 3845 8850
rect 3852 8842 3856 8850
rect 3869 8842 3873 8850
rect 3886 8842 3890 8850
rect 3895 8842 3899 8850
rect 3908 8842 3912 8850
rect 3916 8842 3920 8850
rect 3924 8842 3928 8850
rect 3941 8842 3945 8850
rect 3951 8842 3955 8850
rect 3959 8842 3963 8850
rect 3999 8849 4003 8857
rect 4014 8849 4018 8857
rect 4029 8855 4033 8863
rect 4037 8855 4041 8863
rect 2367 8787 2371 8795
rect 2380 8787 2384 8795
rect 2388 8787 2392 8795
rect 2396 8791 2400 8795
rect 2404 8787 2408 8795
rect 2417 8787 2421 8795
rect 2430 8787 2434 8795
rect 2438 8787 2442 8795
rect 2446 8787 2450 8795
rect 2454 8791 2458 8795
rect 2462 8787 2466 8795
rect 2475 8787 2479 8795
rect 2483 8787 2487 8795
rect 2491 8787 2495 8795
rect 2499 8787 2503 8795
rect 2512 8787 2516 8795
rect 2520 8787 2524 8795
rect 2528 8791 2532 8795
rect 2536 8787 2540 8795
rect 2549 8787 2553 8795
rect 2562 8787 2566 8795
rect 2570 8787 2574 8795
rect 2578 8787 2582 8795
rect 2586 8791 2590 8795
rect 2594 8787 2598 8795
rect 2607 8787 2611 8795
rect 2615 8787 2619 8795
rect 2623 8787 2627 8795
rect 2631 8787 2635 8795
rect 2644 8787 2648 8795
rect 2652 8787 2656 8795
rect 2660 8791 2664 8795
rect 2668 8787 2672 8795
rect 2681 8787 2685 8795
rect 2694 8787 2698 8795
rect 2702 8787 2706 8795
rect 2710 8787 2714 8795
rect 2718 8791 2722 8795
rect 2726 8787 2730 8795
rect 2739 8787 2743 8795
rect 2747 8787 2751 8795
rect 2755 8787 2759 8795
rect 3312 8787 3316 8795
rect 3325 8787 3329 8795
rect 3333 8787 3337 8795
rect 3341 8791 3345 8795
rect 3349 8787 3353 8795
rect 3362 8787 3366 8795
rect 3375 8787 3379 8795
rect 3383 8787 3387 8795
rect 3391 8787 3395 8795
rect 3399 8791 3403 8795
rect 3407 8787 3411 8795
rect 3420 8787 3424 8795
rect 3428 8787 3432 8795
rect 3436 8787 3440 8795
rect 3444 8787 3448 8795
rect 3457 8787 3461 8795
rect 3465 8787 3469 8795
rect 3473 8791 3477 8795
rect 3481 8787 3485 8795
rect 3494 8787 3498 8795
rect 3507 8787 3511 8795
rect 3515 8787 3519 8795
rect 3523 8787 3527 8795
rect 3531 8791 3535 8795
rect 3539 8787 3543 8795
rect 3552 8787 3556 8795
rect 3560 8787 3564 8795
rect 3568 8787 3572 8795
rect 3576 8787 3580 8795
rect 3589 8787 3593 8795
rect 3597 8787 3601 8795
rect 3605 8791 3609 8795
rect 3613 8787 3617 8795
rect 3626 8787 3630 8795
rect 3639 8787 3643 8795
rect 3647 8787 3651 8795
rect 3655 8787 3659 8795
rect 3663 8791 3667 8795
rect 3671 8787 3675 8795
rect 3684 8787 3688 8795
rect 3692 8787 3696 8795
rect 3700 8787 3704 8795
rect 2856 8756 2860 8764
rect 2864 8756 2868 8764
rect 2872 8756 2876 8764
rect 2880 8756 2884 8764
rect 2888 8756 2892 8764
rect 2896 8756 2900 8764
rect 2907 8756 2911 8764
rect 2924 8756 2928 8764
rect 2941 8756 2945 8764
rect 2950 8756 2954 8764
rect 2963 8756 2967 8764
rect 2971 8756 2975 8764
rect 2979 8756 2983 8764
rect 2996 8756 3000 8764
rect 3006 8756 3010 8764
rect 3014 8756 3018 8764
rect 3054 8751 3058 8759
rect 3069 8751 3073 8759
rect 3090 8756 3094 8764
rect 3098 8756 3102 8764
rect 3108 8756 3112 8764
rect 3116 8756 3120 8764
rect 3125 8756 3129 8764
rect 3133 8756 3137 8764
rect 3141 8756 3145 8764
rect 3149 8756 3153 8764
rect 3157 8756 3161 8764
rect 3168 8756 3172 8764
rect 3185 8756 3189 8764
rect 3202 8756 3206 8764
rect 3211 8756 3215 8764
rect 3224 8756 3228 8764
rect 3232 8756 3236 8764
rect 3240 8756 3244 8764
rect 3257 8756 3261 8764
rect 3267 8756 3271 8764
rect 3275 8756 3279 8764
rect 3801 8756 3805 8764
rect 3809 8756 3813 8764
rect 3817 8756 3821 8764
rect 3825 8756 3829 8764
rect 3833 8756 3837 8764
rect 3841 8756 3845 8764
rect 3852 8756 3856 8764
rect 3869 8756 3873 8764
rect 3886 8756 3890 8764
rect 3895 8756 3899 8764
rect 3908 8756 3912 8764
rect 3916 8756 3920 8764
rect 3924 8756 3928 8764
rect 3941 8756 3945 8764
rect 3951 8756 3955 8764
rect 3959 8756 3963 8764
rect 3999 8751 4003 8759
rect 4014 8751 4018 8759
rect 4035 8756 4039 8764
rect 4043 8756 4047 8764
rect 4053 8756 4057 8764
rect 4061 8756 4065 8764
rect 4070 8756 4074 8764
rect 4078 8756 4082 8764
rect 4086 8756 4090 8764
rect 4094 8756 4098 8764
rect 4102 8756 4106 8764
rect 4113 8756 4117 8764
rect 4130 8756 4134 8764
rect 4147 8756 4151 8764
rect 4156 8756 4160 8764
rect 4169 8756 4173 8764
rect 4177 8756 4181 8764
rect 4185 8756 4189 8764
rect 4202 8756 4206 8764
rect 4212 8756 4216 8764
rect 4220 8756 4224 8764
rect 3150 8675 3154 8683
rect 3163 8675 3167 8683
rect 3171 8675 3175 8683
rect 3179 8679 3183 8683
rect 3187 8675 3191 8683
rect 3200 8675 3204 8683
rect 3213 8675 3217 8683
rect 3221 8675 3225 8683
rect 3229 8675 3233 8683
rect 3237 8679 3241 8683
rect 3245 8675 3249 8683
rect 3258 8675 3262 8683
rect 3266 8675 3270 8683
rect 3274 8675 3278 8683
rect 4095 8675 4099 8683
rect 4108 8675 4112 8683
rect 4116 8675 4120 8683
rect 4124 8679 4128 8683
rect 4132 8675 4136 8683
rect 4145 8675 4149 8683
rect 4158 8675 4162 8683
rect 4166 8675 4170 8683
rect 4174 8675 4178 8683
rect 4182 8679 4186 8683
rect 4190 8675 4194 8683
rect 4203 8675 4207 8683
rect 4211 8675 4215 8683
rect 4219 8675 4223 8683
rect 2367 8645 2371 8653
rect 2380 8645 2384 8653
rect 2388 8645 2392 8653
rect 2396 8649 2400 8653
rect 2404 8645 2408 8653
rect 2417 8645 2421 8653
rect 2430 8645 2434 8653
rect 2438 8645 2442 8653
rect 2446 8645 2450 8653
rect 2454 8649 2458 8653
rect 2462 8645 2466 8653
rect 2475 8645 2479 8653
rect 2483 8645 2487 8653
rect 2491 8645 2495 8653
rect 2499 8645 2503 8653
rect 2512 8645 2516 8653
rect 2520 8645 2524 8653
rect 2528 8649 2532 8653
rect 2536 8645 2540 8653
rect 2549 8645 2553 8653
rect 2562 8645 2566 8653
rect 2570 8645 2574 8653
rect 2578 8645 2582 8653
rect 2586 8649 2590 8653
rect 2594 8645 2598 8653
rect 2607 8645 2611 8653
rect 2615 8645 2619 8653
rect 2623 8645 2627 8653
rect 2631 8645 2635 8653
rect 2644 8645 2648 8653
rect 2652 8645 2656 8653
rect 2660 8649 2664 8653
rect 2668 8645 2672 8653
rect 2681 8645 2685 8653
rect 2694 8645 2698 8653
rect 2702 8645 2706 8653
rect 2710 8645 2714 8653
rect 2718 8649 2722 8653
rect 2726 8645 2730 8653
rect 2739 8645 2743 8653
rect 2747 8645 2751 8653
rect 2755 8645 2759 8653
rect 3312 8645 3316 8653
rect 3325 8645 3329 8653
rect 3333 8645 3337 8653
rect 3341 8649 3345 8653
rect 3349 8645 3353 8653
rect 3362 8645 3366 8653
rect 3375 8645 3379 8653
rect 3383 8645 3387 8653
rect 3391 8645 3395 8653
rect 3399 8649 3403 8653
rect 3407 8645 3411 8653
rect 3420 8645 3424 8653
rect 3428 8645 3432 8653
rect 3436 8645 3440 8653
rect 3444 8645 3448 8653
rect 3457 8645 3461 8653
rect 3465 8645 3469 8653
rect 3473 8649 3477 8653
rect 3481 8645 3485 8653
rect 3494 8645 3498 8653
rect 3507 8645 3511 8653
rect 3515 8645 3519 8653
rect 3523 8645 3527 8653
rect 3531 8649 3535 8653
rect 3539 8645 3543 8653
rect 3552 8645 3556 8653
rect 3560 8645 3564 8653
rect 3568 8645 3572 8653
rect 3576 8645 3580 8653
rect 3589 8645 3593 8653
rect 3597 8645 3601 8653
rect 3605 8649 3609 8653
rect 3613 8645 3617 8653
rect 3626 8645 3630 8653
rect 3639 8645 3643 8653
rect 3647 8645 3651 8653
rect 3655 8645 3659 8653
rect 3663 8649 3667 8653
rect 3671 8645 3675 8653
rect 3684 8645 3688 8653
rect 3692 8645 3696 8653
rect 3700 8645 3704 8653
rect 3150 8589 3154 8597
rect 3163 8589 3167 8597
rect 3171 8589 3175 8597
rect 3179 8593 3183 8597
rect 3187 8589 3191 8597
rect 3200 8589 3204 8597
rect 3213 8589 3217 8597
rect 3221 8589 3225 8597
rect 3229 8589 3233 8597
rect 3237 8593 3241 8597
rect 3245 8589 3249 8597
rect 3258 8589 3262 8597
rect 3266 8589 3270 8597
rect 3274 8589 3278 8597
rect 4095 8589 4099 8597
rect 4108 8589 4112 8597
rect 4116 8589 4120 8597
rect 4124 8593 4128 8597
rect 4132 8589 4136 8597
rect 4145 8589 4149 8597
rect 4158 8589 4162 8597
rect 4166 8589 4170 8597
rect 4174 8589 4178 8597
rect 4182 8593 4186 8597
rect 4190 8589 4194 8597
rect 4203 8589 4207 8597
rect 4211 8589 4215 8597
rect 4219 8589 4223 8597
rect 2367 8559 2371 8567
rect 2380 8559 2384 8567
rect 2388 8559 2392 8567
rect 2396 8563 2400 8567
rect 2404 8559 2408 8567
rect 2417 8559 2421 8567
rect 2430 8559 2434 8567
rect 2438 8559 2442 8567
rect 2446 8559 2450 8567
rect 2454 8563 2458 8567
rect 2462 8559 2466 8567
rect 2475 8559 2479 8567
rect 2483 8559 2487 8567
rect 2491 8559 2495 8567
rect 2499 8559 2503 8567
rect 2512 8559 2516 8567
rect 2520 8559 2524 8567
rect 2528 8563 2532 8567
rect 2536 8559 2540 8567
rect 2549 8559 2553 8567
rect 2562 8559 2566 8567
rect 2570 8559 2574 8567
rect 2578 8559 2582 8567
rect 2586 8563 2590 8567
rect 2594 8559 2598 8567
rect 2607 8559 2611 8567
rect 2615 8559 2619 8567
rect 2623 8559 2627 8567
rect 2631 8559 2635 8567
rect 2644 8559 2648 8567
rect 2652 8559 2656 8567
rect 2660 8563 2664 8567
rect 2668 8559 2672 8567
rect 2681 8559 2685 8567
rect 2694 8559 2698 8567
rect 2702 8559 2706 8567
rect 2710 8559 2714 8567
rect 2718 8563 2722 8567
rect 2726 8559 2730 8567
rect 2739 8559 2743 8567
rect 2747 8559 2751 8567
rect 2755 8559 2759 8567
rect 3312 8559 3316 8567
rect 3325 8559 3329 8567
rect 3333 8559 3337 8567
rect 3341 8563 3345 8567
rect 3349 8559 3353 8567
rect 3362 8559 3366 8567
rect 3375 8559 3379 8567
rect 3383 8559 3387 8567
rect 3391 8559 3395 8567
rect 3399 8563 3403 8567
rect 3407 8559 3411 8567
rect 3420 8559 3424 8567
rect 3428 8559 3432 8567
rect 3436 8559 3440 8567
rect 3444 8559 3448 8567
rect 3457 8559 3461 8567
rect 3465 8559 3469 8567
rect 3473 8563 3477 8567
rect 3481 8559 3485 8567
rect 3494 8559 3498 8567
rect 3507 8559 3511 8567
rect 3515 8559 3519 8567
rect 3523 8559 3527 8567
rect 3531 8563 3535 8567
rect 3539 8559 3543 8567
rect 3552 8559 3556 8567
rect 3560 8559 3564 8567
rect 3568 8559 3572 8567
rect 3576 8559 3580 8567
rect 3589 8559 3593 8567
rect 3597 8559 3601 8567
rect 3605 8563 3609 8567
rect 3613 8559 3617 8567
rect 3626 8559 3630 8567
rect 3639 8559 3643 8567
rect 3647 8559 3651 8567
rect 3655 8559 3659 8567
rect 3663 8563 3667 8567
rect 3671 8559 3675 8567
rect 3684 8559 3688 8567
rect 3692 8559 3696 8567
rect 3700 8559 3704 8567
rect 2367 8419 2371 8427
rect 2380 8419 2384 8427
rect 2388 8419 2392 8427
rect 2396 8423 2400 8427
rect 2404 8419 2408 8427
rect 2417 8419 2421 8427
rect 2430 8419 2434 8427
rect 2438 8419 2442 8427
rect 2446 8419 2450 8427
rect 2454 8423 2458 8427
rect 2462 8419 2466 8427
rect 2475 8419 2479 8427
rect 2483 8419 2487 8427
rect 2491 8419 2495 8427
rect 2499 8419 2503 8427
rect 2512 8419 2516 8427
rect 2520 8419 2524 8427
rect 2528 8423 2532 8427
rect 2536 8419 2540 8427
rect 2549 8419 2553 8427
rect 2562 8419 2566 8427
rect 2570 8419 2574 8427
rect 2578 8419 2582 8427
rect 2586 8423 2590 8427
rect 2594 8419 2598 8427
rect 2607 8419 2611 8427
rect 2615 8419 2619 8427
rect 2623 8419 2627 8427
rect 2631 8419 2635 8427
rect 2644 8419 2648 8427
rect 2652 8419 2656 8427
rect 2660 8423 2664 8427
rect 2668 8419 2672 8427
rect 2681 8419 2685 8427
rect 2694 8419 2698 8427
rect 2702 8419 2706 8427
rect 2710 8419 2714 8427
rect 2718 8423 2722 8427
rect 2726 8419 2730 8427
rect 2739 8419 2743 8427
rect 2747 8419 2751 8427
rect 2755 8419 2759 8427
rect 3312 8419 3316 8427
rect 3325 8419 3329 8427
rect 3333 8419 3337 8427
rect 3341 8423 3345 8427
rect 3349 8419 3353 8427
rect 3362 8419 3366 8427
rect 3375 8419 3379 8427
rect 3383 8419 3387 8427
rect 3391 8419 3395 8427
rect 3399 8423 3403 8427
rect 3407 8419 3411 8427
rect 3420 8419 3424 8427
rect 3428 8419 3432 8427
rect 3436 8419 3440 8427
rect 3444 8419 3448 8427
rect 3457 8419 3461 8427
rect 3465 8419 3469 8427
rect 3473 8423 3477 8427
rect 3481 8419 3485 8427
rect 3494 8419 3498 8427
rect 3507 8419 3511 8427
rect 3515 8419 3519 8427
rect 3523 8419 3527 8427
rect 3531 8423 3535 8427
rect 3539 8419 3543 8427
rect 3552 8419 3556 8427
rect 3560 8419 3564 8427
rect 3568 8419 3572 8427
rect 3576 8419 3580 8427
rect 3589 8419 3593 8427
rect 3597 8419 3601 8427
rect 3605 8423 3609 8427
rect 3613 8419 3617 8427
rect 3626 8419 3630 8427
rect 3639 8419 3643 8427
rect 3647 8419 3651 8427
rect 3655 8419 3659 8427
rect 3663 8423 3667 8427
rect 3671 8419 3675 8427
rect 3684 8419 3688 8427
rect 3692 8419 3696 8427
rect 3700 8419 3704 8427
rect 2851 8340 2855 8348
rect 2864 8340 2868 8348
rect 2872 8340 2876 8348
rect 2880 8344 2884 8348
rect 2888 8340 2892 8348
rect 2901 8340 2905 8348
rect 2914 8340 2918 8348
rect 2922 8340 2926 8348
rect 2930 8340 2934 8348
rect 2938 8344 2942 8348
rect 2946 8340 2950 8348
rect 2959 8340 2963 8348
rect 2967 8340 2971 8348
rect 2975 8340 2979 8348
rect 2983 8340 2987 8348
rect 2996 8340 3000 8348
rect 3004 8340 3008 8348
rect 3012 8344 3016 8348
rect 3020 8340 3024 8348
rect 3033 8340 3037 8348
rect 3046 8340 3050 8348
rect 3054 8340 3058 8348
rect 3062 8340 3066 8348
rect 3070 8344 3074 8348
rect 3078 8340 3082 8348
rect 3091 8340 3095 8348
rect 3099 8340 3103 8348
rect 3107 8340 3111 8348
rect 3115 8340 3119 8348
rect 3128 8340 3132 8348
rect 3136 8340 3140 8348
rect 3144 8344 3148 8348
rect 3152 8340 3156 8348
rect 3165 8340 3169 8348
rect 3178 8340 3182 8348
rect 3186 8340 3190 8348
rect 3194 8340 3198 8348
rect 3202 8344 3206 8348
rect 3210 8340 3214 8348
rect 3223 8340 3227 8348
rect 3231 8340 3235 8348
rect 3239 8340 3243 8348
rect 3247 8340 3251 8348
rect 3260 8340 3264 8348
rect 3268 8340 3272 8348
rect 3276 8344 3280 8348
rect 3284 8340 3288 8348
rect 3297 8340 3301 8348
rect 3310 8340 3314 8348
rect 3318 8340 3322 8348
rect 3326 8340 3330 8348
rect 3334 8344 3338 8348
rect 3342 8340 3346 8348
rect 3355 8340 3359 8348
rect 3363 8340 3367 8348
rect 3371 8340 3375 8348
rect 3796 8340 3800 8348
rect 3809 8340 3813 8348
rect 3817 8340 3821 8348
rect 3825 8344 3829 8348
rect 3833 8340 3837 8348
rect 3846 8340 3850 8348
rect 3859 8340 3863 8348
rect 3867 8340 3871 8348
rect 3875 8340 3879 8348
rect 3883 8344 3887 8348
rect 3891 8340 3895 8348
rect 3904 8340 3908 8348
rect 3912 8340 3916 8348
rect 3920 8340 3924 8348
rect 3928 8340 3932 8348
rect 3941 8340 3945 8348
rect 3949 8340 3953 8348
rect 3957 8344 3961 8348
rect 3965 8340 3969 8348
rect 3978 8340 3982 8348
rect 3991 8340 3995 8348
rect 3999 8340 4003 8348
rect 4007 8340 4011 8348
rect 4015 8344 4019 8348
rect 4023 8340 4027 8348
rect 4036 8340 4040 8348
rect 4044 8340 4048 8348
rect 4052 8340 4056 8348
rect 4060 8340 4064 8348
rect 4073 8340 4077 8348
rect 4081 8340 4085 8348
rect 4089 8344 4093 8348
rect 4097 8340 4101 8348
rect 4110 8340 4114 8348
rect 4123 8340 4127 8348
rect 4131 8340 4135 8348
rect 4139 8340 4143 8348
rect 4147 8344 4151 8348
rect 4155 8340 4159 8348
rect 4168 8340 4172 8348
rect 4176 8340 4180 8348
rect 4184 8340 4188 8348
rect 4192 8340 4196 8348
rect 4205 8340 4209 8348
rect 4213 8340 4217 8348
rect 4221 8344 4225 8348
rect 4229 8340 4233 8348
rect 4242 8340 4246 8348
rect 4255 8340 4259 8348
rect 4263 8340 4267 8348
rect 4271 8340 4275 8348
rect 4279 8344 4283 8348
rect 4287 8340 4291 8348
rect 4300 8340 4304 8348
rect 4308 8340 4312 8348
rect 4316 8340 4320 8348
rect 2499 8307 2503 8315
rect 2512 8307 2516 8315
rect 2520 8307 2524 8315
rect 2528 8311 2532 8315
rect 2536 8307 2540 8315
rect 2549 8307 2553 8315
rect 2562 8307 2566 8315
rect 2570 8307 2574 8315
rect 2578 8307 2582 8315
rect 2586 8311 2590 8315
rect 2594 8307 2598 8315
rect 2607 8307 2611 8315
rect 2615 8307 2619 8315
rect 2623 8307 2627 8315
rect 3444 8307 3448 8315
rect 3457 8307 3461 8315
rect 3465 8307 3469 8315
rect 3473 8311 3477 8315
rect 3481 8307 3485 8315
rect 3494 8307 3498 8315
rect 3507 8307 3511 8315
rect 3515 8307 3519 8315
rect 3523 8307 3527 8315
rect 3531 8311 3535 8315
rect 3539 8307 3543 8315
rect 3552 8307 3556 8315
rect 3560 8307 3564 8315
rect 3568 8307 3572 8315
rect 3030 8269 3034 8277
rect 3038 8269 3042 8277
rect 2856 8256 2860 8264
rect 2864 8256 2868 8264
rect 2872 8256 2876 8264
rect 2880 8256 2884 8264
rect 2888 8256 2892 8264
rect 2896 8256 2900 8264
rect 2907 8256 2911 8264
rect 2924 8256 2928 8264
rect 2941 8256 2945 8264
rect 2950 8256 2954 8264
rect 2963 8256 2967 8264
rect 2971 8256 2975 8264
rect 2979 8256 2983 8264
rect 2996 8256 3000 8264
rect 3006 8256 3010 8264
rect 3014 8256 3018 8264
rect 3054 8263 3058 8271
rect 3069 8263 3073 8271
rect 3084 8269 3088 8277
rect 3092 8269 3096 8277
rect 3111 8269 3115 8277
rect 3119 8269 3123 8277
rect 3135 8263 3139 8271
rect 3150 8263 3154 8271
rect 3165 8269 3169 8277
rect 3173 8269 3177 8277
rect 3975 8269 3979 8277
rect 3983 8269 3987 8277
rect 3801 8256 3805 8264
rect 3809 8256 3813 8264
rect 3817 8256 3821 8264
rect 3825 8256 3829 8264
rect 3833 8256 3837 8264
rect 3841 8256 3845 8264
rect 3852 8256 3856 8264
rect 3869 8256 3873 8264
rect 3886 8256 3890 8264
rect 3895 8256 3899 8264
rect 3908 8256 3912 8264
rect 3916 8256 3920 8264
rect 3924 8256 3928 8264
rect 3941 8256 3945 8264
rect 3951 8256 3955 8264
rect 3959 8256 3963 8264
rect 3999 8263 4003 8271
rect 4014 8263 4018 8271
rect 4029 8269 4033 8277
rect 4037 8269 4041 8277
rect 4056 8269 4060 8277
rect 4064 8269 4068 8277
rect 4080 8263 4084 8271
rect 4095 8263 4099 8271
rect 4110 8269 4114 8277
rect 4118 8269 4122 8277
rect 2490 8205 2494 8213
rect 2498 8205 2502 8213
rect 2506 8205 2510 8213
rect 2519 8205 2523 8213
rect 2527 8209 2531 8213
rect 2535 8205 2539 8213
rect 2543 8205 2547 8213
rect 2551 8205 2555 8213
rect 2564 8205 2568 8213
rect 2577 8205 2581 8213
rect 2585 8209 2589 8213
rect 2593 8205 2597 8213
rect 2601 8205 2605 8213
rect 2614 8205 2618 8213
rect 3435 8205 3439 8213
rect 3443 8205 3447 8213
rect 3451 8205 3455 8213
rect 3464 8205 3468 8213
rect 3472 8209 3476 8213
rect 3480 8205 3484 8213
rect 3488 8205 3492 8213
rect 3496 8205 3500 8213
rect 3509 8205 3513 8213
rect 3522 8205 3526 8213
rect 3530 8209 3534 8213
rect 3538 8205 3542 8213
rect 3546 8205 3550 8213
rect 3559 8205 3563 8213
rect 2856 8170 2860 8178
rect 2864 8170 2868 8178
rect 2872 8170 2876 8178
rect 2880 8170 2884 8178
rect 2888 8170 2892 8178
rect 2896 8170 2900 8178
rect 2907 8170 2911 8178
rect 2924 8170 2928 8178
rect 2941 8170 2945 8178
rect 2950 8170 2954 8178
rect 2963 8170 2967 8178
rect 2971 8170 2975 8178
rect 2979 8170 2983 8178
rect 2996 8170 3000 8178
rect 3006 8170 3010 8178
rect 3014 8170 3018 8178
rect 3054 8171 3058 8179
rect 3069 8171 3073 8179
rect 3135 8171 3139 8179
rect 3150 8171 3154 8179
rect 3801 8170 3805 8178
rect 3809 8170 3813 8178
rect 3817 8170 3821 8178
rect 3825 8170 3829 8178
rect 3833 8170 3837 8178
rect 3841 8170 3845 8178
rect 3852 8170 3856 8178
rect 3869 8170 3873 8178
rect 3886 8170 3890 8178
rect 3895 8170 3899 8178
rect 3908 8170 3912 8178
rect 3916 8170 3920 8178
rect 3924 8170 3928 8178
rect 3941 8170 3945 8178
rect 3951 8170 3955 8178
rect 3959 8170 3963 8178
rect 3999 8171 4003 8179
rect 4014 8171 4018 8179
rect 4080 8171 4084 8179
rect 4095 8171 4099 8179
rect 2856 8124 2860 8132
rect 2864 8124 2868 8132
rect 2872 8124 2876 8132
rect 2880 8124 2884 8132
rect 2888 8124 2892 8132
rect 2896 8124 2900 8132
rect 2907 8124 2911 8132
rect 2924 8124 2928 8132
rect 2941 8124 2945 8132
rect 2950 8124 2954 8132
rect 2963 8124 2967 8132
rect 2971 8124 2975 8132
rect 2979 8124 2983 8132
rect 2996 8124 3000 8132
rect 3006 8124 3010 8132
rect 3014 8124 3018 8132
rect 3054 8131 3058 8139
rect 3069 8131 3073 8139
rect 3084 8137 3088 8145
rect 3092 8137 3096 8145
rect 3135 8137 3139 8145
rect 3143 8137 3147 8145
rect 3159 8131 3163 8139
rect 3174 8131 3178 8139
rect 3189 8137 3193 8145
rect 3197 8137 3201 8145
rect 3801 8124 3805 8132
rect 3809 8124 3813 8132
rect 3817 8124 3821 8132
rect 3825 8124 3829 8132
rect 3833 8124 3837 8132
rect 3841 8124 3845 8132
rect 3852 8124 3856 8132
rect 3869 8124 3873 8132
rect 3886 8124 3890 8132
rect 3895 8124 3899 8132
rect 3908 8124 3912 8132
rect 3916 8124 3920 8132
rect 3924 8124 3928 8132
rect 3941 8124 3945 8132
rect 3951 8124 3955 8132
rect 3959 8124 3963 8132
rect 3999 8131 4003 8139
rect 4014 8131 4018 8139
rect 4029 8137 4033 8145
rect 4037 8137 4041 8145
rect 4080 8137 4084 8145
rect 4088 8137 4092 8145
rect 4104 8131 4108 8139
rect 4119 8131 4123 8139
rect 4134 8137 4138 8145
rect 4142 8137 4146 8145
rect 2856 8038 2860 8046
rect 2864 8038 2868 8046
rect 2872 8038 2876 8046
rect 2880 8038 2884 8046
rect 2888 8038 2892 8046
rect 2896 8038 2900 8046
rect 2907 8038 2911 8046
rect 2924 8038 2928 8046
rect 2941 8038 2945 8046
rect 2950 8038 2954 8046
rect 2963 8038 2967 8046
rect 2971 8038 2975 8046
rect 2979 8038 2983 8046
rect 2996 8038 3000 8046
rect 3006 8038 3010 8046
rect 3014 8038 3018 8046
rect 3054 8040 3058 8048
rect 3069 8040 3073 8048
rect 3159 8040 3163 8048
rect 3174 8040 3178 8048
rect 3801 8038 3805 8046
rect 3809 8038 3813 8046
rect 3817 8038 3821 8046
rect 3825 8038 3829 8046
rect 3833 8038 3837 8046
rect 3841 8038 3845 8046
rect 3852 8038 3856 8046
rect 3869 8038 3873 8046
rect 3886 8038 3890 8046
rect 3895 8038 3899 8046
rect 3908 8038 3912 8046
rect 3916 8038 3920 8046
rect 3924 8038 3928 8046
rect 3941 8038 3945 8046
rect 3951 8038 3955 8046
rect 3959 8038 3963 8046
rect 3999 8040 4003 8048
rect 4014 8040 4018 8048
rect 4104 8040 4108 8048
rect 4119 8040 4123 8048
rect 2856 7992 2860 8000
rect 2864 7992 2868 8000
rect 2872 7992 2876 8000
rect 2880 7992 2884 8000
rect 2888 7992 2892 8000
rect 2896 7992 2900 8000
rect 2907 7992 2911 8000
rect 2924 7992 2928 8000
rect 2941 7992 2945 8000
rect 2950 7992 2954 8000
rect 2963 7992 2967 8000
rect 2971 7992 2975 8000
rect 2979 7992 2983 8000
rect 2996 7992 3000 8000
rect 3006 7992 3010 8000
rect 3014 7992 3018 8000
rect 3054 7999 3058 8007
rect 3069 7999 3073 8007
rect 3084 8005 3088 8013
rect 3092 8005 3096 8013
rect 3111 8005 3115 8013
rect 3119 8005 3123 8013
rect 3135 7999 3139 8007
rect 3150 7999 3154 8007
rect 3165 8005 3169 8013
rect 3173 8005 3177 8013
rect 3201 8005 3205 8013
rect 3209 8005 3213 8013
rect 3225 7999 3229 8007
rect 3240 7999 3244 8007
rect 3255 8005 3259 8013
rect 3263 8005 3267 8013
rect 3801 7992 3805 8000
rect 3809 7992 3813 8000
rect 3817 7992 3821 8000
rect 3825 7992 3829 8000
rect 3833 7992 3837 8000
rect 3841 7992 3845 8000
rect 3852 7992 3856 8000
rect 3869 7992 3873 8000
rect 3886 7992 3890 8000
rect 3895 7992 3899 8000
rect 3908 7992 3912 8000
rect 3916 7992 3920 8000
rect 3924 7992 3928 8000
rect 3941 7992 3945 8000
rect 3951 7992 3955 8000
rect 3959 7992 3963 8000
rect 3999 7999 4003 8007
rect 4014 7999 4018 8007
rect 4029 8005 4033 8013
rect 4037 8005 4041 8013
rect 4056 8005 4060 8013
rect 4064 8005 4068 8013
rect 4080 7999 4084 8007
rect 4095 7999 4099 8007
rect 4110 8005 4114 8013
rect 4118 8005 4122 8013
rect 4146 8005 4150 8013
rect 4154 8005 4158 8013
rect 4170 7999 4174 8007
rect 4185 7999 4189 8007
rect 4200 8005 4204 8013
rect 4208 8005 4212 8013
rect 2856 7906 2860 7914
rect 2864 7906 2868 7914
rect 2872 7906 2876 7914
rect 2880 7906 2884 7914
rect 2888 7906 2892 7914
rect 2896 7906 2900 7914
rect 2907 7906 2911 7914
rect 2924 7906 2928 7914
rect 2941 7906 2945 7914
rect 2950 7906 2954 7914
rect 2963 7906 2967 7914
rect 2971 7906 2975 7914
rect 2979 7906 2983 7914
rect 2996 7906 3000 7914
rect 3006 7906 3010 7914
rect 3014 7906 3018 7914
rect 3054 7905 3058 7913
rect 3069 7905 3073 7913
rect 3135 7905 3139 7913
rect 3150 7905 3154 7913
rect 3225 7905 3229 7913
rect 3240 7905 3244 7913
rect 3801 7906 3805 7914
rect 3809 7906 3813 7914
rect 3817 7906 3821 7914
rect 3825 7906 3829 7914
rect 3833 7906 3837 7914
rect 3841 7906 3845 7914
rect 3852 7906 3856 7914
rect 3869 7906 3873 7914
rect 3886 7906 3890 7914
rect 3895 7906 3899 7914
rect 3908 7906 3912 7914
rect 3916 7906 3920 7914
rect 3924 7906 3928 7914
rect 3941 7906 3945 7914
rect 3951 7906 3955 7914
rect 3959 7906 3963 7914
rect 3999 7905 4003 7913
rect 4014 7905 4018 7913
rect 4080 7905 4084 7913
rect 4095 7905 4099 7913
rect 4170 7905 4174 7913
rect 4185 7905 4189 7913
rect 2856 7860 2860 7868
rect 2864 7860 2868 7868
rect 2872 7860 2876 7868
rect 2880 7860 2884 7868
rect 2888 7860 2892 7868
rect 2896 7860 2900 7868
rect 2907 7860 2911 7868
rect 2924 7860 2928 7868
rect 2941 7860 2945 7868
rect 2950 7860 2954 7868
rect 2963 7860 2967 7868
rect 2971 7860 2975 7868
rect 2979 7860 2983 7868
rect 2996 7860 3000 7868
rect 3006 7860 3010 7868
rect 3014 7860 3018 7868
rect 3054 7867 3058 7875
rect 3069 7867 3073 7875
rect 3084 7873 3088 7881
rect 3092 7873 3096 7881
rect 3801 7860 3805 7868
rect 3809 7860 3813 7868
rect 3817 7860 3821 7868
rect 3825 7860 3829 7868
rect 3833 7860 3837 7868
rect 3841 7860 3845 7868
rect 3852 7860 3856 7868
rect 3869 7860 3873 7868
rect 3886 7860 3890 7868
rect 3895 7860 3899 7868
rect 3908 7860 3912 7868
rect 3916 7860 3920 7868
rect 3924 7860 3928 7868
rect 3941 7860 3945 7868
rect 3951 7860 3955 7868
rect 3959 7860 3963 7868
rect 3999 7867 4003 7875
rect 4014 7867 4018 7875
rect 4029 7873 4033 7881
rect 4037 7873 4041 7881
rect 2367 7805 2371 7813
rect 2380 7805 2384 7813
rect 2388 7805 2392 7813
rect 2396 7809 2400 7813
rect 2404 7805 2408 7813
rect 2417 7805 2421 7813
rect 2430 7805 2434 7813
rect 2438 7805 2442 7813
rect 2446 7805 2450 7813
rect 2454 7809 2458 7813
rect 2462 7805 2466 7813
rect 2475 7805 2479 7813
rect 2483 7805 2487 7813
rect 2491 7805 2495 7813
rect 2499 7805 2503 7813
rect 2512 7805 2516 7813
rect 2520 7805 2524 7813
rect 2528 7809 2532 7813
rect 2536 7805 2540 7813
rect 2549 7805 2553 7813
rect 2562 7805 2566 7813
rect 2570 7805 2574 7813
rect 2578 7805 2582 7813
rect 2586 7809 2590 7813
rect 2594 7805 2598 7813
rect 2607 7805 2611 7813
rect 2615 7805 2619 7813
rect 2623 7805 2627 7813
rect 2631 7805 2635 7813
rect 2644 7805 2648 7813
rect 2652 7805 2656 7813
rect 2660 7809 2664 7813
rect 2668 7805 2672 7813
rect 2681 7805 2685 7813
rect 2694 7805 2698 7813
rect 2702 7805 2706 7813
rect 2710 7805 2714 7813
rect 2718 7809 2722 7813
rect 2726 7805 2730 7813
rect 2739 7805 2743 7813
rect 2747 7805 2751 7813
rect 2755 7805 2759 7813
rect 3312 7805 3316 7813
rect 3325 7805 3329 7813
rect 3333 7805 3337 7813
rect 3341 7809 3345 7813
rect 3349 7805 3353 7813
rect 3362 7805 3366 7813
rect 3375 7805 3379 7813
rect 3383 7805 3387 7813
rect 3391 7805 3395 7813
rect 3399 7809 3403 7813
rect 3407 7805 3411 7813
rect 3420 7805 3424 7813
rect 3428 7805 3432 7813
rect 3436 7805 3440 7813
rect 3444 7805 3448 7813
rect 3457 7805 3461 7813
rect 3465 7805 3469 7813
rect 3473 7809 3477 7813
rect 3481 7805 3485 7813
rect 3494 7805 3498 7813
rect 3507 7805 3511 7813
rect 3515 7805 3519 7813
rect 3523 7805 3527 7813
rect 3531 7809 3535 7813
rect 3539 7805 3543 7813
rect 3552 7805 3556 7813
rect 3560 7805 3564 7813
rect 3568 7805 3572 7813
rect 3576 7805 3580 7813
rect 3589 7805 3593 7813
rect 3597 7805 3601 7813
rect 3605 7809 3609 7813
rect 3613 7805 3617 7813
rect 3626 7805 3630 7813
rect 3639 7805 3643 7813
rect 3647 7805 3651 7813
rect 3655 7805 3659 7813
rect 3663 7809 3667 7813
rect 3671 7805 3675 7813
rect 3684 7805 3688 7813
rect 3692 7805 3696 7813
rect 3700 7805 3704 7813
rect 2856 7774 2860 7782
rect 2864 7774 2868 7782
rect 2872 7774 2876 7782
rect 2880 7774 2884 7782
rect 2888 7774 2892 7782
rect 2896 7774 2900 7782
rect 2907 7774 2911 7782
rect 2924 7774 2928 7782
rect 2941 7774 2945 7782
rect 2950 7774 2954 7782
rect 2963 7774 2967 7782
rect 2971 7774 2975 7782
rect 2979 7774 2983 7782
rect 2996 7774 3000 7782
rect 3006 7774 3010 7782
rect 3014 7774 3018 7782
rect 3054 7769 3058 7777
rect 3069 7769 3073 7777
rect 3090 7774 3094 7782
rect 3098 7774 3102 7782
rect 3108 7774 3112 7782
rect 3116 7774 3120 7782
rect 3125 7774 3129 7782
rect 3133 7774 3137 7782
rect 3141 7774 3145 7782
rect 3149 7774 3153 7782
rect 3157 7774 3161 7782
rect 3168 7774 3172 7782
rect 3185 7774 3189 7782
rect 3202 7774 3206 7782
rect 3211 7774 3215 7782
rect 3224 7774 3228 7782
rect 3232 7774 3236 7782
rect 3240 7774 3244 7782
rect 3257 7774 3261 7782
rect 3267 7774 3271 7782
rect 3275 7774 3279 7782
rect 3801 7774 3805 7782
rect 3809 7774 3813 7782
rect 3817 7774 3821 7782
rect 3825 7774 3829 7782
rect 3833 7774 3837 7782
rect 3841 7774 3845 7782
rect 3852 7774 3856 7782
rect 3869 7774 3873 7782
rect 3886 7774 3890 7782
rect 3895 7774 3899 7782
rect 3908 7774 3912 7782
rect 3916 7774 3920 7782
rect 3924 7774 3928 7782
rect 3941 7774 3945 7782
rect 3951 7774 3955 7782
rect 3959 7774 3963 7782
rect 3999 7769 4003 7777
rect 4014 7769 4018 7777
rect 4035 7774 4039 7782
rect 4043 7774 4047 7782
rect 4053 7774 4057 7782
rect 4061 7774 4065 7782
rect 4070 7774 4074 7782
rect 4078 7774 4082 7782
rect 4086 7774 4090 7782
rect 4094 7774 4098 7782
rect 4102 7774 4106 7782
rect 4113 7774 4117 7782
rect 4130 7774 4134 7782
rect 4147 7774 4151 7782
rect 4156 7774 4160 7782
rect 4169 7774 4173 7782
rect 4177 7774 4181 7782
rect 4185 7774 4189 7782
rect 4202 7774 4206 7782
rect 4212 7774 4216 7782
rect 4220 7774 4224 7782
rect 3150 7693 3154 7701
rect 3163 7693 3167 7701
rect 3171 7693 3175 7701
rect 3179 7697 3183 7701
rect 3187 7693 3191 7701
rect 3200 7693 3204 7701
rect 3213 7693 3217 7701
rect 3221 7693 3225 7701
rect 3229 7693 3233 7701
rect 3237 7697 3241 7701
rect 3245 7693 3249 7701
rect 3258 7693 3262 7701
rect 3266 7693 3270 7701
rect 3274 7693 3278 7701
rect 4095 7693 4099 7701
rect 4108 7693 4112 7701
rect 4116 7693 4120 7701
rect 4124 7697 4128 7701
rect 4132 7693 4136 7701
rect 4145 7693 4149 7701
rect 4158 7693 4162 7701
rect 4166 7693 4170 7701
rect 4174 7693 4178 7701
rect 4182 7697 4186 7701
rect 4190 7693 4194 7701
rect 4203 7693 4207 7701
rect 4211 7693 4215 7701
rect 4219 7693 4223 7701
rect 2367 7663 2371 7671
rect 2380 7663 2384 7671
rect 2388 7663 2392 7671
rect 2396 7667 2400 7671
rect 2404 7663 2408 7671
rect 2417 7663 2421 7671
rect 2430 7663 2434 7671
rect 2438 7663 2442 7671
rect 2446 7663 2450 7671
rect 2454 7667 2458 7671
rect 2462 7663 2466 7671
rect 2475 7663 2479 7671
rect 2483 7663 2487 7671
rect 2491 7663 2495 7671
rect 2499 7663 2503 7671
rect 2512 7663 2516 7671
rect 2520 7663 2524 7671
rect 2528 7667 2532 7671
rect 2536 7663 2540 7671
rect 2549 7663 2553 7671
rect 2562 7663 2566 7671
rect 2570 7663 2574 7671
rect 2578 7663 2582 7671
rect 2586 7667 2590 7671
rect 2594 7663 2598 7671
rect 2607 7663 2611 7671
rect 2615 7663 2619 7671
rect 2623 7663 2627 7671
rect 2631 7663 2635 7671
rect 2644 7663 2648 7671
rect 2652 7663 2656 7671
rect 2660 7667 2664 7671
rect 2668 7663 2672 7671
rect 2681 7663 2685 7671
rect 2694 7663 2698 7671
rect 2702 7663 2706 7671
rect 2710 7663 2714 7671
rect 2718 7667 2722 7671
rect 2726 7663 2730 7671
rect 2739 7663 2743 7671
rect 2747 7663 2751 7671
rect 2755 7663 2759 7671
rect 3312 7663 3316 7671
rect 3325 7663 3329 7671
rect 3333 7663 3337 7671
rect 3341 7667 3345 7671
rect 3349 7663 3353 7671
rect 3362 7663 3366 7671
rect 3375 7663 3379 7671
rect 3383 7663 3387 7671
rect 3391 7663 3395 7671
rect 3399 7667 3403 7671
rect 3407 7663 3411 7671
rect 3420 7663 3424 7671
rect 3428 7663 3432 7671
rect 3436 7663 3440 7671
rect 3444 7663 3448 7671
rect 3457 7663 3461 7671
rect 3465 7663 3469 7671
rect 3473 7667 3477 7671
rect 3481 7663 3485 7671
rect 3494 7663 3498 7671
rect 3507 7663 3511 7671
rect 3515 7663 3519 7671
rect 3523 7663 3527 7671
rect 3531 7667 3535 7671
rect 3539 7663 3543 7671
rect 3552 7663 3556 7671
rect 3560 7663 3564 7671
rect 3568 7663 3572 7671
rect 3576 7663 3580 7671
rect 3589 7663 3593 7671
rect 3597 7663 3601 7671
rect 3605 7667 3609 7671
rect 3613 7663 3617 7671
rect 3626 7663 3630 7671
rect 3639 7663 3643 7671
rect 3647 7663 3651 7671
rect 3655 7663 3659 7671
rect 3663 7667 3667 7671
rect 3671 7663 3675 7671
rect 3684 7663 3688 7671
rect 3692 7663 3696 7671
rect 3700 7663 3704 7671
rect 3150 7607 3154 7615
rect 3163 7607 3167 7615
rect 3171 7607 3175 7615
rect 3179 7611 3183 7615
rect 3187 7607 3191 7615
rect 3200 7607 3204 7615
rect 3213 7607 3217 7615
rect 3221 7607 3225 7615
rect 3229 7607 3233 7615
rect 3237 7611 3241 7615
rect 3245 7607 3249 7615
rect 3258 7607 3262 7615
rect 3266 7607 3270 7615
rect 3274 7607 3278 7615
rect 4095 7607 4099 7615
rect 4108 7607 4112 7615
rect 4116 7607 4120 7615
rect 4124 7611 4128 7615
rect 4132 7607 4136 7615
rect 4145 7607 4149 7615
rect 4158 7607 4162 7615
rect 4166 7607 4170 7615
rect 4174 7607 4178 7615
rect 4182 7611 4186 7615
rect 4190 7607 4194 7615
rect 4203 7607 4207 7615
rect 4211 7607 4215 7615
rect 4219 7607 4223 7615
rect 2367 7577 2371 7585
rect 2380 7577 2384 7585
rect 2388 7577 2392 7585
rect 2396 7581 2400 7585
rect 2404 7577 2408 7585
rect 2417 7577 2421 7585
rect 2430 7577 2434 7585
rect 2438 7577 2442 7585
rect 2446 7577 2450 7585
rect 2454 7581 2458 7585
rect 2462 7577 2466 7585
rect 2475 7577 2479 7585
rect 2483 7577 2487 7585
rect 2491 7577 2495 7585
rect 2499 7577 2503 7585
rect 2512 7577 2516 7585
rect 2520 7577 2524 7585
rect 2528 7581 2532 7585
rect 2536 7577 2540 7585
rect 2549 7577 2553 7585
rect 2562 7577 2566 7585
rect 2570 7577 2574 7585
rect 2578 7577 2582 7585
rect 2586 7581 2590 7585
rect 2594 7577 2598 7585
rect 2607 7577 2611 7585
rect 2615 7577 2619 7585
rect 2623 7577 2627 7585
rect 2631 7577 2635 7585
rect 2644 7577 2648 7585
rect 2652 7577 2656 7585
rect 2660 7581 2664 7585
rect 2668 7577 2672 7585
rect 2681 7577 2685 7585
rect 2694 7577 2698 7585
rect 2702 7577 2706 7585
rect 2710 7577 2714 7585
rect 2718 7581 2722 7585
rect 2726 7577 2730 7585
rect 2739 7577 2743 7585
rect 2747 7577 2751 7585
rect 2755 7577 2759 7585
rect 3312 7577 3316 7585
rect 3325 7577 3329 7585
rect 3333 7577 3337 7585
rect 3341 7581 3345 7585
rect 3349 7577 3353 7585
rect 3362 7577 3366 7585
rect 3375 7577 3379 7585
rect 3383 7577 3387 7585
rect 3391 7577 3395 7585
rect 3399 7581 3403 7585
rect 3407 7577 3411 7585
rect 3420 7577 3424 7585
rect 3428 7577 3432 7585
rect 3436 7577 3440 7585
rect 3444 7577 3448 7585
rect 3457 7577 3461 7585
rect 3465 7577 3469 7585
rect 3473 7581 3477 7585
rect 3481 7577 3485 7585
rect 3494 7577 3498 7585
rect 3507 7577 3511 7585
rect 3515 7577 3519 7585
rect 3523 7577 3527 7585
rect 3531 7581 3535 7585
rect 3539 7577 3543 7585
rect 3552 7577 3556 7585
rect 3560 7577 3564 7585
rect 3568 7577 3572 7585
rect 3576 7577 3580 7585
rect 3589 7577 3593 7585
rect 3597 7577 3601 7585
rect 3605 7581 3609 7585
rect 3613 7577 3617 7585
rect 3626 7577 3630 7585
rect 3639 7577 3643 7585
rect 3647 7577 3651 7585
rect 3655 7577 3659 7585
rect 3663 7581 3667 7585
rect 3671 7577 3675 7585
rect 3684 7577 3688 7585
rect 3692 7577 3696 7585
rect 3700 7577 3704 7585
rect 2367 7437 2371 7445
rect 2380 7437 2384 7445
rect 2388 7437 2392 7445
rect 2396 7441 2400 7445
rect 2404 7437 2408 7445
rect 2417 7437 2421 7445
rect 2430 7437 2434 7445
rect 2438 7437 2442 7445
rect 2446 7437 2450 7445
rect 2454 7441 2458 7445
rect 2462 7437 2466 7445
rect 2475 7437 2479 7445
rect 2483 7437 2487 7445
rect 2491 7437 2495 7445
rect 2499 7437 2503 7445
rect 2512 7437 2516 7445
rect 2520 7437 2524 7445
rect 2528 7441 2532 7445
rect 2536 7437 2540 7445
rect 2549 7437 2553 7445
rect 2562 7437 2566 7445
rect 2570 7437 2574 7445
rect 2578 7437 2582 7445
rect 2586 7441 2590 7445
rect 2594 7437 2598 7445
rect 2607 7437 2611 7445
rect 2615 7437 2619 7445
rect 2623 7437 2627 7445
rect 2631 7437 2635 7445
rect 2644 7437 2648 7445
rect 2652 7437 2656 7445
rect 2660 7441 2664 7445
rect 2668 7437 2672 7445
rect 2681 7437 2685 7445
rect 2694 7437 2698 7445
rect 2702 7437 2706 7445
rect 2710 7437 2714 7445
rect 2718 7441 2722 7445
rect 2726 7437 2730 7445
rect 2739 7437 2743 7445
rect 2747 7437 2751 7445
rect 2755 7437 2759 7445
rect 3312 7437 3316 7445
rect 3325 7437 3329 7445
rect 3333 7437 3337 7445
rect 3341 7441 3345 7445
rect 3349 7437 3353 7445
rect 3362 7437 3366 7445
rect 3375 7437 3379 7445
rect 3383 7437 3387 7445
rect 3391 7437 3395 7445
rect 3399 7441 3403 7445
rect 3407 7437 3411 7445
rect 3420 7437 3424 7445
rect 3428 7437 3432 7445
rect 3436 7437 3440 7445
rect 3444 7437 3448 7445
rect 3457 7437 3461 7445
rect 3465 7437 3469 7445
rect 3473 7441 3477 7445
rect 3481 7437 3485 7445
rect 3494 7437 3498 7445
rect 3507 7437 3511 7445
rect 3515 7437 3519 7445
rect 3523 7437 3527 7445
rect 3531 7441 3535 7445
rect 3539 7437 3543 7445
rect 3552 7437 3556 7445
rect 3560 7437 3564 7445
rect 3568 7437 3572 7445
rect 3576 7437 3580 7445
rect 3589 7437 3593 7445
rect 3597 7437 3601 7445
rect 3605 7441 3609 7445
rect 3613 7437 3617 7445
rect 3626 7437 3630 7445
rect 3639 7437 3643 7445
rect 3647 7437 3651 7445
rect 3655 7437 3659 7445
rect 3663 7441 3667 7445
rect 3671 7437 3675 7445
rect 3684 7437 3688 7445
rect 3692 7437 3696 7445
rect 3700 7437 3704 7445
rect 4574 7928 4578 7945
rect 4574 7889 4578 7924
rect 4582 7889 4586 7945
rect 4590 7928 4594 7945
rect 4590 7889 4594 7924
rect 4598 7889 4602 7945
rect 4606 7928 4610 7945
rect 4606 7889 4610 7924
rect 4614 7889 4618 7945
rect 4622 7928 4626 7945
rect 4622 7889 4626 7924
rect 4637 7857 4641 7945
rect 4645 7928 4649 7936
rect 4645 7857 4649 7924
rect 4653 7857 4657 7945
rect 4661 7928 4665 7945
rect 4661 7857 4665 7924
rect 4680 7857 4684 7945
rect 4688 7928 4692 7936
rect 4688 7857 4692 7924
rect 4696 7857 4700 7945
rect 4704 7928 4708 7945
rect 4704 7857 4708 7924
rect 4721 7857 4725 7945
rect 4729 7928 4733 7936
rect 4729 7857 4733 7924
rect 4737 7857 4741 7945
rect 4745 7928 4749 7945
rect 4745 7857 4749 7924
<< psubstratepdiff >>
rect 1383 9965 1455 9967
rect 1383 9961 1385 9965
rect 1389 9961 1392 9965
rect 1396 9961 1397 9965
rect 1401 9961 1402 9965
rect 1406 9961 1407 9965
rect 1411 9961 1412 9965
rect 1416 9961 1417 9965
rect 1421 9961 1422 9965
rect 1426 9961 1427 9965
rect 1431 9961 1432 9965
rect 1436 9961 1437 9965
rect 1441 9961 1442 9965
rect 1446 9961 1449 9965
rect 1453 9961 1455 9965
rect 1383 9959 1455 9961
rect 1383 9958 1391 9959
rect 1383 9954 1385 9958
rect 1389 9954 1391 9958
rect 1383 9953 1391 9954
rect 1447 9958 1455 9959
rect 1447 9954 1449 9958
rect 1453 9954 1455 9958
rect 1447 9953 1455 9954
rect 1383 9949 1385 9953
rect 1389 9949 1391 9953
rect 1383 9948 1391 9949
rect 1383 9944 1385 9948
rect 1389 9944 1391 9948
rect 1383 9943 1391 9944
rect 1383 9939 1385 9943
rect 1389 9939 1391 9943
rect 1383 9938 1391 9939
rect 1383 9934 1385 9938
rect 1389 9934 1391 9938
rect 1383 9933 1391 9934
rect 1383 9929 1385 9933
rect 1389 9929 1391 9933
rect 1383 9928 1391 9929
rect 1383 9924 1385 9928
rect 1389 9924 1391 9928
rect 1383 9923 1391 9924
rect 1383 9919 1385 9923
rect 1389 9919 1391 9923
rect 1383 9918 1391 9919
rect 1383 9914 1385 9918
rect 1389 9914 1391 9918
rect 1383 9913 1391 9914
rect 1383 9909 1385 9913
rect 1389 9909 1391 9913
rect 1383 9908 1391 9909
rect 1383 9904 1385 9908
rect 1389 9904 1391 9908
rect 1383 9903 1391 9904
rect 1383 9899 1385 9903
rect 1389 9899 1391 9903
rect 1383 9898 1391 9899
rect 1383 9894 1385 9898
rect 1389 9894 1391 9898
rect 1383 9893 1391 9894
rect 1383 9889 1385 9893
rect 1389 9889 1391 9893
rect 1383 9888 1391 9889
rect 1383 9884 1385 9888
rect 1389 9884 1391 9888
rect 1383 9883 1391 9884
rect 1383 9879 1385 9883
rect 1389 9879 1391 9883
rect 1383 9878 1391 9879
rect 1383 9874 1385 9878
rect 1389 9874 1391 9878
rect 1383 9873 1391 9874
rect 1383 9869 1385 9873
rect 1389 9869 1391 9873
rect 1383 9868 1391 9869
rect 1383 9864 1385 9868
rect 1389 9864 1391 9868
rect 1447 9949 1449 9953
rect 1453 9949 1455 9953
rect 1447 9948 1455 9949
rect 1447 9944 1449 9948
rect 1453 9944 1455 9948
rect 1447 9943 1455 9944
rect 1447 9939 1449 9943
rect 1453 9939 1455 9943
rect 1447 9938 1455 9939
rect 1447 9934 1449 9938
rect 1453 9934 1455 9938
rect 1447 9933 1455 9934
rect 1447 9929 1449 9933
rect 1453 9929 1455 9933
rect 1447 9928 1455 9929
rect 1447 9924 1449 9928
rect 1453 9924 1455 9928
rect 1447 9923 1455 9924
rect 1447 9919 1449 9923
rect 1453 9919 1455 9923
rect 1447 9918 1455 9919
rect 1447 9914 1449 9918
rect 1453 9914 1455 9918
rect 1447 9913 1455 9914
rect 1447 9909 1449 9913
rect 1453 9909 1455 9913
rect 1447 9908 1455 9909
rect 1447 9904 1449 9908
rect 1453 9904 1455 9908
rect 1447 9903 1455 9904
rect 1447 9899 1449 9903
rect 1453 9899 1455 9903
rect 1447 9898 1455 9899
rect 1447 9894 1449 9898
rect 1453 9894 1455 9898
rect 1447 9893 1455 9894
rect 1447 9889 1449 9893
rect 1453 9889 1455 9893
rect 1447 9888 1455 9889
rect 1447 9884 1449 9888
rect 1453 9884 1455 9888
rect 1447 9883 1455 9884
rect 1447 9879 1449 9883
rect 1453 9879 1455 9883
rect 1447 9878 1455 9879
rect 1447 9874 1449 9878
rect 1453 9874 1455 9878
rect 1447 9873 1455 9874
rect 1447 9869 1449 9873
rect 1453 9869 1455 9873
rect 1447 9868 1455 9869
rect 1447 9864 1449 9868
rect 1453 9864 1455 9868
rect 1383 9863 1391 9864
rect 1383 9859 1385 9863
rect 1389 9859 1391 9863
rect 1383 9858 1391 9859
rect 1447 9863 1455 9864
rect 1447 9859 1449 9863
rect 1453 9859 1455 9863
rect 1447 9858 1455 9859
rect 1383 9856 1455 9858
rect 1383 9852 1385 9856
rect 1389 9852 1392 9856
rect 1396 9852 1397 9856
rect 1401 9852 1402 9856
rect 1406 9852 1407 9856
rect 1411 9852 1412 9856
rect 1416 9852 1417 9856
rect 1421 9852 1422 9856
rect 1426 9852 1427 9856
rect 1431 9852 1432 9856
rect 1436 9852 1437 9856
rect 1441 9852 1442 9856
rect 1446 9852 1449 9856
rect 1453 9852 1455 9856
rect 1383 9850 1455 9852
rect 1531 9978 1627 9979
rect 1531 9974 1532 9978
rect 1536 9974 1537 9978
rect 1541 9974 1542 9978
rect 1546 9974 1547 9978
rect 1551 9974 1552 9978
rect 1556 9974 1557 9978
rect 1561 9974 1562 9978
rect 1566 9974 1567 9978
rect 1571 9974 1572 9978
rect 1576 9974 1577 9978
rect 1581 9974 1582 9978
rect 1586 9974 1587 9978
rect 1591 9974 1592 9978
rect 1596 9974 1597 9978
rect 1601 9974 1602 9978
rect 1606 9974 1607 9978
rect 1611 9974 1612 9978
rect 1616 9974 1617 9978
rect 1621 9974 1622 9978
rect 1626 9974 1627 9978
rect 1531 9973 1627 9974
rect 1531 9969 1532 9973
rect 1536 9969 1537 9973
rect 1531 9968 1537 9969
rect 1531 9964 1532 9968
rect 1536 9964 1537 9968
rect 1621 9969 1622 9973
rect 1626 9969 1627 9973
rect 1621 9968 1627 9969
rect 1531 9963 1537 9964
rect 1531 9959 1532 9963
rect 1536 9959 1537 9963
rect 1531 9958 1537 9959
rect 1531 9954 1532 9958
rect 1536 9954 1537 9958
rect 1531 9953 1537 9954
rect 1531 9949 1532 9953
rect 1536 9949 1537 9953
rect 1531 9948 1537 9949
rect 1531 9944 1532 9948
rect 1536 9944 1537 9948
rect 1531 9943 1537 9944
rect 1531 9939 1532 9943
rect 1536 9939 1537 9943
rect 1531 9938 1537 9939
rect 1531 9934 1532 9938
rect 1536 9934 1537 9938
rect 1531 9933 1537 9934
rect 1531 9929 1532 9933
rect 1536 9929 1537 9933
rect 1531 9928 1537 9929
rect 1531 9924 1532 9928
rect 1536 9924 1537 9928
rect 1531 9923 1537 9924
rect 1531 9919 1532 9923
rect 1536 9919 1537 9923
rect 1531 9918 1537 9919
rect 1531 9914 1532 9918
rect 1536 9914 1537 9918
rect 1531 9913 1537 9914
rect 1531 9909 1532 9913
rect 1536 9909 1537 9913
rect 1531 9908 1537 9909
rect 1531 9904 1532 9908
rect 1536 9904 1537 9908
rect 1531 9903 1537 9904
rect 1531 9899 1532 9903
rect 1536 9899 1537 9903
rect 1531 9898 1537 9899
rect 1531 9894 1532 9898
rect 1536 9894 1537 9898
rect 1531 9893 1537 9894
rect 1531 9889 1532 9893
rect 1536 9889 1537 9893
rect 1531 9888 1537 9889
rect 1531 9884 1532 9888
rect 1536 9884 1537 9888
rect 1531 9883 1537 9884
rect 1531 9879 1532 9883
rect 1536 9879 1537 9883
rect 1531 9878 1537 9879
rect 1531 9874 1532 9878
rect 1536 9874 1537 9878
rect 1531 9873 1537 9874
rect 1531 9869 1532 9873
rect 1536 9869 1537 9873
rect 1531 9868 1537 9869
rect 1531 9864 1532 9868
rect 1536 9864 1537 9868
rect 1531 9863 1537 9864
rect 1531 9859 1532 9863
rect 1536 9859 1537 9863
rect 1531 9858 1537 9859
rect 1531 9854 1532 9858
rect 1536 9854 1537 9858
rect 1531 9853 1537 9854
rect 1531 9849 1532 9853
rect 1536 9849 1537 9853
rect 1621 9964 1622 9968
rect 1626 9964 1627 9968
rect 1621 9963 1627 9964
rect 1621 9959 1622 9963
rect 1626 9959 1627 9963
rect 1621 9958 1627 9959
rect 1621 9954 1622 9958
rect 1626 9954 1627 9958
rect 1621 9953 1627 9954
rect 1621 9949 1622 9953
rect 1626 9949 1627 9953
rect 1621 9948 1627 9949
rect 1621 9944 1622 9948
rect 1626 9944 1627 9948
rect 1621 9943 1627 9944
rect 1621 9939 1622 9943
rect 1626 9939 1627 9943
rect 1621 9938 1627 9939
rect 1621 9934 1622 9938
rect 1626 9934 1627 9938
rect 1621 9933 1627 9934
rect 1621 9929 1622 9933
rect 1626 9929 1627 9933
rect 1621 9928 1627 9929
rect 1621 9924 1622 9928
rect 1626 9924 1627 9928
rect 1621 9923 1627 9924
rect 1621 9919 1622 9923
rect 1626 9919 1627 9923
rect 1621 9918 1627 9919
rect 1621 9914 1622 9918
rect 1626 9914 1627 9918
rect 1621 9913 1627 9914
rect 1621 9909 1622 9913
rect 1626 9909 1627 9913
rect 1621 9908 1627 9909
rect 1621 9904 1622 9908
rect 1626 9904 1627 9908
rect 1621 9903 1627 9904
rect 1621 9899 1622 9903
rect 1626 9899 1627 9903
rect 1621 9898 1627 9899
rect 1621 9894 1622 9898
rect 1626 9894 1627 9898
rect 1621 9893 1627 9894
rect 1621 9889 1622 9893
rect 1626 9889 1627 9893
rect 1621 9888 1627 9889
rect 1621 9884 1622 9888
rect 1626 9884 1627 9888
rect 1621 9883 1627 9884
rect 1621 9879 1622 9883
rect 1626 9879 1627 9883
rect 1621 9878 1627 9879
rect 1621 9874 1622 9878
rect 1626 9874 1627 9878
rect 1621 9873 1627 9874
rect 1621 9869 1622 9873
rect 1626 9869 1627 9873
rect 1621 9868 1627 9869
rect 1621 9864 1622 9868
rect 1626 9864 1627 9868
rect 1621 9863 1627 9864
rect 1621 9859 1622 9863
rect 1626 9859 1627 9863
rect 1621 9858 1627 9859
rect 1621 9854 1622 9858
rect 1626 9854 1627 9858
rect 1621 9853 1627 9854
rect 1531 9848 1537 9849
rect 1531 9844 1532 9848
rect 1536 9844 1537 9848
rect 1621 9849 1622 9853
rect 1626 9849 1627 9853
rect 1621 9848 1627 9849
rect 1621 9844 1622 9848
rect 1626 9844 1627 9848
rect 1531 9843 1627 9844
rect 1531 9839 1532 9843
rect 1536 9839 1537 9843
rect 1541 9839 1542 9843
rect 1546 9839 1547 9843
rect 1551 9839 1552 9843
rect 1556 9839 1557 9843
rect 1561 9839 1562 9843
rect 1566 9839 1567 9843
rect 1571 9839 1572 9843
rect 1576 9839 1577 9843
rect 1581 9839 1582 9843
rect 1586 9839 1587 9843
rect 1591 9839 1592 9843
rect 1596 9839 1597 9843
rect 1601 9839 1602 9843
rect 1606 9839 1607 9843
rect 1611 9839 1612 9843
rect 1616 9839 1617 9843
rect 1621 9839 1622 9843
rect 1626 9839 1627 9843
rect 1531 9838 1627 9839
rect 1692 9965 1764 9967
rect 1692 9961 1694 9965
rect 1698 9961 1701 9965
rect 1705 9961 1706 9965
rect 1710 9961 1711 9965
rect 1715 9961 1716 9965
rect 1720 9961 1721 9965
rect 1725 9961 1726 9965
rect 1730 9961 1731 9965
rect 1735 9961 1736 9965
rect 1740 9961 1741 9965
rect 1745 9961 1746 9965
rect 1750 9961 1751 9965
rect 1755 9961 1758 9965
rect 1762 9961 1764 9965
rect 1692 9959 1764 9961
rect 1692 9958 1700 9959
rect 1692 9954 1694 9958
rect 1698 9954 1700 9958
rect 1692 9953 1700 9954
rect 1756 9958 1764 9959
rect 1756 9954 1758 9958
rect 1762 9954 1764 9958
rect 1756 9953 1764 9954
rect 1692 9949 1694 9953
rect 1698 9949 1700 9953
rect 1692 9948 1700 9949
rect 1692 9944 1694 9948
rect 1698 9944 1700 9948
rect 1692 9943 1700 9944
rect 1692 9939 1694 9943
rect 1698 9939 1700 9943
rect 1692 9938 1700 9939
rect 1692 9934 1694 9938
rect 1698 9934 1700 9938
rect 1692 9933 1700 9934
rect 1692 9929 1694 9933
rect 1698 9929 1700 9933
rect 1692 9928 1700 9929
rect 1692 9924 1694 9928
rect 1698 9924 1700 9928
rect 1692 9923 1700 9924
rect 1692 9919 1694 9923
rect 1698 9919 1700 9923
rect 1692 9918 1700 9919
rect 1692 9914 1694 9918
rect 1698 9914 1700 9918
rect 1692 9913 1700 9914
rect 1692 9909 1694 9913
rect 1698 9909 1700 9913
rect 1692 9908 1700 9909
rect 1692 9904 1694 9908
rect 1698 9904 1700 9908
rect 1692 9903 1700 9904
rect 1692 9899 1694 9903
rect 1698 9899 1700 9903
rect 1692 9898 1700 9899
rect 1692 9894 1694 9898
rect 1698 9894 1700 9898
rect 1692 9893 1700 9894
rect 1692 9889 1694 9893
rect 1698 9889 1700 9893
rect 1692 9888 1700 9889
rect 1692 9884 1694 9888
rect 1698 9884 1700 9888
rect 1692 9883 1700 9884
rect 1692 9879 1694 9883
rect 1698 9879 1700 9883
rect 1692 9878 1700 9879
rect 1692 9874 1694 9878
rect 1698 9874 1700 9878
rect 1692 9873 1700 9874
rect 1692 9869 1694 9873
rect 1698 9869 1700 9873
rect 1692 9868 1700 9869
rect 1692 9864 1694 9868
rect 1698 9864 1700 9868
rect 1756 9949 1758 9953
rect 1762 9949 1764 9953
rect 1756 9948 1764 9949
rect 1756 9944 1758 9948
rect 1762 9944 1764 9948
rect 1756 9943 1764 9944
rect 1756 9939 1758 9943
rect 1762 9939 1764 9943
rect 1756 9938 1764 9939
rect 1756 9934 1758 9938
rect 1762 9934 1764 9938
rect 1756 9933 1764 9934
rect 1756 9929 1758 9933
rect 1762 9929 1764 9933
rect 1756 9928 1764 9929
rect 1756 9924 1758 9928
rect 1762 9924 1764 9928
rect 1756 9923 1764 9924
rect 1756 9919 1758 9923
rect 1762 9919 1764 9923
rect 1756 9918 1764 9919
rect 1756 9914 1758 9918
rect 1762 9914 1764 9918
rect 1756 9913 1764 9914
rect 1756 9909 1758 9913
rect 1762 9909 1764 9913
rect 1756 9908 1764 9909
rect 1756 9904 1758 9908
rect 1762 9904 1764 9908
rect 1756 9903 1764 9904
rect 1756 9899 1758 9903
rect 1762 9899 1764 9903
rect 1756 9898 1764 9899
rect 1756 9894 1758 9898
rect 1762 9894 1764 9898
rect 1756 9893 1764 9894
rect 1756 9889 1758 9893
rect 1762 9889 1764 9893
rect 1756 9888 1764 9889
rect 1756 9884 1758 9888
rect 1762 9884 1764 9888
rect 1756 9883 1764 9884
rect 1756 9879 1758 9883
rect 1762 9879 1764 9883
rect 1756 9878 1764 9879
rect 1756 9874 1758 9878
rect 1762 9874 1764 9878
rect 1756 9873 1764 9874
rect 1756 9869 1758 9873
rect 1762 9869 1764 9873
rect 1756 9868 1764 9869
rect 1756 9864 1758 9868
rect 1762 9864 1764 9868
rect 1692 9863 1700 9864
rect 1692 9859 1694 9863
rect 1698 9859 1700 9863
rect 1692 9858 1700 9859
rect 1756 9863 1764 9864
rect 1756 9859 1758 9863
rect 1762 9859 1764 9863
rect 1756 9858 1764 9859
rect 1692 9856 1764 9858
rect 1692 9852 1694 9856
rect 1698 9852 1701 9856
rect 1705 9852 1706 9856
rect 1710 9852 1711 9856
rect 1715 9852 1716 9856
rect 1720 9852 1721 9856
rect 1725 9852 1726 9856
rect 1730 9852 1731 9856
rect 1735 9852 1736 9856
rect 1740 9852 1741 9856
rect 1745 9852 1746 9856
rect 1750 9852 1751 9856
rect 1755 9852 1758 9856
rect 1762 9852 1764 9856
rect 1692 9850 1764 9852
rect 1840 9978 1936 9979
rect 1840 9974 1841 9978
rect 1845 9974 1846 9978
rect 1850 9974 1851 9978
rect 1855 9974 1856 9978
rect 1860 9974 1861 9978
rect 1865 9974 1866 9978
rect 1870 9974 1871 9978
rect 1875 9974 1876 9978
rect 1880 9974 1881 9978
rect 1885 9974 1886 9978
rect 1890 9974 1891 9978
rect 1895 9974 1896 9978
rect 1900 9974 1901 9978
rect 1905 9974 1906 9978
rect 1910 9974 1911 9978
rect 1915 9974 1916 9978
rect 1920 9974 1921 9978
rect 1925 9974 1926 9978
rect 1930 9974 1931 9978
rect 1935 9974 1936 9978
rect 1840 9973 1936 9974
rect 1840 9969 1841 9973
rect 1845 9969 1846 9973
rect 1840 9968 1846 9969
rect 1840 9964 1841 9968
rect 1845 9964 1846 9968
rect 1930 9969 1931 9973
rect 1935 9969 1936 9973
rect 1930 9968 1936 9969
rect 1840 9963 1846 9964
rect 1840 9959 1841 9963
rect 1845 9959 1846 9963
rect 1840 9958 1846 9959
rect 1840 9954 1841 9958
rect 1845 9954 1846 9958
rect 1840 9953 1846 9954
rect 1840 9949 1841 9953
rect 1845 9949 1846 9953
rect 1840 9948 1846 9949
rect 1840 9944 1841 9948
rect 1845 9944 1846 9948
rect 1840 9943 1846 9944
rect 1840 9939 1841 9943
rect 1845 9939 1846 9943
rect 1840 9938 1846 9939
rect 1840 9934 1841 9938
rect 1845 9934 1846 9938
rect 1840 9933 1846 9934
rect 1840 9929 1841 9933
rect 1845 9929 1846 9933
rect 1840 9928 1846 9929
rect 1840 9924 1841 9928
rect 1845 9924 1846 9928
rect 1840 9923 1846 9924
rect 1840 9919 1841 9923
rect 1845 9919 1846 9923
rect 1840 9918 1846 9919
rect 1840 9914 1841 9918
rect 1845 9914 1846 9918
rect 1840 9913 1846 9914
rect 1840 9909 1841 9913
rect 1845 9909 1846 9913
rect 1840 9908 1846 9909
rect 1840 9904 1841 9908
rect 1845 9904 1846 9908
rect 1840 9903 1846 9904
rect 1840 9899 1841 9903
rect 1845 9899 1846 9903
rect 1840 9898 1846 9899
rect 1840 9894 1841 9898
rect 1845 9894 1846 9898
rect 1840 9893 1846 9894
rect 1840 9889 1841 9893
rect 1845 9889 1846 9893
rect 1840 9888 1846 9889
rect 1840 9884 1841 9888
rect 1845 9884 1846 9888
rect 1840 9883 1846 9884
rect 1840 9879 1841 9883
rect 1845 9879 1846 9883
rect 1840 9878 1846 9879
rect 1840 9874 1841 9878
rect 1845 9874 1846 9878
rect 1840 9873 1846 9874
rect 1840 9869 1841 9873
rect 1845 9869 1846 9873
rect 1840 9868 1846 9869
rect 1840 9864 1841 9868
rect 1845 9864 1846 9868
rect 1840 9863 1846 9864
rect 1840 9859 1841 9863
rect 1845 9859 1846 9863
rect 1840 9858 1846 9859
rect 1840 9854 1841 9858
rect 1845 9854 1846 9858
rect 1840 9853 1846 9854
rect 1840 9849 1841 9853
rect 1845 9849 1846 9853
rect 1930 9964 1931 9968
rect 1935 9964 1936 9968
rect 1930 9963 1936 9964
rect 1930 9959 1931 9963
rect 1935 9959 1936 9963
rect 1930 9958 1936 9959
rect 1930 9954 1931 9958
rect 1935 9954 1936 9958
rect 1930 9953 1936 9954
rect 1930 9949 1931 9953
rect 1935 9949 1936 9953
rect 1930 9948 1936 9949
rect 1930 9944 1931 9948
rect 1935 9944 1936 9948
rect 1930 9943 1936 9944
rect 1930 9939 1931 9943
rect 1935 9939 1936 9943
rect 1930 9938 1936 9939
rect 1930 9934 1931 9938
rect 1935 9934 1936 9938
rect 1930 9933 1936 9934
rect 1930 9929 1931 9933
rect 1935 9929 1936 9933
rect 1930 9928 1936 9929
rect 1930 9924 1931 9928
rect 1935 9924 1936 9928
rect 1930 9923 1936 9924
rect 1930 9919 1931 9923
rect 1935 9919 1936 9923
rect 1930 9918 1936 9919
rect 1930 9914 1931 9918
rect 1935 9914 1936 9918
rect 1930 9913 1936 9914
rect 1930 9909 1931 9913
rect 1935 9909 1936 9913
rect 1930 9908 1936 9909
rect 1930 9904 1931 9908
rect 1935 9904 1936 9908
rect 1930 9903 1936 9904
rect 1930 9899 1931 9903
rect 1935 9899 1936 9903
rect 1930 9898 1936 9899
rect 1930 9894 1931 9898
rect 1935 9894 1936 9898
rect 1930 9893 1936 9894
rect 1930 9889 1931 9893
rect 1935 9889 1936 9893
rect 1930 9888 1936 9889
rect 1930 9884 1931 9888
rect 1935 9884 1936 9888
rect 1930 9883 1936 9884
rect 1930 9879 1931 9883
rect 1935 9879 1936 9883
rect 1930 9878 1936 9879
rect 1930 9874 1931 9878
rect 1935 9874 1936 9878
rect 1930 9873 1936 9874
rect 1930 9869 1931 9873
rect 1935 9869 1936 9873
rect 1930 9868 1936 9869
rect 1930 9864 1931 9868
rect 1935 9864 1936 9868
rect 1930 9863 1936 9864
rect 1930 9859 1931 9863
rect 1935 9859 1936 9863
rect 1930 9858 1936 9859
rect 1930 9854 1931 9858
rect 1935 9854 1936 9858
rect 1930 9853 1936 9854
rect 1840 9848 1846 9849
rect 1840 9844 1841 9848
rect 1845 9844 1846 9848
rect 1930 9849 1931 9853
rect 1935 9849 1936 9853
rect 1930 9848 1936 9849
rect 1930 9844 1931 9848
rect 1935 9844 1936 9848
rect 1840 9843 1936 9844
rect 1840 9839 1841 9843
rect 1845 9839 1846 9843
rect 1850 9839 1851 9843
rect 1855 9839 1856 9843
rect 1860 9839 1861 9843
rect 1865 9839 1866 9843
rect 1870 9839 1871 9843
rect 1875 9839 1876 9843
rect 1880 9839 1881 9843
rect 1885 9839 1886 9843
rect 1890 9839 1891 9843
rect 1895 9839 1896 9843
rect 1900 9839 1901 9843
rect 1905 9839 1906 9843
rect 1910 9839 1911 9843
rect 1915 9839 1916 9843
rect 1920 9839 1921 9843
rect 1925 9839 1926 9843
rect 1930 9839 1931 9843
rect 1935 9839 1936 9843
rect 1840 9838 1936 9839
rect 2001 9965 2073 9967
rect 2001 9961 2003 9965
rect 2007 9961 2010 9965
rect 2014 9961 2015 9965
rect 2019 9961 2020 9965
rect 2024 9961 2025 9965
rect 2029 9961 2030 9965
rect 2034 9961 2035 9965
rect 2039 9961 2040 9965
rect 2044 9961 2045 9965
rect 2049 9961 2050 9965
rect 2054 9961 2055 9965
rect 2059 9961 2060 9965
rect 2064 9961 2067 9965
rect 2071 9961 2073 9965
rect 2001 9959 2073 9961
rect 2001 9958 2009 9959
rect 2001 9954 2003 9958
rect 2007 9954 2009 9958
rect 2001 9953 2009 9954
rect 2065 9958 2073 9959
rect 2065 9954 2067 9958
rect 2071 9954 2073 9958
rect 2065 9953 2073 9954
rect 2001 9949 2003 9953
rect 2007 9949 2009 9953
rect 2001 9948 2009 9949
rect 2001 9944 2003 9948
rect 2007 9944 2009 9948
rect 2001 9943 2009 9944
rect 2001 9939 2003 9943
rect 2007 9939 2009 9943
rect 2001 9938 2009 9939
rect 2001 9934 2003 9938
rect 2007 9934 2009 9938
rect 2001 9933 2009 9934
rect 2001 9929 2003 9933
rect 2007 9929 2009 9933
rect 2001 9928 2009 9929
rect 2001 9924 2003 9928
rect 2007 9924 2009 9928
rect 2001 9923 2009 9924
rect 2001 9919 2003 9923
rect 2007 9919 2009 9923
rect 2001 9918 2009 9919
rect 2001 9914 2003 9918
rect 2007 9914 2009 9918
rect 2001 9913 2009 9914
rect 2001 9909 2003 9913
rect 2007 9909 2009 9913
rect 2001 9908 2009 9909
rect 2001 9904 2003 9908
rect 2007 9904 2009 9908
rect 2001 9903 2009 9904
rect 2001 9899 2003 9903
rect 2007 9899 2009 9903
rect 2001 9898 2009 9899
rect 2001 9894 2003 9898
rect 2007 9894 2009 9898
rect 2001 9893 2009 9894
rect 2001 9889 2003 9893
rect 2007 9889 2009 9893
rect 2001 9888 2009 9889
rect 2001 9884 2003 9888
rect 2007 9884 2009 9888
rect 2001 9883 2009 9884
rect 2001 9879 2003 9883
rect 2007 9879 2009 9883
rect 2001 9878 2009 9879
rect 2001 9874 2003 9878
rect 2007 9874 2009 9878
rect 2001 9873 2009 9874
rect 2001 9869 2003 9873
rect 2007 9869 2009 9873
rect 2001 9868 2009 9869
rect 2001 9864 2003 9868
rect 2007 9864 2009 9868
rect 2065 9949 2067 9953
rect 2071 9949 2073 9953
rect 2065 9948 2073 9949
rect 2065 9944 2067 9948
rect 2071 9944 2073 9948
rect 2065 9943 2073 9944
rect 2065 9939 2067 9943
rect 2071 9939 2073 9943
rect 2065 9938 2073 9939
rect 2065 9934 2067 9938
rect 2071 9934 2073 9938
rect 2065 9933 2073 9934
rect 2065 9929 2067 9933
rect 2071 9929 2073 9933
rect 2065 9928 2073 9929
rect 2065 9924 2067 9928
rect 2071 9924 2073 9928
rect 2065 9923 2073 9924
rect 2065 9919 2067 9923
rect 2071 9919 2073 9923
rect 2065 9918 2073 9919
rect 2065 9914 2067 9918
rect 2071 9914 2073 9918
rect 2065 9913 2073 9914
rect 2065 9909 2067 9913
rect 2071 9909 2073 9913
rect 2065 9908 2073 9909
rect 2065 9904 2067 9908
rect 2071 9904 2073 9908
rect 2065 9903 2073 9904
rect 2065 9899 2067 9903
rect 2071 9899 2073 9903
rect 2065 9898 2073 9899
rect 2065 9894 2067 9898
rect 2071 9894 2073 9898
rect 2065 9893 2073 9894
rect 2065 9889 2067 9893
rect 2071 9889 2073 9893
rect 2065 9888 2073 9889
rect 2065 9884 2067 9888
rect 2071 9884 2073 9888
rect 2065 9883 2073 9884
rect 2065 9879 2067 9883
rect 2071 9879 2073 9883
rect 2065 9878 2073 9879
rect 2065 9874 2067 9878
rect 2071 9874 2073 9878
rect 2065 9873 2073 9874
rect 2065 9869 2067 9873
rect 2071 9869 2073 9873
rect 2065 9868 2073 9869
rect 2065 9864 2067 9868
rect 2071 9864 2073 9868
rect 2001 9863 2009 9864
rect 2001 9859 2003 9863
rect 2007 9859 2009 9863
rect 2001 9858 2009 9859
rect 2065 9863 2073 9864
rect 2065 9859 2067 9863
rect 2071 9859 2073 9863
rect 2065 9858 2073 9859
rect 2001 9856 2073 9858
rect 2001 9852 2003 9856
rect 2007 9852 2010 9856
rect 2014 9852 2015 9856
rect 2019 9852 2020 9856
rect 2024 9852 2025 9856
rect 2029 9852 2030 9856
rect 2034 9852 2035 9856
rect 2039 9852 2040 9856
rect 2044 9852 2045 9856
rect 2049 9852 2050 9856
rect 2054 9852 2055 9856
rect 2059 9852 2060 9856
rect 2064 9852 2067 9856
rect 2071 9852 2073 9856
rect 2001 9850 2073 9852
rect 2149 9978 2245 9979
rect 2149 9974 2150 9978
rect 2154 9974 2155 9978
rect 2159 9974 2160 9978
rect 2164 9974 2165 9978
rect 2169 9974 2170 9978
rect 2174 9974 2175 9978
rect 2179 9974 2180 9978
rect 2184 9974 2185 9978
rect 2189 9974 2190 9978
rect 2194 9974 2195 9978
rect 2199 9974 2200 9978
rect 2204 9974 2205 9978
rect 2209 9974 2210 9978
rect 2214 9974 2215 9978
rect 2219 9974 2220 9978
rect 2224 9974 2225 9978
rect 2229 9974 2230 9978
rect 2234 9974 2235 9978
rect 2239 9974 2240 9978
rect 2244 9974 2245 9978
rect 2149 9973 2245 9974
rect 2149 9969 2150 9973
rect 2154 9969 2155 9973
rect 2149 9968 2155 9969
rect 2149 9964 2150 9968
rect 2154 9964 2155 9968
rect 2239 9969 2240 9973
rect 2244 9969 2245 9973
rect 2239 9968 2245 9969
rect 2149 9963 2155 9964
rect 2149 9959 2150 9963
rect 2154 9959 2155 9963
rect 2149 9958 2155 9959
rect 2149 9954 2150 9958
rect 2154 9954 2155 9958
rect 2149 9953 2155 9954
rect 2149 9949 2150 9953
rect 2154 9949 2155 9953
rect 2149 9948 2155 9949
rect 2149 9944 2150 9948
rect 2154 9944 2155 9948
rect 2149 9943 2155 9944
rect 2149 9939 2150 9943
rect 2154 9939 2155 9943
rect 2149 9938 2155 9939
rect 2149 9934 2150 9938
rect 2154 9934 2155 9938
rect 2149 9933 2155 9934
rect 2149 9929 2150 9933
rect 2154 9929 2155 9933
rect 2149 9928 2155 9929
rect 2149 9924 2150 9928
rect 2154 9924 2155 9928
rect 2149 9923 2155 9924
rect 2149 9919 2150 9923
rect 2154 9919 2155 9923
rect 2149 9918 2155 9919
rect 2149 9914 2150 9918
rect 2154 9914 2155 9918
rect 2149 9913 2155 9914
rect 2149 9909 2150 9913
rect 2154 9909 2155 9913
rect 2149 9908 2155 9909
rect 2149 9904 2150 9908
rect 2154 9904 2155 9908
rect 2149 9903 2155 9904
rect 2149 9899 2150 9903
rect 2154 9899 2155 9903
rect 2149 9898 2155 9899
rect 2149 9894 2150 9898
rect 2154 9894 2155 9898
rect 2149 9893 2155 9894
rect 2149 9889 2150 9893
rect 2154 9889 2155 9893
rect 2149 9888 2155 9889
rect 2149 9884 2150 9888
rect 2154 9884 2155 9888
rect 2149 9883 2155 9884
rect 2149 9879 2150 9883
rect 2154 9879 2155 9883
rect 2149 9878 2155 9879
rect 2149 9874 2150 9878
rect 2154 9874 2155 9878
rect 2149 9873 2155 9874
rect 2149 9869 2150 9873
rect 2154 9869 2155 9873
rect 2149 9868 2155 9869
rect 2149 9864 2150 9868
rect 2154 9864 2155 9868
rect 2149 9863 2155 9864
rect 2149 9859 2150 9863
rect 2154 9859 2155 9863
rect 2149 9858 2155 9859
rect 2149 9854 2150 9858
rect 2154 9854 2155 9858
rect 2149 9853 2155 9854
rect 2149 9849 2150 9853
rect 2154 9849 2155 9853
rect 2239 9964 2240 9968
rect 2244 9964 2245 9968
rect 2239 9963 2245 9964
rect 2239 9959 2240 9963
rect 2244 9959 2245 9963
rect 2239 9958 2245 9959
rect 2239 9954 2240 9958
rect 2244 9954 2245 9958
rect 2239 9953 2245 9954
rect 2239 9949 2240 9953
rect 2244 9949 2245 9953
rect 2239 9948 2245 9949
rect 2239 9944 2240 9948
rect 2244 9944 2245 9948
rect 2239 9943 2245 9944
rect 2239 9939 2240 9943
rect 2244 9939 2245 9943
rect 2239 9938 2245 9939
rect 2239 9934 2240 9938
rect 2244 9934 2245 9938
rect 2239 9933 2245 9934
rect 2239 9929 2240 9933
rect 2244 9929 2245 9933
rect 2239 9928 2245 9929
rect 2239 9924 2240 9928
rect 2244 9924 2245 9928
rect 2239 9923 2245 9924
rect 2239 9919 2240 9923
rect 2244 9919 2245 9923
rect 2239 9918 2245 9919
rect 2239 9914 2240 9918
rect 2244 9914 2245 9918
rect 2239 9913 2245 9914
rect 2239 9909 2240 9913
rect 2244 9909 2245 9913
rect 2239 9908 2245 9909
rect 2239 9904 2240 9908
rect 2244 9904 2245 9908
rect 2239 9903 2245 9904
rect 2239 9899 2240 9903
rect 2244 9899 2245 9903
rect 2239 9898 2245 9899
rect 2239 9894 2240 9898
rect 2244 9894 2245 9898
rect 2239 9893 2245 9894
rect 2239 9889 2240 9893
rect 2244 9889 2245 9893
rect 2239 9888 2245 9889
rect 2239 9884 2240 9888
rect 2244 9884 2245 9888
rect 2239 9883 2245 9884
rect 2239 9879 2240 9883
rect 2244 9879 2245 9883
rect 2239 9878 2245 9879
rect 2239 9874 2240 9878
rect 2244 9874 2245 9878
rect 2239 9873 2245 9874
rect 2239 9869 2240 9873
rect 2244 9869 2245 9873
rect 2239 9868 2245 9869
rect 2239 9864 2240 9868
rect 2244 9864 2245 9868
rect 2239 9863 2245 9864
rect 2239 9859 2240 9863
rect 2244 9859 2245 9863
rect 2239 9858 2245 9859
rect 2239 9854 2240 9858
rect 2244 9854 2245 9858
rect 2239 9853 2245 9854
rect 2149 9848 2155 9849
rect 2149 9844 2150 9848
rect 2154 9844 2155 9848
rect 2239 9849 2240 9853
rect 2244 9849 2245 9853
rect 2239 9848 2245 9849
rect 2239 9844 2240 9848
rect 2244 9844 2245 9848
rect 2149 9843 2245 9844
rect 2149 9839 2150 9843
rect 2154 9839 2155 9843
rect 2159 9839 2160 9843
rect 2164 9839 2165 9843
rect 2169 9839 2170 9843
rect 2174 9839 2175 9843
rect 2179 9839 2180 9843
rect 2184 9839 2185 9843
rect 2189 9839 2190 9843
rect 2194 9839 2195 9843
rect 2199 9839 2200 9843
rect 2204 9839 2205 9843
rect 2209 9839 2210 9843
rect 2214 9839 2215 9843
rect 2219 9839 2220 9843
rect 2224 9839 2225 9843
rect 2229 9839 2230 9843
rect 2234 9839 2235 9843
rect 2239 9839 2240 9843
rect 2244 9839 2245 9843
rect 2149 9838 2245 9839
rect 2310 9965 2382 9967
rect 2310 9961 2312 9965
rect 2316 9961 2319 9965
rect 2323 9961 2324 9965
rect 2328 9961 2329 9965
rect 2333 9961 2334 9965
rect 2338 9961 2339 9965
rect 2343 9961 2344 9965
rect 2348 9961 2349 9965
rect 2353 9961 2354 9965
rect 2358 9961 2359 9965
rect 2363 9961 2364 9965
rect 2368 9961 2369 9965
rect 2373 9961 2376 9965
rect 2380 9961 2382 9965
rect 2310 9959 2382 9961
rect 2310 9958 2318 9959
rect 2310 9954 2312 9958
rect 2316 9954 2318 9958
rect 2310 9953 2318 9954
rect 2374 9958 2382 9959
rect 2374 9954 2376 9958
rect 2380 9954 2382 9958
rect 2374 9953 2382 9954
rect 2310 9949 2312 9953
rect 2316 9949 2318 9953
rect 2310 9948 2318 9949
rect 2310 9944 2312 9948
rect 2316 9944 2318 9948
rect 2310 9943 2318 9944
rect 2310 9939 2312 9943
rect 2316 9939 2318 9943
rect 2310 9938 2318 9939
rect 2310 9934 2312 9938
rect 2316 9934 2318 9938
rect 2310 9933 2318 9934
rect 2310 9929 2312 9933
rect 2316 9929 2318 9933
rect 2310 9928 2318 9929
rect 2310 9924 2312 9928
rect 2316 9924 2318 9928
rect 2310 9923 2318 9924
rect 2310 9919 2312 9923
rect 2316 9919 2318 9923
rect 2310 9918 2318 9919
rect 2310 9914 2312 9918
rect 2316 9914 2318 9918
rect 2310 9913 2318 9914
rect 2310 9909 2312 9913
rect 2316 9909 2318 9913
rect 2310 9908 2318 9909
rect 2310 9904 2312 9908
rect 2316 9904 2318 9908
rect 2310 9903 2318 9904
rect 2310 9899 2312 9903
rect 2316 9899 2318 9903
rect 2310 9898 2318 9899
rect 2310 9894 2312 9898
rect 2316 9894 2318 9898
rect 2310 9893 2318 9894
rect 2310 9889 2312 9893
rect 2316 9889 2318 9893
rect 2310 9888 2318 9889
rect 2310 9884 2312 9888
rect 2316 9884 2318 9888
rect 2310 9883 2318 9884
rect 2310 9879 2312 9883
rect 2316 9879 2318 9883
rect 2310 9878 2318 9879
rect 2310 9874 2312 9878
rect 2316 9874 2318 9878
rect 2310 9873 2318 9874
rect 2310 9869 2312 9873
rect 2316 9869 2318 9873
rect 2310 9868 2318 9869
rect 2310 9864 2312 9868
rect 2316 9864 2318 9868
rect 2374 9949 2376 9953
rect 2380 9949 2382 9953
rect 2374 9948 2382 9949
rect 2374 9944 2376 9948
rect 2380 9944 2382 9948
rect 2374 9943 2382 9944
rect 2374 9939 2376 9943
rect 2380 9939 2382 9943
rect 2374 9938 2382 9939
rect 2374 9934 2376 9938
rect 2380 9934 2382 9938
rect 2374 9933 2382 9934
rect 2374 9929 2376 9933
rect 2380 9929 2382 9933
rect 2374 9928 2382 9929
rect 2374 9924 2376 9928
rect 2380 9924 2382 9928
rect 2374 9923 2382 9924
rect 2374 9919 2376 9923
rect 2380 9919 2382 9923
rect 2374 9918 2382 9919
rect 2374 9914 2376 9918
rect 2380 9914 2382 9918
rect 2374 9913 2382 9914
rect 2374 9909 2376 9913
rect 2380 9909 2382 9913
rect 2374 9908 2382 9909
rect 2374 9904 2376 9908
rect 2380 9904 2382 9908
rect 2374 9903 2382 9904
rect 2374 9899 2376 9903
rect 2380 9899 2382 9903
rect 2374 9898 2382 9899
rect 2374 9894 2376 9898
rect 2380 9894 2382 9898
rect 2374 9893 2382 9894
rect 2374 9889 2376 9893
rect 2380 9889 2382 9893
rect 2374 9888 2382 9889
rect 2374 9884 2376 9888
rect 2380 9884 2382 9888
rect 2374 9883 2382 9884
rect 2374 9879 2376 9883
rect 2380 9879 2382 9883
rect 2374 9878 2382 9879
rect 2374 9874 2376 9878
rect 2380 9874 2382 9878
rect 2374 9873 2382 9874
rect 2374 9869 2376 9873
rect 2380 9869 2382 9873
rect 2374 9868 2382 9869
rect 2374 9864 2376 9868
rect 2380 9864 2382 9868
rect 2310 9863 2318 9864
rect 2310 9859 2312 9863
rect 2316 9859 2318 9863
rect 2310 9858 2318 9859
rect 2374 9863 2382 9864
rect 2374 9859 2376 9863
rect 2380 9859 2382 9863
rect 2374 9858 2382 9859
rect 2310 9856 2382 9858
rect 2310 9852 2312 9856
rect 2316 9852 2319 9856
rect 2323 9852 2324 9856
rect 2328 9852 2329 9856
rect 2333 9852 2334 9856
rect 2338 9852 2339 9856
rect 2343 9852 2344 9856
rect 2348 9852 2349 9856
rect 2353 9852 2354 9856
rect 2358 9852 2359 9856
rect 2363 9852 2364 9856
rect 2368 9852 2369 9856
rect 2373 9852 2376 9856
rect 2380 9852 2382 9856
rect 2310 9850 2382 9852
rect 2458 9978 2554 9979
rect 2458 9974 2459 9978
rect 2463 9974 2464 9978
rect 2468 9974 2469 9978
rect 2473 9974 2474 9978
rect 2478 9974 2479 9978
rect 2483 9974 2484 9978
rect 2488 9974 2489 9978
rect 2493 9974 2494 9978
rect 2498 9974 2499 9978
rect 2503 9974 2504 9978
rect 2508 9974 2509 9978
rect 2513 9974 2514 9978
rect 2518 9974 2519 9978
rect 2523 9974 2524 9978
rect 2528 9974 2529 9978
rect 2533 9974 2534 9978
rect 2538 9974 2539 9978
rect 2543 9974 2544 9978
rect 2548 9974 2549 9978
rect 2553 9974 2554 9978
rect 2458 9973 2554 9974
rect 2458 9969 2459 9973
rect 2463 9969 2464 9973
rect 2458 9968 2464 9969
rect 2458 9964 2459 9968
rect 2463 9964 2464 9968
rect 2548 9969 2549 9973
rect 2553 9969 2554 9973
rect 2548 9968 2554 9969
rect 2458 9963 2464 9964
rect 2458 9959 2459 9963
rect 2463 9959 2464 9963
rect 2458 9958 2464 9959
rect 2458 9954 2459 9958
rect 2463 9954 2464 9958
rect 2458 9953 2464 9954
rect 2458 9949 2459 9953
rect 2463 9949 2464 9953
rect 2458 9948 2464 9949
rect 2458 9944 2459 9948
rect 2463 9944 2464 9948
rect 2458 9943 2464 9944
rect 2458 9939 2459 9943
rect 2463 9939 2464 9943
rect 2458 9938 2464 9939
rect 2458 9934 2459 9938
rect 2463 9934 2464 9938
rect 2458 9933 2464 9934
rect 2458 9929 2459 9933
rect 2463 9929 2464 9933
rect 2458 9928 2464 9929
rect 2458 9924 2459 9928
rect 2463 9924 2464 9928
rect 2458 9923 2464 9924
rect 2458 9919 2459 9923
rect 2463 9919 2464 9923
rect 2458 9918 2464 9919
rect 2458 9914 2459 9918
rect 2463 9914 2464 9918
rect 2458 9913 2464 9914
rect 2458 9909 2459 9913
rect 2463 9909 2464 9913
rect 2458 9908 2464 9909
rect 2458 9904 2459 9908
rect 2463 9904 2464 9908
rect 2458 9903 2464 9904
rect 2458 9899 2459 9903
rect 2463 9899 2464 9903
rect 2458 9898 2464 9899
rect 2458 9894 2459 9898
rect 2463 9894 2464 9898
rect 2458 9893 2464 9894
rect 2458 9889 2459 9893
rect 2463 9889 2464 9893
rect 2458 9888 2464 9889
rect 2458 9884 2459 9888
rect 2463 9884 2464 9888
rect 2458 9883 2464 9884
rect 2458 9879 2459 9883
rect 2463 9879 2464 9883
rect 2458 9878 2464 9879
rect 2458 9874 2459 9878
rect 2463 9874 2464 9878
rect 2458 9873 2464 9874
rect 2458 9869 2459 9873
rect 2463 9869 2464 9873
rect 2458 9868 2464 9869
rect 2458 9864 2459 9868
rect 2463 9864 2464 9868
rect 2458 9863 2464 9864
rect 2458 9859 2459 9863
rect 2463 9859 2464 9863
rect 2458 9858 2464 9859
rect 2458 9854 2459 9858
rect 2463 9854 2464 9858
rect 2458 9853 2464 9854
rect 2458 9849 2459 9853
rect 2463 9849 2464 9853
rect 2548 9964 2549 9968
rect 2553 9964 2554 9968
rect 2548 9963 2554 9964
rect 2548 9959 2549 9963
rect 2553 9959 2554 9963
rect 2548 9958 2554 9959
rect 2548 9954 2549 9958
rect 2553 9954 2554 9958
rect 2548 9953 2554 9954
rect 2548 9949 2549 9953
rect 2553 9949 2554 9953
rect 2548 9948 2554 9949
rect 2548 9944 2549 9948
rect 2553 9944 2554 9948
rect 2548 9943 2554 9944
rect 2548 9939 2549 9943
rect 2553 9939 2554 9943
rect 2548 9938 2554 9939
rect 2548 9934 2549 9938
rect 2553 9934 2554 9938
rect 2548 9933 2554 9934
rect 2548 9929 2549 9933
rect 2553 9929 2554 9933
rect 2548 9928 2554 9929
rect 2548 9924 2549 9928
rect 2553 9924 2554 9928
rect 2548 9923 2554 9924
rect 2548 9919 2549 9923
rect 2553 9919 2554 9923
rect 2548 9918 2554 9919
rect 2548 9914 2549 9918
rect 2553 9914 2554 9918
rect 2548 9913 2554 9914
rect 2548 9909 2549 9913
rect 2553 9909 2554 9913
rect 2548 9908 2554 9909
rect 2548 9904 2549 9908
rect 2553 9904 2554 9908
rect 2548 9903 2554 9904
rect 2548 9899 2549 9903
rect 2553 9899 2554 9903
rect 2548 9898 2554 9899
rect 2548 9894 2549 9898
rect 2553 9894 2554 9898
rect 2548 9893 2554 9894
rect 2548 9889 2549 9893
rect 2553 9889 2554 9893
rect 2548 9888 2554 9889
rect 2548 9884 2549 9888
rect 2553 9884 2554 9888
rect 2548 9883 2554 9884
rect 2548 9879 2549 9883
rect 2553 9879 2554 9883
rect 2548 9878 2554 9879
rect 2548 9874 2549 9878
rect 2553 9874 2554 9878
rect 2548 9873 2554 9874
rect 2548 9869 2549 9873
rect 2553 9869 2554 9873
rect 2548 9868 2554 9869
rect 2548 9864 2549 9868
rect 2553 9864 2554 9868
rect 2548 9863 2554 9864
rect 2548 9859 2549 9863
rect 2553 9859 2554 9863
rect 2548 9858 2554 9859
rect 2548 9854 2549 9858
rect 2553 9854 2554 9858
rect 2548 9853 2554 9854
rect 2458 9848 2464 9849
rect 2458 9844 2459 9848
rect 2463 9844 2464 9848
rect 2548 9849 2549 9853
rect 2553 9849 2554 9853
rect 2548 9848 2554 9849
rect 2548 9844 2549 9848
rect 2553 9844 2554 9848
rect 2458 9843 2554 9844
rect 2458 9839 2459 9843
rect 2463 9839 2464 9843
rect 2468 9839 2469 9843
rect 2473 9839 2474 9843
rect 2478 9839 2479 9843
rect 2483 9839 2484 9843
rect 2488 9839 2489 9843
rect 2493 9839 2494 9843
rect 2498 9839 2499 9843
rect 2503 9839 2504 9843
rect 2508 9839 2509 9843
rect 2513 9839 2514 9843
rect 2518 9839 2519 9843
rect 2523 9839 2524 9843
rect 2528 9839 2529 9843
rect 2533 9839 2534 9843
rect 2538 9839 2539 9843
rect 2543 9839 2544 9843
rect 2548 9839 2549 9843
rect 2553 9839 2554 9843
rect 2458 9838 2554 9839
rect 2619 9965 2691 9967
rect 2619 9961 2621 9965
rect 2625 9961 2628 9965
rect 2632 9961 2633 9965
rect 2637 9961 2638 9965
rect 2642 9961 2643 9965
rect 2647 9961 2648 9965
rect 2652 9961 2653 9965
rect 2657 9961 2658 9965
rect 2662 9961 2663 9965
rect 2667 9961 2668 9965
rect 2672 9961 2673 9965
rect 2677 9961 2678 9965
rect 2682 9961 2685 9965
rect 2689 9961 2691 9965
rect 2619 9959 2691 9961
rect 2619 9958 2627 9959
rect 2619 9954 2621 9958
rect 2625 9954 2627 9958
rect 2619 9953 2627 9954
rect 2683 9958 2691 9959
rect 2683 9954 2685 9958
rect 2689 9954 2691 9958
rect 2683 9953 2691 9954
rect 2619 9949 2621 9953
rect 2625 9949 2627 9953
rect 2619 9948 2627 9949
rect 2619 9944 2621 9948
rect 2625 9944 2627 9948
rect 2619 9943 2627 9944
rect 2619 9939 2621 9943
rect 2625 9939 2627 9943
rect 2619 9938 2627 9939
rect 2619 9934 2621 9938
rect 2625 9934 2627 9938
rect 2619 9933 2627 9934
rect 2619 9929 2621 9933
rect 2625 9929 2627 9933
rect 2619 9928 2627 9929
rect 2619 9924 2621 9928
rect 2625 9924 2627 9928
rect 2619 9923 2627 9924
rect 2619 9919 2621 9923
rect 2625 9919 2627 9923
rect 2619 9918 2627 9919
rect 2619 9914 2621 9918
rect 2625 9914 2627 9918
rect 2619 9913 2627 9914
rect 2619 9909 2621 9913
rect 2625 9909 2627 9913
rect 2619 9908 2627 9909
rect 2619 9904 2621 9908
rect 2625 9904 2627 9908
rect 2619 9903 2627 9904
rect 2619 9899 2621 9903
rect 2625 9899 2627 9903
rect 2619 9898 2627 9899
rect 2619 9894 2621 9898
rect 2625 9894 2627 9898
rect 2619 9893 2627 9894
rect 2619 9889 2621 9893
rect 2625 9889 2627 9893
rect 2619 9888 2627 9889
rect 2619 9884 2621 9888
rect 2625 9884 2627 9888
rect 2619 9883 2627 9884
rect 2619 9879 2621 9883
rect 2625 9879 2627 9883
rect 2619 9878 2627 9879
rect 2619 9874 2621 9878
rect 2625 9874 2627 9878
rect 2619 9873 2627 9874
rect 2619 9869 2621 9873
rect 2625 9869 2627 9873
rect 2619 9868 2627 9869
rect 2619 9864 2621 9868
rect 2625 9864 2627 9868
rect 2683 9949 2685 9953
rect 2689 9949 2691 9953
rect 2683 9948 2691 9949
rect 2683 9944 2685 9948
rect 2689 9944 2691 9948
rect 2683 9943 2691 9944
rect 2683 9939 2685 9943
rect 2689 9939 2691 9943
rect 2683 9938 2691 9939
rect 2683 9934 2685 9938
rect 2689 9934 2691 9938
rect 2683 9933 2691 9934
rect 2683 9929 2685 9933
rect 2689 9929 2691 9933
rect 2683 9928 2691 9929
rect 2683 9924 2685 9928
rect 2689 9924 2691 9928
rect 2683 9923 2691 9924
rect 2683 9919 2685 9923
rect 2689 9919 2691 9923
rect 2683 9918 2691 9919
rect 2683 9914 2685 9918
rect 2689 9914 2691 9918
rect 2683 9913 2691 9914
rect 2683 9909 2685 9913
rect 2689 9909 2691 9913
rect 2683 9908 2691 9909
rect 2683 9904 2685 9908
rect 2689 9904 2691 9908
rect 2683 9903 2691 9904
rect 2683 9899 2685 9903
rect 2689 9899 2691 9903
rect 2683 9898 2691 9899
rect 2683 9894 2685 9898
rect 2689 9894 2691 9898
rect 2683 9893 2691 9894
rect 2683 9889 2685 9893
rect 2689 9889 2691 9893
rect 2683 9888 2691 9889
rect 2683 9884 2685 9888
rect 2689 9884 2691 9888
rect 2683 9883 2691 9884
rect 2683 9879 2685 9883
rect 2689 9879 2691 9883
rect 2683 9878 2691 9879
rect 2683 9874 2685 9878
rect 2689 9874 2691 9878
rect 2683 9873 2691 9874
rect 2683 9869 2685 9873
rect 2689 9869 2691 9873
rect 2683 9868 2691 9869
rect 2683 9864 2685 9868
rect 2689 9864 2691 9868
rect 2619 9863 2627 9864
rect 2619 9859 2621 9863
rect 2625 9859 2627 9863
rect 2619 9858 2627 9859
rect 2683 9863 2691 9864
rect 2683 9859 2685 9863
rect 2689 9859 2691 9863
rect 2683 9858 2691 9859
rect 2619 9856 2691 9858
rect 2619 9852 2621 9856
rect 2625 9852 2628 9856
rect 2632 9852 2633 9856
rect 2637 9852 2638 9856
rect 2642 9852 2643 9856
rect 2647 9852 2648 9856
rect 2652 9852 2653 9856
rect 2657 9852 2658 9856
rect 2662 9852 2663 9856
rect 2667 9852 2668 9856
rect 2672 9852 2673 9856
rect 2677 9852 2678 9856
rect 2682 9852 2685 9856
rect 2689 9852 2691 9856
rect 2619 9850 2691 9852
rect 2767 9978 2863 9979
rect 2767 9974 2768 9978
rect 2772 9974 2773 9978
rect 2777 9974 2778 9978
rect 2782 9974 2783 9978
rect 2787 9974 2788 9978
rect 2792 9974 2793 9978
rect 2797 9974 2798 9978
rect 2802 9974 2803 9978
rect 2807 9974 2808 9978
rect 2812 9974 2813 9978
rect 2817 9974 2818 9978
rect 2822 9974 2823 9978
rect 2827 9974 2828 9978
rect 2832 9974 2833 9978
rect 2837 9974 2838 9978
rect 2842 9974 2843 9978
rect 2847 9974 2848 9978
rect 2852 9974 2853 9978
rect 2857 9974 2858 9978
rect 2862 9974 2863 9978
rect 2767 9973 2863 9974
rect 2767 9969 2768 9973
rect 2772 9969 2773 9973
rect 2767 9968 2773 9969
rect 2767 9964 2768 9968
rect 2772 9964 2773 9968
rect 2857 9969 2858 9973
rect 2862 9969 2863 9973
rect 2857 9968 2863 9969
rect 2767 9963 2773 9964
rect 2767 9959 2768 9963
rect 2772 9959 2773 9963
rect 2767 9958 2773 9959
rect 2767 9954 2768 9958
rect 2772 9954 2773 9958
rect 2767 9953 2773 9954
rect 2767 9949 2768 9953
rect 2772 9949 2773 9953
rect 2767 9948 2773 9949
rect 2767 9944 2768 9948
rect 2772 9944 2773 9948
rect 2767 9943 2773 9944
rect 2767 9939 2768 9943
rect 2772 9939 2773 9943
rect 2767 9938 2773 9939
rect 2767 9934 2768 9938
rect 2772 9934 2773 9938
rect 2767 9933 2773 9934
rect 2767 9929 2768 9933
rect 2772 9929 2773 9933
rect 2767 9928 2773 9929
rect 2767 9924 2768 9928
rect 2772 9924 2773 9928
rect 2767 9923 2773 9924
rect 2767 9919 2768 9923
rect 2772 9919 2773 9923
rect 2767 9918 2773 9919
rect 2767 9914 2768 9918
rect 2772 9914 2773 9918
rect 2767 9913 2773 9914
rect 2767 9909 2768 9913
rect 2772 9909 2773 9913
rect 2767 9908 2773 9909
rect 2767 9904 2768 9908
rect 2772 9904 2773 9908
rect 2767 9903 2773 9904
rect 2767 9899 2768 9903
rect 2772 9899 2773 9903
rect 2767 9898 2773 9899
rect 2767 9894 2768 9898
rect 2772 9894 2773 9898
rect 2767 9893 2773 9894
rect 2767 9889 2768 9893
rect 2772 9889 2773 9893
rect 2767 9888 2773 9889
rect 2767 9884 2768 9888
rect 2772 9884 2773 9888
rect 2767 9883 2773 9884
rect 2767 9879 2768 9883
rect 2772 9879 2773 9883
rect 2767 9878 2773 9879
rect 2767 9874 2768 9878
rect 2772 9874 2773 9878
rect 2767 9873 2773 9874
rect 2767 9869 2768 9873
rect 2772 9869 2773 9873
rect 2767 9868 2773 9869
rect 2767 9864 2768 9868
rect 2772 9864 2773 9868
rect 2767 9863 2773 9864
rect 2767 9859 2768 9863
rect 2772 9859 2773 9863
rect 2767 9858 2773 9859
rect 2767 9854 2768 9858
rect 2772 9854 2773 9858
rect 2767 9853 2773 9854
rect 2767 9849 2768 9853
rect 2772 9849 2773 9853
rect 2857 9964 2858 9968
rect 2862 9964 2863 9968
rect 2857 9963 2863 9964
rect 2857 9959 2858 9963
rect 2862 9959 2863 9963
rect 2857 9958 2863 9959
rect 2857 9954 2858 9958
rect 2862 9954 2863 9958
rect 2857 9953 2863 9954
rect 2857 9949 2858 9953
rect 2862 9949 2863 9953
rect 2857 9948 2863 9949
rect 2857 9944 2858 9948
rect 2862 9944 2863 9948
rect 2857 9943 2863 9944
rect 2857 9939 2858 9943
rect 2862 9939 2863 9943
rect 2857 9938 2863 9939
rect 2857 9934 2858 9938
rect 2862 9934 2863 9938
rect 2857 9933 2863 9934
rect 2857 9929 2858 9933
rect 2862 9929 2863 9933
rect 2857 9928 2863 9929
rect 2857 9924 2858 9928
rect 2862 9924 2863 9928
rect 2857 9923 2863 9924
rect 2857 9919 2858 9923
rect 2862 9919 2863 9923
rect 2857 9918 2863 9919
rect 2857 9914 2858 9918
rect 2862 9914 2863 9918
rect 2857 9913 2863 9914
rect 2857 9909 2858 9913
rect 2862 9909 2863 9913
rect 2857 9908 2863 9909
rect 2857 9904 2858 9908
rect 2862 9904 2863 9908
rect 2857 9903 2863 9904
rect 2857 9899 2858 9903
rect 2862 9899 2863 9903
rect 2857 9898 2863 9899
rect 2857 9894 2858 9898
rect 2862 9894 2863 9898
rect 2857 9893 2863 9894
rect 2857 9889 2858 9893
rect 2862 9889 2863 9893
rect 2857 9888 2863 9889
rect 2857 9884 2858 9888
rect 2862 9884 2863 9888
rect 2857 9883 2863 9884
rect 2857 9879 2858 9883
rect 2862 9879 2863 9883
rect 2857 9878 2863 9879
rect 2857 9874 2858 9878
rect 2862 9874 2863 9878
rect 2857 9873 2863 9874
rect 2857 9869 2858 9873
rect 2862 9869 2863 9873
rect 2857 9868 2863 9869
rect 2857 9864 2858 9868
rect 2862 9864 2863 9868
rect 2857 9863 2863 9864
rect 2857 9859 2858 9863
rect 2862 9859 2863 9863
rect 2857 9858 2863 9859
rect 2857 9854 2858 9858
rect 2862 9854 2863 9858
rect 2857 9853 2863 9854
rect 2767 9848 2773 9849
rect 2767 9844 2768 9848
rect 2772 9844 2773 9848
rect 2857 9849 2858 9853
rect 2862 9849 2863 9853
rect 2857 9848 2863 9849
rect 2857 9844 2858 9848
rect 2862 9844 2863 9848
rect 2767 9843 2863 9844
rect 2767 9839 2768 9843
rect 2772 9839 2773 9843
rect 2777 9839 2778 9843
rect 2782 9839 2783 9843
rect 2787 9839 2788 9843
rect 2792 9839 2793 9843
rect 2797 9839 2798 9843
rect 2802 9839 2803 9843
rect 2807 9839 2808 9843
rect 2812 9839 2813 9843
rect 2817 9839 2818 9843
rect 2822 9839 2823 9843
rect 2827 9839 2828 9843
rect 2832 9839 2833 9843
rect 2837 9839 2838 9843
rect 2842 9839 2843 9843
rect 2847 9839 2848 9843
rect 2852 9839 2853 9843
rect 2857 9839 2858 9843
rect 2862 9839 2863 9843
rect 2767 9838 2863 9839
rect 2928 9965 3000 9967
rect 2928 9961 2930 9965
rect 2934 9961 2937 9965
rect 2941 9961 2942 9965
rect 2946 9961 2947 9965
rect 2951 9961 2952 9965
rect 2956 9961 2957 9965
rect 2961 9961 2962 9965
rect 2966 9961 2967 9965
rect 2971 9961 2972 9965
rect 2976 9961 2977 9965
rect 2981 9961 2982 9965
rect 2986 9961 2987 9965
rect 2991 9961 2994 9965
rect 2998 9961 3000 9965
rect 2928 9959 3000 9961
rect 2928 9958 2936 9959
rect 2928 9954 2930 9958
rect 2934 9954 2936 9958
rect 2928 9953 2936 9954
rect 2992 9958 3000 9959
rect 2992 9954 2994 9958
rect 2998 9954 3000 9958
rect 2992 9953 3000 9954
rect 2928 9949 2930 9953
rect 2934 9949 2936 9953
rect 2928 9948 2936 9949
rect 2928 9944 2930 9948
rect 2934 9944 2936 9948
rect 2928 9943 2936 9944
rect 2928 9939 2930 9943
rect 2934 9939 2936 9943
rect 2928 9938 2936 9939
rect 2928 9934 2930 9938
rect 2934 9934 2936 9938
rect 2928 9933 2936 9934
rect 2928 9929 2930 9933
rect 2934 9929 2936 9933
rect 2928 9928 2936 9929
rect 2928 9924 2930 9928
rect 2934 9924 2936 9928
rect 2928 9923 2936 9924
rect 2928 9919 2930 9923
rect 2934 9919 2936 9923
rect 2928 9918 2936 9919
rect 2928 9914 2930 9918
rect 2934 9914 2936 9918
rect 2928 9913 2936 9914
rect 2928 9909 2930 9913
rect 2934 9909 2936 9913
rect 2928 9908 2936 9909
rect 2928 9904 2930 9908
rect 2934 9904 2936 9908
rect 2928 9903 2936 9904
rect 2928 9899 2930 9903
rect 2934 9899 2936 9903
rect 2928 9898 2936 9899
rect 2928 9894 2930 9898
rect 2934 9894 2936 9898
rect 2928 9893 2936 9894
rect 2928 9889 2930 9893
rect 2934 9889 2936 9893
rect 2928 9888 2936 9889
rect 2928 9884 2930 9888
rect 2934 9884 2936 9888
rect 2928 9883 2936 9884
rect 2928 9879 2930 9883
rect 2934 9879 2936 9883
rect 2928 9878 2936 9879
rect 2928 9874 2930 9878
rect 2934 9874 2936 9878
rect 2928 9873 2936 9874
rect 2928 9869 2930 9873
rect 2934 9869 2936 9873
rect 2928 9868 2936 9869
rect 2928 9864 2930 9868
rect 2934 9864 2936 9868
rect 2992 9949 2994 9953
rect 2998 9949 3000 9953
rect 2992 9948 3000 9949
rect 2992 9944 2994 9948
rect 2998 9944 3000 9948
rect 2992 9943 3000 9944
rect 2992 9939 2994 9943
rect 2998 9939 3000 9943
rect 2992 9938 3000 9939
rect 2992 9934 2994 9938
rect 2998 9934 3000 9938
rect 2992 9933 3000 9934
rect 2992 9929 2994 9933
rect 2998 9929 3000 9933
rect 2992 9928 3000 9929
rect 2992 9924 2994 9928
rect 2998 9924 3000 9928
rect 2992 9923 3000 9924
rect 2992 9919 2994 9923
rect 2998 9919 3000 9923
rect 2992 9918 3000 9919
rect 2992 9914 2994 9918
rect 2998 9914 3000 9918
rect 2992 9913 3000 9914
rect 2992 9909 2994 9913
rect 2998 9909 3000 9913
rect 2992 9908 3000 9909
rect 2992 9904 2994 9908
rect 2998 9904 3000 9908
rect 2992 9903 3000 9904
rect 2992 9899 2994 9903
rect 2998 9899 3000 9903
rect 2992 9898 3000 9899
rect 2992 9894 2994 9898
rect 2998 9894 3000 9898
rect 2992 9893 3000 9894
rect 2992 9889 2994 9893
rect 2998 9889 3000 9893
rect 2992 9888 3000 9889
rect 2992 9884 2994 9888
rect 2998 9884 3000 9888
rect 2992 9883 3000 9884
rect 2992 9879 2994 9883
rect 2998 9879 3000 9883
rect 2992 9878 3000 9879
rect 2992 9874 2994 9878
rect 2998 9874 3000 9878
rect 2992 9873 3000 9874
rect 2992 9869 2994 9873
rect 2998 9869 3000 9873
rect 2992 9868 3000 9869
rect 2992 9864 2994 9868
rect 2998 9864 3000 9868
rect 2928 9863 2936 9864
rect 2928 9859 2930 9863
rect 2934 9859 2936 9863
rect 2928 9858 2936 9859
rect 2992 9863 3000 9864
rect 2992 9859 2994 9863
rect 2998 9859 3000 9863
rect 2992 9858 3000 9859
rect 2928 9856 3000 9858
rect 2928 9852 2930 9856
rect 2934 9852 2937 9856
rect 2941 9852 2942 9856
rect 2946 9852 2947 9856
rect 2951 9852 2952 9856
rect 2956 9852 2957 9856
rect 2961 9852 2962 9856
rect 2966 9852 2967 9856
rect 2971 9852 2972 9856
rect 2976 9852 2977 9856
rect 2981 9852 2982 9856
rect 2986 9852 2987 9856
rect 2991 9852 2994 9856
rect 2998 9852 3000 9856
rect 2928 9850 3000 9852
rect 3076 9978 3172 9979
rect 3076 9974 3077 9978
rect 3081 9974 3082 9978
rect 3086 9974 3087 9978
rect 3091 9974 3092 9978
rect 3096 9974 3097 9978
rect 3101 9974 3102 9978
rect 3106 9974 3107 9978
rect 3111 9974 3112 9978
rect 3116 9974 3117 9978
rect 3121 9974 3122 9978
rect 3126 9974 3127 9978
rect 3131 9974 3132 9978
rect 3136 9974 3137 9978
rect 3141 9974 3142 9978
rect 3146 9974 3147 9978
rect 3151 9974 3152 9978
rect 3156 9974 3157 9978
rect 3161 9974 3162 9978
rect 3166 9974 3167 9978
rect 3171 9974 3172 9978
rect 3076 9973 3172 9974
rect 3076 9969 3077 9973
rect 3081 9969 3082 9973
rect 3076 9968 3082 9969
rect 3076 9964 3077 9968
rect 3081 9964 3082 9968
rect 3166 9969 3167 9973
rect 3171 9969 3172 9973
rect 3166 9968 3172 9969
rect 3076 9963 3082 9964
rect 3076 9959 3077 9963
rect 3081 9959 3082 9963
rect 3076 9958 3082 9959
rect 3076 9954 3077 9958
rect 3081 9954 3082 9958
rect 3076 9953 3082 9954
rect 3076 9949 3077 9953
rect 3081 9949 3082 9953
rect 3076 9948 3082 9949
rect 3076 9944 3077 9948
rect 3081 9944 3082 9948
rect 3076 9943 3082 9944
rect 3076 9939 3077 9943
rect 3081 9939 3082 9943
rect 3076 9938 3082 9939
rect 3076 9934 3077 9938
rect 3081 9934 3082 9938
rect 3076 9933 3082 9934
rect 3076 9929 3077 9933
rect 3081 9929 3082 9933
rect 3076 9928 3082 9929
rect 3076 9924 3077 9928
rect 3081 9924 3082 9928
rect 3076 9923 3082 9924
rect 3076 9919 3077 9923
rect 3081 9919 3082 9923
rect 3076 9918 3082 9919
rect 3076 9914 3077 9918
rect 3081 9914 3082 9918
rect 3076 9913 3082 9914
rect 3076 9909 3077 9913
rect 3081 9909 3082 9913
rect 3076 9908 3082 9909
rect 3076 9904 3077 9908
rect 3081 9904 3082 9908
rect 3076 9903 3082 9904
rect 3076 9899 3077 9903
rect 3081 9899 3082 9903
rect 3076 9898 3082 9899
rect 3076 9894 3077 9898
rect 3081 9894 3082 9898
rect 3076 9893 3082 9894
rect 3076 9889 3077 9893
rect 3081 9889 3082 9893
rect 3076 9888 3082 9889
rect 3076 9884 3077 9888
rect 3081 9884 3082 9888
rect 3076 9883 3082 9884
rect 3076 9879 3077 9883
rect 3081 9879 3082 9883
rect 3076 9878 3082 9879
rect 3076 9874 3077 9878
rect 3081 9874 3082 9878
rect 3076 9873 3082 9874
rect 3076 9869 3077 9873
rect 3081 9869 3082 9873
rect 3076 9868 3082 9869
rect 3076 9864 3077 9868
rect 3081 9864 3082 9868
rect 3076 9863 3082 9864
rect 3076 9859 3077 9863
rect 3081 9859 3082 9863
rect 3076 9858 3082 9859
rect 3076 9854 3077 9858
rect 3081 9854 3082 9858
rect 3076 9853 3082 9854
rect 3076 9849 3077 9853
rect 3081 9849 3082 9853
rect 3166 9964 3167 9968
rect 3171 9964 3172 9968
rect 3166 9963 3172 9964
rect 3166 9959 3167 9963
rect 3171 9959 3172 9963
rect 3166 9958 3172 9959
rect 3166 9954 3167 9958
rect 3171 9954 3172 9958
rect 3166 9953 3172 9954
rect 3166 9949 3167 9953
rect 3171 9949 3172 9953
rect 3166 9948 3172 9949
rect 3166 9944 3167 9948
rect 3171 9944 3172 9948
rect 3166 9943 3172 9944
rect 3166 9939 3167 9943
rect 3171 9939 3172 9943
rect 3166 9938 3172 9939
rect 3166 9934 3167 9938
rect 3171 9934 3172 9938
rect 3166 9933 3172 9934
rect 3166 9929 3167 9933
rect 3171 9929 3172 9933
rect 3166 9928 3172 9929
rect 3166 9924 3167 9928
rect 3171 9924 3172 9928
rect 3166 9923 3172 9924
rect 3166 9919 3167 9923
rect 3171 9919 3172 9923
rect 3166 9918 3172 9919
rect 3166 9914 3167 9918
rect 3171 9914 3172 9918
rect 3166 9913 3172 9914
rect 3166 9909 3167 9913
rect 3171 9909 3172 9913
rect 3166 9908 3172 9909
rect 3166 9904 3167 9908
rect 3171 9904 3172 9908
rect 3166 9903 3172 9904
rect 3166 9899 3167 9903
rect 3171 9899 3172 9903
rect 3166 9898 3172 9899
rect 3166 9894 3167 9898
rect 3171 9894 3172 9898
rect 3166 9893 3172 9894
rect 3166 9889 3167 9893
rect 3171 9889 3172 9893
rect 3166 9888 3172 9889
rect 3166 9884 3167 9888
rect 3171 9884 3172 9888
rect 3166 9883 3172 9884
rect 3166 9879 3167 9883
rect 3171 9879 3172 9883
rect 3166 9878 3172 9879
rect 3166 9874 3167 9878
rect 3171 9874 3172 9878
rect 3166 9873 3172 9874
rect 3166 9869 3167 9873
rect 3171 9869 3172 9873
rect 3166 9868 3172 9869
rect 3166 9864 3167 9868
rect 3171 9864 3172 9868
rect 3166 9863 3172 9864
rect 3166 9859 3167 9863
rect 3171 9859 3172 9863
rect 3166 9858 3172 9859
rect 3166 9854 3167 9858
rect 3171 9854 3172 9858
rect 3166 9853 3172 9854
rect 3076 9848 3082 9849
rect 3076 9844 3077 9848
rect 3081 9844 3082 9848
rect 3166 9849 3167 9853
rect 3171 9849 3172 9853
rect 3166 9848 3172 9849
rect 3166 9844 3167 9848
rect 3171 9844 3172 9848
rect 3076 9843 3172 9844
rect 3076 9839 3077 9843
rect 3081 9839 3082 9843
rect 3086 9839 3087 9843
rect 3091 9839 3092 9843
rect 3096 9839 3097 9843
rect 3101 9839 3102 9843
rect 3106 9839 3107 9843
rect 3111 9839 3112 9843
rect 3116 9839 3117 9843
rect 3121 9839 3122 9843
rect 3126 9839 3127 9843
rect 3131 9839 3132 9843
rect 3136 9839 3137 9843
rect 3141 9839 3142 9843
rect 3146 9839 3147 9843
rect 3151 9839 3152 9843
rect 3156 9839 3157 9843
rect 3161 9839 3162 9843
rect 3166 9839 3167 9843
rect 3171 9839 3172 9843
rect 3076 9838 3172 9839
rect 3237 9965 3309 9967
rect 3237 9961 3239 9965
rect 3243 9961 3246 9965
rect 3250 9961 3251 9965
rect 3255 9961 3256 9965
rect 3260 9961 3261 9965
rect 3265 9961 3266 9965
rect 3270 9961 3271 9965
rect 3275 9961 3276 9965
rect 3280 9961 3281 9965
rect 3285 9961 3286 9965
rect 3290 9961 3291 9965
rect 3295 9961 3296 9965
rect 3300 9961 3303 9965
rect 3307 9961 3309 9965
rect 3237 9959 3309 9961
rect 3237 9958 3245 9959
rect 3237 9954 3239 9958
rect 3243 9954 3245 9958
rect 3237 9953 3245 9954
rect 3301 9958 3309 9959
rect 3301 9954 3303 9958
rect 3307 9954 3309 9958
rect 3301 9953 3309 9954
rect 3237 9949 3239 9953
rect 3243 9949 3245 9953
rect 3237 9948 3245 9949
rect 3237 9944 3239 9948
rect 3243 9944 3245 9948
rect 3237 9943 3245 9944
rect 3237 9939 3239 9943
rect 3243 9939 3245 9943
rect 3237 9938 3245 9939
rect 3237 9934 3239 9938
rect 3243 9934 3245 9938
rect 3237 9933 3245 9934
rect 3237 9929 3239 9933
rect 3243 9929 3245 9933
rect 3237 9928 3245 9929
rect 3237 9924 3239 9928
rect 3243 9924 3245 9928
rect 3237 9923 3245 9924
rect 3237 9919 3239 9923
rect 3243 9919 3245 9923
rect 3237 9918 3245 9919
rect 3237 9914 3239 9918
rect 3243 9914 3245 9918
rect 3237 9913 3245 9914
rect 3237 9909 3239 9913
rect 3243 9909 3245 9913
rect 3237 9908 3245 9909
rect 3237 9904 3239 9908
rect 3243 9904 3245 9908
rect 3237 9903 3245 9904
rect 3237 9899 3239 9903
rect 3243 9899 3245 9903
rect 3237 9898 3245 9899
rect 3237 9894 3239 9898
rect 3243 9894 3245 9898
rect 3237 9893 3245 9894
rect 3237 9889 3239 9893
rect 3243 9889 3245 9893
rect 3237 9888 3245 9889
rect 3237 9884 3239 9888
rect 3243 9884 3245 9888
rect 3237 9883 3245 9884
rect 3237 9879 3239 9883
rect 3243 9879 3245 9883
rect 3237 9878 3245 9879
rect 3237 9874 3239 9878
rect 3243 9874 3245 9878
rect 3237 9873 3245 9874
rect 3237 9869 3239 9873
rect 3243 9869 3245 9873
rect 3237 9868 3245 9869
rect 3237 9864 3239 9868
rect 3243 9864 3245 9868
rect 3301 9949 3303 9953
rect 3307 9949 3309 9953
rect 3301 9948 3309 9949
rect 3301 9944 3303 9948
rect 3307 9944 3309 9948
rect 3301 9943 3309 9944
rect 3301 9939 3303 9943
rect 3307 9939 3309 9943
rect 3301 9938 3309 9939
rect 3301 9934 3303 9938
rect 3307 9934 3309 9938
rect 3301 9933 3309 9934
rect 3301 9929 3303 9933
rect 3307 9929 3309 9933
rect 3301 9928 3309 9929
rect 3301 9924 3303 9928
rect 3307 9924 3309 9928
rect 3301 9923 3309 9924
rect 3301 9919 3303 9923
rect 3307 9919 3309 9923
rect 3301 9918 3309 9919
rect 3301 9914 3303 9918
rect 3307 9914 3309 9918
rect 3301 9913 3309 9914
rect 3301 9909 3303 9913
rect 3307 9909 3309 9913
rect 3301 9908 3309 9909
rect 3301 9904 3303 9908
rect 3307 9904 3309 9908
rect 3301 9903 3309 9904
rect 3301 9899 3303 9903
rect 3307 9899 3309 9903
rect 3301 9898 3309 9899
rect 3301 9894 3303 9898
rect 3307 9894 3309 9898
rect 3301 9893 3309 9894
rect 3301 9889 3303 9893
rect 3307 9889 3309 9893
rect 3301 9888 3309 9889
rect 3301 9884 3303 9888
rect 3307 9884 3309 9888
rect 3301 9883 3309 9884
rect 3301 9879 3303 9883
rect 3307 9879 3309 9883
rect 3301 9878 3309 9879
rect 3301 9874 3303 9878
rect 3307 9874 3309 9878
rect 3301 9873 3309 9874
rect 3301 9869 3303 9873
rect 3307 9869 3309 9873
rect 3301 9868 3309 9869
rect 3301 9864 3303 9868
rect 3307 9864 3309 9868
rect 3237 9863 3245 9864
rect 3237 9859 3239 9863
rect 3243 9859 3245 9863
rect 3237 9858 3245 9859
rect 3301 9863 3309 9864
rect 3301 9859 3303 9863
rect 3307 9859 3309 9863
rect 3301 9858 3309 9859
rect 3237 9856 3309 9858
rect 3237 9852 3239 9856
rect 3243 9852 3246 9856
rect 3250 9852 3251 9856
rect 3255 9852 3256 9856
rect 3260 9852 3261 9856
rect 3265 9852 3266 9856
rect 3270 9852 3271 9856
rect 3275 9852 3276 9856
rect 3280 9852 3281 9856
rect 3285 9852 3286 9856
rect 3290 9852 3291 9856
rect 3295 9852 3296 9856
rect 3300 9852 3303 9856
rect 3307 9852 3309 9856
rect 3237 9850 3309 9852
rect 3385 9978 3481 9979
rect 3385 9974 3386 9978
rect 3390 9974 3391 9978
rect 3395 9974 3396 9978
rect 3400 9974 3401 9978
rect 3405 9974 3406 9978
rect 3410 9974 3411 9978
rect 3415 9974 3416 9978
rect 3420 9974 3421 9978
rect 3425 9974 3426 9978
rect 3430 9974 3431 9978
rect 3435 9974 3436 9978
rect 3440 9974 3441 9978
rect 3445 9974 3446 9978
rect 3450 9974 3451 9978
rect 3455 9974 3456 9978
rect 3460 9974 3461 9978
rect 3465 9974 3466 9978
rect 3470 9974 3471 9978
rect 3475 9974 3476 9978
rect 3480 9974 3481 9978
rect 3385 9973 3481 9974
rect 3385 9969 3386 9973
rect 3390 9969 3391 9973
rect 3385 9968 3391 9969
rect 3385 9964 3386 9968
rect 3390 9964 3391 9968
rect 3475 9969 3476 9973
rect 3480 9969 3481 9973
rect 3475 9968 3481 9969
rect 3385 9963 3391 9964
rect 3385 9959 3386 9963
rect 3390 9959 3391 9963
rect 3385 9958 3391 9959
rect 3385 9954 3386 9958
rect 3390 9954 3391 9958
rect 3385 9953 3391 9954
rect 3385 9949 3386 9953
rect 3390 9949 3391 9953
rect 3385 9948 3391 9949
rect 3385 9944 3386 9948
rect 3390 9944 3391 9948
rect 3385 9943 3391 9944
rect 3385 9939 3386 9943
rect 3390 9939 3391 9943
rect 3385 9938 3391 9939
rect 3385 9934 3386 9938
rect 3390 9934 3391 9938
rect 3385 9933 3391 9934
rect 3385 9929 3386 9933
rect 3390 9929 3391 9933
rect 3385 9928 3391 9929
rect 3385 9924 3386 9928
rect 3390 9924 3391 9928
rect 3385 9923 3391 9924
rect 3385 9919 3386 9923
rect 3390 9919 3391 9923
rect 3385 9918 3391 9919
rect 3385 9914 3386 9918
rect 3390 9914 3391 9918
rect 3385 9913 3391 9914
rect 3385 9909 3386 9913
rect 3390 9909 3391 9913
rect 3385 9908 3391 9909
rect 3385 9904 3386 9908
rect 3390 9904 3391 9908
rect 3385 9903 3391 9904
rect 3385 9899 3386 9903
rect 3390 9899 3391 9903
rect 3385 9898 3391 9899
rect 3385 9894 3386 9898
rect 3390 9894 3391 9898
rect 3385 9893 3391 9894
rect 3385 9889 3386 9893
rect 3390 9889 3391 9893
rect 3385 9888 3391 9889
rect 3385 9884 3386 9888
rect 3390 9884 3391 9888
rect 3385 9883 3391 9884
rect 3385 9879 3386 9883
rect 3390 9879 3391 9883
rect 3385 9878 3391 9879
rect 3385 9874 3386 9878
rect 3390 9874 3391 9878
rect 3385 9873 3391 9874
rect 3385 9869 3386 9873
rect 3390 9869 3391 9873
rect 3385 9868 3391 9869
rect 3385 9864 3386 9868
rect 3390 9864 3391 9868
rect 3385 9863 3391 9864
rect 3385 9859 3386 9863
rect 3390 9859 3391 9863
rect 3385 9858 3391 9859
rect 3385 9854 3386 9858
rect 3390 9854 3391 9858
rect 3385 9853 3391 9854
rect 3385 9849 3386 9853
rect 3390 9849 3391 9853
rect 3475 9964 3476 9968
rect 3480 9964 3481 9968
rect 3475 9963 3481 9964
rect 3475 9959 3476 9963
rect 3480 9959 3481 9963
rect 3475 9958 3481 9959
rect 3475 9954 3476 9958
rect 3480 9954 3481 9958
rect 3475 9953 3481 9954
rect 3475 9949 3476 9953
rect 3480 9949 3481 9953
rect 3475 9948 3481 9949
rect 3475 9944 3476 9948
rect 3480 9944 3481 9948
rect 3475 9943 3481 9944
rect 3475 9939 3476 9943
rect 3480 9939 3481 9943
rect 3475 9938 3481 9939
rect 3475 9934 3476 9938
rect 3480 9934 3481 9938
rect 3475 9933 3481 9934
rect 3475 9929 3476 9933
rect 3480 9929 3481 9933
rect 3475 9928 3481 9929
rect 3475 9924 3476 9928
rect 3480 9924 3481 9928
rect 3475 9923 3481 9924
rect 3475 9919 3476 9923
rect 3480 9919 3481 9923
rect 3475 9918 3481 9919
rect 3475 9914 3476 9918
rect 3480 9914 3481 9918
rect 3475 9913 3481 9914
rect 3475 9909 3476 9913
rect 3480 9909 3481 9913
rect 3475 9908 3481 9909
rect 3475 9904 3476 9908
rect 3480 9904 3481 9908
rect 3475 9903 3481 9904
rect 3475 9899 3476 9903
rect 3480 9899 3481 9903
rect 3475 9898 3481 9899
rect 3475 9894 3476 9898
rect 3480 9894 3481 9898
rect 3475 9893 3481 9894
rect 3475 9889 3476 9893
rect 3480 9889 3481 9893
rect 3475 9888 3481 9889
rect 3475 9884 3476 9888
rect 3480 9884 3481 9888
rect 3475 9883 3481 9884
rect 3475 9879 3476 9883
rect 3480 9879 3481 9883
rect 3475 9878 3481 9879
rect 3475 9874 3476 9878
rect 3480 9874 3481 9878
rect 3475 9873 3481 9874
rect 3475 9869 3476 9873
rect 3480 9869 3481 9873
rect 3475 9868 3481 9869
rect 3475 9864 3476 9868
rect 3480 9864 3481 9868
rect 3475 9863 3481 9864
rect 3475 9859 3476 9863
rect 3480 9859 3481 9863
rect 3475 9858 3481 9859
rect 3475 9854 3476 9858
rect 3480 9854 3481 9858
rect 3475 9853 3481 9854
rect 3385 9848 3391 9849
rect 3385 9844 3386 9848
rect 3390 9844 3391 9848
rect 3475 9849 3476 9853
rect 3480 9849 3481 9853
rect 3475 9848 3481 9849
rect 3475 9844 3476 9848
rect 3480 9844 3481 9848
rect 3385 9843 3481 9844
rect 3385 9839 3386 9843
rect 3390 9839 3391 9843
rect 3395 9839 3396 9843
rect 3400 9839 3401 9843
rect 3405 9839 3406 9843
rect 3410 9839 3411 9843
rect 3415 9839 3416 9843
rect 3420 9839 3421 9843
rect 3425 9839 3426 9843
rect 3430 9839 3431 9843
rect 3435 9839 3436 9843
rect 3440 9839 3441 9843
rect 3445 9839 3446 9843
rect 3450 9839 3451 9843
rect 3455 9839 3456 9843
rect 3460 9839 3461 9843
rect 3465 9839 3466 9843
rect 3470 9839 3471 9843
rect 3475 9839 3476 9843
rect 3480 9839 3481 9843
rect 3385 9838 3481 9839
rect 3546 9965 3618 9967
rect 3546 9961 3548 9965
rect 3552 9961 3555 9965
rect 3559 9961 3560 9965
rect 3564 9961 3565 9965
rect 3569 9961 3570 9965
rect 3574 9961 3575 9965
rect 3579 9961 3580 9965
rect 3584 9961 3585 9965
rect 3589 9961 3590 9965
rect 3594 9961 3595 9965
rect 3599 9961 3600 9965
rect 3604 9961 3605 9965
rect 3609 9961 3612 9965
rect 3616 9961 3618 9965
rect 3546 9959 3618 9961
rect 3546 9958 3554 9959
rect 3546 9954 3548 9958
rect 3552 9954 3554 9958
rect 3546 9953 3554 9954
rect 3610 9958 3618 9959
rect 3610 9954 3612 9958
rect 3616 9954 3618 9958
rect 3610 9953 3618 9954
rect 3546 9949 3548 9953
rect 3552 9949 3554 9953
rect 3546 9948 3554 9949
rect 3546 9944 3548 9948
rect 3552 9944 3554 9948
rect 3546 9943 3554 9944
rect 3546 9939 3548 9943
rect 3552 9939 3554 9943
rect 3546 9938 3554 9939
rect 3546 9934 3548 9938
rect 3552 9934 3554 9938
rect 3546 9933 3554 9934
rect 3546 9929 3548 9933
rect 3552 9929 3554 9933
rect 3546 9928 3554 9929
rect 3546 9924 3548 9928
rect 3552 9924 3554 9928
rect 3546 9923 3554 9924
rect 3546 9919 3548 9923
rect 3552 9919 3554 9923
rect 3546 9918 3554 9919
rect 3546 9914 3548 9918
rect 3552 9914 3554 9918
rect 3546 9913 3554 9914
rect 3546 9909 3548 9913
rect 3552 9909 3554 9913
rect 3546 9908 3554 9909
rect 3546 9904 3548 9908
rect 3552 9904 3554 9908
rect 3546 9903 3554 9904
rect 3546 9899 3548 9903
rect 3552 9899 3554 9903
rect 3546 9898 3554 9899
rect 3546 9894 3548 9898
rect 3552 9894 3554 9898
rect 3546 9893 3554 9894
rect 3546 9889 3548 9893
rect 3552 9889 3554 9893
rect 3546 9888 3554 9889
rect 3546 9884 3548 9888
rect 3552 9884 3554 9888
rect 3546 9883 3554 9884
rect 3546 9879 3548 9883
rect 3552 9879 3554 9883
rect 3546 9878 3554 9879
rect 3546 9874 3548 9878
rect 3552 9874 3554 9878
rect 3546 9873 3554 9874
rect 3546 9869 3548 9873
rect 3552 9869 3554 9873
rect 3546 9868 3554 9869
rect 3546 9864 3548 9868
rect 3552 9864 3554 9868
rect 3610 9949 3612 9953
rect 3616 9949 3618 9953
rect 3610 9948 3618 9949
rect 3610 9944 3612 9948
rect 3616 9944 3618 9948
rect 3610 9943 3618 9944
rect 3610 9939 3612 9943
rect 3616 9939 3618 9943
rect 3610 9938 3618 9939
rect 3610 9934 3612 9938
rect 3616 9934 3618 9938
rect 3610 9933 3618 9934
rect 3610 9929 3612 9933
rect 3616 9929 3618 9933
rect 3610 9928 3618 9929
rect 3610 9924 3612 9928
rect 3616 9924 3618 9928
rect 3610 9923 3618 9924
rect 3610 9919 3612 9923
rect 3616 9919 3618 9923
rect 3610 9918 3618 9919
rect 3610 9914 3612 9918
rect 3616 9914 3618 9918
rect 3610 9913 3618 9914
rect 3610 9909 3612 9913
rect 3616 9909 3618 9913
rect 3610 9908 3618 9909
rect 3610 9904 3612 9908
rect 3616 9904 3618 9908
rect 3610 9903 3618 9904
rect 3610 9899 3612 9903
rect 3616 9899 3618 9903
rect 3610 9898 3618 9899
rect 3610 9894 3612 9898
rect 3616 9894 3618 9898
rect 3610 9893 3618 9894
rect 3610 9889 3612 9893
rect 3616 9889 3618 9893
rect 3610 9888 3618 9889
rect 3610 9884 3612 9888
rect 3616 9884 3618 9888
rect 3610 9883 3618 9884
rect 3610 9879 3612 9883
rect 3616 9879 3618 9883
rect 3610 9878 3618 9879
rect 3610 9874 3612 9878
rect 3616 9874 3618 9878
rect 3610 9873 3618 9874
rect 3610 9869 3612 9873
rect 3616 9869 3618 9873
rect 3610 9868 3618 9869
rect 3610 9864 3612 9868
rect 3616 9864 3618 9868
rect 3546 9863 3554 9864
rect 3546 9859 3548 9863
rect 3552 9859 3554 9863
rect 3546 9858 3554 9859
rect 3610 9863 3618 9864
rect 3610 9859 3612 9863
rect 3616 9859 3618 9863
rect 3610 9858 3618 9859
rect 3546 9856 3618 9858
rect 3546 9852 3548 9856
rect 3552 9852 3555 9856
rect 3559 9852 3560 9856
rect 3564 9852 3565 9856
rect 3569 9852 3570 9856
rect 3574 9852 3575 9856
rect 3579 9852 3580 9856
rect 3584 9852 3585 9856
rect 3589 9852 3590 9856
rect 3594 9852 3595 9856
rect 3599 9852 3600 9856
rect 3604 9852 3605 9856
rect 3609 9852 3612 9856
rect 3616 9852 3618 9856
rect 3546 9850 3618 9852
rect 3694 9978 3790 9979
rect 3694 9974 3695 9978
rect 3699 9974 3700 9978
rect 3704 9974 3705 9978
rect 3709 9974 3710 9978
rect 3714 9974 3715 9978
rect 3719 9974 3720 9978
rect 3724 9974 3725 9978
rect 3729 9974 3730 9978
rect 3734 9974 3735 9978
rect 3739 9974 3740 9978
rect 3744 9974 3745 9978
rect 3749 9974 3750 9978
rect 3754 9974 3755 9978
rect 3759 9974 3760 9978
rect 3764 9974 3765 9978
rect 3769 9974 3770 9978
rect 3774 9974 3775 9978
rect 3779 9974 3780 9978
rect 3784 9974 3785 9978
rect 3789 9974 3790 9978
rect 3694 9973 3790 9974
rect 3694 9969 3695 9973
rect 3699 9969 3700 9973
rect 3694 9968 3700 9969
rect 3694 9964 3695 9968
rect 3699 9964 3700 9968
rect 3784 9969 3785 9973
rect 3789 9969 3790 9973
rect 3784 9968 3790 9969
rect 3694 9963 3700 9964
rect 3694 9959 3695 9963
rect 3699 9959 3700 9963
rect 3694 9958 3700 9959
rect 3694 9954 3695 9958
rect 3699 9954 3700 9958
rect 3694 9953 3700 9954
rect 3694 9949 3695 9953
rect 3699 9949 3700 9953
rect 3694 9948 3700 9949
rect 3694 9944 3695 9948
rect 3699 9944 3700 9948
rect 3694 9943 3700 9944
rect 3694 9939 3695 9943
rect 3699 9939 3700 9943
rect 3694 9938 3700 9939
rect 3694 9934 3695 9938
rect 3699 9934 3700 9938
rect 3694 9933 3700 9934
rect 3694 9929 3695 9933
rect 3699 9929 3700 9933
rect 3694 9928 3700 9929
rect 3694 9924 3695 9928
rect 3699 9924 3700 9928
rect 3694 9923 3700 9924
rect 3694 9919 3695 9923
rect 3699 9919 3700 9923
rect 3694 9918 3700 9919
rect 3694 9914 3695 9918
rect 3699 9914 3700 9918
rect 3694 9913 3700 9914
rect 3694 9909 3695 9913
rect 3699 9909 3700 9913
rect 3694 9908 3700 9909
rect 3694 9904 3695 9908
rect 3699 9904 3700 9908
rect 3694 9903 3700 9904
rect 3694 9899 3695 9903
rect 3699 9899 3700 9903
rect 3694 9898 3700 9899
rect 3694 9894 3695 9898
rect 3699 9894 3700 9898
rect 3694 9893 3700 9894
rect 3694 9889 3695 9893
rect 3699 9889 3700 9893
rect 3694 9888 3700 9889
rect 3694 9884 3695 9888
rect 3699 9884 3700 9888
rect 3694 9883 3700 9884
rect 3694 9879 3695 9883
rect 3699 9879 3700 9883
rect 3694 9878 3700 9879
rect 3694 9874 3695 9878
rect 3699 9874 3700 9878
rect 3694 9873 3700 9874
rect 3694 9869 3695 9873
rect 3699 9869 3700 9873
rect 3694 9868 3700 9869
rect 3694 9864 3695 9868
rect 3699 9864 3700 9868
rect 3694 9863 3700 9864
rect 3694 9859 3695 9863
rect 3699 9859 3700 9863
rect 3694 9858 3700 9859
rect 3694 9854 3695 9858
rect 3699 9854 3700 9858
rect 3694 9853 3700 9854
rect 3694 9849 3695 9853
rect 3699 9849 3700 9853
rect 3784 9964 3785 9968
rect 3789 9964 3790 9968
rect 3784 9963 3790 9964
rect 3784 9959 3785 9963
rect 3789 9959 3790 9963
rect 3784 9958 3790 9959
rect 3784 9954 3785 9958
rect 3789 9954 3790 9958
rect 3784 9953 3790 9954
rect 3784 9949 3785 9953
rect 3789 9949 3790 9953
rect 3784 9948 3790 9949
rect 3784 9944 3785 9948
rect 3789 9944 3790 9948
rect 3784 9943 3790 9944
rect 3784 9939 3785 9943
rect 3789 9939 3790 9943
rect 3784 9938 3790 9939
rect 3784 9934 3785 9938
rect 3789 9934 3790 9938
rect 3784 9933 3790 9934
rect 3784 9929 3785 9933
rect 3789 9929 3790 9933
rect 3784 9928 3790 9929
rect 3784 9924 3785 9928
rect 3789 9924 3790 9928
rect 3784 9923 3790 9924
rect 3784 9919 3785 9923
rect 3789 9919 3790 9923
rect 3784 9918 3790 9919
rect 3784 9914 3785 9918
rect 3789 9914 3790 9918
rect 3784 9913 3790 9914
rect 3784 9909 3785 9913
rect 3789 9909 3790 9913
rect 3784 9908 3790 9909
rect 3784 9904 3785 9908
rect 3789 9904 3790 9908
rect 3784 9903 3790 9904
rect 3784 9899 3785 9903
rect 3789 9899 3790 9903
rect 3784 9898 3790 9899
rect 3784 9894 3785 9898
rect 3789 9894 3790 9898
rect 3784 9893 3790 9894
rect 3784 9889 3785 9893
rect 3789 9889 3790 9893
rect 3784 9888 3790 9889
rect 3784 9884 3785 9888
rect 3789 9884 3790 9888
rect 3784 9883 3790 9884
rect 3784 9879 3785 9883
rect 3789 9879 3790 9883
rect 3784 9878 3790 9879
rect 3784 9874 3785 9878
rect 3789 9874 3790 9878
rect 3784 9873 3790 9874
rect 3784 9869 3785 9873
rect 3789 9869 3790 9873
rect 3784 9868 3790 9869
rect 3784 9864 3785 9868
rect 3789 9864 3790 9868
rect 3784 9863 3790 9864
rect 3784 9859 3785 9863
rect 3789 9859 3790 9863
rect 3784 9858 3790 9859
rect 3784 9854 3785 9858
rect 3789 9854 3790 9858
rect 3784 9853 3790 9854
rect 3694 9848 3700 9849
rect 3694 9844 3695 9848
rect 3699 9844 3700 9848
rect 3784 9849 3785 9853
rect 3789 9849 3790 9853
rect 3784 9848 3790 9849
rect 3784 9844 3785 9848
rect 3789 9844 3790 9848
rect 3694 9843 3790 9844
rect 3694 9839 3695 9843
rect 3699 9839 3700 9843
rect 3704 9839 3705 9843
rect 3709 9839 3710 9843
rect 3714 9839 3715 9843
rect 3719 9839 3720 9843
rect 3724 9839 3725 9843
rect 3729 9839 3730 9843
rect 3734 9839 3735 9843
rect 3739 9839 3740 9843
rect 3744 9839 3745 9843
rect 3749 9839 3750 9843
rect 3754 9839 3755 9843
rect 3759 9839 3760 9843
rect 3764 9839 3765 9843
rect 3769 9839 3770 9843
rect 3774 9839 3775 9843
rect 3779 9839 3780 9843
rect 3784 9839 3785 9843
rect 3789 9839 3790 9843
rect 3694 9838 3790 9839
rect 3855 9965 3927 9967
rect 3855 9961 3857 9965
rect 3861 9961 3864 9965
rect 3868 9961 3869 9965
rect 3873 9961 3874 9965
rect 3878 9961 3879 9965
rect 3883 9961 3884 9965
rect 3888 9961 3889 9965
rect 3893 9961 3894 9965
rect 3898 9961 3899 9965
rect 3903 9961 3904 9965
rect 3908 9961 3909 9965
rect 3913 9961 3914 9965
rect 3918 9961 3921 9965
rect 3925 9961 3927 9965
rect 3855 9959 3927 9961
rect 3855 9958 3863 9959
rect 3855 9954 3857 9958
rect 3861 9954 3863 9958
rect 3855 9953 3863 9954
rect 3919 9958 3927 9959
rect 3919 9954 3921 9958
rect 3925 9954 3927 9958
rect 3919 9953 3927 9954
rect 3855 9949 3857 9953
rect 3861 9949 3863 9953
rect 3855 9948 3863 9949
rect 3855 9944 3857 9948
rect 3861 9944 3863 9948
rect 3855 9943 3863 9944
rect 3855 9939 3857 9943
rect 3861 9939 3863 9943
rect 3855 9938 3863 9939
rect 3855 9934 3857 9938
rect 3861 9934 3863 9938
rect 3855 9933 3863 9934
rect 3855 9929 3857 9933
rect 3861 9929 3863 9933
rect 3855 9928 3863 9929
rect 3855 9924 3857 9928
rect 3861 9924 3863 9928
rect 3855 9923 3863 9924
rect 3855 9919 3857 9923
rect 3861 9919 3863 9923
rect 3855 9918 3863 9919
rect 3855 9914 3857 9918
rect 3861 9914 3863 9918
rect 3855 9913 3863 9914
rect 3855 9909 3857 9913
rect 3861 9909 3863 9913
rect 3855 9908 3863 9909
rect 3855 9904 3857 9908
rect 3861 9904 3863 9908
rect 3855 9903 3863 9904
rect 3855 9899 3857 9903
rect 3861 9899 3863 9903
rect 3855 9898 3863 9899
rect 3855 9894 3857 9898
rect 3861 9894 3863 9898
rect 3855 9893 3863 9894
rect 3855 9889 3857 9893
rect 3861 9889 3863 9893
rect 3855 9888 3863 9889
rect 3855 9884 3857 9888
rect 3861 9884 3863 9888
rect 3855 9883 3863 9884
rect 3855 9879 3857 9883
rect 3861 9879 3863 9883
rect 3855 9878 3863 9879
rect 3855 9874 3857 9878
rect 3861 9874 3863 9878
rect 3855 9873 3863 9874
rect 3855 9869 3857 9873
rect 3861 9869 3863 9873
rect 3855 9868 3863 9869
rect 3855 9864 3857 9868
rect 3861 9864 3863 9868
rect 3919 9949 3921 9953
rect 3925 9949 3927 9953
rect 3919 9948 3927 9949
rect 3919 9944 3921 9948
rect 3925 9944 3927 9948
rect 3919 9943 3927 9944
rect 3919 9939 3921 9943
rect 3925 9939 3927 9943
rect 3919 9938 3927 9939
rect 3919 9934 3921 9938
rect 3925 9934 3927 9938
rect 3919 9933 3927 9934
rect 3919 9929 3921 9933
rect 3925 9929 3927 9933
rect 3919 9928 3927 9929
rect 3919 9924 3921 9928
rect 3925 9924 3927 9928
rect 3919 9923 3927 9924
rect 3919 9919 3921 9923
rect 3925 9919 3927 9923
rect 3919 9918 3927 9919
rect 3919 9914 3921 9918
rect 3925 9914 3927 9918
rect 3919 9913 3927 9914
rect 3919 9909 3921 9913
rect 3925 9909 3927 9913
rect 3919 9908 3927 9909
rect 3919 9904 3921 9908
rect 3925 9904 3927 9908
rect 3919 9903 3927 9904
rect 3919 9899 3921 9903
rect 3925 9899 3927 9903
rect 3919 9898 3927 9899
rect 3919 9894 3921 9898
rect 3925 9894 3927 9898
rect 3919 9893 3927 9894
rect 3919 9889 3921 9893
rect 3925 9889 3927 9893
rect 3919 9888 3927 9889
rect 3919 9884 3921 9888
rect 3925 9884 3927 9888
rect 3919 9883 3927 9884
rect 3919 9879 3921 9883
rect 3925 9879 3927 9883
rect 3919 9878 3927 9879
rect 3919 9874 3921 9878
rect 3925 9874 3927 9878
rect 3919 9873 3927 9874
rect 3919 9869 3921 9873
rect 3925 9869 3927 9873
rect 3919 9868 3927 9869
rect 3919 9864 3921 9868
rect 3925 9864 3927 9868
rect 3855 9863 3863 9864
rect 3855 9859 3857 9863
rect 3861 9859 3863 9863
rect 3855 9858 3863 9859
rect 3919 9863 3927 9864
rect 3919 9859 3921 9863
rect 3925 9859 3927 9863
rect 3919 9858 3927 9859
rect 3855 9856 3927 9858
rect 3855 9852 3857 9856
rect 3861 9852 3864 9856
rect 3868 9852 3869 9856
rect 3873 9852 3874 9856
rect 3878 9852 3879 9856
rect 3883 9852 3884 9856
rect 3888 9852 3889 9856
rect 3893 9852 3894 9856
rect 3898 9852 3899 9856
rect 3903 9852 3904 9856
rect 3908 9852 3909 9856
rect 3913 9852 3914 9856
rect 3918 9852 3921 9856
rect 3925 9852 3927 9856
rect 3855 9850 3927 9852
rect 4003 9978 4099 9979
rect 4003 9974 4004 9978
rect 4008 9974 4009 9978
rect 4013 9974 4014 9978
rect 4018 9974 4019 9978
rect 4023 9974 4024 9978
rect 4028 9974 4029 9978
rect 4033 9974 4034 9978
rect 4038 9974 4039 9978
rect 4043 9974 4044 9978
rect 4048 9974 4049 9978
rect 4053 9974 4054 9978
rect 4058 9974 4059 9978
rect 4063 9974 4064 9978
rect 4068 9974 4069 9978
rect 4073 9974 4074 9978
rect 4078 9974 4079 9978
rect 4083 9974 4084 9978
rect 4088 9974 4089 9978
rect 4093 9974 4094 9978
rect 4098 9974 4099 9978
rect 4003 9973 4099 9974
rect 4003 9969 4004 9973
rect 4008 9969 4009 9973
rect 4003 9968 4009 9969
rect 4003 9964 4004 9968
rect 4008 9964 4009 9968
rect 4093 9969 4094 9973
rect 4098 9969 4099 9973
rect 4093 9968 4099 9969
rect 4003 9963 4009 9964
rect 4003 9959 4004 9963
rect 4008 9959 4009 9963
rect 4003 9958 4009 9959
rect 4003 9954 4004 9958
rect 4008 9954 4009 9958
rect 4003 9953 4009 9954
rect 4003 9949 4004 9953
rect 4008 9949 4009 9953
rect 4003 9948 4009 9949
rect 4003 9944 4004 9948
rect 4008 9944 4009 9948
rect 4003 9943 4009 9944
rect 4003 9939 4004 9943
rect 4008 9939 4009 9943
rect 4003 9938 4009 9939
rect 4003 9934 4004 9938
rect 4008 9934 4009 9938
rect 4003 9933 4009 9934
rect 4003 9929 4004 9933
rect 4008 9929 4009 9933
rect 4003 9928 4009 9929
rect 4003 9924 4004 9928
rect 4008 9924 4009 9928
rect 4003 9923 4009 9924
rect 4003 9919 4004 9923
rect 4008 9919 4009 9923
rect 4003 9918 4009 9919
rect 4003 9914 4004 9918
rect 4008 9914 4009 9918
rect 4003 9913 4009 9914
rect 4003 9909 4004 9913
rect 4008 9909 4009 9913
rect 4003 9908 4009 9909
rect 4003 9904 4004 9908
rect 4008 9904 4009 9908
rect 4003 9903 4009 9904
rect 4003 9899 4004 9903
rect 4008 9899 4009 9903
rect 4003 9898 4009 9899
rect 4003 9894 4004 9898
rect 4008 9894 4009 9898
rect 4003 9893 4009 9894
rect 4003 9889 4004 9893
rect 4008 9889 4009 9893
rect 4003 9888 4009 9889
rect 4003 9884 4004 9888
rect 4008 9884 4009 9888
rect 4003 9883 4009 9884
rect 4003 9879 4004 9883
rect 4008 9879 4009 9883
rect 4003 9878 4009 9879
rect 4003 9874 4004 9878
rect 4008 9874 4009 9878
rect 4003 9873 4009 9874
rect 4003 9869 4004 9873
rect 4008 9869 4009 9873
rect 4003 9868 4009 9869
rect 4003 9864 4004 9868
rect 4008 9864 4009 9868
rect 4003 9863 4009 9864
rect 4003 9859 4004 9863
rect 4008 9859 4009 9863
rect 4003 9858 4009 9859
rect 4003 9854 4004 9858
rect 4008 9854 4009 9858
rect 4003 9853 4009 9854
rect 4003 9849 4004 9853
rect 4008 9849 4009 9853
rect 4093 9964 4094 9968
rect 4098 9964 4099 9968
rect 4093 9963 4099 9964
rect 4093 9959 4094 9963
rect 4098 9959 4099 9963
rect 4093 9958 4099 9959
rect 4093 9954 4094 9958
rect 4098 9954 4099 9958
rect 4093 9953 4099 9954
rect 4093 9949 4094 9953
rect 4098 9949 4099 9953
rect 4093 9948 4099 9949
rect 4093 9944 4094 9948
rect 4098 9944 4099 9948
rect 4093 9943 4099 9944
rect 4093 9939 4094 9943
rect 4098 9939 4099 9943
rect 4093 9938 4099 9939
rect 4093 9934 4094 9938
rect 4098 9934 4099 9938
rect 4093 9933 4099 9934
rect 4093 9929 4094 9933
rect 4098 9929 4099 9933
rect 4093 9928 4099 9929
rect 4093 9924 4094 9928
rect 4098 9924 4099 9928
rect 4093 9923 4099 9924
rect 4093 9919 4094 9923
rect 4098 9919 4099 9923
rect 4093 9918 4099 9919
rect 4093 9914 4094 9918
rect 4098 9914 4099 9918
rect 4093 9913 4099 9914
rect 4093 9909 4094 9913
rect 4098 9909 4099 9913
rect 4093 9908 4099 9909
rect 4093 9904 4094 9908
rect 4098 9904 4099 9908
rect 4093 9903 4099 9904
rect 4093 9899 4094 9903
rect 4098 9899 4099 9903
rect 4093 9898 4099 9899
rect 4093 9894 4094 9898
rect 4098 9894 4099 9898
rect 4093 9893 4099 9894
rect 4093 9889 4094 9893
rect 4098 9889 4099 9893
rect 4093 9888 4099 9889
rect 4093 9884 4094 9888
rect 4098 9884 4099 9888
rect 4093 9883 4099 9884
rect 4093 9879 4094 9883
rect 4098 9879 4099 9883
rect 4093 9878 4099 9879
rect 4093 9874 4094 9878
rect 4098 9874 4099 9878
rect 4093 9873 4099 9874
rect 4093 9869 4094 9873
rect 4098 9869 4099 9873
rect 4093 9868 4099 9869
rect 4093 9864 4094 9868
rect 4098 9864 4099 9868
rect 4093 9863 4099 9864
rect 4093 9859 4094 9863
rect 4098 9859 4099 9863
rect 4093 9858 4099 9859
rect 4093 9854 4094 9858
rect 4098 9854 4099 9858
rect 4093 9853 4099 9854
rect 4003 9848 4009 9849
rect 4003 9844 4004 9848
rect 4008 9844 4009 9848
rect 4093 9849 4094 9853
rect 4098 9849 4099 9853
rect 4093 9848 4099 9849
rect 4093 9844 4094 9848
rect 4098 9844 4099 9848
rect 4003 9843 4099 9844
rect 4003 9839 4004 9843
rect 4008 9839 4009 9843
rect 4013 9839 4014 9843
rect 4018 9839 4019 9843
rect 4023 9839 4024 9843
rect 4028 9839 4029 9843
rect 4033 9839 4034 9843
rect 4038 9839 4039 9843
rect 4043 9839 4044 9843
rect 4048 9839 4049 9843
rect 4053 9839 4054 9843
rect 4058 9839 4059 9843
rect 4063 9839 4064 9843
rect 4068 9839 4069 9843
rect 4073 9839 4074 9843
rect 4078 9839 4079 9843
rect 4083 9839 4084 9843
rect 4088 9839 4089 9843
rect 4093 9839 4094 9843
rect 4098 9839 4099 9843
rect 4003 9838 4099 9839
rect 655 9720 4517 9724
rect 655 9716 802 9720
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 821 9716 831 9720
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 850 9716 860 9720
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 879 9716 889 9720
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 908 9716 918 9720
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 937 9716 1319 9720
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1338 9716 1628 9720
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1647 9716 1937 9720
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1956 9716 2246 9720
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2265 9716 2555 9720
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2574 9716 2864 9720
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2883 9716 3173 9720
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3192 9716 3482 9720
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3501 9716 3791 9720
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3810 9716 4100 9720
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4119 9716 4292 9720
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4311 9716 4318 9720
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4337 9716 4344 9720
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4363 9716 4370 9720
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4389 9716 4396 9720
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4415 9716 4517 9720
rect 655 9710 4517 9716
rect 655 9706 802 9710
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 821 9706 831 9710
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 850 9706 860 9710
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 879 9706 889 9710
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 908 9706 918 9710
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 937 9706 1319 9710
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1338 9706 1628 9710
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1647 9706 1937 9710
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1956 9706 2246 9710
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2265 9706 2555 9710
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2574 9706 2864 9710
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2883 9706 3173 9710
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3192 9706 3482 9710
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3501 9706 3791 9710
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3810 9706 4100 9710
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4119 9706 4292 9710
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4311 9706 4318 9710
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4337 9706 4344 9710
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4363 9706 4370 9710
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4389 9706 4396 9710
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4415 9706 4517 9710
rect 655 9700 4517 9706
rect 655 9696 802 9700
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 821 9696 831 9700
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 850 9696 860 9700
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 879 9696 889 9700
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 908 9696 918 9700
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 937 9696 1319 9700
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1338 9696 1628 9700
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1647 9696 1937 9700
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1956 9696 2246 9700
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2265 9696 2555 9700
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2574 9696 2864 9700
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2883 9696 3173 9700
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3192 9696 3482 9700
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3501 9696 3791 9700
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3810 9696 4100 9700
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4119 9696 4292 9700
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4311 9696 4318 9700
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4337 9696 4344 9700
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4363 9696 4370 9700
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4389 9696 4396 9700
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4415 9696 4517 9700
rect 655 9690 4517 9696
rect 655 9686 802 9690
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 821 9686 831 9690
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 850 9686 860 9690
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 879 9686 889 9690
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 908 9686 918 9690
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 937 9686 1319 9690
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1338 9686 1628 9690
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1647 9686 1937 9690
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 1956 9686 2246 9690
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2265 9686 2555 9690
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2574 9686 2864 9690
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 2883 9686 3173 9690
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3192 9686 3482 9690
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 3501 9686 3791 9690
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 3810 9686 4100 9690
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4119 9686 4292 9690
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4311 9686 4318 9690
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4337 9686 4344 9690
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4363 9686 4370 9690
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4389 9686 4396 9690
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 4415 9686 4517 9690
rect 655 9684 4517 9686
rect 655 9622 695 9684
rect 655 9618 659 9622
rect 663 9618 669 9622
rect 673 9618 679 9622
rect 683 9618 689 9622
rect 693 9618 695 9622
rect 655 9617 695 9618
rect 655 9613 659 9617
rect 663 9613 669 9617
rect 673 9613 679 9617
rect 683 9613 689 9617
rect 693 9613 695 9617
rect 655 9612 695 9613
rect 655 9608 659 9612
rect 663 9608 669 9612
rect 673 9608 679 9612
rect 683 9608 689 9612
rect 693 9608 695 9612
rect 655 9607 695 9608
rect 655 9603 659 9607
rect 663 9603 669 9607
rect 673 9603 679 9607
rect 683 9603 689 9607
rect 693 9603 695 9607
rect 655 9596 695 9603
rect 655 9592 659 9596
rect 663 9592 669 9596
rect 673 9592 679 9596
rect 683 9592 689 9596
rect 693 9592 695 9596
rect 655 9591 695 9592
rect 655 9587 659 9591
rect 663 9587 669 9591
rect 673 9587 679 9591
rect 683 9587 689 9591
rect 693 9587 695 9591
rect 655 9586 695 9587
rect 655 9582 659 9586
rect 663 9582 669 9586
rect 673 9582 679 9586
rect 683 9582 689 9586
rect 693 9582 695 9586
rect 655 9581 695 9582
rect 655 9577 659 9581
rect 663 9577 669 9581
rect 673 9577 679 9581
rect 683 9577 689 9581
rect 693 9577 695 9581
rect 655 9570 695 9577
rect 655 9566 659 9570
rect 663 9566 669 9570
rect 673 9566 679 9570
rect 683 9566 689 9570
rect 693 9566 695 9570
rect 655 9565 695 9566
rect 655 9561 659 9565
rect 663 9561 669 9565
rect 673 9561 679 9565
rect 683 9561 689 9565
rect 693 9561 695 9565
rect 655 9560 695 9561
rect 655 9556 659 9560
rect 663 9556 669 9560
rect 673 9556 679 9560
rect 683 9556 689 9560
rect 693 9556 695 9560
rect 655 9555 695 9556
rect 655 9551 659 9555
rect 663 9551 669 9555
rect 673 9551 679 9555
rect 683 9551 689 9555
rect 693 9551 695 9555
rect 655 9544 695 9551
rect 655 9540 659 9544
rect 663 9540 669 9544
rect 673 9540 679 9544
rect 683 9540 689 9544
rect 693 9540 695 9544
rect 655 9539 695 9540
rect 655 9535 659 9539
rect 663 9535 669 9539
rect 673 9535 679 9539
rect 683 9535 689 9539
rect 693 9535 695 9539
rect 655 9534 695 9535
rect 655 9530 659 9534
rect 663 9530 669 9534
rect 673 9530 679 9534
rect 683 9530 689 9534
rect 693 9530 695 9534
rect 655 9529 695 9530
rect 655 9525 659 9529
rect 663 9525 669 9529
rect 673 9525 679 9529
rect 683 9525 689 9529
rect 693 9525 695 9529
rect 655 9518 695 9525
rect 655 9514 659 9518
rect 663 9514 669 9518
rect 673 9514 679 9518
rect 683 9514 689 9518
rect 693 9514 695 9518
rect 655 9513 695 9514
rect 655 9509 659 9513
rect 663 9509 669 9513
rect 673 9509 679 9513
rect 683 9509 689 9513
rect 693 9509 695 9513
rect 655 9508 695 9509
rect 655 9504 659 9508
rect 663 9504 669 9508
rect 673 9504 679 9508
rect 683 9504 689 9508
rect 693 9504 695 9508
rect 655 9503 695 9504
rect 655 9499 659 9503
rect 663 9499 669 9503
rect 673 9499 679 9503
rect 683 9499 689 9503
rect 693 9499 695 9503
rect 655 9325 695 9499
rect 4477 9577 4517 9684
rect 4477 9573 4479 9577
rect 4483 9573 4489 9577
rect 4493 9573 4499 9577
rect 4503 9573 4509 9577
rect 4513 9573 4517 9577
rect 4477 9572 4517 9573
rect 4477 9568 4479 9572
rect 4483 9568 4489 9572
rect 4493 9568 4499 9572
rect 4503 9568 4509 9572
rect 4513 9568 4517 9572
rect 4477 9567 4517 9568
rect 4477 9563 4479 9567
rect 4483 9563 4489 9567
rect 4493 9563 4499 9567
rect 4503 9563 4509 9567
rect 4513 9563 4517 9567
rect 4477 9562 4517 9563
rect 4477 9558 4479 9562
rect 4483 9558 4489 9562
rect 4493 9558 4499 9562
rect 4503 9558 4509 9562
rect 4513 9558 4517 9562
rect 4477 9548 4517 9558
rect 4477 9544 4479 9548
rect 4483 9544 4489 9548
rect 4493 9544 4499 9548
rect 4503 9544 4509 9548
rect 4513 9544 4517 9548
rect 4477 9543 4517 9544
rect 4477 9539 4479 9543
rect 4483 9539 4489 9543
rect 4493 9539 4499 9543
rect 4503 9539 4509 9543
rect 4513 9539 4517 9543
rect 4477 9538 4517 9539
rect 4477 9534 4479 9538
rect 4483 9534 4489 9538
rect 4493 9534 4499 9538
rect 4503 9534 4509 9538
rect 4513 9534 4517 9538
rect 4477 9533 4517 9534
rect 4477 9529 4479 9533
rect 4483 9529 4489 9533
rect 4493 9529 4499 9533
rect 4503 9529 4509 9533
rect 4513 9529 4517 9533
rect 4477 9519 4517 9529
rect 4477 9515 4479 9519
rect 4483 9515 4489 9519
rect 4493 9515 4499 9519
rect 4503 9515 4509 9519
rect 4513 9515 4517 9519
rect 4477 9514 4517 9515
rect 4477 9510 4479 9514
rect 4483 9510 4489 9514
rect 4493 9510 4499 9514
rect 4503 9510 4509 9514
rect 4513 9510 4517 9514
rect 4477 9509 4517 9510
rect 4477 9505 4479 9509
rect 4483 9505 4489 9509
rect 4493 9505 4499 9509
rect 4503 9505 4509 9509
rect 4513 9505 4517 9509
rect 4477 9504 4517 9505
rect 4477 9500 4479 9504
rect 4483 9500 4489 9504
rect 4493 9500 4499 9504
rect 4503 9500 4509 9504
rect 4513 9500 4517 9504
rect 4477 9490 4517 9500
rect 4477 9486 4479 9490
rect 4483 9486 4489 9490
rect 4493 9486 4499 9490
rect 4503 9486 4509 9490
rect 4513 9486 4517 9490
rect 4477 9485 4517 9486
rect 4477 9481 4479 9485
rect 4483 9481 4489 9485
rect 4493 9481 4499 9485
rect 4503 9481 4509 9485
rect 4513 9481 4517 9485
rect 4477 9480 4517 9481
rect 4477 9476 4479 9480
rect 4483 9476 4489 9480
rect 4493 9476 4499 9480
rect 4503 9476 4509 9480
rect 4513 9476 4517 9480
rect 4477 9475 4517 9476
rect 4477 9471 4479 9475
rect 4483 9471 4489 9475
rect 4493 9471 4499 9475
rect 4503 9471 4509 9475
rect 4513 9471 4517 9475
rect 4477 9461 4517 9471
rect 4477 9457 4479 9461
rect 4483 9457 4489 9461
rect 4493 9457 4499 9461
rect 4503 9457 4509 9461
rect 4513 9457 4517 9461
rect 4477 9456 4517 9457
rect 4477 9452 4479 9456
rect 4483 9452 4489 9456
rect 4493 9452 4499 9456
rect 4503 9452 4509 9456
rect 4513 9452 4517 9456
rect 4477 9451 4517 9452
rect 4477 9447 4479 9451
rect 4483 9447 4489 9451
rect 4493 9447 4499 9451
rect 4503 9447 4509 9451
rect 4513 9447 4517 9451
rect 4477 9446 4517 9447
rect 4477 9442 4479 9446
rect 4483 9442 4489 9446
rect 4493 9442 4499 9446
rect 4503 9442 4509 9446
rect 4513 9442 4517 9446
rect 655 9321 659 9325
rect 663 9321 669 9325
rect 673 9321 679 9325
rect 683 9321 689 9325
rect 693 9321 695 9325
rect 655 9320 695 9321
rect 655 9316 659 9320
rect 663 9316 669 9320
rect 673 9316 679 9320
rect 683 9316 689 9320
rect 693 9316 695 9320
rect 655 9315 695 9316
rect 655 9311 659 9315
rect 663 9311 669 9315
rect 673 9311 679 9315
rect 683 9311 689 9315
rect 693 9311 695 9315
rect 655 9310 695 9311
rect 655 9306 659 9310
rect 663 9306 669 9310
rect 673 9306 679 9310
rect 683 9306 689 9310
rect 693 9306 695 9310
rect 655 9016 695 9306
rect 4477 9060 4517 9442
rect 4477 9056 4479 9060
rect 4483 9056 4489 9060
rect 4493 9056 4499 9060
rect 4503 9056 4509 9060
rect 4513 9056 4517 9060
rect 4477 9055 4517 9056
rect 4477 9051 4479 9055
rect 4483 9051 4489 9055
rect 4493 9051 4499 9055
rect 4503 9051 4509 9055
rect 4513 9051 4517 9055
rect 4477 9050 4517 9051
rect 4477 9046 4479 9050
rect 4483 9046 4489 9050
rect 4493 9046 4499 9050
rect 4503 9046 4509 9050
rect 4513 9046 4517 9050
rect 4477 9045 4517 9046
rect 4477 9041 4479 9045
rect 4483 9041 4489 9045
rect 4493 9041 4499 9045
rect 4503 9041 4509 9045
rect 4513 9041 4517 9045
rect 655 9012 659 9016
rect 663 9012 669 9016
rect 673 9012 679 9016
rect 683 9012 689 9016
rect 693 9012 695 9016
rect 655 9011 695 9012
rect 655 9007 659 9011
rect 663 9007 669 9011
rect 673 9007 679 9011
rect 683 9007 689 9011
rect 693 9007 695 9011
rect 655 9006 695 9007
rect 655 9002 659 9006
rect 663 9002 669 9006
rect 673 9002 679 9006
rect 683 9002 689 9006
rect 693 9002 695 9006
rect 655 9001 695 9002
rect 655 8997 659 9001
rect 663 8997 669 9001
rect 673 8997 679 9001
rect 683 8997 689 9001
rect 693 8997 695 9001
rect 655 8707 695 8997
rect 4477 8751 4517 9041
rect 4477 8747 4479 8751
rect 4483 8747 4489 8751
rect 4493 8747 4499 8751
rect 4503 8747 4509 8751
rect 4513 8747 4517 8751
rect 4477 8746 4517 8747
rect 4477 8742 4479 8746
rect 4483 8742 4489 8746
rect 4493 8742 4499 8746
rect 4503 8742 4509 8746
rect 4513 8742 4517 8746
rect 4477 8741 4517 8742
rect 4477 8737 4479 8741
rect 4483 8737 4489 8741
rect 4493 8737 4499 8741
rect 4503 8737 4509 8741
rect 4513 8737 4517 8741
rect 4477 8736 4517 8737
rect 4477 8732 4479 8736
rect 4483 8732 4489 8736
rect 4493 8732 4499 8736
rect 4503 8732 4509 8736
rect 4513 8732 4517 8736
rect 655 8703 659 8707
rect 663 8703 669 8707
rect 673 8703 679 8707
rect 683 8703 689 8707
rect 693 8703 695 8707
rect 655 8702 695 8703
rect 655 8698 659 8702
rect 663 8698 669 8702
rect 673 8698 679 8702
rect 683 8698 689 8702
rect 693 8698 695 8702
rect 655 8697 695 8698
rect 655 8693 659 8697
rect 663 8693 669 8697
rect 673 8693 679 8697
rect 683 8693 689 8697
rect 693 8693 695 8697
rect 655 8692 695 8693
rect 655 8688 659 8692
rect 663 8688 669 8692
rect 673 8688 679 8692
rect 683 8688 689 8692
rect 693 8688 695 8692
rect 655 8398 695 8688
rect 4477 8442 4517 8732
rect 4477 8438 4479 8442
rect 4483 8438 4489 8442
rect 4493 8438 4499 8442
rect 4503 8438 4509 8442
rect 4513 8438 4517 8442
rect 4477 8437 4517 8438
rect 4477 8433 4479 8437
rect 4483 8433 4489 8437
rect 4493 8433 4499 8437
rect 4503 8433 4509 8437
rect 4513 8433 4517 8437
rect 4477 8432 4517 8433
rect 4477 8428 4479 8432
rect 4483 8428 4489 8432
rect 4493 8428 4499 8432
rect 4503 8428 4509 8432
rect 4513 8428 4517 8432
rect 4477 8427 4517 8428
rect 4477 8423 4479 8427
rect 4483 8423 4489 8427
rect 4493 8423 4499 8427
rect 4503 8423 4509 8427
rect 4513 8423 4517 8427
rect 655 8394 659 8398
rect 663 8394 669 8398
rect 673 8394 679 8398
rect 683 8394 689 8398
rect 693 8394 695 8398
rect 655 8393 695 8394
rect 655 8389 659 8393
rect 663 8389 669 8393
rect 673 8389 679 8393
rect 683 8389 689 8393
rect 693 8389 695 8393
rect 655 8388 695 8389
rect 655 8384 659 8388
rect 663 8384 669 8388
rect 673 8384 679 8388
rect 683 8384 689 8388
rect 693 8384 695 8388
rect 655 8383 695 8384
rect 655 8379 659 8383
rect 663 8379 669 8383
rect 673 8379 679 8383
rect 683 8379 689 8383
rect 693 8379 695 8383
rect 655 8089 695 8379
rect 4477 8133 4517 8423
rect 4477 8129 4479 8133
rect 4483 8129 4489 8133
rect 4493 8129 4499 8133
rect 4503 8129 4509 8133
rect 4513 8129 4517 8133
rect 4477 8128 4517 8129
rect 4477 8124 4479 8128
rect 4483 8124 4489 8128
rect 4493 8124 4499 8128
rect 4503 8124 4509 8128
rect 4513 8124 4517 8128
rect 4477 8123 4517 8124
rect 4477 8119 4479 8123
rect 4483 8119 4489 8123
rect 4493 8119 4499 8123
rect 4503 8119 4509 8123
rect 4513 8119 4517 8123
rect 4477 8118 4517 8119
rect 4477 8114 4479 8118
rect 4483 8114 4489 8118
rect 4493 8114 4499 8118
rect 4503 8114 4509 8118
rect 4513 8114 4517 8118
rect 4477 8102 4517 8114
rect 4477 8098 4479 8102
rect 4483 8098 4489 8102
rect 4493 8098 4499 8102
rect 4503 8098 4509 8102
rect 4513 8098 4517 8102
rect 4477 8097 4517 8098
rect 655 8085 659 8089
rect 663 8085 669 8089
rect 673 8085 679 8089
rect 683 8085 689 8089
rect 693 8085 695 8089
rect 4477 8093 4479 8097
rect 4483 8093 4489 8097
rect 4493 8093 4499 8097
rect 4503 8093 4509 8097
rect 4513 8093 4517 8097
rect 4477 8092 4517 8093
rect 4477 8088 4479 8092
rect 4483 8088 4489 8092
rect 4493 8088 4499 8092
rect 4503 8088 4509 8092
rect 4513 8088 4517 8092
rect 4477 8087 4517 8088
rect 655 8084 695 8085
rect 655 8080 659 8084
rect 663 8080 669 8084
rect 673 8080 679 8084
rect 683 8080 689 8084
rect 693 8080 695 8084
rect 4477 8083 4479 8087
rect 4483 8083 4489 8087
rect 4493 8083 4499 8087
rect 4503 8083 4509 8087
rect 4513 8083 4517 8087
rect 655 8079 695 8080
rect 655 8075 659 8079
rect 663 8075 669 8079
rect 673 8075 679 8079
rect 683 8075 689 8079
rect 693 8075 695 8079
rect 655 8074 695 8075
rect 655 8070 659 8074
rect 663 8070 669 8074
rect 673 8070 679 8074
rect 683 8070 689 8074
rect 693 8070 695 8074
rect 655 7780 695 8070
rect 655 7776 659 7780
rect 663 7776 669 7780
rect 673 7776 679 7780
rect 683 7776 689 7780
rect 693 7776 695 7780
rect 655 7775 695 7776
rect 655 7771 659 7775
rect 663 7771 669 7775
rect 673 7771 679 7775
rect 683 7771 689 7775
rect 693 7771 695 7775
rect 655 7770 695 7771
rect 655 7766 659 7770
rect 663 7766 669 7770
rect 673 7766 679 7770
rect 683 7766 689 7770
rect 693 7766 695 7770
rect 655 7765 695 7766
rect 655 7761 659 7765
rect 663 7761 669 7765
rect 673 7761 679 7765
rect 683 7761 689 7765
rect 693 7761 695 7765
rect 655 7471 695 7761
rect 4477 7793 4517 8083
rect 4477 7789 4479 7793
rect 4483 7789 4489 7793
rect 4493 7789 4499 7793
rect 4503 7789 4509 7793
rect 4513 7789 4517 7793
rect 4477 7788 4517 7789
rect 4477 7784 4479 7788
rect 4483 7784 4489 7788
rect 4493 7784 4499 7788
rect 4503 7784 4509 7788
rect 4513 7784 4517 7788
rect 4477 7783 4517 7784
rect 4477 7779 4479 7783
rect 4483 7779 4489 7783
rect 4493 7779 4499 7783
rect 4503 7779 4509 7783
rect 4513 7779 4517 7783
rect 4477 7778 4517 7779
rect 4477 7774 4479 7778
rect 4483 7774 4489 7778
rect 4493 7774 4499 7778
rect 4503 7774 4509 7778
rect 4513 7774 4517 7778
rect 655 7467 659 7471
rect 663 7467 669 7471
rect 673 7467 679 7471
rect 683 7467 689 7471
rect 693 7467 695 7471
rect 655 7466 695 7467
rect 655 7462 659 7466
rect 663 7462 669 7466
rect 673 7462 679 7466
rect 683 7462 689 7466
rect 693 7462 695 7466
rect 655 7461 695 7462
rect 655 7457 659 7461
rect 663 7457 669 7461
rect 673 7457 679 7461
rect 683 7457 689 7461
rect 693 7457 695 7461
rect 655 7456 695 7457
rect 655 7452 659 7456
rect 663 7452 669 7456
rect 673 7452 679 7456
rect 683 7452 689 7456
rect 693 7452 695 7456
rect 655 7162 695 7452
rect 655 7158 659 7162
rect 663 7158 669 7162
rect 673 7158 679 7162
rect 683 7158 689 7162
rect 693 7158 695 7162
rect 655 7157 695 7158
rect 655 7153 659 7157
rect 663 7153 669 7157
rect 673 7153 679 7157
rect 683 7153 689 7157
rect 693 7153 695 7157
rect 655 7152 695 7153
rect 655 7148 659 7152
rect 663 7148 669 7152
rect 673 7148 679 7152
rect 683 7148 689 7152
rect 693 7148 695 7152
rect 655 7147 695 7148
rect 655 7143 659 7147
rect 663 7143 669 7147
rect 673 7143 679 7147
rect 683 7143 689 7147
rect 693 7143 695 7147
rect 655 6853 695 7143
rect 655 6849 659 6853
rect 663 6849 669 6853
rect 673 6849 679 6853
rect 683 6849 689 6853
rect 693 6849 695 6853
rect 655 6848 695 6849
rect 655 6844 659 6848
rect 663 6844 669 6848
rect 673 6844 679 6848
rect 683 6844 689 6848
rect 693 6844 695 6848
rect 655 6843 695 6844
rect 655 6839 659 6843
rect 663 6839 669 6843
rect 673 6839 679 6843
rect 683 6839 689 6843
rect 693 6839 695 6843
rect 655 6838 695 6839
rect 655 6834 659 6838
rect 663 6834 669 6838
rect 673 6834 679 6838
rect 683 6834 689 6838
rect 693 6834 695 6838
rect 655 6544 695 6834
rect 655 6540 659 6544
rect 663 6540 669 6544
rect 673 6540 679 6544
rect 683 6540 689 6544
rect 693 6540 695 6544
rect 655 6539 695 6540
rect 655 6535 659 6539
rect 663 6535 669 6539
rect 673 6535 679 6539
rect 683 6535 689 6539
rect 693 6535 695 6539
rect 655 6534 695 6535
rect 655 6530 659 6534
rect 663 6530 669 6534
rect 673 6530 679 6534
rect 683 6530 689 6534
rect 693 6530 695 6534
rect 655 6529 695 6530
rect 655 6525 659 6529
rect 663 6525 669 6529
rect 673 6525 679 6529
rect 683 6525 689 6529
rect 693 6525 695 6529
rect 655 6144 695 6525
rect 655 6140 659 6144
rect 663 6140 669 6144
rect 673 6140 679 6144
rect 683 6140 689 6144
rect 693 6140 695 6144
rect 655 6139 695 6140
rect 655 6135 659 6139
rect 663 6135 669 6139
rect 673 6135 679 6139
rect 683 6135 689 6139
rect 693 6135 695 6139
rect 655 6134 695 6135
rect 655 6130 659 6134
rect 663 6130 669 6134
rect 673 6130 679 6134
rect 683 6130 689 6134
rect 693 6130 695 6134
rect 655 6129 695 6130
rect 655 6125 659 6129
rect 663 6125 669 6129
rect 673 6125 679 6129
rect 683 6125 689 6129
rect 693 6125 695 6129
rect 655 6115 695 6125
rect 655 6111 659 6115
rect 663 6111 669 6115
rect 673 6111 679 6115
rect 683 6111 689 6115
rect 693 6111 695 6115
rect 655 6110 695 6111
rect 655 6106 659 6110
rect 663 6106 669 6110
rect 673 6106 679 6110
rect 683 6106 689 6110
rect 693 6106 695 6110
rect 655 6105 695 6106
rect 655 6101 659 6105
rect 663 6101 669 6105
rect 673 6101 679 6105
rect 683 6101 689 6105
rect 693 6101 695 6105
rect 655 6100 695 6101
rect 655 6096 659 6100
rect 663 6096 669 6100
rect 673 6096 679 6100
rect 683 6096 689 6100
rect 693 6096 695 6100
rect 655 6086 695 6096
rect 655 6082 659 6086
rect 663 6082 669 6086
rect 673 6082 679 6086
rect 683 6082 689 6086
rect 693 6082 695 6086
rect 655 6081 695 6082
rect 655 6077 659 6081
rect 663 6077 669 6081
rect 673 6077 679 6081
rect 683 6077 689 6081
rect 693 6077 695 6081
rect 655 6076 695 6077
rect 655 6072 659 6076
rect 663 6072 669 6076
rect 673 6072 679 6076
rect 683 6072 689 6076
rect 693 6072 695 6076
rect 655 6071 695 6072
rect 655 6067 659 6071
rect 663 6067 669 6071
rect 673 6067 679 6071
rect 683 6067 689 6071
rect 693 6067 695 6071
rect 655 6057 695 6067
rect 655 6053 659 6057
rect 663 6053 669 6057
rect 673 6053 679 6057
rect 683 6053 689 6057
rect 693 6053 695 6057
rect 655 6052 695 6053
rect 655 6048 659 6052
rect 663 6048 669 6052
rect 673 6048 679 6052
rect 683 6048 689 6052
rect 693 6048 695 6052
rect 655 6047 695 6048
rect 655 6043 659 6047
rect 663 6043 669 6047
rect 673 6043 679 6047
rect 683 6043 689 6047
rect 693 6043 695 6047
rect 655 6042 695 6043
rect 655 6038 659 6042
rect 663 6038 669 6042
rect 673 6038 679 6042
rect 683 6038 689 6042
rect 693 6038 695 6042
rect 655 6028 695 6038
rect 655 6024 659 6028
rect 663 6024 669 6028
rect 673 6024 679 6028
rect 683 6024 689 6028
rect 693 6024 695 6028
rect 655 6023 695 6024
rect 655 6019 659 6023
rect 663 6019 669 6023
rect 673 6019 679 6023
rect 683 6019 689 6023
rect 693 6019 695 6023
rect 655 6018 695 6019
rect 655 6014 659 6018
rect 663 6014 669 6018
rect 673 6014 679 6018
rect 683 6014 689 6018
rect 693 6014 695 6018
rect 655 6013 695 6014
rect 655 6009 659 6013
rect 663 6009 669 6013
rect 673 6009 679 6013
rect 683 6009 689 6013
rect 693 6009 695 6013
rect 655 5902 695 6009
rect 4477 7206 4517 7774
rect 4477 7202 4479 7206
rect 4483 7202 4489 7206
rect 4493 7202 4499 7206
rect 4503 7202 4509 7206
rect 4513 7202 4517 7206
rect 4477 7201 4517 7202
rect 4477 7197 4479 7201
rect 4483 7197 4489 7201
rect 4493 7197 4499 7201
rect 4503 7197 4509 7201
rect 4513 7197 4517 7201
rect 4477 7196 4517 7197
rect 4477 7192 4479 7196
rect 4483 7192 4489 7196
rect 4493 7192 4499 7196
rect 4503 7192 4509 7196
rect 4513 7192 4517 7196
rect 4477 7191 4517 7192
rect 4477 7187 4479 7191
rect 4483 7187 4489 7191
rect 4493 7187 4499 7191
rect 4503 7187 4509 7191
rect 4513 7187 4517 7191
rect 4477 6897 4517 7187
rect 4477 6893 4479 6897
rect 4483 6893 4489 6897
rect 4493 6893 4499 6897
rect 4503 6893 4509 6897
rect 4513 6893 4517 6897
rect 4477 6892 4517 6893
rect 4477 6888 4479 6892
rect 4483 6888 4489 6892
rect 4493 6888 4499 6892
rect 4503 6888 4509 6892
rect 4513 6888 4517 6892
rect 4477 6887 4517 6888
rect 4477 6883 4479 6887
rect 4483 6883 4489 6887
rect 4493 6883 4499 6887
rect 4503 6883 4509 6887
rect 4513 6883 4517 6887
rect 4477 6882 4517 6883
rect 4477 6878 4479 6882
rect 4483 6878 4489 6882
rect 4493 6878 4499 6882
rect 4503 6878 4509 6882
rect 4513 6878 4517 6882
rect 4477 6588 4517 6878
rect 4477 6584 4479 6588
rect 4483 6584 4489 6588
rect 4493 6584 4499 6588
rect 4503 6584 4509 6588
rect 4513 6584 4517 6588
rect 4477 6583 4517 6584
rect 4477 6579 4479 6583
rect 4483 6579 4489 6583
rect 4493 6579 4499 6583
rect 4503 6579 4509 6583
rect 4513 6579 4517 6583
rect 4477 6578 4517 6579
rect 4477 6574 4479 6578
rect 4483 6574 4489 6578
rect 4493 6574 4499 6578
rect 4503 6574 4509 6578
rect 4513 6574 4517 6578
rect 4477 6573 4517 6574
rect 4477 6569 4479 6573
rect 4483 6569 4489 6573
rect 4493 6569 4499 6573
rect 4503 6569 4509 6573
rect 4513 6569 4517 6573
rect 4477 6279 4517 6569
rect 4477 6275 4479 6279
rect 4483 6275 4489 6279
rect 4493 6275 4499 6279
rect 4503 6275 4509 6279
rect 4513 6275 4517 6279
rect 4477 6274 4517 6275
rect 4477 6270 4479 6274
rect 4483 6270 4489 6274
rect 4493 6270 4499 6274
rect 4503 6270 4509 6274
rect 4513 6270 4517 6274
rect 4477 6269 4517 6270
rect 4477 6265 4479 6269
rect 4483 6265 4489 6269
rect 4493 6265 4499 6269
rect 4503 6265 4509 6269
rect 4513 6265 4517 6269
rect 4477 6264 4517 6265
rect 4477 6260 4479 6264
rect 4483 6260 4489 6264
rect 4493 6260 4499 6264
rect 4503 6260 4509 6264
rect 4513 6260 4517 6264
rect 4477 6087 4517 6260
rect 4477 6083 4479 6087
rect 4483 6083 4489 6087
rect 4493 6083 4499 6087
rect 4503 6083 4509 6087
rect 4513 6083 4517 6087
rect 4477 6082 4517 6083
rect 4477 6078 4479 6082
rect 4483 6078 4489 6082
rect 4493 6078 4499 6082
rect 4503 6078 4509 6082
rect 4513 6078 4517 6082
rect 4477 6077 4517 6078
rect 4477 6073 4479 6077
rect 4483 6073 4489 6077
rect 4493 6073 4499 6077
rect 4503 6073 4509 6077
rect 4513 6073 4517 6077
rect 4477 6072 4517 6073
rect 4477 6068 4479 6072
rect 4483 6068 4489 6072
rect 4493 6068 4499 6072
rect 4503 6068 4509 6072
rect 4513 6068 4517 6072
rect 4477 6061 4517 6068
rect 4477 6057 4479 6061
rect 4483 6057 4489 6061
rect 4493 6057 4499 6061
rect 4503 6057 4509 6061
rect 4513 6057 4517 6061
rect 4477 6056 4517 6057
rect 4477 6052 4479 6056
rect 4483 6052 4489 6056
rect 4493 6052 4499 6056
rect 4503 6052 4509 6056
rect 4513 6052 4517 6056
rect 4477 6051 4517 6052
rect 4477 6047 4479 6051
rect 4483 6047 4489 6051
rect 4493 6047 4499 6051
rect 4503 6047 4509 6051
rect 4513 6047 4517 6051
rect 4477 6046 4517 6047
rect 4477 6042 4479 6046
rect 4483 6042 4489 6046
rect 4493 6042 4499 6046
rect 4503 6042 4509 6046
rect 4513 6042 4517 6046
rect 4477 6035 4517 6042
rect 4477 6031 4479 6035
rect 4483 6031 4489 6035
rect 4493 6031 4499 6035
rect 4503 6031 4509 6035
rect 4513 6031 4517 6035
rect 4477 6030 4517 6031
rect 4477 6026 4479 6030
rect 4483 6026 4489 6030
rect 4493 6026 4499 6030
rect 4503 6026 4509 6030
rect 4513 6026 4517 6030
rect 4477 6025 4517 6026
rect 4477 6021 4479 6025
rect 4483 6021 4489 6025
rect 4493 6021 4499 6025
rect 4503 6021 4509 6025
rect 4513 6021 4517 6025
rect 4477 6020 4517 6021
rect 4477 6016 4479 6020
rect 4483 6016 4489 6020
rect 4493 6016 4499 6020
rect 4503 6016 4509 6020
rect 4513 6016 4517 6020
rect 4477 6009 4517 6016
rect 4477 6005 4479 6009
rect 4483 6005 4489 6009
rect 4493 6005 4499 6009
rect 4503 6005 4509 6009
rect 4513 6005 4517 6009
rect 4477 6004 4517 6005
rect 4477 6000 4479 6004
rect 4483 6000 4489 6004
rect 4493 6000 4499 6004
rect 4503 6000 4509 6004
rect 4513 6000 4517 6004
rect 4477 5999 4517 6000
rect 4477 5995 4479 5999
rect 4483 5995 4489 5999
rect 4493 5995 4499 5999
rect 4503 5995 4509 5999
rect 4513 5995 4517 5999
rect 4477 5994 4517 5995
rect 4477 5990 4479 5994
rect 4483 5990 4489 5994
rect 4493 5990 4499 5994
rect 4503 5990 4509 5994
rect 4513 5990 4517 5994
rect 4477 5983 4517 5990
rect 4477 5979 4479 5983
rect 4483 5979 4489 5983
rect 4493 5979 4499 5983
rect 4503 5979 4509 5983
rect 4513 5979 4517 5983
rect 4477 5978 4517 5979
rect 4477 5974 4479 5978
rect 4483 5974 4489 5978
rect 4493 5974 4499 5978
rect 4503 5974 4509 5978
rect 4513 5974 4517 5978
rect 4477 5973 4517 5974
rect 4477 5969 4479 5973
rect 4483 5969 4489 5973
rect 4493 5969 4499 5973
rect 4503 5969 4509 5973
rect 4513 5969 4517 5973
rect 4477 5968 4517 5969
rect 4477 5964 4479 5968
rect 4483 5964 4489 5968
rect 4493 5964 4499 5968
rect 4503 5964 4509 5968
rect 4513 5964 4517 5968
rect 4477 5902 4517 5964
rect 655 5900 4517 5902
rect 655 5896 757 5900
rect 761 5896 762 5900
rect 766 5896 767 5900
rect 771 5896 772 5900
rect 776 5896 783 5900
rect 787 5896 788 5900
rect 792 5896 793 5900
rect 797 5896 798 5900
rect 802 5896 809 5900
rect 813 5896 814 5900
rect 818 5896 819 5900
rect 823 5896 824 5900
rect 828 5896 835 5900
rect 839 5896 840 5900
rect 844 5896 845 5900
rect 849 5896 850 5900
rect 854 5896 861 5900
rect 865 5896 866 5900
rect 870 5896 871 5900
rect 875 5896 876 5900
rect 880 5896 1054 5900
rect 1058 5896 1059 5900
rect 1063 5896 1064 5900
rect 1068 5896 1069 5900
rect 1073 5896 1363 5900
rect 1367 5896 1368 5900
rect 1372 5896 1373 5900
rect 1377 5896 1378 5900
rect 1382 5896 1672 5900
rect 1676 5896 1677 5900
rect 1681 5896 1682 5900
rect 1686 5896 1687 5900
rect 1691 5896 1981 5900
rect 1985 5896 1986 5900
rect 1990 5896 1991 5900
rect 1995 5896 1996 5900
rect 2000 5896 2290 5900
rect 2294 5896 2295 5900
rect 2299 5896 2300 5900
rect 2304 5896 2305 5900
rect 2309 5896 2599 5900
rect 2603 5896 2604 5900
rect 2608 5896 2609 5900
rect 2613 5896 2614 5900
rect 2618 5896 2908 5900
rect 2912 5896 2913 5900
rect 2917 5896 2918 5900
rect 2922 5896 2923 5900
rect 2927 5896 3217 5900
rect 3221 5896 3222 5900
rect 3226 5896 3227 5900
rect 3231 5896 3232 5900
rect 3236 5896 3526 5900
rect 3530 5896 3531 5900
rect 3535 5896 3536 5900
rect 3540 5896 3541 5900
rect 3545 5896 3835 5900
rect 3839 5896 3840 5900
rect 3844 5896 3845 5900
rect 3849 5896 3850 5900
rect 3854 5896 4235 5900
rect 4239 5896 4240 5900
rect 4244 5896 4245 5900
rect 4249 5896 4250 5900
rect 4254 5896 4264 5900
rect 4268 5896 4269 5900
rect 4273 5896 4274 5900
rect 4278 5896 4279 5900
rect 4283 5896 4293 5900
rect 4297 5896 4298 5900
rect 4302 5896 4303 5900
rect 4307 5896 4308 5900
rect 4312 5896 4322 5900
rect 4326 5896 4327 5900
rect 4331 5896 4332 5900
rect 4336 5896 4337 5900
rect 4341 5896 4351 5900
rect 4355 5896 4356 5900
rect 4360 5896 4361 5900
rect 4365 5896 4366 5900
rect 4370 5896 4517 5900
rect 655 5890 4517 5896
rect 655 5886 757 5890
rect 761 5886 762 5890
rect 766 5886 767 5890
rect 771 5886 772 5890
rect 776 5886 783 5890
rect 787 5886 788 5890
rect 792 5886 793 5890
rect 797 5886 798 5890
rect 802 5886 809 5890
rect 813 5886 814 5890
rect 818 5886 819 5890
rect 823 5886 824 5890
rect 828 5886 835 5890
rect 839 5886 840 5890
rect 844 5886 845 5890
rect 849 5886 850 5890
rect 854 5886 861 5890
rect 865 5886 866 5890
rect 870 5886 871 5890
rect 875 5886 876 5890
rect 880 5886 1054 5890
rect 1058 5886 1059 5890
rect 1063 5886 1064 5890
rect 1068 5886 1069 5890
rect 1073 5886 1363 5890
rect 1367 5886 1368 5890
rect 1372 5886 1373 5890
rect 1377 5886 1378 5890
rect 1382 5886 1672 5890
rect 1676 5886 1677 5890
rect 1681 5886 1682 5890
rect 1686 5886 1687 5890
rect 1691 5886 1981 5890
rect 1985 5886 1986 5890
rect 1990 5886 1991 5890
rect 1995 5886 1996 5890
rect 2000 5886 2290 5890
rect 2294 5886 2295 5890
rect 2299 5886 2300 5890
rect 2304 5886 2305 5890
rect 2309 5886 2599 5890
rect 2603 5886 2604 5890
rect 2608 5886 2609 5890
rect 2613 5886 2614 5890
rect 2618 5886 2908 5890
rect 2912 5886 2913 5890
rect 2917 5886 2918 5890
rect 2922 5886 2923 5890
rect 2927 5886 3217 5890
rect 3221 5886 3222 5890
rect 3226 5886 3227 5890
rect 3231 5886 3232 5890
rect 3236 5886 3526 5890
rect 3530 5886 3531 5890
rect 3535 5886 3536 5890
rect 3540 5886 3541 5890
rect 3545 5886 3835 5890
rect 3839 5886 3840 5890
rect 3844 5886 3845 5890
rect 3849 5886 3850 5890
rect 3854 5886 4235 5890
rect 4239 5886 4240 5890
rect 4244 5886 4245 5890
rect 4249 5886 4250 5890
rect 4254 5886 4264 5890
rect 4268 5886 4269 5890
rect 4273 5886 4274 5890
rect 4278 5886 4279 5890
rect 4283 5886 4293 5890
rect 4297 5886 4298 5890
rect 4302 5886 4303 5890
rect 4307 5886 4308 5890
rect 4312 5886 4322 5890
rect 4326 5886 4327 5890
rect 4331 5886 4332 5890
rect 4336 5886 4337 5890
rect 4341 5886 4351 5890
rect 4355 5886 4356 5890
rect 4360 5886 4361 5890
rect 4365 5886 4366 5890
rect 4370 5886 4517 5890
rect 655 5880 4517 5886
rect 655 5876 757 5880
rect 761 5876 762 5880
rect 766 5876 767 5880
rect 771 5876 772 5880
rect 776 5876 783 5880
rect 787 5876 788 5880
rect 792 5876 793 5880
rect 797 5876 798 5880
rect 802 5876 809 5880
rect 813 5876 814 5880
rect 818 5876 819 5880
rect 823 5876 824 5880
rect 828 5876 835 5880
rect 839 5876 840 5880
rect 844 5876 845 5880
rect 849 5876 850 5880
rect 854 5876 861 5880
rect 865 5876 866 5880
rect 870 5876 871 5880
rect 875 5876 876 5880
rect 880 5876 1054 5880
rect 1058 5876 1059 5880
rect 1063 5876 1064 5880
rect 1068 5876 1069 5880
rect 1073 5876 1363 5880
rect 1367 5876 1368 5880
rect 1372 5876 1373 5880
rect 1377 5876 1378 5880
rect 1382 5876 1672 5880
rect 1676 5876 1677 5880
rect 1681 5876 1682 5880
rect 1686 5876 1687 5880
rect 1691 5876 1981 5880
rect 1985 5876 1986 5880
rect 1990 5876 1991 5880
rect 1995 5876 1996 5880
rect 2000 5876 2290 5880
rect 2294 5876 2295 5880
rect 2299 5876 2300 5880
rect 2304 5876 2305 5880
rect 2309 5876 2599 5880
rect 2603 5876 2604 5880
rect 2608 5876 2609 5880
rect 2613 5876 2614 5880
rect 2618 5876 2908 5880
rect 2912 5876 2913 5880
rect 2917 5876 2918 5880
rect 2922 5876 2923 5880
rect 2927 5876 3217 5880
rect 3221 5876 3222 5880
rect 3226 5876 3227 5880
rect 3231 5876 3232 5880
rect 3236 5876 3526 5880
rect 3530 5876 3531 5880
rect 3535 5876 3536 5880
rect 3540 5876 3541 5880
rect 3545 5876 3835 5880
rect 3839 5876 3840 5880
rect 3844 5876 3845 5880
rect 3849 5876 3850 5880
rect 3854 5876 4235 5880
rect 4239 5876 4240 5880
rect 4244 5876 4245 5880
rect 4249 5876 4250 5880
rect 4254 5876 4264 5880
rect 4268 5876 4269 5880
rect 4273 5876 4274 5880
rect 4278 5876 4279 5880
rect 4283 5876 4293 5880
rect 4297 5876 4298 5880
rect 4302 5876 4303 5880
rect 4307 5876 4308 5880
rect 4312 5876 4322 5880
rect 4326 5876 4327 5880
rect 4331 5876 4332 5880
rect 4336 5876 4337 5880
rect 4341 5876 4351 5880
rect 4355 5876 4356 5880
rect 4360 5876 4361 5880
rect 4365 5876 4366 5880
rect 4370 5876 4517 5880
rect 655 5870 4517 5876
rect 655 5866 757 5870
rect 761 5866 762 5870
rect 766 5866 767 5870
rect 771 5866 772 5870
rect 776 5866 783 5870
rect 787 5866 788 5870
rect 792 5866 793 5870
rect 797 5866 798 5870
rect 802 5866 809 5870
rect 813 5866 814 5870
rect 818 5866 819 5870
rect 823 5866 824 5870
rect 828 5866 835 5870
rect 839 5866 840 5870
rect 844 5866 845 5870
rect 849 5866 850 5870
rect 854 5866 861 5870
rect 865 5866 866 5870
rect 870 5866 871 5870
rect 875 5866 876 5870
rect 880 5866 1054 5870
rect 1058 5866 1059 5870
rect 1063 5866 1064 5870
rect 1068 5866 1069 5870
rect 1073 5866 1363 5870
rect 1367 5866 1368 5870
rect 1372 5866 1373 5870
rect 1377 5866 1378 5870
rect 1382 5866 1672 5870
rect 1676 5866 1677 5870
rect 1681 5866 1682 5870
rect 1686 5866 1687 5870
rect 1691 5866 1981 5870
rect 1985 5866 1986 5870
rect 1990 5866 1991 5870
rect 1995 5866 1996 5870
rect 2000 5866 2290 5870
rect 2294 5866 2295 5870
rect 2299 5866 2300 5870
rect 2304 5866 2305 5870
rect 2309 5866 2599 5870
rect 2603 5866 2604 5870
rect 2608 5866 2609 5870
rect 2613 5866 2614 5870
rect 2618 5866 2908 5870
rect 2912 5866 2913 5870
rect 2917 5866 2918 5870
rect 2922 5866 2923 5870
rect 2927 5866 3217 5870
rect 3221 5866 3222 5870
rect 3226 5866 3227 5870
rect 3231 5866 3232 5870
rect 3236 5866 3526 5870
rect 3530 5866 3531 5870
rect 3535 5866 3536 5870
rect 3540 5866 3541 5870
rect 3545 5866 3835 5870
rect 3839 5866 3840 5870
rect 3844 5866 3845 5870
rect 3849 5866 3850 5870
rect 3854 5866 4235 5870
rect 4239 5866 4240 5870
rect 4244 5866 4245 5870
rect 4249 5866 4250 5870
rect 4254 5866 4264 5870
rect 4268 5866 4269 5870
rect 4273 5866 4274 5870
rect 4278 5866 4279 5870
rect 4283 5866 4293 5870
rect 4297 5866 4298 5870
rect 4302 5866 4303 5870
rect 4307 5866 4308 5870
rect 4312 5866 4322 5870
rect 4326 5866 4327 5870
rect 4331 5866 4332 5870
rect 4336 5866 4337 5870
rect 4341 5866 4351 5870
rect 4355 5866 4356 5870
rect 4360 5866 4361 5870
rect 4365 5866 4366 5870
rect 4370 5866 4517 5870
rect 655 5862 4517 5866
<< nsubstratendiff >>
rect 1371 9978 1467 9979
rect 1371 9974 1372 9978
rect 1376 9974 1377 9978
rect 1381 9974 1382 9978
rect 1386 9974 1387 9978
rect 1391 9974 1392 9978
rect 1396 9974 1397 9978
rect 1401 9974 1402 9978
rect 1406 9974 1407 9978
rect 1411 9974 1412 9978
rect 1416 9974 1417 9978
rect 1421 9974 1422 9978
rect 1426 9974 1427 9978
rect 1431 9974 1432 9978
rect 1436 9974 1437 9978
rect 1441 9974 1442 9978
rect 1446 9974 1447 9978
rect 1451 9974 1452 9978
rect 1456 9974 1457 9978
rect 1461 9974 1462 9978
rect 1466 9974 1467 9978
rect 1371 9973 1467 9974
rect 1371 9969 1372 9973
rect 1376 9969 1377 9973
rect 1371 9968 1377 9969
rect 1371 9964 1372 9968
rect 1376 9964 1377 9968
rect 1461 9969 1462 9973
rect 1466 9969 1467 9973
rect 1461 9968 1467 9969
rect 1371 9963 1377 9964
rect 1371 9959 1372 9963
rect 1376 9959 1377 9963
rect 1371 9958 1377 9959
rect 1371 9954 1372 9958
rect 1376 9954 1377 9958
rect 1371 9953 1377 9954
rect 1371 9949 1372 9953
rect 1376 9949 1377 9953
rect 1371 9948 1377 9949
rect 1371 9944 1372 9948
rect 1376 9944 1377 9948
rect 1371 9943 1377 9944
rect 1371 9939 1372 9943
rect 1376 9939 1377 9943
rect 1371 9938 1377 9939
rect 1371 9934 1372 9938
rect 1376 9934 1377 9938
rect 1371 9933 1377 9934
rect 1371 9929 1372 9933
rect 1376 9929 1377 9933
rect 1371 9928 1377 9929
rect 1371 9924 1372 9928
rect 1376 9924 1377 9928
rect 1371 9923 1377 9924
rect 1371 9919 1372 9923
rect 1376 9919 1377 9923
rect 1371 9918 1377 9919
rect 1371 9914 1372 9918
rect 1376 9914 1377 9918
rect 1371 9913 1377 9914
rect 1371 9909 1372 9913
rect 1376 9909 1377 9913
rect 1371 9908 1377 9909
rect 1371 9904 1372 9908
rect 1376 9904 1377 9908
rect 1371 9903 1377 9904
rect 1371 9899 1372 9903
rect 1376 9899 1377 9903
rect 1371 9898 1377 9899
rect 1371 9894 1372 9898
rect 1376 9894 1377 9898
rect 1371 9893 1377 9894
rect 1371 9889 1372 9893
rect 1376 9889 1377 9893
rect 1371 9888 1377 9889
rect 1371 9884 1372 9888
rect 1376 9884 1377 9888
rect 1371 9883 1377 9884
rect 1371 9879 1372 9883
rect 1376 9879 1377 9883
rect 1371 9878 1377 9879
rect 1371 9874 1372 9878
rect 1376 9874 1377 9878
rect 1371 9873 1377 9874
rect 1371 9869 1372 9873
rect 1376 9869 1377 9873
rect 1371 9868 1377 9869
rect 1371 9864 1372 9868
rect 1376 9864 1377 9868
rect 1371 9863 1377 9864
rect 1371 9859 1372 9863
rect 1376 9859 1377 9863
rect 1371 9858 1377 9859
rect 1371 9854 1372 9858
rect 1376 9854 1377 9858
rect 1371 9853 1377 9854
rect 1371 9849 1372 9853
rect 1376 9849 1377 9853
rect 1461 9964 1462 9968
rect 1466 9964 1467 9968
rect 1461 9963 1467 9964
rect 1461 9959 1462 9963
rect 1466 9959 1467 9963
rect 1461 9958 1467 9959
rect 1461 9954 1462 9958
rect 1466 9954 1467 9958
rect 1461 9953 1467 9954
rect 1461 9949 1462 9953
rect 1466 9949 1467 9953
rect 1461 9948 1467 9949
rect 1461 9944 1462 9948
rect 1466 9944 1467 9948
rect 1461 9943 1467 9944
rect 1461 9939 1462 9943
rect 1466 9939 1467 9943
rect 1461 9938 1467 9939
rect 1461 9934 1462 9938
rect 1466 9934 1467 9938
rect 1461 9933 1467 9934
rect 1461 9929 1462 9933
rect 1466 9929 1467 9933
rect 1461 9928 1467 9929
rect 1461 9924 1462 9928
rect 1466 9924 1467 9928
rect 1461 9923 1467 9924
rect 1461 9919 1462 9923
rect 1466 9919 1467 9923
rect 1461 9918 1467 9919
rect 1461 9914 1462 9918
rect 1466 9914 1467 9918
rect 1461 9913 1467 9914
rect 1461 9909 1462 9913
rect 1466 9909 1467 9913
rect 1461 9908 1467 9909
rect 1461 9904 1462 9908
rect 1466 9904 1467 9908
rect 1461 9903 1467 9904
rect 1461 9899 1462 9903
rect 1466 9899 1467 9903
rect 1461 9898 1467 9899
rect 1461 9894 1462 9898
rect 1466 9894 1467 9898
rect 1461 9893 1467 9894
rect 1461 9889 1462 9893
rect 1466 9889 1467 9893
rect 1461 9888 1467 9889
rect 1461 9884 1462 9888
rect 1466 9884 1467 9888
rect 1461 9883 1467 9884
rect 1461 9879 1462 9883
rect 1466 9879 1467 9883
rect 1461 9878 1467 9879
rect 1461 9874 1462 9878
rect 1466 9874 1467 9878
rect 1461 9873 1467 9874
rect 1461 9869 1462 9873
rect 1466 9869 1467 9873
rect 1461 9868 1467 9869
rect 1461 9864 1462 9868
rect 1466 9864 1467 9868
rect 1461 9863 1467 9864
rect 1461 9859 1462 9863
rect 1466 9859 1467 9863
rect 1461 9858 1467 9859
rect 1461 9854 1462 9858
rect 1466 9854 1467 9858
rect 1461 9853 1467 9854
rect 1371 9848 1377 9849
rect 1371 9844 1372 9848
rect 1376 9844 1377 9848
rect 1461 9849 1462 9853
rect 1466 9849 1467 9853
rect 1461 9848 1467 9849
rect 1461 9844 1462 9848
rect 1466 9844 1467 9848
rect 1371 9843 1467 9844
rect 1371 9839 1372 9843
rect 1376 9839 1377 9843
rect 1381 9839 1382 9843
rect 1386 9839 1387 9843
rect 1391 9839 1392 9843
rect 1396 9839 1397 9843
rect 1401 9839 1402 9843
rect 1406 9839 1407 9843
rect 1411 9839 1412 9843
rect 1416 9839 1417 9843
rect 1421 9839 1422 9843
rect 1426 9839 1427 9843
rect 1431 9839 1432 9843
rect 1436 9839 1437 9843
rect 1441 9839 1442 9843
rect 1446 9839 1447 9843
rect 1451 9839 1452 9843
rect 1456 9839 1457 9843
rect 1461 9839 1462 9843
rect 1466 9839 1467 9843
rect 1371 9838 1467 9839
rect 1543 9965 1615 9967
rect 1543 9961 1545 9965
rect 1549 9961 1552 9965
rect 1556 9961 1557 9965
rect 1561 9961 1562 9965
rect 1566 9961 1567 9965
rect 1571 9961 1572 9965
rect 1576 9961 1577 9965
rect 1581 9961 1582 9965
rect 1586 9961 1587 9965
rect 1591 9961 1592 9965
rect 1596 9961 1597 9965
rect 1601 9961 1602 9965
rect 1606 9961 1609 9965
rect 1613 9961 1615 9965
rect 1543 9959 1615 9961
rect 1543 9958 1551 9959
rect 1543 9954 1545 9958
rect 1549 9954 1551 9958
rect 1543 9953 1551 9954
rect 1607 9958 1615 9959
rect 1607 9954 1609 9958
rect 1613 9954 1615 9958
rect 1607 9953 1615 9954
rect 1543 9949 1545 9953
rect 1549 9949 1551 9953
rect 1543 9948 1551 9949
rect 1543 9944 1545 9948
rect 1549 9944 1551 9948
rect 1543 9943 1551 9944
rect 1543 9939 1545 9943
rect 1549 9939 1551 9943
rect 1543 9938 1551 9939
rect 1543 9934 1545 9938
rect 1549 9934 1551 9938
rect 1543 9933 1551 9934
rect 1543 9929 1545 9933
rect 1549 9929 1551 9933
rect 1543 9928 1551 9929
rect 1543 9924 1545 9928
rect 1549 9924 1551 9928
rect 1543 9923 1551 9924
rect 1543 9919 1545 9923
rect 1549 9919 1551 9923
rect 1543 9918 1551 9919
rect 1543 9914 1545 9918
rect 1549 9914 1551 9918
rect 1543 9913 1551 9914
rect 1543 9909 1545 9913
rect 1549 9909 1551 9913
rect 1543 9908 1551 9909
rect 1543 9904 1545 9908
rect 1549 9904 1551 9908
rect 1543 9903 1551 9904
rect 1543 9899 1545 9903
rect 1549 9899 1551 9903
rect 1543 9898 1551 9899
rect 1543 9894 1545 9898
rect 1549 9894 1551 9898
rect 1543 9893 1551 9894
rect 1543 9889 1545 9893
rect 1549 9889 1551 9893
rect 1543 9888 1551 9889
rect 1543 9884 1545 9888
rect 1549 9884 1551 9888
rect 1543 9883 1551 9884
rect 1543 9879 1545 9883
rect 1549 9879 1551 9883
rect 1543 9878 1551 9879
rect 1543 9874 1545 9878
rect 1549 9874 1551 9878
rect 1543 9873 1551 9874
rect 1543 9869 1545 9873
rect 1549 9869 1551 9873
rect 1543 9868 1551 9869
rect 1543 9864 1545 9868
rect 1549 9864 1551 9868
rect 1607 9949 1609 9953
rect 1613 9949 1615 9953
rect 1607 9948 1615 9949
rect 1607 9944 1609 9948
rect 1613 9944 1615 9948
rect 1607 9943 1615 9944
rect 1607 9939 1609 9943
rect 1613 9939 1615 9943
rect 1607 9938 1615 9939
rect 1607 9934 1609 9938
rect 1613 9934 1615 9938
rect 1607 9933 1615 9934
rect 1607 9929 1609 9933
rect 1613 9929 1615 9933
rect 1607 9928 1615 9929
rect 1607 9924 1609 9928
rect 1613 9924 1615 9928
rect 1607 9923 1615 9924
rect 1607 9919 1609 9923
rect 1613 9919 1615 9923
rect 1607 9918 1615 9919
rect 1607 9914 1609 9918
rect 1613 9914 1615 9918
rect 1607 9913 1615 9914
rect 1607 9909 1609 9913
rect 1613 9909 1615 9913
rect 1607 9908 1615 9909
rect 1607 9904 1609 9908
rect 1613 9904 1615 9908
rect 1607 9903 1615 9904
rect 1607 9899 1609 9903
rect 1613 9899 1615 9903
rect 1607 9898 1615 9899
rect 1607 9894 1609 9898
rect 1613 9894 1615 9898
rect 1607 9893 1615 9894
rect 1607 9889 1609 9893
rect 1613 9889 1615 9893
rect 1607 9888 1615 9889
rect 1607 9884 1609 9888
rect 1613 9884 1615 9888
rect 1607 9883 1615 9884
rect 1607 9879 1609 9883
rect 1613 9879 1615 9883
rect 1607 9878 1615 9879
rect 1607 9874 1609 9878
rect 1613 9874 1615 9878
rect 1607 9873 1615 9874
rect 1607 9869 1609 9873
rect 1613 9869 1615 9873
rect 1607 9868 1615 9869
rect 1607 9864 1609 9868
rect 1613 9864 1615 9868
rect 1543 9863 1551 9864
rect 1543 9859 1545 9863
rect 1549 9859 1551 9863
rect 1543 9858 1551 9859
rect 1607 9863 1615 9864
rect 1607 9859 1609 9863
rect 1613 9859 1615 9863
rect 1607 9858 1615 9859
rect 1543 9856 1615 9858
rect 1543 9852 1545 9856
rect 1549 9852 1552 9856
rect 1556 9852 1557 9856
rect 1561 9852 1562 9856
rect 1566 9852 1567 9856
rect 1571 9852 1572 9856
rect 1576 9852 1577 9856
rect 1581 9852 1582 9856
rect 1586 9852 1587 9856
rect 1591 9852 1592 9856
rect 1596 9852 1597 9856
rect 1601 9852 1602 9856
rect 1606 9852 1609 9856
rect 1613 9852 1615 9856
rect 1543 9850 1615 9852
rect 1680 9978 1776 9979
rect 1680 9974 1681 9978
rect 1685 9974 1686 9978
rect 1690 9974 1691 9978
rect 1695 9974 1696 9978
rect 1700 9974 1701 9978
rect 1705 9974 1706 9978
rect 1710 9974 1711 9978
rect 1715 9974 1716 9978
rect 1720 9974 1721 9978
rect 1725 9974 1726 9978
rect 1730 9974 1731 9978
rect 1735 9974 1736 9978
rect 1740 9974 1741 9978
rect 1745 9974 1746 9978
rect 1750 9974 1751 9978
rect 1755 9974 1756 9978
rect 1760 9974 1761 9978
rect 1765 9974 1766 9978
rect 1770 9974 1771 9978
rect 1775 9974 1776 9978
rect 1680 9973 1776 9974
rect 1680 9969 1681 9973
rect 1685 9969 1686 9973
rect 1680 9968 1686 9969
rect 1680 9964 1681 9968
rect 1685 9964 1686 9968
rect 1770 9969 1771 9973
rect 1775 9969 1776 9973
rect 1770 9968 1776 9969
rect 1680 9963 1686 9964
rect 1680 9959 1681 9963
rect 1685 9959 1686 9963
rect 1680 9958 1686 9959
rect 1680 9954 1681 9958
rect 1685 9954 1686 9958
rect 1680 9953 1686 9954
rect 1680 9949 1681 9953
rect 1685 9949 1686 9953
rect 1680 9948 1686 9949
rect 1680 9944 1681 9948
rect 1685 9944 1686 9948
rect 1680 9943 1686 9944
rect 1680 9939 1681 9943
rect 1685 9939 1686 9943
rect 1680 9938 1686 9939
rect 1680 9934 1681 9938
rect 1685 9934 1686 9938
rect 1680 9933 1686 9934
rect 1680 9929 1681 9933
rect 1685 9929 1686 9933
rect 1680 9928 1686 9929
rect 1680 9924 1681 9928
rect 1685 9924 1686 9928
rect 1680 9923 1686 9924
rect 1680 9919 1681 9923
rect 1685 9919 1686 9923
rect 1680 9918 1686 9919
rect 1680 9914 1681 9918
rect 1685 9914 1686 9918
rect 1680 9913 1686 9914
rect 1680 9909 1681 9913
rect 1685 9909 1686 9913
rect 1680 9908 1686 9909
rect 1680 9904 1681 9908
rect 1685 9904 1686 9908
rect 1680 9903 1686 9904
rect 1680 9899 1681 9903
rect 1685 9899 1686 9903
rect 1680 9898 1686 9899
rect 1680 9894 1681 9898
rect 1685 9894 1686 9898
rect 1680 9893 1686 9894
rect 1680 9889 1681 9893
rect 1685 9889 1686 9893
rect 1680 9888 1686 9889
rect 1680 9884 1681 9888
rect 1685 9884 1686 9888
rect 1680 9883 1686 9884
rect 1680 9879 1681 9883
rect 1685 9879 1686 9883
rect 1680 9878 1686 9879
rect 1680 9874 1681 9878
rect 1685 9874 1686 9878
rect 1680 9873 1686 9874
rect 1680 9869 1681 9873
rect 1685 9869 1686 9873
rect 1680 9868 1686 9869
rect 1680 9864 1681 9868
rect 1685 9864 1686 9868
rect 1680 9863 1686 9864
rect 1680 9859 1681 9863
rect 1685 9859 1686 9863
rect 1680 9858 1686 9859
rect 1680 9854 1681 9858
rect 1685 9854 1686 9858
rect 1680 9853 1686 9854
rect 1680 9849 1681 9853
rect 1685 9849 1686 9853
rect 1770 9964 1771 9968
rect 1775 9964 1776 9968
rect 1770 9963 1776 9964
rect 1770 9959 1771 9963
rect 1775 9959 1776 9963
rect 1770 9958 1776 9959
rect 1770 9954 1771 9958
rect 1775 9954 1776 9958
rect 1770 9953 1776 9954
rect 1770 9949 1771 9953
rect 1775 9949 1776 9953
rect 1770 9948 1776 9949
rect 1770 9944 1771 9948
rect 1775 9944 1776 9948
rect 1770 9943 1776 9944
rect 1770 9939 1771 9943
rect 1775 9939 1776 9943
rect 1770 9938 1776 9939
rect 1770 9934 1771 9938
rect 1775 9934 1776 9938
rect 1770 9933 1776 9934
rect 1770 9929 1771 9933
rect 1775 9929 1776 9933
rect 1770 9928 1776 9929
rect 1770 9924 1771 9928
rect 1775 9924 1776 9928
rect 1770 9923 1776 9924
rect 1770 9919 1771 9923
rect 1775 9919 1776 9923
rect 1770 9918 1776 9919
rect 1770 9914 1771 9918
rect 1775 9914 1776 9918
rect 1770 9913 1776 9914
rect 1770 9909 1771 9913
rect 1775 9909 1776 9913
rect 1770 9908 1776 9909
rect 1770 9904 1771 9908
rect 1775 9904 1776 9908
rect 1770 9903 1776 9904
rect 1770 9899 1771 9903
rect 1775 9899 1776 9903
rect 1770 9898 1776 9899
rect 1770 9894 1771 9898
rect 1775 9894 1776 9898
rect 1770 9893 1776 9894
rect 1770 9889 1771 9893
rect 1775 9889 1776 9893
rect 1770 9888 1776 9889
rect 1770 9884 1771 9888
rect 1775 9884 1776 9888
rect 1770 9883 1776 9884
rect 1770 9879 1771 9883
rect 1775 9879 1776 9883
rect 1770 9878 1776 9879
rect 1770 9874 1771 9878
rect 1775 9874 1776 9878
rect 1770 9873 1776 9874
rect 1770 9869 1771 9873
rect 1775 9869 1776 9873
rect 1770 9868 1776 9869
rect 1770 9864 1771 9868
rect 1775 9864 1776 9868
rect 1770 9863 1776 9864
rect 1770 9859 1771 9863
rect 1775 9859 1776 9863
rect 1770 9858 1776 9859
rect 1770 9854 1771 9858
rect 1775 9854 1776 9858
rect 1770 9853 1776 9854
rect 1680 9848 1686 9849
rect 1680 9844 1681 9848
rect 1685 9844 1686 9848
rect 1770 9849 1771 9853
rect 1775 9849 1776 9853
rect 1770 9848 1776 9849
rect 1770 9844 1771 9848
rect 1775 9844 1776 9848
rect 1680 9843 1776 9844
rect 1680 9839 1681 9843
rect 1685 9839 1686 9843
rect 1690 9839 1691 9843
rect 1695 9839 1696 9843
rect 1700 9839 1701 9843
rect 1705 9839 1706 9843
rect 1710 9839 1711 9843
rect 1715 9839 1716 9843
rect 1720 9839 1721 9843
rect 1725 9839 1726 9843
rect 1730 9839 1731 9843
rect 1735 9839 1736 9843
rect 1740 9839 1741 9843
rect 1745 9839 1746 9843
rect 1750 9839 1751 9843
rect 1755 9839 1756 9843
rect 1760 9839 1761 9843
rect 1765 9839 1766 9843
rect 1770 9839 1771 9843
rect 1775 9839 1776 9843
rect 1680 9838 1776 9839
rect 1852 9965 1924 9967
rect 1852 9961 1854 9965
rect 1858 9961 1861 9965
rect 1865 9961 1866 9965
rect 1870 9961 1871 9965
rect 1875 9961 1876 9965
rect 1880 9961 1881 9965
rect 1885 9961 1886 9965
rect 1890 9961 1891 9965
rect 1895 9961 1896 9965
rect 1900 9961 1901 9965
rect 1905 9961 1906 9965
rect 1910 9961 1911 9965
rect 1915 9961 1918 9965
rect 1922 9961 1924 9965
rect 1852 9959 1924 9961
rect 1852 9958 1860 9959
rect 1852 9954 1854 9958
rect 1858 9954 1860 9958
rect 1852 9953 1860 9954
rect 1916 9958 1924 9959
rect 1916 9954 1918 9958
rect 1922 9954 1924 9958
rect 1916 9953 1924 9954
rect 1852 9949 1854 9953
rect 1858 9949 1860 9953
rect 1852 9948 1860 9949
rect 1852 9944 1854 9948
rect 1858 9944 1860 9948
rect 1852 9943 1860 9944
rect 1852 9939 1854 9943
rect 1858 9939 1860 9943
rect 1852 9938 1860 9939
rect 1852 9934 1854 9938
rect 1858 9934 1860 9938
rect 1852 9933 1860 9934
rect 1852 9929 1854 9933
rect 1858 9929 1860 9933
rect 1852 9928 1860 9929
rect 1852 9924 1854 9928
rect 1858 9924 1860 9928
rect 1852 9923 1860 9924
rect 1852 9919 1854 9923
rect 1858 9919 1860 9923
rect 1852 9918 1860 9919
rect 1852 9914 1854 9918
rect 1858 9914 1860 9918
rect 1852 9913 1860 9914
rect 1852 9909 1854 9913
rect 1858 9909 1860 9913
rect 1852 9908 1860 9909
rect 1852 9904 1854 9908
rect 1858 9904 1860 9908
rect 1852 9903 1860 9904
rect 1852 9899 1854 9903
rect 1858 9899 1860 9903
rect 1852 9898 1860 9899
rect 1852 9894 1854 9898
rect 1858 9894 1860 9898
rect 1852 9893 1860 9894
rect 1852 9889 1854 9893
rect 1858 9889 1860 9893
rect 1852 9888 1860 9889
rect 1852 9884 1854 9888
rect 1858 9884 1860 9888
rect 1852 9883 1860 9884
rect 1852 9879 1854 9883
rect 1858 9879 1860 9883
rect 1852 9878 1860 9879
rect 1852 9874 1854 9878
rect 1858 9874 1860 9878
rect 1852 9873 1860 9874
rect 1852 9869 1854 9873
rect 1858 9869 1860 9873
rect 1852 9868 1860 9869
rect 1852 9864 1854 9868
rect 1858 9864 1860 9868
rect 1916 9949 1918 9953
rect 1922 9949 1924 9953
rect 1916 9948 1924 9949
rect 1916 9944 1918 9948
rect 1922 9944 1924 9948
rect 1916 9943 1924 9944
rect 1916 9939 1918 9943
rect 1922 9939 1924 9943
rect 1916 9938 1924 9939
rect 1916 9934 1918 9938
rect 1922 9934 1924 9938
rect 1916 9933 1924 9934
rect 1916 9929 1918 9933
rect 1922 9929 1924 9933
rect 1916 9928 1924 9929
rect 1916 9924 1918 9928
rect 1922 9924 1924 9928
rect 1916 9923 1924 9924
rect 1916 9919 1918 9923
rect 1922 9919 1924 9923
rect 1916 9918 1924 9919
rect 1916 9914 1918 9918
rect 1922 9914 1924 9918
rect 1916 9913 1924 9914
rect 1916 9909 1918 9913
rect 1922 9909 1924 9913
rect 1916 9908 1924 9909
rect 1916 9904 1918 9908
rect 1922 9904 1924 9908
rect 1916 9903 1924 9904
rect 1916 9899 1918 9903
rect 1922 9899 1924 9903
rect 1916 9898 1924 9899
rect 1916 9894 1918 9898
rect 1922 9894 1924 9898
rect 1916 9893 1924 9894
rect 1916 9889 1918 9893
rect 1922 9889 1924 9893
rect 1916 9888 1924 9889
rect 1916 9884 1918 9888
rect 1922 9884 1924 9888
rect 1916 9883 1924 9884
rect 1916 9879 1918 9883
rect 1922 9879 1924 9883
rect 1916 9878 1924 9879
rect 1916 9874 1918 9878
rect 1922 9874 1924 9878
rect 1916 9873 1924 9874
rect 1916 9869 1918 9873
rect 1922 9869 1924 9873
rect 1916 9868 1924 9869
rect 1916 9864 1918 9868
rect 1922 9864 1924 9868
rect 1852 9863 1860 9864
rect 1852 9859 1854 9863
rect 1858 9859 1860 9863
rect 1852 9858 1860 9859
rect 1916 9863 1924 9864
rect 1916 9859 1918 9863
rect 1922 9859 1924 9863
rect 1916 9858 1924 9859
rect 1852 9856 1924 9858
rect 1852 9852 1854 9856
rect 1858 9852 1861 9856
rect 1865 9852 1866 9856
rect 1870 9852 1871 9856
rect 1875 9852 1876 9856
rect 1880 9852 1881 9856
rect 1885 9852 1886 9856
rect 1890 9852 1891 9856
rect 1895 9852 1896 9856
rect 1900 9852 1901 9856
rect 1905 9852 1906 9856
rect 1910 9852 1911 9856
rect 1915 9852 1918 9856
rect 1922 9852 1924 9856
rect 1852 9850 1924 9852
rect 1989 9978 2085 9979
rect 1989 9974 1990 9978
rect 1994 9974 1995 9978
rect 1999 9974 2000 9978
rect 2004 9974 2005 9978
rect 2009 9974 2010 9978
rect 2014 9974 2015 9978
rect 2019 9974 2020 9978
rect 2024 9974 2025 9978
rect 2029 9974 2030 9978
rect 2034 9974 2035 9978
rect 2039 9974 2040 9978
rect 2044 9974 2045 9978
rect 2049 9974 2050 9978
rect 2054 9974 2055 9978
rect 2059 9974 2060 9978
rect 2064 9974 2065 9978
rect 2069 9974 2070 9978
rect 2074 9974 2075 9978
rect 2079 9974 2080 9978
rect 2084 9974 2085 9978
rect 1989 9973 2085 9974
rect 1989 9969 1990 9973
rect 1994 9969 1995 9973
rect 1989 9968 1995 9969
rect 1989 9964 1990 9968
rect 1994 9964 1995 9968
rect 2079 9969 2080 9973
rect 2084 9969 2085 9973
rect 2079 9968 2085 9969
rect 1989 9963 1995 9964
rect 1989 9959 1990 9963
rect 1994 9959 1995 9963
rect 1989 9958 1995 9959
rect 1989 9954 1990 9958
rect 1994 9954 1995 9958
rect 1989 9953 1995 9954
rect 1989 9949 1990 9953
rect 1994 9949 1995 9953
rect 1989 9948 1995 9949
rect 1989 9944 1990 9948
rect 1994 9944 1995 9948
rect 1989 9943 1995 9944
rect 1989 9939 1990 9943
rect 1994 9939 1995 9943
rect 1989 9938 1995 9939
rect 1989 9934 1990 9938
rect 1994 9934 1995 9938
rect 1989 9933 1995 9934
rect 1989 9929 1990 9933
rect 1994 9929 1995 9933
rect 1989 9928 1995 9929
rect 1989 9924 1990 9928
rect 1994 9924 1995 9928
rect 1989 9923 1995 9924
rect 1989 9919 1990 9923
rect 1994 9919 1995 9923
rect 1989 9918 1995 9919
rect 1989 9914 1990 9918
rect 1994 9914 1995 9918
rect 1989 9913 1995 9914
rect 1989 9909 1990 9913
rect 1994 9909 1995 9913
rect 1989 9908 1995 9909
rect 1989 9904 1990 9908
rect 1994 9904 1995 9908
rect 1989 9903 1995 9904
rect 1989 9899 1990 9903
rect 1994 9899 1995 9903
rect 1989 9898 1995 9899
rect 1989 9894 1990 9898
rect 1994 9894 1995 9898
rect 1989 9893 1995 9894
rect 1989 9889 1990 9893
rect 1994 9889 1995 9893
rect 1989 9888 1995 9889
rect 1989 9884 1990 9888
rect 1994 9884 1995 9888
rect 1989 9883 1995 9884
rect 1989 9879 1990 9883
rect 1994 9879 1995 9883
rect 1989 9878 1995 9879
rect 1989 9874 1990 9878
rect 1994 9874 1995 9878
rect 1989 9873 1995 9874
rect 1989 9869 1990 9873
rect 1994 9869 1995 9873
rect 1989 9868 1995 9869
rect 1989 9864 1990 9868
rect 1994 9864 1995 9868
rect 1989 9863 1995 9864
rect 1989 9859 1990 9863
rect 1994 9859 1995 9863
rect 1989 9858 1995 9859
rect 1989 9854 1990 9858
rect 1994 9854 1995 9858
rect 1989 9853 1995 9854
rect 1989 9849 1990 9853
rect 1994 9849 1995 9853
rect 2079 9964 2080 9968
rect 2084 9964 2085 9968
rect 2079 9963 2085 9964
rect 2079 9959 2080 9963
rect 2084 9959 2085 9963
rect 2079 9958 2085 9959
rect 2079 9954 2080 9958
rect 2084 9954 2085 9958
rect 2079 9953 2085 9954
rect 2079 9949 2080 9953
rect 2084 9949 2085 9953
rect 2079 9948 2085 9949
rect 2079 9944 2080 9948
rect 2084 9944 2085 9948
rect 2079 9943 2085 9944
rect 2079 9939 2080 9943
rect 2084 9939 2085 9943
rect 2079 9938 2085 9939
rect 2079 9934 2080 9938
rect 2084 9934 2085 9938
rect 2079 9933 2085 9934
rect 2079 9929 2080 9933
rect 2084 9929 2085 9933
rect 2079 9928 2085 9929
rect 2079 9924 2080 9928
rect 2084 9924 2085 9928
rect 2079 9923 2085 9924
rect 2079 9919 2080 9923
rect 2084 9919 2085 9923
rect 2079 9918 2085 9919
rect 2079 9914 2080 9918
rect 2084 9914 2085 9918
rect 2079 9913 2085 9914
rect 2079 9909 2080 9913
rect 2084 9909 2085 9913
rect 2079 9908 2085 9909
rect 2079 9904 2080 9908
rect 2084 9904 2085 9908
rect 2079 9903 2085 9904
rect 2079 9899 2080 9903
rect 2084 9899 2085 9903
rect 2079 9898 2085 9899
rect 2079 9894 2080 9898
rect 2084 9894 2085 9898
rect 2079 9893 2085 9894
rect 2079 9889 2080 9893
rect 2084 9889 2085 9893
rect 2079 9888 2085 9889
rect 2079 9884 2080 9888
rect 2084 9884 2085 9888
rect 2079 9883 2085 9884
rect 2079 9879 2080 9883
rect 2084 9879 2085 9883
rect 2079 9878 2085 9879
rect 2079 9874 2080 9878
rect 2084 9874 2085 9878
rect 2079 9873 2085 9874
rect 2079 9869 2080 9873
rect 2084 9869 2085 9873
rect 2079 9868 2085 9869
rect 2079 9864 2080 9868
rect 2084 9864 2085 9868
rect 2079 9863 2085 9864
rect 2079 9859 2080 9863
rect 2084 9859 2085 9863
rect 2079 9858 2085 9859
rect 2079 9854 2080 9858
rect 2084 9854 2085 9858
rect 2079 9853 2085 9854
rect 1989 9848 1995 9849
rect 1989 9844 1990 9848
rect 1994 9844 1995 9848
rect 2079 9849 2080 9853
rect 2084 9849 2085 9853
rect 2079 9848 2085 9849
rect 2079 9844 2080 9848
rect 2084 9844 2085 9848
rect 1989 9843 2085 9844
rect 1989 9839 1990 9843
rect 1994 9839 1995 9843
rect 1999 9839 2000 9843
rect 2004 9839 2005 9843
rect 2009 9839 2010 9843
rect 2014 9839 2015 9843
rect 2019 9839 2020 9843
rect 2024 9839 2025 9843
rect 2029 9839 2030 9843
rect 2034 9839 2035 9843
rect 2039 9839 2040 9843
rect 2044 9839 2045 9843
rect 2049 9839 2050 9843
rect 2054 9839 2055 9843
rect 2059 9839 2060 9843
rect 2064 9839 2065 9843
rect 2069 9839 2070 9843
rect 2074 9839 2075 9843
rect 2079 9839 2080 9843
rect 2084 9839 2085 9843
rect 1989 9838 2085 9839
rect 2161 9965 2233 9967
rect 2161 9961 2163 9965
rect 2167 9961 2170 9965
rect 2174 9961 2175 9965
rect 2179 9961 2180 9965
rect 2184 9961 2185 9965
rect 2189 9961 2190 9965
rect 2194 9961 2195 9965
rect 2199 9961 2200 9965
rect 2204 9961 2205 9965
rect 2209 9961 2210 9965
rect 2214 9961 2215 9965
rect 2219 9961 2220 9965
rect 2224 9961 2227 9965
rect 2231 9961 2233 9965
rect 2161 9959 2233 9961
rect 2161 9958 2169 9959
rect 2161 9954 2163 9958
rect 2167 9954 2169 9958
rect 2161 9953 2169 9954
rect 2225 9958 2233 9959
rect 2225 9954 2227 9958
rect 2231 9954 2233 9958
rect 2225 9953 2233 9954
rect 2161 9949 2163 9953
rect 2167 9949 2169 9953
rect 2161 9948 2169 9949
rect 2161 9944 2163 9948
rect 2167 9944 2169 9948
rect 2161 9943 2169 9944
rect 2161 9939 2163 9943
rect 2167 9939 2169 9943
rect 2161 9938 2169 9939
rect 2161 9934 2163 9938
rect 2167 9934 2169 9938
rect 2161 9933 2169 9934
rect 2161 9929 2163 9933
rect 2167 9929 2169 9933
rect 2161 9928 2169 9929
rect 2161 9924 2163 9928
rect 2167 9924 2169 9928
rect 2161 9923 2169 9924
rect 2161 9919 2163 9923
rect 2167 9919 2169 9923
rect 2161 9918 2169 9919
rect 2161 9914 2163 9918
rect 2167 9914 2169 9918
rect 2161 9913 2169 9914
rect 2161 9909 2163 9913
rect 2167 9909 2169 9913
rect 2161 9908 2169 9909
rect 2161 9904 2163 9908
rect 2167 9904 2169 9908
rect 2161 9903 2169 9904
rect 2161 9899 2163 9903
rect 2167 9899 2169 9903
rect 2161 9898 2169 9899
rect 2161 9894 2163 9898
rect 2167 9894 2169 9898
rect 2161 9893 2169 9894
rect 2161 9889 2163 9893
rect 2167 9889 2169 9893
rect 2161 9888 2169 9889
rect 2161 9884 2163 9888
rect 2167 9884 2169 9888
rect 2161 9883 2169 9884
rect 2161 9879 2163 9883
rect 2167 9879 2169 9883
rect 2161 9878 2169 9879
rect 2161 9874 2163 9878
rect 2167 9874 2169 9878
rect 2161 9873 2169 9874
rect 2161 9869 2163 9873
rect 2167 9869 2169 9873
rect 2161 9868 2169 9869
rect 2161 9864 2163 9868
rect 2167 9864 2169 9868
rect 2225 9949 2227 9953
rect 2231 9949 2233 9953
rect 2225 9948 2233 9949
rect 2225 9944 2227 9948
rect 2231 9944 2233 9948
rect 2225 9943 2233 9944
rect 2225 9939 2227 9943
rect 2231 9939 2233 9943
rect 2225 9938 2233 9939
rect 2225 9934 2227 9938
rect 2231 9934 2233 9938
rect 2225 9933 2233 9934
rect 2225 9929 2227 9933
rect 2231 9929 2233 9933
rect 2225 9928 2233 9929
rect 2225 9924 2227 9928
rect 2231 9924 2233 9928
rect 2225 9923 2233 9924
rect 2225 9919 2227 9923
rect 2231 9919 2233 9923
rect 2225 9918 2233 9919
rect 2225 9914 2227 9918
rect 2231 9914 2233 9918
rect 2225 9913 2233 9914
rect 2225 9909 2227 9913
rect 2231 9909 2233 9913
rect 2225 9908 2233 9909
rect 2225 9904 2227 9908
rect 2231 9904 2233 9908
rect 2225 9903 2233 9904
rect 2225 9899 2227 9903
rect 2231 9899 2233 9903
rect 2225 9898 2233 9899
rect 2225 9894 2227 9898
rect 2231 9894 2233 9898
rect 2225 9893 2233 9894
rect 2225 9889 2227 9893
rect 2231 9889 2233 9893
rect 2225 9888 2233 9889
rect 2225 9884 2227 9888
rect 2231 9884 2233 9888
rect 2225 9883 2233 9884
rect 2225 9879 2227 9883
rect 2231 9879 2233 9883
rect 2225 9878 2233 9879
rect 2225 9874 2227 9878
rect 2231 9874 2233 9878
rect 2225 9873 2233 9874
rect 2225 9869 2227 9873
rect 2231 9869 2233 9873
rect 2225 9868 2233 9869
rect 2225 9864 2227 9868
rect 2231 9864 2233 9868
rect 2161 9863 2169 9864
rect 2161 9859 2163 9863
rect 2167 9859 2169 9863
rect 2161 9858 2169 9859
rect 2225 9863 2233 9864
rect 2225 9859 2227 9863
rect 2231 9859 2233 9863
rect 2225 9858 2233 9859
rect 2161 9856 2233 9858
rect 2161 9852 2163 9856
rect 2167 9852 2170 9856
rect 2174 9852 2175 9856
rect 2179 9852 2180 9856
rect 2184 9852 2185 9856
rect 2189 9852 2190 9856
rect 2194 9852 2195 9856
rect 2199 9852 2200 9856
rect 2204 9852 2205 9856
rect 2209 9852 2210 9856
rect 2214 9852 2215 9856
rect 2219 9852 2220 9856
rect 2224 9852 2227 9856
rect 2231 9852 2233 9856
rect 2161 9850 2233 9852
rect 2298 9978 2394 9979
rect 2298 9974 2299 9978
rect 2303 9974 2304 9978
rect 2308 9974 2309 9978
rect 2313 9974 2314 9978
rect 2318 9974 2319 9978
rect 2323 9974 2324 9978
rect 2328 9974 2329 9978
rect 2333 9974 2334 9978
rect 2338 9974 2339 9978
rect 2343 9974 2344 9978
rect 2348 9974 2349 9978
rect 2353 9974 2354 9978
rect 2358 9974 2359 9978
rect 2363 9974 2364 9978
rect 2368 9974 2369 9978
rect 2373 9974 2374 9978
rect 2378 9974 2379 9978
rect 2383 9974 2384 9978
rect 2388 9974 2389 9978
rect 2393 9974 2394 9978
rect 2298 9973 2394 9974
rect 2298 9969 2299 9973
rect 2303 9969 2304 9973
rect 2298 9968 2304 9969
rect 2298 9964 2299 9968
rect 2303 9964 2304 9968
rect 2388 9969 2389 9973
rect 2393 9969 2394 9973
rect 2388 9968 2394 9969
rect 2298 9963 2304 9964
rect 2298 9959 2299 9963
rect 2303 9959 2304 9963
rect 2298 9958 2304 9959
rect 2298 9954 2299 9958
rect 2303 9954 2304 9958
rect 2298 9953 2304 9954
rect 2298 9949 2299 9953
rect 2303 9949 2304 9953
rect 2298 9948 2304 9949
rect 2298 9944 2299 9948
rect 2303 9944 2304 9948
rect 2298 9943 2304 9944
rect 2298 9939 2299 9943
rect 2303 9939 2304 9943
rect 2298 9938 2304 9939
rect 2298 9934 2299 9938
rect 2303 9934 2304 9938
rect 2298 9933 2304 9934
rect 2298 9929 2299 9933
rect 2303 9929 2304 9933
rect 2298 9928 2304 9929
rect 2298 9924 2299 9928
rect 2303 9924 2304 9928
rect 2298 9923 2304 9924
rect 2298 9919 2299 9923
rect 2303 9919 2304 9923
rect 2298 9918 2304 9919
rect 2298 9914 2299 9918
rect 2303 9914 2304 9918
rect 2298 9913 2304 9914
rect 2298 9909 2299 9913
rect 2303 9909 2304 9913
rect 2298 9908 2304 9909
rect 2298 9904 2299 9908
rect 2303 9904 2304 9908
rect 2298 9903 2304 9904
rect 2298 9899 2299 9903
rect 2303 9899 2304 9903
rect 2298 9898 2304 9899
rect 2298 9894 2299 9898
rect 2303 9894 2304 9898
rect 2298 9893 2304 9894
rect 2298 9889 2299 9893
rect 2303 9889 2304 9893
rect 2298 9888 2304 9889
rect 2298 9884 2299 9888
rect 2303 9884 2304 9888
rect 2298 9883 2304 9884
rect 2298 9879 2299 9883
rect 2303 9879 2304 9883
rect 2298 9878 2304 9879
rect 2298 9874 2299 9878
rect 2303 9874 2304 9878
rect 2298 9873 2304 9874
rect 2298 9869 2299 9873
rect 2303 9869 2304 9873
rect 2298 9868 2304 9869
rect 2298 9864 2299 9868
rect 2303 9864 2304 9868
rect 2298 9863 2304 9864
rect 2298 9859 2299 9863
rect 2303 9859 2304 9863
rect 2298 9858 2304 9859
rect 2298 9854 2299 9858
rect 2303 9854 2304 9858
rect 2298 9853 2304 9854
rect 2298 9849 2299 9853
rect 2303 9849 2304 9853
rect 2388 9964 2389 9968
rect 2393 9964 2394 9968
rect 2388 9963 2394 9964
rect 2388 9959 2389 9963
rect 2393 9959 2394 9963
rect 2388 9958 2394 9959
rect 2388 9954 2389 9958
rect 2393 9954 2394 9958
rect 2388 9953 2394 9954
rect 2388 9949 2389 9953
rect 2393 9949 2394 9953
rect 2388 9948 2394 9949
rect 2388 9944 2389 9948
rect 2393 9944 2394 9948
rect 2388 9943 2394 9944
rect 2388 9939 2389 9943
rect 2393 9939 2394 9943
rect 2388 9938 2394 9939
rect 2388 9934 2389 9938
rect 2393 9934 2394 9938
rect 2388 9933 2394 9934
rect 2388 9929 2389 9933
rect 2393 9929 2394 9933
rect 2388 9928 2394 9929
rect 2388 9924 2389 9928
rect 2393 9924 2394 9928
rect 2388 9923 2394 9924
rect 2388 9919 2389 9923
rect 2393 9919 2394 9923
rect 2388 9918 2394 9919
rect 2388 9914 2389 9918
rect 2393 9914 2394 9918
rect 2388 9913 2394 9914
rect 2388 9909 2389 9913
rect 2393 9909 2394 9913
rect 2388 9908 2394 9909
rect 2388 9904 2389 9908
rect 2393 9904 2394 9908
rect 2388 9903 2394 9904
rect 2388 9899 2389 9903
rect 2393 9899 2394 9903
rect 2388 9898 2394 9899
rect 2388 9894 2389 9898
rect 2393 9894 2394 9898
rect 2388 9893 2394 9894
rect 2388 9889 2389 9893
rect 2393 9889 2394 9893
rect 2388 9888 2394 9889
rect 2388 9884 2389 9888
rect 2393 9884 2394 9888
rect 2388 9883 2394 9884
rect 2388 9879 2389 9883
rect 2393 9879 2394 9883
rect 2388 9878 2394 9879
rect 2388 9874 2389 9878
rect 2393 9874 2394 9878
rect 2388 9873 2394 9874
rect 2388 9869 2389 9873
rect 2393 9869 2394 9873
rect 2388 9868 2394 9869
rect 2388 9864 2389 9868
rect 2393 9864 2394 9868
rect 2388 9863 2394 9864
rect 2388 9859 2389 9863
rect 2393 9859 2394 9863
rect 2388 9858 2394 9859
rect 2388 9854 2389 9858
rect 2393 9854 2394 9858
rect 2388 9853 2394 9854
rect 2298 9848 2304 9849
rect 2298 9844 2299 9848
rect 2303 9844 2304 9848
rect 2388 9849 2389 9853
rect 2393 9849 2394 9853
rect 2388 9848 2394 9849
rect 2388 9844 2389 9848
rect 2393 9844 2394 9848
rect 2298 9843 2394 9844
rect 2298 9839 2299 9843
rect 2303 9839 2304 9843
rect 2308 9839 2309 9843
rect 2313 9839 2314 9843
rect 2318 9839 2319 9843
rect 2323 9839 2324 9843
rect 2328 9839 2329 9843
rect 2333 9839 2334 9843
rect 2338 9839 2339 9843
rect 2343 9839 2344 9843
rect 2348 9839 2349 9843
rect 2353 9839 2354 9843
rect 2358 9839 2359 9843
rect 2363 9839 2364 9843
rect 2368 9839 2369 9843
rect 2373 9839 2374 9843
rect 2378 9839 2379 9843
rect 2383 9839 2384 9843
rect 2388 9839 2389 9843
rect 2393 9839 2394 9843
rect 2298 9838 2394 9839
rect 2470 9965 2542 9967
rect 2470 9961 2472 9965
rect 2476 9961 2479 9965
rect 2483 9961 2484 9965
rect 2488 9961 2489 9965
rect 2493 9961 2494 9965
rect 2498 9961 2499 9965
rect 2503 9961 2504 9965
rect 2508 9961 2509 9965
rect 2513 9961 2514 9965
rect 2518 9961 2519 9965
rect 2523 9961 2524 9965
rect 2528 9961 2529 9965
rect 2533 9961 2536 9965
rect 2540 9961 2542 9965
rect 2470 9959 2542 9961
rect 2470 9958 2478 9959
rect 2470 9954 2472 9958
rect 2476 9954 2478 9958
rect 2470 9953 2478 9954
rect 2534 9958 2542 9959
rect 2534 9954 2536 9958
rect 2540 9954 2542 9958
rect 2534 9953 2542 9954
rect 2470 9949 2472 9953
rect 2476 9949 2478 9953
rect 2470 9948 2478 9949
rect 2470 9944 2472 9948
rect 2476 9944 2478 9948
rect 2470 9943 2478 9944
rect 2470 9939 2472 9943
rect 2476 9939 2478 9943
rect 2470 9938 2478 9939
rect 2470 9934 2472 9938
rect 2476 9934 2478 9938
rect 2470 9933 2478 9934
rect 2470 9929 2472 9933
rect 2476 9929 2478 9933
rect 2470 9928 2478 9929
rect 2470 9924 2472 9928
rect 2476 9924 2478 9928
rect 2470 9923 2478 9924
rect 2470 9919 2472 9923
rect 2476 9919 2478 9923
rect 2470 9918 2478 9919
rect 2470 9914 2472 9918
rect 2476 9914 2478 9918
rect 2470 9913 2478 9914
rect 2470 9909 2472 9913
rect 2476 9909 2478 9913
rect 2470 9908 2478 9909
rect 2470 9904 2472 9908
rect 2476 9904 2478 9908
rect 2470 9903 2478 9904
rect 2470 9899 2472 9903
rect 2476 9899 2478 9903
rect 2470 9898 2478 9899
rect 2470 9894 2472 9898
rect 2476 9894 2478 9898
rect 2470 9893 2478 9894
rect 2470 9889 2472 9893
rect 2476 9889 2478 9893
rect 2470 9888 2478 9889
rect 2470 9884 2472 9888
rect 2476 9884 2478 9888
rect 2470 9883 2478 9884
rect 2470 9879 2472 9883
rect 2476 9879 2478 9883
rect 2470 9878 2478 9879
rect 2470 9874 2472 9878
rect 2476 9874 2478 9878
rect 2470 9873 2478 9874
rect 2470 9869 2472 9873
rect 2476 9869 2478 9873
rect 2470 9868 2478 9869
rect 2470 9864 2472 9868
rect 2476 9864 2478 9868
rect 2534 9949 2536 9953
rect 2540 9949 2542 9953
rect 2534 9948 2542 9949
rect 2534 9944 2536 9948
rect 2540 9944 2542 9948
rect 2534 9943 2542 9944
rect 2534 9939 2536 9943
rect 2540 9939 2542 9943
rect 2534 9938 2542 9939
rect 2534 9934 2536 9938
rect 2540 9934 2542 9938
rect 2534 9933 2542 9934
rect 2534 9929 2536 9933
rect 2540 9929 2542 9933
rect 2534 9928 2542 9929
rect 2534 9924 2536 9928
rect 2540 9924 2542 9928
rect 2534 9923 2542 9924
rect 2534 9919 2536 9923
rect 2540 9919 2542 9923
rect 2534 9918 2542 9919
rect 2534 9914 2536 9918
rect 2540 9914 2542 9918
rect 2534 9913 2542 9914
rect 2534 9909 2536 9913
rect 2540 9909 2542 9913
rect 2534 9908 2542 9909
rect 2534 9904 2536 9908
rect 2540 9904 2542 9908
rect 2534 9903 2542 9904
rect 2534 9899 2536 9903
rect 2540 9899 2542 9903
rect 2534 9898 2542 9899
rect 2534 9894 2536 9898
rect 2540 9894 2542 9898
rect 2534 9893 2542 9894
rect 2534 9889 2536 9893
rect 2540 9889 2542 9893
rect 2534 9888 2542 9889
rect 2534 9884 2536 9888
rect 2540 9884 2542 9888
rect 2534 9883 2542 9884
rect 2534 9879 2536 9883
rect 2540 9879 2542 9883
rect 2534 9878 2542 9879
rect 2534 9874 2536 9878
rect 2540 9874 2542 9878
rect 2534 9873 2542 9874
rect 2534 9869 2536 9873
rect 2540 9869 2542 9873
rect 2534 9868 2542 9869
rect 2534 9864 2536 9868
rect 2540 9864 2542 9868
rect 2470 9863 2478 9864
rect 2470 9859 2472 9863
rect 2476 9859 2478 9863
rect 2470 9858 2478 9859
rect 2534 9863 2542 9864
rect 2534 9859 2536 9863
rect 2540 9859 2542 9863
rect 2534 9858 2542 9859
rect 2470 9856 2542 9858
rect 2470 9852 2472 9856
rect 2476 9852 2479 9856
rect 2483 9852 2484 9856
rect 2488 9852 2489 9856
rect 2493 9852 2494 9856
rect 2498 9852 2499 9856
rect 2503 9852 2504 9856
rect 2508 9852 2509 9856
rect 2513 9852 2514 9856
rect 2518 9852 2519 9856
rect 2523 9852 2524 9856
rect 2528 9852 2529 9856
rect 2533 9852 2536 9856
rect 2540 9852 2542 9856
rect 2470 9850 2542 9852
rect 2607 9978 2703 9979
rect 2607 9974 2608 9978
rect 2612 9974 2613 9978
rect 2617 9974 2618 9978
rect 2622 9974 2623 9978
rect 2627 9974 2628 9978
rect 2632 9974 2633 9978
rect 2637 9974 2638 9978
rect 2642 9974 2643 9978
rect 2647 9974 2648 9978
rect 2652 9974 2653 9978
rect 2657 9974 2658 9978
rect 2662 9974 2663 9978
rect 2667 9974 2668 9978
rect 2672 9974 2673 9978
rect 2677 9974 2678 9978
rect 2682 9974 2683 9978
rect 2687 9974 2688 9978
rect 2692 9974 2693 9978
rect 2697 9974 2698 9978
rect 2702 9974 2703 9978
rect 2607 9973 2703 9974
rect 2607 9969 2608 9973
rect 2612 9969 2613 9973
rect 2607 9968 2613 9969
rect 2607 9964 2608 9968
rect 2612 9964 2613 9968
rect 2697 9969 2698 9973
rect 2702 9969 2703 9973
rect 2697 9968 2703 9969
rect 2607 9963 2613 9964
rect 2607 9959 2608 9963
rect 2612 9959 2613 9963
rect 2607 9958 2613 9959
rect 2607 9954 2608 9958
rect 2612 9954 2613 9958
rect 2607 9953 2613 9954
rect 2607 9949 2608 9953
rect 2612 9949 2613 9953
rect 2607 9948 2613 9949
rect 2607 9944 2608 9948
rect 2612 9944 2613 9948
rect 2607 9943 2613 9944
rect 2607 9939 2608 9943
rect 2612 9939 2613 9943
rect 2607 9938 2613 9939
rect 2607 9934 2608 9938
rect 2612 9934 2613 9938
rect 2607 9933 2613 9934
rect 2607 9929 2608 9933
rect 2612 9929 2613 9933
rect 2607 9928 2613 9929
rect 2607 9924 2608 9928
rect 2612 9924 2613 9928
rect 2607 9923 2613 9924
rect 2607 9919 2608 9923
rect 2612 9919 2613 9923
rect 2607 9918 2613 9919
rect 2607 9914 2608 9918
rect 2612 9914 2613 9918
rect 2607 9913 2613 9914
rect 2607 9909 2608 9913
rect 2612 9909 2613 9913
rect 2607 9908 2613 9909
rect 2607 9904 2608 9908
rect 2612 9904 2613 9908
rect 2607 9903 2613 9904
rect 2607 9899 2608 9903
rect 2612 9899 2613 9903
rect 2607 9898 2613 9899
rect 2607 9894 2608 9898
rect 2612 9894 2613 9898
rect 2607 9893 2613 9894
rect 2607 9889 2608 9893
rect 2612 9889 2613 9893
rect 2607 9888 2613 9889
rect 2607 9884 2608 9888
rect 2612 9884 2613 9888
rect 2607 9883 2613 9884
rect 2607 9879 2608 9883
rect 2612 9879 2613 9883
rect 2607 9878 2613 9879
rect 2607 9874 2608 9878
rect 2612 9874 2613 9878
rect 2607 9873 2613 9874
rect 2607 9869 2608 9873
rect 2612 9869 2613 9873
rect 2607 9868 2613 9869
rect 2607 9864 2608 9868
rect 2612 9864 2613 9868
rect 2607 9863 2613 9864
rect 2607 9859 2608 9863
rect 2612 9859 2613 9863
rect 2607 9858 2613 9859
rect 2607 9854 2608 9858
rect 2612 9854 2613 9858
rect 2607 9853 2613 9854
rect 2607 9849 2608 9853
rect 2612 9849 2613 9853
rect 2697 9964 2698 9968
rect 2702 9964 2703 9968
rect 2697 9963 2703 9964
rect 2697 9959 2698 9963
rect 2702 9959 2703 9963
rect 2697 9958 2703 9959
rect 2697 9954 2698 9958
rect 2702 9954 2703 9958
rect 2697 9953 2703 9954
rect 2697 9949 2698 9953
rect 2702 9949 2703 9953
rect 2697 9948 2703 9949
rect 2697 9944 2698 9948
rect 2702 9944 2703 9948
rect 2697 9943 2703 9944
rect 2697 9939 2698 9943
rect 2702 9939 2703 9943
rect 2697 9938 2703 9939
rect 2697 9934 2698 9938
rect 2702 9934 2703 9938
rect 2697 9933 2703 9934
rect 2697 9929 2698 9933
rect 2702 9929 2703 9933
rect 2697 9928 2703 9929
rect 2697 9924 2698 9928
rect 2702 9924 2703 9928
rect 2697 9923 2703 9924
rect 2697 9919 2698 9923
rect 2702 9919 2703 9923
rect 2697 9918 2703 9919
rect 2697 9914 2698 9918
rect 2702 9914 2703 9918
rect 2697 9913 2703 9914
rect 2697 9909 2698 9913
rect 2702 9909 2703 9913
rect 2697 9908 2703 9909
rect 2697 9904 2698 9908
rect 2702 9904 2703 9908
rect 2697 9903 2703 9904
rect 2697 9899 2698 9903
rect 2702 9899 2703 9903
rect 2697 9898 2703 9899
rect 2697 9894 2698 9898
rect 2702 9894 2703 9898
rect 2697 9893 2703 9894
rect 2697 9889 2698 9893
rect 2702 9889 2703 9893
rect 2697 9888 2703 9889
rect 2697 9884 2698 9888
rect 2702 9884 2703 9888
rect 2697 9883 2703 9884
rect 2697 9879 2698 9883
rect 2702 9879 2703 9883
rect 2697 9878 2703 9879
rect 2697 9874 2698 9878
rect 2702 9874 2703 9878
rect 2697 9873 2703 9874
rect 2697 9869 2698 9873
rect 2702 9869 2703 9873
rect 2697 9868 2703 9869
rect 2697 9864 2698 9868
rect 2702 9864 2703 9868
rect 2697 9863 2703 9864
rect 2697 9859 2698 9863
rect 2702 9859 2703 9863
rect 2697 9858 2703 9859
rect 2697 9854 2698 9858
rect 2702 9854 2703 9858
rect 2697 9853 2703 9854
rect 2607 9848 2613 9849
rect 2607 9844 2608 9848
rect 2612 9844 2613 9848
rect 2697 9849 2698 9853
rect 2702 9849 2703 9853
rect 2697 9848 2703 9849
rect 2697 9844 2698 9848
rect 2702 9844 2703 9848
rect 2607 9843 2703 9844
rect 2607 9839 2608 9843
rect 2612 9839 2613 9843
rect 2617 9839 2618 9843
rect 2622 9839 2623 9843
rect 2627 9839 2628 9843
rect 2632 9839 2633 9843
rect 2637 9839 2638 9843
rect 2642 9839 2643 9843
rect 2647 9839 2648 9843
rect 2652 9839 2653 9843
rect 2657 9839 2658 9843
rect 2662 9839 2663 9843
rect 2667 9839 2668 9843
rect 2672 9839 2673 9843
rect 2677 9839 2678 9843
rect 2682 9839 2683 9843
rect 2687 9839 2688 9843
rect 2692 9839 2693 9843
rect 2697 9839 2698 9843
rect 2702 9839 2703 9843
rect 2607 9838 2703 9839
rect 2779 9965 2851 9967
rect 2779 9961 2781 9965
rect 2785 9961 2788 9965
rect 2792 9961 2793 9965
rect 2797 9961 2798 9965
rect 2802 9961 2803 9965
rect 2807 9961 2808 9965
rect 2812 9961 2813 9965
rect 2817 9961 2818 9965
rect 2822 9961 2823 9965
rect 2827 9961 2828 9965
rect 2832 9961 2833 9965
rect 2837 9961 2838 9965
rect 2842 9961 2845 9965
rect 2849 9961 2851 9965
rect 2779 9959 2851 9961
rect 2779 9958 2787 9959
rect 2779 9954 2781 9958
rect 2785 9954 2787 9958
rect 2779 9953 2787 9954
rect 2843 9958 2851 9959
rect 2843 9954 2845 9958
rect 2849 9954 2851 9958
rect 2843 9953 2851 9954
rect 2779 9949 2781 9953
rect 2785 9949 2787 9953
rect 2779 9948 2787 9949
rect 2779 9944 2781 9948
rect 2785 9944 2787 9948
rect 2779 9943 2787 9944
rect 2779 9939 2781 9943
rect 2785 9939 2787 9943
rect 2779 9938 2787 9939
rect 2779 9934 2781 9938
rect 2785 9934 2787 9938
rect 2779 9933 2787 9934
rect 2779 9929 2781 9933
rect 2785 9929 2787 9933
rect 2779 9928 2787 9929
rect 2779 9924 2781 9928
rect 2785 9924 2787 9928
rect 2779 9923 2787 9924
rect 2779 9919 2781 9923
rect 2785 9919 2787 9923
rect 2779 9918 2787 9919
rect 2779 9914 2781 9918
rect 2785 9914 2787 9918
rect 2779 9913 2787 9914
rect 2779 9909 2781 9913
rect 2785 9909 2787 9913
rect 2779 9908 2787 9909
rect 2779 9904 2781 9908
rect 2785 9904 2787 9908
rect 2779 9903 2787 9904
rect 2779 9899 2781 9903
rect 2785 9899 2787 9903
rect 2779 9898 2787 9899
rect 2779 9894 2781 9898
rect 2785 9894 2787 9898
rect 2779 9893 2787 9894
rect 2779 9889 2781 9893
rect 2785 9889 2787 9893
rect 2779 9888 2787 9889
rect 2779 9884 2781 9888
rect 2785 9884 2787 9888
rect 2779 9883 2787 9884
rect 2779 9879 2781 9883
rect 2785 9879 2787 9883
rect 2779 9878 2787 9879
rect 2779 9874 2781 9878
rect 2785 9874 2787 9878
rect 2779 9873 2787 9874
rect 2779 9869 2781 9873
rect 2785 9869 2787 9873
rect 2779 9868 2787 9869
rect 2779 9864 2781 9868
rect 2785 9864 2787 9868
rect 2843 9949 2845 9953
rect 2849 9949 2851 9953
rect 2843 9948 2851 9949
rect 2843 9944 2845 9948
rect 2849 9944 2851 9948
rect 2843 9943 2851 9944
rect 2843 9939 2845 9943
rect 2849 9939 2851 9943
rect 2843 9938 2851 9939
rect 2843 9934 2845 9938
rect 2849 9934 2851 9938
rect 2843 9933 2851 9934
rect 2843 9929 2845 9933
rect 2849 9929 2851 9933
rect 2843 9928 2851 9929
rect 2843 9924 2845 9928
rect 2849 9924 2851 9928
rect 2843 9923 2851 9924
rect 2843 9919 2845 9923
rect 2849 9919 2851 9923
rect 2843 9918 2851 9919
rect 2843 9914 2845 9918
rect 2849 9914 2851 9918
rect 2843 9913 2851 9914
rect 2843 9909 2845 9913
rect 2849 9909 2851 9913
rect 2843 9908 2851 9909
rect 2843 9904 2845 9908
rect 2849 9904 2851 9908
rect 2843 9903 2851 9904
rect 2843 9899 2845 9903
rect 2849 9899 2851 9903
rect 2843 9898 2851 9899
rect 2843 9894 2845 9898
rect 2849 9894 2851 9898
rect 2843 9893 2851 9894
rect 2843 9889 2845 9893
rect 2849 9889 2851 9893
rect 2843 9888 2851 9889
rect 2843 9884 2845 9888
rect 2849 9884 2851 9888
rect 2843 9883 2851 9884
rect 2843 9879 2845 9883
rect 2849 9879 2851 9883
rect 2843 9878 2851 9879
rect 2843 9874 2845 9878
rect 2849 9874 2851 9878
rect 2843 9873 2851 9874
rect 2843 9869 2845 9873
rect 2849 9869 2851 9873
rect 2843 9868 2851 9869
rect 2843 9864 2845 9868
rect 2849 9864 2851 9868
rect 2779 9863 2787 9864
rect 2779 9859 2781 9863
rect 2785 9859 2787 9863
rect 2779 9858 2787 9859
rect 2843 9863 2851 9864
rect 2843 9859 2845 9863
rect 2849 9859 2851 9863
rect 2843 9858 2851 9859
rect 2779 9856 2851 9858
rect 2779 9852 2781 9856
rect 2785 9852 2788 9856
rect 2792 9852 2793 9856
rect 2797 9852 2798 9856
rect 2802 9852 2803 9856
rect 2807 9852 2808 9856
rect 2812 9852 2813 9856
rect 2817 9852 2818 9856
rect 2822 9852 2823 9856
rect 2827 9852 2828 9856
rect 2832 9852 2833 9856
rect 2837 9852 2838 9856
rect 2842 9852 2845 9856
rect 2849 9852 2851 9856
rect 2779 9850 2851 9852
rect 2916 9978 3012 9979
rect 2916 9974 2917 9978
rect 2921 9974 2922 9978
rect 2926 9974 2927 9978
rect 2931 9974 2932 9978
rect 2936 9974 2937 9978
rect 2941 9974 2942 9978
rect 2946 9974 2947 9978
rect 2951 9974 2952 9978
rect 2956 9974 2957 9978
rect 2961 9974 2962 9978
rect 2966 9974 2967 9978
rect 2971 9974 2972 9978
rect 2976 9974 2977 9978
rect 2981 9974 2982 9978
rect 2986 9974 2987 9978
rect 2991 9974 2992 9978
rect 2996 9974 2997 9978
rect 3001 9974 3002 9978
rect 3006 9974 3007 9978
rect 3011 9974 3012 9978
rect 2916 9973 3012 9974
rect 2916 9969 2917 9973
rect 2921 9969 2922 9973
rect 2916 9968 2922 9969
rect 2916 9964 2917 9968
rect 2921 9964 2922 9968
rect 3006 9969 3007 9973
rect 3011 9969 3012 9973
rect 3006 9968 3012 9969
rect 2916 9963 2922 9964
rect 2916 9959 2917 9963
rect 2921 9959 2922 9963
rect 2916 9958 2922 9959
rect 2916 9954 2917 9958
rect 2921 9954 2922 9958
rect 2916 9953 2922 9954
rect 2916 9949 2917 9953
rect 2921 9949 2922 9953
rect 2916 9948 2922 9949
rect 2916 9944 2917 9948
rect 2921 9944 2922 9948
rect 2916 9943 2922 9944
rect 2916 9939 2917 9943
rect 2921 9939 2922 9943
rect 2916 9938 2922 9939
rect 2916 9934 2917 9938
rect 2921 9934 2922 9938
rect 2916 9933 2922 9934
rect 2916 9929 2917 9933
rect 2921 9929 2922 9933
rect 2916 9928 2922 9929
rect 2916 9924 2917 9928
rect 2921 9924 2922 9928
rect 2916 9923 2922 9924
rect 2916 9919 2917 9923
rect 2921 9919 2922 9923
rect 2916 9918 2922 9919
rect 2916 9914 2917 9918
rect 2921 9914 2922 9918
rect 2916 9913 2922 9914
rect 2916 9909 2917 9913
rect 2921 9909 2922 9913
rect 2916 9908 2922 9909
rect 2916 9904 2917 9908
rect 2921 9904 2922 9908
rect 2916 9903 2922 9904
rect 2916 9899 2917 9903
rect 2921 9899 2922 9903
rect 2916 9898 2922 9899
rect 2916 9894 2917 9898
rect 2921 9894 2922 9898
rect 2916 9893 2922 9894
rect 2916 9889 2917 9893
rect 2921 9889 2922 9893
rect 2916 9888 2922 9889
rect 2916 9884 2917 9888
rect 2921 9884 2922 9888
rect 2916 9883 2922 9884
rect 2916 9879 2917 9883
rect 2921 9879 2922 9883
rect 2916 9878 2922 9879
rect 2916 9874 2917 9878
rect 2921 9874 2922 9878
rect 2916 9873 2922 9874
rect 2916 9869 2917 9873
rect 2921 9869 2922 9873
rect 2916 9868 2922 9869
rect 2916 9864 2917 9868
rect 2921 9864 2922 9868
rect 2916 9863 2922 9864
rect 2916 9859 2917 9863
rect 2921 9859 2922 9863
rect 2916 9858 2922 9859
rect 2916 9854 2917 9858
rect 2921 9854 2922 9858
rect 2916 9853 2922 9854
rect 2916 9849 2917 9853
rect 2921 9849 2922 9853
rect 3006 9964 3007 9968
rect 3011 9964 3012 9968
rect 3006 9963 3012 9964
rect 3006 9959 3007 9963
rect 3011 9959 3012 9963
rect 3006 9958 3012 9959
rect 3006 9954 3007 9958
rect 3011 9954 3012 9958
rect 3006 9953 3012 9954
rect 3006 9949 3007 9953
rect 3011 9949 3012 9953
rect 3006 9948 3012 9949
rect 3006 9944 3007 9948
rect 3011 9944 3012 9948
rect 3006 9943 3012 9944
rect 3006 9939 3007 9943
rect 3011 9939 3012 9943
rect 3006 9938 3012 9939
rect 3006 9934 3007 9938
rect 3011 9934 3012 9938
rect 3006 9933 3012 9934
rect 3006 9929 3007 9933
rect 3011 9929 3012 9933
rect 3006 9928 3012 9929
rect 3006 9924 3007 9928
rect 3011 9924 3012 9928
rect 3006 9923 3012 9924
rect 3006 9919 3007 9923
rect 3011 9919 3012 9923
rect 3006 9918 3012 9919
rect 3006 9914 3007 9918
rect 3011 9914 3012 9918
rect 3006 9913 3012 9914
rect 3006 9909 3007 9913
rect 3011 9909 3012 9913
rect 3006 9908 3012 9909
rect 3006 9904 3007 9908
rect 3011 9904 3012 9908
rect 3006 9903 3012 9904
rect 3006 9899 3007 9903
rect 3011 9899 3012 9903
rect 3006 9898 3012 9899
rect 3006 9894 3007 9898
rect 3011 9894 3012 9898
rect 3006 9893 3012 9894
rect 3006 9889 3007 9893
rect 3011 9889 3012 9893
rect 3006 9888 3012 9889
rect 3006 9884 3007 9888
rect 3011 9884 3012 9888
rect 3006 9883 3012 9884
rect 3006 9879 3007 9883
rect 3011 9879 3012 9883
rect 3006 9878 3012 9879
rect 3006 9874 3007 9878
rect 3011 9874 3012 9878
rect 3006 9873 3012 9874
rect 3006 9869 3007 9873
rect 3011 9869 3012 9873
rect 3006 9868 3012 9869
rect 3006 9864 3007 9868
rect 3011 9864 3012 9868
rect 3006 9863 3012 9864
rect 3006 9859 3007 9863
rect 3011 9859 3012 9863
rect 3006 9858 3012 9859
rect 3006 9854 3007 9858
rect 3011 9854 3012 9858
rect 3006 9853 3012 9854
rect 2916 9848 2922 9849
rect 2916 9844 2917 9848
rect 2921 9844 2922 9848
rect 3006 9849 3007 9853
rect 3011 9849 3012 9853
rect 3006 9848 3012 9849
rect 3006 9844 3007 9848
rect 3011 9844 3012 9848
rect 2916 9843 3012 9844
rect 2916 9839 2917 9843
rect 2921 9839 2922 9843
rect 2926 9839 2927 9843
rect 2931 9839 2932 9843
rect 2936 9839 2937 9843
rect 2941 9839 2942 9843
rect 2946 9839 2947 9843
rect 2951 9839 2952 9843
rect 2956 9839 2957 9843
rect 2961 9839 2962 9843
rect 2966 9839 2967 9843
rect 2971 9839 2972 9843
rect 2976 9839 2977 9843
rect 2981 9839 2982 9843
rect 2986 9839 2987 9843
rect 2991 9839 2992 9843
rect 2996 9839 2997 9843
rect 3001 9839 3002 9843
rect 3006 9839 3007 9843
rect 3011 9839 3012 9843
rect 2916 9838 3012 9839
rect 3088 9965 3160 9967
rect 3088 9961 3090 9965
rect 3094 9961 3097 9965
rect 3101 9961 3102 9965
rect 3106 9961 3107 9965
rect 3111 9961 3112 9965
rect 3116 9961 3117 9965
rect 3121 9961 3122 9965
rect 3126 9961 3127 9965
rect 3131 9961 3132 9965
rect 3136 9961 3137 9965
rect 3141 9961 3142 9965
rect 3146 9961 3147 9965
rect 3151 9961 3154 9965
rect 3158 9961 3160 9965
rect 3088 9959 3160 9961
rect 3088 9958 3096 9959
rect 3088 9954 3090 9958
rect 3094 9954 3096 9958
rect 3088 9953 3096 9954
rect 3152 9958 3160 9959
rect 3152 9954 3154 9958
rect 3158 9954 3160 9958
rect 3152 9953 3160 9954
rect 3088 9949 3090 9953
rect 3094 9949 3096 9953
rect 3088 9948 3096 9949
rect 3088 9944 3090 9948
rect 3094 9944 3096 9948
rect 3088 9943 3096 9944
rect 3088 9939 3090 9943
rect 3094 9939 3096 9943
rect 3088 9938 3096 9939
rect 3088 9934 3090 9938
rect 3094 9934 3096 9938
rect 3088 9933 3096 9934
rect 3088 9929 3090 9933
rect 3094 9929 3096 9933
rect 3088 9928 3096 9929
rect 3088 9924 3090 9928
rect 3094 9924 3096 9928
rect 3088 9923 3096 9924
rect 3088 9919 3090 9923
rect 3094 9919 3096 9923
rect 3088 9918 3096 9919
rect 3088 9914 3090 9918
rect 3094 9914 3096 9918
rect 3088 9913 3096 9914
rect 3088 9909 3090 9913
rect 3094 9909 3096 9913
rect 3088 9908 3096 9909
rect 3088 9904 3090 9908
rect 3094 9904 3096 9908
rect 3088 9903 3096 9904
rect 3088 9899 3090 9903
rect 3094 9899 3096 9903
rect 3088 9898 3096 9899
rect 3088 9894 3090 9898
rect 3094 9894 3096 9898
rect 3088 9893 3096 9894
rect 3088 9889 3090 9893
rect 3094 9889 3096 9893
rect 3088 9888 3096 9889
rect 3088 9884 3090 9888
rect 3094 9884 3096 9888
rect 3088 9883 3096 9884
rect 3088 9879 3090 9883
rect 3094 9879 3096 9883
rect 3088 9878 3096 9879
rect 3088 9874 3090 9878
rect 3094 9874 3096 9878
rect 3088 9873 3096 9874
rect 3088 9869 3090 9873
rect 3094 9869 3096 9873
rect 3088 9868 3096 9869
rect 3088 9864 3090 9868
rect 3094 9864 3096 9868
rect 3152 9949 3154 9953
rect 3158 9949 3160 9953
rect 3152 9948 3160 9949
rect 3152 9944 3154 9948
rect 3158 9944 3160 9948
rect 3152 9943 3160 9944
rect 3152 9939 3154 9943
rect 3158 9939 3160 9943
rect 3152 9938 3160 9939
rect 3152 9934 3154 9938
rect 3158 9934 3160 9938
rect 3152 9933 3160 9934
rect 3152 9929 3154 9933
rect 3158 9929 3160 9933
rect 3152 9928 3160 9929
rect 3152 9924 3154 9928
rect 3158 9924 3160 9928
rect 3152 9923 3160 9924
rect 3152 9919 3154 9923
rect 3158 9919 3160 9923
rect 3152 9918 3160 9919
rect 3152 9914 3154 9918
rect 3158 9914 3160 9918
rect 3152 9913 3160 9914
rect 3152 9909 3154 9913
rect 3158 9909 3160 9913
rect 3152 9908 3160 9909
rect 3152 9904 3154 9908
rect 3158 9904 3160 9908
rect 3152 9903 3160 9904
rect 3152 9899 3154 9903
rect 3158 9899 3160 9903
rect 3152 9898 3160 9899
rect 3152 9894 3154 9898
rect 3158 9894 3160 9898
rect 3152 9893 3160 9894
rect 3152 9889 3154 9893
rect 3158 9889 3160 9893
rect 3152 9888 3160 9889
rect 3152 9884 3154 9888
rect 3158 9884 3160 9888
rect 3152 9883 3160 9884
rect 3152 9879 3154 9883
rect 3158 9879 3160 9883
rect 3152 9878 3160 9879
rect 3152 9874 3154 9878
rect 3158 9874 3160 9878
rect 3152 9873 3160 9874
rect 3152 9869 3154 9873
rect 3158 9869 3160 9873
rect 3152 9868 3160 9869
rect 3152 9864 3154 9868
rect 3158 9864 3160 9868
rect 3088 9863 3096 9864
rect 3088 9859 3090 9863
rect 3094 9859 3096 9863
rect 3088 9858 3096 9859
rect 3152 9863 3160 9864
rect 3152 9859 3154 9863
rect 3158 9859 3160 9863
rect 3152 9858 3160 9859
rect 3088 9856 3160 9858
rect 3088 9852 3090 9856
rect 3094 9852 3097 9856
rect 3101 9852 3102 9856
rect 3106 9852 3107 9856
rect 3111 9852 3112 9856
rect 3116 9852 3117 9856
rect 3121 9852 3122 9856
rect 3126 9852 3127 9856
rect 3131 9852 3132 9856
rect 3136 9852 3137 9856
rect 3141 9852 3142 9856
rect 3146 9852 3147 9856
rect 3151 9852 3154 9856
rect 3158 9852 3160 9856
rect 3088 9850 3160 9852
rect 3225 9978 3321 9979
rect 3225 9974 3226 9978
rect 3230 9974 3231 9978
rect 3235 9974 3236 9978
rect 3240 9974 3241 9978
rect 3245 9974 3246 9978
rect 3250 9974 3251 9978
rect 3255 9974 3256 9978
rect 3260 9974 3261 9978
rect 3265 9974 3266 9978
rect 3270 9974 3271 9978
rect 3275 9974 3276 9978
rect 3280 9974 3281 9978
rect 3285 9974 3286 9978
rect 3290 9974 3291 9978
rect 3295 9974 3296 9978
rect 3300 9974 3301 9978
rect 3305 9974 3306 9978
rect 3310 9974 3311 9978
rect 3315 9974 3316 9978
rect 3320 9974 3321 9978
rect 3225 9973 3321 9974
rect 3225 9969 3226 9973
rect 3230 9969 3231 9973
rect 3225 9968 3231 9969
rect 3225 9964 3226 9968
rect 3230 9964 3231 9968
rect 3315 9969 3316 9973
rect 3320 9969 3321 9973
rect 3315 9968 3321 9969
rect 3225 9963 3231 9964
rect 3225 9959 3226 9963
rect 3230 9959 3231 9963
rect 3225 9958 3231 9959
rect 3225 9954 3226 9958
rect 3230 9954 3231 9958
rect 3225 9953 3231 9954
rect 3225 9949 3226 9953
rect 3230 9949 3231 9953
rect 3225 9948 3231 9949
rect 3225 9944 3226 9948
rect 3230 9944 3231 9948
rect 3225 9943 3231 9944
rect 3225 9939 3226 9943
rect 3230 9939 3231 9943
rect 3225 9938 3231 9939
rect 3225 9934 3226 9938
rect 3230 9934 3231 9938
rect 3225 9933 3231 9934
rect 3225 9929 3226 9933
rect 3230 9929 3231 9933
rect 3225 9928 3231 9929
rect 3225 9924 3226 9928
rect 3230 9924 3231 9928
rect 3225 9923 3231 9924
rect 3225 9919 3226 9923
rect 3230 9919 3231 9923
rect 3225 9918 3231 9919
rect 3225 9914 3226 9918
rect 3230 9914 3231 9918
rect 3225 9913 3231 9914
rect 3225 9909 3226 9913
rect 3230 9909 3231 9913
rect 3225 9908 3231 9909
rect 3225 9904 3226 9908
rect 3230 9904 3231 9908
rect 3225 9903 3231 9904
rect 3225 9899 3226 9903
rect 3230 9899 3231 9903
rect 3225 9898 3231 9899
rect 3225 9894 3226 9898
rect 3230 9894 3231 9898
rect 3225 9893 3231 9894
rect 3225 9889 3226 9893
rect 3230 9889 3231 9893
rect 3225 9888 3231 9889
rect 3225 9884 3226 9888
rect 3230 9884 3231 9888
rect 3225 9883 3231 9884
rect 3225 9879 3226 9883
rect 3230 9879 3231 9883
rect 3225 9878 3231 9879
rect 3225 9874 3226 9878
rect 3230 9874 3231 9878
rect 3225 9873 3231 9874
rect 3225 9869 3226 9873
rect 3230 9869 3231 9873
rect 3225 9868 3231 9869
rect 3225 9864 3226 9868
rect 3230 9864 3231 9868
rect 3225 9863 3231 9864
rect 3225 9859 3226 9863
rect 3230 9859 3231 9863
rect 3225 9858 3231 9859
rect 3225 9854 3226 9858
rect 3230 9854 3231 9858
rect 3225 9853 3231 9854
rect 3225 9849 3226 9853
rect 3230 9849 3231 9853
rect 3315 9964 3316 9968
rect 3320 9964 3321 9968
rect 3315 9963 3321 9964
rect 3315 9959 3316 9963
rect 3320 9959 3321 9963
rect 3315 9958 3321 9959
rect 3315 9954 3316 9958
rect 3320 9954 3321 9958
rect 3315 9953 3321 9954
rect 3315 9949 3316 9953
rect 3320 9949 3321 9953
rect 3315 9948 3321 9949
rect 3315 9944 3316 9948
rect 3320 9944 3321 9948
rect 3315 9943 3321 9944
rect 3315 9939 3316 9943
rect 3320 9939 3321 9943
rect 3315 9938 3321 9939
rect 3315 9934 3316 9938
rect 3320 9934 3321 9938
rect 3315 9933 3321 9934
rect 3315 9929 3316 9933
rect 3320 9929 3321 9933
rect 3315 9928 3321 9929
rect 3315 9924 3316 9928
rect 3320 9924 3321 9928
rect 3315 9923 3321 9924
rect 3315 9919 3316 9923
rect 3320 9919 3321 9923
rect 3315 9918 3321 9919
rect 3315 9914 3316 9918
rect 3320 9914 3321 9918
rect 3315 9913 3321 9914
rect 3315 9909 3316 9913
rect 3320 9909 3321 9913
rect 3315 9908 3321 9909
rect 3315 9904 3316 9908
rect 3320 9904 3321 9908
rect 3315 9903 3321 9904
rect 3315 9899 3316 9903
rect 3320 9899 3321 9903
rect 3315 9898 3321 9899
rect 3315 9894 3316 9898
rect 3320 9894 3321 9898
rect 3315 9893 3321 9894
rect 3315 9889 3316 9893
rect 3320 9889 3321 9893
rect 3315 9888 3321 9889
rect 3315 9884 3316 9888
rect 3320 9884 3321 9888
rect 3315 9883 3321 9884
rect 3315 9879 3316 9883
rect 3320 9879 3321 9883
rect 3315 9878 3321 9879
rect 3315 9874 3316 9878
rect 3320 9874 3321 9878
rect 3315 9873 3321 9874
rect 3315 9869 3316 9873
rect 3320 9869 3321 9873
rect 3315 9868 3321 9869
rect 3315 9864 3316 9868
rect 3320 9864 3321 9868
rect 3315 9863 3321 9864
rect 3315 9859 3316 9863
rect 3320 9859 3321 9863
rect 3315 9858 3321 9859
rect 3315 9854 3316 9858
rect 3320 9854 3321 9858
rect 3315 9853 3321 9854
rect 3225 9848 3231 9849
rect 3225 9844 3226 9848
rect 3230 9844 3231 9848
rect 3315 9849 3316 9853
rect 3320 9849 3321 9853
rect 3315 9848 3321 9849
rect 3315 9844 3316 9848
rect 3320 9844 3321 9848
rect 3225 9843 3321 9844
rect 3225 9839 3226 9843
rect 3230 9839 3231 9843
rect 3235 9839 3236 9843
rect 3240 9839 3241 9843
rect 3245 9839 3246 9843
rect 3250 9839 3251 9843
rect 3255 9839 3256 9843
rect 3260 9839 3261 9843
rect 3265 9839 3266 9843
rect 3270 9839 3271 9843
rect 3275 9839 3276 9843
rect 3280 9839 3281 9843
rect 3285 9839 3286 9843
rect 3290 9839 3291 9843
rect 3295 9839 3296 9843
rect 3300 9839 3301 9843
rect 3305 9839 3306 9843
rect 3310 9839 3311 9843
rect 3315 9839 3316 9843
rect 3320 9839 3321 9843
rect 3225 9838 3321 9839
rect 3397 9965 3469 9967
rect 3397 9961 3399 9965
rect 3403 9961 3406 9965
rect 3410 9961 3411 9965
rect 3415 9961 3416 9965
rect 3420 9961 3421 9965
rect 3425 9961 3426 9965
rect 3430 9961 3431 9965
rect 3435 9961 3436 9965
rect 3440 9961 3441 9965
rect 3445 9961 3446 9965
rect 3450 9961 3451 9965
rect 3455 9961 3456 9965
rect 3460 9961 3463 9965
rect 3467 9961 3469 9965
rect 3397 9959 3469 9961
rect 3397 9958 3405 9959
rect 3397 9954 3399 9958
rect 3403 9954 3405 9958
rect 3397 9953 3405 9954
rect 3461 9958 3469 9959
rect 3461 9954 3463 9958
rect 3467 9954 3469 9958
rect 3461 9953 3469 9954
rect 3397 9949 3399 9953
rect 3403 9949 3405 9953
rect 3397 9948 3405 9949
rect 3397 9944 3399 9948
rect 3403 9944 3405 9948
rect 3397 9943 3405 9944
rect 3397 9939 3399 9943
rect 3403 9939 3405 9943
rect 3397 9938 3405 9939
rect 3397 9934 3399 9938
rect 3403 9934 3405 9938
rect 3397 9933 3405 9934
rect 3397 9929 3399 9933
rect 3403 9929 3405 9933
rect 3397 9928 3405 9929
rect 3397 9924 3399 9928
rect 3403 9924 3405 9928
rect 3397 9923 3405 9924
rect 3397 9919 3399 9923
rect 3403 9919 3405 9923
rect 3397 9918 3405 9919
rect 3397 9914 3399 9918
rect 3403 9914 3405 9918
rect 3397 9913 3405 9914
rect 3397 9909 3399 9913
rect 3403 9909 3405 9913
rect 3397 9908 3405 9909
rect 3397 9904 3399 9908
rect 3403 9904 3405 9908
rect 3397 9903 3405 9904
rect 3397 9899 3399 9903
rect 3403 9899 3405 9903
rect 3397 9898 3405 9899
rect 3397 9894 3399 9898
rect 3403 9894 3405 9898
rect 3397 9893 3405 9894
rect 3397 9889 3399 9893
rect 3403 9889 3405 9893
rect 3397 9888 3405 9889
rect 3397 9884 3399 9888
rect 3403 9884 3405 9888
rect 3397 9883 3405 9884
rect 3397 9879 3399 9883
rect 3403 9879 3405 9883
rect 3397 9878 3405 9879
rect 3397 9874 3399 9878
rect 3403 9874 3405 9878
rect 3397 9873 3405 9874
rect 3397 9869 3399 9873
rect 3403 9869 3405 9873
rect 3397 9868 3405 9869
rect 3397 9864 3399 9868
rect 3403 9864 3405 9868
rect 3461 9949 3463 9953
rect 3467 9949 3469 9953
rect 3461 9948 3469 9949
rect 3461 9944 3463 9948
rect 3467 9944 3469 9948
rect 3461 9943 3469 9944
rect 3461 9939 3463 9943
rect 3467 9939 3469 9943
rect 3461 9938 3469 9939
rect 3461 9934 3463 9938
rect 3467 9934 3469 9938
rect 3461 9933 3469 9934
rect 3461 9929 3463 9933
rect 3467 9929 3469 9933
rect 3461 9928 3469 9929
rect 3461 9924 3463 9928
rect 3467 9924 3469 9928
rect 3461 9923 3469 9924
rect 3461 9919 3463 9923
rect 3467 9919 3469 9923
rect 3461 9918 3469 9919
rect 3461 9914 3463 9918
rect 3467 9914 3469 9918
rect 3461 9913 3469 9914
rect 3461 9909 3463 9913
rect 3467 9909 3469 9913
rect 3461 9908 3469 9909
rect 3461 9904 3463 9908
rect 3467 9904 3469 9908
rect 3461 9903 3469 9904
rect 3461 9899 3463 9903
rect 3467 9899 3469 9903
rect 3461 9898 3469 9899
rect 3461 9894 3463 9898
rect 3467 9894 3469 9898
rect 3461 9893 3469 9894
rect 3461 9889 3463 9893
rect 3467 9889 3469 9893
rect 3461 9888 3469 9889
rect 3461 9884 3463 9888
rect 3467 9884 3469 9888
rect 3461 9883 3469 9884
rect 3461 9879 3463 9883
rect 3467 9879 3469 9883
rect 3461 9878 3469 9879
rect 3461 9874 3463 9878
rect 3467 9874 3469 9878
rect 3461 9873 3469 9874
rect 3461 9869 3463 9873
rect 3467 9869 3469 9873
rect 3461 9868 3469 9869
rect 3461 9864 3463 9868
rect 3467 9864 3469 9868
rect 3397 9863 3405 9864
rect 3397 9859 3399 9863
rect 3403 9859 3405 9863
rect 3397 9858 3405 9859
rect 3461 9863 3469 9864
rect 3461 9859 3463 9863
rect 3467 9859 3469 9863
rect 3461 9858 3469 9859
rect 3397 9856 3469 9858
rect 3397 9852 3399 9856
rect 3403 9852 3406 9856
rect 3410 9852 3411 9856
rect 3415 9852 3416 9856
rect 3420 9852 3421 9856
rect 3425 9852 3426 9856
rect 3430 9852 3431 9856
rect 3435 9852 3436 9856
rect 3440 9852 3441 9856
rect 3445 9852 3446 9856
rect 3450 9852 3451 9856
rect 3455 9852 3456 9856
rect 3460 9852 3463 9856
rect 3467 9852 3469 9856
rect 3397 9850 3469 9852
rect 3534 9978 3630 9979
rect 3534 9974 3535 9978
rect 3539 9974 3540 9978
rect 3544 9974 3545 9978
rect 3549 9974 3550 9978
rect 3554 9974 3555 9978
rect 3559 9974 3560 9978
rect 3564 9974 3565 9978
rect 3569 9974 3570 9978
rect 3574 9974 3575 9978
rect 3579 9974 3580 9978
rect 3584 9974 3585 9978
rect 3589 9974 3590 9978
rect 3594 9974 3595 9978
rect 3599 9974 3600 9978
rect 3604 9974 3605 9978
rect 3609 9974 3610 9978
rect 3614 9974 3615 9978
rect 3619 9974 3620 9978
rect 3624 9974 3625 9978
rect 3629 9974 3630 9978
rect 3534 9973 3630 9974
rect 3534 9969 3535 9973
rect 3539 9969 3540 9973
rect 3534 9968 3540 9969
rect 3534 9964 3535 9968
rect 3539 9964 3540 9968
rect 3624 9969 3625 9973
rect 3629 9969 3630 9973
rect 3624 9968 3630 9969
rect 3534 9963 3540 9964
rect 3534 9959 3535 9963
rect 3539 9959 3540 9963
rect 3534 9958 3540 9959
rect 3534 9954 3535 9958
rect 3539 9954 3540 9958
rect 3534 9953 3540 9954
rect 3534 9949 3535 9953
rect 3539 9949 3540 9953
rect 3534 9948 3540 9949
rect 3534 9944 3535 9948
rect 3539 9944 3540 9948
rect 3534 9943 3540 9944
rect 3534 9939 3535 9943
rect 3539 9939 3540 9943
rect 3534 9938 3540 9939
rect 3534 9934 3535 9938
rect 3539 9934 3540 9938
rect 3534 9933 3540 9934
rect 3534 9929 3535 9933
rect 3539 9929 3540 9933
rect 3534 9928 3540 9929
rect 3534 9924 3535 9928
rect 3539 9924 3540 9928
rect 3534 9923 3540 9924
rect 3534 9919 3535 9923
rect 3539 9919 3540 9923
rect 3534 9918 3540 9919
rect 3534 9914 3535 9918
rect 3539 9914 3540 9918
rect 3534 9913 3540 9914
rect 3534 9909 3535 9913
rect 3539 9909 3540 9913
rect 3534 9908 3540 9909
rect 3534 9904 3535 9908
rect 3539 9904 3540 9908
rect 3534 9903 3540 9904
rect 3534 9899 3535 9903
rect 3539 9899 3540 9903
rect 3534 9898 3540 9899
rect 3534 9894 3535 9898
rect 3539 9894 3540 9898
rect 3534 9893 3540 9894
rect 3534 9889 3535 9893
rect 3539 9889 3540 9893
rect 3534 9888 3540 9889
rect 3534 9884 3535 9888
rect 3539 9884 3540 9888
rect 3534 9883 3540 9884
rect 3534 9879 3535 9883
rect 3539 9879 3540 9883
rect 3534 9878 3540 9879
rect 3534 9874 3535 9878
rect 3539 9874 3540 9878
rect 3534 9873 3540 9874
rect 3534 9869 3535 9873
rect 3539 9869 3540 9873
rect 3534 9868 3540 9869
rect 3534 9864 3535 9868
rect 3539 9864 3540 9868
rect 3534 9863 3540 9864
rect 3534 9859 3535 9863
rect 3539 9859 3540 9863
rect 3534 9858 3540 9859
rect 3534 9854 3535 9858
rect 3539 9854 3540 9858
rect 3534 9853 3540 9854
rect 3534 9849 3535 9853
rect 3539 9849 3540 9853
rect 3624 9964 3625 9968
rect 3629 9964 3630 9968
rect 3624 9963 3630 9964
rect 3624 9959 3625 9963
rect 3629 9959 3630 9963
rect 3624 9958 3630 9959
rect 3624 9954 3625 9958
rect 3629 9954 3630 9958
rect 3624 9953 3630 9954
rect 3624 9949 3625 9953
rect 3629 9949 3630 9953
rect 3624 9948 3630 9949
rect 3624 9944 3625 9948
rect 3629 9944 3630 9948
rect 3624 9943 3630 9944
rect 3624 9939 3625 9943
rect 3629 9939 3630 9943
rect 3624 9938 3630 9939
rect 3624 9934 3625 9938
rect 3629 9934 3630 9938
rect 3624 9933 3630 9934
rect 3624 9929 3625 9933
rect 3629 9929 3630 9933
rect 3624 9928 3630 9929
rect 3624 9924 3625 9928
rect 3629 9924 3630 9928
rect 3624 9923 3630 9924
rect 3624 9919 3625 9923
rect 3629 9919 3630 9923
rect 3624 9918 3630 9919
rect 3624 9914 3625 9918
rect 3629 9914 3630 9918
rect 3624 9913 3630 9914
rect 3624 9909 3625 9913
rect 3629 9909 3630 9913
rect 3624 9908 3630 9909
rect 3624 9904 3625 9908
rect 3629 9904 3630 9908
rect 3624 9903 3630 9904
rect 3624 9899 3625 9903
rect 3629 9899 3630 9903
rect 3624 9898 3630 9899
rect 3624 9894 3625 9898
rect 3629 9894 3630 9898
rect 3624 9893 3630 9894
rect 3624 9889 3625 9893
rect 3629 9889 3630 9893
rect 3624 9888 3630 9889
rect 3624 9884 3625 9888
rect 3629 9884 3630 9888
rect 3624 9883 3630 9884
rect 3624 9879 3625 9883
rect 3629 9879 3630 9883
rect 3624 9878 3630 9879
rect 3624 9874 3625 9878
rect 3629 9874 3630 9878
rect 3624 9873 3630 9874
rect 3624 9869 3625 9873
rect 3629 9869 3630 9873
rect 3624 9868 3630 9869
rect 3624 9864 3625 9868
rect 3629 9864 3630 9868
rect 3624 9863 3630 9864
rect 3624 9859 3625 9863
rect 3629 9859 3630 9863
rect 3624 9858 3630 9859
rect 3624 9854 3625 9858
rect 3629 9854 3630 9858
rect 3624 9853 3630 9854
rect 3534 9848 3540 9849
rect 3534 9844 3535 9848
rect 3539 9844 3540 9848
rect 3624 9849 3625 9853
rect 3629 9849 3630 9853
rect 3624 9848 3630 9849
rect 3624 9844 3625 9848
rect 3629 9844 3630 9848
rect 3534 9843 3630 9844
rect 3534 9839 3535 9843
rect 3539 9839 3540 9843
rect 3544 9839 3545 9843
rect 3549 9839 3550 9843
rect 3554 9839 3555 9843
rect 3559 9839 3560 9843
rect 3564 9839 3565 9843
rect 3569 9839 3570 9843
rect 3574 9839 3575 9843
rect 3579 9839 3580 9843
rect 3584 9839 3585 9843
rect 3589 9839 3590 9843
rect 3594 9839 3595 9843
rect 3599 9839 3600 9843
rect 3604 9839 3605 9843
rect 3609 9839 3610 9843
rect 3614 9839 3615 9843
rect 3619 9839 3620 9843
rect 3624 9839 3625 9843
rect 3629 9839 3630 9843
rect 3534 9838 3630 9839
rect 3706 9965 3778 9967
rect 3706 9961 3708 9965
rect 3712 9961 3715 9965
rect 3719 9961 3720 9965
rect 3724 9961 3725 9965
rect 3729 9961 3730 9965
rect 3734 9961 3735 9965
rect 3739 9961 3740 9965
rect 3744 9961 3745 9965
rect 3749 9961 3750 9965
rect 3754 9961 3755 9965
rect 3759 9961 3760 9965
rect 3764 9961 3765 9965
rect 3769 9961 3772 9965
rect 3776 9961 3778 9965
rect 3706 9959 3778 9961
rect 3706 9958 3714 9959
rect 3706 9954 3708 9958
rect 3712 9954 3714 9958
rect 3706 9953 3714 9954
rect 3770 9958 3778 9959
rect 3770 9954 3772 9958
rect 3776 9954 3778 9958
rect 3770 9953 3778 9954
rect 3706 9949 3708 9953
rect 3712 9949 3714 9953
rect 3706 9948 3714 9949
rect 3706 9944 3708 9948
rect 3712 9944 3714 9948
rect 3706 9943 3714 9944
rect 3706 9939 3708 9943
rect 3712 9939 3714 9943
rect 3706 9938 3714 9939
rect 3706 9934 3708 9938
rect 3712 9934 3714 9938
rect 3706 9933 3714 9934
rect 3706 9929 3708 9933
rect 3712 9929 3714 9933
rect 3706 9928 3714 9929
rect 3706 9924 3708 9928
rect 3712 9924 3714 9928
rect 3706 9923 3714 9924
rect 3706 9919 3708 9923
rect 3712 9919 3714 9923
rect 3706 9918 3714 9919
rect 3706 9914 3708 9918
rect 3712 9914 3714 9918
rect 3706 9913 3714 9914
rect 3706 9909 3708 9913
rect 3712 9909 3714 9913
rect 3706 9908 3714 9909
rect 3706 9904 3708 9908
rect 3712 9904 3714 9908
rect 3706 9903 3714 9904
rect 3706 9899 3708 9903
rect 3712 9899 3714 9903
rect 3706 9898 3714 9899
rect 3706 9894 3708 9898
rect 3712 9894 3714 9898
rect 3706 9893 3714 9894
rect 3706 9889 3708 9893
rect 3712 9889 3714 9893
rect 3706 9888 3714 9889
rect 3706 9884 3708 9888
rect 3712 9884 3714 9888
rect 3706 9883 3714 9884
rect 3706 9879 3708 9883
rect 3712 9879 3714 9883
rect 3706 9878 3714 9879
rect 3706 9874 3708 9878
rect 3712 9874 3714 9878
rect 3706 9873 3714 9874
rect 3706 9869 3708 9873
rect 3712 9869 3714 9873
rect 3706 9868 3714 9869
rect 3706 9864 3708 9868
rect 3712 9864 3714 9868
rect 3770 9949 3772 9953
rect 3776 9949 3778 9953
rect 3770 9948 3778 9949
rect 3770 9944 3772 9948
rect 3776 9944 3778 9948
rect 3770 9943 3778 9944
rect 3770 9939 3772 9943
rect 3776 9939 3778 9943
rect 3770 9938 3778 9939
rect 3770 9934 3772 9938
rect 3776 9934 3778 9938
rect 3770 9933 3778 9934
rect 3770 9929 3772 9933
rect 3776 9929 3778 9933
rect 3770 9928 3778 9929
rect 3770 9924 3772 9928
rect 3776 9924 3778 9928
rect 3770 9923 3778 9924
rect 3770 9919 3772 9923
rect 3776 9919 3778 9923
rect 3770 9918 3778 9919
rect 3770 9914 3772 9918
rect 3776 9914 3778 9918
rect 3770 9913 3778 9914
rect 3770 9909 3772 9913
rect 3776 9909 3778 9913
rect 3770 9908 3778 9909
rect 3770 9904 3772 9908
rect 3776 9904 3778 9908
rect 3770 9903 3778 9904
rect 3770 9899 3772 9903
rect 3776 9899 3778 9903
rect 3770 9898 3778 9899
rect 3770 9894 3772 9898
rect 3776 9894 3778 9898
rect 3770 9893 3778 9894
rect 3770 9889 3772 9893
rect 3776 9889 3778 9893
rect 3770 9888 3778 9889
rect 3770 9884 3772 9888
rect 3776 9884 3778 9888
rect 3770 9883 3778 9884
rect 3770 9879 3772 9883
rect 3776 9879 3778 9883
rect 3770 9878 3778 9879
rect 3770 9874 3772 9878
rect 3776 9874 3778 9878
rect 3770 9873 3778 9874
rect 3770 9869 3772 9873
rect 3776 9869 3778 9873
rect 3770 9868 3778 9869
rect 3770 9864 3772 9868
rect 3776 9864 3778 9868
rect 3706 9863 3714 9864
rect 3706 9859 3708 9863
rect 3712 9859 3714 9863
rect 3706 9858 3714 9859
rect 3770 9863 3778 9864
rect 3770 9859 3772 9863
rect 3776 9859 3778 9863
rect 3770 9858 3778 9859
rect 3706 9856 3778 9858
rect 3706 9852 3708 9856
rect 3712 9852 3715 9856
rect 3719 9852 3720 9856
rect 3724 9852 3725 9856
rect 3729 9852 3730 9856
rect 3734 9852 3735 9856
rect 3739 9852 3740 9856
rect 3744 9852 3745 9856
rect 3749 9852 3750 9856
rect 3754 9852 3755 9856
rect 3759 9852 3760 9856
rect 3764 9852 3765 9856
rect 3769 9852 3772 9856
rect 3776 9852 3778 9856
rect 3706 9850 3778 9852
rect 3843 9978 3939 9979
rect 3843 9974 3844 9978
rect 3848 9974 3849 9978
rect 3853 9974 3854 9978
rect 3858 9974 3859 9978
rect 3863 9974 3864 9978
rect 3868 9974 3869 9978
rect 3873 9974 3874 9978
rect 3878 9974 3879 9978
rect 3883 9974 3884 9978
rect 3888 9974 3889 9978
rect 3893 9974 3894 9978
rect 3898 9974 3899 9978
rect 3903 9974 3904 9978
rect 3908 9974 3909 9978
rect 3913 9974 3914 9978
rect 3918 9974 3919 9978
rect 3923 9974 3924 9978
rect 3928 9974 3929 9978
rect 3933 9974 3934 9978
rect 3938 9974 3939 9978
rect 3843 9973 3939 9974
rect 3843 9969 3844 9973
rect 3848 9969 3849 9973
rect 3843 9968 3849 9969
rect 3843 9964 3844 9968
rect 3848 9964 3849 9968
rect 3933 9969 3934 9973
rect 3938 9969 3939 9973
rect 3933 9968 3939 9969
rect 3843 9963 3849 9964
rect 3843 9959 3844 9963
rect 3848 9959 3849 9963
rect 3843 9958 3849 9959
rect 3843 9954 3844 9958
rect 3848 9954 3849 9958
rect 3843 9953 3849 9954
rect 3843 9949 3844 9953
rect 3848 9949 3849 9953
rect 3843 9948 3849 9949
rect 3843 9944 3844 9948
rect 3848 9944 3849 9948
rect 3843 9943 3849 9944
rect 3843 9939 3844 9943
rect 3848 9939 3849 9943
rect 3843 9938 3849 9939
rect 3843 9934 3844 9938
rect 3848 9934 3849 9938
rect 3843 9933 3849 9934
rect 3843 9929 3844 9933
rect 3848 9929 3849 9933
rect 3843 9928 3849 9929
rect 3843 9924 3844 9928
rect 3848 9924 3849 9928
rect 3843 9923 3849 9924
rect 3843 9919 3844 9923
rect 3848 9919 3849 9923
rect 3843 9918 3849 9919
rect 3843 9914 3844 9918
rect 3848 9914 3849 9918
rect 3843 9913 3849 9914
rect 3843 9909 3844 9913
rect 3848 9909 3849 9913
rect 3843 9908 3849 9909
rect 3843 9904 3844 9908
rect 3848 9904 3849 9908
rect 3843 9903 3849 9904
rect 3843 9899 3844 9903
rect 3848 9899 3849 9903
rect 3843 9898 3849 9899
rect 3843 9894 3844 9898
rect 3848 9894 3849 9898
rect 3843 9893 3849 9894
rect 3843 9889 3844 9893
rect 3848 9889 3849 9893
rect 3843 9888 3849 9889
rect 3843 9884 3844 9888
rect 3848 9884 3849 9888
rect 3843 9883 3849 9884
rect 3843 9879 3844 9883
rect 3848 9879 3849 9883
rect 3843 9878 3849 9879
rect 3843 9874 3844 9878
rect 3848 9874 3849 9878
rect 3843 9873 3849 9874
rect 3843 9869 3844 9873
rect 3848 9869 3849 9873
rect 3843 9868 3849 9869
rect 3843 9864 3844 9868
rect 3848 9864 3849 9868
rect 3843 9863 3849 9864
rect 3843 9859 3844 9863
rect 3848 9859 3849 9863
rect 3843 9858 3849 9859
rect 3843 9854 3844 9858
rect 3848 9854 3849 9858
rect 3843 9853 3849 9854
rect 3843 9849 3844 9853
rect 3848 9849 3849 9853
rect 3933 9964 3934 9968
rect 3938 9964 3939 9968
rect 3933 9963 3939 9964
rect 3933 9959 3934 9963
rect 3938 9959 3939 9963
rect 3933 9958 3939 9959
rect 3933 9954 3934 9958
rect 3938 9954 3939 9958
rect 3933 9953 3939 9954
rect 3933 9949 3934 9953
rect 3938 9949 3939 9953
rect 3933 9948 3939 9949
rect 3933 9944 3934 9948
rect 3938 9944 3939 9948
rect 3933 9943 3939 9944
rect 3933 9939 3934 9943
rect 3938 9939 3939 9943
rect 3933 9938 3939 9939
rect 3933 9934 3934 9938
rect 3938 9934 3939 9938
rect 3933 9933 3939 9934
rect 3933 9929 3934 9933
rect 3938 9929 3939 9933
rect 3933 9928 3939 9929
rect 3933 9924 3934 9928
rect 3938 9924 3939 9928
rect 3933 9923 3939 9924
rect 3933 9919 3934 9923
rect 3938 9919 3939 9923
rect 3933 9918 3939 9919
rect 3933 9914 3934 9918
rect 3938 9914 3939 9918
rect 3933 9913 3939 9914
rect 3933 9909 3934 9913
rect 3938 9909 3939 9913
rect 3933 9908 3939 9909
rect 3933 9904 3934 9908
rect 3938 9904 3939 9908
rect 3933 9903 3939 9904
rect 3933 9899 3934 9903
rect 3938 9899 3939 9903
rect 3933 9898 3939 9899
rect 3933 9894 3934 9898
rect 3938 9894 3939 9898
rect 3933 9893 3939 9894
rect 3933 9889 3934 9893
rect 3938 9889 3939 9893
rect 3933 9888 3939 9889
rect 3933 9884 3934 9888
rect 3938 9884 3939 9888
rect 3933 9883 3939 9884
rect 3933 9879 3934 9883
rect 3938 9879 3939 9883
rect 3933 9878 3939 9879
rect 3933 9874 3934 9878
rect 3938 9874 3939 9878
rect 3933 9873 3939 9874
rect 3933 9869 3934 9873
rect 3938 9869 3939 9873
rect 3933 9868 3939 9869
rect 3933 9864 3934 9868
rect 3938 9864 3939 9868
rect 3933 9863 3939 9864
rect 3933 9859 3934 9863
rect 3938 9859 3939 9863
rect 3933 9858 3939 9859
rect 3933 9854 3934 9858
rect 3938 9854 3939 9858
rect 3933 9853 3939 9854
rect 3843 9848 3849 9849
rect 3843 9844 3844 9848
rect 3848 9844 3849 9848
rect 3933 9849 3934 9853
rect 3938 9849 3939 9853
rect 3933 9848 3939 9849
rect 3933 9844 3934 9848
rect 3938 9844 3939 9848
rect 3843 9843 3939 9844
rect 3843 9839 3844 9843
rect 3848 9839 3849 9843
rect 3853 9839 3854 9843
rect 3858 9839 3859 9843
rect 3863 9839 3864 9843
rect 3868 9839 3869 9843
rect 3873 9839 3874 9843
rect 3878 9839 3879 9843
rect 3883 9839 3884 9843
rect 3888 9839 3889 9843
rect 3893 9839 3894 9843
rect 3898 9839 3899 9843
rect 3903 9839 3904 9843
rect 3908 9839 3909 9843
rect 3913 9839 3914 9843
rect 3918 9839 3919 9843
rect 3923 9839 3924 9843
rect 3928 9839 3929 9843
rect 3933 9839 3934 9843
rect 3938 9839 3939 9843
rect 3843 9838 3939 9839
rect 4015 9965 4087 9967
rect 4015 9961 4017 9965
rect 4021 9961 4024 9965
rect 4028 9961 4029 9965
rect 4033 9961 4034 9965
rect 4038 9961 4039 9965
rect 4043 9961 4044 9965
rect 4048 9961 4049 9965
rect 4053 9961 4054 9965
rect 4058 9961 4059 9965
rect 4063 9961 4064 9965
rect 4068 9961 4069 9965
rect 4073 9961 4074 9965
rect 4078 9961 4081 9965
rect 4085 9961 4087 9965
rect 4015 9959 4087 9961
rect 4015 9958 4023 9959
rect 4015 9954 4017 9958
rect 4021 9954 4023 9958
rect 4015 9953 4023 9954
rect 4079 9958 4087 9959
rect 4079 9954 4081 9958
rect 4085 9954 4087 9958
rect 4079 9953 4087 9954
rect 4015 9949 4017 9953
rect 4021 9949 4023 9953
rect 4015 9948 4023 9949
rect 4015 9944 4017 9948
rect 4021 9944 4023 9948
rect 4015 9943 4023 9944
rect 4015 9939 4017 9943
rect 4021 9939 4023 9943
rect 4015 9938 4023 9939
rect 4015 9934 4017 9938
rect 4021 9934 4023 9938
rect 4015 9933 4023 9934
rect 4015 9929 4017 9933
rect 4021 9929 4023 9933
rect 4015 9928 4023 9929
rect 4015 9924 4017 9928
rect 4021 9924 4023 9928
rect 4015 9923 4023 9924
rect 4015 9919 4017 9923
rect 4021 9919 4023 9923
rect 4015 9918 4023 9919
rect 4015 9914 4017 9918
rect 4021 9914 4023 9918
rect 4015 9913 4023 9914
rect 4015 9909 4017 9913
rect 4021 9909 4023 9913
rect 4015 9908 4023 9909
rect 4015 9904 4017 9908
rect 4021 9904 4023 9908
rect 4015 9903 4023 9904
rect 4015 9899 4017 9903
rect 4021 9899 4023 9903
rect 4015 9898 4023 9899
rect 4015 9894 4017 9898
rect 4021 9894 4023 9898
rect 4015 9893 4023 9894
rect 4015 9889 4017 9893
rect 4021 9889 4023 9893
rect 4015 9888 4023 9889
rect 4015 9884 4017 9888
rect 4021 9884 4023 9888
rect 4015 9883 4023 9884
rect 4015 9879 4017 9883
rect 4021 9879 4023 9883
rect 4015 9878 4023 9879
rect 4015 9874 4017 9878
rect 4021 9874 4023 9878
rect 4015 9873 4023 9874
rect 4015 9869 4017 9873
rect 4021 9869 4023 9873
rect 4015 9868 4023 9869
rect 4015 9864 4017 9868
rect 4021 9864 4023 9868
rect 4079 9949 4081 9953
rect 4085 9949 4087 9953
rect 4079 9948 4087 9949
rect 4079 9944 4081 9948
rect 4085 9944 4087 9948
rect 4079 9943 4087 9944
rect 4079 9939 4081 9943
rect 4085 9939 4087 9943
rect 4079 9938 4087 9939
rect 4079 9934 4081 9938
rect 4085 9934 4087 9938
rect 4079 9933 4087 9934
rect 4079 9929 4081 9933
rect 4085 9929 4087 9933
rect 4079 9928 4087 9929
rect 4079 9924 4081 9928
rect 4085 9924 4087 9928
rect 4079 9923 4087 9924
rect 4079 9919 4081 9923
rect 4085 9919 4087 9923
rect 4079 9918 4087 9919
rect 4079 9914 4081 9918
rect 4085 9914 4087 9918
rect 4079 9913 4087 9914
rect 4079 9909 4081 9913
rect 4085 9909 4087 9913
rect 4079 9908 4087 9909
rect 4079 9904 4081 9908
rect 4085 9904 4087 9908
rect 4079 9903 4087 9904
rect 4079 9899 4081 9903
rect 4085 9899 4087 9903
rect 4079 9898 4087 9899
rect 4079 9894 4081 9898
rect 4085 9894 4087 9898
rect 4079 9893 4087 9894
rect 4079 9889 4081 9893
rect 4085 9889 4087 9893
rect 4079 9888 4087 9889
rect 4079 9884 4081 9888
rect 4085 9884 4087 9888
rect 4079 9883 4087 9884
rect 4079 9879 4081 9883
rect 4085 9879 4087 9883
rect 4079 9878 4087 9879
rect 4079 9874 4081 9878
rect 4085 9874 4087 9878
rect 4079 9873 4087 9874
rect 4079 9869 4081 9873
rect 4085 9869 4087 9873
rect 4079 9868 4087 9869
rect 4079 9864 4081 9868
rect 4085 9864 4087 9868
rect 4015 9863 4023 9864
rect 4015 9859 4017 9863
rect 4021 9859 4023 9863
rect 4015 9858 4023 9859
rect 4079 9863 4087 9864
rect 4079 9859 4081 9863
rect 4085 9859 4087 9863
rect 4079 9858 4087 9859
rect 4015 9856 4087 9858
rect 4015 9852 4017 9856
rect 4021 9852 4024 9856
rect 4028 9852 4029 9856
rect 4033 9852 4034 9856
rect 4038 9852 4039 9856
rect 4043 9852 4044 9856
rect 4048 9852 4049 9856
rect 4053 9852 4054 9856
rect 4058 9852 4059 9856
rect 4063 9852 4064 9856
rect 4068 9852 4069 9856
rect 4073 9852 4074 9856
rect 4078 9852 4081 9856
rect 4085 9852 4087 9856
rect 4015 9850 4087 9852
rect 609 9766 4563 9770
rect 609 9762 802 9766
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 821 9762 831 9766
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 850 9762 860 9766
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 879 9762 889 9766
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 908 9762 918 9766
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 937 9762 1319 9766
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1338 9762 1628 9766
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1647 9762 1937 9766
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1956 9762 2246 9766
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2265 9762 2555 9766
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2574 9762 2864 9766
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2883 9762 3173 9766
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3192 9762 3482 9766
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3501 9762 3791 9766
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3810 9762 4100 9766
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4119 9762 4292 9766
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4311 9762 4318 9766
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4337 9762 4344 9766
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4363 9762 4370 9766
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4389 9762 4396 9766
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4415 9762 4563 9766
rect 609 9756 4563 9762
rect 609 9752 802 9756
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 821 9752 831 9756
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 850 9752 860 9756
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 879 9752 889 9756
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 908 9752 918 9756
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 937 9752 1319 9756
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1338 9752 1628 9756
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1647 9752 1937 9756
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1956 9752 2246 9756
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2265 9752 2555 9756
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2574 9752 2864 9756
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2883 9752 3173 9756
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3192 9752 3482 9756
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3501 9752 3791 9756
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3810 9752 4100 9756
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4119 9752 4292 9756
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4311 9752 4318 9756
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4337 9752 4344 9756
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4363 9752 4370 9756
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4389 9752 4396 9756
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4415 9752 4563 9756
rect 609 9746 4563 9752
rect 609 9742 802 9746
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 821 9742 831 9746
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 850 9742 860 9746
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 879 9742 889 9746
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 908 9742 918 9746
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 937 9742 1319 9746
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1338 9742 1628 9746
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1647 9742 1937 9746
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1956 9742 2246 9746
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2265 9742 2555 9746
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2574 9742 2864 9746
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2883 9742 3173 9746
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3192 9742 3482 9746
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3501 9742 3791 9746
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3810 9742 4100 9746
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4119 9742 4292 9746
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4311 9742 4318 9746
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4337 9742 4344 9746
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4363 9742 4370 9746
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4389 9742 4396 9746
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4415 9742 4563 9746
rect 609 9736 4563 9742
rect 609 9732 802 9736
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 821 9732 831 9736
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 850 9732 860 9736
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 879 9732 889 9736
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 908 9732 918 9736
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 937 9732 1319 9736
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1338 9732 1628 9736
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1647 9732 1937 9736
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1956 9732 2246 9736
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2265 9732 2555 9736
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2574 9732 2864 9736
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2883 9732 3173 9736
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3192 9732 3482 9736
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3501 9732 3791 9736
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3810 9732 4100 9736
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4119 9732 4292 9736
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4311 9732 4318 9736
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4337 9732 4344 9736
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4363 9732 4370 9736
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4389 9732 4396 9736
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 4415 9732 4563 9736
rect 609 9730 4563 9732
rect 609 9622 649 9730
rect 609 9618 613 9622
rect 617 9618 623 9622
rect 627 9618 633 9622
rect 637 9618 643 9622
rect 647 9618 649 9622
rect 609 9617 649 9618
rect 609 9613 613 9617
rect 617 9613 623 9617
rect 627 9613 633 9617
rect 637 9613 643 9617
rect 647 9613 649 9617
rect 609 9612 649 9613
rect 609 9608 613 9612
rect 617 9608 623 9612
rect 627 9608 633 9612
rect 637 9608 643 9612
rect 647 9608 649 9612
rect 609 9607 649 9608
rect 609 9603 613 9607
rect 617 9603 623 9607
rect 627 9603 633 9607
rect 637 9603 643 9607
rect 647 9603 649 9607
rect 609 9596 649 9603
rect 609 9592 613 9596
rect 617 9592 623 9596
rect 627 9592 633 9596
rect 637 9592 643 9596
rect 647 9592 649 9596
rect 609 9591 649 9592
rect 609 9587 613 9591
rect 617 9587 623 9591
rect 627 9587 633 9591
rect 637 9587 643 9591
rect 647 9587 649 9591
rect 609 9586 649 9587
rect 609 9582 613 9586
rect 617 9582 623 9586
rect 627 9582 633 9586
rect 637 9582 643 9586
rect 647 9582 649 9586
rect 609 9581 649 9582
rect 609 9577 613 9581
rect 617 9577 623 9581
rect 627 9577 633 9581
rect 637 9577 643 9581
rect 647 9577 649 9581
rect 609 9570 649 9577
rect 609 9566 613 9570
rect 617 9566 623 9570
rect 627 9566 633 9570
rect 637 9566 643 9570
rect 647 9566 649 9570
rect 609 9565 649 9566
rect 609 9561 613 9565
rect 617 9561 623 9565
rect 627 9561 633 9565
rect 637 9561 643 9565
rect 647 9561 649 9565
rect 609 9560 649 9561
rect 609 9556 613 9560
rect 617 9556 623 9560
rect 627 9556 633 9560
rect 637 9556 643 9560
rect 647 9556 649 9560
rect 609 9555 649 9556
rect 609 9551 613 9555
rect 617 9551 623 9555
rect 627 9551 633 9555
rect 637 9551 643 9555
rect 647 9551 649 9555
rect 609 9544 649 9551
rect 609 9540 613 9544
rect 617 9540 623 9544
rect 627 9540 633 9544
rect 637 9540 643 9544
rect 647 9540 649 9544
rect 609 9539 649 9540
rect 609 9535 613 9539
rect 617 9535 623 9539
rect 627 9535 633 9539
rect 637 9535 643 9539
rect 647 9535 649 9539
rect 609 9534 649 9535
rect 609 9530 613 9534
rect 617 9530 623 9534
rect 627 9530 633 9534
rect 637 9530 643 9534
rect 647 9530 649 9534
rect 609 9529 649 9530
rect 609 9525 613 9529
rect 617 9525 623 9529
rect 627 9525 633 9529
rect 637 9525 643 9529
rect 647 9525 649 9529
rect 609 9518 649 9525
rect 609 9514 613 9518
rect 617 9514 623 9518
rect 627 9514 633 9518
rect 637 9514 643 9518
rect 647 9514 649 9518
rect 609 9513 649 9514
rect 609 9509 613 9513
rect 617 9509 623 9513
rect 627 9509 633 9513
rect 637 9509 643 9513
rect 647 9509 649 9513
rect 609 9508 649 9509
rect 609 9504 613 9508
rect 617 9504 623 9508
rect 627 9504 633 9508
rect 637 9504 643 9508
rect 647 9504 649 9508
rect 609 9503 649 9504
rect 609 9499 613 9503
rect 617 9499 623 9503
rect 627 9499 633 9503
rect 637 9499 643 9503
rect 647 9499 649 9503
rect 609 9325 649 9499
rect 609 9321 613 9325
rect 617 9321 623 9325
rect 627 9321 633 9325
rect 637 9321 643 9325
rect 647 9321 649 9325
rect 609 9320 649 9321
rect 609 9316 613 9320
rect 617 9316 623 9320
rect 627 9316 633 9320
rect 637 9316 643 9320
rect 647 9316 649 9320
rect 609 9315 649 9316
rect 609 9311 613 9315
rect 617 9311 623 9315
rect 627 9311 633 9315
rect 637 9311 643 9315
rect 647 9311 649 9315
rect 609 9310 649 9311
rect 609 9306 613 9310
rect 617 9306 623 9310
rect 627 9306 633 9310
rect 637 9306 643 9310
rect 647 9306 649 9310
rect 609 9016 649 9306
rect 609 9012 613 9016
rect 617 9012 623 9016
rect 627 9012 633 9016
rect 637 9012 643 9016
rect 647 9012 649 9016
rect 609 9011 649 9012
rect 609 9007 613 9011
rect 617 9007 623 9011
rect 627 9007 633 9011
rect 637 9007 643 9011
rect 647 9007 649 9011
rect 609 9006 649 9007
rect 609 9002 613 9006
rect 617 9002 623 9006
rect 627 9002 633 9006
rect 637 9002 643 9006
rect 647 9002 649 9006
rect 609 9001 649 9002
rect 609 8997 613 9001
rect 617 8997 623 9001
rect 627 8997 633 9001
rect 637 8997 643 9001
rect 647 8997 649 9001
rect 609 8707 649 8997
rect 609 8703 613 8707
rect 617 8703 623 8707
rect 627 8703 633 8707
rect 637 8703 643 8707
rect 647 8703 649 8707
rect 609 8702 649 8703
rect 609 8698 613 8702
rect 617 8698 623 8702
rect 627 8698 633 8702
rect 637 8698 643 8702
rect 647 8698 649 8702
rect 609 8697 649 8698
rect 609 8693 613 8697
rect 617 8693 623 8697
rect 627 8693 633 8697
rect 637 8693 643 8697
rect 647 8693 649 8697
rect 609 8692 649 8693
rect 609 8688 613 8692
rect 617 8688 623 8692
rect 627 8688 633 8692
rect 637 8688 643 8692
rect 647 8688 649 8692
rect 609 8398 649 8688
rect 609 8394 613 8398
rect 617 8394 623 8398
rect 627 8394 633 8398
rect 637 8394 643 8398
rect 647 8394 649 8398
rect 609 8393 649 8394
rect 609 8389 613 8393
rect 617 8389 623 8393
rect 627 8389 633 8393
rect 637 8389 643 8393
rect 647 8389 649 8393
rect 609 8388 649 8389
rect 609 8384 613 8388
rect 617 8384 623 8388
rect 627 8384 633 8388
rect 637 8384 643 8388
rect 647 8384 649 8388
rect 609 8383 649 8384
rect 609 8379 613 8383
rect 617 8379 623 8383
rect 627 8379 633 8383
rect 637 8379 643 8383
rect 647 8379 649 8383
rect 609 8089 649 8379
rect 609 8085 613 8089
rect 617 8085 623 8089
rect 627 8085 633 8089
rect 637 8085 643 8089
rect 647 8085 649 8089
rect 609 8084 649 8085
rect 609 8080 613 8084
rect 617 8080 623 8084
rect 627 8080 633 8084
rect 637 8080 643 8084
rect 647 8080 649 8084
rect 609 8079 649 8080
rect 609 8075 613 8079
rect 617 8075 623 8079
rect 627 8075 633 8079
rect 637 8075 643 8079
rect 647 8075 649 8079
rect 609 8074 649 8075
rect 609 8070 613 8074
rect 617 8070 623 8074
rect 627 8070 633 8074
rect 637 8070 643 8074
rect 647 8070 649 8074
rect 609 7780 649 8070
rect 609 7776 613 7780
rect 617 7776 623 7780
rect 627 7776 633 7780
rect 637 7776 643 7780
rect 647 7776 649 7780
rect 609 7775 649 7776
rect 609 7771 613 7775
rect 617 7771 623 7775
rect 627 7771 633 7775
rect 637 7771 643 7775
rect 647 7771 649 7775
rect 609 7770 649 7771
rect 609 7766 613 7770
rect 617 7766 623 7770
rect 627 7766 633 7770
rect 637 7766 643 7770
rect 647 7766 649 7770
rect 609 7765 649 7766
rect 609 7761 613 7765
rect 617 7761 623 7765
rect 627 7761 633 7765
rect 637 7761 643 7765
rect 647 7761 649 7765
rect 609 7471 649 7761
rect 609 7467 613 7471
rect 617 7467 623 7471
rect 627 7467 633 7471
rect 637 7467 643 7471
rect 647 7467 649 7471
rect 609 7466 649 7467
rect 609 7462 613 7466
rect 617 7462 623 7466
rect 627 7462 633 7466
rect 637 7462 643 7466
rect 647 7462 649 7466
rect 609 7461 649 7462
rect 609 7457 613 7461
rect 617 7457 623 7461
rect 627 7457 633 7461
rect 637 7457 643 7461
rect 647 7457 649 7461
rect 609 7456 649 7457
rect 609 7452 613 7456
rect 617 7452 623 7456
rect 627 7452 633 7456
rect 637 7452 643 7456
rect 647 7452 649 7456
rect 609 7162 649 7452
rect 609 7158 613 7162
rect 617 7158 623 7162
rect 627 7158 633 7162
rect 637 7158 643 7162
rect 647 7158 649 7162
rect 609 7157 649 7158
rect 609 7153 613 7157
rect 617 7153 623 7157
rect 627 7153 633 7157
rect 637 7153 643 7157
rect 647 7153 649 7157
rect 609 7152 649 7153
rect 609 7148 613 7152
rect 617 7148 623 7152
rect 627 7148 633 7152
rect 637 7148 643 7152
rect 647 7148 649 7152
rect 609 7147 649 7148
rect 609 7143 613 7147
rect 617 7143 623 7147
rect 627 7143 633 7147
rect 637 7143 643 7147
rect 647 7143 649 7147
rect 609 6853 649 7143
rect 609 6849 613 6853
rect 617 6849 623 6853
rect 627 6849 633 6853
rect 637 6849 643 6853
rect 647 6849 649 6853
rect 609 6848 649 6849
rect 609 6844 613 6848
rect 617 6844 623 6848
rect 627 6844 633 6848
rect 637 6844 643 6848
rect 647 6844 649 6848
rect 609 6843 649 6844
rect 609 6839 613 6843
rect 617 6839 623 6843
rect 627 6839 633 6843
rect 637 6839 643 6843
rect 647 6839 649 6843
rect 609 6838 649 6839
rect 609 6834 613 6838
rect 617 6834 623 6838
rect 627 6834 633 6838
rect 637 6834 643 6838
rect 647 6834 649 6838
rect 609 6544 649 6834
rect 609 6540 613 6544
rect 617 6540 623 6544
rect 627 6540 633 6544
rect 637 6540 643 6544
rect 647 6540 649 6544
rect 609 6539 649 6540
rect 609 6535 613 6539
rect 617 6535 623 6539
rect 627 6535 633 6539
rect 637 6535 643 6539
rect 647 6535 649 6539
rect 609 6534 649 6535
rect 609 6530 613 6534
rect 617 6530 623 6534
rect 627 6530 633 6534
rect 637 6530 643 6534
rect 647 6530 649 6534
rect 609 6529 649 6530
rect 609 6525 613 6529
rect 617 6525 623 6529
rect 627 6525 633 6529
rect 637 6525 643 6529
rect 647 6525 649 6529
rect 609 6144 649 6525
rect 609 6140 613 6144
rect 617 6140 623 6144
rect 627 6140 633 6144
rect 637 6140 643 6144
rect 647 6140 649 6144
rect 609 6139 649 6140
rect 609 6135 613 6139
rect 617 6135 623 6139
rect 627 6135 633 6139
rect 637 6135 643 6139
rect 647 6135 649 6139
rect 609 6134 649 6135
rect 609 6130 613 6134
rect 617 6130 623 6134
rect 627 6130 633 6134
rect 637 6130 643 6134
rect 647 6130 649 6134
rect 609 6129 649 6130
rect 609 6125 613 6129
rect 617 6125 623 6129
rect 627 6125 633 6129
rect 637 6125 643 6129
rect 647 6125 649 6129
rect 609 6115 649 6125
rect 609 6111 613 6115
rect 617 6111 623 6115
rect 627 6111 633 6115
rect 637 6111 643 6115
rect 647 6111 649 6115
rect 609 6110 649 6111
rect 609 6106 613 6110
rect 617 6106 623 6110
rect 627 6106 633 6110
rect 637 6106 643 6110
rect 647 6106 649 6110
rect 609 6105 649 6106
rect 609 6101 613 6105
rect 617 6101 623 6105
rect 627 6101 633 6105
rect 637 6101 643 6105
rect 647 6101 649 6105
rect 609 6100 649 6101
rect 609 6096 613 6100
rect 617 6096 623 6100
rect 627 6096 633 6100
rect 637 6096 643 6100
rect 647 6096 649 6100
rect 609 6086 649 6096
rect 609 6082 613 6086
rect 617 6082 623 6086
rect 627 6082 633 6086
rect 637 6082 643 6086
rect 647 6082 649 6086
rect 609 6081 649 6082
rect 609 6077 613 6081
rect 617 6077 623 6081
rect 627 6077 633 6081
rect 637 6077 643 6081
rect 647 6077 649 6081
rect 609 6076 649 6077
rect 609 6072 613 6076
rect 617 6072 623 6076
rect 627 6072 633 6076
rect 637 6072 643 6076
rect 647 6072 649 6076
rect 609 6071 649 6072
rect 609 6067 613 6071
rect 617 6067 623 6071
rect 627 6067 633 6071
rect 637 6067 643 6071
rect 647 6067 649 6071
rect 609 6057 649 6067
rect 609 6053 613 6057
rect 617 6053 623 6057
rect 627 6053 633 6057
rect 637 6053 643 6057
rect 647 6053 649 6057
rect 609 6052 649 6053
rect 609 6048 613 6052
rect 617 6048 623 6052
rect 627 6048 633 6052
rect 637 6048 643 6052
rect 647 6048 649 6052
rect 609 6047 649 6048
rect 609 6043 613 6047
rect 617 6043 623 6047
rect 627 6043 633 6047
rect 637 6043 643 6047
rect 647 6043 649 6047
rect 609 6042 649 6043
rect 609 6038 613 6042
rect 617 6038 623 6042
rect 627 6038 633 6042
rect 637 6038 643 6042
rect 647 6038 649 6042
rect 609 6028 649 6038
rect 609 6024 613 6028
rect 617 6024 623 6028
rect 627 6024 633 6028
rect 637 6024 643 6028
rect 647 6024 649 6028
rect 609 6023 649 6024
rect 609 6019 613 6023
rect 617 6019 623 6023
rect 627 6019 633 6023
rect 637 6019 643 6023
rect 647 6019 649 6023
rect 609 6018 649 6019
rect 609 6014 613 6018
rect 617 6014 623 6018
rect 627 6014 633 6018
rect 637 6014 643 6018
rect 647 6014 649 6018
rect 609 6013 649 6014
rect 609 6009 613 6013
rect 617 6009 623 6013
rect 627 6009 633 6013
rect 637 6009 643 6013
rect 647 6009 649 6013
rect 609 5856 649 6009
rect 4523 9577 4563 9730
rect 4523 9573 4525 9577
rect 4529 9573 4535 9577
rect 4539 9573 4545 9577
rect 4549 9573 4555 9577
rect 4559 9573 4563 9577
rect 4523 9572 4563 9573
rect 4523 9568 4525 9572
rect 4529 9568 4535 9572
rect 4539 9568 4545 9572
rect 4549 9568 4555 9572
rect 4559 9568 4563 9572
rect 4523 9567 4563 9568
rect 4523 9563 4525 9567
rect 4529 9563 4535 9567
rect 4539 9563 4545 9567
rect 4549 9563 4555 9567
rect 4559 9563 4563 9567
rect 4523 9562 4563 9563
rect 4523 9558 4525 9562
rect 4529 9558 4535 9562
rect 4539 9558 4545 9562
rect 4549 9558 4555 9562
rect 4559 9558 4563 9562
rect 4523 9548 4563 9558
rect 4523 9544 4525 9548
rect 4529 9544 4535 9548
rect 4539 9544 4545 9548
rect 4549 9544 4555 9548
rect 4559 9544 4563 9548
rect 4523 9543 4563 9544
rect 4523 9539 4525 9543
rect 4529 9539 4535 9543
rect 4539 9539 4545 9543
rect 4549 9539 4555 9543
rect 4559 9539 4563 9543
rect 4523 9538 4563 9539
rect 4523 9534 4525 9538
rect 4529 9534 4535 9538
rect 4539 9534 4545 9538
rect 4549 9534 4555 9538
rect 4559 9534 4563 9538
rect 4523 9533 4563 9534
rect 4523 9529 4525 9533
rect 4529 9529 4535 9533
rect 4539 9529 4545 9533
rect 4549 9529 4555 9533
rect 4559 9529 4563 9533
rect 4523 9519 4563 9529
rect 4523 9515 4525 9519
rect 4529 9515 4535 9519
rect 4539 9515 4545 9519
rect 4549 9515 4555 9519
rect 4559 9515 4563 9519
rect 4523 9514 4563 9515
rect 4523 9510 4525 9514
rect 4529 9510 4535 9514
rect 4539 9510 4545 9514
rect 4549 9510 4555 9514
rect 4559 9510 4563 9514
rect 4523 9509 4563 9510
rect 4523 9505 4525 9509
rect 4529 9505 4535 9509
rect 4539 9505 4545 9509
rect 4549 9505 4555 9509
rect 4559 9505 4563 9509
rect 4523 9504 4563 9505
rect 4523 9500 4525 9504
rect 4529 9500 4535 9504
rect 4539 9500 4545 9504
rect 4549 9500 4555 9504
rect 4559 9500 4563 9504
rect 4523 9490 4563 9500
rect 4523 9486 4525 9490
rect 4529 9486 4535 9490
rect 4539 9486 4545 9490
rect 4549 9486 4555 9490
rect 4559 9486 4563 9490
rect 4523 9485 4563 9486
rect 4523 9481 4525 9485
rect 4529 9481 4535 9485
rect 4539 9481 4545 9485
rect 4549 9481 4555 9485
rect 4559 9481 4563 9485
rect 4523 9480 4563 9481
rect 4523 9476 4525 9480
rect 4529 9476 4535 9480
rect 4539 9476 4545 9480
rect 4549 9476 4555 9480
rect 4559 9476 4563 9480
rect 4523 9475 4563 9476
rect 4523 9471 4525 9475
rect 4529 9471 4535 9475
rect 4539 9471 4545 9475
rect 4549 9471 4555 9475
rect 4559 9471 4563 9475
rect 4523 9461 4563 9471
rect 4523 9457 4525 9461
rect 4529 9457 4535 9461
rect 4539 9457 4545 9461
rect 4549 9457 4555 9461
rect 4559 9457 4563 9461
rect 4523 9456 4563 9457
rect 4523 9452 4525 9456
rect 4529 9452 4535 9456
rect 4539 9452 4545 9456
rect 4549 9452 4555 9456
rect 4559 9452 4563 9456
rect 4523 9451 4563 9452
rect 4523 9447 4525 9451
rect 4529 9447 4535 9451
rect 4539 9447 4545 9451
rect 4549 9447 4555 9451
rect 4559 9447 4563 9451
rect 4523 9446 4563 9447
rect 4523 9442 4525 9446
rect 4529 9442 4535 9446
rect 4539 9442 4545 9446
rect 4549 9442 4555 9446
rect 4559 9442 4563 9446
rect 4523 9060 4563 9442
rect 4523 9056 4525 9060
rect 4529 9056 4535 9060
rect 4539 9056 4545 9060
rect 4549 9056 4555 9060
rect 4559 9056 4563 9060
rect 4523 9055 4563 9056
rect 4523 9051 4525 9055
rect 4529 9051 4535 9055
rect 4539 9051 4545 9055
rect 4549 9051 4555 9055
rect 4559 9051 4563 9055
rect 4523 9050 4563 9051
rect 4523 9046 4525 9050
rect 4529 9046 4535 9050
rect 4539 9046 4545 9050
rect 4549 9046 4555 9050
rect 4559 9046 4563 9050
rect 4523 9045 4563 9046
rect 4523 9041 4525 9045
rect 4529 9041 4535 9045
rect 4539 9041 4545 9045
rect 4549 9041 4555 9045
rect 4559 9041 4563 9045
rect 4523 8751 4563 9041
rect 4523 8747 4525 8751
rect 4529 8747 4535 8751
rect 4539 8747 4545 8751
rect 4549 8747 4555 8751
rect 4559 8747 4563 8751
rect 4523 8746 4563 8747
rect 4523 8742 4525 8746
rect 4529 8742 4535 8746
rect 4539 8742 4545 8746
rect 4549 8742 4555 8746
rect 4559 8742 4563 8746
rect 4523 8741 4563 8742
rect 4523 8737 4525 8741
rect 4529 8737 4535 8741
rect 4539 8737 4545 8741
rect 4549 8737 4555 8741
rect 4559 8737 4563 8741
rect 4523 8736 4563 8737
rect 4523 8732 4525 8736
rect 4529 8732 4535 8736
rect 4539 8732 4545 8736
rect 4549 8732 4555 8736
rect 4559 8732 4563 8736
rect 4523 8442 4563 8732
rect 4523 8438 4525 8442
rect 4529 8438 4535 8442
rect 4539 8438 4545 8442
rect 4549 8438 4555 8442
rect 4559 8438 4563 8442
rect 4523 8437 4563 8438
rect 4523 8433 4525 8437
rect 4529 8433 4535 8437
rect 4539 8433 4545 8437
rect 4549 8433 4555 8437
rect 4559 8433 4563 8437
rect 4523 8432 4563 8433
rect 4523 8428 4525 8432
rect 4529 8428 4535 8432
rect 4539 8428 4545 8432
rect 4549 8428 4555 8432
rect 4559 8428 4563 8432
rect 4523 8427 4563 8428
rect 4523 8423 4525 8427
rect 4529 8423 4535 8427
rect 4539 8423 4545 8427
rect 4549 8423 4555 8427
rect 4559 8423 4563 8427
rect 4523 8133 4563 8423
rect 4523 8129 4525 8133
rect 4529 8129 4535 8133
rect 4539 8129 4545 8133
rect 4549 8129 4555 8133
rect 4559 8129 4563 8133
rect 4523 8128 4563 8129
rect 4523 8124 4525 8128
rect 4529 8124 4535 8128
rect 4539 8124 4545 8128
rect 4549 8124 4555 8128
rect 4559 8124 4563 8128
rect 4523 8123 4563 8124
rect 4523 8119 4525 8123
rect 4529 8119 4535 8123
rect 4539 8119 4545 8123
rect 4549 8119 4555 8123
rect 4559 8119 4563 8123
rect 4523 8118 4563 8119
rect 4523 8114 4525 8118
rect 4529 8114 4535 8118
rect 4539 8114 4545 8118
rect 4549 8114 4555 8118
rect 4559 8114 4563 8118
rect 4523 8102 4563 8114
rect 4523 8098 4525 8102
rect 4529 8098 4535 8102
rect 4539 8098 4545 8102
rect 4549 8098 4555 8102
rect 4559 8098 4563 8102
rect 4523 8097 4563 8098
rect 4523 8093 4525 8097
rect 4529 8093 4535 8097
rect 4539 8093 4545 8097
rect 4549 8093 4555 8097
rect 4559 8093 4563 8097
rect 4523 8092 4563 8093
rect 4523 8088 4525 8092
rect 4529 8088 4535 8092
rect 4539 8088 4545 8092
rect 4549 8088 4555 8092
rect 4559 8088 4563 8092
rect 4523 8087 4563 8088
rect 4523 8083 4525 8087
rect 4529 8083 4535 8087
rect 4539 8083 4545 8087
rect 4549 8083 4555 8087
rect 4559 8083 4563 8087
rect 4523 7793 4563 8083
rect 4523 7789 4525 7793
rect 4529 7789 4535 7793
rect 4539 7789 4545 7793
rect 4549 7789 4555 7793
rect 4559 7789 4563 7793
rect 4523 7788 4563 7789
rect 4523 7784 4525 7788
rect 4529 7784 4535 7788
rect 4539 7784 4545 7788
rect 4549 7784 4555 7788
rect 4559 7784 4563 7788
rect 4523 7783 4563 7784
rect 4523 7779 4525 7783
rect 4529 7779 4535 7783
rect 4539 7779 4545 7783
rect 4549 7779 4555 7783
rect 4559 7779 4563 7783
rect 4523 7778 4563 7779
rect 4523 7774 4525 7778
rect 4529 7774 4535 7778
rect 4539 7774 4545 7778
rect 4549 7774 4555 7778
rect 4559 7774 4563 7778
rect 4523 7206 4563 7774
rect 4523 7202 4525 7206
rect 4529 7202 4535 7206
rect 4539 7202 4545 7206
rect 4549 7202 4555 7206
rect 4559 7202 4563 7206
rect 4523 7201 4563 7202
rect 4523 7197 4525 7201
rect 4529 7197 4535 7201
rect 4539 7197 4545 7201
rect 4549 7197 4555 7201
rect 4559 7197 4563 7201
rect 4523 7196 4563 7197
rect 4523 7192 4525 7196
rect 4529 7192 4535 7196
rect 4539 7192 4545 7196
rect 4549 7192 4555 7196
rect 4559 7192 4563 7196
rect 4523 7191 4563 7192
rect 4523 7187 4525 7191
rect 4529 7187 4535 7191
rect 4539 7187 4545 7191
rect 4549 7187 4555 7191
rect 4559 7187 4563 7191
rect 4523 6897 4563 7187
rect 4523 6893 4525 6897
rect 4529 6893 4535 6897
rect 4539 6893 4545 6897
rect 4549 6893 4555 6897
rect 4559 6893 4563 6897
rect 4523 6892 4563 6893
rect 4523 6888 4525 6892
rect 4529 6888 4535 6892
rect 4539 6888 4545 6892
rect 4549 6888 4555 6892
rect 4559 6888 4563 6892
rect 4523 6887 4563 6888
rect 4523 6883 4525 6887
rect 4529 6883 4535 6887
rect 4539 6883 4545 6887
rect 4549 6883 4555 6887
rect 4559 6883 4563 6887
rect 4523 6882 4563 6883
rect 4523 6878 4525 6882
rect 4529 6878 4535 6882
rect 4539 6878 4545 6882
rect 4549 6878 4555 6882
rect 4559 6878 4563 6882
rect 4523 6588 4563 6878
rect 4523 6584 4525 6588
rect 4529 6584 4535 6588
rect 4539 6584 4545 6588
rect 4549 6584 4555 6588
rect 4559 6584 4563 6588
rect 4523 6583 4563 6584
rect 4523 6579 4525 6583
rect 4529 6579 4535 6583
rect 4539 6579 4545 6583
rect 4549 6579 4555 6583
rect 4559 6579 4563 6583
rect 4523 6578 4563 6579
rect 4523 6574 4525 6578
rect 4529 6574 4535 6578
rect 4539 6574 4545 6578
rect 4549 6574 4555 6578
rect 4559 6574 4563 6578
rect 4523 6573 4563 6574
rect 4523 6569 4525 6573
rect 4529 6569 4535 6573
rect 4539 6569 4545 6573
rect 4549 6569 4555 6573
rect 4559 6569 4563 6573
rect 4523 6279 4563 6569
rect 4523 6275 4525 6279
rect 4529 6275 4535 6279
rect 4539 6275 4545 6279
rect 4549 6275 4555 6279
rect 4559 6275 4563 6279
rect 4523 6274 4563 6275
rect 4523 6270 4525 6274
rect 4529 6270 4535 6274
rect 4539 6270 4545 6274
rect 4549 6270 4555 6274
rect 4559 6270 4563 6274
rect 4523 6269 4563 6270
rect 4523 6265 4525 6269
rect 4529 6265 4535 6269
rect 4539 6265 4545 6269
rect 4549 6265 4555 6269
rect 4559 6265 4563 6269
rect 4523 6264 4563 6265
rect 4523 6260 4525 6264
rect 4529 6260 4535 6264
rect 4539 6260 4545 6264
rect 4549 6260 4555 6264
rect 4559 6260 4563 6264
rect 4523 6087 4563 6260
rect 4523 6083 4525 6087
rect 4529 6083 4535 6087
rect 4539 6083 4545 6087
rect 4549 6083 4555 6087
rect 4559 6083 4563 6087
rect 4523 6082 4563 6083
rect 4523 6078 4525 6082
rect 4529 6078 4535 6082
rect 4539 6078 4545 6082
rect 4549 6078 4555 6082
rect 4559 6078 4563 6082
rect 4523 6077 4563 6078
rect 4523 6073 4525 6077
rect 4529 6073 4535 6077
rect 4539 6073 4545 6077
rect 4549 6073 4555 6077
rect 4559 6073 4563 6077
rect 4523 6072 4563 6073
rect 4523 6068 4525 6072
rect 4529 6068 4535 6072
rect 4539 6068 4545 6072
rect 4549 6068 4555 6072
rect 4559 6068 4563 6072
rect 4523 6061 4563 6068
rect 4523 6057 4525 6061
rect 4529 6057 4535 6061
rect 4539 6057 4545 6061
rect 4549 6057 4555 6061
rect 4559 6057 4563 6061
rect 4523 6056 4563 6057
rect 4523 6052 4525 6056
rect 4529 6052 4535 6056
rect 4539 6052 4545 6056
rect 4549 6052 4555 6056
rect 4559 6052 4563 6056
rect 4523 6051 4563 6052
rect 4523 6047 4525 6051
rect 4529 6047 4535 6051
rect 4539 6047 4545 6051
rect 4549 6047 4555 6051
rect 4559 6047 4563 6051
rect 4523 6046 4563 6047
rect 4523 6042 4525 6046
rect 4529 6042 4535 6046
rect 4539 6042 4545 6046
rect 4549 6042 4555 6046
rect 4559 6042 4563 6046
rect 4523 6035 4563 6042
rect 4523 6031 4525 6035
rect 4529 6031 4535 6035
rect 4539 6031 4545 6035
rect 4549 6031 4555 6035
rect 4559 6031 4563 6035
rect 4523 6030 4563 6031
rect 4523 6026 4525 6030
rect 4529 6026 4535 6030
rect 4539 6026 4545 6030
rect 4549 6026 4555 6030
rect 4559 6026 4563 6030
rect 4523 6025 4563 6026
rect 4523 6021 4525 6025
rect 4529 6021 4535 6025
rect 4539 6021 4545 6025
rect 4549 6021 4555 6025
rect 4559 6021 4563 6025
rect 4523 6020 4563 6021
rect 4523 6016 4525 6020
rect 4529 6016 4535 6020
rect 4539 6016 4545 6020
rect 4549 6016 4555 6020
rect 4559 6016 4563 6020
rect 4523 6009 4563 6016
rect 4523 6005 4525 6009
rect 4529 6005 4535 6009
rect 4539 6005 4545 6009
rect 4549 6005 4555 6009
rect 4559 6005 4563 6009
rect 4523 6004 4563 6005
rect 4523 6000 4525 6004
rect 4529 6000 4535 6004
rect 4539 6000 4545 6004
rect 4549 6000 4555 6004
rect 4559 6000 4563 6004
rect 4523 5999 4563 6000
rect 4523 5995 4525 5999
rect 4529 5995 4535 5999
rect 4539 5995 4545 5999
rect 4549 5995 4555 5999
rect 4559 5995 4563 5999
rect 4523 5994 4563 5995
rect 4523 5990 4525 5994
rect 4529 5990 4535 5994
rect 4539 5990 4545 5994
rect 4549 5990 4555 5994
rect 4559 5990 4563 5994
rect 4523 5983 4563 5990
rect 4523 5979 4525 5983
rect 4529 5979 4535 5983
rect 4539 5979 4545 5983
rect 4549 5979 4555 5983
rect 4559 5979 4563 5983
rect 4523 5978 4563 5979
rect 4523 5974 4525 5978
rect 4529 5974 4535 5978
rect 4539 5974 4545 5978
rect 4549 5974 4555 5978
rect 4559 5974 4563 5978
rect 4523 5973 4563 5974
rect 4523 5969 4525 5973
rect 4529 5969 4535 5973
rect 4539 5969 4545 5973
rect 4549 5969 4555 5973
rect 4559 5969 4563 5973
rect 4523 5968 4563 5969
rect 4523 5964 4525 5968
rect 4529 5964 4535 5968
rect 4539 5964 4545 5968
rect 4549 5964 4555 5968
rect 4559 5964 4563 5968
rect 4523 5856 4563 5964
rect 609 5854 4563 5856
rect 609 5850 757 5854
rect 761 5850 762 5854
rect 766 5850 767 5854
rect 771 5850 772 5854
rect 776 5850 783 5854
rect 787 5850 788 5854
rect 792 5850 793 5854
rect 797 5850 798 5854
rect 802 5850 809 5854
rect 813 5850 814 5854
rect 818 5850 819 5854
rect 823 5850 824 5854
rect 828 5850 835 5854
rect 839 5850 840 5854
rect 844 5850 845 5854
rect 849 5850 850 5854
rect 854 5850 861 5854
rect 865 5850 866 5854
rect 870 5850 871 5854
rect 875 5850 876 5854
rect 880 5850 1054 5854
rect 1058 5850 1059 5854
rect 1063 5850 1064 5854
rect 1068 5850 1069 5854
rect 1073 5850 1363 5854
rect 1367 5850 1368 5854
rect 1372 5850 1373 5854
rect 1377 5850 1378 5854
rect 1382 5850 1672 5854
rect 1676 5850 1677 5854
rect 1681 5850 1682 5854
rect 1686 5850 1687 5854
rect 1691 5850 1981 5854
rect 1985 5850 1986 5854
rect 1990 5850 1991 5854
rect 1995 5850 1996 5854
rect 2000 5850 2290 5854
rect 2294 5850 2295 5854
rect 2299 5850 2300 5854
rect 2304 5850 2305 5854
rect 2309 5850 2599 5854
rect 2603 5850 2604 5854
rect 2608 5850 2609 5854
rect 2613 5850 2614 5854
rect 2618 5850 2908 5854
rect 2912 5850 2913 5854
rect 2917 5850 2918 5854
rect 2922 5850 2923 5854
rect 2927 5850 3217 5854
rect 3221 5850 3222 5854
rect 3226 5850 3227 5854
rect 3231 5850 3232 5854
rect 3236 5850 3526 5854
rect 3530 5850 3531 5854
rect 3535 5850 3536 5854
rect 3540 5850 3541 5854
rect 3545 5850 3835 5854
rect 3839 5850 3840 5854
rect 3844 5850 3845 5854
rect 3849 5850 3850 5854
rect 3854 5850 4235 5854
rect 4239 5850 4240 5854
rect 4244 5850 4245 5854
rect 4249 5850 4250 5854
rect 4254 5850 4264 5854
rect 4268 5850 4269 5854
rect 4273 5850 4274 5854
rect 4278 5850 4279 5854
rect 4283 5850 4293 5854
rect 4297 5850 4298 5854
rect 4302 5850 4303 5854
rect 4307 5850 4308 5854
rect 4312 5850 4322 5854
rect 4326 5850 4327 5854
rect 4331 5850 4332 5854
rect 4336 5850 4337 5854
rect 4341 5850 4351 5854
rect 4355 5850 4356 5854
rect 4360 5850 4361 5854
rect 4365 5850 4366 5854
rect 4370 5850 4563 5854
rect 609 5844 4563 5850
rect 609 5840 757 5844
rect 761 5840 762 5844
rect 766 5840 767 5844
rect 771 5840 772 5844
rect 776 5840 783 5844
rect 787 5840 788 5844
rect 792 5840 793 5844
rect 797 5840 798 5844
rect 802 5840 809 5844
rect 813 5840 814 5844
rect 818 5840 819 5844
rect 823 5840 824 5844
rect 828 5840 835 5844
rect 839 5840 840 5844
rect 844 5840 845 5844
rect 849 5840 850 5844
rect 854 5840 861 5844
rect 865 5840 866 5844
rect 870 5840 871 5844
rect 875 5840 876 5844
rect 880 5840 1054 5844
rect 1058 5840 1059 5844
rect 1063 5840 1064 5844
rect 1068 5840 1069 5844
rect 1073 5840 1363 5844
rect 1367 5840 1368 5844
rect 1372 5840 1373 5844
rect 1377 5840 1378 5844
rect 1382 5840 1672 5844
rect 1676 5840 1677 5844
rect 1681 5840 1682 5844
rect 1686 5840 1687 5844
rect 1691 5840 1981 5844
rect 1985 5840 1986 5844
rect 1990 5840 1991 5844
rect 1995 5840 1996 5844
rect 2000 5840 2290 5844
rect 2294 5840 2295 5844
rect 2299 5840 2300 5844
rect 2304 5840 2305 5844
rect 2309 5840 2599 5844
rect 2603 5840 2604 5844
rect 2608 5840 2609 5844
rect 2613 5840 2614 5844
rect 2618 5840 2908 5844
rect 2912 5840 2913 5844
rect 2917 5840 2918 5844
rect 2922 5840 2923 5844
rect 2927 5840 3217 5844
rect 3221 5840 3222 5844
rect 3226 5840 3227 5844
rect 3231 5840 3232 5844
rect 3236 5840 3526 5844
rect 3530 5840 3531 5844
rect 3535 5840 3536 5844
rect 3540 5840 3541 5844
rect 3545 5840 3835 5844
rect 3839 5840 3840 5844
rect 3844 5840 3845 5844
rect 3849 5840 3850 5844
rect 3854 5840 4235 5844
rect 4239 5840 4240 5844
rect 4244 5840 4245 5844
rect 4249 5840 4250 5844
rect 4254 5840 4264 5844
rect 4268 5840 4269 5844
rect 4273 5840 4274 5844
rect 4278 5840 4279 5844
rect 4283 5840 4293 5844
rect 4297 5840 4298 5844
rect 4302 5840 4303 5844
rect 4307 5840 4308 5844
rect 4312 5840 4322 5844
rect 4326 5840 4327 5844
rect 4331 5840 4332 5844
rect 4336 5840 4337 5844
rect 4341 5840 4351 5844
rect 4355 5840 4356 5844
rect 4360 5840 4361 5844
rect 4365 5840 4366 5844
rect 4370 5840 4563 5844
rect 609 5834 4563 5840
rect 609 5830 757 5834
rect 761 5830 762 5834
rect 766 5830 767 5834
rect 771 5830 772 5834
rect 776 5830 783 5834
rect 787 5830 788 5834
rect 792 5830 793 5834
rect 797 5830 798 5834
rect 802 5830 809 5834
rect 813 5830 814 5834
rect 818 5830 819 5834
rect 823 5830 824 5834
rect 828 5830 835 5834
rect 839 5830 840 5834
rect 844 5830 845 5834
rect 849 5830 850 5834
rect 854 5830 861 5834
rect 865 5830 866 5834
rect 870 5830 871 5834
rect 875 5830 876 5834
rect 880 5830 1054 5834
rect 1058 5830 1059 5834
rect 1063 5830 1064 5834
rect 1068 5830 1069 5834
rect 1073 5830 1363 5834
rect 1367 5830 1368 5834
rect 1372 5830 1373 5834
rect 1377 5830 1378 5834
rect 1382 5830 1672 5834
rect 1676 5830 1677 5834
rect 1681 5830 1682 5834
rect 1686 5830 1687 5834
rect 1691 5830 1981 5834
rect 1985 5830 1986 5834
rect 1990 5830 1991 5834
rect 1995 5830 1996 5834
rect 2000 5830 2290 5834
rect 2294 5830 2295 5834
rect 2299 5830 2300 5834
rect 2304 5830 2305 5834
rect 2309 5830 2599 5834
rect 2603 5830 2604 5834
rect 2608 5830 2609 5834
rect 2613 5830 2614 5834
rect 2618 5830 2908 5834
rect 2912 5830 2913 5834
rect 2917 5830 2918 5834
rect 2922 5830 2923 5834
rect 2927 5830 3217 5834
rect 3221 5830 3222 5834
rect 3226 5830 3227 5834
rect 3231 5830 3232 5834
rect 3236 5830 3526 5834
rect 3530 5830 3531 5834
rect 3535 5830 3536 5834
rect 3540 5830 3541 5834
rect 3545 5830 3835 5834
rect 3839 5830 3840 5834
rect 3844 5830 3845 5834
rect 3849 5830 3850 5834
rect 3854 5830 4235 5834
rect 4239 5830 4240 5834
rect 4244 5830 4245 5834
rect 4249 5830 4250 5834
rect 4254 5830 4264 5834
rect 4268 5830 4269 5834
rect 4273 5830 4274 5834
rect 4278 5830 4279 5834
rect 4283 5830 4293 5834
rect 4297 5830 4298 5834
rect 4302 5830 4303 5834
rect 4307 5830 4308 5834
rect 4312 5830 4322 5834
rect 4326 5830 4327 5834
rect 4331 5830 4332 5834
rect 4336 5830 4337 5834
rect 4341 5830 4351 5834
rect 4355 5830 4356 5834
rect 4360 5830 4361 5834
rect 4365 5830 4366 5834
rect 4370 5830 4563 5834
rect 609 5824 4563 5830
rect 609 5820 757 5824
rect 761 5820 762 5824
rect 766 5820 767 5824
rect 771 5820 772 5824
rect 776 5820 783 5824
rect 787 5820 788 5824
rect 792 5820 793 5824
rect 797 5820 798 5824
rect 802 5820 809 5824
rect 813 5820 814 5824
rect 818 5820 819 5824
rect 823 5820 824 5824
rect 828 5820 835 5824
rect 839 5820 840 5824
rect 844 5820 845 5824
rect 849 5820 850 5824
rect 854 5820 861 5824
rect 865 5820 866 5824
rect 870 5820 871 5824
rect 875 5820 876 5824
rect 880 5820 1054 5824
rect 1058 5820 1059 5824
rect 1063 5820 1064 5824
rect 1068 5820 1069 5824
rect 1073 5820 1363 5824
rect 1367 5820 1368 5824
rect 1372 5820 1373 5824
rect 1377 5820 1378 5824
rect 1382 5820 1672 5824
rect 1676 5820 1677 5824
rect 1681 5820 1682 5824
rect 1686 5820 1687 5824
rect 1691 5820 1981 5824
rect 1985 5820 1986 5824
rect 1990 5820 1991 5824
rect 1995 5820 1996 5824
rect 2000 5820 2290 5824
rect 2294 5820 2295 5824
rect 2299 5820 2300 5824
rect 2304 5820 2305 5824
rect 2309 5820 2599 5824
rect 2603 5820 2604 5824
rect 2608 5820 2609 5824
rect 2613 5820 2614 5824
rect 2618 5820 2908 5824
rect 2912 5820 2913 5824
rect 2917 5820 2918 5824
rect 2922 5820 2923 5824
rect 2927 5820 3217 5824
rect 3221 5820 3222 5824
rect 3226 5820 3227 5824
rect 3231 5820 3232 5824
rect 3236 5820 3526 5824
rect 3530 5820 3531 5824
rect 3535 5820 3536 5824
rect 3540 5820 3541 5824
rect 3545 5820 3835 5824
rect 3839 5820 3840 5824
rect 3844 5820 3845 5824
rect 3849 5820 3850 5824
rect 3854 5820 4235 5824
rect 4239 5820 4240 5824
rect 4244 5820 4245 5824
rect 4249 5820 4250 5824
rect 4254 5820 4264 5824
rect 4268 5820 4269 5824
rect 4273 5820 4274 5824
rect 4278 5820 4279 5824
rect 4283 5820 4293 5824
rect 4297 5820 4298 5824
rect 4302 5820 4303 5824
rect 4307 5820 4308 5824
rect 4312 5820 4322 5824
rect 4326 5820 4327 5824
rect 4331 5820 4332 5824
rect 4336 5820 4337 5824
rect 4341 5820 4351 5824
rect 4355 5820 4356 5824
rect 4360 5820 4361 5824
rect 4365 5820 4366 5824
rect 4370 5820 4563 5824
rect 609 5816 4563 5820
<< psubstratepcontact >>
rect 1385 9961 1389 9965
rect 1392 9961 1396 9965
rect 1397 9961 1401 9965
rect 1402 9961 1406 9965
rect 1407 9961 1411 9965
rect 1412 9961 1416 9965
rect 1417 9961 1421 9965
rect 1422 9961 1426 9965
rect 1427 9961 1431 9965
rect 1432 9961 1436 9965
rect 1437 9961 1441 9965
rect 1442 9961 1446 9965
rect 1449 9961 1453 9965
rect 1385 9954 1389 9958
rect 1449 9954 1453 9958
rect 1385 9949 1389 9953
rect 1385 9944 1389 9948
rect 1385 9939 1389 9943
rect 1385 9934 1389 9938
rect 1385 9929 1389 9933
rect 1385 9924 1389 9928
rect 1385 9919 1389 9923
rect 1385 9914 1389 9918
rect 1385 9909 1389 9913
rect 1385 9904 1389 9908
rect 1385 9899 1389 9903
rect 1385 9894 1389 9898
rect 1385 9889 1389 9893
rect 1385 9884 1389 9888
rect 1385 9879 1389 9883
rect 1385 9874 1389 9878
rect 1385 9869 1389 9873
rect 1385 9864 1389 9868
rect 1449 9949 1453 9953
rect 1449 9944 1453 9948
rect 1449 9939 1453 9943
rect 1449 9934 1453 9938
rect 1449 9929 1453 9933
rect 1449 9924 1453 9928
rect 1449 9919 1453 9923
rect 1449 9914 1453 9918
rect 1449 9909 1453 9913
rect 1449 9904 1453 9908
rect 1449 9899 1453 9903
rect 1449 9894 1453 9898
rect 1449 9889 1453 9893
rect 1449 9884 1453 9888
rect 1449 9879 1453 9883
rect 1449 9874 1453 9878
rect 1449 9869 1453 9873
rect 1449 9864 1453 9868
rect 1385 9859 1389 9863
rect 1449 9859 1453 9863
rect 1385 9852 1389 9856
rect 1392 9852 1396 9856
rect 1397 9852 1401 9856
rect 1402 9852 1406 9856
rect 1407 9852 1411 9856
rect 1412 9852 1416 9856
rect 1417 9852 1421 9856
rect 1422 9852 1426 9856
rect 1427 9852 1431 9856
rect 1432 9852 1436 9856
rect 1437 9852 1441 9856
rect 1442 9852 1446 9856
rect 1449 9852 1453 9856
rect 1532 9974 1536 9978
rect 1537 9974 1541 9978
rect 1542 9974 1546 9978
rect 1547 9974 1551 9978
rect 1552 9974 1556 9978
rect 1557 9974 1561 9978
rect 1562 9974 1566 9978
rect 1567 9974 1571 9978
rect 1572 9974 1576 9978
rect 1577 9974 1581 9978
rect 1582 9974 1586 9978
rect 1587 9974 1591 9978
rect 1592 9974 1596 9978
rect 1597 9974 1601 9978
rect 1602 9974 1606 9978
rect 1607 9974 1611 9978
rect 1612 9974 1616 9978
rect 1617 9974 1621 9978
rect 1622 9974 1626 9978
rect 1532 9969 1536 9973
rect 1532 9964 1536 9968
rect 1622 9969 1626 9973
rect 1532 9959 1536 9963
rect 1532 9954 1536 9958
rect 1532 9949 1536 9953
rect 1532 9944 1536 9948
rect 1532 9939 1536 9943
rect 1532 9934 1536 9938
rect 1532 9929 1536 9933
rect 1532 9924 1536 9928
rect 1532 9919 1536 9923
rect 1532 9914 1536 9918
rect 1532 9909 1536 9913
rect 1532 9904 1536 9908
rect 1532 9899 1536 9903
rect 1532 9894 1536 9898
rect 1532 9889 1536 9893
rect 1532 9884 1536 9888
rect 1532 9879 1536 9883
rect 1532 9874 1536 9878
rect 1532 9869 1536 9873
rect 1532 9864 1536 9868
rect 1532 9859 1536 9863
rect 1532 9854 1536 9858
rect 1532 9849 1536 9853
rect 1622 9964 1626 9968
rect 1622 9959 1626 9963
rect 1622 9954 1626 9958
rect 1622 9949 1626 9953
rect 1622 9944 1626 9948
rect 1622 9939 1626 9943
rect 1622 9934 1626 9938
rect 1622 9929 1626 9933
rect 1622 9924 1626 9928
rect 1622 9919 1626 9923
rect 1622 9914 1626 9918
rect 1622 9909 1626 9913
rect 1622 9904 1626 9908
rect 1622 9899 1626 9903
rect 1622 9894 1626 9898
rect 1622 9889 1626 9893
rect 1622 9884 1626 9888
rect 1622 9879 1626 9883
rect 1622 9874 1626 9878
rect 1622 9869 1626 9873
rect 1622 9864 1626 9868
rect 1622 9859 1626 9863
rect 1622 9854 1626 9858
rect 1532 9844 1536 9848
rect 1622 9849 1626 9853
rect 1622 9844 1626 9848
rect 1532 9839 1536 9843
rect 1537 9839 1541 9843
rect 1542 9839 1546 9843
rect 1547 9839 1551 9843
rect 1552 9839 1556 9843
rect 1557 9839 1561 9843
rect 1562 9839 1566 9843
rect 1567 9839 1571 9843
rect 1572 9839 1576 9843
rect 1577 9839 1581 9843
rect 1582 9839 1586 9843
rect 1587 9839 1591 9843
rect 1592 9839 1596 9843
rect 1597 9839 1601 9843
rect 1602 9839 1606 9843
rect 1607 9839 1611 9843
rect 1612 9839 1616 9843
rect 1617 9839 1621 9843
rect 1622 9839 1626 9843
rect 1694 9961 1698 9965
rect 1701 9961 1705 9965
rect 1706 9961 1710 9965
rect 1711 9961 1715 9965
rect 1716 9961 1720 9965
rect 1721 9961 1725 9965
rect 1726 9961 1730 9965
rect 1731 9961 1735 9965
rect 1736 9961 1740 9965
rect 1741 9961 1745 9965
rect 1746 9961 1750 9965
rect 1751 9961 1755 9965
rect 1758 9961 1762 9965
rect 1694 9954 1698 9958
rect 1758 9954 1762 9958
rect 1694 9949 1698 9953
rect 1694 9944 1698 9948
rect 1694 9939 1698 9943
rect 1694 9934 1698 9938
rect 1694 9929 1698 9933
rect 1694 9924 1698 9928
rect 1694 9919 1698 9923
rect 1694 9914 1698 9918
rect 1694 9909 1698 9913
rect 1694 9904 1698 9908
rect 1694 9899 1698 9903
rect 1694 9894 1698 9898
rect 1694 9889 1698 9893
rect 1694 9884 1698 9888
rect 1694 9879 1698 9883
rect 1694 9874 1698 9878
rect 1694 9869 1698 9873
rect 1694 9864 1698 9868
rect 1758 9949 1762 9953
rect 1758 9944 1762 9948
rect 1758 9939 1762 9943
rect 1758 9934 1762 9938
rect 1758 9929 1762 9933
rect 1758 9924 1762 9928
rect 1758 9919 1762 9923
rect 1758 9914 1762 9918
rect 1758 9909 1762 9913
rect 1758 9904 1762 9908
rect 1758 9899 1762 9903
rect 1758 9894 1762 9898
rect 1758 9889 1762 9893
rect 1758 9884 1762 9888
rect 1758 9879 1762 9883
rect 1758 9874 1762 9878
rect 1758 9869 1762 9873
rect 1758 9864 1762 9868
rect 1694 9859 1698 9863
rect 1758 9859 1762 9863
rect 1694 9852 1698 9856
rect 1701 9852 1705 9856
rect 1706 9852 1710 9856
rect 1711 9852 1715 9856
rect 1716 9852 1720 9856
rect 1721 9852 1725 9856
rect 1726 9852 1730 9856
rect 1731 9852 1735 9856
rect 1736 9852 1740 9856
rect 1741 9852 1745 9856
rect 1746 9852 1750 9856
rect 1751 9852 1755 9856
rect 1758 9852 1762 9856
rect 1841 9974 1845 9978
rect 1846 9974 1850 9978
rect 1851 9974 1855 9978
rect 1856 9974 1860 9978
rect 1861 9974 1865 9978
rect 1866 9974 1870 9978
rect 1871 9974 1875 9978
rect 1876 9974 1880 9978
rect 1881 9974 1885 9978
rect 1886 9974 1890 9978
rect 1891 9974 1895 9978
rect 1896 9974 1900 9978
rect 1901 9974 1905 9978
rect 1906 9974 1910 9978
rect 1911 9974 1915 9978
rect 1916 9974 1920 9978
rect 1921 9974 1925 9978
rect 1926 9974 1930 9978
rect 1931 9974 1935 9978
rect 1841 9969 1845 9973
rect 1841 9964 1845 9968
rect 1931 9969 1935 9973
rect 1841 9959 1845 9963
rect 1841 9954 1845 9958
rect 1841 9949 1845 9953
rect 1841 9944 1845 9948
rect 1841 9939 1845 9943
rect 1841 9934 1845 9938
rect 1841 9929 1845 9933
rect 1841 9924 1845 9928
rect 1841 9919 1845 9923
rect 1841 9914 1845 9918
rect 1841 9909 1845 9913
rect 1841 9904 1845 9908
rect 1841 9899 1845 9903
rect 1841 9894 1845 9898
rect 1841 9889 1845 9893
rect 1841 9884 1845 9888
rect 1841 9879 1845 9883
rect 1841 9874 1845 9878
rect 1841 9869 1845 9873
rect 1841 9864 1845 9868
rect 1841 9859 1845 9863
rect 1841 9854 1845 9858
rect 1841 9849 1845 9853
rect 1931 9964 1935 9968
rect 1931 9959 1935 9963
rect 1931 9954 1935 9958
rect 1931 9949 1935 9953
rect 1931 9944 1935 9948
rect 1931 9939 1935 9943
rect 1931 9934 1935 9938
rect 1931 9929 1935 9933
rect 1931 9924 1935 9928
rect 1931 9919 1935 9923
rect 1931 9914 1935 9918
rect 1931 9909 1935 9913
rect 1931 9904 1935 9908
rect 1931 9899 1935 9903
rect 1931 9894 1935 9898
rect 1931 9889 1935 9893
rect 1931 9884 1935 9888
rect 1931 9879 1935 9883
rect 1931 9874 1935 9878
rect 1931 9869 1935 9873
rect 1931 9864 1935 9868
rect 1931 9859 1935 9863
rect 1931 9854 1935 9858
rect 1841 9844 1845 9848
rect 1931 9849 1935 9853
rect 1931 9844 1935 9848
rect 1841 9839 1845 9843
rect 1846 9839 1850 9843
rect 1851 9839 1855 9843
rect 1856 9839 1860 9843
rect 1861 9839 1865 9843
rect 1866 9839 1870 9843
rect 1871 9839 1875 9843
rect 1876 9839 1880 9843
rect 1881 9839 1885 9843
rect 1886 9839 1890 9843
rect 1891 9839 1895 9843
rect 1896 9839 1900 9843
rect 1901 9839 1905 9843
rect 1906 9839 1910 9843
rect 1911 9839 1915 9843
rect 1916 9839 1920 9843
rect 1921 9839 1925 9843
rect 1926 9839 1930 9843
rect 1931 9839 1935 9843
rect 2003 9961 2007 9965
rect 2010 9961 2014 9965
rect 2015 9961 2019 9965
rect 2020 9961 2024 9965
rect 2025 9961 2029 9965
rect 2030 9961 2034 9965
rect 2035 9961 2039 9965
rect 2040 9961 2044 9965
rect 2045 9961 2049 9965
rect 2050 9961 2054 9965
rect 2055 9961 2059 9965
rect 2060 9961 2064 9965
rect 2067 9961 2071 9965
rect 2003 9954 2007 9958
rect 2067 9954 2071 9958
rect 2003 9949 2007 9953
rect 2003 9944 2007 9948
rect 2003 9939 2007 9943
rect 2003 9934 2007 9938
rect 2003 9929 2007 9933
rect 2003 9924 2007 9928
rect 2003 9919 2007 9923
rect 2003 9914 2007 9918
rect 2003 9909 2007 9913
rect 2003 9904 2007 9908
rect 2003 9899 2007 9903
rect 2003 9894 2007 9898
rect 2003 9889 2007 9893
rect 2003 9884 2007 9888
rect 2003 9879 2007 9883
rect 2003 9874 2007 9878
rect 2003 9869 2007 9873
rect 2003 9864 2007 9868
rect 2067 9949 2071 9953
rect 2067 9944 2071 9948
rect 2067 9939 2071 9943
rect 2067 9934 2071 9938
rect 2067 9929 2071 9933
rect 2067 9924 2071 9928
rect 2067 9919 2071 9923
rect 2067 9914 2071 9918
rect 2067 9909 2071 9913
rect 2067 9904 2071 9908
rect 2067 9899 2071 9903
rect 2067 9894 2071 9898
rect 2067 9889 2071 9893
rect 2067 9884 2071 9888
rect 2067 9879 2071 9883
rect 2067 9874 2071 9878
rect 2067 9869 2071 9873
rect 2067 9864 2071 9868
rect 2003 9859 2007 9863
rect 2067 9859 2071 9863
rect 2003 9852 2007 9856
rect 2010 9852 2014 9856
rect 2015 9852 2019 9856
rect 2020 9852 2024 9856
rect 2025 9852 2029 9856
rect 2030 9852 2034 9856
rect 2035 9852 2039 9856
rect 2040 9852 2044 9856
rect 2045 9852 2049 9856
rect 2050 9852 2054 9856
rect 2055 9852 2059 9856
rect 2060 9852 2064 9856
rect 2067 9852 2071 9856
rect 2150 9974 2154 9978
rect 2155 9974 2159 9978
rect 2160 9974 2164 9978
rect 2165 9974 2169 9978
rect 2170 9974 2174 9978
rect 2175 9974 2179 9978
rect 2180 9974 2184 9978
rect 2185 9974 2189 9978
rect 2190 9974 2194 9978
rect 2195 9974 2199 9978
rect 2200 9974 2204 9978
rect 2205 9974 2209 9978
rect 2210 9974 2214 9978
rect 2215 9974 2219 9978
rect 2220 9974 2224 9978
rect 2225 9974 2229 9978
rect 2230 9974 2234 9978
rect 2235 9974 2239 9978
rect 2240 9974 2244 9978
rect 2150 9969 2154 9973
rect 2150 9964 2154 9968
rect 2240 9969 2244 9973
rect 2150 9959 2154 9963
rect 2150 9954 2154 9958
rect 2150 9949 2154 9953
rect 2150 9944 2154 9948
rect 2150 9939 2154 9943
rect 2150 9934 2154 9938
rect 2150 9929 2154 9933
rect 2150 9924 2154 9928
rect 2150 9919 2154 9923
rect 2150 9914 2154 9918
rect 2150 9909 2154 9913
rect 2150 9904 2154 9908
rect 2150 9899 2154 9903
rect 2150 9894 2154 9898
rect 2150 9889 2154 9893
rect 2150 9884 2154 9888
rect 2150 9879 2154 9883
rect 2150 9874 2154 9878
rect 2150 9869 2154 9873
rect 2150 9864 2154 9868
rect 2150 9859 2154 9863
rect 2150 9854 2154 9858
rect 2150 9849 2154 9853
rect 2240 9964 2244 9968
rect 2240 9959 2244 9963
rect 2240 9954 2244 9958
rect 2240 9949 2244 9953
rect 2240 9944 2244 9948
rect 2240 9939 2244 9943
rect 2240 9934 2244 9938
rect 2240 9929 2244 9933
rect 2240 9924 2244 9928
rect 2240 9919 2244 9923
rect 2240 9914 2244 9918
rect 2240 9909 2244 9913
rect 2240 9904 2244 9908
rect 2240 9899 2244 9903
rect 2240 9894 2244 9898
rect 2240 9889 2244 9893
rect 2240 9884 2244 9888
rect 2240 9879 2244 9883
rect 2240 9874 2244 9878
rect 2240 9869 2244 9873
rect 2240 9864 2244 9868
rect 2240 9859 2244 9863
rect 2240 9854 2244 9858
rect 2150 9844 2154 9848
rect 2240 9849 2244 9853
rect 2240 9844 2244 9848
rect 2150 9839 2154 9843
rect 2155 9839 2159 9843
rect 2160 9839 2164 9843
rect 2165 9839 2169 9843
rect 2170 9839 2174 9843
rect 2175 9839 2179 9843
rect 2180 9839 2184 9843
rect 2185 9839 2189 9843
rect 2190 9839 2194 9843
rect 2195 9839 2199 9843
rect 2200 9839 2204 9843
rect 2205 9839 2209 9843
rect 2210 9839 2214 9843
rect 2215 9839 2219 9843
rect 2220 9839 2224 9843
rect 2225 9839 2229 9843
rect 2230 9839 2234 9843
rect 2235 9839 2239 9843
rect 2240 9839 2244 9843
rect 2312 9961 2316 9965
rect 2319 9961 2323 9965
rect 2324 9961 2328 9965
rect 2329 9961 2333 9965
rect 2334 9961 2338 9965
rect 2339 9961 2343 9965
rect 2344 9961 2348 9965
rect 2349 9961 2353 9965
rect 2354 9961 2358 9965
rect 2359 9961 2363 9965
rect 2364 9961 2368 9965
rect 2369 9961 2373 9965
rect 2376 9961 2380 9965
rect 2312 9954 2316 9958
rect 2376 9954 2380 9958
rect 2312 9949 2316 9953
rect 2312 9944 2316 9948
rect 2312 9939 2316 9943
rect 2312 9934 2316 9938
rect 2312 9929 2316 9933
rect 2312 9924 2316 9928
rect 2312 9919 2316 9923
rect 2312 9914 2316 9918
rect 2312 9909 2316 9913
rect 2312 9904 2316 9908
rect 2312 9899 2316 9903
rect 2312 9894 2316 9898
rect 2312 9889 2316 9893
rect 2312 9884 2316 9888
rect 2312 9879 2316 9883
rect 2312 9874 2316 9878
rect 2312 9869 2316 9873
rect 2312 9864 2316 9868
rect 2376 9949 2380 9953
rect 2376 9944 2380 9948
rect 2376 9939 2380 9943
rect 2376 9934 2380 9938
rect 2376 9929 2380 9933
rect 2376 9924 2380 9928
rect 2376 9919 2380 9923
rect 2376 9914 2380 9918
rect 2376 9909 2380 9913
rect 2376 9904 2380 9908
rect 2376 9899 2380 9903
rect 2376 9894 2380 9898
rect 2376 9889 2380 9893
rect 2376 9884 2380 9888
rect 2376 9879 2380 9883
rect 2376 9874 2380 9878
rect 2376 9869 2380 9873
rect 2376 9864 2380 9868
rect 2312 9859 2316 9863
rect 2376 9859 2380 9863
rect 2312 9852 2316 9856
rect 2319 9852 2323 9856
rect 2324 9852 2328 9856
rect 2329 9852 2333 9856
rect 2334 9852 2338 9856
rect 2339 9852 2343 9856
rect 2344 9852 2348 9856
rect 2349 9852 2353 9856
rect 2354 9852 2358 9856
rect 2359 9852 2363 9856
rect 2364 9852 2368 9856
rect 2369 9852 2373 9856
rect 2376 9852 2380 9856
rect 2459 9974 2463 9978
rect 2464 9974 2468 9978
rect 2469 9974 2473 9978
rect 2474 9974 2478 9978
rect 2479 9974 2483 9978
rect 2484 9974 2488 9978
rect 2489 9974 2493 9978
rect 2494 9974 2498 9978
rect 2499 9974 2503 9978
rect 2504 9974 2508 9978
rect 2509 9974 2513 9978
rect 2514 9974 2518 9978
rect 2519 9974 2523 9978
rect 2524 9974 2528 9978
rect 2529 9974 2533 9978
rect 2534 9974 2538 9978
rect 2539 9974 2543 9978
rect 2544 9974 2548 9978
rect 2549 9974 2553 9978
rect 2459 9969 2463 9973
rect 2459 9964 2463 9968
rect 2549 9969 2553 9973
rect 2459 9959 2463 9963
rect 2459 9954 2463 9958
rect 2459 9949 2463 9953
rect 2459 9944 2463 9948
rect 2459 9939 2463 9943
rect 2459 9934 2463 9938
rect 2459 9929 2463 9933
rect 2459 9924 2463 9928
rect 2459 9919 2463 9923
rect 2459 9914 2463 9918
rect 2459 9909 2463 9913
rect 2459 9904 2463 9908
rect 2459 9899 2463 9903
rect 2459 9894 2463 9898
rect 2459 9889 2463 9893
rect 2459 9884 2463 9888
rect 2459 9879 2463 9883
rect 2459 9874 2463 9878
rect 2459 9869 2463 9873
rect 2459 9864 2463 9868
rect 2459 9859 2463 9863
rect 2459 9854 2463 9858
rect 2459 9849 2463 9853
rect 2549 9964 2553 9968
rect 2549 9959 2553 9963
rect 2549 9954 2553 9958
rect 2549 9949 2553 9953
rect 2549 9944 2553 9948
rect 2549 9939 2553 9943
rect 2549 9934 2553 9938
rect 2549 9929 2553 9933
rect 2549 9924 2553 9928
rect 2549 9919 2553 9923
rect 2549 9914 2553 9918
rect 2549 9909 2553 9913
rect 2549 9904 2553 9908
rect 2549 9899 2553 9903
rect 2549 9894 2553 9898
rect 2549 9889 2553 9893
rect 2549 9884 2553 9888
rect 2549 9879 2553 9883
rect 2549 9874 2553 9878
rect 2549 9869 2553 9873
rect 2549 9864 2553 9868
rect 2549 9859 2553 9863
rect 2549 9854 2553 9858
rect 2459 9844 2463 9848
rect 2549 9849 2553 9853
rect 2549 9844 2553 9848
rect 2459 9839 2463 9843
rect 2464 9839 2468 9843
rect 2469 9839 2473 9843
rect 2474 9839 2478 9843
rect 2479 9839 2483 9843
rect 2484 9839 2488 9843
rect 2489 9839 2493 9843
rect 2494 9839 2498 9843
rect 2499 9839 2503 9843
rect 2504 9839 2508 9843
rect 2509 9839 2513 9843
rect 2514 9839 2518 9843
rect 2519 9839 2523 9843
rect 2524 9839 2528 9843
rect 2529 9839 2533 9843
rect 2534 9839 2538 9843
rect 2539 9839 2543 9843
rect 2544 9839 2548 9843
rect 2549 9839 2553 9843
rect 2621 9961 2625 9965
rect 2628 9961 2632 9965
rect 2633 9961 2637 9965
rect 2638 9961 2642 9965
rect 2643 9961 2647 9965
rect 2648 9961 2652 9965
rect 2653 9961 2657 9965
rect 2658 9961 2662 9965
rect 2663 9961 2667 9965
rect 2668 9961 2672 9965
rect 2673 9961 2677 9965
rect 2678 9961 2682 9965
rect 2685 9961 2689 9965
rect 2621 9954 2625 9958
rect 2685 9954 2689 9958
rect 2621 9949 2625 9953
rect 2621 9944 2625 9948
rect 2621 9939 2625 9943
rect 2621 9934 2625 9938
rect 2621 9929 2625 9933
rect 2621 9924 2625 9928
rect 2621 9919 2625 9923
rect 2621 9914 2625 9918
rect 2621 9909 2625 9913
rect 2621 9904 2625 9908
rect 2621 9899 2625 9903
rect 2621 9894 2625 9898
rect 2621 9889 2625 9893
rect 2621 9884 2625 9888
rect 2621 9879 2625 9883
rect 2621 9874 2625 9878
rect 2621 9869 2625 9873
rect 2621 9864 2625 9868
rect 2685 9949 2689 9953
rect 2685 9944 2689 9948
rect 2685 9939 2689 9943
rect 2685 9934 2689 9938
rect 2685 9929 2689 9933
rect 2685 9924 2689 9928
rect 2685 9919 2689 9923
rect 2685 9914 2689 9918
rect 2685 9909 2689 9913
rect 2685 9904 2689 9908
rect 2685 9899 2689 9903
rect 2685 9894 2689 9898
rect 2685 9889 2689 9893
rect 2685 9884 2689 9888
rect 2685 9879 2689 9883
rect 2685 9874 2689 9878
rect 2685 9869 2689 9873
rect 2685 9864 2689 9868
rect 2621 9859 2625 9863
rect 2685 9859 2689 9863
rect 2621 9852 2625 9856
rect 2628 9852 2632 9856
rect 2633 9852 2637 9856
rect 2638 9852 2642 9856
rect 2643 9852 2647 9856
rect 2648 9852 2652 9856
rect 2653 9852 2657 9856
rect 2658 9852 2662 9856
rect 2663 9852 2667 9856
rect 2668 9852 2672 9856
rect 2673 9852 2677 9856
rect 2678 9852 2682 9856
rect 2685 9852 2689 9856
rect 2768 9974 2772 9978
rect 2773 9974 2777 9978
rect 2778 9974 2782 9978
rect 2783 9974 2787 9978
rect 2788 9974 2792 9978
rect 2793 9974 2797 9978
rect 2798 9974 2802 9978
rect 2803 9974 2807 9978
rect 2808 9974 2812 9978
rect 2813 9974 2817 9978
rect 2818 9974 2822 9978
rect 2823 9974 2827 9978
rect 2828 9974 2832 9978
rect 2833 9974 2837 9978
rect 2838 9974 2842 9978
rect 2843 9974 2847 9978
rect 2848 9974 2852 9978
rect 2853 9974 2857 9978
rect 2858 9974 2862 9978
rect 2768 9969 2772 9973
rect 2768 9964 2772 9968
rect 2858 9969 2862 9973
rect 2768 9959 2772 9963
rect 2768 9954 2772 9958
rect 2768 9949 2772 9953
rect 2768 9944 2772 9948
rect 2768 9939 2772 9943
rect 2768 9934 2772 9938
rect 2768 9929 2772 9933
rect 2768 9924 2772 9928
rect 2768 9919 2772 9923
rect 2768 9914 2772 9918
rect 2768 9909 2772 9913
rect 2768 9904 2772 9908
rect 2768 9899 2772 9903
rect 2768 9894 2772 9898
rect 2768 9889 2772 9893
rect 2768 9884 2772 9888
rect 2768 9879 2772 9883
rect 2768 9874 2772 9878
rect 2768 9869 2772 9873
rect 2768 9864 2772 9868
rect 2768 9859 2772 9863
rect 2768 9854 2772 9858
rect 2768 9849 2772 9853
rect 2858 9964 2862 9968
rect 2858 9959 2862 9963
rect 2858 9954 2862 9958
rect 2858 9949 2862 9953
rect 2858 9944 2862 9948
rect 2858 9939 2862 9943
rect 2858 9934 2862 9938
rect 2858 9929 2862 9933
rect 2858 9924 2862 9928
rect 2858 9919 2862 9923
rect 2858 9914 2862 9918
rect 2858 9909 2862 9913
rect 2858 9904 2862 9908
rect 2858 9899 2862 9903
rect 2858 9894 2862 9898
rect 2858 9889 2862 9893
rect 2858 9884 2862 9888
rect 2858 9879 2862 9883
rect 2858 9874 2862 9878
rect 2858 9869 2862 9873
rect 2858 9864 2862 9868
rect 2858 9859 2862 9863
rect 2858 9854 2862 9858
rect 2768 9844 2772 9848
rect 2858 9849 2862 9853
rect 2858 9844 2862 9848
rect 2768 9839 2772 9843
rect 2773 9839 2777 9843
rect 2778 9839 2782 9843
rect 2783 9839 2787 9843
rect 2788 9839 2792 9843
rect 2793 9839 2797 9843
rect 2798 9839 2802 9843
rect 2803 9839 2807 9843
rect 2808 9839 2812 9843
rect 2813 9839 2817 9843
rect 2818 9839 2822 9843
rect 2823 9839 2827 9843
rect 2828 9839 2832 9843
rect 2833 9839 2837 9843
rect 2838 9839 2842 9843
rect 2843 9839 2847 9843
rect 2848 9839 2852 9843
rect 2853 9839 2857 9843
rect 2858 9839 2862 9843
rect 2930 9961 2934 9965
rect 2937 9961 2941 9965
rect 2942 9961 2946 9965
rect 2947 9961 2951 9965
rect 2952 9961 2956 9965
rect 2957 9961 2961 9965
rect 2962 9961 2966 9965
rect 2967 9961 2971 9965
rect 2972 9961 2976 9965
rect 2977 9961 2981 9965
rect 2982 9961 2986 9965
rect 2987 9961 2991 9965
rect 2994 9961 2998 9965
rect 2930 9954 2934 9958
rect 2994 9954 2998 9958
rect 2930 9949 2934 9953
rect 2930 9944 2934 9948
rect 2930 9939 2934 9943
rect 2930 9934 2934 9938
rect 2930 9929 2934 9933
rect 2930 9924 2934 9928
rect 2930 9919 2934 9923
rect 2930 9914 2934 9918
rect 2930 9909 2934 9913
rect 2930 9904 2934 9908
rect 2930 9899 2934 9903
rect 2930 9894 2934 9898
rect 2930 9889 2934 9893
rect 2930 9884 2934 9888
rect 2930 9879 2934 9883
rect 2930 9874 2934 9878
rect 2930 9869 2934 9873
rect 2930 9864 2934 9868
rect 2994 9949 2998 9953
rect 2994 9944 2998 9948
rect 2994 9939 2998 9943
rect 2994 9934 2998 9938
rect 2994 9929 2998 9933
rect 2994 9924 2998 9928
rect 2994 9919 2998 9923
rect 2994 9914 2998 9918
rect 2994 9909 2998 9913
rect 2994 9904 2998 9908
rect 2994 9899 2998 9903
rect 2994 9894 2998 9898
rect 2994 9889 2998 9893
rect 2994 9884 2998 9888
rect 2994 9879 2998 9883
rect 2994 9874 2998 9878
rect 2994 9869 2998 9873
rect 2994 9864 2998 9868
rect 2930 9859 2934 9863
rect 2994 9859 2998 9863
rect 2930 9852 2934 9856
rect 2937 9852 2941 9856
rect 2942 9852 2946 9856
rect 2947 9852 2951 9856
rect 2952 9852 2956 9856
rect 2957 9852 2961 9856
rect 2962 9852 2966 9856
rect 2967 9852 2971 9856
rect 2972 9852 2976 9856
rect 2977 9852 2981 9856
rect 2982 9852 2986 9856
rect 2987 9852 2991 9856
rect 2994 9852 2998 9856
rect 3077 9974 3081 9978
rect 3082 9974 3086 9978
rect 3087 9974 3091 9978
rect 3092 9974 3096 9978
rect 3097 9974 3101 9978
rect 3102 9974 3106 9978
rect 3107 9974 3111 9978
rect 3112 9974 3116 9978
rect 3117 9974 3121 9978
rect 3122 9974 3126 9978
rect 3127 9974 3131 9978
rect 3132 9974 3136 9978
rect 3137 9974 3141 9978
rect 3142 9974 3146 9978
rect 3147 9974 3151 9978
rect 3152 9974 3156 9978
rect 3157 9974 3161 9978
rect 3162 9974 3166 9978
rect 3167 9974 3171 9978
rect 3077 9969 3081 9973
rect 3077 9964 3081 9968
rect 3167 9969 3171 9973
rect 3077 9959 3081 9963
rect 3077 9954 3081 9958
rect 3077 9949 3081 9953
rect 3077 9944 3081 9948
rect 3077 9939 3081 9943
rect 3077 9934 3081 9938
rect 3077 9929 3081 9933
rect 3077 9924 3081 9928
rect 3077 9919 3081 9923
rect 3077 9914 3081 9918
rect 3077 9909 3081 9913
rect 3077 9904 3081 9908
rect 3077 9899 3081 9903
rect 3077 9894 3081 9898
rect 3077 9889 3081 9893
rect 3077 9884 3081 9888
rect 3077 9879 3081 9883
rect 3077 9874 3081 9878
rect 3077 9869 3081 9873
rect 3077 9864 3081 9868
rect 3077 9859 3081 9863
rect 3077 9854 3081 9858
rect 3077 9849 3081 9853
rect 3167 9964 3171 9968
rect 3167 9959 3171 9963
rect 3167 9954 3171 9958
rect 3167 9949 3171 9953
rect 3167 9944 3171 9948
rect 3167 9939 3171 9943
rect 3167 9934 3171 9938
rect 3167 9929 3171 9933
rect 3167 9924 3171 9928
rect 3167 9919 3171 9923
rect 3167 9914 3171 9918
rect 3167 9909 3171 9913
rect 3167 9904 3171 9908
rect 3167 9899 3171 9903
rect 3167 9894 3171 9898
rect 3167 9889 3171 9893
rect 3167 9884 3171 9888
rect 3167 9879 3171 9883
rect 3167 9874 3171 9878
rect 3167 9869 3171 9873
rect 3167 9864 3171 9868
rect 3167 9859 3171 9863
rect 3167 9854 3171 9858
rect 3077 9844 3081 9848
rect 3167 9849 3171 9853
rect 3167 9844 3171 9848
rect 3077 9839 3081 9843
rect 3082 9839 3086 9843
rect 3087 9839 3091 9843
rect 3092 9839 3096 9843
rect 3097 9839 3101 9843
rect 3102 9839 3106 9843
rect 3107 9839 3111 9843
rect 3112 9839 3116 9843
rect 3117 9839 3121 9843
rect 3122 9839 3126 9843
rect 3127 9839 3131 9843
rect 3132 9839 3136 9843
rect 3137 9839 3141 9843
rect 3142 9839 3146 9843
rect 3147 9839 3151 9843
rect 3152 9839 3156 9843
rect 3157 9839 3161 9843
rect 3162 9839 3166 9843
rect 3167 9839 3171 9843
rect 3239 9961 3243 9965
rect 3246 9961 3250 9965
rect 3251 9961 3255 9965
rect 3256 9961 3260 9965
rect 3261 9961 3265 9965
rect 3266 9961 3270 9965
rect 3271 9961 3275 9965
rect 3276 9961 3280 9965
rect 3281 9961 3285 9965
rect 3286 9961 3290 9965
rect 3291 9961 3295 9965
rect 3296 9961 3300 9965
rect 3303 9961 3307 9965
rect 3239 9954 3243 9958
rect 3303 9954 3307 9958
rect 3239 9949 3243 9953
rect 3239 9944 3243 9948
rect 3239 9939 3243 9943
rect 3239 9934 3243 9938
rect 3239 9929 3243 9933
rect 3239 9924 3243 9928
rect 3239 9919 3243 9923
rect 3239 9914 3243 9918
rect 3239 9909 3243 9913
rect 3239 9904 3243 9908
rect 3239 9899 3243 9903
rect 3239 9894 3243 9898
rect 3239 9889 3243 9893
rect 3239 9884 3243 9888
rect 3239 9879 3243 9883
rect 3239 9874 3243 9878
rect 3239 9869 3243 9873
rect 3239 9864 3243 9868
rect 3303 9949 3307 9953
rect 3303 9944 3307 9948
rect 3303 9939 3307 9943
rect 3303 9934 3307 9938
rect 3303 9929 3307 9933
rect 3303 9924 3307 9928
rect 3303 9919 3307 9923
rect 3303 9914 3307 9918
rect 3303 9909 3307 9913
rect 3303 9904 3307 9908
rect 3303 9899 3307 9903
rect 3303 9894 3307 9898
rect 3303 9889 3307 9893
rect 3303 9884 3307 9888
rect 3303 9879 3307 9883
rect 3303 9874 3307 9878
rect 3303 9869 3307 9873
rect 3303 9864 3307 9868
rect 3239 9859 3243 9863
rect 3303 9859 3307 9863
rect 3239 9852 3243 9856
rect 3246 9852 3250 9856
rect 3251 9852 3255 9856
rect 3256 9852 3260 9856
rect 3261 9852 3265 9856
rect 3266 9852 3270 9856
rect 3271 9852 3275 9856
rect 3276 9852 3280 9856
rect 3281 9852 3285 9856
rect 3286 9852 3290 9856
rect 3291 9852 3295 9856
rect 3296 9852 3300 9856
rect 3303 9852 3307 9856
rect 3386 9974 3390 9978
rect 3391 9974 3395 9978
rect 3396 9974 3400 9978
rect 3401 9974 3405 9978
rect 3406 9974 3410 9978
rect 3411 9974 3415 9978
rect 3416 9974 3420 9978
rect 3421 9974 3425 9978
rect 3426 9974 3430 9978
rect 3431 9974 3435 9978
rect 3436 9974 3440 9978
rect 3441 9974 3445 9978
rect 3446 9974 3450 9978
rect 3451 9974 3455 9978
rect 3456 9974 3460 9978
rect 3461 9974 3465 9978
rect 3466 9974 3470 9978
rect 3471 9974 3475 9978
rect 3476 9974 3480 9978
rect 3386 9969 3390 9973
rect 3386 9964 3390 9968
rect 3476 9969 3480 9973
rect 3386 9959 3390 9963
rect 3386 9954 3390 9958
rect 3386 9949 3390 9953
rect 3386 9944 3390 9948
rect 3386 9939 3390 9943
rect 3386 9934 3390 9938
rect 3386 9929 3390 9933
rect 3386 9924 3390 9928
rect 3386 9919 3390 9923
rect 3386 9914 3390 9918
rect 3386 9909 3390 9913
rect 3386 9904 3390 9908
rect 3386 9899 3390 9903
rect 3386 9894 3390 9898
rect 3386 9889 3390 9893
rect 3386 9884 3390 9888
rect 3386 9879 3390 9883
rect 3386 9874 3390 9878
rect 3386 9869 3390 9873
rect 3386 9864 3390 9868
rect 3386 9859 3390 9863
rect 3386 9854 3390 9858
rect 3386 9849 3390 9853
rect 3476 9964 3480 9968
rect 3476 9959 3480 9963
rect 3476 9954 3480 9958
rect 3476 9949 3480 9953
rect 3476 9944 3480 9948
rect 3476 9939 3480 9943
rect 3476 9934 3480 9938
rect 3476 9929 3480 9933
rect 3476 9924 3480 9928
rect 3476 9919 3480 9923
rect 3476 9914 3480 9918
rect 3476 9909 3480 9913
rect 3476 9904 3480 9908
rect 3476 9899 3480 9903
rect 3476 9894 3480 9898
rect 3476 9889 3480 9893
rect 3476 9884 3480 9888
rect 3476 9879 3480 9883
rect 3476 9874 3480 9878
rect 3476 9869 3480 9873
rect 3476 9864 3480 9868
rect 3476 9859 3480 9863
rect 3476 9854 3480 9858
rect 3386 9844 3390 9848
rect 3476 9849 3480 9853
rect 3476 9844 3480 9848
rect 3386 9839 3390 9843
rect 3391 9839 3395 9843
rect 3396 9839 3400 9843
rect 3401 9839 3405 9843
rect 3406 9839 3410 9843
rect 3411 9839 3415 9843
rect 3416 9839 3420 9843
rect 3421 9839 3425 9843
rect 3426 9839 3430 9843
rect 3431 9839 3435 9843
rect 3436 9839 3440 9843
rect 3441 9839 3445 9843
rect 3446 9839 3450 9843
rect 3451 9839 3455 9843
rect 3456 9839 3460 9843
rect 3461 9839 3465 9843
rect 3466 9839 3470 9843
rect 3471 9839 3475 9843
rect 3476 9839 3480 9843
rect 3548 9961 3552 9965
rect 3555 9961 3559 9965
rect 3560 9961 3564 9965
rect 3565 9961 3569 9965
rect 3570 9961 3574 9965
rect 3575 9961 3579 9965
rect 3580 9961 3584 9965
rect 3585 9961 3589 9965
rect 3590 9961 3594 9965
rect 3595 9961 3599 9965
rect 3600 9961 3604 9965
rect 3605 9961 3609 9965
rect 3612 9961 3616 9965
rect 3548 9954 3552 9958
rect 3612 9954 3616 9958
rect 3548 9949 3552 9953
rect 3548 9944 3552 9948
rect 3548 9939 3552 9943
rect 3548 9934 3552 9938
rect 3548 9929 3552 9933
rect 3548 9924 3552 9928
rect 3548 9919 3552 9923
rect 3548 9914 3552 9918
rect 3548 9909 3552 9913
rect 3548 9904 3552 9908
rect 3548 9899 3552 9903
rect 3548 9894 3552 9898
rect 3548 9889 3552 9893
rect 3548 9884 3552 9888
rect 3548 9879 3552 9883
rect 3548 9874 3552 9878
rect 3548 9869 3552 9873
rect 3548 9864 3552 9868
rect 3612 9949 3616 9953
rect 3612 9944 3616 9948
rect 3612 9939 3616 9943
rect 3612 9934 3616 9938
rect 3612 9929 3616 9933
rect 3612 9924 3616 9928
rect 3612 9919 3616 9923
rect 3612 9914 3616 9918
rect 3612 9909 3616 9913
rect 3612 9904 3616 9908
rect 3612 9899 3616 9903
rect 3612 9894 3616 9898
rect 3612 9889 3616 9893
rect 3612 9884 3616 9888
rect 3612 9879 3616 9883
rect 3612 9874 3616 9878
rect 3612 9869 3616 9873
rect 3612 9864 3616 9868
rect 3548 9859 3552 9863
rect 3612 9859 3616 9863
rect 3548 9852 3552 9856
rect 3555 9852 3559 9856
rect 3560 9852 3564 9856
rect 3565 9852 3569 9856
rect 3570 9852 3574 9856
rect 3575 9852 3579 9856
rect 3580 9852 3584 9856
rect 3585 9852 3589 9856
rect 3590 9852 3594 9856
rect 3595 9852 3599 9856
rect 3600 9852 3604 9856
rect 3605 9852 3609 9856
rect 3612 9852 3616 9856
rect 3695 9974 3699 9978
rect 3700 9974 3704 9978
rect 3705 9974 3709 9978
rect 3710 9974 3714 9978
rect 3715 9974 3719 9978
rect 3720 9974 3724 9978
rect 3725 9974 3729 9978
rect 3730 9974 3734 9978
rect 3735 9974 3739 9978
rect 3740 9974 3744 9978
rect 3745 9974 3749 9978
rect 3750 9974 3754 9978
rect 3755 9974 3759 9978
rect 3760 9974 3764 9978
rect 3765 9974 3769 9978
rect 3770 9974 3774 9978
rect 3775 9974 3779 9978
rect 3780 9974 3784 9978
rect 3785 9974 3789 9978
rect 3695 9969 3699 9973
rect 3695 9964 3699 9968
rect 3785 9969 3789 9973
rect 3695 9959 3699 9963
rect 3695 9954 3699 9958
rect 3695 9949 3699 9953
rect 3695 9944 3699 9948
rect 3695 9939 3699 9943
rect 3695 9934 3699 9938
rect 3695 9929 3699 9933
rect 3695 9924 3699 9928
rect 3695 9919 3699 9923
rect 3695 9914 3699 9918
rect 3695 9909 3699 9913
rect 3695 9904 3699 9908
rect 3695 9899 3699 9903
rect 3695 9894 3699 9898
rect 3695 9889 3699 9893
rect 3695 9884 3699 9888
rect 3695 9879 3699 9883
rect 3695 9874 3699 9878
rect 3695 9869 3699 9873
rect 3695 9864 3699 9868
rect 3695 9859 3699 9863
rect 3695 9854 3699 9858
rect 3695 9849 3699 9853
rect 3785 9964 3789 9968
rect 3785 9959 3789 9963
rect 3785 9954 3789 9958
rect 3785 9949 3789 9953
rect 3785 9944 3789 9948
rect 3785 9939 3789 9943
rect 3785 9934 3789 9938
rect 3785 9929 3789 9933
rect 3785 9924 3789 9928
rect 3785 9919 3789 9923
rect 3785 9914 3789 9918
rect 3785 9909 3789 9913
rect 3785 9904 3789 9908
rect 3785 9899 3789 9903
rect 3785 9894 3789 9898
rect 3785 9889 3789 9893
rect 3785 9884 3789 9888
rect 3785 9879 3789 9883
rect 3785 9874 3789 9878
rect 3785 9869 3789 9873
rect 3785 9864 3789 9868
rect 3785 9859 3789 9863
rect 3785 9854 3789 9858
rect 3695 9844 3699 9848
rect 3785 9849 3789 9853
rect 3785 9844 3789 9848
rect 3695 9839 3699 9843
rect 3700 9839 3704 9843
rect 3705 9839 3709 9843
rect 3710 9839 3714 9843
rect 3715 9839 3719 9843
rect 3720 9839 3724 9843
rect 3725 9839 3729 9843
rect 3730 9839 3734 9843
rect 3735 9839 3739 9843
rect 3740 9839 3744 9843
rect 3745 9839 3749 9843
rect 3750 9839 3754 9843
rect 3755 9839 3759 9843
rect 3760 9839 3764 9843
rect 3765 9839 3769 9843
rect 3770 9839 3774 9843
rect 3775 9839 3779 9843
rect 3780 9839 3784 9843
rect 3785 9839 3789 9843
rect 3857 9961 3861 9965
rect 3864 9961 3868 9965
rect 3869 9961 3873 9965
rect 3874 9961 3878 9965
rect 3879 9961 3883 9965
rect 3884 9961 3888 9965
rect 3889 9961 3893 9965
rect 3894 9961 3898 9965
rect 3899 9961 3903 9965
rect 3904 9961 3908 9965
rect 3909 9961 3913 9965
rect 3914 9961 3918 9965
rect 3921 9961 3925 9965
rect 3857 9954 3861 9958
rect 3921 9954 3925 9958
rect 3857 9949 3861 9953
rect 3857 9944 3861 9948
rect 3857 9939 3861 9943
rect 3857 9934 3861 9938
rect 3857 9929 3861 9933
rect 3857 9924 3861 9928
rect 3857 9919 3861 9923
rect 3857 9914 3861 9918
rect 3857 9909 3861 9913
rect 3857 9904 3861 9908
rect 3857 9899 3861 9903
rect 3857 9894 3861 9898
rect 3857 9889 3861 9893
rect 3857 9884 3861 9888
rect 3857 9879 3861 9883
rect 3857 9874 3861 9878
rect 3857 9869 3861 9873
rect 3857 9864 3861 9868
rect 3921 9949 3925 9953
rect 3921 9944 3925 9948
rect 3921 9939 3925 9943
rect 3921 9934 3925 9938
rect 3921 9929 3925 9933
rect 3921 9924 3925 9928
rect 3921 9919 3925 9923
rect 3921 9914 3925 9918
rect 3921 9909 3925 9913
rect 3921 9904 3925 9908
rect 3921 9899 3925 9903
rect 3921 9894 3925 9898
rect 3921 9889 3925 9893
rect 3921 9884 3925 9888
rect 3921 9879 3925 9883
rect 3921 9874 3925 9878
rect 3921 9869 3925 9873
rect 3921 9864 3925 9868
rect 3857 9859 3861 9863
rect 3921 9859 3925 9863
rect 3857 9852 3861 9856
rect 3864 9852 3868 9856
rect 3869 9852 3873 9856
rect 3874 9852 3878 9856
rect 3879 9852 3883 9856
rect 3884 9852 3888 9856
rect 3889 9852 3893 9856
rect 3894 9852 3898 9856
rect 3899 9852 3903 9856
rect 3904 9852 3908 9856
rect 3909 9852 3913 9856
rect 3914 9852 3918 9856
rect 3921 9852 3925 9856
rect 4004 9974 4008 9978
rect 4009 9974 4013 9978
rect 4014 9974 4018 9978
rect 4019 9974 4023 9978
rect 4024 9974 4028 9978
rect 4029 9974 4033 9978
rect 4034 9974 4038 9978
rect 4039 9974 4043 9978
rect 4044 9974 4048 9978
rect 4049 9974 4053 9978
rect 4054 9974 4058 9978
rect 4059 9974 4063 9978
rect 4064 9974 4068 9978
rect 4069 9974 4073 9978
rect 4074 9974 4078 9978
rect 4079 9974 4083 9978
rect 4084 9974 4088 9978
rect 4089 9974 4093 9978
rect 4094 9974 4098 9978
rect 4004 9969 4008 9973
rect 4004 9964 4008 9968
rect 4094 9969 4098 9973
rect 4004 9959 4008 9963
rect 4004 9954 4008 9958
rect 4004 9949 4008 9953
rect 4004 9944 4008 9948
rect 4004 9939 4008 9943
rect 4004 9934 4008 9938
rect 4004 9929 4008 9933
rect 4004 9924 4008 9928
rect 4004 9919 4008 9923
rect 4004 9914 4008 9918
rect 4004 9909 4008 9913
rect 4004 9904 4008 9908
rect 4004 9899 4008 9903
rect 4004 9894 4008 9898
rect 4004 9889 4008 9893
rect 4004 9884 4008 9888
rect 4004 9879 4008 9883
rect 4004 9874 4008 9878
rect 4004 9869 4008 9873
rect 4004 9864 4008 9868
rect 4004 9859 4008 9863
rect 4004 9854 4008 9858
rect 4004 9849 4008 9853
rect 4094 9964 4098 9968
rect 4094 9959 4098 9963
rect 4094 9954 4098 9958
rect 4094 9949 4098 9953
rect 4094 9944 4098 9948
rect 4094 9939 4098 9943
rect 4094 9934 4098 9938
rect 4094 9929 4098 9933
rect 4094 9924 4098 9928
rect 4094 9919 4098 9923
rect 4094 9914 4098 9918
rect 4094 9909 4098 9913
rect 4094 9904 4098 9908
rect 4094 9899 4098 9903
rect 4094 9894 4098 9898
rect 4094 9889 4098 9893
rect 4094 9884 4098 9888
rect 4094 9879 4098 9883
rect 4094 9874 4098 9878
rect 4094 9869 4098 9873
rect 4094 9864 4098 9868
rect 4094 9859 4098 9863
rect 4094 9854 4098 9858
rect 4004 9844 4008 9848
rect 4094 9849 4098 9853
rect 4094 9844 4098 9848
rect 4004 9839 4008 9843
rect 4009 9839 4013 9843
rect 4014 9839 4018 9843
rect 4019 9839 4023 9843
rect 4024 9839 4028 9843
rect 4029 9839 4033 9843
rect 4034 9839 4038 9843
rect 4039 9839 4043 9843
rect 4044 9839 4048 9843
rect 4049 9839 4053 9843
rect 4054 9839 4058 9843
rect 4059 9839 4063 9843
rect 4064 9839 4068 9843
rect 4069 9839 4073 9843
rect 4074 9839 4078 9843
rect 4079 9839 4083 9843
rect 4084 9839 4088 9843
rect 4089 9839 4093 9843
rect 4094 9839 4098 9843
rect 802 9716 806 9720
rect 807 9716 811 9720
rect 812 9716 816 9720
rect 817 9716 821 9720
rect 831 9716 835 9720
rect 836 9716 840 9720
rect 841 9716 845 9720
rect 846 9716 850 9720
rect 860 9716 864 9720
rect 865 9716 869 9720
rect 870 9716 874 9720
rect 875 9716 879 9720
rect 889 9716 893 9720
rect 894 9716 898 9720
rect 899 9716 903 9720
rect 904 9716 908 9720
rect 918 9716 922 9720
rect 923 9716 927 9720
rect 928 9716 932 9720
rect 933 9716 937 9720
rect 1319 9716 1323 9720
rect 1324 9716 1328 9720
rect 1329 9716 1333 9720
rect 1334 9716 1338 9720
rect 1628 9716 1632 9720
rect 1633 9716 1637 9720
rect 1638 9716 1642 9720
rect 1643 9716 1647 9720
rect 1937 9716 1941 9720
rect 1942 9716 1946 9720
rect 1947 9716 1951 9720
rect 1952 9716 1956 9720
rect 2246 9716 2250 9720
rect 2251 9716 2255 9720
rect 2256 9716 2260 9720
rect 2261 9716 2265 9720
rect 2555 9716 2559 9720
rect 2560 9716 2564 9720
rect 2565 9716 2569 9720
rect 2570 9716 2574 9720
rect 2864 9716 2868 9720
rect 2869 9716 2873 9720
rect 2874 9716 2878 9720
rect 2879 9716 2883 9720
rect 3173 9716 3177 9720
rect 3178 9716 3182 9720
rect 3183 9716 3187 9720
rect 3188 9716 3192 9720
rect 3482 9716 3486 9720
rect 3487 9716 3491 9720
rect 3492 9716 3496 9720
rect 3497 9716 3501 9720
rect 3791 9716 3795 9720
rect 3796 9716 3800 9720
rect 3801 9716 3805 9720
rect 3806 9716 3810 9720
rect 4100 9716 4104 9720
rect 4105 9716 4109 9720
rect 4110 9716 4114 9720
rect 4115 9716 4119 9720
rect 4292 9716 4296 9720
rect 4297 9716 4301 9720
rect 4302 9716 4306 9720
rect 4307 9716 4311 9720
rect 4318 9716 4322 9720
rect 4323 9716 4327 9720
rect 4328 9716 4332 9720
rect 4333 9716 4337 9720
rect 4344 9716 4348 9720
rect 4349 9716 4353 9720
rect 4354 9716 4358 9720
rect 4359 9716 4363 9720
rect 4370 9716 4374 9720
rect 4375 9716 4379 9720
rect 4380 9716 4384 9720
rect 4385 9716 4389 9720
rect 4396 9716 4400 9720
rect 4401 9716 4405 9720
rect 4406 9716 4410 9720
rect 4411 9716 4415 9720
rect 802 9706 806 9710
rect 807 9706 811 9710
rect 812 9706 816 9710
rect 817 9706 821 9710
rect 831 9706 835 9710
rect 836 9706 840 9710
rect 841 9706 845 9710
rect 846 9706 850 9710
rect 860 9706 864 9710
rect 865 9706 869 9710
rect 870 9706 874 9710
rect 875 9706 879 9710
rect 889 9706 893 9710
rect 894 9706 898 9710
rect 899 9706 903 9710
rect 904 9706 908 9710
rect 918 9706 922 9710
rect 923 9706 927 9710
rect 928 9706 932 9710
rect 933 9706 937 9710
rect 1319 9706 1323 9710
rect 1324 9706 1328 9710
rect 1329 9706 1333 9710
rect 1334 9706 1338 9710
rect 1628 9706 1632 9710
rect 1633 9706 1637 9710
rect 1638 9706 1642 9710
rect 1643 9706 1647 9710
rect 1937 9706 1941 9710
rect 1942 9706 1946 9710
rect 1947 9706 1951 9710
rect 1952 9706 1956 9710
rect 2246 9706 2250 9710
rect 2251 9706 2255 9710
rect 2256 9706 2260 9710
rect 2261 9706 2265 9710
rect 2555 9706 2559 9710
rect 2560 9706 2564 9710
rect 2565 9706 2569 9710
rect 2570 9706 2574 9710
rect 2864 9706 2868 9710
rect 2869 9706 2873 9710
rect 2874 9706 2878 9710
rect 2879 9706 2883 9710
rect 3173 9706 3177 9710
rect 3178 9706 3182 9710
rect 3183 9706 3187 9710
rect 3188 9706 3192 9710
rect 3482 9706 3486 9710
rect 3487 9706 3491 9710
rect 3492 9706 3496 9710
rect 3497 9706 3501 9710
rect 3791 9706 3795 9710
rect 3796 9706 3800 9710
rect 3801 9706 3805 9710
rect 3806 9706 3810 9710
rect 4100 9706 4104 9710
rect 4105 9706 4109 9710
rect 4110 9706 4114 9710
rect 4115 9706 4119 9710
rect 4292 9706 4296 9710
rect 4297 9706 4301 9710
rect 4302 9706 4306 9710
rect 4307 9706 4311 9710
rect 4318 9706 4322 9710
rect 4323 9706 4327 9710
rect 4328 9706 4332 9710
rect 4333 9706 4337 9710
rect 4344 9706 4348 9710
rect 4349 9706 4353 9710
rect 4354 9706 4358 9710
rect 4359 9706 4363 9710
rect 4370 9706 4374 9710
rect 4375 9706 4379 9710
rect 4380 9706 4384 9710
rect 4385 9706 4389 9710
rect 4396 9706 4400 9710
rect 4401 9706 4405 9710
rect 4406 9706 4410 9710
rect 4411 9706 4415 9710
rect 802 9696 806 9700
rect 807 9696 811 9700
rect 812 9696 816 9700
rect 817 9696 821 9700
rect 831 9696 835 9700
rect 836 9696 840 9700
rect 841 9696 845 9700
rect 846 9696 850 9700
rect 860 9696 864 9700
rect 865 9696 869 9700
rect 870 9696 874 9700
rect 875 9696 879 9700
rect 889 9696 893 9700
rect 894 9696 898 9700
rect 899 9696 903 9700
rect 904 9696 908 9700
rect 918 9696 922 9700
rect 923 9696 927 9700
rect 928 9696 932 9700
rect 933 9696 937 9700
rect 1319 9696 1323 9700
rect 1324 9696 1328 9700
rect 1329 9696 1333 9700
rect 1334 9696 1338 9700
rect 1628 9696 1632 9700
rect 1633 9696 1637 9700
rect 1638 9696 1642 9700
rect 1643 9696 1647 9700
rect 1937 9696 1941 9700
rect 1942 9696 1946 9700
rect 1947 9696 1951 9700
rect 1952 9696 1956 9700
rect 2246 9696 2250 9700
rect 2251 9696 2255 9700
rect 2256 9696 2260 9700
rect 2261 9696 2265 9700
rect 2555 9696 2559 9700
rect 2560 9696 2564 9700
rect 2565 9696 2569 9700
rect 2570 9696 2574 9700
rect 2864 9696 2868 9700
rect 2869 9696 2873 9700
rect 2874 9696 2878 9700
rect 2879 9696 2883 9700
rect 3173 9696 3177 9700
rect 3178 9696 3182 9700
rect 3183 9696 3187 9700
rect 3188 9696 3192 9700
rect 3482 9696 3486 9700
rect 3487 9696 3491 9700
rect 3492 9696 3496 9700
rect 3497 9696 3501 9700
rect 3791 9696 3795 9700
rect 3796 9696 3800 9700
rect 3801 9696 3805 9700
rect 3806 9696 3810 9700
rect 4100 9696 4104 9700
rect 4105 9696 4109 9700
rect 4110 9696 4114 9700
rect 4115 9696 4119 9700
rect 4292 9696 4296 9700
rect 4297 9696 4301 9700
rect 4302 9696 4306 9700
rect 4307 9696 4311 9700
rect 4318 9696 4322 9700
rect 4323 9696 4327 9700
rect 4328 9696 4332 9700
rect 4333 9696 4337 9700
rect 4344 9696 4348 9700
rect 4349 9696 4353 9700
rect 4354 9696 4358 9700
rect 4359 9696 4363 9700
rect 4370 9696 4374 9700
rect 4375 9696 4379 9700
rect 4380 9696 4384 9700
rect 4385 9696 4389 9700
rect 4396 9696 4400 9700
rect 4401 9696 4405 9700
rect 4406 9696 4410 9700
rect 4411 9696 4415 9700
rect 802 9686 806 9690
rect 807 9686 811 9690
rect 812 9686 816 9690
rect 817 9686 821 9690
rect 831 9686 835 9690
rect 836 9686 840 9690
rect 841 9686 845 9690
rect 846 9686 850 9690
rect 860 9686 864 9690
rect 865 9686 869 9690
rect 870 9686 874 9690
rect 875 9686 879 9690
rect 889 9686 893 9690
rect 894 9686 898 9690
rect 899 9686 903 9690
rect 904 9686 908 9690
rect 918 9686 922 9690
rect 923 9686 927 9690
rect 928 9686 932 9690
rect 933 9686 937 9690
rect 1319 9686 1323 9690
rect 1324 9686 1328 9690
rect 1329 9686 1333 9690
rect 1334 9686 1338 9690
rect 1628 9686 1632 9690
rect 1633 9686 1637 9690
rect 1638 9686 1642 9690
rect 1643 9686 1647 9690
rect 1937 9686 1941 9690
rect 1942 9686 1946 9690
rect 1947 9686 1951 9690
rect 1952 9686 1956 9690
rect 2246 9686 2250 9690
rect 2251 9686 2255 9690
rect 2256 9686 2260 9690
rect 2261 9686 2265 9690
rect 2555 9686 2559 9690
rect 2560 9686 2564 9690
rect 2565 9686 2569 9690
rect 2570 9686 2574 9690
rect 2864 9686 2868 9690
rect 2869 9686 2873 9690
rect 2874 9686 2878 9690
rect 2879 9686 2883 9690
rect 3173 9686 3177 9690
rect 3178 9686 3182 9690
rect 3183 9686 3187 9690
rect 3188 9686 3192 9690
rect 3482 9686 3486 9690
rect 3487 9686 3491 9690
rect 3492 9686 3496 9690
rect 3497 9686 3501 9690
rect 3791 9686 3795 9690
rect 3796 9686 3800 9690
rect 3801 9686 3805 9690
rect 3806 9686 3810 9690
rect 4100 9686 4104 9690
rect 4105 9686 4109 9690
rect 4110 9686 4114 9690
rect 4115 9686 4119 9690
rect 4292 9686 4296 9690
rect 4297 9686 4301 9690
rect 4302 9686 4306 9690
rect 4307 9686 4311 9690
rect 4318 9686 4322 9690
rect 4323 9686 4327 9690
rect 4328 9686 4332 9690
rect 4333 9686 4337 9690
rect 4344 9686 4348 9690
rect 4349 9686 4353 9690
rect 4354 9686 4358 9690
rect 4359 9686 4363 9690
rect 4370 9686 4374 9690
rect 4375 9686 4379 9690
rect 4380 9686 4384 9690
rect 4385 9686 4389 9690
rect 4396 9686 4400 9690
rect 4401 9686 4405 9690
rect 4406 9686 4410 9690
rect 4411 9686 4415 9690
rect 659 9618 663 9622
rect 669 9618 673 9622
rect 679 9618 683 9622
rect 689 9618 693 9622
rect 659 9613 663 9617
rect 669 9613 673 9617
rect 679 9613 683 9617
rect 689 9613 693 9617
rect 659 9608 663 9612
rect 669 9608 673 9612
rect 679 9608 683 9612
rect 689 9608 693 9612
rect 659 9603 663 9607
rect 669 9603 673 9607
rect 679 9603 683 9607
rect 689 9603 693 9607
rect 659 9592 663 9596
rect 669 9592 673 9596
rect 679 9592 683 9596
rect 689 9592 693 9596
rect 659 9587 663 9591
rect 669 9587 673 9591
rect 679 9587 683 9591
rect 689 9587 693 9591
rect 659 9582 663 9586
rect 669 9582 673 9586
rect 679 9582 683 9586
rect 689 9582 693 9586
rect 659 9577 663 9581
rect 669 9577 673 9581
rect 679 9577 683 9581
rect 689 9577 693 9581
rect 659 9566 663 9570
rect 669 9566 673 9570
rect 679 9566 683 9570
rect 689 9566 693 9570
rect 659 9561 663 9565
rect 669 9561 673 9565
rect 679 9561 683 9565
rect 689 9561 693 9565
rect 659 9556 663 9560
rect 669 9556 673 9560
rect 679 9556 683 9560
rect 689 9556 693 9560
rect 659 9551 663 9555
rect 669 9551 673 9555
rect 679 9551 683 9555
rect 689 9551 693 9555
rect 659 9540 663 9544
rect 669 9540 673 9544
rect 679 9540 683 9544
rect 689 9540 693 9544
rect 659 9535 663 9539
rect 669 9535 673 9539
rect 679 9535 683 9539
rect 689 9535 693 9539
rect 659 9530 663 9534
rect 669 9530 673 9534
rect 679 9530 683 9534
rect 689 9530 693 9534
rect 659 9525 663 9529
rect 669 9525 673 9529
rect 679 9525 683 9529
rect 689 9525 693 9529
rect 659 9514 663 9518
rect 669 9514 673 9518
rect 679 9514 683 9518
rect 689 9514 693 9518
rect 659 9509 663 9513
rect 669 9509 673 9513
rect 679 9509 683 9513
rect 689 9509 693 9513
rect 659 9504 663 9508
rect 669 9504 673 9508
rect 679 9504 683 9508
rect 689 9504 693 9508
rect 659 9499 663 9503
rect 669 9499 673 9503
rect 679 9499 683 9503
rect 689 9499 693 9503
rect 4479 9573 4483 9577
rect 4489 9573 4493 9577
rect 4499 9573 4503 9577
rect 4509 9573 4513 9577
rect 4479 9568 4483 9572
rect 4489 9568 4493 9572
rect 4499 9568 4503 9572
rect 4509 9568 4513 9572
rect 4479 9563 4483 9567
rect 4489 9563 4493 9567
rect 4499 9563 4503 9567
rect 4509 9563 4513 9567
rect 4479 9558 4483 9562
rect 4489 9558 4493 9562
rect 4499 9558 4503 9562
rect 4509 9558 4513 9562
rect 4479 9544 4483 9548
rect 4489 9544 4493 9548
rect 4499 9544 4503 9548
rect 4509 9544 4513 9548
rect 4479 9539 4483 9543
rect 4489 9539 4493 9543
rect 4499 9539 4503 9543
rect 4509 9539 4513 9543
rect 4479 9534 4483 9538
rect 4489 9534 4493 9538
rect 4499 9534 4503 9538
rect 4509 9534 4513 9538
rect 4479 9529 4483 9533
rect 4489 9529 4493 9533
rect 4499 9529 4503 9533
rect 4509 9529 4513 9533
rect 4479 9515 4483 9519
rect 4489 9515 4493 9519
rect 4499 9515 4503 9519
rect 4509 9515 4513 9519
rect 4479 9510 4483 9514
rect 4489 9510 4493 9514
rect 4499 9510 4503 9514
rect 4509 9510 4513 9514
rect 4479 9505 4483 9509
rect 4489 9505 4493 9509
rect 4499 9505 4503 9509
rect 4509 9505 4513 9509
rect 4479 9500 4483 9504
rect 4489 9500 4493 9504
rect 4499 9500 4503 9504
rect 4509 9500 4513 9504
rect 4479 9486 4483 9490
rect 4489 9486 4493 9490
rect 4499 9486 4503 9490
rect 4509 9486 4513 9490
rect 4479 9481 4483 9485
rect 4489 9481 4493 9485
rect 4499 9481 4503 9485
rect 4509 9481 4513 9485
rect 4479 9476 4483 9480
rect 4489 9476 4493 9480
rect 4499 9476 4503 9480
rect 4509 9476 4513 9480
rect 4479 9471 4483 9475
rect 4489 9471 4493 9475
rect 4499 9471 4503 9475
rect 4509 9471 4513 9475
rect 4479 9457 4483 9461
rect 4489 9457 4493 9461
rect 4499 9457 4503 9461
rect 4509 9457 4513 9461
rect 4479 9452 4483 9456
rect 4489 9452 4493 9456
rect 4499 9452 4503 9456
rect 4509 9452 4513 9456
rect 4479 9447 4483 9451
rect 4489 9447 4493 9451
rect 4499 9447 4503 9451
rect 4509 9447 4513 9451
rect 4479 9442 4483 9446
rect 4489 9442 4493 9446
rect 4499 9442 4503 9446
rect 4509 9442 4513 9446
rect 659 9321 663 9325
rect 669 9321 673 9325
rect 679 9321 683 9325
rect 689 9321 693 9325
rect 659 9316 663 9320
rect 669 9316 673 9320
rect 679 9316 683 9320
rect 689 9316 693 9320
rect 659 9311 663 9315
rect 669 9311 673 9315
rect 679 9311 683 9315
rect 689 9311 693 9315
rect 659 9306 663 9310
rect 669 9306 673 9310
rect 679 9306 683 9310
rect 689 9306 693 9310
rect 2881 9283 2885 9287
rect 2909 9283 2913 9287
rect 2939 9283 2943 9287
rect 3013 9283 3017 9287
rect 3041 9283 3045 9287
rect 3071 9283 3075 9287
rect 3145 9283 3149 9287
rect 3173 9283 3177 9287
rect 3203 9283 3207 9287
rect 3277 9283 3281 9287
rect 3305 9283 3309 9287
rect 3335 9283 3339 9287
rect 3826 9283 3830 9287
rect 3854 9283 3858 9287
rect 3884 9283 3888 9287
rect 3958 9283 3962 9287
rect 3986 9283 3990 9287
rect 4016 9283 4020 9287
rect 4090 9283 4094 9287
rect 4118 9283 4122 9287
rect 4148 9283 4152 9287
rect 4222 9283 4226 9287
rect 4250 9283 4254 9287
rect 4280 9283 4284 9287
rect 2529 9250 2533 9254
rect 2557 9250 2561 9254
rect 2587 9250 2591 9254
rect 3474 9250 3478 9254
rect 3502 9250 3506 9254
rect 3532 9250 3536 9254
rect 2862 9197 2866 9201
rect 2897 9197 2901 9201
rect 3023 9197 3027 9201
rect 3047 9197 3051 9201
rect 3101 9197 3108 9201
rect 3128 9197 3132 9201
rect 3182 9197 3186 9201
rect 3807 9197 3811 9201
rect 3842 9197 3846 9201
rect 3968 9197 3972 9201
rect 3992 9197 3996 9201
rect 4046 9197 4053 9201
rect 4073 9197 4077 9201
rect 4127 9197 4131 9201
rect 2526 9148 2530 9152
rect 2556 9148 2560 9152
rect 2584 9148 2588 9152
rect 3471 9148 3475 9152
rect 3501 9148 3505 9152
rect 3529 9148 3533 9152
rect 2862 9065 2866 9069
rect 2897 9065 2901 9069
rect 3023 9065 3027 9069
rect 3047 9065 3051 9069
rect 3101 9065 3105 9069
rect 3128 9065 3132 9069
rect 3152 9065 3156 9069
rect 3807 9065 3811 9069
rect 3842 9065 3846 9069
rect 3968 9065 3972 9069
rect 3992 9065 3996 9069
rect 4046 9065 4050 9069
rect 4073 9065 4077 9069
rect 4097 9065 4101 9069
rect 4479 9056 4483 9060
rect 4489 9056 4493 9060
rect 4499 9056 4503 9060
rect 4509 9056 4513 9060
rect 4479 9051 4483 9055
rect 4489 9051 4493 9055
rect 4499 9051 4503 9055
rect 4509 9051 4513 9055
rect 4479 9046 4483 9050
rect 4489 9046 4493 9050
rect 4499 9046 4503 9050
rect 4509 9046 4513 9050
rect 4479 9041 4483 9045
rect 4489 9041 4493 9045
rect 4499 9041 4503 9045
rect 4509 9041 4513 9045
rect 3359 9022 3363 9026
rect 3383 9022 3387 9026
rect 3437 9022 3441 9026
rect 3580 9022 3584 9026
rect 659 9012 663 9016
rect 669 9012 673 9016
rect 679 9012 683 9016
rect 689 9012 693 9016
rect 659 9007 663 9011
rect 669 9007 673 9011
rect 679 9007 683 9011
rect 689 9007 693 9011
rect 659 9002 663 9006
rect 669 9002 673 9006
rect 679 9002 683 9006
rect 689 9002 693 9006
rect 659 8997 663 9001
rect 669 8997 673 9001
rect 679 8997 683 9001
rect 689 8997 693 9001
rect 2862 8933 2866 8937
rect 2897 8933 2901 8937
rect 3023 8933 3027 8937
rect 3047 8933 3051 8937
rect 3101 8933 3108 8937
rect 3128 8933 3132 8937
rect 3182 8933 3186 8937
rect 3218 8933 3222 8937
rect 3272 8933 3276 8937
rect 3807 8933 3811 8937
rect 3842 8933 3846 8937
rect 3968 8933 3972 8937
rect 3992 8933 3996 8937
rect 4046 8933 4053 8937
rect 4073 8933 4077 8937
rect 4127 8933 4131 8937
rect 4163 8933 4167 8937
rect 4217 8933 4221 8937
rect 3337 8892 3341 8896
rect 3359 8892 3363 8896
rect 3383 8892 3387 8896
rect 3437 8892 3441 8896
rect 3486 8892 3490 8896
rect 2862 8801 2866 8805
rect 2897 8801 2901 8805
rect 3023 8801 3027 8805
rect 3047 8801 3051 8805
rect 3158 8801 3162 8805
rect 3807 8801 3811 8805
rect 3842 8801 3846 8805
rect 3968 8801 3972 8805
rect 3992 8801 3996 8805
rect 4103 8801 4107 8805
rect 2397 8748 2401 8752
rect 2425 8748 2429 8752
rect 2455 8748 2459 8752
rect 2529 8748 2533 8752
rect 2557 8748 2561 8752
rect 2587 8748 2591 8752
rect 2661 8748 2665 8752
rect 2689 8748 2693 8752
rect 2719 8748 2723 8752
rect 3342 8748 3346 8752
rect 3370 8748 3374 8752
rect 3400 8748 3404 8752
rect 3474 8748 3478 8752
rect 3502 8748 3506 8752
rect 3532 8748 3536 8752
rect 3606 8748 3610 8752
rect 3634 8748 3638 8752
rect 3664 8748 3668 8752
rect 4479 8747 4483 8751
rect 4489 8747 4493 8751
rect 4499 8747 4503 8751
rect 4509 8747 4513 8751
rect 4479 8742 4483 8746
rect 4489 8742 4493 8746
rect 4499 8742 4503 8746
rect 4509 8742 4513 8746
rect 4479 8737 4483 8741
rect 4489 8737 4493 8741
rect 4499 8737 4503 8741
rect 4509 8737 4513 8741
rect 4479 8732 4483 8736
rect 4489 8732 4493 8736
rect 4499 8732 4503 8736
rect 4509 8732 4513 8736
rect 659 8703 663 8707
rect 669 8703 673 8707
rect 679 8703 683 8707
rect 689 8703 693 8707
rect 659 8698 663 8702
rect 669 8698 673 8702
rect 679 8698 683 8702
rect 689 8698 693 8702
rect 659 8693 663 8697
rect 669 8693 673 8697
rect 679 8693 683 8697
rect 689 8693 693 8697
rect 659 8688 663 8692
rect 669 8688 673 8692
rect 679 8688 683 8692
rect 689 8688 693 8692
rect 3180 8636 3184 8640
rect 3208 8636 3212 8640
rect 3238 8636 3242 8640
rect 4125 8636 4129 8640
rect 4153 8636 4157 8640
rect 4183 8636 4187 8640
rect 2397 8606 2401 8610
rect 2425 8606 2429 8610
rect 2455 8606 2459 8610
rect 2529 8606 2533 8610
rect 2557 8606 2561 8610
rect 2587 8606 2591 8610
rect 2661 8606 2665 8610
rect 2689 8606 2693 8610
rect 2719 8606 2723 8610
rect 3342 8606 3346 8610
rect 3370 8606 3374 8610
rect 3400 8606 3404 8610
rect 3474 8606 3478 8610
rect 3502 8606 3506 8610
rect 3532 8606 3536 8610
rect 3606 8606 3610 8610
rect 3634 8606 3638 8610
rect 3664 8606 3668 8610
rect 3180 8550 3184 8554
rect 3208 8550 3212 8554
rect 3238 8550 3242 8554
rect 4125 8550 4129 8554
rect 4153 8550 4157 8554
rect 4183 8550 4187 8554
rect 2397 8520 2401 8524
rect 2425 8520 2429 8524
rect 2455 8520 2459 8524
rect 2529 8520 2533 8524
rect 2557 8520 2561 8524
rect 2587 8520 2591 8524
rect 2661 8520 2665 8524
rect 2689 8520 2693 8524
rect 2719 8520 2723 8524
rect 3342 8520 3346 8524
rect 3370 8520 3374 8524
rect 3400 8520 3404 8524
rect 3474 8520 3478 8524
rect 3502 8520 3506 8524
rect 3532 8520 3536 8524
rect 3606 8520 3610 8524
rect 3634 8520 3638 8524
rect 3664 8520 3668 8524
rect 4479 8438 4483 8442
rect 4489 8438 4493 8442
rect 4499 8438 4503 8442
rect 4509 8438 4513 8442
rect 4479 8433 4483 8437
rect 4489 8433 4493 8437
rect 4499 8433 4503 8437
rect 4509 8433 4513 8437
rect 4479 8428 4483 8432
rect 4489 8428 4493 8432
rect 4499 8428 4503 8432
rect 4509 8428 4513 8432
rect 4479 8423 4483 8427
rect 4489 8423 4493 8427
rect 4499 8423 4503 8427
rect 4509 8423 4513 8427
rect 659 8394 663 8398
rect 669 8394 673 8398
rect 679 8394 683 8398
rect 689 8394 693 8398
rect 659 8389 663 8393
rect 669 8389 673 8393
rect 679 8389 683 8393
rect 689 8389 693 8393
rect 659 8384 663 8388
rect 669 8384 673 8388
rect 679 8384 683 8388
rect 689 8384 693 8388
rect 659 8379 663 8383
rect 669 8379 673 8383
rect 679 8379 683 8383
rect 689 8379 693 8383
rect 2397 8380 2401 8384
rect 2425 8380 2429 8384
rect 2455 8380 2459 8384
rect 2529 8380 2533 8384
rect 2557 8380 2561 8384
rect 2587 8380 2591 8384
rect 2661 8380 2665 8384
rect 2689 8380 2693 8384
rect 2719 8380 2723 8384
rect 3342 8380 3346 8384
rect 3370 8380 3374 8384
rect 3400 8380 3404 8384
rect 3474 8380 3478 8384
rect 3502 8380 3506 8384
rect 3532 8380 3536 8384
rect 3606 8380 3610 8384
rect 3634 8380 3638 8384
rect 3664 8380 3668 8384
rect 2881 8301 2885 8305
rect 2909 8301 2913 8305
rect 2939 8301 2943 8305
rect 3013 8301 3017 8305
rect 3041 8301 3045 8305
rect 3071 8301 3075 8305
rect 3145 8301 3149 8305
rect 3173 8301 3177 8305
rect 3203 8301 3207 8305
rect 3277 8301 3281 8305
rect 3305 8301 3309 8305
rect 3335 8301 3339 8305
rect 3826 8301 3830 8305
rect 3854 8301 3858 8305
rect 3884 8301 3888 8305
rect 3958 8301 3962 8305
rect 3986 8301 3990 8305
rect 4016 8301 4020 8305
rect 4090 8301 4094 8305
rect 4118 8301 4122 8305
rect 4148 8301 4152 8305
rect 4222 8301 4226 8305
rect 4250 8301 4254 8305
rect 4280 8301 4284 8305
rect 2529 8268 2533 8272
rect 2557 8268 2561 8272
rect 2587 8268 2591 8272
rect 3474 8268 3478 8272
rect 3502 8268 3506 8272
rect 3532 8268 3536 8272
rect 2862 8215 2866 8219
rect 2897 8215 2901 8219
rect 3023 8215 3027 8219
rect 3047 8215 3051 8219
rect 3101 8215 3108 8219
rect 3128 8215 3132 8219
rect 3182 8215 3186 8219
rect 3807 8215 3811 8219
rect 3842 8215 3846 8219
rect 3968 8215 3972 8219
rect 3992 8215 3996 8219
rect 4046 8215 4053 8219
rect 4073 8215 4077 8219
rect 4127 8215 4131 8219
rect 2526 8166 2530 8170
rect 2556 8166 2560 8170
rect 2584 8166 2588 8170
rect 3471 8166 3475 8170
rect 3501 8166 3505 8170
rect 3529 8166 3533 8170
rect 4479 8129 4483 8133
rect 4489 8129 4493 8133
rect 4499 8129 4503 8133
rect 4509 8129 4513 8133
rect 4479 8124 4483 8128
rect 4489 8124 4493 8128
rect 4499 8124 4503 8128
rect 4509 8124 4513 8128
rect 4479 8119 4483 8123
rect 4489 8119 4493 8123
rect 4499 8119 4503 8123
rect 4509 8119 4513 8123
rect 4479 8114 4483 8118
rect 4489 8114 4493 8118
rect 4499 8114 4503 8118
rect 4509 8114 4513 8118
rect 4479 8098 4483 8102
rect 4489 8098 4493 8102
rect 4499 8098 4503 8102
rect 4509 8098 4513 8102
rect 659 8085 663 8089
rect 669 8085 673 8089
rect 679 8085 683 8089
rect 689 8085 693 8089
rect 4479 8093 4483 8097
rect 4489 8093 4493 8097
rect 4499 8093 4503 8097
rect 4509 8093 4513 8097
rect 4479 8088 4483 8092
rect 4489 8088 4493 8092
rect 4499 8088 4503 8092
rect 4509 8088 4513 8092
rect 659 8080 663 8084
rect 669 8080 673 8084
rect 679 8080 683 8084
rect 689 8080 693 8084
rect 2862 8083 2866 8087
rect 2897 8083 2901 8087
rect 3023 8083 3027 8087
rect 3047 8083 3051 8087
rect 3101 8083 3105 8087
rect 3128 8083 3132 8087
rect 3152 8083 3156 8087
rect 3807 8083 3811 8087
rect 3842 8083 3846 8087
rect 3968 8083 3972 8087
rect 3992 8083 3996 8087
rect 4046 8083 4050 8087
rect 4073 8083 4077 8087
rect 4097 8083 4101 8087
rect 4479 8083 4483 8087
rect 4489 8083 4493 8087
rect 4499 8083 4503 8087
rect 4509 8083 4513 8087
rect 659 8075 663 8079
rect 669 8075 673 8079
rect 679 8075 683 8079
rect 689 8075 693 8079
rect 659 8070 663 8074
rect 669 8070 673 8074
rect 679 8070 683 8074
rect 689 8070 693 8074
rect 2862 7951 2866 7955
rect 2897 7951 2901 7955
rect 3023 7951 3027 7955
rect 3047 7951 3051 7955
rect 3101 7951 3108 7955
rect 3128 7951 3132 7955
rect 3182 7951 3186 7955
rect 3218 7951 3222 7955
rect 3272 7951 3276 7955
rect 3807 7951 3811 7955
rect 3842 7951 3846 7955
rect 3968 7951 3972 7955
rect 3992 7951 3996 7955
rect 4046 7951 4053 7955
rect 4073 7951 4077 7955
rect 4127 7951 4131 7955
rect 4163 7951 4167 7955
rect 4217 7951 4221 7955
rect 2862 7819 2866 7823
rect 2897 7819 2901 7823
rect 3023 7819 3027 7823
rect 3047 7819 3051 7823
rect 3158 7819 3162 7823
rect 3807 7819 3811 7823
rect 3842 7819 3846 7823
rect 3968 7819 3972 7823
rect 3992 7819 3996 7823
rect 4103 7819 4107 7823
rect 659 7776 663 7780
rect 669 7776 673 7780
rect 679 7776 683 7780
rect 689 7776 693 7780
rect 659 7771 663 7775
rect 669 7771 673 7775
rect 679 7771 683 7775
rect 689 7771 693 7775
rect 659 7766 663 7770
rect 669 7766 673 7770
rect 679 7766 683 7770
rect 689 7766 693 7770
rect 2397 7766 2401 7770
rect 2425 7766 2429 7770
rect 2455 7766 2459 7770
rect 2529 7766 2533 7770
rect 2557 7766 2561 7770
rect 2587 7766 2591 7770
rect 2661 7766 2665 7770
rect 2689 7766 2693 7770
rect 2719 7766 2723 7770
rect 659 7761 663 7765
rect 669 7761 673 7765
rect 679 7761 683 7765
rect 689 7761 693 7765
rect 4479 7789 4483 7793
rect 4489 7789 4493 7793
rect 4499 7789 4503 7793
rect 4509 7789 4513 7793
rect 4479 7784 4483 7788
rect 4489 7784 4493 7788
rect 4499 7784 4503 7788
rect 4509 7784 4513 7788
rect 3342 7766 3346 7770
rect 3370 7766 3374 7770
rect 3400 7766 3404 7770
rect 3474 7766 3478 7770
rect 3502 7766 3506 7770
rect 3532 7766 3536 7770
rect 3606 7766 3610 7770
rect 3634 7766 3638 7770
rect 3664 7766 3668 7770
rect 4479 7779 4483 7783
rect 4489 7779 4493 7783
rect 4499 7779 4503 7783
rect 4509 7779 4513 7783
rect 4479 7774 4483 7778
rect 4489 7774 4493 7778
rect 4499 7774 4503 7778
rect 4509 7774 4513 7778
rect 3180 7654 3184 7658
rect 3208 7654 3212 7658
rect 3238 7654 3242 7658
rect 4125 7654 4129 7658
rect 4153 7654 4157 7658
rect 4183 7654 4187 7658
rect 2397 7624 2401 7628
rect 2425 7624 2429 7628
rect 2455 7624 2459 7628
rect 2529 7624 2533 7628
rect 2557 7624 2561 7628
rect 2587 7624 2591 7628
rect 2661 7624 2665 7628
rect 2689 7624 2693 7628
rect 2719 7624 2723 7628
rect 3342 7624 3346 7628
rect 3370 7624 3374 7628
rect 3400 7624 3404 7628
rect 3474 7624 3478 7628
rect 3502 7624 3506 7628
rect 3532 7624 3536 7628
rect 3606 7624 3610 7628
rect 3634 7624 3638 7628
rect 3664 7624 3668 7628
rect 3180 7568 3184 7572
rect 3208 7568 3212 7572
rect 3238 7568 3242 7572
rect 4125 7568 4129 7572
rect 4153 7568 4157 7572
rect 4183 7568 4187 7572
rect 2397 7538 2401 7542
rect 2425 7538 2429 7542
rect 2455 7538 2459 7542
rect 2529 7538 2533 7542
rect 2557 7538 2561 7542
rect 2587 7538 2591 7542
rect 2661 7538 2665 7542
rect 2689 7538 2693 7542
rect 2719 7538 2723 7542
rect 3342 7538 3346 7542
rect 3370 7538 3374 7542
rect 3400 7538 3404 7542
rect 3474 7538 3478 7542
rect 3502 7538 3506 7542
rect 3532 7538 3536 7542
rect 3606 7538 3610 7542
rect 3634 7538 3638 7542
rect 3664 7538 3668 7542
rect 659 7467 663 7471
rect 669 7467 673 7471
rect 679 7467 683 7471
rect 689 7467 693 7471
rect 659 7462 663 7466
rect 669 7462 673 7466
rect 679 7462 683 7466
rect 689 7462 693 7466
rect 659 7457 663 7461
rect 669 7457 673 7461
rect 679 7457 683 7461
rect 689 7457 693 7461
rect 659 7452 663 7456
rect 669 7452 673 7456
rect 679 7452 683 7456
rect 689 7452 693 7456
rect 2397 7398 2401 7402
rect 2425 7398 2429 7402
rect 2455 7398 2459 7402
rect 2529 7398 2533 7402
rect 2557 7398 2561 7402
rect 2587 7398 2591 7402
rect 2661 7398 2665 7402
rect 2689 7398 2693 7402
rect 2719 7398 2723 7402
rect 3342 7398 3346 7402
rect 3370 7398 3374 7402
rect 3400 7398 3404 7402
rect 3474 7398 3478 7402
rect 3502 7398 3506 7402
rect 3532 7398 3536 7402
rect 3606 7398 3610 7402
rect 3634 7398 3638 7402
rect 3664 7398 3668 7402
rect 659 7158 663 7162
rect 669 7158 673 7162
rect 679 7158 683 7162
rect 689 7158 693 7162
rect 659 7153 663 7157
rect 669 7153 673 7157
rect 679 7153 683 7157
rect 689 7153 693 7157
rect 659 7148 663 7152
rect 669 7148 673 7152
rect 679 7148 683 7152
rect 689 7148 693 7152
rect 659 7143 663 7147
rect 669 7143 673 7147
rect 679 7143 683 7147
rect 689 7143 693 7147
rect 659 6849 663 6853
rect 669 6849 673 6853
rect 679 6849 683 6853
rect 689 6849 693 6853
rect 659 6844 663 6848
rect 669 6844 673 6848
rect 679 6844 683 6848
rect 689 6844 693 6848
rect 659 6839 663 6843
rect 669 6839 673 6843
rect 679 6839 683 6843
rect 689 6839 693 6843
rect 659 6834 663 6838
rect 669 6834 673 6838
rect 679 6834 683 6838
rect 689 6834 693 6838
rect 659 6540 663 6544
rect 669 6540 673 6544
rect 679 6540 683 6544
rect 689 6540 693 6544
rect 659 6535 663 6539
rect 669 6535 673 6539
rect 679 6535 683 6539
rect 689 6535 693 6539
rect 659 6530 663 6534
rect 669 6530 673 6534
rect 679 6530 683 6534
rect 689 6530 693 6534
rect 659 6525 663 6529
rect 669 6525 673 6529
rect 679 6525 683 6529
rect 689 6525 693 6529
rect 659 6140 663 6144
rect 669 6140 673 6144
rect 679 6140 683 6144
rect 689 6140 693 6144
rect 659 6135 663 6139
rect 669 6135 673 6139
rect 679 6135 683 6139
rect 689 6135 693 6139
rect 659 6130 663 6134
rect 669 6130 673 6134
rect 679 6130 683 6134
rect 689 6130 693 6134
rect 659 6125 663 6129
rect 669 6125 673 6129
rect 679 6125 683 6129
rect 689 6125 693 6129
rect 659 6111 663 6115
rect 669 6111 673 6115
rect 679 6111 683 6115
rect 689 6111 693 6115
rect 659 6106 663 6110
rect 669 6106 673 6110
rect 679 6106 683 6110
rect 689 6106 693 6110
rect 659 6101 663 6105
rect 669 6101 673 6105
rect 679 6101 683 6105
rect 689 6101 693 6105
rect 659 6096 663 6100
rect 669 6096 673 6100
rect 679 6096 683 6100
rect 689 6096 693 6100
rect 659 6082 663 6086
rect 669 6082 673 6086
rect 679 6082 683 6086
rect 689 6082 693 6086
rect 659 6077 663 6081
rect 669 6077 673 6081
rect 679 6077 683 6081
rect 689 6077 693 6081
rect 659 6072 663 6076
rect 669 6072 673 6076
rect 679 6072 683 6076
rect 689 6072 693 6076
rect 659 6067 663 6071
rect 669 6067 673 6071
rect 679 6067 683 6071
rect 689 6067 693 6071
rect 659 6053 663 6057
rect 669 6053 673 6057
rect 679 6053 683 6057
rect 689 6053 693 6057
rect 659 6048 663 6052
rect 669 6048 673 6052
rect 679 6048 683 6052
rect 689 6048 693 6052
rect 659 6043 663 6047
rect 669 6043 673 6047
rect 679 6043 683 6047
rect 689 6043 693 6047
rect 659 6038 663 6042
rect 669 6038 673 6042
rect 679 6038 683 6042
rect 689 6038 693 6042
rect 659 6024 663 6028
rect 669 6024 673 6028
rect 679 6024 683 6028
rect 689 6024 693 6028
rect 659 6019 663 6023
rect 669 6019 673 6023
rect 679 6019 683 6023
rect 689 6019 693 6023
rect 659 6014 663 6018
rect 669 6014 673 6018
rect 679 6014 683 6018
rect 689 6014 693 6018
rect 659 6009 663 6013
rect 669 6009 673 6013
rect 679 6009 683 6013
rect 689 6009 693 6013
rect 4479 7202 4483 7206
rect 4489 7202 4493 7206
rect 4499 7202 4503 7206
rect 4509 7202 4513 7206
rect 4479 7197 4483 7201
rect 4489 7197 4493 7201
rect 4499 7197 4503 7201
rect 4509 7197 4513 7201
rect 4479 7192 4483 7196
rect 4489 7192 4493 7196
rect 4499 7192 4503 7196
rect 4509 7192 4513 7196
rect 4479 7187 4483 7191
rect 4489 7187 4493 7191
rect 4499 7187 4503 7191
rect 4509 7187 4513 7191
rect 4479 6893 4483 6897
rect 4489 6893 4493 6897
rect 4499 6893 4503 6897
rect 4509 6893 4513 6897
rect 4479 6888 4483 6892
rect 4489 6888 4493 6892
rect 4499 6888 4503 6892
rect 4509 6888 4513 6892
rect 4479 6883 4483 6887
rect 4489 6883 4493 6887
rect 4499 6883 4503 6887
rect 4509 6883 4513 6887
rect 4479 6878 4483 6882
rect 4489 6878 4493 6882
rect 4499 6878 4503 6882
rect 4509 6878 4513 6882
rect 4479 6584 4483 6588
rect 4489 6584 4493 6588
rect 4499 6584 4503 6588
rect 4509 6584 4513 6588
rect 4479 6579 4483 6583
rect 4489 6579 4493 6583
rect 4499 6579 4503 6583
rect 4509 6579 4513 6583
rect 4479 6574 4483 6578
rect 4489 6574 4493 6578
rect 4499 6574 4503 6578
rect 4509 6574 4513 6578
rect 4479 6569 4483 6573
rect 4489 6569 4493 6573
rect 4499 6569 4503 6573
rect 4509 6569 4513 6573
rect 4479 6275 4483 6279
rect 4489 6275 4493 6279
rect 4499 6275 4503 6279
rect 4509 6275 4513 6279
rect 4479 6270 4483 6274
rect 4489 6270 4493 6274
rect 4499 6270 4503 6274
rect 4509 6270 4513 6274
rect 4479 6265 4483 6269
rect 4489 6265 4493 6269
rect 4499 6265 4503 6269
rect 4509 6265 4513 6269
rect 4479 6260 4483 6264
rect 4489 6260 4493 6264
rect 4499 6260 4503 6264
rect 4509 6260 4513 6264
rect 4479 6083 4483 6087
rect 4489 6083 4493 6087
rect 4499 6083 4503 6087
rect 4509 6083 4513 6087
rect 4479 6078 4483 6082
rect 4489 6078 4493 6082
rect 4499 6078 4503 6082
rect 4509 6078 4513 6082
rect 4479 6073 4483 6077
rect 4489 6073 4493 6077
rect 4499 6073 4503 6077
rect 4509 6073 4513 6077
rect 4479 6068 4483 6072
rect 4489 6068 4493 6072
rect 4499 6068 4503 6072
rect 4509 6068 4513 6072
rect 4479 6057 4483 6061
rect 4489 6057 4493 6061
rect 4499 6057 4503 6061
rect 4509 6057 4513 6061
rect 4479 6052 4483 6056
rect 4489 6052 4493 6056
rect 4499 6052 4503 6056
rect 4509 6052 4513 6056
rect 4479 6047 4483 6051
rect 4489 6047 4493 6051
rect 4499 6047 4503 6051
rect 4509 6047 4513 6051
rect 4479 6042 4483 6046
rect 4489 6042 4493 6046
rect 4499 6042 4503 6046
rect 4509 6042 4513 6046
rect 4479 6031 4483 6035
rect 4489 6031 4493 6035
rect 4499 6031 4503 6035
rect 4509 6031 4513 6035
rect 4479 6026 4483 6030
rect 4489 6026 4493 6030
rect 4499 6026 4503 6030
rect 4509 6026 4513 6030
rect 4479 6021 4483 6025
rect 4489 6021 4493 6025
rect 4499 6021 4503 6025
rect 4509 6021 4513 6025
rect 4479 6016 4483 6020
rect 4489 6016 4493 6020
rect 4499 6016 4503 6020
rect 4509 6016 4513 6020
rect 4479 6005 4483 6009
rect 4489 6005 4493 6009
rect 4499 6005 4503 6009
rect 4509 6005 4513 6009
rect 4479 6000 4483 6004
rect 4489 6000 4493 6004
rect 4499 6000 4503 6004
rect 4509 6000 4513 6004
rect 4479 5995 4483 5999
rect 4489 5995 4493 5999
rect 4499 5995 4503 5999
rect 4509 5995 4513 5999
rect 4479 5990 4483 5994
rect 4489 5990 4493 5994
rect 4499 5990 4503 5994
rect 4509 5990 4513 5994
rect 4479 5979 4483 5983
rect 4489 5979 4493 5983
rect 4499 5979 4503 5983
rect 4509 5979 4513 5983
rect 4479 5974 4483 5978
rect 4489 5974 4493 5978
rect 4499 5974 4503 5978
rect 4509 5974 4513 5978
rect 4479 5969 4483 5973
rect 4489 5969 4493 5973
rect 4499 5969 4503 5973
rect 4509 5969 4513 5973
rect 4479 5964 4483 5968
rect 4489 5964 4493 5968
rect 4499 5964 4503 5968
rect 4509 5964 4513 5968
rect 757 5896 761 5900
rect 762 5896 766 5900
rect 767 5896 771 5900
rect 772 5896 776 5900
rect 783 5896 787 5900
rect 788 5896 792 5900
rect 793 5896 797 5900
rect 798 5896 802 5900
rect 809 5896 813 5900
rect 814 5896 818 5900
rect 819 5896 823 5900
rect 824 5896 828 5900
rect 835 5896 839 5900
rect 840 5896 844 5900
rect 845 5896 849 5900
rect 850 5896 854 5900
rect 861 5896 865 5900
rect 866 5896 870 5900
rect 871 5896 875 5900
rect 876 5896 880 5900
rect 1054 5896 1058 5900
rect 1059 5896 1063 5900
rect 1064 5896 1068 5900
rect 1069 5896 1073 5900
rect 1363 5896 1367 5900
rect 1368 5896 1372 5900
rect 1373 5896 1377 5900
rect 1378 5896 1382 5900
rect 1672 5896 1676 5900
rect 1677 5896 1681 5900
rect 1682 5896 1686 5900
rect 1687 5896 1691 5900
rect 1981 5896 1985 5900
rect 1986 5896 1990 5900
rect 1991 5896 1995 5900
rect 1996 5896 2000 5900
rect 2290 5896 2294 5900
rect 2295 5896 2299 5900
rect 2300 5896 2304 5900
rect 2305 5896 2309 5900
rect 2599 5896 2603 5900
rect 2604 5896 2608 5900
rect 2609 5896 2613 5900
rect 2614 5896 2618 5900
rect 2908 5896 2912 5900
rect 2913 5896 2917 5900
rect 2918 5896 2922 5900
rect 2923 5896 2927 5900
rect 3217 5896 3221 5900
rect 3222 5896 3226 5900
rect 3227 5896 3231 5900
rect 3232 5896 3236 5900
rect 3526 5896 3530 5900
rect 3531 5896 3535 5900
rect 3536 5896 3540 5900
rect 3541 5896 3545 5900
rect 3835 5896 3839 5900
rect 3840 5896 3844 5900
rect 3845 5896 3849 5900
rect 3850 5896 3854 5900
rect 4235 5896 4239 5900
rect 4240 5896 4244 5900
rect 4245 5896 4249 5900
rect 4250 5896 4254 5900
rect 4264 5896 4268 5900
rect 4269 5896 4273 5900
rect 4274 5896 4278 5900
rect 4279 5896 4283 5900
rect 4293 5896 4297 5900
rect 4298 5896 4302 5900
rect 4303 5896 4307 5900
rect 4308 5896 4312 5900
rect 4322 5896 4326 5900
rect 4327 5896 4331 5900
rect 4332 5896 4336 5900
rect 4337 5896 4341 5900
rect 4351 5896 4355 5900
rect 4356 5896 4360 5900
rect 4361 5896 4365 5900
rect 4366 5896 4370 5900
rect 757 5886 761 5890
rect 762 5886 766 5890
rect 767 5886 771 5890
rect 772 5886 776 5890
rect 783 5886 787 5890
rect 788 5886 792 5890
rect 793 5886 797 5890
rect 798 5886 802 5890
rect 809 5886 813 5890
rect 814 5886 818 5890
rect 819 5886 823 5890
rect 824 5886 828 5890
rect 835 5886 839 5890
rect 840 5886 844 5890
rect 845 5886 849 5890
rect 850 5886 854 5890
rect 861 5886 865 5890
rect 866 5886 870 5890
rect 871 5886 875 5890
rect 876 5886 880 5890
rect 1054 5886 1058 5890
rect 1059 5886 1063 5890
rect 1064 5886 1068 5890
rect 1069 5886 1073 5890
rect 1363 5886 1367 5890
rect 1368 5886 1372 5890
rect 1373 5886 1377 5890
rect 1378 5886 1382 5890
rect 1672 5886 1676 5890
rect 1677 5886 1681 5890
rect 1682 5886 1686 5890
rect 1687 5886 1691 5890
rect 1981 5886 1985 5890
rect 1986 5886 1990 5890
rect 1991 5886 1995 5890
rect 1996 5886 2000 5890
rect 2290 5886 2294 5890
rect 2295 5886 2299 5890
rect 2300 5886 2304 5890
rect 2305 5886 2309 5890
rect 2599 5886 2603 5890
rect 2604 5886 2608 5890
rect 2609 5886 2613 5890
rect 2614 5886 2618 5890
rect 2908 5886 2912 5890
rect 2913 5886 2917 5890
rect 2918 5886 2922 5890
rect 2923 5886 2927 5890
rect 3217 5886 3221 5890
rect 3222 5886 3226 5890
rect 3227 5886 3231 5890
rect 3232 5886 3236 5890
rect 3526 5886 3530 5890
rect 3531 5886 3535 5890
rect 3536 5886 3540 5890
rect 3541 5886 3545 5890
rect 3835 5886 3839 5890
rect 3840 5886 3844 5890
rect 3845 5886 3849 5890
rect 3850 5886 3854 5890
rect 4235 5886 4239 5890
rect 4240 5886 4244 5890
rect 4245 5886 4249 5890
rect 4250 5886 4254 5890
rect 4264 5886 4268 5890
rect 4269 5886 4273 5890
rect 4274 5886 4278 5890
rect 4279 5886 4283 5890
rect 4293 5886 4297 5890
rect 4298 5886 4302 5890
rect 4303 5886 4307 5890
rect 4308 5886 4312 5890
rect 4322 5886 4326 5890
rect 4327 5886 4331 5890
rect 4332 5886 4336 5890
rect 4337 5886 4341 5890
rect 4351 5886 4355 5890
rect 4356 5886 4360 5890
rect 4361 5886 4365 5890
rect 4366 5886 4370 5890
rect 757 5876 761 5880
rect 762 5876 766 5880
rect 767 5876 771 5880
rect 772 5876 776 5880
rect 783 5876 787 5880
rect 788 5876 792 5880
rect 793 5876 797 5880
rect 798 5876 802 5880
rect 809 5876 813 5880
rect 814 5876 818 5880
rect 819 5876 823 5880
rect 824 5876 828 5880
rect 835 5876 839 5880
rect 840 5876 844 5880
rect 845 5876 849 5880
rect 850 5876 854 5880
rect 861 5876 865 5880
rect 866 5876 870 5880
rect 871 5876 875 5880
rect 876 5876 880 5880
rect 1054 5876 1058 5880
rect 1059 5876 1063 5880
rect 1064 5876 1068 5880
rect 1069 5876 1073 5880
rect 1363 5876 1367 5880
rect 1368 5876 1372 5880
rect 1373 5876 1377 5880
rect 1378 5876 1382 5880
rect 1672 5876 1676 5880
rect 1677 5876 1681 5880
rect 1682 5876 1686 5880
rect 1687 5876 1691 5880
rect 1981 5876 1985 5880
rect 1986 5876 1990 5880
rect 1991 5876 1995 5880
rect 1996 5876 2000 5880
rect 2290 5876 2294 5880
rect 2295 5876 2299 5880
rect 2300 5876 2304 5880
rect 2305 5876 2309 5880
rect 2599 5876 2603 5880
rect 2604 5876 2608 5880
rect 2609 5876 2613 5880
rect 2614 5876 2618 5880
rect 2908 5876 2912 5880
rect 2913 5876 2917 5880
rect 2918 5876 2922 5880
rect 2923 5876 2927 5880
rect 3217 5876 3221 5880
rect 3222 5876 3226 5880
rect 3227 5876 3231 5880
rect 3232 5876 3236 5880
rect 3526 5876 3530 5880
rect 3531 5876 3535 5880
rect 3536 5876 3540 5880
rect 3541 5876 3545 5880
rect 3835 5876 3839 5880
rect 3840 5876 3844 5880
rect 3845 5876 3849 5880
rect 3850 5876 3854 5880
rect 4235 5876 4239 5880
rect 4240 5876 4244 5880
rect 4245 5876 4249 5880
rect 4250 5876 4254 5880
rect 4264 5876 4268 5880
rect 4269 5876 4273 5880
rect 4274 5876 4278 5880
rect 4279 5876 4283 5880
rect 4293 5876 4297 5880
rect 4298 5876 4302 5880
rect 4303 5876 4307 5880
rect 4308 5876 4312 5880
rect 4322 5876 4326 5880
rect 4327 5876 4331 5880
rect 4332 5876 4336 5880
rect 4337 5876 4341 5880
rect 4351 5876 4355 5880
rect 4356 5876 4360 5880
rect 4361 5876 4365 5880
rect 4366 5876 4370 5880
rect 757 5866 761 5870
rect 762 5866 766 5870
rect 767 5866 771 5870
rect 772 5866 776 5870
rect 783 5866 787 5870
rect 788 5866 792 5870
rect 793 5866 797 5870
rect 798 5866 802 5870
rect 809 5866 813 5870
rect 814 5866 818 5870
rect 819 5866 823 5870
rect 824 5866 828 5870
rect 835 5866 839 5870
rect 840 5866 844 5870
rect 845 5866 849 5870
rect 850 5866 854 5870
rect 861 5866 865 5870
rect 866 5866 870 5870
rect 871 5866 875 5870
rect 876 5866 880 5870
rect 1054 5866 1058 5870
rect 1059 5866 1063 5870
rect 1064 5866 1068 5870
rect 1069 5866 1073 5870
rect 1363 5866 1367 5870
rect 1368 5866 1372 5870
rect 1373 5866 1377 5870
rect 1378 5866 1382 5870
rect 1672 5866 1676 5870
rect 1677 5866 1681 5870
rect 1682 5866 1686 5870
rect 1687 5866 1691 5870
rect 1981 5866 1985 5870
rect 1986 5866 1990 5870
rect 1991 5866 1995 5870
rect 1996 5866 2000 5870
rect 2290 5866 2294 5870
rect 2295 5866 2299 5870
rect 2300 5866 2304 5870
rect 2305 5866 2309 5870
rect 2599 5866 2603 5870
rect 2604 5866 2608 5870
rect 2609 5866 2613 5870
rect 2614 5866 2618 5870
rect 2908 5866 2912 5870
rect 2913 5866 2917 5870
rect 2918 5866 2922 5870
rect 2923 5866 2927 5870
rect 3217 5866 3221 5870
rect 3222 5866 3226 5870
rect 3227 5866 3231 5870
rect 3232 5866 3236 5870
rect 3526 5866 3530 5870
rect 3531 5866 3535 5870
rect 3536 5866 3540 5870
rect 3541 5866 3545 5870
rect 3835 5866 3839 5870
rect 3840 5866 3844 5870
rect 3845 5866 3849 5870
rect 3850 5866 3854 5870
rect 4235 5866 4239 5870
rect 4240 5866 4244 5870
rect 4245 5866 4249 5870
rect 4250 5866 4254 5870
rect 4264 5866 4268 5870
rect 4269 5866 4273 5870
rect 4274 5866 4278 5870
rect 4279 5866 4283 5870
rect 4293 5866 4297 5870
rect 4298 5866 4302 5870
rect 4303 5866 4307 5870
rect 4308 5866 4312 5870
rect 4322 5866 4326 5870
rect 4327 5866 4331 5870
rect 4332 5866 4336 5870
rect 4337 5866 4341 5870
rect 4351 5866 4355 5870
rect 4356 5866 4360 5870
rect 4361 5866 4365 5870
rect 4366 5866 4370 5870
rect 4627 7975 4631 8015
rect 4666 7975 4670 8034
rect 4709 7975 4713 8034
rect 4750 7975 4754 8034
<< nsubstratencontact >>
rect 1372 9974 1376 9978
rect 1377 9974 1381 9978
rect 1382 9974 1386 9978
rect 1387 9974 1391 9978
rect 1392 9974 1396 9978
rect 1397 9974 1401 9978
rect 1402 9974 1406 9978
rect 1407 9974 1411 9978
rect 1412 9974 1416 9978
rect 1417 9974 1421 9978
rect 1422 9974 1426 9978
rect 1427 9974 1431 9978
rect 1432 9974 1436 9978
rect 1437 9974 1441 9978
rect 1442 9974 1446 9978
rect 1447 9974 1451 9978
rect 1452 9974 1456 9978
rect 1457 9974 1461 9978
rect 1462 9974 1466 9978
rect 1372 9969 1376 9973
rect 1372 9964 1376 9968
rect 1462 9969 1466 9973
rect 1372 9959 1376 9963
rect 1372 9954 1376 9958
rect 1372 9949 1376 9953
rect 1372 9944 1376 9948
rect 1372 9939 1376 9943
rect 1372 9934 1376 9938
rect 1372 9929 1376 9933
rect 1372 9924 1376 9928
rect 1372 9919 1376 9923
rect 1372 9914 1376 9918
rect 1372 9909 1376 9913
rect 1372 9904 1376 9908
rect 1372 9899 1376 9903
rect 1372 9894 1376 9898
rect 1372 9889 1376 9893
rect 1372 9884 1376 9888
rect 1372 9879 1376 9883
rect 1372 9874 1376 9878
rect 1372 9869 1376 9873
rect 1372 9864 1376 9868
rect 1372 9859 1376 9863
rect 1372 9854 1376 9858
rect 1372 9849 1376 9853
rect 1462 9964 1466 9968
rect 1462 9959 1466 9963
rect 1462 9954 1466 9958
rect 1462 9949 1466 9953
rect 1462 9944 1466 9948
rect 1462 9939 1466 9943
rect 1462 9934 1466 9938
rect 1462 9929 1466 9933
rect 1462 9924 1466 9928
rect 1462 9919 1466 9923
rect 1462 9914 1466 9918
rect 1462 9909 1466 9913
rect 1462 9904 1466 9908
rect 1462 9899 1466 9903
rect 1462 9894 1466 9898
rect 1462 9889 1466 9893
rect 1462 9884 1466 9888
rect 1462 9879 1466 9883
rect 1462 9874 1466 9878
rect 1462 9869 1466 9873
rect 1462 9864 1466 9868
rect 1462 9859 1466 9863
rect 1462 9854 1466 9858
rect 1372 9844 1376 9848
rect 1462 9849 1466 9853
rect 1462 9844 1466 9848
rect 1372 9839 1376 9843
rect 1377 9839 1381 9843
rect 1382 9839 1386 9843
rect 1387 9839 1391 9843
rect 1392 9839 1396 9843
rect 1397 9839 1401 9843
rect 1402 9839 1406 9843
rect 1407 9839 1411 9843
rect 1412 9839 1416 9843
rect 1417 9839 1421 9843
rect 1422 9839 1426 9843
rect 1427 9839 1431 9843
rect 1432 9839 1436 9843
rect 1437 9839 1441 9843
rect 1442 9839 1446 9843
rect 1447 9839 1451 9843
rect 1452 9839 1456 9843
rect 1457 9839 1461 9843
rect 1462 9839 1466 9843
rect 1545 9961 1549 9965
rect 1552 9961 1556 9965
rect 1557 9961 1561 9965
rect 1562 9961 1566 9965
rect 1567 9961 1571 9965
rect 1572 9961 1576 9965
rect 1577 9961 1581 9965
rect 1582 9961 1586 9965
rect 1587 9961 1591 9965
rect 1592 9961 1596 9965
rect 1597 9961 1601 9965
rect 1602 9961 1606 9965
rect 1609 9961 1613 9965
rect 1545 9954 1549 9958
rect 1609 9954 1613 9958
rect 1545 9949 1549 9953
rect 1545 9944 1549 9948
rect 1545 9939 1549 9943
rect 1545 9934 1549 9938
rect 1545 9929 1549 9933
rect 1545 9924 1549 9928
rect 1545 9919 1549 9923
rect 1545 9914 1549 9918
rect 1545 9909 1549 9913
rect 1545 9904 1549 9908
rect 1545 9899 1549 9903
rect 1545 9894 1549 9898
rect 1545 9889 1549 9893
rect 1545 9884 1549 9888
rect 1545 9879 1549 9883
rect 1545 9874 1549 9878
rect 1545 9869 1549 9873
rect 1545 9864 1549 9868
rect 1609 9949 1613 9953
rect 1609 9944 1613 9948
rect 1609 9939 1613 9943
rect 1609 9934 1613 9938
rect 1609 9929 1613 9933
rect 1609 9924 1613 9928
rect 1609 9919 1613 9923
rect 1609 9914 1613 9918
rect 1609 9909 1613 9913
rect 1609 9904 1613 9908
rect 1609 9899 1613 9903
rect 1609 9894 1613 9898
rect 1609 9889 1613 9893
rect 1609 9884 1613 9888
rect 1609 9879 1613 9883
rect 1609 9874 1613 9878
rect 1609 9869 1613 9873
rect 1609 9864 1613 9868
rect 1545 9859 1549 9863
rect 1609 9859 1613 9863
rect 1545 9852 1549 9856
rect 1552 9852 1556 9856
rect 1557 9852 1561 9856
rect 1562 9852 1566 9856
rect 1567 9852 1571 9856
rect 1572 9852 1576 9856
rect 1577 9852 1581 9856
rect 1582 9852 1586 9856
rect 1587 9852 1591 9856
rect 1592 9852 1596 9856
rect 1597 9852 1601 9856
rect 1602 9852 1606 9856
rect 1609 9852 1613 9856
rect 1681 9974 1685 9978
rect 1686 9974 1690 9978
rect 1691 9974 1695 9978
rect 1696 9974 1700 9978
rect 1701 9974 1705 9978
rect 1706 9974 1710 9978
rect 1711 9974 1715 9978
rect 1716 9974 1720 9978
rect 1721 9974 1725 9978
rect 1726 9974 1730 9978
rect 1731 9974 1735 9978
rect 1736 9974 1740 9978
rect 1741 9974 1745 9978
rect 1746 9974 1750 9978
rect 1751 9974 1755 9978
rect 1756 9974 1760 9978
rect 1761 9974 1765 9978
rect 1766 9974 1770 9978
rect 1771 9974 1775 9978
rect 1681 9969 1685 9973
rect 1681 9964 1685 9968
rect 1771 9969 1775 9973
rect 1681 9959 1685 9963
rect 1681 9954 1685 9958
rect 1681 9949 1685 9953
rect 1681 9944 1685 9948
rect 1681 9939 1685 9943
rect 1681 9934 1685 9938
rect 1681 9929 1685 9933
rect 1681 9924 1685 9928
rect 1681 9919 1685 9923
rect 1681 9914 1685 9918
rect 1681 9909 1685 9913
rect 1681 9904 1685 9908
rect 1681 9899 1685 9903
rect 1681 9894 1685 9898
rect 1681 9889 1685 9893
rect 1681 9884 1685 9888
rect 1681 9879 1685 9883
rect 1681 9874 1685 9878
rect 1681 9869 1685 9873
rect 1681 9864 1685 9868
rect 1681 9859 1685 9863
rect 1681 9854 1685 9858
rect 1681 9849 1685 9853
rect 1771 9964 1775 9968
rect 1771 9959 1775 9963
rect 1771 9954 1775 9958
rect 1771 9949 1775 9953
rect 1771 9944 1775 9948
rect 1771 9939 1775 9943
rect 1771 9934 1775 9938
rect 1771 9929 1775 9933
rect 1771 9924 1775 9928
rect 1771 9919 1775 9923
rect 1771 9914 1775 9918
rect 1771 9909 1775 9913
rect 1771 9904 1775 9908
rect 1771 9899 1775 9903
rect 1771 9894 1775 9898
rect 1771 9889 1775 9893
rect 1771 9884 1775 9888
rect 1771 9879 1775 9883
rect 1771 9874 1775 9878
rect 1771 9869 1775 9873
rect 1771 9864 1775 9868
rect 1771 9859 1775 9863
rect 1771 9854 1775 9858
rect 1681 9844 1685 9848
rect 1771 9849 1775 9853
rect 1771 9844 1775 9848
rect 1681 9839 1685 9843
rect 1686 9839 1690 9843
rect 1691 9839 1695 9843
rect 1696 9839 1700 9843
rect 1701 9839 1705 9843
rect 1706 9839 1710 9843
rect 1711 9839 1715 9843
rect 1716 9839 1720 9843
rect 1721 9839 1725 9843
rect 1726 9839 1730 9843
rect 1731 9839 1735 9843
rect 1736 9839 1740 9843
rect 1741 9839 1745 9843
rect 1746 9839 1750 9843
rect 1751 9839 1755 9843
rect 1756 9839 1760 9843
rect 1761 9839 1765 9843
rect 1766 9839 1770 9843
rect 1771 9839 1775 9843
rect 1854 9961 1858 9965
rect 1861 9961 1865 9965
rect 1866 9961 1870 9965
rect 1871 9961 1875 9965
rect 1876 9961 1880 9965
rect 1881 9961 1885 9965
rect 1886 9961 1890 9965
rect 1891 9961 1895 9965
rect 1896 9961 1900 9965
rect 1901 9961 1905 9965
rect 1906 9961 1910 9965
rect 1911 9961 1915 9965
rect 1918 9961 1922 9965
rect 1854 9954 1858 9958
rect 1918 9954 1922 9958
rect 1854 9949 1858 9953
rect 1854 9944 1858 9948
rect 1854 9939 1858 9943
rect 1854 9934 1858 9938
rect 1854 9929 1858 9933
rect 1854 9924 1858 9928
rect 1854 9919 1858 9923
rect 1854 9914 1858 9918
rect 1854 9909 1858 9913
rect 1854 9904 1858 9908
rect 1854 9899 1858 9903
rect 1854 9894 1858 9898
rect 1854 9889 1858 9893
rect 1854 9884 1858 9888
rect 1854 9879 1858 9883
rect 1854 9874 1858 9878
rect 1854 9869 1858 9873
rect 1854 9864 1858 9868
rect 1918 9949 1922 9953
rect 1918 9944 1922 9948
rect 1918 9939 1922 9943
rect 1918 9934 1922 9938
rect 1918 9929 1922 9933
rect 1918 9924 1922 9928
rect 1918 9919 1922 9923
rect 1918 9914 1922 9918
rect 1918 9909 1922 9913
rect 1918 9904 1922 9908
rect 1918 9899 1922 9903
rect 1918 9894 1922 9898
rect 1918 9889 1922 9893
rect 1918 9884 1922 9888
rect 1918 9879 1922 9883
rect 1918 9874 1922 9878
rect 1918 9869 1922 9873
rect 1918 9864 1922 9868
rect 1854 9859 1858 9863
rect 1918 9859 1922 9863
rect 1854 9852 1858 9856
rect 1861 9852 1865 9856
rect 1866 9852 1870 9856
rect 1871 9852 1875 9856
rect 1876 9852 1880 9856
rect 1881 9852 1885 9856
rect 1886 9852 1890 9856
rect 1891 9852 1895 9856
rect 1896 9852 1900 9856
rect 1901 9852 1905 9856
rect 1906 9852 1910 9856
rect 1911 9852 1915 9856
rect 1918 9852 1922 9856
rect 1990 9974 1994 9978
rect 1995 9974 1999 9978
rect 2000 9974 2004 9978
rect 2005 9974 2009 9978
rect 2010 9974 2014 9978
rect 2015 9974 2019 9978
rect 2020 9974 2024 9978
rect 2025 9974 2029 9978
rect 2030 9974 2034 9978
rect 2035 9974 2039 9978
rect 2040 9974 2044 9978
rect 2045 9974 2049 9978
rect 2050 9974 2054 9978
rect 2055 9974 2059 9978
rect 2060 9974 2064 9978
rect 2065 9974 2069 9978
rect 2070 9974 2074 9978
rect 2075 9974 2079 9978
rect 2080 9974 2084 9978
rect 1990 9969 1994 9973
rect 1990 9964 1994 9968
rect 2080 9969 2084 9973
rect 1990 9959 1994 9963
rect 1990 9954 1994 9958
rect 1990 9949 1994 9953
rect 1990 9944 1994 9948
rect 1990 9939 1994 9943
rect 1990 9934 1994 9938
rect 1990 9929 1994 9933
rect 1990 9924 1994 9928
rect 1990 9919 1994 9923
rect 1990 9914 1994 9918
rect 1990 9909 1994 9913
rect 1990 9904 1994 9908
rect 1990 9899 1994 9903
rect 1990 9894 1994 9898
rect 1990 9889 1994 9893
rect 1990 9884 1994 9888
rect 1990 9879 1994 9883
rect 1990 9874 1994 9878
rect 1990 9869 1994 9873
rect 1990 9864 1994 9868
rect 1990 9859 1994 9863
rect 1990 9854 1994 9858
rect 1990 9849 1994 9853
rect 2080 9964 2084 9968
rect 2080 9959 2084 9963
rect 2080 9954 2084 9958
rect 2080 9949 2084 9953
rect 2080 9944 2084 9948
rect 2080 9939 2084 9943
rect 2080 9934 2084 9938
rect 2080 9929 2084 9933
rect 2080 9924 2084 9928
rect 2080 9919 2084 9923
rect 2080 9914 2084 9918
rect 2080 9909 2084 9913
rect 2080 9904 2084 9908
rect 2080 9899 2084 9903
rect 2080 9894 2084 9898
rect 2080 9889 2084 9893
rect 2080 9884 2084 9888
rect 2080 9879 2084 9883
rect 2080 9874 2084 9878
rect 2080 9869 2084 9873
rect 2080 9864 2084 9868
rect 2080 9859 2084 9863
rect 2080 9854 2084 9858
rect 1990 9844 1994 9848
rect 2080 9849 2084 9853
rect 2080 9844 2084 9848
rect 1990 9839 1994 9843
rect 1995 9839 1999 9843
rect 2000 9839 2004 9843
rect 2005 9839 2009 9843
rect 2010 9839 2014 9843
rect 2015 9839 2019 9843
rect 2020 9839 2024 9843
rect 2025 9839 2029 9843
rect 2030 9839 2034 9843
rect 2035 9839 2039 9843
rect 2040 9839 2044 9843
rect 2045 9839 2049 9843
rect 2050 9839 2054 9843
rect 2055 9839 2059 9843
rect 2060 9839 2064 9843
rect 2065 9839 2069 9843
rect 2070 9839 2074 9843
rect 2075 9839 2079 9843
rect 2080 9839 2084 9843
rect 2163 9961 2167 9965
rect 2170 9961 2174 9965
rect 2175 9961 2179 9965
rect 2180 9961 2184 9965
rect 2185 9961 2189 9965
rect 2190 9961 2194 9965
rect 2195 9961 2199 9965
rect 2200 9961 2204 9965
rect 2205 9961 2209 9965
rect 2210 9961 2214 9965
rect 2215 9961 2219 9965
rect 2220 9961 2224 9965
rect 2227 9961 2231 9965
rect 2163 9954 2167 9958
rect 2227 9954 2231 9958
rect 2163 9949 2167 9953
rect 2163 9944 2167 9948
rect 2163 9939 2167 9943
rect 2163 9934 2167 9938
rect 2163 9929 2167 9933
rect 2163 9924 2167 9928
rect 2163 9919 2167 9923
rect 2163 9914 2167 9918
rect 2163 9909 2167 9913
rect 2163 9904 2167 9908
rect 2163 9899 2167 9903
rect 2163 9894 2167 9898
rect 2163 9889 2167 9893
rect 2163 9884 2167 9888
rect 2163 9879 2167 9883
rect 2163 9874 2167 9878
rect 2163 9869 2167 9873
rect 2163 9864 2167 9868
rect 2227 9949 2231 9953
rect 2227 9944 2231 9948
rect 2227 9939 2231 9943
rect 2227 9934 2231 9938
rect 2227 9929 2231 9933
rect 2227 9924 2231 9928
rect 2227 9919 2231 9923
rect 2227 9914 2231 9918
rect 2227 9909 2231 9913
rect 2227 9904 2231 9908
rect 2227 9899 2231 9903
rect 2227 9894 2231 9898
rect 2227 9889 2231 9893
rect 2227 9884 2231 9888
rect 2227 9879 2231 9883
rect 2227 9874 2231 9878
rect 2227 9869 2231 9873
rect 2227 9864 2231 9868
rect 2163 9859 2167 9863
rect 2227 9859 2231 9863
rect 2163 9852 2167 9856
rect 2170 9852 2174 9856
rect 2175 9852 2179 9856
rect 2180 9852 2184 9856
rect 2185 9852 2189 9856
rect 2190 9852 2194 9856
rect 2195 9852 2199 9856
rect 2200 9852 2204 9856
rect 2205 9852 2209 9856
rect 2210 9852 2214 9856
rect 2215 9852 2219 9856
rect 2220 9852 2224 9856
rect 2227 9852 2231 9856
rect 2299 9974 2303 9978
rect 2304 9974 2308 9978
rect 2309 9974 2313 9978
rect 2314 9974 2318 9978
rect 2319 9974 2323 9978
rect 2324 9974 2328 9978
rect 2329 9974 2333 9978
rect 2334 9974 2338 9978
rect 2339 9974 2343 9978
rect 2344 9974 2348 9978
rect 2349 9974 2353 9978
rect 2354 9974 2358 9978
rect 2359 9974 2363 9978
rect 2364 9974 2368 9978
rect 2369 9974 2373 9978
rect 2374 9974 2378 9978
rect 2379 9974 2383 9978
rect 2384 9974 2388 9978
rect 2389 9974 2393 9978
rect 2299 9969 2303 9973
rect 2299 9964 2303 9968
rect 2389 9969 2393 9973
rect 2299 9959 2303 9963
rect 2299 9954 2303 9958
rect 2299 9949 2303 9953
rect 2299 9944 2303 9948
rect 2299 9939 2303 9943
rect 2299 9934 2303 9938
rect 2299 9929 2303 9933
rect 2299 9924 2303 9928
rect 2299 9919 2303 9923
rect 2299 9914 2303 9918
rect 2299 9909 2303 9913
rect 2299 9904 2303 9908
rect 2299 9899 2303 9903
rect 2299 9894 2303 9898
rect 2299 9889 2303 9893
rect 2299 9884 2303 9888
rect 2299 9879 2303 9883
rect 2299 9874 2303 9878
rect 2299 9869 2303 9873
rect 2299 9864 2303 9868
rect 2299 9859 2303 9863
rect 2299 9854 2303 9858
rect 2299 9849 2303 9853
rect 2389 9964 2393 9968
rect 2389 9959 2393 9963
rect 2389 9954 2393 9958
rect 2389 9949 2393 9953
rect 2389 9944 2393 9948
rect 2389 9939 2393 9943
rect 2389 9934 2393 9938
rect 2389 9929 2393 9933
rect 2389 9924 2393 9928
rect 2389 9919 2393 9923
rect 2389 9914 2393 9918
rect 2389 9909 2393 9913
rect 2389 9904 2393 9908
rect 2389 9899 2393 9903
rect 2389 9894 2393 9898
rect 2389 9889 2393 9893
rect 2389 9884 2393 9888
rect 2389 9879 2393 9883
rect 2389 9874 2393 9878
rect 2389 9869 2393 9873
rect 2389 9864 2393 9868
rect 2389 9859 2393 9863
rect 2389 9854 2393 9858
rect 2299 9844 2303 9848
rect 2389 9849 2393 9853
rect 2389 9844 2393 9848
rect 2299 9839 2303 9843
rect 2304 9839 2308 9843
rect 2309 9839 2313 9843
rect 2314 9839 2318 9843
rect 2319 9839 2323 9843
rect 2324 9839 2328 9843
rect 2329 9839 2333 9843
rect 2334 9839 2338 9843
rect 2339 9839 2343 9843
rect 2344 9839 2348 9843
rect 2349 9839 2353 9843
rect 2354 9839 2358 9843
rect 2359 9839 2363 9843
rect 2364 9839 2368 9843
rect 2369 9839 2373 9843
rect 2374 9839 2378 9843
rect 2379 9839 2383 9843
rect 2384 9839 2388 9843
rect 2389 9839 2393 9843
rect 2472 9961 2476 9965
rect 2479 9961 2483 9965
rect 2484 9961 2488 9965
rect 2489 9961 2493 9965
rect 2494 9961 2498 9965
rect 2499 9961 2503 9965
rect 2504 9961 2508 9965
rect 2509 9961 2513 9965
rect 2514 9961 2518 9965
rect 2519 9961 2523 9965
rect 2524 9961 2528 9965
rect 2529 9961 2533 9965
rect 2536 9961 2540 9965
rect 2472 9954 2476 9958
rect 2536 9954 2540 9958
rect 2472 9949 2476 9953
rect 2472 9944 2476 9948
rect 2472 9939 2476 9943
rect 2472 9934 2476 9938
rect 2472 9929 2476 9933
rect 2472 9924 2476 9928
rect 2472 9919 2476 9923
rect 2472 9914 2476 9918
rect 2472 9909 2476 9913
rect 2472 9904 2476 9908
rect 2472 9899 2476 9903
rect 2472 9894 2476 9898
rect 2472 9889 2476 9893
rect 2472 9884 2476 9888
rect 2472 9879 2476 9883
rect 2472 9874 2476 9878
rect 2472 9869 2476 9873
rect 2472 9864 2476 9868
rect 2536 9949 2540 9953
rect 2536 9944 2540 9948
rect 2536 9939 2540 9943
rect 2536 9934 2540 9938
rect 2536 9929 2540 9933
rect 2536 9924 2540 9928
rect 2536 9919 2540 9923
rect 2536 9914 2540 9918
rect 2536 9909 2540 9913
rect 2536 9904 2540 9908
rect 2536 9899 2540 9903
rect 2536 9894 2540 9898
rect 2536 9889 2540 9893
rect 2536 9884 2540 9888
rect 2536 9879 2540 9883
rect 2536 9874 2540 9878
rect 2536 9869 2540 9873
rect 2536 9864 2540 9868
rect 2472 9859 2476 9863
rect 2536 9859 2540 9863
rect 2472 9852 2476 9856
rect 2479 9852 2483 9856
rect 2484 9852 2488 9856
rect 2489 9852 2493 9856
rect 2494 9852 2498 9856
rect 2499 9852 2503 9856
rect 2504 9852 2508 9856
rect 2509 9852 2513 9856
rect 2514 9852 2518 9856
rect 2519 9852 2523 9856
rect 2524 9852 2528 9856
rect 2529 9852 2533 9856
rect 2536 9852 2540 9856
rect 2608 9974 2612 9978
rect 2613 9974 2617 9978
rect 2618 9974 2622 9978
rect 2623 9974 2627 9978
rect 2628 9974 2632 9978
rect 2633 9974 2637 9978
rect 2638 9974 2642 9978
rect 2643 9974 2647 9978
rect 2648 9974 2652 9978
rect 2653 9974 2657 9978
rect 2658 9974 2662 9978
rect 2663 9974 2667 9978
rect 2668 9974 2672 9978
rect 2673 9974 2677 9978
rect 2678 9974 2682 9978
rect 2683 9974 2687 9978
rect 2688 9974 2692 9978
rect 2693 9974 2697 9978
rect 2698 9974 2702 9978
rect 2608 9969 2612 9973
rect 2608 9964 2612 9968
rect 2698 9969 2702 9973
rect 2608 9959 2612 9963
rect 2608 9954 2612 9958
rect 2608 9949 2612 9953
rect 2608 9944 2612 9948
rect 2608 9939 2612 9943
rect 2608 9934 2612 9938
rect 2608 9929 2612 9933
rect 2608 9924 2612 9928
rect 2608 9919 2612 9923
rect 2608 9914 2612 9918
rect 2608 9909 2612 9913
rect 2608 9904 2612 9908
rect 2608 9899 2612 9903
rect 2608 9894 2612 9898
rect 2608 9889 2612 9893
rect 2608 9884 2612 9888
rect 2608 9879 2612 9883
rect 2608 9874 2612 9878
rect 2608 9869 2612 9873
rect 2608 9864 2612 9868
rect 2608 9859 2612 9863
rect 2608 9854 2612 9858
rect 2608 9849 2612 9853
rect 2698 9964 2702 9968
rect 2698 9959 2702 9963
rect 2698 9954 2702 9958
rect 2698 9949 2702 9953
rect 2698 9944 2702 9948
rect 2698 9939 2702 9943
rect 2698 9934 2702 9938
rect 2698 9929 2702 9933
rect 2698 9924 2702 9928
rect 2698 9919 2702 9923
rect 2698 9914 2702 9918
rect 2698 9909 2702 9913
rect 2698 9904 2702 9908
rect 2698 9899 2702 9903
rect 2698 9894 2702 9898
rect 2698 9889 2702 9893
rect 2698 9884 2702 9888
rect 2698 9879 2702 9883
rect 2698 9874 2702 9878
rect 2698 9869 2702 9873
rect 2698 9864 2702 9868
rect 2698 9859 2702 9863
rect 2698 9854 2702 9858
rect 2608 9844 2612 9848
rect 2698 9849 2702 9853
rect 2698 9844 2702 9848
rect 2608 9839 2612 9843
rect 2613 9839 2617 9843
rect 2618 9839 2622 9843
rect 2623 9839 2627 9843
rect 2628 9839 2632 9843
rect 2633 9839 2637 9843
rect 2638 9839 2642 9843
rect 2643 9839 2647 9843
rect 2648 9839 2652 9843
rect 2653 9839 2657 9843
rect 2658 9839 2662 9843
rect 2663 9839 2667 9843
rect 2668 9839 2672 9843
rect 2673 9839 2677 9843
rect 2678 9839 2682 9843
rect 2683 9839 2687 9843
rect 2688 9839 2692 9843
rect 2693 9839 2697 9843
rect 2698 9839 2702 9843
rect 2781 9961 2785 9965
rect 2788 9961 2792 9965
rect 2793 9961 2797 9965
rect 2798 9961 2802 9965
rect 2803 9961 2807 9965
rect 2808 9961 2812 9965
rect 2813 9961 2817 9965
rect 2818 9961 2822 9965
rect 2823 9961 2827 9965
rect 2828 9961 2832 9965
rect 2833 9961 2837 9965
rect 2838 9961 2842 9965
rect 2845 9961 2849 9965
rect 2781 9954 2785 9958
rect 2845 9954 2849 9958
rect 2781 9949 2785 9953
rect 2781 9944 2785 9948
rect 2781 9939 2785 9943
rect 2781 9934 2785 9938
rect 2781 9929 2785 9933
rect 2781 9924 2785 9928
rect 2781 9919 2785 9923
rect 2781 9914 2785 9918
rect 2781 9909 2785 9913
rect 2781 9904 2785 9908
rect 2781 9899 2785 9903
rect 2781 9894 2785 9898
rect 2781 9889 2785 9893
rect 2781 9884 2785 9888
rect 2781 9879 2785 9883
rect 2781 9874 2785 9878
rect 2781 9869 2785 9873
rect 2781 9864 2785 9868
rect 2845 9949 2849 9953
rect 2845 9944 2849 9948
rect 2845 9939 2849 9943
rect 2845 9934 2849 9938
rect 2845 9929 2849 9933
rect 2845 9924 2849 9928
rect 2845 9919 2849 9923
rect 2845 9914 2849 9918
rect 2845 9909 2849 9913
rect 2845 9904 2849 9908
rect 2845 9899 2849 9903
rect 2845 9894 2849 9898
rect 2845 9889 2849 9893
rect 2845 9884 2849 9888
rect 2845 9879 2849 9883
rect 2845 9874 2849 9878
rect 2845 9869 2849 9873
rect 2845 9864 2849 9868
rect 2781 9859 2785 9863
rect 2845 9859 2849 9863
rect 2781 9852 2785 9856
rect 2788 9852 2792 9856
rect 2793 9852 2797 9856
rect 2798 9852 2802 9856
rect 2803 9852 2807 9856
rect 2808 9852 2812 9856
rect 2813 9852 2817 9856
rect 2818 9852 2822 9856
rect 2823 9852 2827 9856
rect 2828 9852 2832 9856
rect 2833 9852 2837 9856
rect 2838 9852 2842 9856
rect 2845 9852 2849 9856
rect 2917 9974 2921 9978
rect 2922 9974 2926 9978
rect 2927 9974 2931 9978
rect 2932 9974 2936 9978
rect 2937 9974 2941 9978
rect 2942 9974 2946 9978
rect 2947 9974 2951 9978
rect 2952 9974 2956 9978
rect 2957 9974 2961 9978
rect 2962 9974 2966 9978
rect 2967 9974 2971 9978
rect 2972 9974 2976 9978
rect 2977 9974 2981 9978
rect 2982 9974 2986 9978
rect 2987 9974 2991 9978
rect 2992 9974 2996 9978
rect 2997 9974 3001 9978
rect 3002 9974 3006 9978
rect 3007 9974 3011 9978
rect 2917 9969 2921 9973
rect 2917 9964 2921 9968
rect 3007 9969 3011 9973
rect 2917 9959 2921 9963
rect 2917 9954 2921 9958
rect 2917 9949 2921 9953
rect 2917 9944 2921 9948
rect 2917 9939 2921 9943
rect 2917 9934 2921 9938
rect 2917 9929 2921 9933
rect 2917 9924 2921 9928
rect 2917 9919 2921 9923
rect 2917 9914 2921 9918
rect 2917 9909 2921 9913
rect 2917 9904 2921 9908
rect 2917 9899 2921 9903
rect 2917 9894 2921 9898
rect 2917 9889 2921 9893
rect 2917 9884 2921 9888
rect 2917 9879 2921 9883
rect 2917 9874 2921 9878
rect 2917 9869 2921 9873
rect 2917 9864 2921 9868
rect 2917 9859 2921 9863
rect 2917 9854 2921 9858
rect 2917 9849 2921 9853
rect 3007 9964 3011 9968
rect 3007 9959 3011 9963
rect 3007 9954 3011 9958
rect 3007 9949 3011 9953
rect 3007 9944 3011 9948
rect 3007 9939 3011 9943
rect 3007 9934 3011 9938
rect 3007 9929 3011 9933
rect 3007 9924 3011 9928
rect 3007 9919 3011 9923
rect 3007 9914 3011 9918
rect 3007 9909 3011 9913
rect 3007 9904 3011 9908
rect 3007 9899 3011 9903
rect 3007 9894 3011 9898
rect 3007 9889 3011 9893
rect 3007 9884 3011 9888
rect 3007 9879 3011 9883
rect 3007 9874 3011 9878
rect 3007 9869 3011 9873
rect 3007 9864 3011 9868
rect 3007 9859 3011 9863
rect 3007 9854 3011 9858
rect 2917 9844 2921 9848
rect 3007 9849 3011 9853
rect 3007 9844 3011 9848
rect 2917 9839 2921 9843
rect 2922 9839 2926 9843
rect 2927 9839 2931 9843
rect 2932 9839 2936 9843
rect 2937 9839 2941 9843
rect 2942 9839 2946 9843
rect 2947 9839 2951 9843
rect 2952 9839 2956 9843
rect 2957 9839 2961 9843
rect 2962 9839 2966 9843
rect 2967 9839 2971 9843
rect 2972 9839 2976 9843
rect 2977 9839 2981 9843
rect 2982 9839 2986 9843
rect 2987 9839 2991 9843
rect 2992 9839 2996 9843
rect 2997 9839 3001 9843
rect 3002 9839 3006 9843
rect 3007 9839 3011 9843
rect 3090 9961 3094 9965
rect 3097 9961 3101 9965
rect 3102 9961 3106 9965
rect 3107 9961 3111 9965
rect 3112 9961 3116 9965
rect 3117 9961 3121 9965
rect 3122 9961 3126 9965
rect 3127 9961 3131 9965
rect 3132 9961 3136 9965
rect 3137 9961 3141 9965
rect 3142 9961 3146 9965
rect 3147 9961 3151 9965
rect 3154 9961 3158 9965
rect 3090 9954 3094 9958
rect 3154 9954 3158 9958
rect 3090 9949 3094 9953
rect 3090 9944 3094 9948
rect 3090 9939 3094 9943
rect 3090 9934 3094 9938
rect 3090 9929 3094 9933
rect 3090 9924 3094 9928
rect 3090 9919 3094 9923
rect 3090 9914 3094 9918
rect 3090 9909 3094 9913
rect 3090 9904 3094 9908
rect 3090 9899 3094 9903
rect 3090 9894 3094 9898
rect 3090 9889 3094 9893
rect 3090 9884 3094 9888
rect 3090 9879 3094 9883
rect 3090 9874 3094 9878
rect 3090 9869 3094 9873
rect 3090 9864 3094 9868
rect 3154 9949 3158 9953
rect 3154 9944 3158 9948
rect 3154 9939 3158 9943
rect 3154 9934 3158 9938
rect 3154 9929 3158 9933
rect 3154 9924 3158 9928
rect 3154 9919 3158 9923
rect 3154 9914 3158 9918
rect 3154 9909 3158 9913
rect 3154 9904 3158 9908
rect 3154 9899 3158 9903
rect 3154 9894 3158 9898
rect 3154 9889 3158 9893
rect 3154 9884 3158 9888
rect 3154 9879 3158 9883
rect 3154 9874 3158 9878
rect 3154 9869 3158 9873
rect 3154 9864 3158 9868
rect 3090 9859 3094 9863
rect 3154 9859 3158 9863
rect 3090 9852 3094 9856
rect 3097 9852 3101 9856
rect 3102 9852 3106 9856
rect 3107 9852 3111 9856
rect 3112 9852 3116 9856
rect 3117 9852 3121 9856
rect 3122 9852 3126 9856
rect 3127 9852 3131 9856
rect 3132 9852 3136 9856
rect 3137 9852 3141 9856
rect 3142 9852 3146 9856
rect 3147 9852 3151 9856
rect 3154 9852 3158 9856
rect 3226 9974 3230 9978
rect 3231 9974 3235 9978
rect 3236 9974 3240 9978
rect 3241 9974 3245 9978
rect 3246 9974 3250 9978
rect 3251 9974 3255 9978
rect 3256 9974 3260 9978
rect 3261 9974 3265 9978
rect 3266 9974 3270 9978
rect 3271 9974 3275 9978
rect 3276 9974 3280 9978
rect 3281 9974 3285 9978
rect 3286 9974 3290 9978
rect 3291 9974 3295 9978
rect 3296 9974 3300 9978
rect 3301 9974 3305 9978
rect 3306 9974 3310 9978
rect 3311 9974 3315 9978
rect 3316 9974 3320 9978
rect 3226 9969 3230 9973
rect 3226 9964 3230 9968
rect 3316 9969 3320 9973
rect 3226 9959 3230 9963
rect 3226 9954 3230 9958
rect 3226 9949 3230 9953
rect 3226 9944 3230 9948
rect 3226 9939 3230 9943
rect 3226 9934 3230 9938
rect 3226 9929 3230 9933
rect 3226 9924 3230 9928
rect 3226 9919 3230 9923
rect 3226 9914 3230 9918
rect 3226 9909 3230 9913
rect 3226 9904 3230 9908
rect 3226 9899 3230 9903
rect 3226 9894 3230 9898
rect 3226 9889 3230 9893
rect 3226 9884 3230 9888
rect 3226 9879 3230 9883
rect 3226 9874 3230 9878
rect 3226 9869 3230 9873
rect 3226 9864 3230 9868
rect 3226 9859 3230 9863
rect 3226 9854 3230 9858
rect 3226 9849 3230 9853
rect 3316 9964 3320 9968
rect 3316 9959 3320 9963
rect 3316 9954 3320 9958
rect 3316 9949 3320 9953
rect 3316 9944 3320 9948
rect 3316 9939 3320 9943
rect 3316 9934 3320 9938
rect 3316 9929 3320 9933
rect 3316 9924 3320 9928
rect 3316 9919 3320 9923
rect 3316 9914 3320 9918
rect 3316 9909 3320 9913
rect 3316 9904 3320 9908
rect 3316 9899 3320 9903
rect 3316 9894 3320 9898
rect 3316 9889 3320 9893
rect 3316 9884 3320 9888
rect 3316 9879 3320 9883
rect 3316 9874 3320 9878
rect 3316 9869 3320 9873
rect 3316 9864 3320 9868
rect 3316 9859 3320 9863
rect 3316 9854 3320 9858
rect 3226 9844 3230 9848
rect 3316 9849 3320 9853
rect 3316 9844 3320 9848
rect 3226 9839 3230 9843
rect 3231 9839 3235 9843
rect 3236 9839 3240 9843
rect 3241 9839 3245 9843
rect 3246 9839 3250 9843
rect 3251 9839 3255 9843
rect 3256 9839 3260 9843
rect 3261 9839 3265 9843
rect 3266 9839 3270 9843
rect 3271 9839 3275 9843
rect 3276 9839 3280 9843
rect 3281 9839 3285 9843
rect 3286 9839 3290 9843
rect 3291 9839 3295 9843
rect 3296 9839 3300 9843
rect 3301 9839 3305 9843
rect 3306 9839 3310 9843
rect 3311 9839 3315 9843
rect 3316 9839 3320 9843
rect 3399 9961 3403 9965
rect 3406 9961 3410 9965
rect 3411 9961 3415 9965
rect 3416 9961 3420 9965
rect 3421 9961 3425 9965
rect 3426 9961 3430 9965
rect 3431 9961 3435 9965
rect 3436 9961 3440 9965
rect 3441 9961 3445 9965
rect 3446 9961 3450 9965
rect 3451 9961 3455 9965
rect 3456 9961 3460 9965
rect 3463 9961 3467 9965
rect 3399 9954 3403 9958
rect 3463 9954 3467 9958
rect 3399 9949 3403 9953
rect 3399 9944 3403 9948
rect 3399 9939 3403 9943
rect 3399 9934 3403 9938
rect 3399 9929 3403 9933
rect 3399 9924 3403 9928
rect 3399 9919 3403 9923
rect 3399 9914 3403 9918
rect 3399 9909 3403 9913
rect 3399 9904 3403 9908
rect 3399 9899 3403 9903
rect 3399 9894 3403 9898
rect 3399 9889 3403 9893
rect 3399 9884 3403 9888
rect 3399 9879 3403 9883
rect 3399 9874 3403 9878
rect 3399 9869 3403 9873
rect 3399 9864 3403 9868
rect 3463 9949 3467 9953
rect 3463 9944 3467 9948
rect 3463 9939 3467 9943
rect 3463 9934 3467 9938
rect 3463 9929 3467 9933
rect 3463 9924 3467 9928
rect 3463 9919 3467 9923
rect 3463 9914 3467 9918
rect 3463 9909 3467 9913
rect 3463 9904 3467 9908
rect 3463 9899 3467 9903
rect 3463 9894 3467 9898
rect 3463 9889 3467 9893
rect 3463 9884 3467 9888
rect 3463 9879 3467 9883
rect 3463 9874 3467 9878
rect 3463 9869 3467 9873
rect 3463 9864 3467 9868
rect 3399 9859 3403 9863
rect 3463 9859 3467 9863
rect 3399 9852 3403 9856
rect 3406 9852 3410 9856
rect 3411 9852 3415 9856
rect 3416 9852 3420 9856
rect 3421 9852 3425 9856
rect 3426 9852 3430 9856
rect 3431 9852 3435 9856
rect 3436 9852 3440 9856
rect 3441 9852 3445 9856
rect 3446 9852 3450 9856
rect 3451 9852 3455 9856
rect 3456 9852 3460 9856
rect 3463 9852 3467 9856
rect 3535 9974 3539 9978
rect 3540 9974 3544 9978
rect 3545 9974 3549 9978
rect 3550 9974 3554 9978
rect 3555 9974 3559 9978
rect 3560 9974 3564 9978
rect 3565 9974 3569 9978
rect 3570 9974 3574 9978
rect 3575 9974 3579 9978
rect 3580 9974 3584 9978
rect 3585 9974 3589 9978
rect 3590 9974 3594 9978
rect 3595 9974 3599 9978
rect 3600 9974 3604 9978
rect 3605 9974 3609 9978
rect 3610 9974 3614 9978
rect 3615 9974 3619 9978
rect 3620 9974 3624 9978
rect 3625 9974 3629 9978
rect 3535 9969 3539 9973
rect 3535 9964 3539 9968
rect 3625 9969 3629 9973
rect 3535 9959 3539 9963
rect 3535 9954 3539 9958
rect 3535 9949 3539 9953
rect 3535 9944 3539 9948
rect 3535 9939 3539 9943
rect 3535 9934 3539 9938
rect 3535 9929 3539 9933
rect 3535 9924 3539 9928
rect 3535 9919 3539 9923
rect 3535 9914 3539 9918
rect 3535 9909 3539 9913
rect 3535 9904 3539 9908
rect 3535 9899 3539 9903
rect 3535 9894 3539 9898
rect 3535 9889 3539 9893
rect 3535 9884 3539 9888
rect 3535 9879 3539 9883
rect 3535 9874 3539 9878
rect 3535 9869 3539 9873
rect 3535 9864 3539 9868
rect 3535 9859 3539 9863
rect 3535 9854 3539 9858
rect 3535 9849 3539 9853
rect 3625 9964 3629 9968
rect 3625 9959 3629 9963
rect 3625 9954 3629 9958
rect 3625 9949 3629 9953
rect 3625 9944 3629 9948
rect 3625 9939 3629 9943
rect 3625 9934 3629 9938
rect 3625 9929 3629 9933
rect 3625 9924 3629 9928
rect 3625 9919 3629 9923
rect 3625 9914 3629 9918
rect 3625 9909 3629 9913
rect 3625 9904 3629 9908
rect 3625 9899 3629 9903
rect 3625 9894 3629 9898
rect 3625 9889 3629 9893
rect 3625 9884 3629 9888
rect 3625 9879 3629 9883
rect 3625 9874 3629 9878
rect 3625 9869 3629 9873
rect 3625 9864 3629 9868
rect 3625 9859 3629 9863
rect 3625 9854 3629 9858
rect 3535 9844 3539 9848
rect 3625 9849 3629 9853
rect 3625 9844 3629 9848
rect 3535 9839 3539 9843
rect 3540 9839 3544 9843
rect 3545 9839 3549 9843
rect 3550 9839 3554 9843
rect 3555 9839 3559 9843
rect 3560 9839 3564 9843
rect 3565 9839 3569 9843
rect 3570 9839 3574 9843
rect 3575 9839 3579 9843
rect 3580 9839 3584 9843
rect 3585 9839 3589 9843
rect 3590 9839 3594 9843
rect 3595 9839 3599 9843
rect 3600 9839 3604 9843
rect 3605 9839 3609 9843
rect 3610 9839 3614 9843
rect 3615 9839 3619 9843
rect 3620 9839 3624 9843
rect 3625 9839 3629 9843
rect 3708 9961 3712 9965
rect 3715 9961 3719 9965
rect 3720 9961 3724 9965
rect 3725 9961 3729 9965
rect 3730 9961 3734 9965
rect 3735 9961 3739 9965
rect 3740 9961 3744 9965
rect 3745 9961 3749 9965
rect 3750 9961 3754 9965
rect 3755 9961 3759 9965
rect 3760 9961 3764 9965
rect 3765 9961 3769 9965
rect 3772 9961 3776 9965
rect 3708 9954 3712 9958
rect 3772 9954 3776 9958
rect 3708 9949 3712 9953
rect 3708 9944 3712 9948
rect 3708 9939 3712 9943
rect 3708 9934 3712 9938
rect 3708 9929 3712 9933
rect 3708 9924 3712 9928
rect 3708 9919 3712 9923
rect 3708 9914 3712 9918
rect 3708 9909 3712 9913
rect 3708 9904 3712 9908
rect 3708 9899 3712 9903
rect 3708 9894 3712 9898
rect 3708 9889 3712 9893
rect 3708 9884 3712 9888
rect 3708 9879 3712 9883
rect 3708 9874 3712 9878
rect 3708 9869 3712 9873
rect 3708 9864 3712 9868
rect 3772 9949 3776 9953
rect 3772 9944 3776 9948
rect 3772 9939 3776 9943
rect 3772 9934 3776 9938
rect 3772 9929 3776 9933
rect 3772 9924 3776 9928
rect 3772 9919 3776 9923
rect 3772 9914 3776 9918
rect 3772 9909 3776 9913
rect 3772 9904 3776 9908
rect 3772 9899 3776 9903
rect 3772 9894 3776 9898
rect 3772 9889 3776 9893
rect 3772 9884 3776 9888
rect 3772 9879 3776 9883
rect 3772 9874 3776 9878
rect 3772 9869 3776 9873
rect 3772 9864 3776 9868
rect 3708 9859 3712 9863
rect 3772 9859 3776 9863
rect 3708 9852 3712 9856
rect 3715 9852 3719 9856
rect 3720 9852 3724 9856
rect 3725 9852 3729 9856
rect 3730 9852 3734 9856
rect 3735 9852 3739 9856
rect 3740 9852 3744 9856
rect 3745 9852 3749 9856
rect 3750 9852 3754 9856
rect 3755 9852 3759 9856
rect 3760 9852 3764 9856
rect 3765 9852 3769 9856
rect 3772 9852 3776 9856
rect 3844 9974 3848 9978
rect 3849 9974 3853 9978
rect 3854 9974 3858 9978
rect 3859 9974 3863 9978
rect 3864 9974 3868 9978
rect 3869 9974 3873 9978
rect 3874 9974 3878 9978
rect 3879 9974 3883 9978
rect 3884 9974 3888 9978
rect 3889 9974 3893 9978
rect 3894 9974 3898 9978
rect 3899 9974 3903 9978
rect 3904 9974 3908 9978
rect 3909 9974 3913 9978
rect 3914 9974 3918 9978
rect 3919 9974 3923 9978
rect 3924 9974 3928 9978
rect 3929 9974 3933 9978
rect 3934 9974 3938 9978
rect 3844 9969 3848 9973
rect 3844 9964 3848 9968
rect 3934 9969 3938 9973
rect 3844 9959 3848 9963
rect 3844 9954 3848 9958
rect 3844 9949 3848 9953
rect 3844 9944 3848 9948
rect 3844 9939 3848 9943
rect 3844 9934 3848 9938
rect 3844 9929 3848 9933
rect 3844 9924 3848 9928
rect 3844 9919 3848 9923
rect 3844 9914 3848 9918
rect 3844 9909 3848 9913
rect 3844 9904 3848 9908
rect 3844 9899 3848 9903
rect 3844 9894 3848 9898
rect 3844 9889 3848 9893
rect 3844 9884 3848 9888
rect 3844 9879 3848 9883
rect 3844 9874 3848 9878
rect 3844 9869 3848 9873
rect 3844 9864 3848 9868
rect 3844 9859 3848 9863
rect 3844 9854 3848 9858
rect 3844 9849 3848 9853
rect 3934 9964 3938 9968
rect 3934 9959 3938 9963
rect 3934 9954 3938 9958
rect 3934 9949 3938 9953
rect 3934 9944 3938 9948
rect 3934 9939 3938 9943
rect 3934 9934 3938 9938
rect 3934 9929 3938 9933
rect 3934 9924 3938 9928
rect 3934 9919 3938 9923
rect 3934 9914 3938 9918
rect 3934 9909 3938 9913
rect 3934 9904 3938 9908
rect 3934 9899 3938 9903
rect 3934 9894 3938 9898
rect 3934 9889 3938 9893
rect 3934 9884 3938 9888
rect 3934 9879 3938 9883
rect 3934 9874 3938 9878
rect 3934 9869 3938 9873
rect 3934 9864 3938 9868
rect 3934 9859 3938 9863
rect 3934 9854 3938 9858
rect 3844 9844 3848 9848
rect 3934 9849 3938 9853
rect 3934 9844 3938 9848
rect 3844 9839 3848 9843
rect 3849 9839 3853 9843
rect 3854 9839 3858 9843
rect 3859 9839 3863 9843
rect 3864 9839 3868 9843
rect 3869 9839 3873 9843
rect 3874 9839 3878 9843
rect 3879 9839 3883 9843
rect 3884 9839 3888 9843
rect 3889 9839 3893 9843
rect 3894 9839 3898 9843
rect 3899 9839 3903 9843
rect 3904 9839 3908 9843
rect 3909 9839 3913 9843
rect 3914 9839 3918 9843
rect 3919 9839 3923 9843
rect 3924 9839 3928 9843
rect 3929 9839 3933 9843
rect 3934 9839 3938 9843
rect 4017 9961 4021 9965
rect 4024 9961 4028 9965
rect 4029 9961 4033 9965
rect 4034 9961 4038 9965
rect 4039 9961 4043 9965
rect 4044 9961 4048 9965
rect 4049 9961 4053 9965
rect 4054 9961 4058 9965
rect 4059 9961 4063 9965
rect 4064 9961 4068 9965
rect 4069 9961 4073 9965
rect 4074 9961 4078 9965
rect 4081 9961 4085 9965
rect 4017 9954 4021 9958
rect 4081 9954 4085 9958
rect 4017 9949 4021 9953
rect 4017 9944 4021 9948
rect 4017 9939 4021 9943
rect 4017 9934 4021 9938
rect 4017 9929 4021 9933
rect 4017 9924 4021 9928
rect 4017 9919 4021 9923
rect 4017 9914 4021 9918
rect 4017 9909 4021 9913
rect 4017 9904 4021 9908
rect 4017 9899 4021 9903
rect 4017 9894 4021 9898
rect 4017 9889 4021 9893
rect 4017 9884 4021 9888
rect 4017 9879 4021 9883
rect 4017 9874 4021 9878
rect 4017 9869 4021 9873
rect 4017 9864 4021 9868
rect 4081 9949 4085 9953
rect 4081 9944 4085 9948
rect 4081 9939 4085 9943
rect 4081 9934 4085 9938
rect 4081 9929 4085 9933
rect 4081 9924 4085 9928
rect 4081 9919 4085 9923
rect 4081 9914 4085 9918
rect 4081 9909 4085 9913
rect 4081 9904 4085 9908
rect 4081 9899 4085 9903
rect 4081 9894 4085 9898
rect 4081 9889 4085 9893
rect 4081 9884 4085 9888
rect 4081 9879 4085 9883
rect 4081 9874 4085 9878
rect 4081 9869 4085 9873
rect 4081 9864 4085 9868
rect 4017 9859 4021 9863
rect 4081 9859 4085 9863
rect 4017 9852 4021 9856
rect 4024 9852 4028 9856
rect 4029 9852 4033 9856
rect 4034 9852 4038 9856
rect 4039 9852 4043 9856
rect 4044 9852 4048 9856
rect 4049 9852 4053 9856
rect 4054 9852 4058 9856
rect 4059 9852 4063 9856
rect 4064 9852 4068 9856
rect 4069 9852 4073 9856
rect 4074 9852 4078 9856
rect 4081 9852 4085 9856
rect 802 9762 806 9766
rect 807 9762 811 9766
rect 812 9762 816 9766
rect 817 9762 821 9766
rect 831 9762 835 9766
rect 836 9762 840 9766
rect 841 9762 845 9766
rect 846 9762 850 9766
rect 860 9762 864 9766
rect 865 9762 869 9766
rect 870 9762 874 9766
rect 875 9762 879 9766
rect 889 9762 893 9766
rect 894 9762 898 9766
rect 899 9762 903 9766
rect 904 9762 908 9766
rect 918 9762 922 9766
rect 923 9762 927 9766
rect 928 9762 932 9766
rect 933 9762 937 9766
rect 1319 9762 1323 9766
rect 1324 9762 1328 9766
rect 1329 9762 1333 9766
rect 1334 9762 1338 9766
rect 1628 9762 1632 9766
rect 1633 9762 1637 9766
rect 1638 9762 1642 9766
rect 1643 9762 1647 9766
rect 1937 9762 1941 9766
rect 1942 9762 1946 9766
rect 1947 9762 1951 9766
rect 1952 9762 1956 9766
rect 2246 9762 2250 9766
rect 2251 9762 2255 9766
rect 2256 9762 2260 9766
rect 2261 9762 2265 9766
rect 2555 9762 2559 9766
rect 2560 9762 2564 9766
rect 2565 9762 2569 9766
rect 2570 9762 2574 9766
rect 2864 9762 2868 9766
rect 2869 9762 2873 9766
rect 2874 9762 2878 9766
rect 2879 9762 2883 9766
rect 3173 9762 3177 9766
rect 3178 9762 3182 9766
rect 3183 9762 3187 9766
rect 3188 9762 3192 9766
rect 3482 9762 3486 9766
rect 3487 9762 3491 9766
rect 3492 9762 3496 9766
rect 3497 9762 3501 9766
rect 3791 9762 3795 9766
rect 3796 9762 3800 9766
rect 3801 9762 3805 9766
rect 3806 9762 3810 9766
rect 4100 9762 4104 9766
rect 4105 9762 4109 9766
rect 4110 9762 4114 9766
rect 4115 9762 4119 9766
rect 4292 9762 4296 9766
rect 4297 9762 4301 9766
rect 4302 9762 4306 9766
rect 4307 9762 4311 9766
rect 4318 9762 4322 9766
rect 4323 9762 4327 9766
rect 4328 9762 4332 9766
rect 4333 9762 4337 9766
rect 4344 9762 4348 9766
rect 4349 9762 4353 9766
rect 4354 9762 4358 9766
rect 4359 9762 4363 9766
rect 4370 9762 4374 9766
rect 4375 9762 4379 9766
rect 4380 9762 4384 9766
rect 4385 9762 4389 9766
rect 4396 9762 4400 9766
rect 4401 9762 4405 9766
rect 4406 9762 4410 9766
rect 4411 9762 4415 9766
rect 802 9752 806 9756
rect 807 9752 811 9756
rect 812 9752 816 9756
rect 817 9752 821 9756
rect 831 9752 835 9756
rect 836 9752 840 9756
rect 841 9752 845 9756
rect 846 9752 850 9756
rect 860 9752 864 9756
rect 865 9752 869 9756
rect 870 9752 874 9756
rect 875 9752 879 9756
rect 889 9752 893 9756
rect 894 9752 898 9756
rect 899 9752 903 9756
rect 904 9752 908 9756
rect 918 9752 922 9756
rect 923 9752 927 9756
rect 928 9752 932 9756
rect 933 9752 937 9756
rect 1319 9752 1323 9756
rect 1324 9752 1328 9756
rect 1329 9752 1333 9756
rect 1334 9752 1338 9756
rect 1628 9752 1632 9756
rect 1633 9752 1637 9756
rect 1638 9752 1642 9756
rect 1643 9752 1647 9756
rect 1937 9752 1941 9756
rect 1942 9752 1946 9756
rect 1947 9752 1951 9756
rect 1952 9752 1956 9756
rect 2246 9752 2250 9756
rect 2251 9752 2255 9756
rect 2256 9752 2260 9756
rect 2261 9752 2265 9756
rect 2555 9752 2559 9756
rect 2560 9752 2564 9756
rect 2565 9752 2569 9756
rect 2570 9752 2574 9756
rect 2864 9752 2868 9756
rect 2869 9752 2873 9756
rect 2874 9752 2878 9756
rect 2879 9752 2883 9756
rect 3173 9752 3177 9756
rect 3178 9752 3182 9756
rect 3183 9752 3187 9756
rect 3188 9752 3192 9756
rect 3482 9752 3486 9756
rect 3487 9752 3491 9756
rect 3492 9752 3496 9756
rect 3497 9752 3501 9756
rect 3791 9752 3795 9756
rect 3796 9752 3800 9756
rect 3801 9752 3805 9756
rect 3806 9752 3810 9756
rect 4100 9752 4104 9756
rect 4105 9752 4109 9756
rect 4110 9752 4114 9756
rect 4115 9752 4119 9756
rect 4292 9752 4296 9756
rect 4297 9752 4301 9756
rect 4302 9752 4306 9756
rect 4307 9752 4311 9756
rect 4318 9752 4322 9756
rect 4323 9752 4327 9756
rect 4328 9752 4332 9756
rect 4333 9752 4337 9756
rect 4344 9752 4348 9756
rect 4349 9752 4353 9756
rect 4354 9752 4358 9756
rect 4359 9752 4363 9756
rect 4370 9752 4374 9756
rect 4375 9752 4379 9756
rect 4380 9752 4384 9756
rect 4385 9752 4389 9756
rect 4396 9752 4400 9756
rect 4401 9752 4405 9756
rect 4406 9752 4410 9756
rect 4411 9752 4415 9756
rect 802 9742 806 9746
rect 807 9742 811 9746
rect 812 9742 816 9746
rect 817 9742 821 9746
rect 831 9742 835 9746
rect 836 9742 840 9746
rect 841 9742 845 9746
rect 846 9742 850 9746
rect 860 9742 864 9746
rect 865 9742 869 9746
rect 870 9742 874 9746
rect 875 9742 879 9746
rect 889 9742 893 9746
rect 894 9742 898 9746
rect 899 9742 903 9746
rect 904 9742 908 9746
rect 918 9742 922 9746
rect 923 9742 927 9746
rect 928 9742 932 9746
rect 933 9742 937 9746
rect 1319 9742 1323 9746
rect 1324 9742 1328 9746
rect 1329 9742 1333 9746
rect 1334 9742 1338 9746
rect 1628 9742 1632 9746
rect 1633 9742 1637 9746
rect 1638 9742 1642 9746
rect 1643 9742 1647 9746
rect 1937 9742 1941 9746
rect 1942 9742 1946 9746
rect 1947 9742 1951 9746
rect 1952 9742 1956 9746
rect 2246 9742 2250 9746
rect 2251 9742 2255 9746
rect 2256 9742 2260 9746
rect 2261 9742 2265 9746
rect 2555 9742 2559 9746
rect 2560 9742 2564 9746
rect 2565 9742 2569 9746
rect 2570 9742 2574 9746
rect 2864 9742 2868 9746
rect 2869 9742 2873 9746
rect 2874 9742 2878 9746
rect 2879 9742 2883 9746
rect 3173 9742 3177 9746
rect 3178 9742 3182 9746
rect 3183 9742 3187 9746
rect 3188 9742 3192 9746
rect 3482 9742 3486 9746
rect 3487 9742 3491 9746
rect 3492 9742 3496 9746
rect 3497 9742 3501 9746
rect 3791 9742 3795 9746
rect 3796 9742 3800 9746
rect 3801 9742 3805 9746
rect 3806 9742 3810 9746
rect 4100 9742 4104 9746
rect 4105 9742 4109 9746
rect 4110 9742 4114 9746
rect 4115 9742 4119 9746
rect 4292 9742 4296 9746
rect 4297 9742 4301 9746
rect 4302 9742 4306 9746
rect 4307 9742 4311 9746
rect 4318 9742 4322 9746
rect 4323 9742 4327 9746
rect 4328 9742 4332 9746
rect 4333 9742 4337 9746
rect 4344 9742 4348 9746
rect 4349 9742 4353 9746
rect 4354 9742 4358 9746
rect 4359 9742 4363 9746
rect 4370 9742 4374 9746
rect 4375 9742 4379 9746
rect 4380 9742 4384 9746
rect 4385 9742 4389 9746
rect 4396 9742 4400 9746
rect 4401 9742 4405 9746
rect 4406 9742 4410 9746
rect 4411 9742 4415 9746
rect 802 9732 806 9736
rect 807 9732 811 9736
rect 812 9732 816 9736
rect 817 9732 821 9736
rect 831 9732 835 9736
rect 836 9732 840 9736
rect 841 9732 845 9736
rect 846 9732 850 9736
rect 860 9732 864 9736
rect 865 9732 869 9736
rect 870 9732 874 9736
rect 875 9732 879 9736
rect 889 9732 893 9736
rect 894 9732 898 9736
rect 899 9732 903 9736
rect 904 9732 908 9736
rect 918 9732 922 9736
rect 923 9732 927 9736
rect 928 9732 932 9736
rect 933 9732 937 9736
rect 1319 9732 1323 9736
rect 1324 9732 1328 9736
rect 1329 9732 1333 9736
rect 1334 9732 1338 9736
rect 1628 9732 1632 9736
rect 1633 9732 1637 9736
rect 1638 9732 1642 9736
rect 1643 9732 1647 9736
rect 1937 9732 1941 9736
rect 1942 9732 1946 9736
rect 1947 9732 1951 9736
rect 1952 9732 1956 9736
rect 2246 9732 2250 9736
rect 2251 9732 2255 9736
rect 2256 9732 2260 9736
rect 2261 9732 2265 9736
rect 2555 9732 2559 9736
rect 2560 9732 2564 9736
rect 2565 9732 2569 9736
rect 2570 9732 2574 9736
rect 2864 9732 2868 9736
rect 2869 9732 2873 9736
rect 2874 9732 2878 9736
rect 2879 9732 2883 9736
rect 3173 9732 3177 9736
rect 3178 9732 3182 9736
rect 3183 9732 3187 9736
rect 3188 9732 3192 9736
rect 3482 9732 3486 9736
rect 3487 9732 3491 9736
rect 3492 9732 3496 9736
rect 3497 9732 3501 9736
rect 3791 9732 3795 9736
rect 3796 9732 3800 9736
rect 3801 9732 3805 9736
rect 3806 9732 3810 9736
rect 4100 9732 4104 9736
rect 4105 9732 4109 9736
rect 4110 9732 4114 9736
rect 4115 9732 4119 9736
rect 4292 9732 4296 9736
rect 4297 9732 4301 9736
rect 4302 9732 4306 9736
rect 4307 9732 4311 9736
rect 4318 9732 4322 9736
rect 4323 9732 4327 9736
rect 4328 9732 4332 9736
rect 4333 9732 4337 9736
rect 4344 9732 4348 9736
rect 4349 9732 4353 9736
rect 4354 9732 4358 9736
rect 4359 9732 4363 9736
rect 4370 9732 4374 9736
rect 4375 9732 4379 9736
rect 4380 9732 4384 9736
rect 4385 9732 4389 9736
rect 4396 9732 4400 9736
rect 4401 9732 4405 9736
rect 4406 9732 4410 9736
rect 4411 9732 4415 9736
rect 613 9618 617 9622
rect 623 9618 627 9622
rect 633 9618 637 9622
rect 643 9618 647 9622
rect 613 9613 617 9617
rect 623 9613 627 9617
rect 633 9613 637 9617
rect 643 9613 647 9617
rect 613 9608 617 9612
rect 623 9608 627 9612
rect 633 9608 637 9612
rect 643 9608 647 9612
rect 613 9603 617 9607
rect 623 9603 627 9607
rect 633 9603 637 9607
rect 643 9603 647 9607
rect 613 9592 617 9596
rect 623 9592 627 9596
rect 633 9592 637 9596
rect 643 9592 647 9596
rect 613 9587 617 9591
rect 623 9587 627 9591
rect 633 9587 637 9591
rect 643 9587 647 9591
rect 613 9582 617 9586
rect 623 9582 627 9586
rect 633 9582 637 9586
rect 643 9582 647 9586
rect 613 9577 617 9581
rect 623 9577 627 9581
rect 633 9577 637 9581
rect 643 9577 647 9581
rect 613 9566 617 9570
rect 623 9566 627 9570
rect 633 9566 637 9570
rect 643 9566 647 9570
rect 613 9561 617 9565
rect 623 9561 627 9565
rect 633 9561 637 9565
rect 643 9561 647 9565
rect 613 9556 617 9560
rect 623 9556 627 9560
rect 633 9556 637 9560
rect 643 9556 647 9560
rect 613 9551 617 9555
rect 623 9551 627 9555
rect 633 9551 637 9555
rect 643 9551 647 9555
rect 613 9540 617 9544
rect 623 9540 627 9544
rect 633 9540 637 9544
rect 643 9540 647 9544
rect 613 9535 617 9539
rect 623 9535 627 9539
rect 633 9535 637 9539
rect 643 9535 647 9539
rect 613 9530 617 9534
rect 623 9530 627 9534
rect 633 9530 637 9534
rect 643 9530 647 9534
rect 613 9525 617 9529
rect 623 9525 627 9529
rect 633 9525 637 9529
rect 643 9525 647 9529
rect 613 9514 617 9518
rect 623 9514 627 9518
rect 633 9514 637 9518
rect 643 9514 647 9518
rect 613 9509 617 9513
rect 623 9509 627 9513
rect 633 9509 637 9513
rect 643 9509 647 9513
rect 613 9504 617 9508
rect 623 9504 627 9508
rect 633 9504 637 9508
rect 643 9504 647 9508
rect 613 9499 617 9503
rect 623 9499 627 9503
rect 633 9499 637 9503
rect 643 9499 647 9503
rect 613 9321 617 9325
rect 623 9321 627 9325
rect 633 9321 637 9325
rect 643 9321 647 9325
rect 613 9316 617 9320
rect 623 9316 627 9320
rect 633 9316 637 9320
rect 643 9316 647 9320
rect 613 9311 617 9315
rect 623 9311 627 9315
rect 633 9311 637 9315
rect 643 9311 647 9315
rect 613 9306 617 9310
rect 623 9306 627 9310
rect 633 9306 637 9310
rect 643 9306 647 9310
rect 613 9012 617 9016
rect 623 9012 627 9016
rect 633 9012 637 9016
rect 643 9012 647 9016
rect 613 9007 617 9011
rect 623 9007 627 9011
rect 633 9007 637 9011
rect 643 9007 647 9011
rect 613 9002 617 9006
rect 623 9002 627 9006
rect 633 9002 637 9006
rect 643 9002 647 9006
rect 613 8997 617 9001
rect 623 8997 627 9001
rect 633 8997 637 9001
rect 643 8997 647 9001
rect 613 8703 617 8707
rect 623 8703 627 8707
rect 633 8703 637 8707
rect 643 8703 647 8707
rect 613 8698 617 8702
rect 623 8698 627 8702
rect 633 8698 637 8702
rect 643 8698 647 8702
rect 613 8693 617 8697
rect 623 8693 627 8697
rect 633 8693 637 8697
rect 643 8693 647 8697
rect 613 8688 617 8692
rect 623 8688 627 8692
rect 633 8688 637 8692
rect 643 8688 647 8692
rect 613 8394 617 8398
rect 623 8394 627 8398
rect 633 8394 637 8398
rect 643 8394 647 8398
rect 613 8389 617 8393
rect 623 8389 627 8393
rect 633 8389 637 8393
rect 643 8389 647 8393
rect 613 8384 617 8388
rect 623 8384 627 8388
rect 633 8384 637 8388
rect 643 8384 647 8388
rect 613 8379 617 8383
rect 623 8379 627 8383
rect 633 8379 637 8383
rect 643 8379 647 8383
rect 613 8085 617 8089
rect 623 8085 627 8089
rect 633 8085 637 8089
rect 643 8085 647 8089
rect 613 8080 617 8084
rect 623 8080 627 8084
rect 633 8080 637 8084
rect 643 8080 647 8084
rect 613 8075 617 8079
rect 623 8075 627 8079
rect 633 8075 637 8079
rect 643 8075 647 8079
rect 613 8070 617 8074
rect 623 8070 627 8074
rect 633 8070 637 8074
rect 643 8070 647 8074
rect 613 7776 617 7780
rect 623 7776 627 7780
rect 633 7776 637 7780
rect 643 7776 647 7780
rect 613 7771 617 7775
rect 623 7771 627 7775
rect 633 7771 637 7775
rect 643 7771 647 7775
rect 613 7766 617 7770
rect 623 7766 627 7770
rect 633 7766 637 7770
rect 643 7766 647 7770
rect 613 7761 617 7765
rect 623 7761 627 7765
rect 633 7761 637 7765
rect 643 7761 647 7765
rect 613 7467 617 7471
rect 623 7467 627 7471
rect 633 7467 637 7471
rect 643 7467 647 7471
rect 613 7462 617 7466
rect 623 7462 627 7466
rect 633 7462 637 7466
rect 643 7462 647 7466
rect 613 7457 617 7461
rect 623 7457 627 7461
rect 633 7457 637 7461
rect 643 7457 647 7461
rect 613 7452 617 7456
rect 623 7452 627 7456
rect 633 7452 637 7456
rect 643 7452 647 7456
rect 613 7158 617 7162
rect 623 7158 627 7162
rect 633 7158 637 7162
rect 643 7158 647 7162
rect 613 7153 617 7157
rect 623 7153 627 7157
rect 633 7153 637 7157
rect 643 7153 647 7157
rect 613 7148 617 7152
rect 623 7148 627 7152
rect 633 7148 637 7152
rect 643 7148 647 7152
rect 613 7143 617 7147
rect 623 7143 627 7147
rect 633 7143 637 7147
rect 643 7143 647 7147
rect 613 6849 617 6853
rect 623 6849 627 6853
rect 633 6849 637 6853
rect 643 6849 647 6853
rect 613 6844 617 6848
rect 623 6844 627 6848
rect 633 6844 637 6848
rect 643 6844 647 6848
rect 613 6839 617 6843
rect 623 6839 627 6843
rect 633 6839 637 6843
rect 643 6839 647 6843
rect 613 6834 617 6838
rect 623 6834 627 6838
rect 633 6834 637 6838
rect 643 6834 647 6838
rect 613 6540 617 6544
rect 623 6540 627 6544
rect 633 6540 637 6544
rect 643 6540 647 6544
rect 613 6535 617 6539
rect 623 6535 627 6539
rect 633 6535 637 6539
rect 643 6535 647 6539
rect 613 6530 617 6534
rect 623 6530 627 6534
rect 633 6530 637 6534
rect 643 6530 647 6534
rect 613 6525 617 6529
rect 623 6525 627 6529
rect 633 6525 637 6529
rect 643 6525 647 6529
rect 613 6140 617 6144
rect 623 6140 627 6144
rect 633 6140 637 6144
rect 643 6140 647 6144
rect 613 6135 617 6139
rect 623 6135 627 6139
rect 633 6135 637 6139
rect 643 6135 647 6139
rect 613 6130 617 6134
rect 623 6130 627 6134
rect 633 6130 637 6134
rect 643 6130 647 6134
rect 613 6125 617 6129
rect 623 6125 627 6129
rect 633 6125 637 6129
rect 643 6125 647 6129
rect 613 6111 617 6115
rect 623 6111 627 6115
rect 633 6111 637 6115
rect 643 6111 647 6115
rect 613 6106 617 6110
rect 623 6106 627 6110
rect 633 6106 637 6110
rect 643 6106 647 6110
rect 613 6101 617 6105
rect 623 6101 627 6105
rect 633 6101 637 6105
rect 643 6101 647 6105
rect 613 6096 617 6100
rect 623 6096 627 6100
rect 633 6096 637 6100
rect 643 6096 647 6100
rect 613 6082 617 6086
rect 623 6082 627 6086
rect 633 6082 637 6086
rect 643 6082 647 6086
rect 613 6077 617 6081
rect 623 6077 627 6081
rect 633 6077 637 6081
rect 643 6077 647 6081
rect 613 6072 617 6076
rect 623 6072 627 6076
rect 633 6072 637 6076
rect 643 6072 647 6076
rect 613 6067 617 6071
rect 623 6067 627 6071
rect 633 6067 637 6071
rect 643 6067 647 6071
rect 613 6053 617 6057
rect 623 6053 627 6057
rect 633 6053 637 6057
rect 643 6053 647 6057
rect 613 6048 617 6052
rect 623 6048 627 6052
rect 633 6048 637 6052
rect 643 6048 647 6052
rect 613 6043 617 6047
rect 623 6043 627 6047
rect 633 6043 637 6047
rect 643 6043 647 6047
rect 613 6038 617 6042
rect 623 6038 627 6042
rect 633 6038 637 6042
rect 643 6038 647 6042
rect 613 6024 617 6028
rect 623 6024 627 6028
rect 633 6024 637 6028
rect 643 6024 647 6028
rect 613 6019 617 6023
rect 623 6019 627 6023
rect 633 6019 637 6023
rect 643 6019 647 6023
rect 613 6014 617 6018
rect 623 6014 627 6018
rect 633 6014 637 6018
rect 643 6014 647 6018
rect 613 6009 617 6013
rect 623 6009 627 6013
rect 633 6009 637 6013
rect 643 6009 647 6013
rect 2881 9340 2885 9344
rect 2909 9340 2913 9344
rect 2939 9340 2943 9344
rect 2976 9340 2980 9344
rect 3013 9340 3017 9344
rect 3041 9340 3045 9344
rect 3071 9340 3075 9344
rect 3108 9340 3112 9344
rect 3145 9340 3149 9344
rect 3173 9340 3177 9344
rect 3203 9340 3207 9344
rect 3240 9340 3244 9344
rect 3277 9340 3281 9344
rect 3305 9340 3309 9344
rect 3335 9340 3339 9344
rect 3372 9340 3376 9344
rect 3826 9340 3830 9344
rect 3854 9340 3858 9344
rect 3884 9340 3888 9344
rect 3921 9340 3925 9344
rect 3958 9340 3962 9344
rect 3986 9340 3990 9344
rect 4016 9340 4020 9344
rect 4053 9340 4057 9344
rect 4090 9340 4094 9344
rect 4118 9340 4122 9344
rect 4148 9340 4152 9344
rect 4185 9340 4189 9344
rect 4222 9340 4226 9344
rect 4250 9340 4254 9344
rect 4280 9340 4284 9344
rect 4317 9340 4321 9344
rect 2529 9307 2533 9311
rect 2557 9307 2561 9311
rect 2587 9307 2591 9311
rect 2624 9307 2628 9311
rect 3474 9307 3478 9311
rect 3502 9307 3506 9311
rect 3532 9307 3536 9311
rect 3569 9307 3573 9311
rect 2871 9263 2875 9267
rect 2900 9263 2904 9267
rect 2925 9263 2929 9267
rect 2967 9263 2971 9267
rect 3023 9263 3027 9267
rect 3047 9263 3051 9267
rect 3101 9263 3105 9267
rect 3128 9263 3132 9267
rect 3182 9263 3186 9267
rect 3816 9263 3820 9267
rect 3845 9263 3849 9267
rect 3870 9263 3874 9267
rect 3912 9263 3916 9267
rect 3968 9263 3972 9267
rect 3992 9263 3996 9267
rect 4046 9263 4050 9267
rect 4073 9263 4077 9267
rect 4127 9263 4131 9267
rect 2489 9205 2493 9209
rect 2526 9205 2530 9209
rect 2556 9205 2560 9209
rect 2584 9205 2588 9209
rect 3434 9205 3438 9209
rect 3471 9205 3475 9209
rect 3501 9205 3505 9209
rect 3529 9205 3533 9209
rect 2871 9131 2875 9135
rect 2900 9131 2904 9135
rect 2925 9131 2929 9135
rect 2967 9131 2971 9135
rect 3023 9131 3027 9135
rect 3047 9131 3051 9135
rect 3101 9131 3105 9135
rect 3128 9131 3132 9135
rect 3190 9131 3194 9135
rect 3816 9131 3820 9135
rect 3845 9131 3849 9135
rect 3870 9131 3874 9135
rect 3912 9131 3916 9135
rect 3968 9131 3972 9135
rect 3992 9131 3996 9135
rect 4046 9131 4050 9135
rect 4073 9131 4077 9135
rect 4135 9131 4139 9135
rect 3359 9102 3363 9106
rect 3383 9102 3387 9106
rect 3437 9102 3441 9106
rect 3580 9102 3584 9106
rect 2871 8999 2875 9003
rect 2900 8999 2904 9003
rect 2925 8999 2929 9003
rect 2967 8999 2971 9003
rect 3023 8999 3027 9003
rect 3047 8999 3051 9003
rect 3101 8999 3105 9003
rect 3128 8999 3132 9003
rect 3182 8999 3186 9003
rect 3190 8999 3194 9003
rect 3218 8999 3222 9003
rect 3272 8999 3276 9003
rect 3816 8999 3820 9003
rect 3845 8999 3849 9003
rect 3870 8999 3874 9003
rect 3912 8999 3916 9003
rect 3968 8999 3972 9003
rect 3992 8999 3996 9003
rect 4046 8999 4050 9003
rect 4073 8999 4077 9003
rect 4127 8999 4131 9003
rect 4135 8999 4139 9003
rect 4163 8999 4167 9003
rect 4217 8999 4221 9003
rect 3337 8972 3341 8976
rect 3359 8972 3363 8976
rect 3383 8972 3387 8976
rect 3437 8972 3441 8976
rect 3486 8972 3490 8976
rect 2871 8867 2875 8871
rect 2900 8867 2904 8871
rect 2925 8867 2929 8871
rect 2967 8867 2971 8871
rect 3023 8867 3027 8871
rect 3047 8867 3051 8871
rect 3101 8867 3105 8871
rect 3128 8867 3132 8871
rect 3218 8867 3222 8871
rect 3816 8867 3820 8871
rect 3845 8867 3849 8871
rect 3870 8867 3874 8871
rect 3912 8867 3916 8871
rect 3968 8867 3972 8871
rect 3992 8867 3996 8871
rect 4046 8867 4050 8871
rect 4073 8867 4077 8871
rect 4163 8867 4167 8871
rect 3383 8842 3387 8846
rect 2397 8805 2401 8809
rect 2425 8805 2429 8809
rect 2455 8805 2459 8809
rect 2492 8805 2496 8809
rect 2529 8805 2533 8809
rect 2557 8805 2561 8809
rect 2587 8805 2591 8809
rect 2624 8805 2628 8809
rect 2661 8805 2665 8809
rect 2689 8805 2693 8809
rect 2719 8805 2723 8809
rect 2756 8805 2760 8809
rect 3342 8805 3346 8809
rect 3370 8805 3374 8809
rect 3400 8805 3404 8809
rect 3437 8805 3441 8809
rect 3474 8805 3478 8809
rect 3502 8805 3506 8809
rect 3532 8805 3536 8809
rect 3569 8805 3573 8809
rect 3606 8805 3610 8809
rect 3634 8805 3638 8809
rect 3664 8805 3668 8809
rect 3701 8805 3705 8809
rect 2871 8735 2875 8739
rect 2900 8735 2904 8739
rect 2925 8735 2929 8739
rect 2967 8735 2971 8739
rect 3047 8735 3051 8739
rect 3101 8735 3105 8739
rect 3132 8735 3136 8739
rect 3161 8735 3165 8739
rect 3186 8735 3190 8739
rect 3228 8735 3232 8739
rect 3816 8735 3820 8739
rect 3845 8735 3849 8739
rect 3870 8735 3874 8739
rect 3912 8735 3916 8739
rect 3992 8735 3996 8739
rect 4046 8735 4050 8739
rect 4077 8735 4081 8739
rect 4106 8735 4110 8739
rect 4131 8735 4135 8739
rect 4173 8735 4177 8739
rect 3180 8693 3184 8697
rect 3208 8693 3212 8697
rect 3238 8693 3242 8697
rect 3275 8693 3279 8697
rect 4125 8693 4129 8697
rect 4153 8693 4157 8697
rect 4183 8693 4187 8697
rect 4220 8693 4224 8697
rect 2397 8663 2401 8667
rect 2425 8663 2429 8667
rect 2455 8663 2459 8667
rect 2492 8663 2496 8667
rect 2529 8663 2533 8667
rect 2557 8663 2561 8667
rect 2587 8663 2591 8667
rect 2624 8663 2628 8667
rect 2661 8663 2665 8667
rect 2689 8663 2693 8667
rect 2719 8663 2723 8667
rect 2756 8663 2760 8667
rect 3342 8663 3346 8667
rect 3370 8663 3374 8667
rect 3400 8663 3404 8667
rect 3437 8663 3441 8667
rect 3474 8663 3478 8667
rect 3502 8663 3506 8667
rect 3532 8663 3536 8667
rect 3569 8663 3573 8667
rect 3606 8663 3610 8667
rect 3634 8663 3638 8667
rect 3664 8663 3668 8667
rect 3701 8663 3705 8667
rect 3180 8607 3184 8611
rect 3208 8607 3212 8611
rect 3238 8607 3242 8611
rect 3275 8607 3279 8611
rect 4125 8607 4129 8611
rect 4153 8607 4157 8611
rect 4183 8607 4187 8611
rect 4220 8607 4224 8611
rect 2397 8577 2401 8581
rect 2425 8577 2429 8581
rect 2455 8577 2459 8581
rect 2492 8577 2496 8581
rect 2529 8577 2533 8581
rect 2557 8577 2561 8581
rect 2587 8577 2591 8581
rect 2624 8577 2628 8581
rect 2661 8577 2665 8581
rect 2689 8577 2693 8581
rect 2719 8577 2723 8581
rect 2756 8577 2760 8581
rect 3342 8577 3346 8581
rect 3370 8577 3374 8581
rect 3400 8577 3404 8581
rect 3437 8577 3441 8581
rect 3474 8577 3478 8581
rect 3502 8577 3506 8581
rect 3532 8577 3536 8581
rect 3569 8577 3573 8581
rect 3606 8577 3610 8581
rect 3634 8577 3638 8581
rect 3664 8577 3668 8581
rect 3701 8577 3705 8581
rect 2397 8437 2401 8441
rect 2425 8437 2429 8441
rect 2455 8437 2459 8441
rect 2492 8437 2496 8441
rect 2529 8437 2533 8441
rect 2557 8437 2561 8441
rect 2587 8437 2591 8441
rect 2624 8437 2628 8441
rect 2661 8437 2665 8441
rect 2689 8437 2693 8441
rect 2719 8437 2723 8441
rect 2756 8437 2760 8441
rect 3342 8437 3346 8441
rect 3370 8437 3374 8441
rect 3400 8437 3404 8441
rect 3437 8437 3441 8441
rect 3474 8437 3478 8441
rect 3502 8437 3506 8441
rect 3532 8437 3536 8441
rect 3569 8437 3573 8441
rect 3606 8437 3610 8441
rect 3634 8437 3638 8441
rect 3664 8437 3668 8441
rect 3701 8437 3705 8441
rect 2881 8358 2885 8362
rect 2909 8358 2913 8362
rect 2939 8358 2943 8362
rect 2976 8358 2980 8362
rect 3013 8358 3017 8362
rect 3041 8358 3045 8362
rect 3071 8358 3075 8362
rect 3108 8358 3112 8362
rect 3145 8358 3149 8362
rect 3173 8358 3177 8362
rect 3203 8358 3207 8362
rect 3240 8358 3244 8362
rect 3277 8358 3281 8362
rect 3305 8358 3309 8362
rect 3335 8358 3339 8362
rect 3372 8358 3376 8362
rect 3826 8358 3830 8362
rect 3854 8358 3858 8362
rect 3884 8358 3888 8362
rect 3921 8358 3925 8362
rect 3958 8358 3962 8362
rect 3986 8358 3990 8362
rect 4016 8358 4020 8362
rect 4053 8358 4057 8362
rect 4090 8358 4094 8362
rect 4118 8358 4122 8362
rect 4148 8358 4152 8362
rect 4185 8358 4189 8362
rect 4222 8358 4226 8362
rect 4250 8358 4254 8362
rect 4280 8358 4284 8362
rect 4317 8358 4321 8362
rect 2529 8325 2533 8329
rect 2557 8325 2561 8329
rect 2587 8325 2591 8329
rect 2624 8325 2628 8329
rect 3474 8325 3478 8329
rect 3502 8325 3506 8329
rect 3532 8325 3536 8329
rect 3569 8325 3573 8329
rect 2871 8281 2875 8285
rect 2900 8281 2904 8285
rect 2925 8281 2929 8285
rect 2967 8281 2971 8285
rect 3023 8281 3027 8285
rect 3047 8281 3051 8285
rect 3101 8281 3105 8285
rect 3128 8281 3132 8285
rect 3182 8281 3186 8285
rect 3816 8281 3820 8285
rect 3845 8281 3849 8285
rect 3870 8281 3874 8285
rect 3912 8281 3916 8285
rect 3968 8281 3972 8285
rect 3992 8281 3996 8285
rect 4046 8281 4050 8285
rect 4073 8281 4077 8285
rect 4127 8281 4131 8285
rect 2489 8223 2493 8227
rect 2526 8223 2530 8227
rect 2556 8223 2560 8227
rect 2584 8223 2588 8227
rect 3434 8223 3438 8227
rect 3471 8223 3475 8227
rect 3501 8223 3505 8227
rect 3529 8223 3533 8227
rect 2871 8149 2875 8153
rect 2900 8149 2904 8153
rect 2925 8149 2929 8153
rect 2967 8149 2971 8153
rect 3023 8149 3027 8153
rect 3047 8149 3051 8153
rect 3101 8149 3105 8153
rect 3128 8149 3132 8153
rect 3190 8149 3194 8153
rect 3816 8149 3820 8153
rect 3845 8149 3849 8153
rect 3870 8149 3874 8153
rect 3912 8149 3916 8153
rect 3968 8149 3972 8153
rect 3992 8149 3996 8153
rect 4046 8149 4050 8153
rect 4073 8149 4077 8153
rect 4135 8149 4139 8153
rect 2871 8017 2875 8021
rect 2900 8017 2904 8021
rect 2925 8017 2929 8021
rect 2967 8017 2971 8021
rect 3023 8017 3027 8021
rect 3047 8017 3051 8021
rect 3101 8017 3105 8021
rect 3128 8017 3132 8021
rect 3182 8017 3186 8021
rect 3190 8017 3194 8021
rect 3218 8017 3222 8021
rect 3272 8017 3276 8021
rect 3816 8017 3820 8021
rect 3845 8017 3849 8021
rect 3870 8017 3874 8021
rect 3912 8017 3916 8021
rect 3968 8017 3972 8021
rect 3992 8017 3996 8021
rect 4046 8017 4050 8021
rect 4073 8017 4077 8021
rect 4127 8017 4131 8021
rect 4135 8017 4139 8021
rect 4163 8017 4167 8021
rect 4217 8017 4221 8021
rect 2871 7885 2875 7889
rect 2900 7885 2904 7889
rect 2925 7885 2929 7889
rect 2967 7885 2971 7889
rect 3023 7885 3027 7889
rect 3047 7885 3051 7889
rect 3101 7885 3105 7889
rect 3128 7885 3132 7889
rect 3218 7885 3222 7889
rect 3816 7885 3820 7889
rect 3845 7885 3849 7889
rect 3870 7885 3874 7889
rect 3912 7885 3916 7889
rect 3968 7885 3972 7889
rect 3992 7885 3996 7889
rect 4046 7885 4050 7889
rect 4073 7885 4077 7889
rect 4163 7885 4167 7889
rect 2397 7823 2401 7827
rect 2425 7823 2429 7827
rect 2455 7823 2459 7827
rect 2492 7823 2496 7827
rect 2529 7823 2533 7827
rect 2557 7823 2561 7827
rect 2587 7823 2591 7827
rect 2624 7823 2628 7827
rect 2661 7823 2665 7827
rect 2689 7823 2693 7827
rect 2719 7823 2723 7827
rect 2756 7823 2760 7827
rect 3342 7823 3346 7827
rect 3370 7823 3374 7827
rect 3400 7823 3404 7827
rect 3437 7823 3441 7827
rect 3474 7823 3478 7827
rect 3502 7823 3506 7827
rect 3532 7823 3536 7827
rect 3569 7823 3573 7827
rect 3606 7823 3610 7827
rect 3634 7823 3638 7827
rect 3664 7823 3668 7827
rect 3701 7823 3705 7827
rect 2871 7753 2875 7757
rect 2900 7753 2904 7757
rect 2925 7753 2929 7757
rect 2967 7753 2971 7757
rect 3047 7753 3051 7757
rect 3101 7753 3105 7757
rect 3132 7753 3136 7757
rect 3161 7753 3165 7757
rect 3186 7753 3190 7757
rect 3228 7753 3232 7757
rect 3816 7753 3820 7757
rect 3845 7753 3849 7757
rect 3870 7753 3874 7757
rect 3912 7753 3916 7757
rect 3992 7753 3996 7757
rect 4046 7753 4050 7757
rect 4077 7753 4081 7757
rect 4106 7753 4110 7757
rect 4131 7753 4135 7757
rect 4173 7753 4177 7757
rect 3180 7711 3184 7715
rect 3208 7711 3212 7715
rect 3238 7711 3242 7715
rect 3275 7711 3279 7715
rect 4125 7711 4129 7715
rect 4153 7711 4157 7715
rect 4183 7711 4187 7715
rect 4220 7711 4224 7715
rect 2397 7681 2401 7685
rect 2425 7681 2429 7685
rect 2455 7681 2459 7685
rect 2492 7681 2496 7685
rect 2529 7681 2533 7685
rect 2557 7681 2561 7685
rect 2587 7681 2591 7685
rect 2624 7681 2628 7685
rect 2661 7681 2665 7685
rect 2689 7681 2693 7685
rect 2719 7681 2723 7685
rect 2756 7681 2760 7685
rect 3342 7681 3346 7685
rect 3370 7681 3374 7685
rect 3400 7681 3404 7685
rect 3437 7681 3441 7685
rect 3474 7681 3478 7685
rect 3502 7681 3506 7685
rect 3532 7681 3536 7685
rect 3569 7681 3573 7685
rect 3606 7681 3610 7685
rect 3634 7681 3638 7685
rect 3664 7681 3668 7685
rect 3701 7681 3705 7685
rect 3180 7625 3184 7629
rect 3208 7625 3212 7629
rect 3238 7625 3242 7629
rect 3275 7625 3279 7629
rect 4125 7625 4129 7629
rect 4153 7625 4157 7629
rect 4183 7625 4187 7629
rect 4220 7625 4224 7629
rect 2397 7595 2401 7599
rect 2425 7595 2429 7599
rect 2455 7595 2459 7599
rect 2492 7595 2496 7599
rect 2529 7595 2533 7599
rect 2557 7595 2561 7599
rect 2587 7595 2591 7599
rect 2624 7595 2628 7599
rect 2661 7595 2665 7599
rect 2689 7595 2693 7599
rect 2719 7595 2723 7599
rect 2756 7595 2760 7599
rect 3342 7595 3346 7599
rect 3370 7595 3374 7599
rect 3400 7595 3404 7599
rect 3437 7595 3441 7599
rect 3474 7595 3478 7599
rect 3502 7595 3506 7599
rect 3532 7595 3536 7599
rect 3569 7595 3573 7599
rect 3606 7595 3610 7599
rect 3634 7595 3638 7599
rect 3664 7595 3668 7599
rect 3701 7595 3705 7599
rect 2397 7455 2401 7459
rect 2425 7455 2429 7459
rect 2455 7455 2459 7459
rect 2492 7455 2496 7459
rect 2529 7455 2533 7459
rect 2557 7455 2561 7459
rect 2587 7455 2591 7459
rect 2624 7455 2628 7459
rect 2661 7455 2665 7459
rect 2689 7455 2693 7459
rect 2719 7455 2723 7459
rect 2756 7455 2760 7459
rect 3342 7455 3346 7459
rect 3370 7455 3374 7459
rect 3400 7455 3404 7459
rect 3437 7455 3441 7459
rect 3474 7455 3478 7459
rect 3502 7455 3506 7459
rect 3532 7455 3536 7459
rect 3569 7455 3573 7459
rect 3606 7455 3610 7459
rect 3634 7455 3638 7459
rect 3664 7455 3668 7459
rect 3701 7455 3705 7459
rect 4525 9573 4529 9577
rect 4535 9573 4539 9577
rect 4545 9573 4549 9577
rect 4555 9573 4559 9577
rect 4525 9568 4529 9572
rect 4535 9568 4539 9572
rect 4545 9568 4549 9572
rect 4555 9568 4559 9572
rect 4525 9563 4529 9567
rect 4535 9563 4539 9567
rect 4545 9563 4549 9567
rect 4555 9563 4559 9567
rect 4525 9558 4529 9562
rect 4535 9558 4539 9562
rect 4545 9558 4549 9562
rect 4555 9558 4559 9562
rect 4525 9544 4529 9548
rect 4535 9544 4539 9548
rect 4545 9544 4549 9548
rect 4555 9544 4559 9548
rect 4525 9539 4529 9543
rect 4535 9539 4539 9543
rect 4545 9539 4549 9543
rect 4555 9539 4559 9543
rect 4525 9534 4529 9538
rect 4535 9534 4539 9538
rect 4545 9534 4549 9538
rect 4555 9534 4559 9538
rect 4525 9529 4529 9533
rect 4535 9529 4539 9533
rect 4545 9529 4549 9533
rect 4555 9529 4559 9533
rect 4525 9515 4529 9519
rect 4535 9515 4539 9519
rect 4545 9515 4549 9519
rect 4555 9515 4559 9519
rect 4525 9510 4529 9514
rect 4535 9510 4539 9514
rect 4545 9510 4549 9514
rect 4555 9510 4559 9514
rect 4525 9505 4529 9509
rect 4535 9505 4539 9509
rect 4545 9505 4549 9509
rect 4555 9505 4559 9509
rect 4525 9500 4529 9504
rect 4535 9500 4539 9504
rect 4545 9500 4549 9504
rect 4555 9500 4559 9504
rect 4525 9486 4529 9490
rect 4535 9486 4539 9490
rect 4545 9486 4549 9490
rect 4555 9486 4559 9490
rect 4525 9481 4529 9485
rect 4535 9481 4539 9485
rect 4545 9481 4549 9485
rect 4555 9481 4559 9485
rect 4525 9476 4529 9480
rect 4535 9476 4539 9480
rect 4545 9476 4549 9480
rect 4555 9476 4559 9480
rect 4525 9471 4529 9475
rect 4535 9471 4539 9475
rect 4545 9471 4549 9475
rect 4555 9471 4559 9475
rect 4525 9457 4529 9461
rect 4535 9457 4539 9461
rect 4545 9457 4549 9461
rect 4555 9457 4559 9461
rect 4525 9452 4529 9456
rect 4535 9452 4539 9456
rect 4545 9452 4549 9456
rect 4555 9452 4559 9456
rect 4525 9447 4529 9451
rect 4535 9447 4539 9451
rect 4545 9447 4549 9451
rect 4555 9447 4559 9451
rect 4525 9442 4529 9446
rect 4535 9442 4539 9446
rect 4545 9442 4549 9446
rect 4555 9442 4559 9446
rect 4525 9056 4529 9060
rect 4535 9056 4539 9060
rect 4545 9056 4549 9060
rect 4555 9056 4559 9060
rect 4525 9051 4529 9055
rect 4535 9051 4539 9055
rect 4545 9051 4549 9055
rect 4555 9051 4559 9055
rect 4525 9046 4529 9050
rect 4535 9046 4539 9050
rect 4545 9046 4549 9050
rect 4555 9046 4559 9050
rect 4525 9041 4529 9045
rect 4535 9041 4539 9045
rect 4545 9041 4549 9045
rect 4555 9041 4559 9045
rect 4525 8747 4529 8751
rect 4535 8747 4539 8751
rect 4545 8747 4549 8751
rect 4555 8747 4559 8751
rect 4525 8742 4529 8746
rect 4535 8742 4539 8746
rect 4545 8742 4549 8746
rect 4555 8742 4559 8746
rect 4525 8737 4529 8741
rect 4535 8737 4539 8741
rect 4545 8737 4549 8741
rect 4555 8737 4559 8741
rect 4525 8732 4529 8736
rect 4535 8732 4539 8736
rect 4545 8732 4549 8736
rect 4555 8732 4559 8736
rect 4525 8438 4529 8442
rect 4535 8438 4539 8442
rect 4545 8438 4549 8442
rect 4555 8438 4559 8442
rect 4525 8433 4529 8437
rect 4535 8433 4539 8437
rect 4545 8433 4549 8437
rect 4555 8433 4559 8437
rect 4525 8428 4529 8432
rect 4535 8428 4539 8432
rect 4545 8428 4549 8432
rect 4555 8428 4559 8432
rect 4525 8423 4529 8427
rect 4535 8423 4539 8427
rect 4545 8423 4549 8427
rect 4555 8423 4559 8427
rect 4525 8129 4529 8133
rect 4535 8129 4539 8133
rect 4545 8129 4549 8133
rect 4555 8129 4559 8133
rect 4525 8124 4529 8128
rect 4535 8124 4539 8128
rect 4545 8124 4549 8128
rect 4555 8124 4559 8128
rect 4525 8119 4529 8123
rect 4535 8119 4539 8123
rect 4545 8119 4549 8123
rect 4555 8119 4559 8123
rect 4525 8114 4529 8118
rect 4535 8114 4539 8118
rect 4545 8114 4549 8118
rect 4555 8114 4559 8118
rect 4525 8098 4529 8102
rect 4535 8098 4539 8102
rect 4545 8098 4549 8102
rect 4555 8098 4559 8102
rect 4525 8093 4529 8097
rect 4535 8093 4539 8097
rect 4545 8093 4549 8097
rect 4555 8093 4559 8097
rect 4525 8088 4529 8092
rect 4535 8088 4539 8092
rect 4545 8088 4549 8092
rect 4555 8088 4559 8092
rect 4525 8083 4529 8087
rect 4535 8083 4539 8087
rect 4545 8083 4549 8087
rect 4555 8083 4559 8087
rect 4627 7889 4631 7945
rect 4666 7857 4670 7945
rect 4709 7857 4713 7945
rect 4750 7857 4754 7945
rect 4525 7789 4529 7793
rect 4535 7789 4539 7793
rect 4545 7789 4549 7793
rect 4555 7789 4559 7793
rect 4525 7784 4529 7788
rect 4535 7784 4539 7788
rect 4545 7784 4549 7788
rect 4555 7784 4559 7788
rect 4525 7779 4529 7783
rect 4535 7779 4539 7783
rect 4545 7779 4549 7783
rect 4555 7779 4559 7783
rect 4525 7774 4529 7778
rect 4535 7774 4539 7778
rect 4545 7774 4549 7778
rect 4555 7774 4559 7778
rect 4525 7202 4529 7206
rect 4535 7202 4539 7206
rect 4545 7202 4549 7206
rect 4555 7202 4559 7206
rect 4525 7197 4529 7201
rect 4535 7197 4539 7201
rect 4545 7197 4549 7201
rect 4555 7197 4559 7201
rect 4525 7192 4529 7196
rect 4535 7192 4539 7196
rect 4545 7192 4549 7196
rect 4555 7192 4559 7196
rect 4525 7187 4529 7191
rect 4535 7187 4539 7191
rect 4545 7187 4549 7191
rect 4555 7187 4559 7191
rect 4525 6893 4529 6897
rect 4535 6893 4539 6897
rect 4545 6893 4549 6897
rect 4555 6893 4559 6897
rect 4525 6888 4529 6892
rect 4535 6888 4539 6892
rect 4545 6888 4549 6892
rect 4555 6888 4559 6892
rect 4525 6883 4529 6887
rect 4535 6883 4539 6887
rect 4545 6883 4549 6887
rect 4555 6883 4559 6887
rect 4525 6878 4529 6882
rect 4535 6878 4539 6882
rect 4545 6878 4549 6882
rect 4555 6878 4559 6882
rect 4525 6584 4529 6588
rect 4535 6584 4539 6588
rect 4545 6584 4549 6588
rect 4555 6584 4559 6588
rect 4525 6579 4529 6583
rect 4535 6579 4539 6583
rect 4545 6579 4549 6583
rect 4555 6579 4559 6583
rect 4525 6574 4529 6578
rect 4535 6574 4539 6578
rect 4545 6574 4549 6578
rect 4555 6574 4559 6578
rect 4525 6569 4529 6573
rect 4535 6569 4539 6573
rect 4545 6569 4549 6573
rect 4555 6569 4559 6573
rect 4525 6275 4529 6279
rect 4535 6275 4539 6279
rect 4545 6275 4549 6279
rect 4555 6275 4559 6279
rect 4525 6270 4529 6274
rect 4535 6270 4539 6274
rect 4545 6270 4549 6274
rect 4555 6270 4559 6274
rect 4525 6265 4529 6269
rect 4535 6265 4539 6269
rect 4545 6265 4549 6269
rect 4555 6265 4559 6269
rect 4525 6260 4529 6264
rect 4535 6260 4539 6264
rect 4545 6260 4549 6264
rect 4555 6260 4559 6264
rect 4525 6083 4529 6087
rect 4535 6083 4539 6087
rect 4545 6083 4549 6087
rect 4555 6083 4559 6087
rect 4525 6078 4529 6082
rect 4535 6078 4539 6082
rect 4545 6078 4549 6082
rect 4555 6078 4559 6082
rect 4525 6073 4529 6077
rect 4535 6073 4539 6077
rect 4545 6073 4549 6077
rect 4555 6073 4559 6077
rect 4525 6068 4529 6072
rect 4535 6068 4539 6072
rect 4545 6068 4549 6072
rect 4555 6068 4559 6072
rect 4525 6057 4529 6061
rect 4535 6057 4539 6061
rect 4545 6057 4549 6061
rect 4555 6057 4559 6061
rect 4525 6052 4529 6056
rect 4535 6052 4539 6056
rect 4545 6052 4549 6056
rect 4555 6052 4559 6056
rect 4525 6047 4529 6051
rect 4535 6047 4539 6051
rect 4545 6047 4549 6051
rect 4555 6047 4559 6051
rect 4525 6042 4529 6046
rect 4535 6042 4539 6046
rect 4545 6042 4549 6046
rect 4555 6042 4559 6046
rect 4525 6031 4529 6035
rect 4535 6031 4539 6035
rect 4545 6031 4549 6035
rect 4555 6031 4559 6035
rect 4525 6026 4529 6030
rect 4535 6026 4539 6030
rect 4545 6026 4549 6030
rect 4555 6026 4559 6030
rect 4525 6021 4529 6025
rect 4535 6021 4539 6025
rect 4545 6021 4549 6025
rect 4555 6021 4559 6025
rect 4525 6016 4529 6020
rect 4535 6016 4539 6020
rect 4545 6016 4549 6020
rect 4555 6016 4559 6020
rect 4525 6005 4529 6009
rect 4535 6005 4539 6009
rect 4545 6005 4549 6009
rect 4555 6005 4559 6009
rect 4525 6000 4529 6004
rect 4535 6000 4539 6004
rect 4545 6000 4549 6004
rect 4555 6000 4559 6004
rect 4525 5995 4529 5999
rect 4535 5995 4539 5999
rect 4545 5995 4549 5999
rect 4555 5995 4559 5999
rect 4525 5990 4529 5994
rect 4535 5990 4539 5994
rect 4545 5990 4549 5994
rect 4555 5990 4559 5994
rect 4525 5979 4529 5983
rect 4535 5979 4539 5983
rect 4545 5979 4549 5983
rect 4555 5979 4559 5983
rect 4525 5974 4529 5978
rect 4535 5974 4539 5978
rect 4545 5974 4549 5978
rect 4555 5974 4559 5978
rect 4525 5969 4529 5973
rect 4535 5969 4539 5973
rect 4545 5969 4549 5973
rect 4555 5969 4559 5973
rect 4525 5964 4529 5968
rect 4535 5964 4539 5968
rect 4545 5964 4549 5968
rect 4555 5964 4559 5968
rect 757 5850 761 5854
rect 762 5850 766 5854
rect 767 5850 771 5854
rect 772 5850 776 5854
rect 783 5850 787 5854
rect 788 5850 792 5854
rect 793 5850 797 5854
rect 798 5850 802 5854
rect 809 5850 813 5854
rect 814 5850 818 5854
rect 819 5850 823 5854
rect 824 5850 828 5854
rect 835 5850 839 5854
rect 840 5850 844 5854
rect 845 5850 849 5854
rect 850 5850 854 5854
rect 861 5850 865 5854
rect 866 5850 870 5854
rect 871 5850 875 5854
rect 876 5850 880 5854
rect 1054 5850 1058 5854
rect 1059 5850 1063 5854
rect 1064 5850 1068 5854
rect 1069 5850 1073 5854
rect 1363 5850 1367 5854
rect 1368 5850 1372 5854
rect 1373 5850 1377 5854
rect 1378 5850 1382 5854
rect 1672 5850 1676 5854
rect 1677 5850 1681 5854
rect 1682 5850 1686 5854
rect 1687 5850 1691 5854
rect 1981 5850 1985 5854
rect 1986 5850 1990 5854
rect 1991 5850 1995 5854
rect 1996 5850 2000 5854
rect 2290 5850 2294 5854
rect 2295 5850 2299 5854
rect 2300 5850 2304 5854
rect 2305 5850 2309 5854
rect 2599 5850 2603 5854
rect 2604 5850 2608 5854
rect 2609 5850 2613 5854
rect 2614 5850 2618 5854
rect 2908 5850 2912 5854
rect 2913 5850 2917 5854
rect 2918 5850 2922 5854
rect 2923 5850 2927 5854
rect 3217 5850 3221 5854
rect 3222 5850 3226 5854
rect 3227 5850 3231 5854
rect 3232 5850 3236 5854
rect 3526 5850 3530 5854
rect 3531 5850 3535 5854
rect 3536 5850 3540 5854
rect 3541 5850 3545 5854
rect 3835 5850 3839 5854
rect 3840 5850 3844 5854
rect 3845 5850 3849 5854
rect 3850 5850 3854 5854
rect 4235 5850 4239 5854
rect 4240 5850 4244 5854
rect 4245 5850 4249 5854
rect 4250 5850 4254 5854
rect 4264 5850 4268 5854
rect 4269 5850 4273 5854
rect 4274 5850 4278 5854
rect 4279 5850 4283 5854
rect 4293 5850 4297 5854
rect 4298 5850 4302 5854
rect 4303 5850 4307 5854
rect 4308 5850 4312 5854
rect 4322 5850 4326 5854
rect 4327 5850 4331 5854
rect 4332 5850 4336 5854
rect 4337 5850 4341 5854
rect 4351 5850 4355 5854
rect 4356 5850 4360 5854
rect 4361 5850 4365 5854
rect 4366 5850 4370 5854
rect 757 5840 761 5844
rect 762 5840 766 5844
rect 767 5840 771 5844
rect 772 5840 776 5844
rect 783 5840 787 5844
rect 788 5840 792 5844
rect 793 5840 797 5844
rect 798 5840 802 5844
rect 809 5840 813 5844
rect 814 5840 818 5844
rect 819 5840 823 5844
rect 824 5840 828 5844
rect 835 5840 839 5844
rect 840 5840 844 5844
rect 845 5840 849 5844
rect 850 5840 854 5844
rect 861 5840 865 5844
rect 866 5840 870 5844
rect 871 5840 875 5844
rect 876 5840 880 5844
rect 1054 5840 1058 5844
rect 1059 5840 1063 5844
rect 1064 5840 1068 5844
rect 1069 5840 1073 5844
rect 1363 5840 1367 5844
rect 1368 5840 1372 5844
rect 1373 5840 1377 5844
rect 1378 5840 1382 5844
rect 1672 5840 1676 5844
rect 1677 5840 1681 5844
rect 1682 5840 1686 5844
rect 1687 5840 1691 5844
rect 1981 5840 1985 5844
rect 1986 5840 1990 5844
rect 1991 5840 1995 5844
rect 1996 5840 2000 5844
rect 2290 5840 2294 5844
rect 2295 5840 2299 5844
rect 2300 5840 2304 5844
rect 2305 5840 2309 5844
rect 2599 5840 2603 5844
rect 2604 5840 2608 5844
rect 2609 5840 2613 5844
rect 2614 5840 2618 5844
rect 2908 5840 2912 5844
rect 2913 5840 2917 5844
rect 2918 5840 2922 5844
rect 2923 5840 2927 5844
rect 3217 5840 3221 5844
rect 3222 5840 3226 5844
rect 3227 5840 3231 5844
rect 3232 5840 3236 5844
rect 3526 5840 3530 5844
rect 3531 5840 3535 5844
rect 3536 5840 3540 5844
rect 3541 5840 3545 5844
rect 3835 5840 3839 5844
rect 3840 5840 3844 5844
rect 3845 5840 3849 5844
rect 3850 5840 3854 5844
rect 4235 5840 4239 5844
rect 4240 5840 4244 5844
rect 4245 5840 4249 5844
rect 4250 5840 4254 5844
rect 4264 5840 4268 5844
rect 4269 5840 4273 5844
rect 4274 5840 4278 5844
rect 4279 5840 4283 5844
rect 4293 5840 4297 5844
rect 4298 5840 4302 5844
rect 4303 5840 4307 5844
rect 4308 5840 4312 5844
rect 4322 5840 4326 5844
rect 4327 5840 4331 5844
rect 4332 5840 4336 5844
rect 4337 5840 4341 5844
rect 4351 5840 4355 5844
rect 4356 5840 4360 5844
rect 4361 5840 4365 5844
rect 4366 5840 4370 5844
rect 757 5830 761 5834
rect 762 5830 766 5834
rect 767 5830 771 5834
rect 772 5830 776 5834
rect 783 5830 787 5834
rect 788 5830 792 5834
rect 793 5830 797 5834
rect 798 5830 802 5834
rect 809 5830 813 5834
rect 814 5830 818 5834
rect 819 5830 823 5834
rect 824 5830 828 5834
rect 835 5830 839 5834
rect 840 5830 844 5834
rect 845 5830 849 5834
rect 850 5830 854 5834
rect 861 5830 865 5834
rect 866 5830 870 5834
rect 871 5830 875 5834
rect 876 5830 880 5834
rect 1054 5830 1058 5834
rect 1059 5830 1063 5834
rect 1064 5830 1068 5834
rect 1069 5830 1073 5834
rect 1363 5830 1367 5834
rect 1368 5830 1372 5834
rect 1373 5830 1377 5834
rect 1378 5830 1382 5834
rect 1672 5830 1676 5834
rect 1677 5830 1681 5834
rect 1682 5830 1686 5834
rect 1687 5830 1691 5834
rect 1981 5830 1985 5834
rect 1986 5830 1990 5834
rect 1991 5830 1995 5834
rect 1996 5830 2000 5834
rect 2290 5830 2294 5834
rect 2295 5830 2299 5834
rect 2300 5830 2304 5834
rect 2305 5830 2309 5834
rect 2599 5830 2603 5834
rect 2604 5830 2608 5834
rect 2609 5830 2613 5834
rect 2614 5830 2618 5834
rect 2908 5830 2912 5834
rect 2913 5830 2917 5834
rect 2918 5830 2922 5834
rect 2923 5830 2927 5834
rect 3217 5830 3221 5834
rect 3222 5830 3226 5834
rect 3227 5830 3231 5834
rect 3232 5830 3236 5834
rect 3526 5830 3530 5834
rect 3531 5830 3535 5834
rect 3536 5830 3540 5834
rect 3541 5830 3545 5834
rect 3835 5830 3839 5834
rect 3840 5830 3844 5834
rect 3845 5830 3849 5834
rect 3850 5830 3854 5834
rect 4235 5830 4239 5834
rect 4240 5830 4244 5834
rect 4245 5830 4249 5834
rect 4250 5830 4254 5834
rect 4264 5830 4268 5834
rect 4269 5830 4273 5834
rect 4274 5830 4278 5834
rect 4279 5830 4283 5834
rect 4293 5830 4297 5834
rect 4298 5830 4302 5834
rect 4303 5830 4307 5834
rect 4308 5830 4312 5834
rect 4322 5830 4326 5834
rect 4327 5830 4331 5834
rect 4332 5830 4336 5834
rect 4337 5830 4341 5834
rect 4351 5830 4355 5834
rect 4356 5830 4360 5834
rect 4361 5830 4365 5834
rect 4366 5830 4370 5834
rect 757 5820 761 5824
rect 762 5820 766 5824
rect 767 5820 771 5824
rect 772 5820 776 5824
rect 783 5820 787 5824
rect 788 5820 792 5824
rect 793 5820 797 5824
rect 798 5820 802 5824
rect 809 5820 813 5824
rect 814 5820 818 5824
rect 819 5820 823 5824
rect 824 5820 828 5824
rect 835 5820 839 5824
rect 840 5820 844 5824
rect 845 5820 849 5824
rect 850 5820 854 5824
rect 861 5820 865 5824
rect 866 5820 870 5824
rect 871 5820 875 5824
rect 876 5820 880 5824
rect 1054 5820 1058 5824
rect 1059 5820 1063 5824
rect 1064 5820 1068 5824
rect 1069 5820 1073 5824
rect 1363 5820 1367 5824
rect 1368 5820 1372 5824
rect 1373 5820 1377 5824
rect 1378 5820 1382 5824
rect 1672 5820 1676 5824
rect 1677 5820 1681 5824
rect 1682 5820 1686 5824
rect 1687 5820 1691 5824
rect 1981 5820 1985 5824
rect 1986 5820 1990 5824
rect 1991 5820 1995 5824
rect 1996 5820 2000 5824
rect 2290 5820 2294 5824
rect 2295 5820 2299 5824
rect 2300 5820 2304 5824
rect 2305 5820 2309 5824
rect 2599 5820 2603 5824
rect 2604 5820 2608 5824
rect 2609 5820 2613 5824
rect 2614 5820 2618 5824
rect 2908 5820 2912 5824
rect 2913 5820 2917 5824
rect 2918 5820 2922 5824
rect 2923 5820 2927 5824
rect 3217 5820 3221 5824
rect 3222 5820 3226 5824
rect 3227 5820 3231 5824
rect 3232 5820 3236 5824
rect 3526 5820 3530 5824
rect 3531 5820 3535 5824
rect 3536 5820 3540 5824
rect 3541 5820 3545 5824
rect 3835 5820 3839 5824
rect 3840 5820 3844 5824
rect 3845 5820 3849 5824
rect 3850 5820 3854 5824
rect 4235 5820 4239 5824
rect 4240 5820 4244 5824
rect 4245 5820 4249 5824
rect 4250 5820 4254 5824
rect 4264 5820 4268 5824
rect 4269 5820 4273 5824
rect 4274 5820 4278 5824
rect 4279 5820 4283 5824
rect 4293 5820 4297 5824
rect 4298 5820 4302 5824
rect 4303 5820 4307 5824
rect 4308 5820 4312 5824
rect 4322 5820 4326 5824
rect 4327 5820 4331 5824
rect 4332 5820 4336 5824
rect 4337 5820 4341 5824
rect 4351 5820 4355 5824
rect 4356 5820 4360 5824
rect 4361 5820 4365 5824
rect 4366 5820 4370 5824
<< polysilicon >>
rect 118 9786 1024 10280
rect 1797 9883 1818 9952
rect 2106 9883 2127 9952
rect 2415 9883 2436 9952
rect 2724 9883 2745 9952
rect 3033 9883 3054 9952
rect 3960 9883 3981 9952
rect 1803 9826 1812 9827
rect 2112 9826 2121 9827
rect 2421 9826 2430 9827
rect 2730 9826 2739 9827
rect 3039 9826 3048 9827
rect 3966 9826 3975 9827
rect 1741 9824 1743 9826
rect 1799 9824 1829 9826
rect 1869 9824 1871 9826
rect 2050 9824 2052 9826
rect 2108 9824 2138 9826
rect 2178 9824 2180 9826
rect 2359 9824 2361 9826
rect 2417 9824 2447 9826
rect 2487 9824 2489 9826
rect 2668 9824 2670 9826
rect 2726 9824 2756 9826
rect 2796 9824 2798 9826
rect 2977 9824 2979 9826
rect 3035 9824 3065 9826
rect 3105 9824 3107 9826
rect 3904 9824 3906 9826
rect 3962 9824 3992 9826
rect 4032 9824 4034 9826
rect 1806 9818 1808 9824
rect 2115 9818 2117 9824
rect 2424 9818 2426 9824
rect 2733 9818 2735 9824
rect 3042 9818 3044 9824
rect 3969 9818 3971 9824
rect 1741 9816 1743 9818
rect 1799 9816 1829 9818
rect 1869 9816 1871 9818
rect 2050 9816 2052 9818
rect 2108 9816 2138 9818
rect 2178 9816 2180 9818
rect 2359 9816 2361 9818
rect 2417 9816 2447 9818
rect 2487 9816 2489 9818
rect 2668 9816 2670 9818
rect 2726 9816 2756 9818
rect 2796 9816 2798 9818
rect 2977 9816 2979 9818
rect 3035 9816 3065 9818
rect 3105 9816 3107 9818
rect 3904 9816 3906 9818
rect 3962 9816 3992 9818
rect 4032 9816 4034 9818
rect 1740 9808 1743 9810
rect 1799 9808 1813 9810
rect 1819 9808 1829 9810
rect 1869 9808 1872 9810
rect 1740 9802 1742 9808
rect 1800 9806 1828 9808
rect 1800 9802 1802 9806
rect 1740 9800 1743 9802
rect 1799 9800 1802 9802
rect 1740 9794 1742 9800
rect 1800 9794 1802 9800
rect 1740 9792 1743 9794
rect 1799 9792 1802 9794
rect 1740 9786 1742 9792
rect 1800 9786 1802 9792
rect 118 9348 593 9786
rect 1740 9784 1743 9786
rect 1799 9784 1802 9786
rect 1826 9802 1828 9806
rect 1870 9802 1872 9808
rect 1826 9800 1829 9802
rect 1869 9800 1872 9802
rect 1826 9794 1828 9800
rect 1870 9794 1872 9800
rect 1826 9792 1829 9794
rect 1869 9792 1872 9794
rect 1826 9786 1828 9792
rect 1870 9786 1872 9792
rect 1826 9784 1829 9786
rect 1869 9784 1872 9786
rect 2049 9808 2052 9810
rect 2108 9808 2122 9810
rect 2128 9808 2138 9810
rect 2178 9808 2181 9810
rect 2049 9802 2051 9808
rect 2109 9806 2137 9808
rect 2109 9802 2111 9806
rect 2049 9800 2052 9802
rect 2108 9800 2111 9802
rect 2049 9794 2051 9800
rect 2109 9794 2111 9800
rect 2049 9792 2052 9794
rect 2108 9792 2111 9794
rect 2049 9786 2051 9792
rect 2109 9786 2111 9792
rect 2049 9784 2052 9786
rect 2108 9784 2111 9786
rect 2135 9802 2137 9806
rect 2179 9802 2181 9808
rect 2135 9800 2138 9802
rect 2178 9800 2181 9802
rect 2135 9794 2137 9800
rect 2179 9794 2181 9800
rect 2135 9792 2138 9794
rect 2178 9792 2181 9794
rect 2135 9786 2137 9792
rect 2179 9786 2181 9792
rect 2135 9784 2138 9786
rect 2178 9784 2181 9786
rect 2358 9808 2361 9810
rect 2417 9808 2431 9810
rect 2437 9808 2447 9810
rect 2487 9808 2490 9810
rect 2358 9802 2360 9808
rect 2418 9806 2446 9808
rect 2418 9802 2420 9806
rect 2358 9800 2361 9802
rect 2417 9800 2420 9802
rect 2358 9794 2360 9800
rect 2418 9794 2420 9800
rect 2358 9792 2361 9794
rect 2417 9792 2420 9794
rect 2358 9786 2360 9792
rect 2418 9786 2420 9792
rect 2358 9784 2361 9786
rect 2417 9784 2420 9786
rect 2444 9802 2446 9806
rect 2488 9802 2490 9808
rect 2444 9800 2447 9802
rect 2487 9800 2490 9802
rect 2444 9794 2446 9800
rect 2488 9794 2490 9800
rect 2444 9792 2447 9794
rect 2487 9792 2490 9794
rect 2444 9786 2446 9792
rect 2488 9786 2490 9792
rect 2444 9784 2447 9786
rect 2487 9784 2490 9786
rect 2667 9808 2670 9810
rect 2726 9808 2740 9810
rect 2746 9808 2756 9810
rect 2796 9808 2799 9810
rect 2667 9802 2669 9808
rect 2727 9806 2755 9808
rect 2727 9802 2729 9806
rect 2667 9800 2670 9802
rect 2726 9800 2729 9802
rect 2667 9794 2669 9800
rect 2727 9794 2729 9800
rect 2667 9792 2670 9794
rect 2726 9792 2729 9794
rect 2667 9786 2669 9792
rect 2727 9786 2729 9792
rect 2667 9784 2670 9786
rect 2726 9784 2729 9786
rect 2753 9802 2755 9806
rect 2797 9802 2799 9808
rect 2753 9800 2756 9802
rect 2796 9800 2799 9802
rect 2753 9794 2755 9800
rect 2797 9794 2799 9800
rect 2753 9792 2756 9794
rect 2796 9792 2799 9794
rect 2753 9786 2755 9792
rect 2797 9786 2799 9792
rect 2753 9784 2756 9786
rect 2796 9784 2799 9786
rect 2976 9808 2979 9810
rect 3035 9808 3049 9810
rect 3055 9808 3065 9810
rect 3105 9808 3108 9810
rect 2976 9802 2978 9808
rect 3036 9806 3064 9808
rect 3036 9802 3038 9806
rect 2976 9800 2979 9802
rect 3035 9800 3038 9802
rect 2976 9794 2978 9800
rect 3036 9794 3038 9800
rect 2976 9792 2979 9794
rect 3035 9792 3038 9794
rect 2976 9786 2978 9792
rect 3036 9786 3038 9792
rect 2976 9784 2979 9786
rect 3035 9784 3038 9786
rect 3062 9802 3064 9806
rect 3106 9802 3108 9808
rect 3062 9800 3065 9802
rect 3105 9800 3108 9802
rect 3062 9794 3064 9800
rect 3106 9794 3108 9800
rect 3062 9792 3065 9794
rect 3105 9792 3108 9794
rect 3062 9786 3064 9792
rect 3106 9786 3108 9792
rect 3062 9784 3065 9786
rect 3105 9784 3108 9786
rect 3903 9808 3906 9810
rect 3962 9808 3976 9810
rect 3982 9808 3992 9810
rect 4032 9808 4035 9810
rect 3903 9802 3905 9808
rect 3963 9806 3991 9808
rect 3963 9802 3965 9806
rect 3903 9800 3906 9802
rect 3962 9800 3965 9802
rect 3903 9794 3905 9800
rect 3963 9794 3965 9800
rect 3903 9792 3906 9794
rect 3962 9792 3965 9794
rect 3903 9786 3905 9792
rect 3963 9786 3965 9792
rect 3903 9784 3906 9786
rect 3962 9784 3965 9786
rect 3989 9802 3991 9806
rect 4033 9802 4035 9808
rect 3989 9800 3992 9802
rect 4032 9800 4035 9802
rect 3989 9794 3991 9800
rect 4033 9794 4035 9800
rect 3989 9792 3992 9794
rect 4032 9792 4035 9794
rect 3989 9786 3991 9792
rect 4033 9786 4035 9792
rect 4141 9786 5073 10261
rect 3989 9784 3992 9786
rect 4032 9784 4035 9786
rect 99 5800 593 6231
rect 2856 9330 2858 9332
rect 2861 9330 2863 9333
rect 2877 9330 2879 9332
rect 2893 9330 2895 9332
rect 2898 9330 2900 9333
rect 2919 9330 2921 9333
rect 2935 9330 2937 9333
rect 2951 9330 2953 9332
rect 2956 9330 2958 9333
rect 2972 9330 2974 9332
rect 2988 9330 2990 9332
rect 2993 9330 2995 9333
rect 3009 9330 3011 9332
rect 3025 9330 3027 9332
rect 3030 9330 3032 9333
rect 3051 9330 3053 9333
rect 3067 9330 3069 9333
rect 3083 9330 3085 9332
rect 3088 9330 3090 9333
rect 3104 9330 3106 9332
rect 3120 9330 3122 9332
rect 3125 9330 3127 9333
rect 3141 9330 3143 9332
rect 3157 9330 3159 9332
rect 3162 9330 3164 9333
rect 3183 9330 3185 9333
rect 3199 9330 3201 9333
rect 3215 9330 3217 9332
rect 3220 9330 3222 9333
rect 3236 9330 3238 9332
rect 3252 9330 3254 9332
rect 3257 9330 3259 9333
rect 3273 9330 3275 9332
rect 3289 9330 3291 9332
rect 3294 9330 3296 9333
rect 3315 9330 3317 9333
rect 3331 9330 3333 9333
rect 3347 9330 3349 9332
rect 3352 9330 3354 9333
rect 3368 9330 3370 9332
rect 3801 9330 3803 9332
rect 3806 9330 3808 9333
rect 3822 9330 3824 9332
rect 3838 9330 3840 9332
rect 3843 9330 3845 9333
rect 3864 9330 3866 9333
rect 3880 9330 3882 9333
rect 3896 9330 3898 9332
rect 3901 9330 3903 9333
rect 3917 9330 3919 9332
rect 3933 9330 3935 9332
rect 3938 9330 3940 9333
rect 3954 9330 3956 9332
rect 3970 9330 3972 9332
rect 3975 9330 3977 9333
rect 3996 9330 3998 9333
rect 4012 9330 4014 9333
rect 4028 9330 4030 9332
rect 4033 9330 4035 9333
rect 4049 9330 4051 9332
rect 4065 9330 4067 9332
rect 4070 9330 4072 9333
rect 4086 9330 4088 9332
rect 4102 9330 4104 9332
rect 4107 9330 4109 9333
rect 4128 9330 4130 9333
rect 4144 9330 4146 9333
rect 4160 9330 4162 9332
rect 4165 9330 4167 9333
rect 4181 9330 4183 9332
rect 4197 9330 4199 9332
rect 4202 9330 4204 9333
rect 4218 9330 4220 9332
rect 4234 9330 4236 9332
rect 4239 9330 4241 9333
rect 4260 9330 4262 9333
rect 4276 9330 4278 9333
rect 4292 9330 4294 9332
rect 4297 9330 4299 9333
rect 4313 9330 4315 9332
rect 2856 9317 2858 9322
rect 2861 9320 2863 9322
rect 2856 9303 2858 9313
rect 2861 9303 2863 9310
rect 2877 9303 2879 9322
rect 2893 9313 2895 9322
rect 2898 9320 2900 9322
rect 2919 9320 2921 9322
rect 2935 9319 2937 9322
rect 2893 9303 2895 9306
rect 2898 9303 2900 9305
rect 2919 9303 2921 9305
rect 2935 9303 2937 9315
rect 2951 9313 2953 9322
rect 2956 9320 2958 9322
rect 2972 9314 2974 9322
rect 2988 9317 2990 9322
rect 2993 9320 2995 9322
rect 2951 9303 2953 9306
rect 2956 9303 2958 9305
rect 2972 9303 2974 9310
rect 2988 9303 2990 9313
rect 2993 9303 2995 9310
rect 3009 9303 3011 9322
rect 3025 9313 3027 9322
rect 3030 9320 3032 9322
rect 3051 9320 3053 9322
rect 3067 9319 3069 9322
rect 3025 9303 3027 9306
rect 3030 9303 3032 9305
rect 3051 9303 3053 9305
rect 3067 9303 3069 9315
rect 3083 9313 3085 9322
rect 3088 9320 3090 9322
rect 3104 9314 3106 9322
rect 3120 9317 3122 9322
rect 3125 9320 3127 9322
rect 3083 9303 3085 9306
rect 3088 9303 3090 9305
rect 3104 9303 3106 9310
rect 3120 9303 3122 9313
rect 3125 9303 3127 9310
rect 3141 9303 3143 9322
rect 3157 9313 3159 9322
rect 3162 9320 3164 9322
rect 3183 9320 3185 9322
rect 3199 9319 3201 9322
rect 3157 9303 3159 9306
rect 3162 9303 3164 9305
rect 3183 9303 3185 9305
rect 3199 9303 3201 9315
rect 3215 9313 3217 9322
rect 3220 9320 3222 9322
rect 3236 9314 3238 9322
rect 3252 9317 3254 9322
rect 3257 9320 3259 9322
rect 3215 9303 3217 9306
rect 3220 9303 3222 9305
rect 3236 9303 3238 9310
rect 3252 9303 3254 9313
rect 3257 9303 3259 9310
rect 3273 9303 3275 9322
rect 3289 9313 3291 9322
rect 3294 9320 3296 9322
rect 3315 9320 3317 9322
rect 3331 9319 3333 9322
rect 3289 9303 3291 9306
rect 3294 9303 3296 9305
rect 3315 9303 3317 9305
rect 3331 9303 3333 9315
rect 3347 9313 3349 9322
rect 3352 9320 3354 9322
rect 3368 9314 3370 9322
rect 3801 9317 3803 9322
rect 3806 9320 3808 9322
rect 3347 9303 3349 9306
rect 3352 9303 3354 9305
rect 3368 9303 3370 9310
rect 2504 9297 2506 9299
rect 2509 9297 2511 9300
rect 2525 9297 2527 9299
rect 2541 9297 2543 9299
rect 2546 9297 2548 9300
rect 2567 9297 2569 9300
rect 2583 9297 2585 9300
rect 2599 9297 2601 9299
rect 2604 9297 2606 9300
rect 3801 9303 3803 9313
rect 3806 9303 3808 9310
rect 3822 9303 3824 9322
rect 3838 9313 3840 9322
rect 3843 9320 3845 9322
rect 3864 9320 3866 9322
rect 3880 9319 3882 9322
rect 3838 9303 3840 9306
rect 3843 9303 3845 9305
rect 3864 9303 3866 9305
rect 3880 9303 3882 9315
rect 3896 9313 3898 9322
rect 3901 9320 3903 9322
rect 3917 9314 3919 9322
rect 3933 9317 3935 9322
rect 3938 9320 3940 9322
rect 3896 9303 3898 9306
rect 3901 9303 3903 9305
rect 3917 9303 3919 9310
rect 3933 9303 3935 9313
rect 3938 9303 3940 9310
rect 3954 9303 3956 9322
rect 3970 9313 3972 9322
rect 3975 9320 3977 9322
rect 3996 9320 3998 9322
rect 4012 9319 4014 9322
rect 3970 9303 3972 9306
rect 3975 9303 3977 9305
rect 3996 9303 3998 9305
rect 4012 9303 4014 9315
rect 4028 9313 4030 9322
rect 4033 9320 4035 9322
rect 4049 9314 4051 9322
rect 4065 9317 4067 9322
rect 4070 9320 4072 9322
rect 4028 9303 4030 9306
rect 4033 9303 4035 9305
rect 4049 9303 4051 9310
rect 4065 9303 4067 9313
rect 4070 9303 4072 9310
rect 4086 9303 4088 9322
rect 4102 9313 4104 9322
rect 4107 9320 4109 9322
rect 4128 9320 4130 9322
rect 4144 9319 4146 9322
rect 4102 9303 4104 9306
rect 4107 9303 4109 9305
rect 4128 9303 4130 9305
rect 4144 9303 4146 9315
rect 4160 9313 4162 9322
rect 4165 9320 4167 9322
rect 4181 9314 4183 9322
rect 4197 9317 4199 9322
rect 4202 9320 4204 9322
rect 4160 9303 4162 9306
rect 4165 9303 4167 9305
rect 4181 9303 4183 9310
rect 4197 9303 4199 9313
rect 4202 9303 4204 9310
rect 4218 9303 4220 9322
rect 4234 9313 4236 9322
rect 4239 9320 4241 9322
rect 4260 9320 4262 9322
rect 4276 9319 4278 9322
rect 4234 9303 4236 9306
rect 4239 9303 4241 9305
rect 4260 9303 4262 9305
rect 4276 9303 4278 9315
rect 4292 9313 4294 9322
rect 4297 9320 4299 9322
rect 4313 9314 4315 9322
rect 4292 9303 4294 9306
rect 4297 9303 4299 9305
rect 4313 9303 4315 9310
rect 2620 9297 2622 9299
rect 2856 9297 2858 9299
rect 2861 9296 2863 9299
rect 2877 9297 2879 9299
rect 2893 9297 2895 9299
rect 2898 9294 2900 9299
rect 2919 9294 2921 9299
rect 2935 9297 2937 9299
rect 2951 9297 2953 9299
rect 2956 9294 2958 9299
rect 2972 9297 2974 9299
rect 2988 9297 2990 9299
rect 2993 9296 2995 9299
rect 3009 9297 3011 9299
rect 3025 9297 3027 9299
rect 3030 9294 3032 9299
rect 3051 9294 3053 9299
rect 3067 9297 3069 9299
rect 3083 9297 3085 9299
rect 3088 9294 3090 9299
rect 3104 9297 3106 9299
rect 3120 9297 3122 9299
rect 3125 9296 3127 9299
rect 3141 9297 3143 9299
rect 3157 9297 3159 9299
rect 3162 9294 3164 9299
rect 3183 9294 3185 9299
rect 3199 9297 3201 9299
rect 3215 9297 3217 9299
rect 3220 9294 3222 9299
rect 3236 9297 3238 9299
rect 3252 9297 3254 9299
rect 3257 9296 3259 9299
rect 3273 9297 3275 9299
rect 3289 9297 3291 9299
rect 3294 9294 3296 9299
rect 3315 9294 3317 9299
rect 3331 9297 3333 9299
rect 3347 9297 3349 9299
rect 3352 9294 3354 9299
rect 3368 9297 3370 9299
rect 3449 9297 3451 9299
rect 3454 9297 3456 9300
rect 3470 9297 3472 9299
rect 3486 9297 3488 9299
rect 3491 9297 3493 9300
rect 3512 9297 3514 9300
rect 3528 9297 3530 9300
rect 3544 9297 3546 9299
rect 3549 9297 3551 9300
rect 3565 9297 3567 9299
rect 3801 9297 3803 9299
rect 3806 9296 3808 9299
rect 3822 9297 3824 9299
rect 3838 9297 3840 9299
rect 3843 9294 3845 9299
rect 3864 9294 3866 9299
rect 3880 9297 3882 9299
rect 3896 9297 3898 9299
rect 3901 9294 3903 9299
rect 3917 9297 3919 9299
rect 3933 9297 3935 9299
rect 3938 9296 3940 9299
rect 3954 9297 3956 9299
rect 3970 9297 3972 9299
rect 3975 9294 3977 9299
rect 3996 9294 3998 9299
rect 4012 9297 4014 9299
rect 4028 9297 4030 9299
rect 4033 9294 4035 9299
rect 4049 9297 4051 9299
rect 4065 9297 4067 9299
rect 4070 9296 4072 9299
rect 4086 9297 4088 9299
rect 4102 9297 4104 9299
rect 4107 9294 4109 9299
rect 4128 9294 4130 9299
rect 4144 9297 4146 9299
rect 4160 9297 4162 9299
rect 4165 9294 4167 9299
rect 4181 9297 4183 9299
rect 4197 9297 4199 9299
rect 4202 9296 4204 9299
rect 4218 9297 4220 9299
rect 4234 9297 4236 9299
rect 4239 9294 4241 9299
rect 4260 9294 4262 9299
rect 4276 9297 4278 9299
rect 4292 9297 4294 9299
rect 4297 9294 4299 9299
rect 4313 9297 4315 9299
rect 2504 9284 2506 9289
rect 2509 9287 2511 9289
rect 2504 9270 2506 9280
rect 2509 9270 2511 9277
rect 2525 9270 2527 9289
rect 2541 9280 2543 9289
rect 2546 9287 2548 9289
rect 2567 9287 2569 9289
rect 2583 9286 2585 9289
rect 2541 9270 2543 9273
rect 2546 9270 2548 9272
rect 2567 9270 2569 9272
rect 2583 9270 2585 9282
rect 2599 9280 2601 9289
rect 2604 9287 2606 9289
rect 2599 9270 2601 9273
rect 2604 9270 2606 9272
rect 2620 9270 2622 9289
rect 3449 9284 3451 9289
rect 3454 9287 3456 9289
rect 3449 9270 3451 9280
rect 3454 9270 3456 9277
rect 3470 9270 3472 9289
rect 3486 9280 3488 9289
rect 3491 9287 3493 9289
rect 3512 9287 3514 9289
rect 3528 9286 3530 9289
rect 3486 9270 3488 9273
rect 3491 9270 3493 9272
rect 3512 9270 3514 9272
rect 3528 9270 3530 9282
rect 3544 9280 3546 9289
rect 3549 9287 3551 9289
rect 3544 9270 3546 9273
rect 3549 9270 3551 9272
rect 3565 9270 3567 9289
rect 2504 9264 2506 9266
rect 2509 9263 2511 9266
rect 2525 9264 2527 9266
rect 2541 9264 2543 9266
rect 2546 9261 2548 9266
rect 2567 9261 2569 9266
rect 2583 9264 2585 9266
rect 2599 9264 2601 9266
rect 2604 9261 2606 9266
rect 2620 9264 2622 9266
rect 3449 9264 3451 9266
rect 3454 9263 3456 9266
rect 3470 9264 3472 9266
rect 3486 9264 3488 9266
rect 3035 9259 3037 9261
rect 2877 9253 2879 9256
rect 2921 9253 2923 9256
rect 2947 9253 2949 9256
rect 2993 9253 2995 9256
rect 2947 9249 2948 9253
rect 3061 9253 3063 9257
rect 3089 9259 3091 9261
rect 3116 9259 3118 9261
rect 3066 9253 3068 9256
rect 2861 9246 2863 9248
rect 2877 9246 2879 9249
rect 2893 9246 2895 9248
rect 2916 9246 2918 9248
rect 2921 9246 2923 9249
rect 2947 9246 2949 9249
rect 2968 9246 2970 9249
rect 2988 9246 2990 9248
rect 2993 9246 2995 9249
rect 3011 9246 3013 9248
rect 2628 9233 2630 9236
rect 2628 9227 2630 9229
rect 2511 9224 2513 9227
rect 2861 9224 2863 9238
rect 2877 9236 2879 9238
rect 2877 9224 2879 9226
rect 2893 9224 2895 9238
rect 2916 9233 2918 9238
rect 2921 9236 2923 9238
rect 2947 9236 2949 9238
rect 2912 9229 2918 9233
rect 2916 9224 2918 9229
rect 2921 9224 2923 9226
rect 2947 9224 2949 9226
rect 2968 9224 2970 9238
rect 2988 9233 2990 9238
rect 2993 9236 2995 9238
rect 2984 9229 2990 9233
rect 2988 9224 2990 9229
rect 2993 9224 2995 9226
rect 3011 9224 3013 9238
rect 3035 9237 3037 9251
rect 3142 9253 3144 9257
rect 3170 9259 3172 9261
rect 3491 9261 3493 9266
rect 3512 9261 3514 9266
rect 3528 9264 3530 9266
rect 3544 9264 3546 9266
rect 3549 9261 3551 9266
rect 3565 9264 3567 9266
rect 3147 9253 3149 9256
rect 3061 9242 3063 9245
rect 3066 9243 3068 9245
rect 3062 9238 3063 9242
rect 3061 9233 3063 9238
rect 3066 9233 3068 9235
rect 3035 9231 3037 9233
rect 3089 9229 3091 9251
rect 3116 9237 3118 9251
rect 3980 9259 3982 9261
rect 3142 9242 3144 9245
rect 3147 9243 3149 9245
rect 3143 9238 3144 9242
rect 3142 9233 3144 9238
rect 3147 9233 3149 9235
rect 3116 9231 3118 9233
rect 3170 9229 3172 9251
rect 3822 9253 3824 9256
rect 3866 9253 3868 9256
rect 3892 9253 3894 9256
rect 3938 9253 3940 9256
rect 3892 9249 3893 9253
rect 4006 9253 4008 9257
rect 4034 9259 4036 9261
rect 4061 9259 4063 9261
rect 4011 9253 4013 9256
rect 3806 9246 3808 9248
rect 3822 9246 3824 9249
rect 3838 9246 3840 9248
rect 3861 9246 3863 9248
rect 3866 9246 3868 9249
rect 3892 9246 3894 9249
rect 3913 9246 3915 9249
rect 3933 9246 3935 9248
rect 3938 9246 3940 9249
rect 3956 9246 3958 9248
rect 3573 9233 3575 9236
rect 3061 9227 3063 9229
rect 3066 9224 3068 9229
rect 3142 9227 3144 9229
rect 3089 9223 3091 9225
rect 3147 9224 3149 9229
rect 3573 9227 3575 9229
rect 3170 9223 3172 9225
rect 3456 9224 3458 9227
rect 3806 9224 3808 9238
rect 3822 9236 3824 9238
rect 3822 9224 3824 9226
rect 3838 9224 3840 9238
rect 3861 9233 3863 9238
rect 3866 9236 3868 9238
rect 3892 9236 3894 9238
rect 3857 9229 3863 9233
rect 3861 9224 3863 9229
rect 3866 9224 3868 9226
rect 3892 9224 3894 9226
rect 3913 9224 3915 9238
rect 3933 9233 3935 9238
rect 3938 9236 3940 9238
rect 3929 9229 3935 9233
rect 3933 9224 3935 9229
rect 3938 9224 3940 9226
rect 3956 9224 3958 9238
rect 3980 9237 3982 9251
rect 4087 9253 4089 9257
rect 4115 9259 4117 9261
rect 4092 9253 4094 9256
rect 4006 9242 4008 9245
rect 4011 9243 4013 9245
rect 4007 9238 4008 9242
rect 4006 9233 4008 9238
rect 4011 9233 4013 9235
rect 3980 9231 3982 9233
rect 4034 9229 4036 9251
rect 4061 9237 4063 9251
rect 4087 9242 4089 9245
rect 4092 9243 4094 9245
rect 4088 9238 4089 9242
rect 4087 9233 4089 9238
rect 4092 9233 4094 9235
rect 4061 9231 4063 9233
rect 4115 9229 4117 9251
rect 4006 9227 4008 9229
rect 4011 9224 4013 9229
rect 4087 9227 4089 9229
rect 4034 9223 4036 9225
rect 4092 9224 4094 9229
rect 4115 9223 4117 9225
rect 2511 9218 2513 9220
rect 2861 9218 2863 9220
rect 2877 9216 2879 9220
rect 2893 9218 2895 9220
rect 2916 9218 2918 9220
rect 2878 9212 2879 9216
rect 2921 9215 2923 9220
rect 2947 9216 2949 9220
rect 2968 9218 2970 9220
rect 2988 9218 2990 9220
rect 2877 9209 2879 9212
rect 2922 9211 2923 9215
rect 2948 9212 2949 9216
rect 2993 9215 2995 9220
rect 3011 9218 3013 9220
rect 3456 9218 3458 9220
rect 3806 9218 3808 9220
rect 3822 9216 3824 9220
rect 3838 9218 3840 9220
rect 3861 9218 3863 9220
rect 2921 9209 2923 9211
rect 2947 9208 2949 9212
rect 2994 9211 2995 9215
rect 3823 9212 3824 9216
rect 3866 9215 3868 9220
rect 3892 9216 3894 9220
rect 3913 9218 3915 9220
rect 3933 9218 3935 9220
rect 2993 9209 2995 9211
rect 3822 9209 3824 9212
rect 3867 9211 3868 9215
rect 3893 9212 3894 9216
rect 3938 9215 3940 9220
rect 3956 9218 3958 9220
rect 3866 9209 3868 9211
rect 3892 9208 3894 9212
rect 3939 9211 3940 9215
rect 3938 9209 3940 9211
rect 2495 9195 2497 9197
rect 2511 9195 2513 9198
rect 2516 9195 2518 9197
rect 2532 9195 2534 9198
rect 2548 9195 2550 9198
rect 2569 9195 2571 9198
rect 2574 9195 2576 9197
rect 2590 9195 2592 9197
rect 2606 9195 2608 9198
rect 2611 9195 2613 9197
rect 3440 9195 3442 9197
rect 3456 9195 3458 9198
rect 3461 9195 3463 9197
rect 3477 9195 3479 9198
rect 3493 9195 3495 9198
rect 3514 9195 3516 9198
rect 3519 9195 3521 9197
rect 3535 9195 3537 9197
rect 3551 9195 3553 9198
rect 3556 9195 3558 9197
rect 2495 9168 2497 9187
rect 2511 9185 2513 9187
rect 2516 9178 2518 9187
rect 2532 9184 2534 9187
rect 2548 9185 2550 9187
rect 2569 9185 2571 9187
rect 2511 9168 2513 9170
rect 2516 9168 2518 9171
rect 2532 9168 2534 9180
rect 2574 9178 2576 9187
rect 2548 9168 2550 9170
rect 2569 9168 2571 9170
rect 2574 9168 2576 9171
rect 2590 9168 2592 9187
rect 2606 9185 2608 9187
rect 2611 9182 2613 9187
rect 2877 9186 2879 9189
rect 2921 9187 2923 9189
rect 2878 9182 2879 9186
rect 2922 9183 2923 9187
rect 2947 9186 2949 9190
rect 2993 9187 2995 9189
rect 2861 9178 2863 9180
rect 2877 9178 2879 9182
rect 2893 9178 2895 9180
rect 2916 9178 2918 9180
rect 2921 9178 2923 9183
rect 2948 9182 2949 9186
rect 2994 9183 2995 9187
rect 2947 9178 2949 9182
rect 2968 9178 2970 9180
rect 2988 9178 2990 9180
rect 2993 9178 2995 9183
rect 3011 9178 3013 9180
rect 2606 9168 2608 9175
rect 2611 9168 2613 9178
rect 3061 9177 3063 9180
rect 3066 9177 3068 9180
rect 3142 9177 3144 9180
rect 3147 9177 3149 9180
rect 2495 9162 2497 9164
rect 2511 9159 2513 9164
rect 2516 9162 2518 9164
rect 2532 9162 2534 9164
rect 2548 9159 2550 9164
rect 2569 9159 2571 9164
rect 2574 9162 2576 9164
rect 2590 9162 2592 9164
rect 2606 9161 2608 9164
rect 2611 9162 2613 9164
rect 2861 9160 2863 9174
rect 2877 9172 2879 9174
rect 2877 9160 2879 9162
rect 2893 9160 2895 9174
rect 2916 9169 2918 9174
rect 2921 9172 2923 9174
rect 2947 9172 2949 9174
rect 2912 9165 2918 9169
rect 2916 9160 2918 9165
rect 2921 9160 2923 9162
rect 2947 9160 2949 9162
rect 2968 9160 2970 9174
rect 2988 9169 2990 9174
rect 2993 9172 2995 9174
rect 2984 9165 2990 9169
rect 2988 9160 2990 9165
rect 2993 9160 2995 9162
rect 3011 9160 3013 9174
rect 3061 9161 3063 9173
rect 3066 9171 3068 9173
rect 3066 9161 3068 9163
rect 3142 9161 3144 9173
rect 3147 9171 3149 9173
rect 3440 9168 3442 9187
rect 3456 9185 3458 9187
rect 3461 9178 3463 9187
rect 3477 9184 3479 9187
rect 3493 9185 3495 9187
rect 3514 9185 3516 9187
rect 3456 9168 3458 9170
rect 3461 9168 3463 9171
rect 3477 9168 3479 9180
rect 3519 9178 3521 9187
rect 3493 9168 3495 9170
rect 3514 9168 3516 9170
rect 3519 9168 3521 9171
rect 3535 9168 3537 9187
rect 3551 9185 3553 9187
rect 3556 9182 3558 9187
rect 3822 9186 3824 9189
rect 3866 9187 3868 9189
rect 3823 9182 3824 9186
rect 3867 9183 3868 9187
rect 3892 9186 3894 9190
rect 3938 9187 3940 9189
rect 3806 9178 3808 9180
rect 3822 9178 3824 9182
rect 3838 9178 3840 9180
rect 3861 9178 3863 9180
rect 3866 9178 3868 9183
rect 3893 9182 3894 9186
rect 3939 9183 3940 9187
rect 3892 9178 3894 9182
rect 3913 9178 3915 9180
rect 3933 9178 3935 9180
rect 3938 9178 3940 9183
rect 3956 9178 3958 9180
rect 3551 9168 3553 9175
rect 3556 9168 3558 9178
rect 4006 9177 4008 9180
rect 4011 9177 4013 9180
rect 4087 9177 4089 9180
rect 4092 9177 4094 9180
rect 3147 9161 3149 9163
rect 3440 9162 3442 9164
rect 3456 9159 3458 9164
rect 3461 9162 3463 9164
rect 3477 9162 3479 9164
rect 3493 9159 3495 9164
rect 3514 9159 3516 9164
rect 3519 9162 3521 9164
rect 3535 9162 3537 9164
rect 3551 9161 3553 9164
rect 3556 9162 3558 9164
rect 3806 9160 3808 9174
rect 3822 9172 3824 9174
rect 3822 9160 3824 9162
rect 3838 9160 3840 9174
rect 3861 9169 3863 9174
rect 3866 9172 3868 9174
rect 3892 9172 3894 9174
rect 3857 9165 3863 9169
rect 3861 9160 3863 9165
rect 3866 9160 3868 9162
rect 3892 9160 3894 9162
rect 3913 9160 3915 9174
rect 3933 9169 3935 9174
rect 3938 9172 3940 9174
rect 3929 9165 3935 9169
rect 3933 9160 3935 9165
rect 3938 9160 3940 9162
rect 3956 9160 3958 9174
rect 4006 9161 4008 9173
rect 4011 9171 4013 9173
rect 4011 9161 4013 9163
rect 4087 9161 4089 9173
rect 4092 9171 4094 9173
rect 4092 9161 4094 9163
rect 2861 9150 2863 9152
rect 2877 9149 2879 9152
rect 2893 9150 2895 9152
rect 2916 9150 2918 9152
rect 2921 9149 2923 9152
rect 2947 9149 2949 9152
rect 2968 9149 2970 9152
rect 2988 9150 2990 9152
rect 2993 9149 2995 9152
rect 3011 9150 3013 9152
rect 3061 9151 3063 9153
rect 2947 9145 2948 9149
rect 3066 9148 3068 9153
rect 3142 9151 3144 9153
rect 3147 9148 3149 9153
rect 3806 9150 3808 9152
rect 3822 9149 3824 9152
rect 3838 9150 3840 9152
rect 3861 9150 3863 9152
rect 3866 9149 3868 9152
rect 3892 9149 3894 9152
rect 3913 9149 3915 9152
rect 3933 9150 3935 9152
rect 3938 9149 3940 9152
rect 3956 9150 3958 9152
rect 4006 9151 4008 9153
rect 2877 9142 2879 9145
rect 2921 9142 2923 9145
rect 2947 9142 2949 9145
rect 2993 9142 2995 9145
rect 3892 9145 3893 9149
rect 4011 9148 4013 9153
rect 4087 9151 4089 9153
rect 4092 9148 4094 9153
rect 3822 9142 3824 9145
rect 3866 9142 3868 9145
rect 3892 9142 3894 9145
rect 3938 9142 3940 9145
rect 2877 9121 2879 9124
rect 2921 9121 2923 9124
rect 2947 9121 2949 9124
rect 2993 9121 2995 9124
rect 3061 9121 3063 9125
rect 3089 9127 3091 9129
rect 3140 9127 3142 9129
rect 3066 9121 3068 9124
rect 2947 9117 2948 9121
rect 2861 9114 2863 9116
rect 2877 9114 2879 9117
rect 2893 9114 2895 9116
rect 2916 9114 2918 9116
rect 2921 9114 2923 9117
rect 2947 9114 2949 9117
rect 2968 9114 2970 9117
rect 2988 9114 2990 9116
rect 2993 9114 2995 9117
rect 3011 9114 3013 9116
rect 3166 9121 3168 9125
rect 3194 9127 3196 9129
rect 3171 9121 3173 9124
rect 3061 9110 3063 9113
rect 3066 9111 3068 9113
rect 3062 9106 3063 9110
rect 2861 9092 2863 9106
rect 2877 9104 2879 9106
rect 2877 9092 2879 9094
rect 2893 9092 2895 9106
rect 2916 9101 2918 9106
rect 2921 9104 2923 9106
rect 2947 9104 2949 9106
rect 2912 9097 2918 9101
rect 2916 9092 2918 9097
rect 2921 9092 2923 9094
rect 2947 9092 2949 9094
rect 2968 9092 2970 9106
rect 2988 9101 2990 9106
rect 2993 9104 2995 9106
rect 2984 9097 2990 9101
rect 2988 9092 2990 9097
rect 2993 9092 2995 9094
rect 3011 9092 3013 9106
rect 3061 9101 3063 9106
rect 3066 9101 3068 9103
rect 3089 9097 3091 9119
rect 3140 9105 3142 9119
rect 3822 9121 3824 9124
rect 3866 9121 3868 9124
rect 3892 9121 3894 9124
rect 3938 9121 3940 9124
rect 4006 9121 4008 9125
rect 4034 9127 4036 9129
rect 4085 9127 4087 9129
rect 4011 9121 4013 9124
rect 3166 9110 3168 9113
rect 3171 9111 3173 9113
rect 3167 9106 3168 9110
rect 3166 9101 3168 9106
rect 3171 9101 3173 9103
rect 3140 9099 3142 9101
rect 3194 9097 3196 9119
rect 3892 9117 3893 9121
rect 3806 9114 3808 9116
rect 3822 9114 3824 9117
rect 3838 9114 3840 9116
rect 3861 9114 3863 9116
rect 3866 9114 3868 9117
rect 3892 9114 3894 9117
rect 3913 9114 3915 9117
rect 3933 9114 3935 9116
rect 3938 9114 3940 9117
rect 3956 9114 3958 9116
rect 4111 9121 4113 9125
rect 4139 9127 4141 9129
rect 4116 9121 4118 9124
rect 4006 9110 4008 9113
rect 4011 9111 4013 9113
rect 4007 9106 4008 9110
rect 3371 9098 3373 9100
rect 3061 9095 3063 9097
rect 3066 9092 3068 9097
rect 3166 9095 3168 9097
rect 3089 9091 3091 9093
rect 3171 9092 3173 9097
rect 3194 9091 3196 9093
rect 3397 9092 3399 9096
rect 3425 9098 3427 9100
rect 3402 9092 3404 9095
rect 2861 9086 2863 9088
rect 2877 9084 2879 9088
rect 2893 9086 2895 9088
rect 2916 9086 2918 9088
rect 2878 9080 2879 9084
rect 2921 9083 2923 9088
rect 2947 9084 2949 9088
rect 2968 9086 2970 9088
rect 2988 9086 2990 9088
rect 2877 9077 2879 9080
rect 2922 9079 2923 9083
rect 2948 9080 2949 9084
rect 2993 9083 2995 9088
rect 3011 9086 3013 9088
rect 2921 9077 2923 9079
rect 2947 9076 2949 9080
rect 2994 9079 2995 9083
rect 2993 9077 2995 9079
rect 3371 9076 3373 9090
rect 3557 9095 3559 9098
rect 3610 9095 3612 9098
rect 3397 9081 3399 9084
rect 3402 9082 3404 9084
rect 3398 9077 3399 9081
rect 3397 9072 3399 9077
rect 3402 9072 3404 9074
rect 3371 9070 3373 9072
rect 3425 9068 3427 9090
rect 3397 9066 3399 9068
rect 3402 9063 3404 9068
rect 3806 9092 3808 9106
rect 3822 9104 3824 9106
rect 3822 9092 3824 9094
rect 3838 9092 3840 9106
rect 3861 9101 3863 9106
rect 3866 9104 3868 9106
rect 3892 9104 3894 9106
rect 3857 9097 3863 9101
rect 3861 9092 3863 9097
rect 3866 9092 3868 9094
rect 3892 9092 3894 9094
rect 3913 9092 3915 9106
rect 3933 9101 3935 9106
rect 3938 9104 3940 9106
rect 3929 9097 3935 9101
rect 3933 9092 3935 9097
rect 3938 9092 3940 9094
rect 3956 9092 3958 9106
rect 4006 9101 4008 9106
rect 4011 9101 4013 9103
rect 4034 9097 4036 9119
rect 4085 9105 4087 9119
rect 4111 9110 4113 9113
rect 4116 9111 4118 9113
rect 4112 9106 4113 9110
rect 4111 9101 4113 9106
rect 4116 9101 4118 9103
rect 4085 9099 4087 9101
rect 4139 9097 4141 9119
rect 4006 9095 4008 9097
rect 4011 9092 4013 9097
rect 4111 9095 4113 9097
rect 4034 9091 4036 9093
rect 4116 9092 4118 9097
rect 4139 9091 4141 9093
rect 3806 9086 3808 9088
rect 3822 9084 3824 9088
rect 3838 9086 3840 9088
rect 3861 9086 3863 9088
rect 3823 9080 3824 9084
rect 3866 9083 3868 9088
rect 3892 9084 3894 9088
rect 3913 9086 3915 9088
rect 3933 9086 3935 9088
rect 3822 9077 3824 9080
rect 3867 9079 3868 9083
rect 3893 9080 3894 9084
rect 3938 9083 3940 9088
rect 3956 9086 3958 9088
rect 3866 9077 3868 9079
rect 3892 9076 3894 9080
rect 3939 9079 3940 9083
rect 3938 9077 3940 9079
rect 3425 9062 3427 9064
rect 2877 9054 2879 9057
rect 2921 9055 2923 9057
rect 2878 9050 2879 9054
rect 2922 9051 2923 9055
rect 2947 9054 2949 9058
rect 3557 9057 3559 9065
rect 3610 9057 3612 9065
rect 2993 9055 2995 9057
rect 2861 9046 2863 9048
rect 2877 9046 2879 9050
rect 2893 9046 2895 9048
rect 2916 9046 2918 9048
rect 2921 9046 2923 9051
rect 2948 9050 2949 9054
rect 2994 9051 2995 9055
rect 3822 9054 3824 9057
rect 3866 9055 3868 9057
rect 2947 9046 2949 9050
rect 2968 9046 2970 9048
rect 2988 9046 2990 9048
rect 2993 9046 2995 9051
rect 3011 9046 3013 9048
rect 3061 9046 3063 9049
rect 3066 9046 3068 9049
rect 3166 9046 3168 9049
rect 3171 9046 3173 9049
rect 3557 9045 3559 9053
rect 3610 9045 3612 9053
rect 3823 9050 3824 9054
rect 3867 9051 3868 9055
rect 3892 9054 3894 9058
rect 3938 9055 3940 9057
rect 3806 9046 3808 9048
rect 3822 9046 3824 9050
rect 3838 9046 3840 9048
rect 3861 9046 3863 9048
rect 3866 9046 3868 9051
rect 3893 9050 3894 9054
rect 3939 9051 3940 9055
rect 3892 9046 3894 9050
rect 3913 9046 3915 9048
rect 3933 9046 3935 9048
rect 3938 9046 3940 9051
rect 3956 9046 3958 9048
rect 4006 9046 4008 9049
rect 4011 9046 4013 9049
rect 4111 9046 4113 9049
rect 4116 9046 4118 9049
rect 2861 9028 2863 9042
rect 2877 9040 2879 9042
rect 2877 9028 2879 9030
rect 2893 9028 2895 9042
rect 2916 9037 2918 9042
rect 2921 9040 2923 9042
rect 2947 9040 2949 9042
rect 2912 9033 2918 9037
rect 2916 9028 2918 9033
rect 2921 9028 2923 9030
rect 2947 9028 2949 9030
rect 2968 9028 2970 9042
rect 2988 9037 2990 9042
rect 2993 9040 2995 9042
rect 2984 9033 2990 9037
rect 2988 9028 2990 9033
rect 2993 9028 2995 9030
rect 3011 9028 3013 9042
rect 3061 9030 3063 9042
rect 3066 9040 3068 9042
rect 3066 9030 3068 9032
rect 3166 9030 3168 9042
rect 3171 9040 3173 9042
rect 3171 9030 3173 9032
rect 3557 9031 3559 9033
rect 3610 9031 3612 9033
rect 3806 9028 3808 9042
rect 3822 9040 3824 9042
rect 3822 9028 3824 9030
rect 3838 9028 3840 9042
rect 3861 9037 3863 9042
rect 3866 9040 3868 9042
rect 3892 9040 3894 9042
rect 3857 9033 3863 9037
rect 3861 9028 3863 9033
rect 3866 9028 3868 9030
rect 3892 9028 3894 9030
rect 3913 9028 3915 9042
rect 3933 9037 3935 9042
rect 3938 9040 3940 9042
rect 3929 9033 3935 9037
rect 3933 9028 3935 9033
rect 3938 9028 3940 9030
rect 3956 9028 3958 9042
rect 4006 9030 4008 9042
rect 4011 9040 4013 9042
rect 4011 9030 4013 9032
rect 4111 9030 4113 9042
rect 4116 9040 4118 9042
rect 4116 9030 4118 9032
rect 3061 9020 3063 9022
rect 2861 9018 2863 9020
rect 2877 9017 2879 9020
rect 2893 9018 2895 9020
rect 2916 9018 2918 9020
rect 2921 9017 2923 9020
rect 2947 9017 2949 9020
rect 2968 9017 2970 9020
rect 2988 9018 2990 9020
rect 2993 9017 2995 9020
rect 3011 9018 3013 9020
rect 3066 9017 3068 9022
rect 3166 9020 3168 9022
rect 3171 9017 3173 9022
rect 4006 9020 4008 9022
rect 2947 9013 2948 9017
rect 3806 9018 3808 9020
rect 3822 9017 3824 9020
rect 3838 9018 3840 9020
rect 3861 9018 3863 9020
rect 3866 9017 3868 9020
rect 3892 9017 3894 9020
rect 3913 9017 3915 9020
rect 3933 9018 3935 9020
rect 3938 9017 3940 9020
rect 3956 9018 3958 9020
rect 4011 9017 4013 9022
rect 4111 9020 4113 9022
rect 4116 9017 4118 9022
rect 2877 9010 2879 9013
rect 2921 9010 2923 9013
rect 2947 9010 2949 9013
rect 2993 9010 2995 9013
rect 3397 9012 3399 9015
rect 3402 9012 3404 9015
rect 3892 9013 3893 9017
rect 3822 9010 3824 9013
rect 3866 9010 3868 9013
rect 3892 9010 3894 9013
rect 3938 9010 3940 9013
rect 2877 8989 2879 8992
rect 2921 8989 2923 8992
rect 2947 8989 2949 8992
rect 2993 8989 2995 8992
rect 3061 8989 3063 8993
rect 3089 8995 3091 8997
rect 3116 8995 3118 8997
rect 3066 8989 3068 8992
rect 2947 8985 2948 8989
rect 2861 8982 2863 8984
rect 2877 8982 2879 8985
rect 2893 8982 2895 8984
rect 2916 8982 2918 8984
rect 2921 8982 2923 8985
rect 2947 8982 2949 8985
rect 2968 8982 2970 8985
rect 2988 8982 2990 8984
rect 2993 8982 2995 8985
rect 3011 8982 3013 8984
rect 3142 8989 3144 8993
rect 3170 8995 3172 8997
rect 3206 8995 3208 8997
rect 3147 8989 3149 8992
rect 3061 8978 3063 8981
rect 3066 8979 3068 8981
rect 3062 8974 3063 8978
rect 2861 8960 2863 8974
rect 2877 8972 2879 8974
rect 2877 8960 2879 8962
rect 2893 8960 2895 8974
rect 2916 8969 2918 8974
rect 2921 8972 2923 8974
rect 2947 8972 2949 8974
rect 2912 8965 2918 8969
rect 2916 8960 2918 8965
rect 2921 8960 2923 8962
rect 2947 8960 2949 8962
rect 2968 8960 2970 8974
rect 2988 8969 2990 8974
rect 2993 8972 2995 8974
rect 2984 8965 2990 8969
rect 2988 8960 2990 8965
rect 2993 8960 2995 8962
rect 3011 8960 3013 8974
rect 3061 8969 3063 8974
rect 3066 8969 3068 8971
rect 3089 8965 3091 8987
rect 3116 8973 3118 8987
rect 3232 8989 3234 8993
rect 3260 8995 3262 8997
rect 3397 8996 3399 9008
rect 3402 9006 3404 9008
rect 3402 8996 3404 8998
rect 3237 8989 3239 8992
rect 3142 8978 3144 8981
rect 3147 8979 3149 8981
rect 3143 8974 3144 8978
rect 3142 8969 3144 8974
rect 3147 8969 3149 8971
rect 3116 8967 3118 8969
rect 3170 8965 3172 8987
rect 3206 8973 3208 8987
rect 3822 8989 3824 8992
rect 3866 8989 3868 8992
rect 3892 8989 3894 8992
rect 3938 8989 3940 8992
rect 4006 8989 4008 8993
rect 4034 8995 4036 8997
rect 4061 8995 4063 8997
rect 4011 8989 4013 8992
rect 3232 8978 3234 8981
rect 3237 8979 3239 8981
rect 3233 8974 3234 8978
rect 3232 8969 3234 8974
rect 3237 8969 3239 8971
rect 3206 8967 3208 8969
rect 3260 8965 3262 8987
rect 3397 8986 3399 8988
rect 3402 8983 3404 8988
rect 3892 8985 3893 8989
rect 3806 8982 3808 8984
rect 3822 8982 3824 8985
rect 3838 8982 3840 8984
rect 3861 8982 3863 8984
rect 3866 8982 3868 8985
rect 3892 8982 3894 8985
rect 3913 8982 3915 8985
rect 3933 8982 3935 8984
rect 3938 8982 3940 8985
rect 3956 8982 3958 8984
rect 4087 8989 4089 8993
rect 4115 8995 4117 8997
rect 4151 8995 4153 8997
rect 4092 8989 4094 8992
rect 4006 8978 4008 8981
rect 4011 8979 4013 8981
rect 4007 8974 4008 8978
rect 3349 8968 3351 8970
rect 3371 8968 3373 8970
rect 3061 8963 3063 8965
rect 3066 8960 3068 8965
rect 3142 8963 3144 8965
rect 3089 8959 3091 8961
rect 3147 8960 3149 8965
rect 3232 8963 3234 8965
rect 3170 8959 3172 8961
rect 3237 8960 3239 8965
rect 3260 8959 3262 8961
rect 3397 8962 3399 8966
rect 3425 8968 3427 8970
rect 3402 8962 3404 8965
rect 2861 8954 2863 8956
rect 2877 8952 2879 8956
rect 2893 8954 2895 8956
rect 2916 8954 2918 8956
rect 2878 8948 2879 8952
rect 2921 8951 2923 8956
rect 2947 8952 2949 8956
rect 2968 8954 2970 8956
rect 2988 8954 2990 8956
rect 2877 8945 2879 8948
rect 2922 8947 2923 8951
rect 2948 8948 2949 8952
rect 2993 8951 2995 8956
rect 3011 8954 3013 8956
rect 2921 8945 2923 8947
rect 2947 8944 2949 8948
rect 2994 8947 2995 8951
rect 2993 8945 2995 8947
rect 3349 8946 3351 8960
rect 3371 8946 3373 8960
rect 3463 8965 3465 8968
rect 3516 8965 3518 8968
rect 3397 8951 3399 8954
rect 3402 8952 3404 8954
rect 3398 8947 3399 8951
rect 3397 8942 3399 8947
rect 3402 8942 3404 8944
rect 3349 8940 3351 8942
rect 3371 8940 3373 8942
rect 3425 8938 3427 8960
rect 3397 8936 3399 8938
rect 3402 8933 3404 8938
rect 3806 8960 3808 8974
rect 3822 8972 3824 8974
rect 3822 8960 3824 8962
rect 3838 8960 3840 8974
rect 3861 8969 3863 8974
rect 3866 8972 3868 8974
rect 3892 8972 3894 8974
rect 3857 8965 3863 8969
rect 3861 8960 3863 8965
rect 3866 8960 3868 8962
rect 3892 8960 3894 8962
rect 3913 8960 3915 8974
rect 3933 8969 3935 8974
rect 3938 8972 3940 8974
rect 3929 8965 3935 8969
rect 3933 8960 3935 8965
rect 3938 8960 3940 8962
rect 3956 8960 3958 8974
rect 4006 8969 4008 8974
rect 4011 8969 4013 8971
rect 4034 8965 4036 8987
rect 4061 8973 4063 8987
rect 4177 8989 4179 8993
rect 4205 8995 4207 8997
rect 4182 8989 4184 8992
rect 4087 8978 4089 8981
rect 4092 8979 4094 8981
rect 4088 8974 4089 8978
rect 4087 8969 4089 8974
rect 4092 8969 4094 8971
rect 4061 8967 4063 8969
rect 4115 8965 4117 8987
rect 4151 8973 4153 8987
rect 4177 8978 4179 8981
rect 4182 8979 4184 8981
rect 4178 8974 4179 8978
rect 4177 8969 4179 8974
rect 4182 8969 4184 8971
rect 4151 8967 4153 8969
rect 4205 8965 4207 8987
rect 4006 8963 4008 8965
rect 4011 8960 4013 8965
rect 4087 8963 4089 8965
rect 4034 8959 4036 8961
rect 4092 8960 4094 8965
rect 4177 8963 4179 8965
rect 4115 8959 4117 8961
rect 4182 8960 4184 8965
rect 4205 8959 4207 8961
rect 3806 8954 3808 8956
rect 3822 8952 3824 8956
rect 3838 8954 3840 8956
rect 3861 8954 3863 8956
rect 3823 8948 3824 8952
rect 3866 8951 3868 8956
rect 3892 8952 3894 8956
rect 3913 8954 3915 8956
rect 3933 8954 3935 8956
rect 3822 8945 3824 8948
rect 3867 8947 3868 8951
rect 3893 8948 3894 8952
rect 3938 8951 3940 8956
rect 3956 8954 3958 8956
rect 3866 8945 3868 8947
rect 3892 8944 3894 8948
rect 3939 8947 3940 8951
rect 3938 8945 3940 8947
rect 3425 8932 3427 8934
rect 3463 8927 3465 8935
rect 3516 8927 3518 8935
rect 2877 8922 2879 8925
rect 2921 8923 2923 8925
rect 2878 8918 2879 8922
rect 2922 8919 2923 8923
rect 2947 8922 2949 8926
rect 2993 8923 2995 8925
rect 2861 8914 2863 8916
rect 2877 8914 2879 8918
rect 2893 8914 2895 8916
rect 2916 8914 2918 8916
rect 2921 8914 2923 8919
rect 2948 8918 2949 8922
rect 2994 8919 2995 8923
rect 2947 8914 2949 8918
rect 2968 8914 2970 8916
rect 2988 8914 2990 8916
rect 2993 8914 2995 8919
rect 3011 8914 3013 8916
rect 3463 8915 3465 8923
rect 3516 8915 3518 8923
rect 3822 8922 3824 8925
rect 3866 8923 3868 8925
rect 3823 8918 3824 8922
rect 3867 8919 3868 8923
rect 3892 8922 3894 8926
rect 3938 8923 3940 8925
rect 3061 8911 3063 8914
rect 3066 8911 3068 8914
rect 3142 8911 3144 8914
rect 3147 8911 3149 8914
rect 3232 8911 3234 8914
rect 3237 8911 3239 8914
rect 2861 8896 2863 8910
rect 2877 8908 2879 8910
rect 2877 8896 2879 8898
rect 2893 8896 2895 8910
rect 2916 8905 2918 8910
rect 2921 8908 2923 8910
rect 2947 8908 2949 8910
rect 2912 8901 2918 8905
rect 2916 8896 2918 8901
rect 2921 8896 2923 8898
rect 2947 8896 2949 8898
rect 2968 8896 2970 8910
rect 2988 8905 2990 8910
rect 2993 8908 2995 8910
rect 2984 8901 2990 8905
rect 2988 8896 2990 8901
rect 2993 8896 2995 8898
rect 3011 8896 3013 8910
rect 3061 8895 3063 8907
rect 3066 8905 3068 8907
rect 3066 8895 3068 8897
rect 3142 8895 3144 8907
rect 3147 8905 3149 8907
rect 3147 8895 3149 8897
rect 3232 8895 3234 8907
rect 3237 8905 3239 8907
rect 3806 8914 3808 8916
rect 3822 8914 3824 8918
rect 3838 8914 3840 8916
rect 3861 8914 3863 8916
rect 3866 8914 3868 8919
rect 3893 8918 3894 8922
rect 3939 8919 3940 8923
rect 3892 8914 3894 8918
rect 3913 8914 3915 8916
rect 3933 8914 3935 8916
rect 3938 8914 3940 8919
rect 3956 8914 3958 8916
rect 4006 8911 4008 8914
rect 4011 8911 4013 8914
rect 4087 8911 4089 8914
rect 4092 8911 4094 8914
rect 4177 8911 4179 8914
rect 4182 8911 4184 8914
rect 3463 8901 3465 8903
rect 3516 8901 3518 8903
rect 3237 8895 3239 8897
rect 3806 8896 3808 8910
rect 3822 8908 3824 8910
rect 3822 8896 3824 8898
rect 3838 8896 3840 8910
rect 3861 8905 3863 8910
rect 3866 8908 3868 8910
rect 3892 8908 3894 8910
rect 3857 8901 3863 8905
rect 3861 8896 3863 8901
rect 3866 8896 3868 8898
rect 3892 8896 3894 8898
rect 3913 8896 3915 8910
rect 3933 8905 3935 8910
rect 3938 8908 3940 8910
rect 3929 8901 3935 8905
rect 3933 8896 3935 8901
rect 3938 8896 3940 8898
rect 3956 8896 3958 8910
rect 2861 8886 2863 8888
rect 2877 8885 2879 8888
rect 2893 8886 2895 8888
rect 2916 8886 2918 8888
rect 2921 8885 2923 8888
rect 2947 8885 2949 8888
rect 2968 8885 2970 8888
rect 2988 8886 2990 8888
rect 2993 8885 2995 8888
rect 3011 8886 3013 8888
rect 3061 8885 3063 8887
rect 2947 8881 2948 8885
rect 3066 8882 3068 8887
rect 3142 8885 3144 8887
rect 3147 8882 3149 8887
rect 3232 8885 3234 8887
rect 3237 8882 3239 8887
rect 4006 8895 4008 8907
rect 4011 8905 4013 8907
rect 4011 8895 4013 8897
rect 4087 8895 4089 8907
rect 4092 8905 4094 8907
rect 4092 8895 4094 8897
rect 4177 8895 4179 8907
rect 4182 8905 4184 8907
rect 4182 8895 4184 8897
rect 3806 8886 3808 8888
rect 3822 8885 3824 8888
rect 3838 8886 3840 8888
rect 3861 8886 3863 8888
rect 3866 8885 3868 8888
rect 3892 8885 3894 8888
rect 3913 8885 3915 8888
rect 3933 8886 3935 8888
rect 3938 8885 3940 8888
rect 3956 8886 3958 8888
rect 4006 8885 4008 8887
rect 3397 8882 3399 8885
rect 3402 8882 3404 8885
rect 2877 8878 2879 8881
rect 2921 8878 2923 8881
rect 2947 8878 2949 8881
rect 2993 8878 2995 8881
rect 3892 8881 3893 8885
rect 4011 8882 4013 8887
rect 4087 8885 4089 8887
rect 4092 8882 4094 8887
rect 4177 8885 4179 8887
rect 4182 8882 4184 8887
rect 3822 8878 3824 8881
rect 3866 8878 3868 8881
rect 3892 8878 3894 8881
rect 3938 8878 3940 8881
rect 3397 8866 3399 8878
rect 3402 8876 3404 8878
rect 3402 8866 3404 8868
rect 2877 8857 2879 8860
rect 2921 8857 2923 8860
rect 2947 8857 2949 8860
rect 2993 8857 2995 8860
rect 3061 8857 3063 8861
rect 3089 8863 3091 8865
rect 3066 8857 3068 8860
rect 2947 8853 2948 8857
rect 2861 8850 2863 8852
rect 2877 8850 2879 8853
rect 2893 8850 2895 8852
rect 2916 8850 2918 8852
rect 2921 8850 2923 8853
rect 2947 8850 2949 8853
rect 2968 8850 2970 8853
rect 2988 8850 2990 8852
rect 2993 8850 2995 8853
rect 3011 8850 3013 8852
rect 3397 8856 3399 8858
rect 3061 8846 3063 8849
rect 3066 8847 3068 8849
rect 3062 8842 3063 8846
rect 2861 8828 2863 8842
rect 2877 8840 2879 8842
rect 2877 8828 2879 8830
rect 2893 8828 2895 8842
rect 2916 8837 2918 8842
rect 2921 8840 2923 8842
rect 2947 8840 2949 8842
rect 2912 8833 2918 8837
rect 2916 8828 2918 8833
rect 2921 8828 2923 8830
rect 2947 8828 2949 8830
rect 2968 8828 2970 8842
rect 2988 8837 2990 8842
rect 2993 8840 2995 8842
rect 2984 8833 2990 8837
rect 2988 8828 2990 8833
rect 2993 8828 2995 8830
rect 3011 8828 3013 8842
rect 3061 8837 3063 8842
rect 3066 8837 3068 8839
rect 3089 8833 3091 8855
rect 3402 8853 3404 8858
rect 3822 8857 3824 8860
rect 3866 8857 3868 8860
rect 3892 8857 3894 8860
rect 3938 8857 3940 8860
rect 4006 8857 4008 8861
rect 4034 8863 4036 8865
rect 4011 8857 4013 8860
rect 3892 8853 3893 8857
rect 3806 8850 3808 8852
rect 3822 8850 3824 8853
rect 3838 8850 3840 8852
rect 3861 8850 3863 8852
rect 3866 8850 3868 8853
rect 3892 8850 3894 8853
rect 3913 8850 3915 8853
rect 3933 8850 3935 8852
rect 3938 8850 3940 8853
rect 3956 8850 3958 8852
rect 4006 8846 4008 8849
rect 4011 8847 4013 8849
rect 4007 8842 4008 8846
rect 3061 8831 3063 8833
rect 3066 8828 3068 8833
rect 3089 8827 3091 8829
rect 3806 8828 3808 8842
rect 3822 8840 3824 8842
rect 3822 8828 3824 8830
rect 3838 8828 3840 8842
rect 3861 8837 3863 8842
rect 3866 8840 3868 8842
rect 3892 8840 3894 8842
rect 3857 8833 3863 8837
rect 3861 8828 3863 8833
rect 3866 8828 3868 8830
rect 3892 8828 3894 8830
rect 3913 8828 3915 8842
rect 3933 8837 3935 8842
rect 3938 8840 3940 8842
rect 3929 8833 3935 8837
rect 3933 8828 3935 8833
rect 3938 8828 3940 8830
rect 3956 8828 3958 8842
rect 4006 8837 4008 8842
rect 4011 8837 4013 8839
rect 4034 8833 4036 8855
rect 4006 8831 4008 8833
rect 4011 8828 4013 8833
rect 4034 8827 4036 8829
rect 2861 8822 2863 8824
rect 2877 8820 2879 8824
rect 2893 8822 2895 8824
rect 2916 8822 2918 8824
rect 2878 8816 2879 8820
rect 2921 8819 2923 8824
rect 2947 8820 2949 8824
rect 2968 8822 2970 8824
rect 2988 8822 2990 8824
rect 2877 8813 2879 8816
rect 2922 8815 2923 8819
rect 2948 8816 2949 8820
rect 2993 8819 2995 8824
rect 3011 8822 3013 8824
rect 3806 8822 3808 8824
rect 3822 8820 3824 8824
rect 3838 8822 3840 8824
rect 3861 8822 3863 8824
rect 2921 8813 2923 8815
rect 2947 8812 2949 8816
rect 2994 8815 2995 8819
rect 3823 8816 3824 8820
rect 3866 8819 3868 8824
rect 3892 8820 3894 8824
rect 3913 8822 3915 8824
rect 3933 8822 3935 8824
rect 2993 8813 2995 8815
rect 3822 8813 3824 8816
rect 3867 8815 3868 8819
rect 3893 8816 3894 8820
rect 3938 8819 3940 8824
rect 3956 8822 3958 8824
rect 3866 8813 3868 8815
rect 3892 8812 3894 8816
rect 3939 8815 3940 8819
rect 3938 8813 3940 8815
rect 2372 8795 2374 8797
rect 2377 8795 2379 8798
rect 2393 8795 2395 8797
rect 2409 8795 2411 8797
rect 2414 8795 2416 8798
rect 2435 8795 2437 8798
rect 2451 8795 2453 8798
rect 2467 8795 2469 8797
rect 2472 8795 2474 8798
rect 2488 8795 2490 8797
rect 2504 8795 2506 8797
rect 2509 8795 2511 8798
rect 2525 8795 2527 8797
rect 2541 8795 2543 8797
rect 2546 8795 2548 8798
rect 2567 8795 2569 8798
rect 2583 8795 2585 8798
rect 2599 8795 2601 8797
rect 2604 8795 2606 8798
rect 2620 8795 2622 8797
rect 2636 8795 2638 8797
rect 2641 8795 2643 8798
rect 2657 8795 2659 8797
rect 2673 8795 2675 8797
rect 2678 8795 2680 8798
rect 2699 8795 2701 8798
rect 2715 8795 2717 8798
rect 2731 8795 2733 8797
rect 2736 8795 2738 8798
rect 2752 8795 2754 8797
rect 3317 8795 3319 8797
rect 3322 8795 3324 8798
rect 3338 8795 3340 8797
rect 3354 8795 3356 8797
rect 3359 8795 3361 8798
rect 3380 8795 3382 8798
rect 3396 8795 3398 8798
rect 3412 8795 3414 8797
rect 3417 8795 3419 8798
rect 3433 8795 3435 8797
rect 3449 8795 3451 8797
rect 3454 8795 3456 8798
rect 3470 8795 3472 8797
rect 3486 8795 3488 8797
rect 3491 8795 3493 8798
rect 3512 8795 3514 8798
rect 3528 8795 3530 8798
rect 3544 8795 3546 8797
rect 3549 8795 3551 8798
rect 3565 8795 3567 8797
rect 3581 8795 3583 8797
rect 3586 8795 3588 8798
rect 3602 8795 3604 8797
rect 3618 8795 3620 8797
rect 3623 8795 3625 8798
rect 3644 8795 3646 8798
rect 3660 8795 3662 8798
rect 3676 8795 3678 8797
rect 3681 8795 3683 8798
rect 3697 8795 3699 8797
rect 2877 8790 2879 8793
rect 2921 8791 2923 8793
rect 2372 8782 2374 8787
rect 2377 8785 2379 8787
rect 2372 8768 2374 8778
rect 2377 8768 2379 8775
rect 2393 8768 2395 8787
rect 2409 8778 2411 8787
rect 2414 8785 2416 8787
rect 2435 8785 2437 8787
rect 2451 8784 2453 8787
rect 2409 8768 2411 8771
rect 2414 8768 2416 8770
rect 2435 8768 2437 8770
rect 2451 8768 2453 8780
rect 2467 8778 2469 8787
rect 2472 8785 2474 8787
rect 2467 8768 2469 8771
rect 2472 8768 2474 8770
rect 2488 8768 2490 8787
rect 2504 8784 2506 8787
rect 2509 8785 2511 8787
rect 2504 8768 2506 8780
rect 2509 8768 2511 8775
rect 2525 8768 2527 8787
rect 2541 8778 2543 8787
rect 2546 8785 2548 8787
rect 2567 8785 2569 8787
rect 2583 8784 2585 8787
rect 2541 8768 2543 8771
rect 2546 8768 2548 8770
rect 2567 8768 2569 8770
rect 2583 8768 2585 8780
rect 2599 8778 2601 8787
rect 2604 8785 2606 8787
rect 2599 8768 2601 8771
rect 2604 8768 2606 8770
rect 2620 8768 2622 8787
rect 2636 8784 2638 8787
rect 2641 8785 2643 8787
rect 2636 8768 2638 8780
rect 2641 8768 2643 8775
rect 2657 8768 2659 8787
rect 2673 8778 2675 8787
rect 2678 8785 2680 8787
rect 2699 8785 2701 8787
rect 2715 8784 2717 8787
rect 2673 8768 2675 8771
rect 2678 8768 2680 8770
rect 2699 8768 2701 8770
rect 2715 8768 2717 8780
rect 2731 8778 2733 8787
rect 2736 8785 2738 8787
rect 2752 8779 2754 8787
rect 2878 8786 2879 8790
rect 2922 8787 2923 8791
rect 2947 8790 2949 8794
rect 2993 8791 2995 8793
rect 2861 8782 2863 8784
rect 2877 8782 2879 8786
rect 2893 8782 2895 8784
rect 2916 8782 2918 8784
rect 2921 8782 2923 8787
rect 2948 8786 2949 8790
rect 2994 8787 2995 8791
rect 3138 8790 3140 8793
rect 3182 8791 3184 8793
rect 2947 8782 2949 8786
rect 2968 8782 2970 8784
rect 2988 8782 2990 8784
rect 2993 8782 2995 8787
rect 3139 8786 3140 8790
rect 3183 8787 3184 8791
rect 3208 8790 3210 8794
rect 3254 8791 3256 8793
rect 3011 8782 3013 8784
rect 3095 8782 3097 8785
rect 3113 8782 3115 8785
rect 3138 8782 3140 8786
rect 3154 8782 3156 8784
rect 3177 8782 3179 8784
rect 3182 8782 3184 8787
rect 3209 8786 3210 8790
rect 3255 8787 3256 8791
rect 3822 8790 3824 8793
rect 3866 8791 3868 8793
rect 3208 8782 3210 8786
rect 3229 8782 3231 8784
rect 3249 8782 3251 8784
rect 3254 8782 3256 8787
rect 3272 8782 3274 8784
rect 3317 8782 3319 8787
rect 3322 8785 3324 8787
rect 2731 8768 2733 8771
rect 2736 8768 2738 8770
rect 2752 8768 2754 8775
rect 2861 8764 2863 8778
rect 2877 8776 2879 8778
rect 2877 8764 2879 8766
rect 2893 8764 2895 8778
rect 2916 8773 2918 8778
rect 2921 8776 2923 8778
rect 2947 8776 2949 8778
rect 2912 8769 2918 8773
rect 2916 8764 2918 8769
rect 2921 8764 2923 8766
rect 2947 8764 2949 8766
rect 2968 8764 2970 8778
rect 2988 8773 2990 8778
rect 2993 8776 2995 8778
rect 2984 8769 2990 8773
rect 2988 8764 2990 8769
rect 2993 8764 2995 8766
rect 3011 8764 3013 8778
rect 3061 8775 3063 8778
rect 3066 8775 3068 8778
rect 3095 8773 3097 8778
rect 2372 8762 2374 8764
rect 2377 8761 2379 8764
rect 2393 8762 2395 8764
rect 2409 8762 2411 8764
rect 2414 8759 2416 8764
rect 2435 8759 2437 8764
rect 2451 8762 2453 8764
rect 2467 8762 2469 8764
rect 2472 8759 2474 8764
rect 2488 8762 2490 8764
rect 2504 8762 2506 8764
rect 2509 8761 2511 8764
rect 2525 8762 2527 8764
rect 2541 8762 2543 8764
rect 2546 8759 2548 8764
rect 2567 8759 2569 8764
rect 2583 8762 2585 8764
rect 2599 8762 2601 8764
rect 2604 8759 2606 8764
rect 2620 8762 2622 8764
rect 2636 8762 2638 8764
rect 2641 8761 2643 8764
rect 2657 8762 2659 8764
rect 2673 8762 2675 8764
rect 2678 8759 2680 8764
rect 2699 8759 2701 8764
rect 2715 8762 2717 8764
rect 2731 8762 2733 8764
rect 2736 8759 2738 8764
rect 2752 8762 2754 8764
rect 3061 8759 3063 8771
rect 3066 8769 3068 8771
rect 3095 8764 3097 8769
rect 3113 8764 3115 8778
rect 3138 8776 3140 8778
rect 3138 8764 3140 8766
rect 3154 8764 3156 8778
rect 3177 8773 3179 8778
rect 3182 8776 3184 8778
rect 3208 8776 3210 8778
rect 3173 8769 3179 8773
rect 3177 8764 3179 8769
rect 3182 8764 3184 8766
rect 3208 8764 3210 8766
rect 3229 8764 3231 8778
rect 3249 8773 3251 8778
rect 3254 8776 3256 8778
rect 3245 8769 3251 8773
rect 3249 8764 3251 8769
rect 3254 8764 3256 8766
rect 3272 8764 3274 8778
rect 3317 8768 3319 8778
rect 3322 8768 3324 8775
rect 3338 8768 3340 8787
rect 3354 8778 3356 8787
rect 3359 8785 3361 8787
rect 3380 8785 3382 8787
rect 3396 8784 3398 8787
rect 3354 8768 3356 8771
rect 3359 8768 3361 8770
rect 3380 8768 3382 8770
rect 3396 8768 3398 8780
rect 3412 8778 3414 8787
rect 3417 8785 3419 8787
rect 3412 8768 3414 8771
rect 3417 8768 3419 8770
rect 3433 8768 3435 8787
rect 3449 8784 3451 8787
rect 3454 8785 3456 8787
rect 3449 8768 3451 8780
rect 3454 8768 3456 8775
rect 3470 8768 3472 8787
rect 3486 8778 3488 8787
rect 3491 8785 3493 8787
rect 3512 8785 3514 8787
rect 3528 8784 3530 8787
rect 3486 8768 3488 8771
rect 3491 8768 3493 8770
rect 3512 8768 3514 8770
rect 3528 8768 3530 8780
rect 3544 8778 3546 8787
rect 3549 8785 3551 8787
rect 3544 8768 3546 8771
rect 3549 8768 3551 8770
rect 3565 8768 3567 8787
rect 3581 8784 3583 8787
rect 3586 8785 3588 8787
rect 3581 8768 3583 8780
rect 3586 8768 3588 8775
rect 3602 8768 3604 8787
rect 3618 8778 3620 8787
rect 3623 8785 3625 8787
rect 3644 8785 3646 8787
rect 3660 8784 3662 8787
rect 3618 8768 3620 8771
rect 3623 8768 3625 8770
rect 3644 8768 3646 8770
rect 3660 8768 3662 8780
rect 3676 8778 3678 8787
rect 3681 8785 3683 8787
rect 3697 8779 3699 8787
rect 3823 8786 3824 8790
rect 3867 8787 3868 8791
rect 3892 8790 3894 8794
rect 3938 8791 3940 8793
rect 3806 8782 3808 8784
rect 3822 8782 3824 8786
rect 3838 8782 3840 8784
rect 3861 8782 3863 8784
rect 3866 8782 3868 8787
rect 3893 8786 3894 8790
rect 3939 8787 3940 8791
rect 4083 8790 4085 8793
rect 4127 8791 4129 8793
rect 3892 8782 3894 8786
rect 3913 8782 3915 8784
rect 3933 8782 3935 8784
rect 3938 8782 3940 8787
rect 4084 8786 4085 8790
rect 4128 8787 4129 8791
rect 4153 8790 4155 8794
rect 4199 8791 4201 8793
rect 3956 8782 3958 8784
rect 4040 8782 4042 8785
rect 4058 8782 4060 8785
rect 4083 8782 4085 8786
rect 4099 8782 4101 8784
rect 4122 8782 4124 8784
rect 4127 8782 4129 8787
rect 4154 8786 4155 8790
rect 4200 8787 4201 8791
rect 4153 8782 4155 8786
rect 4174 8782 4176 8784
rect 4194 8782 4196 8784
rect 4199 8782 4201 8787
rect 4217 8782 4219 8784
rect 3676 8768 3678 8771
rect 3681 8768 3683 8770
rect 3697 8768 3699 8775
rect 3806 8764 3808 8778
rect 3822 8776 3824 8778
rect 3822 8764 3824 8766
rect 3838 8764 3840 8778
rect 3861 8773 3863 8778
rect 3866 8776 3868 8778
rect 3892 8776 3894 8778
rect 3857 8769 3863 8773
rect 3861 8764 3863 8769
rect 3866 8764 3868 8766
rect 3892 8764 3894 8766
rect 3913 8764 3915 8778
rect 3933 8773 3935 8778
rect 3938 8776 3940 8778
rect 3929 8769 3935 8773
rect 3933 8764 3935 8769
rect 3938 8764 3940 8766
rect 3956 8764 3958 8778
rect 4006 8775 4008 8778
rect 4011 8775 4013 8778
rect 4040 8773 4042 8778
rect 3066 8759 3068 8761
rect 2861 8754 2863 8756
rect 2877 8753 2879 8756
rect 2893 8754 2895 8756
rect 2916 8754 2918 8756
rect 2921 8753 2923 8756
rect 2947 8753 2949 8756
rect 2968 8753 2970 8756
rect 2988 8754 2990 8756
rect 2993 8753 2995 8756
rect 3011 8754 3013 8756
rect 2947 8749 2948 8753
rect 3317 8762 3319 8764
rect 3322 8761 3324 8764
rect 3338 8762 3340 8764
rect 3354 8762 3356 8764
rect 3359 8759 3361 8764
rect 3380 8759 3382 8764
rect 3396 8762 3398 8764
rect 3412 8762 3414 8764
rect 3417 8759 3419 8764
rect 3433 8762 3435 8764
rect 3449 8762 3451 8764
rect 3095 8753 3097 8756
rect 3061 8749 3063 8751
rect 2877 8746 2879 8749
rect 2921 8746 2923 8749
rect 2947 8746 2949 8749
rect 2993 8746 2995 8749
rect 3066 8746 3068 8751
rect 2487 8724 2489 8727
rect 2511 8724 2513 8727
rect 2487 8717 2489 8720
rect 2511 8717 2513 8720
rect 3113 8714 3115 8756
rect 3138 8753 3140 8756
rect 3154 8754 3156 8756
rect 3177 8754 3179 8756
rect 3182 8753 3184 8756
rect 3208 8753 3210 8756
rect 3229 8753 3231 8756
rect 3249 8754 3251 8756
rect 3254 8753 3256 8756
rect 3272 8754 3274 8756
rect 3454 8761 3456 8764
rect 3470 8762 3472 8764
rect 3486 8762 3488 8764
rect 3491 8759 3493 8764
rect 3512 8759 3514 8764
rect 3528 8762 3530 8764
rect 3544 8762 3546 8764
rect 3549 8759 3551 8764
rect 3565 8762 3567 8764
rect 3581 8762 3583 8764
rect 3586 8761 3588 8764
rect 3602 8762 3604 8764
rect 3618 8762 3620 8764
rect 3623 8759 3625 8764
rect 3644 8759 3646 8764
rect 3660 8762 3662 8764
rect 3676 8762 3678 8764
rect 3681 8759 3683 8764
rect 3697 8762 3699 8764
rect 4006 8759 4008 8771
rect 4011 8769 4013 8771
rect 4040 8764 4042 8769
rect 4058 8764 4060 8778
rect 4083 8776 4085 8778
rect 4083 8764 4085 8766
rect 4099 8764 4101 8778
rect 4122 8773 4124 8778
rect 4127 8776 4129 8778
rect 4153 8776 4155 8778
rect 4118 8769 4124 8773
rect 4122 8764 4124 8769
rect 4127 8764 4129 8766
rect 4153 8764 4155 8766
rect 4174 8764 4176 8778
rect 4194 8773 4196 8778
rect 4199 8776 4201 8778
rect 4190 8769 4196 8773
rect 4194 8764 4196 8769
rect 4199 8764 4201 8766
rect 4217 8764 4219 8778
rect 4011 8759 4013 8761
rect 3806 8754 3808 8756
rect 3822 8753 3824 8756
rect 3838 8754 3840 8756
rect 3861 8754 3863 8756
rect 3866 8753 3868 8756
rect 3892 8753 3894 8756
rect 3913 8753 3915 8756
rect 3933 8754 3935 8756
rect 3938 8753 3940 8756
rect 3956 8754 3958 8756
rect 3208 8749 3209 8753
rect 3138 8746 3140 8749
rect 3182 8746 3184 8749
rect 3208 8746 3210 8749
rect 3254 8746 3256 8749
rect 3892 8749 3893 8753
rect 4040 8753 4042 8756
rect 4006 8749 4008 8751
rect 3822 8746 3824 8749
rect 3866 8746 3868 8749
rect 3892 8746 3894 8749
rect 3938 8746 3940 8749
rect 4011 8746 4013 8751
rect 3432 8724 3434 8727
rect 3456 8724 3458 8727
rect 3281 8722 3284 8724
rect 3288 8722 3291 8724
rect 3432 8717 3434 8720
rect 3456 8717 3458 8720
rect 4058 8718 4060 8756
rect 4083 8753 4085 8756
rect 4099 8754 4101 8756
rect 4122 8754 4124 8756
rect 4127 8753 4129 8756
rect 4153 8753 4155 8756
rect 4174 8753 4176 8756
rect 4194 8754 4196 8756
rect 4199 8753 4201 8756
rect 4217 8754 4219 8756
rect 4153 8749 4154 8753
rect 4083 8746 4085 8749
rect 4127 8746 4129 8749
rect 4153 8746 4155 8749
rect 4199 8746 4201 8749
rect 4226 8722 4229 8724
rect 4233 8722 4236 8724
rect 2507 8711 2509 8713
rect 3452 8711 3454 8713
rect 2507 8704 2509 8707
rect 3452 8704 3454 8707
rect 2496 8693 2498 8695
rect 2502 8693 2521 8695
rect 3441 8693 3443 8695
rect 3447 8693 3466 8695
rect 2487 8688 2489 8690
rect 2511 8688 2513 8690
rect 3432 8688 3434 8690
rect 3456 8688 3458 8690
rect 2487 8681 2489 8684
rect 2511 8681 2513 8684
rect 3155 8683 3157 8685
rect 3160 8683 3162 8686
rect 3176 8683 3178 8685
rect 3192 8683 3194 8685
rect 3197 8683 3199 8686
rect 3218 8683 3220 8686
rect 3234 8683 3236 8686
rect 3250 8683 3252 8685
rect 3255 8683 3257 8686
rect 3271 8683 3273 8685
rect 3432 8681 3434 8684
rect 3456 8681 3458 8684
rect 4100 8683 4102 8685
rect 4105 8683 4107 8686
rect 4121 8683 4123 8685
rect 4137 8683 4139 8685
rect 4142 8683 4144 8686
rect 4163 8683 4165 8686
rect 4179 8683 4181 8686
rect 4195 8683 4197 8685
rect 4200 8683 4202 8686
rect 4216 8683 4218 8685
rect 3155 8670 3157 8675
rect 3160 8673 3162 8675
rect 3155 8656 3157 8666
rect 3160 8656 3162 8663
rect 3176 8656 3178 8675
rect 3192 8666 3194 8675
rect 3197 8673 3199 8675
rect 3218 8673 3220 8675
rect 3234 8672 3236 8675
rect 3192 8656 3194 8659
rect 3197 8656 3199 8658
rect 3218 8656 3220 8658
rect 3234 8656 3236 8668
rect 3250 8666 3252 8675
rect 3255 8673 3257 8675
rect 3250 8656 3252 8659
rect 3255 8656 3257 8658
rect 3271 8656 3273 8675
rect 4100 8670 4102 8675
rect 4105 8673 4107 8675
rect 4100 8656 4102 8666
rect 4105 8656 4107 8663
rect 4121 8656 4123 8675
rect 4137 8666 4139 8675
rect 4142 8673 4144 8675
rect 4163 8673 4165 8675
rect 4179 8672 4181 8675
rect 4137 8656 4139 8659
rect 4142 8656 4144 8658
rect 4163 8656 4165 8658
rect 4179 8656 4181 8668
rect 4195 8666 4197 8675
rect 4200 8673 4202 8675
rect 4195 8656 4197 8659
rect 4200 8656 4202 8658
rect 4216 8656 4218 8675
rect 2372 8653 2374 8655
rect 2377 8653 2379 8656
rect 2393 8653 2395 8655
rect 2409 8653 2411 8655
rect 2414 8653 2416 8656
rect 2435 8653 2437 8656
rect 2451 8653 2453 8656
rect 2467 8653 2469 8655
rect 2472 8653 2474 8656
rect 2488 8653 2490 8655
rect 2504 8653 2506 8655
rect 2509 8653 2511 8656
rect 2525 8653 2527 8655
rect 2541 8653 2543 8655
rect 2546 8653 2548 8656
rect 2567 8653 2569 8656
rect 2583 8653 2585 8656
rect 2599 8653 2601 8655
rect 2604 8653 2606 8656
rect 2620 8653 2622 8655
rect 2636 8653 2638 8655
rect 2641 8653 2643 8656
rect 2657 8653 2659 8655
rect 2673 8653 2675 8655
rect 2678 8653 2680 8656
rect 2699 8653 2701 8656
rect 2715 8653 2717 8656
rect 2731 8653 2733 8655
rect 2736 8653 2738 8656
rect 2752 8653 2754 8655
rect 3317 8653 3319 8655
rect 3322 8653 3324 8656
rect 3338 8653 3340 8655
rect 3354 8653 3356 8655
rect 3359 8653 3361 8656
rect 3380 8653 3382 8656
rect 3396 8653 3398 8656
rect 3412 8653 3414 8655
rect 3417 8653 3419 8656
rect 3433 8653 3435 8655
rect 3449 8653 3451 8655
rect 3454 8653 3456 8656
rect 3470 8653 3472 8655
rect 3486 8653 3488 8655
rect 3491 8653 3493 8656
rect 3512 8653 3514 8656
rect 3528 8653 3530 8656
rect 3544 8653 3546 8655
rect 3549 8653 3551 8656
rect 3565 8653 3567 8655
rect 3581 8653 3583 8655
rect 3586 8653 3588 8656
rect 3602 8653 3604 8655
rect 3618 8653 3620 8655
rect 3623 8653 3625 8656
rect 3644 8653 3646 8656
rect 3660 8653 3662 8656
rect 3676 8653 3678 8655
rect 3681 8653 3683 8656
rect 3697 8653 3699 8655
rect 3155 8650 3157 8652
rect 3160 8649 3162 8652
rect 3176 8650 3178 8652
rect 3192 8650 3194 8652
rect 3197 8647 3199 8652
rect 3218 8647 3220 8652
rect 3234 8650 3236 8652
rect 3250 8650 3252 8652
rect 3255 8647 3257 8652
rect 3271 8650 3273 8652
rect 2372 8640 2374 8645
rect 2377 8643 2379 8645
rect 2372 8626 2374 8636
rect 2377 8626 2379 8633
rect 2393 8626 2395 8645
rect 2409 8636 2411 8645
rect 2414 8643 2416 8645
rect 2435 8643 2437 8645
rect 2451 8642 2453 8645
rect 2409 8626 2411 8629
rect 2414 8626 2416 8628
rect 2435 8626 2437 8628
rect 2451 8626 2453 8638
rect 2467 8636 2469 8645
rect 2472 8643 2474 8645
rect 2467 8626 2469 8629
rect 2472 8626 2474 8628
rect 2488 8626 2490 8645
rect 2504 8642 2506 8645
rect 2509 8643 2511 8645
rect 2504 8626 2506 8638
rect 2509 8626 2511 8633
rect 2525 8626 2527 8645
rect 2541 8636 2543 8645
rect 2546 8643 2548 8645
rect 2567 8643 2569 8645
rect 2583 8642 2585 8645
rect 2541 8626 2543 8629
rect 2546 8626 2548 8628
rect 2567 8626 2569 8628
rect 2583 8626 2585 8638
rect 2599 8636 2601 8645
rect 2604 8643 2606 8645
rect 2599 8626 2601 8629
rect 2604 8626 2606 8628
rect 2620 8626 2622 8645
rect 2636 8642 2638 8645
rect 2641 8643 2643 8645
rect 2636 8626 2638 8638
rect 2641 8626 2643 8633
rect 2657 8626 2659 8645
rect 2673 8636 2675 8645
rect 2678 8643 2680 8645
rect 2699 8643 2701 8645
rect 2715 8642 2717 8645
rect 2673 8626 2675 8629
rect 2678 8626 2680 8628
rect 2699 8626 2701 8628
rect 2715 8626 2717 8638
rect 2731 8636 2733 8645
rect 2736 8643 2738 8645
rect 2752 8637 2754 8645
rect 4100 8650 4102 8652
rect 4105 8649 4107 8652
rect 4121 8650 4123 8652
rect 4137 8650 4139 8652
rect 4142 8647 4144 8652
rect 4163 8647 4165 8652
rect 4179 8650 4181 8652
rect 4195 8650 4197 8652
rect 4200 8647 4202 8652
rect 4216 8650 4218 8652
rect 3317 8640 3319 8645
rect 3322 8643 3324 8645
rect 2731 8626 2733 8629
rect 2736 8626 2738 8628
rect 2752 8626 2754 8633
rect 3317 8626 3319 8636
rect 3322 8626 3324 8633
rect 3338 8626 3340 8645
rect 3354 8636 3356 8645
rect 3359 8643 3361 8645
rect 3380 8643 3382 8645
rect 3396 8642 3398 8645
rect 3354 8626 3356 8629
rect 3359 8626 3361 8628
rect 3380 8626 3382 8628
rect 3396 8626 3398 8638
rect 3412 8636 3414 8645
rect 3417 8643 3419 8645
rect 3412 8626 3414 8629
rect 3417 8626 3419 8628
rect 3433 8626 3435 8645
rect 3449 8642 3451 8645
rect 3454 8643 3456 8645
rect 3449 8626 3451 8638
rect 3454 8626 3456 8633
rect 3470 8626 3472 8645
rect 3486 8636 3488 8645
rect 3491 8643 3493 8645
rect 3512 8643 3514 8645
rect 3528 8642 3530 8645
rect 3486 8626 3488 8629
rect 3491 8626 3493 8628
rect 3512 8626 3514 8628
rect 3528 8626 3530 8638
rect 3544 8636 3546 8645
rect 3549 8643 3551 8645
rect 3544 8626 3546 8629
rect 3549 8626 3551 8628
rect 3565 8626 3567 8645
rect 3581 8642 3583 8645
rect 3586 8643 3588 8645
rect 3581 8626 3583 8638
rect 3586 8626 3588 8633
rect 3602 8626 3604 8645
rect 3618 8636 3620 8645
rect 3623 8643 3625 8645
rect 3644 8643 3646 8645
rect 3660 8642 3662 8645
rect 3618 8626 3620 8629
rect 3623 8626 3625 8628
rect 3644 8626 3646 8628
rect 3660 8626 3662 8638
rect 3676 8636 3678 8645
rect 3681 8643 3683 8645
rect 3697 8637 3699 8645
rect 3676 8626 3678 8629
rect 3681 8626 3683 8628
rect 3697 8626 3699 8633
rect 2372 8620 2374 8622
rect 2377 8619 2379 8622
rect 2393 8620 2395 8622
rect 2409 8620 2411 8622
rect 2414 8617 2416 8622
rect 2435 8617 2437 8622
rect 2451 8620 2453 8622
rect 2467 8620 2469 8622
rect 2472 8617 2474 8622
rect 2488 8620 2490 8622
rect 2504 8620 2506 8622
rect 2509 8619 2511 8622
rect 2525 8620 2527 8622
rect 2541 8620 2543 8622
rect 2546 8617 2548 8622
rect 2567 8617 2569 8622
rect 2583 8620 2585 8622
rect 2599 8620 2601 8622
rect 2604 8617 2606 8622
rect 2620 8620 2622 8622
rect 2636 8620 2638 8622
rect 2641 8619 2643 8622
rect 2657 8620 2659 8622
rect 2673 8620 2675 8622
rect 2678 8617 2680 8622
rect 2699 8617 2701 8622
rect 2715 8620 2717 8622
rect 2731 8620 2733 8622
rect 2736 8617 2738 8622
rect 2752 8620 2754 8622
rect 3317 8620 3319 8622
rect 3322 8619 3324 8622
rect 3338 8620 3340 8622
rect 3354 8620 3356 8622
rect 3359 8617 3361 8622
rect 3380 8617 3382 8622
rect 3396 8620 3398 8622
rect 3412 8620 3414 8622
rect 3417 8617 3419 8622
rect 3433 8620 3435 8622
rect 3449 8620 3451 8622
rect 3454 8619 3456 8622
rect 3470 8620 3472 8622
rect 3486 8620 3488 8622
rect 3491 8617 3493 8622
rect 3512 8617 3514 8622
rect 3528 8620 3530 8622
rect 3544 8620 3546 8622
rect 3549 8617 3551 8622
rect 3565 8620 3567 8622
rect 3581 8620 3583 8622
rect 3586 8619 3588 8622
rect 3602 8620 3604 8622
rect 3618 8620 3620 8622
rect 3623 8617 3625 8622
rect 3644 8617 3646 8622
rect 3660 8620 3662 8622
rect 3676 8620 3678 8622
rect 3681 8617 3683 8622
rect 3697 8620 3699 8622
rect 3155 8597 3157 8599
rect 3160 8597 3162 8600
rect 3176 8597 3178 8599
rect 3192 8597 3194 8599
rect 3197 8597 3199 8600
rect 3218 8597 3220 8600
rect 3234 8597 3236 8600
rect 3250 8597 3252 8599
rect 3255 8597 3257 8600
rect 3271 8597 3273 8599
rect 4100 8597 4102 8599
rect 4105 8597 4107 8600
rect 4121 8597 4123 8599
rect 4137 8597 4139 8599
rect 4142 8597 4144 8600
rect 4163 8597 4165 8600
rect 4179 8597 4181 8600
rect 4195 8597 4197 8599
rect 4200 8597 4202 8600
rect 4216 8597 4218 8599
rect 3155 8584 3157 8589
rect 3160 8587 3162 8589
rect 3155 8570 3157 8580
rect 3160 8570 3162 8577
rect 3176 8570 3178 8589
rect 3192 8580 3194 8589
rect 3197 8587 3199 8589
rect 3218 8587 3220 8589
rect 3234 8586 3236 8589
rect 3192 8570 3194 8573
rect 3197 8570 3199 8572
rect 3218 8570 3220 8572
rect 3234 8570 3236 8582
rect 3250 8580 3252 8589
rect 3255 8587 3257 8589
rect 3250 8570 3252 8573
rect 3255 8570 3257 8572
rect 3271 8570 3273 8589
rect 4100 8584 4102 8589
rect 4105 8587 4107 8589
rect 3293 8576 3296 8578
rect 3300 8576 3303 8578
rect 4100 8570 4102 8580
rect 4105 8570 4107 8577
rect 4121 8570 4123 8589
rect 4137 8580 4139 8589
rect 4142 8587 4144 8589
rect 4163 8587 4165 8589
rect 4179 8586 4181 8589
rect 4137 8570 4139 8573
rect 4142 8570 4144 8572
rect 4163 8570 4165 8572
rect 4179 8570 4181 8582
rect 4195 8580 4197 8589
rect 4200 8587 4202 8589
rect 4195 8570 4197 8573
rect 4200 8570 4202 8572
rect 4216 8570 4218 8589
rect 4238 8576 4241 8578
rect 4245 8576 4248 8578
rect 2372 8567 2374 8569
rect 2377 8567 2379 8570
rect 2393 8567 2395 8569
rect 2409 8567 2411 8569
rect 2414 8567 2416 8570
rect 2435 8567 2437 8570
rect 2451 8567 2453 8570
rect 2467 8567 2469 8569
rect 2472 8567 2474 8570
rect 2488 8567 2490 8569
rect 2504 8567 2506 8569
rect 2509 8567 2511 8570
rect 2525 8567 2527 8569
rect 2541 8567 2543 8569
rect 2546 8567 2548 8570
rect 2567 8567 2569 8570
rect 2583 8567 2585 8570
rect 2599 8567 2601 8569
rect 2604 8567 2606 8570
rect 2620 8567 2622 8569
rect 2636 8567 2638 8569
rect 2641 8567 2643 8570
rect 2657 8567 2659 8569
rect 2673 8567 2675 8569
rect 2678 8567 2680 8570
rect 2699 8567 2701 8570
rect 2715 8567 2717 8570
rect 2731 8567 2733 8569
rect 2736 8567 2738 8570
rect 2752 8567 2754 8569
rect 3317 8567 3319 8569
rect 3322 8567 3324 8570
rect 3338 8567 3340 8569
rect 3354 8567 3356 8569
rect 3359 8567 3361 8570
rect 3380 8567 3382 8570
rect 3396 8567 3398 8570
rect 3412 8567 3414 8569
rect 3417 8567 3419 8570
rect 3433 8567 3435 8569
rect 3449 8567 3451 8569
rect 3454 8567 3456 8570
rect 3470 8567 3472 8569
rect 3486 8567 3488 8569
rect 3491 8567 3493 8570
rect 3512 8567 3514 8570
rect 3528 8567 3530 8570
rect 3544 8567 3546 8569
rect 3549 8567 3551 8570
rect 3565 8567 3567 8569
rect 3581 8567 3583 8569
rect 3586 8567 3588 8570
rect 3602 8567 3604 8569
rect 3618 8567 3620 8569
rect 3623 8567 3625 8570
rect 3644 8567 3646 8570
rect 3660 8567 3662 8570
rect 3676 8567 3678 8569
rect 3681 8567 3683 8570
rect 3697 8567 3699 8569
rect 3155 8564 3157 8566
rect 3160 8563 3162 8566
rect 3176 8564 3178 8566
rect 3192 8564 3194 8566
rect 3197 8561 3199 8566
rect 3218 8561 3220 8566
rect 3234 8564 3236 8566
rect 3250 8564 3252 8566
rect 3255 8561 3257 8566
rect 3271 8564 3273 8566
rect 2372 8554 2374 8559
rect 2377 8557 2379 8559
rect 2372 8540 2374 8550
rect 2377 8540 2379 8547
rect 2393 8540 2395 8559
rect 2409 8550 2411 8559
rect 2414 8557 2416 8559
rect 2435 8557 2437 8559
rect 2451 8556 2453 8559
rect 2409 8540 2411 8543
rect 2414 8540 2416 8542
rect 2435 8540 2437 8542
rect 2451 8540 2453 8552
rect 2467 8550 2469 8559
rect 2472 8557 2474 8559
rect 2467 8540 2469 8543
rect 2472 8540 2474 8542
rect 2488 8540 2490 8559
rect 2504 8556 2506 8559
rect 2509 8557 2511 8559
rect 2504 8540 2506 8552
rect 2509 8540 2511 8547
rect 2525 8540 2527 8559
rect 2541 8550 2543 8559
rect 2546 8557 2548 8559
rect 2567 8557 2569 8559
rect 2583 8556 2585 8559
rect 2541 8540 2543 8543
rect 2546 8540 2548 8542
rect 2567 8540 2569 8542
rect 2583 8540 2585 8552
rect 2599 8550 2601 8559
rect 2604 8557 2606 8559
rect 2599 8540 2601 8543
rect 2604 8540 2606 8542
rect 2620 8540 2622 8559
rect 2636 8556 2638 8559
rect 2641 8557 2643 8559
rect 2636 8540 2638 8552
rect 2641 8540 2643 8547
rect 2657 8540 2659 8559
rect 2673 8550 2675 8559
rect 2678 8557 2680 8559
rect 2699 8557 2701 8559
rect 2715 8556 2717 8559
rect 2673 8540 2675 8543
rect 2678 8540 2680 8542
rect 2699 8540 2701 8542
rect 2715 8540 2717 8552
rect 2731 8550 2733 8559
rect 2736 8557 2738 8559
rect 2752 8551 2754 8559
rect 4100 8564 4102 8566
rect 4105 8563 4107 8566
rect 4121 8564 4123 8566
rect 4137 8564 4139 8566
rect 4142 8561 4144 8566
rect 4163 8561 4165 8566
rect 4179 8564 4181 8566
rect 4195 8564 4197 8566
rect 4200 8561 4202 8566
rect 4216 8564 4218 8566
rect 3317 8554 3319 8559
rect 3322 8557 3324 8559
rect 2731 8540 2733 8543
rect 2736 8540 2738 8542
rect 2752 8540 2754 8547
rect 3317 8540 3319 8550
rect 3322 8540 3324 8547
rect 3338 8540 3340 8559
rect 3354 8550 3356 8559
rect 3359 8557 3361 8559
rect 3380 8557 3382 8559
rect 3396 8556 3398 8559
rect 3354 8540 3356 8543
rect 3359 8540 3361 8542
rect 3380 8540 3382 8542
rect 3396 8540 3398 8552
rect 3412 8550 3414 8559
rect 3417 8557 3419 8559
rect 3412 8540 3414 8543
rect 3417 8540 3419 8542
rect 3433 8540 3435 8559
rect 3449 8556 3451 8559
rect 3454 8557 3456 8559
rect 3449 8540 3451 8552
rect 3454 8540 3456 8547
rect 3470 8540 3472 8559
rect 3486 8550 3488 8559
rect 3491 8557 3493 8559
rect 3512 8557 3514 8559
rect 3528 8556 3530 8559
rect 3486 8540 3488 8543
rect 3491 8540 3493 8542
rect 3512 8540 3514 8542
rect 3528 8540 3530 8552
rect 3544 8550 3546 8559
rect 3549 8557 3551 8559
rect 3544 8540 3546 8543
rect 3549 8540 3551 8542
rect 3565 8540 3567 8559
rect 3581 8556 3583 8559
rect 3586 8557 3588 8559
rect 3581 8540 3583 8552
rect 3586 8540 3588 8547
rect 3602 8540 3604 8559
rect 3618 8550 3620 8559
rect 3623 8557 3625 8559
rect 3644 8557 3646 8559
rect 3660 8556 3662 8559
rect 3618 8540 3620 8543
rect 3623 8540 3625 8542
rect 3644 8540 3646 8542
rect 3660 8540 3662 8552
rect 3676 8550 3678 8559
rect 3681 8557 3683 8559
rect 3697 8551 3699 8559
rect 3676 8540 3678 8543
rect 3681 8540 3683 8542
rect 3697 8540 3699 8547
rect 2372 8534 2374 8536
rect 2377 8533 2379 8536
rect 2393 8534 2395 8536
rect 2409 8534 2411 8536
rect 2414 8531 2416 8536
rect 2435 8531 2437 8536
rect 2451 8534 2453 8536
rect 2467 8534 2469 8536
rect 2472 8531 2474 8536
rect 2488 8534 2490 8536
rect 2504 8534 2506 8536
rect 2509 8533 2511 8536
rect 2525 8534 2527 8536
rect 2541 8534 2543 8536
rect 2546 8531 2548 8536
rect 2567 8531 2569 8536
rect 2583 8534 2585 8536
rect 2599 8534 2601 8536
rect 2604 8531 2606 8536
rect 2620 8534 2622 8536
rect 2636 8534 2638 8536
rect 2641 8533 2643 8536
rect 2657 8534 2659 8536
rect 2673 8534 2675 8536
rect 2678 8531 2680 8536
rect 2699 8531 2701 8536
rect 2715 8534 2717 8536
rect 2731 8534 2733 8536
rect 2736 8531 2738 8536
rect 2752 8534 2754 8536
rect 3317 8534 3319 8536
rect 3322 8533 3324 8536
rect 3338 8534 3340 8536
rect 3354 8534 3356 8536
rect 3359 8531 3361 8536
rect 3380 8531 3382 8536
rect 3396 8534 3398 8536
rect 3412 8534 3414 8536
rect 3417 8531 3419 8536
rect 3433 8534 3435 8536
rect 3449 8534 3451 8536
rect 3454 8533 3456 8536
rect 3470 8534 3472 8536
rect 3486 8534 3488 8536
rect 3491 8531 3493 8536
rect 3512 8531 3514 8536
rect 3528 8534 3530 8536
rect 3544 8534 3546 8536
rect 3549 8531 3551 8536
rect 3565 8534 3567 8536
rect 3581 8534 3583 8536
rect 3586 8533 3588 8536
rect 3602 8534 3604 8536
rect 3618 8534 3620 8536
rect 3623 8531 3625 8536
rect 3644 8531 3646 8536
rect 3660 8534 3662 8536
rect 3676 8534 3678 8536
rect 3681 8531 3683 8536
rect 3697 8534 3699 8536
rect 2604 8496 2606 8499
rect 2628 8496 2630 8499
rect 3549 8496 3551 8499
rect 3573 8496 3575 8499
rect 2604 8490 2606 8492
rect 2628 8490 2630 8492
rect 3549 8490 3551 8492
rect 3573 8490 3575 8492
rect 2624 8485 2626 8487
rect 3569 8485 3571 8487
rect 2624 8478 2626 8481
rect 3569 8478 3571 8481
rect 2613 8467 2615 8469
rect 2619 8467 2638 8469
rect 3558 8467 3560 8469
rect 3564 8467 3583 8469
rect 2604 8462 2606 8464
rect 2628 8462 2630 8464
rect 3549 8462 3551 8464
rect 3573 8462 3575 8464
rect 2604 8455 2606 8458
rect 2628 8455 2630 8458
rect 3549 8455 3551 8458
rect 3573 8455 3575 8458
rect 2372 8427 2374 8429
rect 2377 8427 2379 8430
rect 2393 8427 2395 8429
rect 2409 8427 2411 8429
rect 2414 8427 2416 8430
rect 2435 8427 2437 8430
rect 2451 8427 2453 8430
rect 2467 8427 2469 8429
rect 2472 8427 2474 8430
rect 2488 8427 2490 8429
rect 2504 8427 2506 8429
rect 2509 8427 2511 8430
rect 2525 8427 2527 8429
rect 2541 8427 2543 8429
rect 2546 8427 2548 8430
rect 2567 8427 2569 8430
rect 2583 8427 2585 8430
rect 2599 8427 2601 8429
rect 2604 8427 2606 8430
rect 2620 8427 2622 8429
rect 2636 8427 2638 8429
rect 2641 8427 2643 8430
rect 2657 8427 2659 8429
rect 2673 8427 2675 8429
rect 2678 8427 2680 8430
rect 2699 8427 2701 8430
rect 2715 8427 2717 8430
rect 2731 8427 2733 8429
rect 2736 8427 2738 8430
rect 2752 8427 2754 8429
rect 3317 8427 3319 8429
rect 3322 8427 3324 8430
rect 3338 8427 3340 8429
rect 3354 8427 3356 8429
rect 3359 8427 3361 8430
rect 3380 8427 3382 8430
rect 3396 8427 3398 8430
rect 3412 8427 3414 8429
rect 3417 8427 3419 8430
rect 3433 8427 3435 8429
rect 3449 8427 3451 8429
rect 3454 8427 3456 8430
rect 3470 8427 3472 8429
rect 3486 8427 3488 8429
rect 3491 8427 3493 8430
rect 3512 8427 3514 8430
rect 3528 8427 3530 8430
rect 3544 8427 3546 8429
rect 3549 8427 3551 8430
rect 3565 8427 3567 8429
rect 3581 8427 3583 8429
rect 3586 8427 3588 8430
rect 3602 8427 3604 8429
rect 3618 8427 3620 8429
rect 3623 8427 3625 8430
rect 3644 8427 3646 8430
rect 3660 8427 3662 8430
rect 3676 8427 3678 8429
rect 3681 8427 3683 8430
rect 3697 8427 3699 8429
rect 2372 8414 2374 8419
rect 2377 8417 2379 8419
rect 2372 8400 2374 8410
rect 2377 8400 2379 8407
rect 2393 8400 2395 8419
rect 2409 8410 2411 8419
rect 2414 8417 2416 8419
rect 2435 8417 2437 8419
rect 2451 8416 2453 8419
rect 2409 8400 2411 8403
rect 2414 8400 2416 8402
rect 2435 8400 2437 8402
rect 2451 8400 2453 8412
rect 2467 8410 2469 8419
rect 2472 8417 2474 8419
rect 2467 8400 2469 8403
rect 2472 8400 2474 8402
rect 2488 8400 2490 8419
rect 2504 8416 2506 8419
rect 2509 8417 2511 8419
rect 2504 8400 2506 8412
rect 2509 8400 2511 8407
rect 2525 8400 2527 8419
rect 2541 8410 2543 8419
rect 2546 8417 2548 8419
rect 2567 8417 2569 8419
rect 2583 8416 2585 8419
rect 2541 8400 2543 8403
rect 2546 8400 2548 8402
rect 2567 8400 2569 8402
rect 2583 8400 2585 8412
rect 2599 8410 2601 8419
rect 2604 8417 2606 8419
rect 2599 8400 2601 8403
rect 2604 8400 2606 8402
rect 2620 8400 2622 8419
rect 2636 8416 2638 8419
rect 2641 8417 2643 8419
rect 2636 8400 2638 8412
rect 2641 8400 2643 8407
rect 2657 8400 2659 8419
rect 2673 8410 2675 8419
rect 2678 8417 2680 8419
rect 2699 8417 2701 8419
rect 2715 8416 2717 8419
rect 2673 8400 2675 8403
rect 2678 8400 2680 8402
rect 2699 8400 2701 8402
rect 2715 8400 2717 8412
rect 2731 8410 2733 8419
rect 2736 8417 2738 8419
rect 2752 8411 2754 8419
rect 3317 8414 3319 8419
rect 3322 8417 3324 8419
rect 2731 8400 2733 8403
rect 2736 8400 2738 8402
rect 2752 8400 2754 8407
rect 3317 8400 3319 8410
rect 3322 8400 3324 8407
rect 3338 8400 3340 8419
rect 3354 8410 3356 8419
rect 3359 8417 3361 8419
rect 3380 8417 3382 8419
rect 3396 8416 3398 8419
rect 3354 8400 3356 8403
rect 3359 8400 3361 8402
rect 3380 8400 3382 8402
rect 3396 8400 3398 8412
rect 3412 8410 3414 8419
rect 3417 8417 3419 8419
rect 3412 8400 3414 8403
rect 3417 8400 3419 8402
rect 3433 8400 3435 8419
rect 3449 8416 3451 8419
rect 3454 8417 3456 8419
rect 3449 8400 3451 8412
rect 3454 8400 3456 8407
rect 3470 8400 3472 8419
rect 3486 8410 3488 8419
rect 3491 8417 3493 8419
rect 3512 8417 3514 8419
rect 3528 8416 3530 8419
rect 3486 8400 3488 8403
rect 3491 8400 3493 8402
rect 3512 8400 3514 8402
rect 3528 8400 3530 8412
rect 3544 8410 3546 8419
rect 3549 8417 3551 8419
rect 3544 8400 3546 8403
rect 3549 8400 3551 8402
rect 3565 8400 3567 8419
rect 3581 8416 3583 8419
rect 3586 8417 3588 8419
rect 3581 8400 3583 8412
rect 3586 8400 3588 8407
rect 3602 8400 3604 8419
rect 3618 8410 3620 8419
rect 3623 8417 3625 8419
rect 3644 8417 3646 8419
rect 3660 8416 3662 8419
rect 3618 8400 3620 8403
rect 3623 8400 3625 8402
rect 3644 8400 3646 8402
rect 3660 8400 3662 8412
rect 3676 8410 3678 8419
rect 3681 8417 3683 8419
rect 3697 8411 3699 8419
rect 3676 8400 3678 8403
rect 3681 8400 3683 8402
rect 3697 8400 3699 8407
rect 2372 8394 2374 8396
rect 2377 8393 2379 8396
rect 2393 8394 2395 8396
rect 2409 8394 2411 8396
rect 2414 8391 2416 8396
rect 2435 8391 2437 8396
rect 2451 8394 2453 8396
rect 2467 8394 2469 8396
rect 2472 8391 2474 8396
rect 2488 8394 2490 8396
rect 2504 8394 2506 8396
rect 2509 8393 2511 8396
rect 2525 8394 2527 8396
rect 2541 8394 2543 8396
rect 2546 8391 2548 8396
rect 2567 8391 2569 8396
rect 2583 8394 2585 8396
rect 2599 8394 2601 8396
rect 2604 8391 2606 8396
rect 2620 8394 2622 8396
rect 2636 8394 2638 8396
rect 2641 8393 2643 8396
rect 2657 8394 2659 8396
rect 2673 8394 2675 8396
rect 2678 8391 2680 8396
rect 2699 8391 2701 8396
rect 2715 8394 2717 8396
rect 2731 8394 2733 8396
rect 2736 8391 2738 8396
rect 2752 8394 2754 8396
rect 3317 8394 3319 8396
rect 3322 8393 3324 8396
rect 3338 8394 3340 8396
rect 3354 8394 3356 8396
rect 3359 8391 3361 8396
rect 3380 8391 3382 8396
rect 3396 8394 3398 8396
rect 3412 8394 3414 8396
rect 3417 8391 3419 8396
rect 3433 8394 3435 8396
rect 3449 8394 3451 8396
rect 3454 8393 3456 8396
rect 3470 8394 3472 8396
rect 3486 8394 3488 8396
rect 3491 8391 3493 8396
rect 3512 8391 3514 8396
rect 3528 8394 3530 8396
rect 3544 8394 3546 8396
rect 3549 8391 3551 8396
rect 3565 8394 3567 8396
rect 3581 8394 3583 8396
rect 3586 8393 3588 8396
rect 3602 8394 3604 8396
rect 3618 8394 3620 8396
rect 3623 8391 3625 8396
rect 3644 8391 3646 8396
rect 3660 8394 3662 8396
rect 3676 8394 3678 8396
rect 3681 8391 3683 8396
rect 3697 8394 3699 8396
rect 2856 8348 2858 8350
rect 2861 8348 2863 8351
rect 2877 8348 2879 8350
rect 2893 8348 2895 8350
rect 2898 8348 2900 8351
rect 2919 8348 2921 8351
rect 2935 8348 2937 8351
rect 2951 8348 2953 8350
rect 2956 8348 2958 8351
rect 2972 8348 2974 8350
rect 2988 8348 2990 8350
rect 2993 8348 2995 8351
rect 3009 8348 3011 8350
rect 3025 8348 3027 8350
rect 3030 8348 3032 8351
rect 3051 8348 3053 8351
rect 3067 8348 3069 8351
rect 3083 8348 3085 8350
rect 3088 8348 3090 8351
rect 3104 8348 3106 8350
rect 3120 8348 3122 8350
rect 3125 8348 3127 8351
rect 3141 8348 3143 8350
rect 3157 8348 3159 8350
rect 3162 8348 3164 8351
rect 3183 8348 3185 8351
rect 3199 8348 3201 8351
rect 3215 8348 3217 8350
rect 3220 8348 3222 8351
rect 3236 8348 3238 8350
rect 3252 8348 3254 8350
rect 3257 8348 3259 8351
rect 3273 8348 3275 8350
rect 3289 8348 3291 8350
rect 3294 8348 3296 8351
rect 3315 8348 3317 8351
rect 3331 8348 3333 8351
rect 3347 8348 3349 8350
rect 3352 8348 3354 8351
rect 3368 8348 3370 8350
rect 3801 8348 3803 8350
rect 3806 8348 3808 8351
rect 3822 8348 3824 8350
rect 3838 8348 3840 8350
rect 3843 8348 3845 8351
rect 3864 8348 3866 8351
rect 3880 8348 3882 8351
rect 3896 8348 3898 8350
rect 3901 8348 3903 8351
rect 3917 8348 3919 8350
rect 3933 8348 3935 8350
rect 3938 8348 3940 8351
rect 3954 8348 3956 8350
rect 3970 8348 3972 8350
rect 3975 8348 3977 8351
rect 3996 8348 3998 8351
rect 4012 8348 4014 8351
rect 4028 8348 4030 8350
rect 4033 8348 4035 8351
rect 4049 8348 4051 8350
rect 4065 8348 4067 8350
rect 4070 8348 4072 8351
rect 4086 8348 4088 8350
rect 4102 8348 4104 8350
rect 4107 8348 4109 8351
rect 4128 8348 4130 8351
rect 4144 8348 4146 8351
rect 4160 8348 4162 8350
rect 4165 8348 4167 8351
rect 4181 8348 4183 8350
rect 4197 8348 4199 8350
rect 4202 8348 4204 8351
rect 4218 8348 4220 8350
rect 4234 8348 4236 8350
rect 4239 8348 4241 8351
rect 4260 8348 4262 8351
rect 4276 8348 4278 8351
rect 4292 8348 4294 8350
rect 4297 8348 4299 8351
rect 4313 8348 4315 8350
rect 2856 8335 2858 8340
rect 2861 8338 2863 8340
rect 2856 8321 2858 8331
rect 2861 8321 2863 8328
rect 2877 8321 2879 8340
rect 2893 8331 2895 8340
rect 2898 8338 2900 8340
rect 2919 8338 2921 8340
rect 2935 8337 2937 8340
rect 2893 8321 2895 8324
rect 2898 8321 2900 8323
rect 2919 8321 2921 8323
rect 2935 8321 2937 8333
rect 2951 8331 2953 8340
rect 2956 8338 2958 8340
rect 2972 8332 2974 8340
rect 2988 8335 2990 8340
rect 2993 8338 2995 8340
rect 2951 8321 2953 8324
rect 2956 8321 2958 8323
rect 2972 8321 2974 8328
rect 2988 8321 2990 8331
rect 2993 8321 2995 8328
rect 3009 8321 3011 8340
rect 3025 8331 3027 8340
rect 3030 8338 3032 8340
rect 3051 8338 3053 8340
rect 3067 8337 3069 8340
rect 3025 8321 3027 8324
rect 3030 8321 3032 8323
rect 3051 8321 3053 8323
rect 3067 8321 3069 8333
rect 3083 8331 3085 8340
rect 3088 8338 3090 8340
rect 3104 8332 3106 8340
rect 3120 8335 3122 8340
rect 3125 8338 3127 8340
rect 3083 8321 3085 8324
rect 3088 8321 3090 8323
rect 3104 8321 3106 8328
rect 3120 8321 3122 8331
rect 3125 8321 3127 8328
rect 3141 8321 3143 8340
rect 3157 8331 3159 8340
rect 3162 8338 3164 8340
rect 3183 8338 3185 8340
rect 3199 8337 3201 8340
rect 3157 8321 3159 8324
rect 3162 8321 3164 8323
rect 3183 8321 3185 8323
rect 3199 8321 3201 8333
rect 3215 8331 3217 8340
rect 3220 8338 3222 8340
rect 3236 8332 3238 8340
rect 3252 8335 3254 8340
rect 3257 8338 3259 8340
rect 3215 8321 3217 8324
rect 3220 8321 3222 8323
rect 3236 8321 3238 8328
rect 3252 8321 3254 8331
rect 3257 8321 3259 8328
rect 3273 8321 3275 8340
rect 3289 8331 3291 8340
rect 3294 8338 3296 8340
rect 3315 8338 3317 8340
rect 3331 8337 3333 8340
rect 3289 8321 3291 8324
rect 3294 8321 3296 8323
rect 3315 8321 3317 8323
rect 3331 8321 3333 8333
rect 3347 8331 3349 8340
rect 3352 8338 3354 8340
rect 3368 8332 3370 8340
rect 3801 8335 3803 8340
rect 3806 8338 3808 8340
rect 3347 8321 3349 8324
rect 3352 8321 3354 8323
rect 3368 8321 3370 8328
rect 2504 8315 2506 8317
rect 2509 8315 2511 8318
rect 2525 8315 2527 8317
rect 2541 8315 2543 8317
rect 2546 8315 2548 8318
rect 2567 8315 2569 8318
rect 2583 8315 2585 8318
rect 2599 8315 2601 8317
rect 2604 8315 2606 8318
rect 3801 8321 3803 8331
rect 3806 8321 3808 8328
rect 3822 8321 3824 8340
rect 3838 8331 3840 8340
rect 3843 8338 3845 8340
rect 3864 8338 3866 8340
rect 3880 8337 3882 8340
rect 3838 8321 3840 8324
rect 3843 8321 3845 8323
rect 3864 8321 3866 8323
rect 3880 8321 3882 8333
rect 3896 8331 3898 8340
rect 3901 8338 3903 8340
rect 3917 8332 3919 8340
rect 3933 8335 3935 8340
rect 3938 8338 3940 8340
rect 3896 8321 3898 8324
rect 3901 8321 3903 8323
rect 3917 8321 3919 8328
rect 3933 8321 3935 8331
rect 3938 8321 3940 8328
rect 3954 8321 3956 8340
rect 3970 8331 3972 8340
rect 3975 8338 3977 8340
rect 3996 8338 3998 8340
rect 4012 8337 4014 8340
rect 3970 8321 3972 8324
rect 3975 8321 3977 8323
rect 3996 8321 3998 8323
rect 4012 8321 4014 8333
rect 4028 8331 4030 8340
rect 4033 8338 4035 8340
rect 4049 8332 4051 8340
rect 4065 8335 4067 8340
rect 4070 8338 4072 8340
rect 4028 8321 4030 8324
rect 4033 8321 4035 8323
rect 4049 8321 4051 8328
rect 4065 8321 4067 8331
rect 4070 8321 4072 8328
rect 4086 8321 4088 8340
rect 4102 8331 4104 8340
rect 4107 8338 4109 8340
rect 4128 8338 4130 8340
rect 4144 8337 4146 8340
rect 4102 8321 4104 8324
rect 4107 8321 4109 8323
rect 4128 8321 4130 8323
rect 4144 8321 4146 8333
rect 4160 8331 4162 8340
rect 4165 8338 4167 8340
rect 4181 8332 4183 8340
rect 4197 8335 4199 8340
rect 4202 8338 4204 8340
rect 4160 8321 4162 8324
rect 4165 8321 4167 8323
rect 4181 8321 4183 8328
rect 4197 8321 4199 8331
rect 4202 8321 4204 8328
rect 4218 8321 4220 8340
rect 4234 8331 4236 8340
rect 4239 8338 4241 8340
rect 4260 8338 4262 8340
rect 4276 8337 4278 8340
rect 4234 8321 4236 8324
rect 4239 8321 4241 8323
rect 4260 8321 4262 8323
rect 4276 8321 4278 8333
rect 4292 8331 4294 8340
rect 4297 8338 4299 8340
rect 4313 8332 4315 8340
rect 4292 8321 4294 8324
rect 4297 8321 4299 8323
rect 4313 8321 4315 8328
rect 2620 8315 2622 8317
rect 2856 8315 2858 8317
rect 2861 8314 2863 8317
rect 2877 8315 2879 8317
rect 2893 8315 2895 8317
rect 2898 8312 2900 8317
rect 2919 8312 2921 8317
rect 2935 8315 2937 8317
rect 2951 8315 2953 8317
rect 2956 8312 2958 8317
rect 2972 8315 2974 8317
rect 2988 8315 2990 8317
rect 2993 8314 2995 8317
rect 3009 8315 3011 8317
rect 3025 8315 3027 8317
rect 3030 8312 3032 8317
rect 3051 8312 3053 8317
rect 3067 8315 3069 8317
rect 3083 8315 3085 8317
rect 3088 8312 3090 8317
rect 3104 8315 3106 8317
rect 3120 8315 3122 8317
rect 3125 8314 3127 8317
rect 3141 8315 3143 8317
rect 3157 8315 3159 8317
rect 3162 8312 3164 8317
rect 3183 8312 3185 8317
rect 3199 8315 3201 8317
rect 3215 8315 3217 8317
rect 3220 8312 3222 8317
rect 3236 8315 3238 8317
rect 3252 8315 3254 8317
rect 3257 8314 3259 8317
rect 3273 8315 3275 8317
rect 3289 8315 3291 8317
rect 3294 8312 3296 8317
rect 3315 8312 3317 8317
rect 3331 8315 3333 8317
rect 3347 8315 3349 8317
rect 3352 8312 3354 8317
rect 3368 8315 3370 8317
rect 3449 8315 3451 8317
rect 3454 8315 3456 8318
rect 3470 8315 3472 8317
rect 3486 8315 3488 8317
rect 3491 8315 3493 8318
rect 3512 8315 3514 8318
rect 3528 8315 3530 8318
rect 3544 8315 3546 8317
rect 3549 8315 3551 8318
rect 3565 8315 3567 8317
rect 3801 8315 3803 8317
rect 3806 8314 3808 8317
rect 3822 8315 3824 8317
rect 3838 8315 3840 8317
rect 3843 8312 3845 8317
rect 3864 8312 3866 8317
rect 3880 8315 3882 8317
rect 3896 8315 3898 8317
rect 3901 8312 3903 8317
rect 3917 8315 3919 8317
rect 3933 8315 3935 8317
rect 3938 8314 3940 8317
rect 3954 8315 3956 8317
rect 3970 8315 3972 8317
rect 3975 8312 3977 8317
rect 3996 8312 3998 8317
rect 4012 8315 4014 8317
rect 4028 8315 4030 8317
rect 4033 8312 4035 8317
rect 4049 8315 4051 8317
rect 4065 8315 4067 8317
rect 4070 8314 4072 8317
rect 4086 8315 4088 8317
rect 4102 8315 4104 8317
rect 4107 8312 4109 8317
rect 4128 8312 4130 8317
rect 4144 8315 4146 8317
rect 4160 8315 4162 8317
rect 4165 8312 4167 8317
rect 4181 8315 4183 8317
rect 4197 8315 4199 8317
rect 4202 8314 4204 8317
rect 4218 8315 4220 8317
rect 4234 8315 4236 8317
rect 4239 8312 4241 8317
rect 4260 8312 4262 8317
rect 4276 8315 4278 8317
rect 4292 8315 4294 8317
rect 4297 8312 4299 8317
rect 4313 8315 4315 8317
rect 2504 8302 2506 8307
rect 2509 8305 2511 8307
rect 2504 8288 2506 8298
rect 2509 8288 2511 8295
rect 2525 8288 2527 8307
rect 2541 8298 2543 8307
rect 2546 8305 2548 8307
rect 2567 8305 2569 8307
rect 2583 8304 2585 8307
rect 2541 8288 2543 8291
rect 2546 8288 2548 8290
rect 2567 8288 2569 8290
rect 2583 8288 2585 8300
rect 2599 8298 2601 8307
rect 2604 8305 2606 8307
rect 2599 8288 2601 8291
rect 2604 8288 2606 8290
rect 2620 8288 2622 8307
rect 3449 8302 3451 8307
rect 3454 8305 3456 8307
rect 3449 8288 3451 8298
rect 3454 8288 3456 8295
rect 3470 8288 3472 8307
rect 3486 8298 3488 8307
rect 3491 8305 3493 8307
rect 3512 8305 3514 8307
rect 3528 8304 3530 8307
rect 3486 8288 3488 8291
rect 3491 8288 3493 8290
rect 3512 8288 3514 8290
rect 3528 8288 3530 8300
rect 3544 8298 3546 8307
rect 3549 8305 3551 8307
rect 3544 8288 3546 8291
rect 3549 8288 3551 8290
rect 3565 8288 3567 8307
rect 2504 8282 2506 8284
rect 2509 8281 2511 8284
rect 2525 8282 2527 8284
rect 2541 8282 2543 8284
rect 2546 8279 2548 8284
rect 2567 8279 2569 8284
rect 2583 8282 2585 8284
rect 2599 8282 2601 8284
rect 2604 8279 2606 8284
rect 2620 8282 2622 8284
rect 3449 8282 3451 8284
rect 3454 8281 3456 8284
rect 3470 8282 3472 8284
rect 3486 8282 3488 8284
rect 3035 8277 3037 8279
rect 2877 8271 2879 8274
rect 2921 8271 2923 8274
rect 2947 8271 2949 8274
rect 2993 8271 2995 8274
rect 2947 8267 2948 8271
rect 3061 8271 3063 8275
rect 3089 8277 3091 8279
rect 3116 8277 3118 8279
rect 3066 8271 3068 8274
rect 2861 8264 2863 8266
rect 2877 8264 2879 8267
rect 2893 8264 2895 8266
rect 2916 8264 2918 8266
rect 2921 8264 2923 8267
rect 2947 8264 2949 8267
rect 2968 8264 2970 8267
rect 2988 8264 2990 8266
rect 2993 8264 2995 8267
rect 3011 8264 3013 8266
rect 2628 8251 2630 8254
rect 2628 8245 2630 8247
rect 2511 8242 2513 8245
rect 2861 8242 2863 8256
rect 2877 8254 2879 8256
rect 2877 8242 2879 8244
rect 2893 8242 2895 8256
rect 2916 8251 2918 8256
rect 2921 8254 2923 8256
rect 2947 8254 2949 8256
rect 2912 8247 2918 8251
rect 2916 8242 2918 8247
rect 2921 8242 2923 8244
rect 2947 8242 2949 8244
rect 2968 8242 2970 8256
rect 2988 8251 2990 8256
rect 2993 8254 2995 8256
rect 2984 8247 2990 8251
rect 2988 8242 2990 8247
rect 2993 8242 2995 8244
rect 3011 8242 3013 8256
rect 3035 8255 3037 8269
rect 3142 8271 3144 8275
rect 3170 8277 3172 8279
rect 3491 8279 3493 8284
rect 3512 8279 3514 8284
rect 3528 8282 3530 8284
rect 3544 8282 3546 8284
rect 3549 8279 3551 8284
rect 3565 8282 3567 8284
rect 3147 8271 3149 8274
rect 3061 8260 3063 8263
rect 3066 8261 3068 8263
rect 3062 8256 3063 8260
rect 3061 8251 3063 8256
rect 3066 8251 3068 8253
rect 3035 8249 3037 8251
rect 3089 8247 3091 8269
rect 3116 8255 3118 8269
rect 3980 8277 3982 8279
rect 3142 8260 3144 8263
rect 3147 8261 3149 8263
rect 3143 8256 3144 8260
rect 3142 8251 3144 8256
rect 3147 8251 3149 8253
rect 3116 8249 3118 8251
rect 3170 8247 3172 8269
rect 3822 8271 3824 8274
rect 3866 8271 3868 8274
rect 3892 8271 3894 8274
rect 3938 8271 3940 8274
rect 3892 8267 3893 8271
rect 4006 8271 4008 8275
rect 4034 8277 4036 8279
rect 4061 8277 4063 8279
rect 4011 8271 4013 8274
rect 3806 8264 3808 8266
rect 3822 8264 3824 8267
rect 3838 8264 3840 8266
rect 3861 8264 3863 8266
rect 3866 8264 3868 8267
rect 3892 8264 3894 8267
rect 3913 8264 3915 8267
rect 3933 8264 3935 8266
rect 3938 8264 3940 8267
rect 3956 8264 3958 8266
rect 3573 8251 3575 8254
rect 3061 8245 3063 8247
rect 3066 8242 3068 8247
rect 3142 8245 3144 8247
rect 3089 8241 3091 8243
rect 3147 8242 3149 8247
rect 3573 8245 3575 8247
rect 3170 8241 3172 8243
rect 3456 8242 3458 8245
rect 3806 8242 3808 8256
rect 3822 8254 3824 8256
rect 3822 8242 3824 8244
rect 3838 8242 3840 8256
rect 3861 8251 3863 8256
rect 3866 8254 3868 8256
rect 3892 8254 3894 8256
rect 3857 8247 3863 8251
rect 3861 8242 3863 8247
rect 3866 8242 3868 8244
rect 3892 8242 3894 8244
rect 3913 8242 3915 8256
rect 3933 8251 3935 8256
rect 3938 8254 3940 8256
rect 3929 8247 3935 8251
rect 3933 8242 3935 8247
rect 3938 8242 3940 8244
rect 3956 8242 3958 8256
rect 3980 8255 3982 8269
rect 4087 8271 4089 8275
rect 4115 8277 4117 8279
rect 4092 8271 4094 8274
rect 4006 8260 4008 8263
rect 4011 8261 4013 8263
rect 4007 8256 4008 8260
rect 4006 8251 4008 8256
rect 4011 8251 4013 8253
rect 3980 8249 3982 8251
rect 4034 8247 4036 8269
rect 4061 8255 4063 8269
rect 4087 8260 4089 8263
rect 4092 8261 4094 8263
rect 4088 8256 4089 8260
rect 4087 8251 4089 8256
rect 4092 8251 4094 8253
rect 4061 8249 4063 8251
rect 4115 8247 4117 8269
rect 4006 8245 4008 8247
rect 4011 8242 4013 8247
rect 4087 8245 4089 8247
rect 4034 8241 4036 8243
rect 4092 8242 4094 8247
rect 4115 8241 4117 8243
rect 2511 8236 2513 8238
rect 2861 8236 2863 8238
rect 2877 8234 2879 8238
rect 2893 8236 2895 8238
rect 2916 8236 2918 8238
rect 2878 8230 2879 8234
rect 2921 8233 2923 8238
rect 2947 8234 2949 8238
rect 2968 8236 2970 8238
rect 2988 8236 2990 8238
rect 2877 8227 2879 8230
rect 2922 8229 2923 8233
rect 2948 8230 2949 8234
rect 2993 8233 2995 8238
rect 3011 8236 3013 8238
rect 3456 8236 3458 8238
rect 3806 8236 3808 8238
rect 3822 8234 3824 8238
rect 3838 8236 3840 8238
rect 3861 8236 3863 8238
rect 2921 8227 2923 8229
rect 2947 8226 2949 8230
rect 2994 8229 2995 8233
rect 3823 8230 3824 8234
rect 3866 8233 3868 8238
rect 3892 8234 3894 8238
rect 3913 8236 3915 8238
rect 3933 8236 3935 8238
rect 2993 8227 2995 8229
rect 3822 8227 3824 8230
rect 3867 8229 3868 8233
rect 3893 8230 3894 8234
rect 3938 8233 3940 8238
rect 3956 8236 3958 8238
rect 3866 8227 3868 8229
rect 3892 8226 3894 8230
rect 3939 8229 3940 8233
rect 3938 8227 3940 8229
rect 2495 8213 2497 8215
rect 2511 8213 2513 8216
rect 2516 8213 2518 8215
rect 2532 8213 2534 8216
rect 2548 8213 2550 8216
rect 2569 8213 2571 8216
rect 2574 8213 2576 8215
rect 2590 8213 2592 8215
rect 2606 8213 2608 8216
rect 2611 8213 2613 8215
rect 3440 8213 3442 8215
rect 3456 8213 3458 8216
rect 3461 8213 3463 8215
rect 3477 8213 3479 8216
rect 3493 8213 3495 8216
rect 3514 8213 3516 8216
rect 3519 8213 3521 8215
rect 3535 8213 3537 8215
rect 3551 8213 3553 8216
rect 3556 8213 3558 8215
rect 2495 8186 2497 8205
rect 2511 8203 2513 8205
rect 2516 8196 2518 8205
rect 2532 8202 2534 8205
rect 2548 8203 2550 8205
rect 2569 8203 2571 8205
rect 2511 8186 2513 8188
rect 2516 8186 2518 8189
rect 2532 8186 2534 8198
rect 2574 8196 2576 8205
rect 2548 8186 2550 8188
rect 2569 8186 2571 8188
rect 2574 8186 2576 8189
rect 2590 8186 2592 8205
rect 2606 8203 2608 8205
rect 2611 8200 2613 8205
rect 2877 8204 2879 8207
rect 2921 8205 2923 8207
rect 2878 8200 2879 8204
rect 2922 8201 2923 8205
rect 2947 8204 2949 8208
rect 2993 8205 2995 8207
rect 2861 8196 2863 8198
rect 2877 8196 2879 8200
rect 2893 8196 2895 8198
rect 2916 8196 2918 8198
rect 2921 8196 2923 8201
rect 2948 8200 2949 8204
rect 2994 8201 2995 8205
rect 2947 8196 2949 8200
rect 2968 8196 2970 8198
rect 2988 8196 2990 8198
rect 2993 8196 2995 8201
rect 3011 8196 3013 8198
rect 2606 8186 2608 8193
rect 2611 8186 2613 8196
rect 3061 8195 3063 8198
rect 3066 8195 3068 8198
rect 3142 8195 3144 8198
rect 3147 8195 3149 8198
rect 2495 8180 2497 8182
rect 2511 8177 2513 8182
rect 2516 8180 2518 8182
rect 2532 8180 2534 8182
rect 2548 8177 2550 8182
rect 2569 8177 2571 8182
rect 2574 8180 2576 8182
rect 2590 8180 2592 8182
rect 2606 8179 2608 8182
rect 2611 8180 2613 8182
rect 2861 8178 2863 8192
rect 2877 8190 2879 8192
rect 2877 8178 2879 8180
rect 2893 8178 2895 8192
rect 2916 8187 2918 8192
rect 2921 8190 2923 8192
rect 2947 8190 2949 8192
rect 2912 8183 2918 8187
rect 2916 8178 2918 8183
rect 2921 8178 2923 8180
rect 2947 8178 2949 8180
rect 2968 8178 2970 8192
rect 2988 8187 2990 8192
rect 2993 8190 2995 8192
rect 2984 8183 2990 8187
rect 2988 8178 2990 8183
rect 2993 8178 2995 8180
rect 3011 8178 3013 8192
rect 3061 8179 3063 8191
rect 3066 8189 3068 8191
rect 3066 8179 3068 8181
rect 3142 8179 3144 8191
rect 3147 8189 3149 8191
rect 3440 8186 3442 8205
rect 3456 8203 3458 8205
rect 3461 8196 3463 8205
rect 3477 8202 3479 8205
rect 3493 8203 3495 8205
rect 3514 8203 3516 8205
rect 3456 8186 3458 8188
rect 3461 8186 3463 8189
rect 3477 8186 3479 8198
rect 3519 8196 3521 8205
rect 3493 8186 3495 8188
rect 3514 8186 3516 8188
rect 3519 8186 3521 8189
rect 3535 8186 3537 8205
rect 3551 8203 3553 8205
rect 3556 8200 3558 8205
rect 3822 8204 3824 8207
rect 3866 8205 3868 8207
rect 3823 8200 3824 8204
rect 3867 8201 3868 8205
rect 3892 8204 3894 8208
rect 3938 8205 3940 8207
rect 3806 8196 3808 8198
rect 3822 8196 3824 8200
rect 3838 8196 3840 8198
rect 3861 8196 3863 8198
rect 3866 8196 3868 8201
rect 3893 8200 3894 8204
rect 3939 8201 3940 8205
rect 3892 8196 3894 8200
rect 3913 8196 3915 8198
rect 3933 8196 3935 8198
rect 3938 8196 3940 8201
rect 3956 8196 3958 8198
rect 3551 8186 3553 8193
rect 3556 8186 3558 8196
rect 4006 8195 4008 8198
rect 4011 8195 4013 8198
rect 4087 8195 4089 8198
rect 4092 8195 4094 8198
rect 3147 8179 3149 8181
rect 3440 8180 3442 8182
rect 3456 8177 3458 8182
rect 3461 8180 3463 8182
rect 3477 8180 3479 8182
rect 3493 8177 3495 8182
rect 3514 8177 3516 8182
rect 3519 8180 3521 8182
rect 3535 8180 3537 8182
rect 3551 8179 3553 8182
rect 3556 8180 3558 8182
rect 3806 8178 3808 8192
rect 3822 8190 3824 8192
rect 3822 8178 3824 8180
rect 3838 8178 3840 8192
rect 3861 8187 3863 8192
rect 3866 8190 3868 8192
rect 3892 8190 3894 8192
rect 3857 8183 3863 8187
rect 3861 8178 3863 8183
rect 3866 8178 3868 8180
rect 3892 8178 3894 8180
rect 3913 8178 3915 8192
rect 3933 8187 3935 8192
rect 3938 8190 3940 8192
rect 3929 8183 3935 8187
rect 3933 8178 3935 8183
rect 3938 8178 3940 8180
rect 3956 8178 3958 8192
rect 4006 8179 4008 8191
rect 4011 8189 4013 8191
rect 4011 8179 4013 8181
rect 4087 8179 4089 8191
rect 4092 8189 4094 8191
rect 4092 8179 4094 8181
rect 2861 8168 2863 8170
rect 2877 8167 2879 8170
rect 2893 8168 2895 8170
rect 2916 8168 2918 8170
rect 2921 8167 2923 8170
rect 2947 8167 2949 8170
rect 2968 8167 2970 8170
rect 2988 8168 2990 8170
rect 2993 8167 2995 8170
rect 3011 8168 3013 8170
rect 3061 8169 3063 8171
rect 2947 8163 2948 8167
rect 3066 8166 3068 8171
rect 3142 8169 3144 8171
rect 3147 8166 3149 8171
rect 3806 8168 3808 8170
rect 3822 8167 3824 8170
rect 3838 8168 3840 8170
rect 3861 8168 3863 8170
rect 3866 8167 3868 8170
rect 3892 8167 3894 8170
rect 3913 8167 3915 8170
rect 3933 8168 3935 8170
rect 3938 8167 3940 8170
rect 3956 8168 3958 8170
rect 4006 8169 4008 8171
rect 2877 8160 2879 8163
rect 2921 8160 2923 8163
rect 2947 8160 2949 8163
rect 2993 8160 2995 8163
rect 3892 8163 3893 8167
rect 4011 8166 4013 8171
rect 4087 8169 4089 8171
rect 4092 8166 4094 8171
rect 3822 8160 3824 8163
rect 3866 8160 3868 8163
rect 3892 8160 3894 8163
rect 3938 8160 3940 8163
rect 2877 8139 2879 8142
rect 2921 8139 2923 8142
rect 2947 8139 2949 8142
rect 2993 8139 2995 8142
rect 3061 8139 3063 8143
rect 3089 8145 3091 8147
rect 3140 8145 3142 8147
rect 3066 8139 3068 8142
rect 2947 8135 2948 8139
rect 2861 8132 2863 8134
rect 2877 8132 2879 8135
rect 2893 8132 2895 8134
rect 2916 8132 2918 8134
rect 2921 8132 2923 8135
rect 2947 8132 2949 8135
rect 2968 8132 2970 8135
rect 2988 8132 2990 8134
rect 2993 8132 2995 8135
rect 3011 8132 3013 8134
rect 3166 8139 3168 8143
rect 3194 8145 3196 8147
rect 3171 8139 3173 8142
rect 3061 8128 3063 8131
rect 3066 8129 3068 8131
rect 3062 8124 3063 8128
rect 2861 8110 2863 8124
rect 2877 8122 2879 8124
rect 2877 8110 2879 8112
rect 2893 8110 2895 8124
rect 2916 8119 2918 8124
rect 2921 8122 2923 8124
rect 2947 8122 2949 8124
rect 2912 8115 2918 8119
rect 2916 8110 2918 8115
rect 2921 8110 2923 8112
rect 2947 8110 2949 8112
rect 2968 8110 2970 8124
rect 2988 8119 2990 8124
rect 2993 8122 2995 8124
rect 2984 8115 2990 8119
rect 2988 8110 2990 8115
rect 2993 8110 2995 8112
rect 3011 8110 3013 8124
rect 3061 8119 3063 8124
rect 3066 8119 3068 8121
rect 3089 8115 3091 8137
rect 3140 8123 3142 8137
rect 3822 8139 3824 8142
rect 3866 8139 3868 8142
rect 3892 8139 3894 8142
rect 3938 8139 3940 8142
rect 4006 8139 4008 8143
rect 4034 8145 4036 8147
rect 4085 8145 4087 8147
rect 4011 8139 4013 8142
rect 3166 8128 3168 8131
rect 3171 8129 3173 8131
rect 3167 8124 3168 8128
rect 3166 8119 3168 8124
rect 3171 8119 3173 8121
rect 3140 8117 3142 8119
rect 3194 8115 3196 8137
rect 3892 8135 3893 8139
rect 3806 8132 3808 8134
rect 3822 8132 3824 8135
rect 3838 8132 3840 8134
rect 3861 8132 3863 8134
rect 3866 8132 3868 8135
rect 3892 8132 3894 8135
rect 3913 8132 3915 8135
rect 3933 8132 3935 8134
rect 3938 8132 3940 8135
rect 3956 8132 3958 8134
rect 4111 8139 4113 8143
rect 4139 8145 4141 8147
rect 4116 8139 4118 8142
rect 4006 8128 4008 8131
rect 4011 8129 4013 8131
rect 4007 8124 4008 8128
rect 3061 8113 3063 8115
rect 3066 8110 3068 8115
rect 3166 8113 3168 8115
rect 3089 8109 3091 8111
rect 3171 8110 3173 8115
rect 3194 8109 3196 8111
rect 3806 8110 3808 8124
rect 3822 8122 3824 8124
rect 3822 8110 3824 8112
rect 3838 8110 3840 8124
rect 3861 8119 3863 8124
rect 3866 8122 3868 8124
rect 3892 8122 3894 8124
rect 3857 8115 3863 8119
rect 3861 8110 3863 8115
rect 3866 8110 3868 8112
rect 3892 8110 3894 8112
rect 3913 8110 3915 8124
rect 3933 8119 3935 8124
rect 3938 8122 3940 8124
rect 3929 8115 3935 8119
rect 3933 8110 3935 8115
rect 3938 8110 3940 8112
rect 3956 8110 3958 8124
rect 4006 8119 4008 8124
rect 4011 8119 4013 8121
rect 4034 8115 4036 8137
rect 4085 8123 4087 8137
rect 4111 8128 4113 8131
rect 4116 8129 4118 8131
rect 4112 8124 4113 8128
rect 4111 8119 4113 8124
rect 4116 8119 4118 8121
rect 4085 8117 4087 8119
rect 4139 8115 4141 8137
rect 4006 8113 4008 8115
rect 4011 8110 4013 8115
rect 4111 8113 4113 8115
rect 4034 8109 4036 8111
rect 4116 8110 4118 8115
rect 4139 8109 4141 8111
rect 2861 8104 2863 8106
rect 2877 8102 2879 8106
rect 2893 8104 2895 8106
rect 2916 8104 2918 8106
rect 2878 8098 2879 8102
rect 2921 8101 2923 8106
rect 2947 8102 2949 8106
rect 2968 8104 2970 8106
rect 2988 8104 2990 8106
rect 2877 8095 2879 8098
rect 2922 8097 2923 8101
rect 2948 8098 2949 8102
rect 2993 8101 2995 8106
rect 3011 8104 3013 8106
rect 3806 8104 3808 8106
rect 3822 8102 3824 8106
rect 3838 8104 3840 8106
rect 3861 8104 3863 8106
rect 2921 8095 2923 8097
rect 2947 8094 2949 8098
rect 2994 8097 2995 8101
rect 3823 8098 3824 8102
rect 3866 8101 3868 8106
rect 3892 8102 3894 8106
rect 3913 8104 3915 8106
rect 3933 8104 3935 8106
rect 2993 8095 2995 8097
rect 3822 8095 3824 8098
rect 3867 8097 3868 8101
rect 3893 8098 3894 8102
rect 3938 8101 3940 8106
rect 3956 8104 3958 8106
rect 3866 8095 3868 8097
rect 3892 8094 3894 8098
rect 3939 8097 3940 8101
rect 3938 8095 3940 8097
rect 2877 8072 2879 8075
rect 2921 8073 2923 8075
rect 2878 8068 2879 8072
rect 2922 8069 2923 8073
rect 2947 8072 2949 8076
rect 2993 8073 2995 8075
rect 2861 8064 2863 8066
rect 2877 8064 2879 8068
rect 2893 8064 2895 8066
rect 2916 8064 2918 8066
rect 2921 8064 2923 8069
rect 2948 8068 2949 8072
rect 2994 8069 2995 8073
rect 3822 8072 3824 8075
rect 3866 8073 3868 8075
rect 2947 8064 2949 8068
rect 2968 8064 2970 8066
rect 2988 8064 2990 8066
rect 2993 8064 2995 8069
rect 3823 8068 3824 8072
rect 3867 8069 3868 8073
rect 3892 8072 3894 8076
rect 3938 8073 3940 8075
rect 3011 8064 3013 8066
rect 3061 8064 3063 8067
rect 3066 8064 3068 8067
rect 3166 8064 3168 8067
rect 3171 8064 3173 8067
rect 3806 8064 3808 8066
rect 3822 8064 3824 8068
rect 3838 8064 3840 8066
rect 3861 8064 3863 8066
rect 3866 8064 3868 8069
rect 3893 8068 3894 8072
rect 3939 8069 3940 8073
rect 3892 8064 3894 8068
rect 3913 8064 3915 8066
rect 3933 8064 3935 8066
rect 3938 8064 3940 8069
rect 3956 8064 3958 8066
rect 4006 8064 4008 8067
rect 4011 8064 4013 8067
rect 4111 8064 4113 8067
rect 4116 8064 4118 8067
rect 2861 8046 2863 8060
rect 2877 8058 2879 8060
rect 2877 8046 2879 8048
rect 2893 8046 2895 8060
rect 2916 8055 2918 8060
rect 2921 8058 2923 8060
rect 2947 8058 2949 8060
rect 2912 8051 2918 8055
rect 2916 8046 2918 8051
rect 2921 8046 2923 8048
rect 2947 8046 2949 8048
rect 2968 8046 2970 8060
rect 2988 8055 2990 8060
rect 2993 8058 2995 8060
rect 2984 8051 2990 8055
rect 2988 8046 2990 8051
rect 2993 8046 2995 8048
rect 3011 8046 3013 8060
rect 3061 8048 3063 8060
rect 3066 8058 3068 8060
rect 3066 8048 3068 8050
rect 3166 8048 3168 8060
rect 3171 8058 3173 8060
rect 3171 8048 3173 8050
rect 3806 8046 3808 8060
rect 3822 8058 3824 8060
rect 3822 8046 3824 8048
rect 3838 8046 3840 8060
rect 3861 8055 3863 8060
rect 3866 8058 3868 8060
rect 3892 8058 3894 8060
rect 3857 8051 3863 8055
rect 3861 8046 3863 8051
rect 3866 8046 3868 8048
rect 3892 8046 3894 8048
rect 3913 8046 3915 8060
rect 3933 8055 3935 8060
rect 3938 8058 3940 8060
rect 3929 8051 3935 8055
rect 3933 8046 3935 8051
rect 3938 8046 3940 8048
rect 3956 8046 3958 8060
rect 4006 8048 4008 8060
rect 4011 8058 4013 8060
rect 4011 8048 4013 8050
rect 4111 8048 4113 8060
rect 4116 8058 4118 8060
rect 4116 8048 4118 8050
rect 3061 8038 3063 8040
rect 2861 8036 2863 8038
rect 2877 8035 2879 8038
rect 2893 8036 2895 8038
rect 2916 8036 2918 8038
rect 2921 8035 2923 8038
rect 2947 8035 2949 8038
rect 2968 8035 2970 8038
rect 2988 8036 2990 8038
rect 2993 8035 2995 8038
rect 3011 8036 3013 8038
rect 3066 8035 3068 8040
rect 3166 8038 3168 8040
rect 3171 8035 3173 8040
rect 4006 8038 4008 8040
rect 3806 8036 3808 8038
rect 2947 8031 2948 8035
rect 3822 8035 3824 8038
rect 3838 8036 3840 8038
rect 3861 8036 3863 8038
rect 3866 8035 3868 8038
rect 3892 8035 3894 8038
rect 3913 8035 3915 8038
rect 3933 8036 3935 8038
rect 3938 8035 3940 8038
rect 3956 8036 3958 8038
rect 4011 8035 4013 8040
rect 4111 8038 4113 8040
rect 4116 8035 4118 8040
rect 3892 8031 3893 8035
rect 2877 8028 2879 8031
rect 2921 8028 2923 8031
rect 2947 8028 2949 8031
rect 2993 8028 2995 8031
rect 3822 8028 3824 8031
rect 3866 8028 3868 8031
rect 3892 8028 3894 8031
rect 3938 8028 3940 8031
rect 2877 8007 2879 8010
rect 2921 8007 2923 8010
rect 2947 8007 2949 8010
rect 2993 8007 2995 8010
rect 3061 8007 3063 8011
rect 3089 8013 3091 8015
rect 3116 8013 3118 8015
rect 3066 8007 3068 8010
rect 2947 8003 2948 8007
rect 2861 8000 2863 8002
rect 2877 8000 2879 8003
rect 2893 8000 2895 8002
rect 2916 8000 2918 8002
rect 2921 8000 2923 8003
rect 2947 8000 2949 8003
rect 2968 8000 2970 8003
rect 2988 8000 2990 8002
rect 2993 8000 2995 8003
rect 3011 8000 3013 8002
rect 3142 8007 3144 8011
rect 3170 8013 3172 8015
rect 3206 8013 3208 8015
rect 3147 8007 3149 8010
rect 3061 7996 3063 7999
rect 3066 7997 3068 7999
rect 3062 7992 3063 7996
rect 2861 7978 2863 7992
rect 2877 7990 2879 7992
rect 2877 7978 2879 7980
rect 2893 7978 2895 7992
rect 2916 7987 2918 7992
rect 2921 7990 2923 7992
rect 2947 7990 2949 7992
rect 2912 7983 2918 7987
rect 2916 7978 2918 7983
rect 2921 7978 2923 7980
rect 2947 7978 2949 7980
rect 2968 7978 2970 7992
rect 2988 7987 2990 7992
rect 2993 7990 2995 7992
rect 2984 7983 2990 7987
rect 2988 7978 2990 7983
rect 2993 7978 2995 7980
rect 3011 7978 3013 7992
rect 3061 7987 3063 7992
rect 3066 7987 3068 7989
rect 3089 7983 3091 8005
rect 3116 7991 3118 8005
rect 3232 8007 3234 8011
rect 3260 8013 3262 8015
rect 3237 8007 3239 8010
rect 3142 7996 3144 7999
rect 3147 7997 3149 7999
rect 3143 7992 3144 7996
rect 3142 7987 3144 7992
rect 3147 7987 3149 7989
rect 3116 7985 3118 7987
rect 3170 7983 3172 8005
rect 3206 7991 3208 8005
rect 3822 8007 3824 8010
rect 3866 8007 3868 8010
rect 3892 8007 3894 8010
rect 3938 8007 3940 8010
rect 4006 8007 4008 8011
rect 4034 8013 4036 8015
rect 4061 8013 4063 8015
rect 4011 8007 4013 8010
rect 3232 7996 3234 7999
rect 3237 7997 3239 7999
rect 3233 7992 3234 7996
rect 3232 7987 3234 7992
rect 3237 7987 3239 7989
rect 3206 7985 3208 7987
rect 3260 7983 3262 8005
rect 3892 8003 3893 8007
rect 3806 8000 3808 8002
rect 3822 8000 3824 8003
rect 3838 8000 3840 8002
rect 3861 8000 3863 8002
rect 3866 8000 3868 8003
rect 3892 8000 3894 8003
rect 3913 8000 3915 8003
rect 3933 8000 3935 8002
rect 3938 8000 3940 8003
rect 3956 8000 3958 8002
rect 4087 8007 4089 8011
rect 4115 8013 4117 8015
rect 4151 8013 4153 8015
rect 4092 8007 4094 8010
rect 4006 7996 4008 7999
rect 4011 7997 4013 7999
rect 4007 7992 4008 7996
rect 3061 7981 3063 7983
rect 3066 7978 3068 7983
rect 3142 7981 3144 7983
rect 3089 7977 3091 7979
rect 3147 7978 3149 7983
rect 3232 7981 3234 7983
rect 3170 7977 3172 7979
rect 3237 7978 3239 7983
rect 3260 7977 3262 7979
rect 3806 7978 3808 7992
rect 3822 7990 3824 7992
rect 3822 7978 3824 7980
rect 3838 7978 3840 7992
rect 3861 7987 3863 7992
rect 3866 7990 3868 7992
rect 3892 7990 3894 7992
rect 3857 7983 3863 7987
rect 3861 7978 3863 7983
rect 3866 7978 3868 7980
rect 3892 7978 3894 7980
rect 3913 7978 3915 7992
rect 3933 7987 3935 7992
rect 3938 7990 3940 7992
rect 3929 7983 3935 7987
rect 3933 7978 3935 7983
rect 3938 7978 3940 7980
rect 3956 7978 3958 7992
rect 4006 7987 4008 7992
rect 4011 7987 4013 7989
rect 4034 7983 4036 8005
rect 4061 7991 4063 8005
rect 4177 8007 4179 8011
rect 4205 8013 4207 8015
rect 4182 8007 4184 8010
rect 4087 7996 4089 7999
rect 4092 7997 4094 7999
rect 4088 7992 4089 7996
rect 4087 7987 4089 7992
rect 4092 7987 4094 7989
rect 4061 7985 4063 7987
rect 4115 7983 4117 8005
rect 4151 7991 4153 8005
rect 4177 7996 4179 7999
rect 4182 7997 4184 7999
rect 4178 7992 4179 7996
rect 4177 7987 4179 7992
rect 4182 7987 4184 7989
rect 4151 7985 4153 7987
rect 4205 7983 4207 8005
rect 4006 7981 4008 7983
rect 4011 7978 4013 7983
rect 4087 7981 4089 7983
rect 4034 7977 4036 7979
rect 4092 7978 4094 7983
rect 4177 7981 4179 7983
rect 4115 7977 4117 7979
rect 4182 7978 4184 7983
rect 4205 7977 4207 7979
rect 2861 7972 2863 7974
rect 2877 7970 2879 7974
rect 2893 7972 2895 7974
rect 2916 7972 2918 7974
rect 2878 7966 2879 7970
rect 2921 7969 2923 7974
rect 2947 7970 2949 7974
rect 2968 7972 2970 7974
rect 2988 7972 2990 7974
rect 2877 7963 2879 7966
rect 2922 7965 2923 7969
rect 2948 7966 2949 7970
rect 2993 7969 2995 7974
rect 3011 7972 3013 7974
rect 3806 7972 3808 7974
rect 3822 7970 3824 7974
rect 3838 7972 3840 7974
rect 3861 7972 3863 7974
rect 2921 7963 2923 7965
rect 2947 7962 2949 7966
rect 2994 7965 2995 7969
rect 3823 7966 3824 7970
rect 3866 7969 3868 7974
rect 3892 7970 3894 7974
rect 3913 7972 3915 7974
rect 3933 7972 3935 7974
rect 2993 7963 2995 7965
rect 3822 7963 3824 7966
rect 3867 7965 3868 7969
rect 3893 7966 3894 7970
rect 3938 7969 3940 7974
rect 3956 7972 3958 7974
rect 3866 7963 3868 7965
rect 3892 7962 3894 7966
rect 3939 7965 3940 7969
rect 3938 7963 3940 7965
rect 2877 7940 2879 7943
rect 2921 7941 2923 7943
rect 2878 7936 2879 7940
rect 2922 7937 2923 7941
rect 2947 7940 2949 7944
rect 2993 7941 2995 7943
rect 2861 7932 2863 7934
rect 2877 7932 2879 7936
rect 2893 7932 2895 7934
rect 2916 7932 2918 7934
rect 2921 7932 2923 7937
rect 2948 7936 2949 7940
rect 2994 7937 2995 7941
rect 3822 7940 3824 7943
rect 3866 7941 3868 7943
rect 2947 7932 2949 7936
rect 2968 7932 2970 7934
rect 2988 7932 2990 7934
rect 2993 7932 2995 7937
rect 3823 7936 3824 7940
rect 3867 7937 3868 7941
rect 3892 7940 3894 7944
rect 3938 7941 3940 7943
rect 3011 7932 3013 7934
rect 3806 7932 3808 7934
rect 3822 7932 3824 7936
rect 3838 7932 3840 7934
rect 3861 7932 3863 7934
rect 3866 7932 3868 7937
rect 3893 7936 3894 7940
rect 3939 7937 3940 7941
rect 3892 7932 3894 7936
rect 3913 7932 3915 7934
rect 3933 7932 3935 7934
rect 3938 7932 3940 7937
rect 3956 7932 3958 7934
rect 3061 7929 3063 7932
rect 3066 7929 3068 7932
rect 3142 7929 3144 7932
rect 3147 7929 3149 7932
rect 3232 7929 3234 7932
rect 3237 7929 3239 7932
rect 2861 7914 2863 7928
rect 2877 7926 2879 7928
rect 2877 7914 2879 7916
rect 2893 7914 2895 7928
rect 2916 7923 2918 7928
rect 2921 7926 2923 7928
rect 2947 7926 2949 7928
rect 2912 7919 2918 7923
rect 2916 7914 2918 7919
rect 2921 7914 2923 7916
rect 2947 7914 2949 7916
rect 2968 7914 2970 7928
rect 2988 7923 2990 7928
rect 2993 7926 2995 7928
rect 2984 7919 2990 7923
rect 2988 7914 2990 7919
rect 2993 7914 2995 7916
rect 3011 7914 3013 7928
rect 4006 7929 4008 7932
rect 4011 7929 4013 7932
rect 4087 7929 4089 7932
rect 4092 7929 4094 7932
rect 4177 7929 4179 7932
rect 4182 7929 4184 7932
rect 3061 7913 3063 7925
rect 3066 7923 3068 7925
rect 3066 7913 3068 7915
rect 3142 7913 3144 7925
rect 3147 7923 3149 7925
rect 3147 7913 3149 7915
rect 3232 7913 3234 7925
rect 3237 7923 3239 7925
rect 3237 7913 3239 7915
rect 3806 7914 3808 7928
rect 3822 7926 3824 7928
rect 3822 7914 3824 7916
rect 3838 7914 3840 7928
rect 3861 7923 3863 7928
rect 3866 7926 3868 7928
rect 3892 7926 3894 7928
rect 3857 7919 3863 7923
rect 3861 7914 3863 7919
rect 3866 7914 3868 7916
rect 3892 7914 3894 7916
rect 3913 7914 3915 7928
rect 3933 7923 3935 7928
rect 3938 7926 3940 7928
rect 3929 7919 3935 7923
rect 3933 7914 3935 7919
rect 3938 7914 3940 7916
rect 3956 7914 3958 7928
rect 2861 7904 2863 7906
rect 2877 7903 2879 7906
rect 2893 7904 2895 7906
rect 2916 7904 2918 7906
rect 2921 7903 2923 7906
rect 2947 7903 2949 7906
rect 2968 7903 2970 7906
rect 2988 7904 2990 7906
rect 2993 7903 2995 7906
rect 3011 7904 3013 7906
rect 4006 7913 4008 7925
rect 4011 7923 4013 7925
rect 4011 7913 4013 7915
rect 4087 7913 4089 7925
rect 4092 7923 4094 7925
rect 4092 7913 4094 7915
rect 4177 7913 4179 7925
rect 4182 7923 4184 7925
rect 4182 7913 4184 7915
rect 3061 7903 3063 7905
rect 2947 7899 2948 7903
rect 3066 7900 3068 7905
rect 3142 7903 3144 7905
rect 3147 7900 3149 7905
rect 3232 7903 3234 7905
rect 3237 7900 3239 7905
rect 3806 7904 3808 7906
rect 2877 7896 2879 7899
rect 2921 7896 2923 7899
rect 2947 7896 2949 7899
rect 2993 7896 2995 7899
rect 3822 7903 3824 7906
rect 3838 7904 3840 7906
rect 3861 7904 3863 7906
rect 3866 7903 3868 7906
rect 3892 7903 3894 7906
rect 3913 7903 3915 7906
rect 3933 7904 3935 7906
rect 3938 7903 3940 7906
rect 3956 7904 3958 7906
rect 4006 7903 4008 7905
rect 3892 7899 3893 7903
rect 4011 7900 4013 7905
rect 4087 7903 4089 7905
rect 4092 7900 4094 7905
rect 4177 7903 4179 7905
rect 4182 7900 4184 7905
rect 3822 7896 3824 7899
rect 3866 7896 3868 7899
rect 3892 7896 3894 7899
rect 3938 7896 3940 7899
rect 2877 7875 2879 7878
rect 2921 7875 2923 7878
rect 2947 7875 2949 7878
rect 2993 7875 2995 7878
rect 3061 7875 3063 7879
rect 3089 7881 3091 7883
rect 3066 7875 3068 7878
rect 2947 7871 2948 7875
rect 2861 7868 2863 7870
rect 2877 7868 2879 7871
rect 2893 7868 2895 7870
rect 2916 7868 2918 7870
rect 2921 7868 2923 7871
rect 2947 7868 2949 7871
rect 2968 7868 2970 7871
rect 2988 7868 2990 7870
rect 2993 7868 2995 7871
rect 3011 7868 3013 7870
rect 3822 7875 3824 7878
rect 3866 7875 3868 7878
rect 3892 7875 3894 7878
rect 3938 7875 3940 7878
rect 4006 7875 4008 7879
rect 4034 7881 4036 7883
rect 4011 7875 4013 7878
rect 3061 7864 3063 7867
rect 3066 7865 3068 7867
rect 3062 7860 3063 7864
rect 2861 7846 2863 7860
rect 2877 7858 2879 7860
rect 2877 7846 2879 7848
rect 2893 7846 2895 7860
rect 2916 7855 2918 7860
rect 2921 7858 2923 7860
rect 2947 7858 2949 7860
rect 2912 7851 2918 7855
rect 2916 7846 2918 7851
rect 2921 7846 2923 7848
rect 2947 7846 2949 7848
rect 2968 7846 2970 7860
rect 2988 7855 2990 7860
rect 2993 7858 2995 7860
rect 2984 7851 2990 7855
rect 2988 7846 2990 7851
rect 2993 7846 2995 7848
rect 3011 7846 3013 7860
rect 3061 7855 3063 7860
rect 3066 7855 3068 7857
rect 3089 7851 3091 7873
rect 3892 7871 3893 7875
rect 3806 7868 3808 7870
rect 3822 7868 3824 7871
rect 3838 7868 3840 7870
rect 3861 7868 3863 7870
rect 3866 7868 3868 7871
rect 3892 7868 3894 7871
rect 3913 7868 3915 7871
rect 3933 7868 3935 7870
rect 3938 7868 3940 7871
rect 3956 7868 3958 7870
rect 4006 7864 4008 7867
rect 4011 7865 4013 7867
rect 4007 7860 4008 7864
rect 3061 7849 3063 7851
rect 3066 7846 3068 7851
rect 3089 7845 3091 7847
rect 3806 7846 3808 7860
rect 3822 7858 3824 7860
rect 3822 7846 3824 7848
rect 3838 7846 3840 7860
rect 3861 7855 3863 7860
rect 3866 7858 3868 7860
rect 3892 7858 3894 7860
rect 3857 7851 3863 7855
rect 3861 7846 3863 7851
rect 3866 7846 3868 7848
rect 3892 7846 3894 7848
rect 3913 7846 3915 7860
rect 3933 7855 3935 7860
rect 3938 7858 3940 7860
rect 3929 7851 3935 7855
rect 3933 7846 3935 7851
rect 3938 7846 3940 7848
rect 3956 7846 3958 7860
rect 4006 7855 4008 7860
rect 4011 7855 4013 7857
rect 4034 7851 4036 7873
rect 4006 7849 4008 7851
rect 4011 7846 4013 7851
rect 4034 7845 4036 7847
rect 2861 7840 2863 7842
rect 2877 7838 2879 7842
rect 2893 7840 2895 7842
rect 2916 7840 2918 7842
rect 2878 7834 2879 7838
rect 2921 7837 2923 7842
rect 2947 7838 2949 7842
rect 2968 7840 2970 7842
rect 2988 7840 2990 7842
rect 2877 7831 2879 7834
rect 2922 7833 2923 7837
rect 2948 7834 2949 7838
rect 2993 7837 2995 7842
rect 3011 7840 3013 7842
rect 3806 7840 3808 7842
rect 3822 7838 3824 7842
rect 3838 7840 3840 7842
rect 3861 7840 3863 7842
rect 2921 7831 2923 7833
rect 2947 7830 2949 7834
rect 2994 7833 2995 7837
rect 3823 7834 3824 7838
rect 3866 7837 3868 7842
rect 3892 7838 3894 7842
rect 3913 7840 3915 7842
rect 3933 7840 3935 7842
rect 2993 7831 2995 7833
rect 3822 7831 3824 7834
rect 3867 7833 3868 7837
rect 3893 7834 3894 7838
rect 3938 7837 3940 7842
rect 3956 7840 3958 7842
rect 3866 7831 3868 7833
rect 3892 7830 3894 7834
rect 3939 7833 3940 7837
rect 3938 7831 3940 7833
rect 2372 7813 2374 7815
rect 2377 7813 2379 7816
rect 2393 7813 2395 7815
rect 2409 7813 2411 7815
rect 2414 7813 2416 7816
rect 2435 7813 2437 7816
rect 2451 7813 2453 7816
rect 2467 7813 2469 7815
rect 2472 7813 2474 7816
rect 2488 7813 2490 7815
rect 2504 7813 2506 7815
rect 2509 7813 2511 7816
rect 2525 7813 2527 7815
rect 2541 7813 2543 7815
rect 2546 7813 2548 7816
rect 2567 7813 2569 7816
rect 2583 7813 2585 7816
rect 2599 7813 2601 7815
rect 2604 7813 2606 7816
rect 2620 7813 2622 7815
rect 2636 7813 2638 7815
rect 2641 7813 2643 7816
rect 2657 7813 2659 7815
rect 2673 7813 2675 7815
rect 2678 7813 2680 7816
rect 2699 7813 2701 7816
rect 2715 7813 2717 7816
rect 2731 7813 2733 7815
rect 2736 7813 2738 7816
rect 2752 7813 2754 7815
rect 3317 7813 3319 7815
rect 3322 7813 3324 7816
rect 3338 7813 3340 7815
rect 3354 7813 3356 7815
rect 3359 7813 3361 7816
rect 3380 7813 3382 7816
rect 3396 7813 3398 7816
rect 3412 7813 3414 7815
rect 3417 7813 3419 7816
rect 3433 7813 3435 7815
rect 3449 7813 3451 7815
rect 3454 7813 3456 7816
rect 3470 7813 3472 7815
rect 3486 7813 3488 7815
rect 3491 7813 3493 7816
rect 3512 7813 3514 7816
rect 3528 7813 3530 7816
rect 3544 7813 3546 7815
rect 3549 7813 3551 7816
rect 3565 7813 3567 7815
rect 3581 7813 3583 7815
rect 3586 7813 3588 7816
rect 3602 7813 3604 7815
rect 3618 7813 3620 7815
rect 3623 7813 3625 7816
rect 3644 7813 3646 7816
rect 3660 7813 3662 7816
rect 3676 7813 3678 7815
rect 3681 7813 3683 7816
rect 3697 7813 3699 7815
rect 2877 7808 2879 7811
rect 2921 7809 2923 7811
rect 2372 7800 2374 7805
rect 2377 7803 2379 7805
rect 2372 7786 2374 7796
rect 2377 7786 2379 7793
rect 2393 7786 2395 7805
rect 2409 7796 2411 7805
rect 2414 7803 2416 7805
rect 2435 7803 2437 7805
rect 2451 7802 2453 7805
rect 2409 7786 2411 7789
rect 2414 7786 2416 7788
rect 2435 7786 2437 7788
rect 2451 7786 2453 7798
rect 2467 7796 2469 7805
rect 2472 7803 2474 7805
rect 2467 7786 2469 7789
rect 2472 7786 2474 7788
rect 2488 7786 2490 7805
rect 2504 7802 2506 7805
rect 2509 7803 2511 7805
rect 2504 7786 2506 7798
rect 2509 7786 2511 7793
rect 2525 7786 2527 7805
rect 2541 7796 2543 7805
rect 2546 7803 2548 7805
rect 2567 7803 2569 7805
rect 2583 7802 2585 7805
rect 2541 7786 2543 7789
rect 2546 7786 2548 7788
rect 2567 7786 2569 7788
rect 2583 7786 2585 7798
rect 2599 7796 2601 7805
rect 2604 7803 2606 7805
rect 2599 7786 2601 7789
rect 2604 7786 2606 7788
rect 2620 7786 2622 7805
rect 2636 7802 2638 7805
rect 2641 7803 2643 7805
rect 2636 7786 2638 7798
rect 2641 7786 2643 7793
rect 2657 7786 2659 7805
rect 2673 7796 2675 7805
rect 2678 7803 2680 7805
rect 2699 7803 2701 7805
rect 2715 7802 2717 7805
rect 2673 7786 2675 7789
rect 2678 7786 2680 7788
rect 2699 7786 2701 7788
rect 2715 7786 2717 7798
rect 2731 7796 2733 7805
rect 2736 7803 2738 7805
rect 2752 7797 2754 7805
rect 2878 7804 2879 7808
rect 2922 7805 2923 7809
rect 2947 7808 2949 7812
rect 2993 7809 2995 7811
rect 2861 7800 2863 7802
rect 2877 7800 2879 7804
rect 2893 7800 2895 7802
rect 2916 7800 2918 7802
rect 2921 7800 2923 7805
rect 2948 7804 2949 7808
rect 2994 7805 2995 7809
rect 3138 7808 3140 7811
rect 3182 7809 3184 7811
rect 2947 7800 2949 7804
rect 2968 7800 2970 7802
rect 2988 7800 2990 7802
rect 2993 7800 2995 7805
rect 3139 7804 3140 7808
rect 3183 7805 3184 7809
rect 3208 7808 3210 7812
rect 3254 7809 3256 7811
rect 3011 7800 3013 7802
rect 3095 7800 3097 7803
rect 3113 7800 3115 7803
rect 3138 7800 3140 7804
rect 3154 7800 3156 7802
rect 3177 7800 3179 7802
rect 3182 7800 3184 7805
rect 3209 7804 3210 7808
rect 3255 7805 3256 7809
rect 3822 7808 3824 7811
rect 3866 7809 3868 7811
rect 3208 7800 3210 7804
rect 3229 7800 3231 7802
rect 3249 7800 3251 7802
rect 3254 7800 3256 7805
rect 3272 7800 3274 7802
rect 3317 7800 3319 7805
rect 3322 7803 3324 7805
rect 2731 7786 2733 7789
rect 2736 7786 2738 7788
rect 2752 7786 2754 7793
rect 2861 7782 2863 7796
rect 2877 7794 2879 7796
rect 2877 7782 2879 7784
rect 2893 7782 2895 7796
rect 2916 7791 2918 7796
rect 2921 7794 2923 7796
rect 2947 7794 2949 7796
rect 2912 7787 2918 7791
rect 2916 7782 2918 7787
rect 2921 7782 2923 7784
rect 2947 7782 2949 7784
rect 2968 7782 2970 7796
rect 2988 7791 2990 7796
rect 2993 7794 2995 7796
rect 2984 7787 2990 7791
rect 2988 7782 2990 7787
rect 2993 7782 2995 7784
rect 3011 7782 3013 7796
rect 3061 7793 3063 7796
rect 3066 7793 3068 7796
rect 3095 7791 3097 7796
rect 2372 7780 2374 7782
rect 2377 7779 2379 7782
rect 2393 7780 2395 7782
rect 2409 7780 2411 7782
rect 2414 7777 2416 7782
rect 2435 7777 2437 7782
rect 2451 7780 2453 7782
rect 2467 7780 2469 7782
rect 2472 7777 2474 7782
rect 2488 7780 2490 7782
rect 2504 7780 2506 7782
rect 2509 7779 2511 7782
rect 2525 7780 2527 7782
rect 2541 7780 2543 7782
rect 2546 7777 2548 7782
rect 2567 7777 2569 7782
rect 2583 7780 2585 7782
rect 2599 7780 2601 7782
rect 2604 7777 2606 7782
rect 2620 7780 2622 7782
rect 2636 7780 2638 7782
rect 2641 7779 2643 7782
rect 2657 7780 2659 7782
rect 2673 7780 2675 7782
rect 2678 7777 2680 7782
rect 2699 7777 2701 7782
rect 2715 7780 2717 7782
rect 2731 7780 2733 7782
rect 2736 7777 2738 7782
rect 2752 7780 2754 7782
rect 3061 7777 3063 7789
rect 3066 7787 3068 7789
rect 3095 7782 3097 7787
rect 3113 7782 3115 7796
rect 3138 7794 3140 7796
rect 3138 7782 3140 7784
rect 3154 7782 3156 7796
rect 3177 7791 3179 7796
rect 3182 7794 3184 7796
rect 3208 7794 3210 7796
rect 3173 7787 3179 7791
rect 3177 7782 3179 7787
rect 3182 7782 3184 7784
rect 3208 7782 3210 7784
rect 3229 7782 3231 7796
rect 3249 7791 3251 7796
rect 3254 7794 3256 7796
rect 3245 7787 3251 7791
rect 3249 7782 3251 7787
rect 3254 7782 3256 7784
rect 3272 7782 3274 7796
rect 3317 7786 3319 7796
rect 3322 7786 3324 7793
rect 3338 7786 3340 7805
rect 3354 7796 3356 7805
rect 3359 7803 3361 7805
rect 3380 7803 3382 7805
rect 3396 7802 3398 7805
rect 3354 7786 3356 7789
rect 3359 7786 3361 7788
rect 3380 7786 3382 7788
rect 3396 7786 3398 7798
rect 3412 7796 3414 7805
rect 3417 7803 3419 7805
rect 3412 7786 3414 7789
rect 3417 7786 3419 7788
rect 3433 7786 3435 7805
rect 3449 7802 3451 7805
rect 3454 7803 3456 7805
rect 3449 7786 3451 7798
rect 3454 7786 3456 7793
rect 3470 7786 3472 7805
rect 3486 7796 3488 7805
rect 3491 7803 3493 7805
rect 3512 7803 3514 7805
rect 3528 7802 3530 7805
rect 3486 7786 3488 7789
rect 3491 7786 3493 7788
rect 3512 7786 3514 7788
rect 3528 7786 3530 7798
rect 3544 7796 3546 7805
rect 3549 7803 3551 7805
rect 3544 7786 3546 7789
rect 3549 7786 3551 7788
rect 3565 7786 3567 7805
rect 3581 7802 3583 7805
rect 3586 7803 3588 7805
rect 3581 7786 3583 7798
rect 3586 7786 3588 7793
rect 3602 7786 3604 7805
rect 3618 7796 3620 7805
rect 3623 7803 3625 7805
rect 3644 7803 3646 7805
rect 3660 7802 3662 7805
rect 3618 7786 3620 7789
rect 3623 7786 3625 7788
rect 3644 7786 3646 7788
rect 3660 7786 3662 7798
rect 3676 7796 3678 7805
rect 3681 7803 3683 7805
rect 3697 7797 3699 7805
rect 3823 7804 3824 7808
rect 3867 7805 3868 7809
rect 3892 7808 3894 7812
rect 3938 7809 3940 7811
rect 3806 7800 3808 7802
rect 3822 7800 3824 7804
rect 3838 7800 3840 7802
rect 3861 7800 3863 7802
rect 3866 7800 3868 7805
rect 3893 7804 3894 7808
rect 3939 7805 3940 7809
rect 4083 7808 4085 7811
rect 4127 7809 4129 7811
rect 3892 7800 3894 7804
rect 3913 7800 3915 7802
rect 3933 7800 3935 7802
rect 3938 7800 3940 7805
rect 4084 7804 4085 7808
rect 4128 7805 4129 7809
rect 4153 7808 4155 7812
rect 4199 7809 4201 7811
rect 3956 7800 3958 7802
rect 4040 7800 4042 7803
rect 4058 7800 4060 7803
rect 4083 7800 4085 7804
rect 4099 7800 4101 7802
rect 4122 7800 4124 7802
rect 4127 7800 4129 7805
rect 4154 7804 4155 7808
rect 4200 7805 4201 7809
rect 4153 7800 4155 7804
rect 4174 7800 4176 7802
rect 4194 7800 4196 7802
rect 4199 7800 4201 7805
rect 4217 7800 4219 7802
rect 3676 7786 3678 7789
rect 3681 7786 3683 7788
rect 3697 7786 3699 7793
rect 3806 7782 3808 7796
rect 3822 7794 3824 7796
rect 3822 7782 3824 7784
rect 3838 7782 3840 7796
rect 3861 7791 3863 7796
rect 3866 7794 3868 7796
rect 3892 7794 3894 7796
rect 3857 7787 3863 7791
rect 3861 7782 3863 7787
rect 3866 7782 3868 7784
rect 3892 7782 3894 7784
rect 3913 7782 3915 7796
rect 3933 7791 3935 7796
rect 3938 7794 3940 7796
rect 3929 7787 3935 7791
rect 3933 7782 3935 7787
rect 3938 7782 3940 7784
rect 3956 7782 3958 7796
rect 4006 7793 4008 7796
rect 4011 7793 4013 7796
rect 4040 7791 4042 7796
rect 3066 7777 3068 7779
rect 2861 7772 2863 7774
rect 2877 7771 2879 7774
rect 2893 7772 2895 7774
rect 2916 7772 2918 7774
rect 2921 7771 2923 7774
rect 2947 7771 2949 7774
rect 2968 7771 2970 7774
rect 2988 7772 2990 7774
rect 2993 7771 2995 7774
rect 3011 7772 3013 7774
rect 2947 7767 2948 7771
rect 3317 7780 3319 7782
rect 3322 7779 3324 7782
rect 3338 7780 3340 7782
rect 3354 7780 3356 7782
rect 3359 7777 3361 7782
rect 3380 7777 3382 7782
rect 3396 7780 3398 7782
rect 3412 7780 3414 7782
rect 3417 7777 3419 7782
rect 3433 7780 3435 7782
rect 3449 7780 3451 7782
rect 3095 7771 3097 7774
rect 3061 7767 3063 7769
rect 2877 7764 2879 7767
rect 2921 7764 2923 7767
rect 2947 7764 2949 7767
rect 2993 7764 2995 7767
rect 3066 7764 3068 7769
rect 2487 7742 2489 7745
rect 2511 7742 2513 7745
rect 2487 7736 2489 7738
rect 2511 7736 2513 7738
rect 3113 7732 3115 7774
rect 3138 7771 3140 7774
rect 3154 7772 3156 7774
rect 3177 7772 3179 7774
rect 3182 7771 3184 7774
rect 3208 7771 3210 7774
rect 3229 7771 3231 7774
rect 3249 7772 3251 7774
rect 3254 7771 3256 7774
rect 3272 7772 3274 7774
rect 3454 7779 3456 7782
rect 3470 7780 3472 7782
rect 3486 7780 3488 7782
rect 3491 7777 3493 7782
rect 3512 7777 3514 7782
rect 3528 7780 3530 7782
rect 3544 7780 3546 7782
rect 3549 7777 3551 7782
rect 3565 7780 3567 7782
rect 3581 7780 3583 7782
rect 3586 7779 3588 7782
rect 3602 7780 3604 7782
rect 3618 7780 3620 7782
rect 3623 7777 3625 7782
rect 3644 7777 3646 7782
rect 3660 7780 3662 7782
rect 3676 7780 3678 7782
rect 3681 7777 3683 7782
rect 3697 7780 3699 7782
rect 4006 7777 4008 7789
rect 4011 7787 4013 7789
rect 4040 7782 4042 7787
rect 4058 7782 4060 7796
rect 4083 7794 4085 7796
rect 4083 7782 4085 7784
rect 4099 7782 4101 7796
rect 4122 7791 4124 7796
rect 4127 7794 4129 7796
rect 4153 7794 4155 7796
rect 4118 7787 4124 7791
rect 4122 7782 4124 7787
rect 4127 7782 4129 7784
rect 4153 7782 4155 7784
rect 4174 7782 4176 7796
rect 4194 7791 4196 7796
rect 4199 7794 4201 7796
rect 4190 7787 4196 7791
rect 4194 7782 4196 7787
rect 4199 7782 4201 7784
rect 4217 7782 4219 7796
rect 4011 7777 4013 7779
rect 3806 7772 3808 7774
rect 3822 7771 3824 7774
rect 3838 7772 3840 7774
rect 3861 7772 3863 7774
rect 3866 7771 3868 7774
rect 3892 7771 3894 7774
rect 3913 7771 3915 7774
rect 3933 7772 3935 7774
rect 3938 7771 3940 7774
rect 3956 7772 3958 7774
rect 3208 7767 3209 7771
rect 3138 7764 3140 7767
rect 3182 7764 3184 7767
rect 3208 7764 3210 7767
rect 3254 7764 3256 7767
rect 3892 7767 3893 7771
rect 4040 7771 4042 7774
rect 4006 7767 4008 7769
rect 3822 7764 3824 7767
rect 3866 7764 3868 7767
rect 3892 7764 3894 7767
rect 3938 7764 3940 7767
rect 4011 7764 4013 7769
rect 3432 7742 3434 7745
rect 3456 7742 3458 7745
rect 3281 7740 3284 7742
rect 3288 7740 3291 7742
rect 3432 7736 3434 7738
rect 3456 7736 3458 7738
rect 4058 7736 4060 7774
rect 4083 7771 4085 7774
rect 4099 7772 4101 7774
rect 4122 7772 4124 7774
rect 4127 7771 4129 7774
rect 4153 7771 4155 7774
rect 4174 7771 4176 7774
rect 4194 7772 4196 7774
rect 4199 7771 4201 7774
rect 4217 7772 4219 7774
rect 4153 7767 4154 7771
rect 4083 7764 4085 7767
rect 4127 7764 4129 7767
rect 4153 7764 4155 7767
rect 4199 7764 4201 7767
rect 4226 7740 4229 7742
rect 4233 7740 4236 7742
rect 2507 7729 2509 7731
rect 3452 7729 3454 7731
rect 2507 7722 2509 7725
rect 3452 7722 3454 7725
rect 2496 7711 2498 7713
rect 2502 7711 2521 7713
rect 3441 7711 3443 7713
rect 3447 7711 3466 7713
rect 2487 7706 2489 7708
rect 2511 7706 2513 7708
rect 3432 7706 3434 7708
rect 3456 7706 3458 7708
rect 2487 7699 2489 7702
rect 2511 7699 2513 7702
rect 3155 7701 3157 7703
rect 3160 7701 3162 7704
rect 3176 7701 3178 7703
rect 3192 7701 3194 7703
rect 3197 7701 3199 7704
rect 3218 7701 3220 7704
rect 3234 7701 3236 7704
rect 3250 7701 3252 7703
rect 3255 7701 3257 7704
rect 3271 7701 3273 7703
rect 3432 7699 3434 7702
rect 3456 7699 3458 7702
rect 4100 7701 4102 7703
rect 4105 7701 4107 7704
rect 4121 7701 4123 7703
rect 4137 7701 4139 7703
rect 4142 7701 4144 7704
rect 4163 7701 4165 7704
rect 4179 7701 4181 7704
rect 4195 7701 4197 7703
rect 4200 7701 4202 7704
rect 4216 7701 4218 7703
rect 3155 7688 3157 7693
rect 3160 7691 3162 7693
rect 3155 7674 3157 7684
rect 3160 7674 3162 7681
rect 3176 7674 3178 7693
rect 3192 7684 3194 7693
rect 3197 7691 3199 7693
rect 3218 7691 3220 7693
rect 3234 7690 3236 7693
rect 3192 7674 3194 7677
rect 3197 7674 3199 7676
rect 3218 7674 3220 7676
rect 3234 7674 3236 7686
rect 3250 7684 3252 7693
rect 3255 7691 3257 7693
rect 3250 7674 3252 7677
rect 3255 7674 3257 7676
rect 3271 7674 3273 7693
rect 4100 7688 4102 7693
rect 4105 7691 4107 7693
rect 4100 7674 4102 7684
rect 4105 7674 4107 7681
rect 4121 7674 4123 7693
rect 4137 7684 4139 7693
rect 4142 7691 4144 7693
rect 4163 7691 4165 7693
rect 4179 7690 4181 7693
rect 4137 7674 4139 7677
rect 4142 7674 4144 7676
rect 4163 7674 4165 7676
rect 4179 7674 4181 7686
rect 4195 7684 4197 7693
rect 4200 7691 4202 7693
rect 4195 7674 4197 7677
rect 4200 7674 4202 7676
rect 4216 7674 4218 7693
rect 2372 7671 2374 7673
rect 2377 7671 2379 7674
rect 2393 7671 2395 7673
rect 2409 7671 2411 7673
rect 2414 7671 2416 7674
rect 2435 7671 2437 7674
rect 2451 7671 2453 7674
rect 2467 7671 2469 7673
rect 2472 7671 2474 7674
rect 2488 7671 2490 7673
rect 2504 7671 2506 7673
rect 2509 7671 2511 7674
rect 2525 7671 2527 7673
rect 2541 7671 2543 7673
rect 2546 7671 2548 7674
rect 2567 7671 2569 7674
rect 2583 7671 2585 7674
rect 2599 7671 2601 7673
rect 2604 7671 2606 7674
rect 2620 7671 2622 7673
rect 2636 7671 2638 7673
rect 2641 7671 2643 7674
rect 2657 7671 2659 7673
rect 2673 7671 2675 7673
rect 2678 7671 2680 7674
rect 2699 7671 2701 7674
rect 2715 7671 2717 7674
rect 2731 7671 2733 7673
rect 2736 7671 2738 7674
rect 2752 7671 2754 7673
rect 3317 7671 3319 7673
rect 3322 7671 3324 7674
rect 3338 7671 3340 7673
rect 3354 7671 3356 7673
rect 3359 7671 3361 7674
rect 3380 7671 3382 7674
rect 3396 7671 3398 7674
rect 3412 7671 3414 7673
rect 3417 7671 3419 7674
rect 3433 7671 3435 7673
rect 3449 7671 3451 7673
rect 3454 7671 3456 7674
rect 3470 7671 3472 7673
rect 3486 7671 3488 7673
rect 3491 7671 3493 7674
rect 3512 7671 3514 7674
rect 3528 7671 3530 7674
rect 3544 7671 3546 7673
rect 3549 7671 3551 7674
rect 3565 7671 3567 7673
rect 3581 7671 3583 7673
rect 3586 7671 3588 7674
rect 3602 7671 3604 7673
rect 3618 7671 3620 7673
rect 3623 7671 3625 7674
rect 3644 7671 3646 7674
rect 3660 7671 3662 7674
rect 3676 7671 3678 7673
rect 3681 7671 3683 7674
rect 3697 7671 3699 7673
rect 3155 7668 3157 7670
rect 3160 7667 3162 7670
rect 3176 7668 3178 7670
rect 3192 7668 3194 7670
rect 3197 7665 3199 7670
rect 3218 7665 3220 7670
rect 3234 7668 3236 7670
rect 3250 7668 3252 7670
rect 3255 7665 3257 7670
rect 3271 7668 3273 7670
rect 2372 7658 2374 7663
rect 2377 7661 2379 7663
rect 2372 7644 2374 7654
rect 2377 7644 2379 7651
rect 2393 7644 2395 7663
rect 2409 7654 2411 7663
rect 2414 7661 2416 7663
rect 2435 7661 2437 7663
rect 2451 7660 2453 7663
rect 2409 7644 2411 7647
rect 2414 7644 2416 7646
rect 2435 7644 2437 7646
rect 2451 7644 2453 7656
rect 2467 7654 2469 7663
rect 2472 7661 2474 7663
rect 2467 7644 2469 7647
rect 2472 7644 2474 7646
rect 2488 7644 2490 7663
rect 2504 7660 2506 7663
rect 2509 7661 2511 7663
rect 2504 7644 2506 7656
rect 2509 7644 2511 7651
rect 2525 7644 2527 7663
rect 2541 7654 2543 7663
rect 2546 7661 2548 7663
rect 2567 7661 2569 7663
rect 2583 7660 2585 7663
rect 2541 7644 2543 7647
rect 2546 7644 2548 7646
rect 2567 7644 2569 7646
rect 2583 7644 2585 7656
rect 2599 7654 2601 7663
rect 2604 7661 2606 7663
rect 2599 7644 2601 7647
rect 2604 7644 2606 7646
rect 2620 7644 2622 7663
rect 2636 7660 2638 7663
rect 2641 7661 2643 7663
rect 2636 7644 2638 7656
rect 2641 7644 2643 7651
rect 2657 7644 2659 7663
rect 2673 7654 2675 7663
rect 2678 7661 2680 7663
rect 2699 7661 2701 7663
rect 2715 7660 2717 7663
rect 2673 7644 2675 7647
rect 2678 7644 2680 7646
rect 2699 7644 2701 7646
rect 2715 7644 2717 7656
rect 2731 7654 2733 7663
rect 2736 7661 2738 7663
rect 2752 7655 2754 7663
rect 4100 7668 4102 7670
rect 4105 7667 4107 7670
rect 4121 7668 4123 7670
rect 4137 7668 4139 7670
rect 4142 7665 4144 7670
rect 4163 7665 4165 7670
rect 4179 7668 4181 7670
rect 4195 7668 4197 7670
rect 4200 7665 4202 7670
rect 4216 7668 4218 7670
rect 3317 7658 3319 7663
rect 3322 7661 3324 7663
rect 2731 7644 2733 7647
rect 2736 7644 2738 7646
rect 2752 7644 2754 7651
rect 3317 7644 3319 7654
rect 3322 7644 3324 7651
rect 3338 7644 3340 7663
rect 3354 7654 3356 7663
rect 3359 7661 3361 7663
rect 3380 7661 3382 7663
rect 3396 7660 3398 7663
rect 3354 7644 3356 7647
rect 3359 7644 3361 7646
rect 3380 7644 3382 7646
rect 3396 7644 3398 7656
rect 3412 7654 3414 7663
rect 3417 7661 3419 7663
rect 3412 7644 3414 7647
rect 3417 7644 3419 7646
rect 3433 7644 3435 7663
rect 3449 7660 3451 7663
rect 3454 7661 3456 7663
rect 3449 7644 3451 7656
rect 3454 7644 3456 7651
rect 3470 7644 3472 7663
rect 3486 7654 3488 7663
rect 3491 7661 3493 7663
rect 3512 7661 3514 7663
rect 3528 7660 3530 7663
rect 3486 7644 3488 7647
rect 3491 7644 3493 7646
rect 3512 7644 3514 7646
rect 3528 7644 3530 7656
rect 3544 7654 3546 7663
rect 3549 7661 3551 7663
rect 3544 7644 3546 7647
rect 3549 7644 3551 7646
rect 3565 7644 3567 7663
rect 3581 7660 3583 7663
rect 3586 7661 3588 7663
rect 3581 7644 3583 7656
rect 3586 7644 3588 7651
rect 3602 7644 3604 7663
rect 3618 7654 3620 7663
rect 3623 7661 3625 7663
rect 3644 7661 3646 7663
rect 3660 7660 3662 7663
rect 3618 7644 3620 7647
rect 3623 7644 3625 7646
rect 3644 7644 3646 7646
rect 3660 7644 3662 7656
rect 3676 7654 3678 7663
rect 3681 7661 3683 7663
rect 3697 7655 3699 7663
rect 3676 7644 3678 7647
rect 3681 7644 3683 7646
rect 3697 7644 3699 7651
rect 2372 7638 2374 7640
rect 2377 7637 2379 7640
rect 2393 7638 2395 7640
rect 2409 7638 2411 7640
rect 2414 7635 2416 7640
rect 2435 7635 2437 7640
rect 2451 7638 2453 7640
rect 2467 7638 2469 7640
rect 2472 7635 2474 7640
rect 2488 7638 2490 7640
rect 2504 7638 2506 7640
rect 2509 7637 2511 7640
rect 2525 7638 2527 7640
rect 2541 7638 2543 7640
rect 2546 7635 2548 7640
rect 2567 7635 2569 7640
rect 2583 7638 2585 7640
rect 2599 7638 2601 7640
rect 2604 7635 2606 7640
rect 2620 7638 2622 7640
rect 2636 7638 2638 7640
rect 2641 7637 2643 7640
rect 2657 7638 2659 7640
rect 2673 7638 2675 7640
rect 2678 7635 2680 7640
rect 2699 7635 2701 7640
rect 2715 7638 2717 7640
rect 2731 7638 2733 7640
rect 2736 7635 2738 7640
rect 2752 7638 2754 7640
rect 3317 7638 3319 7640
rect 3322 7637 3324 7640
rect 3338 7638 3340 7640
rect 3354 7638 3356 7640
rect 3359 7635 3361 7640
rect 3380 7635 3382 7640
rect 3396 7638 3398 7640
rect 3412 7638 3414 7640
rect 3417 7635 3419 7640
rect 3433 7638 3435 7640
rect 3449 7638 3451 7640
rect 3454 7637 3456 7640
rect 3470 7638 3472 7640
rect 3486 7638 3488 7640
rect 3491 7635 3493 7640
rect 3512 7635 3514 7640
rect 3528 7638 3530 7640
rect 3544 7638 3546 7640
rect 3549 7635 3551 7640
rect 3565 7638 3567 7640
rect 3581 7638 3583 7640
rect 3586 7637 3588 7640
rect 3602 7638 3604 7640
rect 3618 7638 3620 7640
rect 3623 7635 3625 7640
rect 3644 7635 3646 7640
rect 3660 7638 3662 7640
rect 3676 7638 3678 7640
rect 3681 7635 3683 7640
rect 3697 7638 3699 7640
rect 3155 7615 3157 7617
rect 3160 7615 3162 7618
rect 3176 7615 3178 7617
rect 3192 7615 3194 7617
rect 3197 7615 3199 7618
rect 3218 7615 3220 7618
rect 3234 7615 3236 7618
rect 3250 7615 3252 7617
rect 3255 7615 3257 7618
rect 3271 7615 3273 7617
rect 4100 7615 4102 7617
rect 4105 7615 4107 7618
rect 4121 7615 4123 7617
rect 4137 7615 4139 7617
rect 4142 7615 4144 7618
rect 4163 7615 4165 7618
rect 4179 7615 4181 7618
rect 4195 7615 4197 7617
rect 4200 7615 4202 7618
rect 4216 7615 4218 7617
rect 3155 7602 3157 7607
rect 3160 7605 3162 7607
rect 3155 7588 3157 7598
rect 3160 7588 3162 7595
rect 3176 7588 3178 7607
rect 3192 7598 3194 7607
rect 3197 7605 3199 7607
rect 3218 7605 3220 7607
rect 3234 7604 3236 7607
rect 3192 7588 3194 7591
rect 3197 7588 3199 7590
rect 3218 7588 3220 7590
rect 3234 7588 3236 7600
rect 3250 7598 3252 7607
rect 3255 7605 3257 7607
rect 3250 7588 3252 7591
rect 3255 7588 3257 7590
rect 3271 7588 3273 7607
rect 4100 7602 4102 7607
rect 4105 7605 4107 7607
rect 3293 7594 3296 7596
rect 3300 7594 3303 7596
rect 4100 7588 4102 7598
rect 4105 7588 4107 7595
rect 4121 7588 4123 7607
rect 4137 7598 4139 7607
rect 4142 7605 4144 7607
rect 4163 7605 4165 7607
rect 4179 7604 4181 7607
rect 4137 7588 4139 7591
rect 4142 7588 4144 7590
rect 4163 7588 4165 7590
rect 4179 7588 4181 7600
rect 4195 7598 4197 7607
rect 4200 7605 4202 7607
rect 4195 7588 4197 7591
rect 4200 7588 4202 7590
rect 4216 7588 4218 7607
rect 4238 7594 4241 7596
rect 4245 7594 4248 7596
rect 2372 7585 2374 7587
rect 2377 7585 2379 7588
rect 2393 7585 2395 7587
rect 2409 7585 2411 7587
rect 2414 7585 2416 7588
rect 2435 7585 2437 7588
rect 2451 7585 2453 7588
rect 2467 7585 2469 7587
rect 2472 7585 2474 7588
rect 2488 7585 2490 7587
rect 2504 7585 2506 7587
rect 2509 7585 2511 7588
rect 2525 7585 2527 7587
rect 2541 7585 2543 7587
rect 2546 7585 2548 7588
rect 2567 7585 2569 7588
rect 2583 7585 2585 7588
rect 2599 7585 2601 7587
rect 2604 7585 2606 7588
rect 2620 7585 2622 7587
rect 2636 7585 2638 7587
rect 2641 7585 2643 7588
rect 2657 7585 2659 7587
rect 2673 7585 2675 7587
rect 2678 7585 2680 7588
rect 2699 7585 2701 7588
rect 2715 7585 2717 7588
rect 2731 7585 2733 7587
rect 2736 7585 2738 7588
rect 2752 7585 2754 7587
rect 3317 7585 3319 7587
rect 3322 7585 3324 7588
rect 3338 7585 3340 7587
rect 3354 7585 3356 7587
rect 3359 7585 3361 7588
rect 3380 7585 3382 7588
rect 3396 7585 3398 7588
rect 3412 7585 3414 7587
rect 3417 7585 3419 7588
rect 3433 7585 3435 7587
rect 3449 7585 3451 7587
rect 3454 7585 3456 7588
rect 3470 7585 3472 7587
rect 3486 7585 3488 7587
rect 3491 7585 3493 7588
rect 3512 7585 3514 7588
rect 3528 7585 3530 7588
rect 3544 7585 3546 7587
rect 3549 7585 3551 7588
rect 3565 7585 3567 7587
rect 3581 7585 3583 7587
rect 3586 7585 3588 7588
rect 3602 7585 3604 7587
rect 3618 7585 3620 7587
rect 3623 7585 3625 7588
rect 3644 7585 3646 7588
rect 3660 7585 3662 7588
rect 3676 7585 3678 7587
rect 3681 7585 3683 7588
rect 3697 7585 3699 7587
rect 3155 7582 3157 7584
rect 3160 7581 3162 7584
rect 3176 7582 3178 7584
rect 3192 7582 3194 7584
rect 3197 7579 3199 7584
rect 3218 7579 3220 7584
rect 3234 7582 3236 7584
rect 3250 7582 3252 7584
rect 3255 7579 3257 7584
rect 3271 7582 3273 7584
rect 2372 7572 2374 7577
rect 2377 7575 2379 7577
rect 2372 7558 2374 7568
rect 2377 7558 2379 7565
rect 2393 7558 2395 7577
rect 2409 7568 2411 7577
rect 2414 7575 2416 7577
rect 2435 7575 2437 7577
rect 2451 7574 2453 7577
rect 2409 7558 2411 7561
rect 2414 7558 2416 7560
rect 2435 7558 2437 7560
rect 2451 7558 2453 7570
rect 2467 7568 2469 7577
rect 2472 7575 2474 7577
rect 2467 7558 2469 7561
rect 2472 7558 2474 7560
rect 2488 7558 2490 7577
rect 2504 7574 2506 7577
rect 2509 7575 2511 7577
rect 2504 7558 2506 7570
rect 2509 7558 2511 7565
rect 2525 7558 2527 7577
rect 2541 7568 2543 7577
rect 2546 7575 2548 7577
rect 2567 7575 2569 7577
rect 2583 7574 2585 7577
rect 2541 7558 2543 7561
rect 2546 7558 2548 7560
rect 2567 7558 2569 7560
rect 2583 7558 2585 7570
rect 2599 7568 2601 7577
rect 2604 7575 2606 7577
rect 2599 7558 2601 7561
rect 2604 7558 2606 7560
rect 2620 7558 2622 7577
rect 2636 7574 2638 7577
rect 2641 7575 2643 7577
rect 2636 7558 2638 7570
rect 2641 7558 2643 7565
rect 2657 7558 2659 7577
rect 2673 7568 2675 7577
rect 2678 7575 2680 7577
rect 2699 7575 2701 7577
rect 2715 7574 2717 7577
rect 2673 7558 2675 7561
rect 2678 7558 2680 7560
rect 2699 7558 2701 7560
rect 2715 7558 2717 7570
rect 2731 7568 2733 7577
rect 2736 7575 2738 7577
rect 2752 7569 2754 7577
rect 4100 7582 4102 7584
rect 4105 7581 4107 7584
rect 4121 7582 4123 7584
rect 4137 7582 4139 7584
rect 4142 7579 4144 7584
rect 4163 7579 4165 7584
rect 4179 7582 4181 7584
rect 4195 7582 4197 7584
rect 4200 7579 4202 7584
rect 4216 7582 4218 7584
rect 3317 7572 3319 7577
rect 3322 7575 3324 7577
rect 2731 7558 2733 7561
rect 2736 7558 2738 7560
rect 2752 7558 2754 7565
rect 3317 7558 3319 7568
rect 3322 7558 3324 7565
rect 3338 7558 3340 7577
rect 3354 7568 3356 7577
rect 3359 7575 3361 7577
rect 3380 7575 3382 7577
rect 3396 7574 3398 7577
rect 3354 7558 3356 7561
rect 3359 7558 3361 7560
rect 3380 7558 3382 7560
rect 3396 7558 3398 7570
rect 3412 7568 3414 7577
rect 3417 7575 3419 7577
rect 3412 7558 3414 7561
rect 3417 7558 3419 7560
rect 3433 7558 3435 7577
rect 3449 7574 3451 7577
rect 3454 7575 3456 7577
rect 3449 7558 3451 7570
rect 3454 7558 3456 7565
rect 3470 7558 3472 7577
rect 3486 7568 3488 7577
rect 3491 7575 3493 7577
rect 3512 7575 3514 7577
rect 3528 7574 3530 7577
rect 3486 7558 3488 7561
rect 3491 7558 3493 7560
rect 3512 7558 3514 7560
rect 3528 7558 3530 7570
rect 3544 7568 3546 7577
rect 3549 7575 3551 7577
rect 3544 7558 3546 7561
rect 3549 7558 3551 7560
rect 3565 7558 3567 7577
rect 3581 7574 3583 7577
rect 3586 7575 3588 7577
rect 3581 7558 3583 7570
rect 3586 7558 3588 7565
rect 3602 7558 3604 7577
rect 3618 7568 3620 7577
rect 3623 7575 3625 7577
rect 3644 7575 3646 7577
rect 3660 7574 3662 7577
rect 3618 7558 3620 7561
rect 3623 7558 3625 7560
rect 3644 7558 3646 7560
rect 3660 7558 3662 7570
rect 3676 7568 3678 7577
rect 3681 7575 3683 7577
rect 3697 7569 3699 7577
rect 3676 7558 3678 7561
rect 3681 7558 3683 7560
rect 3697 7558 3699 7565
rect 2372 7552 2374 7554
rect 2377 7551 2379 7554
rect 2393 7552 2395 7554
rect 2409 7552 2411 7554
rect 2414 7549 2416 7554
rect 2435 7549 2437 7554
rect 2451 7552 2453 7554
rect 2467 7552 2469 7554
rect 2472 7549 2474 7554
rect 2488 7552 2490 7554
rect 2504 7552 2506 7554
rect 2509 7551 2511 7554
rect 2525 7552 2527 7554
rect 2541 7552 2543 7554
rect 2546 7549 2548 7554
rect 2567 7549 2569 7554
rect 2583 7552 2585 7554
rect 2599 7552 2601 7554
rect 2604 7549 2606 7554
rect 2620 7552 2622 7554
rect 2636 7552 2638 7554
rect 2641 7551 2643 7554
rect 2657 7552 2659 7554
rect 2673 7552 2675 7554
rect 2678 7549 2680 7554
rect 2699 7549 2701 7554
rect 2715 7552 2717 7554
rect 2731 7552 2733 7554
rect 2736 7549 2738 7554
rect 2752 7552 2754 7554
rect 3317 7552 3319 7554
rect 3322 7551 3324 7554
rect 3338 7552 3340 7554
rect 3354 7552 3356 7554
rect 3359 7549 3361 7554
rect 3380 7549 3382 7554
rect 3396 7552 3398 7554
rect 3412 7552 3414 7554
rect 3417 7549 3419 7554
rect 3433 7552 3435 7554
rect 3449 7552 3451 7554
rect 3454 7551 3456 7554
rect 3470 7552 3472 7554
rect 3486 7552 3488 7554
rect 3491 7549 3493 7554
rect 3512 7549 3514 7554
rect 3528 7552 3530 7554
rect 3544 7552 3546 7554
rect 3549 7549 3551 7554
rect 3565 7552 3567 7554
rect 3581 7552 3583 7554
rect 3586 7551 3588 7554
rect 3602 7552 3604 7554
rect 3618 7552 3620 7554
rect 3623 7549 3625 7554
rect 3644 7549 3646 7554
rect 3660 7552 3662 7554
rect 3676 7552 3678 7554
rect 3681 7549 3683 7554
rect 3697 7552 3699 7554
rect 2604 7514 2606 7517
rect 2628 7514 2630 7517
rect 3549 7514 3551 7517
rect 3573 7514 3575 7517
rect 2604 7508 2606 7510
rect 2628 7508 2630 7510
rect 3549 7508 3551 7510
rect 3573 7508 3575 7510
rect 2624 7503 2626 7505
rect 3569 7503 3571 7505
rect 2624 7496 2626 7499
rect 3569 7496 3571 7499
rect 2613 7485 2615 7487
rect 2619 7485 2638 7487
rect 3558 7485 3560 7487
rect 3564 7485 3583 7487
rect 2604 7480 2606 7482
rect 2628 7480 2630 7482
rect 3549 7480 3551 7482
rect 3573 7480 3575 7482
rect 2604 7473 2606 7476
rect 2628 7473 2630 7476
rect 3549 7473 3551 7476
rect 3573 7473 3575 7476
rect 2372 7445 2374 7447
rect 2377 7445 2379 7448
rect 2393 7445 2395 7447
rect 2409 7445 2411 7447
rect 2414 7445 2416 7448
rect 2435 7445 2437 7448
rect 2451 7445 2453 7448
rect 2467 7445 2469 7447
rect 2472 7445 2474 7448
rect 2488 7445 2490 7447
rect 2504 7445 2506 7447
rect 2509 7445 2511 7448
rect 2525 7445 2527 7447
rect 2541 7445 2543 7447
rect 2546 7445 2548 7448
rect 2567 7445 2569 7448
rect 2583 7445 2585 7448
rect 2599 7445 2601 7447
rect 2604 7445 2606 7448
rect 2620 7445 2622 7447
rect 2636 7445 2638 7447
rect 2641 7445 2643 7448
rect 2657 7445 2659 7447
rect 2673 7445 2675 7447
rect 2678 7445 2680 7448
rect 2699 7445 2701 7448
rect 2715 7445 2717 7448
rect 2731 7445 2733 7447
rect 2736 7445 2738 7448
rect 2752 7445 2754 7447
rect 3317 7445 3319 7447
rect 3322 7445 3324 7448
rect 3338 7445 3340 7447
rect 3354 7445 3356 7447
rect 3359 7445 3361 7448
rect 3380 7445 3382 7448
rect 3396 7445 3398 7448
rect 3412 7445 3414 7447
rect 3417 7445 3419 7448
rect 3433 7445 3435 7447
rect 3449 7445 3451 7447
rect 3454 7445 3456 7448
rect 3470 7445 3472 7447
rect 3486 7445 3488 7447
rect 3491 7445 3493 7448
rect 3512 7445 3514 7448
rect 3528 7445 3530 7448
rect 3544 7445 3546 7447
rect 3549 7445 3551 7448
rect 3565 7445 3567 7447
rect 3581 7445 3583 7447
rect 3586 7445 3588 7448
rect 3602 7445 3604 7447
rect 3618 7445 3620 7447
rect 3623 7445 3625 7448
rect 3644 7445 3646 7448
rect 3660 7445 3662 7448
rect 3676 7445 3678 7447
rect 3681 7445 3683 7448
rect 3697 7445 3699 7447
rect 2372 7432 2374 7437
rect 2377 7435 2379 7437
rect 2372 7418 2374 7428
rect 2377 7418 2379 7425
rect 2393 7418 2395 7437
rect 2409 7428 2411 7437
rect 2414 7435 2416 7437
rect 2435 7435 2437 7437
rect 2451 7434 2453 7437
rect 2409 7418 2411 7421
rect 2414 7418 2416 7420
rect 2435 7418 2437 7420
rect 2451 7418 2453 7430
rect 2467 7428 2469 7437
rect 2472 7435 2474 7437
rect 2467 7418 2469 7421
rect 2472 7418 2474 7420
rect 2488 7418 2490 7437
rect 2504 7434 2506 7437
rect 2509 7435 2511 7437
rect 2504 7418 2506 7430
rect 2509 7418 2511 7425
rect 2525 7418 2527 7437
rect 2541 7428 2543 7437
rect 2546 7435 2548 7437
rect 2567 7435 2569 7437
rect 2583 7434 2585 7437
rect 2541 7418 2543 7421
rect 2546 7418 2548 7420
rect 2567 7418 2569 7420
rect 2583 7418 2585 7430
rect 2599 7428 2601 7437
rect 2604 7435 2606 7437
rect 2599 7418 2601 7421
rect 2604 7418 2606 7420
rect 2620 7418 2622 7437
rect 2636 7434 2638 7437
rect 2641 7435 2643 7437
rect 2636 7418 2638 7430
rect 2641 7418 2643 7425
rect 2657 7418 2659 7437
rect 2673 7428 2675 7437
rect 2678 7435 2680 7437
rect 2699 7435 2701 7437
rect 2715 7434 2717 7437
rect 2673 7418 2675 7421
rect 2678 7418 2680 7420
rect 2699 7418 2701 7420
rect 2715 7418 2717 7430
rect 2731 7428 2733 7437
rect 2736 7435 2738 7437
rect 2752 7429 2754 7437
rect 3317 7432 3319 7437
rect 3322 7435 3324 7437
rect 2731 7418 2733 7421
rect 2736 7418 2738 7420
rect 2752 7418 2754 7425
rect 3317 7418 3319 7428
rect 3322 7418 3324 7425
rect 3338 7418 3340 7437
rect 3354 7428 3356 7437
rect 3359 7435 3361 7437
rect 3380 7435 3382 7437
rect 3396 7434 3398 7437
rect 3354 7418 3356 7421
rect 3359 7418 3361 7420
rect 3380 7418 3382 7420
rect 3396 7418 3398 7430
rect 3412 7428 3414 7437
rect 3417 7435 3419 7437
rect 3412 7418 3414 7421
rect 3417 7418 3419 7420
rect 3433 7418 3435 7437
rect 3449 7434 3451 7437
rect 3454 7435 3456 7437
rect 3449 7418 3451 7430
rect 3454 7418 3456 7425
rect 3470 7418 3472 7437
rect 3486 7428 3488 7437
rect 3491 7435 3493 7437
rect 3512 7435 3514 7437
rect 3528 7434 3530 7437
rect 3486 7418 3488 7421
rect 3491 7418 3493 7420
rect 3512 7418 3514 7420
rect 3528 7418 3530 7430
rect 3544 7428 3546 7437
rect 3549 7435 3551 7437
rect 3544 7418 3546 7421
rect 3549 7418 3551 7420
rect 3565 7418 3567 7437
rect 3581 7434 3583 7437
rect 3586 7435 3588 7437
rect 3581 7418 3583 7430
rect 3586 7418 3588 7425
rect 3602 7418 3604 7437
rect 3618 7428 3620 7437
rect 3623 7435 3625 7437
rect 3644 7435 3646 7437
rect 3660 7434 3662 7437
rect 3618 7418 3620 7421
rect 3623 7418 3625 7420
rect 3644 7418 3646 7420
rect 3660 7418 3662 7430
rect 3676 7428 3678 7437
rect 3681 7435 3683 7437
rect 3697 7429 3699 7437
rect 3676 7418 3678 7421
rect 3681 7418 3683 7420
rect 3697 7418 3699 7425
rect 2372 7412 2374 7414
rect 2377 7411 2379 7414
rect 2393 7412 2395 7414
rect 2409 7412 2411 7414
rect 2414 7409 2416 7414
rect 2435 7409 2437 7414
rect 2451 7412 2453 7414
rect 2467 7412 2469 7414
rect 2472 7409 2474 7414
rect 2488 7412 2490 7414
rect 2504 7412 2506 7414
rect 2509 7411 2511 7414
rect 2525 7412 2527 7414
rect 2541 7412 2543 7414
rect 2546 7409 2548 7414
rect 2567 7409 2569 7414
rect 2583 7412 2585 7414
rect 2599 7412 2601 7414
rect 2604 7409 2606 7414
rect 2620 7412 2622 7414
rect 2636 7412 2638 7414
rect 2641 7411 2643 7414
rect 2657 7412 2659 7414
rect 2673 7412 2675 7414
rect 2678 7409 2680 7414
rect 2699 7409 2701 7414
rect 2715 7412 2717 7414
rect 2731 7412 2733 7414
rect 2736 7409 2738 7414
rect 2752 7412 2754 7414
rect 3317 7412 3319 7414
rect 3322 7411 3324 7414
rect 3338 7412 3340 7414
rect 3354 7412 3356 7414
rect 3359 7409 3361 7414
rect 3380 7409 3382 7414
rect 3396 7412 3398 7414
rect 3412 7412 3414 7414
rect 3417 7409 3419 7414
rect 3433 7412 3435 7414
rect 3449 7412 3451 7414
rect 3454 7411 3456 7414
rect 3470 7412 3472 7414
rect 3486 7412 3488 7414
rect 3491 7409 3493 7414
rect 3512 7409 3514 7414
rect 3528 7412 3530 7414
rect 3544 7412 3546 7414
rect 3549 7409 3551 7414
rect 3565 7412 3567 7414
rect 3581 7412 3583 7414
rect 3586 7411 3588 7414
rect 3602 7412 3604 7414
rect 3618 7412 3620 7414
rect 3623 7409 3625 7414
rect 3644 7409 3646 7414
rect 3660 7412 3662 7414
rect 3676 7412 3678 7414
rect 3681 7409 3683 7414
rect 3697 7412 3699 7414
rect 4579 9355 5073 9786
rect 4634 8035 4644 8037
rect 4634 8034 4636 8035
rect 4642 8034 4644 8035
rect 4650 8035 4660 8037
rect 4650 8034 4652 8035
rect 4658 8034 4660 8035
rect 4677 8035 4687 8037
rect 4677 8034 4679 8035
rect 4685 8034 4687 8035
rect 4693 8035 4703 8037
rect 4693 8034 4695 8035
rect 4701 8034 4703 8035
rect 4718 8035 4728 8037
rect 4718 8034 4720 8035
rect 4726 8034 4728 8035
rect 4734 8035 4744 8037
rect 4734 8034 4736 8035
rect 4742 8034 4744 8035
rect 4579 8015 4581 8017
rect 4587 8015 4589 8017
rect 4595 8016 4621 8018
rect 4595 8015 4597 8016
rect 4603 8015 4605 8016
rect 4611 8015 4613 8016
rect 4619 8015 4621 8016
rect 4579 7960 4581 7975
rect 4576 7954 4581 7960
rect 4587 7954 4589 7975
rect 4595 7974 4597 7975
rect 4603 7974 4605 7975
rect 4611 7974 4613 7975
rect 4619 7974 4621 7975
rect 4595 7972 4621 7974
rect 4634 7974 4636 7975
rect 4642 7974 4644 7975
rect 4650 7974 4652 7975
rect 4658 7974 4660 7975
rect 4634 7972 4660 7974
rect 4677 7974 4679 7975
rect 4685 7974 4687 7975
rect 4693 7974 4695 7975
rect 4701 7974 4703 7975
rect 4718 7974 4720 7975
rect 4726 7974 4728 7975
rect 4734 7974 4736 7975
rect 4742 7974 4744 7975
rect 4595 7965 4599 7972
rect 4597 7959 4599 7965
rect 4579 7952 4589 7954
rect 4579 7945 4581 7952
rect 4587 7945 4589 7952
rect 4595 7948 4599 7959
rect 4634 7963 4641 7972
rect 4634 7950 4635 7963
rect 4639 7950 4641 7963
rect 4634 7948 4641 7950
rect 4677 7965 4744 7974
rect 4677 7952 4678 7965
rect 4682 7963 4744 7965
rect 4682 7954 4711 7963
rect 4717 7954 4744 7963
rect 4682 7952 4744 7954
rect 4677 7950 4744 7952
rect 4677 7948 4703 7950
rect 4595 7946 4621 7948
rect 4595 7945 4597 7946
rect 4603 7945 4605 7946
rect 4611 7945 4613 7946
rect 4619 7945 4621 7946
rect 4634 7946 4660 7948
rect 4634 7945 4636 7946
rect 4642 7945 4644 7946
rect 4650 7945 4652 7946
rect 4658 7945 4660 7946
rect 4677 7945 4679 7948
rect 4685 7945 4687 7948
rect 4693 7945 4695 7948
rect 4701 7945 4703 7948
rect 4718 7948 4744 7950
rect 4718 7945 4720 7948
rect 4726 7945 4728 7948
rect 4734 7945 4736 7948
rect 4742 7945 4744 7948
rect 4579 7887 4581 7889
rect 4587 7887 4589 7889
rect 4595 7888 4597 7889
rect 4603 7888 4605 7889
rect 4611 7888 4613 7889
rect 4619 7888 4621 7889
rect 4595 7886 4621 7888
rect 4634 7856 4636 7857
rect 4642 7856 4644 7857
rect 4650 7856 4652 7857
rect 4658 7856 4660 7857
rect 4634 7854 4660 7856
rect 4677 7856 4679 7857
rect 4685 7856 4687 7857
rect 4693 7856 4695 7857
rect 4701 7856 4703 7857
rect 4677 7854 4703 7856
rect 4718 7856 4720 7857
rect 4726 7856 4728 7857
rect 4734 7856 4736 7857
rect 4742 7856 4744 7857
rect 4718 7854 4744 7856
rect 4579 5800 5054 6238
rect 99 5325 1031 5800
rect 4148 5306 5054 5800
<< polycontact >>
rect 1797 9952 1818 9961
rect 1797 9874 1818 9883
rect 2106 9952 2127 9961
rect 2106 9874 2127 9883
rect 2415 9952 2436 9961
rect 2415 9874 2436 9883
rect 2724 9952 2745 9961
rect 2724 9874 2745 9883
rect 3033 9952 3054 9961
rect 3033 9874 3054 9883
rect 3960 9952 3981 9961
rect 3960 9874 3981 9883
rect 1803 9827 1812 9831
rect 2112 9827 2121 9831
rect 2421 9827 2430 9831
rect 2730 9827 2739 9831
rect 3039 9827 3048 9831
rect 3966 9827 3975 9831
rect 1813 9808 1819 9812
rect 2122 9808 2128 9812
rect 2431 9808 2437 9812
rect 2740 9808 2746 9812
rect 3049 9808 3055 9812
rect 3976 9808 3982 9812
rect 2861 9333 2865 9337
rect 2898 9333 2902 9337
rect 2918 9333 2922 9337
rect 2956 9333 2960 9337
rect 2993 9333 2997 9337
rect 3030 9333 3034 9337
rect 3050 9333 3054 9337
rect 3088 9333 3092 9337
rect 3125 9333 3129 9337
rect 3162 9333 3166 9337
rect 3182 9333 3186 9337
rect 3220 9333 3224 9337
rect 3257 9333 3261 9337
rect 3294 9333 3298 9337
rect 3314 9333 3318 9337
rect 3352 9333 3356 9337
rect 3806 9333 3810 9337
rect 3843 9333 3847 9337
rect 3863 9333 3867 9337
rect 3901 9333 3905 9337
rect 3938 9333 3942 9337
rect 3975 9333 3979 9337
rect 3995 9333 3999 9337
rect 4033 9333 4037 9337
rect 4070 9333 4074 9337
rect 4107 9333 4111 9337
rect 4127 9333 4131 9337
rect 4165 9333 4169 9337
rect 4202 9333 4206 9337
rect 4239 9333 4243 9337
rect 4259 9333 4263 9337
rect 4297 9333 4301 9337
rect 2855 9313 2859 9317
rect 2873 9315 2877 9319
rect 2509 9300 2513 9304
rect 2546 9300 2550 9304
rect 2566 9300 2570 9304
rect 2604 9300 2608 9304
rect 2933 9315 2937 9319
rect 2891 9306 2895 9313
rect 2949 9306 2953 9313
rect 2970 9310 2974 9314
rect 2987 9313 2991 9317
rect 3005 9315 3009 9319
rect 3065 9315 3069 9319
rect 3023 9306 3027 9313
rect 3081 9306 3085 9313
rect 3102 9310 3106 9314
rect 3119 9313 3123 9317
rect 3137 9315 3141 9319
rect 3197 9315 3201 9319
rect 3155 9306 3159 9313
rect 3213 9306 3217 9313
rect 3234 9310 3238 9314
rect 3251 9313 3255 9317
rect 3269 9315 3273 9319
rect 3329 9315 3333 9319
rect 3287 9306 3291 9313
rect 3345 9306 3349 9313
rect 3366 9310 3370 9314
rect 3800 9313 3804 9317
rect 3818 9315 3822 9319
rect 3454 9300 3458 9304
rect 3491 9300 3495 9304
rect 3511 9300 3515 9304
rect 3549 9300 3553 9304
rect 3878 9315 3882 9319
rect 3836 9306 3840 9313
rect 3894 9306 3898 9313
rect 3915 9310 3919 9314
rect 3932 9313 3936 9317
rect 3950 9315 3954 9319
rect 4010 9315 4014 9319
rect 3968 9306 3972 9313
rect 4026 9306 4030 9313
rect 4047 9310 4051 9314
rect 4064 9313 4068 9317
rect 4082 9315 4086 9319
rect 4142 9315 4146 9319
rect 4100 9306 4104 9313
rect 4158 9306 4162 9313
rect 4179 9310 4183 9314
rect 4196 9313 4200 9317
rect 4214 9315 4218 9319
rect 4274 9315 4278 9319
rect 4232 9306 4236 9313
rect 4290 9306 4294 9313
rect 4311 9310 4315 9314
rect 2861 9292 2865 9296
rect 2898 9290 2902 9294
rect 2918 9290 2922 9294
rect 2954 9290 2958 9294
rect 2993 9292 2997 9296
rect 3030 9290 3034 9294
rect 3050 9290 3054 9294
rect 3086 9290 3090 9294
rect 3125 9292 3129 9296
rect 3162 9290 3166 9294
rect 3182 9290 3186 9294
rect 3218 9290 3222 9294
rect 3257 9292 3261 9296
rect 3294 9290 3298 9294
rect 3314 9290 3318 9294
rect 3350 9290 3354 9294
rect 3806 9292 3810 9296
rect 3843 9290 3847 9294
rect 3863 9290 3867 9294
rect 3899 9290 3903 9294
rect 3938 9292 3942 9296
rect 3975 9290 3979 9294
rect 3995 9290 3999 9294
rect 4031 9290 4035 9294
rect 4070 9292 4074 9296
rect 4107 9290 4111 9294
rect 4127 9290 4131 9294
rect 4163 9290 4167 9294
rect 4202 9292 4206 9296
rect 4239 9290 4243 9294
rect 4259 9290 4263 9294
rect 4295 9290 4299 9294
rect 2503 9280 2507 9284
rect 2521 9282 2525 9286
rect 2581 9282 2585 9286
rect 2539 9273 2543 9280
rect 2597 9273 2601 9280
rect 2616 9277 2620 9281
rect 3448 9280 3452 9284
rect 3466 9282 3470 9286
rect 3526 9282 3530 9286
rect 3484 9273 3488 9280
rect 3542 9273 3546 9280
rect 3561 9277 3565 9281
rect 2509 9259 2513 9263
rect 2546 9257 2550 9261
rect 2566 9257 2570 9261
rect 2602 9257 2606 9261
rect 2877 9249 2881 9253
rect 2921 9249 2925 9253
rect 2948 9249 2952 9253
rect 2993 9249 2997 9253
rect 3066 9256 3070 9260
rect 2627 9236 2631 9240
rect 3031 9242 3035 9246
rect 2510 9227 2514 9231
rect 2857 9229 2861 9233
rect 2889 9230 2893 9234
rect 2908 9229 2912 9233
rect 2964 9230 2968 9234
rect 2980 9229 2984 9233
rect 3007 9229 3011 9233
rect 3147 9256 3151 9260
rect 3454 9259 3458 9263
rect 3058 9238 3062 9242
rect 3085 9234 3089 9238
rect 3112 9242 3116 9246
rect 3491 9257 3495 9261
rect 3511 9257 3515 9261
rect 3547 9257 3551 9261
rect 3139 9238 3143 9242
rect 3166 9234 3170 9238
rect 3822 9249 3826 9253
rect 3866 9249 3870 9253
rect 3893 9249 3897 9253
rect 3938 9249 3942 9253
rect 4011 9256 4015 9260
rect 3572 9236 3576 9240
rect 3976 9242 3980 9246
rect 3064 9220 3068 9224
rect 3455 9227 3459 9231
rect 3802 9229 3806 9233
rect 3145 9220 3149 9224
rect 3834 9230 3838 9234
rect 3853 9229 3857 9233
rect 3909 9230 3913 9234
rect 3925 9229 3929 9233
rect 3952 9229 3956 9233
rect 4092 9256 4096 9260
rect 4003 9238 4007 9242
rect 4030 9234 4034 9238
rect 4057 9242 4061 9246
rect 4084 9238 4088 9242
rect 4111 9234 4115 9238
rect 4009 9220 4013 9224
rect 4090 9220 4094 9224
rect 2874 9212 2878 9216
rect 2918 9211 2922 9215
rect 2943 9212 2948 9216
rect 2990 9211 2994 9215
rect 3819 9212 3823 9216
rect 3863 9211 3867 9215
rect 3888 9212 3893 9216
rect 3935 9211 3939 9215
rect 2509 9198 2513 9202
rect 2547 9198 2551 9202
rect 2567 9198 2571 9202
rect 2604 9198 2608 9202
rect 3454 9198 3458 9202
rect 3492 9198 3496 9202
rect 3512 9198 3516 9202
rect 3549 9198 3553 9202
rect 2497 9175 2501 9179
rect 2532 9180 2536 9184
rect 2516 9171 2520 9178
rect 2574 9171 2578 9178
rect 2592 9180 2596 9184
rect 2874 9182 2878 9186
rect 2918 9183 2922 9187
rect 2610 9178 2614 9182
rect 2943 9182 2948 9186
rect 2990 9183 2994 9187
rect 3066 9180 3070 9184
rect 3147 9180 3151 9184
rect 2857 9165 2861 9169
rect 2511 9155 2515 9159
rect 2547 9155 2551 9159
rect 2567 9155 2571 9159
rect 2604 9157 2608 9161
rect 2889 9164 2893 9168
rect 2908 9165 2912 9169
rect 2964 9164 2968 9168
rect 2980 9165 2984 9169
rect 3007 9165 3011 9169
rect 3055 9164 3061 9168
rect 3136 9164 3142 9168
rect 3442 9175 3446 9179
rect 3477 9180 3481 9184
rect 3461 9171 3465 9178
rect 3519 9171 3523 9178
rect 3537 9180 3541 9184
rect 3819 9182 3823 9186
rect 3863 9183 3867 9187
rect 3555 9178 3559 9182
rect 3888 9182 3893 9186
rect 3935 9183 3939 9187
rect 4011 9180 4015 9184
rect 4092 9180 4096 9184
rect 3802 9165 3806 9169
rect 3456 9155 3460 9159
rect 3492 9155 3496 9159
rect 3512 9155 3516 9159
rect 3549 9157 3553 9161
rect 3834 9164 3838 9168
rect 3853 9165 3857 9169
rect 3909 9164 3913 9168
rect 3925 9165 3929 9169
rect 3952 9165 3956 9169
rect 4000 9164 4006 9168
rect 4081 9164 4087 9168
rect 2877 9145 2881 9149
rect 2921 9145 2925 9149
rect 2948 9145 2952 9149
rect 2993 9145 2997 9149
rect 3064 9144 3068 9148
rect 3145 9144 3149 9148
rect 3822 9145 3826 9149
rect 3866 9145 3870 9149
rect 3893 9145 3897 9149
rect 3938 9145 3942 9149
rect 4009 9144 4013 9148
rect 4090 9144 4094 9148
rect 3066 9124 3070 9128
rect 2877 9117 2881 9121
rect 2921 9117 2925 9121
rect 2948 9117 2952 9121
rect 2993 9117 2997 9121
rect 3171 9124 3175 9128
rect 3058 9106 3062 9110
rect 2857 9097 2861 9101
rect 2889 9098 2893 9102
rect 2908 9097 2912 9101
rect 2964 9098 2968 9102
rect 2980 9097 2984 9101
rect 3007 9097 3011 9101
rect 3085 9102 3089 9106
rect 3136 9110 3140 9114
rect 4011 9124 4015 9128
rect 3163 9106 3167 9110
rect 3190 9102 3194 9106
rect 3822 9117 3826 9121
rect 3866 9117 3870 9121
rect 3893 9117 3897 9121
rect 3938 9117 3942 9121
rect 4116 9124 4120 9128
rect 4003 9106 4007 9110
rect 3064 9088 3068 9092
rect 3169 9088 3173 9092
rect 3402 9095 3406 9099
rect 2874 9080 2878 9084
rect 2918 9079 2922 9083
rect 2943 9080 2948 9084
rect 2990 9079 2994 9083
rect 3367 9081 3371 9085
rect 3802 9097 3806 9101
rect 3394 9077 3398 9081
rect 3421 9073 3425 9077
rect 3834 9098 3838 9102
rect 3853 9097 3857 9101
rect 3909 9098 3913 9102
rect 3925 9097 3929 9101
rect 3952 9097 3956 9101
rect 4030 9102 4034 9106
rect 4081 9110 4085 9114
rect 4108 9106 4112 9110
rect 4135 9102 4139 9106
rect 4009 9088 4013 9092
rect 4114 9088 4118 9092
rect 3819 9080 3823 9084
rect 3863 9079 3867 9083
rect 3888 9080 3893 9084
rect 3935 9079 3939 9083
rect 3400 9059 3404 9063
rect 2874 9050 2878 9054
rect 2918 9051 2922 9055
rect 2943 9050 2948 9054
rect 2990 9051 2994 9055
rect 3555 9053 3559 9057
rect 3608 9053 3612 9057
rect 3066 9049 3070 9053
rect 3171 9049 3175 9053
rect 3819 9050 3823 9054
rect 3863 9051 3867 9055
rect 3888 9050 3893 9054
rect 3935 9051 3939 9055
rect 4011 9049 4015 9053
rect 4116 9049 4120 9053
rect 2857 9033 2861 9037
rect 2889 9032 2893 9036
rect 2908 9033 2912 9037
rect 2964 9032 2968 9036
rect 2980 9033 2984 9037
rect 3007 9033 3011 9037
rect 3055 9033 3061 9037
rect 3160 9033 3166 9037
rect 3802 9033 3806 9037
rect 3834 9032 3838 9036
rect 3853 9033 3857 9037
rect 3909 9032 3913 9036
rect 3925 9033 3929 9037
rect 3952 9033 3956 9037
rect 4000 9033 4006 9037
rect 4105 9033 4111 9037
rect 2877 9013 2881 9017
rect 2921 9013 2925 9017
rect 2948 9013 2952 9017
rect 2993 9013 2997 9017
rect 3064 9013 3068 9017
rect 3169 9013 3173 9017
rect 3402 9015 3406 9019
rect 3822 9013 3826 9017
rect 3866 9013 3870 9017
rect 3893 9013 3897 9017
rect 3938 9013 3942 9017
rect 4009 9013 4013 9017
rect 4114 9013 4118 9017
rect 3391 8999 3397 9003
rect 3066 8992 3070 8996
rect 2877 8985 2881 8989
rect 2921 8985 2925 8989
rect 2948 8985 2952 8989
rect 2993 8985 2997 8989
rect 3147 8992 3151 8996
rect 3058 8974 3062 8978
rect 2857 8965 2861 8969
rect 2889 8966 2893 8970
rect 2908 8965 2912 8969
rect 2964 8966 2968 8970
rect 2980 8965 2984 8969
rect 3007 8965 3011 8969
rect 3085 8970 3089 8974
rect 3112 8978 3116 8982
rect 3237 8992 3241 8996
rect 3139 8974 3143 8978
rect 3166 8970 3170 8974
rect 3202 8978 3206 8982
rect 4011 8992 4015 8996
rect 3229 8974 3233 8978
rect 3256 8970 3260 8974
rect 3822 8985 3826 8989
rect 3866 8985 3870 8989
rect 3893 8985 3897 8989
rect 3938 8985 3942 8989
rect 3400 8979 3404 8983
rect 4092 8992 4096 8996
rect 4003 8974 4007 8978
rect 3064 8956 3068 8960
rect 3145 8956 3149 8960
rect 3235 8956 3239 8960
rect 3402 8965 3406 8969
rect 2874 8948 2878 8952
rect 2918 8947 2922 8951
rect 2943 8948 2948 8952
rect 3345 8951 3349 8955
rect 2990 8947 2994 8951
rect 3367 8951 3371 8955
rect 3802 8965 3806 8969
rect 3394 8947 3398 8951
rect 3421 8943 3425 8947
rect 3834 8966 3838 8970
rect 3853 8965 3857 8969
rect 3909 8966 3913 8970
rect 3925 8965 3929 8969
rect 3952 8965 3956 8969
rect 4030 8970 4034 8974
rect 4057 8978 4061 8982
rect 4182 8992 4186 8996
rect 4084 8974 4088 8978
rect 4111 8970 4115 8974
rect 4147 8978 4151 8982
rect 4174 8974 4178 8978
rect 4201 8970 4205 8974
rect 4009 8956 4013 8960
rect 4090 8956 4094 8960
rect 4180 8956 4184 8960
rect 3819 8948 3823 8952
rect 3863 8947 3867 8951
rect 3888 8948 3893 8952
rect 3935 8947 3939 8951
rect 3400 8929 3404 8933
rect 2874 8918 2878 8922
rect 2918 8919 2922 8923
rect 3461 8923 3465 8927
rect 3514 8923 3518 8927
rect 2943 8918 2948 8922
rect 2990 8919 2994 8923
rect 3066 8914 3070 8918
rect 3147 8914 3151 8918
rect 3237 8914 3241 8918
rect 3819 8918 3823 8922
rect 3863 8919 3867 8923
rect 2857 8901 2861 8905
rect 2889 8900 2893 8904
rect 2908 8901 2912 8905
rect 2964 8900 2968 8904
rect 2980 8901 2984 8905
rect 3007 8901 3011 8905
rect 3055 8898 3061 8902
rect 3136 8898 3142 8902
rect 3226 8898 3232 8902
rect 3888 8918 3893 8922
rect 3935 8919 3939 8923
rect 4011 8914 4015 8918
rect 4092 8914 4096 8918
rect 4182 8914 4186 8918
rect 3802 8901 3806 8905
rect 3834 8900 3838 8904
rect 3853 8901 3857 8905
rect 3909 8900 3913 8904
rect 3925 8901 3929 8905
rect 3952 8901 3956 8905
rect 4000 8898 4006 8902
rect 2877 8881 2881 8885
rect 2921 8881 2925 8885
rect 2948 8881 2952 8885
rect 2993 8881 2997 8885
rect 3402 8885 3406 8889
rect 4081 8898 4087 8902
rect 4171 8898 4177 8902
rect 3064 8878 3068 8882
rect 3145 8878 3149 8882
rect 3235 8878 3239 8882
rect 3822 8881 3826 8885
rect 3866 8881 3870 8885
rect 3893 8881 3897 8885
rect 3938 8881 3942 8885
rect 4009 8878 4013 8882
rect 4090 8878 4094 8882
rect 4180 8878 4184 8882
rect 3391 8869 3397 8873
rect 3066 8860 3070 8864
rect 2877 8853 2881 8857
rect 2921 8853 2925 8857
rect 2948 8853 2952 8857
rect 2993 8853 2997 8857
rect 3058 8842 3062 8846
rect 2857 8833 2861 8837
rect 2889 8834 2893 8838
rect 2908 8833 2912 8837
rect 2964 8834 2968 8838
rect 2980 8833 2984 8837
rect 3007 8833 3011 8837
rect 3085 8838 3089 8842
rect 3400 8849 3404 8853
rect 4011 8860 4015 8864
rect 3822 8853 3826 8857
rect 3866 8853 3870 8857
rect 3893 8853 3897 8857
rect 3938 8853 3942 8857
rect 4003 8842 4007 8846
rect 3802 8833 3806 8837
rect 3064 8824 3068 8828
rect 3834 8834 3838 8838
rect 3853 8833 3857 8837
rect 3909 8834 3913 8838
rect 3925 8833 3929 8837
rect 3952 8833 3956 8837
rect 4030 8838 4034 8842
rect 4009 8824 4013 8828
rect 2874 8816 2878 8820
rect 2918 8815 2922 8819
rect 2943 8816 2948 8820
rect 2990 8815 2994 8819
rect 3819 8816 3823 8820
rect 3863 8815 3867 8819
rect 3888 8816 3893 8820
rect 3935 8815 3939 8819
rect 2377 8798 2381 8802
rect 2414 8798 2418 8802
rect 2434 8798 2438 8802
rect 2472 8798 2476 8802
rect 2509 8798 2513 8802
rect 2546 8798 2550 8802
rect 2566 8798 2570 8802
rect 2604 8798 2608 8802
rect 2641 8798 2645 8802
rect 2678 8798 2682 8802
rect 2698 8798 2702 8802
rect 2736 8798 2740 8802
rect 3322 8798 3326 8802
rect 3359 8798 3363 8802
rect 3379 8798 3383 8802
rect 3417 8798 3421 8802
rect 3454 8798 3458 8802
rect 3491 8798 3495 8802
rect 3511 8798 3515 8802
rect 3549 8798 3553 8802
rect 3586 8798 3590 8802
rect 3623 8798 3627 8802
rect 3643 8798 3647 8802
rect 3681 8798 3685 8802
rect 2371 8778 2375 8782
rect 2389 8780 2393 8784
rect 2449 8780 2453 8784
rect 2407 8771 2411 8778
rect 2465 8771 2469 8778
rect 2484 8775 2488 8779
rect 2502 8780 2506 8784
rect 2521 8780 2525 8784
rect 2581 8780 2585 8784
rect 2539 8771 2543 8778
rect 2597 8771 2601 8778
rect 2616 8775 2620 8779
rect 2634 8780 2638 8784
rect 2653 8780 2657 8784
rect 2713 8780 2717 8784
rect 2671 8771 2675 8778
rect 2874 8786 2878 8790
rect 2918 8787 2922 8791
rect 2943 8786 2948 8790
rect 2990 8787 2994 8791
rect 3135 8786 3139 8790
rect 3179 8787 3183 8791
rect 3204 8786 3209 8790
rect 3251 8787 3255 8791
rect 2729 8771 2733 8778
rect 2750 8775 2754 8779
rect 3066 8778 3070 8782
rect 3316 8778 3320 8782
rect 3334 8780 3338 8784
rect 2857 8769 2861 8773
rect 2889 8768 2893 8772
rect 2908 8769 2912 8773
rect 2964 8768 2968 8772
rect 2980 8769 2984 8773
rect 3007 8769 3011 8773
rect 2377 8757 2381 8761
rect 2414 8755 2418 8759
rect 2434 8755 2438 8759
rect 2470 8755 2474 8759
rect 2509 8757 2513 8761
rect 2546 8755 2550 8759
rect 2566 8755 2570 8759
rect 2602 8755 2606 8759
rect 2641 8757 2645 8761
rect 2678 8755 2682 8759
rect 2698 8755 2702 8759
rect 2734 8755 2738 8759
rect 3055 8762 3061 8766
rect 3093 8769 3097 8773
rect 3150 8768 3154 8772
rect 3169 8769 3173 8773
rect 3225 8768 3229 8772
rect 3241 8769 3245 8773
rect 3268 8769 3272 8773
rect 3394 8780 3398 8784
rect 3352 8771 3356 8778
rect 3410 8771 3414 8778
rect 3429 8775 3433 8779
rect 3447 8780 3451 8784
rect 3466 8780 3470 8784
rect 3526 8780 3530 8784
rect 3484 8771 3488 8778
rect 3542 8771 3546 8778
rect 3561 8775 3565 8779
rect 3579 8780 3583 8784
rect 3598 8780 3602 8784
rect 3658 8780 3662 8784
rect 3616 8771 3620 8778
rect 3819 8786 3823 8790
rect 3863 8787 3867 8791
rect 3888 8786 3893 8790
rect 3935 8787 3939 8791
rect 4080 8786 4084 8790
rect 4124 8787 4128 8791
rect 4149 8786 4154 8790
rect 4196 8787 4200 8791
rect 3674 8771 3678 8778
rect 3695 8775 3699 8779
rect 4011 8778 4015 8782
rect 3802 8769 3806 8773
rect 3834 8768 3838 8772
rect 3853 8769 3857 8773
rect 3909 8768 3913 8772
rect 3925 8769 3929 8773
rect 3952 8769 3956 8773
rect 2877 8749 2881 8753
rect 2921 8749 2925 8753
rect 2948 8749 2952 8753
rect 2993 8749 2997 8753
rect 3322 8757 3326 8761
rect 3064 8742 3068 8746
rect 2486 8727 2490 8731
rect 2510 8727 2514 8731
rect 3359 8755 3363 8759
rect 3379 8755 3383 8759
rect 3415 8755 3419 8759
rect 3454 8757 3458 8761
rect 3491 8755 3495 8759
rect 3511 8755 3515 8759
rect 3547 8755 3551 8759
rect 3586 8757 3590 8761
rect 3623 8755 3627 8759
rect 3643 8755 3647 8759
rect 3679 8755 3683 8759
rect 4000 8762 4006 8766
rect 4038 8769 4042 8773
rect 4095 8768 4099 8772
rect 4114 8769 4118 8773
rect 4170 8768 4174 8772
rect 4186 8769 4190 8773
rect 4213 8769 4217 8773
rect 3138 8749 3142 8753
rect 3182 8749 3186 8753
rect 3209 8749 3213 8753
rect 3254 8749 3258 8753
rect 3822 8749 3826 8753
rect 3866 8749 3870 8753
rect 3893 8749 3897 8753
rect 3938 8749 3942 8753
rect 4009 8742 4013 8746
rect 3431 8727 3435 8731
rect 3455 8727 3459 8731
rect 3277 8721 3281 8725
rect 3115 8714 3119 8718
rect 4083 8749 4087 8753
rect 4127 8749 4131 8753
rect 4154 8749 4158 8753
rect 4199 8749 4203 8753
rect 4222 8721 4226 8725
rect 4058 8714 4062 8718
rect 2506 8700 2510 8704
rect 3451 8700 3455 8704
rect 2521 8692 2525 8696
rect 3466 8692 3470 8696
rect 3160 8686 3164 8690
rect 3197 8686 3201 8690
rect 3217 8686 3221 8690
rect 3255 8686 3259 8690
rect 4105 8686 4109 8690
rect 4142 8686 4146 8690
rect 4162 8686 4166 8690
rect 4200 8686 4204 8690
rect 2486 8677 2490 8681
rect 2510 8677 2514 8681
rect 3431 8677 3435 8681
rect 3455 8677 3459 8681
rect 3154 8666 3158 8670
rect 3172 8668 3176 8672
rect 2377 8656 2381 8660
rect 2414 8656 2418 8660
rect 2434 8656 2438 8660
rect 2472 8656 2476 8660
rect 2509 8656 2513 8660
rect 2546 8656 2550 8660
rect 2566 8656 2570 8660
rect 2604 8656 2608 8660
rect 2641 8656 2645 8660
rect 2678 8656 2682 8660
rect 2698 8656 2702 8660
rect 2736 8656 2740 8660
rect 3232 8668 3236 8672
rect 3190 8659 3194 8666
rect 3248 8659 3252 8666
rect 3267 8663 3271 8667
rect 4099 8666 4103 8670
rect 4117 8668 4121 8672
rect 3322 8656 3326 8660
rect 3359 8656 3363 8660
rect 3379 8656 3383 8660
rect 3417 8656 3421 8660
rect 3454 8656 3458 8660
rect 3491 8656 3495 8660
rect 3511 8656 3515 8660
rect 3549 8656 3553 8660
rect 3586 8656 3590 8660
rect 3623 8656 3627 8660
rect 3643 8656 3647 8660
rect 3681 8656 3685 8660
rect 4177 8668 4181 8672
rect 4135 8659 4139 8666
rect 4193 8659 4197 8666
rect 4212 8663 4216 8667
rect 3160 8645 3164 8649
rect 2371 8636 2375 8640
rect 2389 8638 2393 8642
rect 2449 8638 2453 8642
rect 2407 8629 2411 8636
rect 2465 8629 2469 8636
rect 2484 8633 2488 8637
rect 2502 8638 2506 8642
rect 2521 8638 2525 8642
rect 2581 8638 2585 8642
rect 2539 8629 2543 8636
rect 2597 8629 2601 8636
rect 2616 8633 2620 8637
rect 2634 8638 2638 8642
rect 2653 8638 2657 8642
rect 2713 8638 2717 8642
rect 2671 8629 2675 8636
rect 3197 8643 3201 8647
rect 3217 8643 3221 8647
rect 3253 8643 3257 8647
rect 4105 8645 4109 8649
rect 2729 8629 2733 8636
rect 2750 8633 2754 8637
rect 3316 8636 3320 8640
rect 3334 8638 3338 8642
rect 3394 8638 3398 8642
rect 3352 8629 3356 8636
rect 3410 8629 3414 8636
rect 3429 8633 3433 8637
rect 3447 8638 3451 8642
rect 3466 8638 3470 8642
rect 3526 8638 3530 8642
rect 3484 8629 3488 8636
rect 3542 8629 3546 8636
rect 3561 8633 3565 8637
rect 3579 8638 3583 8642
rect 3598 8638 3602 8642
rect 3658 8638 3662 8642
rect 3616 8629 3620 8636
rect 4142 8643 4146 8647
rect 4162 8643 4166 8647
rect 4198 8643 4202 8647
rect 3674 8629 3678 8636
rect 3695 8633 3699 8637
rect 2377 8615 2381 8619
rect 2414 8613 2418 8617
rect 2434 8613 2438 8617
rect 2470 8613 2474 8617
rect 2509 8615 2513 8619
rect 2546 8613 2550 8617
rect 2566 8613 2570 8617
rect 2602 8613 2606 8617
rect 2641 8615 2645 8619
rect 2678 8613 2682 8617
rect 2698 8613 2702 8617
rect 2734 8613 2738 8617
rect 3322 8615 3326 8619
rect 3359 8613 3363 8617
rect 3379 8613 3383 8617
rect 3415 8613 3419 8617
rect 3454 8615 3458 8619
rect 3491 8613 3495 8617
rect 3511 8613 3515 8617
rect 3547 8613 3551 8617
rect 3586 8615 3590 8619
rect 3623 8613 3627 8617
rect 3643 8613 3647 8617
rect 3679 8613 3683 8617
rect 3160 8600 3164 8604
rect 3197 8600 3201 8604
rect 3217 8600 3221 8604
rect 3255 8600 3259 8604
rect 4105 8600 4109 8604
rect 4142 8600 4146 8604
rect 4162 8600 4166 8604
rect 4200 8600 4204 8604
rect 3154 8580 3158 8584
rect 3172 8582 3176 8586
rect 2377 8570 2381 8574
rect 2414 8570 2418 8574
rect 2434 8570 2438 8574
rect 2472 8570 2476 8574
rect 2509 8570 2513 8574
rect 2546 8570 2550 8574
rect 2566 8570 2570 8574
rect 2604 8570 2608 8574
rect 2641 8570 2645 8574
rect 2678 8570 2682 8574
rect 2698 8570 2702 8574
rect 2736 8570 2740 8574
rect 3232 8582 3236 8586
rect 3190 8573 3194 8580
rect 3248 8573 3252 8580
rect 3267 8577 3271 8581
rect 3289 8575 3293 8579
rect 4099 8580 4103 8584
rect 4117 8582 4121 8586
rect 3322 8570 3326 8574
rect 3359 8570 3363 8574
rect 3379 8570 3383 8574
rect 3417 8570 3421 8574
rect 3454 8570 3458 8574
rect 3491 8570 3495 8574
rect 3511 8570 3515 8574
rect 3549 8570 3553 8574
rect 3586 8570 3590 8574
rect 3623 8570 3627 8574
rect 3643 8570 3647 8574
rect 3681 8570 3685 8574
rect 4177 8582 4181 8586
rect 4135 8573 4139 8580
rect 4193 8573 4197 8580
rect 4212 8577 4216 8581
rect 4234 8575 4238 8579
rect 3160 8559 3164 8563
rect 2371 8550 2375 8554
rect 2389 8552 2393 8556
rect 2449 8552 2453 8556
rect 2407 8543 2411 8550
rect 2465 8543 2469 8550
rect 2484 8547 2488 8551
rect 2502 8552 2506 8556
rect 2521 8552 2525 8556
rect 2581 8552 2585 8556
rect 2539 8543 2543 8550
rect 2597 8543 2601 8550
rect 2616 8547 2620 8551
rect 2634 8552 2638 8556
rect 2653 8552 2657 8556
rect 2713 8552 2717 8556
rect 2671 8543 2675 8550
rect 3197 8557 3201 8561
rect 3217 8557 3221 8561
rect 3253 8557 3257 8561
rect 4105 8559 4109 8563
rect 2729 8543 2733 8550
rect 2750 8547 2754 8551
rect 3316 8550 3320 8554
rect 3334 8552 3338 8556
rect 3394 8552 3398 8556
rect 3352 8543 3356 8550
rect 3410 8543 3414 8550
rect 3429 8547 3433 8551
rect 3447 8552 3451 8556
rect 3466 8552 3470 8556
rect 3526 8552 3530 8556
rect 3484 8543 3488 8550
rect 3542 8543 3546 8550
rect 3561 8547 3565 8551
rect 3579 8552 3583 8556
rect 3598 8552 3602 8556
rect 3658 8552 3662 8556
rect 3616 8543 3620 8550
rect 4142 8557 4146 8561
rect 4162 8557 4166 8561
rect 4198 8557 4202 8561
rect 3674 8543 3678 8550
rect 3695 8547 3699 8551
rect 2377 8529 2381 8533
rect 2414 8527 2418 8531
rect 2434 8527 2438 8531
rect 2470 8527 2474 8531
rect 2509 8529 2513 8533
rect 2546 8527 2550 8531
rect 2566 8527 2570 8531
rect 2602 8527 2606 8531
rect 2641 8529 2645 8533
rect 2678 8527 2682 8531
rect 2698 8527 2702 8531
rect 2734 8527 2738 8531
rect 3322 8529 3326 8533
rect 3359 8527 3363 8531
rect 3379 8527 3383 8531
rect 3415 8527 3419 8531
rect 3454 8529 3458 8533
rect 3491 8527 3495 8531
rect 3511 8527 3515 8531
rect 3547 8527 3551 8531
rect 3586 8529 3590 8533
rect 3623 8527 3627 8531
rect 3643 8527 3647 8531
rect 3679 8527 3683 8531
rect 2603 8499 2607 8503
rect 2627 8499 2631 8503
rect 3548 8499 3552 8503
rect 3572 8499 3576 8503
rect 2623 8474 2627 8478
rect 3568 8474 3572 8478
rect 2638 8466 2642 8470
rect 3583 8466 3587 8470
rect 2603 8451 2607 8455
rect 2627 8451 2631 8455
rect 3548 8451 3552 8455
rect 3572 8451 3576 8455
rect 2377 8430 2381 8434
rect 2414 8430 2418 8434
rect 2434 8430 2438 8434
rect 2472 8430 2476 8434
rect 2509 8430 2513 8434
rect 2546 8430 2550 8434
rect 2566 8430 2570 8434
rect 2604 8430 2608 8434
rect 2641 8430 2645 8434
rect 2678 8430 2682 8434
rect 2698 8430 2702 8434
rect 2736 8430 2740 8434
rect 3322 8430 3326 8434
rect 3359 8430 3363 8434
rect 3379 8430 3383 8434
rect 3417 8430 3421 8434
rect 3454 8430 3458 8434
rect 3491 8430 3495 8434
rect 3511 8430 3515 8434
rect 3549 8430 3553 8434
rect 3586 8430 3590 8434
rect 3623 8430 3627 8434
rect 3643 8430 3647 8434
rect 3681 8430 3685 8434
rect 2371 8410 2375 8414
rect 2389 8412 2393 8416
rect 2449 8412 2453 8416
rect 2407 8403 2411 8410
rect 2465 8403 2469 8410
rect 2484 8407 2488 8411
rect 2502 8412 2506 8416
rect 2521 8412 2525 8416
rect 2581 8412 2585 8416
rect 2539 8403 2543 8410
rect 2597 8403 2601 8410
rect 2616 8407 2620 8411
rect 2634 8412 2638 8416
rect 2653 8412 2657 8416
rect 2713 8412 2717 8416
rect 2671 8403 2675 8410
rect 2729 8403 2733 8410
rect 2750 8407 2754 8411
rect 3316 8410 3320 8414
rect 3334 8412 3338 8416
rect 3394 8412 3398 8416
rect 3352 8403 3356 8410
rect 3410 8403 3414 8410
rect 3429 8407 3433 8411
rect 3447 8412 3451 8416
rect 3466 8412 3470 8416
rect 3526 8412 3530 8416
rect 3484 8403 3488 8410
rect 3542 8403 3546 8410
rect 3561 8407 3565 8411
rect 3579 8412 3583 8416
rect 3598 8412 3602 8416
rect 3658 8412 3662 8416
rect 3616 8403 3620 8410
rect 3674 8403 3678 8410
rect 3695 8407 3699 8411
rect 2377 8389 2381 8393
rect 2414 8387 2418 8391
rect 2434 8387 2438 8391
rect 2470 8387 2474 8391
rect 2509 8389 2513 8393
rect 2546 8387 2550 8391
rect 2566 8387 2570 8391
rect 2602 8387 2606 8391
rect 2641 8389 2645 8393
rect 2678 8387 2682 8391
rect 2698 8387 2702 8391
rect 2734 8387 2738 8391
rect 3322 8389 3326 8393
rect 3359 8387 3363 8391
rect 3379 8387 3383 8391
rect 3415 8387 3419 8391
rect 3454 8389 3458 8393
rect 3491 8387 3495 8391
rect 3511 8387 3515 8391
rect 3547 8387 3551 8391
rect 3586 8389 3590 8393
rect 3623 8387 3627 8391
rect 3643 8387 3647 8391
rect 3679 8387 3683 8391
rect 2861 8351 2865 8355
rect 2898 8351 2902 8355
rect 2918 8351 2922 8355
rect 2956 8351 2960 8355
rect 2993 8351 2997 8355
rect 3030 8351 3034 8355
rect 3050 8351 3054 8355
rect 3088 8351 3092 8355
rect 3125 8351 3129 8355
rect 3162 8351 3166 8355
rect 3182 8351 3186 8355
rect 3220 8351 3224 8355
rect 3257 8351 3261 8355
rect 3294 8351 3298 8355
rect 3314 8351 3318 8355
rect 3352 8351 3356 8355
rect 3806 8351 3810 8355
rect 3843 8351 3847 8355
rect 3863 8351 3867 8355
rect 3901 8351 3905 8355
rect 3938 8351 3942 8355
rect 3975 8351 3979 8355
rect 3995 8351 3999 8355
rect 4033 8351 4037 8355
rect 4070 8351 4074 8355
rect 4107 8351 4111 8355
rect 4127 8351 4131 8355
rect 4165 8351 4169 8355
rect 4202 8351 4206 8355
rect 4239 8351 4243 8355
rect 4259 8351 4263 8355
rect 4297 8351 4301 8355
rect 2855 8331 2859 8335
rect 2873 8333 2877 8337
rect 2509 8318 2513 8322
rect 2546 8318 2550 8322
rect 2566 8318 2570 8322
rect 2604 8318 2608 8322
rect 2933 8333 2937 8337
rect 2891 8324 2895 8331
rect 2949 8324 2953 8331
rect 2970 8328 2974 8332
rect 2987 8331 2991 8335
rect 3005 8333 3009 8337
rect 3065 8333 3069 8337
rect 3023 8324 3027 8331
rect 3081 8324 3085 8331
rect 3102 8328 3106 8332
rect 3119 8331 3123 8335
rect 3137 8333 3141 8337
rect 3197 8333 3201 8337
rect 3155 8324 3159 8331
rect 3213 8324 3217 8331
rect 3234 8328 3238 8332
rect 3251 8331 3255 8335
rect 3269 8333 3273 8337
rect 3329 8333 3333 8337
rect 3287 8324 3291 8331
rect 3345 8324 3349 8331
rect 3366 8328 3370 8332
rect 3800 8331 3804 8335
rect 3818 8333 3822 8337
rect 3454 8318 3458 8322
rect 3491 8318 3495 8322
rect 3511 8318 3515 8322
rect 3549 8318 3553 8322
rect 3878 8333 3882 8337
rect 3836 8324 3840 8331
rect 3894 8324 3898 8331
rect 3915 8328 3919 8332
rect 3932 8331 3936 8335
rect 3950 8333 3954 8337
rect 4010 8333 4014 8337
rect 3968 8324 3972 8331
rect 4026 8324 4030 8331
rect 4047 8328 4051 8332
rect 4064 8331 4068 8335
rect 4082 8333 4086 8337
rect 4142 8333 4146 8337
rect 4100 8324 4104 8331
rect 4158 8324 4162 8331
rect 4179 8328 4183 8332
rect 4196 8331 4200 8335
rect 4214 8333 4218 8337
rect 4274 8333 4278 8337
rect 4232 8324 4236 8331
rect 4290 8324 4294 8331
rect 4311 8328 4315 8332
rect 2861 8310 2865 8314
rect 2898 8308 2902 8312
rect 2918 8308 2922 8312
rect 2954 8308 2958 8312
rect 2993 8310 2997 8314
rect 3030 8308 3034 8312
rect 3050 8308 3054 8312
rect 3086 8308 3090 8312
rect 3125 8310 3129 8314
rect 3162 8308 3166 8312
rect 3182 8308 3186 8312
rect 3218 8308 3222 8312
rect 3257 8310 3261 8314
rect 3294 8308 3298 8312
rect 3314 8308 3318 8312
rect 3350 8308 3354 8312
rect 3806 8310 3810 8314
rect 3843 8308 3847 8312
rect 3863 8308 3867 8312
rect 3899 8308 3903 8312
rect 3938 8310 3942 8314
rect 3975 8308 3979 8312
rect 3995 8308 3999 8312
rect 4031 8308 4035 8312
rect 4070 8310 4074 8314
rect 4107 8308 4111 8312
rect 4127 8308 4131 8312
rect 4163 8308 4167 8312
rect 4202 8310 4206 8314
rect 4239 8308 4243 8312
rect 4259 8308 4263 8312
rect 4295 8308 4299 8312
rect 2503 8298 2507 8302
rect 2521 8300 2525 8304
rect 2581 8300 2585 8304
rect 2539 8291 2543 8298
rect 2597 8291 2601 8298
rect 2616 8295 2620 8299
rect 3448 8298 3452 8302
rect 3466 8300 3470 8304
rect 3526 8300 3530 8304
rect 3484 8291 3488 8298
rect 3542 8291 3546 8298
rect 3561 8295 3565 8299
rect 2509 8277 2513 8281
rect 2546 8275 2550 8279
rect 2566 8275 2570 8279
rect 2602 8275 2606 8279
rect 2877 8267 2881 8271
rect 2921 8267 2925 8271
rect 2948 8267 2952 8271
rect 2993 8267 2997 8271
rect 3066 8274 3070 8278
rect 2627 8254 2631 8258
rect 3031 8260 3035 8264
rect 2510 8245 2514 8249
rect 2857 8247 2861 8251
rect 2889 8248 2893 8252
rect 2908 8247 2912 8251
rect 2964 8248 2968 8252
rect 2980 8247 2984 8251
rect 3007 8247 3011 8251
rect 3147 8274 3151 8278
rect 3454 8277 3458 8281
rect 3058 8256 3062 8260
rect 3085 8252 3089 8256
rect 3112 8260 3116 8264
rect 3491 8275 3495 8279
rect 3511 8275 3515 8279
rect 3547 8275 3551 8279
rect 3139 8256 3143 8260
rect 3166 8252 3170 8256
rect 3822 8267 3826 8271
rect 3866 8267 3870 8271
rect 3893 8267 3897 8271
rect 3938 8267 3942 8271
rect 4011 8274 4015 8278
rect 3572 8254 3576 8258
rect 3976 8260 3980 8264
rect 3064 8238 3068 8242
rect 3455 8245 3459 8249
rect 3802 8247 3806 8251
rect 3145 8238 3149 8242
rect 3834 8248 3838 8252
rect 3853 8247 3857 8251
rect 3909 8248 3913 8252
rect 3925 8247 3929 8251
rect 3952 8247 3956 8251
rect 4092 8274 4096 8278
rect 4003 8256 4007 8260
rect 4030 8252 4034 8256
rect 4057 8260 4061 8264
rect 4084 8256 4088 8260
rect 4111 8252 4115 8256
rect 4009 8238 4013 8242
rect 4090 8238 4094 8242
rect 2874 8230 2878 8234
rect 2918 8229 2922 8233
rect 2943 8230 2948 8234
rect 2990 8229 2994 8233
rect 3819 8230 3823 8234
rect 3863 8229 3867 8233
rect 3888 8230 3893 8234
rect 3935 8229 3939 8233
rect 2509 8216 2513 8220
rect 2547 8216 2551 8220
rect 2567 8216 2571 8220
rect 2604 8216 2608 8220
rect 3454 8216 3458 8220
rect 3492 8216 3496 8220
rect 3512 8216 3516 8220
rect 3549 8216 3553 8220
rect 2497 8193 2501 8197
rect 2532 8198 2536 8202
rect 2516 8189 2520 8196
rect 2574 8189 2578 8196
rect 2592 8198 2596 8202
rect 2874 8200 2878 8204
rect 2918 8201 2922 8205
rect 2610 8196 2614 8200
rect 2943 8200 2948 8204
rect 2990 8201 2994 8205
rect 3066 8198 3070 8202
rect 3147 8198 3151 8202
rect 2857 8183 2861 8187
rect 2511 8173 2515 8177
rect 2547 8173 2551 8177
rect 2567 8173 2571 8177
rect 2604 8175 2608 8179
rect 2889 8182 2893 8186
rect 2908 8183 2912 8187
rect 2964 8182 2968 8186
rect 2980 8183 2984 8187
rect 3007 8183 3011 8187
rect 3055 8182 3061 8186
rect 3136 8182 3142 8186
rect 3442 8193 3446 8197
rect 3477 8198 3481 8202
rect 3461 8189 3465 8196
rect 3519 8189 3523 8196
rect 3537 8198 3541 8202
rect 3819 8200 3823 8204
rect 3863 8201 3867 8205
rect 3555 8196 3559 8200
rect 3888 8200 3893 8204
rect 3935 8201 3939 8205
rect 4011 8198 4015 8202
rect 4092 8198 4096 8202
rect 3802 8183 3806 8187
rect 3456 8173 3460 8177
rect 3492 8173 3496 8177
rect 3512 8173 3516 8177
rect 3549 8175 3553 8179
rect 3834 8182 3838 8186
rect 3853 8183 3857 8187
rect 3909 8182 3913 8186
rect 3925 8183 3929 8187
rect 3952 8183 3956 8187
rect 4000 8182 4006 8186
rect 4081 8182 4087 8186
rect 2877 8163 2881 8167
rect 2921 8163 2925 8167
rect 2948 8163 2952 8167
rect 2993 8163 2997 8167
rect 3064 8162 3068 8166
rect 3145 8162 3149 8166
rect 3822 8163 3826 8167
rect 3866 8163 3870 8167
rect 3893 8163 3897 8167
rect 3938 8163 3942 8167
rect 4009 8162 4013 8166
rect 4090 8162 4094 8166
rect 3066 8142 3070 8146
rect 2877 8135 2881 8139
rect 2921 8135 2925 8139
rect 2948 8135 2952 8139
rect 2993 8135 2997 8139
rect 3171 8142 3175 8146
rect 3058 8124 3062 8128
rect 2857 8115 2861 8119
rect 2889 8116 2893 8120
rect 2908 8115 2912 8119
rect 2964 8116 2968 8120
rect 2980 8115 2984 8119
rect 3007 8115 3011 8119
rect 3085 8120 3089 8124
rect 3136 8128 3140 8132
rect 4011 8142 4015 8146
rect 3163 8124 3167 8128
rect 3190 8120 3194 8124
rect 3822 8135 3826 8139
rect 3866 8135 3870 8139
rect 3893 8135 3897 8139
rect 3938 8135 3942 8139
rect 4116 8142 4120 8146
rect 4003 8124 4007 8128
rect 3802 8115 3806 8119
rect 3064 8106 3068 8110
rect 3169 8106 3173 8110
rect 3834 8116 3838 8120
rect 3853 8115 3857 8119
rect 3909 8116 3913 8120
rect 3925 8115 3929 8119
rect 3952 8115 3956 8119
rect 4030 8120 4034 8124
rect 4081 8128 4085 8132
rect 4108 8124 4112 8128
rect 4135 8120 4139 8124
rect 4009 8106 4013 8110
rect 4114 8106 4118 8110
rect 2874 8098 2878 8102
rect 2918 8097 2922 8101
rect 2943 8098 2948 8102
rect 2990 8097 2994 8101
rect 3819 8098 3823 8102
rect 3863 8097 3867 8101
rect 3888 8098 3893 8102
rect 3935 8097 3939 8101
rect 2874 8068 2878 8072
rect 2918 8069 2922 8073
rect 2943 8068 2948 8072
rect 2990 8069 2994 8073
rect 3066 8067 3070 8071
rect 3171 8067 3175 8071
rect 3819 8068 3823 8072
rect 3863 8069 3867 8073
rect 3888 8068 3893 8072
rect 3935 8069 3939 8073
rect 4011 8067 4015 8071
rect 4116 8067 4120 8071
rect 2857 8051 2861 8055
rect 2889 8050 2893 8054
rect 2908 8051 2912 8055
rect 2964 8050 2968 8054
rect 2980 8051 2984 8055
rect 3007 8051 3011 8055
rect 3055 8051 3061 8055
rect 3160 8051 3166 8055
rect 3802 8051 3806 8055
rect 3834 8050 3838 8054
rect 3853 8051 3857 8055
rect 3909 8050 3913 8054
rect 3925 8051 3929 8055
rect 3952 8051 3956 8055
rect 4000 8051 4006 8055
rect 4105 8051 4111 8055
rect 2877 8031 2881 8035
rect 2921 8031 2925 8035
rect 2948 8031 2952 8035
rect 2993 8031 2997 8035
rect 3064 8031 3068 8035
rect 3169 8031 3173 8035
rect 3822 8031 3826 8035
rect 3866 8031 3870 8035
rect 3893 8031 3897 8035
rect 3938 8031 3942 8035
rect 4009 8031 4013 8035
rect 4114 8031 4118 8035
rect 3066 8010 3070 8014
rect 2877 8003 2881 8007
rect 2921 8003 2925 8007
rect 2948 8003 2952 8007
rect 2993 8003 2997 8007
rect 3147 8010 3151 8014
rect 3058 7992 3062 7996
rect 2857 7983 2861 7987
rect 2889 7984 2893 7988
rect 2908 7983 2912 7987
rect 2964 7984 2968 7988
rect 2980 7983 2984 7987
rect 3007 7983 3011 7987
rect 3085 7988 3089 7992
rect 3112 7996 3116 8000
rect 3237 8010 3241 8014
rect 3139 7992 3143 7996
rect 3166 7988 3170 7992
rect 3202 7996 3206 8000
rect 4011 8010 4015 8014
rect 3229 7992 3233 7996
rect 3256 7988 3260 7992
rect 3822 8003 3826 8007
rect 3866 8003 3870 8007
rect 3893 8003 3897 8007
rect 3938 8003 3942 8007
rect 4092 8010 4096 8014
rect 4003 7992 4007 7996
rect 3802 7983 3806 7987
rect 3064 7974 3068 7978
rect 3145 7974 3149 7978
rect 3235 7974 3239 7978
rect 3834 7984 3838 7988
rect 3853 7983 3857 7987
rect 3909 7984 3913 7988
rect 3925 7983 3929 7987
rect 3952 7983 3956 7987
rect 4030 7988 4034 7992
rect 4057 7996 4061 8000
rect 4182 8010 4186 8014
rect 4084 7992 4088 7996
rect 4111 7988 4115 7992
rect 4147 7996 4151 8000
rect 4174 7992 4178 7996
rect 4201 7988 4205 7992
rect 4009 7974 4013 7978
rect 4090 7974 4094 7978
rect 4180 7974 4184 7978
rect 2874 7966 2878 7970
rect 2918 7965 2922 7969
rect 2943 7966 2948 7970
rect 2990 7965 2994 7969
rect 3819 7966 3823 7970
rect 3863 7965 3867 7969
rect 3888 7966 3893 7970
rect 3935 7965 3939 7969
rect 2874 7936 2878 7940
rect 2918 7937 2922 7941
rect 2943 7936 2948 7940
rect 2990 7937 2994 7941
rect 3819 7936 3823 7940
rect 3863 7937 3867 7941
rect 3066 7932 3070 7936
rect 3147 7932 3151 7936
rect 3237 7932 3241 7936
rect 3888 7936 3893 7940
rect 3935 7937 3939 7941
rect 4011 7932 4015 7936
rect 4092 7932 4096 7936
rect 4182 7932 4186 7936
rect 2857 7919 2861 7923
rect 2889 7918 2893 7922
rect 2908 7919 2912 7923
rect 2964 7918 2968 7922
rect 2980 7919 2984 7923
rect 3007 7919 3011 7923
rect 3055 7916 3061 7920
rect 3136 7916 3142 7920
rect 3226 7916 3232 7920
rect 3802 7919 3806 7923
rect 3834 7918 3838 7922
rect 3853 7919 3857 7923
rect 3909 7918 3913 7922
rect 3925 7919 3929 7923
rect 3952 7919 3956 7923
rect 4000 7916 4006 7920
rect 4081 7916 4087 7920
rect 4171 7916 4177 7920
rect 2877 7899 2881 7903
rect 2921 7899 2925 7903
rect 2948 7899 2952 7903
rect 2993 7899 2997 7903
rect 3064 7896 3068 7900
rect 3145 7896 3149 7900
rect 3235 7896 3239 7900
rect 3822 7899 3826 7903
rect 3866 7899 3870 7903
rect 3893 7899 3897 7903
rect 3938 7899 3942 7903
rect 4009 7896 4013 7900
rect 4090 7896 4094 7900
rect 4180 7896 4184 7900
rect 3066 7878 3070 7882
rect 2877 7871 2881 7875
rect 2921 7871 2925 7875
rect 2948 7871 2952 7875
rect 2993 7871 2997 7875
rect 4011 7878 4015 7882
rect 3058 7860 3062 7864
rect 2857 7851 2861 7855
rect 2889 7852 2893 7856
rect 2908 7851 2912 7855
rect 2964 7852 2968 7856
rect 2980 7851 2984 7855
rect 3007 7851 3011 7855
rect 3085 7856 3089 7860
rect 3822 7871 3826 7875
rect 3866 7871 3870 7875
rect 3893 7871 3897 7875
rect 3938 7871 3942 7875
rect 4003 7860 4007 7864
rect 3802 7851 3806 7855
rect 3064 7842 3068 7846
rect 3834 7852 3838 7856
rect 3853 7851 3857 7855
rect 3909 7852 3913 7856
rect 3925 7851 3929 7855
rect 3952 7851 3956 7855
rect 4030 7856 4034 7860
rect 4009 7842 4013 7846
rect 2874 7834 2878 7838
rect 2918 7833 2922 7837
rect 2943 7834 2948 7838
rect 2990 7833 2994 7837
rect 3819 7834 3823 7838
rect 3863 7833 3867 7837
rect 3888 7834 3893 7838
rect 3935 7833 3939 7837
rect 2377 7816 2381 7820
rect 2414 7816 2418 7820
rect 2434 7816 2438 7820
rect 2472 7816 2476 7820
rect 2509 7816 2513 7820
rect 2546 7816 2550 7820
rect 2566 7816 2570 7820
rect 2604 7816 2608 7820
rect 2641 7816 2645 7820
rect 2678 7816 2682 7820
rect 2698 7816 2702 7820
rect 2736 7816 2740 7820
rect 3322 7816 3326 7820
rect 3359 7816 3363 7820
rect 3379 7816 3383 7820
rect 3417 7816 3421 7820
rect 3454 7816 3458 7820
rect 3491 7816 3495 7820
rect 3511 7816 3515 7820
rect 3549 7816 3553 7820
rect 3586 7816 3590 7820
rect 3623 7816 3627 7820
rect 3643 7816 3647 7820
rect 3681 7816 3685 7820
rect 2371 7796 2375 7800
rect 2389 7798 2393 7802
rect 2449 7798 2453 7802
rect 2407 7789 2411 7796
rect 2465 7789 2469 7796
rect 2484 7793 2488 7797
rect 2502 7798 2506 7802
rect 2521 7798 2525 7802
rect 2581 7798 2585 7802
rect 2539 7789 2543 7796
rect 2597 7789 2601 7796
rect 2616 7793 2620 7797
rect 2634 7798 2638 7802
rect 2653 7798 2657 7802
rect 2713 7798 2717 7802
rect 2671 7789 2675 7796
rect 2874 7804 2878 7808
rect 2918 7805 2922 7809
rect 2943 7804 2948 7808
rect 2990 7805 2994 7809
rect 3135 7804 3139 7808
rect 3179 7805 3183 7809
rect 3204 7804 3209 7808
rect 3251 7805 3255 7809
rect 2729 7789 2733 7796
rect 2750 7793 2754 7797
rect 3066 7796 3070 7800
rect 3316 7796 3320 7800
rect 3334 7798 3338 7802
rect 2857 7787 2861 7791
rect 2889 7786 2893 7790
rect 2908 7787 2912 7791
rect 2964 7786 2968 7790
rect 2980 7787 2984 7791
rect 3007 7787 3011 7791
rect 2377 7775 2381 7779
rect 2414 7773 2418 7777
rect 2434 7773 2438 7777
rect 2470 7773 2474 7777
rect 2509 7775 2513 7779
rect 2546 7773 2550 7777
rect 2566 7773 2570 7777
rect 2602 7773 2606 7777
rect 2641 7775 2645 7779
rect 2678 7773 2682 7777
rect 2698 7773 2702 7777
rect 2734 7773 2738 7777
rect 3055 7780 3061 7784
rect 3093 7787 3097 7791
rect 3150 7786 3154 7790
rect 3169 7787 3173 7791
rect 3225 7786 3229 7790
rect 3241 7787 3245 7791
rect 3268 7787 3272 7791
rect 3394 7798 3398 7802
rect 3352 7789 3356 7796
rect 3410 7789 3414 7796
rect 3429 7793 3433 7797
rect 3447 7798 3451 7802
rect 3466 7798 3470 7802
rect 3526 7798 3530 7802
rect 3484 7789 3488 7796
rect 3542 7789 3546 7796
rect 3561 7793 3565 7797
rect 3579 7798 3583 7802
rect 3598 7798 3602 7802
rect 3658 7798 3662 7802
rect 3616 7789 3620 7796
rect 3819 7804 3823 7808
rect 3863 7805 3867 7809
rect 3888 7804 3893 7808
rect 3935 7805 3939 7809
rect 4080 7804 4084 7808
rect 4124 7805 4128 7809
rect 4149 7804 4154 7808
rect 4196 7805 4200 7809
rect 3674 7789 3678 7796
rect 3695 7793 3699 7797
rect 4011 7796 4015 7800
rect 3802 7787 3806 7791
rect 3834 7786 3838 7790
rect 3853 7787 3857 7791
rect 3909 7786 3913 7790
rect 3925 7787 3929 7791
rect 3952 7787 3956 7791
rect 2877 7767 2881 7771
rect 2921 7767 2925 7771
rect 2948 7767 2952 7771
rect 2993 7767 2997 7771
rect 3322 7775 3326 7779
rect 3064 7760 3068 7764
rect 2486 7745 2490 7749
rect 2510 7745 2514 7749
rect 3359 7773 3363 7777
rect 3379 7773 3383 7777
rect 3415 7773 3419 7777
rect 3454 7775 3458 7779
rect 3491 7773 3495 7777
rect 3511 7773 3515 7777
rect 3547 7773 3551 7777
rect 3586 7775 3590 7779
rect 3623 7773 3627 7777
rect 3643 7773 3647 7777
rect 3679 7773 3683 7777
rect 4000 7780 4006 7784
rect 4038 7787 4042 7791
rect 4095 7786 4099 7790
rect 4114 7787 4118 7791
rect 4170 7786 4174 7790
rect 4186 7787 4190 7791
rect 4213 7787 4217 7791
rect 3138 7767 3142 7771
rect 3182 7767 3186 7771
rect 3209 7767 3213 7771
rect 3254 7767 3258 7771
rect 3822 7767 3826 7771
rect 3866 7767 3870 7771
rect 3893 7767 3897 7771
rect 3938 7767 3942 7771
rect 4009 7760 4013 7764
rect 3431 7745 3435 7749
rect 3455 7745 3459 7749
rect 3277 7739 3281 7743
rect 3115 7732 3119 7736
rect 4083 7767 4087 7771
rect 4127 7767 4131 7771
rect 4154 7767 4158 7771
rect 4199 7767 4203 7771
rect 4222 7739 4226 7743
rect 4058 7732 4062 7736
rect 2506 7718 2510 7722
rect 3451 7718 3455 7722
rect 2521 7710 2525 7714
rect 3466 7710 3470 7714
rect 3160 7704 3164 7708
rect 3197 7704 3201 7708
rect 3217 7704 3221 7708
rect 3255 7704 3259 7708
rect 4105 7704 4109 7708
rect 4142 7704 4146 7708
rect 4162 7704 4166 7708
rect 4200 7704 4204 7708
rect 2486 7695 2490 7699
rect 2510 7695 2514 7699
rect 3431 7695 3435 7699
rect 3455 7695 3459 7699
rect 3154 7684 3158 7688
rect 3172 7686 3176 7690
rect 2377 7674 2381 7678
rect 2414 7674 2418 7678
rect 2434 7674 2438 7678
rect 2472 7674 2476 7678
rect 2509 7674 2513 7678
rect 2546 7674 2550 7678
rect 2566 7674 2570 7678
rect 2604 7674 2608 7678
rect 2641 7674 2645 7678
rect 2678 7674 2682 7678
rect 2698 7674 2702 7678
rect 2736 7674 2740 7678
rect 3232 7686 3236 7690
rect 3190 7677 3194 7684
rect 3248 7677 3252 7684
rect 3267 7681 3271 7685
rect 4099 7684 4103 7688
rect 4117 7686 4121 7690
rect 3322 7674 3326 7678
rect 3359 7674 3363 7678
rect 3379 7674 3383 7678
rect 3417 7674 3421 7678
rect 3454 7674 3458 7678
rect 3491 7674 3495 7678
rect 3511 7674 3515 7678
rect 3549 7674 3553 7678
rect 3586 7674 3590 7678
rect 3623 7674 3627 7678
rect 3643 7674 3647 7678
rect 3681 7674 3685 7678
rect 4177 7686 4181 7690
rect 4135 7677 4139 7684
rect 4193 7677 4197 7684
rect 4212 7681 4216 7685
rect 3160 7663 3164 7667
rect 2371 7654 2375 7658
rect 2389 7656 2393 7660
rect 2449 7656 2453 7660
rect 2407 7647 2411 7654
rect 2465 7647 2469 7654
rect 2484 7651 2488 7655
rect 2502 7656 2506 7660
rect 2521 7656 2525 7660
rect 2581 7656 2585 7660
rect 2539 7647 2543 7654
rect 2597 7647 2601 7654
rect 2616 7651 2620 7655
rect 2634 7656 2638 7660
rect 2653 7656 2657 7660
rect 2713 7656 2717 7660
rect 2671 7647 2675 7654
rect 3197 7661 3201 7665
rect 3217 7661 3221 7665
rect 3253 7661 3257 7665
rect 4105 7663 4109 7667
rect 2729 7647 2733 7654
rect 2750 7651 2754 7655
rect 3316 7654 3320 7658
rect 3334 7656 3338 7660
rect 3394 7656 3398 7660
rect 3352 7647 3356 7654
rect 3410 7647 3414 7654
rect 3429 7651 3433 7655
rect 3447 7656 3451 7660
rect 3466 7656 3470 7660
rect 3526 7656 3530 7660
rect 3484 7647 3488 7654
rect 3542 7647 3546 7654
rect 3561 7651 3565 7655
rect 3579 7656 3583 7660
rect 3598 7656 3602 7660
rect 3658 7656 3662 7660
rect 3616 7647 3620 7654
rect 4142 7661 4146 7665
rect 4162 7661 4166 7665
rect 4198 7661 4202 7665
rect 3674 7647 3678 7654
rect 3695 7651 3699 7655
rect 2377 7633 2381 7637
rect 2414 7631 2418 7635
rect 2434 7631 2438 7635
rect 2470 7631 2474 7635
rect 2509 7633 2513 7637
rect 2546 7631 2550 7635
rect 2566 7631 2570 7635
rect 2602 7631 2606 7635
rect 2641 7633 2645 7637
rect 2678 7631 2682 7635
rect 2698 7631 2702 7635
rect 2734 7631 2738 7635
rect 3322 7633 3326 7637
rect 3359 7631 3363 7635
rect 3379 7631 3383 7635
rect 3415 7631 3419 7635
rect 3454 7633 3458 7637
rect 3491 7631 3495 7635
rect 3511 7631 3515 7635
rect 3547 7631 3551 7635
rect 3586 7633 3590 7637
rect 3623 7631 3627 7635
rect 3643 7631 3647 7635
rect 3679 7631 3683 7635
rect 3160 7618 3164 7622
rect 3197 7618 3201 7622
rect 3217 7618 3221 7622
rect 3255 7618 3259 7622
rect 4105 7618 4109 7622
rect 4142 7618 4146 7622
rect 4162 7618 4166 7622
rect 4200 7618 4204 7622
rect 3154 7598 3158 7602
rect 3172 7600 3176 7604
rect 2377 7588 2381 7592
rect 2414 7588 2418 7592
rect 2434 7588 2438 7592
rect 2472 7588 2476 7592
rect 2509 7588 2513 7592
rect 2546 7588 2550 7592
rect 2566 7588 2570 7592
rect 2604 7588 2608 7592
rect 2641 7588 2645 7592
rect 2678 7588 2682 7592
rect 2698 7588 2702 7592
rect 2736 7588 2740 7592
rect 3232 7600 3236 7604
rect 3190 7591 3194 7598
rect 3248 7591 3252 7598
rect 3267 7595 3271 7599
rect 3289 7593 3293 7597
rect 4099 7598 4103 7602
rect 4117 7600 4121 7604
rect 3322 7588 3326 7592
rect 3359 7588 3363 7592
rect 3379 7588 3383 7592
rect 3417 7588 3421 7592
rect 3454 7588 3458 7592
rect 3491 7588 3495 7592
rect 3511 7588 3515 7592
rect 3549 7588 3553 7592
rect 3586 7588 3590 7592
rect 3623 7588 3627 7592
rect 3643 7588 3647 7592
rect 3681 7588 3685 7592
rect 4177 7600 4181 7604
rect 4135 7591 4139 7598
rect 4193 7591 4197 7598
rect 4212 7595 4216 7599
rect 4234 7593 4238 7597
rect 3160 7577 3164 7581
rect 2371 7568 2375 7572
rect 2389 7570 2393 7574
rect 2449 7570 2453 7574
rect 2407 7561 2411 7568
rect 2465 7561 2469 7568
rect 2484 7565 2488 7569
rect 2502 7570 2506 7574
rect 2521 7570 2525 7574
rect 2581 7570 2585 7574
rect 2539 7561 2543 7568
rect 2597 7561 2601 7568
rect 2616 7565 2620 7569
rect 2634 7570 2638 7574
rect 2653 7570 2657 7574
rect 2713 7570 2717 7574
rect 2671 7561 2675 7568
rect 3197 7575 3201 7579
rect 3217 7575 3221 7579
rect 3253 7575 3257 7579
rect 4105 7577 4109 7581
rect 2729 7561 2733 7568
rect 2750 7565 2754 7569
rect 3316 7568 3320 7572
rect 3334 7570 3338 7574
rect 3394 7570 3398 7574
rect 3352 7561 3356 7568
rect 3410 7561 3414 7568
rect 3429 7565 3433 7569
rect 3447 7570 3451 7574
rect 3466 7570 3470 7574
rect 3526 7570 3530 7574
rect 3484 7561 3488 7568
rect 3542 7561 3546 7568
rect 3561 7565 3565 7569
rect 3579 7570 3583 7574
rect 3598 7570 3602 7574
rect 3658 7570 3662 7574
rect 3616 7561 3620 7568
rect 4142 7575 4146 7579
rect 4162 7575 4166 7579
rect 4198 7575 4202 7579
rect 3674 7561 3678 7568
rect 3695 7565 3699 7569
rect 2377 7547 2381 7551
rect 2414 7545 2418 7549
rect 2434 7545 2438 7549
rect 2470 7545 2474 7549
rect 2509 7547 2513 7551
rect 2546 7545 2550 7549
rect 2566 7545 2570 7549
rect 2602 7545 2606 7549
rect 2641 7547 2645 7551
rect 2678 7545 2682 7549
rect 2698 7545 2702 7549
rect 2734 7545 2738 7549
rect 3322 7547 3326 7551
rect 3359 7545 3363 7549
rect 3379 7545 3383 7549
rect 3415 7545 3419 7549
rect 3454 7547 3458 7551
rect 3491 7545 3495 7549
rect 3511 7545 3515 7549
rect 3547 7545 3551 7549
rect 3586 7547 3590 7551
rect 3623 7545 3627 7549
rect 3643 7545 3647 7549
rect 3679 7545 3683 7549
rect 2603 7517 2607 7521
rect 2627 7517 2631 7521
rect 3548 7517 3552 7521
rect 3572 7517 3576 7521
rect 2623 7492 2627 7496
rect 3568 7492 3572 7496
rect 2638 7484 2642 7488
rect 3583 7484 3587 7488
rect 2603 7469 2607 7473
rect 2627 7469 2631 7473
rect 3548 7469 3552 7473
rect 3572 7469 3576 7473
rect 2377 7448 2381 7452
rect 2414 7448 2418 7452
rect 2434 7448 2438 7452
rect 2472 7448 2476 7452
rect 2509 7448 2513 7452
rect 2546 7448 2550 7452
rect 2566 7448 2570 7452
rect 2604 7448 2608 7452
rect 2641 7448 2645 7452
rect 2678 7448 2682 7452
rect 2698 7448 2702 7452
rect 2736 7448 2740 7452
rect 3322 7448 3326 7452
rect 3359 7448 3363 7452
rect 3379 7448 3383 7452
rect 3417 7448 3421 7452
rect 3454 7448 3458 7452
rect 3491 7448 3495 7452
rect 3511 7448 3515 7452
rect 3549 7448 3553 7452
rect 3586 7448 3590 7452
rect 3623 7448 3627 7452
rect 3643 7448 3647 7452
rect 3681 7448 3685 7452
rect 2371 7428 2375 7432
rect 2389 7430 2393 7434
rect 2449 7430 2453 7434
rect 2407 7421 2411 7428
rect 2465 7421 2469 7428
rect 2484 7425 2488 7429
rect 2502 7430 2506 7434
rect 2521 7430 2525 7434
rect 2581 7430 2585 7434
rect 2539 7421 2543 7428
rect 2597 7421 2601 7428
rect 2616 7425 2620 7429
rect 2634 7430 2638 7434
rect 2653 7430 2657 7434
rect 2713 7430 2717 7434
rect 2671 7421 2675 7428
rect 2729 7421 2733 7428
rect 2750 7425 2754 7429
rect 3316 7428 3320 7432
rect 3334 7430 3338 7434
rect 3394 7430 3398 7434
rect 3352 7421 3356 7428
rect 3410 7421 3414 7428
rect 3429 7425 3433 7429
rect 3447 7430 3451 7434
rect 3466 7430 3470 7434
rect 3526 7430 3530 7434
rect 3484 7421 3488 7428
rect 3542 7421 3546 7428
rect 3561 7425 3565 7429
rect 3579 7430 3583 7434
rect 3598 7430 3602 7434
rect 3658 7430 3662 7434
rect 3616 7421 3620 7428
rect 3674 7421 3678 7428
rect 3695 7425 3699 7429
rect 2377 7407 2381 7411
rect 2414 7405 2418 7409
rect 2434 7405 2438 7409
rect 2470 7405 2474 7409
rect 2509 7407 2513 7411
rect 2546 7405 2550 7409
rect 2566 7405 2570 7409
rect 2602 7405 2606 7409
rect 2641 7407 2645 7411
rect 2678 7405 2682 7409
rect 2698 7405 2702 7409
rect 2734 7405 2738 7409
rect 3322 7407 3326 7411
rect 3359 7405 3363 7409
rect 3379 7405 3383 7409
rect 3415 7405 3419 7409
rect 3454 7407 3458 7411
rect 3491 7405 3495 7409
rect 3511 7405 3515 7409
rect 3547 7405 3551 7409
rect 3586 7407 3590 7411
rect 3623 7405 3627 7409
rect 3643 7405 3647 7409
rect 3679 7405 3683 7409
rect 4572 7954 4576 7960
rect 4593 7959 4597 7965
rect 4635 7950 4639 7963
rect 4678 7952 4682 7965
rect 4711 7954 4717 7963
<< metal1 >>
rect 1060 10290 1320 10293
rect 118 9786 1024 10280
rect 1060 10036 1063 10290
rect 1317 10036 1320 10290
rect 1060 10033 1320 10036
rect 1369 10290 1629 10293
rect 1369 10036 1372 10290
rect 1462 10138 1546 10223
rect 1626 10036 1629 10290
rect 1369 10033 1629 10036
rect 1678 10290 1938 10293
rect 1678 10036 1681 10290
rect 1765 10113 1843 10202
rect 1935 10036 1938 10290
rect 1678 10033 1938 10036
rect 1987 10290 2247 10293
rect 1987 10036 1990 10290
rect 2072 10118 2150 10207
rect 2244 10036 2247 10290
rect 1987 10033 2247 10036
rect 2296 10290 2556 10293
rect 2296 10036 2299 10290
rect 2389 10118 2467 10207
rect 2553 10036 2556 10290
rect 2296 10033 2556 10036
rect 2605 10290 2865 10293
rect 2605 10036 2608 10290
rect 2700 10120 2778 10209
rect 2862 10036 2865 10290
rect 2605 10033 2865 10036
rect 2914 10290 3174 10293
rect 2914 10036 2917 10290
rect 3004 10110 3082 10199
rect 3171 10036 3174 10290
rect 2914 10033 3174 10036
rect 3223 10290 3483 10293
rect 3223 10036 3226 10290
rect 3318 10118 3396 10207
rect 3480 10036 3483 10290
rect 3223 10033 3483 10036
rect 3532 10290 3792 10293
rect 3532 10036 3535 10290
rect 3608 10103 3720 10217
rect 3789 10036 3792 10290
rect 3532 10033 3792 10036
rect 3841 10290 4101 10293
rect 3841 10036 3844 10290
rect 4098 10036 4101 10290
rect 3841 10033 4101 10036
rect 1102 10023 1278 10033
rect 1411 10023 1587 10033
rect 1720 10023 1896 10033
rect 2029 10023 2205 10033
rect 2338 10023 2514 10033
rect 2647 10023 2823 10033
rect 2956 10023 3132 10033
rect 3265 10023 3441 10033
rect 3574 10023 3750 10033
rect 3883 10023 4059 10033
rect 1112 10013 1268 10023
rect 1421 10013 1577 10023
rect 1730 10013 1886 10023
rect 2039 10013 2195 10023
rect 2348 10013 2504 10023
rect 2657 10013 2813 10023
rect 2966 10013 3122 10023
rect 3275 10013 3431 10023
rect 3584 10013 3740 10023
rect 3893 10013 4049 10023
rect 1122 10003 1258 10013
rect 1431 10003 1567 10013
rect 1740 10003 1876 10013
rect 2049 10003 2185 10013
rect 2358 10003 2494 10013
rect 2667 10003 2803 10013
rect 2976 10003 3112 10013
rect 3285 10003 3421 10013
rect 3594 10003 3730 10013
rect 3903 10003 4039 10013
rect 1132 9993 1248 10003
rect 1441 10001 1557 10003
rect 1441 9997 1454 10001
rect 1458 9997 1461 10001
rect 1465 9997 1468 10001
rect 1472 9997 1475 10001
rect 1479 9997 1482 10001
rect 1486 9997 1489 10001
rect 1493 9997 1496 10001
rect 1500 9997 1503 10001
rect 1507 9997 1510 10001
rect 1514 9997 1517 10001
rect 1521 9997 1524 10001
rect 1528 9997 1531 10001
rect 1535 9997 1538 10001
rect 1542 9997 1557 10001
rect 1441 9996 1557 9997
rect 1441 9993 1454 9996
rect 118 9348 593 9786
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 802 9761 821 9762
rect 806 9757 807 9761
rect 811 9757 812 9761
rect 816 9757 817 9761
rect 802 9756 821 9757
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 802 9751 821 9752
rect 806 9747 807 9751
rect 811 9747 812 9751
rect 816 9747 817 9751
rect 802 9746 821 9747
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 802 9741 821 9742
rect 806 9737 807 9741
rect 811 9737 812 9741
rect 816 9737 817 9741
rect 802 9736 821 9737
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 831 9761 850 9762
rect 835 9757 836 9761
rect 840 9757 841 9761
rect 845 9757 846 9761
rect 831 9756 850 9757
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 831 9751 850 9752
rect 835 9747 836 9751
rect 840 9747 841 9751
rect 845 9747 846 9751
rect 831 9746 850 9747
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 831 9741 850 9742
rect 835 9737 836 9741
rect 840 9737 841 9741
rect 845 9737 846 9741
rect 831 9736 850 9737
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 860 9761 879 9762
rect 864 9757 865 9761
rect 869 9757 870 9761
rect 874 9757 875 9761
rect 860 9756 879 9757
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 860 9751 879 9752
rect 864 9747 865 9751
rect 869 9747 870 9751
rect 874 9747 875 9751
rect 860 9746 879 9747
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 860 9741 879 9742
rect 864 9737 865 9741
rect 869 9737 870 9741
rect 874 9737 875 9741
rect 860 9736 879 9737
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 889 9761 908 9762
rect 893 9757 894 9761
rect 898 9757 899 9761
rect 903 9757 904 9761
rect 889 9756 908 9757
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 889 9751 908 9752
rect 893 9747 894 9751
rect 898 9747 899 9751
rect 903 9747 904 9751
rect 889 9746 908 9747
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 889 9741 908 9742
rect 893 9737 894 9741
rect 898 9737 899 9741
rect 903 9737 904 9741
rect 889 9736 908 9737
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 918 9761 937 9762
rect 922 9757 923 9761
rect 927 9757 928 9761
rect 932 9757 933 9761
rect 918 9756 937 9757
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 918 9751 937 9752
rect 922 9747 923 9751
rect 927 9747 928 9751
rect 932 9747 933 9751
rect 918 9746 937 9747
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 918 9741 937 9742
rect 922 9737 923 9741
rect 927 9737 928 9741
rect 932 9737 933 9741
rect 918 9736 937 9737
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 802 9715 821 9716
rect 806 9711 807 9715
rect 811 9711 812 9715
rect 816 9711 817 9715
rect 802 9710 821 9711
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 802 9705 821 9706
rect 806 9701 807 9705
rect 811 9701 812 9705
rect 816 9701 817 9705
rect 802 9700 821 9701
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 802 9695 821 9696
rect 806 9691 807 9695
rect 811 9691 812 9695
rect 816 9691 817 9695
rect 802 9690 821 9691
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 831 9715 850 9716
rect 835 9711 836 9715
rect 840 9711 841 9715
rect 845 9711 846 9715
rect 831 9710 850 9711
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 831 9705 850 9706
rect 835 9701 836 9705
rect 840 9701 841 9705
rect 845 9701 846 9705
rect 831 9700 850 9701
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 831 9695 850 9696
rect 835 9691 836 9695
rect 840 9691 841 9695
rect 845 9691 846 9695
rect 831 9690 850 9691
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 860 9715 879 9716
rect 864 9711 865 9715
rect 869 9711 870 9715
rect 874 9711 875 9715
rect 860 9710 879 9711
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 860 9705 879 9706
rect 864 9701 865 9705
rect 869 9701 870 9705
rect 874 9701 875 9705
rect 860 9700 879 9701
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 860 9695 879 9696
rect 864 9691 865 9695
rect 869 9691 870 9695
rect 874 9691 875 9695
rect 860 9690 879 9691
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 889 9715 908 9716
rect 893 9711 894 9715
rect 898 9711 899 9715
rect 903 9711 904 9715
rect 889 9710 908 9711
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 889 9705 908 9706
rect 893 9701 894 9705
rect 898 9701 899 9705
rect 903 9701 904 9705
rect 889 9700 908 9701
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 889 9695 908 9696
rect 893 9691 894 9695
rect 898 9691 899 9695
rect 903 9691 904 9695
rect 889 9690 908 9691
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 918 9715 937 9716
rect 922 9711 923 9715
rect 927 9711 928 9715
rect 932 9711 933 9715
rect 918 9710 937 9711
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 918 9705 937 9706
rect 922 9701 923 9705
rect 927 9701 928 9705
rect 932 9701 933 9705
rect 918 9700 937 9701
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 918 9695 937 9696
rect 922 9691 923 9695
rect 927 9691 928 9695
rect 932 9691 933 9695
rect 918 9690 937 9691
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 617 9618 618 9622
rect 622 9618 623 9622
rect 627 9618 628 9622
rect 632 9618 633 9622
rect 637 9618 638 9622
rect 642 9618 643 9622
rect 613 9617 647 9618
rect 617 9613 618 9617
rect 622 9613 623 9617
rect 627 9613 628 9617
rect 632 9613 633 9617
rect 637 9613 638 9617
rect 642 9613 643 9617
rect 613 9612 647 9613
rect 617 9608 618 9612
rect 622 9608 623 9612
rect 627 9608 628 9612
rect 632 9608 633 9612
rect 637 9608 638 9612
rect 642 9608 643 9612
rect 613 9607 647 9608
rect 617 9603 618 9607
rect 622 9603 623 9607
rect 627 9603 628 9607
rect 632 9603 633 9607
rect 637 9603 638 9607
rect 642 9603 643 9607
rect 663 9618 664 9622
rect 668 9618 669 9622
rect 673 9618 674 9622
rect 678 9618 679 9622
rect 683 9618 684 9622
rect 688 9618 689 9622
rect 659 9617 693 9618
rect 663 9613 664 9617
rect 668 9613 669 9617
rect 673 9613 674 9617
rect 678 9613 679 9617
rect 683 9613 684 9617
rect 688 9613 689 9617
rect 659 9612 693 9613
rect 663 9608 664 9612
rect 668 9608 669 9612
rect 673 9608 674 9612
rect 678 9608 679 9612
rect 683 9608 684 9612
rect 688 9608 689 9612
rect 1142 9610 1238 9993
rect 1451 9992 1454 9993
rect 1458 9992 1461 9996
rect 1465 9992 1468 9996
rect 1472 9992 1475 9996
rect 1479 9992 1482 9996
rect 1486 9992 1489 9996
rect 1493 9992 1496 9996
rect 1500 9992 1503 9996
rect 1507 9992 1510 9996
rect 1514 9992 1517 9996
rect 1521 9992 1524 9996
rect 1528 9992 1531 9996
rect 1535 9992 1538 9996
rect 1542 9993 1557 9996
rect 1750 10001 1866 10003
rect 1750 9997 1763 10001
rect 1767 9997 1770 10001
rect 1774 9997 1777 10001
rect 1781 9997 1784 10001
rect 1788 9997 1791 10001
rect 1795 9997 1798 10001
rect 1802 9997 1805 10001
rect 1809 9997 1812 10001
rect 1816 9997 1819 10001
rect 1823 9997 1826 10001
rect 1830 9997 1833 10001
rect 1837 9997 1840 10001
rect 1844 9997 1847 10001
rect 1851 9997 1866 10001
rect 1750 9996 1866 9997
rect 1750 9993 1763 9996
rect 1542 9992 1547 9993
rect 1451 9991 1547 9992
rect 1451 9987 1454 9991
rect 1458 9987 1461 9991
rect 1465 9987 1468 9991
rect 1472 9987 1475 9991
rect 1479 9987 1482 9991
rect 1486 9987 1489 9991
rect 1493 9987 1496 9991
rect 1500 9987 1503 9991
rect 1507 9987 1510 9991
rect 1514 9987 1517 9991
rect 1521 9987 1524 9991
rect 1528 9987 1531 9991
rect 1535 9987 1538 9991
rect 1542 9987 1547 9991
rect 1451 9986 1547 9987
rect 1451 9982 1454 9986
rect 1458 9982 1461 9986
rect 1465 9982 1468 9986
rect 1472 9982 1475 9986
rect 1479 9982 1482 9986
rect 1486 9982 1489 9986
rect 1493 9982 1496 9986
rect 1500 9982 1503 9986
rect 1507 9982 1510 9986
rect 1514 9982 1517 9986
rect 1521 9982 1524 9986
rect 1528 9982 1531 9986
rect 1535 9982 1538 9986
rect 1542 9982 1547 9986
rect 1451 9981 1547 9982
rect 1760 9992 1763 9993
rect 1767 9992 1770 9996
rect 1774 9992 1777 9996
rect 1781 9992 1784 9996
rect 1788 9992 1791 9996
rect 1795 9992 1798 9996
rect 1802 9992 1805 9996
rect 1809 9992 1812 9996
rect 1816 9992 1819 9996
rect 1823 9992 1826 9996
rect 1830 9992 1833 9996
rect 1837 9992 1840 9996
rect 1844 9992 1847 9996
rect 1851 9993 1866 9996
rect 2059 10001 2175 10003
rect 2059 9997 2072 10001
rect 2076 9997 2079 10001
rect 2083 9997 2086 10001
rect 2090 9997 2093 10001
rect 2097 9997 2100 10001
rect 2104 9997 2107 10001
rect 2111 9997 2114 10001
rect 2118 9997 2121 10001
rect 2125 9997 2128 10001
rect 2132 9997 2135 10001
rect 2139 9997 2142 10001
rect 2146 9997 2149 10001
rect 2153 9997 2156 10001
rect 2160 9997 2175 10001
rect 2059 9996 2175 9997
rect 2059 9993 2072 9996
rect 1851 9992 1856 9993
rect 1760 9991 1856 9992
rect 1760 9987 1763 9991
rect 1767 9987 1770 9991
rect 1774 9987 1777 9991
rect 1781 9987 1784 9991
rect 1788 9987 1791 9991
rect 1795 9987 1798 9991
rect 1802 9987 1805 9991
rect 1809 9987 1812 9991
rect 1816 9987 1819 9991
rect 1823 9987 1826 9991
rect 1830 9987 1833 9991
rect 1837 9987 1840 9991
rect 1844 9987 1847 9991
rect 1851 9987 1856 9991
rect 1760 9986 1856 9987
rect 1760 9982 1763 9986
rect 1767 9982 1770 9986
rect 1774 9982 1777 9986
rect 1781 9982 1784 9986
rect 1788 9982 1791 9986
rect 1795 9982 1798 9986
rect 1802 9982 1805 9986
rect 1809 9982 1812 9986
rect 1816 9982 1819 9986
rect 1823 9982 1826 9986
rect 1830 9982 1833 9986
rect 1837 9982 1840 9986
rect 1844 9982 1847 9986
rect 1851 9982 1856 9986
rect 1760 9981 1856 9982
rect 2069 9992 2072 9993
rect 2076 9992 2079 9996
rect 2083 9992 2086 9996
rect 2090 9992 2093 9996
rect 2097 9992 2100 9996
rect 2104 9992 2107 9996
rect 2111 9992 2114 9996
rect 2118 9992 2121 9996
rect 2125 9992 2128 9996
rect 2132 9992 2135 9996
rect 2139 9992 2142 9996
rect 2146 9992 2149 9996
rect 2153 9992 2156 9996
rect 2160 9993 2175 9996
rect 2368 10001 2484 10003
rect 2368 9997 2381 10001
rect 2385 9997 2388 10001
rect 2392 9997 2395 10001
rect 2399 9997 2402 10001
rect 2406 9997 2409 10001
rect 2413 9997 2416 10001
rect 2420 9997 2423 10001
rect 2427 9997 2430 10001
rect 2434 9997 2437 10001
rect 2441 9997 2444 10001
rect 2448 9997 2451 10001
rect 2455 9997 2458 10001
rect 2462 9997 2465 10001
rect 2469 9997 2484 10001
rect 2368 9996 2484 9997
rect 2368 9993 2381 9996
rect 2160 9992 2165 9993
rect 2069 9991 2165 9992
rect 2069 9987 2072 9991
rect 2076 9987 2079 9991
rect 2083 9987 2086 9991
rect 2090 9987 2093 9991
rect 2097 9987 2100 9991
rect 2104 9987 2107 9991
rect 2111 9987 2114 9991
rect 2118 9987 2121 9991
rect 2125 9987 2128 9991
rect 2132 9987 2135 9991
rect 2139 9987 2142 9991
rect 2146 9987 2149 9991
rect 2153 9987 2156 9991
rect 2160 9987 2165 9991
rect 2069 9986 2165 9987
rect 2069 9982 2072 9986
rect 2076 9982 2079 9986
rect 2083 9982 2086 9986
rect 2090 9982 2093 9986
rect 2097 9982 2100 9986
rect 2104 9982 2107 9986
rect 2111 9982 2114 9986
rect 2118 9982 2121 9986
rect 2125 9982 2128 9986
rect 2132 9982 2135 9986
rect 2139 9982 2142 9986
rect 2146 9982 2149 9986
rect 2153 9982 2156 9986
rect 2160 9982 2165 9986
rect 2069 9981 2165 9982
rect 2378 9992 2381 9993
rect 2385 9992 2388 9996
rect 2392 9992 2395 9996
rect 2399 9992 2402 9996
rect 2406 9992 2409 9996
rect 2413 9992 2416 9996
rect 2420 9992 2423 9996
rect 2427 9992 2430 9996
rect 2434 9992 2437 9996
rect 2441 9992 2444 9996
rect 2448 9992 2451 9996
rect 2455 9992 2458 9996
rect 2462 9992 2465 9996
rect 2469 9993 2484 9996
rect 2677 10001 2793 10003
rect 2677 9997 2690 10001
rect 2694 9997 2697 10001
rect 2701 9997 2704 10001
rect 2708 9997 2711 10001
rect 2715 9997 2718 10001
rect 2722 9997 2725 10001
rect 2729 9997 2732 10001
rect 2736 9997 2739 10001
rect 2743 9997 2746 10001
rect 2750 9997 2753 10001
rect 2757 9997 2760 10001
rect 2764 9997 2767 10001
rect 2771 9997 2774 10001
rect 2778 9997 2793 10001
rect 2677 9996 2793 9997
rect 2677 9993 2690 9996
rect 2469 9992 2474 9993
rect 2378 9991 2474 9992
rect 2378 9987 2381 9991
rect 2385 9987 2388 9991
rect 2392 9987 2395 9991
rect 2399 9987 2402 9991
rect 2406 9987 2409 9991
rect 2413 9987 2416 9991
rect 2420 9987 2423 9991
rect 2427 9987 2430 9991
rect 2434 9987 2437 9991
rect 2441 9987 2444 9991
rect 2448 9987 2451 9991
rect 2455 9987 2458 9991
rect 2462 9987 2465 9991
rect 2469 9987 2474 9991
rect 2378 9986 2474 9987
rect 2378 9982 2381 9986
rect 2385 9982 2388 9986
rect 2392 9982 2395 9986
rect 2399 9982 2402 9986
rect 2406 9982 2409 9986
rect 2413 9982 2416 9986
rect 2420 9982 2423 9986
rect 2427 9982 2430 9986
rect 2434 9982 2437 9986
rect 2441 9982 2444 9986
rect 2448 9982 2451 9986
rect 2455 9982 2458 9986
rect 2462 9982 2465 9986
rect 2469 9982 2474 9986
rect 2378 9981 2474 9982
rect 2687 9992 2690 9993
rect 2694 9992 2697 9996
rect 2701 9992 2704 9996
rect 2708 9992 2711 9996
rect 2715 9992 2718 9996
rect 2722 9992 2725 9996
rect 2729 9992 2732 9996
rect 2736 9992 2739 9996
rect 2743 9992 2746 9996
rect 2750 9992 2753 9996
rect 2757 9992 2760 9996
rect 2764 9992 2767 9996
rect 2771 9992 2774 9996
rect 2778 9993 2793 9996
rect 2986 10001 3102 10003
rect 2986 9997 2999 10001
rect 3003 9997 3006 10001
rect 3010 9997 3013 10001
rect 3017 9997 3020 10001
rect 3024 9997 3027 10001
rect 3031 9997 3034 10001
rect 3038 9997 3041 10001
rect 3045 9997 3048 10001
rect 3052 9997 3055 10001
rect 3059 9997 3062 10001
rect 3066 9997 3069 10001
rect 3073 9997 3076 10001
rect 3080 9997 3083 10001
rect 3087 9997 3102 10001
rect 2986 9996 3102 9997
rect 2986 9993 2999 9996
rect 2778 9992 2783 9993
rect 2687 9991 2783 9992
rect 2687 9987 2690 9991
rect 2694 9987 2697 9991
rect 2701 9987 2704 9991
rect 2708 9987 2711 9991
rect 2715 9987 2718 9991
rect 2722 9987 2725 9991
rect 2729 9987 2732 9991
rect 2736 9987 2739 9991
rect 2743 9987 2746 9991
rect 2750 9987 2753 9991
rect 2757 9987 2760 9991
rect 2764 9987 2767 9991
rect 2771 9987 2774 9991
rect 2778 9987 2783 9991
rect 2687 9986 2783 9987
rect 2687 9982 2690 9986
rect 2694 9982 2697 9986
rect 2701 9982 2704 9986
rect 2708 9982 2711 9986
rect 2715 9982 2718 9986
rect 2722 9982 2725 9986
rect 2729 9982 2732 9986
rect 2736 9982 2739 9986
rect 2743 9982 2746 9986
rect 2750 9982 2753 9986
rect 2757 9982 2760 9986
rect 2764 9982 2767 9986
rect 2771 9982 2774 9986
rect 2778 9982 2783 9986
rect 2687 9981 2783 9982
rect 2996 9992 2999 9993
rect 3003 9992 3006 9996
rect 3010 9992 3013 9996
rect 3017 9992 3020 9996
rect 3024 9992 3027 9996
rect 3031 9992 3034 9996
rect 3038 9992 3041 9996
rect 3045 9992 3048 9996
rect 3052 9992 3055 9996
rect 3059 9992 3062 9996
rect 3066 9992 3069 9996
rect 3073 9992 3076 9996
rect 3080 9992 3083 9996
rect 3087 9993 3102 9996
rect 3295 10001 3411 10003
rect 3295 9997 3308 10001
rect 3312 9997 3315 10001
rect 3319 9997 3322 10001
rect 3326 9997 3329 10001
rect 3333 9997 3336 10001
rect 3340 9997 3343 10001
rect 3347 9997 3350 10001
rect 3354 9997 3357 10001
rect 3361 9997 3364 10001
rect 3368 9997 3371 10001
rect 3375 9997 3378 10001
rect 3382 9997 3385 10001
rect 3389 9997 3392 10001
rect 3396 9997 3411 10001
rect 3295 9996 3411 9997
rect 3295 9993 3308 9996
rect 3087 9992 3092 9993
rect 2996 9991 3092 9992
rect 2996 9987 2999 9991
rect 3003 9987 3006 9991
rect 3010 9987 3013 9991
rect 3017 9987 3020 9991
rect 3024 9987 3027 9991
rect 3031 9987 3034 9991
rect 3038 9987 3041 9991
rect 3045 9987 3048 9991
rect 3052 9987 3055 9991
rect 3059 9987 3062 9991
rect 3066 9987 3069 9991
rect 3073 9987 3076 9991
rect 3080 9987 3083 9991
rect 3087 9987 3092 9991
rect 2996 9986 3092 9987
rect 2996 9982 2999 9986
rect 3003 9982 3006 9986
rect 3010 9982 3013 9986
rect 3017 9982 3020 9986
rect 3024 9982 3027 9986
rect 3031 9982 3034 9986
rect 3038 9982 3041 9986
rect 3045 9982 3048 9986
rect 3052 9982 3055 9986
rect 3059 9982 3062 9986
rect 3066 9982 3069 9986
rect 3073 9982 3076 9986
rect 3080 9982 3083 9986
rect 3087 9982 3092 9986
rect 2996 9981 3092 9982
rect 3305 9992 3308 9993
rect 3312 9992 3315 9996
rect 3319 9992 3322 9996
rect 3326 9992 3329 9996
rect 3333 9992 3336 9996
rect 3340 9992 3343 9996
rect 3347 9992 3350 9996
rect 3354 9992 3357 9996
rect 3361 9992 3364 9996
rect 3368 9992 3371 9996
rect 3375 9992 3378 9996
rect 3382 9992 3385 9996
rect 3389 9992 3392 9996
rect 3396 9993 3411 9996
rect 3604 10001 3720 10003
rect 3604 9997 3617 10001
rect 3621 9997 3624 10001
rect 3628 9997 3631 10001
rect 3635 9997 3638 10001
rect 3642 9997 3645 10001
rect 3649 9997 3652 10001
rect 3656 9997 3659 10001
rect 3663 9997 3666 10001
rect 3670 9997 3673 10001
rect 3677 9997 3680 10001
rect 3684 9997 3687 10001
rect 3691 9997 3694 10001
rect 3698 9997 3701 10001
rect 3705 9997 3720 10001
rect 3604 9996 3720 9997
rect 3604 9993 3617 9996
rect 3396 9992 3401 9993
rect 3305 9991 3401 9992
rect 3305 9987 3308 9991
rect 3312 9987 3315 9991
rect 3319 9987 3322 9991
rect 3326 9987 3329 9991
rect 3333 9987 3336 9991
rect 3340 9987 3343 9991
rect 3347 9987 3350 9991
rect 3354 9987 3357 9991
rect 3361 9987 3364 9991
rect 3368 9987 3371 9991
rect 3375 9987 3378 9991
rect 3382 9987 3385 9991
rect 3389 9987 3392 9991
rect 3396 9987 3401 9991
rect 3305 9986 3401 9987
rect 3305 9982 3308 9986
rect 3312 9982 3315 9986
rect 3319 9982 3322 9986
rect 3326 9982 3329 9986
rect 3333 9982 3336 9986
rect 3340 9982 3343 9986
rect 3347 9982 3350 9986
rect 3354 9982 3357 9986
rect 3361 9982 3364 9986
rect 3368 9982 3371 9986
rect 3375 9982 3378 9986
rect 3382 9982 3385 9986
rect 3389 9982 3392 9986
rect 3396 9982 3401 9986
rect 3305 9981 3401 9982
rect 3614 9992 3617 9993
rect 3621 9992 3624 9996
rect 3628 9992 3631 9996
rect 3635 9992 3638 9996
rect 3642 9992 3645 9996
rect 3649 9992 3652 9996
rect 3656 9992 3659 9996
rect 3663 9992 3666 9996
rect 3670 9992 3673 9996
rect 3677 9992 3680 9996
rect 3684 9992 3687 9996
rect 3691 9992 3694 9996
rect 3698 9992 3701 9996
rect 3705 9993 3720 9996
rect 3913 10001 4029 10003
rect 3913 9997 3926 10001
rect 3930 9997 3933 10001
rect 3937 9997 3940 10001
rect 3944 9997 3947 10001
rect 3951 9997 3954 10001
rect 3958 9997 3961 10001
rect 3965 9997 3968 10001
rect 3972 9997 3975 10001
rect 3979 9997 3982 10001
rect 3986 9997 3989 10001
rect 3993 9997 3996 10001
rect 4000 9997 4003 10001
rect 4007 9997 4010 10001
rect 4014 9997 4029 10001
rect 3913 9996 4029 9997
rect 3913 9993 3926 9996
rect 3705 9992 3710 9993
rect 3614 9991 3710 9992
rect 3614 9987 3617 9991
rect 3621 9987 3624 9991
rect 3628 9987 3631 9991
rect 3635 9987 3638 9991
rect 3642 9987 3645 9991
rect 3649 9987 3652 9991
rect 3656 9987 3659 9991
rect 3663 9987 3666 9991
rect 3670 9987 3673 9991
rect 3677 9987 3680 9991
rect 3684 9987 3687 9991
rect 3691 9987 3694 9991
rect 3698 9987 3701 9991
rect 3705 9987 3710 9991
rect 3614 9986 3710 9987
rect 3614 9982 3617 9986
rect 3621 9982 3624 9986
rect 3628 9982 3631 9986
rect 3635 9982 3638 9986
rect 3642 9982 3645 9986
rect 3649 9982 3652 9986
rect 3656 9982 3659 9986
rect 3663 9982 3666 9986
rect 3670 9982 3673 9986
rect 3677 9982 3680 9986
rect 3684 9982 3687 9986
rect 3691 9982 3694 9986
rect 3698 9982 3701 9986
rect 3705 9982 3710 9986
rect 3614 9981 3710 9982
rect 3923 9992 3926 9993
rect 3930 9992 3933 9996
rect 3937 9992 3940 9996
rect 3944 9992 3947 9996
rect 3951 9992 3954 9996
rect 3958 9992 3961 9996
rect 3965 9992 3968 9996
rect 3972 9992 3975 9996
rect 3979 9992 3982 9996
rect 3986 9992 3989 9996
rect 3993 9992 3996 9996
rect 4000 9992 4003 9996
rect 4007 9992 4010 9996
rect 4014 9993 4029 9996
rect 4014 9992 4019 9993
rect 3923 9991 4019 9992
rect 3923 9987 3926 9991
rect 3930 9987 3933 9991
rect 3937 9987 3940 9991
rect 3944 9987 3947 9991
rect 3951 9987 3954 9991
rect 3958 9987 3961 9991
rect 3965 9987 3968 9991
rect 3972 9987 3975 9991
rect 3979 9987 3982 9991
rect 3986 9987 3989 9991
rect 3993 9987 3996 9991
rect 4000 9987 4003 9991
rect 4007 9987 4010 9991
rect 4014 9987 4019 9991
rect 3923 9986 4019 9987
rect 3923 9982 3926 9986
rect 3930 9982 3933 9986
rect 3937 9982 3940 9986
rect 3944 9982 3947 9986
rect 3951 9982 3954 9986
rect 3958 9982 3961 9986
rect 3965 9982 3968 9986
rect 3972 9982 3975 9986
rect 3979 9982 3982 9986
rect 3986 9982 3989 9986
rect 3993 9982 3996 9986
rect 4000 9982 4003 9986
rect 4007 9982 4010 9986
rect 4014 9982 4019 9986
rect 3923 9981 4019 9982
rect 1376 9974 1377 9978
rect 1381 9974 1382 9978
rect 1386 9974 1387 9978
rect 1391 9974 1392 9978
rect 1396 9974 1397 9978
rect 1401 9974 1402 9978
rect 1406 9974 1407 9978
rect 1411 9974 1412 9978
rect 1416 9974 1417 9978
rect 1421 9974 1422 9978
rect 1426 9974 1427 9978
rect 1431 9974 1432 9978
rect 1436 9974 1437 9978
rect 1441 9974 1442 9978
rect 1446 9974 1447 9978
rect 1451 9974 1452 9978
rect 1456 9974 1457 9978
rect 1461 9974 1462 9978
rect 1372 9973 1376 9974
rect 1372 9968 1376 9969
rect 1462 9973 1466 9974
rect 1462 9968 1466 9969
rect 1372 9963 1376 9964
rect 1372 9958 1376 9959
rect 1372 9953 1376 9954
rect 1372 9948 1376 9949
rect 1372 9943 1376 9944
rect 1372 9938 1376 9939
rect 1372 9933 1376 9934
rect 1372 9928 1376 9929
rect 1372 9923 1376 9924
rect 1372 9918 1376 9919
rect 1372 9913 1376 9914
rect 1372 9908 1376 9909
rect 1372 9903 1376 9904
rect 1372 9898 1376 9899
rect 1372 9893 1376 9894
rect 1372 9888 1376 9889
rect 1372 9883 1376 9884
rect 1372 9878 1376 9879
rect 1372 9873 1376 9874
rect 1372 9868 1376 9869
rect 1372 9863 1376 9864
rect 1372 9858 1376 9859
rect 1372 9853 1376 9854
rect 1372 9848 1376 9849
rect 1389 9961 1392 9965
rect 1396 9961 1397 9965
rect 1401 9961 1402 9965
rect 1406 9961 1407 9965
rect 1411 9961 1412 9965
rect 1416 9961 1417 9965
rect 1421 9961 1422 9965
rect 1426 9961 1427 9965
rect 1431 9961 1432 9965
rect 1436 9961 1437 9965
rect 1441 9961 1442 9965
rect 1446 9961 1449 9965
rect 1385 9958 1389 9961
rect 1385 9953 1389 9954
rect 1449 9958 1453 9961
rect 1449 9953 1453 9954
rect 1385 9948 1389 9949
rect 1385 9943 1389 9944
rect 1385 9938 1389 9939
rect 1385 9933 1389 9934
rect 1385 9928 1389 9929
rect 1385 9923 1389 9924
rect 1385 9918 1389 9919
rect 1385 9913 1389 9914
rect 1385 9908 1389 9909
rect 1385 9903 1389 9904
rect 1385 9898 1389 9899
rect 1385 9893 1389 9894
rect 1385 9888 1389 9889
rect 1385 9883 1389 9884
rect 1385 9878 1389 9879
rect 1385 9873 1389 9874
rect 1385 9868 1389 9869
rect 1401 9949 1402 9953
rect 1406 9949 1407 9953
rect 1411 9949 1412 9953
rect 1416 9949 1417 9953
rect 1421 9949 1422 9953
rect 1426 9949 1427 9953
rect 1431 9949 1432 9953
rect 1436 9949 1437 9953
rect 1397 9948 1441 9949
rect 1401 9944 1402 9948
rect 1406 9944 1407 9948
rect 1411 9944 1412 9948
rect 1416 9944 1417 9948
rect 1421 9944 1422 9948
rect 1426 9944 1427 9948
rect 1431 9944 1432 9948
rect 1436 9944 1437 9948
rect 1397 9943 1441 9944
rect 1401 9939 1402 9943
rect 1406 9939 1407 9943
rect 1411 9939 1412 9943
rect 1416 9939 1417 9943
rect 1421 9939 1422 9943
rect 1426 9939 1427 9943
rect 1431 9939 1432 9943
rect 1436 9939 1437 9943
rect 1397 9938 1441 9939
rect 1401 9934 1402 9938
rect 1406 9934 1407 9938
rect 1411 9934 1412 9938
rect 1416 9934 1417 9938
rect 1421 9934 1422 9938
rect 1426 9934 1427 9938
rect 1431 9934 1432 9938
rect 1436 9934 1437 9938
rect 1397 9933 1441 9934
rect 1401 9929 1402 9933
rect 1406 9929 1407 9933
rect 1411 9929 1412 9933
rect 1416 9929 1417 9933
rect 1421 9929 1422 9933
rect 1426 9929 1427 9933
rect 1431 9929 1432 9933
rect 1436 9929 1437 9933
rect 1397 9928 1441 9929
rect 1401 9924 1402 9928
rect 1406 9924 1407 9928
rect 1411 9924 1412 9928
rect 1416 9924 1417 9928
rect 1421 9924 1422 9928
rect 1426 9924 1427 9928
rect 1431 9924 1432 9928
rect 1436 9924 1437 9928
rect 1397 9923 1441 9924
rect 1401 9919 1402 9923
rect 1406 9919 1407 9923
rect 1411 9919 1412 9923
rect 1416 9919 1417 9923
rect 1421 9919 1422 9923
rect 1426 9919 1427 9923
rect 1431 9919 1432 9923
rect 1436 9919 1437 9923
rect 1397 9918 1441 9919
rect 1401 9914 1402 9918
rect 1406 9914 1407 9918
rect 1411 9914 1412 9918
rect 1416 9914 1417 9918
rect 1421 9914 1422 9918
rect 1426 9914 1427 9918
rect 1431 9914 1432 9918
rect 1436 9914 1437 9918
rect 1397 9913 1441 9914
rect 1401 9909 1402 9913
rect 1406 9909 1407 9913
rect 1411 9909 1412 9913
rect 1416 9909 1417 9913
rect 1421 9909 1422 9913
rect 1426 9909 1427 9913
rect 1431 9909 1432 9913
rect 1436 9909 1437 9913
rect 1397 9908 1441 9909
rect 1401 9904 1402 9908
rect 1406 9904 1407 9908
rect 1411 9904 1412 9908
rect 1416 9904 1417 9908
rect 1421 9904 1422 9908
rect 1426 9904 1427 9908
rect 1431 9904 1432 9908
rect 1436 9904 1437 9908
rect 1397 9903 1441 9904
rect 1401 9899 1402 9903
rect 1406 9899 1407 9903
rect 1411 9899 1412 9903
rect 1416 9899 1417 9903
rect 1421 9899 1422 9903
rect 1426 9899 1427 9903
rect 1431 9899 1432 9903
rect 1436 9899 1437 9903
rect 1397 9898 1441 9899
rect 1401 9894 1402 9898
rect 1406 9894 1407 9898
rect 1411 9894 1412 9898
rect 1416 9894 1417 9898
rect 1421 9894 1422 9898
rect 1426 9894 1427 9898
rect 1431 9894 1432 9898
rect 1436 9894 1437 9898
rect 1397 9893 1441 9894
rect 1401 9889 1402 9893
rect 1406 9889 1407 9893
rect 1411 9889 1412 9893
rect 1416 9889 1417 9893
rect 1421 9889 1422 9893
rect 1426 9889 1427 9893
rect 1431 9889 1432 9893
rect 1436 9889 1437 9893
rect 1397 9888 1441 9889
rect 1401 9884 1402 9888
rect 1406 9884 1407 9888
rect 1411 9884 1412 9888
rect 1416 9884 1417 9888
rect 1421 9884 1422 9888
rect 1426 9884 1427 9888
rect 1431 9884 1432 9888
rect 1436 9884 1437 9888
rect 1397 9883 1441 9884
rect 1401 9879 1402 9883
rect 1406 9879 1407 9883
rect 1411 9879 1412 9883
rect 1416 9879 1417 9883
rect 1421 9879 1422 9883
rect 1426 9879 1427 9883
rect 1431 9879 1432 9883
rect 1436 9879 1437 9883
rect 1397 9878 1441 9879
rect 1401 9874 1402 9878
rect 1406 9874 1407 9878
rect 1411 9874 1412 9878
rect 1416 9874 1417 9878
rect 1421 9874 1422 9878
rect 1426 9874 1427 9878
rect 1431 9874 1432 9878
rect 1436 9874 1437 9878
rect 1397 9873 1441 9874
rect 1401 9869 1402 9873
rect 1406 9869 1407 9873
rect 1411 9869 1412 9873
rect 1416 9869 1417 9873
rect 1421 9869 1422 9873
rect 1426 9869 1427 9873
rect 1431 9869 1432 9873
rect 1436 9869 1437 9873
rect 1397 9868 1441 9869
rect 1401 9864 1402 9868
rect 1406 9864 1407 9868
rect 1411 9864 1412 9868
rect 1416 9864 1417 9868
rect 1421 9864 1422 9868
rect 1426 9864 1427 9868
rect 1431 9864 1432 9868
rect 1436 9864 1437 9868
rect 1449 9948 1453 9949
rect 1449 9943 1453 9944
rect 1449 9938 1453 9939
rect 1449 9933 1453 9934
rect 1449 9928 1453 9929
rect 1449 9923 1453 9924
rect 1449 9918 1453 9919
rect 1449 9913 1453 9914
rect 1449 9908 1453 9909
rect 1449 9903 1453 9904
rect 1449 9898 1453 9899
rect 1449 9893 1453 9894
rect 1449 9888 1453 9889
rect 1449 9883 1453 9884
rect 1449 9878 1453 9879
rect 1449 9873 1453 9874
rect 1449 9868 1453 9869
rect 1385 9863 1389 9864
rect 1385 9856 1389 9859
rect 1449 9863 1453 9864
rect 1449 9856 1453 9859
rect 1389 9848 1392 9856
rect 1396 9848 1397 9856
rect 1401 9848 1402 9856
rect 1406 9848 1407 9856
rect 1411 9848 1412 9856
rect 1416 9848 1417 9856
rect 1421 9848 1422 9856
rect 1426 9848 1427 9856
rect 1431 9848 1432 9856
rect 1436 9848 1437 9856
rect 1441 9848 1442 9856
rect 1446 9848 1449 9856
rect 1462 9963 1466 9964
rect 1462 9958 1466 9959
rect 1462 9953 1466 9954
rect 1462 9948 1466 9949
rect 1462 9943 1466 9944
rect 1462 9938 1466 9939
rect 1462 9933 1466 9934
rect 1462 9928 1466 9929
rect 1462 9923 1466 9924
rect 1462 9918 1466 9919
rect 1462 9913 1466 9914
rect 1462 9908 1466 9909
rect 1462 9903 1466 9904
rect 1462 9898 1466 9899
rect 1462 9893 1466 9894
rect 1462 9888 1466 9889
rect 1462 9883 1466 9884
rect 1462 9878 1466 9879
rect 1462 9873 1466 9874
rect 1462 9868 1466 9869
rect 1462 9863 1466 9864
rect 1462 9858 1466 9859
rect 1462 9853 1466 9854
rect 1462 9848 1466 9849
rect 1372 9843 1376 9844
rect 1462 9843 1466 9844
rect 1376 9839 1377 9843
rect 1381 9839 1382 9843
rect 1386 9839 1387 9843
rect 1391 9839 1392 9843
rect 1396 9839 1397 9843
rect 1401 9839 1402 9843
rect 1406 9839 1407 9843
rect 1411 9839 1412 9843
rect 1416 9839 1417 9843
rect 1421 9839 1422 9843
rect 1426 9839 1427 9843
rect 1431 9839 1432 9843
rect 1436 9839 1437 9843
rect 1441 9839 1442 9843
rect 1446 9839 1447 9843
rect 1451 9839 1452 9843
rect 1456 9839 1457 9843
rect 1461 9839 1462 9843
rect 1375 9802 1431 9839
rect 1363 9800 1431 9802
rect 1363 9796 1364 9800
rect 1368 9796 1369 9800
rect 1373 9796 1431 9800
rect 1363 9795 1431 9796
rect 1363 9791 1364 9795
rect 1368 9791 1369 9795
rect 1373 9791 1431 9795
rect 1363 9790 1431 9791
rect 1363 9786 1364 9790
rect 1368 9786 1369 9790
rect 1373 9786 1431 9790
rect 1363 9785 1431 9786
rect 1363 9781 1364 9785
rect 1368 9781 1369 9785
rect 1373 9781 1431 9785
rect 1363 9780 1431 9781
rect 1363 9776 1364 9780
rect 1368 9776 1369 9780
rect 1373 9776 1431 9780
rect 1363 9775 1431 9776
rect 1363 9771 1364 9775
rect 1368 9771 1369 9775
rect 1373 9771 1431 9775
rect 1363 9770 1431 9771
rect 1363 9766 1364 9770
rect 1368 9766 1369 9770
rect 1373 9766 1431 9770
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1319 9761 1338 9762
rect 1323 9757 1324 9761
rect 1328 9757 1329 9761
rect 1333 9757 1334 9761
rect 1319 9756 1338 9757
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1319 9751 1338 9752
rect 1323 9747 1324 9751
rect 1328 9747 1329 9751
rect 1333 9747 1334 9751
rect 1319 9746 1338 9747
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1319 9741 1338 9742
rect 1323 9737 1324 9741
rect 1328 9737 1329 9741
rect 1333 9737 1334 9741
rect 1319 9736 1338 9737
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1363 9765 1431 9766
rect 1363 9761 1364 9765
rect 1368 9761 1369 9765
rect 1373 9761 1431 9765
rect 1363 9760 1431 9761
rect 1363 9756 1364 9760
rect 1368 9756 1369 9760
rect 1373 9756 1431 9760
rect 1363 9755 1431 9756
rect 1363 9751 1364 9755
rect 1368 9751 1369 9755
rect 1373 9751 1431 9755
rect 1363 9750 1431 9751
rect 1363 9746 1364 9750
rect 1368 9746 1369 9750
rect 1373 9746 1431 9750
rect 1363 9745 1431 9746
rect 1363 9741 1364 9745
rect 1368 9741 1369 9745
rect 1373 9741 1431 9745
rect 1363 9740 1431 9741
rect 1363 9736 1364 9740
rect 1368 9736 1369 9740
rect 1373 9736 1431 9740
rect 1363 9734 1431 9736
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1319 9715 1338 9716
rect 1323 9711 1324 9715
rect 1328 9711 1329 9715
rect 1333 9711 1334 9715
rect 1319 9710 1338 9711
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1319 9705 1338 9706
rect 1323 9701 1324 9705
rect 1328 9701 1329 9705
rect 1333 9701 1334 9705
rect 1319 9700 1338 9701
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1319 9695 1338 9696
rect 1323 9691 1324 9695
rect 1328 9691 1329 9695
rect 1333 9691 1334 9695
rect 1319 9690 1338 9691
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1473 9715 1525 9981
rect 1536 9974 1537 9978
rect 1541 9974 1542 9978
rect 1546 9974 1547 9978
rect 1551 9974 1552 9978
rect 1556 9974 1557 9978
rect 1561 9974 1562 9978
rect 1566 9974 1567 9978
rect 1571 9974 1572 9978
rect 1576 9974 1577 9978
rect 1581 9974 1582 9978
rect 1586 9974 1587 9978
rect 1591 9974 1592 9978
rect 1596 9974 1597 9978
rect 1601 9974 1602 9978
rect 1606 9974 1607 9978
rect 1611 9974 1612 9978
rect 1616 9974 1617 9978
rect 1621 9974 1622 9978
rect 1532 9973 1536 9974
rect 1532 9968 1536 9969
rect 1622 9973 1626 9974
rect 1622 9968 1626 9969
rect 1532 9963 1536 9964
rect 1532 9958 1536 9959
rect 1532 9953 1536 9954
rect 1532 9948 1536 9949
rect 1532 9943 1536 9944
rect 1532 9938 1536 9939
rect 1532 9933 1536 9934
rect 1532 9928 1536 9929
rect 1532 9923 1536 9924
rect 1532 9918 1536 9919
rect 1532 9913 1536 9914
rect 1532 9908 1536 9909
rect 1532 9903 1536 9904
rect 1532 9898 1536 9899
rect 1532 9893 1536 9894
rect 1532 9888 1536 9889
rect 1532 9883 1536 9884
rect 1532 9878 1536 9879
rect 1532 9873 1536 9874
rect 1532 9868 1536 9869
rect 1532 9863 1536 9864
rect 1532 9858 1536 9859
rect 1532 9853 1536 9854
rect 1532 9848 1536 9849
rect 1549 9961 1552 9965
rect 1556 9961 1557 9965
rect 1561 9961 1562 9965
rect 1566 9961 1567 9965
rect 1571 9961 1572 9965
rect 1576 9961 1577 9965
rect 1581 9961 1582 9965
rect 1586 9961 1587 9965
rect 1591 9961 1592 9965
rect 1596 9961 1597 9965
rect 1601 9961 1602 9965
rect 1606 9961 1609 9965
rect 1545 9958 1549 9961
rect 1545 9953 1549 9954
rect 1609 9958 1613 9961
rect 1609 9953 1613 9954
rect 1545 9948 1549 9949
rect 1545 9943 1549 9944
rect 1545 9938 1549 9939
rect 1545 9933 1549 9934
rect 1545 9928 1549 9929
rect 1545 9923 1549 9924
rect 1545 9918 1549 9919
rect 1545 9913 1549 9914
rect 1545 9908 1549 9909
rect 1545 9903 1549 9904
rect 1545 9898 1549 9899
rect 1545 9893 1549 9894
rect 1545 9888 1549 9889
rect 1545 9883 1549 9884
rect 1545 9878 1549 9879
rect 1545 9873 1549 9874
rect 1545 9868 1549 9869
rect 1556 9949 1557 9953
rect 1561 9949 1562 9953
rect 1566 9949 1567 9953
rect 1571 9949 1572 9953
rect 1576 9949 1577 9953
rect 1581 9949 1582 9953
rect 1586 9949 1587 9953
rect 1591 9949 1592 9953
rect 1596 9949 1597 9953
rect 1556 9948 1601 9949
rect 1556 9944 1557 9948
rect 1561 9944 1562 9948
rect 1566 9944 1567 9948
rect 1571 9944 1572 9948
rect 1576 9944 1577 9948
rect 1581 9944 1582 9948
rect 1586 9944 1587 9948
rect 1591 9944 1592 9948
rect 1596 9944 1597 9948
rect 1556 9943 1601 9944
rect 1556 9939 1557 9943
rect 1561 9939 1562 9943
rect 1566 9939 1567 9943
rect 1571 9939 1572 9943
rect 1576 9939 1577 9943
rect 1581 9939 1582 9943
rect 1586 9939 1587 9943
rect 1591 9939 1592 9943
rect 1596 9939 1597 9943
rect 1556 9938 1601 9939
rect 1556 9934 1557 9938
rect 1561 9934 1562 9938
rect 1566 9934 1567 9938
rect 1571 9934 1572 9938
rect 1576 9934 1577 9938
rect 1581 9934 1582 9938
rect 1586 9934 1587 9938
rect 1591 9934 1592 9938
rect 1596 9934 1597 9938
rect 1556 9933 1601 9934
rect 1556 9929 1557 9933
rect 1561 9929 1562 9933
rect 1566 9929 1567 9933
rect 1571 9929 1572 9933
rect 1576 9929 1577 9933
rect 1581 9929 1582 9933
rect 1586 9929 1587 9933
rect 1591 9929 1592 9933
rect 1596 9929 1597 9933
rect 1556 9928 1601 9929
rect 1556 9924 1557 9928
rect 1561 9924 1562 9928
rect 1566 9924 1567 9928
rect 1571 9924 1572 9928
rect 1576 9924 1577 9928
rect 1581 9924 1582 9928
rect 1586 9924 1587 9928
rect 1591 9924 1592 9928
rect 1596 9924 1597 9928
rect 1556 9923 1601 9924
rect 1556 9919 1557 9923
rect 1561 9919 1562 9923
rect 1566 9919 1567 9923
rect 1571 9919 1572 9923
rect 1576 9919 1577 9923
rect 1581 9919 1582 9923
rect 1586 9919 1587 9923
rect 1591 9919 1592 9923
rect 1596 9919 1597 9923
rect 1556 9918 1601 9919
rect 1556 9914 1557 9918
rect 1561 9914 1562 9918
rect 1566 9914 1567 9918
rect 1571 9914 1572 9918
rect 1576 9914 1577 9918
rect 1581 9914 1582 9918
rect 1586 9914 1587 9918
rect 1591 9914 1592 9918
rect 1596 9914 1597 9918
rect 1556 9913 1601 9914
rect 1556 9909 1557 9913
rect 1561 9909 1562 9913
rect 1566 9909 1567 9913
rect 1571 9909 1572 9913
rect 1576 9909 1577 9913
rect 1581 9909 1582 9913
rect 1586 9909 1587 9913
rect 1591 9909 1592 9913
rect 1596 9909 1597 9913
rect 1556 9908 1601 9909
rect 1556 9904 1557 9908
rect 1561 9904 1562 9908
rect 1566 9904 1567 9908
rect 1571 9904 1572 9908
rect 1576 9904 1577 9908
rect 1581 9904 1582 9908
rect 1586 9904 1587 9908
rect 1591 9904 1592 9908
rect 1596 9904 1597 9908
rect 1556 9903 1601 9904
rect 1556 9899 1557 9903
rect 1561 9899 1562 9903
rect 1566 9899 1567 9903
rect 1571 9899 1572 9903
rect 1576 9899 1577 9903
rect 1581 9899 1582 9903
rect 1586 9899 1587 9903
rect 1591 9899 1592 9903
rect 1596 9899 1597 9903
rect 1556 9898 1601 9899
rect 1556 9894 1557 9898
rect 1561 9894 1562 9898
rect 1566 9894 1567 9898
rect 1571 9894 1572 9898
rect 1576 9894 1577 9898
rect 1581 9894 1582 9898
rect 1586 9894 1587 9898
rect 1591 9894 1592 9898
rect 1596 9894 1597 9898
rect 1556 9893 1601 9894
rect 1556 9889 1557 9893
rect 1561 9889 1562 9893
rect 1566 9889 1567 9893
rect 1571 9889 1572 9893
rect 1576 9889 1577 9893
rect 1581 9889 1582 9893
rect 1586 9889 1587 9893
rect 1591 9889 1592 9893
rect 1596 9889 1597 9893
rect 1556 9888 1601 9889
rect 1556 9884 1557 9888
rect 1561 9884 1562 9888
rect 1566 9884 1567 9888
rect 1571 9884 1572 9888
rect 1576 9884 1577 9888
rect 1581 9884 1582 9888
rect 1586 9884 1587 9888
rect 1591 9884 1592 9888
rect 1596 9884 1597 9888
rect 1556 9883 1601 9884
rect 1556 9879 1557 9883
rect 1561 9879 1562 9883
rect 1566 9879 1567 9883
rect 1571 9879 1572 9883
rect 1576 9879 1577 9883
rect 1581 9879 1582 9883
rect 1586 9879 1587 9883
rect 1591 9879 1592 9883
rect 1596 9879 1597 9883
rect 1556 9878 1601 9879
rect 1556 9874 1557 9878
rect 1561 9874 1562 9878
rect 1566 9874 1567 9878
rect 1571 9874 1572 9878
rect 1576 9874 1577 9878
rect 1581 9874 1582 9878
rect 1586 9874 1587 9878
rect 1591 9874 1592 9878
rect 1596 9874 1597 9878
rect 1556 9873 1601 9874
rect 1556 9869 1557 9873
rect 1561 9869 1562 9873
rect 1566 9869 1567 9873
rect 1571 9869 1572 9873
rect 1576 9869 1577 9873
rect 1581 9869 1582 9873
rect 1586 9869 1587 9873
rect 1591 9869 1592 9873
rect 1596 9869 1597 9873
rect 1556 9868 1601 9869
rect 1556 9864 1557 9868
rect 1561 9864 1562 9868
rect 1566 9864 1567 9868
rect 1571 9864 1572 9868
rect 1576 9864 1577 9868
rect 1581 9864 1582 9868
rect 1586 9864 1587 9868
rect 1591 9864 1592 9868
rect 1596 9864 1597 9868
rect 1609 9948 1613 9949
rect 1609 9943 1613 9944
rect 1609 9938 1613 9939
rect 1609 9933 1613 9934
rect 1609 9928 1613 9929
rect 1609 9923 1613 9924
rect 1609 9918 1613 9919
rect 1609 9913 1613 9914
rect 1609 9908 1613 9909
rect 1609 9903 1613 9904
rect 1609 9898 1613 9899
rect 1609 9893 1613 9894
rect 1609 9888 1613 9889
rect 1609 9883 1613 9884
rect 1609 9878 1613 9879
rect 1609 9873 1613 9874
rect 1609 9868 1613 9869
rect 1545 9863 1549 9864
rect 1545 9856 1549 9859
rect 1609 9863 1613 9864
rect 1609 9856 1613 9859
rect 1549 9848 1552 9856
rect 1556 9848 1557 9856
rect 1561 9848 1562 9856
rect 1566 9848 1567 9856
rect 1571 9848 1572 9856
rect 1576 9848 1577 9856
rect 1581 9848 1582 9856
rect 1586 9848 1587 9856
rect 1591 9848 1592 9856
rect 1596 9848 1597 9856
rect 1601 9848 1602 9856
rect 1606 9848 1609 9856
rect 1622 9963 1626 9964
rect 1622 9958 1626 9959
rect 1622 9953 1626 9954
rect 1622 9948 1626 9949
rect 1622 9943 1626 9944
rect 1622 9938 1626 9939
rect 1622 9933 1626 9934
rect 1622 9928 1626 9929
rect 1622 9923 1626 9924
rect 1622 9918 1626 9919
rect 1622 9913 1626 9914
rect 1622 9908 1626 9909
rect 1622 9903 1626 9904
rect 1622 9898 1626 9899
rect 1622 9893 1626 9894
rect 1622 9888 1626 9889
rect 1622 9883 1626 9884
rect 1622 9878 1626 9879
rect 1622 9873 1626 9874
rect 1622 9868 1626 9869
rect 1622 9863 1626 9864
rect 1622 9858 1626 9859
rect 1622 9853 1626 9854
rect 1622 9848 1626 9849
rect 1532 9843 1536 9844
rect 1622 9843 1626 9844
rect 1536 9839 1537 9843
rect 1541 9839 1542 9843
rect 1546 9839 1547 9843
rect 1551 9839 1552 9843
rect 1556 9839 1557 9843
rect 1561 9839 1562 9843
rect 1566 9839 1567 9843
rect 1571 9839 1572 9843
rect 1576 9839 1577 9843
rect 1581 9839 1582 9843
rect 1586 9839 1587 9843
rect 1591 9839 1592 9843
rect 1596 9839 1597 9843
rect 1601 9839 1602 9843
rect 1606 9839 1607 9843
rect 1611 9839 1612 9843
rect 1616 9839 1617 9843
rect 1621 9839 1622 9843
rect 1685 9974 1686 9978
rect 1690 9974 1691 9978
rect 1695 9974 1696 9978
rect 1700 9974 1701 9978
rect 1705 9974 1706 9978
rect 1710 9974 1711 9978
rect 1715 9974 1716 9978
rect 1720 9974 1721 9978
rect 1725 9974 1726 9978
rect 1730 9974 1731 9978
rect 1735 9974 1736 9978
rect 1740 9974 1741 9978
rect 1745 9974 1746 9978
rect 1750 9974 1751 9978
rect 1755 9974 1756 9978
rect 1760 9974 1761 9978
rect 1765 9974 1766 9978
rect 1770 9974 1771 9978
rect 1681 9973 1685 9974
rect 1681 9968 1685 9969
rect 1771 9973 1775 9974
rect 1771 9968 1775 9969
rect 1681 9963 1685 9964
rect 1681 9958 1685 9959
rect 1681 9953 1685 9954
rect 1681 9948 1685 9949
rect 1681 9943 1685 9944
rect 1681 9938 1685 9939
rect 1681 9933 1685 9934
rect 1681 9928 1685 9929
rect 1681 9923 1685 9924
rect 1681 9918 1685 9919
rect 1681 9913 1685 9914
rect 1681 9908 1685 9909
rect 1681 9903 1685 9904
rect 1681 9898 1685 9899
rect 1681 9893 1685 9894
rect 1681 9888 1685 9889
rect 1681 9883 1685 9884
rect 1681 9878 1685 9879
rect 1681 9873 1685 9874
rect 1681 9868 1685 9869
rect 1681 9863 1685 9864
rect 1681 9858 1685 9859
rect 1681 9853 1685 9854
rect 1681 9848 1685 9849
rect 1698 9961 1701 9965
rect 1705 9961 1706 9965
rect 1710 9961 1711 9965
rect 1715 9961 1716 9965
rect 1720 9961 1721 9965
rect 1725 9961 1726 9965
rect 1730 9961 1731 9965
rect 1735 9961 1736 9965
rect 1740 9961 1741 9965
rect 1745 9961 1746 9965
rect 1750 9961 1751 9965
rect 1755 9961 1758 9965
rect 1694 9958 1698 9961
rect 1694 9953 1698 9954
rect 1758 9958 1762 9961
rect 1758 9953 1762 9954
rect 1694 9948 1698 9949
rect 1694 9943 1698 9944
rect 1694 9938 1698 9939
rect 1694 9933 1698 9934
rect 1694 9928 1698 9929
rect 1694 9923 1698 9924
rect 1694 9918 1698 9919
rect 1694 9913 1698 9914
rect 1694 9908 1698 9909
rect 1694 9903 1698 9904
rect 1694 9898 1698 9899
rect 1694 9893 1698 9894
rect 1694 9888 1698 9889
rect 1694 9883 1698 9884
rect 1694 9878 1698 9879
rect 1694 9873 1698 9874
rect 1694 9868 1698 9869
rect 1710 9949 1711 9953
rect 1715 9949 1716 9953
rect 1720 9949 1721 9953
rect 1725 9949 1726 9953
rect 1730 9949 1731 9953
rect 1735 9949 1736 9953
rect 1740 9949 1741 9953
rect 1745 9949 1746 9953
rect 1706 9948 1750 9949
rect 1710 9944 1711 9948
rect 1715 9944 1716 9948
rect 1720 9944 1721 9948
rect 1725 9944 1726 9948
rect 1730 9944 1731 9948
rect 1735 9944 1736 9948
rect 1740 9944 1741 9948
rect 1745 9944 1746 9948
rect 1706 9943 1750 9944
rect 1710 9939 1711 9943
rect 1715 9939 1716 9943
rect 1720 9939 1721 9943
rect 1725 9939 1726 9943
rect 1730 9939 1731 9943
rect 1735 9939 1736 9943
rect 1740 9939 1741 9943
rect 1745 9939 1746 9943
rect 1706 9938 1750 9939
rect 1710 9934 1711 9938
rect 1715 9934 1716 9938
rect 1720 9934 1721 9938
rect 1725 9934 1726 9938
rect 1730 9934 1731 9938
rect 1735 9934 1736 9938
rect 1740 9934 1741 9938
rect 1745 9934 1746 9938
rect 1706 9933 1750 9934
rect 1710 9929 1711 9933
rect 1715 9929 1716 9933
rect 1720 9929 1721 9933
rect 1725 9929 1726 9933
rect 1730 9929 1731 9933
rect 1735 9929 1736 9933
rect 1740 9929 1741 9933
rect 1745 9929 1746 9933
rect 1706 9928 1750 9929
rect 1710 9924 1711 9928
rect 1715 9924 1716 9928
rect 1720 9924 1721 9928
rect 1725 9924 1726 9928
rect 1730 9924 1731 9928
rect 1735 9924 1736 9928
rect 1740 9924 1741 9928
rect 1745 9924 1746 9928
rect 1706 9923 1750 9924
rect 1710 9919 1711 9923
rect 1715 9919 1716 9923
rect 1720 9919 1721 9923
rect 1725 9919 1726 9923
rect 1730 9919 1731 9923
rect 1735 9919 1736 9923
rect 1740 9919 1741 9923
rect 1745 9919 1746 9923
rect 1706 9918 1750 9919
rect 1710 9914 1711 9918
rect 1715 9914 1716 9918
rect 1720 9914 1721 9918
rect 1725 9914 1726 9918
rect 1730 9914 1731 9918
rect 1735 9914 1736 9918
rect 1740 9914 1741 9918
rect 1745 9914 1746 9918
rect 1706 9913 1750 9914
rect 1710 9909 1711 9913
rect 1715 9909 1716 9913
rect 1720 9909 1721 9913
rect 1725 9909 1726 9913
rect 1730 9909 1731 9913
rect 1735 9909 1736 9913
rect 1740 9909 1741 9913
rect 1745 9909 1746 9913
rect 1706 9908 1750 9909
rect 1710 9904 1711 9908
rect 1715 9904 1716 9908
rect 1720 9904 1721 9908
rect 1725 9904 1726 9908
rect 1730 9904 1731 9908
rect 1735 9904 1736 9908
rect 1740 9904 1741 9908
rect 1745 9904 1746 9908
rect 1706 9903 1750 9904
rect 1710 9899 1711 9903
rect 1715 9899 1716 9903
rect 1720 9899 1721 9903
rect 1725 9899 1726 9903
rect 1730 9899 1731 9903
rect 1735 9899 1736 9903
rect 1740 9899 1741 9903
rect 1745 9899 1746 9903
rect 1706 9898 1750 9899
rect 1710 9894 1711 9898
rect 1715 9894 1716 9898
rect 1720 9894 1721 9898
rect 1725 9894 1726 9898
rect 1730 9894 1731 9898
rect 1735 9894 1736 9898
rect 1740 9894 1741 9898
rect 1745 9894 1746 9898
rect 1706 9893 1750 9894
rect 1710 9889 1711 9893
rect 1715 9889 1716 9893
rect 1720 9889 1721 9893
rect 1725 9889 1726 9893
rect 1730 9889 1731 9893
rect 1735 9889 1736 9893
rect 1740 9889 1741 9893
rect 1745 9889 1746 9893
rect 1706 9888 1750 9889
rect 1710 9884 1711 9888
rect 1715 9884 1716 9888
rect 1720 9884 1721 9888
rect 1725 9884 1726 9888
rect 1730 9884 1731 9888
rect 1735 9884 1736 9888
rect 1740 9884 1741 9888
rect 1745 9884 1746 9888
rect 1706 9883 1750 9884
rect 1710 9879 1711 9883
rect 1715 9879 1716 9883
rect 1720 9879 1721 9883
rect 1725 9879 1726 9883
rect 1730 9879 1731 9883
rect 1735 9879 1736 9883
rect 1740 9879 1741 9883
rect 1745 9879 1746 9883
rect 1706 9878 1750 9879
rect 1710 9874 1711 9878
rect 1715 9874 1716 9878
rect 1720 9874 1721 9878
rect 1725 9874 1726 9878
rect 1730 9874 1731 9878
rect 1735 9874 1736 9878
rect 1740 9874 1741 9878
rect 1745 9874 1746 9878
rect 1706 9873 1750 9874
rect 1710 9869 1711 9873
rect 1715 9869 1716 9873
rect 1720 9869 1721 9873
rect 1725 9869 1726 9873
rect 1730 9869 1731 9873
rect 1735 9869 1736 9873
rect 1740 9869 1741 9873
rect 1745 9869 1746 9873
rect 1706 9868 1750 9869
rect 1710 9864 1711 9868
rect 1715 9864 1716 9868
rect 1720 9864 1721 9868
rect 1725 9864 1726 9868
rect 1730 9864 1731 9868
rect 1735 9864 1736 9868
rect 1740 9864 1741 9868
rect 1745 9864 1746 9868
rect 1758 9948 1762 9949
rect 1758 9943 1762 9944
rect 1758 9938 1762 9939
rect 1758 9933 1762 9934
rect 1758 9928 1762 9929
rect 1758 9923 1762 9924
rect 1758 9918 1762 9919
rect 1758 9913 1762 9914
rect 1758 9908 1762 9909
rect 1758 9903 1762 9904
rect 1758 9898 1762 9899
rect 1758 9893 1762 9894
rect 1758 9888 1762 9889
rect 1758 9883 1762 9884
rect 1758 9878 1762 9879
rect 1758 9873 1762 9874
rect 1758 9868 1762 9869
rect 1694 9863 1698 9864
rect 1694 9856 1698 9859
rect 1758 9863 1762 9864
rect 1758 9856 1762 9859
rect 1698 9848 1701 9856
rect 1705 9848 1706 9856
rect 1710 9848 1711 9856
rect 1715 9848 1716 9856
rect 1720 9848 1721 9856
rect 1725 9848 1726 9856
rect 1730 9848 1731 9856
rect 1735 9848 1736 9856
rect 1740 9848 1741 9856
rect 1745 9848 1746 9856
rect 1750 9848 1751 9856
rect 1755 9848 1758 9856
rect 1771 9963 1775 9964
rect 1771 9958 1775 9959
rect 1771 9953 1775 9954
rect 1797 9961 1818 9981
rect 1845 9974 1846 9978
rect 1850 9974 1851 9978
rect 1855 9974 1856 9978
rect 1860 9974 1861 9978
rect 1865 9974 1866 9978
rect 1870 9974 1871 9978
rect 1875 9974 1876 9978
rect 1880 9974 1881 9978
rect 1885 9974 1886 9978
rect 1890 9974 1891 9978
rect 1895 9974 1896 9978
rect 1900 9974 1901 9978
rect 1905 9974 1906 9978
rect 1910 9974 1911 9978
rect 1915 9974 1916 9978
rect 1920 9974 1921 9978
rect 1925 9974 1926 9978
rect 1930 9974 1931 9978
rect 1841 9973 1845 9974
rect 1841 9968 1845 9969
rect 1931 9973 1935 9974
rect 1931 9968 1935 9969
rect 1841 9963 1845 9964
rect 1841 9958 1845 9959
rect 1841 9953 1845 9954
rect 1771 9948 1775 9949
rect 1771 9943 1775 9944
rect 1771 9938 1775 9939
rect 1771 9933 1775 9934
rect 1771 9928 1775 9929
rect 1771 9923 1775 9924
rect 1771 9918 1775 9919
rect 1771 9913 1775 9914
rect 1771 9908 1775 9909
rect 1771 9903 1775 9904
rect 1771 9898 1775 9899
rect 1771 9893 1775 9894
rect 1771 9888 1775 9889
rect 1771 9883 1775 9884
rect 1841 9948 1845 9949
rect 1841 9943 1845 9944
rect 1841 9938 1845 9939
rect 1841 9933 1845 9934
rect 1841 9928 1845 9929
rect 1841 9923 1845 9924
rect 1841 9918 1845 9919
rect 1841 9913 1845 9914
rect 1841 9908 1845 9909
rect 1841 9903 1845 9904
rect 1841 9898 1845 9899
rect 1841 9893 1845 9894
rect 1841 9888 1845 9889
rect 1841 9883 1845 9884
rect 1771 9878 1775 9879
rect 1771 9873 1775 9874
rect 1771 9868 1775 9869
rect 1771 9863 1775 9864
rect 1771 9858 1775 9859
rect 1771 9853 1775 9854
rect 1771 9848 1775 9849
rect 1681 9843 1685 9844
rect 1797 9846 1818 9874
rect 1841 9878 1845 9879
rect 1841 9873 1845 9874
rect 1841 9868 1845 9869
rect 1841 9863 1845 9864
rect 1841 9858 1845 9859
rect 1841 9853 1845 9854
rect 1841 9848 1845 9849
rect 1858 9961 1861 9965
rect 1865 9961 1866 9965
rect 1870 9961 1871 9965
rect 1875 9961 1876 9965
rect 1880 9961 1881 9965
rect 1885 9961 1886 9965
rect 1890 9961 1891 9965
rect 1895 9961 1896 9965
rect 1900 9961 1901 9965
rect 1905 9961 1906 9965
rect 1910 9961 1911 9965
rect 1915 9961 1918 9965
rect 1854 9958 1858 9961
rect 1854 9953 1858 9954
rect 1918 9958 1922 9961
rect 1918 9953 1922 9954
rect 1854 9948 1858 9949
rect 1854 9943 1858 9944
rect 1854 9938 1858 9939
rect 1854 9933 1858 9934
rect 1854 9928 1858 9929
rect 1854 9923 1858 9924
rect 1854 9918 1858 9919
rect 1854 9913 1858 9914
rect 1854 9908 1858 9909
rect 1854 9903 1858 9904
rect 1854 9898 1858 9899
rect 1854 9893 1858 9894
rect 1854 9888 1858 9889
rect 1854 9883 1858 9884
rect 1854 9878 1858 9879
rect 1854 9873 1858 9874
rect 1854 9868 1858 9869
rect 1865 9949 1866 9953
rect 1870 9949 1871 9953
rect 1875 9949 1876 9953
rect 1880 9949 1881 9953
rect 1885 9949 1886 9953
rect 1890 9949 1891 9953
rect 1895 9949 1896 9953
rect 1900 9949 1901 9953
rect 1905 9949 1906 9953
rect 1865 9948 1910 9949
rect 1865 9944 1866 9948
rect 1870 9944 1871 9948
rect 1875 9944 1876 9948
rect 1880 9944 1881 9948
rect 1885 9944 1886 9948
rect 1890 9944 1891 9948
rect 1895 9944 1896 9948
rect 1900 9944 1901 9948
rect 1905 9944 1906 9948
rect 1865 9943 1910 9944
rect 1865 9939 1866 9943
rect 1870 9939 1871 9943
rect 1875 9939 1876 9943
rect 1880 9939 1881 9943
rect 1885 9939 1886 9943
rect 1890 9939 1891 9943
rect 1895 9939 1896 9943
rect 1900 9939 1901 9943
rect 1905 9939 1906 9943
rect 1865 9938 1910 9939
rect 1865 9934 1866 9938
rect 1870 9934 1871 9938
rect 1875 9934 1876 9938
rect 1880 9934 1881 9938
rect 1885 9934 1886 9938
rect 1890 9934 1891 9938
rect 1895 9934 1896 9938
rect 1900 9934 1901 9938
rect 1905 9934 1906 9938
rect 1865 9933 1910 9934
rect 1865 9929 1866 9933
rect 1870 9929 1871 9933
rect 1875 9929 1876 9933
rect 1880 9929 1881 9933
rect 1885 9929 1886 9933
rect 1890 9929 1891 9933
rect 1895 9929 1896 9933
rect 1900 9929 1901 9933
rect 1905 9929 1906 9933
rect 1865 9928 1910 9929
rect 1865 9924 1866 9928
rect 1870 9924 1871 9928
rect 1875 9924 1876 9928
rect 1880 9924 1881 9928
rect 1885 9924 1886 9928
rect 1890 9924 1891 9928
rect 1895 9924 1896 9928
rect 1900 9924 1901 9928
rect 1905 9924 1906 9928
rect 1865 9923 1910 9924
rect 1865 9919 1866 9923
rect 1870 9919 1871 9923
rect 1875 9919 1876 9923
rect 1880 9919 1881 9923
rect 1885 9919 1886 9923
rect 1890 9919 1891 9923
rect 1895 9919 1896 9923
rect 1900 9919 1901 9923
rect 1905 9919 1906 9923
rect 1865 9918 1910 9919
rect 1865 9914 1866 9918
rect 1870 9914 1871 9918
rect 1875 9914 1876 9918
rect 1880 9914 1881 9918
rect 1885 9914 1886 9918
rect 1890 9914 1891 9918
rect 1895 9914 1896 9918
rect 1900 9914 1901 9918
rect 1905 9914 1906 9918
rect 1865 9913 1910 9914
rect 1865 9909 1866 9913
rect 1870 9909 1871 9913
rect 1875 9909 1876 9913
rect 1880 9909 1881 9913
rect 1885 9909 1886 9913
rect 1890 9909 1891 9913
rect 1895 9909 1896 9913
rect 1900 9909 1901 9913
rect 1905 9909 1906 9913
rect 1865 9908 1910 9909
rect 1865 9904 1866 9908
rect 1870 9904 1871 9908
rect 1875 9904 1876 9908
rect 1880 9904 1881 9908
rect 1885 9904 1886 9908
rect 1890 9904 1891 9908
rect 1895 9904 1896 9908
rect 1900 9904 1901 9908
rect 1905 9904 1906 9908
rect 1865 9903 1910 9904
rect 1865 9899 1866 9903
rect 1870 9899 1871 9903
rect 1875 9899 1876 9903
rect 1880 9899 1881 9903
rect 1885 9899 1886 9903
rect 1890 9899 1891 9903
rect 1895 9899 1896 9903
rect 1900 9899 1901 9903
rect 1905 9899 1906 9903
rect 1865 9898 1910 9899
rect 1865 9894 1866 9898
rect 1870 9894 1871 9898
rect 1875 9894 1876 9898
rect 1880 9894 1881 9898
rect 1885 9894 1886 9898
rect 1890 9894 1891 9898
rect 1895 9894 1896 9898
rect 1900 9894 1901 9898
rect 1905 9894 1906 9898
rect 1865 9893 1910 9894
rect 1865 9889 1866 9893
rect 1870 9889 1871 9893
rect 1875 9889 1876 9893
rect 1880 9889 1881 9893
rect 1885 9889 1886 9893
rect 1890 9889 1891 9893
rect 1895 9889 1896 9893
rect 1900 9889 1901 9893
rect 1905 9889 1906 9893
rect 1865 9888 1910 9889
rect 1865 9884 1866 9888
rect 1870 9884 1871 9888
rect 1875 9884 1876 9888
rect 1880 9884 1881 9888
rect 1885 9884 1886 9888
rect 1890 9884 1891 9888
rect 1895 9884 1896 9888
rect 1900 9884 1901 9888
rect 1905 9884 1906 9888
rect 1865 9883 1910 9884
rect 1865 9879 1866 9883
rect 1870 9879 1871 9883
rect 1875 9879 1876 9883
rect 1880 9879 1881 9883
rect 1885 9879 1886 9883
rect 1890 9879 1891 9883
rect 1895 9879 1896 9883
rect 1900 9879 1901 9883
rect 1905 9879 1906 9883
rect 1865 9878 1910 9879
rect 1865 9874 1866 9878
rect 1870 9874 1871 9878
rect 1875 9874 1876 9878
rect 1880 9874 1881 9878
rect 1885 9874 1886 9878
rect 1890 9874 1891 9878
rect 1895 9874 1896 9878
rect 1900 9874 1901 9878
rect 1905 9874 1906 9878
rect 1865 9873 1910 9874
rect 1865 9869 1866 9873
rect 1870 9869 1871 9873
rect 1875 9869 1876 9873
rect 1880 9869 1881 9873
rect 1885 9869 1886 9873
rect 1890 9869 1891 9873
rect 1895 9869 1896 9873
rect 1900 9869 1901 9873
rect 1905 9869 1906 9873
rect 1865 9868 1910 9869
rect 1865 9864 1866 9868
rect 1870 9864 1871 9868
rect 1875 9864 1876 9868
rect 1880 9864 1881 9868
rect 1885 9864 1886 9868
rect 1890 9864 1891 9868
rect 1895 9864 1896 9868
rect 1900 9864 1901 9868
rect 1905 9864 1906 9868
rect 1918 9948 1922 9949
rect 1918 9943 1922 9944
rect 1918 9938 1922 9939
rect 1918 9933 1922 9934
rect 1918 9928 1922 9929
rect 1918 9923 1922 9924
rect 1918 9918 1922 9919
rect 1918 9913 1922 9914
rect 1918 9908 1922 9909
rect 1918 9903 1922 9904
rect 1918 9898 1922 9899
rect 1918 9893 1922 9894
rect 1918 9888 1922 9889
rect 1918 9883 1922 9884
rect 1918 9878 1922 9879
rect 1918 9873 1922 9874
rect 1918 9868 1922 9869
rect 1854 9863 1858 9864
rect 1854 9856 1858 9859
rect 1918 9863 1922 9864
rect 1918 9856 1922 9859
rect 1858 9848 1861 9856
rect 1865 9848 1866 9856
rect 1870 9848 1871 9856
rect 1875 9848 1876 9856
rect 1880 9848 1881 9856
rect 1885 9848 1886 9856
rect 1890 9848 1891 9856
rect 1895 9848 1896 9856
rect 1900 9848 1901 9856
rect 1905 9848 1906 9856
rect 1910 9848 1911 9856
rect 1915 9848 1918 9856
rect 1931 9963 1935 9964
rect 1931 9958 1935 9959
rect 1931 9953 1935 9954
rect 1931 9948 1935 9949
rect 1931 9943 1935 9944
rect 1931 9938 1935 9939
rect 1931 9933 1935 9934
rect 1931 9928 1935 9929
rect 1931 9923 1935 9924
rect 1931 9918 1935 9919
rect 1931 9913 1935 9914
rect 1931 9908 1935 9909
rect 1931 9903 1935 9904
rect 1931 9898 1935 9899
rect 1931 9893 1935 9894
rect 1931 9888 1935 9889
rect 1931 9883 1935 9884
rect 1931 9878 1935 9879
rect 1931 9873 1935 9874
rect 1931 9868 1935 9869
rect 1931 9863 1935 9864
rect 1931 9858 1935 9859
rect 1931 9853 1935 9854
rect 1931 9848 1935 9849
rect 1799 9844 1816 9846
rect 1771 9843 1775 9844
rect 1685 9839 1686 9843
rect 1690 9839 1691 9843
rect 1695 9839 1696 9843
rect 1700 9839 1701 9843
rect 1705 9839 1706 9843
rect 1710 9839 1711 9843
rect 1715 9839 1716 9843
rect 1720 9839 1721 9843
rect 1725 9839 1726 9843
rect 1730 9839 1731 9843
rect 1735 9839 1736 9843
rect 1740 9839 1741 9843
rect 1745 9839 1746 9843
rect 1750 9839 1751 9843
rect 1755 9839 1756 9843
rect 1760 9839 1761 9843
rect 1765 9839 1766 9843
rect 1770 9839 1771 9843
rect 1801 9842 1814 9844
rect 1841 9843 1845 9844
rect 1931 9843 1935 9844
rect 1473 9711 1499 9715
rect 1503 9711 1504 9715
rect 1508 9711 1525 9715
rect 1569 9722 1625 9839
rect 1684 9831 1740 9839
rect 1803 9831 1812 9842
rect 1845 9839 1846 9843
rect 1850 9839 1851 9843
rect 1855 9839 1856 9843
rect 1860 9839 1861 9843
rect 1865 9839 1866 9843
rect 1870 9839 1871 9843
rect 1875 9839 1876 9843
rect 1880 9839 1881 9843
rect 1885 9839 1886 9843
rect 1890 9839 1891 9843
rect 1895 9839 1896 9843
rect 1900 9839 1901 9843
rect 1905 9839 1906 9843
rect 1910 9839 1911 9843
rect 1915 9839 1916 9843
rect 1920 9839 1921 9843
rect 1925 9839 1926 9843
rect 1930 9839 1931 9843
rect 1994 9974 1995 9978
rect 1999 9974 2000 9978
rect 2004 9974 2005 9978
rect 2009 9974 2010 9978
rect 2014 9974 2015 9978
rect 2019 9974 2020 9978
rect 2024 9974 2025 9978
rect 2029 9974 2030 9978
rect 2034 9974 2035 9978
rect 2039 9974 2040 9978
rect 2044 9974 2045 9978
rect 2049 9974 2050 9978
rect 2054 9974 2055 9978
rect 2059 9974 2060 9978
rect 2064 9974 2065 9978
rect 2069 9974 2070 9978
rect 2074 9974 2075 9978
rect 2079 9974 2080 9978
rect 1990 9973 1994 9974
rect 1990 9968 1994 9969
rect 2080 9973 2084 9974
rect 2080 9968 2084 9969
rect 1990 9963 1994 9964
rect 1990 9958 1994 9959
rect 1990 9953 1994 9954
rect 1990 9948 1994 9949
rect 1990 9943 1994 9944
rect 1990 9938 1994 9939
rect 1990 9933 1994 9934
rect 1990 9928 1994 9929
rect 1990 9923 1994 9924
rect 1990 9918 1994 9919
rect 1990 9913 1994 9914
rect 1990 9908 1994 9909
rect 1990 9903 1994 9904
rect 1990 9898 1994 9899
rect 1990 9893 1994 9894
rect 1990 9888 1994 9889
rect 1990 9883 1994 9884
rect 1990 9878 1994 9879
rect 1990 9873 1994 9874
rect 1990 9868 1994 9869
rect 1990 9863 1994 9864
rect 1990 9858 1994 9859
rect 1990 9853 1994 9854
rect 1990 9848 1994 9849
rect 2007 9961 2010 9965
rect 2014 9961 2015 9965
rect 2019 9961 2020 9965
rect 2024 9961 2025 9965
rect 2029 9961 2030 9965
rect 2034 9961 2035 9965
rect 2039 9961 2040 9965
rect 2044 9961 2045 9965
rect 2049 9961 2050 9965
rect 2054 9961 2055 9965
rect 2059 9961 2060 9965
rect 2064 9961 2067 9965
rect 2003 9958 2007 9961
rect 2003 9953 2007 9954
rect 2067 9958 2071 9961
rect 2067 9953 2071 9954
rect 2003 9948 2007 9949
rect 2003 9943 2007 9944
rect 2003 9938 2007 9939
rect 2003 9933 2007 9934
rect 2003 9928 2007 9929
rect 2003 9923 2007 9924
rect 2003 9918 2007 9919
rect 2003 9913 2007 9914
rect 2003 9908 2007 9909
rect 2003 9903 2007 9904
rect 2003 9898 2007 9899
rect 2003 9893 2007 9894
rect 2003 9888 2007 9889
rect 2003 9883 2007 9884
rect 2003 9878 2007 9879
rect 2003 9873 2007 9874
rect 2003 9868 2007 9869
rect 2019 9949 2020 9953
rect 2024 9949 2025 9953
rect 2029 9949 2030 9953
rect 2034 9949 2035 9953
rect 2039 9949 2040 9953
rect 2044 9949 2045 9953
rect 2049 9949 2050 9953
rect 2054 9949 2055 9953
rect 2015 9948 2059 9949
rect 2019 9944 2020 9948
rect 2024 9944 2025 9948
rect 2029 9944 2030 9948
rect 2034 9944 2035 9948
rect 2039 9944 2040 9948
rect 2044 9944 2045 9948
rect 2049 9944 2050 9948
rect 2054 9944 2055 9948
rect 2015 9943 2059 9944
rect 2019 9939 2020 9943
rect 2024 9939 2025 9943
rect 2029 9939 2030 9943
rect 2034 9939 2035 9943
rect 2039 9939 2040 9943
rect 2044 9939 2045 9943
rect 2049 9939 2050 9943
rect 2054 9939 2055 9943
rect 2015 9938 2059 9939
rect 2019 9934 2020 9938
rect 2024 9934 2025 9938
rect 2029 9934 2030 9938
rect 2034 9934 2035 9938
rect 2039 9934 2040 9938
rect 2044 9934 2045 9938
rect 2049 9934 2050 9938
rect 2054 9934 2055 9938
rect 2015 9933 2059 9934
rect 2019 9929 2020 9933
rect 2024 9929 2025 9933
rect 2029 9929 2030 9933
rect 2034 9929 2035 9933
rect 2039 9929 2040 9933
rect 2044 9929 2045 9933
rect 2049 9929 2050 9933
rect 2054 9929 2055 9933
rect 2015 9928 2059 9929
rect 2019 9924 2020 9928
rect 2024 9924 2025 9928
rect 2029 9924 2030 9928
rect 2034 9924 2035 9928
rect 2039 9924 2040 9928
rect 2044 9924 2045 9928
rect 2049 9924 2050 9928
rect 2054 9924 2055 9928
rect 2015 9923 2059 9924
rect 2019 9919 2020 9923
rect 2024 9919 2025 9923
rect 2029 9919 2030 9923
rect 2034 9919 2035 9923
rect 2039 9919 2040 9923
rect 2044 9919 2045 9923
rect 2049 9919 2050 9923
rect 2054 9919 2055 9923
rect 2015 9918 2059 9919
rect 2019 9914 2020 9918
rect 2024 9914 2025 9918
rect 2029 9914 2030 9918
rect 2034 9914 2035 9918
rect 2039 9914 2040 9918
rect 2044 9914 2045 9918
rect 2049 9914 2050 9918
rect 2054 9914 2055 9918
rect 2015 9913 2059 9914
rect 2019 9909 2020 9913
rect 2024 9909 2025 9913
rect 2029 9909 2030 9913
rect 2034 9909 2035 9913
rect 2039 9909 2040 9913
rect 2044 9909 2045 9913
rect 2049 9909 2050 9913
rect 2054 9909 2055 9913
rect 2015 9908 2059 9909
rect 2019 9904 2020 9908
rect 2024 9904 2025 9908
rect 2029 9904 2030 9908
rect 2034 9904 2035 9908
rect 2039 9904 2040 9908
rect 2044 9904 2045 9908
rect 2049 9904 2050 9908
rect 2054 9904 2055 9908
rect 2015 9903 2059 9904
rect 2019 9899 2020 9903
rect 2024 9899 2025 9903
rect 2029 9899 2030 9903
rect 2034 9899 2035 9903
rect 2039 9899 2040 9903
rect 2044 9899 2045 9903
rect 2049 9899 2050 9903
rect 2054 9899 2055 9903
rect 2015 9898 2059 9899
rect 2019 9894 2020 9898
rect 2024 9894 2025 9898
rect 2029 9894 2030 9898
rect 2034 9894 2035 9898
rect 2039 9894 2040 9898
rect 2044 9894 2045 9898
rect 2049 9894 2050 9898
rect 2054 9894 2055 9898
rect 2015 9893 2059 9894
rect 2019 9889 2020 9893
rect 2024 9889 2025 9893
rect 2029 9889 2030 9893
rect 2034 9889 2035 9893
rect 2039 9889 2040 9893
rect 2044 9889 2045 9893
rect 2049 9889 2050 9893
rect 2054 9889 2055 9893
rect 2015 9888 2059 9889
rect 2019 9884 2020 9888
rect 2024 9884 2025 9888
rect 2029 9884 2030 9888
rect 2034 9884 2035 9888
rect 2039 9884 2040 9888
rect 2044 9884 2045 9888
rect 2049 9884 2050 9888
rect 2054 9884 2055 9888
rect 2015 9883 2059 9884
rect 2019 9879 2020 9883
rect 2024 9879 2025 9883
rect 2029 9879 2030 9883
rect 2034 9879 2035 9883
rect 2039 9879 2040 9883
rect 2044 9879 2045 9883
rect 2049 9879 2050 9883
rect 2054 9879 2055 9883
rect 2015 9878 2059 9879
rect 2019 9874 2020 9878
rect 2024 9874 2025 9878
rect 2029 9874 2030 9878
rect 2034 9874 2035 9878
rect 2039 9874 2040 9878
rect 2044 9874 2045 9878
rect 2049 9874 2050 9878
rect 2054 9874 2055 9878
rect 2015 9873 2059 9874
rect 2019 9869 2020 9873
rect 2024 9869 2025 9873
rect 2029 9869 2030 9873
rect 2034 9869 2035 9873
rect 2039 9869 2040 9873
rect 2044 9869 2045 9873
rect 2049 9869 2050 9873
rect 2054 9869 2055 9873
rect 2015 9868 2059 9869
rect 2019 9864 2020 9868
rect 2024 9864 2025 9868
rect 2029 9864 2030 9868
rect 2034 9864 2035 9868
rect 2039 9864 2040 9868
rect 2044 9864 2045 9868
rect 2049 9864 2050 9868
rect 2054 9864 2055 9868
rect 2067 9948 2071 9949
rect 2067 9943 2071 9944
rect 2067 9938 2071 9939
rect 2067 9933 2071 9934
rect 2067 9928 2071 9929
rect 2067 9923 2071 9924
rect 2067 9918 2071 9919
rect 2067 9913 2071 9914
rect 2067 9908 2071 9909
rect 2067 9903 2071 9904
rect 2067 9898 2071 9899
rect 2067 9893 2071 9894
rect 2067 9888 2071 9889
rect 2067 9883 2071 9884
rect 2067 9878 2071 9879
rect 2067 9873 2071 9874
rect 2067 9868 2071 9869
rect 2003 9863 2007 9864
rect 2003 9856 2007 9859
rect 2067 9863 2071 9864
rect 2067 9856 2071 9859
rect 2007 9848 2010 9856
rect 2014 9848 2015 9856
rect 2019 9848 2020 9856
rect 2024 9848 2025 9856
rect 2029 9848 2030 9856
rect 2034 9848 2035 9856
rect 2039 9848 2040 9856
rect 2044 9848 2045 9856
rect 2049 9848 2050 9856
rect 2054 9848 2055 9856
rect 2059 9848 2060 9856
rect 2064 9848 2067 9856
rect 2080 9963 2084 9964
rect 2080 9958 2084 9959
rect 2080 9953 2084 9954
rect 2106 9961 2127 9981
rect 2154 9974 2155 9978
rect 2159 9974 2160 9978
rect 2164 9974 2165 9978
rect 2169 9974 2170 9978
rect 2174 9974 2175 9978
rect 2179 9974 2180 9978
rect 2184 9974 2185 9978
rect 2189 9974 2190 9978
rect 2194 9974 2195 9978
rect 2199 9974 2200 9978
rect 2204 9974 2205 9978
rect 2209 9974 2210 9978
rect 2214 9974 2215 9978
rect 2219 9974 2220 9978
rect 2224 9974 2225 9978
rect 2229 9974 2230 9978
rect 2234 9974 2235 9978
rect 2239 9974 2240 9978
rect 2150 9973 2154 9974
rect 2150 9968 2154 9969
rect 2240 9973 2244 9974
rect 2240 9968 2244 9969
rect 2150 9963 2154 9964
rect 2150 9958 2154 9959
rect 2150 9953 2154 9954
rect 2080 9948 2084 9949
rect 2080 9943 2084 9944
rect 2080 9938 2084 9939
rect 2080 9933 2084 9934
rect 2080 9928 2084 9929
rect 2080 9923 2084 9924
rect 2080 9918 2084 9919
rect 2080 9913 2084 9914
rect 2080 9908 2084 9909
rect 2080 9903 2084 9904
rect 2080 9898 2084 9899
rect 2080 9893 2084 9894
rect 2080 9888 2084 9889
rect 2080 9883 2084 9884
rect 2150 9948 2154 9949
rect 2150 9943 2154 9944
rect 2150 9938 2154 9939
rect 2150 9933 2154 9934
rect 2150 9928 2154 9929
rect 2150 9923 2154 9924
rect 2150 9918 2154 9919
rect 2150 9913 2154 9914
rect 2150 9908 2154 9909
rect 2150 9903 2154 9904
rect 2150 9898 2154 9899
rect 2150 9893 2154 9894
rect 2150 9888 2154 9889
rect 2150 9883 2154 9884
rect 2080 9878 2084 9879
rect 2080 9873 2084 9874
rect 2080 9868 2084 9869
rect 2080 9863 2084 9864
rect 2080 9858 2084 9859
rect 2080 9853 2084 9854
rect 2080 9848 2084 9849
rect 1990 9843 1994 9844
rect 2106 9846 2127 9874
rect 2150 9878 2154 9879
rect 2150 9873 2154 9874
rect 2150 9868 2154 9869
rect 2150 9863 2154 9864
rect 2150 9858 2154 9859
rect 2150 9853 2154 9854
rect 2150 9848 2154 9849
rect 2167 9961 2170 9965
rect 2174 9961 2175 9965
rect 2179 9961 2180 9965
rect 2184 9961 2185 9965
rect 2189 9961 2190 9965
rect 2194 9961 2195 9965
rect 2199 9961 2200 9965
rect 2204 9961 2205 9965
rect 2209 9961 2210 9965
rect 2214 9961 2215 9965
rect 2219 9961 2220 9965
rect 2224 9961 2227 9965
rect 2163 9958 2167 9961
rect 2163 9953 2167 9954
rect 2227 9958 2231 9961
rect 2227 9953 2231 9954
rect 2163 9948 2167 9949
rect 2163 9943 2167 9944
rect 2163 9938 2167 9939
rect 2163 9933 2167 9934
rect 2163 9928 2167 9929
rect 2163 9923 2167 9924
rect 2163 9918 2167 9919
rect 2163 9913 2167 9914
rect 2163 9908 2167 9909
rect 2163 9903 2167 9904
rect 2163 9898 2167 9899
rect 2163 9893 2167 9894
rect 2163 9888 2167 9889
rect 2163 9883 2167 9884
rect 2163 9878 2167 9879
rect 2163 9873 2167 9874
rect 2163 9868 2167 9869
rect 2174 9949 2175 9953
rect 2179 9949 2180 9953
rect 2184 9949 2185 9953
rect 2189 9949 2190 9953
rect 2194 9949 2195 9953
rect 2199 9949 2200 9953
rect 2204 9949 2205 9953
rect 2209 9949 2210 9953
rect 2214 9949 2215 9953
rect 2174 9948 2219 9949
rect 2174 9944 2175 9948
rect 2179 9944 2180 9948
rect 2184 9944 2185 9948
rect 2189 9944 2190 9948
rect 2194 9944 2195 9948
rect 2199 9944 2200 9948
rect 2204 9944 2205 9948
rect 2209 9944 2210 9948
rect 2214 9944 2215 9948
rect 2174 9943 2219 9944
rect 2174 9939 2175 9943
rect 2179 9939 2180 9943
rect 2184 9939 2185 9943
rect 2189 9939 2190 9943
rect 2194 9939 2195 9943
rect 2199 9939 2200 9943
rect 2204 9939 2205 9943
rect 2209 9939 2210 9943
rect 2214 9939 2215 9943
rect 2174 9938 2219 9939
rect 2174 9934 2175 9938
rect 2179 9934 2180 9938
rect 2184 9934 2185 9938
rect 2189 9934 2190 9938
rect 2194 9934 2195 9938
rect 2199 9934 2200 9938
rect 2204 9934 2205 9938
rect 2209 9934 2210 9938
rect 2214 9934 2215 9938
rect 2174 9933 2219 9934
rect 2174 9929 2175 9933
rect 2179 9929 2180 9933
rect 2184 9929 2185 9933
rect 2189 9929 2190 9933
rect 2194 9929 2195 9933
rect 2199 9929 2200 9933
rect 2204 9929 2205 9933
rect 2209 9929 2210 9933
rect 2214 9929 2215 9933
rect 2174 9928 2219 9929
rect 2174 9924 2175 9928
rect 2179 9924 2180 9928
rect 2184 9924 2185 9928
rect 2189 9924 2190 9928
rect 2194 9924 2195 9928
rect 2199 9924 2200 9928
rect 2204 9924 2205 9928
rect 2209 9924 2210 9928
rect 2214 9924 2215 9928
rect 2174 9923 2219 9924
rect 2174 9919 2175 9923
rect 2179 9919 2180 9923
rect 2184 9919 2185 9923
rect 2189 9919 2190 9923
rect 2194 9919 2195 9923
rect 2199 9919 2200 9923
rect 2204 9919 2205 9923
rect 2209 9919 2210 9923
rect 2214 9919 2215 9923
rect 2174 9918 2219 9919
rect 2174 9914 2175 9918
rect 2179 9914 2180 9918
rect 2184 9914 2185 9918
rect 2189 9914 2190 9918
rect 2194 9914 2195 9918
rect 2199 9914 2200 9918
rect 2204 9914 2205 9918
rect 2209 9914 2210 9918
rect 2214 9914 2215 9918
rect 2174 9913 2219 9914
rect 2174 9909 2175 9913
rect 2179 9909 2180 9913
rect 2184 9909 2185 9913
rect 2189 9909 2190 9913
rect 2194 9909 2195 9913
rect 2199 9909 2200 9913
rect 2204 9909 2205 9913
rect 2209 9909 2210 9913
rect 2214 9909 2215 9913
rect 2174 9908 2219 9909
rect 2174 9904 2175 9908
rect 2179 9904 2180 9908
rect 2184 9904 2185 9908
rect 2189 9904 2190 9908
rect 2194 9904 2195 9908
rect 2199 9904 2200 9908
rect 2204 9904 2205 9908
rect 2209 9904 2210 9908
rect 2214 9904 2215 9908
rect 2174 9903 2219 9904
rect 2174 9899 2175 9903
rect 2179 9899 2180 9903
rect 2184 9899 2185 9903
rect 2189 9899 2190 9903
rect 2194 9899 2195 9903
rect 2199 9899 2200 9903
rect 2204 9899 2205 9903
rect 2209 9899 2210 9903
rect 2214 9899 2215 9903
rect 2174 9898 2219 9899
rect 2174 9894 2175 9898
rect 2179 9894 2180 9898
rect 2184 9894 2185 9898
rect 2189 9894 2190 9898
rect 2194 9894 2195 9898
rect 2199 9894 2200 9898
rect 2204 9894 2205 9898
rect 2209 9894 2210 9898
rect 2214 9894 2215 9898
rect 2174 9893 2219 9894
rect 2174 9889 2175 9893
rect 2179 9889 2180 9893
rect 2184 9889 2185 9893
rect 2189 9889 2190 9893
rect 2194 9889 2195 9893
rect 2199 9889 2200 9893
rect 2204 9889 2205 9893
rect 2209 9889 2210 9893
rect 2214 9889 2215 9893
rect 2174 9888 2219 9889
rect 2174 9884 2175 9888
rect 2179 9884 2180 9888
rect 2184 9884 2185 9888
rect 2189 9884 2190 9888
rect 2194 9884 2195 9888
rect 2199 9884 2200 9888
rect 2204 9884 2205 9888
rect 2209 9884 2210 9888
rect 2214 9884 2215 9888
rect 2174 9883 2219 9884
rect 2174 9879 2175 9883
rect 2179 9879 2180 9883
rect 2184 9879 2185 9883
rect 2189 9879 2190 9883
rect 2194 9879 2195 9883
rect 2199 9879 2200 9883
rect 2204 9879 2205 9883
rect 2209 9879 2210 9883
rect 2214 9879 2215 9883
rect 2174 9878 2219 9879
rect 2174 9874 2175 9878
rect 2179 9874 2180 9878
rect 2184 9874 2185 9878
rect 2189 9874 2190 9878
rect 2194 9874 2195 9878
rect 2199 9874 2200 9878
rect 2204 9874 2205 9878
rect 2209 9874 2210 9878
rect 2214 9874 2215 9878
rect 2174 9873 2219 9874
rect 2174 9869 2175 9873
rect 2179 9869 2180 9873
rect 2184 9869 2185 9873
rect 2189 9869 2190 9873
rect 2194 9869 2195 9873
rect 2199 9869 2200 9873
rect 2204 9869 2205 9873
rect 2209 9869 2210 9873
rect 2214 9869 2215 9873
rect 2174 9868 2219 9869
rect 2174 9864 2175 9868
rect 2179 9864 2180 9868
rect 2184 9864 2185 9868
rect 2189 9864 2190 9868
rect 2194 9864 2195 9868
rect 2199 9864 2200 9868
rect 2204 9864 2205 9868
rect 2209 9864 2210 9868
rect 2214 9864 2215 9868
rect 2227 9948 2231 9949
rect 2227 9943 2231 9944
rect 2227 9938 2231 9939
rect 2227 9933 2231 9934
rect 2227 9928 2231 9929
rect 2227 9923 2231 9924
rect 2227 9918 2231 9919
rect 2227 9913 2231 9914
rect 2227 9908 2231 9909
rect 2227 9903 2231 9904
rect 2227 9898 2231 9899
rect 2227 9893 2231 9894
rect 2227 9888 2231 9889
rect 2227 9883 2231 9884
rect 2227 9878 2231 9879
rect 2227 9873 2231 9874
rect 2227 9868 2231 9869
rect 2163 9863 2167 9864
rect 2163 9856 2167 9859
rect 2227 9863 2231 9864
rect 2227 9856 2231 9859
rect 2167 9848 2170 9856
rect 2174 9848 2175 9856
rect 2179 9848 2180 9856
rect 2184 9848 2185 9856
rect 2189 9848 2190 9856
rect 2194 9848 2195 9856
rect 2199 9848 2200 9856
rect 2204 9848 2205 9856
rect 2209 9848 2210 9856
rect 2214 9848 2215 9856
rect 2219 9848 2220 9856
rect 2224 9848 2227 9856
rect 2240 9963 2244 9964
rect 2240 9958 2244 9959
rect 2240 9953 2244 9954
rect 2240 9948 2244 9949
rect 2240 9943 2244 9944
rect 2240 9938 2244 9939
rect 2240 9933 2244 9934
rect 2240 9928 2244 9929
rect 2240 9923 2244 9924
rect 2240 9918 2244 9919
rect 2240 9913 2244 9914
rect 2240 9908 2244 9909
rect 2240 9903 2244 9904
rect 2240 9898 2244 9899
rect 2240 9893 2244 9894
rect 2240 9888 2244 9889
rect 2240 9883 2244 9884
rect 2240 9878 2244 9879
rect 2240 9873 2244 9874
rect 2240 9868 2244 9869
rect 2240 9863 2244 9864
rect 2240 9858 2244 9859
rect 2240 9853 2244 9854
rect 2240 9848 2244 9849
rect 2108 9844 2125 9846
rect 2080 9843 2084 9844
rect 1994 9839 1995 9843
rect 1999 9839 2000 9843
rect 2004 9839 2005 9843
rect 2009 9839 2010 9843
rect 2014 9839 2015 9843
rect 2019 9839 2020 9843
rect 2024 9839 2025 9843
rect 2029 9839 2030 9843
rect 2034 9839 2035 9843
rect 2039 9839 2040 9843
rect 2044 9839 2045 9843
rect 2049 9839 2050 9843
rect 2054 9839 2055 9843
rect 2059 9839 2060 9843
rect 2064 9839 2065 9843
rect 2069 9839 2070 9843
rect 2074 9839 2075 9843
rect 2079 9839 2080 9843
rect 2110 9842 2123 9844
rect 2150 9843 2154 9844
rect 2240 9843 2244 9844
rect 1878 9831 1934 9839
rect 1684 9827 1743 9831
rect 1869 9827 1934 9831
rect 1684 9815 1740 9827
rect 1799 9819 1829 9823
rect 1684 9811 1743 9815
rect 1813 9812 1817 9819
rect 1878 9815 1934 9827
rect 1684 9802 1740 9811
rect 1869 9811 1934 9815
rect 1799 9803 1810 9807
rect 1672 9800 1740 9802
rect 1672 9796 1673 9800
rect 1677 9796 1678 9800
rect 1682 9799 1740 9800
rect 1803 9800 1810 9803
rect 1822 9803 1829 9807
rect 1822 9800 1826 9803
rect 1682 9796 1743 9799
rect 1672 9795 1743 9796
rect 1672 9791 1673 9795
rect 1677 9791 1678 9795
rect 1682 9791 1740 9795
rect 1803 9791 1826 9800
rect 1878 9799 1934 9811
rect 1993 9831 2049 9839
rect 2112 9831 2121 9842
rect 2154 9839 2155 9843
rect 2159 9839 2160 9843
rect 2164 9839 2165 9843
rect 2169 9839 2170 9843
rect 2174 9839 2175 9843
rect 2179 9839 2180 9843
rect 2184 9839 2185 9843
rect 2189 9839 2190 9843
rect 2194 9839 2195 9843
rect 2199 9839 2200 9843
rect 2204 9839 2205 9843
rect 2209 9839 2210 9843
rect 2214 9839 2215 9843
rect 2219 9839 2220 9843
rect 2224 9839 2225 9843
rect 2229 9839 2230 9843
rect 2234 9839 2235 9843
rect 2239 9839 2240 9843
rect 2303 9974 2304 9978
rect 2308 9974 2309 9978
rect 2313 9974 2314 9978
rect 2318 9974 2319 9978
rect 2323 9974 2324 9978
rect 2328 9974 2329 9978
rect 2333 9974 2334 9978
rect 2338 9974 2339 9978
rect 2343 9974 2344 9978
rect 2348 9974 2349 9978
rect 2353 9974 2354 9978
rect 2358 9974 2359 9978
rect 2363 9974 2364 9978
rect 2368 9974 2369 9978
rect 2373 9974 2374 9978
rect 2378 9974 2379 9978
rect 2383 9974 2384 9978
rect 2388 9974 2389 9978
rect 2299 9973 2303 9974
rect 2299 9968 2303 9969
rect 2389 9973 2393 9974
rect 2389 9968 2393 9969
rect 2299 9963 2303 9964
rect 2299 9958 2303 9959
rect 2299 9953 2303 9954
rect 2299 9948 2303 9949
rect 2299 9943 2303 9944
rect 2299 9938 2303 9939
rect 2299 9933 2303 9934
rect 2299 9928 2303 9929
rect 2299 9923 2303 9924
rect 2299 9918 2303 9919
rect 2299 9913 2303 9914
rect 2299 9908 2303 9909
rect 2299 9903 2303 9904
rect 2299 9898 2303 9899
rect 2299 9893 2303 9894
rect 2299 9888 2303 9889
rect 2299 9883 2303 9884
rect 2299 9878 2303 9879
rect 2299 9873 2303 9874
rect 2299 9868 2303 9869
rect 2299 9863 2303 9864
rect 2299 9858 2303 9859
rect 2299 9853 2303 9854
rect 2299 9848 2303 9849
rect 2316 9961 2319 9965
rect 2323 9961 2324 9965
rect 2328 9961 2329 9965
rect 2333 9961 2334 9965
rect 2338 9961 2339 9965
rect 2343 9961 2344 9965
rect 2348 9961 2349 9965
rect 2353 9961 2354 9965
rect 2358 9961 2359 9965
rect 2363 9961 2364 9965
rect 2368 9961 2369 9965
rect 2373 9961 2376 9965
rect 2312 9958 2316 9961
rect 2312 9953 2316 9954
rect 2376 9958 2380 9961
rect 2376 9953 2380 9954
rect 2312 9948 2316 9949
rect 2312 9943 2316 9944
rect 2312 9938 2316 9939
rect 2312 9933 2316 9934
rect 2312 9928 2316 9929
rect 2312 9923 2316 9924
rect 2312 9918 2316 9919
rect 2312 9913 2316 9914
rect 2312 9908 2316 9909
rect 2312 9903 2316 9904
rect 2312 9898 2316 9899
rect 2312 9893 2316 9894
rect 2312 9888 2316 9889
rect 2312 9883 2316 9884
rect 2312 9878 2316 9879
rect 2312 9873 2316 9874
rect 2312 9868 2316 9869
rect 2328 9949 2329 9953
rect 2333 9949 2334 9953
rect 2338 9949 2339 9953
rect 2343 9949 2344 9953
rect 2348 9949 2349 9953
rect 2353 9949 2354 9953
rect 2358 9949 2359 9953
rect 2363 9949 2364 9953
rect 2324 9948 2368 9949
rect 2328 9944 2329 9948
rect 2333 9944 2334 9948
rect 2338 9944 2339 9948
rect 2343 9944 2344 9948
rect 2348 9944 2349 9948
rect 2353 9944 2354 9948
rect 2358 9944 2359 9948
rect 2363 9944 2364 9948
rect 2324 9943 2368 9944
rect 2328 9939 2329 9943
rect 2333 9939 2334 9943
rect 2338 9939 2339 9943
rect 2343 9939 2344 9943
rect 2348 9939 2349 9943
rect 2353 9939 2354 9943
rect 2358 9939 2359 9943
rect 2363 9939 2364 9943
rect 2324 9938 2368 9939
rect 2328 9934 2329 9938
rect 2333 9934 2334 9938
rect 2338 9934 2339 9938
rect 2343 9934 2344 9938
rect 2348 9934 2349 9938
rect 2353 9934 2354 9938
rect 2358 9934 2359 9938
rect 2363 9934 2364 9938
rect 2324 9933 2368 9934
rect 2328 9929 2329 9933
rect 2333 9929 2334 9933
rect 2338 9929 2339 9933
rect 2343 9929 2344 9933
rect 2348 9929 2349 9933
rect 2353 9929 2354 9933
rect 2358 9929 2359 9933
rect 2363 9929 2364 9933
rect 2324 9928 2368 9929
rect 2328 9924 2329 9928
rect 2333 9924 2334 9928
rect 2338 9924 2339 9928
rect 2343 9924 2344 9928
rect 2348 9924 2349 9928
rect 2353 9924 2354 9928
rect 2358 9924 2359 9928
rect 2363 9924 2364 9928
rect 2324 9923 2368 9924
rect 2328 9919 2329 9923
rect 2333 9919 2334 9923
rect 2338 9919 2339 9923
rect 2343 9919 2344 9923
rect 2348 9919 2349 9923
rect 2353 9919 2354 9923
rect 2358 9919 2359 9923
rect 2363 9919 2364 9923
rect 2324 9918 2368 9919
rect 2328 9914 2329 9918
rect 2333 9914 2334 9918
rect 2338 9914 2339 9918
rect 2343 9914 2344 9918
rect 2348 9914 2349 9918
rect 2353 9914 2354 9918
rect 2358 9914 2359 9918
rect 2363 9914 2364 9918
rect 2324 9913 2368 9914
rect 2328 9909 2329 9913
rect 2333 9909 2334 9913
rect 2338 9909 2339 9913
rect 2343 9909 2344 9913
rect 2348 9909 2349 9913
rect 2353 9909 2354 9913
rect 2358 9909 2359 9913
rect 2363 9909 2364 9913
rect 2324 9908 2368 9909
rect 2328 9904 2329 9908
rect 2333 9904 2334 9908
rect 2338 9904 2339 9908
rect 2343 9904 2344 9908
rect 2348 9904 2349 9908
rect 2353 9904 2354 9908
rect 2358 9904 2359 9908
rect 2363 9904 2364 9908
rect 2324 9903 2368 9904
rect 2328 9899 2329 9903
rect 2333 9899 2334 9903
rect 2338 9899 2339 9903
rect 2343 9899 2344 9903
rect 2348 9899 2349 9903
rect 2353 9899 2354 9903
rect 2358 9899 2359 9903
rect 2363 9899 2364 9903
rect 2324 9898 2368 9899
rect 2328 9894 2329 9898
rect 2333 9894 2334 9898
rect 2338 9894 2339 9898
rect 2343 9894 2344 9898
rect 2348 9894 2349 9898
rect 2353 9894 2354 9898
rect 2358 9894 2359 9898
rect 2363 9894 2364 9898
rect 2324 9893 2368 9894
rect 2328 9889 2329 9893
rect 2333 9889 2334 9893
rect 2338 9889 2339 9893
rect 2343 9889 2344 9893
rect 2348 9889 2349 9893
rect 2353 9889 2354 9893
rect 2358 9889 2359 9893
rect 2363 9889 2364 9893
rect 2324 9888 2368 9889
rect 2328 9884 2329 9888
rect 2333 9884 2334 9888
rect 2338 9884 2339 9888
rect 2343 9884 2344 9888
rect 2348 9884 2349 9888
rect 2353 9884 2354 9888
rect 2358 9884 2359 9888
rect 2363 9884 2364 9888
rect 2324 9883 2368 9884
rect 2328 9879 2329 9883
rect 2333 9879 2334 9883
rect 2338 9879 2339 9883
rect 2343 9879 2344 9883
rect 2348 9879 2349 9883
rect 2353 9879 2354 9883
rect 2358 9879 2359 9883
rect 2363 9879 2364 9883
rect 2324 9878 2368 9879
rect 2328 9874 2329 9878
rect 2333 9874 2334 9878
rect 2338 9874 2339 9878
rect 2343 9874 2344 9878
rect 2348 9874 2349 9878
rect 2353 9874 2354 9878
rect 2358 9874 2359 9878
rect 2363 9874 2364 9878
rect 2324 9873 2368 9874
rect 2328 9869 2329 9873
rect 2333 9869 2334 9873
rect 2338 9869 2339 9873
rect 2343 9869 2344 9873
rect 2348 9869 2349 9873
rect 2353 9869 2354 9873
rect 2358 9869 2359 9873
rect 2363 9869 2364 9873
rect 2324 9868 2368 9869
rect 2328 9864 2329 9868
rect 2333 9864 2334 9868
rect 2338 9864 2339 9868
rect 2343 9864 2344 9868
rect 2348 9864 2349 9868
rect 2353 9864 2354 9868
rect 2358 9864 2359 9868
rect 2363 9864 2364 9868
rect 2376 9948 2380 9949
rect 2376 9943 2380 9944
rect 2376 9938 2380 9939
rect 2376 9933 2380 9934
rect 2376 9928 2380 9929
rect 2376 9923 2380 9924
rect 2376 9918 2380 9919
rect 2376 9913 2380 9914
rect 2376 9908 2380 9909
rect 2376 9903 2380 9904
rect 2376 9898 2380 9899
rect 2376 9893 2380 9894
rect 2376 9888 2380 9889
rect 2376 9883 2380 9884
rect 2376 9878 2380 9879
rect 2376 9873 2380 9874
rect 2376 9868 2380 9869
rect 2312 9863 2316 9864
rect 2312 9856 2316 9859
rect 2376 9863 2380 9864
rect 2376 9856 2380 9859
rect 2316 9848 2319 9856
rect 2323 9848 2324 9856
rect 2328 9848 2329 9856
rect 2333 9848 2334 9856
rect 2338 9848 2339 9856
rect 2343 9848 2344 9856
rect 2348 9848 2349 9856
rect 2353 9848 2354 9856
rect 2358 9848 2359 9856
rect 2363 9848 2364 9856
rect 2368 9848 2369 9856
rect 2373 9848 2376 9856
rect 2389 9963 2393 9964
rect 2389 9958 2393 9959
rect 2389 9953 2393 9954
rect 2415 9961 2436 9981
rect 2463 9974 2464 9978
rect 2468 9974 2469 9978
rect 2473 9974 2474 9978
rect 2478 9974 2479 9978
rect 2483 9974 2484 9978
rect 2488 9974 2489 9978
rect 2493 9974 2494 9978
rect 2498 9974 2499 9978
rect 2503 9974 2504 9978
rect 2508 9974 2509 9978
rect 2513 9974 2514 9978
rect 2518 9974 2519 9978
rect 2523 9974 2524 9978
rect 2528 9974 2529 9978
rect 2533 9974 2534 9978
rect 2538 9974 2539 9978
rect 2543 9974 2544 9978
rect 2548 9974 2549 9978
rect 2459 9973 2463 9974
rect 2459 9968 2463 9969
rect 2549 9973 2553 9974
rect 2549 9968 2553 9969
rect 2459 9963 2463 9964
rect 2459 9958 2463 9959
rect 2459 9953 2463 9954
rect 2389 9948 2393 9949
rect 2389 9943 2393 9944
rect 2389 9938 2393 9939
rect 2389 9933 2393 9934
rect 2389 9928 2393 9929
rect 2389 9923 2393 9924
rect 2389 9918 2393 9919
rect 2389 9913 2393 9914
rect 2389 9908 2393 9909
rect 2389 9903 2393 9904
rect 2389 9898 2393 9899
rect 2389 9893 2393 9894
rect 2389 9888 2393 9889
rect 2389 9883 2393 9884
rect 2459 9948 2463 9949
rect 2459 9943 2463 9944
rect 2459 9938 2463 9939
rect 2459 9933 2463 9934
rect 2459 9928 2463 9929
rect 2459 9923 2463 9924
rect 2459 9918 2463 9919
rect 2459 9913 2463 9914
rect 2459 9908 2463 9909
rect 2459 9903 2463 9904
rect 2459 9898 2463 9899
rect 2459 9893 2463 9894
rect 2459 9888 2463 9889
rect 2459 9883 2463 9884
rect 2389 9878 2393 9879
rect 2389 9873 2393 9874
rect 2389 9868 2393 9869
rect 2389 9863 2393 9864
rect 2389 9858 2393 9859
rect 2389 9853 2393 9854
rect 2389 9848 2393 9849
rect 2299 9843 2303 9844
rect 2415 9846 2436 9874
rect 2459 9878 2463 9879
rect 2459 9873 2463 9874
rect 2459 9868 2463 9869
rect 2459 9863 2463 9864
rect 2459 9858 2463 9859
rect 2459 9853 2463 9854
rect 2459 9848 2463 9849
rect 2476 9961 2479 9965
rect 2483 9961 2484 9965
rect 2488 9961 2489 9965
rect 2493 9961 2494 9965
rect 2498 9961 2499 9965
rect 2503 9961 2504 9965
rect 2508 9961 2509 9965
rect 2513 9961 2514 9965
rect 2518 9961 2519 9965
rect 2523 9961 2524 9965
rect 2528 9961 2529 9965
rect 2533 9961 2536 9965
rect 2472 9958 2476 9961
rect 2472 9953 2476 9954
rect 2536 9958 2540 9961
rect 2536 9953 2540 9954
rect 2472 9948 2476 9949
rect 2472 9943 2476 9944
rect 2472 9938 2476 9939
rect 2472 9933 2476 9934
rect 2472 9928 2476 9929
rect 2472 9923 2476 9924
rect 2472 9918 2476 9919
rect 2472 9913 2476 9914
rect 2472 9908 2476 9909
rect 2472 9903 2476 9904
rect 2472 9898 2476 9899
rect 2472 9893 2476 9894
rect 2472 9888 2476 9889
rect 2472 9883 2476 9884
rect 2472 9878 2476 9879
rect 2472 9873 2476 9874
rect 2472 9868 2476 9869
rect 2483 9949 2484 9953
rect 2488 9949 2489 9953
rect 2493 9949 2494 9953
rect 2498 9949 2499 9953
rect 2503 9949 2504 9953
rect 2508 9949 2509 9953
rect 2513 9949 2514 9953
rect 2518 9949 2519 9953
rect 2523 9949 2524 9953
rect 2483 9948 2528 9949
rect 2483 9944 2484 9948
rect 2488 9944 2489 9948
rect 2493 9944 2494 9948
rect 2498 9944 2499 9948
rect 2503 9944 2504 9948
rect 2508 9944 2509 9948
rect 2513 9944 2514 9948
rect 2518 9944 2519 9948
rect 2523 9944 2524 9948
rect 2483 9943 2528 9944
rect 2483 9939 2484 9943
rect 2488 9939 2489 9943
rect 2493 9939 2494 9943
rect 2498 9939 2499 9943
rect 2503 9939 2504 9943
rect 2508 9939 2509 9943
rect 2513 9939 2514 9943
rect 2518 9939 2519 9943
rect 2523 9939 2524 9943
rect 2483 9938 2528 9939
rect 2483 9934 2484 9938
rect 2488 9934 2489 9938
rect 2493 9934 2494 9938
rect 2498 9934 2499 9938
rect 2503 9934 2504 9938
rect 2508 9934 2509 9938
rect 2513 9934 2514 9938
rect 2518 9934 2519 9938
rect 2523 9934 2524 9938
rect 2483 9933 2528 9934
rect 2483 9929 2484 9933
rect 2488 9929 2489 9933
rect 2493 9929 2494 9933
rect 2498 9929 2499 9933
rect 2503 9929 2504 9933
rect 2508 9929 2509 9933
rect 2513 9929 2514 9933
rect 2518 9929 2519 9933
rect 2523 9929 2524 9933
rect 2483 9928 2528 9929
rect 2483 9924 2484 9928
rect 2488 9924 2489 9928
rect 2493 9924 2494 9928
rect 2498 9924 2499 9928
rect 2503 9924 2504 9928
rect 2508 9924 2509 9928
rect 2513 9924 2514 9928
rect 2518 9924 2519 9928
rect 2523 9924 2524 9928
rect 2483 9923 2528 9924
rect 2483 9919 2484 9923
rect 2488 9919 2489 9923
rect 2493 9919 2494 9923
rect 2498 9919 2499 9923
rect 2503 9919 2504 9923
rect 2508 9919 2509 9923
rect 2513 9919 2514 9923
rect 2518 9919 2519 9923
rect 2523 9919 2524 9923
rect 2483 9918 2528 9919
rect 2483 9914 2484 9918
rect 2488 9914 2489 9918
rect 2493 9914 2494 9918
rect 2498 9914 2499 9918
rect 2503 9914 2504 9918
rect 2508 9914 2509 9918
rect 2513 9914 2514 9918
rect 2518 9914 2519 9918
rect 2523 9914 2524 9918
rect 2483 9913 2528 9914
rect 2483 9909 2484 9913
rect 2488 9909 2489 9913
rect 2493 9909 2494 9913
rect 2498 9909 2499 9913
rect 2503 9909 2504 9913
rect 2508 9909 2509 9913
rect 2513 9909 2514 9913
rect 2518 9909 2519 9913
rect 2523 9909 2524 9913
rect 2483 9908 2528 9909
rect 2483 9904 2484 9908
rect 2488 9904 2489 9908
rect 2493 9904 2494 9908
rect 2498 9904 2499 9908
rect 2503 9904 2504 9908
rect 2508 9904 2509 9908
rect 2513 9904 2514 9908
rect 2518 9904 2519 9908
rect 2523 9904 2524 9908
rect 2483 9903 2528 9904
rect 2483 9899 2484 9903
rect 2488 9899 2489 9903
rect 2493 9899 2494 9903
rect 2498 9899 2499 9903
rect 2503 9899 2504 9903
rect 2508 9899 2509 9903
rect 2513 9899 2514 9903
rect 2518 9899 2519 9903
rect 2523 9899 2524 9903
rect 2483 9898 2528 9899
rect 2483 9894 2484 9898
rect 2488 9894 2489 9898
rect 2493 9894 2494 9898
rect 2498 9894 2499 9898
rect 2503 9894 2504 9898
rect 2508 9894 2509 9898
rect 2513 9894 2514 9898
rect 2518 9894 2519 9898
rect 2523 9894 2524 9898
rect 2483 9893 2528 9894
rect 2483 9889 2484 9893
rect 2488 9889 2489 9893
rect 2493 9889 2494 9893
rect 2498 9889 2499 9893
rect 2503 9889 2504 9893
rect 2508 9889 2509 9893
rect 2513 9889 2514 9893
rect 2518 9889 2519 9893
rect 2523 9889 2524 9893
rect 2483 9888 2528 9889
rect 2483 9884 2484 9888
rect 2488 9884 2489 9888
rect 2493 9884 2494 9888
rect 2498 9884 2499 9888
rect 2503 9884 2504 9888
rect 2508 9884 2509 9888
rect 2513 9884 2514 9888
rect 2518 9884 2519 9888
rect 2523 9884 2524 9888
rect 2483 9883 2528 9884
rect 2483 9879 2484 9883
rect 2488 9879 2489 9883
rect 2493 9879 2494 9883
rect 2498 9879 2499 9883
rect 2503 9879 2504 9883
rect 2508 9879 2509 9883
rect 2513 9879 2514 9883
rect 2518 9879 2519 9883
rect 2523 9879 2524 9883
rect 2483 9878 2528 9879
rect 2483 9874 2484 9878
rect 2488 9874 2489 9878
rect 2493 9874 2494 9878
rect 2498 9874 2499 9878
rect 2503 9874 2504 9878
rect 2508 9874 2509 9878
rect 2513 9874 2514 9878
rect 2518 9874 2519 9878
rect 2523 9874 2524 9878
rect 2483 9873 2528 9874
rect 2483 9869 2484 9873
rect 2488 9869 2489 9873
rect 2493 9869 2494 9873
rect 2498 9869 2499 9873
rect 2503 9869 2504 9873
rect 2508 9869 2509 9873
rect 2513 9869 2514 9873
rect 2518 9869 2519 9873
rect 2523 9869 2524 9873
rect 2483 9868 2528 9869
rect 2483 9864 2484 9868
rect 2488 9864 2489 9868
rect 2493 9864 2494 9868
rect 2498 9864 2499 9868
rect 2503 9864 2504 9868
rect 2508 9864 2509 9868
rect 2513 9864 2514 9868
rect 2518 9864 2519 9868
rect 2523 9864 2524 9868
rect 2536 9948 2540 9949
rect 2536 9943 2540 9944
rect 2536 9938 2540 9939
rect 2536 9933 2540 9934
rect 2536 9928 2540 9929
rect 2536 9923 2540 9924
rect 2536 9918 2540 9919
rect 2536 9913 2540 9914
rect 2536 9908 2540 9909
rect 2536 9903 2540 9904
rect 2536 9898 2540 9899
rect 2536 9893 2540 9894
rect 2536 9888 2540 9889
rect 2536 9883 2540 9884
rect 2536 9878 2540 9879
rect 2536 9873 2540 9874
rect 2536 9868 2540 9869
rect 2472 9863 2476 9864
rect 2472 9856 2476 9859
rect 2536 9863 2540 9864
rect 2536 9856 2540 9859
rect 2476 9848 2479 9856
rect 2483 9848 2484 9856
rect 2488 9848 2489 9856
rect 2493 9848 2494 9856
rect 2498 9848 2499 9856
rect 2503 9848 2504 9856
rect 2508 9848 2509 9856
rect 2513 9848 2514 9856
rect 2518 9848 2519 9856
rect 2523 9848 2524 9856
rect 2528 9848 2529 9856
rect 2533 9848 2536 9856
rect 2549 9963 2553 9964
rect 2549 9958 2553 9959
rect 2549 9953 2553 9954
rect 2549 9948 2553 9949
rect 2549 9943 2553 9944
rect 2549 9938 2553 9939
rect 2549 9933 2553 9934
rect 2549 9928 2553 9929
rect 2549 9923 2553 9924
rect 2549 9918 2553 9919
rect 2549 9913 2553 9914
rect 2549 9908 2553 9909
rect 2549 9903 2553 9904
rect 2549 9898 2553 9899
rect 2549 9893 2553 9894
rect 2549 9888 2553 9889
rect 2549 9883 2553 9884
rect 2549 9878 2553 9879
rect 2549 9873 2553 9874
rect 2549 9868 2553 9869
rect 2549 9863 2553 9864
rect 2549 9858 2553 9859
rect 2549 9853 2553 9854
rect 2549 9848 2553 9849
rect 2417 9844 2434 9846
rect 2389 9843 2393 9844
rect 2303 9839 2304 9843
rect 2308 9839 2309 9843
rect 2313 9839 2314 9843
rect 2318 9839 2319 9843
rect 2323 9839 2324 9843
rect 2328 9839 2329 9843
rect 2333 9839 2334 9843
rect 2338 9839 2339 9843
rect 2343 9839 2344 9843
rect 2348 9839 2349 9843
rect 2353 9839 2354 9843
rect 2358 9839 2359 9843
rect 2363 9839 2364 9843
rect 2368 9839 2369 9843
rect 2373 9839 2374 9843
rect 2378 9839 2379 9843
rect 2383 9839 2384 9843
rect 2388 9839 2389 9843
rect 2419 9842 2432 9844
rect 2459 9843 2463 9844
rect 2549 9843 2553 9844
rect 2187 9831 2243 9839
rect 1993 9827 2052 9831
rect 2178 9827 2243 9831
rect 1993 9815 2049 9827
rect 2108 9819 2138 9823
rect 1993 9811 2052 9815
rect 2122 9812 2126 9819
rect 2187 9815 2243 9827
rect 1993 9802 2049 9811
rect 2178 9811 2243 9815
rect 2108 9803 2119 9807
rect 1869 9795 1934 9799
rect 1672 9790 1740 9791
rect 1672 9786 1673 9790
rect 1677 9786 1678 9790
rect 1682 9786 1740 9790
rect 1799 9787 1829 9791
rect 1672 9785 1740 9786
rect 1672 9781 1673 9785
rect 1677 9781 1678 9785
rect 1682 9783 1740 9785
rect 1682 9781 1743 9783
rect 1672 9780 1743 9781
rect 1672 9776 1673 9780
rect 1677 9776 1678 9780
rect 1682 9779 1743 9780
rect 1682 9776 1740 9779
rect 1672 9775 1740 9776
rect 1672 9771 1673 9775
rect 1677 9771 1678 9775
rect 1682 9771 1740 9775
rect 1672 9770 1740 9771
rect 1672 9766 1673 9770
rect 1677 9766 1678 9770
rect 1682 9766 1740 9770
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1628 9761 1647 9762
rect 1632 9757 1633 9761
rect 1637 9757 1638 9761
rect 1642 9757 1643 9761
rect 1628 9756 1647 9757
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1628 9751 1647 9752
rect 1632 9747 1633 9751
rect 1637 9747 1638 9751
rect 1642 9747 1643 9751
rect 1628 9746 1647 9747
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1628 9741 1647 9742
rect 1632 9737 1633 9741
rect 1637 9737 1638 9741
rect 1642 9737 1643 9741
rect 1628 9736 1647 9737
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1672 9765 1740 9766
rect 1672 9761 1673 9765
rect 1677 9761 1678 9765
rect 1682 9761 1740 9765
rect 1672 9760 1740 9761
rect 1672 9756 1673 9760
rect 1677 9756 1678 9760
rect 1682 9756 1740 9760
rect 1672 9755 1740 9756
rect 1672 9751 1673 9755
rect 1677 9751 1678 9755
rect 1682 9751 1740 9755
rect 1672 9750 1740 9751
rect 1672 9746 1673 9750
rect 1677 9746 1678 9750
rect 1682 9746 1740 9750
rect 1672 9745 1740 9746
rect 1672 9741 1673 9745
rect 1677 9741 1678 9745
rect 1682 9741 1740 9745
rect 1672 9740 1740 9741
rect 1672 9736 1673 9740
rect 1677 9736 1678 9740
rect 1682 9736 1740 9740
rect 1672 9734 1740 9736
rect 1573 9718 1574 9722
rect 1578 9718 1579 9722
rect 1583 9718 1584 9722
rect 1588 9718 1589 9722
rect 1593 9718 1594 9722
rect 1598 9718 1599 9722
rect 1603 9718 1604 9722
rect 1608 9718 1609 9722
rect 1613 9718 1614 9722
rect 1618 9718 1619 9722
rect 1623 9718 1625 9722
rect 1569 9717 1625 9718
rect 1573 9713 1574 9717
rect 1578 9713 1579 9717
rect 1583 9713 1584 9717
rect 1588 9713 1589 9717
rect 1593 9713 1594 9717
rect 1598 9713 1599 9717
rect 1603 9713 1604 9717
rect 1608 9713 1609 9717
rect 1613 9713 1614 9717
rect 1618 9713 1619 9717
rect 1623 9713 1625 9717
rect 1569 9712 1625 9713
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1628 9715 1647 9716
rect 1473 9710 1525 9711
rect 1473 9706 1499 9710
rect 1503 9706 1504 9710
rect 1508 9706 1525 9710
rect 1473 9705 1525 9706
rect 1473 9701 1499 9705
rect 1503 9701 1504 9705
rect 1508 9701 1525 9705
rect 1473 9700 1525 9701
rect 1473 9696 1499 9700
rect 1503 9696 1504 9700
rect 1508 9696 1525 9700
rect 1473 9695 1525 9696
rect 1473 9691 1499 9695
rect 1503 9691 1504 9695
rect 1508 9691 1525 9695
rect 1473 9690 1525 9691
rect 1473 9686 1499 9690
rect 1503 9686 1504 9690
rect 1508 9686 1525 9690
rect 1632 9711 1633 9715
rect 1637 9711 1638 9715
rect 1642 9711 1643 9715
rect 1628 9710 1647 9711
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1628 9705 1647 9706
rect 1632 9701 1633 9705
rect 1637 9701 1638 9705
rect 1642 9701 1643 9705
rect 1628 9700 1647 9701
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1628 9695 1647 9696
rect 1632 9691 1633 9695
rect 1637 9691 1638 9695
rect 1642 9691 1643 9695
rect 1628 9690 1647 9691
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1473 9685 1525 9686
rect 1473 9681 1499 9685
rect 1503 9681 1504 9685
rect 1508 9681 1525 9685
rect 1473 9680 1525 9681
rect 1473 9676 1499 9680
rect 1503 9676 1504 9680
rect 1508 9676 1525 9680
rect 1473 9675 1525 9676
rect 1473 9671 1499 9675
rect 1503 9671 1504 9675
rect 1508 9671 1525 9675
rect 1473 9670 1525 9671
rect 1473 9666 1499 9670
rect 1503 9666 1504 9670
rect 1508 9666 1525 9670
rect 1473 9665 1525 9666
rect 1473 9661 1499 9665
rect 1503 9661 1504 9665
rect 1508 9661 1525 9665
rect 1473 9610 1525 9661
rect 659 9607 693 9608
rect 663 9603 664 9607
rect 668 9603 669 9607
rect 673 9603 674 9607
rect 678 9603 679 9607
rect 683 9603 684 9607
rect 688 9603 689 9607
rect 617 9592 618 9596
rect 622 9592 623 9596
rect 627 9592 628 9596
rect 632 9592 633 9596
rect 637 9592 638 9596
rect 642 9592 643 9596
rect 613 9591 647 9592
rect 617 9587 618 9591
rect 622 9587 623 9591
rect 627 9587 628 9591
rect 632 9587 633 9591
rect 637 9587 638 9591
rect 642 9587 643 9591
rect 613 9586 647 9587
rect 617 9582 618 9586
rect 622 9582 623 9586
rect 627 9582 628 9586
rect 632 9582 633 9586
rect 637 9582 638 9586
rect 642 9582 643 9586
rect 613 9581 647 9582
rect 617 9577 618 9581
rect 622 9577 623 9581
rect 627 9577 628 9581
rect 632 9577 633 9581
rect 637 9577 638 9581
rect 642 9577 643 9581
rect 663 9592 664 9596
rect 668 9592 669 9596
rect 673 9592 674 9596
rect 678 9592 679 9596
rect 683 9592 684 9596
rect 688 9592 689 9596
rect 1804 9593 1817 9787
rect 1878 9783 1934 9795
rect 1869 9779 1934 9783
rect 1878 9722 1934 9779
rect 1981 9800 2049 9802
rect 1981 9796 1982 9800
rect 1986 9796 1987 9800
rect 1991 9799 2049 9800
rect 2112 9800 2119 9803
rect 2131 9803 2138 9807
rect 2131 9800 2135 9803
rect 1991 9796 2052 9799
rect 1981 9795 2052 9796
rect 1981 9791 1982 9795
rect 1986 9791 1987 9795
rect 1991 9791 2049 9795
rect 2112 9791 2135 9800
rect 2187 9799 2243 9811
rect 2302 9831 2358 9839
rect 2421 9831 2430 9842
rect 2463 9839 2464 9843
rect 2468 9839 2469 9843
rect 2473 9839 2474 9843
rect 2478 9839 2479 9843
rect 2483 9839 2484 9843
rect 2488 9839 2489 9843
rect 2493 9839 2494 9843
rect 2498 9839 2499 9843
rect 2503 9839 2504 9843
rect 2508 9839 2509 9843
rect 2513 9839 2514 9843
rect 2518 9839 2519 9843
rect 2523 9839 2524 9843
rect 2528 9839 2529 9843
rect 2533 9839 2534 9843
rect 2538 9839 2539 9843
rect 2543 9839 2544 9843
rect 2548 9839 2549 9843
rect 2612 9974 2613 9978
rect 2617 9974 2618 9978
rect 2622 9974 2623 9978
rect 2627 9974 2628 9978
rect 2632 9974 2633 9978
rect 2637 9974 2638 9978
rect 2642 9974 2643 9978
rect 2647 9974 2648 9978
rect 2652 9974 2653 9978
rect 2657 9974 2658 9978
rect 2662 9974 2663 9978
rect 2667 9974 2668 9978
rect 2672 9974 2673 9978
rect 2677 9974 2678 9978
rect 2682 9974 2683 9978
rect 2687 9974 2688 9978
rect 2692 9974 2693 9978
rect 2697 9974 2698 9978
rect 2608 9973 2612 9974
rect 2608 9968 2612 9969
rect 2698 9973 2702 9974
rect 2698 9968 2702 9969
rect 2608 9963 2612 9964
rect 2608 9958 2612 9959
rect 2608 9953 2612 9954
rect 2608 9948 2612 9949
rect 2608 9943 2612 9944
rect 2608 9938 2612 9939
rect 2608 9933 2612 9934
rect 2608 9928 2612 9929
rect 2608 9923 2612 9924
rect 2608 9918 2612 9919
rect 2608 9913 2612 9914
rect 2608 9908 2612 9909
rect 2608 9903 2612 9904
rect 2608 9898 2612 9899
rect 2608 9893 2612 9894
rect 2608 9888 2612 9889
rect 2608 9883 2612 9884
rect 2608 9878 2612 9879
rect 2608 9873 2612 9874
rect 2608 9868 2612 9869
rect 2608 9863 2612 9864
rect 2608 9858 2612 9859
rect 2608 9853 2612 9854
rect 2608 9848 2612 9849
rect 2625 9961 2628 9965
rect 2632 9961 2633 9965
rect 2637 9961 2638 9965
rect 2642 9961 2643 9965
rect 2647 9961 2648 9965
rect 2652 9961 2653 9965
rect 2657 9961 2658 9965
rect 2662 9961 2663 9965
rect 2667 9961 2668 9965
rect 2672 9961 2673 9965
rect 2677 9961 2678 9965
rect 2682 9961 2685 9965
rect 2621 9958 2625 9961
rect 2621 9953 2625 9954
rect 2685 9958 2689 9961
rect 2685 9953 2689 9954
rect 2621 9948 2625 9949
rect 2621 9943 2625 9944
rect 2621 9938 2625 9939
rect 2621 9933 2625 9934
rect 2621 9928 2625 9929
rect 2621 9923 2625 9924
rect 2621 9918 2625 9919
rect 2621 9913 2625 9914
rect 2621 9908 2625 9909
rect 2621 9903 2625 9904
rect 2621 9898 2625 9899
rect 2621 9893 2625 9894
rect 2621 9888 2625 9889
rect 2621 9883 2625 9884
rect 2621 9878 2625 9879
rect 2621 9873 2625 9874
rect 2621 9868 2625 9869
rect 2637 9949 2638 9953
rect 2642 9949 2643 9953
rect 2647 9949 2648 9953
rect 2652 9949 2653 9953
rect 2657 9949 2658 9953
rect 2662 9949 2663 9953
rect 2667 9949 2668 9953
rect 2672 9949 2673 9953
rect 2633 9948 2677 9949
rect 2637 9944 2638 9948
rect 2642 9944 2643 9948
rect 2647 9944 2648 9948
rect 2652 9944 2653 9948
rect 2657 9944 2658 9948
rect 2662 9944 2663 9948
rect 2667 9944 2668 9948
rect 2672 9944 2673 9948
rect 2633 9943 2677 9944
rect 2637 9939 2638 9943
rect 2642 9939 2643 9943
rect 2647 9939 2648 9943
rect 2652 9939 2653 9943
rect 2657 9939 2658 9943
rect 2662 9939 2663 9943
rect 2667 9939 2668 9943
rect 2672 9939 2673 9943
rect 2633 9938 2677 9939
rect 2637 9934 2638 9938
rect 2642 9934 2643 9938
rect 2647 9934 2648 9938
rect 2652 9934 2653 9938
rect 2657 9934 2658 9938
rect 2662 9934 2663 9938
rect 2667 9934 2668 9938
rect 2672 9934 2673 9938
rect 2633 9933 2677 9934
rect 2637 9929 2638 9933
rect 2642 9929 2643 9933
rect 2647 9929 2648 9933
rect 2652 9929 2653 9933
rect 2657 9929 2658 9933
rect 2662 9929 2663 9933
rect 2667 9929 2668 9933
rect 2672 9929 2673 9933
rect 2633 9928 2677 9929
rect 2637 9924 2638 9928
rect 2642 9924 2643 9928
rect 2647 9924 2648 9928
rect 2652 9924 2653 9928
rect 2657 9924 2658 9928
rect 2662 9924 2663 9928
rect 2667 9924 2668 9928
rect 2672 9924 2673 9928
rect 2633 9923 2677 9924
rect 2637 9919 2638 9923
rect 2642 9919 2643 9923
rect 2647 9919 2648 9923
rect 2652 9919 2653 9923
rect 2657 9919 2658 9923
rect 2662 9919 2663 9923
rect 2667 9919 2668 9923
rect 2672 9919 2673 9923
rect 2633 9918 2677 9919
rect 2637 9914 2638 9918
rect 2642 9914 2643 9918
rect 2647 9914 2648 9918
rect 2652 9914 2653 9918
rect 2657 9914 2658 9918
rect 2662 9914 2663 9918
rect 2667 9914 2668 9918
rect 2672 9914 2673 9918
rect 2633 9913 2677 9914
rect 2637 9909 2638 9913
rect 2642 9909 2643 9913
rect 2647 9909 2648 9913
rect 2652 9909 2653 9913
rect 2657 9909 2658 9913
rect 2662 9909 2663 9913
rect 2667 9909 2668 9913
rect 2672 9909 2673 9913
rect 2633 9908 2677 9909
rect 2637 9904 2638 9908
rect 2642 9904 2643 9908
rect 2647 9904 2648 9908
rect 2652 9904 2653 9908
rect 2657 9904 2658 9908
rect 2662 9904 2663 9908
rect 2667 9904 2668 9908
rect 2672 9904 2673 9908
rect 2633 9903 2677 9904
rect 2637 9899 2638 9903
rect 2642 9899 2643 9903
rect 2647 9899 2648 9903
rect 2652 9899 2653 9903
rect 2657 9899 2658 9903
rect 2662 9899 2663 9903
rect 2667 9899 2668 9903
rect 2672 9899 2673 9903
rect 2633 9898 2677 9899
rect 2637 9894 2638 9898
rect 2642 9894 2643 9898
rect 2647 9894 2648 9898
rect 2652 9894 2653 9898
rect 2657 9894 2658 9898
rect 2662 9894 2663 9898
rect 2667 9894 2668 9898
rect 2672 9894 2673 9898
rect 2633 9893 2677 9894
rect 2637 9889 2638 9893
rect 2642 9889 2643 9893
rect 2647 9889 2648 9893
rect 2652 9889 2653 9893
rect 2657 9889 2658 9893
rect 2662 9889 2663 9893
rect 2667 9889 2668 9893
rect 2672 9889 2673 9893
rect 2633 9888 2677 9889
rect 2637 9884 2638 9888
rect 2642 9884 2643 9888
rect 2647 9884 2648 9888
rect 2652 9884 2653 9888
rect 2657 9884 2658 9888
rect 2662 9884 2663 9888
rect 2667 9884 2668 9888
rect 2672 9884 2673 9888
rect 2633 9883 2677 9884
rect 2637 9879 2638 9883
rect 2642 9879 2643 9883
rect 2647 9879 2648 9883
rect 2652 9879 2653 9883
rect 2657 9879 2658 9883
rect 2662 9879 2663 9883
rect 2667 9879 2668 9883
rect 2672 9879 2673 9883
rect 2633 9878 2677 9879
rect 2637 9874 2638 9878
rect 2642 9874 2643 9878
rect 2647 9874 2648 9878
rect 2652 9874 2653 9878
rect 2657 9874 2658 9878
rect 2662 9874 2663 9878
rect 2667 9874 2668 9878
rect 2672 9874 2673 9878
rect 2633 9873 2677 9874
rect 2637 9869 2638 9873
rect 2642 9869 2643 9873
rect 2647 9869 2648 9873
rect 2652 9869 2653 9873
rect 2657 9869 2658 9873
rect 2662 9869 2663 9873
rect 2667 9869 2668 9873
rect 2672 9869 2673 9873
rect 2633 9868 2677 9869
rect 2637 9864 2638 9868
rect 2642 9864 2643 9868
rect 2647 9864 2648 9868
rect 2652 9864 2653 9868
rect 2657 9864 2658 9868
rect 2662 9864 2663 9868
rect 2667 9864 2668 9868
rect 2672 9864 2673 9868
rect 2685 9948 2689 9949
rect 2685 9943 2689 9944
rect 2685 9938 2689 9939
rect 2685 9933 2689 9934
rect 2685 9928 2689 9929
rect 2685 9923 2689 9924
rect 2685 9918 2689 9919
rect 2685 9913 2689 9914
rect 2685 9908 2689 9909
rect 2685 9903 2689 9904
rect 2685 9898 2689 9899
rect 2685 9893 2689 9894
rect 2685 9888 2689 9889
rect 2685 9883 2689 9884
rect 2685 9878 2689 9879
rect 2685 9873 2689 9874
rect 2685 9868 2689 9869
rect 2621 9863 2625 9864
rect 2621 9856 2625 9859
rect 2685 9863 2689 9864
rect 2685 9856 2689 9859
rect 2625 9848 2628 9856
rect 2632 9848 2633 9856
rect 2637 9848 2638 9856
rect 2642 9848 2643 9856
rect 2647 9848 2648 9856
rect 2652 9848 2653 9856
rect 2657 9848 2658 9856
rect 2662 9848 2663 9856
rect 2667 9848 2668 9856
rect 2672 9848 2673 9856
rect 2677 9848 2678 9856
rect 2682 9848 2685 9856
rect 2698 9963 2702 9964
rect 2698 9958 2702 9959
rect 2698 9953 2702 9954
rect 2724 9961 2745 9981
rect 2772 9974 2773 9978
rect 2777 9974 2778 9978
rect 2782 9974 2783 9978
rect 2787 9974 2788 9978
rect 2792 9974 2793 9978
rect 2797 9974 2798 9978
rect 2802 9974 2803 9978
rect 2807 9974 2808 9978
rect 2812 9974 2813 9978
rect 2817 9974 2818 9978
rect 2822 9974 2823 9978
rect 2827 9974 2828 9978
rect 2832 9974 2833 9978
rect 2837 9974 2838 9978
rect 2842 9974 2843 9978
rect 2847 9974 2848 9978
rect 2852 9974 2853 9978
rect 2857 9974 2858 9978
rect 2768 9973 2772 9974
rect 2768 9968 2772 9969
rect 2858 9973 2862 9974
rect 2858 9968 2862 9969
rect 2768 9963 2772 9964
rect 2768 9958 2772 9959
rect 2768 9953 2772 9954
rect 2698 9948 2702 9949
rect 2698 9943 2702 9944
rect 2698 9938 2702 9939
rect 2698 9933 2702 9934
rect 2698 9928 2702 9929
rect 2698 9923 2702 9924
rect 2698 9918 2702 9919
rect 2698 9913 2702 9914
rect 2698 9908 2702 9909
rect 2698 9903 2702 9904
rect 2698 9898 2702 9899
rect 2698 9893 2702 9894
rect 2698 9888 2702 9889
rect 2698 9883 2702 9884
rect 2768 9948 2772 9949
rect 2768 9943 2772 9944
rect 2768 9938 2772 9939
rect 2768 9933 2772 9934
rect 2768 9928 2772 9929
rect 2768 9923 2772 9924
rect 2768 9918 2772 9919
rect 2768 9913 2772 9914
rect 2768 9908 2772 9909
rect 2768 9903 2772 9904
rect 2768 9898 2772 9899
rect 2768 9893 2772 9894
rect 2768 9888 2772 9889
rect 2768 9883 2772 9884
rect 2698 9878 2702 9879
rect 2698 9873 2702 9874
rect 2698 9868 2702 9869
rect 2698 9863 2702 9864
rect 2698 9858 2702 9859
rect 2698 9853 2702 9854
rect 2698 9848 2702 9849
rect 2608 9843 2612 9844
rect 2724 9846 2745 9874
rect 2768 9878 2772 9879
rect 2768 9873 2772 9874
rect 2768 9868 2772 9869
rect 2768 9863 2772 9864
rect 2768 9858 2772 9859
rect 2768 9853 2772 9854
rect 2768 9848 2772 9849
rect 2785 9961 2788 9965
rect 2792 9961 2793 9965
rect 2797 9961 2798 9965
rect 2802 9961 2803 9965
rect 2807 9961 2808 9965
rect 2812 9961 2813 9965
rect 2817 9961 2818 9965
rect 2822 9961 2823 9965
rect 2827 9961 2828 9965
rect 2832 9961 2833 9965
rect 2837 9961 2838 9965
rect 2842 9961 2845 9965
rect 2781 9958 2785 9961
rect 2781 9953 2785 9954
rect 2845 9958 2849 9961
rect 2845 9953 2849 9954
rect 2781 9948 2785 9949
rect 2781 9943 2785 9944
rect 2781 9938 2785 9939
rect 2781 9933 2785 9934
rect 2781 9928 2785 9929
rect 2781 9923 2785 9924
rect 2781 9918 2785 9919
rect 2781 9913 2785 9914
rect 2781 9908 2785 9909
rect 2781 9903 2785 9904
rect 2781 9898 2785 9899
rect 2781 9893 2785 9894
rect 2781 9888 2785 9889
rect 2781 9883 2785 9884
rect 2781 9878 2785 9879
rect 2781 9873 2785 9874
rect 2781 9868 2785 9869
rect 2792 9949 2793 9953
rect 2797 9949 2798 9953
rect 2802 9949 2803 9953
rect 2807 9949 2808 9953
rect 2812 9949 2813 9953
rect 2817 9949 2818 9953
rect 2822 9949 2823 9953
rect 2827 9949 2828 9953
rect 2832 9949 2833 9953
rect 2792 9948 2837 9949
rect 2792 9944 2793 9948
rect 2797 9944 2798 9948
rect 2802 9944 2803 9948
rect 2807 9944 2808 9948
rect 2812 9944 2813 9948
rect 2817 9944 2818 9948
rect 2822 9944 2823 9948
rect 2827 9944 2828 9948
rect 2832 9944 2833 9948
rect 2792 9943 2837 9944
rect 2792 9939 2793 9943
rect 2797 9939 2798 9943
rect 2802 9939 2803 9943
rect 2807 9939 2808 9943
rect 2812 9939 2813 9943
rect 2817 9939 2818 9943
rect 2822 9939 2823 9943
rect 2827 9939 2828 9943
rect 2832 9939 2833 9943
rect 2792 9938 2837 9939
rect 2792 9934 2793 9938
rect 2797 9934 2798 9938
rect 2802 9934 2803 9938
rect 2807 9934 2808 9938
rect 2812 9934 2813 9938
rect 2817 9934 2818 9938
rect 2822 9934 2823 9938
rect 2827 9934 2828 9938
rect 2832 9934 2833 9938
rect 2792 9933 2837 9934
rect 2792 9929 2793 9933
rect 2797 9929 2798 9933
rect 2802 9929 2803 9933
rect 2807 9929 2808 9933
rect 2812 9929 2813 9933
rect 2817 9929 2818 9933
rect 2822 9929 2823 9933
rect 2827 9929 2828 9933
rect 2832 9929 2833 9933
rect 2792 9928 2837 9929
rect 2792 9924 2793 9928
rect 2797 9924 2798 9928
rect 2802 9924 2803 9928
rect 2807 9924 2808 9928
rect 2812 9924 2813 9928
rect 2817 9924 2818 9928
rect 2822 9924 2823 9928
rect 2827 9924 2828 9928
rect 2832 9924 2833 9928
rect 2792 9923 2837 9924
rect 2792 9919 2793 9923
rect 2797 9919 2798 9923
rect 2802 9919 2803 9923
rect 2807 9919 2808 9923
rect 2812 9919 2813 9923
rect 2817 9919 2818 9923
rect 2822 9919 2823 9923
rect 2827 9919 2828 9923
rect 2832 9919 2833 9923
rect 2792 9918 2837 9919
rect 2792 9914 2793 9918
rect 2797 9914 2798 9918
rect 2802 9914 2803 9918
rect 2807 9914 2808 9918
rect 2812 9914 2813 9918
rect 2817 9914 2818 9918
rect 2822 9914 2823 9918
rect 2827 9914 2828 9918
rect 2832 9914 2833 9918
rect 2792 9913 2837 9914
rect 2792 9909 2793 9913
rect 2797 9909 2798 9913
rect 2802 9909 2803 9913
rect 2807 9909 2808 9913
rect 2812 9909 2813 9913
rect 2817 9909 2818 9913
rect 2822 9909 2823 9913
rect 2827 9909 2828 9913
rect 2832 9909 2833 9913
rect 2792 9908 2837 9909
rect 2792 9904 2793 9908
rect 2797 9904 2798 9908
rect 2802 9904 2803 9908
rect 2807 9904 2808 9908
rect 2812 9904 2813 9908
rect 2817 9904 2818 9908
rect 2822 9904 2823 9908
rect 2827 9904 2828 9908
rect 2832 9904 2833 9908
rect 2792 9903 2837 9904
rect 2792 9899 2793 9903
rect 2797 9899 2798 9903
rect 2802 9899 2803 9903
rect 2807 9899 2808 9903
rect 2812 9899 2813 9903
rect 2817 9899 2818 9903
rect 2822 9899 2823 9903
rect 2827 9899 2828 9903
rect 2832 9899 2833 9903
rect 2792 9898 2837 9899
rect 2792 9894 2793 9898
rect 2797 9894 2798 9898
rect 2802 9894 2803 9898
rect 2807 9894 2808 9898
rect 2812 9894 2813 9898
rect 2817 9894 2818 9898
rect 2822 9894 2823 9898
rect 2827 9894 2828 9898
rect 2832 9894 2833 9898
rect 2792 9893 2837 9894
rect 2792 9889 2793 9893
rect 2797 9889 2798 9893
rect 2802 9889 2803 9893
rect 2807 9889 2808 9893
rect 2812 9889 2813 9893
rect 2817 9889 2818 9893
rect 2822 9889 2823 9893
rect 2827 9889 2828 9893
rect 2832 9889 2833 9893
rect 2792 9888 2837 9889
rect 2792 9884 2793 9888
rect 2797 9884 2798 9888
rect 2802 9884 2803 9888
rect 2807 9884 2808 9888
rect 2812 9884 2813 9888
rect 2817 9884 2818 9888
rect 2822 9884 2823 9888
rect 2827 9884 2828 9888
rect 2832 9884 2833 9888
rect 2792 9883 2837 9884
rect 2792 9879 2793 9883
rect 2797 9879 2798 9883
rect 2802 9879 2803 9883
rect 2807 9879 2808 9883
rect 2812 9879 2813 9883
rect 2817 9879 2818 9883
rect 2822 9879 2823 9883
rect 2827 9879 2828 9883
rect 2832 9879 2833 9883
rect 2792 9878 2837 9879
rect 2792 9874 2793 9878
rect 2797 9874 2798 9878
rect 2802 9874 2803 9878
rect 2807 9874 2808 9878
rect 2812 9874 2813 9878
rect 2817 9874 2818 9878
rect 2822 9874 2823 9878
rect 2827 9874 2828 9878
rect 2832 9874 2833 9878
rect 2792 9873 2837 9874
rect 2792 9869 2793 9873
rect 2797 9869 2798 9873
rect 2802 9869 2803 9873
rect 2807 9869 2808 9873
rect 2812 9869 2813 9873
rect 2817 9869 2818 9873
rect 2822 9869 2823 9873
rect 2827 9869 2828 9873
rect 2832 9869 2833 9873
rect 2792 9868 2837 9869
rect 2792 9864 2793 9868
rect 2797 9864 2798 9868
rect 2802 9864 2803 9868
rect 2807 9864 2808 9868
rect 2812 9864 2813 9868
rect 2817 9864 2818 9868
rect 2822 9864 2823 9868
rect 2827 9864 2828 9868
rect 2832 9864 2833 9868
rect 2845 9948 2849 9949
rect 2845 9943 2849 9944
rect 2845 9938 2849 9939
rect 2845 9933 2849 9934
rect 2845 9928 2849 9929
rect 2845 9923 2849 9924
rect 2845 9918 2849 9919
rect 2845 9913 2849 9914
rect 2845 9908 2849 9909
rect 2845 9903 2849 9904
rect 2845 9898 2849 9899
rect 2845 9893 2849 9894
rect 2845 9888 2849 9889
rect 2845 9883 2849 9884
rect 2845 9878 2849 9879
rect 2845 9873 2849 9874
rect 2845 9868 2849 9869
rect 2781 9863 2785 9864
rect 2781 9856 2785 9859
rect 2845 9863 2849 9864
rect 2845 9856 2849 9859
rect 2785 9848 2788 9856
rect 2792 9848 2793 9856
rect 2797 9848 2798 9856
rect 2802 9848 2803 9856
rect 2807 9848 2808 9856
rect 2812 9848 2813 9856
rect 2817 9848 2818 9856
rect 2822 9848 2823 9856
rect 2827 9848 2828 9856
rect 2832 9848 2833 9856
rect 2837 9848 2838 9856
rect 2842 9848 2845 9856
rect 2858 9963 2862 9964
rect 2858 9958 2862 9959
rect 2858 9953 2862 9954
rect 2858 9948 2862 9949
rect 2858 9943 2862 9944
rect 2858 9938 2862 9939
rect 2858 9933 2862 9934
rect 2858 9928 2862 9929
rect 2858 9923 2862 9924
rect 2858 9918 2862 9919
rect 2858 9913 2862 9914
rect 2858 9908 2862 9909
rect 2858 9903 2862 9904
rect 2858 9898 2862 9899
rect 2858 9893 2862 9894
rect 2858 9888 2862 9889
rect 2858 9883 2862 9884
rect 2858 9878 2862 9879
rect 2858 9873 2862 9874
rect 2858 9868 2862 9869
rect 2858 9863 2862 9864
rect 2858 9858 2862 9859
rect 2858 9853 2862 9854
rect 2858 9848 2862 9849
rect 2726 9844 2743 9846
rect 2698 9843 2702 9844
rect 2612 9839 2613 9843
rect 2617 9839 2618 9843
rect 2622 9839 2623 9843
rect 2627 9839 2628 9843
rect 2632 9839 2633 9843
rect 2637 9839 2638 9843
rect 2642 9839 2643 9843
rect 2647 9839 2648 9843
rect 2652 9839 2653 9843
rect 2657 9839 2658 9843
rect 2662 9839 2663 9843
rect 2667 9839 2668 9843
rect 2672 9839 2673 9843
rect 2677 9839 2678 9843
rect 2682 9839 2683 9843
rect 2687 9839 2688 9843
rect 2692 9839 2693 9843
rect 2697 9839 2698 9843
rect 2728 9842 2741 9844
rect 2768 9843 2772 9844
rect 2858 9843 2862 9844
rect 2496 9831 2552 9839
rect 2302 9827 2361 9831
rect 2487 9827 2552 9831
rect 2302 9815 2358 9827
rect 2417 9819 2447 9823
rect 2302 9811 2361 9815
rect 2431 9812 2435 9819
rect 2496 9815 2552 9827
rect 2302 9802 2358 9811
rect 2487 9811 2552 9815
rect 2417 9803 2428 9807
rect 2178 9795 2243 9799
rect 1981 9790 2049 9791
rect 1981 9786 1982 9790
rect 1986 9786 1987 9790
rect 1991 9786 2049 9790
rect 2108 9787 2138 9791
rect 1981 9785 2049 9786
rect 1981 9781 1982 9785
rect 1986 9781 1987 9785
rect 1991 9783 2049 9785
rect 1991 9781 2052 9783
rect 1981 9780 2052 9781
rect 1981 9776 1982 9780
rect 1986 9776 1987 9780
rect 1991 9779 2052 9780
rect 1991 9776 2049 9779
rect 1981 9775 2049 9776
rect 1981 9771 1982 9775
rect 1986 9771 1987 9775
rect 1991 9771 2049 9775
rect 1981 9770 2049 9771
rect 1981 9766 1982 9770
rect 1986 9766 1987 9770
rect 1991 9766 2049 9770
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1937 9761 1956 9762
rect 1941 9757 1942 9761
rect 1946 9757 1947 9761
rect 1951 9757 1952 9761
rect 1937 9756 1956 9757
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1937 9751 1956 9752
rect 1941 9747 1942 9751
rect 1946 9747 1947 9751
rect 1951 9747 1952 9751
rect 1937 9746 1956 9747
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1937 9741 1956 9742
rect 1941 9737 1942 9741
rect 1946 9737 1947 9741
rect 1951 9737 1952 9741
rect 1937 9736 1956 9737
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1981 9765 2049 9766
rect 1981 9761 1982 9765
rect 1986 9761 1987 9765
rect 1991 9761 2049 9765
rect 1981 9760 2049 9761
rect 1981 9756 1982 9760
rect 1986 9756 1987 9760
rect 1991 9756 2049 9760
rect 1981 9755 2049 9756
rect 1981 9751 1982 9755
rect 1986 9751 1987 9755
rect 1991 9751 2049 9755
rect 1981 9750 2049 9751
rect 1981 9746 1982 9750
rect 1986 9746 1987 9750
rect 1991 9746 2049 9750
rect 1981 9745 2049 9746
rect 1981 9741 1982 9745
rect 1986 9741 1987 9745
rect 1991 9741 2049 9745
rect 1981 9740 2049 9741
rect 1981 9736 1982 9740
rect 1986 9736 1987 9740
rect 1991 9736 2049 9740
rect 1981 9734 2049 9736
rect 1882 9718 1883 9722
rect 1887 9718 1888 9722
rect 1892 9718 1893 9722
rect 1897 9718 1898 9722
rect 1902 9718 1903 9722
rect 1907 9718 1908 9722
rect 1912 9718 1913 9722
rect 1917 9718 1918 9722
rect 1922 9718 1923 9722
rect 1927 9718 1928 9722
rect 1932 9718 1934 9722
rect 1878 9717 1934 9718
rect 1882 9713 1883 9717
rect 1887 9713 1888 9717
rect 1892 9713 1893 9717
rect 1897 9713 1898 9717
rect 1902 9713 1903 9717
rect 1907 9713 1908 9717
rect 1912 9713 1913 9717
rect 1917 9713 1918 9717
rect 1922 9713 1923 9717
rect 1927 9713 1928 9717
rect 1932 9713 1934 9717
rect 1878 9712 1934 9713
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1937 9715 1956 9716
rect 1941 9711 1942 9715
rect 1946 9711 1947 9715
rect 1951 9711 1952 9715
rect 1937 9710 1956 9711
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1937 9705 1956 9706
rect 1941 9701 1942 9705
rect 1946 9701 1947 9705
rect 1951 9701 1952 9705
rect 1937 9700 1956 9701
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1937 9695 1956 9696
rect 1941 9691 1942 9695
rect 1946 9691 1947 9695
rect 1951 9691 1952 9695
rect 1937 9690 1956 9691
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 2113 9597 2126 9787
rect 2187 9783 2243 9795
rect 2178 9779 2243 9783
rect 2187 9722 2243 9779
rect 2290 9800 2358 9802
rect 2290 9796 2291 9800
rect 2295 9796 2296 9800
rect 2300 9799 2358 9800
rect 2421 9800 2428 9803
rect 2440 9803 2447 9807
rect 2440 9800 2444 9803
rect 2300 9796 2361 9799
rect 2290 9795 2361 9796
rect 2290 9791 2291 9795
rect 2295 9791 2296 9795
rect 2300 9791 2358 9795
rect 2421 9791 2444 9800
rect 2496 9799 2552 9811
rect 2611 9831 2667 9839
rect 2730 9831 2739 9842
rect 2772 9839 2773 9843
rect 2777 9839 2778 9843
rect 2782 9839 2783 9843
rect 2787 9839 2788 9843
rect 2792 9839 2793 9843
rect 2797 9839 2798 9843
rect 2802 9839 2803 9843
rect 2807 9839 2808 9843
rect 2812 9839 2813 9843
rect 2817 9839 2818 9843
rect 2822 9839 2823 9843
rect 2827 9839 2828 9843
rect 2832 9839 2833 9843
rect 2837 9839 2838 9843
rect 2842 9839 2843 9843
rect 2847 9839 2848 9843
rect 2852 9839 2853 9843
rect 2857 9839 2858 9843
rect 2921 9974 2922 9978
rect 2926 9974 2927 9978
rect 2931 9974 2932 9978
rect 2936 9974 2937 9978
rect 2941 9974 2942 9978
rect 2946 9974 2947 9978
rect 2951 9974 2952 9978
rect 2956 9974 2957 9978
rect 2961 9974 2962 9978
rect 2966 9974 2967 9978
rect 2971 9974 2972 9978
rect 2976 9974 2977 9978
rect 2981 9974 2982 9978
rect 2986 9974 2987 9978
rect 2991 9974 2992 9978
rect 2996 9974 2997 9978
rect 3001 9974 3002 9978
rect 3006 9974 3007 9978
rect 2917 9973 2921 9974
rect 2917 9968 2921 9969
rect 3007 9973 3011 9974
rect 3007 9968 3011 9969
rect 2917 9963 2921 9964
rect 2917 9958 2921 9959
rect 2917 9953 2921 9954
rect 2917 9948 2921 9949
rect 2917 9943 2921 9944
rect 2917 9938 2921 9939
rect 2917 9933 2921 9934
rect 2917 9928 2921 9929
rect 2917 9923 2921 9924
rect 2917 9918 2921 9919
rect 2917 9913 2921 9914
rect 2917 9908 2921 9909
rect 2917 9903 2921 9904
rect 2917 9898 2921 9899
rect 2917 9893 2921 9894
rect 2917 9888 2921 9889
rect 2917 9883 2921 9884
rect 2917 9878 2921 9879
rect 2917 9873 2921 9874
rect 2917 9868 2921 9869
rect 2917 9863 2921 9864
rect 2917 9858 2921 9859
rect 2917 9853 2921 9854
rect 2917 9848 2921 9849
rect 2934 9961 2937 9965
rect 2941 9961 2942 9965
rect 2946 9961 2947 9965
rect 2951 9961 2952 9965
rect 2956 9961 2957 9965
rect 2961 9961 2962 9965
rect 2966 9961 2967 9965
rect 2971 9961 2972 9965
rect 2976 9961 2977 9965
rect 2981 9961 2982 9965
rect 2986 9961 2987 9965
rect 2991 9961 2994 9965
rect 2930 9958 2934 9961
rect 2930 9953 2934 9954
rect 2994 9958 2998 9961
rect 2994 9953 2998 9954
rect 2930 9948 2934 9949
rect 2930 9943 2934 9944
rect 2930 9938 2934 9939
rect 2930 9933 2934 9934
rect 2930 9928 2934 9929
rect 2930 9923 2934 9924
rect 2930 9918 2934 9919
rect 2930 9913 2934 9914
rect 2930 9908 2934 9909
rect 2930 9903 2934 9904
rect 2930 9898 2934 9899
rect 2930 9893 2934 9894
rect 2930 9888 2934 9889
rect 2930 9883 2934 9884
rect 2930 9878 2934 9879
rect 2930 9873 2934 9874
rect 2930 9868 2934 9869
rect 2946 9949 2947 9953
rect 2951 9949 2952 9953
rect 2956 9949 2957 9953
rect 2961 9949 2962 9953
rect 2966 9949 2967 9953
rect 2971 9949 2972 9953
rect 2976 9949 2977 9953
rect 2981 9949 2982 9953
rect 2942 9948 2986 9949
rect 2946 9944 2947 9948
rect 2951 9944 2952 9948
rect 2956 9944 2957 9948
rect 2961 9944 2962 9948
rect 2966 9944 2967 9948
rect 2971 9944 2972 9948
rect 2976 9944 2977 9948
rect 2981 9944 2982 9948
rect 2942 9943 2986 9944
rect 2946 9939 2947 9943
rect 2951 9939 2952 9943
rect 2956 9939 2957 9943
rect 2961 9939 2962 9943
rect 2966 9939 2967 9943
rect 2971 9939 2972 9943
rect 2976 9939 2977 9943
rect 2981 9939 2982 9943
rect 2942 9938 2986 9939
rect 2946 9934 2947 9938
rect 2951 9934 2952 9938
rect 2956 9934 2957 9938
rect 2961 9934 2962 9938
rect 2966 9934 2967 9938
rect 2971 9934 2972 9938
rect 2976 9934 2977 9938
rect 2981 9934 2982 9938
rect 2942 9933 2986 9934
rect 2946 9929 2947 9933
rect 2951 9929 2952 9933
rect 2956 9929 2957 9933
rect 2961 9929 2962 9933
rect 2966 9929 2967 9933
rect 2971 9929 2972 9933
rect 2976 9929 2977 9933
rect 2981 9929 2982 9933
rect 2942 9928 2986 9929
rect 2946 9924 2947 9928
rect 2951 9924 2952 9928
rect 2956 9924 2957 9928
rect 2961 9924 2962 9928
rect 2966 9924 2967 9928
rect 2971 9924 2972 9928
rect 2976 9924 2977 9928
rect 2981 9924 2982 9928
rect 2942 9923 2986 9924
rect 2946 9919 2947 9923
rect 2951 9919 2952 9923
rect 2956 9919 2957 9923
rect 2961 9919 2962 9923
rect 2966 9919 2967 9923
rect 2971 9919 2972 9923
rect 2976 9919 2977 9923
rect 2981 9919 2982 9923
rect 2942 9918 2986 9919
rect 2946 9914 2947 9918
rect 2951 9914 2952 9918
rect 2956 9914 2957 9918
rect 2961 9914 2962 9918
rect 2966 9914 2967 9918
rect 2971 9914 2972 9918
rect 2976 9914 2977 9918
rect 2981 9914 2982 9918
rect 2942 9913 2986 9914
rect 2946 9909 2947 9913
rect 2951 9909 2952 9913
rect 2956 9909 2957 9913
rect 2961 9909 2962 9913
rect 2966 9909 2967 9913
rect 2971 9909 2972 9913
rect 2976 9909 2977 9913
rect 2981 9909 2982 9913
rect 2942 9908 2986 9909
rect 2946 9904 2947 9908
rect 2951 9904 2952 9908
rect 2956 9904 2957 9908
rect 2961 9904 2962 9908
rect 2966 9904 2967 9908
rect 2971 9904 2972 9908
rect 2976 9904 2977 9908
rect 2981 9904 2982 9908
rect 2942 9903 2986 9904
rect 2946 9899 2947 9903
rect 2951 9899 2952 9903
rect 2956 9899 2957 9903
rect 2961 9899 2962 9903
rect 2966 9899 2967 9903
rect 2971 9899 2972 9903
rect 2976 9899 2977 9903
rect 2981 9899 2982 9903
rect 2942 9898 2986 9899
rect 2946 9894 2947 9898
rect 2951 9894 2952 9898
rect 2956 9894 2957 9898
rect 2961 9894 2962 9898
rect 2966 9894 2967 9898
rect 2971 9894 2972 9898
rect 2976 9894 2977 9898
rect 2981 9894 2982 9898
rect 2942 9893 2986 9894
rect 2946 9889 2947 9893
rect 2951 9889 2952 9893
rect 2956 9889 2957 9893
rect 2961 9889 2962 9893
rect 2966 9889 2967 9893
rect 2971 9889 2972 9893
rect 2976 9889 2977 9893
rect 2981 9889 2982 9893
rect 2942 9888 2986 9889
rect 2946 9884 2947 9888
rect 2951 9884 2952 9888
rect 2956 9884 2957 9888
rect 2961 9884 2962 9888
rect 2966 9884 2967 9888
rect 2971 9884 2972 9888
rect 2976 9884 2977 9888
rect 2981 9884 2982 9888
rect 2942 9883 2986 9884
rect 2946 9879 2947 9883
rect 2951 9879 2952 9883
rect 2956 9879 2957 9883
rect 2961 9879 2962 9883
rect 2966 9879 2967 9883
rect 2971 9879 2972 9883
rect 2976 9879 2977 9883
rect 2981 9879 2982 9883
rect 2942 9878 2986 9879
rect 2946 9874 2947 9878
rect 2951 9874 2952 9878
rect 2956 9874 2957 9878
rect 2961 9874 2962 9878
rect 2966 9874 2967 9878
rect 2971 9874 2972 9878
rect 2976 9874 2977 9878
rect 2981 9874 2982 9878
rect 2942 9873 2986 9874
rect 2946 9869 2947 9873
rect 2951 9869 2952 9873
rect 2956 9869 2957 9873
rect 2961 9869 2962 9873
rect 2966 9869 2967 9873
rect 2971 9869 2972 9873
rect 2976 9869 2977 9873
rect 2981 9869 2982 9873
rect 2942 9868 2986 9869
rect 2946 9864 2947 9868
rect 2951 9864 2952 9868
rect 2956 9864 2957 9868
rect 2961 9864 2962 9868
rect 2966 9864 2967 9868
rect 2971 9864 2972 9868
rect 2976 9864 2977 9868
rect 2981 9864 2982 9868
rect 2994 9948 2998 9949
rect 2994 9943 2998 9944
rect 2994 9938 2998 9939
rect 2994 9933 2998 9934
rect 2994 9928 2998 9929
rect 2994 9923 2998 9924
rect 2994 9918 2998 9919
rect 2994 9913 2998 9914
rect 2994 9908 2998 9909
rect 2994 9903 2998 9904
rect 2994 9898 2998 9899
rect 2994 9893 2998 9894
rect 2994 9888 2998 9889
rect 2994 9883 2998 9884
rect 2994 9878 2998 9879
rect 2994 9873 2998 9874
rect 2994 9868 2998 9869
rect 2930 9863 2934 9864
rect 2930 9856 2934 9859
rect 2994 9863 2998 9864
rect 2994 9856 2998 9859
rect 2934 9848 2937 9856
rect 2941 9848 2942 9856
rect 2946 9848 2947 9856
rect 2951 9848 2952 9856
rect 2956 9848 2957 9856
rect 2961 9848 2962 9856
rect 2966 9848 2967 9856
rect 2971 9848 2972 9856
rect 2976 9848 2977 9856
rect 2981 9848 2982 9856
rect 2986 9848 2987 9856
rect 2991 9848 2994 9856
rect 3007 9963 3011 9964
rect 3007 9958 3011 9959
rect 3007 9953 3011 9954
rect 3033 9961 3054 9981
rect 3081 9974 3082 9978
rect 3086 9974 3087 9978
rect 3091 9974 3092 9978
rect 3096 9974 3097 9978
rect 3101 9974 3102 9978
rect 3106 9974 3107 9978
rect 3111 9974 3112 9978
rect 3116 9974 3117 9978
rect 3121 9974 3122 9978
rect 3126 9974 3127 9978
rect 3131 9974 3132 9978
rect 3136 9974 3137 9978
rect 3141 9974 3142 9978
rect 3146 9974 3147 9978
rect 3151 9974 3152 9978
rect 3156 9974 3157 9978
rect 3161 9974 3162 9978
rect 3166 9974 3167 9978
rect 3077 9973 3081 9974
rect 3077 9968 3081 9969
rect 3167 9973 3171 9974
rect 3167 9968 3171 9969
rect 3077 9963 3081 9964
rect 3077 9958 3081 9959
rect 3077 9953 3081 9954
rect 3007 9948 3011 9949
rect 3007 9943 3011 9944
rect 3007 9938 3011 9939
rect 3007 9933 3011 9934
rect 3007 9928 3011 9929
rect 3007 9923 3011 9924
rect 3007 9918 3011 9919
rect 3007 9913 3011 9914
rect 3007 9908 3011 9909
rect 3007 9903 3011 9904
rect 3007 9898 3011 9899
rect 3007 9893 3011 9894
rect 3007 9888 3011 9889
rect 3007 9883 3011 9884
rect 3077 9948 3081 9949
rect 3077 9943 3081 9944
rect 3077 9938 3081 9939
rect 3077 9933 3081 9934
rect 3077 9928 3081 9929
rect 3077 9923 3081 9924
rect 3077 9918 3081 9919
rect 3077 9913 3081 9914
rect 3077 9908 3081 9909
rect 3077 9903 3081 9904
rect 3077 9898 3081 9899
rect 3077 9893 3081 9894
rect 3077 9888 3081 9889
rect 3077 9883 3081 9884
rect 3007 9878 3011 9879
rect 3007 9873 3011 9874
rect 3007 9868 3011 9869
rect 3007 9863 3011 9864
rect 3007 9858 3011 9859
rect 3007 9853 3011 9854
rect 3007 9848 3011 9849
rect 2917 9843 2921 9844
rect 3033 9846 3054 9874
rect 3077 9878 3081 9879
rect 3077 9873 3081 9874
rect 3077 9868 3081 9869
rect 3077 9863 3081 9864
rect 3077 9858 3081 9859
rect 3077 9853 3081 9854
rect 3077 9848 3081 9849
rect 3094 9961 3097 9965
rect 3101 9961 3102 9965
rect 3106 9961 3107 9965
rect 3111 9961 3112 9965
rect 3116 9961 3117 9965
rect 3121 9961 3122 9965
rect 3126 9961 3127 9965
rect 3131 9961 3132 9965
rect 3136 9961 3137 9965
rect 3141 9961 3142 9965
rect 3146 9961 3147 9965
rect 3151 9961 3154 9965
rect 3090 9958 3094 9961
rect 3090 9953 3094 9954
rect 3154 9958 3158 9961
rect 3154 9953 3158 9954
rect 3090 9948 3094 9949
rect 3090 9943 3094 9944
rect 3090 9938 3094 9939
rect 3090 9933 3094 9934
rect 3090 9928 3094 9929
rect 3090 9923 3094 9924
rect 3090 9918 3094 9919
rect 3090 9913 3094 9914
rect 3090 9908 3094 9909
rect 3090 9903 3094 9904
rect 3090 9898 3094 9899
rect 3090 9893 3094 9894
rect 3090 9888 3094 9889
rect 3090 9883 3094 9884
rect 3090 9878 3094 9879
rect 3090 9873 3094 9874
rect 3090 9868 3094 9869
rect 3101 9949 3102 9953
rect 3106 9949 3107 9953
rect 3111 9949 3112 9953
rect 3116 9949 3117 9953
rect 3121 9949 3122 9953
rect 3126 9949 3127 9953
rect 3131 9949 3132 9953
rect 3136 9949 3137 9953
rect 3141 9949 3142 9953
rect 3101 9948 3146 9949
rect 3101 9944 3102 9948
rect 3106 9944 3107 9948
rect 3111 9944 3112 9948
rect 3116 9944 3117 9948
rect 3121 9944 3122 9948
rect 3126 9944 3127 9948
rect 3131 9944 3132 9948
rect 3136 9944 3137 9948
rect 3141 9944 3142 9948
rect 3101 9943 3146 9944
rect 3101 9939 3102 9943
rect 3106 9939 3107 9943
rect 3111 9939 3112 9943
rect 3116 9939 3117 9943
rect 3121 9939 3122 9943
rect 3126 9939 3127 9943
rect 3131 9939 3132 9943
rect 3136 9939 3137 9943
rect 3141 9939 3142 9943
rect 3101 9938 3146 9939
rect 3101 9934 3102 9938
rect 3106 9934 3107 9938
rect 3111 9934 3112 9938
rect 3116 9934 3117 9938
rect 3121 9934 3122 9938
rect 3126 9934 3127 9938
rect 3131 9934 3132 9938
rect 3136 9934 3137 9938
rect 3141 9934 3142 9938
rect 3101 9933 3146 9934
rect 3101 9929 3102 9933
rect 3106 9929 3107 9933
rect 3111 9929 3112 9933
rect 3116 9929 3117 9933
rect 3121 9929 3122 9933
rect 3126 9929 3127 9933
rect 3131 9929 3132 9933
rect 3136 9929 3137 9933
rect 3141 9929 3142 9933
rect 3101 9928 3146 9929
rect 3101 9924 3102 9928
rect 3106 9924 3107 9928
rect 3111 9924 3112 9928
rect 3116 9924 3117 9928
rect 3121 9924 3122 9928
rect 3126 9924 3127 9928
rect 3131 9924 3132 9928
rect 3136 9924 3137 9928
rect 3141 9924 3142 9928
rect 3101 9923 3146 9924
rect 3101 9919 3102 9923
rect 3106 9919 3107 9923
rect 3111 9919 3112 9923
rect 3116 9919 3117 9923
rect 3121 9919 3122 9923
rect 3126 9919 3127 9923
rect 3131 9919 3132 9923
rect 3136 9919 3137 9923
rect 3141 9919 3142 9923
rect 3101 9918 3146 9919
rect 3101 9914 3102 9918
rect 3106 9914 3107 9918
rect 3111 9914 3112 9918
rect 3116 9914 3117 9918
rect 3121 9914 3122 9918
rect 3126 9914 3127 9918
rect 3131 9914 3132 9918
rect 3136 9914 3137 9918
rect 3141 9914 3142 9918
rect 3101 9913 3146 9914
rect 3101 9909 3102 9913
rect 3106 9909 3107 9913
rect 3111 9909 3112 9913
rect 3116 9909 3117 9913
rect 3121 9909 3122 9913
rect 3126 9909 3127 9913
rect 3131 9909 3132 9913
rect 3136 9909 3137 9913
rect 3141 9909 3142 9913
rect 3101 9908 3146 9909
rect 3101 9904 3102 9908
rect 3106 9904 3107 9908
rect 3111 9904 3112 9908
rect 3116 9904 3117 9908
rect 3121 9904 3122 9908
rect 3126 9904 3127 9908
rect 3131 9904 3132 9908
rect 3136 9904 3137 9908
rect 3141 9904 3142 9908
rect 3101 9903 3146 9904
rect 3101 9899 3102 9903
rect 3106 9899 3107 9903
rect 3111 9899 3112 9903
rect 3116 9899 3117 9903
rect 3121 9899 3122 9903
rect 3126 9899 3127 9903
rect 3131 9899 3132 9903
rect 3136 9899 3137 9903
rect 3141 9899 3142 9903
rect 3101 9898 3146 9899
rect 3101 9894 3102 9898
rect 3106 9894 3107 9898
rect 3111 9894 3112 9898
rect 3116 9894 3117 9898
rect 3121 9894 3122 9898
rect 3126 9894 3127 9898
rect 3131 9894 3132 9898
rect 3136 9894 3137 9898
rect 3141 9894 3142 9898
rect 3101 9893 3146 9894
rect 3101 9889 3102 9893
rect 3106 9889 3107 9893
rect 3111 9889 3112 9893
rect 3116 9889 3117 9893
rect 3121 9889 3122 9893
rect 3126 9889 3127 9893
rect 3131 9889 3132 9893
rect 3136 9889 3137 9893
rect 3141 9889 3142 9893
rect 3101 9888 3146 9889
rect 3101 9884 3102 9888
rect 3106 9884 3107 9888
rect 3111 9884 3112 9888
rect 3116 9884 3117 9888
rect 3121 9884 3122 9888
rect 3126 9884 3127 9888
rect 3131 9884 3132 9888
rect 3136 9884 3137 9888
rect 3141 9884 3142 9888
rect 3101 9883 3146 9884
rect 3101 9879 3102 9883
rect 3106 9879 3107 9883
rect 3111 9879 3112 9883
rect 3116 9879 3117 9883
rect 3121 9879 3122 9883
rect 3126 9879 3127 9883
rect 3131 9879 3132 9883
rect 3136 9879 3137 9883
rect 3141 9879 3142 9883
rect 3101 9878 3146 9879
rect 3101 9874 3102 9878
rect 3106 9874 3107 9878
rect 3111 9874 3112 9878
rect 3116 9874 3117 9878
rect 3121 9874 3122 9878
rect 3126 9874 3127 9878
rect 3131 9874 3132 9878
rect 3136 9874 3137 9878
rect 3141 9874 3142 9878
rect 3101 9873 3146 9874
rect 3101 9869 3102 9873
rect 3106 9869 3107 9873
rect 3111 9869 3112 9873
rect 3116 9869 3117 9873
rect 3121 9869 3122 9873
rect 3126 9869 3127 9873
rect 3131 9869 3132 9873
rect 3136 9869 3137 9873
rect 3141 9869 3142 9873
rect 3101 9868 3146 9869
rect 3101 9864 3102 9868
rect 3106 9864 3107 9868
rect 3111 9864 3112 9868
rect 3116 9864 3117 9868
rect 3121 9864 3122 9868
rect 3126 9864 3127 9868
rect 3131 9864 3132 9868
rect 3136 9864 3137 9868
rect 3141 9864 3142 9868
rect 3154 9948 3158 9949
rect 3154 9943 3158 9944
rect 3154 9938 3158 9939
rect 3154 9933 3158 9934
rect 3154 9928 3158 9929
rect 3154 9923 3158 9924
rect 3154 9918 3158 9919
rect 3154 9913 3158 9914
rect 3154 9908 3158 9909
rect 3154 9903 3158 9904
rect 3154 9898 3158 9899
rect 3154 9893 3158 9894
rect 3154 9888 3158 9889
rect 3154 9883 3158 9884
rect 3154 9878 3158 9879
rect 3154 9873 3158 9874
rect 3154 9868 3158 9869
rect 3090 9863 3094 9864
rect 3090 9856 3094 9859
rect 3154 9863 3158 9864
rect 3154 9856 3158 9859
rect 3094 9848 3097 9856
rect 3101 9848 3102 9856
rect 3106 9848 3107 9856
rect 3111 9848 3112 9856
rect 3116 9848 3117 9856
rect 3121 9848 3122 9856
rect 3126 9848 3127 9856
rect 3131 9848 3132 9856
rect 3136 9848 3137 9856
rect 3141 9848 3142 9856
rect 3146 9848 3147 9856
rect 3151 9848 3154 9856
rect 3167 9963 3171 9964
rect 3167 9958 3171 9959
rect 3167 9953 3171 9954
rect 3167 9948 3171 9949
rect 3167 9943 3171 9944
rect 3167 9938 3171 9939
rect 3167 9933 3171 9934
rect 3167 9928 3171 9929
rect 3167 9923 3171 9924
rect 3167 9918 3171 9919
rect 3167 9913 3171 9914
rect 3167 9908 3171 9909
rect 3167 9903 3171 9904
rect 3167 9898 3171 9899
rect 3167 9893 3171 9894
rect 3167 9888 3171 9889
rect 3167 9883 3171 9884
rect 3167 9878 3171 9879
rect 3167 9873 3171 9874
rect 3167 9868 3171 9869
rect 3167 9863 3171 9864
rect 3167 9858 3171 9859
rect 3167 9853 3171 9854
rect 3167 9848 3171 9849
rect 3035 9844 3052 9846
rect 3007 9843 3011 9844
rect 2921 9839 2922 9843
rect 2926 9839 2927 9843
rect 2931 9839 2932 9843
rect 2936 9839 2937 9843
rect 2941 9839 2942 9843
rect 2946 9839 2947 9843
rect 2951 9839 2952 9843
rect 2956 9839 2957 9843
rect 2961 9839 2962 9843
rect 2966 9839 2967 9843
rect 2971 9839 2972 9843
rect 2976 9839 2977 9843
rect 2981 9839 2982 9843
rect 2986 9839 2987 9843
rect 2991 9839 2992 9843
rect 2996 9839 2997 9843
rect 3001 9839 3002 9843
rect 3006 9839 3007 9843
rect 3037 9842 3050 9844
rect 3077 9843 3081 9844
rect 3167 9843 3171 9844
rect 2805 9831 2861 9839
rect 2611 9827 2670 9831
rect 2796 9827 2861 9831
rect 2611 9815 2667 9827
rect 2726 9819 2756 9823
rect 2611 9811 2670 9815
rect 2740 9812 2744 9819
rect 2805 9815 2861 9827
rect 2611 9802 2667 9811
rect 2796 9811 2861 9815
rect 2726 9803 2737 9807
rect 2487 9795 2552 9799
rect 2290 9790 2358 9791
rect 2290 9786 2291 9790
rect 2295 9786 2296 9790
rect 2300 9786 2358 9790
rect 2417 9787 2447 9791
rect 2290 9785 2358 9786
rect 2290 9781 2291 9785
rect 2295 9781 2296 9785
rect 2300 9783 2358 9785
rect 2300 9781 2361 9783
rect 2290 9780 2361 9781
rect 2290 9776 2291 9780
rect 2295 9776 2296 9780
rect 2300 9779 2361 9780
rect 2300 9776 2358 9779
rect 2290 9775 2358 9776
rect 2290 9771 2291 9775
rect 2295 9771 2296 9775
rect 2300 9771 2358 9775
rect 2290 9770 2358 9771
rect 2290 9766 2291 9770
rect 2295 9766 2296 9770
rect 2300 9766 2358 9770
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2246 9761 2265 9762
rect 2250 9757 2251 9761
rect 2255 9757 2256 9761
rect 2260 9757 2261 9761
rect 2246 9756 2265 9757
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2246 9751 2265 9752
rect 2250 9747 2251 9751
rect 2255 9747 2256 9751
rect 2260 9747 2261 9751
rect 2246 9746 2265 9747
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2246 9741 2265 9742
rect 2250 9737 2251 9741
rect 2255 9737 2256 9741
rect 2260 9737 2261 9741
rect 2246 9736 2265 9737
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2290 9765 2358 9766
rect 2290 9761 2291 9765
rect 2295 9761 2296 9765
rect 2300 9761 2358 9765
rect 2290 9760 2358 9761
rect 2290 9756 2291 9760
rect 2295 9756 2296 9760
rect 2300 9756 2358 9760
rect 2290 9755 2358 9756
rect 2290 9751 2291 9755
rect 2295 9751 2296 9755
rect 2300 9751 2358 9755
rect 2290 9750 2358 9751
rect 2290 9746 2291 9750
rect 2295 9746 2296 9750
rect 2300 9746 2358 9750
rect 2290 9745 2358 9746
rect 2290 9741 2291 9745
rect 2295 9741 2296 9745
rect 2300 9741 2358 9745
rect 2290 9740 2358 9741
rect 2290 9736 2291 9740
rect 2295 9736 2296 9740
rect 2300 9736 2358 9740
rect 2290 9734 2358 9736
rect 2191 9718 2192 9722
rect 2196 9718 2197 9722
rect 2201 9718 2202 9722
rect 2206 9718 2207 9722
rect 2211 9718 2212 9722
rect 2216 9718 2217 9722
rect 2221 9718 2222 9722
rect 2226 9718 2227 9722
rect 2231 9718 2232 9722
rect 2236 9718 2237 9722
rect 2241 9718 2243 9722
rect 2187 9717 2243 9718
rect 2191 9713 2192 9717
rect 2196 9713 2197 9717
rect 2201 9713 2202 9717
rect 2206 9713 2207 9717
rect 2211 9713 2212 9717
rect 2216 9713 2217 9717
rect 2221 9713 2222 9717
rect 2226 9713 2227 9717
rect 2231 9713 2232 9717
rect 2236 9713 2237 9717
rect 2241 9713 2243 9717
rect 2187 9712 2243 9713
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2246 9715 2265 9716
rect 2250 9711 2251 9715
rect 2255 9711 2256 9715
rect 2260 9711 2261 9715
rect 2246 9710 2265 9711
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2246 9705 2265 9706
rect 2250 9701 2251 9705
rect 2255 9701 2256 9705
rect 2260 9701 2261 9705
rect 2246 9700 2265 9701
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2246 9695 2265 9696
rect 2250 9691 2251 9695
rect 2255 9691 2256 9695
rect 2260 9691 2261 9695
rect 2246 9690 2265 9691
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2422 9597 2435 9787
rect 2496 9783 2552 9795
rect 2487 9779 2552 9783
rect 2496 9722 2552 9779
rect 2599 9800 2667 9802
rect 2599 9796 2600 9800
rect 2604 9796 2605 9800
rect 2609 9799 2667 9800
rect 2730 9800 2737 9803
rect 2749 9803 2756 9807
rect 2749 9800 2753 9803
rect 2609 9796 2670 9799
rect 2599 9795 2670 9796
rect 2599 9791 2600 9795
rect 2604 9791 2605 9795
rect 2609 9791 2667 9795
rect 2730 9791 2753 9800
rect 2805 9799 2861 9811
rect 2920 9831 2976 9839
rect 3039 9831 3048 9842
rect 3081 9839 3082 9843
rect 3086 9839 3087 9843
rect 3091 9839 3092 9843
rect 3096 9839 3097 9843
rect 3101 9839 3102 9843
rect 3106 9839 3107 9843
rect 3111 9839 3112 9843
rect 3116 9839 3117 9843
rect 3121 9839 3122 9843
rect 3126 9839 3127 9843
rect 3131 9839 3132 9843
rect 3136 9839 3137 9843
rect 3141 9839 3142 9843
rect 3146 9839 3147 9843
rect 3151 9839 3152 9843
rect 3156 9839 3157 9843
rect 3161 9839 3162 9843
rect 3166 9839 3167 9843
rect 3230 9974 3231 9978
rect 3235 9974 3236 9978
rect 3240 9974 3241 9978
rect 3245 9974 3246 9978
rect 3250 9974 3251 9978
rect 3255 9974 3256 9978
rect 3260 9974 3261 9978
rect 3265 9974 3266 9978
rect 3270 9974 3271 9978
rect 3275 9974 3276 9978
rect 3280 9974 3281 9978
rect 3285 9974 3286 9978
rect 3290 9974 3291 9978
rect 3295 9974 3296 9978
rect 3300 9974 3301 9978
rect 3305 9974 3306 9978
rect 3310 9974 3311 9978
rect 3315 9974 3316 9978
rect 3226 9973 3230 9974
rect 3226 9968 3230 9969
rect 3316 9973 3320 9974
rect 3316 9968 3320 9969
rect 3226 9963 3230 9964
rect 3226 9958 3230 9959
rect 3226 9953 3230 9954
rect 3226 9948 3230 9949
rect 3226 9943 3230 9944
rect 3226 9938 3230 9939
rect 3226 9933 3230 9934
rect 3226 9928 3230 9929
rect 3226 9923 3230 9924
rect 3226 9918 3230 9919
rect 3226 9913 3230 9914
rect 3226 9908 3230 9909
rect 3226 9903 3230 9904
rect 3226 9898 3230 9899
rect 3226 9893 3230 9894
rect 3226 9888 3230 9889
rect 3226 9883 3230 9884
rect 3226 9878 3230 9879
rect 3226 9873 3230 9874
rect 3226 9868 3230 9869
rect 3226 9863 3230 9864
rect 3226 9858 3230 9859
rect 3226 9853 3230 9854
rect 3226 9848 3230 9849
rect 3243 9961 3246 9965
rect 3250 9961 3251 9965
rect 3255 9961 3256 9965
rect 3260 9961 3261 9965
rect 3265 9961 3266 9965
rect 3270 9961 3271 9965
rect 3275 9961 3276 9965
rect 3280 9961 3281 9965
rect 3285 9961 3286 9965
rect 3290 9961 3291 9965
rect 3295 9961 3296 9965
rect 3300 9961 3303 9965
rect 3239 9958 3243 9961
rect 3239 9953 3243 9954
rect 3303 9958 3307 9961
rect 3303 9953 3307 9954
rect 3239 9948 3243 9949
rect 3239 9943 3243 9944
rect 3239 9938 3243 9939
rect 3239 9933 3243 9934
rect 3239 9928 3243 9929
rect 3239 9923 3243 9924
rect 3239 9918 3243 9919
rect 3239 9913 3243 9914
rect 3239 9908 3243 9909
rect 3239 9903 3243 9904
rect 3239 9898 3243 9899
rect 3239 9893 3243 9894
rect 3239 9888 3243 9889
rect 3239 9883 3243 9884
rect 3239 9878 3243 9879
rect 3239 9873 3243 9874
rect 3239 9868 3243 9869
rect 3255 9949 3256 9953
rect 3260 9949 3261 9953
rect 3265 9949 3266 9953
rect 3270 9949 3271 9953
rect 3275 9949 3276 9953
rect 3280 9949 3281 9953
rect 3285 9949 3286 9953
rect 3290 9949 3291 9953
rect 3251 9948 3295 9949
rect 3255 9944 3256 9948
rect 3260 9944 3261 9948
rect 3265 9944 3266 9948
rect 3270 9944 3271 9948
rect 3275 9944 3276 9948
rect 3280 9944 3281 9948
rect 3285 9944 3286 9948
rect 3290 9944 3291 9948
rect 3251 9943 3295 9944
rect 3255 9939 3256 9943
rect 3260 9939 3261 9943
rect 3265 9939 3266 9943
rect 3270 9939 3271 9943
rect 3275 9939 3276 9943
rect 3280 9939 3281 9943
rect 3285 9939 3286 9943
rect 3290 9939 3291 9943
rect 3251 9938 3295 9939
rect 3255 9934 3256 9938
rect 3260 9934 3261 9938
rect 3265 9934 3266 9938
rect 3270 9934 3271 9938
rect 3275 9934 3276 9938
rect 3280 9934 3281 9938
rect 3285 9934 3286 9938
rect 3290 9934 3291 9938
rect 3251 9933 3295 9934
rect 3255 9929 3256 9933
rect 3260 9929 3261 9933
rect 3265 9929 3266 9933
rect 3270 9929 3271 9933
rect 3275 9929 3276 9933
rect 3280 9929 3281 9933
rect 3285 9929 3286 9933
rect 3290 9929 3291 9933
rect 3251 9928 3295 9929
rect 3255 9924 3256 9928
rect 3260 9924 3261 9928
rect 3265 9924 3266 9928
rect 3270 9924 3271 9928
rect 3275 9924 3276 9928
rect 3280 9924 3281 9928
rect 3285 9924 3286 9928
rect 3290 9924 3291 9928
rect 3251 9923 3295 9924
rect 3255 9919 3256 9923
rect 3260 9919 3261 9923
rect 3265 9919 3266 9923
rect 3270 9919 3271 9923
rect 3275 9919 3276 9923
rect 3280 9919 3281 9923
rect 3285 9919 3286 9923
rect 3290 9919 3291 9923
rect 3251 9918 3295 9919
rect 3255 9914 3256 9918
rect 3260 9914 3261 9918
rect 3265 9914 3266 9918
rect 3270 9914 3271 9918
rect 3275 9914 3276 9918
rect 3280 9914 3281 9918
rect 3285 9914 3286 9918
rect 3290 9914 3291 9918
rect 3251 9913 3295 9914
rect 3255 9909 3256 9913
rect 3260 9909 3261 9913
rect 3265 9909 3266 9913
rect 3270 9909 3271 9913
rect 3275 9909 3276 9913
rect 3280 9909 3281 9913
rect 3285 9909 3286 9913
rect 3290 9909 3291 9913
rect 3251 9908 3295 9909
rect 3255 9904 3256 9908
rect 3260 9904 3261 9908
rect 3265 9904 3266 9908
rect 3270 9904 3271 9908
rect 3275 9904 3276 9908
rect 3280 9904 3281 9908
rect 3285 9904 3286 9908
rect 3290 9904 3291 9908
rect 3251 9903 3295 9904
rect 3255 9899 3256 9903
rect 3260 9899 3261 9903
rect 3265 9899 3266 9903
rect 3270 9899 3271 9903
rect 3275 9899 3276 9903
rect 3280 9899 3281 9903
rect 3285 9899 3286 9903
rect 3290 9899 3291 9903
rect 3251 9898 3295 9899
rect 3255 9894 3256 9898
rect 3260 9894 3261 9898
rect 3265 9894 3266 9898
rect 3270 9894 3271 9898
rect 3275 9894 3276 9898
rect 3280 9894 3281 9898
rect 3285 9894 3286 9898
rect 3290 9894 3291 9898
rect 3251 9893 3295 9894
rect 3255 9889 3256 9893
rect 3260 9889 3261 9893
rect 3265 9889 3266 9893
rect 3270 9889 3271 9893
rect 3275 9889 3276 9893
rect 3280 9889 3281 9893
rect 3285 9889 3286 9893
rect 3290 9889 3291 9893
rect 3251 9888 3295 9889
rect 3255 9884 3256 9888
rect 3260 9884 3261 9888
rect 3265 9884 3266 9888
rect 3270 9884 3271 9888
rect 3275 9884 3276 9888
rect 3280 9884 3281 9888
rect 3285 9884 3286 9888
rect 3290 9884 3291 9888
rect 3251 9883 3295 9884
rect 3255 9879 3256 9883
rect 3260 9879 3261 9883
rect 3265 9879 3266 9883
rect 3270 9879 3271 9883
rect 3275 9879 3276 9883
rect 3280 9879 3281 9883
rect 3285 9879 3286 9883
rect 3290 9879 3291 9883
rect 3251 9878 3295 9879
rect 3255 9874 3256 9878
rect 3260 9874 3261 9878
rect 3265 9874 3266 9878
rect 3270 9874 3271 9878
rect 3275 9874 3276 9878
rect 3280 9874 3281 9878
rect 3285 9874 3286 9878
rect 3290 9874 3291 9878
rect 3251 9873 3295 9874
rect 3255 9869 3256 9873
rect 3260 9869 3261 9873
rect 3265 9869 3266 9873
rect 3270 9869 3271 9873
rect 3275 9869 3276 9873
rect 3280 9869 3281 9873
rect 3285 9869 3286 9873
rect 3290 9869 3291 9873
rect 3251 9868 3295 9869
rect 3255 9864 3256 9868
rect 3260 9864 3261 9868
rect 3265 9864 3266 9868
rect 3270 9864 3271 9868
rect 3275 9864 3276 9868
rect 3280 9864 3281 9868
rect 3285 9864 3286 9868
rect 3290 9864 3291 9868
rect 3303 9948 3307 9949
rect 3303 9943 3307 9944
rect 3303 9938 3307 9939
rect 3303 9933 3307 9934
rect 3303 9928 3307 9929
rect 3303 9923 3307 9924
rect 3303 9918 3307 9919
rect 3303 9913 3307 9914
rect 3303 9908 3307 9909
rect 3303 9903 3307 9904
rect 3303 9898 3307 9899
rect 3303 9893 3307 9894
rect 3303 9888 3307 9889
rect 3303 9883 3307 9884
rect 3303 9878 3307 9879
rect 3303 9873 3307 9874
rect 3303 9868 3307 9869
rect 3239 9863 3243 9864
rect 3239 9856 3243 9859
rect 3303 9863 3307 9864
rect 3303 9856 3307 9859
rect 3243 9848 3246 9856
rect 3250 9848 3251 9856
rect 3255 9848 3256 9856
rect 3260 9848 3261 9856
rect 3265 9848 3266 9856
rect 3270 9848 3271 9856
rect 3275 9848 3276 9856
rect 3280 9848 3281 9856
rect 3285 9848 3286 9856
rect 3290 9848 3291 9856
rect 3295 9848 3296 9856
rect 3300 9848 3303 9856
rect 3316 9963 3320 9964
rect 3316 9958 3320 9959
rect 3316 9953 3320 9954
rect 3316 9948 3320 9949
rect 3316 9943 3320 9944
rect 3316 9938 3320 9939
rect 3316 9933 3320 9934
rect 3316 9928 3320 9929
rect 3316 9923 3320 9924
rect 3316 9918 3320 9919
rect 3316 9913 3320 9914
rect 3316 9908 3320 9909
rect 3316 9903 3320 9904
rect 3316 9898 3320 9899
rect 3316 9893 3320 9894
rect 3316 9888 3320 9889
rect 3316 9883 3320 9884
rect 3316 9878 3320 9879
rect 3316 9873 3320 9874
rect 3316 9868 3320 9869
rect 3316 9863 3320 9864
rect 3316 9858 3320 9859
rect 3316 9853 3320 9854
rect 3316 9848 3320 9849
rect 3226 9843 3230 9844
rect 3316 9843 3320 9844
rect 3230 9839 3231 9843
rect 3235 9839 3236 9843
rect 3240 9839 3241 9843
rect 3245 9839 3246 9843
rect 3250 9839 3251 9843
rect 3255 9839 3256 9843
rect 3260 9839 3261 9843
rect 3265 9839 3266 9843
rect 3270 9839 3271 9843
rect 3275 9839 3276 9843
rect 3280 9839 3281 9843
rect 3285 9839 3286 9843
rect 3290 9839 3291 9843
rect 3295 9839 3296 9843
rect 3300 9839 3301 9843
rect 3305 9839 3306 9843
rect 3310 9839 3311 9843
rect 3315 9839 3316 9843
rect 3114 9831 3170 9839
rect 2920 9827 2979 9831
rect 3105 9827 3170 9831
rect 2920 9815 2976 9827
rect 3035 9819 3065 9823
rect 2920 9811 2979 9815
rect 3049 9812 3053 9819
rect 3114 9815 3170 9827
rect 2920 9802 2976 9811
rect 3105 9811 3170 9815
rect 3035 9803 3046 9807
rect 2796 9795 2861 9799
rect 2599 9790 2667 9791
rect 2599 9786 2600 9790
rect 2604 9786 2605 9790
rect 2609 9786 2667 9790
rect 2726 9787 2756 9791
rect 2599 9785 2667 9786
rect 2599 9781 2600 9785
rect 2604 9781 2605 9785
rect 2609 9783 2667 9785
rect 2609 9781 2670 9783
rect 2599 9780 2670 9781
rect 2599 9776 2600 9780
rect 2604 9776 2605 9780
rect 2609 9779 2670 9780
rect 2609 9776 2667 9779
rect 2599 9775 2667 9776
rect 2599 9771 2600 9775
rect 2604 9771 2605 9775
rect 2609 9771 2667 9775
rect 2599 9770 2667 9771
rect 2599 9766 2600 9770
rect 2604 9766 2605 9770
rect 2609 9766 2667 9770
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2555 9761 2574 9762
rect 2559 9757 2560 9761
rect 2564 9757 2565 9761
rect 2569 9757 2570 9761
rect 2555 9756 2574 9757
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2555 9751 2574 9752
rect 2559 9747 2560 9751
rect 2564 9747 2565 9751
rect 2569 9747 2570 9751
rect 2555 9746 2574 9747
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2555 9741 2574 9742
rect 2559 9737 2560 9741
rect 2564 9737 2565 9741
rect 2569 9737 2570 9741
rect 2555 9736 2574 9737
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2599 9765 2667 9766
rect 2599 9761 2600 9765
rect 2604 9761 2605 9765
rect 2609 9761 2667 9765
rect 2599 9760 2667 9761
rect 2599 9756 2600 9760
rect 2604 9756 2605 9760
rect 2609 9756 2667 9760
rect 2599 9755 2667 9756
rect 2599 9751 2600 9755
rect 2604 9751 2605 9755
rect 2609 9751 2667 9755
rect 2599 9750 2667 9751
rect 2599 9746 2600 9750
rect 2604 9746 2605 9750
rect 2609 9746 2667 9750
rect 2599 9745 2667 9746
rect 2599 9741 2600 9745
rect 2604 9741 2605 9745
rect 2609 9741 2667 9745
rect 2599 9740 2667 9741
rect 2599 9736 2600 9740
rect 2604 9736 2605 9740
rect 2609 9736 2667 9740
rect 2599 9734 2667 9736
rect 2500 9718 2501 9722
rect 2505 9718 2506 9722
rect 2510 9718 2511 9722
rect 2515 9718 2516 9722
rect 2520 9718 2521 9722
rect 2525 9718 2526 9722
rect 2530 9718 2531 9722
rect 2535 9718 2536 9722
rect 2540 9718 2541 9722
rect 2545 9718 2546 9722
rect 2550 9718 2552 9722
rect 2496 9717 2552 9718
rect 2500 9713 2501 9717
rect 2505 9713 2506 9717
rect 2510 9713 2511 9717
rect 2515 9713 2516 9717
rect 2520 9713 2521 9717
rect 2525 9713 2526 9717
rect 2530 9713 2531 9717
rect 2535 9713 2536 9717
rect 2540 9713 2541 9717
rect 2545 9713 2546 9717
rect 2550 9713 2552 9717
rect 2496 9712 2552 9713
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2555 9715 2574 9716
rect 2559 9711 2560 9715
rect 2564 9711 2565 9715
rect 2569 9711 2570 9715
rect 2555 9710 2574 9711
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2555 9705 2574 9706
rect 2559 9701 2560 9705
rect 2564 9701 2565 9705
rect 2569 9701 2570 9705
rect 2555 9700 2574 9701
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2555 9695 2574 9696
rect 2559 9691 2560 9695
rect 2564 9691 2565 9695
rect 2569 9691 2570 9695
rect 2555 9690 2574 9691
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2731 9609 2744 9787
rect 2805 9783 2861 9795
rect 2796 9779 2861 9783
rect 2805 9722 2861 9779
rect 2908 9800 2976 9802
rect 2908 9796 2909 9800
rect 2913 9796 2914 9800
rect 2918 9799 2976 9800
rect 3039 9800 3046 9803
rect 3058 9803 3065 9807
rect 3058 9800 3062 9803
rect 2918 9796 2979 9799
rect 2908 9795 2979 9796
rect 2908 9791 2909 9795
rect 2913 9791 2914 9795
rect 2918 9791 2976 9795
rect 3039 9791 3062 9800
rect 3114 9799 3170 9811
rect 3229 9802 3285 9839
rect 3105 9795 3170 9799
rect 2908 9790 2976 9791
rect 2908 9786 2909 9790
rect 2913 9786 2914 9790
rect 2918 9786 2976 9790
rect 3035 9787 3065 9791
rect 2908 9785 2976 9786
rect 2908 9781 2909 9785
rect 2913 9781 2914 9785
rect 2918 9783 2976 9785
rect 2918 9781 2979 9783
rect 2908 9780 2979 9781
rect 2908 9776 2909 9780
rect 2913 9776 2914 9780
rect 2918 9779 2979 9780
rect 2918 9776 2976 9779
rect 2908 9775 2976 9776
rect 2908 9771 2909 9775
rect 2913 9771 2914 9775
rect 2918 9771 2976 9775
rect 2908 9770 2976 9771
rect 2908 9766 2909 9770
rect 2913 9766 2914 9770
rect 2918 9766 2976 9770
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2864 9761 2883 9762
rect 2868 9757 2869 9761
rect 2873 9757 2874 9761
rect 2878 9757 2879 9761
rect 2864 9756 2883 9757
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2864 9751 2883 9752
rect 2868 9747 2869 9751
rect 2873 9747 2874 9751
rect 2878 9747 2879 9751
rect 2864 9746 2883 9747
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2864 9741 2883 9742
rect 2868 9737 2869 9741
rect 2873 9737 2874 9741
rect 2878 9737 2879 9741
rect 2864 9736 2883 9737
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2908 9765 2976 9766
rect 2908 9761 2909 9765
rect 2913 9761 2914 9765
rect 2918 9761 2976 9765
rect 2908 9760 2976 9761
rect 2908 9756 2909 9760
rect 2913 9756 2914 9760
rect 2918 9756 2976 9760
rect 2908 9755 2976 9756
rect 2908 9751 2909 9755
rect 2913 9751 2914 9755
rect 2918 9751 2976 9755
rect 2908 9750 2976 9751
rect 2908 9746 2909 9750
rect 2913 9746 2914 9750
rect 2918 9746 2976 9750
rect 2908 9745 2976 9746
rect 2908 9741 2909 9745
rect 2913 9741 2914 9745
rect 2918 9741 2976 9745
rect 2908 9740 2976 9741
rect 2908 9736 2909 9740
rect 2913 9736 2914 9740
rect 2918 9736 2976 9740
rect 2908 9734 2976 9736
rect 2809 9718 2810 9722
rect 2814 9718 2815 9722
rect 2819 9718 2820 9722
rect 2824 9718 2825 9722
rect 2829 9718 2830 9722
rect 2834 9718 2835 9722
rect 2839 9718 2840 9722
rect 2844 9718 2845 9722
rect 2849 9718 2850 9722
rect 2854 9718 2855 9722
rect 2859 9718 2861 9722
rect 2805 9717 2861 9718
rect 2809 9713 2810 9717
rect 2814 9713 2815 9717
rect 2819 9713 2820 9717
rect 2824 9713 2825 9717
rect 2829 9713 2830 9717
rect 2834 9713 2835 9717
rect 2839 9713 2840 9717
rect 2844 9713 2845 9717
rect 2849 9713 2850 9717
rect 2854 9713 2855 9717
rect 2859 9713 2861 9717
rect 2805 9712 2861 9713
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2864 9715 2883 9716
rect 2868 9711 2869 9715
rect 2873 9711 2874 9715
rect 2878 9711 2879 9715
rect 2864 9710 2883 9711
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2864 9705 2883 9706
rect 2868 9701 2869 9705
rect 2873 9701 2874 9705
rect 2878 9701 2879 9705
rect 2864 9700 2883 9701
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2864 9695 2883 9696
rect 2868 9691 2869 9695
rect 2873 9691 2874 9695
rect 2878 9691 2879 9695
rect 2864 9690 2883 9691
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 3040 9611 3053 9787
rect 3114 9783 3170 9795
rect 3105 9779 3170 9783
rect 3114 9722 3170 9779
rect 3217 9800 3285 9802
rect 3217 9796 3218 9800
rect 3222 9796 3223 9800
rect 3227 9796 3285 9800
rect 3217 9795 3285 9796
rect 3217 9791 3218 9795
rect 3222 9791 3223 9795
rect 3227 9791 3285 9795
rect 3217 9790 3285 9791
rect 3217 9786 3218 9790
rect 3222 9786 3223 9790
rect 3227 9786 3285 9790
rect 3217 9785 3285 9786
rect 3217 9781 3218 9785
rect 3222 9781 3223 9785
rect 3227 9781 3285 9785
rect 3217 9780 3285 9781
rect 3217 9776 3218 9780
rect 3222 9776 3223 9780
rect 3227 9776 3285 9780
rect 3217 9775 3285 9776
rect 3217 9771 3218 9775
rect 3222 9771 3223 9775
rect 3227 9771 3285 9775
rect 3217 9770 3285 9771
rect 3217 9766 3218 9770
rect 3222 9766 3223 9770
rect 3227 9766 3285 9770
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3173 9761 3192 9762
rect 3177 9757 3178 9761
rect 3182 9757 3183 9761
rect 3187 9757 3188 9761
rect 3173 9756 3192 9757
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3173 9751 3192 9752
rect 3177 9747 3178 9751
rect 3182 9747 3183 9751
rect 3187 9747 3188 9751
rect 3173 9746 3192 9747
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3173 9741 3192 9742
rect 3177 9737 3178 9741
rect 3182 9737 3183 9741
rect 3187 9737 3188 9741
rect 3173 9736 3192 9737
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3217 9765 3285 9766
rect 3217 9761 3218 9765
rect 3222 9761 3223 9765
rect 3227 9761 3285 9765
rect 3217 9760 3285 9761
rect 3217 9756 3218 9760
rect 3222 9756 3223 9760
rect 3227 9756 3285 9760
rect 3217 9755 3285 9756
rect 3217 9751 3218 9755
rect 3222 9751 3223 9755
rect 3227 9751 3285 9755
rect 3217 9750 3285 9751
rect 3217 9746 3218 9750
rect 3222 9746 3223 9750
rect 3227 9746 3285 9750
rect 3217 9745 3285 9746
rect 3217 9741 3218 9745
rect 3222 9741 3223 9745
rect 3227 9741 3285 9745
rect 3217 9740 3285 9741
rect 3217 9736 3218 9740
rect 3222 9736 3223 9740
rect 3227 9736 3285 9740
rect 3217 9734 3285 9736
rect 3118 9718 3119 9722
rect 3123 9718 3124 9722
rect 3128 9718 3129 9722
rect 3133 9718 3134 9722
rect 3138 9718 3139 9722
rect 3143 9718 3144 9722
rect 3148 9718 3149 9722
rect 3153 9718 3154 9722
rect 3158 9718 3159 9722
rect 3163 9718 3164 9722
rect 3168 9718 3170 9722
rect 3114 9717 3170 9718
rect 3118 9713 3119 9717
rect 3123 9713 3124 9717
rect 3128 9713 3129 9717
rect 3133 9713 3134 9717
rect 3138 9713 3139 9717
rect 3143 9713 3144 9717
rect 3148 9713 3149 9717
rect 3153 9713 3154 9717
rect 3158 9713 3159 9717
rect 3163 9713 3164 9717
rect 3168 9713 3170 9717
rect 3114 9712 3170 9713
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3173 9715 3192 9716
rect 3177 9711 3178 9715
rect 3182 9711 3183 9715
rect 3187 9711 3188 9715
rect 3173 9710 3192 9711
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3173 9705 3192 9706
rect 3177 9701 3178 9705
rect 3182 9701 3183 9705
rect 3187 9701 3188 9705
rect 3173 9700 3192 9701
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3173 9695 3192 9696
rect 3177 9691 3178 9695
rect 3182 9691 3183 9695
rect 3187 9691 3188 9695
rect 3173 9690 3192 9691
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3327 9715 3379 9981
rect 3390 9974 3391 9978
rect 3395 9974 3396 9978
rect 3400 9974 3401 9978
rect 3405 9974 3406 9978
rect 3410 9974 3411 9978
rect 3415 9974 3416 9978
rect 3420 9974 3421 9978
rect 3425 9974 3426 9978
rect 3430 9974 3431 9978
rect 3435 9974 3436 9978
rect 3440 9974 3441 9978
rect 3445 9974 3446 9978
rect 3450 9974 3451 9978
rect 3455 9974 3456 9978
rect 3460 9974 3461 9978
rect 3465 9974 3466 9978
rect 3470 9974 3471 9978
rect 3475 9974 3476 9978
rect 3386 9973 3390 9974
rect 3386 9968 3390 9969
rect 3476 9973 3480 9974
rect 3476 9968 3480 9969
rect 3386 9963 3390 9964
rect 3386 9958 3390 9959
rect 3386 9953 3390 9954
rect 3386 9948 3390 9949
rect 3386 9943 3390 9944
rect 3386 9938 3390 9939
rect 3386 9933 3390 9934
rect 3386 9928 3390 9929
rect 3386 9923 3390 9924
rect 3386 9918 3390 9919
rect 3386 9913 3390 9914
rect 3386 9908 3390 9909
rect 3386 9903 3390 9904
rect 3386 9898 3390 9899
rect 3386 9893 3390 9894
rect 3386 9888 3390 9889
rect 3386 9883 3390 9884
rect 3386 9878 3390 9879
rect 3386 9873 3390 9874
rect 3386 9868 3390 9869
rect 3386 9863 3390 9864
rect 3386 9858 3390 9859
rect 3386 9853 3390 9854
rect 3386 9848 3390 9849
rect 3403 9961 3406 9965
rect 3410 9961 3411 9965
rect 3415 9961 3416 9965
rect 3420 9961 3421 9965
rect 3425 9961 3426 9965
rect 3430 9961 3431 9965
rect 3435 9961 3436 9965
rect 3440 9961 3441 9965
rect 3445 9961 3446 9965
rect 3450 9961 3451 9965
rect 3455 9961 3456 9965
rect 3460 9961 3463 9965
rect 3399 9958 3403 9961
rect 3399 9953 3403 9954
rect 3463 9958 3467 9961
rect 3463 9953 3467 9954
rect 3399 9948 3403 9949
rect 3399 9943 3403 9944
rect 3399 9938 3403 9939
rect 3399 9933 3403 9934
rect 3399 9928 3403 9929
rect 3399 9923 3403 9924
rect 3399 9918 3403 9919
rect 3399 9913 3403 9914
rect 3399 9908 3403 9909
rect 3399 9903 3403 9904
rect 3399 9898 3403 9899
rect 3399 9893 3403 9894
rect 3399 9888 3403 9889
rect 3399 9883 3403 9884
rect 3399 9878 3403 9879
rect 3399 9873 3403 9874
rect 3399 9868 3403 9869
rect 3410 9949 3411 9953
rect 3415 9949 3416 9953
rect 3420 9949 3421 9953
rect 3425 9949 3426 9953
rect 3430 9949 3431 9953
rect 3435 9949 3436 9953
rect 3440 9949 3441 9953
rect 3445 9949 3446 9953
rect 3450 9949 3451 9953
rect 3410 9948 3455 9949
rect 3410 9944 3411 9948
rect 3415 9944 3416 9948
rect 3420 9944 3421 9948
rect 3425 9944 3426 9948
rect 3430 9944 3431 9948
rect 3435 9944 3436 9948
rect 3440 9944 3441 9948
rect 3445 9944 3446 9948
rect 3450 9944 3451 9948
rect 3410 9943 3455 9944
rect 3410 9939 3411 9943
rect 3415 9939 3416 9943
rect 3420 9939 3421 9943
rect 3425 9939 3426 9943
rect 3430 9939 3431 9943
rect 3435 9939 3436 9943
rect 3440 9939 3441 9943
rect 3445 9939 3446 9943
rect 3450 9939 3451 9943
rect 3410 9938 3455 9939
rect 3410 9934 3411 9938
rect 3415 9934 3416 9938
rect 3420 9934 3421 9938
rect 3425 9934 3426 9938
rect 3430 9934 3431 9938
rect 3435 9934 3436 9938
rect 3440 9934 3441 9938
rect 3445 9934 3446 9938
rect 3450 9934 3451 9938
rect 3410 9933 3455 9934
rect 3410 9929 3411 9933
rect 3415 9929 3416 9933
rect 3420 9929 3421 9933
rect 3425 9929 3426 9933
rect 3430 9929 3431 9933
rect 3435 9929 3436 9933
rect 3440 9929 3441 9933
rect 3445 9929 3446 9933
rect 3450 9929 3451 9933
rect 3410 9928 3455 9929
rect 3410 9924 3411 9928
rect 3415 9924 3416 9928
rect 3420 9924 3421 9928
rect 3425 9924 3426 9928
rect 3430 9924 3431 9928
rect 3435 9924 3436 9928
rect 3440 9924 3441 9928
rect 3445 9924 3446 9928
rect 3450 9924 3451 9928
rect 3410 9923 3455 9924
rect 3410 9919 3411 9923
rect 3415 9919 3416 9923
rect 3420 9919 3421 9923
rect 3425 9919 3426 9923
rect 3430 9919 3431 9923
rect 3435 9919 3436 9923
rect 3440 9919 3441 9923
rect 3445 9919 3446 9923
rect 3450 9919 3451 9923
rect 3410 9918 3455 9919
rect 3410 9914 3411 9918
rect 3415 9914 3416 9918
rect 3420 9914 3421 9918
rect 3425 9914 3426 9918
rect 3430 9914 3431 9918
rect 3435 9914 3436 9918
rect 3440 9914 3441 9918
rect 3445 9914 3446 9918
rect 3450 9914 3451 9918
rect 3410 9913 3455 9914
rect 3410 9909 3411 9913
rect 3415 9909 3416 9913
rect 3420 9909 3421 9913
rect 3425 9909 3426 9913
rect 3430 9909 3431 9913
rect 3435 9909 3436 9913
rect 3440 9909 3441 9913
rect 3445 9909 3446 9913
rect 3450 9909 3451 9913
rect 3410 9908 3455 9909
rect 3410 9904 3411 9908
rect 3415 9904 3416 9908
rect 3420 9904 3421 9908
rect 3425 9904 3426 9908
rect 3430 9904 3431 9908
rect 3435 9904 3436 9908
rect 3440 9904 3441 9908
rect 3445 9904 3446 9908
rect 3450 9904 3451 9908
rect 3410 9903 3455 9904
rect 3410 9899 3411 9903
rect 3415 9899 3416 9903
rect 3420 9899 3421 9903
rect 3425 9899 3426 9903
rect 3430 9899 3431 9903
rect 3435 9899 3436 9903
rect 3440 9899 3441 9903
rect 3445 9899 3446 9903
rect 3450 9899 3451 9903
rect 3410 9898 3455 9899
rect 3410 9894 3411 9898
rect 3415 9894 3416 9898
rect 3420 9894 3421 9898
rect 3425 9894 3426 9898
rect 3430 9894 3431 9898
rect 3435 9894 3436 9898
rect 3440 9894 3441 9898
rect 3445 9894 3446 9898
rect 3450 9894 3451 9898
rect 3410 9893 3455 9894
rect 3410 9889 3411 9893
rect 3415 9889 3416 9893
rect 3420 9889 3421 9893
rect 3425 9889 3426 9893
rect 3430 9889 3431 9893
rect 3435 9889 3436 9893
rect 3440 9889 3441 9893
rect 3445 9889 3446 9893
rect 3450 9889 3451 9893
rect 3410 9888 3455 9889
rect 3410 9884 3411 9888
rect 3415 9884 3416 9888
rect 3420 9884 3421 9888
rect 3425 9884 3426 9888
rect 3430 9884 3431 9888
rect 3435 9884 3436 9888
rect 3440 9884 3441 9888
rect 3445 9884 3446 9888
rect 3450 9884 3451 9888
rect 3410 9883 3455 9884
rect 3410 9879 3411 9883
rect 3415 9879 3416 9883
rect 3420 9879 3421 9883
rect 3425 9879 3426 9883
rect 3430 9879 3431 9883
rect 3435 9879 3436 9883
rect 3440 9879 3441 9883
rect 3445 9879 3446 9883
rect 3450 9879 3451 9883
rect 3410 9878 3455 9879
rect 3410 9874 3411 9878
rect 3415 9874 3416 9878
rect 3420 9874 3421 9878
rect 3425 9874 3426 9878
rect 3430 9874 3431 9878
rect 3435 9874 3436 9878
rect 3440 9874 3441 9878
rect 3445 9874 3446 9878
rect 3450 9874 3451 9878
rect 3410 9873 3455 9874
rect 3410 9869 3411 9873
rect 3415 9869 3416 9873
rect 3420 9869 3421 9873
rect 3425 9869 3426 9873
rect 3430 9869 3431 9873
rect 3435 9869 3436 9873
rect 3440 9869 3441 9873
rect 3445 9869 3446 9873
rect 3450 9869 3451 9873
rect 3410 9868 3455 9869
rect 3410 9864 3411 9868
rect 3415 9864 3416 9868
rect 3420 9864 3421 9868
rect 3425 9864 3426 9868
rect 3430 9864 3431 9868
rect 3435 9864 3436 9868
rect 3440 9864 3441 9868
rect 3445 9864 3446 9868
rect 3450 9864 3451 9868
rect 3463 9948 3467 9949
rect 3463 9943 3467 9944
rect 3463 9938 3467 9939
rect 3463 9933 3467 9934
rect 3463 9928 3467 9929
rect 3463 9923 3467 9924
rect 3463 9918 3467 9919
rect 3463 9913 3467 9914
rect 3463 9908 3467 9909
rect 3463 9903 3467 9904
rect 3463 9898 3467 9899
rect 3463 9893 3467 9894
rect 3463 9888 3467 9889
rect 3463 9883 3467 9884
rect 3463 9878 3467 9879
rect 3463 9873 3467 9874
rect 3463 9868 3467 9869
rect 3399 9863 3403 9864
rect 3399 9856 3403 9859
rect 3463 9863 3467 9864
rect 3463 9856 3467 9859
rect 3403 9848 3406 9856
rect 3410 9848 3411 9856
rect 3415 9848 3416 9856
rect 3420 9848 3421 9856
rect 3425 9848 3426 9856
rect 3430 9848 3431 9856
rect 3435 9848 3436 9856
rect 3440 9848 3441 9856
rect 3445 9848 3446 9856
rect 3450 9848 3451 9856
rect 3455 9848 3456 9856
rect 3460 9848 3463 9856
rect 3476 9963 3480 9964
rect 3476 9958 3480 9959
rect 3476 9953 3480 9954
rect 3476 9948 3480 9949
rect 3476 9943 3480 9944
rect 3476 9938 3480 9939
rect 3476 9933 3480 9934
rect 3476 9928 3480 9929
rect 3476 9923 3480 9924
rect 3476 9918 3480 9919
rect 3476 9913 3480 9914
rect 3476 9908 3480 9909
rect 3476 9903 3480 9904
rect 3476 9898 3480 9899
rect 3476 9893 3480 9894
rect 3476 9888 3480 9889
rect 3476 9883 3480 9884
rect 3476 9878 3480 9879
rect 3476 9873 3480 9874
rect 3476 9868 3480 9869
rect 3476 9863 3480 9864
rect 3476 9858 3480 9859
rect 3476 9853 3480 9854
rect 3476 9848 3480 9849
rect 3386 9843 3390 9844
rect 3476 9843 3480 9844
rect 3390 9839 3391 9843
rect 3395 9839 3396 9843
rect 3400 9839 3401 9843
rect 3405 9839 3406 9843
rect 3410 9839 3411 9843
rect 3415 9839 3416 9843
rect 3420 9839 3421 9843
rect 3425 9839 3426 9843
rect 3430 9839 3431 9843
rect 3435 9839 3436 9843
rect 3440 9839 3441 9843
rect 3445 9839 3446 9843
rect 3450 9839 3451 9843
rect 3455 9839 3456 9843
rect 3460 9839 3461 9843
rect 3465 9839 3466 9843
rect 3470 9839 3471 9843
rect 3475 9839 3476 9843
rect 3539 9974 3540 9978
rect 3544 9974 3545 9978
rect 3549 9974 3550 9978
rect 3554 9974 3555 9978
rect 3559 9974 3560 9978
rect 3564 9974 3565 9978
rect 3569 9974 3570 9978
rect 3574 9974 3575 9978
rect 3579 9974 3580 9978
rect 3584 9974 3585 9978
rect 3589 9974 3590 9978
rect 3594 9974 3595 9978
rect 3599 9974 3600 9978
rect 3604 9974 3605 9978
rect 3609 9974 3610 9978
rect 3614 9974 3615 9978
rect 3619 9974 3620 9978
rect 3624 9974 3625 9978
rect 3535 9973 3539 9974
rect 3535 9968 3539 9969
rect 3625 9973 3629 9974
rect 3625 9968 3629 9969
rect 3535 9963 3539 9964
rect 3535 9958 3539 9959
rect 3535 9953 3539 9954
rect 3535 9948 3539 9949
rect 3535 9943 3539 9944
rect 3535 9938 3539 9939
rect 3535 9933 3539 9934
rect 3535 9928 3539 9929
rect 3535 9923 3539 9924
rect 3535 9918 3539 9919
rect 3535 9913 3539 9914
rect 3535 9908 3539 9909
rect 3535 9903 3539 9904
rect 3535 9898 3539 9899
rect 3535 9893 3539 9894
rect 3535 9888 3539 9889
rect 3535 9883 3539 9884
rect 3535 9878 3539 9879
rect 3535 9873 3539 9874
rect 3535 9868 3539 9869
rect 3535 9863 3539 9864
rect 3535 9858 3539 9859
rect 3535 9853 3539 9854
rect 3535 9848 3539 9849
rect 3552 9961 3555 9965
rect 3559 9961 3560 9965
rect 3564 9961 3565 9965
rect 3569 9961 3570 9965
rect 3574 9961 3575 9965
rect 3579 9961 3580 9965
rect 3584 9961 3585 9965
rect 3589 9961 3590 9965
rect 3594 9961 3595 9965
rect 3599 9961 3600 9965
rect 3604 9961 3605 9965
rect 3609 9961 3612 9965
rect 3548 9958 3552 9961
rect 3548 9953 3552 9954
rect 3612 9958 3616 9961
rect 3612 9953 3616 9954
rect 3548 9948 3552 9949
rect 3548 9943 3552 9944
rect 3548 9938 3552 9939
rect 3548 9933 3552 9934
rect 3548 9928 3552 9929
rect 3548 9923 3552 9924
rect 3548 9918 3552 9919
rect 3548 9913 3552 9914
rect 3548 9908 3552 9909
rect 3548 9903 3552 9904
rect 3548 9898 3552 9899
rect 3548 9893 3552 9894
rect 3548 9888 3552 9889
rect 3548 9883 3552 9884
rect 3548 9878 3552 9879
rect 3548 9873 3552 9874
rect 3548 9868 3552 9869
rect 3564 9949 3565 9953
rect 3569 9949 3570 9953
rect 3574 9949 3575 9953
rect 3579 9949 3580 9953
rect 3584 9949 3585 9953
rect 3589 9949 3590 9953
rect 3594 9949 3595 9953
rect 3599 9949 3600 9953
rect 3560 9948 3604 9949
rect 3564 9944 3565 9948
rect 3569 9944 3570 9948
rect 3574 9944 3575 9948
rect 3579 9944 3580 9948
rect 3584 9944 3585 9948
rect 3589 9944 3590 9948
rect 3594 9944 3595 9948
rect 3599 9944 3600 9948
rect 3560 9943 3604 9944
rect 3564 9939 3565 9943
rect 3569 9939 3570 9943
rect 3574 9939 3575 9943
rect 3579 9939 3580 9943
rect 3584 9939 3585 9943
rect 3589 9939 3590 9943
rect 3594 9939 3595 9943
rect 3599 9939 3600 9943
rect 3560 9938 3604 9939
rect 3564 9934 3565 9938
rect 3569 9934 3570 9938
rect 3574 9934 3575 9938
rect 3579 9934 3580 9938
rect 3584 9934 3585 9938
rect 3589 9934 3590 9938
rect 3594 9934 3595 9938
rect 3599 9934 3600 9938
rect 3560 9933 3604 9934
rect 3564 9929 3565 9933
rect 3569 9929 3570 9933
rect 3574 9929 3575 9933
rect 3579 9929 3580 9933
rect 3584 9929 3585 9933
rect 3589 9929 3590 9933
rect 3594 9929 3595 9933
rect 3599 9929 3600 9933
rect 3560 9928 3604 9929
rect 3564 9924 3565 9928
rect 3569 9924 3570 9928
rect 3574 9924 3575 9928
rect 3579 9924 3580 9928
rect 3584 9924 3585 9928
rect 3589 9924 3590 9928
rect 3594 9924 3595 9928
rect 3599 9924 3600 9928
rect 3560 9923 3604 9924
rect 3564 9919 3565 9923
rect 3569 9919 3570 9923
rect 3574 9919 3575 9923
rect 3579 9919 3580 9923
rect 3584 9919 3585 9923
rect 3589 9919 3590 9923
rect 3594 9919 3595 9923
rect 3599 9919 3600 9923
rect 3560 9918 3604 9919
rect 3564 9914 3565 9918
rect 3569 9914 3570 9918
rect 3574 9914 3575 9918
rect 3579 9914 3580 9918
rect 3584 9914 3585 9918
rect 3589 9914 3590 9918
rect 3594 9914 3595 9918
rect 3599 9914 3600 9918
rect 3560 9913 3604 9914
rect 3564 9909 3565 9913
rect 3569 9909 3570 9913
rect 3574 9909 3575 9913
rect 3579 9909 3580 9913
rect 3584 9909 3585 9913
rect 3589 9909 3590 9913
rect 3594 9909 3595 9913
rect 3599 9909 3600 9913
rect 3560 9908 3604 9909
rect 3564 9904 3565 9908
rect 3569 9904 3570 9908
rect 3574 9904 3575 9908
rect 3579 9904 3580 9908
rect 3584 9904 3585 9908
rect 3589 9904 3590 9908
rect 3594 9904 3595 9908
rect 3599 9904 3600 9908
rect 3560 9903 3604 9904
rect 3564 9899 3565 9903
rect 3569 9899 3570 9903
rect 3574 9899 3575 9903
rect 3579 9899 3580 9903
rect 3584 9899 3585 9903
rect 3589 9899 3590 9903
rect 3594 9899 3595 9903
rect 3599 9899 3600 9903
rect 3560 9898 3604 9899
rect 3564 9894 3565 9898
rect 3569 9894 3570 9898
rect 3574 9894 3575 9898
rect 3579 9894 3580 9898
rect 3584 9894 3585 9898
rect 3589 9894 3590 9898
rect 3594 9894 3595 9898
rect 3599 9894 3600 9898
rect 3560 9893 3604 9894
rect 3564 9889 3565 9893
rect 3569 9889 3570 9893
rect 3574 9889 3575 9893
rect 3579 9889 3580 9893
rect 3584 9889 3585 9893
rect 3589 9889 3590 9893
rect 3594 9889 3595 9893
rect 3599 9889 3600 9893
rect 3560 9888 3604 9889
rect 3564 9884 3565 9888
rect 3569 9884 3570 9888
rect 3574 9884 3575 9888
rect 3579 9884 3580 9888
rect 3584 9884 3585 9888
rect 3589 9884 3590 9888
rect 3594 9884 3595 9888
rect 3599 9884 3600 9888
rect 3560 9883 3604 9884
rect 3564 9879 3565 9883
rect 3569 9879 3570 9883
rect 3574 9879 3575 9883
rect 3579 9879 3580 9883
rect 3584 9879 3585 9883
rect 3589 9879 3590 9883
rect 3594 9879 3595 9883
rect 3599 9879 3600 9883
rect 3560 9878 3604 9879
rect 3564 9874 3565 9878
rect 3569 9874 3570 9878
rect 3574 9874 3575 9878
rect 3579 9874 3580 9878
rect 3584 9874 3585 9878
rect 3589 9874 3590 9878
rect 3594 9874 3595 9878
rect 3599 9874 3600 9878
rect 3560 9873 3604 9874
rect 3564 9869 3565 9873
rect 3569 9869 3570 9873
rect 3574 9869 3575 9873
rect 3579 9869 3580 9873
rect 3584 9869 3585 9873
rect 3589 9869 3590 9873
rect 3594 9869 3595 9873
rect 3599 9869 3600 9873
rect 3560 9868 3604 9869
rect 3564 9864 3565 9868
rect 3569 9864 3570 9868
rect 3574 9864 3575 9868
rect 3579 9864 3580 9868
rect 3584 9864 3585 9868
rect 3589 9864 3590 9868
rect 3594 9864 3595 9868
rect 3599 9864 3600 9868
rect 3612 9948 3616 9949
rect 3612 9943 3616 9944
rect 3612 9938 3616 9939
rect 3612 9933 3616 9934
rect 3612 9928 3616 9929
rect 3612 9923 3616 9924
rect 3612 9918 3616 9919
rect 3612 9913 3616 9914
rect 3612 9908 3616 9909
rect 3612 9903 3616 9904
rect 3612 9898 3616 9899
rect 3612 9893 3616 9894
rect 3612 9888 3616 9889
rect 3612 9883 3616 9884
rect 3612 9878 3616 9879
rect 3612 9873 3616 9874
rect 3612 9868 3616 9869
rect 3548 9863 3552 9864
rect 3548 9856 3552 9859
rect 3612 9863 3616 9864
rect 3612 9856 3616 9859
rect 3552 9848 3555 9856
rect 3559 9848 3560 9856
rect 3564 9848 3565 9856
rect 3569 9848 3570 9856
rect 3574 9848 3575 9856
rect 3579 9848 3580 9856
rect 3584 9848 3585 9856
rect 3589 9848 3590 9856
rect 3594 9848 3595 9856
rect 3599 9848 3600 9856
rect 3604 9848 3605 9856
rect 3609 9848 3612 9856
rect 3625 9963 3629 9964
rect 3625 9958 3629 9959
rect 3625 9953 3629 9954
rect 3625 9948 3629 9949
rect 3625 9943 3629 9944
rect 3625 9938 3629 9939
rect 3625 9933 3629 9934
rect 3625 9928 3629 9929
rect 3625 9923 3629 9924
rect 3625 9918 3629 9919
rect 3625 9913 3629 9914
rect 3625 9908 3629 9909
rect 3625 9903 3629 9904
rect 3625 9898 3629 9899
rect 3625 9893 3629 9894
rect 3625 9888 3629 9889
rect 3625 9883 3629 9884
rect 3625 9878 3629 9879
rect 3625 9873 3629 9874
rect 3625 9868 3629 9869
rect 3625 9863 3629 9864
rect 3625 9858 3629 9859
rect 3625 9853 3629 9854
rect 3625 9848 3629 9849
rect 3535 9843 3539 9844
rect 3625 9843 3629 9844
rect 3539 9839 3540 9843
rect 3544 9839 3545 9843
rect 3549 9839 3550 9843
rect 3554 9839 3555 9843
rect 3559 9839 3560 9843
rect 3564 9839 3565 9843
rect 3569 9839 3570 9843
rect 3574 9839 3575 9843
rect 3579 9839 3580 9843
rect 3584 9839 3585 9843
rect 3589 9839 3590 9843
rect 3594 9839 3595 9843
rect 3599 9839 3600 9843
rect 3604 9839 3605 9843
rect 3609 9839 3610 9843
rect 3614 9839 3615 9843
rect 3619 9839 3620 9843
rect 3624 9839 3625 9843
rect 3327 9711 3353 9715
rect 3357 9711 3358 9715
rect 3362 9711 3379 9715
rect 3423 9722 3479 9839
rect 3538 9802 3594 9839
rect 3526 9800 3594 9802
rect 3526 9796 3527 9800
rect 3531 9796 3532 9800
rect 3536 9796 3594 9800
rect 3526 9795 3594 9796
rect 3526 9791 3527 9795
rect 3531 9791 3532 9795
rect 3536 9791 3594 9795
rect 3526 9790 3594 9791
rect 3526 9786 3527 9790
rect 3531 9786 3532 9790
rect 3536 9786 3594 9790
rect 3526 9785 3594 9786
rect 3526 9781 3527 9785
rect 3531 9781 3532 9785
rect 3536 9781 3594 9785
rect 3526 9780 3594 9781
rect 3526 9776 3527 9780
rect 3531 9776 3532 9780
rect 3536 9776 3594 9780
rect 3526 9775 3594 9776
rect 3526 9771 3527 9775
rect 3531 9771 3532 9775
rect 3536 9771 3594 9775
rect 3526 9770 3594 9771
rect 3526 9766 3527 9770
rect 3531 9766 3532 9770
rect 3536 9766 3594 9770
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3482 9761 3501 9762
rect 3486 9757 3487 9761
rect 3491 9757 3492 9761
rect 3496 9757 3497 9761
rect 3482 9756 3501 9757
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3482 9751 3501 9752
rect 3486 9747 3487 9751
rect 3491 9747 3492 9751
rect 3496 9747 3497 9751
rect 3482 9746 3501 9747
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3482 9741 3501 9742
rect 3486 9737 3487 9741
rect 3491 9737 3492 9741
rect 3496 9737 3497 9741
rect 3482 9736 3501 9737
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3526 9765 3594 9766
rect 3526 9761 3527 9765
rect 3531 9761 3532 9765
rect 3536 9761 3594 9765
rect 3526 9760 3594 9761
rect 3526 9756 3527 9760
rect 3531 9756 3532 9760
rect 3536 9756 3594 9760
rect 3526 9755 3594 9756
rect 3526 9751 3527 9755
rect 3531 9751 3532 9755
rect 3536 9751 3594 9755
rect 3526 9750 3594 9751
rect 3526 9746 3527 9750
rect 3531 9746 3532 9750
rect 3536 9746 3594 9750
rect 3526 9745 3594 9746
rect 3526 9741 3527 9745
rect 3531 9741 3532 9745
rect 3536 9741 3594 9745
rect 3526 9740 3594 9741
rect 3526 9736 3527 9740
rect 3531 9736 3532 9740
rect 3536 9736 3594 9740
rect 3526 9734 3594 9736
rect 3634 9795 3688 9981
rect 3699 9974 3700 9978
rect 3704 9974 3705 9978
rect 3709 9974 3710 9978
rect 3714 9974 3715 9978
rect 3719 9974 3720 9978
rect 3724 9974 3725 9978
rect 3729 9974 3730 9978
rect 3734 9974 3735 9978
rect 3739 9974 3740 9978
rect 3744 9974 3745 9978
rect 3749 9974 3750 9978
rect 3754 9974 3755 9978
rect 3759 9974 3760 9978
rect 3764 9974 3765 9978
rect 3769 9974 3770 9978
rect 3774 9974 3775 9978
rect 3779 9974 3780 9978
rect 3784 9974 3785 9978
rect 3695 9973 3699 9974
rect 3695 9968 3699 9969
rect 3785 9973 3789 9974
rect 3785 9968 3789 9969
rect 3695 9963 3699 9964
rect 3695 9958 3699 9959
rect 3695 9953 3699 9954
rect 3695 9948 3699 9949
rect 3695 9943 3699 9944
rect 3695 9938 3699 9939
rect 3695 9933 3699 9934
rect 3695 9928 3699 9929
rect 3695 9923 3699 9924
rect 3695 9918 3699 9919
rect 3695 9913 3699 9914
rect 3695 9908 3699 9909
rect 3695 9903 3699 9904
rect 3695 9898 3699 9899
rect 3695 9893 3699 9894
rect 3695 9888 3699 9889
rect 3695 9883 3699 9884
rect 3695 9878 3699 9879
rect 3695 9873 3699 9874
rect 3695 9868 3699 9869
rect 3695 9863 3699 9864
rect 3695 9858 3699 9859
rect 3695 9853 3699 9854
rect 3695 9848 3699 9849
rect 3712 9961 3715 9965
rect 3719 9961 3720 9965
rect 3724 9961 3725 9965
rect 3729 9961 3730 9965
rect 3734 9961 3735 9965
rect 3739 9961 3740 9965
rect 3744 9961 3745 9965
rect 3749 9961 3750 9965
rect 3754 9961 3755 9965
rect 3759 9961 3760 9965
rect 3764 9961 3765 9965
rect 3769 9961 3772 9965
rect 3708 9958 3712 9961
rect 3708 9953 3712 9954
rect 3772 9958 3776 9961
rect 3772 9953 3776 9954
rect 3708 9948 3712 9949
rect 3708 9943 3712 9944
rect 3708 9938 3712 9939
rect 3708 9933 3712 9934
rect 3708 9928 3712 9929
rect 3708 9923 3712 9924
rect 3708 9918 3712 9919
rect 3708 9913 3712 9914
rect 3708 9908 3712 9909
rect 3708 9903 3712 9904
rect 3708 9898 3712 9899
rect 3708 9893 3712 9894
rect 3708 9888 3712 9889
rect 3708 9883 3712 9884
rect 3708 9878 3712 9879
rect 3708 9873 3712 9874
rect 3708 9868 3712 9869
rect 3719 9949 3720 9953
rect 3724 9949 3725 9953
rect 3729 9949 3730 9953
rect 3734 9949 3735 9953
rect 3739 9949 3740 9953
rect 3744 9949 3745 9953
rect 3749 9949 3750 9953
rect 3754 9949 3755 9953
rect 3759 9949 3760 9953
rect 3719 9948 3764 9949
rect 3719 9944 3720 9948
rect 3724 9944 3725 9948
rect 3729 9944 3730 9948
rect 3734 9944 3735 9948
rect 3739 9944 3740 9948
rect 3744 9944 3745 9948
rect 3749 9944 3750 9948
rect 3754 9944 3755 9948
rect 3759 9944 3760 9948
rect 3719 9943 3764 9944
rect 3719 9939 3720 9943
rect 3724 9939 3725 9943
rect 3729 9939 3730 9943
rect 3734 9939 3735 9943
rect 3739 9939 3740 9943
rect 3744 9939 3745 9943
rect 3749 9939 3750 9943
rect 3754 9939 3755 9943
rect 3759 9939 3760 9943
rect 3719 9938 3764 9939
rect 3719 9934 3720 9938
rect 3724 9934 3725 9938
rect 3729 9934 3730 9938
rect 3734 9934 3735 9938
rect 3739 9934 3740 9938
rect 3744 9934 3745 9938
rect 3749 9934 3750 9938
rect 3754 9934 3755 9938
rect 3759 9934 3760 9938
rect 3719 9933 3764 9934
rect 3719 9929 3720 9933
rect 3724 9929 3725 9933
rect 3729 9929 3730 9933
rect 3734 9929 3735 9933
rect 3739 9929 3740 9933
rect 3744 9929 3745 9933
rect 3749 9929 3750 9933
rect 3754 9929 3755 9933
rect 3759 9929 3760 9933
rect 3719 9928 3764 9929
rect 3719 9924 3720 9928
rect 3724 9924 3725 9928
rect 3729 9924 3730 9928
rect 3734 9924 3735 9928
rect 3739 9924 3740 9928
rect 3744 9924 3745 9928
rect 3749 9924 3750 9928
rect 3754 9924 3755 9928
rect 3759 9924 3760 9928
rect 3719 9923 3764 9924
rect 3719 9919 3720 9923
rect 3724 9919 3725 9923
rect 3729 9919 3730 9923
rect 3734 9919 3735 9923
rect 3739 9919 3740 9923
rect 3744 9919 3745 9923
rect 3749 9919 3750 9923
rect 3754 9919 3755 9923
rect 3759 9919 3760 9923
rect 3719 9918 3764 9919
rect 3719 9914 3720 9918
rect 3724 9914 3725 9918
rect 3729 9914 3730 9918
rect 3734 9914 3735 9918
rect 3739 9914 3740 9918
rect 3744 9914 3745 9918
rect 3749 9914 3750 9918
rect 3754 9914 3755 9918
rect 3759 9914 3760 9918
rect 3719 9913 3764 9914
rect 3719 9909 3720 9913
rect 3724 9909 3725 9913
rect 3729 9909 3730 9913
rect 3734 9909 3735 9913
rect 3739 9909 3740 9913
rect 3744 9909 3745 9913
rect 3749 9909 3750 9913
rect 3754 9909 3755 9913
rect 3759 9909 3760 9913
rect 3719 9908 3764 9909
rect 3719 9904 3720 9908
rect 3724 9904 3725 9908
rect 3729 9904 3730 9908
rect 3734 9904 3735 9908
rect 3739 9904 3740 9908
rect 3744 9904 3745 9908
rect 3749 9904 3750 9908
rect 3754 9904 3755 9908
rect 3759 9904 3760 9908
rect 3719 9903 3764 9904
rect 3719 9899 3720 9903
rect 3724 9899 3725 9903
rect 3729 9899 3730 9903
rect 3734 9899 3735 9903
rect 3739 9899 3740 9903
rect 3744 9899 3745 9903
rect 3749 9899 3750 9903
rect 3754 9899 3755 9903
rect 3759 9899 3760 9903
rect 3719 9898 3764 9899
rect 3719 9894 3720 9898
rect 3724 9894 3725 9898
rect 3729 9894 3730 9898
rect 3734 9894 3735 9898
rect 3739 9894 3740 9898
rect 3744 9894 3745 9898
rect 3749 9894 3750 9898
rect 3754 9894 3755 9898
rect 3759 9894 3760 9898
rect 3719 9893 3764 9894
rect 3719 9889 3720 9893
rect 3724 9889 3725 9893
rect 3729 9889 3730 9893
rect 3734 9889 3735 9893
rect 3739 9889 3740 9893
rect 3744 9889 3745 9893
rect 3749 9889 3750 9893
rect 3754 9889 3755 9893
rect 3759 9889 3760 9893
rect 3719 9888 3764 9889
rect 3719 9884 3720 9888
rect 3724 9884 3725 9888
rect 3729 9884 3730 9888
rect 3734 9884 3735 9888
rect 3739 9884 3740 9888
rect 3744 9884 3745 9888
rect 3749 9884 3750 9888
rect 3754 9884 3755 9888
rect 3759 9884 3760 9888
rect 3719 9883 3764 9884
rect 3719 9879 3720 9883
rect 3724 9879 3725 9883
rect 3729 9879 3730 9883
rect 3734 9879 3735 9883
rect 3739 9879 3740 9883
rect 3744 9879 3745 9883
rect 3749 9879 3750 9883
rect 3754 9879 3755 9883
rect 3759 9879 3760 9883
rect 3719 9878 3764 9879
rect 3719 9874 3720 9878
rect 3724 9874 3725 9878
rect 3729 9874 3730 9878
rect 3734 9874 3735 9878
rect 3739 9874 3740 9878
rect 3744 9874 3745 9878
rect 3749 9874 3750 9878
rect 3754 9874 3755 9878
rect 3759 9874 3760 9878
rect 3719 9873 3764 9874
rect 3719 9869 3720 9873
rect 3724 9869 3725 9873
rect 3729 9869 3730 9873
rect 3734 9869 3735 9873
rect 3739 9869 3740 9873
rect 3744 9869 3745 9873
rect 3749 9869 3750 9873
rect 3754 9869 3755 9873
rect 3759 9869 3760 9873
rect 3719 9868 3764 9869
rect 3719 9864 3720 9868
rect 3724 9864 3725 9868
rect 3729 9864 3730 9868
rect 3734 9864 3735 9868
rect 3739 9864 3740 9868
rect 3744 9864 3745 9868
rect 3749 9864 3750 9868
rect 3754 9864 3755 9868
rect 3759 9864 3760 9868
rect 3772 9948 3776 9949
rect 3772 9943 3776 9944
rect 3772 9938 3776 9939
rect 3772 9933 3776 9934
rect 3772 9928 3776 9929
rect 3772 9923 3776 9924
rect 3772 9918 3776 9919
rect 3772 9913 3776 9914
rect 3772 9908 3776 9909
rect 3772 9903 3776 9904
rect 3772 9898 3776 9899
rect 3772 9893 3776 9894
rect 3772 9888 3776 9889
rect 3772 9883 3776 9884
rect 3772 9878 3776 9879
rect 3772 9873 3776 9874
rect 3772 9868 3776 9869
rect 3708 9863 3712 9864
rect 3708 9856 3712 9859
rect 3772 9863 3776 9864
rect 3772 9856 3776 9859
rect 3712 9848 3715 9856
rect 3719 9848 3720 9856
rect 3724 9848 3725 9856
rect 3729 9848 3730 9856
rect 3734 9848 3735 9856
rect 3739 9848 3740 9856
rect 3744 9848 3745 9856
rect 3749 9848 3750 9856
rect 3754 9848 3755 9856
rect 3759 9848 3760 9856
rect 3764 9848 3765 9856
rect 3769 9848 3772 9856
rect 3785 9963 3789 9964
rect 3785 9958 3789 9959
rect 3785 9953 3789 9954
rect 3785 9948 3789 9949
rect 3785 9943 3789 9944
rect 3785 9938 3789 9939
rect 3785 9933 3789 9934
rect 3785 9928 3789 9929
rect 3785 9923 3789 9924
rect 3785 9918 3789 9919
rect 3785 9913 3789 9914
rect 3785 9908 3789 9909
rect 3785 9903 3789 9904
rect 3785 9898 3789 9899
rect 3785 9893 3789 9894
rect 3785 9888 3789 9889
rect 3785 9883 3789 9884
rect 3785 9878 3789 9879
rect 3785 9873 3789 9874
rect 3785 9868 3789 9869
rect 3785 9863 3789 9864
rect 3785 9858 3789 9859
rect 3785 9853 3789 9854
rect 3785 9848 3789 9849
rect 3695 9843 3699 9844
rect 3785 9843 3789 9844
rect 3699 9839 3700 9843
rect 3704 9839 3705 9843
rect 3709 9839 3710 9843
rect 3714 9839 3715 9843
rect 3719 9839 3720 9843
rect 3724 9839 3725 9843
rect 3729 9839 3730 9843
rect 3734 9839 3735 9843
rect 3739 9839 3740 9843
rect 3744 9839 3745 9843
rect 3749 9839 3750 9843
rect 3754 9839 3755 9843
rect 3759 9839 3760 9843
rect 3764 9839 3765 9843
rect 3769 9839 3770 9843
rect 3774 9839 3775 9843
rect 3779 9839 3780 9843
rect 3784 9839 3785 9843
rect 3848 9974 3849 9978
rect 3853 9974 3854 9978
rect 3858 9974 3859 9978
rect 3863 9974 3864 9978
rect 3868 9974 3869 9978
rect 3873 9974 3874 9978
rect 3878 9974 3879 9978
rect 3883 9974 3884 9978
rect 3888 9974 3889 9978
rect 3893 9974 3894 9978
rect 3898 9974 3899 9978
rect 3903 9974 3904 9978
rect 3908 9974 3909 9978
rect 3913 9974 3914 9978
rect 3918 9974 3919 9978
rect 3923 9974 3924 9978
rect 3928 9974 3929 9978
rect 3933 9974 3934 9978
rect 3844 9973 3848 9974
rect 3844 9968 3848 9969
rect 3934 9973 3938 9974
rect 3934 9968 3938 9969
rect 3844 9963 3848 9964
rect 3844 9958 3848 9959
rect 3844 9953 3848 9954
rect 3844 9948 3848 9949
rect 3844 9943 3848 9944
rect 3844 9938 3848 9939
rect 3844 9933 3848 9934
rect 3844 9928 3848 9929
rect 3844 9923 3848 9924
rect 3844 9918 3848 9919
rect 3844 9913 3848 9914
rect 3844 9908 3848 9909
rect 3844 9903 3848 9904
rect 3844 9898 3848 9899
rect 3844 9893 3848 9894
rect 3844 9888 3848 9889
rect 3844 9883 3848 9884
rect 3844 9878 3848 9879
rect 3844 9873 3848 9874
rect 3844 9868 3848 9869
rect 3844 9863 3848 9864
rect 3844 9858 3848 9859
rect 3844 9853 3848 9854
rect 3844 9848 3848 9849
rect 3861 9961 3864 9965
rect 3868 9961 3869 9965
rect 3873 9961 3874 9965
rect 3878 9961 3879 9965
rect 3883 9961 3884 9965
rect 3888 9961 3889 9965
rect 3893 9961 3894 9965
rect 3898 9961 3899 9965
rect 3903 9961 3904 9965
rect 3908 9961 3909 9965
rect 3913 9961 3914 9965
rect 3918 9961 3921 9965
rect 3857 9958 3861 9961
rect 3857 9953 3861 9954
rect 3921 9958 3925 9961
rect 3921 9953 3925 9954
rect 3857 9948 3861 9949
rect 3857 9943 3861 9944
rect 3857 9938 3861 9939
rect 3857 9933 3861 9934
rect 3857 9928 3861 9929
rect 3857 9923 3861 9924
rect 3857 9918 3861 9919
rect 3857 9913 3861 9914
rect 3857 9908 3861 9909
rect 3857 9903 3861 9904
rect 3857 9898 3861 9899
rect 3857 9893 3861 9894
rect 3857 9888 3861 9889
rect 3857 9883 3861 9884
rect 3857 9878 3861 9879
rect 3857 9873 3861 9874
rect 3857 9868 3861 9869
rect 3873 9949 3874 9953
rect 3878 9949 3879 9953
rect 3883 9949 3884 9953
rect 3888 9949 3889 9953
rect 3893 9949 3894 9953
rect 3898 9949 3899 9953
rect 3903 9949 3904 9953
rect 3908 9949 3909 9953
rect 3869 9948 3913 9949
rect 3873 9944 3874 9948
rect 3878 9944 3879 9948
rect 3883 9944 3884 9948
rect 3888 9944 3889 9948
rect 3893 9944 3894 9948
rect 3898 9944 3899 9948
rect 3903 9944 3904 9948
rect 3908 9944 3909 9948
rect 3869 9943 3913 9944
rect 3873 9939 3874 9943
rect 3878 9939 3879 9943
rect 3883 9939 3884 9943
rect 3888 9939 3889 9943
rect 3893 9939 3894 9943
rect 3898 9939 3899 9943
rect 3903 9939 3904 9943
rect 3908 9939 3909 9943
rect 3869 9938 3913 9939
rect 3873 9934 3874 9938
rect 3878 9934 3879 9938
rect 3883 9934 3884 9938
rect 3888 9934 3889 9938
rect 3893 9934 3894 9938
rect 3898 9934 3899 9938
rect 3903 9934 3904 9938
rect 3908 9934 3909 9938
rect 3869 9933 3913 9934
rect 3873 9929 3874 9933
rect 3878 9929 3879 9933
rect 3883 9929 3884 9933
rect 3888 9929 3889 9933
rect 3893 9929 3894 9933
rect 3898 9929 3899 9933
rect 3903 9929 3904 9933
rect 3908 9929 3909 9933
rect 3869 9928 3913 9929
rect 3873 9924 3874 9928
rect 3878 9924 3879 9928
rect 3883 9924 3884 9928
rect 3888 9924 3889 9928
rect 3893 9924 3894 9928
rect 3898 9924 3899 9928
rect 3903 9924 3904 9928
rect 3908 9924 3909 9928
rect 3869 9923 3913 9924
rect 3873 9919 3874 9923
rect 3878 9919 3879 9923
rect 3883 9919 3884 9923
rect 3888 9919 3889 9923
rect 3893 9919 3894 9923
rect 3898 9919 3899 9923
rect 3903 9919 3904 9923
rect 3908 9919 3909 9923
rect 3869 9918 3913 9919
rect 3873 9914 3874 9918
rect 3878 9914 3879 9918
rect 3883 9914 3884 9918
rect 3888 9914 3889 9918
rect 3893 9914 3894 9918
rect 3898 9914 3899 9918
rect 3903 9914 3904 9918
rect 3908 9914 3909 9918
rect 3869 9913 3913 9914
rect 3873 9909 3874 9913
rect 3878 9909 3879 9913
rect 3883 9909 3884 9913
rect 3888 9909 3889 9913
rect 3893 9909 3894 9913
rect 3898 9909 3899 9913
rect 3903 9909 3904 9913
rect 3908 9909 3909 9913
rect 3869 9908 3913 9909
rect 3873 9904 3874 9908
rect 3878 9904 3879 9908
rect 3883 9904 3884 9908
rect 3888 9904 3889 9908
rect 3893 9904 3894 9908
rect 3898 9904 3899 9908
rect 3903 9904 3904 9908
rect 3908 9904 3909 9908
rect 3869 9903 3913 9904
rect 3873 9899 3874 9903
rect 3878 9899 3879 9903
rect 3883 9899 3884 9903
rect 3888 9899 3889 9903
rect 3893 9899 3894 9903
rect 3898 9899 3899 9903
rect 3903 9899 3904 9903
rect 3908 9899 3909 9903
rect 3869 9898 3913 9899
rect 3873 9894 3874 9898
rect 3878 9894 3879 9898
rect 3883 9894 3884 9898
rect 3888 9894 3889 9898
rect 3893 9894 3894 9898
rect 3898 9894 3899 9898
rect 3903 9894 3904 9898
rect 3908 9894 3909 9898
rect 3869 9893 3913 9894
rect 3873 9889 3874 9893
rect 3878 9889 3879 9893
rect 3883 9889 3884 9893
rect 3888 9889 3889 9893
rect 3893 9889 3894 9893
rect 3898 9889 3899 9893
rect 3903 9889 3904 9893
rect 3908 9889 3909 9893
rect 3869 9888 3913 9889
rect 3873 9884 3874 9888
rect 3878 9884 3879 9888
rect 3883 9884 3884 9888
rect 3888 9884 3889 9888
rect 3893 9884 3894 9888
rect 3898 9884 3899 9888
rect 3903 9884 3904 9888
rect 3908 9884 3909 9888
rect 3869 9883 3913 9884
rect 3873 9879 3874 9883
rect 3878 9879 3879 9883
rect 3883 9879 3884 9883
rect 3888 9879 3889 9883
rect 3893 9879 3894 9883
rect 3898 9879 3899 9883
rect 3903 9879 3904 9883
rect 3908 9879 3909 9883
rect 3869 9878 3913 9879
rect 3873 9874 3874 9878
rect 3878 9874 3879 9878
rect 3883 9874 3884 9878
rect 3888 9874 3889 9878
rect 3893 9874 3894 9878
rect 3898 9874 3899 9878
rect 3903 9874 3904 9878
rect 3908 9874 3909 9878
rect 3869 9873 3913 9874
rect 3873 9869 3874 9873
rect 3878 9869 3879 9873
rect 3883 9869 3884 9873
rect 3888 9869 3889 9873
rect 3893 9869 3894 9873
rect 3898 9869 3899 9873
rect 3903 9869 3904 9873
rect 3908 9869 3909 9873
rect 3869 9868 3913 9869
rect 3873 9864 3874 9868
rect 3878 9864 3879 9868
rect 3883 9864 3884 9868
rect 3888 9864 3889 9868
rect 3893 9864 3894 9868
rect 3898 9864 3899 9868
rect 3903 9864 3904 9868
rect 3908 9864 3909 9868
rect 3921 9948 3925 9949
rect 3921 9943 3925 9944
rect 3921 9938 3925 9939
rect 3921 9933 3925 9934
rect 3921 9928 3925 9929
rect 3921 9923 3925 9924
rect 3921 9918 3925 9919
rect 3921 9913 3925 9914
rect 3921 9908 3925 9909
rect 3921 9903 3925 9904
rect 3921 9898 3925 9899
rect 3921 9893 3925 9894
rect 3921 9888 3925 9889
rect 3921 9883 3925 9884
rect 3921 9878 3925 9879
rect 3921 9873 3925 9874
rect 3921 9868 3925 9869
rect 3857 9863 3861 9864
rect 3857 9856 3861 9859
rect 3921 9863 3925 9864
rect 3921 9856 3925 9859
rect 3861 9848 3864 9856
rect 3868 9848 3869 9856
rect 3873 9848 3874 9856
rect 3878 9848 3879 9856
rect 3883 9848 3884 9856
rect 3888 9848 3889 9856
rect 3893 9848 3894 9856
rect 3898 9848 3899 9856
rect 3903 9848 3904 9856
rect 3908 9848 3909 9856
rect 3913 9848 3914 9856
rect 3918 9848 3921 9856
rect 3934 9963 3938 9964
rect 3934 9958 3938 9959
rect 3934 9953 3938 9954
rect 3960 9961 3981 9981
rect 4008 9974 4009 9978
rect 4013 9974 4014 9978
rect 4018 9974 4019 9978
rect 4023 9974 4024 9978
rect 4028 9974 4029 9978
rect 4033 9974 4034 9978
rect 4038 9974 4039 9978
rect 4043 9974 4044 9978
rect 4048 9974 4049 9978
rect 4053 9974 4054 9978
rect 4058 9974 4059 9978
rect 4063 9974 4064 9978
rect 4068 9974 4069 9978
rect 4073 9974 4074 9978
rect 4078 9974 4079 9978
rect 4083 9974 4084 9978
rect 4088 9974 4089 9978
rect 4093 9974 4094 9978
rect 4004 9973 4008 9974
rect 4004 9968 4008 9969
rect 4094 9973 4098 9974
rect 4094 9968 4098 9969
rect 4004 9963 4008 9964
rect 4004 9958 4008 9959
rect 4004 9953 4008 9954
rect 3934 9948 3938 9949
rect 3934 9943 3938 9944
rect 3934 9938 3938 9939
rect 3934 9933 3938 9934
rect 3934 9928 3938 9929
rect 3934 9923 3938 9924
rect 3934 9918 3938 9919
rect 3934 9913 3938 9914
rect 3934 9908 3938 9909
rect 3934 9903 3938 9904
rect 3934 9898 3938 9899
rect 3934 9893 3938 9894
rect 3934 9888 3938 9889
rect 3934 9883 3938 9884
rect 4004 9948 4008 9949
rect 4004 9943 4008 9944
rect 4004 9938 4008 9939
rect 4004 9933 4008 9934
rect 4004 9928 4008 9929
rect 4004 9923 4008 9924
rect 4004 9918 4008 9919
rect 4004 9913 4008 9914
rect 4004 9908 4008 9909
rect 4004 9903 4008 9904
rect 4004 9898 4008 9899
rect 4004 9893 4008 9894
rect 4004 9888 4008 9889
rect 4004 9883 4008 9884
rect 3934 9878 3938 9879
rect 3934 9873 3938 9874
rect 3934 9868 3938 9869
rect 3934 9863 3938 9864
rect 3934 9858 3938 9859
rect 3934 9853 3938 9854
rect 3934 9848 3938 9849
rect 3844 9843 3848 9844
rect 3960 9846 3981 9874
rect 4004 9878 4008 9879
rect 4004 9873 4008 9874
rect 4004 9868 4008 9869
rect 4004 9863 4008 9864
rect 4004 9858 4008 9859
rect 4004 9853 4008 9854
rect 4004 9848 4008 9849
rect 4021 9961 4024 9965
rect 4028 9961 4029 9965
rect 4033 9961 4034 9965
rect 4038 9961 4039 9965
rect 4043 9961 4044 9965
rect 4048 9961 4049 9965
rect 4053 9961 4054 9965
rect 4058 9961 4059 9965
rect 4063 9961 4064 9965
rect 4068 9961 4069 9965
rect 4073 9961 4074 9965
rect 4078 9961 4081 9965
rect 4017 9958 4021 9961
rect 4017 9953 4021 9954
rect 4081 9958 4085 9961
rect 4081 9953 4085 9954
rect 4017 9948 4021 9949
rect 4017 9943 4021 9944
rect 4017 9938 4021 9939
rect 4017 9933 4021 9934
rect 4017 9928 4021 9929
rect 4017 9923 4021 9924
rect 4017 9918 4021 9919
rect 4017 9913 4021 9914
rect 4017 9908 4021 9909
rect 4017 9903 4021 9904
rect 4017 9898 4021 9899
rect 4017 9893 4021 9894
rect 4017 9888 4021 9889
rect 4017 9883 4021 9884
rect 4017 9878 4021 9879
rect 4017 9873 4021 9874
rect 4017 9868 4021 9869
rect 4028 9949 4029 9953
rect 4033 9949 4034 9953
rect 4038 9949 4039 9953
rect 4043 9949 4044 9953
rect 4048 9949 4049 9953
rect 4053 9949 4054 9953
rect 4058 9949 4059 9953
rect 4063 9949 4064 9953
rect 4068 9949 4069 9953
rect 4028 9948 4073 9949
rect 4028 9944 4029 9948
rect 4033 9944 4034 9948
rect 4038 9944 4039 9948
rect 4043 9944 4044 9948
rect 4048 9944 4049 9948
rect 4053 9944 4054 9948
rect 4058 9944 4059 9948
rect 4063 9944 4064 9948
rect 4068 9944 4069 9948
rect 4028 9943 4073 9944
rect 4028 9939 4029 9943
rect 4033 9939 4034 9943
rect 4038 9939 4039 9943
rect 4043 9939 4044 9943
rect 4048 9939 4049 9943
rect 4053 9939 4054 9943
rect 4058 9939 4059 9943
rect 4063 9939 4064 9943
rect 4068 9939 4069 9943
rect 4028 9938 4073 9939
rect 4028 9934 4029 9938
rect 4033 9934 4034 9938
rect 4038 9934 4039 9938
rect 4043 9934 4044 9938
rect 4048 9934 4049 9938
rect 4053 9934 4054 9938
rect 4058 9934 4059 9938
rect 4063 9934 4064 9938
rect 4068 9934 4069 9938
rect 4028 9933 4073 9934
rect 4028 9929 4029 9933
rect 4033 9929 4034 9933
rect 4038 9929 4039 9933
rect 4043 9929 4044 9933
rect 4048 9929 4049 9933
rect 4053 9929 4054 9933
rect 4058 9929 4059 9933
rect 4063 9929 4064 9933
rect 4068 9929 4069 9933
rect 4028 9928 4073 9929
rect 4028 9924 4029 9928
rect 4033 9924 4034 9928
rect 4038 9924 4039 9928
rect 4043 9924 4044 9928
rect 4048 9924 4049 9928
rect 4053 9924 4054 9928
rect 4058 9924 4059 9928
rect 4063 9924 4064 9928
rect 4068 9924 4069 9928
rect 4028 9923 4073 9924
rect 4028 9919 4029 9923
rect 4033 9919 4034 9923
rect 4038 9919 4039 9923
rect 4043 9919 4044 9923
rect 4048 9919 4049 9923
rect 4053 9919 4054 9923
rect 4058 9919 4059 9923
rect 4063 9919 4064 9923
rect 4068 9919 4069 9923
rect 4028 9918 4073 9919
rect 4028 9914 4029 9918
rect 4033 9914 4034 9918
rect 4038 9914 4039 9918
rect 4043 9914 4044 9918
rect 4048 9914 4049 9918
rect 4053 9914 4054 9918
rect 4058 9914 4059 9918
rect 4063 9914 4064 9918
rect 4068 9914 4069 9918
rect 4028 9913 4073 9914
rect 4028 9909 4029 9913
rect 4033 9909 4034 9913
rect 4038 9909 4039 9913
rect 4043 9909 4044 9913
rect 4048 9909 4049 9913
rect 4053 9909 4054 9913
rect 4058 9909 4059 9913
rect 4063 9909 4064 9913
rect 4068 9909 4069 9913
rect 4028 9908 4073 9909
rect 4028 9904 4029 9908
rect 4033 9904 4034 9908
rect 4038 9904 4039 9908
rect 4043 9904 4044 9908
rect 4048 9904 4049 9908
rect 4053 9904 4054 9908
rect 4058 9904 4059 9908
rect 4063 9904 4064 9908
rect 4068 9904 4069 9908
rect 4028 9903 4073 9904
rect 4028 9899 4029 9903
rect 4033 9899 4034 9903
rect 4038 9899 4039 9903
rect 4043 9899 4044 9903
rect 4048 9899 4049 9903
rect 4053 9899 4054 9903
rect 4058 9899 4059 9903
rect 4063 9899 4064 9903
rect 4068 9899 4069 9903
rect 4028 9898 4073 9899
rect 4028 9894 4029 9898
rect 4033 9894 4034 9898
rect 4038 9894 4039 9898
rect 4043 9894 4044 9898
rect 4048 9894 4049 9898
rect 4053 9894 4054 9898
rect 4058 9894 4059 9898
rect 4063 9894 4064 9898
rect 4068 9894 4069 9898
rect 4028 9893 4073 9894
rect 4028 9889 4029 9893
rect 4033 9889 4034 9893
rect 4038 9889 4039 9893
rect 4043 9889 4044 9893
rect 4048 9889 4049 9893
rect 4053 9889 4054 9893
rect 4058 9889 4059 9893
rect 4063 9889 4064 9893
rect 4068 9889 4069 9893
rect 4028 9888 4073 9889
rect 4028 9884 4029 9888
rect 4033 9884 4034 9888
rect 4038 9884 4039 9888
rect 4043 9884 4044 9888
rect 4048 9884 4049 9888
rect 4053 9884 4054 9888
rect 4058 9884 4059 9888
rect 4063 9884 4064 9888
rect 4068 9884 4069 9888
rect 4028 9883 4073 9884
rect 4028 9879 4029 9883
rect 4033 9879 4034 9883
rect 4038 9879 4039 9883
rect 4043 9879 4044 9883
rect 4048 9879 4049 9883
rect 4053 9879 4054 9883
rect 4058 9879 4059 9883
rect 4063 9879 4064 9883
rect 4068 9879 4069 9883
rect 4028 9878 4073 9879
rect 4028 9874 4029 9878
rect 4033 9874 4034 9878
rect 4038 9874 4039 9878
rect 4043 9874 4044 9878
rect 4048 9874 4049 9878
rect 4053 9874 4054 9878
rect 4058 9874 4059 9878
rect 4063 9874 4064 9878
rect 4068 9874 4069 9878
rect 4028 9873 4073 9874
rect 4028 9869 4029 9873
rect 4033 9869 4034 9873
rect 4038 9869 4039 9873
rect 4043 9869 4044 9873
rect 4048 9869 4049 9873
rect 4053 9869 4054 9873
rect 4058 9869 4059 9873
rect 4063 9869 4064 9873
rect 4068 9869 4069 9873
rect 4028 9868 4073 9869
rect 4028 9864 4029 9868
rect 4033 9864 4034 9868
rect 4038 9864 4039 9868
rect 4043 9864 4044 9868
rect 4048 9864 4049 9868
rect 4053 9864 4054 9868
rect 4058 9864 4059 9868
rect 4063 9864 4064 9868
rect 4068 9864 4069 9868
rect 4081 9948 4085 9949
rect 4081 9943 4085 9944
rect 4081 9938 4085 9939
rect 4081 9933 4085 9934
rect 4081 9928 4085 9929
rect 4081 9923 4085 9924
rect 4081 9918 4085 9919
rect 4081 9913 4085 9914
rect 4081 9908 4085 9909
rect 4081 9903 4085 9904
rect 4081 9898 4085 9899
rect 4081 9893 4085 9894
rect 4081 9888 4085 9889
rect 4081 9883 4085 9884
rect 4081 9878 4085 9879
rect 4081 9873 4085 9874
rect 4081 9868 4085 9869
rect 4017 9863 4021 9864
rect 4017 9856 4021 9859
rect 4081 9863 4085 9864
rect 4081 9856 4085 9859
rect 4021 9848 4024 9856
rect 4028 9848 4029 9856
rect 4033 9848 4034 9856
rect 4038 9848 4039 9856
rect 4043 9848 4044 9856
rect 4048 9848 4049 9856
rect 4053 9848 4054 9856
rect 4058 9848 4059 9856
rect 4063 9848 4064 9856
rect 4068 9848 4069 9856
rect 4073 9848 4074 9856
rect 4078 9848 4081 9856
rect 4094 9963 4098 9964
rect 4094 9958 4098 9959
rect 4094 9953 4098 9954
rect 4094 9948 4098 9949
rect 4094 9943 4098 9944
rect 4094 9938 4098 9939
rect 4094 9933 4098 9934
rect 4094 9928 4098 9929
rect 4094 9923 4098 9924
rect 4094 9918 4098 9919
rect 4094 9913 4098 9914
rect 4094 9908 4098 9909
rect 4094 9903 4098 9904
rect 4094 9898 4098 9899
rect 4094 9893 4098 9894
rect 4094 9888 4098 9889
rect 4094 9883 4098 9884
rect 4094 9878 4098 9879
rect 4094 9873 4098 9874
rect 4094 9868 4098 9869
rect 4094 9863 4098 9864
rect 4094 9858 4098 9859
rect 4094 9853 4098 9854
rect 4094 9848 4098 9849
rect 3962 9844 3979 9846
rect 3934 9843 3938 9844
rect 3848 9839 3849 9843
rect 3853 9839 3854 9843
rect 3858 9839 3859 9843
rect 3863 9839 3864 9843
rect 3868 9839 3869 9843
rect 3873 9839 3874 9843
rect 3878 9839 3879 9843
rect 3883 9839 3884 9843
rect 3888 9839 3889 9843
rect 3893 9839 3894 9843
rect 3898 9839 3899 9843
rect 3903 9839 3904 9843
rect 3908 9839 3909 9843
rect 3913 9839 3914 9843
rect 3918 9839 3919 9843
rect 3923 9839 3924 9843
rect 3928 9839 3929 9843
rect 3933 9839 3934 9843
rect 3964 9842 3977 9844
rect 4004 9843 4008 9844
rect 4094 9843 4098 9844
rect 3634 9791 3662 9795
rect 3666 9791 3667 9795
rect 3671 9791 3688 9795
rect 3634 9790 3688 9791
rect 3634 9786 3662 9790
rect 3666 9786 3667 9790
rect 3671 9786 3688 9790
rect 3634 9785 3688 9786
rect 3634 9781 3662 9785
rect 3666 9781 3667 9785
rect 3671 9781 3688 9785
rect 3634 9780 3688 9781
rect 3634 9776 3662 9780
rect 3666 9776 3667 9780
rect 3671 9776 3688 9780
rect 3634 9775 3688 9776
rect 3634 9771 3662 9775
rect 3666 9771 3667 9775
rect 3671 9771 3688 9775
rect 3634 9770 3688 9771
rect 3634 9766 3662 9770
rect 3666 9766 3667 9770
rect 3671 9766 3688 9770
rect 3634 9765 3688 9766
rect 3634 9761 3662 9765
rect 3666 9761 3667 9765
rect 3671 9761 3688 9765
rect 3634 9760 3688 9761
rect 3634 9756 3662 9760
rect 3666 9756 3667 9760
rect 3671 9756 3688 9760
rect 3634 9755 3688 9756
rect 3634 9751 3662 9755
rect 3666 9751 3667 9755
rect 3671 9751 3688 9755
rect 3634 9750 3688 9751
rect 3634 9746 3662 9750
rect 3666 9746 3667 9750
rect 3671 9746 3688 9750
rect 3634 9745 3688 9746
rect 3634 9741 3662 9745
rect 3666 9741 3667 9745
rect 3671 9741 3688 9745
rect 3427 9718 3428 9722
rect 3432 9718 3433 9722
rect 3437 9718 3438 9722
rect 3442 9718 3443 9722
rect 3447 9718 3448 9722
rect 3452 9718 3453 9722
rect 3457 9718 3458 9722
rect 3462 9718 3463 9722
rect 3467 9718 3468 9722
rect 3472 9718 3473 9722
rect 3477 9718 3479 9722
rect 3423 9717 3479 9718
rect 3427 9713 3428 9717
rect 3432 9713 3433 9717
rect 3437 9713 3438 9717
rect 3442 9713 3443 9717
rect 3447 9713 3448 9717
rect 3452 9713 3453 9717
rect 3457 9713 3458 9717
rect 3462 9713 3463 9717
rect 3467 9713 3468 9717
rect 3472 9713 3473 9717
rect 3477 9713 3479 9717
rect 3423 9712 3479 9713
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3482 9715 3501 9716
rect 3327 9710 3379 9711
rect 3327 9706 3353 9710
rect 3357 9706 3358 9710
rect 3362 9706 3379 9710
rect 3327 9705 3379 9706
rect 3327 9701 3353 9705
rect 3357 9701 3358 9705
rect 3362 9701 3379 9705
rect 3327 9700 3379 9701
rect 3327 9696 3353 9700
rect 3357 9696 3358 9700
rect 3362 9696 3379 9700
rect 3327 9695 3379 9696
rect 3327 9691 3353 9695
rect 3357 9691 3358 9695
rect 3362 9691 3379 9695
rect 3327 9690 3379 9691
rect 3327 9686 3353 9690
rect 3357 9686 3358 9690
rect 3362 9686 3379 9690
rect 3486 9711 3487 9715
rect 3491 9711 3492 9715
rect 3496 9711 3497 9715
rect 3482 9710 3501 9711
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3482 9705 3501 9706
rect 3486 9701 3487 9705
rect 3491 9701 3492 9705
rect 3496 9701 3497 9705
rect 3482 9700 3501 9701
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3482 9695 3501 9696
rect 3486 9691 3487 9695
rect 3491 9691 3492 9695
rect 3496 9691 3497 9695
rect 3482 9690 3501 9691
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 2731 9605 3021 9609
rect 3327 9685 3379 9686
rect 3327 9681 3353 9685
rect 3357 9681 3358 9685
rect 3362 9681 3379 9685
rect 3327 9680 3379 9681
rect 3327 9676 3353 9680
rect 3357 9676 3358 9680
rect 3362 9676 3379 9680
rect 3327 9675 3379 9676
rect 3327 9671 3353 9675
rect 3357 9671 3358 9675
rect 3362 9671 3379 9675
rect 3327 9670 3379 9671
rect 3327 9666 3353 9670
rect 3357 9666 3358 9670
rect 3362 9666 3379 9670
rect 3327 9665 3379 9666
rect 3327 9661 3353 9665
rect 3357 9661 3358 9665
rect 3362 9661 3379 9665
rect 3327 9610 3379 9661
rect 3634 9629 3688 9741
rect 3732 9722 3788 9839
rect 3847 9831 3903 9839
rect 3966 9831 3975 9842
rect 4008 9839 4009 9843
rect 4013 9839 4014 9843
rect 4018 9839 4019 9843
rect 4023 9839 4024 9843
rect 4028 9839 4029 9843
rect 4033 9839 4034 9843
rect 4038 9839 4039 9843
rect 4043 9839 4044 9843
rect 4048 9839 4049 9843
rect 4053 9839 4054 9843
rect 4058 9839 4059 9843
rect 4063 9839 4064 9843
rect 4068 9839 4069 9843
rect 4073 9839 4074 9843
rect 4078 9839 4079 9843
rect 4083 9839 4084 9843
rect 4088 9839 4089 9843
rect 4093 9839 4094 9843
rect 4041 9831 4097 9839
rect 3847 9827 3906 9831
rect 4032 9827 4097 9831
rect 3847 9815 3903 9827
rect 3962 9819 3992 9823
rect 3847 9811 3906 9815
rect 3976 9812 3980 9819
rect 4041 9815 4097 9827
rect 3847 9802 3903 9811
rect 4032 9811 4097 9815
rect 3962 9803 3973 9807
rect 3835 9800 3903 9802
rect 3835 9796 3836 9800
rect 3840 9796 3841 9800
rect 3845 9799 3903 9800
rect 3966 9800 3973 9803
rect 3985 9803 3992 9807
rect 3985 9800 3989 9803
rect 3845 9796 3906 9799
rect 3835 9795 3906 9796
rect 3835 9791 3836 9795
rect 3840 9791 3841 9795
rect 3845 9791 3903 9795
rect 3966 9791 3989 9800
rect 4041 9799 4097 9811
rect 4032 9795 4097 9799
rect 3835 9790 3903 9791
rect 3835 9786 3836 9790
rect 3840 9786 3841 9790
rect 3845 9786 3903 9790
rect 3962 9787 3992 9791
rect 3835 9785 3903 9786
rect 3835 9781 3836 9785
rect 3840 9781 3841 9785
rect 3845 9783 3903 9785
rect 3845 9781 3906 9783
rect 3835 9780 3906 9781
rect 3835 9776 3836 9780
rect 3840 9776 3841 9780
rect 3845 9779 3906 9780
rect 3845 9776 3903 9779
rect 3835 9775 3903 9776
rect 3835 9771 3836 9775
rect 3840 9771 3841 9775
rect 3845 9771 3903 9775
rect 3835 9770 3903 9771
rect 3835 9766 3836 9770
rect 3840 9766 3841 9770
rect 3845 9766 3903 9770
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3791 9761 3810 9762
rect 3795 9757 3796 9761
rect 3800 9757 3801 9761
rect 3805 9757 3806 9761
rect 3791 9756 3810 9757
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3791 9751 3810 9752
rect 3795 9747 3796 9751
rect 3800 9747 3801 9751
rect 3805 9747 3806 9751
rect 3791 9746 3810 9747
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3791 9741 3810 9742
rect 3795 9737 3796 9741
rect 3800 9737 3801 9741
rect 3805 9737 3806 9741
rect 3791 9736 3810 9737
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3835 9765 3903 9766
rect 3835 9761 3836 9765
rect 3840 9761 3841 9765
rect 3845 9761 3903 9765
rect 3835 9760 3903 9761
rect 3835 9756 3836 9760
rect 3840 9756 3841 9760
rect 3845 9756 3903 9760
rect 3835 9755 3903 9756
rect 3835 9751 3836 9755
rect 3840 9751 3841 9755
rect 3845 9751 3903 9755
rect 3835 9750 3903 9751
rect 3835 9746 3836 9750
rect 3840 9746 3841 9750
rect 3845 9746 3903 9750
rect 3835 9745 3903 9746
rect 3835 9741 3836 9745
rect 3840 9741 3841 9745
rect 3845 9741 3903 9745
rect 3835 9740 3903 9741
rect 3835 9736 3836 9740
rect 3840 9736 3841 9740
rect 3845 9736 3903 9740
rect 3835 9734 3903 9736
rect 3736 9718 3737 9722
rect 3741 9718 3742 9722
rect 3746 9718 3747 9722
rect 3751 9718 3752 9722
rect 3756 9718 3757 9722
rect 3761 9718 3762 9722
rect 3766 9718 3767 9722
rect 3771 9718 3772 9722
rect 3776 9718 3777 9722
rect 3781 9718 3782 9722
rect 3786 9718 3788 9722
rect 3732 9717 3788 9718
rect 3736 9713 3737 9717
rect 3741 9713 3742 9717
rect 3746 9713 3747 9717
rect 3751 9713 3752 9717
rect 3756 9713 3757 9717
rect 3761 9713 3762 9717
rect 3766 9713 3767 9717
rect 3771 9713 3772 9717
rect 3776 9713 3777 9717
rect 3781 9713 3782 9717
rect 3786 9713 3788 9717
rect 3732 9712 3788 9713
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3791 9715 3810 9716
rect 3795 9711 3796 9715
rect 3800 9711 3801 9715
rect 3805 9711 3806 9715
rect 3791 9710 3810 9711
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3791 9705 3810 9706
rect 3795 9701 3796 9705
rect 3800 9701 3801 9705
rect 3805 9701 3806 9705
rect 3791 9700 3810 9701
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3791 9695 3810 9696
rect 3795 9691 3796 9695
rect 3800 9691 3801 9695
rect 3805 9691 3806 9695
rect 3791 9690 3810 9691
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 3634 9609 3690 9629
rect 2731 9604 2997 9605
rect 659 9591 693 9592
rect 663 9587 664 9591
rect 668 9587 669 9591
rect 673 9587 674 9591
rect 678 9587 679 9591
rect 683 9587 684 9591
rect 688 9587 689 9591
rect 659 9586 693 9587
rect 663 9582 664 9586
rect 668 9582 669 9586
rect 673 9582 674 9586
rect 678 9582 679 9586
rect 683 9582 684 9586
rect 688 9582 689 9586
rect 659 9581 693 9582
rect 663 9577 664 9581
rect 668 9577 669 9581
rect 673 9577 674 9581
rect 678 9577 679 9581
rect 683 9577 684 9581
rect 688 9577 689 9581
rect 2435 9575 2497 9597
rect 3967 9574 3980 9787
rect 4041 9783 4097 9795
rect 4141 9786 5073 10261
rect 4032 9779 4097 9783
rect 4041 9722 4097 9779
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4100 9761 4119 9762
rect 4104 9757 4105 9761
rect 4109 9757 4110 9761
rect 4114 9757 4115 9761
rect 4100 9756 4119 9757
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4100 9751 4119 9752
rect 4104 9747 4105 9751
rect 4109 9747 4110 9751
rect 4114 9747 4115 9751
rect 4100 9746 4119 9747
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4100 9741 4119 9742
rect 4104 9737 4105 9741
rect 4109 9737 4110 9741
rect 4114 9737 4115 9741
rect 4100 9736 4119 9737
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4292 9761 4311 9762
rect 4296 9757 4297 9761
rect 4301 9757 4302 9761
rect 4306 9757 4307 9761
rect 4292 9756 4311 9757
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4292 9751 4311 9752
rect 4296 9747 4297 9751
rect 4301 9747 4302 9751
rect 4306 9747 4307 9751
rect 4292 9746 4311 9747
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4292 9741 4311 9742
rect 4296 9737 4297 9741
rect 4301 9737 4302 9741
rect 4306 9737 4307 9741
rect 4292 9736 4311 9737
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4318 9761 4337 9762
rect 4322 9757 4323 9761
rect 4327 9757 4328 9761
rect 4332 9757 4333 9761
rect 4318 9756 4337 9757
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4318 9751 4337 9752
rect 4322 9747 4323 9751
rect 4327 9747 4328 9751
rect 4332 9747 4333 9751
rect 4318 9746 4337 9747
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4318 9741 4337 9742
rect 4322 9737 4323 9741
rect 4327 9737 4328 9741
rect 4332 9737 4333 9741
rect 4318 9736 4337 9737
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4344 9761 4363 9762
rect 4348 9757 4349 9761
rect 4353 9757 4354 9761
rect 4358 9757 4359 9761
rect 4344 9756 4363 9757
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4344 9751 4363 9752
rect 4348 9747 4349 9751
rect 4353 9747 4354 9751
rect 4358 9747 4359 9751
rect 4344 9746 4363 9747
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4344 9741 4363 9742
rect 4348 9737 4349 9741
rect 4353 9737 4354 9741
rect 4358 9737 4359 9741
rect 4344 9736 4363 9737
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4370 9761 4389 9762
rect 4374 9757 4375 9761
rect 4379 9757 4380 9761
rect 4384 9757 4385 9761
rect 4370 9756 4389 9757
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4370 9751 4389 9752
rect 4374 9747 4375 9751
rect 4379 9747 4380 9751
rect 4384 9747 4385 9751
rect 4370 9746 4389 9747
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4370 9741 4389 9742
rect 4374 9737 4375 9741
rect 4379 9737 4380 9741
rect 4384 9737 4385 9741
rect 4370 9736 4389 9737
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4396 9761 4415 9762
rect 4400 9757 4401 9761
rect 4405 9757 4406 9761
rect 4410 9757 4411 9761
rect 4396 9756 4415 9757
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4396 9751 4415 9752
rect 4400 9747 4401 9751
rect 4405 9747 4406 9751
rect 4410 9747 4411 9751
rect 4396 9746 4415 9747
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4396 9741 4415 9742
rect 4400 9737 4401 9741
rect 4405 9737 4406 9741
rect 4410 9737 4411 9741
rect 4396 9736 4415 9737
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 4045 9718 4046 9722
rect 4050 9718 4051 9722
rect 4055 9718 4056 9722
rect 4060 9718 4061 9722
rect 4065 9718 4066 9722
rect 4070 9718 4071 9722
rect 4075 9718 4076 9722
rect 4080 9718 4081 9722
rect 4085 9718 4086 9722
rect 4090 9718 4091 9722
rect 4095 9718 4097 9722
rect 4041 9717 4097 9718
rect 4045 9713 4046 9717
rect 4050 9713 4051 9717
rect 4055 9713 4056 9717
rect 4060 9713 4061 9717
rect 4065 9713 4066 9717
rect 4070 9713 4071 9717
rect 4075 9713 4076 9717
rect 4080 9713 4081 9717
rect 4085 9713 4086 9717
rect 4090 9713 4091 9717
rect 4095 9713 4097 9717
rect 4041 9712 4097 9713
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4100 9715 4119 9716
rect 4104 9711 4105 9715
rect 4109 9711 4110 9715
rect 4114 9711 4115 9715
rect 4100 9710 4119 9711
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4100 9705 4119 9706
rect 4104 9701 4105 9705
rect 4109 9701 4110 9705
rect 4114 9701 4115 9705
rect 4100 9700 4119 9701
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4100 9695 4119 9696
rect 4104 9691 4105 9695
rect 4109 9691 4110 9695
rect 4114 9691 4115 9695
rect 4100 9690 4119 9691
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4292 9715 4311 9716
rect 4296 9711 4297 9715
rect 4301 9711 4302 9715
rect 4306 9711 4307 9715
rect 4292 9710 4311 9711
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4292 9705 4311 9706
rect 4296 9701 4297 9705
rect 4301 9701 4302 9705
rect 4306 9701 4307 9705
rect 4292 9700 4311 9701
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4292 9695 4311 9696
rect 4296 9691 4297 9695
rect 4301 9691 4302 9695
rect 4306 9691 4307 9695
rect 4292 9690 4311 9691
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4318 9715 4337 9716
rect 4322 9711 4323 9715
rect 4327 9711 4328 9715
rect 4332 9711 4333 9715
rect 4318 9710 4337 9711
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4318 9705 4337 9706
rect 4322 9701 4323 9705
rect 4327 9701 4328 9705
rect 4332 9701 4333 9705
rect 4318 9700 4337 9701
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4318 9695 4337 9696
rect 4322 9691 4323 9695
rect 4327 9691 4328 9695
rect 4332 9691 4333 9695
rect 4318 9690 4337 9691
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4344 9715 4363 9716
rect 4348 9711 4349 9715
rect 4353 9711 4354 9715
rect 4358 9711 4359 9715
rect 4344 9710 4363 9711
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4344 9705 4363 9706
rect 4348 9701 4349 9705
rect 4353 9701 4354 9705
rect 4358 9701 4359 9705
rect 4344 9700 4363 9701
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4344 9695 4363 9696
rect 4348 9691 4349 9695
rect 4353 9691 4354 9695
rect 4358 9691 4359 9695
rect 4344 9690 4363 9691
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4370 9715 4389 9716
rect 4374 9711 4375 9715
rect 4379 9711 4380 9715
rect 4384 9711 4385 9715
rect 4370 9710 4389 9711
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4370 9705 4389 9706
rect 4374 9701 4375 9705
rect 4379 9701 4380 9705
rect 4384 9701 4385 9705
rect 4370 9700 4389 9701
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4370 9695 4389 9696
rect 4374 9691 4375 9695
rect 4379 9691 4380 9695
rect 4384 9691 4385 9695
rect 4370 9690 4389 9691
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4396 9715 4415 9716
rect 4400 9711 4401 9715
rect 4405 9711 4406 9715
rect 4410 9711 4411 9715
rect 4396 9710 4415 9711
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4396 9705 4415 9706
rect 4400 9701 4401 9705
rect 4405 9701 4406 9705
rect 4410 9701 4411 9705
rect 4396 9700 4415 9701
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4396 9695 4415 9696
rect 4400 9691 4401 9695
rect 4405 9691 4406 9695
rect 4410 9691 4411 9695
rect 4396 9690 4415 9691
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 617 9566 618 9570
rect 622 9566 623 9570
rect 627 9566 628 9570
rect 632 9566 633 9570
rect 637 9566 638 9570
rect 642 9566 643 9570
rect 613 9565 647 9566
rect 617 9561 618 9565
rect 622 9561 623 9565
rect 627 9561 628 9565
rect 632 9561 633 9565
rect 637 9561 638 9565
rect 642 9561 643 9565
rect 613 9560 647 9561
rect 617 9556 618 9560
rect 622 9556 623 9560
rect 627 9556 628 9560
rect 632 9556 633 9560
rect 637 9556 638 9560
rect 642 9556 643 9560
rect 613 9555 647 9556
rect 617 9551 618 9555
rect 622 9551 623 9555
rect 627 9551 628 9555
rect 632 9551 633 9555
rect 637 9551 638 9555
rect 642 9551 643 9555
rect 663 9566 664 9570
rect 668 9566 669 9570
rect 673 9566 674 9570
rect 678 9566 679 9570
rect 683 9566 684 9570
rect 688 9566 689 9570
rect 659 9565 693 9566
rect 663 9561 664 9565
rect 668 9561 669 9565
rect 673 9561 674 9565
rect 678 9561 679 9565
rect 683 9561 684 9565
rect 688 9561 689 9565
rect 659 9560 693 9561
rect 663 9556 664 9560
rect 668 9556 669 9560
rect 673 9556 674 9560
rect 678 9556 679 9560
rect 683 9556 684 9560
rect 688 9556 689 9560
rect 659 9555 693 9556
rect 663 9551 664 9555
rect 668 9551 669 9555
rect 673 9551 674 9555
rect 678 9551 679 9555
rect 683 9551 684 9555
rect 688 9551 689 9555
rect 2134 9549 2401 9571
rect 2414 9549 2476 9571
rect 2134 9547 2416 9549
rect 617 9540 618 9544
rect 622 9540 623 9544
rect 627 9540 628 9544
rect 632 9540 633 9544
rect 637 9540 638 9544
rect 642 9540 643 9544
rect 613 9539 647 9540
rect 617 9535 618 9539
rect 622 9535 623 9539
rect 627 9535 628 9539
rect 632 9535 633 9539
rect 637 9535 638 9539
rect 642 9535 643 9539
rect 613 9534 647 9535
rect 617 9530 618 9534
rect 622 9530 623 9534
rect 627 9530 628 9534
rect 632 9530 633 9534
rect 637 9530 638 9534
rect 642 9530 643 9534
rect 613 9529 647 9530
rect 617 9525 618 9529
rect 622 9525 623 9529
rect 627 9525 628 9529
rect 632 9525 633 9529
rect 637 9525 638 9529
rect 642 9525 643 9529
rect 663 9540 664 9544
rect 668 9540 669 9544
rect 673 9540 674 9544
rect 678 9540 679 9544
rect 683 9540 684 9544
rect 688 9540 689 9544
rect 659 9539 693 9540
rect 663 9535 664 9539
rect 668 9535 669 9539
rect 673 9535 674 9539
rect 678 9535 679 9539
rect 683 9535 684 9539
rect 688 9535 689 9539
rect 659 9534 693 9535
rect 663 9530 664 9534
rect 668 9530 669 9534
rect 673 9530 674 9534
rect 678 9530 679 9534
rect 683 9530 684 9534
rect 688 9530 689 9534
rect 659 9529 693 9530
rect 663 9525 664 9529
rect 668 9525 669 9529
rect 673 9525 674 9529
rect 678 9525 679 9529
rect 683 9525 684 9529
rect 688 9525 689 9529
rect 617 9514 618 9518
rect 622 9514 623 9518
rect 627 9514 628 9518
rect 632 9514 633 9518
rect 637 9514 638 9518
rect 642 9514 643 9518
rect 613 9513 647 9514
rect 617 9509 618 9513
rect 622 9509 623 9513
rect 627 9509 628 9513
rect 632 9509 633 9513
rect 637 9509 638 9513
rect 642 9509 643 9513
rect 613 9508 647 9509
rect 617 9504 618 9508
rect 622 9504 623 9508
rect 627 9504 628 9508
rect 632 9504 633 9508
rect 637 9504 638 9508
rect 642 9504 643 9508
rect 613 9503 647 9504
rect 617 9499 618 9503
rect 622 9499 623 9503
rect 627 9499 628 9503
rect 632 9499 633 9503
rect 637 9499 638 9503
rect 642 9499 643 9503
rect 663 9514 664 9518
rect 668 9514 669 9518
rect 673 9514 674 9518
rect 678 9514 679 9518
rect 683 9514 684 9518
rect 688 9514 689 9518
rect 659 9513 693 9514
rect 663 9509 664 9513
rect 668 9509 669 9513
rect 673 9509 674 9513
rect 678 9509 679 9513
rect 683 9509 684 9513
rect 688 9509 689 9513
rect 659 9508 693 9509
rect 663 9504 664 9508
rect 668 9504 669 9508
rect 673 9504 674 9508
rect 678 9504 679 9508
rect 683 9504 684 9508
rect 688 9504 689 9508
rect 659 9503 693 9504
rect 663 9499 664 9503
rect 668 9499 669 9503
rect 673 9499 674 9503
rect 678 9499 679 9503
rect 683 9499 684 9503
rect 688 9499 689 9503
rect 2830 9497 3769 9501
rect 2818 9489 3757 9493
rect 2806 9482 3745 9486
rect 2794 9475 3733 9479
rect 2782 9467 3327 9471
rect 3382 9467 3721 9471
rect 3727 9467 3788 9471
rect 3692 9463 3709 9464
rect 2770 9459 3635 9463
rect 3690 9460 3709 9463
rect 3715 9460 3788 9464
rect 3690 9459 3698 9460
rect 3968 9456 3980 9574
rect 4483 9573 4484 9577
rect 4488 9573 4489 9577
rect 4493 9573 4494 9577
rect 4498 9573 4499 9577
rect 4503 9573 4504 9577
rect 4508 9573 4509 9577
rect 4479 9572 4513 9573
rect 4483 9568 4484 9572
rect 4488 9568 4489 9572
rect 4493 9568 4494 9572
rect 4498 9568 4499 9572
rect 4503 9568 4504 9572
rect 4508 9568 4509 9572
rect 4479 9567 4513 9568
rect 4483 9563 4484 9567
rect 4488 9563 4489 9567
rect 4493 9563 4494 9567
rect 4498 9563 4499 9567
rect 4503 9563 4504 9567
rect 4508 9563 4509 9567
rect 4479 9562 4513 9563
rect 4483 9558 4484 9562
rect 4488 9558 4489 9562
rect 4493 9558 4494 9562
rect 4498 9558 4499 9562
rect 4503 9558 4504 9562
rect 4508 9558 4509 9562
rect 4529 9573 4530 9577
rect 4534 9573 4535 9577
rect 4539 9573 4540 9577
rect 4544 9573 4545 9577
rect 4549 9573 4550 9577
rect 4554 9573 4555 9577
rect 4525 9572 4559 9573
rect 4529 9568 4530 9572
rect 4534 9568 4535 9572
rect 4539 9568 4540 9572
rect 4544 9568 4545 9572
rect 4549 9568 4550 9572
rect 4554 9568 4555 9572
rect 4525 9567 4559 9568
rect 4529 9563 4530 9567
rect 4534 9563 4535 9567
rect 4539 9563 4540 9567
rect 4544 9563 4545 9567
rect 4549 9563 4550 9567
rect 4554 9563 4555 9567
rect 4525 9562 4559 9563
rect 4529 9558 4530 9562
rect 4534 9558 4535 9562
rect 4539 9558 4540 9562
rect 4544 9558 4545 9562
rect 4549 9558 4550 9562
rect 4554 9558 4555 9562
rect 4483 9544 4484 9548
rect 4488 9544 4489 9548
rect 4493 9544 4494 9548
rect 4498 9544 4499 9548
rect 4503 9544 4504 9548
rect 4508 9544 4509 9548
rect 4479 9543 4513 9544
rect 4483 9539 4484 9543
rect 4488 9539 4489 9543
rect 4493 9539 4494 9543
rect 4498 9539 4499 9543
rect 4503 9539 4504 9543
rect 4508 9539 4509 9543
rect 4479 9538 4513 9539
rect 4483 9534 4484 9538
rect 4488 9534 4489 9538
rect 4493 9534 4494 9538
rect 4498 9534 4499 9538
rect 4503 9534 4504 9538
rect 4508 9534 4509 9538
rect 4479 9533 4513 9534
rect 4483 9529 4484 9533
rect 4488 9529 4489 9533
rect 4493 9529 4494 9533
rect 4498 9529 4499 9533
rect 4503 9529 4504 9533
rect 4508 9529 4509 9533
rect 4529 9544 4530 9548
rect 4534 9544 4535 9548
rect 4539 9544 4540 9548
rect 4544 9544 4545 9548
rect 4549 9544 4550 9548
rect 4554 9544 4555 9548
rect 4525 9543 4559 9544
rect 4529 9539 4530 9543
rect 4534 9539 4535 9543
rect 4539 9539 4540 9543
rect 4544 9539 4545 9543
rect 4549 9539 4550 9543
rect 4554 9539 4555 9543
rect 4525 9538 4559 9539
rect 4529 9534 4530 9538
rect 4534 9534 4535 9538
rect 4539 9534 4540 9538
rect 4544 9534 4545 9538
rect 4549 9534 4550 9538
rect 4554 9534 4555 9538
rect 4525 9533 4559 9534
rect 4529 9529 4530 9533
rect 4534 9529 4535 9533
rect 4539 9529 4540 9533
rect 4544 9529 4545 9533
rect 4549 9529 4550 9533
rect 4554 9529 4555 9533
rect 4483 9515 4484 9519
rect 4488 9515 4489 9519
rect 4493 9515 4494 9519
rect 4498 9515 4499 9519
rect 4503 9515 4504 9519
rect 4508 9515 4509 9519
rect 4479 9514 4513 9515
rect 4483 9510 4484 9514
rect 4488 9510 4489 9514
rect 4493 9510 4494 9514
rect 4498 9510 4499 9514
rect 4503 9510 4504 9514
rect 4508 9510 4509 9514
rect 4479 9509 4513 9510
rect 4483 9505 4484 9509
rect 4488 9505 4489 9509
rect 4493 9505 4494 9509
rect 4498 9505 4499 9509
rect 4503 9505 4504 9509
rect 4508 9505 4509 9509
rect 4479 9504 4513 9505
rect 4483 9500 4484 9504
rect 4488 9500 4489 9504
rect 4493 9500 4494 9504
rect 4498 9500 4499 9504
rect 4503 9500 4504 9504
rect 4508 9500 4509 9504
rect 4529 9515 4530 9519
rect 4534 9515 4535 9519
rect 4539 9515 4540 9519
rect 4544 9515 4545 9519
rect 4549 9515 4550 9519
rect 4554 9515 4555 9519
rect 4525 9514 4559 9515
rect 4529 9510 4530 9514
rect 4534 9510 4535 9514
rect 4539 9510 4540 9514
rect 4544 9510 4545 9514
rect 4549 9510 4550 9514
rect 4554 9510 4555 9514
rect 4525 9509 4559 9510
rect 4529 9505 4530 9509
rect 4534 9505 4535 9509
rect 4539 9505 4540 9509
rect 4544 9505 4545 9509
rect 4549 9505 4550 9509
rect 4554 9505 4555 9509
rect 4525 9504 4559 9505
rect 4529 9500 4530 9504
rect 4534 9500 4535 9504
rect 4539 9500 4540 9504
rect 4544 9500 4545 9504
rect 4549 9500 4550 9504
rect 4554 9500 4555 9504
rect 4483 9486 4484 9490
rect 4488 9486 4489 9490
rect 4493 9486 4494 9490
rect 4498 9486 4499 9490
rect 4503 9486 4504 9490
rect 4508 9486 4509 9490
rect 4479 9485 4513 9486
rect 4483 9481 4484 9485
rect 4488 9481 4489 9485
rect 4493 9481 4494 9485
rect 4498 9481 4499 9485
rect 4503 9481 4504 9485
rect 4508 9481 4509 9485
rect 4479 9480 4513 9481
rect 4483 9476 4484 9480
rect 4488 9476 4489 9480
rect 4493 9476 4494 9480
rect 4498 9476 4499 9480
rect 4503 9476 4504 9480
rect 4508 9476 4509 9480
rect 4479 9475 4513 9476
rect 4483 9471 4484 9475
rect 4488 9471 4489 9475
rect 4493 9471 4494 9475
rect 4498 9471 4499 9475
rect 4503 9471 4504 9475
rect 4508 9471 4509 9475
rect 4529 9486 4530 9490
rect 4534 9486 4535 9490
rect 4539 9486 4540 9490
rect 4544 9486 4545 9490
rect 4549 9486 4550 9490
rect 4554 9486 4555 9490
rect 4525 9485 4559 9486
rect 4529 9481 4530 9485
rect 4534 9481 4535 9485
rect 4539 9481 4540 9485
rect 4544 9481 4545 9485
rect 4549 9481 4550 9485
rect 4554 9481 4555 9485
rect 4525 9480 4559 9481
rect 4529 9476 4530 9480
rect 4534 9476 4535 9480
rect 4539 9476 4540 9480
rect 4544 9476 4545 9480
rect 4549 9476 4550 9480
rect 4554 9476 4555 9480
rect 4525 9475 4559 9476
rect 4529 9471 4530 9475
rect 4534 9471 4535 9475
rect 4539 9471 4540 9475
rect 4544 9471 4545 9475
rect 4549 9471 4550 9475
rect 4554 9471 4555 9475
rect 2842 9452 3781 9456
rect 3787 9452 3980 9456
rect 4483 9457 4484 9461
rect 4488 9457 4489 9461
rect 4493 9457 4494 9461
rect 4498 9457 4499 9461
rect 4503 9457 4504 9461
rect 4508 9457 4509 9461
rect 4479 9456 4513 9457
rect 4483 9452 4484 9456
rect 4488 9452 4489 9456
rect 4493 9452 4494 9456
rect 4498 9452 4499 9456
rect 4503 9452 4504 9456
rect 4508 9452 4509 9456
rect 4479 9451 4513 9452
rect 3053 9444 3423 9448
rect 4483 9447 4484 9451
rect 4488 9447 4489 9451
rect 4493 9447 4494 9451
rect 4498 9447 4499 9451
rect 4503 9447 4504 9451
rect 4508 9447 4509 9451
rect 4479 9446 4513 9447
rect 4483 9442 4484 9446
rect 4488 9442 4489 9446
rect 4493 9442 4494 9446
rect 4498 9442 4499 9446
rect 4503 9442 4504 9446
rect 4508 9442 4509 9446
rect 4529 9457 4530 9461
rect 4534 9457 4535 9461
rect 4539 9457 4540 9461
rect 4544 9457 4545 9461
rect 4549 9457 4550 9461
rect 4554 9457 4555 9461
rect 4525 9456 4559 9457
rect 4529 9452 4530 9456
rect 4534 9452 4535 9456
rect 4539 9452 4540 9456
rect 4544 9452 4545 9456
rect 4549 9452 4550 9456
rect 4554 9452 4555 9456
rect 4525 9451 4559 9452
rect 4529 9447 4530 9451
rect 4534 9447 4535 9451
rect 4539 9447 4540 9451
rect 4544 9447 4545 9451
rect 4549 9447 4550 9451
rect 4554 9447 4555 9451
rect 4525 9446 4559 9447
rect 4529 9442 4530 9446
rect 4534 9442 4535 9446
rect 4539 9442 4540 9446
rect 4544 9442 4545 9446
rect 4549 9442 4550 9446
rect 4554 9442 4555 9446
rect 3026 9434 3411 9438
rect 4579 9355 5073 9786
rect 2830 9347 2857 9351
rect 2861 9347 2893 9351
rect 2897 9347 2960 9351
rect 2964 9347 2989 9351
rect 2993 9347 3025 9351
rect 3029 9347 3092 9351
rect 3096 9347 3121 9351
rect 3125 9347 3157 9351
rect 3161 9347 3224 9351
rect 3228 9347 3253 9351
rect 3257 9347 3289 9351
rect 3293 9347 3356 9351
rect 3360 9347 3376 9351
rect 3775 9347 3802 9351
rect 3806 9347 3838 9351
rect 3842 9347 3905 9351
rect 3909 9347 3934 9351
rect 3938 9347 3970 9351
rect 3974 9347 4037 9351
rect 4041 9347 4066 9351
rect 4070 9347 4102 9351
rect 4106 9347 4169 9351
rect 4173 9347 4198 9351
rect 4202 9347 4234 9351
rect 4238 9347 4301 9351
rect 4305 9347 4321 9351
rect 2770 9340 2881 9344
rect 2885 9340 2909 9344
rect 2913 9340 2939 9344
rect 2943 9340 2976 9344
rect 2980 9340 3013 9344
rect 3017 9340 3041 9344
rect 3045 9340 3071 9344
rect 3075 9340 3108 9344
rect 3112 9340 3145 9344
rect 3149 9340 3173 9344
rect 3177 9340 3203 9344
rect 3207 9340 3240 9344
rect 3244 9340 3277 9344
rect 3281 9340 3305 9344
rect 3309 9340 3335 9344
rect 3339 9340 3372 9344
rect 3715 9340 3826 9344
rect 3830 9340 3854 9344
rect 3858 9340 3884 9344
rect 3888 9340 3921 9344
rect 3925 9340 3958 9344
rect 3962 9340 3986 9344
rect 3990 9340 4016 9344
rect 4020 9340 4053 9344
rect 4057 9340 4090 9344
rect 4094 9340 4118 9344
rect 4122 9340 4148 9344
rect 4152 9340 4185 9344
rect 4189 9340 4222 9344
rect 4226 9340 4250 9344
rect 4254 9340 4280 9344
rect 4284 9340 4317 9344
rect 2851 9330 2854 9340
rect 2872 9330 2875 9340
rect 2888 9330 2891 9340
rect 2902 9333 2907 9337
rect 2911 9333 2918 9337
rect 2930 9330 2933 9340
rect 2946 9330 2949 9340
rect 2967 9330 2970 9340
rect 2983 9330 2986 9340
rect 3004 9330 3007 9340
rect 3020 9330 3023 9340
rect 3034 9333 3039 9337
rect 3043 9333 3050 9337
rect 3062 9330 3065 9340
rect 3078 9330 3081 9340
rect 3099 9330 3102 9340
rect 3115 9330 3118 9340
rect 3136 9330 3139 9340
rect 3152 9330 3155 9340
rect 3166 9333 3171 9337
rect 3175 9333 3182 9337
rect 3194 9330 3197 9340
rect 3210 9330 3213 9340
rect 3231 9330 3234 9340
rect 3247 9330 3250 9340
rect 3268 9330 3271 9340
rect 3284 9330 3287 9340
rect 3298 9333 3303 9337
rect 3307 9333 3314 9337
rect 3326 9330 3329 9340
rect 3342 9330 3345 9340
rect 3363 9330 3366 9340
rect 3796 9330 3799 9340
rect 3817 9330 3820 9340
rect 3833 9330 3836 9340
rect 3847 9333 3852 9337
rect 3856 9333 3863 9337
rect 3875 9330 3878 9340
rect 3891 9330 3894 9340
rect 3912 9330 3915 9340
rect 3928 9330 3931 9340
rect 3949 9330 3952 9340
rect 3965 9330 3968 9340
rect 3979 9333 3984 9337
rect 3988 9333 3995 9337
rect 4007 9330 4010 9340
rect 4023 9330 4026 9340
rect 4044 9330 4047 9340
rect 4060 9330 4063 9340
rect 4081 9330 4084 9340
rect 4097 9330 4100 9340
rect 4111 9333 4116 9337
rect 4120 9333 4127 9337
rect 4139 9330 4142 9340
rect 4155 9330 4158 9340
rect 4176 9330 4179 9340
rect 4192 9330 4195 9340
rect 4213 9330 4216 9340
rect 4229 9330 4232 9340
rect 4243 9333 4248 9337
rect 4252 9333 4259 9337
rect 4271 9330 4274 9340
rect 4287 9330 4290 9340
rect 4308 9330 4311 9340
rect 617 9321 618 9325
rect 622 9321 623 9325
rect 627 9321 628 9325
rect 632 9321 633 9325
rect 637 9321 638 9325
rect 642 9321 643 9325
rect 613 9320 647 9321
rect 617 9316 618 9320
rect 622 9316 623 9320
rect 627 9316 628 9320
rect 632 9316 633 9320
rect 637 9316 638 9320
rect 642 9316 643 9320
rect 613 9315 647 9316
rect 617 9311 618 9315
rect 622 9311 623 9315
rect 627 9311 628 9315
rect 632 9311 633 9315
rect 637 9311 638 9315
rect 642 9311 643 9315
rect 613 9310 647 9311
rect 86 9304 346 9307
rect 617 9306 618 9310
rect 622 9306 623 9310
rect 627 9306 628 9310
rect 632 9306 633 9310
rect 637 9306 638 9310
rect 642 9306 643 9310
rect 663 9321 664 9325
rect 668 9321 669 9325
rect 673 9321 674 9325
rect 678 9321 679 9325
rect 683 9321 684 9325
rect 688 9321 689 9325
rect 659 9320 693 9321
rect 663 9316 664 9320
rect 668 9316 669 9320
rect 673 9316 674 9320
rect 678 9316 679 9320
rect 683 9316 684 9320
rect 688 9316 689 9320
rect 659 9315 693 9316
rect 663 9311 664 9315
rect 668 9311 669 9315
rect 673 9311 674 9315
rect 678 9311 679 9315
rect 683 9311 684 9315
rect 688 9311 689 9315
rect 2496 9314 2505 9318
rect 2509 9314 2541 9318
rect 2545 9314 2608 9318
rect 2612 9314 2824 9318
rect 2868 9316 2873 9319
rect 2877 9316 2901 9319
rect 2926 9316 2933 9319
rect 2937 9316 2959 9319
rect 659 9310 693 9311
rect 663 9306 664 9310
rect 668 9306 669 9310
rect 673 9306 674 9310
rect 678 9306 679 9310
rect 683 9306 684 9310
rect 688 9306 689 9310
rect 2496 9307 2529 9311
rect 2533 9307 2557 9311
rect 2561 9307 2587 9311
rect 2591 9307 2624 9311
rect 2628 9307 2764 9311
rect 86 9050 89 9304
rect 343 9265 346 9304
rect 2499 9297 2502 9307
rect 2520 9297 2523 9307
rect 2536 9297 2539 9307
rect 2550 9300 2555 9304
rect 2559 9300 2566 9304
rect 2578 9297 2581 9307
rect 2594 9297 2597 9307
rect 2615 9297 2618 9307
rect 2884 9306 2891 9309
rect 2895 9310 2914 9313
rect 2914 9303 2917 9309
rect 2942 9306 2949 9309
rect 2953 9310 2970 9313
rect 3000 9316 3005 9319
rect 3009 9316 3033 9319
rect 3058 9316 3065 9319
rect 3069 9316 3091 9319
rect 3016 9306 3023 9309
rect 3027 9310 3046 9313
rect 3046 9303 3049 9309
rect 3074 9306 3081 9309
rect 3085 9310 3102 9313
rect 3132 9316 3137 9319
rect 3141 9316 3165 9319
rect 3190 9316 3197 9319
rect 3201 9316 3223 9319
rect 3148 9306 3155 9309
rect 3159 9310 3178 9313
rect 3178 9303 3181 9309
rect 3206 9306 3213 9309
rect 3217 9310 3234 9313
rect 3264 9316 3269 9319
rect 3273 9316 3297 9319
rect 3322 9316 3329 9319
rect 3333 9316 3355 9319
rect 3441 9314 3450 9318
rect 3454 9314 3486 9318
rect 3490 9314 3553 9318
rect 3557 9314 3769 9318
rect 3280 9306 3287 9309
rect 3291 9310 3310 9313
rect 2494 9280 2503 9284
rect 2516 9283 2521 9286
rect 2525 9283 2549 9286
rect 2574 9283 2581 9286
rect 2585 9283 2607 9286
rect 2851 9287 2854 9299
rect 2872 9287 2875 9299
rect 2888 9287 2891 9299
rect 2902 9290 2914 9293
rect 2930 9287 2933 9299
rect 2946 9287 2949 9299
rect 2967 9287 2970 9299
rect 2983 9287 2986 9299
rect 3004 9287 3007 9299
rect 3020 9287 3023 9299
rect 3034 9290 3046 9293
rect 3062 9287 3065 9299
rect 3078 9287 3081 9299
rect 3099 9287 3102 9299
rect 3115 9287 3118 9299
rect 3136 9287 3139 9299
rect 3152 9287 3155 9299
rect 3166 9290 3178 9293
rect 3194 9287 3197 9299
rect 3210 9287 3213 9299
rect 3231 9287 3234 9299
rect 3310 9303 3313 9309
rect 3338 9306 3345 9309
rect 3349 9310 3366 9313
rect 3813 9316 3818 9319
rect 3822 9316 3846 9319
rect 3871 9316 3878 9319
rect 3882 9316 3904 9319
rect 3441 9307 3474 9311
rect 3478 9307 3502 9311
rect 3506 9307 3532 9311
rect 3536 9307 3569 9311
rect 3573 9307 3709 9311
rect 3247 9287 3250 9299
rect 3268 9287 3271 9299
rect 3284 9287 3287 9299
rect 3298 9290 3310 9293
rect 3326 9287 3329 9299
rect 3342 9287 3345 9299
rect 3363 9287 3366 9299
rect 3444 9297 3447 9307
rect 3465 9297 3468 9307
rect 3481 9297 3484 9307
rect 3495 9300 3500 9304
rect 3504 9300 3511 9304
rect 3523 9297 3526 9307
rect 3539 9297 3542 9307
rect 3560 9297 3563 9307
rect 3829 9306 3836 9309
rect 3840 9310 3859 9313
rect 3859 9303 3862 9309
rect 3887 9306 3894 9309
rect 3898 9310 3915 9313
rect 3945 9316 3950 9319
rect 3954 9316 3978 9319
rect 4003 9316 4010 9319
rect 4014 9316 4036 9319
rect 3961 9306 3968 9309
rect 3972 9310 3991 9313
rect 3991 9303 3994 9309
rect 4019 9306 4026 9309
rect 4030 9310 4047 9313
rect 4077 9316 4082 9319
rect 4086 9316 4110 9319
rect 4135 9316 4142 9319
rect 4146 9316 4168 9319
rect 4093 9306 4100 9309
rect 4104 9310 4123 9313
rect 4123 9303 4126 9309
rect 4151 9306 4158 9309
rect 4162 9310 4179 9313
rect 4209 9316 4214 9319
rect 4218 9316 4242 9319
rect 4267 9316 4274 9319
rect 4278 9316 4300 9319
rect 4826 9316 5086 9319
rect 4225 9306 4232 9309
rect 4236 9310 4255 9313
rect 2782 9283 2881 9287
rect 2885 9283 2909 9287
rect 2913 9283 2939 9287
rect 2943 9283 3013 9287
rect 3017 9283 3041 9287
rect 3045 9283 3071 9287
rect 3075 9283 3145 9287
rect 3149 9283 3173 9287
rect 3177 9283 3203 9287
rect 3207 9283 3277 9287
rect 3281 9283 3305 9287
rect 3309 9283 3335 9287
rect 3339 9283 3376 9287
rect 2532 9273 2539 9276
rect 2543 9277 2562 9280
rect 2562 9270 2565 9276
rect 2590 9273 2597 9276
rect 2601 9277 2616 9280
rect 3439 9280 3448 9284
rect 3461 9283 3466 9286
rect 3470 9283 3494 9286
rect 3519 9283 3526 9286
rect 3530 9283 3552 9286
rect 3796 9287 3799 9299
rect 3817 9287 3820 9299
rect 3833 9287 3836 9299
rect 3847 9290 3859 9293
rect 3875 9287 3878 9299
rect 3891 9287 3894 9299
rect 3912 9287 3915 9299
rect 3928 9287 3931 9299
rect 3949 9287 3952 9299
rect 3965 9287 3968 9299
rect 3979 9290 3991 9293
rect 4007 9287 4010 9299
rect 4023 9287 4026 9299
rect 4044 9287 4047 9299
rect 4060 9287 4063 9299
rect 4081 9287 4084 9299
rect 4097 9287 4100 9299
rect 4111 9290 4123 9293
rect 4139 9287 4142 9299
rect 4155 9287 4158 9299
rect 4176 9287 4179 9299
rect 4255 9303 4258 9309
rect 4283 9306 4290 9309
rect 4294 9310 4311 9313
rect 4192 9287 4195 9299
rect 4213 9287 4216 9299
rect 4229 9287 4232 9299
rect 4243 9290 4255 9293
rect 4271 9287 4274 9299
rect 4287 9287 4290 9299
rect 4308 9287 4311 9299
rect 3727 9283 3826 9287
rect 3830 9283 3854 9287
rect 3858 9283 3884 9287
rect 3888 9283 3958 9287
rect 3962 9283 3986 9287
rect 3990 9283 4016 9287
rect 4020 9283 4090 9287
rect 4094 9283 4118 9287
rect 4122 9283 4148 9287
rect 4152 9283 4222 9287
rect 4226 9283 4250 9287
rect 4254 9283 4280 9287
rect 4284 9283 4321 9287
rect 2818 9276 2857 9280
rect 2861 9276 2908 9280
rect 2912 9276 2958 9280
rect 2962 9276 2989 9280
rect 2993 9276 3040 9280
rect 3044 9276 3090 9280
rect 3094 9276 3121 9280
rect 3125 9276 3172 9280
rect 3176 9276 3222 9280
rect 3226 9276 3253 9280
rect 3257 9276 3304 9280
rect 3308 9276 3354 9280
rect 3358 9276 3376 9280
rect 3477 9273 3484 9276
rect 3488 9277 3507 9280
rect 343 9255 356 9265
rect 343 9245 366 9255
rect 2499 9254 2502 9266
rect 2520 9254 2523 9266
rect 2536 9254 2539 9266
rect 2550 9257 2562 9260
rect 2578 9254 2581 9266
rect 2594 9254 2597 9266
rect 2615 9254 2618 9266
rect 2770 9263 2855 9267
rect 2859 9263 2871 9267
rect 2875 9263 2889 9267
rect 2893 9263 2900 9267
rect 2904 9263 2906 9267
rect 2910 9263 2925 9267
rect 2929 9263 2962 9267
rect 2966 9263 2967 9267
rect 2971 9263 2979 9267
rect 2983 9263 3007 9267
rect 3011 9263 3023 9267
rect 3027 9263 3047 9267
rect 3051 9263 3101 9267
rect 3105 9263 3128 9267
rect 3132 9263 3182 9267
rect 3186 9263 3205 9267
rect 3507 9270 3510 9276
rect 3535 9273 3542 9276
rect 3546 9277 3561 9280
rect 3763 9276 3802 9280
rect 3806 9276 3853 9280
rect 3857 9276 3903 9280
rect 3907 9276 3934 9280
rect 3938 9276 3985 9280
rect 3989 9276 4035 9280
rect 4039 9276 4066 9280
rect 4070 9276 4117 9280
rect 4121 9276 4167 9280
rect 4171 9276 4198 9280
rect 4202 9276 4249 9280
rect 4253 9276 4299 9280
rect 4303 9276 4321 9280
rect 4826 9277 4829 9316
rect 4816 9267 4829 9277
rect 2806 9256 2882 9260
rect 2886 9256 2913 9260
rect 2917 9256 2935 9260
rect 2939 9256 3000 9260
rect 3004 9256 3018 9260
rect 3030 9259 3033 9263
rect 2496 9250 2529 9254
rect 2533 9250 2557 9254
rect 2561 9250 2587 9254
rect 2591 9250 2776 9254
rect 343 9235 376 9245
rect 2496 9243 2505 9247
rect 2509 9243 2556 9247
rect 2560 9243 2606 9247
rect 2610 9243 2812 9247
rect 2925 9249 2928 9253
rect 2952 9249 2953 9253
rect 2997 9249 2999 9253
rect 3039 9246 3042 9251
rect 3054 9253 3057 9263
rect 3084 9259 3087 9263
rect 3111 9259 3114 9263
rect 343 9225 386 9235
rect 2494 9227 2510 9231
rect 2619 9229 2623 9233
rect 2635 9229 2639 9233
rect 2643 9229 2857 9233
rect 2865 9232 2868 9238
rect 2872 9232 2875 9238
rect 2865 9229 2875 9232
rect 343 9129 769 9225
rect 2865 9224 2868 9229
rect 2502 9220 2506 9224
rect 2518 9220 2639 9224
rect 2872 9224 2875 9229
rect 2881 9234 2884 9238
rect 2881 9230 2883 9234
rect 2887 9230 2889 9234
rect 2897 9233 2900 9238
rect 2925 9235 2928 9238
rect 2897 9231 2908 9233
rect 2881 9224 2884 9230
rect 2897 9229 2903 9231
rect 2897 9224 2900 9229
rect 2907 9229 2908 9231
rect 2926 9231 2928 9235
rect 2925 9224 2928 9231
rect 3028 9242 3031 9245
rect 3070 9242 3073 9245
rect 2941 9234 2944 9238
rect 2951 9234 2954 9238
rect 2951 9230 2960 9234
rect 2972 9233 2975 9238
rect 2997 9234 3000 9238
rect 2941 9224 2944 9230
rect 2951 9224 2954 9230
rect 2972 9229 2973 9233
rect 2977 9229 2980 9232
rect 2999 9230 3000 9234
rect 3015 9233 3018 9238
rect 3039 9237 3042 9242
rect 3047 9238 3058 9241
rect 3070 9239 3078 9242
rect 2972 9224 2975 9229
rect 2997 9224 3000 9230
rect 3015 9224 3018 9229
rect 2489 9212 2505 9216
rect 2509 9212 2572 9216
rect 2576 9212 2608 9216
rect 2612 9212 2824 9216
rect 2917 9211 2918 9215
rect 2942 9212 2943 9216
rect 2989 9211 2990 9215
rect 2493 9205 2526 9209
rect 2530 9205 2556 9209
rect 2560 9205 2584 9209
rect 2588 9205 2764 9209
rect 2499 9195 2502 9205
rect 2520 9195 2523 9205
rect 2536 9195 2539 9205
rect 2551 9198 2558 9202
rect 2562 9198 2567 9202
rect 2578 9195 2581 9205
rect 2594 9195 2597 9205
rect 2615 9195 2618 9205
rect 2794 9204 2870 9208
rect 2874 9204 2929 9208
rect 2933 9204 2954 9208
rect 2958 9204 2985 9208
rect 2989 9204 3018 9208
rect 3030 9201 3033 9233
rect 3047 9232 3050 9238
rect 3070 9233 3073 9239
rect 3082 9234 3085 9237
rect 3093 9237 3096 9251
rect 3120 9246 3123 9251
rect 3135 9253 3138 9263
rect 3165 9259 3168 9263
rect 3104 9242 3105 9245
rect 3109 9242 3112 9245
rect 3151 9242 3154 9245
rect 3093 9234 3101 9237
rect 3120 9237 3123 9242
rect 3093 9229 3096 9234
rect 3101 9230 3105 9234
rect 3128 9238 3139 9241
rect 3151 9239 3159 9242
rect 3045 9223 3050 9228
rect 3054 9201 3057 9229
rect 3084 9201 3087 9225
rect 3111 9201 3114 9233
rect 3128 9232 3131 9238
rect 3151 9233 3154 9239
rect 3163 9234 3166 9237
rect 3174 9237 3177 9251
rect 3328 9250 3411 9258
rect 3444 9254 3447 9266
rect 3465 9254 3468 9266
rect 3481 9254 3484 9266
rect 3495 9257 3507 9260
rect 3523 9254 3526 9266
rect 3539 9254 3542 9266
rect 3560 9254 3563 9266
rect 3715 9263 3800 9267
rect 3804 9263 3816 9267
rect 3820 9263 3834 9267
rect 3838 9263 3845 9267
rect 3849 9263 3851 9267
rect 3855 9263 3870 9267
rect 3874 9263 3907 9267
rect 3911 9263 3912 9267
rect 3916 9263 3924 9267
rect 3928 9263 3952 9267
rect 3956 9263 3968 9267
rect 3972 9263 3992 9267
rect 3996 9263 4046 9267
rect 4050 9263 4073 9267
rect 4077 9263 4127 9267
rect 4131 9263 4150 9267
rect 3751 9256 3827 9260
rect 3831 9256 3858 9260
rect 3862 9256 3880 9260
rect 3884 9256 3945 9260
rect 3949 9256 3963 9260
rect 3975 9259 3978 9263
rect 3441 9250 3474 9254
rect 3478 9250 3502 9254
rect 3506 9250 3532 9254
rect 3536 9250 3721 9254
rect 3365 9241 3423 9245
rect 3441 9243 3450 9247
rect 3454 9243 3501 9247
rect 3505 9243 3551 9247
rect 3555 9243 3757 9247
rect 3870 9249 3873 9253
rect 3897 9249 3898 9253
rect 3942 9249 3944 9253
rect 3984 9246 3987 9251
rect 3999 9253 4002 9263
rect 4029 9259 4032 9263
rect 4056 9259 4059 9263
rect 3174 9234 3186 9237
rect 3174 9229 3177 9234
rect 3126 9223 3131 9228
rect 3135 9201 3138 9229
rect 3439 9227 3455 9231
rect 3564 9229 3568 9233
rect 3580 9229 3584 9233
rect 3588 9229 3793 9233
rect 3797 9229 3802 9233
rect 3810 9232 3813 9238
rect 3817 9232 3820 9238
rect 3810 9229 3820 9232
rect 3165 9201 3168 9225
rect 3810 9224 3813 9229
rect 3447 9220 3451 9224
rect 3463 9220 3584 9224
rect 3817 9224 3820 9229
rect 3826 9234 3829 9238
rect 3826 9230 3828 9234
rect 3832 9230 3834 9234
rect 3842 9233 3845 9238
rect 3870 9235 3873 9238
rect 3842 9231 3853 9233
rect 3826 9224 3829 9230
rect 3842 9229 3848 9231
rect 3842 9224 3845 9229
rect 3852 9229 3853 9231
rect 3871 9231 3873 9235
rect 3870 9224 3873 9231
rect 3973 9242 3976 9245
rect 4015 9242 4018 9245
rect 3886 9234 3889 9238
rect 3896 9234 3899 9238
rect 3896 9230 3905 9234
rect 3917 9233 3920 9238
rect 3942 9234 3945 9238
rect 3886 9224 3889 9230
rect 3896 9224 3899 9230
rect 3917 9229 3918 9233
rect 3922 9229 3925 9232
rect 3944 9230 3945 9234
rect 3960 9233 3963 9238
rect 3984 9237 3987 9242
rect 3992 9238 4003 9241
rect 4015 9239 4023 9242
rect 3917 9224 3920 9229
rect 3942 9224 3945 9230
rect 3960 9224 3963 9229
rect 3434 9212 3450 9216
rect 3454 9212 3517 9216
rect 3521 9212 3553 9216
rect 3557 9212 3769 9216
rect 3862 9211 3863 9215
rect 3887 9212 3888 9216
rect 3934 9211 3935 9215
rect 3438 9205 3471 9209
rect 3475 9205 3501 9209
rect 3505 9205 3529 9209
rect 3533 9205 3709 9209
rect 2782 9197 2856 9201
rect 2860 9197 2862 9201
rect 2866 9197 2870 9201
rect 2874 9197 2888 9201
rect 2892 9197 2897 9201
rect 2901 9197 2906 9201
rect 2910 9197 2929 9201
rect 2933 9197 2963 9201
rect 2967 9197 2978 9201
rect 2982 9197 3006 9201
rect 3010 9197 3023 9201
rect 3027 9197 3047 9201
rect 3051 9197 3101 9201
rect 3108 9197 3128 9201
rect 3132 9197 3182 9201
rect 2510 9181 2532 9184
rect 2536 9181 2543 9184
rect 2794 9190 2870 9194
rect 2874 9190 2929 9194
rect 2933 9190 2954 9194
rect 2958 9190 2985 9194
rect 2989 9190 3018 9194
rect 2568 9181 2592 9184
rect 2596 9181 2601 9184
rect 2917 9183 2918 9187
rect 2942 9182 2943 9186
rect 2989 9183 2990 9187
rect 2614 9178 2623 9182
rect 2501 9175 2516 9178
rect 2555 9175 2574 9178
rect 2520 9171 2527 9174
rect 2552 9168 2555 9174
rect 2578 9171 2585 9174
rect 2865 9169 2868 9174
rect 2872 9169 2875 9174
rect 2855 9166 2857 9169
rect 2865 9166 2875 9169
rect 2499 9152 2502 9164
rect 2520 9152 2523 9164
rect 2536 9152 2539 9164
rect 2555 9155 2567 9158
rect 2578 9152 2581 9164
rect 2594 9152 2597 9164
rect 2615 9152 2618 9164
rect 2865 9160 2868 9166
rect 2872 9160 2875 9166
rect 2881 9168 2884 9174
rect 2897 9169 2900 9174
rect 2881 9164 2883 9168
rect 2887 9164 2889 9168
rect 2897 9167 2903 9169
rect 2907 9167 2908 9169
rect 2897 9165 2908 9167
rect 2925 9167 2928 9174
rect 2881 9160 2884 9164
rect 2897 9160 2900 9165
rect 2926 9163 2928 9167
rect 2925 9160 2928 9163
rect 2941 9168 2944 9174
rect 2951 9168 2954 9174
rect 2972 9169 2975 9174
rect 2951 9164 2960 9168
rect 2972 9165 2973 9169
rect 2977 9166 2980 9169
rect 2997 9168 3000 9174
rect 3015 9169 3018 9174
rect 3054 9177 3057 9197
rect 3135 9177 3138 9197
rect 3444 9195 3447 9205
rect 3465 9195 3468 9205
rect 3481 9195 3484 9205
rect 3496 9198 3503 9202
rect 3507 9198 3512 9202
rect 3523 9195 3526 9205
rect 3539 9195 3542 9205
rect 3560 9195 3563 9205
rect 3739 9204 3815 9208
rect 3819 9204 3874 9208
rect 3878 9204 3899 9208
rect 3903 9204 3930 9208
rect 3934 9204 3963 9208
rect 3975 9201 3978 9233
rect 3992 9232 3995 9238
rect 4015 9233 4018 9239
rect 4027 9234 4030 9237
rect 4038 9237 4041 9251
rect 4065 9246 4068 9251
rect 4080 9253 4083 9263
rect 4110 9259 4113 9263
rect 4049 9242 4050 9245
rect 4054 9242 4057 9245
rect 4806 9257 4829 9267
rect 4096 9242 4099 9245
rect 4038 9234 4046 9237
rect 4065 9237 4068 9242
rect 4038 9229 4041 9234
rect 4046 9230 4050 9234
rect 4073 9238 4084 9241
rect 4096 9239 4104 9242
rect 3990 9223 3995 9228
rect 3999 9201 4002 9229
rect 4029 9201 4032 9225
rect 4056 9201 4059 9233
rect 4073 9232 4076 9238
rect 4096 9233 4099 9239
rect 4108 9234 4111 9237
rect 4119 9237 4122 9251
rect 4796 9247 4829 9257
rect 4119 9234 4131 9237
rect 4786 9237 4829 9247
rect 4119 9229 4122 9234
rect 4071 9223 4076 9228
rect 4080 9201 4083 9229
rect 4110 9201 4113 9225
rect 3727 9197 3801 9201
rect 3805 9197 3807 9201
rect 3811 9197 3815 9201
rect 3819 9197 3833 9201
rect 3837 9197 3842 9201
rect 3846 9197 3851 9201
rect 3855 9197 3874 9201
rect 3878 9197 3908 9201
rect 3912 9197 3923 9201
rect 3927 9197 3951 9201
rect 3955 9197 3968 9201
rect 3972 9197 3992 9201
rect 3996 9197 4046 9201
rect 4053 9197 4073 9201
rect 4077 9197 4127 9201
rect 3455 9181 3477 9184
rect 3481 9181 3488 9184
rect 3739 9190 3815 9194
rect 3819 9190 3874 9194
rect 3878 9190 3899 9194
rect 3903 9190 3930 9194
rect 3934 9190 3963 9194
rect 3513 9181 3537 9184
rect 3541 9181 3546 9184
rect 3862 9183 3863 9187
rect 3887 9182 3888 9186
rect 3934 9183 3935 9187
rect 3559 9178 3568 9182
rect 3446 9175 3461 9178
rect 2941 9160 2944 9164
rect 2951 9160 2954 9164
rect 2972 9160 2975 9165
rect 2999 9164 3000 9168
rect 2997 9160 3000 9164
rect 3015 9160 3018 9165
rect 3045 9164 3050 9169
rect 3054 9165 3055 9168
rect 3070 9167 3073 9173
rect 3070 9164 3078 9167
rect 3125 9164 3130 9169
rect 3134 9165 3136 9168
rect 3151 9167 3154 9173
rect 3500 9175 3519 9178
rect 3465 9171 3472 9174
rect 3497 9168 3500 9174
rect 3151 9164 3159 9167
rect 3523 9171 3530 9174
rect 3810 9169 3813 9174
rect 3817 9169 3820 9174
rect 3800 9166 3802 9169
rect 3810 9166 3820 9169
rect 3070 9161 3073 9164
rect 3151 9161 3154 9164
rect 2489 9148 2526 9152
rect 2530 9148 2556 9152
rect 2560 9148 2584 9152
rect 2588 9148 2776 9152
rect 2925 9145 2928 9149
rect 2952 9145 2953 9149
rect 2997 9145 2999 9149
rect 2489 9141 2507 9145
rect 2511 9141 2557 9145
rect 2561 9141 2608 9145
rect 2612 9141 2812 9145
rect 2870 9138 2882 9142
rect 2886 9138 2913 9142
rect 2917 9138 2935 9142
rect 2939 9138 3000 9142
rect 3004 9138 3018 9142
rect 3054 9135 3057 9153
rect 3135 9135 3138 9153
rect 3444 9152 3447 9164
rect 3465 9152 3468 9164
rect 3481 9152 3484 9164
rect 3500 9155 3512 9158
rect 3523 9152 3526 9164
rect 3539 9152 3542 9164
rect 3560 9152 3563 9164
rect 3810 9160 3813 9166
rect 3817 9160 3820 9166
rect 3826 9168 3829 9174
rect 3842 9169 3845 9174
rect 3826 9164 3828 9168
rect 3832 9164 3834 9168
rect 3842 9167 3848 9169
rect 3852 9167 3853 9169
rect 3842 9165 3853 9167
rect 3870 9167 3873 9174
rect 3826 9160 3829 9164
rect 3842 9160 3845 9165
rect 3871 9163 3873 9167
rect 3870 9160 3873 9163
rect 3886 9168 3889 9174
rect 3896 9168 3899 9174
rect 3917 9169 3920 9174
rect 3896 9164 3905 9168
rect 3917 9165 3918 9169
rect 3922 9166 3925 9169
rect 3942 9168 3945 9174
rect 3960 9169 3963 9174
rect 3999 9177 4002 9197
rect 4080 9177 4083 9197
rect 3886 9160 3889 9164
rect 3896 9160 3899 9164
rect 3917 9160 3920 9165
rect 3944 9164 3945 9168
rect 3942 9160 3945 9164
rect 3960 9160 3963 9165
rect 3990 9164 3995 9169
rect 3999 9165 4000 9168
rect 4015 9167 4018 9173
rect 4015 9164 4023 9167
rect 4070 9164 4075 9169
rect 4079 9165 4081 9168
rect 4096 9167 4099 9173
rect 4096 9164 4104 9167
rect 4015 9161 4018 9164
rect 4096 9161 4099 9164
rect 3434 9148 3471 9152
rect 3475 9148 3501 9152
rect 3505 9148 3529 9152
rect 3533 9148 3721 9152
rect 3870 9145 3873 9149
rect 3897 9145 3898 9149
rect 3942 9145 3944 9149
rect 3434 9141 3452 9145
rect 3456 9141 3502 9145
rect 3506 9141 3553 9145
rect 3557 9141 3757 9145
rect 3815 9138 3827 9142
rect 3831 9138 3858 9142
rect 3862 9138 3880 9142
rect 3884 9138 3945 9142
rect 3949 9138 3963 9142
rect 3999 9135 4002 9153
rect 4080 9135 4083 9153
rect 4403 9141 4829 9237
rect 2770 9131 2855 9135
rect 2859 9131 2871 9135
rect 2875 9131 2889 9135
rect 2893 9131 2900 9135
rect 2904 9131 2906 9135
rect 2910 9131 2925 9135
rect 2929 9131 2962 9135
rect 2966 9131 2967 9135
rect 2971 9131 2979 9135
rect 2983 9131 3007 9135
rect 3011 9131 3023 9135
rect 3027 9131 3047 9135
rect 3051 9131 3101 9135
rect 3105 9131 3128 9135
rect 3132 9131 3190 9135
rect 3194 9131 3205 9135
rect 3715 9131 3800 9135
rect 3804 9131 3816 9135
rect 3820 9131 3834 9135
rect 3838 9131 3845 9135
rect 3849 9131 3851 9135
rect 3855 9131 3870 9135
rect 3874 9131 3907 9135
rect 3911 9131 3912 9135
rect 3916 9131 3924 9135
rect 3928 9131 3952 9135
rect 3956 9131 3968 9135
rect 3972 9131 3992 9135
rect 3996 9131 4046 9135
rect 4050 9131 4073 9135
rect 4077 9131 4135 9135
rect 4139 9131 4150 9135
rect 4786 9131 4829 9141
rect 343 9119 386 9129
rect 2806 9124 2866 9128
rect 2870 9124 2882 9128
rect 2886 9124 2913 9128
rect 2917 9124 2935 9128
rect 2939 9124 3000 9128
rect 3004 9124 3018 9128
rect 3054 9121 3057 9131
rect 3084 9127 3087 9131
rect 3135 9127 3138 9131
rect 343 9109 376 9119
rect 2925 9117 2928 9121
rect 2952 9117 2953 9121
rect 2997 9117 2999 9121
rect 343 9099 366 9109
rect 343 9089 356 9099
rect 2854 9097 2857 9100
rect 2865 9100 2868 9106
rect 2872 9100 2875 9106
rect 2865 9097 2875 9100
rect 2865 9092 2868 9097
rect 343 9050 346 9089
rect 2872 9092 2875 9097
rect 2881 9102 2884 9106
rect 2881 9098 2883 9102
rect 2887 9098 2889 9102
rect 2897 9101 2900 9106
rect 2925 9103 2928 9106
rect 2897 9099 2908 9101
rect 2881 9092 2884 9098
rect 2897 9097 2903 9099
rect 2897 9092 2900 9097
rect 2907 9097 2908 9099
rect 2926 9099 2928 9103
rect 2925 9092 2928 9099
rect 3070 9110 3073 9113
rect 2941 9102 2944 9106
rect 2951 9102 2954 9106
rect 2951 9098 2960 9102
rect 2972 9101 2975 9106
rect 2997 9102 3000 9106
rect 2941 9092 2944 9098
rect 2951 9092 2954 9098
rect 2972 9097 2973 9101
rect 2977 9097 2980 9100
rect 2999 9098 3000 9102
rect 3015 9101 3018 9106
rect 3047 9106 3058 9109
rect 3070 9107 3078 9110
rect 2972 9092 2975 9097
rect 2997 9092 3000 9098
rect 3047 9100 3050 9106
rect 3070 9101 3073 9107
rect 3082 9102 3085 9105
rect 3093 9105 3096 9119
rect 3144 9114 3147 9119
rect 3159 9121 3162 9131
rect 3189 9127 3192 9131
rect 3128 9110 3129 9113
rect 3133 9110 3136 9113
rect 3365 9120 3621 9125
rect 3751 9124 3811 9128
rect 3815 9124 3827 9128
rect 3831 9124 3858 9128
rect 3862 9124 3880 9128
rect 3884 9124 3945 9128
rect 3949 9124 3963 9128
rect 3999 9121 4002 9131
rect 4029 9127 4032 9131
rect 4080 9127 4083 9131
rect 3175 9110 3178 9113
rect 3101 9105 3106 9110
rect 3144 9105 3147 9110
rect 3093 9102 3101 9105
rect 3015 9092 3018 9097
rect 3093 9097 3096 9102
rect 3152 9106 3163 9109
rect 3175 9107 3183 9110
rect 3045 9091 3050 9096
rect 2917 9079 2918 9083
rect 2942 9080 2943 9084
rect 2989 9079 2990 9083
rect 2794 9072 2870 9076
rect 2874 9072 2929 9076
rect 2933 9072 2954 9076
rect 2958 9072 2985 9076
rect 2989 9072 3018 9076
rect 3054 9069 3057 9097
rect 3084 9069 3087 9093
rect 3135 9069 3138 9101
rect 3152 9100 3155 9106
rect 3175 9101 3178 9107
rect 3187 9102 3190 9105
rect 3198 9105 3201 9119
rect 3870 9117 3873 9121
rect 3897 9117 3898 9121
rect 3942 9117 3944 9121
rect 3198 9102 3204 9105
rect 3363 9102 3383 9106
rect 3387 9102 3437 9106
rect 3441 9102 3580 9106
rect 3584 9102 3668 9106
rect 3198 9097 3201 9102
rect 3150 9091 3155 9096
rect 3159 9069 3162 9097
rect 3366 9098 3369 9102
rect 3189 9069 3192 9093
rect 3375 9085 3378 9090
rect 3390 9092 3393 9102
rect 3420 9098 3423 9102
rect 3359 9081 3360 9084
rect 3364 9081 3367 9084
rect 3406 9081 3409 9084
rect 3375 9076 3378 9081
rect 3383 9077 3394 9080
rect 3406 9078 3414 9081
rect 3406 9072 3409 9078
rect 3418 9073 3421 9076
rect 3429 9076 3432 9090
rect 3540 9095 3543 9102
rect 3593 9095 3596 9102
rect 3799 9097 3802 9100
rect 3810 9100 3813 9106
rect 3817 9100 3820 9106
rect 3810 9097 3820 9100
rect 3429 9073 3441 9076
rect 2782 9065 2856 9069
rect 2860 9065 2862 9069
rect 2866 9065 2870 9069
rect 2874 9065 2888 9069
rect 2892 9065 2897 9069
rect 2901 9065 2906 9069
rect 2910 9065 2929 9069
rect 2933 9065 2963 9069
rect 2967 9065 2978 9069
rect 2982 9065 3006 9069
rect 3010 9065 3023 9069
rect 3027 9065 3047 9069
rect 3051 9065 3101 9069
rect 3105 9065 3128 9069
rect 3132 9065 3152 9069
rect 3156 9065 3204 9069
rect 2794 9058 2870 9062
rect 2874 9058 2929 9062
rect 2933 9058 2954 9062
rect 2958 9058 2985 9062
rect 2989 9058 3018 9062
rect 2917 9051 2918 9055
rect 2942 9050 2943 9054
rect 2989 9051 2990 9055
rect 86 9047 346 9050
rect 3054 9046 3057 9065
rect 3159 9046 3162 9065
rect 2865 9037 2868 9042
rect 2872 9037 2875 9042
rect 2855 9034 2857 9037
rect 2865 9034 2875 9037
rect 2865 9028 2868 9034
rect 2872 9028 2875 9034
rect 2881 9036 2884 9042
rect 2897 9037 2900 9042
rect 2881 9032 2883 9036
rect 2887 9032 2889 9036
rect 2897 9035 2903 9037
rect 2907 9035 2908 9037
rect 2897 9033 2908 9035
rect 2925 9035 2928 9042
rect 2881 9028 2884 9032
rect 2897 9028 2900 9033
rect 2926 9031 2928 9035
rect 2925 9028 2928 9031
rect 2941 9036 2944 9042
rect 2951 9036 2954 9042
rect 2972 9037 2975 9042
rect 2951 9032 2960 9036
rect 2972 9033 2973 9037
rect 2977 9034 2980 9037
rect 2997 9036 3000 9042
rect 3015 9037 3018 9042
rect 2941 9028 2944 9032
rect 2951 9028 2954 9032
rect 2972 9028 2975 9033
rect 2999 9032 3000 9036
rect 3044 9033 3049 9038
rect 3053 9034 3055 9037
rect 3070 9036 3073 9042
rect 3070 9033 3078 9036
rect 3150 9033 3155 9038
rect 3159 9034 3160 9037
rect 3175 9036 3178 9042
rect 3175 9033 3183 9036
rect 2997 9028 3000 9032
rect 3015 9028 3018 9033
rect 3070 9030 3073 9033
rect 3175 9030 3178 9033
rect 3366 9026 3369 9072
rect 3429 9068 3432 9073
rect 3390 9026 3393 9068
rect 3420 9026 3423 9064
rect 3438 9058 3441 9073
rect 3810 9092 3813 9097
rect 3817 9092 3820 9097
rect 3826 9102 3829 9106
rect 3826 9098 3828 9102
rect 3832 9098 3834 9102
rect 3842 9101 3845 9106
rect 3870 9103 3873 9106
rect 3842 9099 3853 9101
rect 3826 9092 3829 9098
rect 3842 9097 3848 9099
rect 3842 9092 3845 9097
rect 3852 9097 3853 9099
rect 3871 9099 3873 9103
rect 3870 9092 3873 9099
rect 4015 9110 4018 9113
rect 3886 9102 3889 9106
rect 3896 9102 3899 9106
rect 3896 9098 3905 9102
rect 3917 9101 3920 9106
rect 3942 9102 3945 9106
rect 3886 9092 3889 9098
rect 3896 9092 3899 9098
rect 3917 9097 3918 9101
rect 3922 9097 3925 9100
rect 3944 9098 3945 9102
rect 3960 9101 3963 9106
rect 3992 9106 4003 9109
rect 4015 9107 4023 9110
rect 3917 9092 3920 9097
rect 3942 9092 3945 9098
rect 3992 9100 3995 9106
rect 4015 9101 4018 9107
rect 4027 9102 4030 9105
rect 4038 9105 4041 9119
rect 4089 9114 4092 9119
rect 4104 9121 4107 9131
rect 4134 9127 4137 9131
rect 4073 9110 4074 9113
rect 4078 9110 4081 9113
rect 4796 9121 4829 9131
rect 4120 9110 4123 9113
rect 4046 9105 4051 9110
rect 4089 9105 4092 9110
rect 4038 9102 4046 9105
rect 3960 9092 3963 9097
rect 4038 9097 4041 9102
rect 4097 9106 4108 9109
rect 4120 9107 4128 9110
rect 3990 9091 3995 9096
rect 3862 9079 3863 9083
rect 3887 9080 3888 9084
rect 3934 9079 3935 9083
rect 3739 9072 3815 9076
rect 3819 9072 3874 9076
rect 3878 9072 3899 9076
rect 3903 9072 3930 9076
rect 3934 9072 3963 9076
rect 3999 9069 4002 9097
rect 4029 9069 4032 9093
rect 4080 9069 4083 9101
rect 4097 9100 4100 9106
rect 4120 9101 4123 9107
rect 4132 9102 4135 9105
rect 4143 9105 4146 9119
rect 4806 9111 4829 9121
rect 4143 9102 4149 9105
rect 4143 9097 4146 9102
rect 4816 9101 4829 9111
rect 4095 9091 4100 9096
rect 4104 9069 4107 9097
rect 4134 9069 4137 9093
rect 3727 9065 3801 9069
rect 3805 9065 3807 9069
rect 3811 9065 3815 9069
rect 3819 9065 3833 9069
rect 3837 9065 3842 9069
rect 3846 9065 3851 9069
rect 3855 9065 3874 9069
rect 3878 9065 3908 9069
rect 3912 9065 3923 9069
rect 3927 9065 3951 9069
rect 3955 9065 3968 9069
rect 3972 9065 3992 9069
rect 3996 9065 4046 9069
rect 4050 9065 4073 9069
rect 4077 9065 4097 9069
rect 4101 9065 4149 9069
rect 3438 9053 3555 9058
rect 3573 9057 3576 9065
rect 3573 9053 3593 9057
rect 3597 9053 3608 9057
rect 3573 9045 3576 9053
rect 3626 9049 3629 9065
rect 3739 9058 3815 9062
rect 3819 9058 3874 9062
rect 3878 9058 3899 9062
rect 3903 9058 3930 9062
rect 3934 9058 3963 9062
rect 3862 9051 3863 9055
rect 3887 9050 3888 9054
rect 3934 9051 3935 9055
rect 3630 9045 3745 9049
rect 3999 9046 4002 9065
rect 4104 9046 4107 9065
rect 4826 9062 4829 9101
rect 5083 9062 5086 9316
rect 4483 9056 4484 9060
rect 4488 9056 4489 9060
rect 4493 9056 4494 9060
rect 4498 9056 4499 9060
rect 4503 9056 4504 9060
rect 4508 9056 4509 9060
rect 4479 9055 4513 9056
rect 4483 9051 4484 9055
rect 4488 9051 4489 9055
rect 4493 9051 4494 9055
rect 4498 9051 4499 9055
rect 4503 9051 4504 9055
rect 4508 9051 4509 9055
rect 4479 9050 4513 9051
rect 4483 9046 4484 9050
rect 4488 9046 4489 9050
rect 4493 9046 4494 9050
rect 4498 9046 4499 9050
rect 4503 9046 4504 9050
rect 4508 9046 4509 9050
rect 3672 9033 3709 9037
rect 3810 9037 3813 9042
rect 3817 9037 3820 9042
rect 3800 9034 3802 9037
rect 3810 9034 3820 9037
rect 3540 9026 3543 9033
rect 3593 9026 3596 9033
rect 3660 9026 3721 9030
rect 3810 9028 3813 9034
rect 3363 9022 3383 9026
rect 3387 9022 3437 9026
rect 3441 9022 3580 9026
rect 3584 9022 3660 9026
rect 617 9012 618 9016
rect 622 9012 623 9016
rect 627 9012 628 9016
rect 632 9012 633 9016
rect 637 9012 638 9016
rect 642 9012 643 9016
rect 613 9011 647 9012
rect 617 9007 618 9011
rect 622 9007 623 9011
rect 627 9007 628 9011
rect 632 9007 633 9011
rect 637 9007 638 9011
rect 642 9007 643 9011
rect 613 9006 647 9007
rect 617 9002 618 9006
rect 622 9002 623 9006
rect 627 9002 628 9006
rect 632 9002 633 9006
rect 637 9002 638 9006
rect 642 9002 643 9006
rect 613 9001 647 9002
rect 86 8995 346 8998
rect 617 8997 618 9001
rect 622 8997 623 9001
rect 627 8997 628 9001
rect 632 8997 633 9001
rect 637 8997 638 9001
rect 642 8997 643 9001
rect 663 9012 664 9016
rect 668 9012 669 9016
rect 673 9012 674 9016
rect 678 9012 679 9016
rect 683 9012 684 9016
rect 688 9012 689 9016
rect 2925 9013 2928 9017
rect 2952 9013 2953 9017
rect 2997 9013 2999 9017
rect 659 9011 693 9012
rect 663 9007 664 9011
rect 668 9007 669 9011
rect 673 9007 674 9011
rect 678 9007 679 9011
rect 683 9007 684 9011
rect 688 9007 689 9011
rect 659 9006 693 9007
rect 2806 9006 2882 9010
rect 2886 9006 2913 9010
rect 2917 9006 2935 9010
rect 2939 9006 3000 9010
rect 3004 9006 3018 9010
rect 663 9002 664 9006
rect 668 9002 669 9006
rect 673 9002 674 9006
rect 678 9002 679 9006
rect 683 9002 684 9006
rect 688 9002 689 9006
rect 3054 9003 3057 9022
rect 3159 9003 3162 9022
rect 3390 9012 3393 9022
rect 3680 9017 3781 9021
rect 3817 9028 3820 9034
rect 3826 9036 3829 9042
rect 3842 9037 3845 9042
rect 3826 9032 3828 9036
rect 3832 9032 3834 9036
rect 3842 9035 3848 9037
rect 3852 9035 3853 9037
rect 3842 9033 3853 9035
rect 3870 9035 3873 9042
rect 3826 9028 3829 9032
rect 3842 9028 3845 9033
rect 3871 9031 3873 9035
rect 3870 9028 3873 9031
rect 3886 9036 3889 9042
rect 3896 9036 3899 9042
rect 3917 9037 3920 9042
rect 3896 9032 3905 9036
rect 3917 9033 3918 9037
rect 3922 9034 3925 9037
rect 3942 9036 3945 9042
rect 3960 9037 3963 9042
rect 3886 9028 3889 9032
rect 3896 9028 3899 9032
rect 3917 9028 3920 9033
rect 3944 9032 3945 9036
rect 3989 9033 3994 9038
rect 3998 9034 4000 9037
rect 4015 9036 4018 9042
rect 4015 9033 4023 9036
rect 4095 9033 4100 9038
rect 4104 9034 4105 9037
rect 4120 9036 4123 9042
rect 4479 9045 4513 9046
rect 4483 9041 4484 9045
rect 4488 9041 4489 9045
rect 4493 9041 4494 9045
rect 4498 9041 4499 9045
rect 4503 9041 4504 9045
rect 4508 9041 4509 9045
rect 4529 9056 4530 9060
rect 4534 9056 4535 9060
rect 4539 9056 4540 9060
rect 4544 9056 4545 9060
rect 4549 9056 4550 9060
rect 4554 9056 4555 9060
rect 4826 9059 5086 9062
rect 4525 9055 4559 9056
rect 4529 9051 4530 9055
rect 4534 9051 4535 9055
rect 4539 9051 4540 9055
rect 4544 9051 4545 9055
rect 4549 9051 4550 9055
rect 4554 9051 4555 9055
rect 4525 9050 4559 9051
rect 4529 9046 4530 9050
rect 4534 9046 4535 9050
rect 4539 9046 4540 9050
rect 4544 9046 4545 9050
rect 4549 9046 4550 9050
rect 4554 9046 4555 9050
rect 4525 9045 4559 9046
rect 4529 9041 4530 9045
rect 4534 9041 4535 9045
rect 4539 9041 4540 9045
rect 4544 9041 4545 9045
rect 4549 9041 4550 9045
rect 4554 9041 4555 9045
rect 4120 9033 4128 9036
rect 3942 9028 3945 9032
rect 3960 9028 3963 9033
rect 4015 9030 4018 9033
rect 4120 9030 4123 9033
rect 3870 9013 3873 9017
rect 3897 9013 3898 9017
rect 3942 9013 3944 9017
rect 3598 9008 3733 9012
rect 659 9001 693 9002
rect 663 8997 664 9001
rect 668 8997 669 9001
rect 673 8997 674 9001
rect 678 8997 679 9001
rect 683 8997 684 9001
rect 688 8997 689 9001
rect 2770 8999 2855 9003
rect 2859 8999 2871 9003
rect 2875 8999 2889 9003
rect 2893 8999 2900 9003
rect 2904 8999 2906 9003
rect 2910 8999 2925 9003
rect 2929 8999 2962 9003
rect 2966 8999 2967 9003
rect 2971 8999 2979 9003
rect 2983 8999 3007 9003
rect 3011 8999 3023 9003
rect 3027 8999 3047 9003
rect 3051 8999 3101 9003
rect 3105 8999 3128 9003
rect 3132 8999 3182 9003
rect 3186 8999 3190 9003
rect 3194 8999 3218 9003
rect 3222 8999 3272 9003
rect 3330 9000 3391 9003
rect 3406 9002 3409 9008
rect 3751 9006 3827 9010
rect 3831 9006 3858 9010
rect 3862 9006 3880 9010
rect 3884 9006 3945 9010
rect 3949 9006 3963 9010
rect 3999 9003 4002 9022
rect 4104 9003 4107 9022
rect 4826 9007 5086 9010
rect 3406 8999 3414 9002
rect 3715 8999 3800 9003
rect 3804 8999 3816 9003
rect 3820 8999 3834 9003
rect 3838 8999 3845 9003
rect 3849 8999 3851 9003
rect 3855 8999 3870 9003
rect 3874 8999 3907 9003
rect 3911 8999 3912 9003
rect 3916 8999 3924 9003
rect 3928 8999 3952 9003
rect 3956 8999 3968 9003
rect 3972 8999 3992 9003
rect 3996 8999 4046 9003
rect 4050 8999 4073 9003
rect 4077 8999 4127 9003
rect 4131 8999 4135 9003
rect 4139 8999 4163 9003
rect 4167 8999 4217 9003
rect 86 8741 89 8995
rect 343 8956 346 8995
rect 2806 8992 2882 8996
rect 2886 8992 2913 8996
rect 2917 8992 2935 8996
rect 2939 8992 3000 8996
rect 3004 8992 3018 8996
rect 3054 8989 3057 8999
rect 3084 8995 3087 8999
rect 3111 8995 3114 8999
rect 2925 8985 2928 8989
rect 2952 8985 2953 8989
rect 2997 8985 2999 8989
rect 2854 8965 2857 8968
rect 2865 8968 2868 8974
rect 2872 8968 2875 8974
rect 2865 8965 2875 8968
rect 2865 8960 2868 8965
rect 2872 8960 2875 8965
rect 2881 8970 2884 8974
rect 2881 8966 2883 8970
rect 2887 8966 2889 8970
rect 2897 8969 2900 8974
rect 2925 8971 2928 8974
rect 2897 8967 2908 8969
rect 2881 8960 2884 8966
rect 2897 8965 2903 8967
rect 2897 8960 2900 8965
rect 2907 8965 2908 8967
rect 2926 8967 2928 8971
rect 2925 8960 2928 8967
rect 3070 8978 3073 8981
rect 2941 8970 2944 8974
rect 2951 8970 2954 8974
rect 2951 8966 2960 8970
rect 2972 8969 2975 8974
rect 2997 8970 3000 8974
rect 2941 8960 2944 8966
rect 2951 8960 2954 8966
rect 2972 8965 2973 8969
rect 2977 8965 2980 8968
rect 2999 8966 3000 8970
rect 3015 8969 3018 8974
rect 3047 8974 3058 8977
rect 3070 8975 3078 8978
rect 2972 8960 2975 8965
rect 2997 8960 3000 8966
rect 3047 8968 3050 8974
rect 3070 8969 3073 8975
rect 3082 8970 3085 8973
rect 3093 8973 3096 8987
rect 3120 8982 3123 8987
rect 3135 8989 3138 8999
rect 3165 8995 3168 8999
rect 3201 8995 3204 8999
rect 3104 8978 3105 8981
rect 3109 8978 3112 8981
rect 3151 8978 3154 8981
rect 3093 8970 3101 8973
rect 3120 8973 3123 8978
rect 3015 8960 3018 8965
rect 3093 8965 3096 8970
rect 3101 8966 3105 8970
rect 3128 8974 3139 8977
rect 3151 8975 3159 8978
rect 3045 8959 3050 8964
rect 343 8946 356 8956
rect 2917 8947 2918 8951
rect 2942 8948 2943 8952
rect 2989 8947 2990 8951
rect 343 8936 366 8946
rect 2794 8940 2870 8944
rect 2874 8940 2929 8944
rect 2933 8940 2954 8944
rect 2958 8940 2985 8944
rect 2989 8940 3018 8944
rect 3054 8937 3057 8965
rect 3084 8937 3087 8961
rect 3111 8937 3114 8969
rect 3128 8968 3131 8974
rect 3151 8969 3154 8975
rect 3163 8970 3166 8973
rect 3174 8973 3177 8987
rect 3210 8982 3213 8987
rect 3225 8989 3228 8999
rect 3255 8995 3258 8999
rect 3406 8996 3409 8999
rect 3199 8978 3202 8981
rect 3241 8978 3244 8981
rect 3174 8970 3183 8973
rect 3210 8973 3213 8978
rect 3174 8965 3177 8970
rect 3126 8959 3131 8964
rect 3135 8937 3138 8965
rect 3217 8976 3229 8977
rect 3221 8974 3229 8976
rect 3241 8975 3249 8978
rect 3241 8969 3244 8975
rect 3253 8970 3256 8973
rect 3264 8973 3267 8987
rect 3751 8992 3827 8996
rect 3831 8992 3858 8996
rect 3862 8992 3880 8996
rect 3884 8992 3945 8996
rect 3949 8992 3963 8996
rect 3999 8989 4002 8999
rect 4029 8995 4032 8999
rect 4056 8995 4059 8999
rect 3390 8976 3393 8988
rect 3870 8985 3873 8989
rect 3897 8985 3898 8989
rect 3942 8985 3944 8989
rect 3264 8970 3284 8973
rect 3165 8937 3168 8961
rect 3201 8937 3204 8969
rect 3264 8965 3267 8970
rect 3341 8972 3359 8976
rect 3363 8972 3383 8976
rect 3387 8972 3437 8976
rect 3441 8972 3486 8976
rect 3490 8972 3668 8976
rect 3225 8937 3228 8965
rect 3344 8968 3347 8972
rect 3366 8968 3369 8972
rect 3255 8937 3258 8961
rect 3353 8955 3356 8960
rect 3375 8955 3378 8960
rect 3390 8962 3393 8972
rect 3420 8968 3423 8972
rect 3337 8951 3338 8954
rect 3342 8951 3345 8954
rect 3357 8951 3360 8955
rect 3364 8951 3367 8954
rect 3406 8951 3409 8954
rect 3353 8946 3356 8951
rect 3375 8946 3378 8951
rect 3383 8947 3394 8950
rect 3406 8948 3414 8951
rect 3406 8942 3409 8948
rect 3418 8943 3421 8946
rect 3429 8946 3432 8960
rect 3446 8965 3449 8972
rect 3499 8965 3502 8972
rect 3799 8965 3802 8968
rect 3810 8968 3813 8974
rect 3817 8968 3820 8974
rect 3810 8965 3820 8968
rect 3429 8943 3441 8946
rect 343 8926 376 8936
rect 2782 8933 2856 8937
rect 2860 8933 2862 8937
rect 2866 8933 2870 8937
rect 2874 8933 2888 8937
rect 2892 8933 2897 8937
rect 2901 8933 2906 8937
rect 2910 8933 2929 8937
rect 2933 8933 2963 8937
rect 2967 8933 2978 8937
rect 2982 8933 3006 8937
rect 3010 8933 3023 8937
rect 3027 8933 3047 8937
rect 3051 8933 3101 8937
rect 3108 8933 3128 8937
rect 3132 8933 3182 8937
rect 3186 8933 3218 8937
rect 3222 8933 3272 8937
rect 2794 8926 2870 8930
rect 2874 8926 2929 8930
rect 2933 8926 2954 8930
rect 2958 8926 2985 8930
rect 2989 8926 3018 8930
rect 343 8916 386 8926
rect 2917 8919 2918 8923
rect 2942 8918 2943 8922
rect 2989 8919 2990 8923
rect 343 8820 769 8916
rect 2865 8905 2868 8910
rect 2872 8905 2875 8910
rect 2855 8902 2857 8905
rect 2865 8902 2875 8905
rect 2865 8896 2868 8902
rect 2872 8896 2875 8902
rect 2881 8904 2884 8910
rect 2897 8905 2900 8910
rect 2881 8900 2883 8904
rect 2887 8900 2889 8904
rect 2897 8903 2903 8905
rect 2907 8903 2908 8905
rect 2897 8901 2908 8903
rect 2925 8903 2928 8910
rect 2881 8896 2884 8900
rect 2897 8896 2900 8901
rect 2926 8899 2928 8903
rect 2925 8896 2928 8899
rect 2941 8904 2944 8910
rect 2951 8904 2954 8910
rect 2972 8905 2975 8910
rect 2951 8900 2960 8904
rect 2972 8901 2973 8905
rect 2977 8902 2980 8905
rect 2997 8904 3000 8910
rect 3015 8905 3018 8910
rect 3054 8911 3057 8933
rect 3135 8911 3138 8933
rect 3225 8911 3228 8933
rect 2941 8896 2944 8900
rect 2951 8896 2954 8900
rect 2972 8896 2975 8901
rect 2999 8900 3000 8904
rect 2997 8896 3000 8900
rect 3015 8896 3018 8901
rect 3045 8898 3050 8903
rect 3054 8899 3055 8902
rect 3070 8901 3073 8907
rect 3070 8898 3078 8901
rect 3125 8898 3130 8903
rect 3134 8899 3136 8902
rect 3151 8901 3154 8907
rect 3151 8898 3159 8901
rect 3218 8899 3226 8902
rect 3241 8901 3244 8907
rect 3241 8898 3249 8901
rect 3070 8895 3073 8898
rect 3151 8895 3154 8898
rect 3241 8895 3244 8898
rect 3344 8896 3347 8942
rect 3366 8896 3369 8942
rect 3429 8938 3432 8943
rect 3390 8896 3393 8938
rect 3420 8896 3423 8934
rect 3438 8928 3441 8943
rect 3810 8960 3813 8965
rect 3817 8960 3820 8965
rect 3826 8970 3829 8974
rect 3826 8966 3828 8970
rect 3832 8966 3834 8970
rect 3842 8969 3845 8974
rect 3870 8971 3873 8974
rect 3842 8967 3853 8969
rect 3826 8960 3829 8966
rect 3842 8965 3848 8967
rect 3842 8960 3845 8965
rect 3852 8965 3853 8967
rect 3871 8967 3873 8971
rect 3870 8960 3873 8967
rect 4015 8978 4018 8981
rect 3886 8970 3889 8974
rect 3896 8970 3899 8974
rect 3896 8966 3905 8970
rect 3917 8969 3920 8974
rect 3942 8970 3945 8974
rect 3886 8960 3889 8966
rect 3896 8960 3899 8966
rect 3917 8965 3918 8969
rect 3922 8965 3925 8968
rect 3944 8966 3945 8970
rect 3960 8969 3963 8974
rect 3992 8974 4003 8977
rect 4015 8975 4023 8978
rect 3917 8960 3920 8965
rect 3942 8960 3945 8966
rect 3992 8968 3995 8974
rect 4015 8969 4018 8975
rect 4027 8970 4030 8973
rect 4038 8973 4041 8987
rect 4065 8982 4068 8987
rect 4080 8989 4083 8999
rect 4110 8995 4113 8999
rect 4146 8995 4149 8999
rect 4049 8978 4050 8981
rect 4054 8978 4057 8981
rect 4096 8978 4099 8981
rect 4038 8970 4046 8973
rect 4065 8973 4068 8978
rect 3960 8960 3963 8965
rect 4038 8965 4041 8970
rect 4046 8966 4050 8970
rect 4073 8974 4084 8977
rect 4096 8975 4104 8978
rect 3990 8959 3995 8964
rect 3862 8947 3863 8951
rect 3887 8948 3888 8952
rect 3934 8947 3935 8951
rect 3739 8940 3815 8944
rect 3819 8940 3874 8944
rect 3878 8940 3899 8944
rect 3903 8940 3930 8944
rect 3934 8940 3963 8944
rect 3999 8937 4002 8965
rect 4029 8937 4032 8961
rect 4056 8937 4059 8969
rect 4073 8968 4076 8974
rect 4096 8969 4099 8975
rect 4108 8970 4111 8973
rect 4119 8973 4122 8987
rect 4155 8982 4158 8987
rect 4170 8989 4173 8999
rect 4200 8995 4203 8999
rect 4144 8978 4147 8981
rect 4186 8978 4189 8981
rect 4119 8970 4128 8973
rect 4155 8973 4158 8978
rect 4119 8965 4122 8970
rect 4071 8959 4076 8964
rect 4080 8937 4083 8965
rect 4162 8976 4174 8977
rect 4166 8974 4174 8976
rect 4186 8975 4194 8978
rect 4186 8969 4189 8975
rect 4198 8970 4201 8973
rect 4209 8973 4212 8987
rect 4209 8970 4229 8973
rect 4110 8937 4113 8961
rect 4146 8937 4149 8969
rect 4209 8965 4212 8970
rect 4826 8968 4829 9007
rect 4170 8937 4173 8965
rect 4200 8937 4203 8961
rect 4816 8958 4829 8968
rect 4806 8948 4829 8958
rect 4796 8938 4829 8948
rect 3438 8923 3461 8928
rect 3479 8927 3482 8935
rect 3479 8923 3488 8927
rect 3492 8923 3514 8927
rect 3479 8915 3482 8923
rect 3532 8919 3535 8935
rect 3727 8933 3801 8937
rect 3805 8933 3807 8937
rect 3811 8933 3815 8937
rect 3819 8933 3833 8937
rect 3837 8933 3842 8937
rect 3846 8933 3851 8937
rect 3855 8933 3874 8937
rect 3878 8933 3908 8937
rect 3912 8933 3923 8937
rect 3927 8933 3951 8937
rect 3955 8933 3968 8937
rect 3972 8933 3992 8937
rect 3996 8933 4046 8937
rect 4053 8933 4073 8937
rect 4077 8933 4127 8937
rect 4131 8933 4163 8937
rect 4167 8933 4217 8937
rect 3739 8926 3815 8930
rect 3819 8926 3874 8930
rect 3878 8926 3899 8930
rect 3903 8926 3930 8930
rect 3934 8926 3963 8930
rect 3862 8919 3863 8923
rect 3887 8918 3888 8922
rect 3934 8919 3935 8923
rect 3536 8915 3769 8916
rect 3535 8912 3769 8915
rect 3446 8896 3449 8903
rect 3499 8896 3502 8903
rect 3810 8905 3813 8910
rect 3817 8905 3820 8910
rect 3800 8902 3802 8905
rect 3810 8902 3820 8905
rect 3810 8896 3813 8902
rect 2925 8881 2928 8885
rect 2952 8881 2953 8885
rect 2997 8881 2999 8885
rect 3341 8892 3359 8896
rect 3363 8892 3383 8896
rect 3387 8892 3437 8896
rect 3441 8892 3486 8896
rect 3490 8892 3660 8896
rect 2806 8874 2882 8878
rect 2886 8874 2913 8878
rect 2917 8874 2935 8878
rect 2939 8874 3000 8878
rect 3004 8874 3018 8878
rect 3054 8871 3057 8887
rect 3135 8871 3138 8887
rect 3225 8871 3228 8887
rect 3390 8882 3393 8892
rect 3817 8896 3820 8902
rect 3826 8904 3829 8910
rect 3842 8905 3845 8910
rect 3826 8900 3828 8904
rect 3832 8900 3834 8904
rect 3842 8903 3848 8905
rect 3852 8903 3853 8905
rect 3842 8901 3853 8903
rect 3870 8903 3873 8910
rect 3826 8896 3829 8900
rect 3842 8896 3845 8901
rect 3871 8899 3873 8903
rect 3870 8896 3873 8899
rect 3886 8904 3889 8910
rect 3896 8904 3899 8910
rect 3917 8905 3920 8910
rect 3896 8900 3905 8904
rect 3917 8901 3918 8905
rect 3922 8902 3925 8905
rect 3942 8904 3945 8910
rect 3960 8905 3963 8910
rect 3999 8911 4002 8933
rect 4080 8911 4083 8933
rect 4170 8911 4173 8933
rect 4786 8928 4829 8938
rect 3886 8896 3889 8900
rect 3896 8896 3899 8900
rect 3917 8896 3920 8901
rect 3944 8900 3945 8904
rect 3942 8896 3945 8900
rect 3960 8896 3963 8901
rect 3990 8898 3995 8903
rect 3999 8899 4000 8902
rect 4015 8901 4018 8907
rect 4015 8898 4023 8901
rect 4070 8898 4075 8903
rect 4079 8899 4081 8902
rect 4096 8901 4099 8907
rect 4096 8898 4104 8901
rect 4163 8899 4171 8902
rect 4186 8901 4189 8907
rect 4186 8898 4194 8901
rect 4015 8895 4018 8898
rect 4096 8895 4099 8898
rect 4186 8895 4189 8898
rect 3492 8882 3757 8886
rect 3870 8881 3873 8885
rect 3897 8881 3898 8885
rect 3942 8881 3944 8885
rect 2770 8867 2855 8871
rect 2859 8867 2871 8871
rect 2875 8867 2889 8871
rect 2893 8867 2900 8871
rect 2904 8867 2906 8871
rect 2910 8867 2925 8871
rect 2929 8867 2962 8871
rect 2966 8867 2967 8871
rect 2971 8867 2979 8871
rect 2983 8867 3007 8871
rect 3011 8867 3023 8871
rect 3027 8867 3047 8871
rect 3051 8867 3101 8871
rect 3105 8867 3128 8871
rect 3132 8867 3218 8871
rect 3222 8867 3276 8871
rect 3332 8870 3391 8873
rect 3406 8872 3409 8878
rect 3751 8874 3827 8878
rect 3831 8874 3858 8878
rect 3862 8874 3880 8878
rect 3884 8874 3945 8878
rect 3949 8874 3963 8878
rect 3406 8869 3414 8872
rect 3999 8871 4002 8887
rect 4080 8871 4083 8887
rect 4170 8871 4173 8887
rect 2806 8860 2882 8864
rect 2886 8860 2913 8864
rect 2917 8860 2935 8864
rect 2939 8860 3000 8864
rect 3004 8860 3018 8864
rect 3054 8857 3057 8867
rect 3084 8863 3087 8867
rect 3406 8866 3409 8869
rect 3715 8867 3800 8871
rect 3804 8867 3816 8871
rect 3820 8867 3834 8871
rect 3838 8867 3845 8871
rect 3849 8867 3851 8871
rect 3855 8867 3870 8871
rect 3874 8867 3907 8871
rect 3911 8867 3912 8871
rect 3916 8867 3924 8871
rect 3928 8867 3952 8871
rect 3956 8867 3968 8871
rect 3972 8867 3992 8871
rect 3996 8867 4046 8871
rect 4050 8867 4073 8871
rect 4077 8867 4163 8871
rect 4167 8867 4221 8871
rect 2925 8853 2928 8857
rect 2952 8853 2953 8857
rect 2997 8853 2999 8857
rect 2854 8833 2857 8836
rect 2865 8836 2868 8842
rect 2872 8836 2875 8842
rect 2865 8833 2875 8836
rect 2865 8828 2868 8833
rect 2872 8828 2875 8833
rect 2881 8838 2884 8842
rect 2881 8834 2883 8838
rect 2887 8834 2889 8838
rect 2897 8837 2900 8842
rect 2925 8839 2928 8842
rect 2897 8835 2908 8837
rect 2881 8828 2884 8834
rect 2897 8833 2903 8835
rect 2897 8828 2900 8833
rect 2907 8833 2908 8835
rect 2926 8835 2928 8839
rect 2925 8828 2928 8835
rect 3070 8846 3073 8849
rect 2941 8838 2944 8842
rect 2951 8838 2954 8842
rect 2951 8834 2960 8838
rect 2972 8837 2975 8842
rect 2997 8838 3000 8842
rect 2941 8828 2944 8834
rect 2951 8828 2954 8834
rect 2972 8833 2973 8837
rect 2977 8833 2980 8836
rect 2999 8834 3000 8838
rect 3015 8837 3018 8842
rect 3047 8842 3058 8845
rect 3070 8843 3078 8846
rect 2972 8828 2975 8833
rect 2997 8828 3000 8834
rect 3047 8836 3050 8842
rect 3070 8837 3073 8843
rect 3082 8838 3085 8841
rect 3093 8841 3096 8855
rect 3751 8860 3827 8864
rect 3831 8860 3858 8864
rect 3862 8860 3880 8864
rect 3884 8860 3945 8864
rect 3949 8860 3963 8864
rect 3390 8846 3393 8858
rect 3999 8857 4002 8867
rect 4029 8863 4032 8867
rect 3870 8853 3873 8857
rect 3897 8853 3898 8857
rect 3942 8853 3944 8857
rect 3101 8841 3106 8846
rect 3359 8842 3383 8846
rect 3387 8842 3668 8846
rect 3093 8838 3101 8841
rect 3015 8828 3018 8833
rect 3093 8833 3096 8838
rect 3799 8833 3802 8836
rect 3810 8836 3813 8842
rect 3817 8836 3820 8842
rect 3810 8833 3820 8836
rect 3045 8827 3050 8832
rect 343 8810 386 8820
rect 2355 8819 2476 8823
rect 2364 8812 2373 8816
rect 2377 8812 2409 8816
rect 2413 8812 2476 8816
rect 2480 8812 2505 8816
rect 2509 8812 2541 8816
rect 2545 8812 2608 8816
rect 2612 8812 2637 8816
rect 2641 8812 2673 8816
rect 2677 8812 2740 8816
rect 2744 8812 2824 8816
rect 2917 8815 2918 8819
rect 2942 8816 2943 8820
rect 2989 8815 2990 8819
rect 343 8800 376 8810
rect 2364 8805 2397 8809
rect 2401 8805 2425 8809
rect 2429 8805 2455 8809
rect 2459 8805 2492 8809
rect 2496 8805 2529 8809
rect 2533 8805 2557 8809
rect 2561 8805 2587 8809
rect 2591 8805 2624 8809
rect 2628 8805 2661 8809
rect 2665 8805 2689 8809
rect 2693 8805 2719 8809
rect 2723 8805 2756 8809
rect 2760 8805 2764 8809
rect 2849 8808 2870 8812
rect 2874 8808 2879 8812
rect 2883 8808 2929 8812
rect 2933 8808 2954 8812
rect 2958 8808 2985 8812
rect 2989 8808 3018 8812
rect 3054 8805 3057 8833
rect 3084 8805 3087 8829
rect 3810 8828 3813 8833
rect 3817 8828 3820 8833
rect 3826 8838 3829 8842
rect 3826 8834 3828 8838
rect 3832 8834 3834 8838
rect 3842 8837 3845 8842
rect 3870 8839 3873 8842
rect 3842 8835 3853 8837
rect 3826 8828 3829 8834
rect 3842 8833 3848 8835
rect 3842 8828 3845 8833
rect 3852 8833 3853 8835
rect 3871 8835 3873 8839
rect 3870 8828 3873 8835
rect 4015 8846 4018 8849
rect 3886 8838 3889 8842
rect 3896 8838 3899 8842
rect 3896 8834 3905 8838
rect 3917 8837 3920 8842
rect 3942 8838 3945 8842
rect 3886 8828 3889 8834
rect 3896 8828 3899 8834
rect 3917 8833 3918 8837
rect 3922 8833 3925 8836
rect 3944 8834 3945 8838
rect 3960 8837 3963 8842
rect 3992 8842 4003 8845
rect 4015 8843 4023 8846
rect 3917 8828 3920 8833
rect 3942 8828 3945 8834
rect 3992 8836 3995 8842
rect 4015 8837 4018 8843
rect 4027 8838 4030 8841
rect 4038 8841 4041 8855
rect 4046 8841 4051 8846
rect 4038 8838 4046 8841
rect 3960 8828 3963 8833
rect 4038 8833 4041 8838
rect 3990 8827 3995 8832
rect 3309 8812 3318 8816
rect 3322 8812 3354 8816
rect 3358 8812 3421 8816
rect 3425 8812 3450 8816
rect 3454 8812 3486 8816
rect 3490 8812 3553 8816
rect 3557 8812 3582 8816
rect 3586 8812 3618 8816
rect 3622 8812 3685 8816
rect 3689 8812 3769 8816
rect 3862 8815 3863 8819
rect 3887 8816 3888 8820
rect 3934 8815 3935 8819
rect 3309 8805 3342 8809
rect 3346 8805 3370 8809
rect 3374 8805 3400 8809
rect 3404 8805 3437 8809
rect 3441 8805 3474 8809
rect 3478 8805 3502 8809
rect 3506 8805 3532 8809
rect 3536 8805 3569 8809
rect 3573 8805 3606 8809
rect 3610 8805 3634 8809
rect 3638 8805 3664 8809
rect 3668 8805 3701 8809
rect 3705 8805 3709 8809
rect 3794 8808 3815 8812
rect 3819 8808 3824 8812
rect 3828 8808 3874 8812
rect 3878 8808 3899 8812
rect 3903 8808 3930 8812
rect 3934 8808 3963 8812
rect 3999 8805 4002 8833
rect 4403 8832 4829 8928
rect 4029 8805 4032 8829
rect 4786 8822 4829 8832
rect 4796 8812 4829 8822
rect 343 8790 366 8800
rect 2367 8795 2370 8805
rect 2388 8795 2391 8805
rect 2404 8795 2407 8805
rect 2418 8798 2423 8802
rect 2427 8798 2434 8802
rect 2446 8795 2449 8805
rect 2462 8795 2465 8805
rect 2483 8795 2486 8805
rect 2499 8795 2502 8805
rect 2520 8795 2523 8805
rect 2536 8795 2539 8805
rect 2550 8798 2555 8802
rect 2559 8798 2566 8802
rect 2578 8795 2581 8805
rect 2594 8795 2597 8805
rect 2615 8795 2618 8805
rect 2631 8795 2634 8805
rect 2652 8795 2655 8805
rect 2668 8795 2671 8805
rect 2682 8798 2687 8802
rect 2691 8798 2698 8802
rect 2710 8795 2713 8805
rect 2726 8795 2729 8805
rect 2747 8795 2750 8805
rect 2782 8801 2856 8805
rect 2860 8801 2862 8805
rect 2866 8801 2870 8805
rect 2874 8801 2888 8805
rect 2892 8801 2897 8805
rect 2901 8801 2906 8805
rect 2910 8801 2929 8805
rect 2933 8801 2963 8805
rect 2967 8801 2978 8805
rect 2982 8801 3006 8805
rect 3010 8801 3023 8805
rect 3027 8801 3047 8805
rect 3051 8801 3131 8805
rect 3135 8801 3149 8805
rect 3153 8801 3158 8805
rect 3162 8801 3167 8805
rect 3171 8801 3190 8805
rect 3194 8801 3224 8805
rect 3228 8801 3239 8805
rect 3243 8801 3267 8805
rect 3271 8801 3280 8805
rect 343 8780 356 8790
rect 343 8741 346 8780
rect 2384 8781 2389 8784
rect 2393 8781 2417 8784
rect 2442 8781 2449 8784
rect 2453 8781 2475 8784
rect 2495 8781 2502 8784
rect 2516 8781 2521 8784
rect 2525 8781 2549 8784
rect 2574 8781 2581 8784
rect 2585 8781 2607 8784
rect 2627 8781 2634 8784
rect 2648 8781 2653 8784
rect 2657 8781 2681 8784
rect 2794 8794 2870 8798
rect 2874 8794 2879 8798
rect 2883 8794 2929 8798
rect 2933 8794 2954 8798
rect 2958 8794 2985 8798
rect 2989 8794 3018 8798
rect 2706 8781 2713 8784
rect 2717 8781 2739 8784
rect 2917 8787 2918 8791
rect 2942 8786 2943 8790
rect 2989 8787 2990 8791
rect 2400 8771 2407 8774
rect 2411 8775 2430 8778
rect 2430 8768 2433 8774
rect 2458 8771 2465 8774
rect 2469 8775 2484 8778
rect 2532 8771 2539 8774
rect 2543 8775 2562 8778
rect 2562 8768 2565 8774
rect 2590 8771 2597 8774
rect 2601 8775 2616 8778
rect 2664 8771 2671 8774
rect 2675 8775 2694 8778
rect 2694 8768 2697 8774
rect 2722 8771 2729 8774
rect 2733 8775 2750 8778
rect 2865 8773 2868 8778
rect 2872 8773 2875 8778
rect 2855 8770 2857 8773
rect 2865 8770 2875 8773
rect 2865 8764 2868 8770
rect 2367 8752 2370 8764
rect 2388 8752 2391 8764
rect 2404 8752 2407 8764
rect 2418 8755 2430 8758
rect 2446 8752 2449 8764
rect 2462 8752 2465 8764
rect 2483 8752 2486 8764
rect 2499 8752 2502 8764
rect 2520 8752 2523 8764
rect 2536 8752 2539 8764
rect 2550 8755 2562 8758
rect 2578 8752 2581 8764
rect 2594 8752 2597 8764
rect 2615 8752 2618 8764
rect 2631 8752 2634 8764
rect 2652 8752 2655 8764
rect 2668 8752 2671 8764
rect 2682 8755 2694 8758
rect 2710 8752 2713 8764
rect 2726 8752 2729 8764
rect 2747 8752 2750 8764
rect 2872 8764 2875 8770
rect 2881 8772 2884 8778
rect 2897 8773 2900 8778
rect 2881 8768 2883 8772
rect 2887 8768 2889 8772
rect 2897 8771 2903 8773
rect 2907 8771 2908 8773
rect 2897 8769 2908 8771
rect 2925 8771 2928 8778
rect 2881 8764 2884 8768
rect 2897 8764 2900 8769
rect 2926 8767 2928 8771
rect 2925 8764 2928 8767
rect 2941 8772 2944 8778
rect 2951 8772 2954 8778
rect 2972 8773 2975 8778
rect 2951 8768 2960 8772
rect 2972 8769 2973 8773
rect 2977 8770 2980 8773
rect 2997 8772 3000 8778
rect 3015 8773 3018 8778
rect 3054 8775 3057 8801
rect 3090 8794 3109 8798
rect 3113 8794 3131 8798
rect 3135 8794 3190 8798
rect 3194 8794 3215 8798
rect 3219 8794 3246 8798
rect 3250 8794 3279 8798
rect 3312 8795 3315 8805
rect 3333 8795 3336 8805
rect 3349 8795 3352 8805
rect 3363 8798 3368 8802
rect 3372 8798 3379 8802
rect 3391 8795 3394 8805
rect 3407 8795 3410 8805
rect 3428 8795 3431 8805
rect 3444 8795 3447 8805
rect 3465 8795 3468 8805
rect 3481 8795 3484 8805
rect 3495 8798 3500 8802
rect 3504 8798 3511 8802
rect 3523 8795 3526 8805
rect 3539 8795 3542 8805
rect 3560 8795 3563 8805
rect 3576 8795 3579 8805
rect 3597 8795 3600 8805
rect 3613 8795 3616 8805
rect 3627 8798 3632 8802
rect 3636 8798 3643 8802
rect 3655 8795 3658 8805
rect 3671 8795 3674 8805
rect 3692 8795 3695 8805
rect 3727 8801 3801 8805
rect 3805 8801 3807 8805
rect 3811 8801 3815 8805
rect 3819 8801 3833 8805
rect 3837 8801 3842 8805
rect 3846 8801 3851 8805
rect 3855 8801 3874 8805
rect 3878 8801 3908 8805
rect 3912 8801 3923 8805
rect 3927 8801 3951 8805
rect 3955 8801 3968 8805
rect 3972 8801 3992 8805
rect 3996 8801 4076 8805
rect 4080 8801 4094 8805
rect 4098 8801 4103 8805
rect 4107 8801 4112 8805
rect 4116 8801 4135 8805
rect 4139 8801 4169 8805
rect 4173 8801 4184 8805
rect 4188 8801 4212 8805
rect 4216 8801 4225 8805
rect 4806 8802 4829 8812
rect 3090 8782 3093 8794
rect 3178 8787 3179 8791
rect 3203 8786 3204 8790
rect 3250 8787 3251 8791
rect 2941 8764 2944 8768
rect 2951 8764 2954 8768
rect 2972 8764 2975 8769
rect 2999 8768 3000 8772
rect 3117 8773 3120 8778
rect 3126 8773 3129 8778
rect 3133 8773 3136 8778
rect 2997 8764 3000 8768
rect 3015 8764 3018 8769
rect 3044 8762 3049 8767
rect 3053 8763 3055 8766
rect 3070 8765 3073 8771
rect 3102 8770 3136 8773
rect 3070 8762 3078 8765
rect 3070 8759 3073 8762
rect 2364 8748 2397 8752
rect 2401 8748 2425 8752
rect 2429 8748 2455 8752
rect 2459 8748 2529 8752
rect 2533 8748 2557 8752
rect 2561 8748 2587 8752
rect 2591 8748 2661 8752
rect 2665 8748 2689 8752
rect 2693 8748 2719 8752
rect 2723 8748 2776 8752
rect 2925 8749 2928 8753
rect 2952 8749 2953 8753
rect 2997 8749 2999 8753
rect 3102 8756 3105 8770
rect 3126 8764 3129 8770
rect 3133 8764 3136 8770
rect 3142 8772 3145 8778
rect 3158 8773 3161 8778
rect 3142 8768 3144 8772
rect 3148 8768 3150 8772
rect 3158 8771 3164 8773
rect 3168 8771 3169 8773
rect 3158 8769 3169 8771
rect 3186 8771 3189 8778
rect 3142 8764 3145 8768
rect 3158 8764 3161 8769
rect 3187 8767 3189 8771
rect 3186 8764 3189 8767
rect 3329 8781 3334 8784
rect 3338 8781 3362 8784
rect 3387 8781 3394 8784
rect 3398 8781 3420 8784
rect 3440 8781 3447 8784
rect 3461 8781 3466 8784
rect 3470 8781 3494 8784
rect 3519 8781 3526 8784
rect 3530 8781 3552 8784
rect 3572 8781 3579 8784
rect 3593 8781 3598 8784
rect 3602 8781 3626 8784
rect 3739 8794 3815 8798
rect 3819 8794 3824 8798
rect 3828 8794 3874 8798
rect 3878 8794 3899 8798
rect 3903 8794 3930 8798
rect 3934 8794 3963 8798
rect 3651 8781 3658 8784
rect 3662 8781 3684 8784
rect 3862 8787 3863 8791
rect 3887 8786 3888 8790
rect 3934 8787 3935 8791
rect 3202 8772 3205 8778
rect 3212 8772 3215 8778
rect 3233 8773 3236 8778
rect 3212 8768 3221 8772
rect 3233 8769 3234 8773
rect 3238 8770 3241 8773
rect 3258 8772 3261 8778
rect 3276 8773 3279 8778
rect 3202 8764 3205 8768
rect 3212 8764 3215 8768
rect 3233 8764 3236 8769
rect 3260 8768 3261 8772
rect 3258 8764 3261 8768
rect 3276 8764 3279 8769
rect 3345 8771 3352 8774
rect 3356 8775 3375 8778
rect 3375 8768 3378 8774
rect 3403 8771 3410 8774
rect 3414 8775 3429 8778
rect 3477 8771 3484 8774
rect 3488 8775 3507 8778
rect 3507 8768 3510 8774
rect 3535 8771 3542 8774
rect 3546 8775 3561 8778
rect 3609 8771 3616 8774
rect 3620 8775 3639 8778
rect 3639 8768 3642 8774
rect 3667 8771 3674 8774
rect 3678 8775 3695 8778
rect 3810 8773 3813 8778
rect 3817 8773 3820 8778
rect 3800 8770 3802 8773
rect 3810 8770 3820 8773
rect 3810 8764 3813 8770
rect 2364 8741 2373 8745
rect 2377 8741 2424 8745
rect 2428 8741 2474 8745
rect 2478 8741 2505 8745
rect 2509 8741 2556 8745
rect 2560 8741 2606 8745
rect 2610 8741 2637 8745
rect 2641 8741 2688 8745
rect 2692 8741 2738 8745
rect 2742 8742 2812 8745
rect 2868 8742 2882 8746
rect 2886 8742 2913 8746
rect 2917 8742 2935 8746
rect 2939 8742 3000 8746
rect 3004 8742 3018 8746
rect 86 8738 346 8741
rect 3054 8739 3057 8751
rect 3186 8749 3189 8753
rect 3213 8749 3214 8753
rect 3258 8749 3260 8753
rect 3312 8752 3315 8764
rect 3333 8752 3336 8764
rect 3349 8752 3352 8764
rect 3363 8755 3375 8758
rect 3391 8752 3394 8764
rect 3407 8752 3410 8764
rect 3428 8752 3431 8764
rect 3444 8752 3447 8764
rect 3465 8752 3468 8764
rect 3481 8752 3484 8764
rect 3495 8755 3507 8758
rect 3523 8752 3526 8764
rect 3539 8752 3542 8764
rect 3560 8752 3563 8764
rect 3576 8752 3579 8764
rect 3597 8752 3600 8764
rect 3613 8752 3616 8764
rect 3627 8755 3639 8758
rect 3655 8752 3658 8764
rect 3671 8752 3674 8764
rect 3692 8752 3695 8764
rect 3817 8764 3820 8770
rect 3826 8772 3829 8778
rect 3842 8773 3845 8778
rect 3826 8768 3828 8772
rect 3832 8768 3834 8772
rect 3842 8771 3848 8773
rect 3852 8771 3853 8773
rect 3842 8769 3853 8771
rect 3870 8771 3873 8778
rect 3826 8764 3829 8768
rect 3842 8764 3845 8769
rect 3871 8767 3873 8771
rect 3870 8764 3873 8767
rect 3886 8772 3889 8778
rect 3896 8772 3899 8778
rect 3917 8773 3920 8778
rect 3896 8768 3905 8772
rect 3917 8769 3918 8773
rect 3922 8770 3925 8773
rect 3942 8772 3945 8778
rect 3960 8773 3963 8778
rect 3999 8775 4002 8801
rect 4035 8794 4054 8798
rect 4058 8794 4076 8798
rect 4080 8794 4135 8798
rect 4139 8794 4160 8798
rect 4164 8794 4191 8798
rect 4195 8794 4224 8798
rect 4035 8782 4038 8794
rect 4816 8792 4829 8802
rect 4123 8787 4124 8791
rect 4148 8786 4149 8790
rect 4195 8787 4196 8791
rect 3886 8764 3889 8768
rect 3896 8764 3899 8768
rect 3917 8764 3920 8769
rect 3944 8768 3945 8772
rect 4062 8773 4065 8778
rect 4071 8773 4074 8778
rect 4078 8773 4081 8778
rect 3942 8764 3945 8768
rect 3960 8764 3963 8769
rect 3989 8762 3994 8767
rect 3998 8763 4000 8766
rect 4015 8765 4018 8771
rect 4047 8770 4081 8773
rect 4015 8762 4023 8765
rect 4015 8759 4018 8762
rect 3309 8748 3342 8752
rect 3346 8748 3370 8752
rect 3374 8748 3400 8752
rect 3404 8748 3474 8752
rect 3478 8748 3502 8752
rect 3506 8748 3532 8752
rect 3536 8748 3606 8752
rect 3610 8748 3634 8752
rect 3638 8748 3664 8752
rect 3668 8748 3721 8752
rect 3870 8749 3873 8753
rect 3897 8749 3898 8753
rect 3942 8749 3944 8753
rect 4047 8756 4050 8770
rect 4071 8764 4074 8770
rect 4078 8764 4081 8770
rect 4087 8772 4090 8778
rect 4103 8773 4106 8778
rect 4087 8768 4089 8772
rect 4093 8768 4095 8772
rect 4103 8771 4109 8773
rect 4113 8771 4114 8773
rect 4103 8769 4114 8771
rect 4131 8771 4134 8778
rect 4087 8764 4090 8768
rect 4103 8764 4106 8769
rect 4132 8767 4134 8771
rect 4131 8764 4134 8767
rect 4147 8772 4150 8778
rect 4157 8772 4160 8778
rect 4178 8773 4181 8778
rect 4157 8768 4166 8772
rect 4178 8769 4179 8773
rect 4183 8770 4186 8773
rect 4203 8772 4206 8778
rect 4221 8773 4224 8778
rect 4147 8764 4150 8768
rect 4157 8764 4160 8768
rect 4178 8764 4181 8769
rect 4205 8768 4206 8772
rect 4203 8764 4206 8768
rect 4221 8764 4224 8769
rect 3094 8742 3099 8746
rect 3103 8742 3143 8746
rect 3147 8742 3174 8746
rect 3178 8742 3196 8746
rect 3200 8742 3261 8746
rect 3265 8742 3279 8746
rect 3309 8741 3318 8745
rect 3322 8741 3369 8745
rect 3373 8741 3419 8745
rect 3423 8741 3450 8745
rect 3454 8741 3501 8745
rect 3505 8741 3551 8745
rect 3555 8741 3582 8745
rect 3586 8741 3633 8745
rect 3637 8741 3683 8745
rect 3687 8742 3757 8745
rect 3813 8742 3827 8746
rect 3831 8742 3858 8746
rect 3862 8742 3880 8746
rect 3884 8742 3945 8746
rect 3949 8742 3963 8746
rect 3999 8739 4002 8751
rect 4131 8749 4134 8753
rect 4158 8749 4159 8753
rect 4203 8749 4205 8753
rect 4826 8753 4829 8792
rect 5083 8753 5086 9007
rect 4483 8747 4484 8751
rect 4488 8747 4489 8751
rect 4493 8747 4494 8751
rect 4498 8747 4499 8751
rect 4503 8747 4504 8751
rect 4508 8747 4509 8751
rect 4479 8746 4513 8747
rect 4039 8742 4044 8746
rect 4048 8742 4088 8746
rect 4092 8742 4119 8746
rect 4123 8742 4141 8746
rect 4145 8742 4206 8746
rect 4210 8742 4224 8746
rect 4483 8742 4484 8746
rect 4488 8742 4489 8746
rect 4493 8742 4494 8746
rect 4498 8742 4499 8746
rect 4503 8742 4504 8746
rect 4508 8742 4509 8746
rect 4479 8741 4513 8742
rect 2371 8735 2755 8738
rect 2770 8735 2855 8739
rect 2859 8735 2871 8739
rect 2875 8735 2889 8739
rect 2893 8735 2900 8739
rect 2904 8735 2906 8739
rect 2910 8735 2925 8739
rect 2929 8735 2962 8739
rect 2966 8735 2967 8739
rect 2971 8735 2979 8739
rect 2983 8735 3007 8739
rect 3011 8735 3047 8739
rect 3051 8735 3090 8739
rect 3094 8735 3101 8739
rect 3105 8735 3116 8739
rect 3120 8735 3132 8739
rect 3136 8735 3150 8739
rect 3154 8735 3161 8739
rect 3165 8735 3167 8739
rect 3171 8735 3186 8739
rect 3190 8735 3223 8739
rect 3227 8735 3228 8739
rect 3232 8735 3240 8739
rect 3244 8735 3268 8739
rect 3272 8735 3280 8739
rect 3316 8735 3700 8738
rect 3715 8735 3800 8739
rect 3804 8735 3816 8739
rect 3820 8735 3834 8739
rect 3838 8735 3845 8739
rect 3849 8735 3851 8739
rect 3855 8735 3870 8739
rect 3874 8735 3907 8739
rect 3911 8735 3912 8739
rect 3916 8735 3924 8739
rect 3928 8735 3952 8739
rect 3956 8735 3992 8739
rect 3996 8735 4035 8739
rect 4039 8735 4046 8739
rect 4050 8735 4061 8739
rect 4065 8735 4077 8739
rect 4081 8735 4095 8739
rect 4099 8735 4106 8739
rect 4110 8735 4112 8739
rect 4116 8735 4131 8739
rect 4135 8735 4168 8739
rect 4172 8735 4173 8739
rect 4177 8735 4185 8739
rect 4189 8735 4213 8739
rect 4217 8735 4225 8739
rect 4483 8737 4484 8741
rect 4488 8737 4489 8741
rect 4493 8737 4494 8741
rect 4498 8737 4499 8741
rect 4503 8737 4504 8741
rect 4508 8737 4509 8741
rect 4479 8736 4513 8737
rect 2514 8728 2623 8731
rect 2806 8728 2864 8732
rect 2868 8728 3098 8731
rect 3288 8729 3296 8733
rect 3459 8728 3568 8731
rect 3751 8728 3809 8732
rect 3813 8728 4043 8731
rect 4233 8729 4241 8733
rect 4483 8732 4484 8736
rect 4488 8732 4489 8736
rect 4493 8732 4494 8736
rect 4498 8732 4499 8736
rect 4503 8732 4504 8736
rect 4508 8732 4509 8736
rect 4529 8747 4530 8751
rect 4534 8747 4535 8751
rect 4539 8747 4540 8751
rect 4544 8747 4545 8751
rect 4549 8747 4550 8751
rect 4554 8747 4555 8751
rect 4826 8750 5086 8753
rect 4525 8746 4559 8747
rect 4529 8742 4530 8746
rect 4534 8742 4535 8746
rect 4539 8742 4540 8746
rect 4544 8742 4545 8746
rect 4549 8742 4550 8746
rect 4554 8742 4555 8746
rect 4525 8741 4559 8742
rect 4529 8737 4530 8741
rect 4534 8737 4535 8741
rect 4539 8737 4540 8741
rect 4544 8737 4545 8741
rect 4549 8737 4550 8741
rect 4554 8737 4555 8741
rect 4525 8736 4559 8737
rect 4529 8732 4530 8736
rect 4534 8732 4535 8736
rect 4539 8732 4540 8736
rect 4544 8732 4545 8736
rect 4549 8732 4550 8736
rect 4554 8732 4555 8736
rect 2494 8720 2498 8724
rect 2502 8720 2506 8724
rect 2794 8721 3108 8724
rect 2482 8719 2486 8720
rect 2514 8719 2518 8720
rect 2842 8714 3115 8717
rect 3284 8711 3288 8716
rect 3439 8720 3443 8724
rect 3447 8720 3451 8724
rect 3739 8721 4053 8724
rect 3427 8719 3431 8720
rect 3459 8719 3463 8720
rect 3787 8714 4058 8718
rect 4229 8711 4233 8716
rect 2355 8707 2482 8711
rect 2486 8707 2502 8711
rect 2518 8707 3427 8711
rect 3431 8707 3447 8711
rect 3463 8707 4321 8711
rect 617 8703 618 8707
rect 622 8703 623 8707
rect 627 8703 628 8707
rect 632 8703 633 8707
rect 637 8703 638 8707
rect 642 8703 643 8707
rect 613 8702 647 8703
rect 617 8698 618 8702
rect 622 8698 623 8702
rect 627 8698 628 8702
rect 632 8698 633 8702
rect 637 8698 638 8702
rect 642 8698 643 8702
rect 613 8697 647 8698
rect 617 8693 618 8697
rect 622 8693 623 8697
rect 627 8693 628 8697
rect 632 8693 633 8697
rect 637 8693 638 8697
rect 642 8693 643 8697
rect 613 8692 647 8693
rect 86 8686 346 8689
rect 617 8688 618 8692
rect 622 8688 623 8692
rect 627 8688 628 8692
rect 632 8688 633 8692
rect 637 8688 638 8692
rect 642 8688 643 8692
rect 663 8703 664 8707
rect 668 8703 669 8707
rect 673 8703 674 8707
rect 678 8703 679 8707
rect 683 8703 684 8707
rect 688 8703 689 8707
rect 659 8702 693 8703
rect 663 8698 664 8702
rect 668 8698 669 8702
rect 673 8698 674 8702
rect 678 8698 679 8702
rect 683 8698 684 8702
rect 688 8698 689 8702
rect 659 8697 693 8698
rect 663 8693 664 8697
rect 668 8693 669 8697
rect 673 8693 674 8697
rect 678 8693 679 8697
rect 683 8693 684 8697
rect 688 8693 689 8697
rect 2510 8700 2755 8703
rect 2830 8700 3156 8704
rect 3160 8700 3192 8704
rect 3196 8700 3259 8704
rect 3263 8700 3279 8704
rect 3455 8700 3700 8703
rect 3775 8700 4101 8704
rect 4105 8700 4137 8704
rect 4141 8700 4204 8704
rect 4208 8700 4224 8704
rect 659 8692 693 8693
rect 2525 8693 2755 8696
rect 2770 8693 3142 8697
rect 3146 8693 3180 8697
rect 3184 8693 3208 8697
rect 3212 8693 3238 8697
rect 3242 8693 3275 8697
rect 4826 8698 5086 8701
rect 663 8688 664 8692
rect 668 8688 669 8692
rect 673 8688 674 8692
rect 678 8688 679 8692
rect 683 8688 684 8692
rect 688 8688 689 8692
rect 86 8432 89 8686
rect 343 8647 346 8686
rect 2494 8684 2498 8688
rect 2502 8684 2506 8688
rect 3150 8683 3153 8693
rect 3171 8683 3174 8693
rect 3187 8683 3190 8693
rect 3201 8686 3206 8690
rect 3210 8686 3217 8690
rect 3229 8683 3232 8693
rect 3245 8683 3248 8693
rect 3266 8683 3269 8693
rect 3470 8693 3700 8696
rect 3715 8693 4087 8697
rect 4091 8693 4125 8697
rect 4129 8693 4153 8697
rect 4157 8693 4183 8697
rect 4187 8693 4220 8697
rect 3439 8684 3443 8688
rect 3447 8684 3451 8688
rect 4095 8683 4098 8693
rect 4116 8683 4119 8693
rect 4132 8683 4135 8693
rect 4146 8686 4151 8690
rect 4155 8686 4162 8690
rect 4174 8683 4177 8693
rect 4190 8683 4193 8693
rect 4211 8683 4214 8693
rect 2514 8677 2624 8680
rect 2364 8670 2373 8674
rect 2377 8670 2409 8674
rect 2413 8670 2476 8674
rect 2480 8670 2505 8674
rect 2509 8670 2541 8674
rect 2545 8670 2608 8674
rect 2612 8670 2637 8674
rect 2641 8670 2673 8674
rect 2677 8670 2740 8674
rect 2744 8670 2824 8674
rect 2364 8663 2397 8667
rect 2401 8663 2425 8667
rect 2429 8663 2455 8667
rect 2459 8663 2492 8667
rect 2496 8663 2529 8667
rect 2533 8663 2557 8667
rect 2561 8663 2587 8667
rect 2591 8663 2624 8667
rect 2628 8663 2661 8667
rect 2665 8663 2689 8667
rect 2693 8663 2719 8667
rect 2723 8663 2756 8667
rect 2760 8663 2764 8667
rect 3167 8669 3172 8672
rect 3176 8669 3200 8672
rect 3459 8677 3569 8680
rect 3225 8669 3232 8672
rect 3236 8669 3258 8672
rect 3309 8670 3318 8674
rect 3322 8670 3354 8674
rect 3358 8670 3421 8674
rect 3425 8670 3450 8674
rect 3454 8670 3486 8674
rect 3490 8670 3553 8674
rect 3557 8670 3582 8674
rect 3586 8670 3618 8674
rect 3622 8670 3685 8674
rect 3689 8670 3769 8674
rect 2367 8653 2370 8663
rect 2388 8653 2391 8663
rect 2404 8653 2407 8663
rect 2418 8656 2423 8660
rect 2427 8656 2434 8660
rect 2446 8653 2449 8663
rect 2462 8653 2465 8663
rect 2483 8653 2486 8663
rect 2499 8653 2502 8663
rect 2520 8653 2523 8663
rect 2536 8653 2539 8663
rect 2550 8656 2555 8660
rect 2559 8656 2566 8660
rect 2578 8653 2581 8663
rect 2594 8653 2597 8663
rect 2615 8653 2618 8663
rect 2631 8653 2634 8663
rect 2652 8653 2655 8663
rect 2668 8653 2671 8663
rect 2682 8656 2687 8660
rect 2691 8656 2698 8660
rect 2710 8653 2713 8663
rect 2726 8653 2729 8663
rect 2747 8653 2750 8663
rect 3183 8659 3190 8662
rect 3194 8663 3213 8666
rect 343 8637 356 8647
rect 343 8627 366 8637
rect 2384 8639 2389 8642
rect 2393 8639 2417 8642
rect 2442 8639 2449 8642
rect 2453 8639 2475 8642
rect 2495 8639 2502 8642
rect 2516 8639 2521 8642
rect 2525 8639 2549 8642
rect 2574 8639 2581 8642
rect 2585 8639 2607 8642
rect 2627 8639 2634 8642
rect 2648 8639 2653 8642
rect 2657 8639 2681 8642
rect 2706 8639 2713 8642
rect 2717 8639 2739 8642
rect 3213 8656 3216 8662
rect 3241 8659 3248 8662
rect 3252 8663 3267 8666
rect 3309 8663 3342 8667
rect 3346 8663 3370 8667
rect 3374 8663 3400 8667
rect 3404 8663 3437 8667
rect 3441 8663 3474 8667
rect 3478 8663 3502 8667
rect 3506 8663 3532 8667
rect 3536 8663 3569 8667
rect 3573 8663 3606 8667
rect 3610 8663 3634 8667
rect 3638 8663 3664 8667
rect 3668 8663 3701 8667
rect 3705 8663 3709 8667
rect 4112 8669 4117 8672
rect 4121 8669 4145 8672
rect 4170 8669 4177 8672
rect 4181 8669 4203 8672
rect 3312 8653 3315 8663
rect 3333 8653 3336 8663
rect 3349 8653 3352 8663
rect 3363 8656 3368 8660
rect 3372 8656 3379 8660
rect 3391 8653 3394 8663
rect 3407 8653 3410 8663
rect 3428 8653 3431 8663
rect 3444 8653 3447 8663
rect 3465 8653 3468 8663
rect 3481 8653 3484 8663
rect 3495 8656 3500 8660
rect 3504 8656 3511 8660
rect 3523 8653 3526 8663
rect 3539 8653 3542 8663
rect 3560 8653 3563 8663
rect 3576 8653 3579 8663
rect 3597 8653 3600 8663
rect 3613 8653 3616 8663
rect 3627 8656 3632 8660
rect 3636 8656 3643 8660
rect 3655 8653 3658 8663
rect 3671 8653 3674 8663
rect 3692 8653 3695 8663
rect 4128 8659 4135 8662
rect 4139 8663 4158 8666
rect 3150 8640 3153 8652
rect 3171 8640 3174 8652
rect 3187 8640 3190 8652
rect 3201 8643 3213 8646
rect 3229 8640 3232 8652
rect 3245 8640 3248 8652
rect 3266 8640 3269 8652
rect 343 8617 376 8627
rect 2400 8629 2407 8632
rect 2411 8633 2430 8636
rect 2430 8626 2433 8632
rect 2458 8629 2465 8632
rect 2469 8633 2484 8636
rect 2532 8629 2539 8632
rect 2543 8633 2562 8636
rect 2562 8626 2565 8632
rect 2590 8629 2597 8632
rect 2601 8633 2616 8636
rect 2664 8629 2671 8632
rect 2675 8633 2694 8636
rect 2694 8626 2697 8632
rect 2722 8629 2729 8632
rect 2733 8633 2750 8636
rect 2782 8636 3180 8640
rect 3184 8636 3208 8640
rect 3212 8636 3238 8640
rect 3242 8636 3279 8640
rect 3329 8639 3334 8642
rect 3338 8639 3362 8642
rect 3387 8639 3394 8642
rect 3398 8639 3420 8642
rect 3440 8639 3447 8642
rect 3461 8639 3466 8642
rect 3470 8639 3494 8642
rect 3519 8639 3526 8642
rect 3530 8639 3552 8642
rect 3572 8639 3579 8642
rect 3593 8639 3598 8642
rect 3602 8639 3626 8642
rect 3651 8639 3658 8642
rect 3662 8639 3684 8642
rect 4158 8656 4161 8662
rect 4186 8659 4193 8662
rect 4197 8663 4212 8666
rect 4826 8659 4829 8698
rect 4095 8640 4098 8652
rect 4116 8640 4119 8652
rect 4132 8640 4135 8652
rect 4146 8643 4158 8646
rect 4174 8640 4177 8652
rect 4190 8640 4193 8652
rect 4211 8640 4214 8652
rect 4816 8649 4829 8659
rect 2818 8629 3156 8633
rect 3160 8629 3207 8633
rect 3211 8629 3257 8633
rect 3261 8629 3279 8633
rect 3345 8629 3352 8632
rect 3356 8633 3375 8636
rect 343 8607 386 8617
rect 2367 8610 2370 8622
rect 2388 8610 2391 8622
rect 2404 8610 2407 8622
rect 2418 8613 2430 8616
rect 2446 8610 2449 8622
rect 2462 8610 2465 8622
rect 2483 8610 2486 8622
rect 2499 8610 2502 8622
rect 2520 8610 2523 8622
rect 2536 8610 2539 8622
rect 2550 8613 2562 8616
rect 2578 8610 2581 8622
rect 2594 8610 2597 8622
rect 2615 8610 2618 8622
rect 2631 8610 2634 8622
rect 2652 8610 2655 8622
rect 2668 8610 2671 8622
rect 2682 8613 2694 8616
rect 2710 8610 2713 8622
rect 2726 8610 2729 8622
rect 2747 8610 2750 8622
rect 3153 8622 3274 8625
rect 3375 8626 3378 8632
rect 3403 8629 3410 8632
rect 3414 8633 3429 8636
rect 3477 8629 3484 8632
rect 3488 8633 3507 8636
rect 3507 8626 3510 8632
rect 3535 8629 3542 8632
rect 3546 8633 3561 8636
rect 3609 8629 3616 8632
rect 3620 8633 3639 8636
rect 3639 8626 3642 8632
rect 3667 8629 3674 8632
rect 3678 8633 3695 8636
rect 3727 8636 4125 8640
rect 4129 8636 4153 8640
rect 4157 8636 4183 8640
rect 4187 8636 4224 8640
rect 4806 8639 4829 8649
rect 3763 8629 4101 8633
rect 4105 8629 4152 8633
rect 4156 8629 4202 8633
rect 4206 8629 4224 8633
rect 4796 8629 4829 8639
rect 2830 8614 3156 8618
rect 3160 8614 3192 8618
rect 3196 8614 3259 8618
rect 3263 8614 3279 8618
rect 343 8511 769 8607
rect 2364 8606 2397 8610
rect 2401 8606 2425 8610
rect 2429 8606 2455 8610
rect 2459 8606 2529 8610
rect 2533 8606 2557 8610
rect 2561 8606 2587 8610
rect 2591 8606 2661 8610
rect 2665 8606 2689 8610
rect 2693 8606 2719 8610
rect 2723 8606 2776 8610
rect 3146 8607 3180 8611
rect 3184 8607 3208 8611
rect 3212 8607 3238 8611
rect 3242 8607 3275 8611
rect 3312 8610 3315 8622
rect 3333 8610 3336 8622
rect 3349 8610 3352 8622
rect 3363 8613 3375 8616
rect 3391 8610 3394 8622
rect 3407 8610 3410 8622
rect 3428 8610 3431 8622
rect 3444 8610 3447 8622
rect 3465 8610 3468 8622
rect 3481 8610 3484 8622
rect 3495 8613 3507 8616
rect 3523 8610 3526 8622
rect 3539 8610 3542 8622
rect 3560 8610 3563 8622
rect 3576 8610 3579 8622
rect 3597 8610 3600 8622
rect 3613 8610 3616 8622
rect 3627 8613 3639 8616
rect 3655 8610 3658 8622
rect 3671 8610 3674 8622
rect 3692 8610 3695 8622
rect 4098 8622 4219 8625
rect 4786 8619 4829 8629
rect 3775 8614 4101 8618
rect 4105 8614 4137 8618
rect 4141 8614 4204 8618
rect 4208 8614 4224 8618
rect 2364 8599 2373 8603
rect 2377 8599 2424 8603
rect 2428 8599 2474 8603
rect 2478 8599 2505 8603
rect 2509 8599 2556 8603
rect 2560 8599 2606 8603
rect 2610 8599 2637 8603
rect 2641 8599 2688 8603
rect 2692 8599 2738 8603
rect 2742 8599 2812 8603
rect 3150 8597 3153 8607
rect 3171 8597 3174 8607
rect 3187 8597 3190 8607
rect 3201 8600 3206 8604
rect 3210 8600 3217 8604
rect 3229 8597 3232 8607
rect 3245 8597 3248 8607
rect 3266 8597 3269 8607
rect 3309 8606 3342 8610
rect 3346 8606 3370 8610
rect 3374 8606 3400 8610
rect 3404 8606 3474 8610
rect 3478 8606 3502 8610
rect 3506 8606 3532 8610
rect 3536 8606 3606 8610
rect 3610 8606 3634 8610
rect 3638 8606 3664 8610
rect 3668 8606 3721 8610
rect 4091 8607 4125 8611
rect 4129 8607 4153 8611
rect 4157 8607 4183 8611
rect 4187 8607 4220 8611
rect 3309 8599 3318 8603
rect 3322 8599 3369 8603
rect 3373 8599 3419 8603
rect 3423 8599 3450 8603
rect 3454 8599 3501 8603
rect 3505 8599 3551 8603
rect 3555 8599 3582 8603
rect 3586 8599 3633 8603
rect 3637 8599 3683 8603
rect 3687 8599 3757 8603
rect 4095 8597 4098 8607
rect 4116 8597 4119 8607
rect 4132 8597 4135 8607
rect 4146 8600 4151 8604
rect 4155 8600 4162 8604
rect 4174 8597 4177 8607
rect 4190 8597 4193 8607
rect 4211 8597 4214 8607
rect 2370 8592 2755 8595
rect 2364 8584 2373 8588
rect 2377 8584 2409 8588
rect 2413 8584 2476 8588
rect 2480 8584 2505 8588
rect 2509 8584 2541 8588
rect 2545 8584 2608 8588
rect 2612 8584 2637 8588
rect 2641 8584 2673 8588
rect 2677 8584 2740 8588
rect 2744 8584 2824 8588
rect 2364 8577 2397 8581
rect 2401 8577 2425 8581
rect 2429 8577 2455 8581
rect 2459 8577 2492 8581
rect 2496 8577 2529 8581
rect 2533 8577 2557 8581
rect 2561 8577 2587 8581
rect 2591 8577 2624 8581
rect 2628 8577 2661 8581
rect 2665 8577 2689 8581
rect 2693 8577 2719 8581
rect 2723 8577 2756 8581
rect 2760 8577 2764 8581
rect 3167 8583 3172 8586
rect 3176 8583 3200 8586
rect 3315 8592 3700 8595
rect 3225 8583 3232 8586
rect 3236 8583 3258 8586
rect 3309 8584 3318 8588
rect 3322 8584 3354 8588
rect 3358 8584 3421 8588
rect 3425 8584 3450 8588
rect 3454 8584 3486 8588
rect 3490 8584 3553 8588
rect 3557 8584 3582 8588
rect 3586 8584 3618 8588
rect 3622 8584 3685 8588
rect 3689 8584 3769 8588
rect 2367 8567 2370 8577
rect 2388 8567 2391 8577
rect 2404 8567 2407 8577
rect 2418 8570 2423 8574
rect 2427 8570 2434 8574
rect 2446 8567 2449 8577
rect 2462 8567 2465 8577
rect 2483 8567 2486 8577
rect 2499 8567 2502 8577
rect 2520 8567 2523 8577
rect 2536 8567 2539 8577
rect 2550 8570 2555 8574
rect 2559 8570 2566 8574
rect 2578 8567 2581 8577
rect 2594 8567 2597 8577
rect 2615 8567 2618 8577
rect 2631 8567 2634 8577
rect 2652 8567 2655 8577
rect 2668 8567 2671 8577
rect 2682 8570 2687 8574
rect 2691 8570 2698 8574
rect 2710 8567 2713 8577
rect 2726 8567 2729 8577
rect 2747 8567 2750 8577
rect 3183 8573 3190 8576
rect 3194 8577 3213 8580
rect 2384 8553 2389 8556
rect 2393 8553 2417 8556
rect 2442 8553 2449 8556
rect 2453 8553 2475 8556
rect 2495 8553 2502 8556
rect 2516 8553 2521 8556
rect 2525 8553 2549 8556
rect 2574 8553 2581 8556
rect 2585 8553 2607 8556
rect 2627 8553 2634 8556
rect 2648 8553 2653 8556
rect 2657 8553 2681 8556
rect 2706 8553 2713 8556
rect 2717 8553 2739 8556
rect 3213 8570 3216 8576
rect 3241 8573 3248 8576
rect 3252 8577 3267 8580
rect 3278 8575 3289 8579
rect 3309 8577 3342 8581
rect 3346 8577 3370 8581
rect 3374 8577 3400 8581
rect 3404 8577 3437 8581
rect 3441 8577 3474 8581
rect 3478 8577 3502 8581
rect 3506 8577 3532 8581
rect 3536 8577 3569 8581
rect 3573 8577 3606 8581
rect 3610 8577 3634 8581
rect 3638 8577 3664 8581
rect 3668 8577 3701 8581
rect 3705 8577 3709 8581
rect 4112 8583 4117 8586
rect 4121 8583 4145 8586
rect 4170 8583 4177 8586
rect 4181 8583 4203 8586
rect 3312 8567 3315 8577
rect 3333 8567 3336 8577
rect 3349 8567 3352 8577
rect 3363 8570 3368 8574
rect 3372 8570 3379 8574
rect 3391 8567 3394 8577
rect 3407 8567 3410 8577
rect 3428 8567 3431 8577
rect 3444 8567 3447 8577
rect 3465 8567 3468 8577
rect 3481 8567 3484 8577
rect 3495 8570 3500 8574
rect 3504 8570 3511 8574
rect 3523 8567 3526 8577
rect 3539 8567 3542 8577
rect 3560 8567 3563 8577
rect 3576 8567 3579 8577
rect 3597 8567 3600 8577
rect 3613 8567 3616 8577
rect 3627 8570 3632 8574
rect 3636 8570 3643 8574
rect 3655 8567 3658 8577
rect 3671 8567 3674 8577
rect 3692 8567 3695 8577
rect 4128 8573 4135 8576
rect 4139 8577 4158 8580
rect 3150 8554 3153 8566
rect 3171 8554 3174 8566
rect 3187 8554 3190 8566
rect 3201 8557 3213 8560
rect 3229 8554 3232 8566
rect 3245 8554 3248 8566
rect 3266 8554 3269 8566
rect 2400 8543 2407 8546
rect 2411 8547 2430 8550
rect 2430 8540 2433 8546
rect 2458 8543 2465 8546
rect 2469 8547 2484 8550
rect 2532 8543 2539 8546
rect 2543 8547 2562 8550
rect 2562 8540 2565 8546
rect 2590 8543 2597 8546
rect 2601 8547 2616 8550
rect 2664 8543 2671 8546
rect 2675 8547 2694 8550
rect 2694 8540 2697 8546
rect 2722 8543 2729 8546
rect 2733 8547 2750 8550
rect 2782 8550 3180 8554
rect 3184 8550 3208 8554
rect 3212 8550 3238 8554
rect 3242 8550 3279 8554
rect 3329 8553 3334 8556
rect 3338 8553 3362 8556
rect 3387 8553 3394 8556
rect 3398 8553 3420 8556
rect 3440 8553 3447 8556
rect 3461 8553 3466 8556
rect 3470 8553 3494 8556
rect 3519 8553 3526 8556
rect 3530 8553 3552 8556
rect 3572 8553 3579 8556
rect 3593 8553 3598 8556
rect 3602 8553 3626 8556
rect 3651 8553 3658 8556
rect 3662 8553 3684 8556
rect 4158 8570 4161 8576
rect 4186 8573 4193 8576
rect 4197 8577 4212 8580
rect 4223 8575 4234 8579
rect 4095 8554 4098 8566
rect 4116 8554 4119 8566
rect 4132 8554 4135 8566
rect 4146 8557 4158 8560
rect 4174 8554 4177 8566
rect 4190 8554 4193 8566
rect 4211 8554 4214 8566
rect 2818 8543 3156 8547
rect 3160 8543 3207 8547
rect 3211 8543 3257 8547
rect 3261 8543 3279 8547
rect 3345 8543 3352 8546
rect 3356 8547 3375 8550
rect 3375 8540 3378 8546
rect 3403 8543 3410 8546
rect 3414 8547 3429 8550
rect 3477 8543 3484 8546
rect 3488 8547 3507 8550
rect 3507 8540 3510 8546
rect 3535 8543 3542 8546
rect 3546 8547 3561 8550
rect 3609 8543 3616 8546
rect 3620 8547 3639 8550
rect 3639 8540 3642 8546
rect 3667 8543 3674 8546
rect 3678 8547 3695 8550
rect 3727 8550 4125 8554
rect 4129 8550 4153 8554
rect 4157 8550 4183 8554
rect 4187 8550 4224 8554
rect 3763 8543 4101 8547
rect 4105 8543 4152 8547
rect 4156 8543 4202 8547
rect 4206 8543 4224 8547
rect 2367 8524 2370 8536
rect 2388 8524 2391 8536
rect 2404 8524 2407 8536
rect 2418 8527 2430 8530
rect 2446 8524 2449 8536
rect 2462 8524 2465 8536
rect 2483 8524 2486 8536
rect 2499 8524 2502 8536
rect 2520 8524 2523 8536
rect 2536 8524 2539 8536
rect 2550 8527 2562 8530
rect 2578 8524 2581 8536
rect 2594 8524 2597 8536
rect 2615 8524 2618 8536
rect 2631 8524 2634 8536
rect 2652 8524 2655 8536
rect 2668 8524 2671 8536
rect 2682 8527 2694 8530
rect 2710 8524 2713 8536
rect 2726 8524 2729 8536
rect 2747 8524 2750 8536
rect 3312 8524 3315 8536
rect 3333 8524 3336 8536
rect 3349 8524 3352 8536
rect 3363 8527 3375 8530
rect 3391 8524 3394 8536
rect 3407 8524 3410 8536
rect 3428 8524 3431 8536
rect 3444 8524 3447 8536
rect 3465 8524 3468 8536
rect 3481 8524 3484 8536
rect 3495 8527 3507 8530
rect 3523 8524 3526 8536
rect 3539 8524 3542 8536
rect 3560 8524 3563 8536
rect 3576 8524 3579 8536
rect 3597 8524 3600 8536
rect 3613 8524 3616 8536
rect 3627 8527 3639 8530
rect 3655 8524 3658 8536
rect 3671 8524 3674 8536
rect 3692 8524 3695 8536
rect 2364 8520 2397 8524
rect 2401 8520 2425 8524
rect 2429 8520 2455 8524
rect 2459 8520 2529 8524
rect 2533 8520 2557 8524
rect 2561 8520 2587 8524
rect 2591 8520 2661 8524
rect 2665 8520 2689 8524
rect 2693 8520 2719 8524
rect 2723 8520 2776 8524
rect 3309 8520 3342 8524
rect 3346 8520 3370 8524
rect 3374 8520 3400 8524
rect 3404 8520 3474 8524
rect 3478 8520 3502 8524
rect 3506 8520 3532 8524
rect 3536 8520 3606 8524
rect 3610 8520 3634 8524
rect 3638 8520 3664 8524
rect 3668 8520 3721 8524
rect 4403 8523 4829 8619
rect 2364 8513 2373 8517
rect 2377 8513 2424 8517
rect 2428 8513 2474 8517
rect 2478 8513 2505 8517
rect 2509 8513 2556 8517
rect 2560 8513 2606 8517
rect 2610 8513 2637 8517
rect 2641 8513 2688 8517
rect 2692 8513 2738 8517
rect 2742 8513 2812 8517
rect 3309 8513 3318 8517
rect 3322 8513 3369 8517
rect 3373 8513 3419 8517
rect 3423 8513 3450 8517
rect 3454 8513 3501 8517
rect 3505 8513 3551 8517
rect 3555 8513 3582 8517
rect 3586 8513 3633 8517
rect 3637 8513 3683 8517
rect 3687 8513 3757 8517
rect 4786 8513 4829 8523
rect 343 8501 386 8511
rect 2370 8507 2755 8510
rect 3315 8507 3700 8510
rect 4796 8503 4829 8513
rect 343 8491 376 8501
rect 2495 8500 2599 8503
rect 3440 8500 3544 8503
rect 2611 8492 2615 8496
rect 2619 8492 2623 8496
rect 343 8481 366 8491
rect 3556 8492 3560 8496
rect 3564 8492 3568 8496
rect 4806 8493 4829 8503
rect 2354 8481 2599 8485
rect 2603 8481 2619 8485
rect 2635 8481 3296 8485
rect 3300 8481 3544 8485
rect 3548 8481 3564 8485
rect 3580 8481 4241 8485
rect 4245 8481 4323 8485
rect 4816 8483 4829 8493
rect 343 8471 356 8481
rect 2627 8474 2755 8477
rect 3572 8474 3700 8477
rect 343 8432 346 8471
rect 2642 8467 2755 8470
rect 3587 8467 3700 8470
rect 2611 8458 2615 8462
rect 2619 8458 2623 8462
rect 3556 8458 3560 8462
rect 3564 8458 3568 8462
rect 2495 8451 2599 8454
rect 3440 8451 3544 8454
rect 2364 8444 2373 8448
rect 2377 8444 2409 8448
rect 2413 8444 2476 8448
rect 2480 8444 2505 8448
rect 2509 8444 2541 8448
rect 2545 8444 2608 8448
rect 2612 8444 2637 8448
rect 2641 8444 2673 8448
rect 2677 8444 2740 8448
rect 2744 8444 2824 8448
rect 3309 8444 3318 8448
rect 3322 8444 3354 8448
rect 3358 8444 3421 8448
rect 3425 8444 3450 8448
rect 3454 8444 3486 8448
rect 3490 8444 3553 8448
rect 3557 8444 3582 8448
rect 3586 8444 3618 8448
rect 3622 8444 3685 8448
rect 3689 8444 3769 8448
rect 4826 8444 4829 8483
rect 5083 8444 5086 8698
rect 2364 8437 2397 8441
rect 2401 8437 2425 8441
rect 2429 8437 2455 8441
rect 2459 8437 2492 8441
rect 2496 8437 2529 8441
rect 2533 8437 2557 8441
rect 2561 8437 2587 8441
rect 2591 8437 2624 8441
rect 2628 8437 2661 8441
rect 2665 8437 2689 8441
rect 2693 8437 2719 8441
rect 2723 8437 2756 8441
rect 2760 8437 2764 8441
rect 3309 8437 3342 8441
rect 3346 8437 3370 8441
rect 3374 8437 3400 8441
rect 3404 8437 3437 8441
rect 3441 8437 3474 8441
rect 3478 8437 3502 8441
rect 3506 8437 3532 8441
rect 3536 8437 3569 8441
rect 3573 8437 3606 8441
rect 3610 8437 3634 8441
rect 3638 8437 3664 8441
rect 3668 8437 3701 8441
rect 3705 8437 3709 8441
rect 4483 8438 4484 8442
rect 4488 8438 4489 8442
rect 4493 8438 4494 8442
rect 4498 8438 4499 8442
rect 4503 8438 4504 8442
rect 4508 8438 4509 8442
rect 4479 8437 4513 8438
rect 86 8429 346 8432
rect 2367 8427 2370 8437
rect 2388 8427 2391 8437
rect 2404 8427 2407 8437
rect 2418 8430 2423 8434
rect 2427 8430 2434 8434
rect 2446 8427 2449 8437
rect 2462 8427 2465 8437
rect 2483 8427 2486 8437
rect 2499 8427 2502 8437
rect 2520 8427 2523 8437
rect 2536 8427 2539 8437
rect 2550 8430 2555 8434
rect 2559 8430 2566 8434
rect 2578 8427 2581 8437
rect 2594 8427 2597 8437
rect 2615 8427 2618 8437
rect 2631 8427 2634 8437
rect 2652 8427 2655 8437
rect 2668 8427 2671 8437
rect 2682 8430 2687 8434
rect 2691 8430 2698 8434
rect 2710 8427 2713 8437
rect 2726 8427 2729 8437
rect 2747 8427 2750 8437
rect 3312 8427 3315 8437
rect 3333 8427 3336 8437
rect 3349 8427 3352 8437
rect 3363 8430 3368 8434
rect 3372 8430 3379 8434
rect 3391 8427 3394 8437
rect 3407 8427 3410 8437
rect 3428 8427 3431 8437
rect 3444 8427 3447 8437
rect 3465 8427 3468 8437
rect 3481 8427 3484 8437
rect 3495 8430 3500 8434
rect 3504 8430 3511 8434
rect 3523 8427 3526 8437
rect 3539 8427 3542 8437
rect 3560 8427 3563 8437
rect 3576 8427 3579 8437
rect 3597 8427 3600 8437
rect 3613 8427 3616 8437
rect 3627 8430 3632 8434
rect 3636 8430 3643 8434
rect 3655 8427 3658 8437
rect 3671 8427 3674 8437
rect 3692 8427 3695 8437
rect 4483 8433 4484 8437
rect 4488 8433 4489 8437
rect 4493 8433 4494 8437
rect 4498 8433 4499 8437
rect 4503 8433 4504 8437
rect 4508 8433 4509 8437
rect 4479 8432 4513 8433
rect 4483 8428 4484 8432
rect 4488 8428 4489 8432
rect 4493 8428 4494 8432
rect 4498 8428 4499 8432
rect 4503 8428 4504 8432
rect 4508 8428 4509 8432
rect 4479 8427 4513 8428
rect 2384 8413 2389 8416
rect 2393 8413 2417 8416
rect 2442 8413 2449 8416
rect 2453 8413 2475 8416
rect 2495 8413 2502 8416
rect 2516 8413 2521 8416
rect 2525 8413 2549 8416
rect 2574 8413 2581 8416
rect 2585 8413 2607 8416
rect 2627 8413 2634 8416
rect 2648 8413 2653 8416
rect 2657 8413 2681 8416
rect 2706 8413 2713 8416
rect 2717 8413 2739 8416
rect 2400 8403 2407 8406
rect 2411 8407 2430 8410
rect 617 8394 618 8398
rect 622 8394 623 8398
rect 627 8394 628 8398
rect 632 8394 633 8398
rect 637 8394 638 8398
rect 642 8394 643 8398
rect 613 8393 647 8394
rect 617 8389 618 8393
rect 622 8389 623 8393
rect 627 8389 628 8393
rect 632 8389 633 8393
rect 637 8389 638 8393
rect 642 8389 643 8393
rect 613 8388 647 8389
rect 617 8384 618 8388
rect 622 8384 623 8388
rect 627 8384 628 8388
rect 632 8384 633 8388
rect 637 8384 638 8388
rect 642 8384 643 8388
rect 613 8383 647 8384
rect 86 8377 346 8380
rect 617 8379 618 8383
rect 622 8379 623 8383
rect 627 8379 628 8383
rect 632 8379 633 8383
rect 637 8379 638 8383
rect 642 8379 643 8383
rect 663 8394 664 8398
rect 668 8394 669 8398
rect 673 8394 674 8398
rect 678 8394 679 8398
rect 683 8394 684 8398
rect 688 8394 689 8398
rect 659 8393 693 8394
rect 663 8389 664 8393
rect 668 8389 669 8393
rect 673 8389 674 8393
rect 678 8389 679 8393
rect 683 8389 684 8393
rect 688 8389 689 8393
rect 659 8388 693 8389
rect 663 8384 664 8388
rect 668 8384 669 8388
rect 673 8384 674 8388
rect 678 8384 679 8388
rect 683 8384 684 8388
rect 688 8384 689 8388
rect 2430 8400 2433 8406
rect 2458 8403 2465 8406
rect 2469 8407 2484 8410
rect 2532 8403 2539 8406
rect 2543 8407 2562 8410
rect 2562 8400 2565 8406
rect 2590 8403 2597 8406
rect 2601 8407 2616 8410
rect 2664 8403 2671 8406
rect 2675 8407 2694 8410
rect 2694 8400 2697 8406
rect 2722 8403 2729 8406
rect 2733 8407 2750 8410
rect 3329 8413 3334 8416
rect 3338 8413 3362 8416
rect 3387 8413 3394 8416
rect 3398 8413 3420 8416
rect 3440 8413 3447 8416
rect 3461 8413 3466 8416
rect 3470 8413 3494 8416
rect 3519 8413 3526 8416
rect 3530 8413 3552 8416
rect 3572 8413 3579 8416
rect 3593 8413 3598 8416
rect 3602 8413 3626 8416
rect 4483 8423 4484 8427
rect 4488 8423 4489 8427
rect 4493 8423 4494 8427
rect 4498 8423 4499 8427
rect 4503 8423 4504 8427
rect 4508 8423 4509 8427
rect 4529 8438 4530 8442
rect 4534 8438 4535 8442
rect 4539 8438 4540 8442
rect 4544 8438 4545 8442
rect 4549 8438 4550 8442
rect 4554 8438 4555 8442
rect 4826 8441 5086 8444
rect 4525 8437 4559 8438
rect 4529 8433 4530 8437
rect 4534 8433 4535 8437
rect 4539 8433 4540 8437
rect 4544 8433 4545 8437
rect 4549 8433 4550 8437
rect 4554 8433 4555 8437
rect 4525 8432 4559 8433
rect 4529 8428 4530 8432
rect 4534 8428 4535 8432
rect 4539 8428 4540 8432
rect 4544 8428 4545 8432
rect 4549 8428 4550 8432
rect 4554 8428 4555 8432
rect 4525 8427 4559 8428
rect 4529 8423 4530 8427
rect 4534 8423 4535 8427
rect 4539 8423 4540 8427
rect 4544 8423 4545 8427
rect 4549 8423 4550 8427
rect 4554 8423 4555 8427
rect 3651 8413 3658 8416
rect 3662 8413 3684 8416
rect 3345 8403 3352 8406
rect 3356 8407 3375 8410
rect 3375 8400 3378 8406
rect 3403 8403 3410 8406
rect 3414 8407 3429 8410
rect 3477 8403 3484 8406
rect 3488 8407 3507 8410
rect 3507 8400 3510 8406
rect 3535 8403 3542 8406
rect 3546 8407 3561 8410
rect 3609 8403 3616 8406
rect 3620 8407 3639 8410
rect 3639 8400 3642 8406
rect 3667 8403 3674 8406
rect 3678 8407 3695 8410
rect 2367 8384 2370 8396
rect 2388 8384 2391 8396
rect 2404 8384 2407 8396
rect 2418 8387 2430 8390
rect 2446 8384 2449 8396
rect 2462 8384 2465 8396
rect 2483 8384 2486 8396
rect 2499 8384 2502 8396
rect 2520 8384 2523 8396
rect 2536 8384 2539 8396
rect 2550 8387 2562 8390
rect 2578 8384 2581 8396
rect 2594 8384 2597 8396
rect 2615 8384 2618 8396
rect 2631 8384 2634 8396
rect 2652 8384 2655 8396
rect 2668 8384 2671 8396
rect 2682 8387 2694 8390
rect 2710 8384 2713 8396
rect 2726 8384 2729 8396
rect 2747 8384 2750 8396
rect 3312 8384 3315 8396
rect 3333 8384 3336 8396
rect 3349 8384 3352 8396
rect 3363 8387 3375 8390
rect 3391 8384 3394 8396
rect 3407 8384 3410 8396
rect 3428 8384 3431 8396
rect 3444 8384 3447 8396
rect 3465 8384 3468 8396
rect 3481 8384 3484 8396
rect 3495 8387 3507 8390
rect 3523 8384 3526 8396
rect 3539 8384 3542 8396
rect 3560 8384 3563 8396
rect 3576 8384 3579 8396
rect 3597 8384 3600 8396
rect 3613 8384 3616 8396
rect 3627 8387 3639 8390
rect 3655 8384 3658 8396
rect 3671 8384 3674 8396
rect 3692 8384 3695 8396
rect 4826 8389 5086 8392
rect 659 8383 693 8384
rect 663 8379 664 8383
rect 668 8379 669 8383
rect 673 8379 674 8383
rect 678 8379 679 8383
rect 683 8379 684 8383
rect 688 8379 689 8383
rect 2364 8380 2397 8384
rect 2401 8380 2425 8384
rect 2429 8380 2455 8384
rect 2459 8380 2529 8384
rect 2533 8380 2557 8384
rect 2561 8380 2587 8384
rect 2591 8380 2661 8384
rect 2665 8380 2689 8384
rect 2693 8380 2719 8384
rect 2723 8380 2776 8384
rect 3309 8380 3342 8384
rect 3346 8380 3370 8384
rect 3374 8380 3400 8384
rect 3404 8380 3474 8384
rect 3478 8380 3502 8384
rect 3506 8380 3532 8384
rect 3536 8380 3606 8384
rect 3610 8380 3634 8384
rect 3638 8380 3664 8384
rect 3668 8380 3721 8384
rect 86 8123 89 8377
rect 343 8338 346 8377
rect 2364 8373 2373 8377
rect 2377 8373 2424 8377
rect 2428 8373 2474 8377
rect 2478 8373 2505 8377
rect 2509 8373 2556 8377
rect 2560 8373 2606 8377
rect 2610 8373 2637 8377
rect 2641 8373 2688 8377
rect 2692 8373 2738 8377
rect 2742 8373 2812 8377
rect 3309 8373 3318 8377
rect 3322 8373 3369 8377
rect 3373 8373 3419 8377
rect 3423 8373 3450 8377
rect 3454 8373 3501 8377
rect 3505 8373 3551 8377
rect 3555 8373 3582 8377
rect 3586 8373 3633 8377
rect 3637 8373 3683 8377
rect 3687 8373 3757 8377
rect 2830 8365 2857 8369
rect 2861 8365 2893 8369
rect 2897 8365 2960 8369
rect 2964 8365 2989 8369
rect 2993 8365 3025 8369
rect 3029 8365 3092 8369
rect 3096 8365 3121 8369
rect 3125 8365 3157 8369
rect 3161 8365 3224 8369
rect 3228 8365 3253 8369
rect 3257 8365 3289 8369
rect 3293 8365 3356 8369
rect 3360 8365 3376 8369
rect 3775 8365 3802 8369
rect 3806 8365 3838 8369
rect 3842 8365 3905 8369
rect 3909 8365 3934 8369
rect 3938 8365 3970 8369
rect 3974 8365 4037 8369
rect 4041 8365 4066 8369
rect 4070 8365 4102 8369
rect 4106 8365 4169 8369
rect 4173 8365 4198 8369
rect 4202 8365 4234 8369
rect 4238 8365 4301 8369
rect 4305 8365 4321 8369
rect 2770 8358 2881 8362
rect 2885 8358 2909 8362
rect 2913 8358 2939 8362
rect 2943 8358 2976 8362
rect 2980 8358 3013 8362
rect 3017 8358 3041 8362
rect 3045 8358 3071 8362
rect 3075 8358 3108 8362
rect 3112 8358 3145 8362
rect 3149 8358 3173 8362
rect 3177 8358 3203 8362
rect 3207 8358 3240 8362
rect 3244 8358 3277 8362
rect 3281 8358 3305 8362
rect 3309 8358 3335 8362
rect 3339 8358 3372 8362
rect 3715 8358 3826 8362
rect 3830 8358 3854 8362
rect 3858 8358 3884 8362
rect 3888 8358 3921 8362
rect 3925 8358 3958 8362
rect 3962 8358 3986 8362
rect 3990 8358 4016 8362
rect 4020 8358 4053 8362
rect 4057 8358 4090 8362
rect 4094 8358 4118 8362
rect 4122 8358 4148 8362
rect 4152 8358 4185 8362
rect 4189 8358 4222 8362
rect 4226 8358 4250 8362
rect 4254 8358 4280 8362
rect 4284 8358 4317 8362
rect 2851 8348 2854 8358
rect 2872 8348 2875 8358
rect 2888 8348 2891 8358
rect 2902 8351 2907 8355
rect 2911 8351 2918 8355
rect 2930 8348 2933 8358
rect 2946 8348 2949 8358
rect 2967 8348 2970 8358
rect 2983 8348 2986 8358
rect 3004 8348 3007 8358
rect 3020 8348 3023 8358
rect 3034 8351 3039 8355
rect 3043 8351 3050 8355
rect 3062 8348 3065 8358
rect 3078 8348 3081 8358
rect 3099 8348 3102 8358
rect 3115 8348 3118 8358
rect 3136 8348 3139 8358
rect 3152 8348 3155 8358
rect 3166 8351 3171 8355
rect 3175 8351 3182 8355
rect 3194 8348 3197 8358
rect 3210 8348 3213 8358
rect 3231 8348 3234 8358
rect 3247 8348 3250 8358
rect 3268 8348 3271 8358
rect 3284 8348 3287 8358
rect 3298 8351 3303 8355
rect 3307 8351 3314 8355
rect 3326 8348 3329 8358
rect 3342 8348 3345 8358
rect 3363 8348 3366 8358
rect 3796 8348 3799 8358
rect 3817 8348 3820 8358
rect 3833 8348 3836 8358
rect 3847 8351 3852 8355
rect 3856 8351 3863 8355
rect 3875 8348 3878 8358
rect 3891 8348 3894 8358
rect 3912 8348 3915 8358
rect 3928 8348 3931 8358
rect 3949 8348 3952 8358
rect 3965 8348 3968 8358
rect 3979 8351 3984 8355
rect 3988 8351 3995 8355
rect 4007 8348 4010 8358
rect 4023 8348 4026 8358
rect 4044 8348 4047 8358
rect 4060 8348 4063 8358
rect 4081 8348 4084 8358
rect 4097 8348 4100 8358
rect 4111 8351 4116 8355
rect 4120 8351 4127 8355
rect 4139 8348 4142 8358
rect 4155 8348 4158 8358
rect 4176 8348 4179 8358
rect 4192 8348 4195 8358
rect 4213 8348 4216 8358
rect 4229 8348 4232 8358
rect 4243 8351 4248 8355
rect 4252 8351 4259 8355
rect 4271 8348 4274 8358
rect 4287 8348 4290 8358
rect 4308 8348 4311 8358
rect 4826 8350 4829 8389
rect 343 8328 356 8338
rect 2496 8332 2505 8336
rect 2509 8332 2541 8336
rect 2545 8332 2608 8336
rect 2612 8332 2824 8336
rect 2868 8334 2873 8337
rect 2877 8334 2901 8337
rect 2926 8334 2933 8337
rect 2937 8334 2959 8337
rect 343 8318 366 8328
rect 2496 8325 2529 8329
rect 2533 8325 2557 8329
rect 2561 8325 2587 8329
rect 2591 8325 2624 8329
rect 2628 8325 2764 8329
rect 343 8308 376 8318
rect 2499 8315 2502 8325
rect 2520 8315 2523 8325
rect 2536 8315 2539 8325
rect 2550 8318 2555 8322
rect 2559 8318 2566 8322
rect 2578 8315 2581 8325
rect 2594 8315 2597 8325
rect 2615 8315 2618 8325
rect 2884 8324 2891 8327
rect 2895 8328 2914 8331
rect 2914 8321 2917 8327
rect 2942 8324 2949 8327
rect 2953 8328 2970 8331
rect 3000 8334 3005 8337
rect 3009 8334 3033 8337
rect 3058 8334 3065 8337
rect 3069 8334 3091 8337
rect 3016 8324 3023 8327
rect 3027 8328 3046 8331
rect 3046 8321 3049 8327
rect 3074 8324 3081 8327
rect 3085 8328 3102 8331
rect 3132 8334 3137 8337
rect 3141 8334 3165 8337
rect 3190 8334 3197 8337
rect 3201 8334 3223 8337
rect 3148 8324 3155 8327
rect 3159 8328 3178 8331
rect 3178 8321 3181 8327
rect 3206 8324 3213 8327
rect 3217 8328 3234 8331
rect 3264 8334 3269 8337
rect 3273 8334 3297 8337
rect 3322 8334 3329 8337
rect 3333 8334 3355 8337
rect 3441 8332 3450 8336
rect 3454 8332 3486 8336
rect 3490 8332 3553 8336
rect 3557 8332 3769 8336
rect 3280 8324 3287 8327
rect 3291 8328 3310 8331
rect 343 8298 386 8308
rect 2494 8298 2503 8302
rect 2516 8301 2521 8304
rect 2525 8301 2549 8304
rect 2574 8301 2581 8304
rect 2585 8301 2607 8304
rect 2851 8305 2854 8317
rect 2872 8305 2875 8317
rect 2888 8305 2891 8317
rect 2902 8308 2914 8311
rect 2930 8305 2933 8317
rect 2946 8305 2949 8317
rect 2967 8305 2970 8317
rect 2983 8305 2986 8317
rect 3004 8305 3007 8317
rect 3020 8305 3023 8317
rect 3034 8308 3046 8311
rect 3062 8305 3065 8317
rect 3078 8305 3081 8317
rect 3099 8305 3102 8317
rect 3115 8305 3118 8317
rect 3136 8305 3139 8317
rect 3152 8305 3155 8317
rect 3166 8308 3178 8311
rect 3194 8305 3197 8317
rect 3210 8305 3213 8317
rect 3231 8305 3234 8317
rect 3310 8321 3313 8327
rect 3338 8324 3345 8327
rect 3349 8328 3366 8331
rect 3813 8334 3818 8337
rect 3822 8334 3846 8337
rect 3871 8334 3878 8337
rect 3882 8334 3904 8337
rect 3441 8325 3474 8329
rect 3478 8325 3502 8329
rect 3506 8325 3532 8329
rect 3536 8325 3569 8329
rect 3573 8325 3709 8329
rect 3247 8305 3250 8317
rect 3268 8305 3271 8317
rect 3284 8305 3287 8317
rect 3298 8308 3310 8311
rect 3326 8305 3329 8317
rect 3342 8305 3345 8317
rect 3363 8305 3366 8317
rect 3444 8315 3447 8325
rect 3465 8315 3468 8325
rect 3481 8315 3484 8325
rect 3495 8318 3500 8322
rect 3504 8318 3511 8322
rect 3523 8315 3526 8325
rect 3539 8315 3542 8325
rect 3560 8315 3563 8325
rect 3829 8324 3836 8327
rect 3840 8328 3859 8331
rect 3859 8321 3862 8327
rect 3887 8324 3894 8327
rect 3898 8328 3915 8331
rect 3945 8334 3950 8337
rect 3954 8334 3978 8337
rect 4003 8334 4010 8337
rect 4014 8334 4036 8337
rect 3961 8324 3968 8327
rect 3972 8328 3991 8331
rect 3991 8321 3994 8327
rect 4019 8324 4026 8327
rect 4030 8328 4047 8331
rect 4077 8334 4082 8337
rect 4086 8334 4110 8337
rect 4135 8334 4142 8337
rect 4146 8334 4168 8337
rect 4093 8324 4100 8327
rect 4104 8328 4123 8331
rect 4123 8321 4126 8327
rect 4151 8324 4158 8327
rect 4162 8328 4179 8331
rect 4209 8334 4214 8337
rect 4218 8334 4242 8337
rect 4816 8340 4829 8350
rect 4267 8334 4274 8337
rect 4278 8334 4300 8337
rect 4225 8324 4232 8327
rect 4236 8328 4255 8331
rect 2782 8301 2881 8305
rect 2885 8301 2909 8305
rect 2913 8301 2939 8305
rect 2943 8301 3013 8305
rect 3017 8301 3041 8305
rect 3045 8301 3071 8305
rect 3075 8301 3145 8305
rect 3149 8301 3173 8305
rect 3177 8301 3203 8305
rect 3207 8301 3277 8305
rect 3281 8301 3305 8305
rect 3309 8301 3335 8305
rect 3339 8301 3376 8305
rect 343 8202 769 8298
rect 2532 8291 2539 8294
rect 2543 8295 2562 8298
rect 2562 8288 2565 8294
rect 2590 8291 2597 8294
rect 2601 8295 2616 8298
rect 3439 8298 3448 8302
rect 3461 8301 3466 8304
rect 3470 8301 3494 8304
rect 3519 8301 3526 8304
rect 3530 8301 3552 8304
rect 3796 8305 3799 8317
rect 3817 8305 3820 8317
rect 3833 8305 3836 8317
rect 3847 8308 3859 8311
rect 3875 8305 3878 8317
rect 3891 8305 3894 8317
rect 3912 8305 3915 8317
rect 3928 8305 3931 8317
rect 3949 8305 3952 8317
rect 3965 8305 3968 8317
rect 3979 8308 3991 8311
rect 4007 8305 4010 8317
rect 4023 8305 4026 8317
rect 4044 8305 4047 8317
rect 4060 8305 4063 8317
rect 4081 8305 4084 8317
rect 4097 8305 4100 8317
rect 4111 8308 4123 8311
rect 4139 8305 4142 8317
rect 4155 8305 4158 8317
rect 4176 8305 4179 8317
rect 4255 8321 4258 8327
rect 4283 8324 4290 8327
rect 4294 8328 4311 8331
rect 4806 8330 4829 8340
rect 4796 8320 4829 8330
rect 4192 8305 4195 8317
rect 4213 8305 4216 8317
rect 4229 8305 4232 8317
rect 4243 8308 4255 8311
rect 4271 8305 4274 8317
rect 4287 8305 4290 8317
rect 4308 8305 4311 8317
rect 4786 8310 4829 8320
rect 3727 8301 3826 8305
rect 3830 8301 3854 8305
rect 3858 8301 3884 8305
rect 3888 8301 3958 8305
rect 3962 8301 3986 8305
rect 3990 8301 4016 8305
rect 4020 8301 4090 8305
rect 4094 8301 4118 8305
rect 4122 8301 4148 8305
rect 4152 8301 4222 8305
rect 4226 8301 4250 8305
rect 4254 8301 4280 8305
rect 4284 8301 4321 8305
rect 2818 8294 2857 8298
rect 2861 8294 2908 8298
rect 2912 8294 2958 8298
rect 2962 8294 2989 8298
rect 2993 8294 3040 8298
rect 3044 8294 3090 8298
rect 3094 8294 3121 8298
rect 3125 8294 3172 8298
rect 3176 8294 3222 8298
rect 3226 8294 3253 8298
rect 3257 8294 3304 8298
rect 3308 8294 3354 8298
rect 3358 8294 3376 8298
rect 3477 8291 3484 8294
rect 3488 8295 3507 8298
rect 2499 8272 2502 8284
rect 2520 8272 2523 8284
rect 2536 8272 2539 8284
rect 2550 8275 2562 8278
rect 2578 8272 2581 8284
rect 2594 8272 2597 8284
rect 2615 8272 2618 8284
rect 2770 8281 2855 8285
rect 2859 8281 2871 8285
rect 2875 8281 2889 8285
rect 2893 8281 2900 8285
rect 2904 8281 2906 8285
rect 2910 8281 2925 8285
rect 2929 8281 2962 8285
rect 2966 8281 2967 8285
rect 2971 8281 2979 8285
rect 2983 8281 3007 8285
rect 3011 8281 3023 8285
rect 3027 8281 3047 8285
rect 3051 8281 3101 8285
rect 3105 8281 3128 8285
rect 3132 8281 3182 8285
rect 3186 8281 3205 8285
rect 3507 8288 3510 8294
rect 3535 8291 3542 8294
rect 3546 8295 3561 8298
rect 3763 8294 3802 8298
rect 3806 8294 3853 8298
rect 3857 8294 3903 8298
rect 3907 8294 3934 8298
rect 3938 8294 3985 8298
rect 3989 8294 4035 8298
rect 4039 8294 4066 8298
rect 4070 8294 4117 8298
rect 4121 8294 4167 8298
rect 4171 8294 4198 8298
rect 4202 8294 4249 8298
rect 4253 8294 4299 8298
rect 4303 8294 4321 8298
rect 2806 8274 2882 8278
rect 2886 8274 2913 8278
rect 2917 8274 2935 8278
rect 2939 8274 3000 8278
rect 3004 8274 3018 8278
rect 3030 8277 3033 8281
rect 2496 8268 2529 8272
rect 2533 8268 2557 8272
rect 2561 8268 2587 8272
rect 2591 8268 2776 8272
rect 2496 8261 2505 8265
rect 2509 8261 2556 8265
rect 2560 8261 2606 8265
rect 2610 8261 2812 8265
rect 2925 8267 2928 8271
rect 2952 8267 2953 8271
rect 2997 8267 2999 8271
rect 3039 8264 3042 8269
rect 3054 8271 3057 8281
rect 3084 8277 3087 8281
rect 3111 8277 3114 8281
rect 2494 8245 2510 8249
rect 2619 8247 2623 8251
rect 2635 8247 2639 8251
rect 2643 8247 2849 8251
rect 2853 8247 2857 8251
rect 2865 8250 2868 8256
rect 2872 8250 2875 8256
rect 2865 8247 2875 8250
rect 2865 8242 2868 8247
rect 2502 8238 2506 8242
rect 2518 8238 2639 8242
rect 2872 8242 2875 8247
rect 2881 8252 2884 8256
rect 2881 8248 2883 8252
rect 2887 8248 2889 8252
rect 2897 8251 2900 8256
rect 2925 8253 2928 8256
rect 2897 8249 2908 8251
rect 2881 8242 2884 8248
rect 2897 8247 2903 8249
rect 2897 8242 2900 8247
rect 2907 8247 2908 8249
rect 2926 8249 2928 8253
rect 2925 8242 2928 8249
rect 3028 8260 3031 8263
rect 3070 8260 3073 8263
rect 2941 8252 2944 8256
rect 2951 8252 2954 8256
rect 2951 8248 2960 8252
rect 2972 8251 2975 8256
rect 2997 8252 3000 8256
rect 2941 8242 2944 8248
rect 2951 8242 2954 8248
rect 2972 8247 2973 8251
rect 2977 8247 2980 8250
rect 2999 8248 3000 8252
rect 3015 8251 3018 8256
rect 3039 8255 3042 8260
rect 3047 8256 3058 8259
rect 3070 8257 3078 8260
rect 2972 8242 2975 8247
rect 2997 8242 3000 8248
rect 3015 8242 3018 8247
rect 2489 8230 2505 8234
rect 2509 8230 2572 8234
rect 2576 8230 2608 8234
rect 2612 8230 2824 8234
rect 2917 8229 2918 8233
rect 2942 8230 2943 8234
rect 2989 8229 2990 8233
rect 2493 8223 2526 8227
rect 2530 8223 2556 8227
rect 2560 8223 2584 8227
rect 2588 8223 2764 8227
rect 2499 8213 2502 8223
rect 2520 8213 2523 8223
rect 2536 8213 2539 8223
rect 2551 8216 2558 8220
rect 2562 8216 2567 8220
rect 2578 8213 2581 8223
rect 2594 8213 2597 8223
rect 2615 8213 2618 8223
rect 2794 8222 2870 8226
rect 2874 8222 2929 8226
rect 2933 8222 2954 8226
rect 2958 8222 2985 8226
rect 2989 8222 3018 8226
rect 3030 8219 3033 8251
rect 3047 8250 3050 8256
rect 3070 8251 3073 8257
rect 3082 8252 3085 8255
rect 3093 8255 3096 8269
rect 3120 8264 3123 8269
rect 3135 8271 3138 8281
rect 3165 8277 3168 8281
rect 3104 8260 3105 8263
rect 3109 8260 3112 8263
rect 3444 8272 3447 8284
rect 3465 8272 3468 8284
rect 3481 8272 3484 8284
rect 3495 8275 3507 8278
rect 3523 8272 3526 8284
rect 3539 8272 3542 8284
rect 3560 8272 3563 8284
rect 3715 8281 3800 8285
rect 3804 8281 3816 8285
rect 3820 8281 3834 8285
rect 3838 8281 3845 8285
rect 3849 8281 3851 8285
rect 3855 8281 3870 8285
rect 3874 8281 3907 8285
rect 3911 8281 3912 8285
rect 3916 8281 3924 8285
rect 3928 8281 3952 8285
rect 3956 8281 3968 8285
rect 3972 8281 3992 8285
rect 3996 8281 4046 8285
rect 4050 8281 4073 8285
rect 4077 8281 4127 8285
rect 4131 8281 4150 8285
rect 3751 8274 3827 8278
rect 3831 8274 3858 8278
rect 3862 8274 3880 8278
rect 3884 8274 3945 8278
rect 3949 8274 3963 8278
rect 3975 8277 3978 8281
rect 3151 8260 3154 8263
rect 3093 8252 3101 8255
rect 3120 8255 3123 8260
rect 3093 8247 3096 8252
rect 3101 8248 3105 8252
rect 3128 8256 3139 8259
rect 3151 8257 3159 8260
rect 3045 8241 3050 8246
rect 3054 8219 3057 8247
rect 3084 8219 3087 8243
rect 3111 8219 3114 8251
rect 3128 8250 3131 8256
rect 3151 8251 3154 8257
rect 3163 8252 3166 8255
rect 3174 8255 3177 8269
rect 3441 8268 3474 8272
rect 3478 8268 3502 8272
rect 3506 8268 3532 8272
rect 3536 8268 3721 8272
rect 3441 8261 3450 8265
rect 3454 8261 3501 8265
rect 3505 8261 3551 8265
rect 3555 8261 3757 8265
rect 3870 8267 3873 8271
rect 3897 8267 3898 8271
rect 3942 8267 3944 8271
rect 3984 8264 3987 8269
rect 3999 8271 4002 8281
rect 4029 8277 4032 8281
rect 4056 8277 4059 8281
rect 3174 8252 3186 8255
rect 3174 8247 3177 8252
rect 3126 8241 3131 8246
rect 3135 8219 3138 8247
rect 3439 8245 3455 8249
rect 3564 8247 3568 8251
rect 3580 8247 3584 8251
rect 3588 8247 3794 8251
rect 3798 8247 3802 8251
rect 3810 8250 3813 8256
rect 3817 8250 3820 8256
rect 3810 8247 3820 8250
rect 3165 8219 3168 8243
rect 3810 8242 3813 8247
rect 3447 8238 3451 8242
rect 3463 8238 3584 8242
rect 3817 8242 3820 8247
rect 3826 8252 3829 8256
rect 3826 8248 3828 8252
rect 3832 8248 3834 8252
rect 3842 8251 3845 8256
rect 3870 8253 3873 8256
rect 3842 8249 3853 8251
rect 3826 8242 3829 8248
rect 3842 8247 3848 8249
rect 3842 8242 3845 8247
rect 3852 8247 3853 8249
rect 3871 8249 3873 8253
rect 3870 8242 3873 8249
rect 3973 8260 3976 8263
rect 4015 8260 4018 8263
rect 3886 8252 3889 8256
rect 3896 8252 3899 8256
rect 3896 8248 3905 8252
rect 3917 8251 3920 8256
rect 3942 8252 3945 8256
rect 3886 8242 3889 8248
rect 3896 8242 3899 8248
rect 3917 8247 3918 8251
rect 3922 8247 3925 8250
rect 3944 8248 3945 8252
rect 3960 8251 3963 8256
rect 3984 8255 3987 8260
rect 3992 8256 4003 8259
rect 4015 8257 4023 8260
rect 3917 8242 3920 8247
rect 3942 8242 3945 8248
rect 3960 8242 3963 8247
rect 3434 8230 3450 8234
rect 3454 8230 3517 8234
rect 3521 8230 3553 8234
rect 3557 8230 3769 8234
rect 3862 8229 3863 8233
rect 3887 8230 3888 8234
rect 3934 8229 3935 8233
rect 3438 8223 3471 8227
rect 3475 8223 3501 8227
rect 3505 8223 3529 8227
rect 3533 8223 3709 8227
rect 2782 8215 2856 8219
rect 2860 8215 2862 8219
rect 2866 8215 2870 8219
rect 2874 8215 2888 8219
rect 2892 8215 2897 8219
rect 2901 8215 2906 8219
rect 2910 8215 2929 8219
rect 2933 8215 2963 8219
rect 2967 8215 2978 8219
rect 2982 8215 3006 8219
rect 3010 8215 3023 8219
rect 3027 8215 3047 8219
rect 3051 8215 3101 8219
rect 3108 8215 3128 8219
rect 3132 8215 3182 8219
rect 343 8192 386 8202
rect 2510 8199 2532 8202
rect 2536 8199 2543 8202
rect 2794 8208 2870 8212
rect 2874 8208 2929 8212
rect 2933 8208 2954 8212
rect 2958 8208 2985 8212
rect 2989 8208 3018 8212
rect 2568 8199 2592 8202
rect 2596 8199 2601 8202
rect 2917 8201 2918 8205
rect 2942 8200 2943 8204
rect 2989 8201 2990 8205
rect 2614 8196 2623 8200
rect 2501 8193 2516 8196
rect 343 8182 376 8192
rect 2555 8193 2574 8196
rect 2520 8189 2527 8192
rect 2552 8186 2555 8192
rect 2578 8189 2585 8192
rect 2865 8187 2868 8192
rect 2872 8187 2875 8192
rect 2855 8184 2857 8187
rect 2865 8184 2875 8187
rect 343 8172 366 8182
rect 343 8162 356 8172
rect 2499 8170 2502 8182
rect 2520 8170 2523 8182
rect 2536 8170 2539 8182
rect 2555 8173 2567 8176
rect 2578 8170 2581 8182
rect 2594 8170 2597 8182
rect 2615 8170 2618 8182
rect 2865 8178 2868 8184
rect 2872 8178 2875 8184
rect 2881 8186 2884 8192
rect 2897 8187 2900 8192
rect 2881 8182 2883 8186
rect 2887 8182 2889 8186
rect 2897 8185 2903 8187
rect 2907 8185 2908 8187
rect 2897 8183 2908 8185
rect 2925 8185 2928 8192
rect 2881 8178 2884 8182
rect 2897 8178 2900 8183
rect 2926 8181 2928 8185
rect 2925 8178 2928 8181
rect 2941 8186 2944 8192
rect 2951 8186 2954 8192
rect 2972 8187 2975 8192
rect 2951 8182 2960 8186
rect 2972 8183 2973 8187
rect 2977 8184 2980 8187
rect 2997 8186 3000 8192
rect 3015 8187 3018 8192
rect 3054 8195 3057 8215
rect 3135 8195 3138 8215
rect 3444 8213 3447 8223
rect 3465 8213 3468 8223
rect 3481 8213 3484 8223
rect 3496 8216 3503 8220
rect 3507 8216 3512 8220
rect 3523 8213 3526 8223
rect 3539 8213 3542 8223
rect 3560 8213 3563 8223
rect 3739 8222 3815 8226
rect 3819 8222 3874 8226
rect 3878 8222 3899 8226
rect 3903 8222 3930 8226
rect 3934 8222 3963 8226
rect 3975 8219 3978 8251
rect 3992 8250 3995 8256
rect 4015 8251 4018 8257
rect 4027 8252 4030 8255
rect 4038 8255 4041 8269
rect 4065 8264 4068 8269
rect 4080 8271 4083 8281
rect 4110 8277 4113 8281
rect 4049 8260 4050 8263
rect 4054 8260 4057 8263
rect 4096 8260 4099 8263
rect 4038 8252 4046 8255
rect 4065 8255 4068 8260
rect 4038 8247 4041 8252
rect 4046 8248 4050 8252
rect 4073 8256 4084 8259
rect 4096 8257 4104 8260
rect 3990 8241 3995 8246
rect 3999 8219 4002 8247
rect 4029 8219 4032 8243
rect 4056 8219 4059 8251
rect 4073 8250 4076 8256
rect 4096 8251 4099 8257
rect 4108 8252 4111 8255
rect 4119 8255 4122 8269
rect 4119 8252 4131 8255
rect 4119 8247 4122 8252
rect 4071 8241 4076 8246
rect 4080 8219 4083 8247
rect 4110 8219 4113 8243
rect 3727 8215 3801 8219
rect 3805 8215 3807 8219
rect 3811 8215 3815 8219
rect 3819 8215 3833 8219
rect 3837 8215 3842 8219
rect 3846 8215 3851 8219
rect 3855 8215 3874 8219
rect 3878 8215 3908 8219
rect 3912 8215 3923 8219
rect 3927 8215 3951 8219
rect 3955 8215 3968 8219
rect 3972 8215 3992 8219
rect 3996 8215 4046 8219
rect 4053 8215 4073 8219
rect 4077 8215 4127 8219
rect 3455 8199 3477 8202
rect 3481 8199 3488 8202
rect 3739 8208 3815 8212
rect 3819 8208 3874 8212
rect 3878 8208 3899 8212
rect 3903 8208 3930 8212
rect 3934 8208 3963 8212
rect 3513 8199 3537 8202
rect 3541 8199 3546 8202
rect 3862 8201 3863 8205
rect 3887 8200 3888 8204
rect 3934 8201 3935 8205
rect 3559 8196 3568 8200
rect 3446 8193 3461 8196
rect 2941 8178 2944 8182
rect 2951 8178 2954 8182
rect 2972 8178 2975 8183
rect 2999 8182 3000 8186
rect 2997 8178 3000 8182
rect 3015 8178 3018 8183
rect 3045 8182 3050 8187
rect 3054 8183 3055 8186
rect 3070 8185 3073 8191
rect 3070 8182 3078 8185
rect 3125 8182 3130 8187
rect 3134 8183 3136 8186
rect 3151 8185 3154 8191
rect 3500 8193 3519 8196
rect 3465 8189 3472 8192
rect 3497 8186 3500 8192
rect 3151 8182 3159 8185
rect 3523 8189 3530 8192
rect 3810 8187 3813 8192
rect 3817 8187 3820 8192
rect 3800 8184 3802 8187
rect 3810 8184 3820 8187
rect 3070 8179 3073 8182
rect 3151 8179 3154 8182
rect 2489 8166 2526 8170
rect 2530 8166 2556 8170
rect 2560 8166 2584 8170
rect 2588 8166 2776 8170
rect 2925 8163 2928 8167
rect 2952 8163 2953 8167
rect 2997 8163 2999 8167
rect 343 8123 346 8162
rect 2489 8159 2507 8163
rect 2511 8159 2557 8163
rect 2561 8159 2608 8163
rect 2612 8159 2812 8163
rect 2870 8156 2882 8160
rect 2886 8156 2913 8160
rect 2917 8156 2935 8160
rect 2939 8156 3000 8160
rect 3004 8156 3018 8160
rect 3054 8153 3057 8171
rect 3135 8153 3138 8171
rect 3444 8170 3447 8182
rect 3465 8170 3468 8182
rect 3481 8170 3484 8182
rect 3500 8173 3512 8176
rect 3523 8170 3526 8182
rect 3539 8170 3542 8182
rect 3560 8170 3563 8182
rect 3810 8178 3813 8184
rect 3817 8178 3820 8184
rect 3826 8186 3829 8192
rect 3842 8187 3845 8192
rect 3826 8182 3828 8186
rect 3832 8182 3834 8186
rect 3842 8185 3848 8187
rect 3852 8185 3853 8187
rect 3842 8183 3853 8185
rect 3870 8185 3873 8192
rect 3826 8178 3829 8182
rect 3842 8178 3845 8183
rect 3871 8181 3873 8185
rect 3870 8178 3873 8181
rect 3886 8186 3889 8192
rect 3896 8186 3899 8192
rect 3917 8187 3920 8192
rect 3896 8182 3905 8186
rect 3917 8183 3918 8187
rect 3922 8184 3925 8187
rect 3942 8186 3945 8192
rect 3960 8187 3963 8192
rect 3999 8195 4002 8215
rect 4080 8195 4083 8215
rect 4403 8214 4829 8310
rect 4786 8204 4829 8214
rect 4796 8194 4829 8204
rect 3886 8178 3889 8182
rect 3896 8178 3899 8182
rect 3917 8178 3920 8183
rect 3944 8182 3945 8186
rect 3942 8178 3945 8182
rect 3960 8178 3963 8183
rect 3990 8182 3995 8187
rect 3999 8183 4000 8186
rect 4015 8185 4018 8191
rect 4015 8182 4023 8185
rect 4070 8182 4075 8187
rect 4079 8183 4081 8186
rect 4096 8185 4099 8191
rect 4096 8182 4104 8185
rect 4806 8184 4829 8194
rect 4015 8179 4018 8182
rect 4096 8179 4099 8182
rect 4816 8174 4829 8184
rect 3434 8166 3471 8170
rect 3475 8166 3501 8170
rect 3505 8166 3529 8170
rect 3533 8166 3721 8170
rect 3870 8163 3873 8167
rect 3897 8163 3898 8167
rect 3942 8163 3944 8167
rect 3434 8159 3452 8163
rect 3456 8159 3502 8163
rect 3506 8159 3553 8163
rect 3557 8159 3757 8163
rect 3815 8156 3827 8160
rect 3831 8156 3858 8160
rect 3862 8156 3880 8160
rect 3884 8156 3945 8160
rect 3949 8156 3963 8160
rect 3999 8153 4002 8171
rect 4080 8153 4083 8171
rect 2770 8149 2855 8153
rect 2859 8149 2871 8153
rect 2875 8149 2889 8153
rect 2893 8149 2900 8153
rect 2904 8149 2906 8153
rect 2910 8149 2925 8153
rect 2929 8149 2962 8153
rect 2966 8149 2967 8153
rect 2971 8149 2979 8153
rect 2983 8149 3007 8153
rect 3011 8149 3023 8153
rect 3027 8149 3047 8153
rect 3051 8149 3101 8153
rect 3105 8149 3128 8153
rect 3132 8149 3190 8153
rect 3194 8149 3205 8153
rect 3715 8149 3800 8153
rect 3804 8149 3816 8153
rect 3820 8149 3834 8153
rect 3838 8149 3845 8153
rect 3849 8149 3851 8153
rect 3855 8149 3870 8153
rect 3874 8149 3907 8153
rect 3911 8149 3912 8153
rect 3916 8149 3924 8153
rect 3928 8149 3952 8153
rect 3956 8149 3968 8153
rect 3972 8149 3992 8153
rect 3996 8149 4046 8153
rect 4050 8149 4073 8153
rect 4077 8149 4135 8153
rect 4139 8149 4150 8153
rect 2806 8142 2866 8146
rect 2870 8142 2882 8146
rect 2886 8142 2913 8146
rect 2917 8142 2935 8146
rect 2939 8142 3000 8146
rect 3004 8142 3018 8146
rect 3054 8139 3057 8149
rect 3084 8145 3087 8149
rect 3135 8145 3138 8149
rect 2925 8135 2928 8139
rect 2952 8135 2953 8139
rect 2997 8135 2999 8139
rect 86 8120 346 8123
rect 2854 8115 2857 8118
rect 2865 8118 2868 8124
rect 2872 8118 2875 8124
rect 2865 8115 2875 8118
rect 2865 8110 2868 8115
rect 2872 8110 2875 8115
rect 2881 8120 2884 8124
rect 2881 8116 2883 8120
rect 2887 8116 2889 8120
rect 2897 8119 2900 8124
rect 2925 8121 2928 8124
rect 2897 8117 2908 8119
rect 2881 8110 2884 8116
rect 2897 8115 2903 8117
rect 2897 8110 2900 8115
rect 2907 8115 2908 8117
rect 2926 8117 2928 8121
rect 2925 8110 2928 8117
rect 3070 8128 3073 8131
rect 2941 8120 2944 8124
rect 2951 8120 2954 8124
rect 2951 8116 2960 8120
rect 2972 8119 2975 8124
rect 2997 8120 3000 8124
rect 2941 8110 2944 8116
rect 2951 8110 2954 8116
rect 2972 8115 2973 8119
rect 2977 8115 2980 8118
rect 2999 8116 3000 8120
rect 3015 8119 3018 8124
rect 3047 8124 3058 8127
rect 3070 8125 3078 8128
rect 2972 8110 2975 8115
rect 2997 8110 3000 8116
rect 3047 8118 3050 8124
rect 3070 8119 3073 8125
rect 3082 8120 3085 8123
rect 3093 8123 3096 8137
rect 3144 8132 3147 8137
rect 3159 8139 3162 8149
rect 3189 8145 3192 8149
rect 3128 8128 3129 8131
rect 3133 8128 3136 8131
rect 3751 8142 3811 8146
rect 3815 8142 3827 8146
rect 3831 8142 3858 8146
rect 3862 8142 3880 8146
rect 3884 8142 3945 8146
rect 3949 8142 3963 8146
rect 3999 8139 4002 8149
rect 4029 8145 4032 8149
rect 4080 8145 4083 8149
rect 3175 8128 3178 8131
rect 3101 8123 3106 8128
rect 3144 8123 3147 8128
rect 3093 8120 3101 8123
rect 3015 8110 3018 8115
rect 3093 8115 3096 8120
rect 3152 8124 3163 8127
rect 3175 8125 3183 8128
rect 3045 8109 3050 8114
rect 2917 8097 2918 8101
rect 2942 8098 2943 8102
rect 2989 8097 2990 8101
rect 2794 8090 2870 8094
rect 2874 8090 2929 8094
rect 2933 8090 2954 8094
rect 2958 8090 2985 8094
rect 2989 8090 3018 8094
rect 617 8085 618 8089
rect 622 8085 623 8089
rect 627 8085 628 8089
rect 632 8085 633 8089
rect 637 8085 638 8089
rect 642 8085 643 8089
rect 613 8084 647 8085
rect 617 8080 618 8084
rect 622 8080 623 8084
rect 627 8080 628 8084
rect 632 8080 633 8084
rect 637 8080 638 8084
rect 642 8080 643 8084
rect 613 8079 647 8080
rect 617 8075 618 8079
rect 622 8075 623 8079
rect 627 8075 628 8079
rect 632 8075 633 8079
rect 637 8075 638 8079
rect 642 8075 643 8079
rect 613 8074 647 8075
rect 86 8068 346 8071
rect 617 8070 618 8074
rect 622 8070 623 8074
rect 627 8070 628 8074
rect 632 8070 633 8074
rect 637 8070 638 8074
rect 642 8070 643 8074
rect 663 8085 664 8089
rect 668 8085 669 8089
rect 673 8085 674 8089
rect 678 8085 679 8089
rect 683 8085 684 8089
rect 688 8085 689 8089
rect 3054 8087 3057 8115
rect 3084 8087 3087 8111
rect 3135 8087 3138 8119
rect 3152 8118 3155 8124
rect 3175 8119 3178 8125
rect 3187 8120 3190 8123
rect 3198 8123 3201 8137
rect 3870 8135 3873 8139
rect 3897 8135 3898 8139
rect 3942 8135 3944 8139
rect 3198 8120 3204 8123
rect 3198 8115 3201 8120
rect 3799 8115 3802 8118
rect 3810 8118 3813 8124
rect 3817 8118 3820 8124
rect 3810 8115 3820 8118
rect 3150 8109 3155 8114
rect 3159 8087 3162 8115
rect 3189 8087 3192 8111
rect 3810 8110 3813 8115
rect 3817 8110 3820 8115
rect 3826 8120 3829 8124
rect 3826 8116 3828 8120
rect 3832 8116 3834 8120
rect 3842 8119 3845 8124
rect 3870 8121 3873 8124
rect 3842 8117 3853 8119
rect 3826 8110 3829 8116
rect 3842 8115 3848 8117
rect 3842 8110 3845 8115
rect 3852 8115 3853 8117
rect 3871 8117 3873 8121
rect 3870 8110 3873 8117
rect 4015 8128 4018 8131
rect 3886 8120 3889 8124
rect 3896 8120 3899 8124
rect 3896 8116 3905 8120
rect 3917 8119 3920 8124
rect 3942 8120 3945 8124
rect 3886 8110 3889 8116
rect 3896 8110 3899 8116
rect 3917 8115 3918 8119
rect 3922 8115 3925 8118
rect 3944 8116 3945 8120
rect 3960 8119 3963 8124
rect 3992 8124 4003 8127
rect 4015 8125 4023 8128
rect 3917 8110 3920 8115
rect 3942 8110 3945 8116
rect 3992 8118 3995 8124
rect 4015 8119 4018 8125
rect 4027 8120 4030 8123
rect 4038 8123 4041 8137
rect 4089 8132 4092 8137
rect 4104 8139 4107 8149
rect 4134 8145 4137 8149
rect 4073 8128 4074 8131
rect 4078 8128 4081 8131
rect 4120 8128 4123 8131
rect 4046 8123 4051 8128
rect 4089 8123 4092 8128
rect 4038 8120 4046 8123
rect 3960 8110 3963 8115
rect 4038 8115 4041 8120
rect 4097 8124 4108 8127
rect 4120 8125 4128 8128
rect 3990 8109 3995 8114
rect 3862 8097 3863 8101
rect 3887 8098 3888 8102
rect 3934 8097 3935 8101
rect 3739 8090 3815 8094
rect 3819 8090 3874 8094
rect 3878 8090 3899 8094
rect 3903 8090 3930 8094
rect 3934 8090 3963 8094
rect 3999 8087 4002 8115
rect 4029 8087 4032 8111
rect 4080 8087 4083 8119
rect 4097 8118 4100 8124
rect 4120 8119 4123 8125
rect 4132 8120 4135 8123
rect 4143 8123 4146 8137
rect 4826 8135 4829 8174
rect 5083 8135 5086 8389
rect 4483 8129 4484 8133
rect 4488 8129 4489 8133
rect 4493 8129 4494 8133
rect 4498 8129 4499 8133
rect 4503 8129 4504 8133
rect 4508 8129 4509 8133
rect 4479 8128 4513 8129
rect 4483 8124 4484 8128
rect 4488 8124 4489 8128
rect 4493 8124 4494 8128
rect 4498 8124 4499 8128
rect 4503 8124 4504 8128
rect 4508 8124 4509 8128
rect 4143 8120 4149 8123
rect 4479 8123 4513 8124
rect 4143 8115 4146 8120
rect 4095 8109 4100 8114
rect 4104 8087 4107 8115
rect 4483 8119 4484 8123
rect 4488 8119 4489 8123
rect 4493 8119 4494 8123
rect 4498 8119 4499 8123
rect 4503 8119 4504 8123
rect 4508 8119 4509 8123
rect 4479 8118 4513 8119
rect 4483 8114 4484 8118
rect 4488 8114 4489 8118
rect 4493 8114 4494 8118
rect 4498 8114 4499 8118
rect 4503 8114 4504 8118
rect 4508 8114 4509 8118
rect 4529 8129 4530 8133
rect 4534 8129 4535 8133
rect 4539 8129 4540 8133
rect 4544 8129 4545 8133
rect 4549 8129 4550 8133
rect 4554 8129 4555 8133
rect 4826 8132 5086 8135
rect 4525 8128 4559 8129
rect 4529 8124 4530 8128
rect 4534 8124 4535 8128
rect 4539 8124 4540 8128
rect 4544 8124 4545 8128
rect 4549 8124 4550 8128
rect 4554 8124 4555 8128
rect 4525 8123 4559 8124
rect 4529 8119 4530 8123
rect 4534 8119 4535 8123
rect 4539 8119 4540 8123
rect 4544 8119 4545 8123
rect 4549 8119 4550 8123
rect 4554 8119 4555 8123
rect 4525 8118 4559 8119
rect 4529 8114 4530 8118
rect 4534 8114 4535 8118
rect 4539 8114 4540 8118
rect 4544 8114 4545 8118
rect 4549 8114 4550 8118
rect 4554 8114 4555 8118
rect 4134 8087 4137 8111
rect 4483 8098 4484 8102
rect 4488 8098 4489 8102
rect 4493 8098 4494 8102
rect 4498 8098 4499 8102
rect 4503 8098 4504 8102
rect 4508 8098 4509 8102
rect 4479 8097 4513 8098
rect 4483 8093 4484 8097
rect 4488 8093 4489 8097
rect 4493 8093 4494 8097
rect 4498 8093 4499 8097
rect 4503 8093 4504 8097
rect 4508 8093 4509 8097
rect 4479 8092 4513 8093
rect 4483 8088 4484 8092
rect 4488 8088 4489 8092
rect 4493 8088 4494 8092
rect 4498 8088 4499 8092
rect 4503 8088 4504 8092
rect 4508 8088 4509 8092
rect 4479 8087 4513 8088
rect 659 8084 693 8085
rect 663 8080 664 8084
rect 668 8080 669 8084
rect 673 8080 674 8084
rect 678 8080 679 8084
rect 683 8080 684 8084
rect 688 8080 689 8084
rect 2782 8083 2856 8087
rect 2860 8083 2862 8087
rect 2866 8083 2870 8087
rect 2874 8083 2888 8087
rect 2892 8083 2897 8087
rect 2901 8083 2906 8087
rect 2910 8083 2929 8087
rect 2933 8083 2963 8087
rect 2967 8083 2978 8087
rect 2982 8083 3006 8087
rect 3010 8083 3023 8087
rect 3027 8083 3047 8087
rect 3051 8083 3101 8087
rect 3105 8083 3128 8087
rect 3132 8083 3152 8087
rect 3156 8083 3204 8087
rect 3727 8083 3801 8087
rect 3805 8083 3807 8087
rect 3811 8083 3815 8087
rect 3819 8083 3833 8087
rect 3837 8083 3842 8087
rect 3846 8083 3851 8087
rect 3855 8083 3874 8087
rect 3878 8083 3908 8087
rect 3912 8083 3923 8087
rect 3927 8083 3951 8087
rect 3955 8083 3968 8087
rect 3972 8083 3992 8087
rect 3996 8083 4046 8087
rect 4050 8083 4073 8087
rect 4077 8083 4097 8087
rect 4101 8083 4149 8087
rect 4483 8083 4484 8087
rect 4488 8083 4489 8087
rect 4493 8083 4494 8087
rect 4498 8083 4499 8087
rect 4503 8083 4504 8087
rect 4508 8083 4509 8087
rect 4529 8098 4530 8102
rect 4534 8098 4535 8102
rect 4539 8098 4540 8102
rect 4544 8098 4545 8102
rect 4549 8098 4550 8102
rect 4554 8098 4555 8102
rect 4525 8097 4559 8098
rect 4529 8093 4530 8097
rect 4534 8093 4535 8097
rect 4539 8093 4540 8097
rect 4544 8093 4545 8097
rect 4549 8093 4550 8097
rect 4554 8093 4555 8097
rect 4525 8092 4559 8093
rect 4529 8088 4530 8092
rect 4534 8088 4535 8092
rect 4539 8088 4540 8092
rect 4544 8088 4545 8092
rect 4549 8088 4550 8092
rect 4554 8088 4555 8092
rect 4525 8087 4559 8088
rect 4529 8083 4530 8087
rect 4534 8083 4535 8087
rect 4539 8083 4540 8087
rect 4544 8083 4545 8087
rect 4549 8083 4550 8087
rect 4554 8083 4555 8087
rect 659 8079 693 8080
rect 663 8075 664 8079
rect 668 8075 669 8079
rect 673 8075 674 8079
rect 678 8075 679 8079
rect 683 8075 684 8079
rect 688 8075 689 8079
rect 2794 8076 2870 8080
rect 2874 8076 2929 8080
rect 2933 8076 2954 8080
rect 2958 8076 2985 8080
rect 2989 8076 3018 8080
rect 659 8074 693 8075
rect 663 8070 664 8074
rect 668 8070 669 8074
rect 673 8070 674 8074
rect 678 8070 679 8074
rect 683 8070 684 8074
rect 688 8070 689 8074
rect 2917 8069 2918 8073
rect 2942 8068 2943 8072
rect 2989 8069 2990 8073
rect 86 7814 89 8068
rect 343 8029 346 8068
rect 3054 8064 3057 8083
rect 3159 8064 3162 8083
rect 3739 8076 3815 8080
rect 3819 8076 3874 8080
rect 3878 8076 3899 8080
rect 3903 8076 3930 8080
rect 3934 8076 3963 8080
rect 3862 8069 3863 8073
rect 3887 8068 3888 8072
rect 3934 8069 3935 8073
rect 3999 8064 4002 8083
rect 4104 8064 4107 8083
rect 4826 8081 5086 8084
rect 4505 8078 4754 8080
rect 4505 8074 4506 8078
rect 4510 8074 4511 8078
rect 4515 8074 4754 8078
rect 4505 8073 4754 8074
rect 4505 8069 4506 8073
rect 4510 8069 4511 8073
rect 4515 8069 4754 8073
rect 4505 8068 4754 8069
rect 4505 8064 4506 8068
rect 4510 8064 4511 8068
rect 4515 8064 4754 8068
rect 2865 8055 2868 8060
rect 2872 8055 2875 8060
rect 2855 8052 2857 8055
rect 2865 8052 2875 8055
rect 2865 8046 2868 8052
rect 2872 8046 2875 8052
rect 2881 8054 2884 8060
rect 2897 8055 2900 8060
rect 2881 8050 2883 8054
rect 2887 8050 2889 8054
rect 2897 8053 2903 8055
rect 2907 8053 2908 8055
rect 2897 8051 2908 8053
rect 2925 8053 2928 8060
rect 2881 8046 2884 8050
rect 2897 8046 2900 8051
rect 2926 8049 2928 8053
rect 2925 8046 2928 8049
rect 2941 8054 2944 8060
rect 2951 8054 2954 8060
rect 2972 8055 2975 8060
rect 2951 8050 2960 8054
rect 2972 8051 2973 8055
rect 2977 8052 2980 8055
rect 2997 8054 3000 8060
rect 3015 8055 3018 8060
rect 2941 8046 2944 8050
rect 2951 8046 2954 8050
rect 2972 8046 2975 8051
rect 2999 8050 3000 8054
rect 3044 8051 3049 8056
rect 3053 8052 3055 8055
rect 3070 8054 3073 8060
rect 3070 8051 3078 8054
rect 3150 8051 3155 8056
rect 3159 8052 3160 8055
rect 3175 8054 3178 8060
rect 3175 8051 3183 8054
rect 3810 8055 3813 8060
rect 3817 8055 3820 8060
rect 3800 8052 3802 8055
rect 3810 8052 3820 8055
rect 2997 8046 3000 8050
rect 3015 8046 3018 8051
rect 3070 8048 3073 8051
rect 3175 8048 3178 8051
rect 3810 8046 3813 8052
rect 2925 8031 2928 8035
rect 2952 8031 2953 8035
rect 2997 8031 2999 8035
rect 343 8019 356 8029
rect 2806 8024 2882 8028
rect 2886 8024 2913 8028
rect 2917 8024 2935 8028
rect 2939 8024 3000 8028
rect 3004 8024 3018 8028
rect 3054 8021 3057 8040
rect 3159 8021 3162 8040
rect 3817 8046 3820 8052
rect 3826 8054 3829 8060
rect 3842 8055 3845 8060
rect 3826 8050 3828 8054
rect 3832 8050 3834 8054
rect 3842 8053 3848 8055
rect 3852 8053 3853 8055
rect 3842 8051 3853 8053
rect 3870 8053 3873 8060
rect 3826 8046 3829 8050
rect 3842 8046 3845 8051
rect 3871 8049 3873 8053
rect 3870 8046 3873 8049
rect 3886 8054 3889 8060
rect 3896 8054 3899 8060
rect 3917 8055 3920 8060
rect 3896 8050 3905 8054
rect 3917 8051 3918 8055
rect 3922 8052 3925 8055
rect 3942 8054 3945 8060
rect 3960 8055 3963 8060
rect 3886 8046 3889 8050
rect 3896 8046 3899 8050
rect 3917 8046 3920 8051
rect 3944 8050 3945 8054
rect 3989 8051 3994 8056
rect 3998 8052 4000 8055
rect 4015 8054 4018 8060
rect 4015 8051 4023 8054
rect 4095 8051 4100 8056
rect 4104 8052 4105 8055
rect 4120 8054 4123 8060
rect 4505 8063 4754 8064
rect 4505 8059 4506 8063
rect 4510 8059 4511 8063
rect 4515 8059 4754 8063
rect 4505 8058 4754 8059
rect 4120 8051 4128 8054
rect 4505 8054 4506 8058
rect 4510 8054 4511 8058
rect 4515 8054 4754 8058
rect 4505 8053 4754 8054
rect 3942 8046 3945 8050
rect 3960 8046 3963 8051
rect 4015 8048 4018 8051
rect 4120 8048 4123 8051
rect 4505 8049 4506 8053
rect 4510 8049 4511 8053
rect 4515 8049 4754 8053
rect 4505 8048 4754 8049
rect 4505 8044 4506 8048
rect 4510 8044 4511 8048
rect 4515 8044 4754 8048
rect 4505 8043 4754 8044
rect 3870 8031 3873 8035
rect 3897 8031 3898 8035
rect 3942 8031 3944 8035
rect 3751 8024 3827 8028
rect 3831 8024 3858 8028
rect 3862 8024 3880 8028
rect 3884 8024 3945 8028
rect 3949 8024 3963 8028
rect 3999 8021 4002 8040
rect 4104 8021 4107 8040
rect 4505 8039 4506 8043
rect 4510 8039 4511 8043
rect 4515 8039 4754 8043
rect 4826 8042 4829 8081
rect 4505 8038 4670 8039
rect 4505 8034 4506 8038
rect 4510 8034 4511 8038
rect 4515 8037 4670 8038
rect 4515 8034 4626 8037
rect 4645 8034 4649 8037
rect 4661 8034 4670 8037
rect 4688 8034 4692 8039
rect 4704 8034 4713 8039
rect 4729 8034 4733 8039
rect 4745 8034 4754 8039
rect 4505 8033 4626 8034
rect 4505 8029 4506 8033
rect 4510 8029 4511 8033
rect 4515 8029 4626 8033
rect 4505 8028 4626 8029
rect 4505 8024 4506 8028
rect 4510 8024 4511 8028
rect 4515 8024 4626 8028
rect 343 8009 366 8019
rect 2770 8017 2855 8021
rect 2859 8017 2871 8021
rect 2875 8017 2889 8021
rect 2893 8017 2900 8021
rect 2904 8017 2906 8021
rect 2910 8017 2925 8021
rect 2929 8017 2962 8021
rect 2966 8017 2967 8021
rect 2971 8017 2979 8021
rect 2983 8017 3007 8021
rect 3011 8017 3023 8021
rect 3027 8017 3047 8021
rect 3051 8017 3101 8021
rect 3105 8017 3128 8021
rect 3132 8017 3182 8021
rect 3186 8017 3190 8021
rect 3194 8017 3218 8021
rect 3222 8017 3272 8021
rect 3715 8017 3800 8021
rect 3804 8017 3816 8021
rect 3820 8017 3834 8021
rect 3838 8017 3845 8021
rect 3849 8017 3851 8021
rect 3855 8017 3870 8021
rect 3874 8017 3907 8021
rect 3911 8017 3912 8021
rect 3916 8017 3924 8021
rect 3928 8017 3952 8021
rect 3956 8017 3968 8021
rect 3972 8017 3992 8021
rect 3996 8017 4046 8021
rect 4050 8017 4073 8021
rect 4077 8017 4127 8021
rect 4131 8017 4135 8021
rect 4139 8017 4163 8021
rect 4167 8017 4217 8021
rect 2806 8010 2882 8014
rect 2886 8010 2913 8014
rect 2917 8010 2935 8014
rect 2939 8010 3000 8014
rect 3004 8010 3018 8014
rect 343 7999 376 8009
rect 3054 8007 3057 8017
rect 3084 8013 3087 8017
rect 3111 8013 3114 8017
rect 2925 8003 2928 8007
rect 2952 8003 2953 8007
rect 2997 8003 2999 8007
rect 343 7989 386 7999
rect 343 7893 769 7989
rect 2854 7983 2857 7986
rect 2865 7986 2868 7992
rect 2872 7986 2875 7992
rect 2865 7983 2875 7986
rect 2865 7978 2868 7983
rect 2872 7978 2875 7983
rect 2881 7988 2884 7992
rect 2881 7984 2883 7988
rect 2887 7984 2889 7988
rect 2897 7987 2900 7992
rect 2925 7989 2928 7992
rect 2897 7985 2908 7987
rect 2881 7978 2884 7984
rect 2897 7983 2903 7985
rect 2897 7978 2900 7983
rect 2907 7983 2908 7985
rect 2926 7985 2928 7989
rect 2925 7978 2928 7985
rect 3070 7996 3073 7999
rect 2941 7988 2944 7992
rect 2951 7988 2954 7992
rect 2951 7984 2960 7988
rect 2972 7987 2975 7992
rect 2997 7988 3000 7992
rect 2941 7978 2944 7984
rect 2951 7978 2954 7984
rect 2972 7983 2973 7987
rect 2977 7983 2980 7986
rect 2999 7984 3000 7988
rect 3015 7987 3018 7992
rect 3047 7992 3058 7995
rect 3070 7993 3078 7996
rect 2972 7978 2975 7983
rect 2997 7978 3000 7984
rect 3047 7986 3050 7992
rect 3070 7987 3073 7993
rect 3082 7988 3085 7991
rect 3093 7991 3096 8005
rect 3120 8000 3123 8005
rect 3135 8007 3138 8017
rect 3165 8013 3168 8017
rect 3201 8013 3204 8017
rect 3104 7996 3105 7999
rect 3109 7996 3112 7999
rect 3151 7996 3154 7999
rect 3093 7988 3101 7991
rect 3120 7991 3123 7996
rect 3015 7978 3018 7983
rect 3093 7983 3096 7988
rect 3101 7984 3105 7988
rect 3128 7992 3139 7995
rect 3151 7993 3159 7996
rect 3045 7977 3050 7982
rect 2917 7965 2918 7969
rect 2942 7966 2943 7970
rect 2989 7965 2990 7969
rect 2794 7958 2870 7962
rect 2874 7958 2929 7962
rect 2933 7958 2954 7962
rect 2958 7958 2985 7962
rect 2989 7958 3018 7962
rect 3054 7955 3057 7983
rect 3084 7955 3087 7979
rect 3111 7955 3114 7987
rect 3128 7986 3131 7992
rect 3151 7987 3154 7993
rect 3163 7988 3166 7991
rect 3174 7991 3177 8005
rect 3210 8000 3213 8005
rect 3225 8007 3228 8017
rect 3255 8013 3258 8017
rect 3199 7996 3202 7999
rect 3751 8010 3827 8014
rect 3831 8010 3858 8014
rect 3862 8010 3880 8014
rect 3884 8010 3945 8014
rect 3949 8010 3963 8014
rect 3999 8007 4002 8017
rect 4029 8013 4032 8017
rect 4056 8013 4059 8017
rect 3241 7996 3244 7999
rect 3174 7988 3183 7991
rect 3210 7991 3213 7996
rect 3174 7983 3177 7988
rect 3126 7977 3131 7982
rect 3135 7955 3138 7983
rect 3217 7994 3229 7995
rect 3221 7992 3229 7994
rect 3241 7993 3249 7996
rect 3241 7987 3244 7993
rect 3253 7988 3256 7991
rect 3264 7991 3267 8005
rect 3870 8003 3873 8007
rect 3897 8003 3898 8007
rect 3942 8003 3944 8007
rect 3264 7988 3284 7991
rect 3165 7955 3168 7979
rect 3201 7955 3204 7987
rect 3264 7983 3267 7988
rect 3799 7983 3802 7986
rect 3810 7986 3813 7992
rect 3817 7986 3820 7992
rect 3810 7983 3820 7986
rect 3225 7955 3228 7983
rect 3255 7955 3258 7979
rect 3810 7978 3813 7983
rect 3817 7978 3820 7983
rect 3826 7988 3829 7992
rect 3826 7984 3828 7988
rect 3832 7984 3834 7988
rect 3842 7987 3845 7992
rect 3870 7989 3873 7992
rect 3842 7985 3853 7987
rect 3826 7978 3829 7984
rect 3842 7983 3848 7985
rect 3842 7978 3845 7983
rect 3852 7983 3853 7985
rect 3871 7985 3873 7989
rect 3870 7978 3873 7985
rect 4015 7996 4018 7999
rect 3886 7988 3889 7992
rect 3896 7988 3899 7992
rect 3896 7984 3905 7988
rect 3917 7987 3920 7992
rect 3942 7988 3945 7992
rect 3886 7978 3889 7984
rect 3896 7978 3899 7984
rect 3917 7983 3918 7987
rect 3922 7983 3925 7986
rect 3944 7984 3945 7988
rect 3960 7987 3963 7992
rect 3992 7992 4003 7995
rect 4015 7993 4023 7996
rect 3917 7978 3920 7983
rect 3942 7978 3945 7984
rect 3992 7986 3995 7992
rect 4015 7987 4018 7993
rect 4027 7988 4030 7991
rect 4038 7991 4041 8005
rect 4065 8000 4068 8005
rect 4080 8007 4083 8017
rect 4110 8013 4113 8017
rect 4146 8013 4149 8017
rect 4049 7996 4050 7999
rect 4054 7996 4057 7999
rect 4096 7996 4099 7999
rect 4038 7988 4046 7991
rect 4065 7991 4068 7996
rect 3960 7978 3963 7983
rect 4038 7983 4041 7988
rect 4046 7984 4050 7988
rect 4073 7992 4084 7995
rect 4096 7993 4104 7996
rect 3990 7977 3995 7982
rect 3862 7965 3863 7969
rect 3887 7966 3888 7970
rect 3934 7965 3935 7969
rect 3739 7958 3815 7962
rect 3819 7958 3874 7962
rect 3878 7958 3899 7962
rect 3903 7958 3930 7962
rect 3934 7958 3963 7962
rect 3999 7955 4002 7983
rect 4029 7955 4032 7979
rect 4056 7955 4059 7987
rect 4073 7986 4076 7992
rect 4096 7987 4099 7993
rect 4108 7988 4111 7991
rect 4119 7991 4122 8005
rect 4155 8000 4158 8005
rect 4170 8007 4173 8017
rect 4200 8013 4203 8017
rect 4574 8015 4578 8024
rect 4590 8015 4594 8024
rect 4606 8015 4610 8024
rect 4622 8015 4626 8024
rect 4144 7996 4147 7999
rect 4186 7996 4189 7999
rect 4119 7988 4128 7991
rect 4155 7991 4158 7996
rect 4119 7983 4122 7988
rect 4071 7977 4076 7982
rect 4080 7955 4083 7983
rect 4162 7994 4174 7995
rect 4166 7992 4174 7994
rect 4186 7993 4194 7996
rect 4186 7987 4189 7993
rect 4198 7988 4201 7991
rect 4209 7991 4212 8005
rect 4328 7991 4377 7992
rect 4209 7988 4229 7991
rect 4110 7955 4113 7979
rect 4146 7955 4149 7987
rect 4209 7983 4212 7988
rect 4233 7987 4377 7991
rect 4170 7955 4173 7983
rect 4200 7955 4203 7979
rect 4626 7975 4627 8015
rect 4665 7975 4666 8034
rect 4582 7963 4586 7975
rect 4598 7972 4602 7975
rect 4614 7972 4618 7975
rect 4598 7968 4618 7972
rect 4637 7972 4641 7975
rect 4653 7972 4657 7975
rect 4637 7968 4657 7972
rect 4680 7974 4684 7975
rect 4708 7975 4709 8034
rect 4749 7975 4750 8034
rect 4816 8032 4829 8042
rect 4806 8022 4829 8032
rect 4796 8012 4829 8022
rect 4786 8002 4829 8012
rect 4696 7974 4700 7975
rect 4680 7972 4700 7974
rect 4721 7972 4741 7975
rect 4680 7970 4741 7972
rect 4774 7970 4829 8002
rect 2782 7951 2856 7955
rect 2860 7951 2862 7955
rect 2866 7951 2870 7955
rect 2874 7951 2888 7955
rect 2892 7951 2897 7955
rect 2901 7951 2906 7955
rect 2910 7951 2929 7955
rect 2933 7951 2963 7955
rect 2967 7951 2978 7955
rect 2982 7951 3006 7955
rect 3010 7951 3023 7955
rect 3027 7951 3047 7955
rect 3051 7951 3101 7955
rect 3108 7951 3128 7955
rect 3132 7951 3182 7955
rect 3186 7951 3218 7955
rect 3222 7951 3272 7955
rect 3727 7951 3801 7955
rect 3805 7951 3807 7955
rect 3811 7951 3815 7955
rect 3819 7951 3833 7955
rect 3837 7951 3842 7955
rect 3846 7951 3851 7955
rect 3855 7951 3874 7955
rect 3878 7951 3908 7955
rect 3912 7951 3923 7955
rect 3927 7951 3951 7955
rect 3955 7951 3968 7955
rect 3972 7951 3992 7955
rect 3996 7951 4046 7955
rect 4053 7951 4073 7955
rect 4077 7951 4127 7955
rect 4131 7951 4163 7955
rect 4167 7951 4217 7955
rect 2794 7944 2870 7948
rect 2874 7944 2929 7948
rect 2933 7944 2954 7948
rect 2958 7944 2985 7948
rect 2989 7944 3018 7948
rect 2917 7937 2918 7941
rect 2942 7936 2943 7940
rect 2989 7937 2990 7941
rect 2865 7923 2868 7928
rect 2872 7923 2875 7928
rect 2855 7920 2857 7923
rect 2865 7920 2875 7923
rect 2865 7914 2868 7920
rect 2872 7914 2875 7920
rect 2881 7922 2884 7928
rect 2897 7923 2900 7928
rect 2881 7918 2883 7922
rect 2887 7918 2889 7922
rect 2897 7921 2903 7923
rect 2907 7921 2908 7923
rect 2897 7919 2908 7921
rect 2925 7921 2928 7928
rect 2881 7914 2884 7918
rect 2897 7914 2900 7919
rect 2926 7917 2928 7921
rect 2925 7914 2928 7917
rect 2941 7922 2944 7928
rect 2951 7922 2954 7928
rect 2972 7923 2975 7928
rect 2951 7918 2960 7922
rect 2972 7919 2973 7923
rect 2977 7920 2980 7923
rect 2997 7922 3000 7928
rect 3015 7923 3018 7928
rect 3054 7929 3057 7951
rect 3135 7929 3138 7951
rect 3225 7929 3228 7951
rect 3739 7944 3815 7948
rect 3819 7944 3874 7948
rect 3878 7944 3899 7948
rect 3903 7944 3930 7948
rect 3934 7944 3963 7948
rect 3862 7937 3863 7941
rect 3887 7936 3888 7940
rect 3934 7937 3935 7941
rect 2941 7914 2944 7918
rect 2951 7914 2954 7918
rect 2972 7914 2975 7919
rect 2999 7918 3000 7922
rect 2997 7914 3000 7918
rect 3015 7914 3018 7919
rect 3045 7916 3050 7921
rect 3054 7917 3055 7920
rect 3070 7919 3073 7925
rect 3070 7916 3078 7919
rect 3125 7916 3130 7921
rect 3134 7917 3136 7920
rect 3151 7919 3154 7925
rect 3151 7916 3159 7919
rect 3218 7917 3226 7920
rect 3241 7919 3244 7925
rect 3810 7923 3813 7928
rect 3817 7923 3820 7928
rect 3800 7920 3802 7923
rect 3241 7916 3249 7919
rect 3810 7920 3820 7923
rect 3070 7913 3073 7916
rect 3151 7913 3154 7916
rect 3241 7913 3244 7916
rect 3810 7914 3813 7920
rect 2925 7899 2928 7903
rect 2952 7899 2953 7903
rect 2997 7899 2999 7903
rect 3817 7914 3820 7920
rect 3826 7922 3829 7928
rect 3842 7923 3845 7928
rect 3826 7918 3828 7922
rect 3832 7918 3834 7922
rect 3842 7921 3848 7923
rect 3852 7921 3853 7923
rect 3842 7919 3853 7921
rect 3870 7921 3873 7928
rect 3826 7914 3829 7918
rect 3842 7914 3845 7919
rect 3871 7917 3873 7921
rect 3870 7914 3873 7917
rect 3886 7922 3889 7928
rect 3896 7922 3899 7928
rect 3917 7923 3920 7928
rect 3896 7918 3905 7922
rect 3917 7919 3918 7923
rect 3922 7920 3925 7923
rect 3942 7922 3945 7928
rect 3960 7923 3963 7928
rect 3999 7929 4002 7951
rect 4080 7929 4083 7951
rect 4170 7929 4173 7951
rect 4386 7950 4572 7963
rect 4582 7959 4593 7963
rect 4605 7963 4618 7968
rect 4648 7965 4657 7968
rect 4691 7966 4829 7970
rect 4648 7963 4678 7965
rect 4582 7945 4586 7959
rect 4605 7956 4635 7963
rect 4598 7950 4635 7956
rect 4639 7950 4640 7963
rect 4648 7954 4659 7963
rect 4667 7954 4678 7963
rect 4648 7952 4678 7954
rect 4682 7952 4683 7965
rect 4598 7949 4618 7950
rect 4598 7945 4602 7949
rect 4614 7945 4618 7949
rect 4648 7945 4657 7952
rect 4691 7945 4700 7966
rect 4721 7952 4829 7966
rect 4721 7945 4741 7952
rect 3886 7914 3889 7918
rect 3896 7914 3899 7918
rect 3917 7914 3920 7919
rect 3944 7918 3945 7922
rect 3942 7914 3945 7918
rect 3960 7914 3963 7919
rect 3990 7916 3995 7921
rect 3999 7917 4000 7920
rect 4015 7919 4018 7925
rect 4015 7916 4023 7919
rect 4070 7916 4075 7921
rect 4079 7917 4081 7920
rect 4096 7919 4099 7925
rect 4096 7916 4104 7919
rect 4163 7917 4171 7920
rect 4186 7919 4189 7925
rect 4186 7916 4194 7919
rect 4015 7913 4018 7916
rect 4096 7913 4099 7916
rect 4186 7913 4189 7916
rect 343 7883 386 7893
rect 2806 7892 2882 7896
rect 2886 7892 2913 7896
rect 2917 7892 2935 7896
rect 2939 7892 3000 7896
rect 3004 7892 3018 7896
rect 3054 7889 3057 7905
rect 3135 7889 3138 7905
rect 3225 7889 3228 7905
rect 3870 7899 3873 7903
rect 3897 7899 3898 7903
rect 3942 7899 3944 7903
rect 3751 7892 3827 7896
rect 3831 7892 3858 7896
rect 3862 7892 3880 7896
rect 3884 7892 3945 7896
rect 3949 7892 3963 7896
rect 3999 7889 4002 7905
rect 4080 7889 4083 7905
rect 4170 7889 4173 7905
rect 4626 7889 4627 7945
rect 2770 7885 2855 7889
rect 2859 7885 2871 7889
rect 2875 7885 2889 7889
rect 2893 7885 2900 7889
rect 2904 7885 2906 7889
rect 2910 7885 2925 7889
rect 2929 7885 2962 7889
rect 2966 7885 2967 7889
rect 2971 7885 2979 7889
rect 2983 7885 3007 7889
rect 3011 7885 3023 7889
rect 3027 7885 3047 7889
rect 3051 7885 3101 7889
rect 3105 7885 3128 7889
rect 3132 7885 3218 7889
rect 3222 7885 3276 7889
rect 3715 7885 3800 7889
rect 3804 7885 3816 7889
rect 3820 7885 3834 7889
rect 3838 7885 3845 7889
rect 3849 7885 3851 7889
rect 3855 7885 3870 7889
rect 3874 7885 3907 7889
rect 3911 7885 3912 7889
rect 3916 7885 3924 7889
rect 3928 7885 3952 7889
rect 3956 7885 3968 7889
rect 3972 7885 3992 7889
rect 3996 7885 4046 7889
rect 4050 7885 4073 7889
rect 4077 7885 4163 7889
rect 4167 7885 4221 7889
rect 4574 7886 4578 7889
rect 4590 7886 4594 7889
rect 4606 7886 4610 7889
rect 4622 7886 4626 7889
rect 343 7873 376 7883
rect 2806 7878 2882 7882
rect 2886 7878 2913 7882
rect 2917 7878 2935 7882
rect 2939 7878 3000 7882
rect 3004 7878 3018 7882
rect 3054 7875 3057 7885
rect 3084 7881 3087 7885
rect 343 7863 366 7873
rect 2925 7871 2928 7875
rect 2952 7871 2953 7875
rect 2997 7871 2999 7875
rect 343 7853 356 7863
rect 343 7814 346 7853
rect 2854 7851 2857 7854
rect 2865 7854 2868 7860
rect 2872 7854 2875 7860
rect 2865 7851 2875 7854
rect 2865 7846 2868 7851
rect 2872 7846 2875 7851
rect 2881 7856 2884 7860
rect 2881 7852 2883 7856
rect 2887 7852 2889 7856
rect 2897 7855 2900 7860
rect 2925 7857 2928 7860
rect 2897 7853 2908 7855
rect 2881 7846 2884 7852
rect 2897 7851 2903 7853
rect 2897 7846 2900 7851
rect 2907 7851 2908 7853
rect 2926 7853 2928 7857
rect 2925 7846 2928 7853
rect 3751 7878 3827 7882
rect 3831 7878 3858 7882
rect 3862 7878 3880 7882
rect 3884 7878 3945 7882
rect 3949 7878 3963 7882
rect 3999 7875 4002 7885
rect 4029 7881 4032 7885
rect 3070 7864 3073 7867
rect 2941 7856 2944 7860
rect 2951 7856 2954 7860
rect 2951 7852 2960 7856
rect 2972 7855 2975 7860
rect 2997 7856 3000 7860
rect 2941 7846 2944 7852
rect 2951 7846 2954 7852
rect 2972 7851 2973 7855
rect 2977 7851 2980 7854
rect 2999 7852 3000 7856
rect 3015 7855 3018 7860
rect 3047 7860 3058 7863
rect 3070 7861 3078 7864
rect 2972 7846 2975 7851
rect 2997 7846 3000 7852
rect 3047 7854 3050 7860
rect 3070 7855 3073 7861
rect 3082 7856 3085 7859
rect 3093 7859 3096 7873
rect 3870 7871 3873 7875
rect 3897 7871 3898 7875
rect 3942 7871 3944 7875
rect 3101 7859 3106 7864
rect 3093 7856 3101 7859
rect 3015 7846 3018 7851
rect 3093 7851 3096 7856
rect 3799 7851 3802 7854
rect 3810 7854 3813 7860
rect 3817 7854 3820 7860
rect 3810 7851 3820 7854
rect 3045 7845 3050 7850
rect 2364 7830 2373 7834
rect 2377 7830 2409 7834
rect 2413 7830 2476 7834
rect 2480 7830 2505 7834
rect 2509 7830 2541 7834
rect 2545 7830 2608 7834
rect 2612 7830 2637 7834
rect 2641 7830 2673 7834
rect 2677 7830 2740 7834
rect 2744 7830 2824 7834
rect 2917 7833 2918 7837
rect 2942 7834 2943 7838
rect 2989 7833 2990 7837
rect 2364 7823 2397 7827
rect 2401 7823 2425 7827
rect 2429 7823 2455 7827
rect 2459 7823 2492 7827
rect 2496 7823 2529 7827
rect 2533 7823 2557 7827
rect 2561 7823 2587 7827
rect 2591 7823 2624 7827
rect 2628 7823 2661 7827
rect 2665 7823 2689 7827
rect 2693 7823 2719 7827
rect 2723 7823 2756 7827
rect 2760 7823 2764 7827
rect 2849 7826 2870 7830
rect 2874 7826 2879 7830
rect 2883 7826 2929 7830
rect 2933 7826 2954 7830
rect 2958 7826 2985 7830
rect 2989 7826 3018 7830
rect 3054 7823 3057 7851
rect 3084 7823 3087 7847
rect 3810 7846 3813 7851
rect 3817 7846 3820 7851
rect 3826 7856 3829 7860
rect 3826 7852 3828 7856
rect 3832 7852 3834 7856
rect 3842 7855 3845 7860
rect 3870 7857 3873 7860
rect 3842 7853 3853 7855
rect 3826 7846 3829 7852
rect 3842 7851 3848 7853
rect 3842 7846 3845 7851
rect 3852 7851 3853 7853
rect 3871 7853 3873 7857
rect 3870 7846 3873 7853
rect 4015 7864 4018 7867
rect 3886 7856 3889 7860
rect 3896 7856 3899 7860
rect 3896 7852 3905 7856
rect 3917 7855 3920 7860
rect 3942 7856 3945 7860
rect 3886 7846 3889 7852
rect 3896 7846 3899 7852
rect 3917 7851 3918 7855
rect 3922 7851 3925 7854
rect 3944 7852 3945 7856
rect 3960 7855 3963 7860
rect 3992 7860 4003 7863
rect 4015 7861 4023 7864
rect 3917 7846 3920 7851
rect 3942 7846 3945 7852
rect 3992 7854 3995 7860
rect 4015 7855 4018 7861
rect 4027 7856 4030 7859
rect 4038 7859 4041 7873
rect 4046 7859 4051 7864
rect 4038 7856 4046 7859
rect 3960 7846 3963 7851
rect 4038 7851 4041 7856
rect 3990 7845 3995 7850
rect 3309 7830 3318 7834
rect 3322 7830 3354 7834
rect 3358 7830 3421 7834
rect 3425 7830 3450 7834
rect 3454 7830 3486 7834
rect 3490 7830 3553 7834
rect 3557 7830 3582 7834
rect 3586 7830 3618 7834
rect 3622 7830 3685 7834
rect 3689 7830 3769 7834
rect 3862 7833 3863 7837
rect 3887 7834 3888 7838
rect 3934 7833 3935 7837
rect 3309 7823 3342 7827
rect 3346 7823 3370 7827
rect 3374 7823 3400 7827
rect 3404 7823 3437 7827
rect 3441 7823 3474 7827
rect 3478 7823 3502 7827
rect 3506 7823 3532 7827
rect 3536 7823 3569 7827
rect 3573 7823 3606 7827
rect 3610 7823 3634 7827
rect 3638 7823 3664 7827
rect 3668 7823 3701 7827
rect 3705 7823 3709 7827
rect 3794 7826 3815 7830
rect 3819 7826 3824 7830
rect 3828 7826 3874 7830
rect 3878 7826 3899 7830
rect 3903 7826 3930 7830
rect 3934 7826 3963 7830
rect 3999 7823 4002 7851
rect 4527 7854 4626 7886
rect 4641 7939 4653 7945
rect 4665 7857 4666 7945
rect 4684 7939 4696 7945
rect 4708 7857 4709 7945
rect 4725 7939 4737 7945
rect 4749 7857 4750 7945
rect 4774 7906 4829 7952
rect 4786 7896 4829 7906
rect 4796 7886 4829 7896
rect 4806 7876 4829 7886
rect 4816 7866 4829 7876
rect 4645 7854 4649 7857
rect 4661 7854 4670 7857
rect 4688 7854 4692 7857
rect 4704 7854 4713 7857
rect 4729 7854 4733 7857
rect 4745 7854 4754 7857
rect 4029 7823 4032 7847
rect 4527 7830 4754 7854
rect 4527 7828 4595 7830
rect 4527 7824 4529 7828
rect 4533 7824 4534 7828
rect 4538 7824 4539 7828
rect 4543 7824 4544 7828
rect 4548 7824 4549 7828
rect 4553 7824 4554 7828
rect 4558 7824 4559 7828
rect 4563 7824 4564 7828
rect 4568 7824 4569 7828
rect 4573 7824 4574 7828
rect 4578 7824 4579 7828
rect 4583 7824 4584 7828
rect 4588 7824 4589 7828
rect 4593 7824 4595 7828
rect 4826 7827 4829 7866
rect 5083 7827 5086 8081
rect 4826 7824 5086 7827
rect 4527 7823 4595 7824
rect 86 7811 346 7814
rect 2367 7813 2370 7823
rect 2388 7813 2391 7823
rect 2404 7813 2407 7823
rect 2418 7816 2423 7820
rect 2427 7816 2434 7820
rect 2446 7813 2449 7823
rect 2462 7813 2465 7823
rect 2483 7813 2486 7823
rect 2499 7813 2502 7823
rect 2520 7813 2523 7823
rect 2536 7813 2539 7823
rect 2550 7816 2555 7820
rect 2559 7816 2566 7820
rect 2578 7813 2581 7823
rect 2594 7813 2597 7823
rect 2615 7813 2618 7823
rect 2631 7813 2634 7823
rect 2652 7813 2655 7823
rect 2668 7813 2671 7823
rect 2682 7816 2687 7820
rect 2691 7816 2698 7820
rect 2710 7813 2713 7823
rect 2726 7813 2729 7823
rect 2747 7813 2750 7823
rect 2782 7819 2856 7823
rect 2860 7819 2862 7823
rect 2866 7819 2870 7823
rect 2874 7819 2888 7823
rect 2892 7819 2897 7823
rect 2901 7819 2906 7823
rect 2910 7819 2929 7823
rect 2933 7819 2963 7823
rect 2967 7819 2978 7823
rect 2982 7819 3006 7823
rect 3010 7819 3023 7823
rect 3027 7819 3047 7823
rect 3051 7819 3131 7823
rect 3135 7819 3149 7823
rect 3153 7819 3158 7823
rect 3162 7819 3167 7823
rect 3171 7819 3190 7823
rect 3194 7819 3224 7823
rect 3228 7819 3239 7823
rect 3243 7819 3267 7823
rect 3271 7819 3280 7823
rect 2384 7799 2389 7802
rect 2393 7799 2417 7802
rect 2442 7799 2449 7802
rect 2453 7799 2475 7802
rect 2495 7799 2502 7802
rect 2516 7799 2521 7802
rect 2525 7799 2549 7802
rect 2574 7799 2581 7802
rect 2585 7799 2607 7802
rect 2627 7799 2634 7802
rect 2648 7799 2653 7802
rect 2657 7799 2681 7802
rect 2794 7812 2870 7816
rect 2874 7812 2879 7816
rect 2883 7812 2929 7816
rect 2933 7812 2954 7816
rect 2958 7812 2985 7816
rect 2989 7812 3018 7816
rect 2706 7799 2713 7802
rect 2717 7799 2739 7802
rect 2917 7805 2918 7809
rect 2942 7804 2943 7808
rect 2989 7805 2990 7809
rect 2400 7789 2407 7792
rect 2411 7793 2430 7796
rect 2430 7786 2433 7792
rect 2458 7789 2465 7792
rect 2469 7793 2484 7796
rect 2532 7789 2539 7792
rect 2543 7793 2562 7796
rect 2562 7786 2565 7792
rect 2590 7789 2597 7792
rect 2601 7793 2616 7796
rect 2664 7789 2671 7792
rect 2675 7793 2694 7796
rect 2694 7786 2697 7792
rect 2722 7789 2729 7792
rect 2733 7793 2750 7796
rect 2865 7791 2868 7796
rect 2872 7791 2875 7796
rect 2855 7788 2857 7791
rect 2865 7788 2875 7791
rect 2865 7782 2868 7788
rect 617 7776 618 7780
rect 622 7776 623 7780
rect 627 7776 628 7780
rect 632 7776 633 7780
rect 637 7776 638 7780
rect 642 7776 643 7780
rect 613 7775 647 7776
rect 617 7771 618 7775
rect 622 7771 623 7775
rect 627 7771 628 7775
rect 632 7771 633 7775
rect 637 7771 638 7775
rect 642 7771 643 7775
rect 613 7770 647 7771
rect 617 7766 618 7770
rect 622 7766 623 7770
rect 627 7766 628 7770
rect 632 7766 633 7770
rect 637 7766 638 7770
rect 642 7766 643 7770
rect 613 7765 647 7766
rect 86 7759 346 7762
rect 617 7761 618 7765
rect 622 7761 623 7765
rect 627 7761 628 7765
rect 632 7761 633 7765
rect 637 7761 638 7765
rect 642 7761 643 7765
rect 663 7776 664 7780
rect 668 7776 669 7780
rect 673 7776 674 7780
rect 678 7776 679 7780
rect 683 7776 684 7780
rect 688 7776 689 7780
rect 659 7775 693 7776
rect 663 7771 664 7775
rect 668 7771 669 7775
rect 673 7771 674 7775
rect 678 7771 679 7775
rect 683 7771 684 7775
rect 688 7771 689 7775
rect 659 7770 693 7771
rect 2367 7770 2370 7782
rect 2388 7770 2391 7782
rect 2404 7770 2407 7782
rect 2418 7773 2430 7776
rect 2446 7770 2449 7782
rect 2462 7770 2465 7782
rect 2483 7770 2486 7782
rect 2499 7770 2502 7782
rect 2520 7770 2523 7782
rect 2536 7770 2539 7782
rect 2550 7773 2562 7776
rect 2578 7770 2581 7782
rect 2594 7770 2597 7782
rect 2615 7770 2618 7782
rect 2631 7770 2634 7782
rect 2652 7770 2655 7782
rect 2668 7770 2671 7782
rect 2682 7773 2694 7776
rect 2710 7770 2713 7782
rect 2726 7770 2729 7782
rect 2747 7770 2750 7782
rect 2872 7782 2875 7788
rect 2881 7790 2884 7796
rect 2897 7791 2900 7796
rect 2881 7786 2883 7790
rect 2887 7786 2889 7790
rect 2897 7789 2903 7791
rect 2907 7789 2908 7791
rect 2897 7787 2908 7789
rect 2925 7789 2928 7796
rect 2881 7782 2884 7786
rect 2897 7782 2900 7787
rect 2926 7785 2928 7789
rect 2925 7782 2928 7785
rect 2941 7790 2944 7796
rect 2951 7790 2954 7796
rect 2972 7791 2975 7796
rect 2951 7786 2960 7790
rect 2972 7787 2973 7791
rect 2977 7788 2980 7791
rect 2997 7790 3000 7796
rect 3015 7791 3018 7796
rect 3054 7793 3057 7819
rect 3090 7812 3109 7816
rect 3113 7812 3131 7816
rect 3135 7812 3190 7816
rect 3194 7812 3215 7816
rect 3219 7812 3246 7816
rect 3250 7812 3279 7816
rect 3312 7813 3315 7823
rect 3333 7813 3336 7823
rect 3349 7813 3352 7823
rect 3363 7816 3368 7820
rect 3372 7816 3379 7820
rect 3391 7813 3394 7823
rect 3407 7813 3410 7823
rect 3428 7813 3431 7823
rect 3444 7813 3447 7823
rect 3465 7813 3468 7823
rect 3481 7813 3484 7823
rect 3495 7816 3500 7820
rect 3504 7816 3511 7820
rect 3523 7813 3526 7823
rect 3539 7813 3542 7823
rect 3560 7813 3563 7823
rect 3576 7813 3579 7823
rect 3597 7813 3600 7823
rect 3613 7813 3616 7823
rect 3627 7816 3632 7820
rect 3636 7816 3643 7820
rect 3655 7813 3658 7823
rect 3671 7813 3674 7823
rect 3692 7813 3695 7823
rect 3727 7819 3801 7823
rect 3805 7819 3807 7823
rect 3811 7819 3815 7823
rect 3819 7819 3833 7823
rect 3837 7819 3842 7823
rect 3846 7819 3851 7823
rect 3855 7819 3874 7823
rect 3878 7819 3908 7823
rect 3912 7819 3923 7823
rect 3927 7819 3951 7823
rect 3955 7819 3968 7823
rect 3972 7819 3992 7823
rect 3996 7819 4076 7823
rect 4080 7819 4094 7823
rect 4098 7819 4103 7823
rect 4107 7819 4112 7823
rect 4116 7819 4135 7823
rect 4139 7819 4169 7823
rect 4173 7819 4184 7823
rect 4188 7819 4212 7823
rect 4216 7819 4225 7823
rect 4527 7819 4529 7823
rect 4533 7819 4534 7823
rect 4538 7819 4539 7823
rect 4543 7819 4544 7823
rect 4548 7819 4549 7823
rect 4553 7819 4554 7823
rect 4558 7819 4559 7823
rect 4563 7819 4564 7823
rect 4568 7819 4569 7823
rect 4573 7819 4574 7823
rect 4578 7819 4579 7823
rect 4583 7819 4584 7823
rect 4588 7819 4589 7823
rect 4593 7819 4595 7823
rect 3090 7800 3093 7812
rect 3178 7805 3179 7809
rect 3203 7804 3204 7808
rect 3250 7805 3251 7809
rect 2941 7782 2944 7786
rect 2951 7782 2954 7786
rect 2972 7782 2975 7787
rect 2999 7786 3000 7790
rect 3117 7791 3120 7796
rect 3126 7791 3129 7796
rect 3133 7791 3136 7796
rect 2997 7782 3000 7786
rect 3015 7782 3018 7787
rect 3044 7780 3049 7785
rect 3053 7781 3055 7784
rect 3070 7783 3073 7789
rect 3102 7788 3136 7791
rect 3070 7780 3078 7783
rect 3070 7777 3073 7780
rect 663 7766 664 7770
rect 668 7766 669 7770
rect 673 7766 674 7770
rect 678 7766 679 7770
rect 683 7766 684 7770
rect 688 7766 689 7770
rect 2364 7766 2397 7770
rect 2401 7766 2425 7770
rect 2429 7766 2455 7770
rect 2459 7766 2529 7770
rect 2533 7766 2557 7770
rect 2561 7766 2587 7770
rect 2591 7766 2661 7770
rect 2665 7766 2689 7770
rect 2693 7766 2719 7770
rect 2723 7766 2776 7770
rect 2925 7767 2928 7771
rect 2952 7767 2953 7771
rect 2997 7767 2999 7771
rect 3102 7774 3105 7788
rect 3126 7782 3129 7788
rect 3133 7782 3136 7788
rect 3142 7790 3145 7796
rect 3158 7791 3161 7796
rect 3142 7786 3144 7790
rect 3148 7786 3150 7790
rect 3158 7789 3164 7791
rect 3168 7789 3169 7791
rect 3158 7787 3169 7789
rect 3186 7789 3189 7796
rect 3142 7782 3145 7786
rect 3158 7782 3161 7787
rect 3187 7785 3189 7789
rect 3186 7782 3189 7785
rect 3329 7799 3334 7802
rect 3338 7799 3362 7802
rect 3387 7799 3394 7802
rect 3398 7799 3420 7802
rect 3440 7799 3447 7802
rect 3461 7799 3466 7802
rect 3470 7799 3494 7802
rect 3519 7799 3526 7802
rect 3530 7799 3552 7802
rect 3572 7799 3579 7802
rect 3593 7799 3598 7802
rect 3602 7799 3626 7802
rect 3739 7812 3815 7816
rect 3819 7812 3824 7816
rect 3828 7812 3874 7816
rect 3878 7812 3899 7816
rect 3903 7812 3930 7816
rect 3934 7812 3963 7816
rect 3651 7799 3658 7802
rect 3662 7799 3684 7802
rect 3862 7805 3863 7809
rect 3887 7804 3888 7808
rect 3934 7805 3935 7809
rect 3202 7790 3205 7796
rect 3212 7790 3215 7796
rect 3233 7791 3236 7796
rect 3212 7786 3221 7790
rect 3233 7787 3234 7791
rect 3238 7788 3241 7791
rect 3258 7790 3261 7796
rect 3276 7791 3279 7796
rect 3202 7782 3205 7786
rect 3212 7782 3215 7786
rect 3233 7782 3236 7787
rect 3260 7786 3261 7790
rect 3258 7782 3261 7786
rect 3276 7782 3279 7787
rect 3345 7789 3352 7792
rect 3356 7793 3375 7796
rect 3375 7786 3378 7792
rect 3403 7789 3410 7792
rect 3414 7793 3429 7796
rect 3477 7789 3484 7792
rect 3488 7793 3507 7796
rect 3507 7786 3510 7792
rect 3535 7789 3542 7792
rect 3546 7793 3561 7796
rect 3609 7789 3616 7792
rect 3620 7793 3639 7796
rect 3639 7786 3642 7792
rect 3667 7789 3674 7792
rect 3678 7793 3695 7796
rect 3810 7791 3813 7796
rect 3817 7791 3820 7796
rect 3800 7788 3802 7791
rect 3810 7788 3820 7791
rect 3810 7782 3813 7788
rect 659 7765 693 7766
rect 663 7761 664 7765
rect 668 7761 669 7765
rect 673 7761 674 7765
rect 678 7761 679 7765
rect 683 7761 684 7765
rect 688 7761 689 7765
rect 2364 7759 2373 7763
rect 2377 7759 2424 7763
rect 2428 7759 2474 7763
rect 2478 7759 2505 7763
rect 2509 7759 2556 7763
rect 2560 7759 2606 7763
rect 2610 7759 2637 7763
rect 2641 7759 2688 7763
rect 2692 7759 2738 7763
rect 2742 7760 2812 7763
rect 2868 7760 2882 7764
rect 2886 7760 2913 7764
rect 2917 7760 2935 7764
rect 2939 7760 3000 7764
rect 3004 7760 3018 7764
rect 86 7505 89 7759
rect 343 7720 346 7759
rect 3054 7757 3057 7769
rect 3186 7767 3189 7771
rect 3213 7767 3214 7771
rect 3258 7767 3260 7771
rect 3312 7770 3315 7782
rect 3333 7770 3336 7782
rect 3349 7770 3352 7782
rect 3363 7773 3375 7776
rect 3391 7770 3394 7782
rect 3407 7770 3410 7782
rect 3428 7770 3431 7782
rect 3444 7770 3447 7782
rect 3465 7770 3468 7782
rect 3481 7770 3484 7782
rect 3495 7773 3507 7776
rect 3523 7770 3526 7782
rect 3539 7770 3542 7782
rect 3560 7770 3563 7782
rect 3576 7770 3579 7782
rect 3597 7770 3600 7782
rect 3613 7770 3616 7782
rect 3627 7773 3639 7776
rect 3655 7770 3658 7782
rect 3671 7770 3674 7782
rect 3692 7770 3695 7782
rect 3817 7782 3820 7788
rect 3826 7790 3829 7796
rect 3842 7791 3845 7796
rect 3826 7786 3828 7790
rect 3832 7786 3834 7790
rect 3842 7789 3848 7791
rect 3852 7789 3853 7791
rect 3842 7787 3853 7789
rect 3870 7789 3873 7796
rect 3826 7782 3829 7786
rect 3842 7782 3845 7787
rect 3871 7785 3873 7789
rect 3870 7782 3873 7785
rect 3886 7790 3889 7796
rect 3896 7790 3899 7796
rect 3917 7791 3920 7796
rect 3896 7786 3905 7790
rect 3917 7787 3918 7791
rect 3922 7788 3925 7791
rect 3942 7790 3945 7796
rect 3960 7791 3963 7796
rect 3999 7793 4002 7819
rect 4527 7818 4595 7819
rect 4035 7812 4054 7816
rect 4058 7812 4076 7816
rect 4080 7812 4135 7816
rect 4139 7812 4160 7816
rect 4164 7812 4191 7816
rect 4195 7812 4224 7816
rect 4035 7800 4038 7812
rect 4123 7805 4124 7809
rect 4148 7804 4149 7808
rect 4195 7805 4196 7809
rect 3886 7782 3889 7786
rect 3896 7782 3899 7786
rect 3917 7782 3920 7787
rect 3944 7786 3945 7790
rect 4062 7791 4065 7796
rect 4071 7791 4074 7796
rect 4078 7791 4081 7796
rect 3942 7782 3945 7786
rect 3960 7782 3963 7787
rect 3989 7780 3994 7785
rect 3998 7781 4000 7784
rect 4015 7783 4018 7789
rect 4047 7788 4081 7791
rect 4015 7780 4023 7783
rect 4015 7777 4018 7780
rect 3309 7766 3342 7770
rect 3346 7766 3370 7770
rect 3374 7766 3400 7770
rect 3404 7766 3474 7770
rect 3478 7766 3502 7770
rect 3506 7766 3532 7770
rect 3536 7766 3606 7770
rect 3610 7766 3634 7770
rect 3638 7766 3664 7770
rect 3668 7766 3721 7770
rect 3870 7767 3873 7771
rect 3897 7767 3898 7771
rect 3942 7767 3944 7771
rect 4047 7774 4050 7788
rect 4071 7782 4074 7788
rect 4078 7782 4081 7788
rect 4087 7790 4090 7796
rect 4103 7791 4106 7796
rect 4087 7786 4089 7790
rect 4093 7786 4095 7790
rect 4103 7789 4109 7791
rect 4113 7789 4114 7791
rect 4103 7787 4114 7789
rect 4131 7789 4134 7796
rect 4087 7782 4090 7786
rect 4103 7782 4106 7787
rect 4132 7785 4134 7789
rect 4131 7782 4134 7785
rect 4147 7790 4150 7796
rect 4157 7790 4160 7796
rect 4178 7791 4181 7796
rect 4157 7786 4166 7790
rect 4178 7787 4179 7791
rect 4183 7788 4186 7791
rect 4203 7790 4206 7796
rect 4221 7791 4224 7796
rect 4147 7782 4150 7786
rect 4157 7782 4160 7786
rect 4178 7782 4181 7787
rect 4205 7786 4206 7790
rect 4483 7789 4484 7793
rect 4488 7789 4489 7793
rect 4493 7789 4494 7793
rect 4498 7789 4499 7793
rect 4503 7789 4504 7793
rect 4508 7789 4509 7793
rect 4479 7788 4513 7789
rect 4203 7782 4206 7786
rect 4221 7782 4224 7787
rect 4483 7784 4484 7788
rect 4488 7784 4489 7788
rect 4493 7784 4494 7788
rect 4498 7784 4499 7788
rect 4503 7784 4504 7788
rect 4508 7784 4509 7788
rect 4479 7783 4513 7784
rect 4483 7779 4484 7783
rect 4488 7779 4489 7783
rect 4493 7779 4494 7783
rect 4498 7779 4499 7783
rect 4503 7779 4504 7783
rect 4508 7779 4509 7783
rect 4479 7778 4513 7779
rect 4483 7774 4484 7778
rect 4488 7774 4489 7778
rect 4493 7774 4494 7778
rect 4498 7774 4499 7778
rect 4503 7774 4504 7778
rect 4508 7774 4509 7778
rect 4529 7789 4530 7793
rect 4534 7789 4535 7793
rect 4539 7789 4540 7793
rect 4544 7789 4545 7793
rect 4549 7789 4550 7793
rect 4554 7789 4555 7793
rect 4525 7788 4559 7789
rect 4529 7784 4530 7788
rect 4534 7784 4535 7788
rect 4539 7784 4540 7788
rect 4544 7784 4545 7788
rect 4549 7784 4550 7788
rect 4554 7784 4555 7788
rect 4525 7783 4559 7784
rect 4529 7779 4530 7783
rect 4534 7779 4535 7783
rect 4539 7779 4540 7783
rect 4544 7779 4545 7783
rect 4549 7779 4550 7783
rect 4554 7779 4555 7783
rect 4525 7778 4559 7779
rect 4529 7774 4530 7778
rect 4534 7774 4535 7778
rect 4539 7774 4540 7778
rect 4544 7774 4545 7778
rect 4549 7774 4550 7778
rect 4554 7774 4555 7778
rect 3094 7760 3099 7764
rect 3103 7760 3143 7764
rect 3147 7760 3174 7764
rect 3178 7760 3196 7764
rect 3200 7760 3261 7764
rect 3265 7760 3279 7764
rect 3309 7759 3318 7763
rect 3322 7759 3369 7763
rect 3373 7759 3419 7763
rect 3423 7759 3450 7763
rect 3454 7759 3501 7763
rect 3505 7759 3551 7763
rect 3555 7759 3582 7763
rect 3586 7759 3633 7763
rect 3637 7759 3683 7763
rect 3687 7760 3757 7763
rect 3813 7760 3827 7764
rect 3831 7760 3858 7764
rect 3862 7760 3880 7764
rect 3884 7760 3945 7764
rect 3949 7760 3963 7764
rect 3999 7757 4002 7769
rect 4131 7767 4134 7771
rect 4158 7767 4159 7771
rect 4203 7767 4205 7771
rect 4826 7772 5086 7775
rect 4039 7760 4044 7764
rect 4048 7760 4088 7764
rect 4092 7760 4119 7764
rect 4123 7760 4141 7764
rect 4145 7760 4206 7764
rect 4210 7760 4224 7764
rect 2371 7753 2755 7756
rect 2770 7753 2855 7757
rect 2859 7753 2871 7757
rect 2875 7753 2889 7757
rect 2893 7753 2900 7757
rect 2904 7753 2906 7757
rect 2910 7753 2925 7757
rect 2929 7753 2962 7757
rect 2966 7753 2967 7757
rect 2971 7753 2979 7757
rect 2983 7753 3007 7757
rect 3011 7753 3047 7757
rect 3051 7753 3090 7757
rect 3094 7753 3101 7757
rect 3105 7753 3116 7757
rect 3120 7753 3132 7757
rect 3136 7753 3150 7757
rect 3154 7753 3161 7757
rect 3165 7753 3167 7757
rect 3171 7753 3186 7757
rect 3190 7753 3223 7757
rect 3227 7753 3228 7757
rect 3232 7753 3240 7757
rect 3244 7753 3268 7757
rect 3272 7753 3280 7757
rect 3316 7753 3700 7756
rect 3715 7753 3800 7757
rect 3804 7753 3816 7757
rect 3820 7753 3834 7757
rect 3838 7753 3845 7757
rect 3849 7753 3851 7757
rect 3855 7753 3870 7757
rect 3874 7753 3907 7757
rect 3911 7753 3912 7757
rect 3916 7753 3924 7757
rect 3928 7753 3952 7757
rect 3956 7753 3992 7757
rect 3996 7753 4035 7757
rect 4039 7753 4046 7757
rect 4050 7753 4061 7757
rect 4065 7753 4077 7757
rect 4081 7753 4095 7757
rect 4099 7753 4106 7757
rect 4110 7753 4112 7757
rect 4116 7753 4131 7757
rect 4135 7753 4168 7757
rect 4172 7753 4173 7757
rect 4177 7753 4185 7757
rect 4189 7753 4213 7757
rect 4217 7753 4225 7757
rect 2514 7746 2623 7749
rect 2806 7746 2864 7750
rect 2868 7746 3098 7749
rect 3288 7747 3296 7751
rect 3459 7746 3568 7749
rect 3751 7746 3809 7750
rect 3813 7746 4043 7749
rect 4233 7747 4241 7751
rect 2494 7738 2498 7742
rect 2502 7738 2506 7742
rect 2794 7739 3108 7742
rect 2842 7732 3115 7736
rect 3284 7729 3288 7735
rect 3439 7738 3443 7742
rect 3447 7738 3451 7742
rect 3739 7739 4053 7742
rect 3787 7732 4058 7736
rect 4229 7729 4233 7735
rect 4826 7733 4829 7772
rect 2350 7725 2482 7729
rect 2486 7725 2502 7729
rect 2518 7725 3427 7729
rect 3431 7725 3447 7729
rect 3463 7725 4321 7729
rect 4816 7723 4829 7733
rect 343 7710 356 7720
rect 2510 7718 2755 7721
rect 2830 7718 3156 7722
rect 3160 7718 3192 7722
rect 3196 7718 3259 7722
rect 3263 7718 3279 7722
rect 3455 7718 3700 7721
rect 3775 7718 4101 7722
rect 4105 7718 4137 7722
rect 4141 7718 4204 7722
rect 4208 7718 4224 7722
rect 2525 7711 2755 7714
rect 2770 7711 3142 7715
rect 3146 7711 3180 7715
rect 3184 7711 3208 7715
rect 3212 7711 3238 7715
rect 3242 7711 3275 7715
rect 343 7700 366 7710
rect 2494 7702 2498 7706
rect 2502 7702 2506 7706
rect 3150 7701 3153 7711
rect 3171 7701 3174 7711
rect 3187 7701 3190 7711
rect 3201 7704 3206 7708
rect 3210 7704 3217 7708
rect 3229 7701 3232 7711
rect 3245 7701 3248 7711
rect 3266 7701 3269 7711
rect 3470 7711 3700 7714
rect 3715 7711 4087 7715
rect 4091 7711 4125 7715
rect 4129 7711 4153 7715
rect 4157 7711 4183 7715
rect 4187 7711 4220 7715
rect 4806 7713 4829 7723
rect 3439 7702 3443 7706
rect 3447 7702 3451 7706
rect 4095 7701 4098 7711
rect 4116 7701 4119 7711
rect 4132 7701 4135 7711
rect 4146 7704 4151 7708
rect 4155 7704 4162 7708
rect 4174 7701 4177 7711
rect 4190 7701 4193 7711
rect 4211 7701 4214 7711
rect 4796 7703 4829 7713
rect 343 7690 376 7700
rect 2514 7695 2624 7698
rect 343 7680 386 7690
rect 2364 7688 2373 7692
rect 2377 7688 2409 7692
rect 2413 7688 2476 7692
rect 2480 7688 2505 7692
rect 2509 7688 2541 7692
rect 2545 7688 2608 7692
rect 2612 7688 2637 7692
rect 2641 7688 2673 7692
rect 2677 7688 2740 7692
rect 2744 7688 2824 7692
rect 2364 7681 2397 7685
rect 2401 7681 2425 7685
rect 2429 7681 2455 7685
rect 2459 7681 2492 7685
rect 2496 7681 2529 7685
rect 2533 7681 2557 7685
rect 2561 7681 2587 7685
rect 2591 7681 2624 7685
rect 2628 7681 2661 7685
rect 2665 7681 2689 7685
rect 2693 7681 2719 7685
rect 2723 7681 2756 7685
rect 2760 7681 2764 7685
rect 3167 7687 3172 7690
rect 3176 7687 3200 7690
rect 3459 7695 3569 7698
rect 3225 7687 3232 7690
rect 3236 7687 3258 7690
rect 3309 7688 3318 7692
rect 3322 7688 3354 7692
rect 3358 7688 3421 7692
rect 3425 7688 3450 7692
rect 3454 7688 3486 7692
rect 3490 7688 3553 7692
rect 3557 7688 3582 7692
rect 3586 7688 3618 7692
rect 3622 7688 3685 7692
rect 3689 7688 3769 7692
rect 343 7584 769 7680
rect 2367 7671 2370 7681
rect 2388 7671 2391 7681
rect 2404 7671 2407 7681
rect 2418 7674 2423 7678
rect 2427 7674 2434 7678
rect 2446 7671 2449 7681
rect 2462 7671 2465 7681
rect 2483 7671 2486 7681
rect 2499 7671 2502 7681
rect 2520 7671 2523 7681
rect 2536 7671 2539 7681
rect 2550 7674 2555 7678
rect 2559 7674 2566 7678
rect 2578 7671 2581 7681
rect 2594 7671 2597 7681
rect 2615 7671 2618 7681
rect 2631 7671 2634 7681
rect 2652 7671 2655 7681
rect 2668 7671 2671 7681
rect 2682 7674 2687 7678
rect 2691 7674 2698 7678
rect 2710 7671 2713 7681
rect 2726 7671 2729 7681
rect 2747 7671 2750 7681
rect 3183 7677 3190 7680
rect 3194 7681 3213 7684
rect 2384 7657 2389 7660
rect 2393 7657 2417 7660
rect 2442 7657 2449 7660
rect 2453 7657 2475 7660
rect 2495 7657 2502 7660
rect 2516 7657 2521 7660
rect 2525 7657 2549 7660
rect 2574 7657 2581 7660
rect 2585 7657 2607 7660
rect 2627 7657 2634 7660
rect 2648 7657 2653 7660
rect 2657 7657 2681 7660
rect 2706 7657 2713 7660
rect 2717 7657 2739 7660
rect 3213 7674 3216 7680
rect 3241 7677 3248 7680
rect 3252 7681 3267 7684
rect 3309 7681 3342 7685
rect 3346 7681 3370 7685
rect 3374 7681 3400 7685
rect 3404 7681 3437 7685
rect 3441 7681 3474 7685
rect 3478 7681 3502 7685
rect 3506 7681 3532 7685
rect 3536 7681 3569 7685
rect 3573 7681 3606 7685
rect 3610 7681 3634 7685
rect 3638 7681 3664 7685
rect 3668 7681 3701 7685
rect 3705 7681 3709 7685
rect 4112 7687 4117 7690
rect 4121 7687 4145 7690
rect 4786 7693 4829 7703
rect 4170 7687 4177 7690
rect 4181 7687 4203 7690
rect 3312 7671 3315 7681
rect 3333 7671 3336 7681
rect 3349 7671 3352 7681
rect 3363 7674 3368 7678
rect 3372 7674 3379 7678
rect 3391 7671 3394 7681
rect 3407 7671 3410 7681
rect 3428 7671 3431 7681
rect 3444 7671 3447 7681
rect 3465 7671 3468 7681
rect 3481 7671 3484 7681
rect 3495 7674 3500 7678
rect 3504 7674 3511 7678
rect 3523 7671 3526 7681
rect 3539 7671 3542 7681
rect 3560 7671 3563 7681
rect 3576 7671 3579 7681
rect 3597 7671 3600 7681
rect 3613 7671 3616 7681
rect 3627 7674 3632 7678
rect 3636 7674 3643 7678
rect 3655 7671 3658 7681
rect 3671 7671 3674 7681
rect 3692 7671 3695 7681
rect 4128 7677 4135 7680
rect 4139 7681 4158 7684
rect 3150 7658 3153 7670
rect 3171 7658 3174 7670
rect 3187 7658 3190 7670
rect 3201 7661 3213 7664
rect 3229 7658 3232 7670
rect 3245 7658 3248 7670
rect 3266 7658 3269 7670
rect 2400 7647 2407 7650
rect 2411 7651 2430 7654
rect 2430 7644 2433 7650
rect 2458 7647 2465 7650
rect 2469 7651 2484 7654
rect 2532 7647 2539 7650
rect 2543 7651 2562 7654
rect 2562 7644 2565 7650
rect 2590 7647 2597 7650
rect 2601 7651 2616 7654
rect 2664 7647 2671 7650
rect 2675 7651 2694 7654
rect 2694 7644 2697 7650
rect 2722 7647 2729 7650
rect 2733 7651 2750 7654
rect 2782 7654 3180 7658
rect 3184 7654 3208 7658
rect 3212 7654 3238 7658
rect 3242 7654 3279 7658
rect 3329 7657 3334 7660
rect 3338 7657 3362 7660
rect 3387 7657 3394 7660
rect 3398 7657 3420 7660
rect 3440 7657 3447 7660
rect 3461 7657 3466 7660
rect 3470 7657 3494 7660
rect 3519 7657 3526 7660
rect 3530 7657 3552 7660
rect 3572 7657 3579 7660
rect 3593 7657 3598 7660
rect 3602 7657 3626 7660
rect 3651 7657 3658 7660
rect 3662 7657 3684 7660
rect 4158 7674 4161 7680
rect 4186 7677 4193 7680
rect 4197 7681 4212 7684
rect 4095 7658 4098 7670
rect 4116 7658 4119 7670
rect 4132 7658 4135 7670
rect 4146 7661 4158 7664
rect 4174 7658 4177 7670
rect 4190 7658 4193 7670
rect 4211 7658 4214 7670
rect 2818 7647 3156 7651
rect 3160 7647 3207 7651
rect 3211 7647 3257 7651
rect 3261 7647 3279 7651
rect 3345 7647 3352 7650
rect 3356 7651 3375 7654
rect 2367 7628 2370 7640
rect 2388 7628 2391 7640
rect 2404 7628 2407 7640
rect 2418 7631 2430 7634
rect 2446 7628 2449 7640
rect 2462 7628 2465 7640
rect 2483 7628 2486 7640
rect 2499 7628 2502 7640
rect 2520 7628 2523 7640
rect 2536 7628 2539 7640
rect 2550 7631 2562 7634
rect 2578 7628 2581 7640
rect 2594 7628 2597 7640
rect 2615 7628 2618 7640
rect 2631 7628 2634 7640
rect 2652 7628 2655 7640
rect 2668 7628 2671 7640
rect 2682 7631 2694 7634
rect 2710 7628 2713 7640
rect 2726 7628 2729 7640
rect 2747 7628 2750 7640
rect 3153 7640 3274 7643
rect 3375 7644 3378 7650
rect 3403 7647 3410 7650
rect 3414 7651 3429 7654
rect 3477 7647 3484 7650
rect 3488 7651 3507 7654
rect 3507 7644 3510 7650
rect 3535 7647 3542 7650
rect 3546 7651 3561 7654
rect 3609 7647 3616 7650
rect 3620 7651 3639 7654
rect 3639 7644 3642 7650
rect 3667 7647 3674 7650
rect 3678 7651 3695 7654
rect 3727 7654 4125 7658
rect 4129 7654 4153 7658
rect 4157 7654 4183 7658
rect 4187 7654 4224 7658
rect 3763 7647 4101 7651
rect 4105 7647 4152 7651
rect 4156 7647 4202 7651
rect 4206 7647 4224 7651
rect 4403 7648 4829 7693
rect 2830 7632 3156 7636
rect 3160 7632 3192 7636
rect 3196 7632 3259 7636
rect 3263 7632 3279 7636
rect 2364 7624 2397 7628
rect 2401 7624 2425 7628
rect 2429 7624 2455 7628
rect 2459 7624 2529 7628
rect 2533 7624 2557 7628
rect 2561 7624 2587 7628
rect 2591 7624 2661 7628
rect 2665 7624 2689 7628
rect 2693 7624 2719 7628
rect 2723 7624 2776 7628
rect 3146 7625 3180 7629
rect 3184 7625 3208 7629
rect 3212 7625 3238 7629
rect 3242 7625 3275 7629
rect 3312 7628 3315 7640
rect 3333 7628 3336 7640
rect 3349 7628 3352 7640
rect 3363 7631 3375 7634
rect 3391 7628 3394 7640
rect 3407 7628 3410 7640
rect 3428 7628 3431 7640
rect 3444 7628 3447 7640
rect 3465 7628 3468 7640
rect 3481 7628 3484 7640
rect 3495 7631 3507 7634
rect 3523 7628 3526 7640
rect 3539 7628 3542 7640
rect 3560 7628 3563 7640
rect 3576 7628 3579 7640
rect 3597 7628 3600 7640
rect 3613 7628 3616 7640
rect 3627 7631 3639 7634
rect 3655 7628 3658 7640
rect 3671 7628 3674 7640
rect 3692 7628 3695 7640
rect 4098 7640 4219 7643
rect 3775 7632 4101 7636
rect 4105 7632 4137 7636
rect 4141 7632 4204 7636
rect 4208 7632 4224 7636
rect 4384 7635 4829 7648
rect 2364 7617 2373 7621
rect 2377 7617 2424 7621
rect 2428 7617 2474 7621
rect 2478 7617 2505 7621
rect 2509 7617 2556 7621
rect 2560 7617 2606 7621
rect 2610 7617 2637 7621
rect 2641 7617 2688 7621
rect 2692 7617 2738 7621
rect 2742 7617 2812 7621
rect 3150 7615 3153 7625
rect 3171 7615 3174 7625
rect 3187 7615 3190 7625
rect 3201 7618 3206 7622
rect 3210 7618 3217 7622
rect 3229 7615 3232 7625
rect 3245 7615 3248 7625
rect 3266 7615 3269 7625
rect 3309 7624 3342 7628
rect 3346 7624 3370 7628
rect 3374 7624 3400 7628
rect 3404 7624 3474 7628
rect 3478 7624 3502 7628
rect 3506 7624 3532 7628
rect 3536 7624 3606 7628
rect 3610 7624 3634 7628
rect 3638 7624 3664 7628
rect 3668 7624 3721 7628
rect 4091 7625 4125 7629
rect 4129 7625 4153 7629
rect 4157 7625 4183 7629
rect 4187 7625 4220 7629
rect 3309 7617 3318 7621
rect 3322 7617 3369 7621
rect 3373 7617 3419 7621
rect 3423 7617 3450 7621
rect 3454 7617 3501 7621
rect 3505 7617 3551 7621
rect 3555 7617 3582 7621
rect 3586 7617 3633 7621
rect 3637 7617 3683 7621
rect 3687 7617 3757 7621
rect 4095 7615 4098 7625
rect 4116 7615 4119 7625
rect 4132 7615 4135 7625
rect 4146 7618 4151 7622
rect 4155 7618 4162 7622
rect 4174 7615 4177 7625
rect 4190 7615 4193 7625
rect 4211 7615 4214 7625
rect 2370 7610 2755 7613
rect 2364 7602 2373 7606
rect 2377 7602 2409 7606
rect 2413 7602 2476 7606
rect 2480 7602 2505 7606
rect 2509 7602 2541 7606
rect 2545 7602 2608 7606
rect 2612 7602 2637 7606
rect 2641 7602 2673 7606
rect 2677 7602 2740 7606
rect 2744 7602 2824 7606
rect 2364 7595 2397 7599
rect 2401 7595 2425 7599
rect 2429 7595 2455 7599
rect 2459 7595 2492 7599
rect 2496 7595 2529 7599
rect 2533 7595 2557 7599
rect 2561 7595 2587 7599
rect 2591 7595 2624 7599
rect 2628 7595 2661 7599
rect 2665 7595 2689 7599
rect 2693 7595 2719 7599
rect 2723 7595 2756 7599
rect 2760 7595 2764 7599
rect 3167 7601 3172 7604
rect 3176 7601 3200 7604
rect 3315 7610 3700 7613
rect 3225 7601 3232 7604
rect 3236 7601 3258 7604
rect 3309 7602 3318 7606
rect 3322 7602 3354 7606
rect 3358 7602 3421 7606
rect 3425 7602 3450 7606
rect 3454 7602 3486 7606
rect 3490 7602 3553 7606
rect 3557 7602 3582 7606
rect 3586 7602 3618 7606
rect 3622 7602 3685 7606
rect 3689 7602 3769 7606
rect 2367 7585 2370 7595
rect 2388 7585 2391 7595
rect 2404 7585 2407 7595
rect 2418 7588 2423 7592
rect 2427 7588 2434 7592
rect 2446 7585 2449 7595
rect 2462 7585 2465 7595
rect 2483 7585 2486 7595
rect 2499 7585 2502 7595
rect 2520 7585 2523 7595
rect 2536 7585 2539 7595
rect 2550 7588 2555 7592
rect 2559 7588 2566 7592
rect 2578 7585 2581 7595
rect 2594 7585 2597 7595
rect 2615 7585 2618 7595
rect 2631 7585 2634 7595
rect 2652 7585 2655 7595
rect 2668 7585 2671 7595
rect 2682 7588 2687 7592
rect 2691 7588 2698 7592
rect 2710 7585 2713 7595
rect 2726 7585 2729 7595
rect 2747 7585 2750 7595
rect 3183 7591 3190 7594
rect 3194 7595 3213 7598
rect 343 7574 386 7584
rect 343 7564 376 7574
rect 2384 7571 2389 7574
rect 2393 7571 2417 7574
rect 2442 7571 2449 7574
rect 2453 7571 2475 7574
rect 2495 7571 2502 7574
rect 2516 7571 2521 7574
rect 2525 7571 2549 7574
rect 2574 7571 2581 7574
rect 2585 7571 2607 7574
rect 2627 7571 2634 7574
rect 2648 7571 2653 7574
rect 2657 7571 2681 7574
rect 2706 7571 2713 7574
rect 2717 7571 2739 7574
rect 3213 7588 3216 7594
rect 3241 7591 3248 7594
rect 3252 7595 3267 7598
rect 3278 7593 3289 7597
rect 3309 7595 3342 7599
rect 3346 7595 3370 7599
rect 3374 7595 3400 7599
rect 3404 7595 3437 7599
rect 3441 7595 3474 7599
rect 3478 7595 3502 7599
rect 3506 7595 3532 7599
rect 3536 7595 3569 7599
rect 3573 7595 3606 7599
rect 3610 7595 3634 7599
rect 3638 7595 3664 7599
rect 3668 7595 3701 7599
rect 3705 7595 3709 7599
rect 4112 7601 4117 7604
rect 4121 7601 4145 7604
rect 4170 7601 4177 7604
rect 4181 7601 4203 7604
rect 3312 7585 3315 7595
rect 3333 7585 3336 7595
rect 3349 7585 3352 7595
rect 3363 7588 3368 7592
rect 3372 7588 3379 7592
rect 3391 7585 3394 7595
rect 3407 7585 3410 7595
rect 3428 7585 3431 7595
rect 3444 7585 3447 7595
rect 3465 7585 3468 7595
rect 3481 7585 3484 7595
rect 3495 7588 3500 7592
rect 3504 7588 3511 7592
rect 3523 7585 3526 7595
rect 3539 7585 3542 7595
rect 3560 7585 3563 7595
rect 3576 7585 3579 7595
rect 3597 7585 3600 7595
rect 3613 7585 3616 7595
rect 3627 7588 3632 7592
rect 3636 7588 3643 7592
rect 3655 7585 3658 7595
rect 3671 7585 3674 7595
rect 3692 7585 3695 7595
rect 4128 7591 4135 7594
rect 4139 7595 4158 7598
rect 3150 7572 3153 7584
rect 3171 7572 3174 7584
rect 3187 7572 3190 7584
rect 3201 7575 3213 7578
rect 3229 7572 3232 7584
rect 3245 7572 3248 7584
rect 3266 7572 3269 7584
rect 343 7554 366 7564
rect 2400 7561 2407 7564
rect 2411 7565 2430 7568
rect 2430 7558 2433 7564
rect 2458 7561 2465 7564
rect 2469 7565 2484 7568
rect 2532 7561 2539 7564
rect 2543 7565 2562 7568
rect 2562 7558 2565 7564
rect 2590 7561 2597 7564
rect 2601 7565 2616 7568
rect 2664 7561 2671 7564
rect 2675 7565 2694 7568
rect 2694 7558 2697 7564
rect 2722 7561 2729 7564
rect 2733 7565 2750 7568
rect 2782 7568 3180 7572
rect 3184 7568 3208 7572
rect 3212 7568 3238 7572
rect 3242 7568 3279 7572
rect 3329 7571 3334 7574
rect 3338 7571 3362 7574
rect 3387 7571 3394 7574
rect 3398 7571 3420 7574
rect 3440 7571 3447 7574
rect 3461 7571 3466 7574
rect 3470 7571 3494 7574
rect 3519 7571 3526 7574
rect 3530 7571 3552 7574
rect 3572 7571 3579 7574
rect 3593 7571 3598 7574
rect 3602 7571 3626 7574
rect 3651 7571 3658 7574
rect 3662 7571 3684 7574
rect 4158 7588 4161 7594
rect 4186 7591 4193 7594
rect 4197 7595 4212 7598
rect 4403 7597 4829 7635
rect 4223 7593 4234 7597
rect 4786 7587 4829 7597
rect 4095 7572 4098 7584
rect 4116 7572 4119 7584
rect 4132 7572 4135 7584
rect 4146 7575 4158 7578
rect 4174 7572 4177 7584
rect 4190 7572 4193 7584
rect 4211 7572 4214 7584
rect 4796 7577 4829 7587
rect 2818 7561 3156 7565
rect 3160 7561 3207 7565
rect 3211 7561 3257 7565
rect 3261 7561 3279 7565
rect 3345 7561 3352 7564
rect 3356 7565 3375 7568
rect 3375 7558 3378 7564
rect 3403 7561 3410 7564
rect 3414 7565 3429 7568
rect 3477 7561 3484 7564
rect 3488 7565 3507 7568
rect 3507 7558 3510 7564
rect 3535 7561 3542 7564
rect 3546 7565 3561 7568
rect 3609 7561 3616 7564
rect 3620 7565 3639 7568
rect 3639 7558 3642 7564
rect 3667 7561 3674 7564
rect 3678 7565 3695 7568
rect 3727 7568 4125 7572
rect 4129 7568 4153 7572
rect 4157 7568 4183 7572
rect 4187 7568 4224 7572
rect 4806 7567 4829 7577
rect 3763 7561 4101 7565
rect 4105 7561 4152 7565
rect 4156 7561 4202 7565
rect 4206 7561 4224 7565
rect 4816 7557 4829 7567
rect 343 7544 356 7554
rect 343 7505 346 7544
rect 2367 7542 2370 7554
rect 2388 7542 2391 7554
rect 2404 7542 2407 7554
rect 2418 7545 2430 7548
rect 2446 7542 2449 7554
rect 2462 7542 2465 7554
rect 2483 7542 2486 7554
rect 2499 7542 2502 7554
rect 2520 7542 2523 7554
rect 2536 7542 2539 7554
rect 2550 7545 2562 7548
rect 2578 7542 2581 7554
rect 2594 7542 2597 7554
rect 2615 7542 2618 7554
rect 2631 7542 2634 7554
rect 2652 7542 2655 7554
rect 2668 7542 2671 7554
rect 2682 7545 2694 7548
rect 2710 7542 2713 7554
rect 2726 7542 2729 7554
rect 2747 7542 2750 7554
rect 3312 7542 3315 7554
rect 3333 7542 3336 7554
rect 3349 7542 3352 7554
rect 3363 7545 3375 7548
rect 3391 7542 3394 7554
rect 3407 7542 3410 7554
rect 3428 7542 3431 7554
rect 3444 7542 3447 7554
rect 3465 7542 3468 7554
rect 3481 7542 3484 7554
rect 3495 7545 3507 7548
rect 3523 7542 3526 7554
rect 3539 7542 3542 7554
rect 3560 7542 3563 7554
rect 3576 7542 3579 7554
rect 3597 7542 3600 7554
rect 3613 7542 3616 7554
rect 3627 7545 3639 7548
rect 3655 7542 3658 7554
rect 3671 7542 3674 7554
rect 3692 7542 3695 7554
rect 2364 7538 2397 7542
rect 2401 7538 2425 7542
rect 2429 7538 2455 7542
rect 2459 7538 2529 7542
rect 2533 7538 2557 7542
rect 2561 7538 2587 7542
rect 2591 7538 2661 7542
rect 2665 7538 2689 7542
rect 2693 7538 2719 7542
rect 2723 7538 2776 7542
rect 3309 7538 3342 7542
rect 3346 7538 3370 7542
rect 3374 7538 3400 7542
rect 3404 7538 3474 7542
rect 3478 7538 3502 7542
rect 3506 7538 3532 7542
rect 3536 7538 3606 7542
rect 3610 7538 3634 7542
rect 3638 7538 3664 7542
rect 3668 7538 3721 7542
rect 2364 7531 2373 7535
rect 2377 7531 2424 7535
rect 2428 7531 2474 7535
rect 2478 7531 2505 7535
rect 2509 7531 2556 7535
rect 2560 7531 2606 7535
rect 2610 7531 2637 7535
rect 2641 7531 2688 7535
rect 2692 7531 2738 7535
rect 2742 7531 2812 7535
rect 3309 7531 3318 7535
rect 3322 7531 3369 7535
rect 3373 7531 3419 7535
rect 3423 7531 3450 7535
rect 3454 7531 3501 7535
rect 3505 7531 3551 7535
rect 3555 7531 3582 7535
rect 3586 7531 3633 7535
rect 3637 7531 3683 7535
rect 3687 7531 3757 7535
rect 2370 7525 2755 7528
rect 3315 7525 3700 7528
rect 2495 7518 2599 7521
rect 3440 7518 3544 7521
rect 4826 7518 4829 7557
rect 5083 7518 5086 7772
rect 4826 7515 5086 7518
rect 2611 7510 2615 7514
rect 2619 7510 2623 7514
rect 3556 7510 3560 7514
rect 3564 7510 3568 7514
rect 86 7502 346 7505
rect 2347 7499 2599 7503
rect 2603 7499 2619 7503
rect 2635 7499 3296 7503
rect 3300 7499 3544 7503
rect 3548 7499 3564 7503
rect 3580 7499 4241 7503
rect 4245 7499 4328 7503
rect 2627 7492 2755 7495
rect 3572 7492 3700 7495
rect 2642 7485 2755 7488
rect 3587 7485 3700 7488
rect 2611 7476 2615 7480
rect 2619 7476 2623 7480
rect 3556 7476 3560 7480
rect 3564 7476 3568 7480
rect 617 7467 618 7471
rect 622 7467 623 7471
rect 627 7467 628 7471
rect 632 7467 633 7471
rect 637 7467 638 7471
rect 642 7467 643 7471
rect 613 7466 647 7467
rect 617 7462 618 7466
rect 622 7462 623 7466
rect 627 7462 628 7466
rect 632 7462 633 7466
rect 637 7462 638 7466
rect 642 7462 643 7466
rect 613 7461 647 7462
rect 617 7457 618 7461
rect 622 7457 623 7461
rect 627 7457 628 7461
rect 632 7457 633 7461
rect 637 7457 638 7461
rect 642 7457 643 7461
rect 613 7456 647 7457
rect 86 7450 346 7453
rect 617 7452 618 7456
rect 622 7452 623 7456
rect 627 7452 628 7456
rect 632 7452 633 7456
rect 637 7452 638 7456
rect 642 7452 643 7456
rect 663 7467 664 7471
rect 668 7467 669 7471
rect 673 7467 674 7471
rect 678 7467 679 7471
rect 683 7467 684 7471
rect 688 7467 689 7471
rect 2495 7469 2599 7472
rect 3440 7469 3544 7472
rect 659 7466 693 7467
rect 663 7462 664 7466
rect 668 7462 669 7466
rect 673 7462 674 7466
rect 678 7462 679 7466
rect 683 7462 684 7466
rect 688 7462 689 7466
rect 2364 7462 2373 7466
rect 2377 7462 2409 7466
rect 2413 7462 2476 7466
rect 2480 7462 2505 7466
rect 2509 7462 2541 7466
rect 2545 7462 2608 7466
rect 2612 7462 2637 7466
rect 2641 7462 2673 7466
rect 2677 7462 2740 7466
rect 2744 7462 2824 7466
rect 3309 7462 3318 7466
rect 3322 7462 3354 7466
rect 3358 7462 3421 7466
rect 3425 7462 3450 7466
rect 3454 7462 3486 7466
rect 3490 7462 3553 7466
rect 3557 7462 3582 7466
rect 3586 7462 3618 7466
rect 3622 7462 3685 7466
rect 3689 7462 3769 7466
rect 4826 7462 5086 7465
rect 659 7461 693 7462
rect 663 7457 664 7461
rect 668 7457 669 7461
rect 673 7457 674 7461
rect 678 7457 679 7461
rect 683 7457 684 7461
rect 688 7457 689 7461
rect 659 7456 693 7457
rect 663 7452 664 7456
rect 668 7452 669 7456
rect 673 7452 674 7456
rect 678 7452 679 7456
rect 683 7452 684 7456
rect 688 7452 689 7456
rect 2364 7455 2397 7459
rect 2401 7455 2425 7459
rect 2429 7455 2455 7459
rect 2459 7455 2492 7459
rect 2496 7455 2529 7459
rect 2533 7455 2557 7459
rect 2561 7455 2587 7459
rect 2591 7455 2624 7459
rect 2628 7455 2661 7459
rect 2665 7455 2689 7459
rect 2693 7455 2719 7459
rect 2723 7455 2756 7459
rect 2760 7455 2764 7459
rect 3309 7455 3342 7459
rect 3346 7455 3370 7459
rect 3374 7455 3400 7459
rect 3404 7455 3437 7459
rect 3441 7455 3474 7459
rect 3478 7455 3502 7459
rect 3506 7455 3532 7459
rect 3536 7455 3569 7459
rect 3573 7455 3606 7459
rect 3610 7455 3634 7459
rect 3638 7455 3664 7459
rect 3668 7455 3701 7459
rect 3705 7455 3709 7459
rect 86 7196 89 7450
rect 343 7411 346 7450
rect 2367 7445 2370 7455
rect 2388 7445 2391 7455
rect 2404 7445 2407 7455
rect 2418 7448 2423 7452
rect 2427 7448 2434 7452
rect 2446 7445 2449 7455
rect 2462 7445 2465 7455
rect 2483 7445 2486 7455
rect 2499 7445 2502 7455
rect 2520 7445 2523 7455
rect 2536 7445 2539 7455
rect 2550 7448 2555 7452
rect 2559 7448 2566 7452
rect 2578 7445 2581 7455
rect 2594 7445 2597 7455
rect 2615 7445 2618 7455
rect 2631 7445 2634 7455
rect 2652 7445 2655 7455
rect 2668 7445 2671 7455
rect 2682 7448 2687 7452
rect 2691 7448 2698 7452
rect 2710 7445 2713 7455
rect 2726 7445 2729 7455
rect 2747 7445 2750 7455
rect 3312 7445 3315 7455
rect 3333 7445 3336 7455
rect 3349 7445 3352 7455
rect 3363 7448 3368 7452
rect 3372 7448 3379 7452
rect 3391 7445 3394 7455
rect 3407 7445 3410 7455
rect 3428 7445 3431 7455
rect 3444 7445 3447 7455
rect 3465 7445 3468 7455
rect 3481 7445 3484 7455
rect 3495 7448 3500 7452
rect 3504 7448 3511 7452
rect 3523 7445 3526 7455
rect 3539 7445 3542 7455
rect 3560 7445 3563 7455
rect 3576 7445 3579 7455
rect 3597 7445 3600 7455
rect 3613 7445 3616 7455
rect 3627 7448 3632 7452
rect 3636 7448 3643 7452
rect 3655 7445 3658 7455
rect 3671 7445 3674 7455
rect 3692 7445 3695 7455
rect 2384 7431 2389 7434
rect 2393 7431 2417 7434
rect 2442 7431 2449 7434
rect 2453 7431 2475 7434
rect 2495 7431 2502 7434
rect 2516 7431 2521 7434
rect 2525 7431 2549 7434
rect 2574 7431 2581 7434
rect 2585 7431 2607 7434
rect 2627 7431 2634 7434
rect 2648 7431 2653 7434
rect 2657 7431 2681 7434
rect 2706 7431 2713 7434
rect 2717 7431 2739 7434
rect 2400 7421 2407 7424
rect 2411 7425 2430 7428
rect 2430 7418 2433 7424
rect 2458 7421 2465 7424
rect 2469 7425 2484 7428
rect 2532 7421 2539 7424
rect 2543 7425 2562 7428
rect 2562 7418 2565 7424
rect 2590 7421 2597 7424
rect 2601 7425 2616 7428
rect 2664 7421 2671 7424
rect 2675 7425 2694 7428
rect 2694 7418 2697 7424
rect 2722 7421 2729 7424
rect 2733 7425 2750 7428
rect 3329 7431 3334 7434
rect 3338 7431 3362 7434
rect 3387 7431 3394 7434
rect 3398 7431 3420 7434
rect 3440 7431 3447 7434
rect 3461 7431 3466 7434
rect 3470 7431 3494 7434
rect 3519 7431 3526 7434
rect 3530 7431 3552 7434
rect 3572 7431 3579 7434
rect 3593 7431 3598 7434
rect 3602 7431 3626 7434
rect 3651 7431 3658 7434
rect 3662 7431 3684 7434
rect 3345 7421 3352 7424
rect 3356 7425 3375 7428
rect 3375 7418 3378 7424
rect 3403 7421 3410 7424
rect 3414 7425 3429 7428
rect 3477 7421 3484 7424
rect 3488 7425 3507 7428
rect 3507 7418 3510 7424
rect 3535 7421 3542 7424
rect 3546 7425 3561 7428
rect 3609 7421 3616 7424
rect 3620 7425 3639 7428
rect 3639 7418 3642 7424
rect 3667 7421 3674 7424
rect 3678 7425 3695 7428
rect 4826 7423 4829 7462
rect 343 7401 356 7411
rect 2367 7402 2370 7414
rect 2388 7402 2391 7414
rect 2404 7402 2407 7414
rect 2418 7405 2430 7408
rect 2446 7402 2449 7414
rect 2462 7402 2465 7414
rect 2483 7402 2486 7414
rect 2499 7402 2502 7414
rect 2520 7402 2523 7414
rect 2536 7402 2539 7414
rect 2550 7405 2562 7408
rect 2578 7402 2581 7414
rect 2594 7402 2597 7414
rect 2615 7402 2618 7414
rect 2631 7402 2634 7414
rect 2652 7402 2655 7414
rect 2668 7402 2671 7414
rect 2682 7405 2694 7408
rect 2710 7402 2713 7414
rect 2726 7402 2729 7414
rect 2747 7402 2750 7414
rect 3312 7402 3315 7414
rect 3333 7402 3336 7414
rect 3349 7402 3352 7414
rect 3363 7405 3375 7408
rect 3391 7402 3394 7414
rect 3407 7402 3410 7414
rect 3428 7402 3431 7414
rect 3444 7402 3447 7414
rect 3465 7402 3468 7414
rect 3481 7402 3484 7414
rect 3495 7405 3507 7408
rect 3523 7402 3526 7414
rect 3539 7402 3542 7414
rect 3560 7402 3563 7414
rect 3576 7402 3579 7414
rect 3597 7402 3600 7414
rect 3613 7402 3616 7414
rect 3627 7405 3639 7408
rect 3655 7402 3658 7414
rect 3671 7402 3674 7414
rect 3692 7402 3695 7414
rect 4816 7413 4829 7423
rect 4806 7403 4829 7413
rect 343 7391 366 7401
rect 2364 7398 2397 7402
rect 2401 7398 2425 7402
rect 2429 7398 2455 7402
rect 2459 7398 2529 7402
rect 2533 7398 2557 7402
rect 2561 7398 2587 7402
rect 2591 7398 2661 7402
rect 2665 7398 2689 7402
rect 2693 7398 2719 7402
rect 2723 7398 2776 7402
rect 3309 7398 3342 7402
rect 3346 7398 3370 7402
rect 3374 7398 3400 7402
rect 3404 7398 3474 7402
rect 3478 7398 3502 7402
rect 3506 7398 3532 7402
rect 3536 7398 3606 7402
rect 3610 7398 3634 7402
rect 3638 7398 3664 7402
rect 3668 7398 3721 7402
rect 2364 7391 2373 7395
rect 2377 7391 2424 7395
rect 2428 7391 2474 7395
rect 2478 7391 2505 7395
rect 2509 7391 2556 7395
rect 2560 7391 2606 7395
rect 2610 7391 2637 7395
rect 2641 7391 2688 7395
rect 2692 7391 2738 7395
rect 2742 7391 2812 7395
rect 3309 7391 3318 7395
rect 3322 7391 3369 7395
rect 3373 7391 3419 7395
rect 3423 7391 3450 7395
rect 3454 7391 3501 7395
rect 3505 7391 3551 7395
rect 3555 7391 3582 7395
rect 3586 7391 3633 7395
rect 3637 7391 3683 7395
rect 3687 7391 3757 7395
rect 4796 7393 4829 7403
rect 343 7381 376 7391
rect 4786 7383 4829 7393
rect 343 7371 386 7381
rect 343 7275 769 7371
rect 4403 7287 4829 7383
rect 4786 7277 4829 7287
rect 343 7265 386 7275
rect 4796 7267 4829 7277
rect 343 7255 376 7265
rect 4806 7257 4829 7267
rect 343 7245 366 7255
rect 4816 7247 4829 7257
rect 343 7235 356 7245
rect 343 7196 346 7235
rect 4826 7208 4829 7247
rect 5083 7208 5086 7462
rect 86 7193 346 7196
rect 4483 7202 4484 7206
rect 4488 7202 4489 7206
rect 4493 7202 4494 7206
rect 4498 7202 4499 7206
rect 4503 7202 4504 7206
rect 4508 7202 4509 7206
rect 4479 7201 4513 7202
rect 4483 7197 4484 7201
rect 4488 7197 4489 7201
rect 4493 7197 4494 7201
rect 4498 7197 4499 7201
rect 4503 7197 4504 7201
rect 4508 7197 4509 7201
rect 4479 7196 4513 7197
rect 4483 7192 4484 7196
rect 4488 7192 4489 7196
rect 4493 7192 4494 7196
rect 4498 7192 4499 7196
rect 4503 7192 4504 7196
rect 4508 7192 4509 7196
rect 4479 7191 4513 7192
rect 4483 7187 4484 7191
rect 4488 7187 4489 7191
rect 4493 7187 4494 7191
rect 4498 7187 4499 7191
rect 4503 7187 4504 7191
rect 4508 7187 4509 7191
rect 4529 7202 4530 7206
rect 4534 7202 4535 7206
rect 4539 7202 4540 7206
rect 4544 7202 4545 7206
rect 4549 7202 4550 7206
rect 4554 7202 4555 7206
rect 4826 7205 5086 7208
rect 4525 7201 4559 7202
rect 4529 7197 4530 7201
rect 4534 7197 4535 7201
rect 4539 7197 4540 7201
rect 4544 7197 4545 7201
rect 4549 7197 4550 7201
rect 4554 7197 4555 7201
rect 4525 7196 4559 7197
rect 4529 7192 4530 7196
rect 4534 7192 4535 7196
rect 4539 7192 4540 7196
rect 4544 7192 4545 7196
rect 4549 7192 4550 7196
rect 4554 7192 4555 7196
rect 4525 7191 4559 7192
rect 4529 7187 4530 7191
rect 4534 7187 4535 7191
rect 4539 7187 4540 7191
rect 4544 7187 4545 7191
rect 4549 7187 4550 7191
rect 4554 7187 4555 7191
rect 617 7158 618 7162
rect 622 7158 623 7162
rect 627 7158 628 7162
rect 632 7158 633 7162
rect 637 7158 638 7162
rect 642 7158 643 7162
rect 613 7157 647 7158
rect 617 7153 618 7157
rect 622 7153 623 7157
rect 627 7153 628 7157
rect 632 7153 633 7157
rect 637 7153 638 7157
rect 642 7153 643 7157
rect 613 7152 647 7153
rect 617 7148 618 7152
rect 622 7148 623 7152
rect 627 7148 628 7152
rect 632 7148 633 7152
rect 637 7148 638 7152
rect 642 7148 643 7152
rect 613 7147 647 7148
rect 86 7141 346 7144
rect 617 7143 618 7147
rect 622 7143 623 7147
rect 627 7143 628 7147
rect 632 7143 633 7147
rect 637 7143 638 7147
rect 642 7143 643 7147
rect 663 7158 664 7162
rect 668 7158 669 7162
rect 673 7158 674 7162
rect 678 7158 679 7162
rect 683 7158 684 7162
rect 688 7158 689 7162
rect 659 7157 693 7158
rect 663 7153 664 7157
rect 668 7153 669 7157
rect 673 7153 674 7157
rect 678 7153 679 7157
rect 683 7153 684 7157
rect 688 7153 689 7157
rect 659 7152 693 7153
rect 663 7148 664 7152
rect 668 7148 669 7152
rect 673 7148 674 7152
rect 678 7148 679 7152
rect 683 7148 684 7152
rect 688 7148 689 7152
rect 659 7147 693 7148
rect 663 7143 664 7147
rect 668 7143 669 7147
rect 673 7143 674 7147
rect 678 7143 679 7147
rect 683 7143 684 7147
rect 688 7143 689 7147
rect 4826 7153 5086 7156
rect 86 6887 89 7141
rect 343 7102 346 7141
rect 4826 7114 4829 7153
rect 4816 7104 4829 7114
rect 343 7092 356 7102
rect 4806 7094 4829 7104
rect 343 7082 366 7092
rect 4796 7084 4829 7094
rect 343 7072 376 7082
rect 4786 7074 4829 7084
rect 343 7062 386 7072
rect 343 6966 769 7062
rect 4403 6978 4829 7074
rect 4786 6968 4829 6978
rect 343 6956 386 6966
rect 4796 6958 4829 6968
rect 343 6946 376 6956
rect 4806 6948 4829 6958
rect 343 6936 366 6946
rect 4816 6938 4829 6948
rect 343 6926 356 6936
rect 343 6887 346 6926
rect 4826 6899 4829 6938
rect 5083 6899 5086 7153
rect 86 6884 346 6887
rect 4483 6893 4484 6897
rect 4488 6893 4489 6897
rect 4493 6893 4494 6897
rect 4498 6893 4499 6897
rect 4503 6893 4504 6897
rect 4508 6893 4509 6897
rect 4479 6892 4513 6893
rect 4483 6888 4484 6892
rect 4488 6888 4489 6892
rect 4493 6888 4494 6892
rect 4498 6888 4499 6892
rect 4503 6888 4504 6892
rect 4508 6888 4509 6892
rect 4479 6887 4513 6888
rect 4483 6883 4484 6887
rect 4488 6883 4489 6887
rect 4493 6883 4494 6887
rect 4498 6883 4499 6887
rect 4503 6883 4504 6887
rect 4508 6883 4509 6887
rect 4479 6882 4513 6883
rect 4483 6878 4484 6882
rect 4488 6878 4489 6882
rect 4493 6878 4494 6882
rect 4498 6878 4499 6882
rect 4503 6878 4504 6882
rect 4508 6878 4509 6882
rect 4529 6893 4530 6897
rect 4534 6893 4535 6897
rect 4539 6893 4540 6897
rect 4544 6893 4545 6897
rect 4549 6893 4550 6897
rect 4554 6893 4555 6897
rect 4826 6896 5086 6899
rect 4525 6892 4559 6893
rect 4529 6888 4530 6892
rect 4534 6888 4535 6892
rect 4539 6888 4540 6892
rect 4544 6888 4545 6892
rect 4549 6888 4550 6892
rect 4554 6888 4555 6892
rect 4525 6887 4559 6888
rect 4529 6883 4530 6887
rect 4534 6883 4535 6887
rect 4539 6883 4540 6887
rect 4544 6883 4545 6887
rect 4549 6883 4550 6887
rect 4554 6883 4555 6887
rect 4525 6882 4559 6883
rect 4529 6878 4530 6882
rect 4534 6878 4535 6882
rect 4539 6878 4540 6882
rect 4544 6878 4545 6882
rect 4549 6878 4550 6882
rect 4554 6878 4555 6882
rect 617 6849 618 6853
rect 622 6849 623 6853
rect 627 6849 628 6853
rect 632 6849 633 6853
rect 637 6849 638 6853
rect 642 6849 643 6853
rect 613 6848 647 6849
rect 617 6844 618 6848
rect 622 6844 623 6848
rect 627 6844 628 6848
rect 632 6844 633 6848
rect 637 6844 638 6848
rect 642 6844 643 6848
rect 613 6843 647 6844
rect 617 6839 618 6843
rect 622 6839 623 6843
rect 627 6839 628 6843
rect 632 6839 633 6843
rect 637 6839 638 6843
rect 642 6839 643 6843
rect 613 6838 647 6839
rect 86 6832 346 6835
rect 617 6834 618 6838
rect 622 6834 623 6838
rect 627 6834 628 6838
rect 632 6834 633 6838
rect 637 6834 638 6838
rect 642 6834 643 6838
rect 663 6849 664 6853
rect 668 6849 669 6853
rect 673 6849 674 6853
rect 678 6849 679 6853
rect 683 6849 684 6853
rect 688 6849 689 6853
rect 659 6848 693 6849
rect 663 6844 664 6848
rect 668 6844 669 6848
rect 673 6844 674 6848
rect 678 6844 679 6848
rect 683 6844 684 6848
rect 688 6844 689 6848
rect 659 6843 693 6844
rect 663 6839 664 6843
rect 668 6839 669 6843
rect 673 6839 674 6843
rect 678 6839 679 6843
rect 683 6839 684 6843
rect 688 6839 689 6843
rect 659 6838 693 6839
rect 663 6834 664 6838
rect 668 6834 669 6838
rect 673 6834 674 6838
rect 678 6834 679 6838
rect 683 6834 684 6838
rect 688 6834 689 6838
rect 4826 6844 5086 6847
rect 86 6578 89 6832
rect 343 6793 346 6832
rect 4826 6805 4829 6844
rect 4816 6795 4829 6805
rect 343 6783 356 6793
rect 4806 6785 4829 6795
rect 343 6773 366 6783
rect 4796 6775 4829 6785
rect 343 6763 376 6773
rect 4786 6765 4829 6775
rect 343 6753 386 6763
rect 343 6657 769 6753
rect 4403 6669 4829 6765
rect 4786 6659 4829 6669
rect 343 6647 386 6657
rect 4796 6649 4829 6659
rect 343 6637 376 6647
rect 4806 6639 4829 6649
rect 343 6627 366 6637
rect 4816 6629 4829 6639
rect 343 6617 356 6627
rect 343 6578 346 6617
rect 4826 6590 4829 6629
rect 5083 6590 5086 6844
rect 86 6575 346 6578
rect 4483 6584 4484 6588
rect 4488 6584 4489 6588
rect 4493 6584 4494 6588
rect 4498 6584 4499 6588
rect 4503 6584 4504 6588
rect 4508 6584 4509 6588
rect 4479 6583 4513 6584
rect 4483 6579 4484 6583
rect 4488 6579 4489 6583
rect 4493 6579 4494 6583
rect 4498 6579 4499 6583
rect 4503 6579 4504 6583
rect 4508 6579 4509 6583
rect 4479 6578 4513 6579
rect 4483 6574 4484 6578
rect 4488 6574 4489 6578
rect 4493 6574 4494 6578
rect 4498 6574 4499 6578
rect 4503 6574 4504 6578
rect 4508 6574 4509 6578
rect 4479 6573 4513 6574
rect 4483 6569 4484 6573
rect 4488 6569 4489 6573
rect 4493 6569 4494 6573
rect 4498 6569 4499 6573
rect 4503 6569 4504 6573
rect 4508 6569 4509 6573
rect 4529 6584 4530 6588
rect 4534 6584 4535 6588
rect 4539 6584 4540 6588
rect 4544 6584 4545 6588
rect 4549 6584 4550 6588
rect 4554 6584 4555 6588
rect 4826 6587 5086 6590
rect 4525 6583 4559 6584
rect 4529 6579 4530 6583
rect 4534 6579 4535 6583
rect 4539 6579 4540 6583
rect 4544 6579 4545 6583
rect 4549 6579 4550 6583
rect 4554 6579 4555 6583
rect 4525 6578 4559 6579
rect 4529 6574 4530 6578
rect 4534 6574 4535 6578
rect 4539 6574 4540 6578
rect 4544 6574 4545 6578
rect 4549 6574 4550 6578
rect 4554 6574 4555 6578
rect 4525 6573 4559 6574
rect 4529 6569 4530 6573
rect 4534 6569 4535 6573
rect 4539 6569 4540 6573
rect 4544 6569 4545 6573
rect 4549 6569 4550 6573
rect 4554 6569 4555 6573
rect 617 6540 618 6544
rect 622 6540 623 6544
rect 627 6540 628 6544
rect 632 6540 633 6544
rect 637 6540 638 6544
rect 642 6540 643 6544
rect 613 6539 647 6540
rect 617 6535 618 6539
rect 622 6535 623 6539
rect 627 6535 628 6539
rect 632 6535 633 6539
rect 637 6535 638 6539
rect 642 6535 643 6539
rect 613 6534 647 6535
rect 617 6530 618 6534
rect 622 6530 623 6534
rect 627 6530 628 6534
rect 632 6530 633 6534
rect 637 6530 638 6534
rect 642 6530 643 6534
rect 613 6529 647 6530
rect 86 6523 346 6526
rect 617 6525 618 6529
rect 622 6525 623 6529
rect 627 6525 628 6529
rect 632 6525 633 6529
rect 637 6525 638 6529
rect 642 6525 643 6529
rect 663 6540 664 6544
rect 668 6540 669 6544
rect 673 6540 674 6544
rect 678 6540 679 6544
rect 683 6540 684 6544
rect 688 6540 689 6544
rect 659 6539 693 6540
rect 663 6535 664 6539
rect 668 6535 669 6539
rect 673 6535 674 6539
rect 678 6535 679 6539
rect 683 6535 684 6539
rect 688 6535 689 6539
rect 659 6534 693 6535
rect 663 6530 664 6534
rect 668 6530 669 6534
rect 673 6530 674 6534
rect 678 6530 679 6534
rect 683 6530 684 6534
rect 688 6530 689 6534
rect 659 6529 693 6530
rect 663 6525 664 6529
rect 668 6525 669 6529
rect 673 6525 674 6529
rect 678 6525 679 6529
rect 683 6525 684 6529
rect 688 6525 689 6529
rect 4826 6535 5086 6538
rect 86 6269 89 6523
rect 343 6484 346 6523
rect 4826 6496 4829 6535
rect 4816 6486 4829 6496
rect 343 6474 356 6484
rect 4806 6476 4829 6486
rect 343 6464 366 6474
rect 4796 6466 4829 6476
rect 343 6454 376 6464
rect 4786 6456 4829 6466
rect 343 6444 386 6454
rect 343 6348 769 6444
rect 4403 6360 4829 6456
rect 4786 6350 4829 6360
rect 343 6338 386 6348
rect 4796 6340 4829 6350
rect 343 6328 376 6338
rect 4806 6330 4829 6340
rect 343 6318 366 6328
rect 4816 6320 4829 6330
rect 343 6308 356 6318
rect 343 6269 346 6308
rect 4826 6281 4829 6320
rect 5083 6281 5086 6535
rect 86 6266 346 6269
rect 4483 6275 4484 6279
rect 4488 6275 4489 6279
rect 4493 6275 4494 6279
rect 4498 6275 4499 6279
rect 4503 6275 4504 6279
rect 4508 6275 4509 6279
rect 4479 6274 4513 6275
rect 4483 6270 4484 6274
rect 4488 6270 4489 6274
rect 4493 6270 4494 6274
rect 4498 6270 4499 6274
rect 4503 6270 4504 6274
rect 4508 6270 4509 6274
rect 4479 6269 4513 6270
rect 4483 6265 4484 6269
rect 4488 6265 4489 6269
rect 4493 6265 4494 6269
rect 4498 6265 4499 6269
rect 4503 6265 4504 6269
rect 4508 6265 4509 6269
rect 4479 6264 4513 6265
rect 4483 6260 4484 6264
rect 4488 6260 4489 6264
rect 4493 6260 4494 6264
rect 4498 6260 4499 6264
rect 4503 6260 4504 6264
rect 4508 6260 4509 6264
rect 4529 6275 4530 6279
rect 4534 6275 4535 6279
rect 4539 6275 4540 6279
rect 4544 6275 4545 6279
rect 4549 6275 4550 6279
rect 4554 6275 4555 6279
rect 4826 6278 5086 6281
rect 4525 6274 4559 6275
rect 4529 6270 4530 6274
rect 4534 6270 4535 6274
rect 4539 6270 4540 6274
rect 4544 6270 4545 6274
rect 4549 6270 4550 6274
rect 4554 6270 4555 6274
rect 4525 6269 4559 6270
rect 4529 6265 4530 6269
rect 4534 6265 4535 6269
rect 4539 6265 4540 6269
rect 4544 6265 4545 6269
rect 4549 6265 4550 6269
rect 4554 6265 4555 6269
rect 4525 6264 4559 6265
rect 4529 6260 4530 6264
rect 4534 6260 4535 6264
rect 4539 6260 4540 6264
rect 4544 6260 4545 6264
rect 4549 6260 4550 6264
rect 4554 6260 4555 6264
rect 99 5800 593 6231
rect 617 6140 618 6144
rect 622 6140 623 6144
rect 627 6140 628 6144
rect 632 6140 633 6144
rect 637 6140 638 6144
rect 642 6140 643 6144
rect 613 6139 647 6140
rect 617 6135 618 6139
rect 622 6135 623 6139
rect 627 6135 628 6139
rect 632 6135 633 6139
rect 637 6135 638 6139
rect 642 6135 643 6139
rect 613 6134 647 6135
rect 617 6130 618 6134
rect 622 6130 623 6134
rect 627 6130 628 6134
rect 632 6130 633 6134
rect 637 6130 638 6134
rect 642 6130 643 6134
rect 613 6129 647 6130
rect 617 6125 618 6129
rect 622 6125 623 6129
rect 627 6125 628 6129
rect 632 6125 633 6129
rect 637 6125 638 6129
rect 642 6125 643 6129
rect 663 6140 664 6144
rect 668 6140 669 6144
rect 673 6140 674 6144
rect 678 6140 679 6144
rect 683 6140 684 6144
rect 688 6140 689 6144
rect 659 6139 693 6140
rect 663 6135 664 6139
rect 668 6135 669 6139
rect 673 6135 674 6139
rect 678 6135 679 6139
rect 683 6135 684 6139
rect 688 6135 689 6139
rect 659 6134 693 6135
rect 663 6130 664 6134
rect 668 6130 669 6134
rect 673 6130 674 6134
rect 678 6130 679 6134
rect 683 6130 684 6134
rect 688 6130 689 6134
rect 659 6129 693 6130
rect 663 6125 664 6129
rect 668 6125 669 6129
rect 673 6125 674 6129
rect 678 6125 679 6129
rect 683 6125 684 6129
rect 688 6125 689 6129
rect 617 6111 618 6115
rect 622 6111 623 6115
rect 627 6111 628 6115
rect 632 6111 633 6115
rect 637 6111 638 6115
rect 642 6111 643 6115
rect 613 6110 647 6111
rect 617 6106 618 6110
rect 622 6106 623 6110
rect 627 6106 628 6110
rect 632 6106 633 6110
rect 637 6106 638 6110
rect 642 6106 643 6110
rect 613 6105 647 6106
rect 617 6101 618 6105
rect 622 6101 623 6105
rect 627 6101 628 6105
rect 632 6101 633 6105
rect 637 6101 638 6105
rect 642 6101 643 6105
rect 613 6100 647 6101
rect 617 6096 618 6100
rect 622 6096 623 6100
rect 627 6096 628 6100
rect 632 6096 633 6100
rect 637 6096 638 6100
rect 642 6096 643 6100
rect 663 6111 664 6115
rect 668 6111 669 6115
rect 673 6111 674 6115
rect 678 6111 679 6115
rect 683 6111 684 6115
rect 688 6111 689 6115
rect 659 6110 693 6111
rect 663 6106 664 6110
rect 668 6106 669 6110
rect 673 6106 674 6110
rect 678 6106 679 6110
rect 683 6106 684 6110
rect 688 6106 689 6110
rect 659 6105 693 6106
rect 663 6101 664 6105
rect 668 6101 669 6105
rect 673 6101 674 6105
rect 678 6101 679 6105
rect 683 6101 684 6105
rect 688 6101 689 6105
rect 659 6100 693 6101
rect 663 6096 664 6100
rect 668 6096 669 6100
rect 673 6096 674 6100
rect 678 6096 679 6100
rect 683 6096 684 6100
rect 688 6096 689 6100
rect 617 6082 618 6086
rect 622 6082 623 6086
rect 627 6082 628 6086
rect 632 6082 633 6086
rect 637 6082 638 6086
rect 642 6082 643 6086
rect 613 6081 647 6082
rect 617 6077 618 6081
rect 622 6077 623 6081
rect 627 6077 628 6081
rect 632 6077 633 6081
rect 637 6077 638 6081
rect 642 6077 643 6081
rect 613 6076 647 6077
rect 617 6072 618 6076
rect 622 6072 623 6076
rect 627 6072 628 6076
rect 632 6072 633 6076
rect 637 6072 638 6076
rect 642 6072 643 6076
rect 613 6071 647 6072
rect 617 6067 618 6071
rect 622 6067 623 6071
rect 627 6067 628 6071
rect 632 6067 633 6071
rect 637 6067 638 6071
rect 642 6067 643 6071
rect 663 6082 664 6086
rect 668 6082 669 6086
rect 673 6082 674 6086
rect 678 6082 679 6086
rect 683 6082 684 6086
rect 688 6082 689 6086
rect 659 6081 693 6082
rect 663 6077 664 6081
rect 668 6077 669 6081
rect 673 6077 674 6081
rect 678 6077 679 6081
rect 683 6077 684 6081
rect 688 6077 689 6081
rect 659 6076 693 6077
rect 663 6072 664 6076
rect 668 6072 669 6076
rect 673 6072 674 6076
rect 678 6072 679 6076
rect 683 6072 684 6076
rect 688 6072 689 6076
rect 659 6071 693 6072
rect 663 6067 664 6071
rect 668 6067 669 6071
rect 673 6067 674 6071
rect 678 6067 679 6071
rect 683 6067 684 6071
rect 688 6067 689 6071
rect 4483 6083 4484 6087
rect 4488 6083 4489 6087
rect 4493 6083 4494 6087
rect 4498 6083 4499 6087
rect 4503 6083 4504 6087
rect 4508 6083 4509 6087
rect 4479 6082 4513 6083
rect 4483 6078 4484 6082
rect 4488 6078 4489 6082
rect 4493 6078 4494 6082
rect 4498 6078 4499 6082
rect 4503 6078 4504 6082
rect 4508 6078 4509 6082
rect 4479 6077 4513 6078
rect 4483 6073 4484 6077
rect 4488 6073 4489 6077
rect 4493 6073 4494 6077
rect 4498 6073 4499 6077
rect 4503 6073 4504 6077
rect 4508 6073 4509 6077
rect 4479 6072 4513 6073
rect 4483 6068 4484 6072
rect 4488 6068 4489 6072
rect 4493 6068 4494 6072
rect 4498 6068 4499 6072
rect 4503 6068 4504 6072
rect 4508 6068 4509 6072
rect 4529 6083 4530 6087
rect 4534 6083 4535 6087
rect 4539 6083 4540 6087
rect 4544 6083 4545 6087
rect 4549 6083 4550 6087
rect 4554 6083 4555 6087
rect 4525 6082 4559 6083
rect 4529 6078 4530 6082
rect 4534 6078 4535 6082
rect 4539 6078 4540 6082
rect 4544 6078 4545 6082
rect 4549 6078 4550 6082
rect 4554 6078 4555 6082
rect 4525 6077 4559 6078
rect 4529 6073 4530 6077
rect 4534 6073 4535 6077
rect 4539 6073 4540 6077
rect 4544 6073 4545 6077
rect 4549 6073 4550 6077
rect 4554 6073 4555 6077
rect 4525 6072 4559 6073
rect 4529 6068 4530 6072
rect 4534 6068 4535 6072
rect 4539 6068 4540 6072
rect 4544 6068 4545 6072
rect 4549 6068 4550 6072
rect 4554 6068 4555 6072
rect 4483 6057 4484 6061
rect 4488 6057 4489 6061
rect 4493 6057 4494 6061
rect 4498 6057 4499 6061
rect 4503 6057 4504 6061
rect 4508 6057 4509 6061
rect 617 6053 618 6057
rect 622 6053 623 6057
rect 627 6053 628 6057
rect 632 6053 633 6057
rect 637 6053 638 6057
rect 642 6053 643 6057
rect 613 6052 647 6053
rect 617 6048 618 6052
rect 622 6048 623 6052
rect 627 6048 628 6052
rect 632 6048 633 6052
rect 637 6048 638 6052
rect 642 6048 643 6052
rect 613 6047 647 6048
rect 617 6043 618 6047
rect 622 6043 623 6047
rect 627 6043 628 6047
rect 632 6043 633 6047
rect 637 6043 638 6047
rect 642 6043 643 6047
rect 613 6042 647 6043
rect 617 6038 618 6042
rect 622 6038 623 6042
rect 627 6038 628 6042
rect 632 6038 633 6042
rect 637 6038 638 6042
rect 642 6038 643 6042
rect 663 6053 664 6057
rect 668 6053 669 6057
rect 673 6053 674 6057
rect 678 6053 679 6057
rect 683 6053 684 6057
rect 688 6053 689 6057
rect 659 6052 693 6053
rect 663 6048 664 6052
rect 668 6048 669 6052
rect 673 6048 674 6052
rect 678 6048 679 6052
rect 683 6048 684 6052
rect 688 6048 689 6052
rect 659 6047 693 6048
rect 663 6043 664 6047
rect 668 6043 669 6047
rect 673 6043 674 6047
rect 678 6043 679 6047
rect 683 6043 684 6047
rect 688 6043 689 6047
rect 659 6042 693 6043
rect 4479 6056 4513 6057
rect 4483 6052 4484 6056
rect 4488 6052 4489 6056
rect 4493 6052 4494 6056
rect 4498 6052 4499 6056
rect 4503 6052 4504 6056
rect 4508 6052 4509 6056
rect 4479 6051 4513 6052
rect 4483 6047 4484 6051
rect 4488 6047 4489 6051
rect 4493 6047 4494 6051
rect 4498 6047 4499 6051
rect 4503 6047 4504 6051
rect 4508 6047 4509 6051
rect 4479 6046 4513 6047
rect 4483 6042 4484 6046
rect 4488 6042 4489 6046
rect 4493 6042 4494 6046
rect 4498 6042 4499 6046
rect 4503 6042 4504 6046
rect 4508 6042 4509 6046
rect 4529 6057 4530 6061
rect 4534 6057 4535 6061
rect 4539 6057 4540 6061
rect 4544 6057 4545 6061
rect 4549 6057 4550 6061
rect 4554 6057 4555 6061
rect 4525 6056 4559 6057
rect 4529 6052 4530 6056
rect 4534 6052 4535 6056
rect 4539 6052 4540 6056
rect 4544 6052 4545 6056
rect 4549 6052 4550 6056
rect 4554 6052 4555 6056
rect 4525 6051 4559 6052
rect 4529 6047 4530 6051
rect 4534 6047 4535 6051
rect 4539 6047 4540 6051
rect 4544 6047 4545 6051
rect 4549 6047 4550 6051
rect 4554 6047 4555 6051
rect 4525 6046 4559 6047
rect 4529 6042 4530 6046
rect 4534 6042 4535 6046
rect 4539 6042 4540 6046
rect 4544 6042 4545 6046
rect 4549 6042 4550 6046
rect 4554 6042 4555 6046
rect 663 6038 664 6042
rect 668 6038 669 6042
rect 673 6038 674 6042
rect 678 6038 679 6042
rect 683 6038 684 6042
rect 688 6038 689 6042
rect 4483 6031 4484 6035
rect 4488 6031 4489 6035
rect 4493 6031 4494 6035
rect 4498 6031 4499 6035
rect 4503 6031 4504 6035
rect 4508 6031 4509 6035
rect 4479 6030 4513 6031
rect 617 6024 618 6028
rect 622 6024 623 6028
rect 627 6024 628 6028
rect 632 6024 633 6028
rect 637 6024 638 6028
rect 642 6024 643 6028
rect 613 6023 647 6024
rect 617 6019 618 6023
rect 622 6019 623 6023
rect 627 6019 628 6023
rect 632 6019 633 6023
rect 637 6019 638 6023
rect 642 6019 643 6023
rect 613 6018 647 6019
rect 617 6014 618 6018
rect 622 6014 623 6018
rect 627 6014 628 6018
rect 632 6014 633 6018
rect 637 6014 638 6018
rect 642 6014 643 6018
rect 613 6013 647 6014
rect 617 6009 618 6013
rect 622 6009 623 6013
rect 627 6009 628 6013
rect 632 6009 633 6013
rect 637 6009 638 6013
rect 642 6009 643 6013
rect 663 6024 664 6028
rect 668 6024 669 6028
rect 673 6024 674 6028
rect 678 6024 679 6028
rect 683 6024 684 6028
rect 688 6024 689 6028
rect 659 6023 693 6024
rect 663 6019 664 6023
rect 668 6019 669 6023
rect 673 6019 674 6023
rect 678 6019 679 6023
rect 683 6019 684 6023
rect 688 6019 689 6023
rect 659 6018 693 6019
rect 663 6014 664 6018
rect 668 6014 669 6018
rect 673 6014 674 6018
rect 678 6014 679 6018
rect 683 6014 684 6018
rect 688 6014 689 6018
rect 4483 6026 4484 6030
rect 4488 6026 4489 6030
rect 4493 6026 4494 6030
rect 4498 6026 4499 6030
rect 4503 6026 4504 6030
rect 4508 6026 4509 6030
rect 4479 6025 4513 6026
rect 4483 6021 4484 6025
rect 4488 6021 4489 6025
rect 4493 6021 4494 6025
rect 4498 6021 4499 6025
rect 4503 6021 4504 6025
rect 4508 6021 4509 6025
rect 4479 6020 4513 6021
rect 4483 6016 4484 6020
rect 4488 6016 4489 6020
rect 4493 6016 4494 6020
rect 4498 6016 4499 6020
rect 4503 6016 4504 6020
rect 4508 6016 4509 6020
rect 4529 6031 4530 6035
rect 4534 6031 4535 6035
rect 4539 6031 4540 6035
rect 4544 6031 4545 6035
rect 4549 6031 4550 6035
rect 4554 6031 4555 6035
rect 4525 6030 4559 6031
rect 4529 6026 4530 6030
rect 4534 6026 4535 6030
rect 4539 6026 4540 6030
rect 4544 6026 4545 6030
rect 4549 6026 4550 6030
rect 4554 6026 4555 6030
rect 4525 6025 4559 6026
rect 4529 6021 4530 6025
rect 4534 6021 4535 6025
rect 4539 6021 4540 6025
rect 4544 6021 4545 6025
rect 4549 6021 4550 6025
rect 4554 6021 4555 6025
rect 4525 6020 4559 6021
rect 4529 6016 4530 6020
rect 4534 6016 4535 6020
rect 4539 6016 4540 6020
rect 4544 6016 4545 6020
rect 4549 6016 4550 6020
rect 4554 6016 4555 6020
rect 659 6013 693 6014
rect 663 6009 664 6013
rect 668 6009 669 6013
rect 673 6009 674 6013
rect 678 6009 679 6013
rect 683 6009 684 6013
rect 688 6009 689 6013
rect 4483 6005 4484 6009
rect 4488 6005 4489 6009
rect 4493 6005 4494 6009
rect 4498 6005 4499 6009
rect 4503 6005 4504 6009
rect 4508 6005 4509 6009
rect 4479 6004 4513 6005
rect 4483 6000 4484 6004
rect 4488 6000 4489 6004
rect 4493 6000 4494 6004
rect 4498 6000 4499 6004
rect 4503 6000 4504 6004
rect 4508 6000 4509 6004
rect 4479 5999 4513 6000
rect 4483 5995 4484 5999
rect 4488 5995 4489 5999
rect 4493 5995 4494 5999
rect 4498 5995 4499 5999
rect 4503 5995 4504 5999
rect 4508 5995 4509 5999
rect 4479 5994 4513 5995
rect 4483 5990 4484 5994
rect 4488 5990 4489 5994
rect 4493 5990 4494 5994
rect 4498 5990 4499 5994
rect 4503 5990 4504 5994
rect 4508 5990 4509 5994
rect 4529 6005 4530 6009
rect 4534 6005 4535 6009
rect 4539 6005 4540 6009
rect 4544 6005 4545 6009
rect 4549 6005 4550 6009
rect 4554 6005 4555 6009
rect 4525 6004 4559 6005
rect 4529 6000 4530 6004
rect 4534 6000 4535 6004
rect 4539 6000 4540 6004
rect 4544 6000 4545 6004
rect 4549 6000 4550 6004
rect 4554 6000 4555 6004
rect 4525 5999 4559 6000
rect 4529 5995 4530 5999
rect 4534 5995 4535 5999
rect 4539 5995 4540 5999
rect 4544 5995 4545 5999
rect 4549 5995 4550 5999
rect 4554 5995 4555 5999
rect 4525 5994 4559 5995
rect 4529 5990 4530 5994
rect 4534 5990 4535 5994
rect 4539 5990 4540 5994
rect 4544 5990 4545 5994
rect 4549 5990 4550 5994
rect 4554 5990 4555 5994
rect 4483 5979 4484 5983
rect 4488 5979 4489 5983
rect 4493 5979 4494 5983
rect 4498 5979 4499 5983
rect 4503 5979 4504 5983
rect 4508 5979 4509 5983
rect 4479 5978 4513 5979
rect 761 5896 762 5900
rect 766 5896 767 5900
rect 771 5896 772 5900
rect 757 5895 776 5896
rect 761 5891 762 5895
rect 766 5891 767 5895
rect 771 5891 772 5895
rect 757 5890 776 5891
rect 761 5886 762 5890
rect 766 5886 767 5890
rect 771 5886 772 5890
rect 757 5885 776 5886
rect 761 5881 762 5885
rect 766 5881 767 5885
rect 771 5881 772 5885
rect 757 5880 776 5881
rect 761 5876 762 5880
rect 766 5876 767 5880
rect 771 5876 772 5880
rect 757 5875 776 5876
rect 761 5871 762 5875
rect 766 5871 767 5875
rect 771 5871 772 5875
rect 757 5870 776 5871
rect 761 5866 762 5870
rect 766 5866 767 5870
rect 771 5866 772 5870
rect 787 5896 788 5900
rect 792 5896 793 5900
rect 797 5896 798 5900
rect 783 5895 802 5896
rect 787 5891 788 5895
rect 792 5891 793 5895
rect 797 5891 798 5895
rect 783 5890 802 5891
rect 787 5886 788 5890
rect 792 5886 793 5890
rect 797 5886 798 5890
rect 783 5885 802 5886
rect 787 5881 788 5885
rect 792 5881 793 5885
rect 797 5881 798 5885
rect 783 5880 802 5881
rect 787 5876 788 5880
rect 792 5876 793 5880
rect 797 5876 798 5880
rect 783 5875 802 5876
rect 787 5871 788 5875
rect 792 5871 793 5875
rect 797 5871 798 5875
rect 783 5870 802 5871
rect 787 5866 788 5870
rect 792 5866 793 5870
rect 797 5866 798 5870
rect 813 5896 814 5900
rect 818 5896 819 5900
rect 823 5896 824 5900
rect 809 5895 828 5896
rect 813 5891 814 5895
rect 818 5891 819 5895
rect 823 5891 824 5895
rect 809 5890 828 5891
rect 813 5886 814 5890
rect 818 5886 819 5890
rect 823 5886 824 5890
rect 809 5885 828 5886
rect 813 5881 814 5885
rect 818 5881 819 5885
rect 823 5881 824 5885
rect 809 5880 828 5881
rect 813 5876 814 5880
rect 818 5876 819 5880
rect 823 5876 824 5880
rect 809 5875 828 5876
rect 813 5871 814 5875
rect 818 5871 819 5875
rect 823 5871 824 5875
rect 809 5870 828 5871
rect 813 5866 814 5870
rect 818 5866 819 5870
rect 823 5866 824 5870
rect 839 5896 840 5900
rect 844 5896 845 5900
rect 849 5896 850 5900
rect 835 5895 854 5896
rect 839 5891 840 5895
rect 844 5891 845 5895
rect 849 5891 850 5895
rect 835 5890 854 5891
rect 839 5886 840 5890
rect 844 5886 845 5890
rect 849 5886 850 5890
rect 835 5885 854 5886
rect 839 5881 840 5885
rect 844 5881 845 5885
rect 849 5881 850 5885
rect 835 5880 854 5881
rect 839 5876 840 5880
rect 844 5876 845 5880
rect 849 5876 850 5880
rect 835 5875 854 5876
rect 839 5871 840 5875
rect 844 5871 845 5875
rect 849 5871 850 5875
rect 835 5870 854 5871
rect 839 5866 840 5870
rect 844 5866 845 5870
rect 849 5866 850 5870
rect 865 5896 866 5900
rect 870 5896 871 5900
rect 875 5896 876 5900
rect 861 5895 880 5896
rect 865 5891 866 5895
rect 870 5891 871 5895
rect 875 5891 876 5895
rect 861 5890 880 5891
rect 865 5886 866 5890
rect 870 5886 871 5890
rect 875 5886 876 5890
rect 861 5885 880 5886
rect 865 5881 866 5885
rect 870 5881 871 5885
rect 875 5881 876 5885
rect 861 5880 880 5881
rect 865 5876 866 5880
rect 870 5876 871 5880
rect 875 5876 876 5880
rect 861 5875 880 5876
rect 865 5871 866 5875
rect 870 5871 871 5875
rect 875 5871 876 5875
rect 861 5870 880 5871
rect 865 5866 866 5870
rect 870 5866 871 5870
rect 875 5866 876 5870
rect 1058 5896 1059 5900
rect 1063 5896 1064 5900
rect 1068 5896 1069 5900
rect 1054 5895 1073 5896
rect 1058 5891 1059 5895
rect 1063 5891 1064 5895
rect 1068 5891 1069 5895
rect 1054 5890 1073 5891
rect 1058 5886 1059 5890
rect 1063 5886 1064 5890
rect 1068 5886 1069 5890
rect 1054 5885 1073 5886
rect 1058 5881 1059 5885
rect 1063 5881 1064 5885
rect 1068 5881 1069 5885
rect 1054 5880 1073 5881
rect 1058 5876 1059 5880
rect 1063 5876 1064 5880
rect 1068 5876 1069 5880
rect 1054 5875 1073 5876
rect 1058 5871 1059 5875
rect 1063 5871 1064 5875
rect 1068 5871 1069 5875
rect 1054 5870 1073 5871
rect 1058 5866 1059 5870
rect 1063 5866 1064 5870
rect 1068 5866 1069 5870
rect 761 5850 762 5854
rect 766 5850 767 5854
rect 771 5850 772 5854
rect 757 5849 776 5850
rect 761 5845 762 5849
rect 766 5845 767 5849
rect 771 5845 772 5849
rect 757 5844 776 5845
rect 761 5840 762 5844
rect 766 5840 767 5844
rect 771 5840 772 5844
rect 757 5839 776 5840
rect 761 5835 762 5839
rect 766 5835 767 5839
rect 771 5835 772 5839
rect 757 5834 776 5835
rect 761 5830 762 5834
rect 766 5830 767 5834
rect 771 5830 772 5834
rect 757 5829 776 5830
rect 761 5825 762 5829
rect 766 5825 767 5829
rect 771 5825 772 5829
rect 757 5824 776 5825
rect 761 5820 762 5824
rect 766 5820 767 5824
rect 771 5820 772 5824
rect 787 5850 788 5854
rect 792 5850 793 5854
rect 797 5850 798 5854
rect 783 5849 802 5850
rect 787 5845 788 5849
rect 792 5845 793 5849
rect 797 5845 798 5849
rect 783 5844 802 5845
rect 787 5840 788 5844
rect 792 5840 793 5844
rect 797 5840 798 5844
rect 783 5839 802 5840
rect 787 5835 788 5839
rect 792 5835 793 5839
rect 797 5835 798 5839
rect 783 5834 802 5835
rect 787 5830 788 5834
rect 792 5830 793 5834
rect 797 5830 798 5834
rect 783 5829 802 5830
rect 787 5825 788 5829
rect 792 5825 793 5829
rect 797 5825 798 5829
rect 783 5824 802 5825
rect 787 5820 788 5824
rect 792 5820 793 5824
rect 797 5820 798 5824
rect 813 5850 814 5854
rect 818 5850 819 5854
rect 823 5850 824 5854
rect 809 5849 828 5850
rect 813 5845 814 5849
rect 818 5845 819 5849
rect 823 5845 824 5849
rect 809 5844 828 5845
rect 813 5840 814 5844
rect 818 5840 819 5844
rect 823 5840 824 5844
rect 809 5839 828 5840
rect 813 5835 814 5839
rect 818 5835 819 5839
rect 823 5835 824 5839
rect 809 5834 828 5835
rect 813 5830 814 5834
rect 818 5830 819 5834
rect 823 5830 824 5834
rect 809 5829 828 5830
rect 813 5825 814 5829
rect 818 5825 819 5829
rect 823 5825 824 5829
rect 809 5824 828 5825
rect 813 5820 814 5824
rect 818 5820 819 5824
rect 823 5820 824 5824
rect 839 5850 840 5854
rect 844 5850 845 5854
rect 849 5850 850 5854
rect 835 5849 854 5850
rect 839 5845 840 5849
rect 844 5845 845 5849
rect 849 5845 850 5849
rect 835 5844 854 5845
rect 839 5840 840 5844
rect 844 5840 845 5844
rect 849 5840 850 5844
rect 835 5839 854 5840
rect 839 5835 840 5839
rect 844 5835 845 5839
rect 849 5835 850 5839
rect 835 5834 854 5835
rect 839 5830 840 5834
rect 844 5830 845 5834
rect 849 5830 850 5834
rect 835 5829 854 5830
rect 839 5825 840 5829
rect 844 5825 845 5829
rect 849 5825 850 5829
rect 835 5824 854 5825
rect 839 5820 840 5824
rect 844 5820 845 5824
rect 849 5820 850 5824
rect 865 5850 866 5854
rect 870 5850 871 5854
rect 875 5850 876 5854
rect 861 5849 880 5850
rect 865 5845 866 5849
rect 870 5845 871 5849
rect 875 5845 876 5849
rect 861 5844 880 5845
rect 865 5840 866 5844
rect 870 5840 871 5844
rect 875 5840 876 5844
rect 861 5839 880 5840
rect 865 5835 866 5839
rect 870 5835 871 5839
rect 875 5835 876 5839
rect 861 5834 880 5835
rect 865 5830 866 5834
rect 870 5830 871 5834
rect 875 5830 876 5834
rect 861 5829 880 5830
rect 865 5825 866 5829
rect 870 5825 871 5829
rect 875 5825 876 5829
rect 861 5824 880 5825
rect 865 5820 866 5824
rect 870 5820 871 5824
rect 875 5820 876 5824
rect 1058 5850 1059 5854
rect 1063 5850 1064 5854
rect 1068 5850 1069 5854
rect 1054 5849 1073 5850
rect 1058 5845 1059 5849
rect 1063 5845 1064 5849
rect 1068 5845 1069 5849
rect 1054 5844 1073 5845
rect 1058 5840 1059 5844
rect 1063 5840 1064 5844
rect 1068 5840 1069 5844
rect 1054 5839 1073 5840
rect 1058 5835 1059 5839
rect 1063 5835 1064 5839
rect 1068 5835 1069 5839
rect 1054 5834 1073 5835
rect 1058 5830 1059 5834
rect 1063 5830 1064 5834
rect 1068 5830 1069 5834
rect 1054 5829 1073 5830
rect 1058 5825 1059 5829
rect 1063 5825 1064 5829
rect 1068 5825 1069 5829
rect 1054 5824 1073 5825
rect 1058 5820 1059 5824
rect 1063 5820 1064 5824
rect 1068 5820 1069 5824
rect 99 5325 1031 5800
rect 1154 5593 1250 5976
rect 1367 5896 1368 5900
rect 1372 5896 1373 5900
rect 1377 5896 1378 5900
rect 1363 5895 1382 5896
rect 1367 5891 1368 5895
rect 1372 5891 1373 5895
rect 1377 5891 1378 5895
rect 1363 5890 1382 5891
rect 1367 5886 1368 5890
rect 1372 5886 1373 5890
rect 1377 5886 1378 5890
rect 1363 5885 1382 5886
rect 1367 5881 1368 5885
rect 1372 5881 1373 5885
rect 1377 5881 1378 5885
rect 1363 5880 1382 5881
rect 1367 5876 1368 5880
rect 1372 5876 1373 5880
rect 1377 5876 1378 5880
rect 1363 5875 1382 5876
rect 1367 5871 1368 5875
rect 1372 5871 1373 5875
rect 1377 5871 1378 5875
rect 1363 5870 1382 5871
rect 1367 5866 1368 5870
rect 1372 5866 1373 5870
rect 1377 5866 1378 5870
rect 1367 5850 1368 5854
rect 1372 5850 1373 5854
rect 1377 5850 1378 5854
rect 1363 5849 1382 5850
rect 1367 5845 1368 5849
rect 1372 5845 1373 5849
rect 1377 5845 1378 5849
rect 1363 5844 1382 5845
rect 1367 5840 1368 5844
rect 1372 5840 1373 5844
rect 1377 5840 1378 5844
rect 1363 5839 1382 5840
rect 1367 5835 1368 5839
rect 1372 5835 1373 5839
rect 1377 5835 1378 5839
rect 1363 5834 1382 5835
rect 1367 5830 1368 5834
rect 1372 5830 1373 5834
rect 1377 5830 1378 5834
rect 1363 5829 1382 5830
rect 1367 5825 1368 5829
rect 1372 5825 1373 5829
rect 1377 5825 1378 5829
rect 1363 5824 1382 5825
rect 1367 5820 1368 5824
rect 1372 5820 1373 5824
rect 1377 5820 1378 5824
rect 1463 5593 1559 5976
rect 1676 5896 1677 5900
rect 1681 5896 1682 5900
rect 1686 5896 1687 5900
rect 1672 5895 1691 5896
rect 1676 5891 1677 5895
rect 1681 5891 1682 5895
rect 1686 5891 1687 5895
rect 1672 5890 1691 5891
rect 1676 5886 1677 5890
rect 1681 5886 1682 5890
rect 1686 5886 1687 5890
rect 1672 5885 1691 5886
rect 1676 5881 1677 5885
rect 1681 5881 1682 5885
rect 1686 5881 1687 5885
rect 1672 5880 1691 5881
rect 1676 5876 1677 5880
rect 1681 5876 1682 5880
rect 1686 5876 1687 5880
rect 1672 5875 1691 5876
rect 1676 5871 1677 5875
rect 1681 5871 1682 5875
rect 1686 5871 1687 5875
rect 1672 5870 1691 5871
rect 1676 5866 1677 5870
rect 1681 5866 1682 5870
rect 1686 5866 1687 5870
rect 1676 5850 1677 5854
rect 1681 5850 1682 5854
rect 1686 5850 1687 5854
rect 1672 5849 1691 5850
rect 1676 5845 1677 5849
rect 1681 5845 1682 5849
rect 1686 5845 1687 5849
rect 1672 5844 1691 5845
rect 1676 5840 1677 5844
rect 1681 5840 1682 5844
rect 1686 5840 1687 5844
rect 1672 5839 1691 5840
rect 1676 5835 1677 5839
rect 1681 5835 1682 5839
rect 1686 5835 1687 5839
rect 1672 5834 1691 5835
rect 1676 5830 1677 5834
rect 1681 5830 1682 5834
rect 1686 5830 1687 5834
rect 1672 5829 1691 5830
rect 1676 5825 1677 5829
rect 1681 5825 1682 5829
rect 1686 5825 1687 5829
rect 1672 5824 1691 5825
rect 1676 5820 1677 5824
rect 1681 5820 1682 5824
rect 1686 5820 1687 5824
rect 1772 5593 1868 5976
rect 1985 5896 1986 5900
rect 1990 5896 1991 5900
rect 1995 5896 1996 5900
rect 1981 5895 2000 5896
rect 1985 5891 1986 5895
rect 1990 5891 1991 5895
rect 1995 5891 1996 5895
rect 1981 5890 2000 5891
rect 1985 5886 1986 5890
rect 1990 5886 1991 5890
rect 1995 5886 1996 5890
rect 1981 5885 2000 5886
rect 1985 5881 1986 5885
rect 1990 5881 1991 5885
rect 1995 5881 1996 5885
rect 1981 5880 2000 5881
rect 1985 5876 1986 5880
rect 1990 5876 1991 5880
rect 1995 5876 1996 5880
rect 1981 5875 2000 5876
rect 1985 5871 1986 5875
rect 1990 5871 1991 5875
rect 1995 5871 1996 5875
rect 1981 5870 2000 5871
rect 1985 5866 1986 5870
rect 1990 5866 1991 5870
rect 1995 5866 1996 5870
rect 1985 5850 1986 5854
rect 1990 5850 1991 5854
rect 1995 5850 1996 5854
rect 1981 5849 2000 5850
rect 1985 5845 1986 5849
rect 1990 5845 1991 5849
rect 1995 5845 1996 5849
rect 1981 5844 2000 5845
rect 1985 5840 1986 5844
rect 1990 5840 1991 5844
rect 1995 5840 1996 5844
rect 1981 5839 2000 5840
rect 1985 5835 1986 5839
rect 1990 5835 1991 5839
rect 1995 5835 1996 5839
rect 1981 5834 2000 5835
rect 1985 5830 1986 5834
rect 1990 5830 1991 5834
rect 1995 5830 1996 5834
rect 1981 5829 2000 5830
rect 1985 5825 1986 5829
rect 1990 5825 1991 5829
rect 1995 5825 1996 5829
rect 1981 5824 2000 5825
rect 1985 5820 1986 5824
rect 1990 5820 1991 5824
rect 1995 5820 1996 5824
rect 2081 5593 2177 5976
rect 2294 5896 2295 5900
rect 2299 5896 2300 5900
rect 2304 5896 2305 5900
rect 2290 5895 2309 5896
rect 2294 5891 2295 5895
rect 2299 5891 2300 5895
rect 2304 5891 2305 5895
rect 2290 5890 2309 5891
rect 2294 5886 2295 5890
rect 2299 5886 2300 5890
rect 2304 5886 2305 5890
rect 2290 5885 2309 5886
rect 2294 5881 2295 5885
rect 2299 5881 2300 5885
rect 2304 5881 2305 5885
rect 2290 5880 2309 5881
rect 2294 5876 2295 5880
rect 2299 5876 2300 5880
rect 2304 5876 2305 5880
rect 2290 5875 2309 5876
rect 2294 5871 2295 5875
rect 2299 5871 2300 5875
rect 2304 5871 2305 5875
rect 2290 5870 2309 5871
rect 2294 5866 2295 5870
rect 2299 5866 2300 5870
rect 2304 5866 2305 5870
rect 2294 5850 2295 5854
rect 2299 5850 2300 5854
rect 2304 5850 2305 5854
rect 2290 5849 2309 5850
rect 2294 5845 2295 5849
rect 2299 5845 2300 5849
rect 2304 5845 2305 5849
rect 2290 5844 2309 5845
rect 2294 5840 2295 5844
rect 2299 5840 2300 5844
rect 2304 5840 2305 5844
rect 2290 5839 2309 5840
rect 2294 5835 2295 5839
rect 2299 5835 2300 5839
rect 2304 5835 2305 5839
rect 2290 5834 2309 5835
rect 2294 5830 2295 5834
rect 2299 5830 2300 5834
rect 2304 5830 2305 5834
rect 2290 5829 2309 5830
rect 2294 5825 2295 5829
rect 2299 5825 2300 5829
rect 2304 5825 2305 5829
rect 2290 5824 2309 5825
rect 2294 5820 2295 5824
rect 2299 5820 2300 5824
rect 2304 5820 2305 5824
rect 2390 5593 2486 5976
rect 2603 5896 2604 5900
rect 2608 5896 2609 5900
rect 2613 5896 2614 5900
rect 2599 5895 2618 5896
rect 2603 5891 2604 5895
rect 2608 5891 2609 5895
rect 2613 5891 2614 5895
rect 2599 5890 2618 5891
rect 2603 5886 2604 5890
rect 2608 5886 2609 5890
rect 2613 5886 2614 5890
rect 2599 5885 2618 5886
rect 2603 5881 2604 5885
rect 2608 5881 2609 5885
rect 2613 5881 2614 5885
rect 2599 5880 2618 5881
rect 2603 5876 2604 5880
rect 2608 5876 2609 5880
rect 2613 5876 2614 5880
rect 2599 5875 2618 5876
rect 2603 5871 2604 5875
rect 2608 5871 2609 5875
rect 2613 5871 2614 5875
rect 2599 5870 2618 5871
rect 2603 5866 2604 5870
rect 2608 5866 2609 5870
rect 2613 5866 2614 5870
rect 2603 5850 2604 5854
rect 2608 5850 2609 5854
rect 2613 5850 2614 5854
rect 2599 5849 2618 5850
rect 2603 5845 2604 5849
rect 2608 5845 2609 5849
rect 2613 5845 2614 5849
rect 2599 5844 2618 5845
rect 2603 5840 2604 5844
rect 2608 5840 2609 5844
rect 2613 5840 2614 5844
rect 2599 5839 2618 5840
rect 2603 5835 2604 5839
rect 2608 5835 2609 5839
rect 2613 5835 2614 5839
rect 2599 5834 2618 5835
rect 2603 5830 2604 5834
rect 2608 5830 2609 5834
rect 2613 5830 2614 5834
rect 2599 5829 2618 5830
rect 2603 5825 2604 5829
rect 2608 5825 2609 5829
rect 2613 5825 2614 5829
rect 2599 5824 2618 5825
rect 2603 5820 2604 5824
rect 2608 5820 2609 5824
rect 2613 5820 2614 5824
rect 2699 5593 2795 5976
rect 2912 5896 2913 5900
rect 2917 5896 2918 5900
rect 2922 5896 2923 5900
rect 2908 5895 2927 5896
rect 2912 5891 2913 5895
rect 2917 5891 2918 5895
rect 2922 5891 2923 5895
rect 2908 5890 2927 5891
rect 2912 5886 2913 5890
rect 2917 5886 2918 5890
rect 2922 5886 2923 5890
rect 2908 5885 2927 5886
rect 2912 5881 2913 5885
rect 2917 5881 2918 5885
rect 2922 5881 2923 5885
rect 2908 5880 2927 5881
rect 2912 5876 2913 5880
rect 2917 5876 2918 5880
rect 2922 5876 2923 5880
rect 2908 5875 2927 5876
rect 2912 5871 2913 5875
rect 2917 5871 2918 5875
rect 2922 5871 2923 5875
rect 2908 5870 2927 5871
rect 2912 5866 2913 5870
rect 2917 5866 2918 5870
rect 2922 5866 2923 5870
rect 2912 5850 2913 5854
rect 2917 5850 2918 5854
rect 2922 5850 2923 5854
rect 2908 5849 2927 5850
rect 2912 5845 2913 5849
rect 2917 5845 2918 5849
rect 2922 5845 2923 5849
rect 2908 5844 2927 5845
rect 2912 5840 2913 5844
rect 2917 5840 2918 5844
rect 2922 5840 2923 5844
rect 2908 5839 2927 5840
rect 2912 5835 2913 5839
rect 2917 5835 2918 5839
rect 2922 5835 2923 5839
rect 2908 5834 2927 5835
rect 2912 5830 2913 5834
rect 2917 5830 2918 5834
rect 2922 5830 2923 5834
rect 2908 5829 2927 5830
rect 2912 5825 2913 5829
rect 2917 5825 2918 5829
rect 2922 5825 2923 5829
rect 2908 5824 2927 5825
rect 2912 5820 2913 5824
rect 2917 5820 2918 5824
rect 2922 5820 2923 5824
rect 3008 5593 3104 5976
rect 3221 5896 3222 5900
rect 3226 5896 3227 5900
rect 3231 5896 3232 5900
rect 3217 5895 3236 5896
rect 3221 5891 3222 5895
rect 3226 5891 3227 5895
rect 3231 5891 3232 5895
rect 3217 5890 3236 5891
rect 3221 5886 3222 5890
rect 3226 5886 3227 5890
rect 3231 5886 3232 5890
rect 3217 5885 3236 5886
rect 3221 5881 3222 5885
rect 3226 5881 3227 5885
rect 3231 5881 3232 5885
rect 3217 5880 3236 5881
rect 3221 5876 3222 5880
rect 3226 5876 3227 5880
rect 3231 5876 3232 5880
rect 3217 5875 3236 5876
rect 3221 5871 3222 5875
rect 3226 5871 3227 5875
rect 3231 5871 3232 5875
rect 3217 5870 3236 5871
rect 3221 5866 3222 5870
rect 3226 5866 3227 5870
rect 3231 5866 3232 5870
rect 3221 5850 3222 5854
rect 3226 5850 3227 5854
rect 3231 5850 3232 5854
rect 3217 5849 3236 5850
rect 3221 5845 3222 5849
rect 3226 5845 3227 5849
rect 3231 5845 3232 5849
rect 3217 5844 3236 5845
rect 3221 5840 3222 5844
rect 3226 5840 3227 5844
rect 3231 5840 3232 5844
rect 3217 5839 3236 5840
rect 3221 5835 3222 5839
rect 3226 5835 3227 5839
rect 3231 5835 3232 5839
rect 3217 5834 3236 5835
rect 3221 5830 3222 5834
rect 3226 5830 3227 5834
rect 3231 5830 3232 5834
rect 3217 5829 3236 5830
rect 3221 5825 3222 5829
rect 3226 5825 3227 5829
rect 3231 5825 3232 5829
rect 3217 5824 3236 5825
rect 3221 5820 3222 5824
rect 3226 5820 3227 5824
rect 3231 5820 3232 5824
rect 3317 5593 3413 5976
rect 3530 5896 3531 5900
rect 3535 5896 3536 5900
rect 3540 5896 3541 5900
rect 3526 5895 3545 5896
rect 3530 5891 3531 5895
rect 3535 5891 3536 5895
rect 3540 5891 3541 5895
rect 3526 5890 3545 5891
rect 3530 5886 3531 5890
rect 3535 5886 3536 5890
rect 3540 5886 3541 5890
rect 3526 5885 3545 5886
rect 3530 5881 3531 5885
rect 3535 5881 3536 5885
rect 3540 5881 3541 5885
rect 3526 5880 3545 5881
rect 3530 5876 3531 5880
rect 3535 5876 3536 5880
rect 3540 5876 3541 5880
rect 3526 5875 3545 5876
rect 3530 5871 3531 5875
rect 3535 5871 3536 5875
rect 3540 5871 3541 5875
rect 3526 5870 3545 5871
rect 3530 5866 3531 5870
rect 3535 5866 3536 5870
rect 3540 5866 3541 5870
rect 3530 5850 3531 5854
rect 3535 5850 3536 5854
rect 3540 5850 3541 5854
rect 3526 5849 3545 5850
rect 3530 5845 3531 5849
rect 3535 5845 3536 5849
rect 3540 5845 3541 5849
rect 3526 5844 3545 5845
rect 3530 5840 3531 5844
rect 3535 5840 3536 5844
rect 3540 5840 3541 5844
rect 3526 5839 3545 5840
rect 3530 5835 3531 5839
rect 3535 5835 3536 5839
rect 3540 5835 3541 5839
rect 3526 5834 3545 5835
rect 3530 5830 3531 5834
rect 3535 5830 3536 5834
rect 3540 5830 3541 5834
rect 3526 5829 3545 5830
rect 3530 5825 3531 5829
rect 3535 5825 3536 5829
rect 3540 5825 3541 5829
rect 3526 5824 3545 5825
rect 3530 5820 3531 5824
rect 3535 5820 3536 5824
rect 3540 5820 3541 5824
rect 3626 5593 3722 5976
rect 3839 5896 3840 5900
rect 3844 5896 3845 5900
rect 3849 5896 3850 5900
rect 3835 5895 3854 5896
rect 3839 5891 3840 5895
rect 3844 5891 3845 5895
rect 3849 5891 3850 5895
rect 3835 5890 3854 5891
rect 3839 5886 3840 5890
rect 3844 5886 3845 5890
rect 3849 5886 3850 5890
rect 3835 5885 3854 5886
rect 3839 5881 3840 5885
rect 3844 5881 3845 5885
rect 3849 5881 3850 5885
rect 3835 5880 3854 5881
rect 3839 5876 3840 5880
rect 3844 5876 3845 5880
rect 3849 5876 3850 5880
rect 3835 5875 3854 5876
rect 3839 5871 3840 5875
rect 3844 5871 3845 5875
rect 3849 5871 3850 5875
rect 3835 5870 3854 5871
rect 3839 5866 3840 5870
rect 3844 5866 3845 5870
rect 3849 5866 3850 5870
rect 3839 5850 3840 5854
rect 3844 5850 3845 5854
rect 3849 5850 3850 5854
rect 3835 5849 3854 5850
rect 3839 5845 3840 5849
rect 3844 5845 3845 5849
rect 3849 5845 3850 5849
rect 3835 5844 3854 5845
rect 3839 5840 3840 5844
rect 3844 5840 3845 5844
rect 3849 5840 3850 5844
rect 3835 5839 3854 5840
rect 3839 5835 3840 5839
rect 3844 5835 3845 5839
rect 3849 5835 3850 5839
rect 3835 5834 3854 5835
rect 3839 5830 3840 5834
rect 3844 5830 3845 5834
rect 3849 5830 3850 5834
rect 3835 5829 3854 5830
rect 3839 5825 3840 5829
rect 3844 5825 3845 5829
rect 3849 5825 3850 5829
rect 3835 5824 3854 5825
rect 3839 5820 3840 5824
rect 3844 5820 3845 5824
rect 3849 5820 3850 5824
rect 3935 5593 4031 5976
rect 4483 5974 4484 5978
rect 4488 5974 4489 5978
rect 4493 5974 4494 5978
rect 4498 5974 4499 5978
rect 4503 5974 4504 5978
rect 4508 5974 4509 5978
rect 4479 5973 4513 5974
rect 4483 5969 4484 5973
rect 4488 5969 4489 5973
rect 4493 5969 4494 5973
rect 4498 5969 4499 5973
rect 4503 5969 4504 5973
rect 4508 5969 4509 5973
rect 4479 5968 4513 5969
rect 4483 5964 4484 5968
rect 4488 5964 4489 5968
rect 4493 5964 4494 5968
rect 4498 5964 4499 5968
rect 4503 5964 4504 5968
rect 4508 5964 4509 5968
rect 4529 5979 4530 5983
rect 4534 5979 4535 5983
rect 4539 5979 4540 5983
rect 4544 5979 4545 5983
rect 4549 5979 4550 5983
rect 4554 5979 4555 5983
rect 4525 5978 4559 5979
rect 4529 5974 4530 5978
rect 4534 5974 4535 5978
rect 4539 5974 4540 5978
rect 4544 5974 4545 5978
rect 4549 5974 4550 5978
rect 4554 5974 4555 5978
rect 4525 5973 4559 5974
rect 4529 5969 4530 5973
rect 4534 5969 4535 5973
rect 4539 5969 4540 5973
rect 4544 5969 4545 5973
rect 4549 5969 4550 5973
rect 4554 5969 4555 5973
rect 4525 5968 4559 5969
rect 4529 5964 4530 5968
rect 4534 5964 4535 5968
rect 4539 5964 4540 5968
rect 4544 5964 4545 5968
rect 4549 5964 4550 5968
rect 4554 5964 4555 5968
rect 4239 5896 4240 5900
rect 4244 5896 4245 5900
rect 4249 5896 4250 5900
rect 4235 5895 4254 5896
rect 4239 5891 4240 5895
rect 4244 5891 4245 5895
rect 4249 5891 4250 5895
rect 4235 5890 4254 5891
rect 4239 5886 4240 5890
rect 4244 5886 4245 5890
rect 4249 5886 4250 5890
rect 4235 5885 4254 5886
rect 4239 5881 4240 5885
rect 4244 5881 4245 5885
rect 4249 5881 4250 5885
rect 4235 5880 4254 5881
rect 4239 5876 4240 5880
rect 4244 5876 4245 5880
rect 4249 5876 4250 5880
rect 4235 5875 4254 5876
rect 4239 5871 4240 5875
rect 4244 5871 4245 5875
rect 4249 5871 4250 5875
rect 4235 5870 4254 5871
rect 4239 5866 4240 5870
rect 4244 5866 4245 5870
rect 4249 5866 4250 5870
rect 4268 5896 4269 5900
rect 4273 5896 4274 5900
rect 4278 5896 4279 5900
rect 4264 5895 4283 5896
rect 4268 5891 4269 5895
rect 4273 5891 4274 5895
rect 4278 5891 4279 5895
rect 4264 5890 4283 5891
rect 4268 5886 4269 5890
rect 4273 5886 4274 5890
rect 4278 5886 4279 5890
rect 4264 5885 4283 5886
rect 4268 5881 4269 5885
rect 4273 5881 4274 5885
rect 4278 5881 4279 5885
rect 4264 5880 4283 5881
rect 4268 5876 4269 5880
rect 4273 5876 4274 5880
rect 4278 5876 4279 5880
rect 4264 5875 4283 5876
rect 4268 5871 4269 5875
rect 4273 5871 4274 5875
rect 4278 5871 4279 5875
rect 4264 5870 4283 5871
rect 4268 5866 4269 5870
rect 4273 5866 4274 5870
rect 4278 5866 4279 5870
rect 4297 5896 4298 5900
rect 4302 5896 4303 5900
rect 4307 5896 4308 5900
rect 4293 5895 4312 5896
rect 4297 5891 4298 5895
rect 4302 5891 4303 5895
rect 4307 5891 4308 5895
rect 4293 5890 4312 5891
rect 4297 5886 4298 5890
rect 4302 5886 4303 5890
rect 4307 5886 4308 5890
rect 4293 5885 4312 5886
rect 4297 5881 4298 5885
rect 4302 5881 4303 5885
rect 4307 5881 4308 5885
rect 4293 5880 4312 5881
rect 4297 5876 4298 5880
rect 4302 5876 4303 5880
rect 4307 5876 4308 5880
rect 4293 5875 4312 5876
rect 4297 5871 4298 5875
rect 4302 5871 4303 5875
rect 4307 5871 4308 5875
rect 4293 5870 4312 5871
rect 4297 5866 4298 5870
rect 4302 5866 4303 5870
rect 4307 5866 4308 5870
rect 4326 5896 4327 5900
rect 4331 5896 4332 5900
rect 4336 5896 4337 5900
rect 4322 5895 4341 5896
rect 4326 5891 4327 5895
rect 4331 5891 4332 5895
rect 4336 5891 4337 5895
rect 4322 5890 4341 5891
rect 4326 5886 4327 5890
rect 4331 5886 4332 5890
rect 4336 5886 4337 5890
rect 4322 5885 4341 5886
rect 4326 5881 4327 5885
rect 4331 5881 4332 5885
rect 4336 5881 4337 5885
rect 4322 5880 4341 5881
rect 4326 5876 4327 5880
rect 4331 5876 4332 5880
rect 4336 5876 4337 5880
rect 4322 5875 4341 5876
rect 4326 5871 4327 5875
rect 4331 5871 4332 5875
rect 4336 5871 4337 5875
rect 4322 5870 4341 5871
rect 4326 5866 4327 5870
rect 4331 5866 4332 5870
rect 4336 5866 4337 5870
rect 4355 5896 4356 5900
rect 4360 5896 4361 5900
rect 4365 5896 4366 5900
rect 4351 5895 4370 5896
rect 4355 5891 4356 5895
rect 4360 5891 4361 5895
rect 4365 5891 4366 5895
rect 4351 5890 4370 5891
rect 4355 5886 4356 5890
rect 4360 5886 4361 5890
rect 4365 5886 4366 5890
rect 4351 5885 4370 5886
rect 4355 5881 4356 5885
rect 4360 5881 4361 5885
rect 4365 5881 4366 5885
rect 4351 5880 4370 5881
rect 4355 5876 4356 5880
rect 4360 5876 4361 5880
rect 4365 5876 4366 5880
rect 4351 5875 4370 5876
rect 4355 5871 4356 5875
rect 4360 5871 4361 5875
rect 4365 5871 4366 5875
rect 4351 5870 4370 5871
rect 4355 5866 4356 5870
rect 4360 5866 4361 5870
rect 4365 5866 4366 5870
rect 4239 5850 4240 5854
rect 4244 5850 4245 5854
rect 4249 5850 4250 5854
rect 4235 5849 4254 5850
rect 4239 5845 4240 5849
rect 4244 5845 4245 5849
rect 4249 5845 4250 5849
rect 4235 5844 4254 5845
rect 4239 5840 4240 5844
rect 4244 5840 4245 5844
rect 4249 5840 4250 5844
rect 4235 5839 4254 5840
rect 4239 5835 4240 5839
rect 4244 5835 4245 5839
rect 4249 5835 4250 5839
rect 4235 5834 4254 5835
rect 4239 5830 4240 5834
rect 4244 5830 4245 5834
rect 4249 5830 4250 5834
rect 4235 5829 4254 5830
rect 4239 5825 4240 5829
rect 4244 5825 4245 5829
rect 4249 5825 4250 5829
rect 4235 5824 4254 5825
rect 4239 5820 4240 5824
rect 4244 5820 4245 5824
rect 4249 5820 4250 5824
rect 4268 5850 4269 5854
rect 4273 5850 4274 5854
rect 4278 5850 4279 5854
rect 4264 5849 4283 5850
rect 4268 5845 4269 5849
rect 4273 5845 4274 5849
rect 4278 5845 4279 5849
rect 4264 5844 4283 5845
rect 4268 5840 4269 5844
rect 4273 5840 4274 5844
rect 4278 5840 4279 5844
rect 4264 5839 4283 5840
rect 4268 5835 4269 5839
rect 4273 5835 4274 5839
rect 4278 5835 4279 5839
rect 4264 5834 4283 5835
rect 4268 5830 4269 5834
rect 4273 5830 4274 5834
rect 4278 5830 4279 5834
rect 4264 5829 4283 5830
rect 4268 5825 4269 5829
rect 4273 5825 4274 5829
rect 4278 5825 4279 5829
rect 4264 5824 4283 5825
rect 4268 5820 4269 5824
rect 4273 5820 4274 5824
rect 4278 5820 4279 5824
rect 4297 5850 4298 5854
rect 4302 5850 4303 5854
rect 4307 5850 4308 5854
rect 4293 5849 4312 5850
rect 4297 5845 4298 5849
rect 4302 5845 4303 5849
rect 4307 5845 4308 5849
rect 4293 5844 4312 5845
rect 4297 5840 4298 5844
rect 4302 5840 4303 5844
rect 4307 5840 4308 5844
rect 4293 5839 4312 5840
rect 4297 5835 4298 5839
rect 4302 5835 4303 5839
rect 4307 5835 4308 5839
rect 4293 5834 4312 5835
rect 4297 5830 4298 5834
rect 4302 5830 4303 5834
rect 4307 5830 4308 5834
rect 4293 5829 4312 5830
rect 4297 5825 4298 5829
rect 4302 5825 4303 5829
rect 4307 5825 4308 5829
rect 4293 5824 4312 5825
rect 4297 5820 4298 5824
rect 4302 5820 4303 5824
rect 4307 5820 4308 5824
rect 4326 5850 4327 5854
rect 4331 5850 4332 5854
rect 4336 5850 4337 5854
rect 4322 5849 4341 5850
rect 4326 5845 4327 5849
rect 4331 5845 4332 5849
rect 4336 5845 4337 5849
rect 4322 5844 4341 5845
rect 4326 5840 4327 5844
rect 4331 5840 4332 5844
rect 4336 5840 4337 5844
rect 4322 5839 4341 5840
rect 4326 5835 4327 5839
rect 4331 5835 4332 5839
rect 4336 5835 4337 5839
rect 4322 5834 4341 5835
rect 4326 5830 4327 5834
rect 4331 5830 4332 5834
rect 4336 5830 4337 5834
rect 4322 5829 4341 5830
rect 4326 5825 4327 5829
rect 4331 5825 4332 5829
rect 4336 5825 4337 5829
rect 4322 5824 4341 5825
rect 4326 5820 4327 5824
rect 4331 5820 4332 5824
rect 4336 5820 4337 5824
rect 4355 5850 4356 5854
rect 4360 5850 4361 5854
rect 4365 5850 4366 5854
rect 4351 5849 4370 5850
rect 4355 5845 4356 5849
rect 4360 5845 4361 5849
rect 4365 5845 4366 5849
rect 4351 5844 4370 5845
rect 4355 5840 4356 5844
rect 4360 5840 4361 5844
rect 4365 5840 4366 5844
rect 4351 5839 4370 5840
rect 4355 5835 4356 5839
rect 4360 5835 4361 5839
rect 4365 5835 4366 5839
rect 4351 5834 4370 5835
rect 4355 5830 4356 5834
rect 4360 5830 4361 5834
rect 4365 5830 4366 5834
rect 4351 5829 4370 5830
rect 4355 5825 4356 5829
rect 4360 5825 4361 5829
rect 4365 5825 4366 5829
rect 4351 5824 4370 5825
rect 4355 5820 4356 5824
rect 4360 5820 4361 5824
rect 4365 5820 4366 5824
rect 4579 5800 5054 6238
rect 1144 5583 1260 5593
rect 1453 5583 1569 5593
rect 1762 5583 1878 5593
rect 2071 5583 2187 5593
rect 2380 5583 2496 5593
rect 2689 5583 2805 5593
rect 2998 5583 3114 5593
rect 3307 5583 3423 5593
rect 3616 5583 3732 5593
rect 3925 5583 4041 5593
rect 1134 5573 1270 5583
rect 1443 5573 1579 5583
rect 1752 5573 1888 5583
rect 2061 5573 2197 5583
rect 2370 5573 2506 5583
rect 2679 5573 2815 5583
rect 2988 5573 3124 5583
rect 3297 5573 3433 5583
rect 3606 5573 3742 5583
rect 3915 5573 4051 5583
rect 1124 5563 1280 5573
rect 1433 5563 1589 5573
rect 1742 5563 1898 5573
rect 2051 5563 2207 5573
rect 2360 5563 2516 5573
rect 2669 5563 2825 5573
rect 2978 5563 3134 5573
rect 3287 5563 3443 5573
rect 3596 5563 3752 5573
rect 3905 5563 4061 5573
rect 1114 5553 1290 5563
rect 1423 5553 1599 5563
rect 1732 5553 1908 5563
rect 2041 5553 2217 5563
rect 2350 5553 2526 5563
rect 2659 5553 2835 5563
rect 2968 5553 3144 5563
rect 3277 5553 3453 5563
rect 3586 5553 3762 5563
rect 3895 5553 4071 5563
rect 1072 5550 1332 5553
rect 1072 5296 1075 5550
rect 1329 5296 1332 5550
rect 1072 5293 1332 5296
rect 1381 5550 1641 5553
rect 1381 5296 1384 5550
rect 1638 5296 1641 5550
rect 1381 5293 1641 5296
rect 1690 5550 1950 5553
rect 1690 5296 1693 5550
rect 1947 5296 1950 5550
rect 1690 5293 1950 5296
rect 1999 5550 2259 5553
rect 1999 5296 2002 5550
rect 2256 5296 2259 5550
rect 1999 5293 2259 5296
rect 2308 5550 2568 5553
rect 2308 5296 2311 5550
rect 2565 5296 2568 5550
rect 2308 5293 2568 5296
rect 2617 5550 2877 5553
rect 2617 5296 2620 5550
rect 2874 5296 2877 5550
rect 2617 5293 2877 5296
rect 2926 5550 3186 5553
rect 2926 5296 2929 5550
rect 3183 5296 3186 5550
rect 2926 5293 3186 5296
rect 3235 5550 3495 5553
rect 3235 5296 3238 5550
rect 3492 5296 3495 5550
rect 3235 5293 3495 5296
rect 3544 5550 3804 5553
rect 3544 5296 3547 5550
rect 3801 5296 3804 5550
rect 3544 5293 3804 5296
rect 3853 5550 4113 5553
rect 3853 5296 3856 5550
rect 4110 5296 4113 5550
rect 4148 5306 5054 5800
rect 3853 5293 4113 5296
<< m2contact >>
rect 1454 9997 1458 10001
rect 1461 9997 1465 10001
rect 1468 9997 1472 10001
rect 1475 9997 1479 10001
rect 1482 9997 1486 10001
rect 1489 9997 1493 10001
rect 1496 9997 1500 10001
rect 1503 9997 1507 10001
rect 1510 9997 1514 10001
rect 1517 9997 1521 10001
rect 1524 9997 1528 10001
rect 1531 9997 1535 10001
rect 1538 9997 1542 10001
rect 802 9757 806 9761
rect 807 9757 811 9761
rect 812 9757 816 9761
rect 817 9757 821 9761
rect 802 9747 806 9751
rect 807 9747 811 9751
rect 812 9747 816 9751
rect 817 9747 821 9751
rect 802 9737 806 9741
rect 807 9737 811 9741
rect 812 9737 816 9741
rect 817 9737 821 9741
rect 831 9757 835 9761
rect 836 9757 840 9761
rect 841 9757 845 9761
rect 846 9757 850 9761
rect 831 9747 835 9751
rect 836 9747 840 9751
rect 841 9747 845 9751
rect 846 9747 850 9751
rect 831 9737 835 9741
rect 836 9737 840 9741
rect 841 9737 845 9741
rect 846 9737 850 9741
rect 860 9757 864 9761
rect 865 9757 869 9761
rect 870 9757 874 9761
rect 875 9757 879 9761
rect 860 9747 864 9751
rect 865 9747 869 9751
rect 870 9747 874 9751
rect 875 9747 879 9751
rect 860 9737 864 9741
rect 865 9737 869 9741
rect 870 9737 874 9741
rect 875 9737 879 9741
rect 889 9757 893 9761
rect 894 9757 898 9761
rect 899 9757 903 9761
rect 904 9757 908 9761
rect 889 9747 893 9751
rect 894 9747 898 9751
rect 899 9747 903 9751
rect 904 9747 908 9751
rect 889 9737 893 9741
rect 894 9737 898 9741
rect 899 9737 903 9741
rect 904 9737 908 9741
rect 918 9757 922 9761
rect 923 9757 927 9761
rect 928 9757 932 9761
rect 933 9757 937 9761
rect 918 9747 922 9751
rect 923 9747 927 9751
rect 928 9747 932 9751
rect 933 9747 937 9751
rect 918 9737 922 9741
rect 923 9737 927 9741
rect 928 9737 932 9741
rect 933 9737 937 9741
rect 802 9711 806 9715
rect 807 9711 811 9715
rect 812 9711 816 9715
rect 817 9711 821 9715
rect 802 9701 806 9705
rect 807 9701 811 9705
rect 812 9701 816 9705
rect 817 9701 821 9705
rect 802 9691 806 9695
rect 807 9691 811 9695
rect 812 9691 816 9695
rect 817 9691 821 9695
rect 831 9711 835 9715
rect 836 9711 840 9715
rect 841 9711 845 9715
rect 846 9711 850 9715
rect 831 9701 835 9705
rect 836 9701 840 9705
rect 841 9701 845 9705
rect 846 9701 850 9705
rect 831 9691 835 9695
rect 836 9691 840 9695
rect 841 9691 845 9695
rect 846 9691 850 9695
rect 860 9711 864 9715
rect 865 9711 869 9715
rect 870 9711 874 9715
rect 875 9711 879 9715
rect 860 9701 864 9705
rect 865 9701 869 9705
rect 870 9701 874 9705
rect 875 9701 879 9705
rect 860 9691 864 9695
rect 865 9691 869 9695
rect 870 9691 874 9695
rect 875 9691 879 9695
rect 889 9711 893 9715
rect 894 9711 898 9715
rect 899 9711 903 9715
rect 904 9711 908 9715
rect 889 9701 893 9705
rect 894 9701 898 9705
rect 899 9701 903 9705
rect 904 9701 908 9705
rect 889 9691 893 9695
rect 894 9691 898 9695
rect 899 9691 903 9695
rect 904 9691 908 9695
rect 918 9711 922 9715
rect 923 9711 927 9715
rect 928 9711 932 9715
rect 933 9711 937 9715
rect 918 9701 922 9705
rect 923 9701 927 9705
rect 928 9701 932 9705
rect 933 9701 937 9705
rect 918 9691 922 9695
rect 923 9691 927 9695
rect 928 9691 932 9695
rect 933 9691 937 9695
rect 618 9618 622 9622
rect 628 9618 632 9622
rect 638 9618 642 9622
rect 618 9613 622 9617
rect 628 9613 632 9617
rect 638 9613 642 9617
rect 618 9608 622 9612
rect 628 9608 632 9612
rect 638 9608 642 9612
rect 618 9603 622 9607
rect 628 9603 632 9607
rect 638 9603 642 9607
rect 664 9618 668 9622
rect 674 9618 678 9622
rect 684 9618 688 9622
rect 664 9613 668 9617
rect 674 9613 678 9617
rect 684 9613 688 9617
rect 664 9608 668 9612
rect 674 9608 678 9612
rect 684 9608 688 9612
rect 1454 9992 1458 9996
rect 1461 9992 1465 9996
rect 1468 9992 1472 9996
rect 1475 9992 1479 9996
rect 1482 9992 1486 9996
rect 1489 9992 1493 9996
rect 1496 9992 1500 9996
rect 1503 9992 1507 9996
rect 1510 9992 1514 9996
rect 1517 9992 1521 9996
rect 1524 9992 1528 9996
rect 1531 9992 1535 9996
rect 1538 9992 1542 9996
rect 1763 9997 1767 10001
rect 1770 9997 1774 10001
rect 1777 9997 1781 10001
rect 1784 9997 1788 10001
rect 1791 9997 1795 10001
rect 1798 9997 1802 10001
rect 1805 9997 1809 10001
rect 1812 9997 1816 10001
rect 1819 9997 1823 10001
rect 1826 9997 1830 10001
rect 1833 9997 1837 10001
rect 1840 9997 1844 10001
rect 1847 9997 1851 10001
rect 1454 9987 1458 9991
rect 1461 9987 1465 9991
rect 1468 9987 1472 9991
rect 1475 9987 1479 9991
rect 1482 9987 1486 9991
rect 1489 9987 1493 9991
rect 1496 9987 1500 9991
rect 1503 9987 1507 9991
rect 1510 9987 1514 9991
rect 1517 9987 1521 9991
rect 1524 9987 1528 9991
rect 1531 9987 1535 9991
rect 1538 9987 1542 9991
rect 1454 9982 1458 9986
rect 1461 9982 1465 9986
rect 1468 9982 1472 9986
rect 1475 9982 1479 9986
rect 1482 9982 1486 9986
rect 1489 9982 1493 9986
rect 1496 9982 1500 9986
rect 1503 9982 1507 9986
rect 1510 9982 1514 9986
rect 1517 9982 1521 9986
rect 1524 9982 1528 9986
rect 1531 9982 1535 9986
rect 1538 9982 1542 9986
rect 1763 9992 1767 9996
rect 1770 9992 1774 9996
rect 1777 9992 1781 9996
rect 1784 9992 1788 9996
rect 1791 9992 1795 9996
rect 1798 9992 1802 9996
rect 1805 9992 1809 9996
rect 1812 9992 1816 9996
rect 1819 9992 1823 9996
rect 1826 9992 1830 9996
rect 1833 9992 1837 9996
rect 1840 9992 1844 9996
rect 1847 9992 1851 9996
rect 2072 9997 2076 10001
rect 2079 9997 2083 10001
rect 2086 9997 2090 10001
rect 2093 9997 2097 10001
rect 2100 9997 2104 10001
rect 2107 9997 2111 10001
rect 2114 9997 2118 10001
rect 2121 9997 2125 10001
rect 2128 9997 2132 10001
rect 2135 9997 2139 10001
rect 2142 9997 2146 10001
rect 2149 9997 2153 10001
rect 2156 9997 2160 10001
rect 1763 9987 1767 9991
rect 1770 9987 1774 9991
rect 1777 9987 1781 9991
rect 1784 9987 1788 9991
rect 1791 9987 1795 9991
rect 1798 9987 1802 9991
rect 1805 9987 1809 9991
rect 1812 9987 1816 9991
rect 1819 9987 1823 9991
rect 1826 9987 1830 9991
rect 1833 9987 1837 9991
rect 1840 9987 1844 9991
rect 1847 9987 1851 9991
rect 1763 9982 1767 9986
rect 1770 9982 1774 9986
rect 1777 9982 1781 9986
rect 1784 9982 1788 9986
rect 1791 9982 1795 9986
rect 1798 9982 1802 9986
rect 1805 9982 1809 9986
rect 1812 9982 1816 9986
rect 1819 9982 1823 9986
rect 1826 9982 1830 9986
rect 1833 9982 1837 9986
rect 1840 9982 1844 9986
rect 1847 9982 1851 9986
rect 2072 9992 2076 9996
rect 2079 9992 2083 9996
rect 2086 9992 2090 9996
rect 2093 9992 2097 9996
rect 2100 9992 2104 9996
rect 2107 9992 2111 9996
rect 2114 9992 2118 9996
rect 2121 9992 2125 9996
rect 2128 9992 2132 9996
rect 2135 9992 2139 9996
rect 2142 9992 2146 9996
rect 2149 9992 2153 9996
rect 2156 9992 2160 9996
rect 2381 9997 2385 10001
rect 2388 9997 2392 10001
rect 2395 9997 2399 10001
rect 2402 9997 2406 10001
rect 2409 9997 2413 10001
rect 2416 9997 2420 10001
rect 2423 9997 2427 10001
rect 2430 9997 2434 10001
rect 2437 9997 2441 10001
rect 2444 9997 2448 10001
rect 2451 9997 2455 10001
rect 2458 9997 2462 10001
rect 2465 9997 2469 10001
rect 2072 9987 2076 9991
rect 2079 9987 2083 9991
rect 2086 9987 2090 9991
rect 2093 9987 2097 9991
rect 2100 9987 2104 9991
rect 2107 9987 2111 9991
rect 2114 9987 2118 9991
rect 2121 9987 2125 9991
rect 2128 9987 2132 9991
rect 2135 9987 2139 9991
rect 2142 9987 2146 9991
rect 2149 9987 2153 9991
rect 2156 9987 2160 9991
rect 2072 9982 2076 9986
rect 2079 9982 2083 9986
rect 2086 9982 2090 9986
rect 2093 9982 2097 9986
rect 2100 9982 2104 9986
rect 2107 9982 2111 9986
rect 2114 9982 2118 9986
rect 2121 9982 2125 9986
rect 2128 9982 2132 9986
rect 2135 9982 2139 9986
rect 2142 9982 2146 9986
rect 2149 9982 2153 9986
rect 2156 9982 2160 9986
rect 2381 9992 2385 9996
rect 2388 9992 2392 9996
rect 2395 9992 2399 9996
rect 2402 9992 2406 9996
rect 2409 9992 2413 9996
rect 2416 9992 2420 9996
rect 2423 9992 2427 9996
rect 2430 9992 2434 9996
rect 2437 9992 2441 9996
rect 2444 9992 2448 9996
rect 2451 9992 2455 9996
rect 2458 9992 2462 9996
rect 2465 9992 2469 9996
rect 2690 9997 2694 10001
rect 2697 9997 2701 10001
rect 2704 9997 2708 10001
rect 2711 9997 2715 10001
rect 2718 9997 2722 10001
rect 2725 9997 2729 10001
rect 2732 9997 2736 10001
rect 2739 9997 2743 10001
rect 2746 9997 2750 10001
rect 2753 9997 2757 10001
rect 2760 9997 2764 10001
rect 2767 9997 2771 10001
rect 2774 9997 2778 10001
rect 2381 9987 2385 9991
rect 2388 9987 2392 9991
rect 2395 9987 2399 9991
rect 2402 9987 2406 9991
rect 2409 9987 2413 9991
rect 2416 9987 2420 9991
rect 2423 9987 2427 9991
rect 2430 9987 2434 9991
rect 2437 9987 2441 9991
rect 2444 9987 2448 9991
rect 2451 9987 2455 9991
rect 2458 9987 2462 9991
rect 2465 9987 2469 9991
rect 2381 9982 2385 9986
rect 2388 9982 2392 9986
rect 2395 9982 2399 9986
rect 2402 9982 2406 9986
rect 2409 9982 2413 9986
rect 2416 9982 2420 9986
rect 2423 9982 2427 9986
rect 2430 9982 2434 9986
rect 2437 9982 2441 9986
rect 2444 9982 2448 9986
rect 2451 9982 2455 9986
rect 2458 9982 2462 9986
rect 2465 9982 2469 9986
rect 2690 9992 2694 9996
rect 2697 9992 2701 9996
rect 2704 9992 2708 9996
rect 2711 9992 2715 9996
rect 2718 9992 2722 9996
rect 2725 9992 2729 9996
rect 2732 9992 2736 9996
rect 2739 9992 2743 9996
rect 2746 9992 2750 9996
rect 2753 9992 2757 9996
rect 2760 9992 2764 9996
rect 2767 9992 2771 9996
rect 2774 9992 2778 9996
rect 2999 9997 3003 10001
rect 3006 9997 3010 10001
rect 3013 9997 3017 10001
rect 3020 9997 3024 10001
rect 3027 9997 3031 10001
rect 3034 9997 3038 10001
rect 3041 9997 3045 10001
rect 3048 9997 3052 10001
rect 3055 9997 3059 10001
rect 3062 9997 3066 10001
rect 3069 9997 3073 10001
rect 3076 9997 3080 10001
rect 3083 9997 3087 10001
rect 2690 9987 2694 9991
rect 2697 9987 2701 9991
rect 2704 9987 2708 9991
rect 2711 9987 2715 9991
rect 2718 9987 2722 9991
rect 2725 9987 2729 9991
rect 2732 9987 2736 9991
rect 2739 9987 2743 9991
rect 2746 9987 2750 9991
rect 2753 9987 2757 9991
rect 2760 9987 2764 9991
rect 2767 9987 2771 9991
rect 2774 9987 2778 9991
rect 2690 9982 2694 9986
rect 2697 9982 2701 9986
rect 2704 9982 2708 9986
rect 2711 9982 2715 9986
rect 2718 9982 2722 9986
rect 2725 9982 2729 9986
rect 2732 9982 2736 9986
rect 2739 9982 2743 9986
rect 2746 9982 2750 9986
rect 2753 9982 2757 9986
rect 2760 9982 2764 9986
rect 2767 9982 2771 9986
rect 2774 9982 2778 9986
rect 2999 9992 3003 9996
rect 3006 9992 3010 9996
rect 3013 9992 3017 9996
rect 3020 9992 3024 9996
rect 3027 9992 3031 9996
rect 3034 9992 3038 9996
rect 3041 9992 3045 9996
rect 3048 9992 3052 9996
rect 3055 9992 3059 9996
rect 3062 9992 3066 9996
rect 3069 9992 3073 9996
rect 3076 9992 3080 9996
rect 3083 9992 3087 9996
rect 3308 9997 3312 10001
rect 3315 9997 3319 10001
rect 3322 9997 3326 10001
rect 3329 9997 3333 10001
rect 3336 9997 3340 10001
rect 3343 9997 3347 10001
rect 3350 9997 3354 10001
rect 3357 9997 3361 10001
rect 3364 9997 3368 10001
rect 3371 9997 3375 10001
rect 3378 9997 3382 10001
rect 3385 9997 3389 10001
rect 3392 9997 3396 10001
rect 2999 9987 3003 9991
rect 3006 9987 3010 9991
rect 3013 9987 3017 9991
rect 3020 9987 3024 9991
rect 3027 9987 3031 9991
rect 3034 9987 3038 9991
rect 3041 9987 3045 9991
rect 3048 9987 3052 9991
rect 3055 9987 3059 9991
rect 3062 9987 3066 9991
rect 3069 9987 3073 9991
rect 3076 9987 3080 9991
rect 3083 9987 3087 9991
rect 2999 9982 3003 9986
rect 3006 9982 3010 9986
rect 3013 9982 3017 9986
rect 3020 9982 3024 9986
rect 3027 9982 3031 9986
rect 3034 9982 3038 9986
rect 3041 9982 3045 9986
rect 3048 9982 3052 9986
rect 3055 9982 3059 9986
rect 3062 9982 3066 9986
rect 3069 9982 3073 9986
rect 3076 9982 3080 9986
rect 3083 9982 3087 9986
rect 3308 9992 3312 9996
rect 3315 9992 3319 9996
rect 3322 9992 3326 9996
rect 3329 9992 3333 9996
rect 3336 9992 3340 9996
rect 3343 9992 3347 9996
rect 3350 9992 3354 9996
rect 3357 9992 3361 9996
rect 3364 9992 3368 9996
rect 3371 9992 3375 9996
rect 3378 9992 3382 9996
rect 3385 9992 3389 9996
rect 3392 9992 3396 9996
rect 3617 9997 3621 10001
rect 3624 9997 3628 10001
rect 3631 9997 3635 10001
rect 3638 9997 3642 10001
rect 3645 9997 3649 10001
rect 3652 9997 3656 10001
rect 3659 9997 3663 10001
rect 3666 9997 3670 10001
rect 3673 9997 3677 10001
rect 3680 9997 3684 10001
rect 3687 9997 3691 10001
rect 3694 9997 3698 10001
rect 3701 9997 3705 10001
rect 3308 9987 3312 9991
rect 3315 9987 3319 9991
rect 3322 9987 3326 9991
rect 3329 9987 3333 9991
rect 3336 9987 3340 9991
rect 3343 9987 3347 9991
rect 3350 9987 3354 9991
rect 3357 9987 3361 9991
rect 3364 9987 3368 9991
rect 3371 9987 3375 9991
rect 3378 9987 3382 9991
rect 3385 9987 3389 9991
rect 3392 9987 3396 9991
rect 3308 9982 3312 9986
rect 3315 9982 3319 9986
rect 3322 9982 3326 9986
rect 3329 9982 3333 9986
rect 3336 9982 3340 9986
rect 3343 9982 3347 9986
rect 3350 9982 3354 9986
rect 3357 9982 3361 9986
rect 3364 9982 3368 9986
rect 3371 9982 3375 9986
rect 3378 9982 3382 9986
rect 3385 9982 3389 9986
rect 3392 9982 3396 9986
rect 3617 9992 3621 9996
rect 3624 9992 3628 9996
rect 3631 9992 3635 9996
rect 3638 9992 3642 9996
rect 3645 9992 3649 9996
rect 3652 9992 3656 9996
rect 3659 9992 3663 9996
rect 3666 9992 3670 9996
rect 3673 9992 3677 9996
rect 3680 9992 3684 9996
rect 3687 9992 3691 9996
rect 3694 9992 3698 9996
rect 3701 9992 3705 9996
rect 3926 9997 3930 10001
rect 3933 9997 3937 10001
rect 3940 9997 3944 10001
rect 3947 9997 3951 10001
rect 3954 9997 3958 10001
rect 3961 9997 3965 10001
rect 3968 9997 3972 10001
rect 3975 9997 3979 10001
rect 3982 9997 3986 10001
rect 3989 9997 3993 10001
rect 3996 9997 4000 10001
rect 4003 9997 4007 10001
rect 4010 9997 4014 10001
rect 3617 9987 3621 9991
rect 3624 9987 3628 9991
rect 3631 9987 3635 9991
rect 3638 9987 3642 9991
rect 3645 9987 3649 9991
rect 3652 9987 3656 9991
rect 3659 9987 3663 9991
rect 3666 9987 3670 9991
rect 3673 9987 3677 9991
rect 3680 9987 3684 9991
rect 3687 9987 3691 9991
rect 3694 9987 3698 9991
rect 3701 9987 3705 9991
rect 3617 9982 3621 9986
rect 3624 9982 3628 9986
rect 3631 9982 3635 9986
rect 3638 9982 3642 9986
rect 3645 9982 3649 9986
rect 3652 9982 3656 9986
rect 3659 9982 3663 9986
rect 3666 9982 3670 9986
rect 3673 9982 3677 9986
rect 3680 9982 3684 9986
rect 3687 9982 3691 9986
rect 3694 9982 3698 9986
rect 3701 9982 3705 9986
rect 3926 9992 3930 9996
rect 3933 9992 3937 9996
rect 3940 9992 3944 9996
rect 3947 9992 3951 9996
rect 3954 9992 3958 9996
rect 3961 9992 3965 9996
rect 3968 9992 3972 9996
rect 3975 9992 3979 9996
rect 3982 9992 3986 9996
rect 3989 9992 3993 9996
rect 3996 9992 4000 9996
rect 4003 9992 4007 9996
rect 4010 9992 4014 9996
rect 3926 9987 3930 9991
rect 3933 9987 3937 9991
rect 3940 9987 3944 9991
rect 3947 9987 3951 9991
rect 3954 9987 3958 9991
rect 3961 9987 3965 9991
rect 3968 9987 3972 9991
rect 3975 9987 3979 9991
rect 3982 9987 3986 9991
rect 3989 9987 3993 9991
rect 3996 9987 4000 9991
rect 4003 9987 4007 9991
rect 4010 9987 4014 9991
rect 3926 9982 3930 9986
rect 3933 9982 3937 9986
rect 3940 9982 3944 9986
rect 3947 9982 3951 9986
rect 3954 9982 3958 9986
rect 3961 9982 3965 9986
rect 3968 9982 3972 9986
rect 3975 9982 3979 9986
rect 3982 9982 3986 9986
rect 3989 9982 3993 9986
rect 3996 9982 4000 9986
rect 4003 9982 4007 9986
rect 4010 9982 4014 9986
rect 1397 9949 1401 9953
rect 1407 9949 1411 9953
rect 1417 9949 1421 9953
rect 1427 9949 1431 9953
rect 1437 9949 1441 9953
rect 1402 9944 1406 9948
rect 1412 9944 1416 9948
rect 1422 9944 1426 9948
rect 1432 9944 1436 9948
rect 1397 9939 1401 9943
rect 1407 9939 1411 9943
rect 1417 9939 1421 9943
rect 1427 9939 1431 9943
rect 1437 9939 1441 9943
rect 1402 9934 1406 9938
rect 1412 9934 1416 9938
rect 1422 9934 1426 9938
rect 1432 9934 1436 9938
rect 1397 9929 1401 9933
rect 1407 9929 1411 9933
rect 1417 9929 1421 9933
rect 1427 9929 1431 9933
rect 1437 9929 1441 9933
rect 1402 9924 1406 9928
rect 1412 9924 1416 9928
rect 1422 9924 1426 9928
rect 1432 9924 1436 9928
rect 1397 9919 1401 9923
rect 1407 9919 1411 9923
rect 1417 9919 1421 9923
rect 1427 9919 1431 9923
rect 1437 9919 1441 9923
rect 1402 9914 1406 9918
rect 1412 9914 1416 9918
rect 1422 9914 1426 9918
rect 1432 9914 1436 9918
rect 1397 9909 1401 9913
rect 1407 9909 1411 9913
rect 1417 9909 1421 9913
rect 1427 9909 1431 9913
rect 1437 9909 1441 9913
rect 1402 9904 1406 9908
rect 1412 9904 1416 9908
rect 1422 9904 1426 9908
rect 1432 9904 1436 9908
rect 1397 9899 1401 9903
rect 1407 9899 1411 9903
rect 1417 9899 1421 9903
rect 1427 9899 1431 9903
rect 1437 9899 1441 9903
rect 1402 9894 1406 9898
rect 1412 9894 1416 9898
rect 1422 9894 1426 9898
rect 1432 9894 1436 9898
rect 1397 9889 1401 9893
rect 1407 9889 1411 9893
rect 1417 9889 1421 9893
rect 1427 9889 1431 9893
rect 1437 9889 1441 9893
rect 1402 9884 1406 9888
rect 1412 9884 1416 9888
rect 1422 9884 1426 9888
rect 1432 9884 1436 9888
rect 1397 9879 1401 9883
rect 1407 9879 1411 9883
rect 1417 9879 1421 9883
rect 1427 9879 1431 9883
rect 1437 9879 1441 9883
rect 1402 9874 1406 9878
rect 1412 9874 1416 9878
rect 1422 9874 1426 9878
rect 1432 9874 1436 9878
rect 1397 9869 1401 9873
rect 1407 9869 1411 9873
rect 1417 9869 1421 9873
rect 1427 9869 1431 9873
rect 1437 9869 1441 9873
rect 1402 9864 1406 9868
rect 1412 9864 1416 9868
rect 1422 9864 1426 9868
rect 1432 9864 1436 9868
rect 1385 9848 1389 9852
rect 1392 9848 1396 9852
rect 1397 9848 1401 9852
rect 1402 9848 1406 9852
rect 1407 9848 1411 9852
rect 1412 9848 1416 9852
rect 1417 9848 1421 9852
rect 1422 9848 1426 9852
rect 1427 9848 1431 9852
rect 1432 9848 1436 9852
rect 1437 9848 1441 9852
rect 1442 9848 1446 9852
rect 1449 9848 1453 9852
rect 1364 9796 1368 9800
rect 1369 9796 1373 9800
rect 1364 9791 1368 9795
rect 1369 9791 1373 9795
rect 1364 9786 1368 9790
rect 1369 9786 1373 9790
rect 1364 9781 1368 9785
rect 1369 9781 1373 9785
rect 1364 9776 1368 9780
rect 1369 9776 1373 9780
rect 1364 9771 1368 9775
rect 1369 9771 1373 9775
rect 1364 9766 1368 9770
rect 1369 9766 1373 9770
rect 1319 9757 1323 9761
rect 1324 9757 1328 9761
rect 1329 9757 1333 9761
rect 1334 9757 1338 9761
rect 1319 9747 1323 9751
rect 1324 9747 1328 9751
rect 1329 9747 1333 9751
rect 1334 9747 1338 9751
rect 1319 9737 1323 9741
rect 1324 9737 1328 9741
rect 1329 9737 1333 9741
rect 1334 9737 1338 9741
rect 1364 9761 1368 9765
rect 1369 9761 1373 9765
rect 1364 9756 1368 9760
rect 1369 9756 1373 9760
rect 1364 9751 1368 9755
rect 1369 9751 1373 9755
rect 1364 9746 1368 9750
rect 1369 9746 1373 9750
rect 1364 9741 1368 9745
rect 1369 9741 1373 9745
rect 1364 9736 1368 9740
rect 1369 9736 1373 9740
rect 1319 9711 1323 9715
rect 1324 9711 1328 9715
rect 1329 9711 1333 9715
rect 1334 9711 1338 9715
rect 1319 9701 1323 9705
rect 1324 9701 1328 9705
rect 1329 9701 1333 9705
rect 1334 9701 1338 9705
rect 1319 9691 1323 9695
rect 1324 9691 1328 9695
rect 1329 9691 1333 9695
rect 1334 9691 1338 9695
rect 1557 9949 1561 9953
rect 1567 9949 1571 9953
rect 1577 9949 1581 9953
rect 1587 9949 1591 9953
rect 1597 9949 1601 9953
rect 1562 9944 1566 9948
rect 1572 9944 1576 9948
rect 1582 9944 1586 9948
rect 1592 9944 1596 9948
rect 1557 9939 1561 9943
rect 1567 9939 1571 9943
rect 1577 9939 1581 9943
rect 1587 9939 1591 9943
rect 1597 9939 1601 9943
rect 1562 9934 1566 9938
rect 1572 9934 1576 9938
rect 1582 9934 1586 9938
rect 1592 9934 1596 9938
rect 1557 9929 1561 9933
rect 1567 9929 1571 9933
rect 1577 9929 1581 9933
rect 1587 9929 1591 9933
rect 1597 9929 1601 9933
rect 1562 9924 1566 9928
rect 1572 9924 1576 9928
rect 1582 9924 1586 9928
rect 1592 9924 1596 9928
rect 1557 9919 1561 9923
rect 1567 9919 1571 9923
rect 1577 9919 1581 9923
rect 1587 9919 1591 9923
rect 1597 9919 1601 9923
rect 1562 9914 1566 9918
rect 1572 9914 1576 9918
rect 1582 9914 1586 9918
rect 1592 9914 1596 9918
rect 1557 9909 1561 9913
rect 1567 9909 1571 9913
rect 1577 9909 1581 9913
rect 1587 9909 1591 9913
rect 1597 9909 1601 9913
rect 1562 9904 1566 9908
rect 1572 9904 1576 9908
rect 1582 9904 1586 9908
rect 1592 9904 1596 9908
rect 1557 9899 1561 9903
rect 1567 9899 1571 9903
rect 1577 9899 1581 9903
rect 1587 9899 1591 9903
rect 1597 9899 1601 9903
rect 1562 9894 1566 9898
rect 1572 9894 1576 9898
rect 1582 9894 1586 9898
rect 1592 9894 1596 9898
rect 1557 9889 1561 9893
rect 1567 9889 1571 9893
rect 1577 9889 1581 9893
rect 1587 9889 1591 9893
rect 1597 9889 1601 9893
rect 1562 9884 1566 9888
rect 1572 9884 1576 9888
rect 1582 9884 1586 9888
rect 1592 9884 1596 9888
rect 1557 9879 1561 9883
rect 1567 9879 1571 9883
rect 1577 9879 1581 9883
rect 1587 9879 1591 9883
rect 1597 9879 1601 9883
rect 1562 9874 1566 9878
rect 1572 9874 1576 9878
rect 1582 9874 1586 9878
rect 1592 9874 1596 9878
rect 1557 9869 1561 9873
rect 1567 9869 1571 9873
rect 1577 9869 1581 9873
rect 1587 9869 1591 9873
rect 1597 9869 1601 9873
rect 1562 9864 1566 9868
rect 1572 9864 1576 9868
rect 1582 9864 1586 9868
rect 1592 9864 1596 9868
rect 1545 9848 1549 9852
rect 1552 9848 1556 9852
rect 1557 9848 1561 9852
rect 1562 9848 1566 9852
rect 1567 9848 1571 9852
rect 1572 9848 1576 9852
rect 1577 9848 1581 9852
rect 1582 9848 1586 9852
rect 1587 9848 1591 9852
rect 1592 9848 1596 9852
rect 1597 9848 1601 9852
rect 1602 9848 1606 9852
rect 1609 9848 1613 9852
rect 1706 9949 1710 9953
rect 1716 9949 1720 9953
rect 1726 9949 1730 9953
rect 1736 9949 1740 9953
rect 1746 9949 1750 9953
rect 1711 9944 1715 9948
rect 1721 9944 1725 9948
rect 1731 9944 1735 9948
rect 1741 9944 1745 9948
rect 1706 9939 1710 9943
rect 1716 9939 1720 9943
rect 1726 9939 1730 9943
rect 1736 9939 1740 9943
rect 1746 9939 1750 9943
rect 1711 9934 1715 9938
rect 1721 9934 1725 9938
rect 1731 9934 1735 9938
rect 1741 9934 1745 9938
rect 1706 9929 1710 9933
rect 1716 9929 1720 9933
rect 1726 9929 1730 9933
rect 1736 9929 1740 9933
rect 1746 9929 1750 9933
rect 1711 9924 1715 9928
rect 1721 9924 1725 9928
rect 1731 9924 1735 9928
rect 1741 9924 1745 9928
rect 1706 9919 1710 9923
rect 1716 9919 1720 9923
rect 1726 9919 1730 9923
rect 1736 9919 1740 9923
rect 1746 9919 1750 9923
rect 1711 9914 1715 9918
rect 1721 9914 1725 9918
rect 1731 9914 1735 9918
rect 1741 9914 1745 9918
rect 1706 9909 1710 9913
rect 1716 9909 1720 9913
rect 1726 9909 1730 9913
rect 1736 9909 1740 9913
rect 1746 9909 1750 9913
rect 1711 9904 1715 9908
rect 1721 9904 1725 9908
rect 1731 9904 1735 9908
rect 1741 9904 1745 9908
rect 1706 9899 1710 9903
rect 1716 9899 1720 9903
rect 1726 9899 1730 9903
rect 1736 9899 1740 9903
rect 1746 9899 1750 9903
rect 1711 9894 1715 9898
rect 1721 9894 1725 9898
rect 1731 9894 1735 9898
rect 1741 9894 1745 9898
rect 1706 9889 1710 9893
rect 1716 9889 1720 9893
rect 1726 9889 1730 9893
rect 1736 9889 1740 9893
rect 1746 9889 1750 9893
rect 1711 9884 1715 9888
rect 1721 9884 1725 9888
rect 1731 9884 1735 9888
rect 1741 9884 1745 9888
rect 1706 9879 1710 9883
rect 1716 9879 1720 9883
rect 1726 9879 1730 9883
rect 1736 9879 1740 9883
rect 1746 9879 1750 9883
rect 1711 9874 1715 9878
rect 1721 9874 1725 9878
rect 1731 9874 1735 9878
rect 1741 9874 1745 9878
rect 1706 9869 1710 9873
rect 1716 9869 1720 9873
rect 1726 9869 1730 9873
rect 1736 9869 1740 9873
rect 1746 9869 1750 9873
rect 1711 9864 1715 9868
rect 1721 9864 1725 9868
rect 1731 9864 1735 9868
rect 1741 9864 1745 9868
rect 1694 9848 1698 9852
rect 1701 9848 1705 9852
rect 1706 9848 1710 9852
rect 1711 9848 1715 9852
rect 1716 9848 1720 9852
rect 1721 9848 1725 9852
rect 1726 9848 1730 9852
rect 1731 9848 1735 9852
rect 1736 9848 1740 9852
rect 1741 9848 1745 9852
rect 1746 9848 1750 9852
rect 1751 9848 1755 9852
rect 1758 9848 1762 9852
rect 1866 9949 1870 9953
rect 1876 9949 1880 9953
rect 1886 9949 1890 9953
rect 1896 9949 1900 9953
rect 1906 9949 1910 9953
rect 1871 9944 1875 9948
rect 1881 9944 1885 9948
rect 1891 9944 1895 9948
rect 1901 9944 1905 9948
rect 1866 9939 1870 9943
rect 1876 9939 1880 9943
rect 1886 9939 1890 9943
rect 1896 9939 1900 9943
rect 1906 9939 1910 9943
rect 1871 9934 1875 9938
rect 1881 9934 1885 9938
rect 1891 9934 1895 9938
rect 1901 9934 1905 9938
rect 1866 9929 1870 9933
rect 1876 9929 1880 9933
rect 1886 9929 1890 9933
rect 1896 9929 1900 9933
rect 1906 9929 1910 9933
rect 1871 9924 1875 9928
rect 1881 9924 1885 9928
rect 1891 9924 1895 9928
rect 1901 9924 1905 9928
rect 1866 9919 1870 9923
rect 1876 9919 1880 9923
rect 1886 9919 1890 9923
rect 1896 9919 1900 9923
rect 1906 9919 1910 9923
rect 1871 9914 1875 9918
rect 1881 9914 1885 9918
rect 1891 9914 1895 9918
rect 1901 9914 1905 9918
rect 1866 9909 1870 9913
rect 1876 9909 1880 9913
rect 1886 9909 1890 9913
rect 1896 9909 1900 9913
rect 1906 9909 1910 9913
rect 1871 9904 1875 9908
rect 1881 9904 1885 9908
rect 1891 9904 1895 9908
rect 1901 9904 1905 9908
rect 1866 9899 1870 9903
rect 1876 9899 1880 9903
rect 1886 9899 1890 9903
rect 1896 9899 1900 9903
rect 1906 9899 1910 9903
rect 1871 9894 1875 9898
rect 1881 9894 1885 9898
rect 1891 9894 1895 9898
rect 1901 9894 1905 9898
rect 1866 9889 1870 9893
rect 1876 9889 1880 9893
rect 1886 9889 1890 9893
rect 1896 9889 1900 9893
rect 1906 9889 1910 9893
rect 1871 9884 1875 9888
rect 1881 9884 1885 9888
rect 1891 9884 1895 9888
rect 1901 9884 1905 9888
rect 1866 9879 1870 9883
rect 1876 9879 1880 9883
rect 1886 9879 1890 9883
rect 1896 9879 1900 9883
rect 1906 9879 1910 9883
rect 1871 9874 1875 9878
rect 1881 9874 1885 9878
rect 1891 9874 1895 9878
rect 1901 9874 1905 9878
rect 1866 9869 1870 9873
rect 1876 9869 1880 9873
rect 1886 9869 1890 9873
rect 1896 9869 1900 9873
rect 1906 9869 1910 9873
rect 1871 9864 1875 9868
rect 1881 9864 1885 9868
rect 1891 9864 1895 9868
rect 1901 9864 1905 9868
rect 1854 9848 1858 9852
rect 1861 9848 1865 9852
rect 1866 9848 1870 9852
rect 1871 9848 1875 9852
rect 1876 9848 1880 9852
rect 1881 9848 1885 9852
rect 1886 9848 1890 9852
rect 1891 9848 1895 9852
rect 1896 9848 1900 9852
rect 1901 9848 1905 9852
rect 1906 9848 1910 9852
rect 1911 9848 1915 9852
rect 1918 9848 1922 9852
rect 1499 9711 1503 9715
rect 1504 9711 1508 9715
rect 2015 9949 2019 9953
rect 2025 9949 2029 9953
rect 2035 9949 2039 9953
rect 2045 9949 2049 9953
rect 2055 9949 2059 9953
rect 2020 9944 2024 9948
rect 2030 9944 2034 9948
rect 2040 9944 2044 9948
rect 2050 9944 2054 9948
rect 2015 9939 2019 9943
rect 2025 9939 2029 9943
rect 2035 9939 2039 9943
rect 2045 9939 2049 9943
rect 2055 9939 2059 9943
rect 2020 9934 2024 9938
rect 2030 9934 2034 9938
rect 2040 9934 2044 9938
rect 2050 9934 2054 9938
rect 2015 9929 2019 9933
rect 2025 9929 2029 9933
rect 2035 9929 2039 9933
rect 2045 9929 2049 9933
rect 2055 9929 2059 9933
rect 2020 9924 2024 9928
rect 2030 9924 2034 9928
rect 2040 9924 2044 9928
rect 2050 9924 2054 9928
rect 2015 9919 2019 9923
rect 2025 9919 2029 9923
rect 2035 9919 2039 9923
rect 2045 9919 2049 9923
rect 2055 9919 2059 9923
rect 2020 9914 2024 9918
rect 2030 9914 2034 9918
rect 2040 9914 2044 9918
rect 2050 9914 2054 9918
rect 2015 9909 2019 9913
rect 2025 9909 2029 9913
rect 2035 9909 2039 9913
rect 2045 9909 2049 9913
rect 2055 9909 2059 9913
rect 2020 9904 2024 9908
rect 2030 9904 2034 9908
rect 2040 9904 2044 9908
rect 2050 9904 2054 9908
rect 2015 9899 2019 9903
rect 2025 9899 2029 9903
rect 2035 9899 2039 9903
rect 2045 9899 2049 9903
rect 2055 9899 2059 9903
rect 2020 9894 2024 9898
rect 2030 9894 2034 9898
rect 2040 9894 2044 9898
rect 2050 9894 2054 9898
rect 2015 9889 2019 9893
rect 2025 9889 2029 9893
rect 2035 9889 2039 9893
rect 2045 9889 2049 9893
rect 2055 9889 2059 9893
rect 2020 9884 2024 9888
rect 2030 9884 2034 9888
rect 2040 9884 2044 9888
rect 2050 9884 2054 9888
rect 2015 9879 2019 9883
rect 2025 9879 2029 9883
rect 2035 9879 2039 9883
rect 2045 9879 2049 9883
rect 2055 9879 2059 9883
rect 2020 9874 2024 9878
rect 2030 9874 2034 9878
rect 2040 9874 2044 9878
rect 2050 9874 2054 9878
rect 2015 9869 2019 9873
rect 2025 9869 2029 9873
rect 2035 9869 2039 9873
rect 2045 9869 2049 9873
rect 2055 9869 2059 9873
rect 2020 9864 2024 9868
rect 2030 9864 2034 9868
rect 2040 9864 2044 9868
rect 2050 9864 2054 9868
rect 2003 9848 2007 9852
rect 2010 9848 2014 9852
rect 2015 9848 2019 9852
rect 2020 9848 2024 9852
rect 2025 9848 2029 9852
rect 2030 9848 2034 9852
rect 2035 9848 2039 9852
rect 2040 9848 2044 9852
rect 2045 9848 2049 9852
rect 2050 9848 2054 9852
rect 2055 9848 2059 9852
rect 2060 9848 2064 9852
rect 2067 9848 2071 9852
rect 2175 9949 2179 9953
rect 2185 9949 2189 9953
rect 2195 9949 2199 9953
rect 2205 9949 2209 9953
rect 2215 9949 2219 9953
rect 2180 9944 2184 9948
rect 2190 9944 2194 9948
rect 2200 9944 2204 9948
rect 2210 9944 2214 9948
rect 2175 9939 2179 9943
rect 2185 9939 2189 9943
rect 2195 9939 2199 9943
rect 2205 9939 2209 9943
rect 2215 9939 2219 9943
rect 2180 9934 2184 9938
rect 2190 9934 2194 9938
rect 2200 9934 2204 9938
rect 2210 9934 2214 9938
rect 2175 9929 2179 9933
rect 2185 9929 2189 9933
rect 2195 9929 2199 9933
rect 2205 9929 2209 9933
rect 2215 9929 2219 9933
rect 2180 9924 2184 9928
rect 2190 9924 2194 9928
rect 2200 9924 2204 9928
rect 2210 9924 2214 9928
rect 2175 9919 2179 9923
rect 2185 9919 2189 9923
rect 2195 9919 2199 9923
rect 2205 9919 2209 9923
rect 2215 9919 2219 9923
rect 2180 9914 2184 9918
rect 2190 9914 2194 9918
rect 2200 9914 2204 9918
rect 2210 9914 2214 9918
rect 2175 9909 2179 9913
rect 2185 9909 2189 9913
rect 2195 9909 2199 9913
rect 2205 9909 2209 9913
rect 2215 9909 2219 9913
rect 2180 9904 2184 9908
rect 2190 9904 2194 9908
rect 2200 9904 2204 9908
rect 2210 9904 2214 9908
rect 2175 9899 2179 9903
rect 2185 9899 2189 9903
rect 2195 9899 2199 9903
rect 2205 9899 2209 9903
rect 2215 9899 2219 9903
rect 2180 9894 2184 9898
rect 2190 9894 2194 9898
rect 2200 9894 2204 9898
rect 2210 9894 2214 9898
rect 2175 9889 2179 9893
rect 2185 9889 2189 9893
rect 2195 9889 2199 9893
rect 2205 9889 2209 9893
rect 2215 9889 2219 9893
rect 2180 9884 2184 9888
rect 2190 9884 2194 9888
rect 2200 9884 2204 9888
rect 2210 9884 2214 9888
rect 2175 9879 2179 9883
rect 2185 9879 2189 9883
rect 2195 9879 2199 9883
rect 2205 9879 2209 9883
rect 2215 9879 2219 9883
rect 2180 9874 2184 9878
rect 2190 9874 2194 9878
rect 2200 9874 2204 9878
rect 2210 9874 2214 9878
rect 2175 9869 2179 9873
rect 2185 9869 2189 9873
rect 2195 9869 2199 9873
rect 2205 9869 2209 9873
rect 2215 9869 2219 9873
rect 2180 9864 2184 9868
rect 2190 9864 2194 9868
rect 2200 9864 2204 9868
rect 2210 9864 2214 9868
rect 2163 9848 2167 9852
rect 2170 9848 2174 9852
rect 2175 9848 2179 9852
rect 2180 9848 2184 9852
rect 2185 9848 2189 9852
rect 2190 9848 2194 9852
rect 2195 9848 2199 9852
rect 2200 9848 2204 9852
rect 2205 9848 2209 9852
rect 2210 9848 2214 9852
rect 2215 9848 2219 9852
rect 2220 9848 2224 9852
rect 2227 9848 2231 9852
rect 1778 9827 1782 9831
rect 1836 9827 1840 9831
rect 1778 9811 1782 9815
rect 1836 9811 1840 9815
rect 1673 9796 1677 9800
rect 1678 9796 1682 9800
rect 1778 9795 1782 9799
rect 1673 9791 1677 9795
rect 1678 9791 1682 9795
rect 2324 9949 2328 9953
rect 2334 9949 2338 9953
rect 2344 9949 2348 9953
rect 2354 9949 2358 9953
rect 2364 9949 2368 9953
rect 2329 9944 2333 9948
rect 2339 9944 2343 9948
rect 2349 9944 2353 9948
rect 2359 9944 2363 9948
rect 2324 9939 2328 9943
rect 2334 9939 2338 9943
rect 2344 9939 2348 9943
rect 2354 9939 2358 9943
rect 2364 9939 2368 9943
rect 2329 9934 2333 9938
rect 2339 9934 2343 9938
rect 2349 9934 2353 9938
rect 2359 9934 2363 9938
rect 2324 9929 2328 9933
rect 2334 9929 2338 9933
rect 2344 9929 2348 9933
rect 2354 9929 2358 9933
rect 2364 9929 2368 9933
rect 2329 9924 2333 9928
rect 2339 9924 2343 9928
rect 2349 9924 2353 9928
rect 2359 9924 2363 9928
rect 2324 9919 2328 9923
rect 2334 9919 2338 9923
rect 2344 9919 2348 9923
rect 2354 9919 2358 9923
rect 2364 9919 2368 9923
rect 2329 9914 2333 9918
rect 2339 9914 2343 9918
rect 2349 9914 2353 9918
rect 2359 9914 2363 9918
rect 2324 9909 2328 9913
rect 2334 9909 2338 9913
rect 2344 9909 2348 9913
rect 2354 9909 2358 9913
rect 2364 9909 2368 9913
rect 2329 9904 2333 9908
rect 2339 9904 2343 9908
rect 2349 9904 2353 9908
rect 2359 9904 2363 9908
rect 2324 9899 2328 9903
rect 2334 9899 2338 9903
rect 2344 9899 2348 9903
rect 2354 9899 2358 9903
rect 2364 9899 2368 9903
rect 2329 9894 2333 9898
rect 2339 9894 2343 9898
rect 2349 9894 2353 9898
rect 2359 9894 2363 9898
rect 2324 9889 2328 9893
rect 2334 9889 2338 9893
rect 2344 9889 2348 9893
rect 2354 9889 2358 9893
rect 2364 9889 2368 9893
rect 2329 9884 2333 9888
rect 2339 9884 2343 9888
rect 2349 9884 2353 9888
rect 2359 9884 2363 9888
rect 2324 9879 2328 9883
rect 2334 9879 2338 9883
rect 2344 9879 2348 9883
rect 2354 9879 2358 9883
rect 2364 9879 2368 9883
rect 2329 9874 2333 9878
rect 2339 9874 2343 9878
rect 2349 9874 2353 9878
rect 2359 9874 2363 9878
rect 2324 9869 2328 9873
rect 2334 9869 2338 9873
rect 2344 9869 2348 9873
rect 2354 9869 2358 9873
rect 2364 9869 2368 9873
rect 2329 9864 2333 9868
rect 2339 9864 2343 9868
rect 2349 9864 2353 9868
rect 2359 9864 2363 9868
rect 2312 9848 2316 9852
rect 2319 9848 2323 9852
rect 2324 9848 2328 9852
rect 2329 9848 2333 9852
rect 2334 9848 2338 9852
rect 2339 9848 2343 9852
rect 2344 9848 2348 9852
rect 2349 9848 2353 9852
rect 2354 9848 2358 9852
rect 2359 9848 2363 9852
rect 2364 9848 2368 9852
rect 2369 9848 2373 9852
rect 2376 9848 2380 9852
rect 2484 9949 2488 9953
rect 2494 9949 2498 9953
rect 2504 9949 2508 9953
rect 2514 9949 2518 9953
rect 2524 9949 2528 9953
rect 2489 9944 2493 9948
rect 2499 9944 2503 9948
rect 2509 9944 2513 9948
rect 2519 9944 2523 9948
rect 2484 9939 2488 9943
rect 2494 9939 2498 9943
rect 2504 9939 2508 9943
rect 2514 9939 2518 9943
rect 2524 9939 2528 9943
rect 2489 9934 2493 9938
rect 2499 9934 2503 9938
rect 2509 9934 2513 9938
rect 2519 9934 2523 9938
rect 2484 9929 2488 9933
rect 2494 9929 2498 9933
rect 2504 9929 2508 9933
rect 2514 9929 2518 9933
rect 2524 9929 2528 9933
rect 2489 9924 2493 9928
rect 2499 9924 2503 9928
rect 2509 9924 2513 9928
rect 2519 9924 2523 9928
rect 2484 9919 2488 9923
rect 2494 9919 2498 9923
rect 2504 9919 2508 9923
rect 2514 9919 2518 9923
rect 2524 9919 2528 9923
rect 2489 9914 2493 9918
rect 2499 9914 2503 9918
rect 2509 9914 2513 9918
rect 2519 9914 2523 9918
rect 2484 9909 2488 9913
rect 2494 9909 2498 9913
rect 2504 9909 2508 9913
rect 2514 9909 2518 9913
rect 2524 9909 2528 9913
rect 2489 9904 2493 9908
rect 2499 9904 2503 9908
rect 2509 9904 2513 9908
rect 2519 9904 2523 9908
rect 2484 9899 2488 9903
rect 2494 9899 2498 9903
rect 2504 9899 2508 9903
rect 2514 9899 2518 9903
rect 2524 9899 2528 9903
rect 2489 9894 2493 9898
rect 2499 9894 2503 9898
rect 2509 9894 2513 9898
rect 2519 9894 2523 9898
rect 2484 9889 2488 9893
rect 2494 9889 2498 9893
rect 2504 9889 2508 9893
rect 2514 9889 2518 9893
rect 2524 9889 2528 9893
rect 2489 9884 2493 9888
rect 2499 9884 2503 9888
rect 2509 9884 2513 9888
rect 2519 9884 2523 9888
rect 2484 9879 2488 9883
rect 2494 9879 2498 9883
rect 2504 9879 2508 9883
rect 2514 9879 2518 9883
rect 2524 9879 2528 9883
rect 2489 9874 2493 9878
rect 2499 9874 2503 9878
rect 2509 9874 2513 9878
rect 2519 9874 2523 9878
rect 2484 9869 2488 9873
rect 2494 9869 2498 9873
rect 2504 9869 2508 9873
rect 2514 9869 2518 9873
rect 2524 9869 2528 9873
rect 2489 9864 2493 9868
rect 2499 9864 2503 9868
rect 2509 9864 2513 9868
rect 2519 9864 2523 9868
rect 2472 9848 2476 9852
rect 2479 9848 2483 9852
rect 2484 9848 2488 9852
rect 2489 9848 2493 9852
rect 2494 9848 2498 9852
rect 2499 9848 2503 9852
rect 2504 9848 2508 9852
rect 2509 9848 2513 9852
rect 2514 9848 2518 9852
rect 2519 9848 2523 9852
rect 2524 9848 2528 9852
rect 2529 9848 2533 9852
rect 2536 9848 2540 9852
rect 2087 9827 2091 9831
rect 2145 9827 2149 9831
rect 2087 9811 2091 9815
rect 2145 9811 2149 9815
rect 1836 9795 1840 9799
rect 1673 9786 1677 9790
rect 1678 9786 1682 9790
rect 1673 9781 1677 9785
rect 1678 9781 1682 9785
rect 1673 9776 1677 9780
rect 1678 9776 1682 9780
rect 1778 9779 1782 9783
rect 1673 9771 1677 9775
rect 1678 9771 1682 9775
rect 1673 9766 1677 9770
rect 1678 9766 1682 9770
rect 1628 9757 1632 9761
rect 1633 9757 1637 9761
rect 1638 9757 1642 9761
rect 1643 9757 1647 9761
rect 1628 9747 1632 9751
rect 1633 9747 1637 9751
rect 1638 9747 1642 9751
rect 1643 9747 1647 9751
rect 1628 9737 1632 9741
rect 1633 9737 1637 9741
rect 1638 9737 1642 9741
rect 1643 9737 1647 9741
rect 1673 9761 1677 9765
rect 1678 9761 1682 9765
rect 1673 9756 1677 9760
rect 1678 9756 1682 9760
rect 1673 9751 1677 9755
rect 1678 9751 1682 9755
rect 1673 9746 1677 9750
rect 1678 9746 1682 9750
rect 1673 9741 1677 9745
rect 1678 9741 1682 9745
rect 1673 9736 1677 9740
rect 1678 9736 1682 9740
rect 1569 9718 1573 9722
rect 1574 9718 1578 9722
rect 1579 9718 1583 9722
rect 1584 9718 1588 9722
rect 1589 9718 1593 9722
rect 1594 9718 1598 9722
rect 1599 9718 1603 9722
rect 1604 9718 1608 9722
rect 1609 9718 1613 9722
rect 1614 9718 1618 9722
rect 1619 9718 1623 9722
rect 1569 9713 1573 9717
rect 1574 9713 1578 9717
rect 1579 9713 1583 9717
rect 1584 9713 1588 9717
rect 1589 9713 1593 9717
rect 1594 9713 1598 9717
rect 1599 9713 1603 9717
rect 1604 9713 1608 9717
rect 1609 9713 1613 9717
rect 1614 9713 1618 9717
rect 1619 9713 1623 9717
rect 1499 9706 1503 9710
rect 1504 9706 1508 9710
rect 1499 9701 1503 9705
rect 1504 9701 1508 9705
rect 1499 9696 1503 9700
rect 1504 9696 1508 9700
rect 1499 9691 1503 9695
rect 1504 9691 1508 9695
rect 1499 9686 1503 9690
rect 1504 9686 1508 9690
rect 1628 9711 1632 9715
rect 1633 9711 1637 9715
rect 1638 9711 1642 9715
rect 1643 9711 1647 9715
rect 1628 9701 1632 9705
rect 1633 9701 1637 9705
rect 1638 9701 1642 9705
rect 1643 9701 1647 9705
rect 1628 9691 1632 9695
rect 1633 9691 1637 9695
rect 1638 9691 1642 9695
rect 1643 9691 1647 9695
rect 1499 9681 1503 9685
rect 1504 9681 1508 9685
rect 1499 9676 1503 9680
rect 1504 9676 1508 9680
rect 1499 9671 1503 9675
rect 1504 9671 1508 9675
rect 1499 9666 1503 9670
rect 1504 9666 1508 9670
rect 1499 9661 1503 9665
rect 1504 9661 1508 9665
rect 664 9603 668 9607
rect 674 9603 678 9607
rect 684 9603 688 9607
rect 618 9592 622 9596
rect 628 9592 632 9596
rect 638 9592 642 9596
rect 618 9587 622 9591
rect 628 9587 632 9591
rect 638 9587 642 9591
rect 618 9582 622 9586
rect 628 9582 632 9586
rect 638 9582 642 9586
rect 618 9577 622 9581
rect 628 9577 632 9581
rect 638 9577 642 9581
rect 664 9592 668 9596
rect 674 9592 678 9596
rect 684 9592 688 9596
rect 1836 9779 1840 9783
rect 1982 9796 1986 9800
rect 1987 9796 1991 9800
rect 2087 9795 2091 9799
rect 1982 9791 1986 9795
rect 1987 9791 1991 9795
rect 2633 9949 2637 9953
rect 2643 9949 2647 9953
rect 2653 9949 2657 9953
rect 2663 9949 2667 9953
rect 2673 9949 2677 9953
rect 2638 9944 2642 9948
rect 2648 9944 2652 9948
rect 2658 9944 2662 9948
rect 2668 9944 2672 9948
rect 2633 9939 2637 9943
rect 2643 9939 2647 9943
rect 2653 9939 2657 9943
rect 2663 9939 2667 9943
rect 2673 9939 2677 9943
rect 2638 9934 2642 9938
rect 2648 9934 2652 9938
rect 2658 9934 2662 9938
rect 2668 9934 2672 9938
rect 2633 9929 2637 9933
rect 2643 9929 2647 9933
rect 2653 9929 2657 9933
rect 2663 9929 2667 9933
rect 2673 9929 2677 9933
rect 2638 9924 2642 9928
rect 2648 9924 2652 9928
rect 2658 9924 2662 9928
rect 2668 9924 2672 9928
rect 2633 9919 2637 9923
rect 2643 9919 2647 9923
rect 2653 9919 2657 9923
rect 2663 9919 2667 9923
rect 2673 9919 2677 9923
rect 2638 9914 2642 9918
rect 2648 9914 2652 9918
rect 2658 9914 2662 9918
rect 2668 9914 2672 9918
rect 2633 9909 2637 9913
rect 2643 9909 2647 9913
rect 2653 9909 2657 9913
rect 2663 9909 2667 9913
rect 2673 9909 2677 9913
rect 2638 9904 2642 9908
rect 2648 9904 2652 9908
rect 2658 9904 2662 9908
rect 2668 9904 2672 9908
rect 2633 9899 2637 9903
rect 2643 9899 2647 9903
rect 2653 9899 2657 9903
rect 2663 9899 2667 9903
rect 2673 9899 2677 9903
rect 2638 9894 2642 9898
rect 2648 9894 2652 9898
rect 2658 9894 2662 9898
rect 2668 9894 2672 9898
rect 2633 9889 2637 9893
rect 2643 9889 2647 9893
rect 2653 9889 2657 9893
rect 2663 9889 2667 9893
rect 2673 9889 2677 9893
rect 2638 9884 2642 9888
rect 2648 9884 2652 9888
rect 2658 9884 2662 9888
rect 2668 9884 2672 9888
rect 2633 9879 2637 9883
rect 2643 9879 2647 9883
rect 2653 9879 2657 9883
rect 2663 9879 2667 9883
rect 2673 9879 2677 9883
rect 2638 9874 2642 9878
rect 2648 9874 2652 9878
rect 2658 9874 2662 9878
rect 2668 9874 2672 9878
rect 2633 9869 2637 9873
rect 2643 9869 2647 9873
rect 2653 9869 2657 9873
rect 2663 9869 2667 9873
rect 2673 9869 2677 9873
rect 2638 9864 2642 9868
rect 2648 9864 2652 9868
rect 2658 9864 2662 9868
rect 2668 9864 2672 9868
rect 2621 9848 2625 9852
rect 2628 9848 2632 9852
rect 2633 9848 2637 9852
rect 2638 9848 2642 9852
rect 2643 9848 2647 9852
rect 2648 9848 2652 9852
rect 2653 9848 2657 9852
rect 2658 9848 2662 9852
rect 2663 9848 2667 9852
rect 2668 9848 2672 9852
rect 2673 9848 2677 9852
rect 2678 9848 2682 9852
rect 2685 9848 2689 9852
rect 2793 9949 2797 9953
rect 2803 9949 2807 9953
rect 2813 9949 2817 9953
rect 2823 9949 2827 9953
rect 2833 9949 2837 9953
rect 2798 9944 2802 9948
rect 2808 9944 2812 9948
rect 2818 9944 2822 9948
rect 2828 9944 2832 9948
rect 2793 9939 2797 9943
rect 2803 9939 2807 9943
rect 2813 9939 2817 9943
rect 2823 9939 2827 9943
rect 2833 9939 2837 9943
rect 2798 9934 2802 9938
rect 2808 9934 2812 9938
rect 2818 9934 2822 9938
rect 2828 9934 2832 9938
rect 2793 9929 2797 9933
rect 2803 9929 2807 9933
rect 2813 9929 2817 9933
rect 2823 9929 2827 9933
rect 2833 9929 2837 9933
rect 2798 9924 2802 9928
rect 2808 9924 2812 9928
rect 2818 9924 2822 9928
rect 2828 9924 2832 9928
rect 2793 9919 2797 9923
rect 2803 9919 2807 9923
rect 2813 9919 2817 9923
rect 2823 9919 2827 9923
rect 2833 9919 2837 9923
rect 2798 9914 2802 9918
rect 2808 9914 2812 9918
rect 2818 9914 2822 9918
rect 2828 9914 2832 9918
rect 2793 9909 2797 9913
rect 2803 9909 2807 9913
rect 2813 9909 2817 9913
rect 2823 9909 2827 9913
rect 2833 9909 2837 9913
rect 2798 9904 2802 9908
rect 2808 9904 2812 9908
rect 2818 9904 2822 9908
rect 2828 9904 2832 9908
rect 2793 9899 2797 9903
rect 2803 9899 2807 9903
rect 2813 9899 2817 9903
rect 2823 9899 2827 9903
rect 2833 9899 2837 9903
rect 2798 9894 2802 9898
rect 2808 9894 2812 9898
rect 2818 9894 2822 9898
rect 2828 9894 2832 9898
rect 2793 9889 2797 9893
rect 2803 9889 2807 9893
rect 2813 9889 2817 9893
rect 2823 9889 2827 9893
rect 2833 9889 2837 9893
rect 2798 9884 2802 9888
rect 2808 9884 2812 9888
rect 2818 9884 2822 9888
rect 2828 9884 2832 9888
rect 2793 9879 2797 9883
rect 2803 9879 2807 9883
rect 2813 9879 2817 9883
rect 2823 9879 2827 9883
rect 2833 9879 2837 9883
rect 2798 9874 2802 9878
rect 2808 9874 2812 9878
rect 2818 9874 2822 9878
rect 2828 9874 2832 9878
rect 2793 9869 2797 9873
rect 2803 9869 2807 9873
rect 2813 9869 2817 9873
rect 2823 9869 2827 9873
rect 2833 9869 2837 9873
rect 2798 9864 2802 9868
rect 2808 9864 2812 9868
rect 2818 9864 2822 9868
rect 2828 9864 2832 9868
rect 2781 9848 2785 9852
rect 2788 9848 2792 9852
rect 2793 9848 2797 9852
rect 2798 9848 2802 9852
rect 2803 9848 2807 9852
rect 2808 9848 2812 9852
rect 2813 9848 2817 9852
rect 2818 9848 2822 9852
rect 2823 9848 2827 9852
rect 2828 9848 2832 9852
rect 2833 9848 2837 9852
rect 2838 9848 2842 9852
rect 2845 9848 2849 9852
rect 2396 9827 2400 9831
rect 2454 9827 2458 9831
rect 2396 9811 2400 9815
rect 2454 9811 2458 9815
rect 2145 9795 2149 9799
rect 1982 9786 1986 9790
rect 1987 9786 1991 9790
rect 1982 9781 1986 9785
rect 1987 9781 1991 9785
rect 1982 9776 1986 9780
rect 1987 9776 1991 9780
rect 2087 9779 2091 9783
rect 1982 9771 1986 9775
rect 1987 9771 1991 9775
rect 1982 9766 1986 9770
rect 1987 9766 1991 9770
rect 1937 9757 1941 9761
rect 1942 9757 1946 9761
rect 1947 9757 1951 9761
rect 1952 9757 1956 9761
rect 1937 9747 1941 9751
rect 1942 9747 1946 9751
rect 1947 9747 1951 9751
rect 1952 9747 1956 9751
rect 1937 9737 1941 9741
rect 1942 9737 1946 9741
rect 1947 9737 1951 9741
rect 1952 9737 1956 9741
rect 1982 9761 1986 9765
rect 1987 9761 1991 9765
rect 1982 9756 1986 9760
rect 1987 9756 1991 9760
rect 1982 9751 1986 9755
rect 1987 9751 1991 9755
rect 1982 9746 1986 9750
rect 1987 9746 1991 9750
rect 1982 9741 1986 9745
rect 1987 9741 1991 9745
rect 1982 9736 1986 9740
rect 1987 9736 1991 9740
rect 1878 9718 1882 9722
rect 1883 9718 1887 9722
rect 1888 9718 1892 9722
rect 1893 9718 1897 9722
rect 1898 9718 1902 9722
rect 1903 9718 1907 9722
rect 1908 9718 1912 9722
rect 1913 9718 1917 9722
rect 1918 9718 1922 9722
rect 1923 9718 1927 9722
rect 1928 9718 1932 9722
rect 1878 9713 1882 9717
rect 1883 9713 1887 9717
rect 1888 9713 1892 9717
rect 1893 9713 1897 9717
rect 1898 9713 1902 9717
rect 1903 9713 1907 9717
rect 1908 9713 1912 9717
rect 1913 9713 1917 9717
rect 1918 9713 1922 9717
rect 1923 9713 1927 9717
rect 1928 9713 1932 9717
rect 1937 9711 1941 9715
rect 1942 9711 1946 9715
rect 1947 9711 1951 9715
rect 1952 9711 1956 9715
rect 1937 9701 1941 9705
rect 1942 9701 1946 9705
rect 1947 9701 1951 9705
rect 1952 9701 1956 9705
rect 1937 9691 1941 9695
rect 1942 9691 1946 9695
rect 1947 9691 1951 9695
rect 1952 9691 1956 9695
rect 2145 9779 2149 9783
rect 2291 9796 2295 9800
rect 2296 9796 2300 9800
rect 2396 9795 2400 9799
rect 2291 9791 2295 9795
rect 2296 9791 2300 9795
rect 2942 9949 2946 9953
rect 2952 9949 2956 9953
rect 2962 9949 2966 9953
rect 2972 9949 2976 9953
rect 2982 9949 2986 9953
rect 2947 9944 2951 9948
rect 2957 9944 2961 9948
rect 2967 9944 2971 9948
rect 2977 9944 2981 9948
rect 2942 9939 2946 9943
rect 2952 9939 2956 9943
rect 2962 9939 2966 9943
rect 2972 9939 2976 9943
rect 2982 9939 2986 9943
rect 2947 9934 2951 9938
rect 2957 9934 2961 9938
rect 2967 9934 2971 9938
rect 2977 9934 2981 9938
rect 2942 9929 2946 9933
rect 2952 9929 2956 9933
rect 2962 9929 2966 9933
rect 2972 9929 2976 9933
rect 2982 9929 2986 9933
rect 2947 9924 2951 9928
rect 2957 9924 2961 9928
rect 2967 9924 2971 9928
rect 2977 9924 2981 9928
rect 2942 9919 2946 9923
rect 2952 9919 2956 9923
rect 2962 9919 2966 9923
rect 2972 9919 2976 9923
rect 2982 9919 2986 9923
rect 2947 9914 2951 9918
rect 2957 9914 2961 9918
rect 2967 9914 2971 9918
rect 2977 9914 2981 9918
rect 2942 9909 2946 9913
rect 2952 9909 2956 9913
rect 2962 9909 2966 9913
rect 2972 9909 2976 9913
rect 2982 9909 2986 9913
rect 2947 9904 2951 9908
rect 2957 9904 2961 9908
rect 2967 9904 2971 9908
rect 2977 9904 2981 9908
rect 2942 9899 2946 9903
rect 2952 9899 2956 9903
rect 2962 9899 2966 9903
rect 2972 9899 2976 9903
rect 2982 9899 2986 9903
rect 2947 9894 2951 9898
rect 2957 9894 2961 9898
rect 2967 9894 2971 9898
rect 2977 9894 2981 9898
rect 2942 9889 2946 9893
rect 2952 9889 2956 9893
rect 2962 9889 2966 9893
rect 2972 9889 2976 9893
rect 2982 9889 2986 9893
rect 2947 9884 2951 9888
rect 2957 9884 2961 9888
rect 2967 9884 2971 9888
rect 2977 9884 2981 9888
rect 2942 9879 2946 9883
rect 2952 9879 2956 9883
rect 2962 9879 2966 9883
rect 2972 9879 2976 9883
rect 2982 9879 2986 9883
rect 2947 9874 2951 9878
rect 2957 9874 2961 9878
rect 2967 9874 2971 9878
rect 2977 9874 2981 9878
rect 2942 9869 2946 9873
rect 2952 9869 2956 9873
rect 2962 9869 2966 9873
rect 2972 9869 2976 9873
rect 2982 9869 2986 9873
rect 2947 9864 2951 9868
rect 2957 9864 2961 9868
rect 2967 9864 2971 9868
rect 2977 9864 2981 9868
rect 2930 9848 2934 9852
rect 2937 9848 2941 9852
rect 2942 9848 2946 9852
rect 2947 9848 2951 9852
rect 2952 9848 2956 9852
rect 2957 9848 2961 9852
rect 2962 9848 2966 9852
rect 2967 9848 2971 9852
rect 2972 9848 2976 9852
rect 2977 9848 2981 9852
rect 2982 9848 2986 9852
rect 2987 9848 2991 9852
rect 2994 9848 2998 9852
rect 3102 9949 3106 9953
rect 3112 9949 3116 9953
rect 3122 9949 3126 9953
rect 3132 9949 3136 9953
rect 3142 9949 3146 9953
rect 3107 9944 3111 9948
rect 3117 9944 3121 9948
rect 3127 9944 3131 9948
rect 3137 9944 3141 9948
rect 3102 9939 3106 9943
rect 3112 9939 3116 9943
rect 3122 9939 3126 9943
rect 3132 9939 3136 9943
rect 3142 9939 3146 9943
rect 3107 9934 3111 9938
rect 3117 9934 3121 9938
rect 3127 9934 3131 9938
rect 3137 9934 3141 9938
rect 3102 9929 3106 9933
rect 3112 9929 3116 9933
rect 3122 9929 3126 9933
rect 3132 9929 3136 9933
rect 3142 9929 3146 9933
rect 3107 9924 3111 9928
rect 3117 9924 3121 9928
rect 3127 9924 3131 9928
rect 3137 9924 3141 9928
rect 3102 9919 3106 9923
rect 3112 9919 3116 9923
rect 3122 9919 3126 9923
rect 3132 9919 3136 9923
rect 3142 9919 3146 9923
rect 3107 9914 3111 9918
rect 3117 9914 3121 9918
rect 3127 9914 3131 9918
rect 3137 9914 3141 9918
rect 3102 9909 3106 9913
rect 3112 9909 3116 9913
rect 3122 9909 3126 9913
rect 3132 9909 3136 9913
rect 3142 9909 3146 9913
rect 3107 9904 3111 9908
rect 3117 9904 3121 9908
rect 3127 9904 3131 9908
rect 3137 9904 3141 9908
rect 3102 9899 3106 9903
rect 3112 9899 3116 9903
rect 3122 9899 3126 9903
rect 3132 9899 3136 9903
rect 3142 9899 3146 9903
rect 3107 9894 3111 9898
rect 3117 9894 3121 9898
rect 3127 9894 3131 9898
rect 3137 9894 3141 9898
rect 3102 9889 3106 9893
rect 3112 9889 3116 9893
rect 3122 9889 3126 9893
rect 3132 9889 3136 9893
rect 3142 9889 3146 9893
rect 3107 9884 3111 9888
rect 3117 9884 3121 9888
rect 3127 9884 3131 9888
rect 3137 9884 3141 9888
rect 3102 9879 3106 9883
rect 3112 9879 3116 9883
rect 3122 9879 3126 9883
rect 3132 9879 3136 9883
rect 3142 9879 3146 9883
rect 3107 9874 3111 9878
rect 3117 9874 3121 9878
rect 3127 9874 3131 9878
rect 3137 9874 3141 9878
rect 3102 9869 3106 9873
rect 3112 9869 3116 9873
rect 3122 9869 3126 9873
rect 3132 9869 3136 9873
rect 3142 9869 3146 9873
rect 3107 9864 3111 9868
rect 3117 9864 3121 9868
rect 3127 9864 3131 9868
rect 3137 9864 3141 9868
rect 3090 9848 3094 9852
rect 3097 9848 3101 9852
rect 3102 9848 3106 9852
rect 3107 9848 3111 9852
rect 3112 9848 3116 9852
rect 3117 9848 3121 9852
rect 3122 9848 3126 9852
rect 3127 9848 3131 9852
rect 3132 9848 3136 9852
rect 3137 9848 3141 9852
rect 3142 9848 3146 9852
rect 3147 9848 3151 9852
rect 3154 9848 3158 9852
rect 2705 9827 2709 9831
rect 2763 9827 2767 9831
rect 2705 9811 2709 9815
rect 2763 9811 2767 9815
rect 2454 9795 2458 9799
rect 2291 9786 2295 9790
rect 2296 9786 2300 9790
rect 2291 9781 2295 9785
rect 2296 9781 2300 9785
rect 2291 9776 2295 9780
rect 2296 9776 2300 9780
rect 2396 9779 2400 9783
rect 2291 9771 2295 9775
rect 2296 9771 2300 9775
rect 2291 9766 2295 9770
rect 2296 9766 2300 9770
rect 2246 9757 2250 9761
rect 2251 9757 2255 9761
rect 2256 9757 2260 9761
rect 2261 9757 2265 9761
rect 2246 9747 2250 9751
rect 2251 9747 2255 9751
rect 2256 9747 2260 9751
rect 2261 9747 2265 9751
rect 2246 9737 2250 9741
rect 2251 9737 2255 9741
rect 2256 9737 2260 9741
rect 2261 9737 2265 9741
rect 2291 9761 2295 9765
rect 2296 9761 2300 9765
rect 2291 9756 2295 9760
rect 2296 9756 2300 9760
rect 2291 9751 2295 9755
rect 2296 9751 2300 9755
rect 2291 9746 2295 9750
rect 2296 9746 2300 9750
rect 2291 9741 2295 9745
rect 2296 9741 2300 9745
rect 2291 9736 2295 9740
rect 2296 9736 2300 9740
rect 2187 9718 2191 9722
rect 2192 9718 2196 9722
rect 2197 9718 2201 9722
rect 2202 9718 2206 9722
rect 2207 9718 2211 9722
rect 2212 9718 2216 9722
rect 2217 9718 2221 9722
rect 2222 9718 2226 9722
rect 2227 9718 2231 9722
rect 2232 9718 2236 9722
rect 2237 9718 2241 9722
rect 2187 9713 2191 9717
rect 2192 9713 2196 9717
rect 2197 9713 2201 9717
rect 2202 9713 2206 9717
rect 2207 9713 2211 9717
rect 2212 9713 2216 9717
rect 2217 9713 2221 9717
rect 2222 9713 2226 9717
rect 2227 9713 2231 9717
rect 2232 9713 2236 9717
rect 2237 9713 2241 9717
rect 2246 9711 2250 9715
rect 2251 9711 2255 9715
rect 2256 9711 2260 9715
rect 2261 9711 2265 9715
rect 2246 9701 2250 9705
rect 2251 9701 2255 9705
rect 2256 9701 2260 9705
rect 2261 9701 2265 9705
rect 2246 9691 2250 9695
rect 2251 9691 2255 9695
rect 2256 9691 2260 9695
rect 2261 9691 2265 9695
rect 2113 9593 2126 9597
rect 2454 9779 2458 9783
rect 2600 9796 2604 9800
rect 2605 9796 2609 9800
rect 2705 9795 2709 9799
rect 2600 9791 2604 9795
rect 2605 9791 2609 9795
rect 3251 9949 3255 9953
rect 3261 9949 3265 9953
rect 3271 9949 3275 9953
rect 3281 9949 3285 9953
rect 3291 9949 3295 9953
rect 3256 9944 3260 9948
rect 3266 9944 3270 9948
rect 3276 9944 3280 9948
rect 3286 9944 3290 9948
rect 3251 9939 3255 9943
rect 3261 9939 3265 9943
rect 3271 9939 3275 9943
rect 3281 9939 3285 9943
rect 3291 9939 3295 9943
rect 3256 9934 3260 9938
rect 3266 9934 3270 9938
rect 3276 9934 3280 9938
rect 3286 9934 3290 9938
rect 3251 9929 3255 9933
rect 3261 9929 3265 9933
rect 3271 9929 3275 9933
rect 3281 9929 3285 9933
rect 3291 9929 3295 9933
rect 3256 9924 3260 9928
rect 3266 9924 3270 9928
rect 3276 9924 3280 9928
rect 3286 9924 3290 9928
rect 3251 9919 3255 9923
rect 3261 9919 3265 9923
rect 3271 9919 3275 9923
rect 3281 9919 3285 9923
rect 3291 9919 3295 9923
rect 3256 9914 3260 9918
rect 3266 9914 3270 9918
rect 3276 9914 3280 9918
rect 3286 9914 3290 9918
rect 3251 9909 3255 9913
rect 3261 9909 3265 9913
rect 3271 9909 3275 9913
rect 3281 9909 3285 9913
rect 3291 9909 3295 9913
rect 3256 9904 3260 9908
rect 3266 9904 3270 9908
rect 3276 9904 3280 9908
rect 3286 9904 3290 9908
rect 3251 9899 3255 9903
rect 3261 9899 3265 9903
rect 3271 9899 3275 9903
rect 3281 9899 3285 9903
rect 3291 9899 3295 9903
rect 3256 9894 3260 9898
rect 3266 9894 3270 9898
rect 3276 9894 3280 9898
rect 3286 9894 3290 9898
rect 3251 9889 3255 9893
rect 3261 9889 3265 9893
rect 3271 9889 3275 9893
rect 3281 9889 3285 9893
rect 3291 9889 3295 9893
rect 3256 9884 3260 9888
rect 3266 9884 3270 9888
rect 3276 9884 3280 9888
rect 3286 9884 3290 9888
rect 3251 9879 3255 9883
rect 3261 9879 3265 9883
rect 3271 9879 3275 9883
rect 3281 9879 3285 9883
rect 3291 9879 3295 9883
rect 3256 9874 3260 9878
rect 3266 9874 3270 9878
rect 3276 9874 3280 9878
rect 3286 9874 3290 9878
rect 3251 9869 3255 9873
rect 3261 9869 3265 9873
rect 3271 9869 3275 9873
rect 3281 9869 3285 9873
rect 3291 9869 3295 9873
rect 3256 9864 3260 9868
rect 3266 9864 3270 9868
rect 3276 9864 3280 9868
rect 3286 9864 3290 9868
rect 3239 9848 3243 9852
rect 3246 9848 3250 9852
rect 3251 9848 3255 9852
rect 3256 9848 3260 9852
rect 3261 9848 3265 9852
rect 3266 9848 3270 9852
rect 3271 9848 3275 9852
rect 3276 9848 3280 9852
rect 3281 9848 3285 9852
rect 3286 9848 3290 9852
rect 3291 9848 3295 9852
rect 3296 9848 3300 9852
rect 3303 9848 3307 9852
rect 3014 9827 3018 9831
rect 3072 9827 3076 9831
rect 3014 9811 3018 9815
rect 3072 9811 3076 9815
rect 2763 9795 2767 9799
rect 2600 9786 2604 9790
rect 2605 9786 2609 9790
rect 2600 9781 2604 9785
rect 2605 9781 2609 9785
rect 2600 9776 2604 9780
rect 2605 9776 2609 9780
rect 2705 9779 2709 9783
rect 2600 9771 2604 9775
rect 2605 9771 2609 9775
rect 2600 9766 2604 9770
rect 2605 9766 2609 9770
rect 2555 9757 2559 9761
rect 2560 9757 2564 9761
rect 2565 9757 2569 9761
rect 2570 9757 2574 9761
rect 2555 9747 2559 9751
rect 2560 9747 2564 9751
rect 2565 9747 2569 9751
rect 2570 9747 2574 9751
rect 2555 9737 2559 9741
rect 2560 9737 2564 9741
rect 2565 9737 2569 9741
rect 2570 9737 2574 9741
rect 2600 9761 2604 9765
rect 2605 9761 2609 9765
rect 2600 9756 2604 9760
rect 2605 9756 2609 9760
rect 2600 9751 2604 9755
rect 2605 9751 2609 9755
rect 2600 9746 2604 9750
rect 2605 9746 2609 9750
rect 2600 9741 2604 9745
rect 2605 9741 2609 9745
rect 2600 9736 2604 9740
rect 2605 9736 2609 9740
rect 2496 9718 2500 9722
rect 2501 9718 2505 9722
rect 2506 9718 2510 9722
rect 2511 9718 2515 9722
rect 2516 9718 2520 9722
rect 2521 9718 2525 9722
rect 2526 9718 2530 9722
rect 2531 9718 2535 9722
rect 2536 9718 2540 9722
rect 2541 9718 2545 9722
rect 2546 9718 2550 9722
rect 2496 9713 2500 9717
rect 2501 9713 2505 9717
rect 2506 9713 2510 9717
rect 2511 9713 2515 9717
rect 2516 9713 2520 9717
rect 2521 9713 2525 9717
rect 2526 9713 2530 9717
rect 2531 9713 2535 9717
rect 2536 9713 2540 9717
rect 2541 9713 2545 9717
rect 2546 9713 2550 9717
rect 2555 9711 2559 9715
rect 2560 9711 2564 9715
rect 2565 9711 2569 9715
rect 2570 9711 2574 9715
rect 2555 9701 2559 9705
rect 2560 9701 2564 9705
rect 2565 9701 2569 9705
rect 2570 9701 2574 9705
rect 2555 9691 2559 9695
rect 2560 9691 2564 9695
rect 2565 9691 2569 9695
rect 2570 9691 2574 9695
rect 2763 9779 2767 9783
rect 2909 9796 2913 9800
rect 2914 9796 2918 9800
rect 3014 9795 3018 9799
rect 2909 9791 2913 9795
rect 2914 9791 2918 9795
rect 3072 9795 3076 9799
rect 2909 9786 2913 9790
rect 2914 9786 2918 9790
rect 2909 9781 2913 9785
rect 2914 9781 2918 9785
rect 2909 9776 2913 9780
rect 2914 9776 2918 9780
rect 3014 9779 3018 9783
rect 2909 9771 2913 9775
rect 2914 9771 2918 9775
rect 2909 9766 2913 9770
rect 2914 9766 2918 9770
rect 2864 9757 2868 9761
rect 2869 9757 2873 9761
rect 2874 9757 2878 9761
rect 2879 9757 2883 9761
rect 2864 9747 2868 9751
rect 2869 9747 2873 9751
rect 2874 9747 2878 9751
rect 2879 9747 2883 9751
rect 2864 9737 2868 9741
rect 2869 9737 2873 9741
rect 2874 9737 2878 9741
rect 2879 9737 2883 9741
rect 2909 9761 2913 9765
rect 2914 9761 2918 9765
rect 2909 9756 2913 9760
rect 2914 9756 2918 9760
rect 2909 9751 2913 9755
rect 2914 9751 2918 9755
rect 2909 9746 2913 9750
rect 2914 9746 2918 9750
rect 2909 9741 2913 9745
rect 2914 9741 2918 9745
rect 2909 9736 2913 9740
rect 2914 9736 2918 9740
rect 2805 9718 2809 9722
rect 2810 9718 2814 9722
rect 2815 9718 2819 9722
rect 2820 9718 2824 9722
rect 2825 9718 2829 9722
rect 2830 9718 2834 9722
rect 2835 9718 2839 9722
rect 2840 9718 2844 9722
rect 2845 9718 2849 9722
rect 2850 9718 2854 9722
rect 2855 9718 2859 9722
rect 2805 9713 2809 9717
rect 2810 9713 2814 9717
rect 2815 9713 2819 9717
rect 2820 9713 2824 9717
rect 2825 9713 2829 9717
rect 2830 9713 2834 9717
rect 2835 9713 2839 9717
rect 2840 9713 2844 9717
rect 2845 9713 2849 9717
rect 2850 9713 2854 9717
rect 2855 9713 2859 9717
rect 2864 9711 2868 9715
rect 2869 9711 2873 9715
rect 2874 9711 2878 9715
rect 2879 9711 2883 9715
rect 2864 9701 2868 9705
rect 2869 9701 2873 9705
rect 2874 9701 2878 9705
rect 2879 9701 2883 9705
rect 2864 9691 2868 9695
rect 2869 9691 2873 9695
rect 2874 9691 2878 9695
rect 2879 9691 2883 9695
rect 3072 9779 3076 9783
rect 3218 9796 3222 9800
rect 3223 9796 3227 9800
rect 3218 9791 3222 9795
rect 3223 9791 3227 9795
rect 3218 9786 3222 9790
rect 3223 9786 3227 9790
rect 3218 9781 3222 9785
rect 3223 9781 3227 9785
rect 3218 9776 3222 9780
rect 3223 9776 3227 9780
rect 3218 9771 3222 9775
rect 3223 9771 3227 9775
rect 3218 9766 3222 9770
rect 3223 9766 3227 9770
rect 3173 9757 3177 9761
rect 3178 9757 3182 9761
rect 3183 9757 3187 9761
rect 3188 9757 3192 9761
rect 3173 9747 3177 9751
rect 3178 9747 3182 9751
rect 3183 9747 3187 9751
rect 3188 9747 3192 9751
rect 3173 9737 3177 9741
rect 3178 9737 3182 9741
rect 3183 9737 3187 9741
rect 3188 9737 3192 9741
rect 3218 9761 3222 9765
rect 3223 9761 3227 9765
rect 3218 9756 3222 9760
rect 3223 9756 3227 9760
rect 3218 9751 3222 9755
rect 3223 9751 3227 9755
rect 3218 9746 3222 9750
rect 3223 9746 3227 9750
rect 3218 9741 3222 9745
rect 3223 9741 3227 9745
rect 3218 9736 3222 9740
rect 3223 9736 3227 9740
rect 3114 9718 3118 9722
rect 3119 9718 3123 9722
rect 3124 9718 3128 9722
rect 3129 9718 3133 9722
rect 3134 9718 3138 9722
rect 3139 9718 3143 9722
rect 3144 9718 3148 9722
rect 3149 9718 3153 9722
rect 3154 9718 3158 9722
rect 3159 9718 3163 9722
rect 3164 9718 3168 9722
rect 3114 9713 3118 9717
rect 3119 9713 3123 9717
rect 3124 9713 3128 9717
rect 3129 9713 3133 9717
rect 3134 9713 3138 9717
rect 3139 9713 3143 9717
rect 3144 9713 3148 9717
rect 3149 9713 3153 9717
rect 3154 9713 3158 9717
rect 3159 9713 3163 9717
rect 3164 9713 3168 9717
rect 3173 9711 3177 9715
rect 3178 9711 3182 9715
rect 3183 9711 3187 9715
rect 3188 9711 3192 9715
rect 3173 9701 3177 9705
rect 3178 9701 3182 9705
rect 3183 9701 3187 9705
rect 3188 9701 3192 9705
rect 3173 9691 3177 9695
rect 3178 9691 3182 9695
rect 3183 9691 3187 9695
rect 3188 9691 3192 9695
rect 3411 9949 3415 9953
rect 3421 9949 3425 9953
rect 3431 9949 3435 9953
rect 3441 9949 3445 9953
rect 3451 9949 3455 9953
rect 3416 9944 3420 9948
rect 3426 9944 3430 9948
rect 3436 9944 3440 9948
rect 3446 9944 3450 9948
rect 3411 9939 3415 9943
rect 3421 9939 3425 9943
rect 3431 9939 3435 9943
rect 3441 9939 3445 9943
rect 3451 9939 3455 9943
rect 3416 9934 3420 9938
rect 3426 9934 3430 9938
rect 3436 9934 3440 9938
rect 3446 9934 3450 9938
rect 3411 9929 3415 9933
rect 3421 9929 3425 9933
rect 3431 9929 3435 9933
rect 3441 9929 3445 9933
rect 3451 9929 3455 9933
rect 3416 9924 3420 9928
rect 3426 9924 3430 9928
rect 3436 9924 3440 9928
rect 3446 9924 3450 9928
rect 3411 9919 3415 9923
rect 3421 9919 3425 9923
rect 3431 9919 3435 9923
rect 3441 9919 3445 9923
rect 3451 9919 3455 9923
rect 3416 9914 3420 9918
rect 3426 9914 3430 9918
rect 3436 9914 3440 9918
rect 3446 9914 3450 9918
rect 3411 9909 3415 9913
rect 3421 9909 3425 9913
rect 3431 9909 3435 9913
rect 3441 9909 3445 9913
rect 3451 9909 3455 9913
rect 3416 9904 3420 9908
rect 3426 9904 3430 9908
rect 3436 9904 3440 9908
rect 3446 9904 3450 9908
rect 3411 9899 3415 9903
rect 3421 9899 3425 9903
rect 3431 9899 3435 9903
rect 3441 9899 3445 9903
rect 3451 9899 3455 9903
rect 3416 9894 3420 9898
rect 3426 9894 3430 9898
rect 3436 9894 3440 9898
rect 3446 9894 3450 9898
rect 3411 9889 3415 9893
rect 3421 9889 3425 9893
rect 3431 9889 3435 9893
rect 3441 9889 3445 9893
rect 3451 9889 3455 9893
rect 3416 9884 3420 9888
rect 3426 9884 3430 9888
rect 3436 9884 3440 9888
rect 3446 9884 3450 9888
rect 3411 9879 3415 9883
rect 3421 9879 3425 9883
rect 3431 9879 3435 9883
rect 3441 9879 3445 9883
rect 3451 9879 3455 9883
rect 3416 9874 3420 9878
rect 3426 9874 3430 9878
rect 3436 9874 3440 9878
rect 3446 9874 3450 9878
rect 3411 9869 3415 9873
rect 3421 9869 3425 9873
rect 3431 9869 3435 9873
rect 3441 9869 3445 9873
rect 3451 9869 3455 9873
rect 3416 9864 3420 9868
rect 3426 9864 3430 9868
rect 3436 9864 3440 9868
rect 3446 9864 3450 9868
rect 3399 9848 3403 9852
rect 3406 9848 3410 9852
rect 3411 9848 3415 9852
rect 3416 9848 3420 9852
rect 3421 9848 3425 9852
rect 3426 9848 3430 9852
rect 3431 9848 3435 9852
rect 3436 9848 3440 9852
rect 3441 9848 3445 9852
rect 3446 9848 3450 9852
rect 3451 9848 3455 9852
rect 3456 9848 3460 9852
rect 3463 9848 3467 9852
rect 3560 9949 3564 9953
rect 3570 9949 3574 9953
rect 3580 9949 3584 9953
rect 3590 9949 3594 9953
rect 3600 9949 3604 9953
rect 3565 9944 3569 9948
rect 3575 9944 3579 9948
rect 3585 9944 3589 9948
rect 3595 9944 3599 9948
rect 3560 9939 3564 9943
rect 3570 9939 3574 9943
rect 3580 9939 3584 9943
rect 3590 9939 3594 9943
rect 3600 9939 3604 9943
rect 3565 9934 3569 9938
rect 3575 9934 3579 9938
rect 3585 9934 3589 9938
rect 3595 9934 3599 9938
rect 3560 9929 3564 9933
rect 3570 9929 3574 9933
rect 3580 9929 3584 9933
rect 3590 9929 3594 9933
rect 3600 9929 3604 9933
rect 3565 9924 3569 9928
rect 3575 9924 3579 9928
rect 3585 9924 3589 9928
rect 3595 9924 3599 9928
rect 3560 9919 3564 9923
rect 3570 9919 3574 9923
rect 3580 9919 3584 9923
rect 3590 9919 3594 9923
rect 3600 9919 3604 9923
rect 3565 9914 3569 9918
rect 3575 9914 3579 9918
rect 3585 9914 3589 9918
rect 3595 9914 3599 9918
rect 3560 9909 3564 9913
rect 3570 9909 3574 9913
rect 3580 9909 3584 9913
rect 3590 9909 3594 9913
rect 3600 9909 3604 9913
rect 3565 9904 3569 9908
rect 3575 9904 3579 9908
rect 3585 9904 3589 9908
rect 3595 9904 3599 9908
rect 3560 9899 3564 9903
rect 3570 9899 3574 9903
rect 3580 9899 3584 9903
rect 3590 9899 3594 9903
rect 3600 9899 3604 9903
rect 3565 9894 3569 9898
rect 3575 9894 3579 9898
rect 3585 9894 3589 9898
rect 3595 9894 3599 9898
rect 3560 9889 3564 9893
rect 3570 9889 3574 9893
rect 3580 9889 3584 9893
rect 3590 9889 3594 9893
rect 3600 9889 3604 9893
rect 3565 9884 3569 9888
rect 3575 9884 3579 9888
rect 3585 9884 3589 9888
rect 3595 9884 3599 9888
rect 3560 9879 3564 9883
rect 3570 9879 3574 9883
rect 3580 9879 3584 9883
rect 3590 9879 3594 9883
rect 3600 9879 3604 9883
rect 3565 9874 3569 9878
rect 3575 9874 3579 9878
rect 3585 9874 3589 9878
rect 3595 9874 3599 9878
rect 3560 9869 3564 9873
rect 3570 9869 3574 9873
rect 3580 9869 3584 9873
rect 3590 9869 3594 9873
rect 3600 9869 3604 9873
rect 3565 9864 3569 9868
rect 3575 9864 3579 9868
rect 3585 9864 3589 9868
rect 3595 9864 3599 9868
rect 3548 9848 3552 9852
rect 3555 9848 3559 9852
rect 3560 9848 3564 9852
rect 3565 9848 3569 9852
rect 3570 9848 3574 9852
rect 3575 9848 3579 9852
rect 3580 9848 3584 9852
rect 3585 9848 3589 9852
rect 3590 9848 3594 9852
rect 3595 9848 3599 9852
rect 3600 9848 3604 9852
rect 3605 9848 3609 9852
rect 3612 9848 3616 9852
rect 3353 9711 3357 9715
rect 3358 9711 3362 9715
rect 3527 9796 3531 9800
rect 3532 9796 3536 9800
rect 3527 9791 3531 9795
rect 3532 9791 3536 9795
rect 3527 9786 3531 9790
rect 3532 9786 3536 9790
rect 3527 9781 3531 9785
rect 3532 9781 3536 9785
rect 3527 9776 3531 9780
rect 3532 9776 3536 9780
rect 3527 9771 3531 9775
rect 3532 9771 3536 9775
rect 3527 9766 3531 9770
rect 3532 9766 3536 9770
rect 3482 9757 3486 9761
rect 3487 9757 3491 9761
rect 3492 9757 3496 9761
rect 3497 9757 3501 9761
rect 3482 9747 3486 9751
rect 3487 9747 3491 9751
rect 3492 9747 3496 9751
rect 3497 9747 3501 9751
rect 3482 9737 3486 9741
rect 3487 9737 3491 9741
rect 3492 9737 3496 9741
rect 3497 9737 3501 9741
rect 3527 9761 3531 9765
rect 3532 9761 3536 9765
rect 3527 9756 3531 9760
rect 3532 9756 3536 9760
rect 3527 9751 3531 9755
rect 3532 9751 3536 9755
rect 3527 9746 3531 9750
rect 3532 9746 3536 9750
rect 3527 9741 3531 9745
rect 3532 9741 3536 9745
rect 3527 9736 3531 9740
rect 3532 9736 3536 9740
rect 3720 9949 3724 9953
rect 3730 9949 3734 9953
rect 3740 9949 3744 9953
rect 3750 9949 3754 9953
rect 3760 9949 3764 9953
rect 3725 9944 3729 9948
rect 3735 9944 3739 9948
rect 3745 9944 3749 9948
rect 3755 9944 3759 9948
rect 3720 9939 3724 9943
rect 3730 9939 3734 9943
rect 3740 9939 3744 9943
rect 3750 9939 3754 9943
rect 3760 9939 3764 9943
rect 3725 9934 3729 9938
rect 3735 9934 3739 9938
rect 3745 9934 3749 9938
rect 3755 9934 3759 9938
rect 3720 9929 3724 9933
rect 3730 9929 3734 9933
rect 3740 9929 3744 9933
rect 3750 9929 3754 9933
rect 3760 9929 3764 9933
rect 3725 9924 3729 9928
rect 3735 9924 3739 9928
rect 3745 9924 3749 9928
rect 3755 9924 3759 9928
rect 3720 9919 3724 9923
rect 3730 9919 3734 9923
rect 3740 9919 3744 9923
rect 3750 9919 3754 9923
rect 3760 9919 3764 9923
rect 3725 9914 3729 9918
rect 3735 9914 3739 9918
rect 3745 9914 3749 9918
rect 3755 9914 3759 9918
rect 3720 9909 3724 9913
rect 3730 9909 3734 9913
rect 3740 9909 3744 9913
rect 3750 9909 3754 9913
rect 3760 9909 3764 9913
rect 3725 9904 3729 9908
rect 3735 9904 3739 9908
rect 3745 9904 3749 9908
rect 3755 9904 3759 9908
rect 3720 9899 3724 9903
rect 3730 9899 3734 9903
rect 3740 9899 3744 9903
rect 3750 9899 3754 9903
rect 3760 9899 3764 9903
rect 3725 9894 3729 9898
rect 3735 9894 3739 9898
rect 3745 9894 3749 9898
rect 3755 9894 3759 9898
rect 3720 9889 3724 9893
rect 3730 9889 3734 9893
rect 3740 9889 3744 9893
rect 3750 9889 3754 9893
rect 3760 9889 3764 9893
rect 3725 9884 3729 9888
rect 3735 9884 3739 9888
rect 3745 9884 3749 9888
rect 3755 9884 3759 9888
rect 3720 9879 3724 9883
rect 3730 9879 3734 9883
rect 3740 9879 3744 9883
rect 3750 9879 3754 9883
rect 3760 9879 3764 9883
rect 3725 9874 3729 9878
rect 3735 9874 3739 9878
rect 3745 9874 3749 9878
rect 3755 9874 3759 9878
rect 3720 9869 3724 9873
rect 3730 9869 3734 9873
rect 3740 9869 3744 9873
rect 3750 9869 3754 9873
rect 3760 9869 3764 9873
rect 3725 9864 3729 9868
rect 3735 9864 3739 9868
rect 3745 9864 3749 9868
rect 3755 9864 3759 9868
rect 3708 9848 3712 9852
rect 3715 9848 3719 9852
rect 3720 9848 3724 9852
rect 3725 9848 3729 9852
rect 3730 9848 3734 9852
rect 3735 9848 3739 9852
rect 3740 9848 3744 9852
rect 3745 9848 3749 9852
rect 3750 9848 3754 9852
rect 3755 9848 3759 9852
rect 3760 9848 3764 9852
rect 3765 9848 3769 9852
rect 3772 9848 3776 9852
rect 3869 9949 3873 9953
rect 3879 9949 3883 9953
rect 3889 9949 3893 9953
rect 3899 9949 3903 9953
rect 3909 9949 3913 9953
rect 3874 9944 3878 9948
rect 3884 9944 3888 9948
rect 3894 9944 3898 9948
rect 3904 9944 3908 9948
rect 3869 9939 3873 9943
rect 3879 9939 3883 9943
rect 3889 9939 3893 9943
rect 3899 9939 3903 9943
rect 3909 9939 3913 9943
rect 3874 9934 3878 9938
rect 3884 9934 3888 9938
rect 3894 9934 3898 9938
rect 3904 9934 3908 9938
rect 3869 9929 3873 9933
rect 3879 9929 3883 9933
rect 3889 9929 3893 9933
rect 3899 9929 3903 9933
rect 3909 9929 3913 9933
rect 3874 9924 3878 9928
rect 3884 9924 3888 9928
rect 3894 9924 3898 9928
rect 3904 9924 3908 9928
rect 3869 9919 3873 9923
rect 3879 9919 3883 9923
rect 3889 9919 3893 9923
rect 3899 9919 3903 9923
rect 3909 9919 3913 9923
rect 3874 9914 3878 9918
rect 3884 9914 3888 9918
rect 3894 9914 3898 9918
rect 3904 9914 3908 9918
rect 3869 9909 3873 9913
rect 3879 9909 3883 9913
rect 3889 9909 3893 9913
rect 3899 9909 3903 9913
rect 3909 9909 3913 9913
rect 3874 9904 3878 9908
rect 3884 9904 3888 9908
rect 3894 9904 3898 9908
rect 3904 9904 3908 9908
rect 3869 9899 3873 9903
rect 3879 9899 3883 9903
rect 3889 9899 3893 9903
rect 3899 9899 3903 9903
rect 3909 9899 3913 9903
rect 3874 9894 3878 9898
rect 3884 9894 3888 9898
rect 3894 9894 3898 9898
rect 3904 9894 3908 9898
rect 3869 9889 3873 9893
rect 3879 9889 3883 9893
rect 3889 9889 3893 9893
rect 3899 9889 3903 9893
rect 3909 9889 3913 9893
rect 3874 9884 3878 9888
rect 3884 9884 3888 9888
rect 3894 9884 3898 9888
rect 3904 9884 3908 9888
rect 3869 9879 3873 9883
rect 3879 9879 3883 9883
rect 3889 9879 3893 9883
rect 3899 9879 3903 9883
rect 3909 9879 3913 9883
rect 3874 9874 3878 9878
rect 3884 9874 3888 9878
rect 3894 9874 3898 9878
rect 3904 9874 3908 9878
rect 3869 9869 3873 9873
rect 3879 9869 3883 9873
rect 3889 9869 3893 9873
rect 3899 9869 3903 9873
rect 3909 9869 3913 9873
rect 3874 9864 3878 9868
rect 3884 9864 3888 9868
rect 3894 9864 3898 9868
rect 3904 9864 3908 9868
rect 3857 9848 3861 9852
rect 3864 9848 3868 9852
rect 3869 9848 3873 9852
rect 3874 9848 3878 9852
rect 3879 9848 3883 9852
rect 3884 9848 3888 9852
rect 3889 9848 3893 9852
rect 3894 9848 3898 9852
rect 3899 9848 3903 9852
rect 3904 9848 3908 9852
rect 3909 9848 3913 9852
rect 3914 9848 3918 9852
rect 3921 9848 3925 9852
rect 4029 9949 4033 9953
rect 4039 9949 4043 9953
rect 4049 9949 4053 9953
rect 4059 9949 4063 9953
rect 4069 9949 4073 9953
rect 4034 9944 4038 9948
rect 4044 9944 4048 9948
rect 4054 9944 4058 9948
rect 4064 9944 4068 9948
rect 4029 9939 4033 9943
rect 4039 9939 4043 9943
rect 4049 9939 4053 9943
rect 4059 9939 4063 9943
rect 4069 9939 4073 9943
rect 4034 9934 4038 9938
rect 4044 9934 4048 9938
rect 4054 9934 4058 9938
rect 4064 9934 4068 9938
rect 4029 9929 4033 9933
rect 4039 9929 4043 9933
rect 4049 9929 4053 9933
rect 4059 9929 4063 9933
rect 4069 9929 4073 9933
rect 4034 9924 4038 9928
rect 4044 9924 4048 9928
rect 4054 9924 4058 9928
rect 4064 9924 4068 9928
rect 4029 9919 4033 9923
rect 4039 9919 4043 9923
rect 4049 9919 4053 9923
rect 4059 9919 4063 9923
rect 4069 9919 4073 9923
rect 4034 9914 4038 9918
rect 4044 9914 4048 9918
rect 4054 9914 4058 9918
rect 4064 9914 4068 9918
rect 4029 9909 4033 9913
rect 4039 9909 4043 9913
rect 4049 9909 4053 9913
rect 4059 9909 4063 9913
rect 4069 9909 4073 9913
rect 4034 9904 4038 9908
rect 4044 9904 4048 9908
rect 4054 9904 4058 9908
rect 4064 9904 4068 9908
rect 4029 9899 4033 9903
rect 4039 9899 4043 9903
rect 4049 9899 4053 9903
rect 4059 9899 4063 9903
rect 4069 9899 4073 9903
rect 4034 9894 4038 9898
rect 4044 9894 4048 9898
rect 4054 9894 4058 9898
rect 4064 9894 4068 9898
rect 4029 9889 4033 9893
rect 4039 9889 4043 9893
rect 4049 9889 4053 9893
rect 4059 9889 4063 9893
rect 4069 9889 4073 9893
rect 4034 9884 4038 9888
rect 4044 9884 4048 9888
rect 4054 9884 4058 9888
rect 4064 9884 4068 9888
rect 4029 9879 4033 9883
rect 4039 9879 4043 9883
rect 4049 9879 4053 9883
rect 4059 9879 4063 9883
rect 4069 9879 4073 9883
rect 4034 9874 4038 9878
rect 4044 9874 4048 9878
rect 4054 9874 4058 9878
rect 4064 9874 4068 9878
rect 4029 9869 4033 9873
rect 4039 9869 4043 9873
rect 4049 9869 4053 9873
rect 4059 9869 4063 9873
rect 4069 9869 4073 9873
rect 4034 9864 4038 9868
rect 4044 9864 4048 9868
rect 4054 9864 4058 9868
rect 4064 9864 4068 9868
rect 4017 9848 4021 9852
rect 4024 9848 4028 9852
rect 4029 9848 4033 9852
rect 4034 9848 4038 9852
rect 4039 9848 4043 9852
rect 4044 9848 4048 9852
rect 4049 9848 4053 9852
rect 4054 9848 4058 9852
rect 4059 9848 4063 9852
rect 4064 9848 4068 9852
rect 4069 9848 4073 9852
rect 4074 9848 4078 9852
rect 4081 9848 4085 9852
rect 3662 9791 3666 9795
rect 3667 9791 3671 9795
rect 3662 9786 3666 9790
rect 3667 9786 3671 9790
rect 3662 9781 3666 9785
rect 3667 9781 3671 9785
rect 3662 9776 3666 9780
rect 3667 9776 3671 9780
rect 3662 9771 3666 9775
rect 3667 9771 3671 9775
rect 3662 9766 3666 9770
rect 3667 9766 3671 9770
rect 3662 9761 3666 9765
rect 3667 9761 3671 9765
rect 3662 9756 3666 9760
rect 3667 9756 3671 9760
rect 3662 9751 3666 9755
rect 3667 9751 3671 9755
rect 3662 9746 3666 9750
rect 3667 9746 3671 9750
rect 3662 9741 3666 9745
rect 3667 9741 3671 9745
rect 3423 9718 3427 9722
rect 3428 9718 3432 9722
rect 3433 9718 3437 9722
rect 3438 9718 3442 9722
rect 3443 9718 3447 9722
rect 3448 9718 3452 9722
rect 3453 9718 3457 9722
rect 3458 9718 3462 9722
rect 3463 9718 3467 9722
rect 3468 9718 3472 9722
rect 3473 9718 3477 9722
rect 3423 9713 3427 9717
rect 3428 9713 3432 9717
rect 3433 9713 3437 9717
rect 3438 9713 3442 9717
rect 3443 9713 3447 9717
rect 3448 9713 3452 9717
rect 3453 9713 3457 9717
rect 3458 9713 3462 9717
rect 3463 9713 3467 9717
rect 3468 9713 3472 9717
rect 3473 9713 3477 9717
rect 3353 9706 3357 9710
rect 3358 9706 3362 9710
rect 3353 9701 3357 9705
rect 3358 9701 3362 9705
rect 3353 9696 3357 9700
rect 3358 9696 3362 9700
rect 3353 9691 3357 9695
rect 3358 9691 3362 9695
rect 3353 9686 3357 9690
rect 3358 9686 3362 9690
rect 3482 9711 3486 9715
rect 3487 9711 3491 9715
rect 3492 9711 3496 9715
rect 3497 9711 3501 9715
rect 3482 9701 3486 9705
rect 3487 9701 3491 9705
rect 3492 9701 3496 9705
rect 3497 9701 3501 9705
rect 3482 9691 3486 9695
rect 3487 9691 3491 9695
rect 3492 9691 3496 9695
rect 3497 9691 3501 9695
rect 3021 9605 3026 9609
rect 3040 9607 3053 9611
rect 3353 9681 3357 9685
rect 3358 9681 3362 9685
rect 3353 9676 3357 9680
rect 3358 9676 3362 9680
rect 3353 9671 3357 9675
rect 3358 9671 3362 9675
rect 3353 9666 3357 9670
rect 3358 9666 3362 9670
rect 3353 9661 3357 9665
rect 3358 9661 3362 9665
rect 3327 9606 3379 9610
rect 3941 9827 3945 9831
rect 3999 9827 4003 9831
rect 3941 9811 3945 9815
rect 3999 9811 4003 9815
rect 3836 9796 3840 9800
rect 3841 9796 3845 9800
rect 3941 9795 3945 9799
rect 3836 9791 3840 9795
rect 3841 9791 3845 9795
rect 3999 9795 4003 9799
rect 3836 9786 3840 9790
rect 3841 9786 3845 9790
rect 3836 9781 3840 9785
rect 3841 9781 3845 9785
rect 3836 9776 3840 9780
rect 3841 9776 3845 9780
rect 3941 9779 3945 9783
rect 3836 9771 3840 9775
rect 3841 9771 3845 9775
rect 3836 9766 3840 9770
rect 3841 9766 3845 9770
rect 3791 9757 3795 9761
rect 3796 9757 3800 9761
rect 3801 9757 3805 9761
rect 3806 9757 3810 9761
rect 3791 9747 3795 9751
rect 3796 9747 3800 9751
rect 3801 9747 3805 9751
rect 3806 9747 3810 9751
rect 3791 9737 3795 9741
rect 3796 9737 3800 9741
rect 3801 9737 3805 9741
rect 3806 9737 3810 9741
rect 3836 9761 3840 9765
rect 3841 9761 3845 9765
rect 3836 9756 3840 9760
rect 3841 9756 3845 9760
rect 3836 9751 3840 9755
rect 3841 9751 3845 9755
rect 3836 9746 3840 9750
rect 3841 9746 3845 9750
rect 3836 9741 3840 9745
rect 3841 9741 3845 9745
rect 3836 9736 3840 9740
rect 3841 9736 3845 9740
rect 3732 9718 3736 9722
rect 3737 9718 3741 9722
rect 3742 9718 3746 9722
rect 3747 9718 3751 9722
rect 3752 9718 3756 9722
rect 3757 9718 3761 9722
rect 3762 9718 3766 9722
rect 3767 9718 3771 9722
rect 3772 9718 3776 9722
rect 3777 9718 3781 9722
rect 3782 9718 3786 9722
rect 3732 9713 3736 9717
rect 3737 9713 3741 9717
rect 3742 9713 3746 9717
rect 3747 9713 3751 9717
rect 3752 9713 3756 9717
rect 3757 9713 3761 9717
rect 3762 9713 3766 9717
rect 3767 9713 3771 9717
rect 3772 9713 3776 9717
rect 3777 9713 3781 9717
rect 3782 9713 3786 9717
rect 3791 9711 3795 9715
rect 3796 9711 3800 9715
rect 3801 9711 3805 9715
rect 3806 9711 3810 9715
rect 3791 9701 3795 9705
rect 3796 9701 3800 9705
rect 3801 9701 3805 9705
rect 3806 9701 3810 9705
rect 3791 9691 3795 9695
rect 3796 9691 3800 9695
rect 3801 9691 3805 9695
rect 3806 9691 3810 9695
rect 3634 9604 3690 9609
rect 664 9587 668 9591
rect 674 9587 678 9591
rect 684 9587 688 9591
rect 664 9582 668 9586
rect 674 9582 678 9586
rect 684 9582 688 9586
rect 664 9577 668 9581
rect 674 9577 678 9581
rect 684 9577 688 9581
rect 2422 9575 2435 9597
rect 2497 9575 2502 9597
rect 3999 9779 4003 9783
rect 4100 9757 4104 9761
rect 4105 9757 4109 9761
rect 4110 9757 4114 9761
rect 4115 9757 4119 9761
rect 4100 9747 4104 9751
rect 4105 9747 4109 9751
rect 4110 9747 4114 9751
rect 4115 9747 4119 9751
rect 4100 9737 4104 9741
rect 4105 9737 4109 9741
rect 4110 9737 4114 9741
rect 4115 9737 4119 9741
rect 4292 9757 4296 9761
rect 4297 9757 4301 9761
rect 4302 9757 4306 9761
rect 4307 9757 4311 9761
rect 4292 9747 4296 9751
rect 4297 9747 4301 9751
rect 4302 9747 4306 9751
rect 4307 9747 4311 9751
rect 4292 9737 4296 9741
rect 4297 9737 4301 9741
rect 4302 9737 4306 9741
rect 4307 9737 4311 9741
rect 4318 9757 4322 9761
rect 4323 9757 4327 9761
rect 4328 9757 4332 9761
rect 4333 9757 4337 9761
rect 4318 9747 4322 9751
rect 4323 9747 4327 9751
rect 4328 9747 4332 9751
rect 4333 9747 4337 9751
rect 4318 9737 4322 9741
rect 4323 9737 4327 9741
rect 4328 9737 4332 9741
rect 4333 9737 4337 9741
rect 4344 9757 4348 9761
rect 4349 9757 4353 9761
rect 4354 9757 4358 9761
rect 4359 9757 4363 9761
rect 4344 9747 4348 9751
rect 4349 9747 4353 9751
rect 4354 9747 4358 9751
rect 4359 9747 4363 9751
rect 4344 9737 4348 9741
rect 4349 9737 4353 9741
rect 4354 9737 4358 9741
rect 4359 9737 4363 9741
rect 4370 9757 4374 9761
rect 4375 9757 4379 9761
rect 4380 9757 4384 9761
rect 4385 9757 4389 9761
rect 4370 9747 4374 9751
rect 4375 9747 4379 9751
rect 4380 9747 4384 9751
rect 4385 9747 4389 9751
rect 4370 9737 4374 9741
rect 4375 9737 4379 9741
rect 4380 9737 4384 9741
rect 4385 9737 4389 9741
rect 4396 9757 4400 9761
rect 4401 9757 4405 9761
rect 4406 9757 4410 9761
rect 4411 9757 4415 9761
rect 4396 9747 4400 9751
rect 4401 9747 4405 9751
rect 4406 9747 4410 9751
rect 4411 9747 4415 9751
rect 4396 9737 4400 9741
rect 4401 9737 4405 9741
rect 4406 9737 4410 9741
rect 4411 9737 4415 9741
rect 4041 9718 4045 9722
rect 4046 9718 4050 9722
rect 4051 9718 4055 9722
rect 4056 9718 4060 9722
rect 4061 9718 4065 9722
rect 4066 9718 4070 9722
rect 4071 9718 4075 9722
rect 4076 9718 4080 9722
rect 4081 9718 4085 9722
rect 4086 9718 4090 9722
rect 4091 9718 4095 9722
rect 4041 9713 4045 9717
rect 4046 9713 4050 9717
rect 4051 9713 4055 9717
rect 4056 9713 4060 9717
rect 4061 9713 4065 9717
rect 4066 9713 4070 9717
rect 4071 9713 4075 9717
rect 4076 9713 4080 9717
rect 4081 9713 4085 9717
rect 4086 9713 4090 9717
rect 4091 9713 4095 9717
rect 4100 9711 4104 9715
rect 4105 9711 4109 9715
rect 4110 9711 4114 9715
rect 4115 9711 4119 9715
rect 4100 9701 4104 9705
rect 4105 9701 4109 9705
rect 4110 9701 4114 9705
rect 4115 9701 4119 9705
rect 4100 9691 4104 9695
rect 4105 9691 4109 9695
rect 4110 9691 4114 9695
rect 4115 9691 4119 9695
rect 4292 9711 4296 9715
rect 4297 9711 4301 9715
rect 4302 9711 4306 9715
rect 4307 9711 4311 9715
rect 4292 9701 4296 9705
rect 4297 9701 4301 9705
rect 4302 9701 4306 9705
rect 4307 9701 4311 9705
rect 4292 9691 4296 9695
rect 4297 9691 4301 9695
rect 4302 9691 4306 9695
rect 4307 9691 4311 9695
rect 4318 9711 4322 9715
rect 4323 9711 4327 9715
rect 4328 9711 4332 9715
rect 4333 9711 4337 9715
rect 4318 9701 4322 9705
rect 4323 9701 4327 9705
rect 4328 9701 4332 9705
rect 4333 9701 4337 9705
rect 4318 9691 4322 9695
rect 4323 9691 4327 9695
rect 4328 9691 4332 9695
rect 4333 9691 4337 9695
rect 4344 9711 4348 9715
rect 4349 9711 4353 9715
rect 4354 9711 4358 9715
rect 4359 9711 4363 9715
rect 4344 9701 4348 9705
rect 4349 9701 4353 9705
rect 4354 9701 4358 9705
rect 4359 9701 4363 9705
rect 4344 9691 4348 9695
rect 4349 9691 4353 9695
rect 4354 9691 4358 9695
rect 4359 9691 4363 9695
rect 4370 9711 4374 9715
rect 4375 9711 4379 9715
rect 4380 9711 4384 9715
rect 4385 9711 4389 9715
rect 4370 9701 4374 9705
rect 4375 9701 4379 9705
rect 4380 9701 4384 9705
rect 4385 9701 4389 9705
rect 4370 9691 4374 9695
rect 4375 9691 4379 9695
rect 4380 9691 4384 9695
rect 4385 9691 4389 9695
rect 4396 9711 4400 9715
rect 4401 9711 4405 9715
rect 4406 9711 4410 9715
rect 4411 9711 4415 9715
rect 4396 9701 4400 9705
rect 4401 9701 4405 9705
rect 4406 9701 4410 9705
rect 4411 9701 4415 9705
rect 4396 9691 4400 9695
rect 4401 9691 4405 9695
rect 4406 9691 4410 9695
rect 4411 9691 4415 9695
rect 618 9566 622 9570
rect 628 9566 632 9570
rect 638 9566 642 9570
rect 618 9561 622 9565
rect 628 9561 632 9565
rect 638 9561 642 9565
rect 618 9556 622 9560
rect 628 9556 632 9560
rect 638 9556 642 9560
rect 618 9551 622 9555
rect 628 9551 632 9555
rect 638 9551 642 9555
rect 664 9566 668 9570
rect 674 9566 678 9570
rect 684 9566 688 9570
rect 664 9561 668 9565
rect 674 9561 678 9565
rect 684 9561 688 9565
rect 664 9556 668 9560
rect 674 9556 678 9560
rect 684 9556 688 9560
rect 664 9551 668 9555
rect 674 9551 678 9555
rect 684 9551 688 9555
rect 2113 9547 2134 9572
rect 2401 9549 2414 9571
rect 2476 9549 2481 9571
rect 618 9540 622 9544
rect 628 9540 632 9544
rect 638 9540 642 9544
rect 618 9535 622 9539
rect 628 9535 632 9539
rect 638 9535 642 9539
rect 618 9530 622 9534
rect 628 9530 632 9534
rect 638 9530 642 9534
rect 618 9525 622 9529
rect 628 9525 632 9529
rect 638 9525 642 9529
rect 664 9540 668 9544
rect 674 9540 678 9544
rect 684 9540 688 9544
rect 664 9535 668 9539
rect 674 9535 678 9539
rect 684 9535 688 9539
rect 664 9530 668 9534
rect 674 9530 678 9534
rect 684 9530 688 9534
rect 664 9525 668 9529
rect 674 9525 678 9529
rect 684 9525 688 9529
rect 618 9514 622 9518
rect 628 9514 632 9518
rect 638 9514 642 9518
rect 618 9509 622 9513
rect 628 9509 632 9513
rect 638 9509 642 9513
rect 618 9504 622 9508
rect 628 9504 632 9508
rect 638 9504 642 9508
rect 618 9499 622 9503
rect 628 9499 632 9503
rect 638 9499 642 9503
rect 664 9514 668 9518
rect 674 9514 678 9518
rect 684 9514 688 9518
rect 664 9509 668 9513
rect 674 9509 678 9513
rect 684 9509 688 9513
rect 664 9504 668 9508
rect 674 9504 678 9508
rect 684 9504 688 9508
rect 664 9499 668 9503
rect 674 9499 678 9503
rect 684 9499 688 9503
rect 2824 9497 2830 9501
rect 3769 9497 3775 9501
rect 2812 9489 2818 9493
rect 3757 9489 3763 9493
rect 2800 9482 2806 9486
rect 3745 9482 3751 9486
rect 2788 9475 2794 9479
rect 3733 9475 3739 9479
rect 2776 9466 2782 9471
rect 3327 9467 3382 9471
rect 3721 9467 3727 9471
rect 2764 9459 2770 9463
rect 3635 9459 3690 9463
rect 3709 9460 3715 9464
rect 4484 9573 4488 9577
rect 4494 9573 4498 9577
rect 4504 9573 4508 9577
rect 4484 9568 4488 9572
rect 4494 9568 4498 9572
rect 4504 9568 4508 9572
rect 4484 9563 4488 9567
rect 4494 9563 4498 9567
rect 4504 9563 4508 9567
rect 4484 9558 4488 9562
rect 4494 9558 4498 9562
rect 4504 9558 4508 9562
rect 4530 9573 4534 9577
rect 4540 9573 4544 9577
rect 4550 9573 4554 9577
rect 4530 9568 4534 9572
rect 4540 9568 4544 9572
rect 4550 9568 4554 9572
rect 4530 9563 4534 9567
rect 4540 9563 4544 9567
rect 4550 9563 4554 9567
rect 4530 9558 4534 9562
rect 4540 9558 4544 9562
rect 4550 9558 4554 9562
rect 4484 9544 4488 9548
rect 4494 9544 4498 9548
rect 4504 9544 4508 9548
rect 4484 9539 4488 9543
rect 4494 9539 4498 9543
rect 4504 9539 4508 9543
rect 4484 9534 4488 9538
rect 4494 9534 4498 9538
rect 4504 9534 4508 9538
rect 4484 9529 4488 9533
rect 4494 9529 4498 9533
rect 4504 9529 4508 9533
rect 4530 9544 4534 9548
rect 4540 9544 4544 9548
rect 4550 9544 4554 9548
rect 4530 9539 4534 9543
rect 4540 9539 4544 9543
rect 4550 9539 4554 9543
rect 4530 9534 4534 9538
rect 4540 9534 4544 9538
rect 4550 9534 4554 9538
rect 4530 9529 4534 9533
rect 4540 9529 4544 9533
rect 4550 9529 4554 9533
rect 4484 9515 4488 9519
rect 4494 9515 4498 9519
rect 4504 9515 4508 9519
rect 4484 9510 4488 9514
rect 4494 9510 4498 9514
rect 4504 9510 4508 9514
rect 4484 9505 4488 9509
rect 4494 9505 4498 9509
rect 4504 9505 4508 9509
rect 4484 9500 4488 9504
rect 4494 9500 4498 9504
rect 4504 9500 4508 9504
rect 4530 9515 4534 9519
rect 4540 9515 4544 9519
rect 4550 9515 4554 9519
rect 4530 9510 4534 9514
rect 4540 9510 4544 9514
rect 4550 9510 4554 9514
rect 4530 9505 4534 9509
rect 4540 9505 4544 9509
rect 4550 9505 4554 9509
rect 4530 9500 4534 9504
rect 4540 9500 4544 9504
rect 4550 9500 4554 9504
rect 4484 9486 4488 9490
rect 4494 9486 4498 9490
rect 4504 9486 4508 9490
rect 4484 9481 4488 9485
rect 4494 9481 4498 9485
rect 4504 9481 4508 9485
rect 4484 9476 4488 9480
rect 4494 9476 4498 9480
rect 4504 9476 4508 9480
rect 4484 9471 4488 9475
rect 4494 9471 4498 9475
rect 4504 9471 4508 9475
rect 4530 9486 4534 9490
rect 4540 9486 4544 9490
rect 4550 9486 4554 9490
rect 4530 9481 4534 9485
rect 4540 9481 4544 9485
rect 4550 9481 4554 9485
rect 4530 9476 4534 9480
rect 4540 9476 4544 9480
rect 4550 9476 4554 9480
rect 4530 9471 4534 9475
rect 4540 9471 4544 9475
rect 4550 9471 4554 9475
rect 2836 9452 2842 9456
rect 3781 9452 3787 9456
rect 4484 9457 4488 9461
rect 4494 9457 4498 9461
rect 4504 9457 4508 9461
rect 4484 9452 4488 9456
rect 4494 9452 4498 9456
rect 4504 9452 4508 9456
rect 3040 9444 3053 9448
rect 3423 9444 3427 9448
rect 4484 9447 4488 9451
rect 4494 9447 4498 9451
rect 4504 9447 4508 9451
rect 4484 9442 4488 9446
rect 4494 9442 4498 9446
rect 4504 9442 4508 9446
rect 4530 9457 4534 9461
rect 4540 9457 4544 9461
rect 4550 9457 4554 9461
rect 4530 9452 4534 9456
rect 4540 9452 4544 9456
rect 4550 9452 4554 9456
rect 4530 9447 4534 9451
rect 4540 9447 4544 9451
rect 4550 9447 4554 9451
rect 4530 9442 4534 9446
rect 4540 9442 4544 9446
rect 4550 9442 4554 9446
rect 3021 9434 3026 9438
rect 3411 9434 3416 9438
rect 3757 9412 3763 9416
rect 3745 9404 3751 9408
rect 3733 9396 3739 9400
rect 3721 9388 3727 9392
rect 3709 9380 3715 9384
rect 2824 9347 2830 9351
rect 2857 9347 2861 9351
rect 2893 9347 2897 9351
rect 2960 9347 2964 9351
rect 2989 9347 2993 9351
rect 3025 9347 3029 9351
rect 3092 9347 3096 9351
rect 3121 9347 3125 9351
rect 3157 9347 3161 9351
rect 3224 9347 3228 9351
rect 3253 9347 3257 9351
rect 3289 9347 3293 9351
rect 3356 9347 3360 9351
rect 3769 9347 3775 9351
rect 3802 9347 3806 9351
rect 3838 9347 3842 9351
rect 3905 9347 3909 9351
rect 3934 9347 3938 9351
rect 3970 9347 3974 9351
rect 4037 9347 4041 9351
rect 4066 9347 4070 9351
rect 4102 9347 4106 9351
rect 4169 9347 4173 9351
rect 4198 9347 4202 9351
rect 4234 9347 4238 9351
rect 4301 9347 4305 9351
rect 2764 9340 2770 9344
rect 3709 9340 3715 9344
rect 2857 9333 2861 9337
rect 2907 9333 2911 9337
rect 2960 9333 2964 9337
rect 2989 9333 2993 9337
rect 3039 9333 3043 9337
rect 3092 9333 3096 9337
rect 3121 9333 3125 9337
rect 3171 9333 3175 9337
rect 3224 9333 3228 9337
rect 3253 9333 3257 9337
rect 3303 9333 3307 9337
rect 3356 9333 3360 9337
rect 3802 9333 3806 9337
rect 3852 9333 3856 9337
rect 3905 9333 3909 9337
rect 3934 9333 3938 9337
rect 3984 9333 3988 9337
rect 4037 9333 4041 9337
rect 4066 9333 4070 9337
rect 4116 9333 4120 9337
rect 4169 9333 4173 9337
rect 4198 9333 4202 9337
rect 4248 9333 4252 9337
rect 4301 9333 4305 9337
rect 618 9321 622 9325
rect 628 9321 632 9325
rect 638 9321 642 9325
rect 618 9316 622 9320
rect 628 9316 632 9320
rect 638 9316 642 9320
rect 618 9311 622 9315
rect 628 9311 632 9315
rect 638 9311 642 9315
rect 618 9306 622 9310
rect 628 9306 632 9310
rect 638 9306 642 9310
rect 664 9321 668 9325
rect 674 9321 678 9325
rect 684 9321 688 9325
rect 2880 9322 2884 9326
rect 664 9316 668 9320
rect 674 9316 678 9320
rect 684 9316 688 9320
rect 664 9311 668 9315
rect 674 9311 678 9315
rect 684 9311 688 9315
rect 2505 9314 2509 9318
rect 2541 9314 2545 9318
rect 2608 9314 2612 9318
rect 2824 9314 2830 9318
rect 2851 9313 2855 9317
rect 2864 9316 2868 9322
rect 2901 9316 2905 9322
rect 2914 9318 2918 9322
rect 2938 9322 2942 9326
rect 3012 9322 3016 9326
rect 2922 9316 2926 9322
rect 2959 9316 2963 9322
rect 2975 9318 2979 9322
rect 664 9306 668 9310
rect 674 9306 678 9310
rect 684 9306 688 9310
rect 2764 9307 2770 9311
rect 2505 9300 2509 9304
rect 2555 9300 2559 9304
rect 2608 9300 2612 9304
rect 2864 9303 2868 9307
rect 2880 9303 2884 9309
rect 2914 9309 2918 9313
rect 2901 9303 2905 9307
rect 2922 9303 2926 9307
rect 2938 9303 2942 9309
rect 2983 9313 2987 9317
rect 2996 9316 3000 9322
rect 3033 9316 3037 9322
rect 3046 9318 3050 9322
rect 3070 9322 3074 9326
rect 3144 9322 3148 9326
rect 3054 9316 3058 9322
rect 3091 9316 3095 9322
rect 3107 9318 3111 9322
rect 2959 9303 2963 9307
rect 2975 9303 2979 9307
rect 2996 9303 3000 9307
rect 3012 9303 3016 9309
rect 3046 9309 3050 9313
rect 3033 9303 3037 9307
rect 3054 9303 3058 9307
rect 3070 9303 3074 9309
rect 3115 9313 3119 9317
rect 3128 9316 3132 9322
rect 3165 9316 3169 9322
rect 3178 9318 3182 9322
rect 3202 9322 3206 9326
rect 3276 9322 3280 9326
rect 3186 9316 3190 9322
rect 3223 9316 3227 9322
rect 3239 9318 3243 9322
rect 3091 9303 3095 9307
rect 3107 9303 3111 9307
rect 3128 9303 3132 9307
rect 3144 9303 3148 9309
rect 3178 9309 3182 9313
rect 3165 9303 3169 9307
rect 3186 9303 3190 9307
rect 3202 9303 3206 9309
rect 3247 9313 3251 9317
rect 3260 9316 3264 9322
rect 3297 9316 3301 9322
rect 3310 9318 3314 9322
rect 3334 9322 3338 9326
rect 3825 9322 3829 9326
rect 3318 9316 3322 9322
rect 3355 9316 3359 9322
rect 3371 9318 3375 9322
rect 3450 9314 3454 9318
rect 3486 9314 3490 9318
rect 3553 9314 3557 9318
rect 3769 9314 3775 9318
rect 3223 9303 3227 9307
rect 3239 9303 3243 9307
rect 3260 9303 3264 9307
rect 3276 9303 3280 9309
rect 3310 9309 3314 9313
rect 3297 9303 3301 9307
rect 2528 9289 2532 9293
rect 2490 9280 2494 9284
rect 2512 9283 2516 9289
rect 2549 9283 2553 9289
rect 2562 9285 2566 9289
rect 2586 9289 2590 9293
rect 2570 9283 2574 9289
rect 2607 9283 2611 9289
rect 2623 9283 2627 9289
rect 2857 9292 2861 9296
rect 2894 9290 2898 9294
rect 2914 9290 2918 9294
rect 2958 9290 2962 9294
rect 2989 9292 2993 9296
rect 3026 9290 3030 9294
rect 3046 9290 3050 9294
rect 3090 9290 3094 9294
rect 3121 9292 3125 9296
rect 3158 9290 3162 9294
rect 3178 9290 3182 9294
rect 3222 9290 3226 9294
rect 3239 9295 3243 9299
rect 3318 9303 3322 9307
rect 3334 9303 3338 9309
rect 3796 9313 3800 9317
rect 3809 9316 3813 9322
rect 3846 9316 3850 9322
rect 3859 9318 3863 9322
rect 3883 9322 3887 9326
rect 3957 9322 3961 9326
rect 3867 9316 3871 9322
rect 3904 9316 3908 9322
rect 3920 9318 3924 9322
rect 3709 9307 3715 9311
rect 3355 9303 3359 9307
rect 3371 9303 3375 9307
rect 3253 9292 3257 9296
rect 3290 9290 3294 9294
rect 3310 9290 3314 9294
rect 3354 9290 3358 9294
rect 3371 9295 3375 9299
rect 3450 9300 3454 9304
rect 3500 9300 3504 9304
rect 3553 9300 3557 9304
rect 3809 9303 3813 9307
rect 3825 9303 3829 9309
rect 3859 9309 3863 9313
rect 3846 9303 3850 9307
rect 3867 9303 3871 9307
rect 3883 9303 3887 9309
rect 3928 9313 3932 9317
rect 3941 9316 3945 9322
rect 3978 9316 3982 9322
rect 3991 9318 3995 9322
rect 4015 9322 4019 9326
rect 4089 9322 4093 9326
rect 3999 9316 4003 9322
rect 4036 9316 4040 9322
rect 4052 9318 4056 9322
rect 3904 9303 3908 9307
rect 3920 9303 3924 9307
rect 3941 9303 3945 9307
rect 3957 9303 3961 9309
rect 3991 9309 3995 9313
rect 3978 9303 3982 9307
rect 3999 9303 4003 9307
rect 4015 9303 4019 9309
rect 4060 9313 4064 9317
rect 4073 9316 4077 9322
rect 4110 9316 4114 9322
rect 4123 9318 4127 9322
rect 4147 9322 4151 9326
rect 4221 9322 4225 9326
rect 4131 9316 4135 9322
rect 4168 9316 4172 9322
rect 4184 9318 4188 9322
rect 4036 9303 4040 9307
rect 4052 9303 4056 9307
rect 4073 9303 4077 9307
rect 4089 9303 4093 9309
rect 4123 9309 4127 9313
rect 4110 9303 4114 9307
rect 4131 9303 4135 9307
rect 4147 9303 4151 9309
rect 4192 9313 4196 9317
rect 4205 9316 4209 9322
rect 4242 9316 4246 9322
rect 4255 9318 4259 9322
rect 4279 9322 4283 9326
rect 4263 9316 4267 9322
rect 4300 9316 4304 9322
rect 4316 9318 4320 9322
rect 4168 9303 4172 9307
rect 4184 9303 4188 9307
rect 4205 9303 4209 9307
rect 4221 9303 4225 9309
rect 4255 9309 4259 9313
rect 4242 9303 4246 9307
rect 3473 9289 3477 9293
rect 2776 9283 2782 9287
rect 2512 9270 2516 9274
rect 2528 9270 2532 9276
rect 2562 9276 2566 9280
rect 2549 9270 2553 9274
rect 2570 9270 2574 9274
rect 2586 9270 2590 9276
rect 3435 9280 3439 9284
rect 3457 9283 3461 9289
rect 3494 9283 3498 9289
rect 3507 9285 3511 9289
rect 3531 9289 3535 9293
rect 3515 9283 3519 9289
rect 3552 9283 3556 9289
rect 3568 9283 3572 9289
rect 3802 9292 3806 9296
rect 3839 9290 3843 9294
rect 3859 9290 3863 9294
rect 3903 9290 3907 9294
rect 3934 9292 3938 9296
rect 3971 9290 3975 9294
rect 3991 9290 3995 9294
rect 4035 9290 4039 9294
rect 4066 9292 4070 9296
rect 4103 9290 4107 9294
rect 4123 9290 4127 9294
rect 4167 9290 4171 9294
rect 4184 9295 4188 9299
rect 4263 9303 4267 9307
rect 4279 9303 4283 9309
rect 4300 9303 4304 9307
rect 4316 9303 4320 9307
rect 4198 9292 4202 9296
rect 4235 9290 4239 9294
rect 4255 9290 4259 9294
rect 4299 9290 4303 9294
rect 4316 9295 4320 9299
rect 3721 9283 3727 9287
rect 2812 9276 2818 9280
rect 2857 9276 2861 9280
rect 2908 9276 2912 9280
rect 2958 9276 2962 9280
rect 2989 9276 2993 9280
rect 3040 9276 3044 9280
rect 3090 9276 3094 9280
rect 3121 9276 3125 9280
rect 3172 9276 3176 9280
rect 3222 9276 3226 9280
rect 3253 9276 3257 9280
rect 3304 9276 3308 9280
rect 3354 9276 3358 9280
rect 2607 9270 2611 9274
rect 2623 9270 2627 9274
rect 3457 9270 3461 9274
rect 3473 9270 3477 9276
rect 3507 9276 3511 9280
rect 3494 9270 3498 9274
rect 2505 9259 2509 9263
rect 2542 9257 2546 9261
rect 2562 9257 2566 9261
rect 2606 9257 2610 9261
rect 2764 9263 2770 9267
rect 2855 9263 2859 9267
rect 2889 9263 2893 9267
rect 2906 9263 2910 9267
rect 2962 9263 2966 9267
rect 2979 9263 2983 9267
rect 3007 9263 3011 9267
rect 3515 9270 3519 9274
rect 3531 9270 3535 9276
rect 3757 9276 3763 9280
rect 3802 9276 3806 9280
rect 3853 9276 3857 9280
rect 3903 9276 3907 9280
rect 3934 9276 3938 9280
rect 3985 9276 3989 9280
rect 4035 9276 4039 9280
rect 4066 9276 4070 9280
rect 4117 9276 4121 9280
rect 4167 9276 4171 9280
rect 4198 9276 4202 9280
rect 4249 9276 4253 9280
rect 4299 9276 4303 9280
rect 3552 9270 3556 9274
rect 3568 9270 3572 9274
rect 2800 9256 2806 9260
rect 2882 9256 2886 9260
rect 2913 9256 2917 9260
rect 2935 9256 2939 9260
rect 3000 9256 3004 9260
rect 2776 9250 2782 9254
rect 2505 9243 2509 9247
rect 2556 9243 2560 9247
rect 2606 9243 2610 9247
rect 2812 9243 2818 9247
rect 2856 9246 2860 9250
rect 2881 9249 2885 9253
rect 2888 9246 2892 9250
rect 2906 9246 2910 9250
rect 2928 9249 2932 9253
rect 2953 9249 2957 9253
rect 2963 9246 2967 9250
rect 2979 9246 2983 9250
rect 2999 9249 3003 9253
rect 3006 9246 3010 9250
rect 3070 9256 3074 9260
rect 2623 9236 2627 9240
rect 2490 9227 2494 9231
rect 2615 9229 2619 9233
rect 2639 9229 2643 9233
rect 2498 9220 2502 9224
rect 2639 9220 2643 9224
rect 2883 9230 2887 9234
rect 2903 9227 2907 9231
rect 2922 9231 2926 9235
rect 3024 9242 3028 9246
rect 3039 9242 3043 9246
rect 2941 9230 2945 9234
rect 2960 9230 2964 9234
rect 2973 9229 2977 9233
rect 2995 9230 2999 9234
rect 3003 9229 3007 9233
rect 3015 9229 3019 9233
rect 2856 9216 2860 9220
rect 2888 9216 2892 9220
rect 2906 9216 2910 9220
rect 2963 9216 2967 9220
rect 2978 9216 2982 9220
rect 3006 9216 3010 9220
rect 2505 9212 2509 9216
rect 2572 9212 2576 9216
rect 2608 9212 2612 9216
rect 2824 9212 2830 9216
rect 2870 9212 2874 9216
rect 2913 9211 2917 9215
rect 2935 9212 2942 9216
rect 2985 9211 2989 9215
rect 2764 9205 2770 9209
rect 2505 9198 2509 9202
rect 2558 9198 2562 9202
rect 2608 9198 2612 9202
rect 2788 9204 2794 9208
rect 2870 9204 2874 9208
rect 2929 9204 2933 9208
rect 2954 9204 2958 9208
rect 2985 9204 2989 9208
rect 3078 9234 3082 9242
rect 3151 9256 3155 9260
rect 3105 9242 3109 9246
rect 3120 9242 3124 9246
rect 3101 9234 3105 9238
rect 3047 9228 3051 9232
rect 3060 9220 3064 9224
rect 3159 9234 3163 9242
rect 3315 9250 3328 9258
rect 3411 9250 3416 9258
rect 3450 9259 3454 9263
rect 3487 9257 3491 9261
rect 3507 9257 3511 9261
rect 3551 9257 3555 9261
rect 3709 9263 3715 9267
rect 3800 9263 3804 9267
rect 3834 9263 3838 9267
rect 3851 9263 3855 9267
rect 3907 9263 3911 9267
rect 3924 9263 3928 9267
rect 3952 9263 3956 9267
rect 3745 9256 3751 9260
rect 3827 9256 3831 9260
rect 3858 9256 3862 9260
rect 3880 9256 3884 9260
rect 3945 9256 3949 9260
rect 3721 9250 3727 9254
rect 3361 9241 3365 9245
rect 3423 9241 3427 9245
rect 3450 9243 3454 9247
rect 3501 9243 3505 9247
rect 3551 9243 3555 9247
rect 3757 9243 3763 9247
rect 3801 9246 3805 9250
rect 3826 9249 3830 9253
rect 3833 9246 3837 9250
rect 3851 9246 3855 9250
rect 3873 9249 3877 9253
rect 3898 9249 3902 9253
rect 3908 9246 3912 9250
rect 3924 9246 3928 9250
rect 3944 9249 3948 9253
rect 3951 9246 3955 9250
rect 4015 9256 4019 9260
rect 3186 9234 3190 9238
rect 3568 9236 3572 9240
rect 3128 9228 3132 9232
rect 3435 9227 3439 9231
rect 3560 9229 3564 9233
rect 3584 9229 3588 9233
rect 3793 9229 3797 9233
rect 3141 9220 3145 9224
rect 3443 9220 3447 9224
rect 3584 9220 3588 9224
rect 3828 9230 3832 9234
rect 3848 9227 3852 9231
rect 3867 9231 3871 9235
rect 3969 9242 3973 9246
rect 3984 9242 3988 9246
rect 3886 9230 3890 9234
rect 3905 9230 3909 9234
rect 3918 9229 3922 9233
rect 3940 9230 3944 9234
rect 3948 9229 3952 9233
rect 3960 9229 3964 9233
rect 3801 9216 3805 9220
rect 3833 9216 3837 9220
rect 3851 9216 3855 9220
rect 3908 9216 3912 9220
rect 3923 9216 3927 9220
rect 3951 9216 3955 9220
rect 3450 9212 3454 9216
rect 3517 9212 3521 9216
rect 3553 9212 3557 9216
rect 3769 9212 3775 9216
rect 3815 9212 3819 9216
rect 3858 9211 3862 9215
rect 3880 9212 3887 9216
rect 3930 9211 3934 9215
rect 3709 9205 3715 9209
rect 2776 9197 2782 9201
rect 2856 9197 2860 9201
rect 2870 9197 2874 9201
rect 2888 9197 2892 9201
rect 2906 9197 2910 9201
rect 2929 9197 2933 9201
rect 2963 9197 2967 9201
rect 2978 9197 2982 9201
rect 3006 9197 3010 9201
rect 2527 9187 2531 9191
rect 2490 9181 2494 9187
rect 2506 9181 2510 9187
rect 2543 9181 2547 9187
rect 2551 9183 2555 9187
rect 2585 9187 2589 9191
rect 2788 9190 2794 9194
rect 2870 9190 2874 9194
rect 2929 9190 2933 9194
rect 2954 9190 2958 9194
rect 2985 9190 2989 9194
rect 2564 9181 2568 9187
rect 2601 9181 2605 9187
rect 2870 9182 2874 9186
rect 2913 9183 2917 9187
rect 2935 9182 2942 9186
rect 2985 9183 2989 9187
rect 2623 9178 2627 9182
rect 2856 9178 2860 9182
rect 2888 9178 2892 9182
rect 2906 9178 2910 9182
rect 2963 9178 2967 9182
rect 2978 9178 2982 9182
rect 3006 9178 3010 9182
rect 2490 9168 2494 9172
rect 2506 9168 2510 9172
rect 2551 9174 2555 9178
rect 2527 9168 2531 9174
rect 2543 9168 2547 9172
rect 2564 9168 2568 9172
rect 2585 9168 2589 9174
rect 2601 9168 2605 9172
rect 2851 9166 2855 9170
rect 2507 9155 2511 9159
rect 2551 9155 2555 9159
rect 2571 9155 2575 9159
rect 2608 9157 2612 9161
rect 2883 9164 2887 9168
rect 2903 9167 2907 9171
rect 2922 9163 2926 9167
rect 2941 9164 2945 9168
rect 2960 9164 2964 9168
rect 2973 9165 2977 9169
rect 3070 9180 3074 9184
rect 3450 9198 3454 9202
rect 3503 9198 3507 9202
rect 3553 9198 3557 9202
rect 3733 9204 3739 9208
rect 3815 9204 3819 9208
rect 3874 9204 3878 9208
rect 3899 9204 3903 9208
rect 3930 9204 3934 9208
rect 4023 9234 4027 9242
rect 4096 9256 4100 9260
rect 4050 9242 4054 9246
rect 4065 9242 4069 9246
rect 4046 9234 4050 9238
rect 3992 9228 3996 9232
rect 4005 9220 4009 9224
rect 4104 9234 4108 9242
rect 4131 9234 4135 9238
rect 4073 9228 4077 9232
rect 4086 9220 4090 9224
rect 3721 9197 3727 9201
rect 3801 9197 3805 9201
rect 3815 9197 3819 9201
rect 3833 9197 3837 9201
rect 3851 9197 3855 9201
rect 3874 9197 3878 9201
rect 3908 9197 3912 9201
rect 3923 9197 3927 9201
rect 3951 9197 3955 9201
rect 3472 9187 3476 9191
rect 3151 9180 3155 9184
rect 3435 9181 3439 9187
rect 3451 9181 3455 9187
rect 3488 9181 3492 9187
rect 3496 9183 3500 9187
rect 3530 9187 3534 9191
rect 3733 9190 3739 9194
rect 3815 9190 3819 9194
rect 3874 9190 3878 9194
rect 3899 9190 3903 9194
rect 3930 9190 3934 9194
rect 3509 9181 3513 9187
rect 3546 9181 3550 9187
rect 3815 9182 3819 9186
rect 3858 9183 3862 9187
rect 3880 9182 3887 9186
rect 3930 9183 3934 9187
rect 3568 9178 3572 9182
rect 3801 9178 3805 9182
rect 3833 9178 3837 9182
rect 3851 9178 3855 9182
rect 3908 9178 3912 9182
rect 3923 9178 3927 9182
rect 3951 9178 3955 9182
rect 2995 9164 2999 9168
rect 3003 9165 3007 9169
rect 3015 9165 3019 9169
rect 3050 9165 3054 9169
rect 3078 9164 3082 9168
rect 3130 9165 3134 9169
rect 3435 9168 3439 9172
rect 3451 9168 3455 9172
rect 3496 9174 3500 9178
rect 3472 9168 3476 9174
rect 3488 9168 3492 9172
rect 3159 9164 3163 9168
rect 3509 9168 3513 9172
rect 3530 9168 3534 9174
rect 3546 9168 3550 9172
rect 3796 9166 3800 9170
rect 2776 9148 2782 9152
rect 2856 9148 2860 9152
rect 2881 9145 2885 9149
rect 2888 9148 2892 9152
rect 2906 9148 2910 9152
rect 2928 9145 2932 9149
rect 2953 9145 2957 9149
rect 2963 9148 2967 9152
rect 2979 9148 2983 9152
rect 2999 9145 3003 9149
rect 3006 9148 3010 9152
rect 2507 9141 2511 9145
rect 2557 9141 2561 9145
rect 2608 9141 2612 9145
rect 2812 9141 2818 9145
rect 2866 9138 2870 9142
rect 2882 9138 2886 9142
rect 2913 9138 2917 9142
rect 2935 9138 2939 9142
rect 3000 9138 3004 9142
rect 3060 9144 3064 9148
rect 3452 9155 3456 9159
rect 3496 9155 3500 9159
rect 3516 9155 3520 9159
rect 3553 9157 3557 9161
rect 3828 9164 3832 9168
rect 3848 9167 3852 9171
rect 3867 9163 3871 9167
rect 3886 9164 3890 9168
rect 3905 9164 3909 9168
rect 3918 9165 3922 9169
rect 4015 9180 4019 9184
rect 4096 9180 4100 9184
rect 3940 9164 3944 9168
rect 3948 9165 3952 9169
rect 3960 9165 3964 9169
rect 3995 9165 3999 9169
rect 4023 9164 4027 9168
rect 4075 9165 4079 9169
rect 4104 9164 4108 9168
rect 3721 9148 3727 9152
rect 3801 9148 3805 9152
rect 3141 9144 3145 9148
rect 3826 9145 3830 9149
rect 3833 9148 3837 9152
rect 3851 9148 3855 9152
rect 3873 9145 3877 9149
rect 3898 9145 3902 9149
rect 3908 9148 3912 9152
rect 3924 9148 3928 9152
rect 3944 9145 3948 9149
rect 3951 9148 3955 9152
rect 3452 9141 3456 9145
rect 3502 9141 3506 9145
rect 3553 9141 3557 9145
rect 3757 9141 3763 9145
rect 3811 9138 3815 9142
rect 3827 9138 3831 9142
rect 3858 9138 3862 9142
rect 3880 9138 3884 9142
rect 3945 9138 3949 9142
rect 4005 9144 4009 9148
rect 4086 9144 4090 9148
rect 2764 9131 2770 9135
rect 2855 9131 2859 9135
rect 2889 9131 2893 9135
rect 2906 9131 2910 9135
rect 2962 9131 2966 9135
rect 2979 9131 2983 9135
rect 3007 9131 3011 9135
rect 3709 9131 3715 9135
rect 3800 9131 3804 9135
rect 3834 9131 3838 9135
rect 3851 9131 3855 9135
rect 3907 9131 3911 9135
rect 3924 9131 3928 9135
rect 3952 9131 3956 9135
rect 2800 9124 2806 9128
rect 2866 9124 2870 9128
rect 2882 9124 2886 9128
rect 2913 9124 2917 9128
rect 2935 9124 2939 9128
rect 3000 9124 3004 9128
rect 3070 9124 3074 9128
rect 2856 9114 2860 9118
rect 2881 9117 2885 9121
rect 2888 9114 2892 9118
rect 2906 9114 2910 9118
rect 2928 9117 2932 9121
rect 2953 9117 2957 9121
rect 2963 9114 2967 9118
rect 2979 9114 2983 9118
rect 2999 9117 3003 9121
rect 3006 9114 3010 9118
rect 2850 9097 2854 9101
rect 2883 9098 2887 9102
rect 2903 9095 2907 9099
rect 2922 9099 2926 9103
rect 2941 9098 2945 9102
rect 2960 9098 2964 9102
rect 2973 9097 2977 9101
rect 2995 9098 2999 9102
rect 3003 9097 3007 9101
rect 3015 9097 3019 9101
rect 3078 9102 3082 9110
rect 3175 9124 3179 9128
rect 3129 9110 3133 9114
rect 3144 9110 3148 9114
rect 3361 9120 3365 9124
rect 3745 9124 3751 9128
rect 3811 9124 3815 9128
rect 3827 9124 3831 9128
rect 3858 9124 3862 9128
rect 3880 9124 3884 9128
rect 3945 9124 3949 9128
rect 4015 9124 4019 9128
rect 3047 9096 3051 9100
rect 3101 9101 3105 9105
rect 2856 9084 2860 9088
rect 2888 9084 2892 9088
rect 2906 9084 2910 9088
rect 2963 9084 2967 9088
rect 2978 9084 2982 9088
rect 3006 9084 3010 9088
rect 2870 9080 2874 9084
rect 2913 9079 2917 9083
rect 2935 9080 2942 9084
rect 2985 9079 2989 9083
rect 2788 9072 2794 9076
rect 2870 9072 2874 9076
rect 2929 9072 2933 9076
rect 2954 9072 2958 9076
rect 2985 9072 2989 9076
rect 3060 9088 3064 9092
rect 3183 9102 3187 9110
rect 3801 9114 3805 9118
rect 3826 9117 3830 9121
rect 3833 9114 3837 9118
rect 3851 9114 3855 9118
rect 3873 9117 3877 9121
rect 3898 9117 3902 9121
rect 3908 9114 3912 9118
rect 3924 9114 3928 9118
rect 3944 9117 3948 9121
rect 3951 9114 3955 9118
rect 3204 9102 3208 9106
rect 3668 9102 3672 9106
rect 3152 9096 3156 9100
rect 3165 9088 3169 9092
rect 3406 9095 3410 9099
rect 3360 9081 3364 9085
rect 3375 9081 3379 9085
rect 3383 9073 3387 9077
rect 3414 9073 3418 9081
rect 3795 9097 3799 9101
rect 2776 9065 2782 9069
rect 2856 9065 2860 9069
rect 2870 9065 2874 9069
rect 2888 9065 2892 9069
rect 2906 9065 2910 9069
rect 2929 9065 2933 9069
rect 2963 9065 2967 9069
rect 2978 9065 2982 9069
rect 3006 9065 3010 9069
rect 2788 9058 2794 9062
rect 2870 9058 2874 9062
rect 2929 9058 2933 9062
rect 2954 9058 2958 9062
rect 2985 9058 2989 9062
rect 2870 9050 2874 9054
rect 2913 9051 2917 9055
rect 2935 9050 2942 9054
rect 2985 9051 2989 9055
rect 2856 9046 2860 9050
rect 2888 9046 2892 9050
rect 2906 9046 2910 9050
rect 2963 9046 2967 9050
rect 2978 9046 2982 9050
rect 3006 9046 3010 9050
rect 3070 9049 3074 9053
rect 3175 9049 3179 9053
rect 2851 9034 2855 9038
rect 2883 9032 2887 9036
rect 2903 9035 2907 9039
rect 2922 9031 2926 9035
rect 2941 9032 2945 9036
rect 2960 9032 2964 9036
rect 2973 9033 2977 9037
rect 2995 9032 2999 9036
rect 3003 9033 3007 9037
rect 3015 9033 3019 9037
rect 3049 9034 3053 9038
rect 3078 9033 3082 9037
rect 3155 9034 3159 9038
rect 3183 9033 3187 9037
rect 3396 9059 3400 9063
rect 3828 9098 3832 9102
rect 3848 9095 3852 9099
rect 3867 9099 3871 9103
rect 3886 9098 3890 9102
rect 3905 9098 3909 9102
rect 3918 9097 3922 9101
rect 3940 9098 3944 9102
rect 3948 9097 3952 9101
rect 3960 9097 3964 9101
rect 4023 9102 4027 9110
rect 4120 9124 4124 9128
rect 4074 9110 4078 9114
rect 4089 9110 4093 9114
rect 3992 9096 3996 9100
rect 4046 9101 4050 9105
rect 3801 9084 3805 9088
rect 3833 9084 3837 9088
rect 3851 9084 3855 9088
rect 3908 9084 3912 9088
rect 3923 9084 3927 9088
rect 3951 9084 3955 9088
rect 3815 9080 3819 9084
rect 3858 9079 3862 9083
rect 3880 9080 3887 9084
rect 3930 9079 3934 9083
rect 3733 9072 3739 9076
rect 3815 9072 3819 9076
rect 3874 9072 3878 9076
rect 3899 9072 3903 9076
rect 3930 9072 3934 9076
rect 4005 9088 4009 9092
rect 4128 9102 4132 9110
rect 4149 9102 4153 9106
rect 4097 9096 4101 9100
rect 4110 9088 4114 9092
rect 3721 9065 3727 9069
rect 3801 9065 3805 9069
rect 3815 9065 3819 9069
rect 3833 9065 3837 9069
rect 3851 9065 3855 9069
rect 3874 9065 3878 9069
rect 3908 9065 3912 9069
rect 3923 9065 3927 9069
rect 3951 9065 3955 9069
rect 3593 9053 3597 9057
rect 3733 9058 3739 9062
rect 3815 9058 3819 9062
rect 3874 9058 3878 9062
rect 3899 9058 3903 9062
rect 3930 9058 3934 9062
rect 3815 9050 3819 9054
rect 3858 9051 3862 9055
rect 3880 9050 3887 9054
rect 3930 9051 3934 9055
rect 3626 9045 3630 9049
rect 3745 9045 3751 9049
rect 3801 9046 3805 9050
rect 3833 9046 3837 9050
rect 3851 9046 3855 9050
rect 3908 9046 3912 9050
rect 3923 9046 3927 9050
rect 3951 9046 3955 9050
rect 4015 9049 4019 9053
rect 4484 9056 4488 9060
rect 4494 9056 4498 9060
rect 4504 9056 4508 9060
rect 4120 9049 4124 9053
rect 4484 9051 4488 9055
rect 4494 9051 4498 9055
rect 4504 9051 4508 9055
rect 4484 9046 4488 9050
rect 4494 9046 4498 9050
rect 4504 9046 4508 9050
rect 3668 9033 3672 9037
rect 3709 9033 3715 9037
rect 3796 9034 3800 9038
rect 3721 9026 3727 9030
rect 3660 9022 3665 9026
rect 2856 9016 2860 9020
rect 618 9012 622 9016
rect 628 9012 632 9016
rect 638 9012 642 9016
rect 618 9007 622 9011
rect 628 9007 632 9011
rect 638 9007 642 9011
rect 618 9002 622 9006
rect 628 9002 632 9006
rect 638 9002 642 9006
rect 618 8997 622 9001
rect 628 8997 632 9001
rect 638 8997 642 9001
rect 664 9012 668 9016
rect 674 9012 678 9016
rect 684 9012 688 9016
rect 2881 9013 2885 9017
rect 2888 9016 2892 9020
rect 2906 9016 2910 9020
rect 2928 9013 2932 9017
rect 2953 9013 2957 9017
rect 2963 9016 2967 9020
rect 2979 9016 2983 9020
rect 2999 9013 3003 9017
rect 3006 9016 3010 9020
rect 664 9007 668 9011
rect 674 9007 678 9011
rect 684 9007 688 9011
rect 2800 9006 2806 9010
rect 2882 9006 2886 9010
rect 2913 9006 2917 9010
rect 2935 9006 2939 9010
rect 3000 9006 3004 9010
rect 664 9002 668 9006
rect 674 9002 678 9006
rect 684 9002 688 9006
rect 3060 9013 3064 9017
rect 3165 9013 3169 9017
rect 3406 9015 3410 9019
rect 3676 9017 3680 9021
rect 3781 9017 3787 9021
rect 3828 9032 3832 9036
rect 3848 9035 3852 9039
rect 3867 9031 3871 9035
rect 3886 9032 3890 9036
rect 3905 9032 3909 9036
rect 3918 9033 3922 9037
rect 3940 9032 3944 9036
rect 3948 9033 3952 9037
rect 3960 9033 3964 9037
rect 3994 9034 3998 9038
rect 4023 9033 4027 9037
rect 4100 9034 4104 9038
rect 4484 9041 4488 9045
rect 4494 9041 4498 9045
rect 4504 9041 4508 9045
rect 4530 9056 4534 9060
rect 4540 9056 4544 9060
rect 4550 9056 4554 9060
rect 4530 9051 4534 9055
rect 4540 9051 4544 9055
rect 4550 9051 4554 9055
rect 4530 9046 4534 9050
rect 4540 9046 4544 9050
rect 4550 9046 4554 9050
rect 4530 9041 4534 9045
rect 4540 9041 4544 9045
rect 4550 9041 4554 9045
rect 4128 9033 4132 9037
rect 3801 9016 3805 9020
rect 3826 9013 3830 9017
rect 3833 9016 3837 9020
rect 3851 9016 3855 9020
rect 3873 9013 3877 9017
rect 3898 9013 3902 9017
rect 3908 9016 3912 9020
rect 3924 9016 3928 9020
rect 3944 9013 3948 9017
rect 3951 9016 3955 9020
rect 3593 9008 3598 9012
rect 3733 9008 3739 9012
rect 664 8997 668 9001
rect 674 8997 678 9001
rect 684 8997 688 9001
rect 2764 8999 2770 9003
rect 2855 8999 2859 9003
rect 2889 8999 2893 9003
rect 2906 8999 2910 9003
rect 2962 8999 2966 9003
rect 2979 8999 2983 9003
rect 3007 8999 3011 9003
rect 3326 9000 3330 9004
rect 3745 9006 3751 9010
rect 3827 9006 3831 9010
rect 3858 9006 3862 9010
rect 3880 9006 3884 9010
rect 3945 9006 3949 9010
rect 4005 9013 4009 9017
rect 4110 9013 4114 9017
rect 3414 8999 3418 9003
rect 3709 8999 3715 9003
rect 3800 8999 3804 9003
rect 3834 8999 3838 9003
rect 3851 8999 3855 9003
rect 3907 8999 3911 9003
rect 3924 8999 3928 9003
rect 3952 8999 3956 9003
rect 2800 8992 2806 8996
rect 2882 8992 2886 8996
rect 2913 8992 2917 8996
rect 2935 8992 2939 8996
rect 3000 8992 3004 8996
rect 3070 8992 3074 8996
rect 2856 8982 2860 8986
rect 2881 8985 2885 8989
rect 2888 8982 2892 8986
rect 2906 8982 2910 8986
rect 2928 8985 2932 8989
rect 2953 8985 2957 8989
rect 2963 8982 2967 8986
rect 2979 8982 2983 8986
rect 2999 8985 3003 8989
rect 3006 8982 3010 8986
rect 2850 8965 2854 8969
rect 2883 8966 2887 8970
rect 2903 8963 2907 8967
rect 2922 8967 2926 8971
rect 2941 8966 2945 8970
rect 2960 8966 2964 8970
rect 2973 8965 2977 8969
rect 2995 8966 2999 8970
rect 3003 8965 3007 8969
rect 3015 8965 3019 8969
rect 3078 8970 3082 8978
rect 3151 8992 3155 8996
rect 3105 8978 3109 8982
rect 3120 8978 3124 8982
rect 3101 8970 3105 8974
rect 3047 8964 3051 8968
rect 2856 8952 2860 8956
rect 2888 8952 2892 8956
rect 2906 8952 2910 8956
rect 2963 8952 2967 8956
rect 2978 8952 2982 8956
rect 3006 8952 3010 8956
rect 2870 8948 2874 8952
rect 2913 8947 2917 8951
rect 2935 8948 2942 8952
rect 2985 8947 2989 8951
rect 2788 8940 2794 8944
rect 2870 8940 2874 8944
rect 2929 8940 2933 8944
rect 2954 8940 2958 8944
rect 2985 8940 2989 8944
rect 3060 8956 3064 8960
rect 3159 8970 3163 8978
rect 3241 8992 3245 8996
rect 3195 8978 3199 8982
rect 3210 8978 3214 8982
rect 3183 8970 3187 8974
rect 3128 8964 3132 8968
rect 3217 8972 3221 8976
rect 3249 8970 3253 8978
rect 3745 8992 3751 8996
rect 3827 8992 3831 8996
rect 3858 8992 3862 8996
rect 3880 8992 3884 8996
rect 3945 8992 3949 8996
rect 4015 8992 4019 8996
rect 3396 8979 3400 8983
rect 3801 8982 3805 8986
rect 3826 8985 3830 8989
rect 3833 8982 3837 8986
rect 3851 8982 3855 8986
rect 3873 8985 3877 8989
rect 3898 8985 3902 8989
rect 3908 8982 3912 8986
rect 3924 8982 3928 8986
rect 3944 8985 3948 8989
rect 3951 8982 3955 8986
rect 3141 8956 3145 8960
rect 3284 8969 3288 8973
rect 3668 8972 3672 8976
rect 3231 8956 3235 8960
rect 3406 8965 3410 8969
rect 3338 8951 3342 8955
rect 3353 8951 3357 8955
rect 3360 8951 3364 8955
rect 3375 8951 3379 8955
rect 3383 8943 3387 8947
rect 3414 8943 3418 8951
rect 3795 8965 3799 8969
rect 2776 8933 2782 8937
rect 2856 8933 2860 8937
rect 2870 8933 2874 8937
rect 2888 8933 2892 8937
rect 2906 8933 2910 8937
rect 2929 8933 2933 8937
rect 2963 8933 2967 8937
rect 2978 8933 2982 8937
rect 3006 8933 3010 8937
rect 2788 8926 2794 8930
rect 2870 8926 2874 8930
rect 2929 8926 2933 8930
rect 2954 8926 2958 8930
rect 2985 8926 2989 8930
rect 2870 8918 2874 8922
rect 2913 8919 2917 8923
rect 2935 8918 2942 8922
rect 2985 8919 2989 8923
rect 2856 8914 2860 8918
rect 2888 8914 2892 8918
rect 2906 8914 2910 8918
rect 2963 8914 2967 8918
rect 2978 8914 2982 8918
rect 3006 8914 3010 8918
rect 2851 8902 2855 8906
rect 2883 8900 2887 8904
rect 2903 8903 2907 8907
rect 2922 8899 2926 8903
rect 2941 8900 2945 8904
rect 2960 8900 2964 8904
rect 2973 8901 2977 8905
rect 3070 8914 3074 8918
rect 3151 8914 3155 8918
rect 3241 8914 3245 8918
rect 2995 8900 2999 8904
rect 3003 8901 3007 8905
rect 3015 8901 3019 8905
rect 3050 8899 3054 8903
rect 3078 8898 3082 8902
rect 3130 8899 3134 8903
rect 3159 8898 3163 8902
rect 3214 8899 3218 8903
rect 3249 8898 3253 8902
rect 3396 8929 3400 8933
rect 3828 8966 3832 8970
rect 3848 8963 3852 8967
rect 3867 8967 3871 8971
rect 3886 8966 3890 8970
rect 3905 8966 3909 8970
rect 3918 8965 3922 8969
rect 3940 8966 3944 8970
rect 3948 8965 3952 8969
rect 3960 8965 3964 8969
rect 4023 8970 4027 8978
rect 4096 8992 4100 8996
rect 4050 8978 4054 8982
rect 4065 8978 4069 8982
rect 4046 8970 4050 8974
rect 3992 8964 3996 8968
rect 3801 8952 3805 8956
rect 3833 8952 3837 8956
rect 3851 8952 3855 8956
rect 3908 8952 3912 8956
rect 3923 8952 3927 8956
rect 3951 8952 3955 8956
rect 3815 8948 3819 8952
rect 3858 8947 3862 8951
rect 3880 8948 3887 8952
rect 3930 8947 3934 8951
rect 3733 8940 3739 8944
rect 3815 8940 3819 8944
rect 3874 8940 3878 8944
rect 3899 8940 3903 8944
rect 3930 8940 3934 8944
rect 4005 8956 4009 8960
rect 4104 8970 4108 8978
rect 4186 8992 4190 8996
rect 4140 8978 4144 8982
rect 4155 8978 4159 8982
rect 4128 8970 4132 8974
rect 4073 8964 4077 8968
rect 4162 8972 4166 8976
rect 4194 8970 4198 8978
rect 4086 8956 4090 8960
rect 4229 8969 4233 8973
rect 4176 8956 4180 8960
rect 3488 8923 3492 8927
rect 3721 8933 3727 8937
rect 3801 8933 3805 8937
rect 3815 8933 3819 8937
rect 3833 8933 3837 8937
rect 3851 8933 3855 8937
rect 3874 8933 3878 8937
rect 3908 8933 3912 8937
rect 3923 8933 3927 8937
rect 3951 8933 3955 8937
rect 3733 8926 3739 8930
rect 3815 8926 3819 8930
rect 3874 8926 3878 8930
rect 3899 8926 3903 8930
rect 3930 8926 3934 8930
rect 3532 8915 3536 8919
rect 3815 8918 3819 8922
rect 3858 8919 3862 8923
rect 3880 8918 3887 8922
rect 3930 8919 3934 8923
rect 3769 8912 3775 8916
rect 3801 8914 3805 8918
rect 3833 8914 3837 8918
rect 3851 8914 3855 8918
rect 3908 8914 3912 8918
rect 3923 8914 3927 8918
rect 3951 8914 3955 8918
rect 3796 8902 3800 8906
rect 2856 8884 2860 8888
rect 2881 8881 2885 8885
rect 2888 8884 2892 8888
rect 2906 8884 2910 8888
rect 2928 8881 2932 8885
rect 2953 8881 2957 8885
rect 2963 8884 2967 8888
rect 2979 8884 2983 8888
rect 2999 8881 3003 8885
rect 3006 8884 3010 8888
rect 3660 8892 3665 8896
rect 2800 8874 2806 8878
rect 2882 8874 2886 8878
rect 2913 8874 2917 8878
rect 2935 8874 2939 8878
rect 3000 8874 3004 8878
rect 3060 8878 3064 8882
rect 3141 8878 3145 8882
rect 3406 8885 3410 8889
rect 3828 8900 3832 8904
rect 3848 8903 3852 8907
rect 3867 8899 3871 8903
rect 3886 8900 3890 8904
rect 3905 8900 3909 8904
rect 3918 8901 3922 8905
rect 4015 8914 4019 8918
rect 4096 8914 4100 8918
rect 4186 8914 4190 8918
rect 3940 8900 3944 8904
rect 3948 8901 3952 8905
rect 3960 8901 3964 8905
rect 3995 8899 3999 8903
rect 4023 8898 4027 8902
rect 4075 8899 4079 8903
rect 4104 8898 4108 8902
rect 4159 8899 4163 8903
rect 4194 8898 4198 8902
rect 3488 8882 3492 8886
rect 3757 8882 3763 8886
rect 3801 8884 3805 8888
rect 3231 8878 3235 8882
rect 3826 8881 3830 8885
rect 3833 8884 3837 8888
rect 3851 8884 3855 8888
rect 3873 8881 3877 8885
rect 3898 8881 3902 8885
rect 3908 8884 3912 8888
rect 3924 8884 3928 8888
rect 3944 8881 3948 8885
rect 3951 8884 3955 8888
rect 2764 8867 2770 8871
rect 2855 8867 2859 8871
rect 2889 8867 2893 8871
rect 2906 8867 2910 8871
rect 2962 8867 2966 8871
rect 2979 8867 2983 8871
rect 3007 8867 3011 8871
rect 3328 8870 3332 8874
rect 3745 8874 3751 8878
rect 3827 8874 3831 8878
rect 3858 8874 3862 8878
rect 3880 8874 3884 8878
rect 3945 8874 3949 8878
rect 3414 8869 3418 8873
rect 4005 8878 4009 8882
rect 4086 8878 4090 8882
rect 4176 8878 4180 8882
rect 2800 8860 2806 8864
rect 2882 8860 2886 8864
rect 2913 8860 2917 8864
rect 2935 8860 2939 8864
rect 3000 8860 3004 8864
rect 3070 8860 3074 8864
rect 3709 8867 3715 8871
rect 3800 8867 3804 8871
rect 3834 8867 3838 8871
rect 3851 8867 3855 8871
rect 3907 8867 3911 8871
rect 3924 8867 3928 8871
rect 3952 8867 3956 8871
rect 2856 8850 2860 8854
rect 2881 8853 2885 8857
rect 2888 8850 2892 8854
rect 2906 8850 2910 8854
rect 2928 8853 2932 8857
rect 2953 8853 2957 8857
rect 2963 8850 2967 8854
rect 2979 8850 2983 8854
rect 2999 8853 3003 8857
rect 3006 8850 3010 8854
rect 2850 8833 2854 8837
rect 2883 8834 2887 8838
rect 2903 8831 2907 8835
rect 2922 8835 2926 8839
rect 2941 8834 2945 8838
rect 2960 8834 2964 8838
rect 2973 8833 2977 8837
rect 2995 8834 2999 8838
rect 3003 8833 3007 8837
rect 3015 8833 3019 8837
rect 3078 8838 3082 8846
rect 3745 8860 3751 8864
rect 3827 8860 3831 8864
rect 3858 8860 3862 8864
rect 3880 8860 3884 8864
rect 3945 8860 3949 8864
rect 4015 8860 4019 8864
rect 3396 8849 3400 8853
rect 3801 8850 3805 8854
rect 3826 8853 3830 8857
rect 3833 8850 3837 8854
rect 3851 8850 3855 8854
rect 3873 8853 3877 8857
rect 3898 8853 3902 8857
rect 3908 8850 3912 8854
rect 3924 8850 3928 8854
rect 3944 8853 3948 8857
rect 3951 8850 3955 8854
rect 3668 8842 3672 8846
rect 3047 8832 3051 8836
rect 3101 8837 3105 8841
rect 3795 8833 3799 8837
rect 2351 8819 2355 8823
rect 2476 8819 2480 8823
rect 2856 8820 2860 8824
rect 2888 8820 2892 8824
rect 2906 8820 2910 8824
rect 2963 8820 2967 8824
rect 2978 8820 2982 8824
rect 3006 8820 3010 8824
rect 2870 8816 2874 8820
rect 2373 8812 2377 8816
rect 2409 8812 2413 8816
rect 2476 8812 2480 8816
rect 2505 8812 2509 8816
rect 2541 8812 2545 8816
rect 2608 8812 2612 8816
rect 2637 8812 2641 8816
rect 2673 8812 2677 8816
rect 2740 8812 2744 8816
rect 2824 8812 2830 8816
rect 2913 8815 2917 8819
rect 2935 8816 2942 8820
rect 2985 8815 2989 8819
rect 2764 8805 2770 8809
rect 2870 8808 2874 8812
rect 2879 8808 2883 8812
rect 2929 8808 2933 8812
rect 2954 8808 2958 8812
rect 2985 8808 2989 8812
rect 3060 8824 3064 8828
rect 3828 8834 3832 8838
rect 3848 8831 3852 8835
rect 3867 8835 3871 8839
rect 3886 8834 3890 8838
rect 3905 8834 3909 8838
rect 3918 8833 3922 8837
rect 3940 8834 3944 8838
rect 3948 8833 3952 8837
rect 3960 8833 3964 8837
rect 4023 8838 4027 8846
rect 3992 8832 3996 8836
rect 4046 8837 4050 8841
rect 3801 8820 3805 8824
rect 3833 8820 3837 8824
rect 3851 8820 3855 8824
rect 3908 8820 3912 8824
rect 3923 8820 3927 8824
rect 3951 8820 3955 8824
rect 3815 8816 3819 8820
rect 3318 8812 3322 8816
rect 3354 8812 3358 8816
rect 3421 8812 3425 8816
rect 3450 8812 3454 8816
rect 3486 8812 3490 8816
rect 3553 8812 3557 8816
rect 3582 8812 3586 8816
rect 3618 8812 3622 8816
rect 3685 8812 3689 8816
rect 3769 8812 3775 8816
rect 3858 8815 3862 8819
rect 3880 8816 3887 8820
rect 3930 8815 3934 8819
rect 3709 8805 3715 8809
rect 3815 8808 3819 8812
rect 3824 8808 3828 8812
rect 3874 8808 3878 8812
rect 3899 8808 3903 8812
rect 3930 8808 3934 8812
rect 4005 8824 4009 8828
rect 2373 8798 2377 8802
rect 2423 8798 2427 8802
rect 2476 8798 2480 8802
rect 2505 8798 2509 8802
rect 2555 8798 2559 8802
rect 2608 8798 2612 8802
rect 2637 8798 2641 8802
rect 2687 8798 2691 8802
rect 2740 8798 2744 8802
rect 2776 8801 2782 8805
rect 2856 8801 2860 8805
rect 2870 8801 2874 8805
rect 2888 8801 2892 8805
rect 2906 8801 2910 8805
rect 2929 8801 2933 8805
rect 2963 8801 2967 8805
rect 2978 8801 2982 8805
rect 3006 8801 3010 8805
rect 3131 8801 3135 8805
rect 3149 8801 3153 8805
rect 3167 8801 3171 8805
rect 3190 8801 3194 8805
rect 3224 8801 3228 8805
rect 3239 8801 3243 8805
rect 3267 8801 3271 8805
rect 2396 8787 2400 8791
rect 2367 8778 2371 8782
rect 2380 8781 2384 8787
rect 2417 8781 2421 8787
rect 2430 8783 2434 8787
rect 2454 8787 2458 8791
rect 2528 8787 2532 8791
rect 2438 8781 2442 8787
rect 2475 8781 2479 8787
rect 2491 8781 2495 8787
rect 2512 8781 2516 8787
rect 2549 8781 2553 8787
rect 2562 8783 2566 8787
rect 2586 8787 2590 8791
rect 2660 8787 2664 8791
rect 2570 8781 2574 8787
rect 2607 8781 2611 8787
rect 2623 8781 2627 8787
rect 2644 8781 2648 8787
rect 2681 8781 2685 8787
rect 2694 8783 2698 8787
rect 2718 8787 2722 8791
rect 2788 8794 2794 8798
rect 2870 8794 2874 8798
rect 2879 8794 2883 8798
rect 2929 8794 2933 8798
rect 2954 8794 2958 8798
rect 2985 8794 2989 8798
rect 2702 8781 2706 8787
rect 2739 8781 2743 8787
rect 2755 8783 2759 8787
rect 2870 8786 2874 8790
rect 2913 8787 2917 8791
rect 2935 8786 2942 8790
rect 2985 8787 2989 8791
rect 2856 8782 2860 8786
rect 2888 8782 2892 8786
rect 2906 8782 2910 8786
rect 2963 8782 2967 8786
rect 2978 8782 2982 8786
rect 3006 8782 3010 8786
rect 2380 8768 2384 8772
rect 2396 8768 2400 8774
rect 2430 8774 2434 8778
rect 2417 8768 2421 8772
rect 2438 8768 2442 8772
rect 2454 8768 2458 8774
rect 2475 8768 2479 8772
rect 2491 8768 2495 8772
rect 2512 8768 2516 8772
rect 2528 8768 2532 8774
rect 2562 8774 2566 8778
rect 2549 8768 2553 8772
rect 2570 8768 2574 8772
rect 2586 8768 2590 8774
rect 2607 8768 2611 8772
rect 2623 8768 2627 8772
rect 2644 8768 2648 8772
rect 2660 8768 2664 8774
rect 2694 8774 2698 8778
rect 2681 8768 2685 8772
rect 2702 8768 2706 8772
rect 2718 8768 2722 8774
rect 2739 8768 2743 8772
rect 2755 8768 2759 8772
rect 2851 8770 2855 8774
rect 2373 8757 2377 8761
rect 2410 8755 2414 8759
rect 2430 8755 2434 8759
rect 2474 8755 2478 8759
rect 2505 8757 2509 8761
rect 2542 8755 2546 8759
rect 2562 8755 2566 8759
rect 2606 8755 2610 8759
rect 2637 8757 2641 8761
rect 2674 8755 2678 8759
rect 2694 8755 2698 8759
rect 2738 8755 2742 8759
rect 2883 8768 2887 8772
rect 2903 8771 2907 8775
rect 2922 8767 2926 8771
rect 2941 8768 2945 8772
rect 2960 8768 2964 8772
rect 2973 8769 2977 8773
rect 3109 8794 3113 8798
rect 3131 8794 3135 8798
rect 3190 8794 3194 8798
rect 3215 8794 3219 8798
rect 3246 8794 3250 8798
rect 3318 8798 3322 8802
rect 3368 8798 3372 8802
rect 3421 8798 3425 8802
rect 3450 8798 3454 8802
rect 3500 8798 3504 8802
rect 3553 8798 3557 8802
rect 3582 8798 3586 8802
rect 3632 8798 3636 8802
rect 3685 8798 3689 8802
rect 3721 8801 3727 8805
rect 3801 8801 3805 8805
rect 3815 8801 3819 8805
rect 3833 8801 3837 8805
rect 3851 8801 3855 8805
rect 3874 8801 3878 8805
rect 3908 8801 3912 8805
rect 3923 8801 3927 8805
rect 3951 8801 3955 8805
rect 4076 8801 4080 8805
rect 4094 8801 4098 8805
rect 4112 8801 4116 8805
rect 4135 8801 4139 8805
rect 4169 8801 4173 8805
rect 4184 8801 4188 8805
rect 4212 8801 4216 8805
rect 3131 8786 3135 8790
rect 3174 8787 3178 8791
rect 3196 8786 3203 8790
rect 3246 8787 3250 8791
rect 3341 8787 3345 8791
rect 3149 8782 3153 8786
rect 3167 8782 3171 8786
rect 3224 8782 3228 8786
rect 3239 8782 3243 8786
rect 3267 8782 3271 8786
rect 3070 8778 3074 8782
rect 2995 8768 2999 8772
rect 3003 8769 3007 8773
rect 3015 8769 3019 8773
rect 3049 8763 3053 8767
rect 3089 8769 3093 8773
rect 3078 8762 3082 8766
rect 2856 8752 2860 8756
rect 2776 8748 2782 8752
rect 2881 8749 2885 8753
rect 2888 8752 2892 8756
rect 2906 8752 2910 8756
rect 2928 8749 2932 8753
rect 2953 8749 2957 8753
rect 2963 8752 2967 8756
rect 2979 8752 2983 8756
rect 2999 8749 3003 8753
rect 3006 8752 3010 8756
rect 3144 8768 3148 8772
rect 3164 8771 3168 8775
rect 3183 8767 3187 8771
rect 3312 8778 3316 8782
rect 3325 8781 3329 8787
rect 3362 8781 3366 8787
rect 3375 8783 3379 8787
rect 3399 8787 3403 8791
rect 3473 8787 3477 8791
rect 3383 8781 3387 8787
rect 3420 8781 3424 8787
rect 3436 8781 3440 8787
rect 3457 8781 3461 8787
rect 3494 8781 3498 8787
rect 3507 8783 3511 8787
rect 3531 8787 3535 8791
rect 3605 8787 3609 8791
rect 3515 8781 3519 8787
rect 3552 8781 3556 8787
rect 3568 8781 3572 8787
rect 3589 8781 3593 8787
rect 3626 8781 3630 8787
rect 3639 8783 3643 8787
rect 3663 8787 3667 8791
rect 3733 8794 3739 8798
rect 3815 8794 3819 8798
rect 3824 8794 3828 8798
rect 3874 8794 3878 8798
rect 3899 8794 3903 8798
rect 3930 8794 3934 8798
rect 3647 8781 3651 8787
rect 3684 8781 3688 8787
rect 3700 8783 3704 8787
rect 3815 8786 3819 8790
rect 3858 8787 3862 8791
rect 3880 8786 3887 8790
rect 3930 8787 3934 8791
rect 3801 8782 3805 8786
rect 3833 8782 3837 8786
rect 3851 8782 3855 8786
rect 3908 8782 3912 8786
rect 3923 8782 3927 8786
rect 3951 8782 3955 8786
rect 3202 8768 3206 8772
rect 3221 8768 3225 8772
rect 3234 8769 3238 8773
rect 3256 8768 3260 8772
rect 3264 8769 3268 8773
rect 3276 8769 3280 8773
rect 3325 8768 3329 8772
rect 3341 8768 3345 8774
rect 3375 8774 3379 8778
rect 3362 8768 3366 8772
rect 3383 8768 3387 8772
rect 3399 8768 3403 8774
rect 3420 8768 3424 8772
rect 3436 8768 3440 8772
rect 3457 8768 3461 8772
rect 3473 8768 3477 8774
rect 3507 8774 3511 8778
rect 3494 8768 3498 8772
rect 3515 8768 3519 8772
rect 3531 8768 3535 8774
rect 3552 8768 3556 8772
rect 3568 8768 3572 8772
rect 3589 8768 3593 8772
rect 3605 8768 3609 8774
rect 3639 8774 3643 8778
rect 3626 8768 3630 8772
rect 3647 8768 3651 8772
rect 3663 8768 3667 8774
rect 3684 8768 3688 8772
rect 3700 8768 3704 8772
rect 3796 8770 3800 8774
rect 3090 8752 3094 8756
rect 3116 8752 3120 8756
rect 2373 8741 2377 8745
rect 2424 8741 2428 8745
rect 2474 8741 2478 8745
rect 2505 8741 2509 8745
rect 2556 8741 2560 8745
rect 2606 8741 2610 8745
rect 2637 8741 2641 8745
rect 2688 8741 2692 8745
rect 2738 8741 2742 8745
rect 2812 8742 2818 8746
rect 2864 8742 2868 8746
rect 2882 8742 2886 8746
rect 2913 8742 2917 8746
rect 2935 8742 2939 8746
rect 3000 8742 3004 8746
rect 3142 8749 3146 8753
rect 3149 8752 3153 8756
rect 3167 8752 3171 8756
rect 3189 8749 3193 8753
rect 3214 8749 3218 8753
rect 3224 8752 3228 8756
rect 3240 8752 3244 8756
rect 3260 8749 3264 8753
rect 3267 8752 3271 8756
rect 3318 8757 3322 8761
rect 3355 8755 3359 8759
rect 3375 8755 3379 8759
rect 3419 8755 3423 8759
rect 3450 8757 3454 8761
rect 3487 8755 3491 8759
rect 3507 8755 3511 8759
rect 3551 8755 3555 8759
rect 3582 8757 3586 8761
rect 3619 8755 3623 8759
rect 3639 8755 3643 8759
rect 3683 8755 3687 8759
rect 3828 8768 3832 8772
rect 3848 8771 3852 8775
rect 3867 8767 3871 8771
rect 3886 8768 3890 8772
rect 3905 8768 3909 8772
rect 3918 8769 3922 8773
rect 4054 8794 4058 8798
rect 4076 8794 4080 8798
rect 4135 8794 4139 8798
rect 4160 8794 4164 8798
rect 4191 8794 4195 8798
rect 4076 8786 4080 8790
rect 4119 8787 4123 8791
rect 4141 8786 4148 8790
rect 4191 8787 4195 8791
rect 4094 8782 4098 8786
rect 4112 8782 4116 8786
rect 4169 8782 4173 8786
rect 4184 8782 4188 8786
rect 4212 8782 4216 8786
rect 4015 8778 4019 8782
rect 3940 8768 3944 8772
rect 3948 8769 3952 8773
rect 3960 8769 3964 8773
rect 3994 8763 3998 8767
rect 4034 8769 4038 8773
rect 4023 8762 4027 8766
rect 3801 8752 3805 8756
rect 3721 8748 3727 8752
rect 3826 8749 3830 8753
rect 3833 8752 3837 8756
rect 3851 8752 3855 8756
rect 3873 8749 3877 8753
rect 3898 8749 3902 8753
rect 3908 8752 3912 8756
rect 3924 8752 3928 8756
rect 3944 8749 3948 8753
rect 3951 8752 3955 8756
rect 4089 8768 4093 8772
rect 4109 8771 4113 8775
rect 4128 8767 4132 8771
rect 4147 8768 4151 8772
rect 4166 8768 4170 8772
rect 4179 8769 4183 8773
rect 4201 8768 4205 8772
rect 4209 8769 4213 8773
rect 4221 8769 4225 8773
rect 4035 8752 4039 8756
rect 4061 8752 4065 8756
rect 3060 8742 3064 8746
rect 3099 8742 3103 8746
rect 3143 8742 3147 8746
rect 3174 8742 3178 8746
rect 3196 8742 3200 8746
rect 3261 8742 3265 8746
rect 3318 8741 3322 8745
rect 3369 8741 3373 8745
rect 3419 8741 3423 8745
rect 3450 8741 3454 8745
rect 3501 8741 3505 8745
rect 3551 8741 3555 8745
rect 3582 8741 3586 8745
rect 3633 8741 3637 8745
rect 3683 8741 3687 8745
rect 3757 8742 3763 8746
rect 3809 8742 3813 8746
rect 3827 8742 3831 8746
rect 3858 8742 3862 8746
rect 3880 8742 3884 8746
rect 3945 8742 3949 8746
rect 4087 8749 4091 8753
rect 4094 8752 4098 8756
rect 4112 8752 4116 8756
rect 4134 8749 4138 8753
rect 4159 8749 4163 8753
rect 4169 8752 4173 8756
rect 4185 8752 4189 8756
rect 4205 8749 4209 8753
rect 4212 8752 4216 8756
rect 4484 8747 4488 8751
rect 4494 8747 4498 8751
rect 4504 8747 4508 8751
rect 4005 8742 4009 8746
rect 4044 8742 4048 8746
rect 4088 8742 4092 8746
rect 4119 8742 4123 8746
rect 4141 8742 4145 8746
rect 4206 8742 4210 8746
rect 4484 8742 4488 8746
rect 4494 8742 4498 8746
rect 4504 8742 4508 8746
rect 2367 8734 2371 8738
rect 2755 8734 2759 8738
rect 2764 8735 2770 8739
rect 2855 8735 2859 8739
rect 2889 8735 2893 8739
rect 2906 8735 2910 8739
rect 2962 8735 2966 8739
rect 2979 8735 2983 8739
rect 3007 8735 3011 8739
rect 3090 8735 3094 8739
rect 3116 8735 3120 8739
rect 3150 8735 3154 8739
rect 3167 8735 3171 8739
rect 3223 8735 3227 8739
rect 3240 8735 3244 8739
rect 3268 8735 3272 8739
rect 3312 8734 3316 8738
rect 3700 8734 3704 8738
rect 3709 8735 3715 8739
rect 3800 8735 3804 8739
rect 3834 8735 3838 8739
rect 3851 8735 3855 8739
rect 3907 8735 3911 8739
rect 3924 8735 3928 8739
rect 3952 8735 3956 8739
rect 4035 8735 4039 8739
rect 4061 8735 4065 8739
rect 4095 8735 4099 8739
rect 4112 8735 4116 8739
rect 4168 8735 4172 8739
rect 4185 8735 4189 8739
rect 4213 8735 4217 8739
rect 4484 8737 4488 8741
rect 4494 8737 4498 8741
rect 4504 8737 4508 8741
rect 2490 8727 2495 8731
rect 2623 8727 2627 8731
rect 2800 8728 2806 8732
rect 2864 8728 2868 8732
rect 3098 8728 3102 8732
rect 3284 8729 3288 8733
rect 3296 8729 3300 8733
rect 3435 8727 3440 8731
rect 3568 8727 3572 8731
rect 3745 8728 3751 8732
rect 3809 8728 3813 8732
rect 4043 8728 4047 8732
rect 4229 8729 4233 8733
rect 4241 8729 4245 8733
rect 4484 8732 4488 8736
rect 4494 8732 4498 8736
rect 4504 8732 4508 8736
rect 4530 8747 4534 8751
rect 4540 8747 4544 8751
rect 4550 8747 4554 8751
rect 4530 8742 4534 8746
rect 4540 8742 4544 8746
rect 4550 8742 4554 8746
rect 4530 8737 4534 8741
rect 4540 8737 4544 8741
rect 4550 8737 4554 8741
rect 4530 8732 4534 8736
rect 4540 8732 4544 8736
rect 4550 8732 4554 8736
rect 2498 8720 2502 8724
rect 2788 8720 2794 8724
rect 3108 8721 3112 8725
rect 3273 8721 3277 8725
rect 2482 8715 2486 8719
rect 2514 8715 2518 8719
rect 2836 8714 2842 8718
rect 3443 8720 3447 8724
rect 3733 8720 3739 8724
rect 4053 8721 4057 8725
rect 4218 8721 4222 8725
rect 3427 8715 3431 8719
rect 3459 8715 3463 8719
rect 3781 8714 3787 8718
rect 2351 8707 2355 8711
rect 2482 8707 2486 8711
rect 2514 8707 2518 8711
rect 3427 8707 3431 8711
rect 3459 8707 3463 8711
rect 618 8703 622 8707
rect 628 8703 632 8707
rect 638 8703 642 8707
rect 618 8698 622 8702
rect 628 8698 632 8702
rect 638 8698 642 8702
rect 618 8693 622 8697
rect 628 8693 632 8697
rect 638 8693 642 8697
rect 618 8688 622 8692
rect 628 8688 632 8692
rect 638 8688 642 8692
rect 664 8703 668 8707
rect 674 8703 678 8707
rect 684 8703 688 8707
rect 664 8698 668 8702
rect 674 8698 678 8702
rect 684 8698 688 8702
rect 664 8693 668 8697
rect 674 8693 678 8697
rect 684 8693 688 8697
rect 2498 8700 2502 8704
rect 2755 8700 2759 8704
rect 2824 8700 2830 8704
rect 3156 8700 3160 8704
rect 3192 8700 3196 8704
rect 3259 8700 3263 8704
rect 3443 8700 3447 8704
rect 3700 8700 3704 8704
rect 3769 8700 3775 8704
rect 4101 8700 4105 8704
rect 4137 8700 4141 8704
rect 4204 8700 4208 8704
rect 2755 8692 2759 8696
rect 2764 8693 2770 8697
rect 3142 8693 3146 8697
rect 664 8688 668 8692
rect 674 8688 678 8692
rect 684 8688 688 8692
rect 2482 8688 2486 8692
rect 2514 8688 2518 8692
rect 2498 8684 2502 8688
rect 3156 8686 3160 8690
rect 3206 8686 3210 8690
rect 3259 8686 3263 8690
rect 3700 8692 3704 8696
rect 3709 8693 3715 8697
rect 4087 8693 4091 8697
rect 3427 8688 3431 8692
rect 3459 8688 3463 8692
rect 3443 8684 3447 8688
rect 4101 8686 4105 8690
rect 4151 8686 4155 8690
rect 4204 8686 4208 8690
rect 2490 8677 2495 8681
rect 2624 8677 2628 8681
rect 3179 8675 3183 8679
rect 2373 8670 2377 8674
rect 2409 8670 2413 8674
rect 2476 8670 2480 8674
rect 2505 8670 2509 8674
rect 2541 8670 2545 8674
rect 2608 8670 2612 8674
rect 2637 8670 2641 8674
rect 2673 8670 2677 8674
rect 2740 8670 2744 8674
rect 2824 8670 2830 8674
rect 2764 8663 2770 8667
rect 3150 8666 3154 8670
rect 3163 8669 3167 8675
rect 3200 8669 3204 8675
rect 3213 8671 3217 8675
rect 3237 8675 3241 8679
rect 3435 8677 3440 8681
rect 3569 8677 3573 8681
rect 4124 8675 4128 8679
rect 3221 8669 3225 8675
rect 3258 8669 3262 8675
rect 3274 8669 3278 8675
rect 3318 8670 3322 8674
rect 3354 8670 3358 8674
rect 3421 8670 3425 8674
rect 3450 8670 3454 8674
rect 3486 8670 3490 8674
rect 3553 8670 3557 8674
rect 3582 8670 3586 8674
rect 3618 8670 3622 8674
rect 3685 8670 3689 8674
rect 3769 8670 3775 8674
rect 2373 8656 2377 8660
rect 2423 8656 2427 8660
rect 2476 8656 2480 8660
rect 2505 8656 2509 8660
rect 2555 8656 2559 8660
rect 2608 8656 2612 8660
rect 2637 8656 2641 8660
rect 2687 8656 2691 8660
rect 2740 8656 2744 8660
rect 3163 8656 3167 8660
rect 3179 8656 3183 8662
rect 3213 8662 3217 8666
rect 3200 8656 3204 8660
rect 2396 8645 2400 8649
rect 2367 8636 2371 8640
rect 2380 8639 2384 8645
rect 2417 8639 2421 8645
rect 2430 8641 2434 8645
rect 2454 8645 2458 8649
rect 2528 8645 2532 8649
rect 2438 8639 2442 8645
rect 2475 8639 2479 8645
rect 2491 8639 2495 8645
rect 2512 8639 2516 8645
rect 2549 8639 2553 8645
rect 2562 8641 2566 8645
rect 2586 8645 2590 8649
rect 2660 8645 2664 8649
rect 2570 8639 2574 8645
rect 2607 8639 2611 8645
rect 2623 8639 2627 8645
rect 2644 8639 2648 8645
rect 2681 8639 2685 8645
rect 2694 8641 2698 8645
rect 2718 8645 2722 8649
rect 2702 8639 2706 8645
rect 2739 8639 2743 8645
rect 2755 8641 2759 8645
rect 3221 8656 3225 8660
rect 3237 8656 3241 8662
rect 3709 8663 3715 8667
rect 4095 8666 4099 8670
rect 4108 8669 4112 8675
rect 4145 8669 4149 8675
rect 4158 8671 4162 8675
rect 4182 8675 4186 8679
rect 4166 8669 4170 8675
rect 4203 8669 4207 8675
rect 4219 8669 4223 8675
rect 3258 8656 3262 8660
rect 3274 8656 3278 8660
rect 3318 8656 3322 8660
rect 3368 8656 3372 8660
rect 3421 8656 3425 8660
rect 3450 8656 3454 8660
rect 3500 8656 3504 8660
rect 3553 8656 3557 8660
rect 3582 8656 3586 8660
rect 3632 8656 3636 8660
rect 3685 8656 3689 8660
rect 4108 8656 4112 8660
rect 4124 8656 4128 8662
rect 4158 8662 4162 8666
rect 4145 8656 4149 8660
rect 3156 8645 3160 8649
rect 3193 8643 3197 8647
rect 3213 8643 3217 8647
rect 3257 8643 3261 8647
rect 3341 8645 3345 8649
rect 2380 8626 2384 8630
rect 2396 8626 2400 8632
rect 2430 8632 2434 8636
rect 2417 8626 2421 8630
rect 2438 8626 2442 8630
rect 2454 8626 2458 8632
rect 2475 8626 2479 8630
rect 2491 8626 2495 8630
rect 2512 8626 2516 8630
rect 2528 8626 2532 8632
rect 2562 8632 2566 8636
rect 2549 8626 2553 8630
rect 2570 8626 2574 8630
rect 2586 8626 2590 8632
rect 2607 8626 2611 8630
rect 2623 8626 2627 8630
rect 2644 8626 2648 8630
rect 2660 8626 2664 8632
rect 2694 8632 2698 8636
rect 2681 8626 2685 8630
rect 2702 8626 2706 8630
rect 2718 8626 2722 8632
rect 2776 8636 2782 8640
rect 3312 8636 3316 8640
rect 3325 8639 3329 8645
rect 3362 8639 3366 8645
rect 3375 8641 3379 8645
rect 3399 8645 3403 8649
rect 3473 8645 3477 8649
rect 3383 8639 3387 8645
rect 3420 8639 3424 8645
rect 3436 8639 3440 8645
rect 3457 8639 3461 8645
rect 3494 8639 3498 8645
rect 3507 8641 3511 8645
rect 3531 8645 3535 8649
rect 3605 8645 3609 8649
rect 3515 8639 3519 8645
rect 3552 8639 3556 8645
rect 3568 8639 3572 8645
rect 3589 8639 3593 8645
rect 3626 8639 3630 8645
rect 3639 8641 3643 8645
rect 3663 8645 3667 8649
rect 3647 8639 3651 8645
rect 3684 8639 3688 8645
rect 3700 8641 3704 8645
rect 4166 8656 4170 8660
rect 4182 8656 4186 8662
rect 4203 8656 4207 8660
rect 4219 8656 4223 8660
rect 4101 8645 4105 8649
rect 4138 8643 4142 8647
rect 4158 8643 4162 8647
rect 4202 8643 4206 8647
rect 2739 8626 2743 8630
rect 2755 8626 2759 8630
rect 2812 8629 2818 8633
rect 3156 8629 3160 8633
rect 3207 8629 3211 8633
rect 3257 8629 3261 8633
rect 3325 8626 3329 8630
rect 3341 8626 3345 8632
rect 3375 8632 3379 8636
rect 3362 8626 3366 8630
rect 2373 8615 2377 8619
rect 2410 8613 2414 8617
rect 2430 8613 2434 8617
rect 2474 8613 2478 8617
rect 2505 8615 2509 8619
rect 2542 8613 2546 8617
rect 2562 8613 2566 8617
rect 2606 8613 2610 8617
rect 2637 8615 2641 8619
rect 2674 8613 2678 8617
rect 2694 8613 2698 8617
rect 2738 8613 2742 8617
rect 3149 8621 3153 8625
rect 3274 8622 3278 8626
rect 3383 8626 3387 8630
rect 3399 8626 3403 8632
rect 3420 8626 3424 8630
rect 3436 8626 3440 8630
rect 3457 8626 3461 8630
rect 3473 8626 3477 8632
rect 3507 8632 3511 8636
rect 3494 8626 3498 8630
rect 3515 8626 3519 8630
rect 3531 8626 3535 8632
rect 3552 8626 3556 8630
rect 3568 8626 3572 8630
rect 3589 8626 3593 8630
rect 3605 8626 3609 8632
rect 3639 8632 3643 8636
rect 3626 8626 3630 8630
rect 3647 8626 3651 8630
rect 3663 8626 3667 8632
rect 3721 8636 3727 8640
rect 3684 8626 3688 8630
rect 3700 8626 3704 8630
rect 3757 8629 3763 8633
rect 4101 8629 4105 8633
rect 4152 8629 4156 8633
rect 4202 8629 4206 8633
rect 2824 8614 2830 8618
rect 3156 8614 3160 8618
rect 3192 8614 3196 8618
rect 3259 8614 3263 8618
rect 2776 8606 2782 8610
rect 3142 8607 3146 8611
rect 3318 8615 3322 8619
rect 3355 8613 3359 8617
rect 3375 8613 3379 8617
rect 3419 8613 3423 8617
rect 3450 8615 3454 8619
rect 3487 8613 3491 8617
rect 3507 8613 3511 8617
rect 3551 8613 3555 8617
rect 3582 8615 3586 8619
rect 3619 8613 3623 8617
rect 3639 8613 3643 8617
rect 3683 8613 3687 8617
rect 4094 8621 4098 8625
rect 4219 8622 4223 8626
rect 3769 8614 3775 8618
rect 4101 8614 4105 8618
rect 4137 8614 4141 8618
rect 4204 8614 4208 8618
rect 2373 8599 2377 8603
rect 2424 8599 2428 8603
rect 2474 8599 2478 8603
rect 2505 8599 2509 8603
rect 2556 8599 2560 8603
rect 2606 8599 2610 8603
rect 2637 8599 2641 8603
rect 2688 8599 2692 8603
rect 2738 8599 2742 8603
rect 2812 8599 2818 8603
rect 3156 8600 3160 8604
rect 3206 8600 3210 8604
rect 3259 8600 3263 8604
rect 3721 8606 3727 8610
rect 4087 8607 4091 8611
rect 3318 8599 3322 8603
rect 3369 8599 3373 8603
rect 3419 8599 3423 8603
rect 3450 8599 3454 8603
rect 3501 8599 3505 8603
rect 3551 8599 3555 8603
rect 3582 8599 3586 8603
rect 3633 8599 3637 8603
rect 3683 8599 3687 8603
rect 3757 8599 3763 8603
rect 4101 8600 4105 8604
rect 4151 8600 4155 8604
rect 4204 8600 4208 8604
rect 2366 8592 2370 8596
rect 2755 8592 2759 8596
rect 3179 8589 3183 8593
rect 2373 8584 2377 8588
rect 2409 8584 2413 8588
rect 2476 8584 2480 8588
rect 2505 8584 2509 8588
rect 2541 8584 2545 8588
rect 2608 8584 2612 8588
rect 2637 8584 2641 8588
rect 2673 8584 2677 8588
rect 2740 8584 2744 8588
rect 2824 8584 2830 8588
rect 2764 8577 2770 8581
rect 3150 8580 3154 8584
rect 3163 8583 3167 8589
rect 3200 8583 3204 8589
rect 3213 8585 3217 8589
rect 3237 8589 3241 8593
rect 3311 8592 3315 8596
rect 3700 8592 3704 8596
rect 4124 8589 4128 8593
rect 3221 8583 3225 8589
rect 3258 8583 3262 8589
rect 3274 8585 3278 8589
rect 3296 8583 3300 8587
rect 3318 8584 3322 8588
rect 3354 8584 3358 8588
rect 3421 8584 3425 8588
rect 3450 8584 3454 8588
rect 3486 8584 3490 8588
rect 3553 8584 3557 8588
rect 3582 8584 3586 8588
rect 3618 8584 3622 8588
rect 3685 8584 3689 8588
rect 3769 8584 3775 8588
rect 2373 8570 2377 8574
rect 2423 8570 2427 8574
rect 2476 8570 2480 8574
rect 2505 8570 2509 8574
rect 2555 8570 2559 8574
rect 2608 8570 2612 8574
rect 2637 8570 2641 8574
rect 2687 8570 2691 8574
rect 2740 8570 2744 8574
rect 3163 8570 3167 8574
rect 3179 8570 3183 8576
rect 3213 8576 3217 8580
rect 3200 8570 3204 8574
rect 2396 8559 2400 8563
rect 2367 8550 2371 8554
rect 2380 8553 2384 8559
rect 2417 8553 2421 8559
rect 2430 8555 2434 8559
rect 2454 8559 2458 8563
rect 2528 8559 2532 8563
rect 2438 8553 2442 8559
rect 2475 8553 2479 8559
rect 2491 8553 2495 8559
rect 2512 8553 2516 8559
rect 2549 8553 2553 8559
rect 2562 8555 2566 8559
rect 2586 8559 2590 8563
rect 2660 8559 2664 8563
rect 2570 8553 2574 8559
rect 2607 8553 2611 8559
rect 2623 8553 2627 8559
rect 2644 8553 2648 8559
rect 2681 8553 2685 8559
rect 2694 8555 2698 8559
rect 2718 8559 2722 8563
rect 2702 8553 2706 8559
rect 2739 8553 2743 8559
rect 2755 8555 2759 8559
rect 3221 8570 3225 8574
rect 3237 8570 3241 8576
rect 3258 8570 3262 8574
rect 3274 8570 3278 8579
rect 3709 8577 3715 8581
rect 4095 8580 4099 8584
rect 4108 8583 4112 8589
rect 4145 8583 4149 8589
rect 4158 8585 4162 8589
rect 4182 8589 4186 8593
rect 4166 8583 4170 8589
rect 4203 8583 4207 8589
rect 4219 8585 4223 8589
rect 4241 8583 4245 8587
rect 3296 8567 3300 8571
rect 3318 8570 3322 8574
rect 3368 8570 3372 8574
rect 3421 8570 3425 8574
rect 3450 8570 3454 8574
rect 3500 8570 3504 8574
rect 3553 8570 3557 8574
rect 3582 8570 3586 8574
rect 3632 8570 3636 8574
rect 3685 8570 3689 8574
rect 4108 8570 4112 8574
rect 4124 8570 4128 8576
rect 4158 8576 4162 8580
rect 4145 8570 4149 8574
rect 3156 8559 3160 8563
rect 3193 8557 3197 8561
rect 3213 8557 3217 8561
rect 3257 8557 3261 8561
rect 3341 8559 3345 8563
rect 2380 8540 2384 8544
rect 2396 8540 2400 8546
rect 2430 8546 2434 8550
rect 2417 8540 2421 8544
rect 2438 8540 2442 8544
rect 2454 8540 2458 8546
rect 2475 8540 2479 8544
rect 2491 8540 2495 8544
rect 2512 8540 2516 8544
rect 2528 8540 2532 8546
rect 2562 8546 2566 8550
rect 2549 8540 2553 8544
rect 2570 8540 2574 8544
rect 2586 8540 2590 8546
rect 2607 8540 2611 8544
rect 2623 8540 2627 8544
rect 2644 8540 2648 8544
rect 2660 8540 2664 8546
rect 2694 8546 2698 8550
rect 2681 8540 2685 8544
rect 2702 8540 2706 8544
rect 2718 8540 2722 8546
rect 2776 8550 2782 8554
rect 3312 8550 3316 8554
rect 3325 8553 3329 8559
rect 3362 8553 3366 8559
rect 3375 8555 3379 8559
rect 3399 8559 3403 8563
rect 3473 8559 3477 8563
rect 3383 8553 3387 8559
rect 3420 8553 3424 8559
rect 3436 8553 3440 8559
rect 3457 8553 3461 8559
rect 3494 8553 3498 8559
rect 3507 8555 3511 8559
rect 3531 8559 3535 8563
rect 3605 8559 3609 8563
rect 3515 8553 3519 8559
rect 3552 8553 3556 8559
rect 3568 8553 3572 8559
rect 3589 8553 3593 8559
rect 3626 8553 3630 8559
rect 3639 8555 3643 8559
rect 3663 8559 3667 8563
rect 3647 8553 3651 8559
rect 3684 8553 3688 8559
rect 3700 8555 3704 8559
rect 4166 8570 4170 8574
rect 4182 8570 4186 8576
rect 4203 8570 4207 8574
rect 4219 8570 4223 8579
rect 4241 8567 4245 8571
rect 4101 8559 4105 8563
rect 4138 8557 4142 8561
rect 4158 8557 4162 8561
rect 4202 8557 4206 8561
rect 2739 8540 2743 8544
rect 2755 8540 2759 8544
rect 2812 8543 2818 8547
rect 3156 8543 3160 8547
rect 3207 8543 3211 8547
rect 3257 8543 3261 8547
rect 3325 8540 3329 8544
rect 3341 8540 3345 8546
rect 3375 8546 3379 8550
rect 3362 8540 3366 8544
rect 3383 8540 3387 8544
rect 3399 8540 3403 8546
rect 3420 8540 3424 8544
rect 3436 8540 3440 8544
rect 3457 8540 3461 8544
rect 3473 8540 3477 8546
rect 3507 8546 3511 8550
rect 3494 8540 3498 8544
rect 3515 8540 3519 8544
rect 3531 8540 3535 8546
rect 3552 8540 3556 8544
rect 3568 8540 3572 8544
rect 3589 8540 3593 8544
rect 3605 8540 3609 8546
rect 3639 8546 3643 8550
rect 3626 8540 3630 8544
rect 3647 8540 3651 8544
rect 3663 8540 3667 8546
rect 3721 8550 3727 8554
rect 3684 8540 3688 8544
rect 3700 8540 3704 8544
rect 3757 8543 3763 8547
rect 4101 8543 4105 8547
rect 4152 8543 4156 8547
rect 4202 8543 4206 8547
rect 2373 8529 2377 8533
rect 2410 8527 2414 8531
rect 2430 8527 2434 8531
rect 2474 8527 2478 8531
rect 2505 8529 2509 8533
rect 2542 8527 2546 8531
rect 2562 8527 2566 8531
rect 2606 8527 2610 8531
rect 2637 8529 2641 8533
rect 2674 8527 2678 8531
rect 2694 8527 2698 8531
rect 2738 8527 2742 8531
rect 3318 8529 3322 8533
rect 3355 8527 3359 8531
rect 3375 8527 3379 8531
rect 3419 8527 3423 8531
rect 3450 8529 3454 8533
rect 3487 8527 3491 8531
rect 3507 8527 3511 8531
rect 3551 8527 3555 8531
rect 3582 8529 3586 8533
rect 3619 8527 3623 8531
rect 3639 8527 3643 8531
rect 3683 8527 3687 8531
rect 2776 8520 2782 8524
rect 3721 8520 3727 8524
rect 2373 8513 2377 8517
rect 2424 8513 2428 8517
rect 2474 8513 2478 8517
rect 2505 8513 2509 8517
rect 2556 8513 2560 8517
rect 2606 8513 2610 8517
rect 2637 8513 2641 8517
rect 2688 8513 2692 8517
rect 2738 8513 2742 8517
rect 2812 8513 2818 8517
rect 3318 8513 3322 8517
rect 3369 8513 3373 8517
rect 3419 8513 3423 8517
rect 3450 8513 3454 8517
rect 3501 8513 3505 8517
rect 3551 8513 3555 8517
rect 3582 8513 3586 8517
rect 3633 8513 3637 8517
rect 3683 8513 3687 8517
rect 3757 8513 3763 8517
rect 2366 8506 2370 8510
rect 2755 8506 2759 8510
rect 3311 8506 3315 8510
rect 3700 8506 3704 8510
rect 2491 8499 2495 8503
rect 2599 8499 2603 8503
rect 2623 8499 2627 8503
rect 3436 8499 3440 8503
rect 3544 8499 3548 8503
rect 3568 8499 3572 8503
rect 2615 8492 2619 8496
rect 2599 8488 2603 8492
rect 2631 8488 2635 8492
rect 3560 8492 3564 8496
rect 3544 8488 3548 8492
rect 3576 8488 3580 8492
rect 2599 8481 2603 8485
rect 2631 8481 2635 8485
rect 3296 8481 3300 8485
rect 3544 8481 3548 8485
rect 3576 8481 3580 8485
rect 4241 8481 4245 8485
rect 2615 8474 2619 8478
rect 2755 8474 2759 8478
rect 3560 8474 3564 8478
rect 3700 8474 3704 8478
rect 2755 8466 2759 8470
rect 3700 8466 3704 8470
rect 2599 8462 2603 8466
rect 2631 8462 2635 8466
rect 2615 8458 2619 8462
rect 3544 8462 3548 8466
rect 3576 8462 3580 8466
rect 3560 8458 3564 8462
rect 2491 8451 2495 8455
rect 2599 8451 2603 8455
rect 2623 8451 2627 8455
rect 3436 8451 3440 8455
rect 3544 8451 3548 8455
rect 3568 8451 3572 8455
rect 2373 8444 2377 8448
rect 2409 8444 2413 8448
rect 2476 8444 2480 8448
rect 2505 8444 2509 8448
rect 2541 8444 2545 8448
rect 2608 8444 2612 8448
rect 2637 8444 2641 8448
rect 2673 8444 2677 8448
rect 2740 8444 2744 8448
rect 2824 8444 2830 8448
rect 3318 8444 3322 8448
rect 3354 8444 3358 8448
rect 3421 8444 3425 8448
rect 3450 8444 3454 8448
rect 3486 8444 3490 8448
rect 3553 8444 3557 8448
rect 3582 8444 3586 8448
rect 3618 8444 3622 8448
rect 3685 8444 3689 8448
rect 3769 8444 3775 8448
rect 2764 8437 2770 8441
rect 3709 8437 3715 8441
rect 4484 8438 4488 8442
rect 4494 8438 4498 8442
rect 4504 8438 4508 8442
rect 2373 8430 2377 8434
rect 2423 8430 2427 8434
rect 2476 8430 2480 8434
rect 2505 8430 2509 8434
rect 2555 8430 2559 8434
rect 2608 8430 2612 8434
rect 2637 8430 2641 8434
rect 2687 8430 2691 8434
rect 2740 8430 2744 8434
rect 3318 8430 3322 8434
rect 3368 8430 3372 8434
rect 3421 8430 3425 8434
rect 3450 8430 3454 8434
rect 3500 8430 3504 8434
rect 3553 8430 3557 8434
rect 3582 8430 3586 8434
rect 3632 8430 3636 8434
rect 3685 8430 3689 8434
rect 4484 8433 4488 8437
rect 4494 8433 4498 8437
rect 4504 8433 4508 8437
rect 4484 8428 4488 8432
rect 4494 8428 4498 8432
rect 4504 8428 4508 8432
rect 2396 8419 2400 8423
rect 2367 8410 2371 8414
rect 2380 8413 2384 8419
rect 2417 8413 2421 8419
rect 2430 8415 2434 8419
rect 2454 8419 2458 8423
rect 2528 8419 2532 8423
rect 2438 8413 2442 8419
rect 2475 8413 2479 8419
rect 2491 8413 2495 8419
rect 2512 8413 2516 8419
rect 2549 8413 2553 8419
rect 2562 8415 2566 8419
rect 2586 8419 2590 8423
rect 2660 8419 2664 8423
rect 2570 8413 2574 8419
rect 2607 8413 2611 8419
rect 2623 8413 2627 8419
rect 2644 8413 2648 8419
rect 2681 8413 2685 8419
rect 2694 8415 2698 8419
rect 2718 8419 2722 8423
rect 3341 8419 3345 8423
rect 2702 8413 2706 8419
rect 2739 8413 2743 8419
rect 2755 8415 2759 8419
rect 2380 8400 2384 8404
rect 2396 8400 2400 8406
rect 2430 8406 2434 8410
rect 2417 8400 2421 8404
rect 618 8394 622 8398
rect 628 8394 632 8398
rect 638 8394 642 8398
rect 618 8389 622 8393
rect 628 8389 632 8393
rect 638 8389 642 8393
rect 618 8384 622 8388
rect 628 8384 632 8388
rect 638 8384 642 8388
rect 618 8379 622 8383
rect 628 8379 632 8383
rect 638 8379 642 8383
rect 664 8394 668 8398
rect 674 8394 678 8398
rect 684 8394 688 8398
rect 664 8389 668 8393
rect 674 8389 678 8393
rect 684 8389 688 8393
rect 664 8384 668 8388
rect 674 8384 678 8388
rect 684 8384 688 8388
rect 2438 8400 2442 8404
rect 2454 8400 2458 8406
rect 2475 8400 2479 8404
rect 2491 8400 2495 8404
rect 2512 8400 2516 8404
rect 2528 8400 2532 8406
rect 2562 8406 2566 8410
rect 2549 8400 2553 8404
rect 2570 8400 2574 8404
rect 2586 8400 2590 8406
rect 2607 8400 2611 8404
rect 2623 8400 2627 8404
rect 2644 8400 2648 8404
rect 2660 8400 2664 8406
rect 2694 8406 2698 8410
rect 2681 8400 2685 8404
rect 2702 8400 2706 8404
rect 2718 8400 2722 8406
rect 3312 8410 3316 8414
rect 3325 8413 3329 8419
rect 3362 8413 3366 8419
rect 3375 8415 3379 8419
rect 3399 8419 3403 8423
rect 3473 8419 3477 8423
rect 3383 8413 3387 8419
rect 3420 8413 3424 8419
rect 3436 8413 3440 8419
rect 3457 8413 3461 8419
rect 3494 8413 3498 8419
rect 3507 8415 3511 8419
rect 3531 8419 3535 8423
rect 3605 8419 3609 8423
rect 3515 8413 3519 8419
rect 3552 8413 3556 8419
rect 3568 8413 3572 8419
rect 3589 8413 3593 8419
rect 3626 8413 3630 8419
rect 3639 8415 3643 8419
rect 3663 8419 3667 8423
rect 4484 8423 4488 8427
rect 4494 8423 4498 8427
rect 4504 8423 4508 8427
rect 4530 8438 4534 8442
rect 4540 8438 4544 8442
rect 4550 8438 4554 8442
rect 4530 8433 4534 8437
rect 4540 8433 4544 8437
rect 4550 8433 4554 8437
rect 4530 8428 4534 8432
rect 4540 8428 4544 8432
rect 4550 8428 4554 8432
rect 4530 8423 4534 8427
rect 4540 8423 4544 8427
rect 4550 8423 4554 8427
rect 3647 8413 3651 8419
rect 3684 8413 3688 8419
rect 3700 8415 3704 8419
rect 2739 8400 2743 8404
rect 2755 8400 2759 8404
rect 3325 8400 3329 8404
rect 3341 8400 3345 8406
rect 3375 8406 3379 8410
rect 3362 8400 3366 8404
rect 3383 8400 3387 8404
rect 3399 8400 3403 8406
rect 3420 8400 3424 8404
rect 3436 8400 3440 8404
rect 3457 8400 3461 8404
rect 3473 8400 3477 8406
rect 3507 8406 3511 8410
rect 3494 8400 3498 8404
rect 3515 8400 3519 8404
rect 3531 8400 3535 8406
rect 3552 8400 3556 8404
rect 3568 8400 3572 8404
rect 3589 8400 3593 8404
rect 3605 8400 3609 8406
rect 3639 8406 3643 8410
rect 3626 8400 3630 8404
rect 3647 8400 3651 8404
rect 3663 8400 3667 8406
rect 3684 8400 3688 8404
rect 3700 8400 3704 8404
rect 2373 8389 2377 8393
rect 2410 8387 2414 8391
rect 2430 8387 2434 8391
rect 2474 8387 2478 8391
rect 2505 8389 2509 8393
rect 2542 8387 2546 8391
rect 2562 8387 2566 8391
rect 2606 8387 2610 8391
rect 2637 8389 2641 8393
rect 2674 8387 2678 8391
rect 2694 8387 2698 8391
rect 2738 8387 2742 8391
rect 3318 8389 3322 8393
rect 3355 8387 3359 8391
rect 3375 8387 3379 8391
rect 3419 8387 3423 8391
rect 3450 8389 3454 8393
rect 3487 8387 3491 8391
rect 3507 8387 3511 8391
rect 3551 8387 3555 8391
rect 3582 8389 3586 8393
rect 3619 8387 3623 8391
rect 3639 8387 3643 8391
rect 3683 8387 3687 8391
rect 664 8379 668 8383
rect 674 8379 678 8383
rect 684 8379 688 8383
rect 2776 8380 2782 8384
rect 3721 8380 3727 8384
rect 2373 8373 2377 8377
rect 2424 8373 2428 8377
rect 2474 8373 2478 8377
rect 2505 8373 2509 8377
rect 2556 8373 2560 8377
rect 2606 8373 2610 8377
rect 2637 8373 2641 8377
rect 2688 8373 2692 8377
rect 2738 8373 2742 8377
rect 2812 8373 2818 8377
rect 3318 8373 3322 8377
rect 3369 8373 3373 8377
rect 3419 8373 3423 8377
rect 3450 8373 3454 8377
rect 3501 8373 3505 8377
rect 3551 8373 3555 8377
rect 3582 8373 3586 8377
rect 3633 8373 3637 8377
rect 3683 8373 3687 8377
rect 3757 8373 3763 8377
rect 2824 8365 2830 8369
rect 2857 8365 2861 8369
rect 2893 8365 2897 8369
rect 2960 8365 2964 8369
rect 2989 8365 2993 8369
rect 3025 8365 3029 8369
rect 3092 8365 3096 8369
rect 3121 8365 3125 8369
rect 3157 8365 3161 8369
rect 3224 8365 3228 8369
rect 3253 8365 3257 8369
rect 3289 8365 3293 8369
rect 3356 8365 3360 8369
rect 3769 8365 3775 8369
rect 3802 8365 3806 8369
rect 3838 8365 3842 8369
rect 3905 8365 3909 8369
rect 3934 8365 3938 8369
rect 3970 8365 3974 8369
rect 4037 8365 4041 8369
rect 4066 8365 4070 8369
rect 4102 8365 4106 8369
rect 4169 8365 4173 8369
rect 4198 8365 4202 8369
rect 4234 8365 4238 8369
rect 4301 8365 4305 8369
rect 2764 8358 2770 8362
rect 3709 8358 3715 8362
rect 2857 8351 2861 8355
rect 2907 8351 2911 8355
rect 2960 8351 2964 8355
rect 2989 8351 2993 8355
rect 3039 8351 3043 8355
rect 3092 8351 3096 8355
rect 3121 8351 3125 8355
rect 3171 8351 3175 8355
rect 3224 8351 3228 8355
rect 3253 8351 3257 8355
rect 3303 8351 3307 8355
rect 3356 8351 3360 8355
rect 3802 8351 3806 8355
rect 3852 8351 3856 8355
rect 3905 8351 3909 8355
rect 3934 8351 3938 8355
rect 3984 8351 3988 8355
rect 4037 8351 4041 8355
rect 4066 8351 4070 8355
rect 4116 8351 4120 8355
rect 4169 8351 4173 8355
rect 4198 8351 4202 8355
rect 4248 8351 4252 8355
rect 4301 8351 4305 8355
rect 2880 8340 2884 8344
rect 2505 8332 2509 8336
rect 2541 8332 2545 8336
rect 2608 8332 2612 8336
rect 2824 8332 2830 8336
rect 2851 8331 2855 8335
rect 2864 8334 2868 8340
rect 2901 8334 2905 8340
rect 2914 8336 2918 8340
rect 2938 8340 2942 8344
rect 3012 8340 3016 8344
rect 2922 8334 2926 8340
rect 2959 8334 2963 8340
rect 2975 8336 2979 8340
rect 2764 8325 2770 8329
rect 2505 8318 2509 8322
rect 2555 8318 2559 8322
rect 2608 8318 2612 8322
rect 2864 8321 2868 8325
rect 2880 8321 2884 8327
rect 2914 8327 2918 8331
rect 2901 8321 2905 8325
rect 2922 8321 2926 8325
rect 2938 8321 2942 8327
rect 2983 8331 2987 8335
rect 2996 8334 3000 8340
rect 3033 8334 3037 8340
rect 3046 8336 3050 8340
rect 3070 8340 3074 8344
rect 3144 8340 3148 8344
rect 3054 8334 3058 8340
rect 3091 8334 3095 8340
rect 3107 8336 3111 8340
rect 2959 8321 2963 8325
rect 2975 8321 2979 8325
rect 2996 8321 3000 8325
rect 3012 8321 3016 8327
rect 3046 8327 3050 8331
rect 3033 8321 3037 8325
rect 3054 8321 3058 8325
rect 3070 8321 3074 8327
rect 3115 8331 3119 8335
rect 3128 8334 3132 8340
rect 3165 8334 3169 8340
rect 3178 8336 3182 8340
rect 3202 8340 3206 8344
rect 3276 8340 3280 8344
rect 3186 8334 3190 8340
rect 3223 8334 3227 8340
rect 3239 8336 3243 8340
rect 3091 8321 3095 8325
rect 3107 8321 3111 8325
rect 3128 8321 3132 8325
rect 3144 8321 3148 8327
rect 3178 8327 3182 8331
rect 3165 8321 3169 8325
rect 3186 8321 3190 8325
rect 3202 8321 3206 8327
rect 3247 8331 3251 8335
rect 3260 8334 3264 8340
rect 3297 8334 3301 8340
rect 3310 8336 3314 8340
rect 3334 8340 3338 8344
rect 3825 8340 3829 8344
rect 3318 8334 3322 8340
rect 3355 8334 3359 8340
rect 3371 8336 3375 8340
rect 3450 8332 3454 8336
rect 3486 8332 3490 8336
rect 3553 8332 3557 8336
rect 3769 8332 3775 8336
rect 3223 8321 3227 8325
rect 3239 8321 3243 8325
rect 3260 8321 3264 8325
rect 3276 8321 3280 8327
rect 3310 8327 3314 8331
rect 3297 8321 3301 8325
rect 2528 8307 2532 8311
rect 2490 8298 2494 8302
rect 2512 8301 2516 8307
rect 2549 8301 2553 8307
rect 2562 8303 2566 8307
rect 2586 8307 2590 8311
rect 2570 8301 2574 8307
rect 2607 8301 2611 8307
rect 2623 8301 2627 8307
rect 2857 8310 2861 8314
rect 2894 8308 2898 8312
rect 2914 8308 2918 8312
rect 2958 8308 2962 8312
rect 2989 8310 2993 8314
rect 3026 8308 3030 8312
rect 3046 8308 3050 8312
rect 3090 8308 3094 8312
rect 3121 8310 3125 8314
rect 3158 8308 3162 8312
rect 3178 8308 3182 8312
rect 3222 8308 3226 8312
rect 3239 8313 3243 8317
rect 3318 8321 3322 8325
rect 3334 8321 3338 8327
rect 3796 8331 3800 8335
rect 3809 8334 3813 8340
rect 3846 8334 3850 8340
rect 3859 8336 3863 8340
rect 3883 8340 3887 8344
rect 3957 8340 3961 8344
rect 3867 8334 3871 8340
rect 3904 8334 3908 8340
rect 3920 8336 3924 8340
rect 3709 8325 3715 8329
rect 3355 8321 3359 8325
rect 3371 8321 3375 8325
rect 3253 8310 3257 8314
rect 3290 8308 3294 8312
rect 3310 8308 3314 8312
rect 3354 8308 3358 8312
rect 3371 8313 3375 8317
rect 3450 8318 3454 8322
rect 3500 8318 3504 8322
rect 3553 8318 3557 8322
rect 3809 8321 3813 8325
rect 3825 8321 3829 8327
rect 3859 8327 3863 8331
rect 3846 8321 3850 8325
rect 3867 8321 3871 8325
rect 3883 8321 3887 8327
rect 3928 8331 3932 8335
rect 3941 8334 3945 8340
rect 3978 8334 3982 8340
rect 3991 8336 3995 8340
rect 4015 8340 4019 8344
rect 4089 8340 4093 8344
rect 3999 8334 4003 8340
rect 4036 8334 4040 8340
rect 4052 8336 4056 8340
rect 3904 8321 3908 8325
rect 3920 8321 3924 8325
rect 3941 8321 3945 8325
rect 3957 8321 3961 8327
rect 3991 8327 3995 8331
rect 3978 8321 3982 8325
rect 3999 8321 4003 8325
rect 4015 8321 4019 8327
rect 4060 8331 4064 8335
rect 4073 8334 4077 8340
rect 4110 8334 4114 8340
rect 4123 8336 4127 8340
rect 4147 8340 4151 8344
rect 4221 8340 4225 8344
rect 4131 8334 4135 8340
rect 4168 8334 4172 8340
rect 4184 8336 4188 8340
rect 4036 8321 4040 8325
rect 4052 8321 4056 8325
rect 4073 8321 4077 8325
rect 4089 8321 4093 8327
rect 4123 8327 4127 8331
rect 4110 8321 4114 8325
rect 4131 8321 4135 8325
rect 4147 8321 4151 8327
rect 4192 8331 4196 8335
rect 4205 8334 4209 8340
rect 4242 8334 4246 8340
rect 4255 8336 4259 8340
rect 4279 8340 4283 8344
rect 4263 8334 4267 8340
rect 4300 8334 4304 8340
rect 4316 8336 4320 8340
rect 4168 8321 4172 8325
rect 4184 8321 4188 8325
rect 4205 8321 4209 8325
rect 4221 8321 4225 8327
rect 4255 8327 4259 8331
rect 4242 8321 4246 8325
rect 3473 8307 3477 8311
rect 2776 8301 2782 8305
rect 2512 8288 2516 8292
rect 2528 8288 2532 8294
rect 2562 8294 2566 8298
rect 2549 8288 2553 8292
rect 2570 8288 2574 8292
rect 2586 8288 2590 8294
rect 3435 8298 3439 8302
rect 3457 8301 3461 8307
rect 3494 8301 3498 8307
rect 3507 8303 3511 8307
rect 3531 8307 3535 8311
rect 3515 8301 3519 8307
rect 3552 8301 3556 8307
rect 3568 8301 3572 8307
rect 3802 8310 3806 8314
rect 3839 8308 3843 8312
rect 3859 8308 3863 8312
rect 3903 8308 3907 8312
rect 3934 8310 3938 8314
rect 3971 8308 3975 8312
rect 3991 8308 3995 8312
rect 4035 8308 4039 8312
rect 4066 8310 4070 8314
rect 4103 8308 4107 8312
rect 4123 8308 4127 8312
rect 4167 8308 4171 8312
rect 4184 8313 4188 8317
rect 4263 8321 4267 8325
rect 4279 8321 4283 8327
rect 4300 8321 4304 8325
rect 4316 8321 4320 8325
rect 4198 8310 4202 8314
rect 4235 8308 4239 8312
rect 4255 8308 4259 8312
rect 4299 8308 4303 8312
rect 4316 8313 4320 8317
rect 3721 8301 3727 8305
rect 2812 8294 2818 8298
rect 2857 8294 2861 8298
rect 2908 8294 2912 8298
rect 2958 8294 2962 8298
rect 2989 8294 2993 8298
rect 3040 8294 3044 8298
rect 3090 8294 3094 8298
rect 3121 8294 3125 8298
rect 3172 8294 3176 8298
rect 3222 8294 3226 8298
rect 3253 8294 3257 8298
rect 3304 8294 3308 8298
rect 3354 8294 3358 8298
rect 2607 8288 2611 8292
rect 2623 8288 2627 8292
rect 3457 8288 3461 8292
rect 3473 8288 3477 8294
rect 3507 8294 3511 8298
rect 3494 8288 3498 8292
rect 2505 8277 2509 8281
rect 2542 8275 2546 8279
rect 2562 8275 2566 8279
rect 2606 8275 2610 8279
rect 2764 8281 2770 8285
rect 2855 8281 2859 8285
rect 2889 8281 2893 8285
rect 2906 8281 2910 8285
rect 2962 8281 2966 8285
rect 2979 8281 2983 8285
rect 3007 8281 3011 8285
rect 3515 8288 3519 8292
rect 3531 8288 3535 8294
rect 3757 8294 3763 8298
rect 3802 8294 3806 8298
rect 3853 8294 3857 8298
rect 3903 8294 3907 8298
rect 3934 8294 3938 8298
rect 3985 8294 3989 8298
rect 4035 8294 4039 8298
rect 4066 8294 4070 8298
rect 4117 8294 4121 8298
rect 4167 8294 4171 8298
rect 4198 8294 4202 8298
rect 4249 8294 4253 8298
rect 4299 8294 4303 8298
rect 3552 8288 3556 8292
rect 3568 8288 3572 8292
rect 2800 8274 2806 8278
rect 2882 8274 2886 8278
rect 2913 8274 2917 8278
rect 2935 8274 2939 8278
rect 3000 8274 3004 8278
rect 2776 8268 2782 8272
rect 2505 8261 2509 8265
rect 2556 8261 2560 8265
rect 2606 8261 2610 8265
rect 2812 8261 2818 8265
rect 2856 8264 2860 8268
rect 2881 8267 2885 8271
rect 2888 8264 2892 8268
rect 2906 8264 2910 8268
rect 2928 8267 2932 8271
rect 2953 8267 2957 8271
rect 2963 8264 2967 8268
rect 2979 8264 2983 8268
rect 2999 8267 3003 8271
rect 3006 8264 3010 8268
rect 3070 8274 3074 8278
rect 2623 8254 2627 8258
rect 2490 8245 2494 8249
rect 2615 8247 2619 8251
rect 2639 8247 2643 8251
rect 2849 8247 2853 8251
rect 2498 8238 2502 8242
rect 2639 8238 2643 8242
rect 2883 8248 2887 8252
rect 2903 8245 2907 8249
rect 2922 8249 2926 8253
rect 3024 8260 3028 8264
rect 3039 8260 3043 8264
rect 2941 8248 2945 8252
rect 2960 8248 2964 8252
rect 2973 8247 2977 8251
rect 2995 8248 2999 8252
rect 3003 8247 3007 8251
rect 3015 8247 3019 8251
rect 2856 8234 2860 8238
rect 2888 8234 2892 8238
rect 2906 8234 2910 8238
rect 2963 8234 2967 8238
rect 2978 8234 2982 8238
rect 3006 8234 3010 8238
rect 2505 8230 2509 8234
rect 2572 8230 2576 8234
rect 2608 8230 2612 8234
rect 2824 8230 2830 8234
rect 2870 8230 2874 8234
rect 2913 8229 2917 8233
rect 2935 8230 2942 8234
rect 2985 8229 2989 8233
rect 2764 8223 2770 8227
rect 2505 8216 2509 8220
rect 2558 8216 2562 8220
rect 2608 8216 2612 8220
rect 2788 8222 2794 8226
rect 2870 8222 2874 8226
rect 2929 8222 2933 8226
rect 2954 8222 2958 8226
rect 2985 8222 2989 8226
rect 3078 8252 3082 8260
rect 3151 8274 3155 8278
rect 3105 8260 3109 8264
rect 3120 8260 3124 8264
rect 3450 8277 3454 8281
rect 3487 8275 3491 8279
rect 3507 8275 3511 8279
rect 3551 8275 3555 8279
rect 3709 8281 3715 8285
rect 3800 8281 3804 8285
rect 3834 8281 3838 8285
rect 3851 8281 3855 8285
rect 3907 8281 3911 8285
rect 3924 8281 3928 8285
rect 3952 8281 3956 8285
rect 3745 8274 3751 8278
rect 3827 8274 3831 8278
rect 3858 8274 3862 8278
rect 3880 8274 3884 8278
rect 3945 8274 3949 8278
rect 3101 8252 3105 8256
rect 3047 8246 3051 8250
rect 3060 8238 3064 8242
rect 3159 8252 3163 8260
rect 3721 8268 3727 8272
rect 3450 8261 3454 8265
rect 3501 8261 3505 8265
rect 3551 8261 3555 8265
rect 3757 8261 3763 8265
rect 3801 8264 3805 8268
rect 3826 8267 3830 8271
rect 3833 8264 3837 8268
rect 3851 8264 3855 8268
rect 3873 8267 3877 8271
rect 3898 8267 3902 8271
rect 3908 8264 3912 8268
rect 3924 8264 3928 8268
rect 3944 8267 3948 8271
rect 3951 8264 3955 8268
rect 4015 8274 4019 8278
rect 3186 8252 3190 8256
rect 3568 8254 3572 8258
rect 3128 8246 3132 8250
rect 3435 8245 3439 8249
rect 3560 8247 3564 8251
rect 3584 8247 3588 8251
rect 3794 8247 3798 8251
rect 3141 8238 3145 8242
rect 3443 8238 3447 8242
rect 3584 8238 3588 8242
rect 3828 8248 3832 8252
rect 3848 8245 3852 8249
rect 3867 8249 3871 8253
rect 3969 8260 3973 8264
rect 3984 8260 3988 8264
rect 3886 8248 3890 8252
rect 3905 8248 3909 8252
rect 3918 8247 3922 8251
rect 3940 8248 3944 8252
rect 3948 8247 3952 8251
rect 3960 8247 3964 8251
rect 3801 8234 3805 8238
rect 3833 8234 3837 8238
rect 3851 8234 3855 8238
rect 3908 8234 3912 8238
rect 3923 8234 3927 8238
rect 3951 8234 3955 8238
rect 3450 8230 3454 8234
rect 3517 8230 3521 8234
rect 3553 8230 3557 8234
rect 3769 8230 3775 8234
rect 3815 8230 3819 8234
rect 3858 8229 3862 8233
rect 3880 8230 3887 8234
rect 3930 8229 3934 8233
rect 3709 8223 3715 8227
rect 2776 8215 2782 8219
rect 2856 8215 2860 8219
rect 2870 8215 2874 8219
rect 2888 8215 2892 8219
rect 2906 8215 2910 8219
rect 2929 8215 2933 8219
rect 2963 8215 2967 8219
rect 2978 8215 2982 8219
rect 3006 8215 3010 8219
rect 2527 8205 2531 8209
rect 2490 8199 2494 8205
rect 2506 8199 2510 8205
rect 2543 8199 2547 8205
rect 2551 8201 2555 8205
rect 2585 8205 2589 8209
rect 2788 8208 2794 8212
rect 2870 8208 2874 8212
rect 2929 8208 2933 8212
rect 2954 8208 2958 8212
rect 2985 8208 2989 8212
rect 2564 8199 2568 8205
rect 2601 8199 2605 8205
rect 2870 8200 2874 8204
rect 2913 8201 2917 8205
rect 2935 8200 2942 8204
rect 2985 8201 2989 8205
rect 2623 8196 2627 8200
rect 2856 8196 2860 8200
rect 2888 8196 2892 8200
rect 2906 8196 2910 8200
rect 2963 8196 2967 8200
rect 2978 8196 2982 8200
rect 3006 8196 3010 8200
rect 2490 8186 2494 8190
rect 2506 8186 2510 8190
rect 2551 8192 2555 8196
rect 2527 8186 2531 8192
rect 2543 8186 2547 8190
rect 2564 8186 2568 8190
rect 2585 8186 2589 8192
rect 2601 8186 2605 8190
rect 2851 8184 2855 8188
rect 2507 8173 2511 8177
rect 2551 8173 2555 8177
rect 2571 8173 2575 8177
rect 2608 8175 2612 8179
rect 2883 8182 2887 8186
rect 2903 8185 2907 8189
rect 2922 8181 2926 8185
rect 2941 8182 2945 8186
rect 2960 8182 2964 8186
rect 2973 8183 2977 8187
rect 3070 8198 3074 8202
rect 3450 8216 3454 8220
rect 3503 8216 3507 8220
rect 3553 8216 3557 8220
rect 3733 8222 3739 8226
rect 3815 8222 3819 8226
rect 3874 8222 3878 8226
rect 3899 8222 3903 8226
rect 3930 8222 3934 8226
rect 4023 8252 4027 8260
rect 4096 8274 4100 8278
rect 4050 8260 4054 8264
rect 4065 8260 4069 8264
rect 4046 8252 4050 8256
rect 3992 8246 3996 8250
rect 4005 8238 4009 8242
rect 4104 8252 4108 8260
rect 4131 8252 4135 8256
rect 4073 8246 4077 8250
rect 4086 8238 4090 8242
rect 3721 8215 3727 8219
rect 3801 8215 3805 8219
rect 3815 8215 3819 8219
rect 3833 8215 3837 8219
rect 3851 8215 3855 8219
rect 3874 8215 3878 8219
rect 3908 8215 3912 8219
rect 3923 8215 3927 8219
rect 3951 8215 3955 8219
rect 3472 8205 3476 8209
rect 3151 8198 3155 8202
rect 3435 8199 3439 8205
rect 3451 8199 3455 8205
rect 3488 8199 3492 8205
rect 3496 8201 3500 8205
rect 3530 8205 3534 8209
rect 3733 8208 3739 8212
rect 3815 8208 3819 8212
rect 3874 8208 3878 8212
rect 3899 8208 3903 8212
rect 3930 8208 3934 8212
rect 3509 8199 3513 8205
rect 3546 8199 3550 8205
rect 3815 8200 3819 8204
rect 3858 8201 3862 8205
rect 3880 8200 3887 8204
rect 3930 8201 3934 8205
rect 3568 8196 3572 8200
rect 3801 8196 3805 8200
rect 3833 8196 3837 8200
rect 3851 8196 3855 8200
rect 3908 8196 3912 8200
rect 3923 8196 3927 8200
rect 3951 8196 3955 8200
rect 2995 8182 2999 8186
rect 3003 8183 3007 8187
rect 3015 8183 3019 8187
rect 3050 8183 3054 8187
rect 3078 8182 3082 8186
rect 3130 8183 3134 8187
rect 3435 8186 3439 8190
rect 3451 8186 3455 8190
rect 3496 8192 3500 8196
rect 3472 8186 3476 8192
rect 3488 8186 3492 8190
rect 3159 8182 3163 8186
rect 3509 8186 3513 8190
rect 3530 8186 3534 8192
rect 3546 8186 3550 8190
rect 3796 8184 3800 8188
rect 2776 8166 2782 8170
rect 2856 8166 2860 8170
rect 2881 8163 2885 8167
rect 2888 8166 2892 8170
rect 2906 8166 2910 8170
rect 2928 8163 2932 8167
rect 2953 8163 2957 8167
rect 2963 8166 2967 8170
rect 2979 8166 2983 8170
rect 2999 8163 3003 8167
rect 3006 8166 3010 8170
rect 2507 8159 2511 8163
rect 2557 8159 2561 8163
rect 2608 8159 2612 8163
rect 2812 8159 2818 8163
rect 2866 8156 2870 8160
rect 2882 8156 2886 8160
rect 2913 8156 2917 8160
rect 2935 8156 2939 8160
rect 3000 8156 3004 8160
rect 3060 8162 3064 8166
rect 3452 8173 3456 8177
rect 3496 8173 3500 8177
rect 3516 8173 3520 8177
rect 3553 8175 3557 8179
rect 3828 8182 3832 8186
rect 3848 8185 3852 8189
rect 3867 8181 3871 8185
rect 3886 8182 3890 8186
rect 3905 8182 3909 8186
rect 3918 8183 3922 8187
rect 4015 8198 4019 8202
rect 4096 8198 4100 8202
rect 3940 8182 3944 8186
rect 3948 8183 3952 8187
rect 3960 8183 3964 8187
rect 3995 8183 3999 8187
rect 4023 8182 4027 8186
rect 4075 8183 4079 8187
rect 4104 8182 4108 8186
rect 3721 8166 3727 8170
rect 3801 8166 3805 8170
rect 3141 8162 3145 8166
rect 3826 8163 3830 8167
rect 3833 8166 3837 8170
rect 3851 8166 3855 8170
rect 3873 8163 3877 8167
rect 3898 8163 3902 8167
rect 3908 8166 3912 8170
rect 3924 8166 3928 8170
rect 3944 8163 3948 8167
rect 3951 8166 3955 8170
rect 3452 8159 3456 8163
rect 3502 8159 3506 8163
rect 3553 8159 3557 8163
rect 3757 8159 3763 8163
rect 3811 8156 3815 8160
rect 3827 8156 3831 8160
rect 3858 8156 3862 8160
rect 3880 8156 3884 8160
rect 3945 8156 3949 8160
rect 4005 8162 4009 8166
rect 4086 8162 4090 8166
rect 2764 8149 2770 8153
rect 2855 8149 2859 8153
rect 2889 8149 2893 8153
rect 2906 8149 2910 8153
rect 2962 8149 2966 8153
rect 2979 8149 2983 8153
rect 3007 8149 3011 8153
rect 3709 8149 3715 8153
rect 3800 8149 3804 8153
rect 3834 8149 3838 8153
rect 3851 8149 3855 8153
rect 3907 8149 3911 8153
rect 3924 8149 3928 8153
rect 3952 8149 3956 8153
rect 2800 8142 2806 8146
rect 2866 8142 2870 8146
rect 2882 8142 2886 8146
rect 2913 8142 2917 8146
rect 2935 8142 2939 8146
rect 3000 8142 3004 8146
rect 3070 8142 3074 8146
rect 2856 8132 2860 8136
rect 2881 8135 2885 8139
rect 2888 8132 2892 8136
rect 2906 8132 2910 8136
rect 2928 8135 2932 8139
rect 2953 8135 2957 8139
rect 2963 8132 2967 8136
rect 2979 8132 2983 8136
rect 2999 8135 3003 8139
rect 3006 8132 3010 8136
rect 2850 8115 2854 8119
rect 2883 8116 2887 8120
rect 2903 8113 2907 8117
rect 2922 8117 2926 8121
rect 2941 8116 2945 8120
rect 2960 8116 2964 8120
rect 2973 8115 2977 8119
rect 2995 8116 2999 8120
rect 3003 8115 3007 8119
rect 3015 8115 3019 8119
rect 3078 8120 3082 8128
rect 3175 8142 3179 8146
rect 3129 8128 3133 8132
rect 3144 8128 3148 8132
rect 3745 8142 3751 8146
rect 3811 8142 3815 8146
rect 3827 8142 3831 8146
rect 3858 8142 3862 8146
rect 3880 8142 3884 8146
rect 3945 8142 3949 8146
rect 4015 8142 4019 8146
rect 3047 8114 3051 8118
rect 3101 8119 3105 8123
rect 2856 8102 2860 8106
rect 2888 8102 2892 8106
rect 2906 8102 2910 8106
rect 2963 8102 2967 8106
rect 2978 8102 2982 8106
rect 3006 8102 3010 8106
rect 2870 8098 2874 8102
rect 2913 8097 2917 8101
rect 2935 8098 2942 8102
rect 2985 8097 2989 8101
rect 2788 8090 2794 8094
rect 2870 8090 2874 8094
rect 2929 8090 2933 8094
rect 2954 8090 2958 8094
rect 2985 8090 2989 8094
rect 618 8085 622 8089
rect 628 8085 632 8089
rect 638 8085 642 8089
rect 618 8080 622 8084
rect 628 8080 632 8084
rect 638 8080 642 8084
rect 618 8075 622 8079
rect 628 8075 632 8079
rect 638 8075 642 8079
rect 618 8070 622 8074
rect 628 8070 632 8074
rect 638 8070 642 8074
rect 664 8085 668 8089
rect 674 8085 678 8089
rect 684 8085 688 8089
rect 3060 8106 3064 8110
rect 3183 8120 3187 8128
rect 3801 8132 3805 8136
rect 3826 8135 3830 8139
rect 3833 8132 3837 8136
rect 3851 8132 3855 8136
rect 3873 8135 3877 8139
rect 3898 8135 3902 8139
rect 3908 8132 3912 8136
rect 3924 8132 3928 8136
rect 3944 8135 3948 8139
rect 3951 8132 3955 8136
rect 3204 8120 3208 8124
rect 3152 8114 3156 8118
rect 3795 8115 3799 8119
rect 3165 8106 3169 8110
rect 3828 8116 3832 8120
rect 3848 8113 3852 8117
rect 3867 8117 3871 8121
rect 3886 8116 3890 8120
rect 3905 8116 3909 8120
rect 3918 8115 3922 8119
rect 3940 8116 3944 8120
rect 3948 8115 3952 8119
rect 3960 8115 3964 8119
rect 4023 8120 4027 8128
rect 4120 8142 4124 8146
rect 4074 8128 4078 8132
rect 4089 8128 4093 8132
rect 3992 8114 3996 8118
rect 4046 8119 4050 8123
rect 3801 8102 3805 8106
rect 3833 8102 3837 8106
rect 3851 8102 3855 8106
rect 3908 8102 3912 8106
rect 3923 8102 3927 8106
rect 3951 8102 3955 8106
rect 3815 8098 3819 8102
rect 3858 8097 3862 8101
rect 3880 8098 3887 8102
rect 3930 8097 3934 8101
rect 3733 8090 3739 8094
rect 3815 8090 3819 8094
rect 3874 8090 3878 8094
rect 3899 8090 3903 8094
rect 3930 8090 3934 8094
rect 4005 8106 4009 8110
rect 4128 8120 4132 8128
rect 4484 8129 4488 8133
rect 4494 8129 4498 8133
rect 4504 8129 4508 8133
rect 4484 8124 4488 8128
rect 4494 8124 4498 8128
rect 4504 8124 4508 8128
rect 4149 8120 4153 8124
rect 4097 8114 4101 8118
rect 4484 8119 4488 8123
rect 4494 8119 4498 8123
rect 4504 8119 4508 8123
rect 4484 8114 4488 8118
rect 4494 8114 4498 8118
rect 4504 8114 4508 8118
rect 4530 8129 4534 8133
rect 4540 8129 4544 8133
rect 4550 8129 4554 8133
rect 4530 8124 4534 8128
rect 4540 8124 4544 8128
rect 4550 8124 4554 8128
rect 4530 8119 4534 8123
rect 4540 8119 4544 8123
rect 4550 8119 4554 8123
rect 4530 8114 4534 8118
rect 4540 8114 4544 8118
rect 4550 8114 4554 8118
rect 4110 8106 4114 8110
rect 4484 8098 4488 8102
rect 4494 8098 4498 8102
rect 4504 8098 4508 8102
rect 4484 8093 4488 8097
rect 4494 8093 4498 8097
rect 4504 8093 4508 8097
rect 4484 8088 4488 8092
rect 4494 8088 4498 8092
rect 4504 8088 4508 8092
rect 664 8080 668 8084
rect 674 8080 678 8084
rect 684 8080 688 8084
rect 2776 8083 2782 8087
rect 2856 8083 2860 8087
rect 2870 8083 2874 8087
rect 2888 8083 2892 8087
rect 2906 8083 2910 8087
rect 2929 8083 2933 8087
rect 2963 8083 2967 8087
rect 2978 8083 2982 8087
rect 3006 8083 3010 8087
rect 3721 8083 3727 8087
rect 3801 8083 3805 8087
rect 3815 8083 3819 8087
rect 3833 8083 3837 8087
rect 3851 8083 3855 8087
rect 3874 8083 3878 8087
rect 3908 8083 3912 8087
rect 3923 8083 3927 8087
rect 3951 8083 3955 8087
rect 4484 8083 4488 8087
rect 4494 8083 4498 8087
rect 4504 8083 4508 8087
rect 4530 8098 4534 8102
rect 4540 8098 4544 8102
rect 4550 8098 4554 8102
rect 4530 8093 4534 8097
rect 4540 8093 4544 8097
rect 4550 8093 4554 8097
rect 4530 8088 4534 8092
rect 4540 8088 4544 8092
rect 4550 8088 4554 8092
rect 4530 8083 4534 8087
rect 4540 8083 4544 8087
rect 4550 8083 4554 8087
rect 664 8075 668 8079
rect 674 8075 678 8079
rect 684 8075 688 8079
rect 2788 8076 2794 8080
rect 2870 8076 2874 8080
rect 2929 8076 2933 8080
rect 2954 8076 2958 8080
rect 2985 8076 2989 8080
rect 664 8070 668 8074
rect 674 8070 678 8074
rect 684 8070 688 8074
rect 2870 8068 2874 8072
rect 2913 8069 2917 8073
rect 2935 8068 2942 8072
rect 2985 8069 2989 8073
rect 2856 8064 2860 8068
rect 2888 8064 2892 8068
rect 2906 8064 2910 8068
rect 2963 8064 2967 8068
rect 2978 8064 2982 8068
rect 3006 8064 3010 8068
rect 3070 8067 3074 8071
rect 3733 8076 3739 8080
rect 3815 8076 3819 8080
rect 3874 8076 3878 8080
rect 3899 8076 3903 8080
rect 3930 8076 3934 8080
rect 3175 8067 3179 8071
rect 3815 8068 3819 8072
rect 3858 8069 3862 8073
rect 3880 8068 3887 8072
rect 3930 8069 3934 8073
rect 3801 8064 3805 8068
rect 3833 8064 3837 8068
rect 3851 8064 3855 8068
rect 3908 8064 3912 8068
rect 3923 8064 3927 8068
rect 3951 8064 3955 8068
rect 4015 8067 4019 8071
rect 4506 8074 4510 8078
rect 4511 8074 4515 8078
rect 4120 8067 4124 8071
rect 4506 8069 4510 8073
rect 4511 8069 4515 8073
rect 4506 8064 4510 8068
rect 4511 8064 4515 8068
rect 2851 8052 2855 8056
rect 2883 8050 2887 8054
rect 2903 8053 2907 8057
rect 2922 8049 2926 8053
rect 2941 8050 2945 8054
rect 2960 8050 2964 8054
rect 2973 8051 2977 8055
rect 2995 8050 2999 8054
rect 3003 8051 3007 8055
rect 3015 8051 3019 8055
rect 3049 8052 3053 8056
rect 3078 8051 3082 8055
rect 3155 8052 3159 8056
rect 3183 8051 3187 8055
rect 3796 8052 3800 8056
rect 2856 8034 2860 8038
rect 2881 8031 2885 8035
rect 2888 8034 2892 8038
rect 2906 8034 2910 8038
rect 2928 8031 2932 8035
rect 2953 8031 2957 8035
rect 2963 8034 2967 8038
rect 2979 8034 2983 8038
rect 2999 8031 3003 8035
rect 3006 8034 3010 8038
rect 2800 8024 2806 8028
rect 2882 8024 2886 8028
rect 2913 8024 2917 8028
rect 2935 8024 2939 8028
rect 3000 8024 3004 8028
rect 3060 8031 3064 8035
rect 3828 8050 3832 8054
rect 3848 8053 3852 8057
rect 3867 8049 3871 8053
rect 3886 8050 3890 8054
rect 3905 8050 3909 8054
rect 3918 8051 3922 8055
rect 3940 8050 3944 8054
rect 3948 8051 3952 8055
rect 3960 8051 3964 8055
rect 3994 8052 3998 8056
rect 4023 8051 4027 8055
rect 4100 8052 4104 8056
rect 4506 8059 4510 8063
rect 4511 8059 4515 8063
rect 4128 8051 4132 8055
rect 4506 8054 4510 8058
rect 4511 8054 4515 8058
rect 4506 8049 4510 8053
rect 4511 8049 4515 8053
rect 4506 8044 4510 8048
rect 4511 8044 4515 8048
rect 3165 8031 3169 8035
rect 3801 8034 3805 8038
rect 3826 8031 3830 8035
rect 3833 8034 3837 8038
rect 3851 8034 3855 8038
rect 3873 8031 3877 8035
rect 3898 8031 3902 8035
rect 3908 8034 3912 8038
rect 3924 8034 3928 8038
rect 3944 8031 3948 8035
rect 3951 8034 3955 8038
rect 3745 8024 3751 8028
rect 3827 8024 3831 8028
rect 3858 8024 3862 8028
rect 3880 8024 3884 8028
rect 3945 8024 3949 8028
rect 4005 8031 4009 8035
rect 4506 8039 4510 8043
rect 4511 8039 4515 8043
rect 4110 8031 4114 8035
rect 4506 8034 4510 8038
rect 4511 8034 4515 8038
rect 4506 8029 4510 8033
rect 4511 8029 4515 8033
rect 4506 8024 4510 8028
rect 4511 8024 4515 8028
rect 2764 8017 2770 8021
rect 2855 8017 2859 8021
rect 2889 8017 2893 8021
rect 2906 8017 2910 8021
rect 2962 8017 2966 8021
rect 2979 8017 2983 8021
rect 3007 8017 3011 8021
rect 3709 8017 3715 8021
rect 3800 8017 3804 8021
rect 3834 8017 3838 8021
rect 3851 8017 3855 8021
rect 3907 8017 3911 8021
rect 3924 8017 3928 8021
rect 3952 8017 3956 8021
rect 2800 8010 2806 8014
rect 2882 8010 2886 8014
rect 2913 8010 2917 8014
rect 2935 8010 2939 8014
rect 3000 8010 3004 8014
rect 3070 8010 3074 8014
rect 2856 8000 2860 8004
rect 2881 8003 2885 8007
rect 2888 8000 2892 8004
rect 2906 8000 2910 8004
rect 2928 8003 2932 8007
rect 2953 8003 2957 8007
rect 2963 8000 2967 8004
rect 2979 8000 2983 8004
rect 2999 8003 3003 8007
rect 3006 8000 3010 8004
rect 2850 7983 2854 7987
rect 2883 7984 2887 7988
rect 2903 7981 2907 7985
rect 2922 7985 2926 7989
rect 2941 7984 2945 7988
rect 2960 7984 2964 7988
rect 2973 7983 2977 7987
rect 2995 7984 2999 7988
rect 3003 7983 3007 7987
rect 3015 7983 3019 7987
rect 3078 7988 3082 7996
rect 3151 8010 3155 8014
rect 3105 7996 3109 8000
rect 3120 7996 3124 8000
rect 3101 7988 3105 7992
rect 3047 7982 3051 7986
rect 2856 7970 2860 7974
rect 2888 7970 2892 7974
rect 2906 7970 2910 7974
rect 2963 7970 2967 7974
rect 2978 7970 2982 7974
rect 3006 7970 3010 7974
rect 2870 7966 2874 7970
rect 2913 7965 2917 7969
rect 2935 7966 2942 7970
rect 2985 7965 2989 7969
rect 2788 7958 2794 7962
rect 2870 7958 2874 7962
rect 2929 7958 2933 7962
rect 2954 7958 2958 7962
rect 2985 7958 2989 7962
rect 3060 7974 3064 7978
rect 3159 7988 3163 7996
rect 3241 8010 3245 8014
rect 3195 7996 3199 8000
rect 3210 7996 3214 8000
rect 3745 8010 3751 8014
rect 3827 8010 3831 8014
rect 3858 8010 3862 8014
rect 3880 8010 3884 8014
rect 3945 8010 3949 8014
rect 4015 8010 4019 8014
rect 3183 7988 3187 7992
rect 3128 7982 3132 7986
rect 3217 7990 3221 7994
rect 3249 7988 3253 7996
rect 3801 8000 3805 8004
rect 3826 8003 3830 8007
rect 3833 8000 3837 8004
rect 3851 8000 3855 8004
rect 3873 8003 3877 8007
rect 3898 8003 3902 8007
rect 3908 8000 3912 8004
rect 3924 8000 3928 8004
rect 3944 8003 3948 8007
rect 3951 8000 3955 8004
rect 3141 7974 3145 7978
rect 3284 7987 3288 7991
rect 3795 7983 3799 7987
rect 3231 7974 3235 7978
rect 3828 7984 3832 7988
rect 3848 7981 3852 7985
rect 3867 7985 3871 7989
rect 3886 7984 3890 7988
rect 3905 7984 3909 7988
rect 3918 7983 3922 7987
rect 3940 7984 3944 7988
rect 3948 7983 3952 7987
rect 3960 7983 3964 7987
rect 4023 7988 4027 7996
rect 4096 8010 4100 8014
rect 4050 7996 4054 8000
rect 4065 7996 4069 8000
rect 4046 7988 4050 7992
rect 3992 7982 3996 7986
rect 3801 7970 3805 7974
rect 3833 7970 3837 7974
rect 3851 7970 3855 7974
rect 3908 7970 3912 7974
rect 3923 7970 3927 7974
rect 3951 7970 3955 7974
rect 3815 7966 3819 7970
rect 3858 7965 3862 7969
rect 3880 7966 3887 7970
rect 3930 7965 3934 7969
rect 3733 7958 3739 7962
rect 3815 7958 3819 7962
rect 3874 7958 3878 7962
rect 3899 7958 3903 7962
rect 3930 7958 3934 7962
rect 4005 7974 4009 7978
rect 4104 7988 4108 7996
rect 4186 8010 4190 8014
rect 4140 7996 4144 8000
rect 4155 7996 4159 8000
rect 4128 7988 4132 7992
rect 4073 7982 4077 7986
rect 4162 7990 4166 7994
rect 4194 7988 4198 7996
rect 4086 7974 4090 7978
rect 4229 7987 4233 7991
rect 4377 7987 4386 7992
rect 4574 7982 4578 7986
rect 4176 7974 4180 7978
rect 4590 7982 4594 7986
rect 4606 7982 4610 7986
rect 4622 7982 4626 7986
rect 4645 7982 4649 7986
rect 4661 7982 4665 7986
rect 4688 7982 4692 7986
rect 4704 7982 4708 7986
rect 4729 7982 4733 7986
rect 4745 7982 4749 7986
rect 2776 7951 2782 7955
rect 2856 7951 2860 7955
rect 2870 7951 2874 7955
rect 2888 7951 2892 7955
rect 2906 7951 2910 7955
rect 2929 7951 2933 7955
rect 2963 7951 2967 7955
rect 2978 7951 2982 7955
rect 3006 7951 3010 7955
rect 3721 7951 3727 7955
rect 3801 7951 3805 7955
rect 3815 7951 3819 7955
rect 3833 7951 3837 7955
rect 3851 7951 3855 7955
rect 3874 7951 3878 7955
rect 3908 7951 3912 7955
rect 3923 7951 3927 7955
rect 3951 7951 3955 7955
rect 2788 7944 2794 7948
rect 2870 7944 2874 7948
rect 2929 7944 2933 7948
rect 2954 7944 2958 7948
rect 2985 7944 2989 7948
rect 2870 7936 2874 7940
rect 2913 7937 2917 7941
rect 2935 7936 2942 7940
rect 2985 7937 2989 7941
rect 2856 7932 2860 7936
rect 2888 7932 2892 7936
rect 2906 7932 2910 7936
rect 2963 7932 2967 7936
rect 2978 7932 2982 7936
rect 3006 7932 3010 7936
rect 2851 7920 2855 7924
rect 2883 7918 2887 7922
rect 2903 7921 2907 7925
rect 2922 7917 2926 7921
rect 2941 7918 2945 7922
rect 2960 7918 2964 7922
rect 2973 7919 2977 7923
rect 3070 7932 3074 7936
rect 3151 7932 3155 7936
rect 3733 7944 3739 7948
rect 3815 7944 3819 7948
rect 3874 7944 3878 7948
rect 3899 7944 3903 7948
rect 3930 7944 3934 7948
rect 3815 7936 3819 7940
rect 3858 7937 3862 7941
rect 3880 7936 3887 7940
rect 3930 7937 3934 7941
rect 3241 7932 3245 7936
rect 3801 7932 3805 7936
rect 3833 7932 3837 7936
rect 3851 7932 3855 7936
rect 3908 7932 3912 7936
rect 3923 7932 3927 7936
rect 3951 7932 3955 7936
rect 2995 7918 2999 7922
rect 3003 7919 3007 7923
rect 3015 7919 3019 7923
rect 3050 7917 3054 7921
rect 3078 7916 3082 7920
rect 3130 7917 3134 7921
rect 3159 7916 3163 7920
rect 3214 7917 3218 7921
rect 3796 7920 3800 7924
rect 3249 7916 3253 7920
rect 2856 7902 2860 7906
rect 2881 7899 2885 7903
rect 2888 7902 2892 7906
rect 2906 7902 2910 7906
rect 2928 7899 2932 7903
rect 2953 7899 2957 7903
rect 2963 7902 2967 7906
rect 2979 7902 2983 7906
rect 2999 7899 3003 7903
rect 3006 7902 3010 7906
rect 3828 7918 3832 7922
rect 3848 7921 3852 7925
rect 3867 7917 3871 7921
rect 3886 7918 3890 7922
rect 3905 7918 3909 7922
rect 3918 7919 3922 7923
rect 4015 7932 4019 7936
rect 4096 7932 4100 7936
rect 4377 7950 4386 7963
rect 4659 7954 4667 7963
rect 4703 7954 4711 7963
rect 4186 7932 4190 7936
rect 3940 7918 3944 7922
rect 3948 7919 3952 7923
rect 3960 7919 3964 7923
rect 3995 7917 3999 7921
rect 4023 7916 4027 7920
rect 4075 7917 4079 7921
rect 4104 7916 4108 7920
rect 4159 7917 4163 7921
rect 4574 7924 4578 7928
rect 4194 7916 4198 7920
rect 2800 7892 2806 7896
rect 2882 7892 2886 7896
rect 2913 7892 2917 7896
rect 2935 7892 2939 7896
rect 3000 7892 3004 7896
rect 3060 7896 3064 7900
rect 3141 7896 3145 7900
rect 3801 7902 3805 7906
rect 3231 7896 3235 7900
rect 3826 7899 3830 7903
rect 3833 7902 3837 7906
rect 3851 7902 3855 7906
rect 3873 7899 3877 7903
rect 3898 7899 3902 7903
rect 3908 7902 3912 7906
rect 3924 7902 3928 7906
rect 3944 7899 3948 7903
rect 3951 7902 3955 7906
rect 3745 7892 3751 7896
rect 3827 7892 3831 7896
rect 3858 7892 3862 7896
rect 3880 7892 3884 7896
rect 3945 7892 3949 7896
rect 4005 7896 4009 7900
rect 4086 7896 4090 7900
rect 4176 7896 4180 7900
rect 4590 7924 4594 7928
rect 4606 7924 4610 7928
rect 4622 7924 4626 7928
rect 2764 7885 2770 7889
rect 2855 7885 2859 7889
rect 2889 7885 2893 7889
rect 2906 7885 2910 7889
rect 2962 7885 2966 7889
rect 2979 7885 2983 7889
rect 3007 7885 3011 7889
rect 3709 7885 3715 7889
rect 3800 7885 3804 7889
rect 3834 7885 3838 7889
rect 3851 7885 3855 7889
rect 3907 7885 3911 7889
rect 3924 7885 3928 7889
rect 3952 7885 3956 7889
rect 2800 7878 2806 7882
rect 2882 7878 2886 7882
rect 2913 7878 2917 7882
rect 2935 7878 2939 7882
rect 3000 7878 3004 7882
rect 3070 7878 3074 7882
rect 2856 7868 2860 7872
rect 2881 7871 2885 7875
rect 2888 7868 2892 7872
rect 2906 7868 2910 7872
rect 2928 7871 2932 7875
rect 2953 7871 2957 7875
rect 2963 7868 2967 7872
rect 2979 7868 2983 7872
rect 2999 7871 3003 7875
rect 3006 7868 3010 7872
rect 2850 7851 2854 7855
rect 2883 7852 2887 7856
rect 2903 7849 2907 7853
rect 2922 7853 2926 7857
rect 3745 7878 3751 7882
rect 3827 7878 3831 7882
rect 3858 7878 3862 7882
rect 3880 7878 3884 7882
rect 3945 7878 3949 7882
rect 4015 7878 4019 7882
rect 2941 7852 2945 7856
rect 2960 7852 2964 7856
rect 2973 7851 2977 7855
rect 2995 7852 2999 7856
rect 3003 7851 3007 7855
rect 3015 7851 3019 7855
rect 3078 7856 3082 7864
rect 3801 7868 3805 7872
rect 3826 7871 3830 7875
rect 3833 7868 3837 7872
rect 3851 7868 3855 7872
rect 3873 7871 3877 7875
rect 3898 7871 3902 7875
rect 3908 7868 3912 7872
rect 3924 7868 3928 7872
rect 3944 7871 3948 7875
rect 3951 7868 3955 7872
rect 3047 7850 3051 7854
rect 3101 7855 3105 7859
rect 3795 7851 3799 7855
rect 2856 7838 2860 7842
rect 2888 7838 2892 7842
rect 2906 7838 2910 7842
rect 2963 7838 2967 7842
rect 2978 7838 2982 7842
rect 3006 7838 3010 7842
rect 2870 7834 2874 7838
rect 2373 7830 2377 7834
rect 2409 7830 2413 7834
rect 2476 7830 2480 7834
rect 2505 7830 2509 7834
rect 2541 7830 2545 7834
rect 2608 7830 2612 7834
rect 2637 7830 2641 7834
rect 2673 7830 2677 7834
rect 2740 7830 2744 7834
rect 2824 7830 2830 7834
rect 2913 7833 2917 7837
rect 2935 7834 2942 7838
rect 2985 7833 2989 7837
rect 2764 7823 2770 7827
rect 2870 7826 2874 7830
rect 2879 7826 2883 7830
rect 2929 7826 2933 7830
rect 2954 7826 2958 7830
rect 2985 7826 2989 7830
rect 3060 7842 3064 7846
rect 3828 7852 3832 7856
rect 3848 7849 3852 7853
rect 3867 7853 3871 7857
rect 3886 7852 3890 7856
rect 3905 7852 3909 7856
rect 3918 7851 3922 7855
rect 3940 7852 3944 7856
rect 3948 7851 3952 7855
rect 3960 7851 3964 7855
rect 4023 7856 4027 7864
rect 3992 7850 3996 7854
rect 4046 7855 4050 7859
rect 3801 7838 3805 7842
rect 3833 7838 3837 7842
rect 3851 7838 3855 7842
rect 3908 7838 3912 7842
rect 3923 7838 3927 7842
rect 3951 7838 3955 7842
rect 3815 7834 3819 7838
rect 3318 7830 3322 7834
rect 3354 7830 3358 7834
rect 3421 7830 3425 7834
rect 3450 7830 3454 7834
rect 3486 7830 3490 7834
rect 3553 7830 3557 7834
rect 3582 7830 3586 7834
rect 3618 7830 3622 7834
rect 3685 7830 3689 7834
rect 3769 7830 3775 7834
rect 3858 7833 3862 7837
rect 3880 7834 3887 7838
rect 3930 7833 3934 7837
rect 3709 7823 3715 7827
rect 3815 7826 3819 7830
rect 3824 7826 3828 7830
rect 3874 7826 3878 7830
rect 3899 7826 3903 7830
rect 3930 7826 3934 7830
rect 4645 7924 4649 7928
rect 4661 7924 4665 7928
rect 4688 7924 4692 7928
rect 4704 7924 4708 7928
rect 4729 7924 4733 7928
rect 4745 7924 4749 7928
rect 4005 7842 4009 7846
rect 4529 7824 4533 7828
rect 4534 7824 4538 7828
rect 4539 7824 4543 7828
rect 4544 7824 4548 7828
rect 4549 7824 4553 7828
rect 4554 7824 4558 7828
rect 4559 7824 4563 7828
rect 4564 7824 4568 7828
rect 4569 7824 4573 7828
rect 4574 7824 4578 7828
rect 4579 7824 4583 7828
rect 4584 7824 4588 7828
rect 4589 7824 4593 7828
rect 2373 7816 2377 7820
rect 2423 7816 2427 7820
rect 2476 7816 2480 7820
rect 2505 7816 2509 7820
rect 2555 7816 2559 7820
rect 2608 7816 2612 7820
rect 2637 7816 2641 7820
rect 2687 7816 2691 7820
rect 2740 7816 2744 7820
rect 2776 7819 2782 7823
rect 2856 7819 2860 7823
rect 2870 7819 2874 7823
rect 2888 7819 2892 7823
rect 2906 7819 2910 7823
rect 2929 7819 2933 7823
rect 2963 7819 2967 7823
rect 2978 7819 2982 7823
rect 3006 7819 3010 7823
rect 3131 7819 3135 7823
rect 3149 7819 3153 7823
rect 3167 7819 3171 7823
rect 3190 7819 3194 7823
rect 3224 7819 3228 7823
rect 3239 7819 3243 7823
rect 3267 7819 3271 7823
rect 2396 7805 2400 7809
rect 2367 7796 2371 7800
rect 2380 7799 2384 7805
rect 2417 7799 2421 7805
rect 2430 7801 2434 7805
rect 2454 7805 2458 7809
rect 2528 7805 2532 7809
rect 2438 7799 2442 7805
rect 2475 7799 2479 7805
rect 2491 7799 2495 7805
rect 2512 7799 2516 7805
rect 2549 7799 2553 7805
rect 2562 7801 2566 7805
rect 2586 7805 2590 7809
rect 2660 7805 2664 7809
rect 2570 7799 2574 7805
rect 2607 7799 2611 7805
rect 2623 7799 2627 7805
rect 2644 7799 2648 7805
rect 2681 7799 2685 7805
rect 2694 7801 2698 7805
rect 2718 7805 2722 7809
rect 2788 7812 2794 7816
rect 2870 7812 2874 7816
rect 2879 7812 2883 7816
rect 2929 7812 2933 7816
rect 2954 7812 2958 7816
rect 2985 7812 2989 7816
rect 2702 7799 2706 7805
rect 2739 7799 2743 7805
rect 2755 7801 2759 7805
rect 2870 7804 2874 7808
rect 2913 7805 2917 7809
rect 2935 7804 2942 7808
rect 2985 7805 2989 7809
rect 2856 7800 2860 7804
rect 2888 7800 2892 7804
rect 2906 7800 2910 7804
rect 2963 7800 2967 7804
rect 2978 7800 2982 7804
rect 3006 7800 3010 7804
rect 2380 7786 2384 7790
rect 2396 7786 2400 7792
rect 2430 7792 2434 7796
rect 2417 7786 2421 7790
rect 2438 7786 2442 7790
rect 2454 7786 2458 7792
rect 2475 7786 2479 7790
rect 2491 7786 2495 7790
rect 2512 7786 2516 7790
rect 2528 7786 2532 7792
rect 2562 7792 2566 7796
rect 2549 7786 2553 7790
rect 2570 7786 2574 7790
rect 2586 7786 2590 7792
rect 2607 7786 2611 7790
rect 2623 7786 2627 7790
rect 2644 7786 2648 7790
rect 2660 7786 2664 7792
rect 2694 7792 2698 7796
rect 2681 7786 2685 7790
rect 2702 7786 2706 7790
rect 2718 7786 2722 7792
rect 2739 7786 2743 7790
rect 2755 7786 2759 7790
rect 2851 7788 2855 7792
rect 618 7776 622 7780
rect 628 7776 632 7780
rect 638 7776 642 7780
rect 618 7771 622 7775
rect 628 7771 632 7775
rect 638 7771 642 7775
rect 618 7766 622 7770
rect 628 7766 632 7770
rect 638 7766 642 7770
rect 618 7761 622 7765
rect 628 7761 632 7765
rect 638 7761 642 7765
rect 664 7776 668 7780
rect 674 7776 678 7780
rect 684 7776 688 7780
rect 664 7771 668 7775
rect 674 7771 678 7775
rect 684 7771 688 7775
rect 2373 7775 2377 7779
rect 2410 7773 2414 7777
rect 2430 7773 2434 7777
rect 2474 7773 2478 7777
rect 2505 7775 2509 7779
rect 2542 7773 2546 7777
rect 2562 7773 2566 7777
rect 2606 7773 2610 7777
rect 2637 7775 2641 7779
rect 2674 7773 2678 7777
rect 2694 7773 2698 7777
rect 2738 7773 2742 7777
rect 2883 7786 2887 7790
rect 2903 7789 2907 7793
rect 2922 7785 2926 7789
rect 2941 7786 2945 7790
rect 2960 7786 2964 7790
rect 2973 7787 2977 7791
rect 3109 7812 3113 7816
rect 3131 7812 3135 7816
rect 3190 7812 3194 7816
rect 3215 7812 3219 7816
rect 3246 7812 3250 7816
rect 3318 7816 3322 7820
rect 3368 7816 3372 7820
rect 3421 7816 3425 7820
rect 3450 7816 3454 7820
rect 3500 7816 3504 7820
rect 3553 7816 3557 7820
rect 3582 7816 3586 7820
rect 3632 7816 3636 7820
rect 3685 7816 3689 7820
rect 3721 7819 3727 7823
rect 3801 7819 3805 7823
rect 3815 7819 3819 7823
rect 3833 7819 3837 7823
rect 3851 7819 3855 7823
rect 3874 7819 3878 7823
rect 3908 7819 3912 7823
rect 3923 7819 3927 7823
rect 3951 7819 3955 7823
rect 4076 7819 4080 7823
rect 4094 7819 4098 7823
rect 4112 7819 4116 7823
rect 4135 7819 4139 7823
rect 4169 7819 4173 7823
rect 4184 7819 4188 7823
rect 4212 7819 4216 7823
rect 4529 7819 4533 7823
rect 4534 7819 4538 7823
rect 4539 7819 4543 7823
rect 4544 7819 4548 7823
rect 4549 7819 4553 7823
rect 4554 7819 4558 7823
rect 4559 7819 4563 7823
rect 4564 7819 4568 7823
rect 4569 7819 4573 7823
rect 4574 7819 4578 7823
rect 4579 7819 4583 7823
rect 4584 7819 4588 7823
rect 4589 7819 4593 7823
rect 3131 7804 3135 7808
rect 3174 7805 3178 7809
rect 3196 7804 3203 7808
rect 3246 7805 3250 7809
rect 3341 7805 3345 7809
rect 3149 7800 3153 7804
rect 3167 7800 3171 7804
rect 3224 7800 3228 7804
rect 3239 7800 3243 7804
rect 3267 7800 3271 7804
rect 3070 7796 3074 7800
rect 2995 7786 2999 7790
rect 3003 7787 3007 7791
rect 3015 7787 3019 7791
rect 3049 7781 3053 7785
rect 3089 7787 3093 7791
rect 3078 7780 3082 7784
rect 2856 7770 2860 7774
rect 664 7766 668 7770
rect 674 7766 678 7770
rect 684 7766 688 7770
rect 2776 7766 2782 7770
rect 2881 7767 2885 7771
rect 2888 7770 2892 7774
rect 2906 7770 2910 7774
rect 2928 7767 2932 7771
rect 2953 7767 2957 7771
rect 2963 7770 2967 7774
rect 2979 7770 2983 7774
rect 2999 7767 3003 7771
rect 3006 7770 3010 7774
rect 3144 7786 3148 7790
rect 3164 7789 3168 7793
rect 3183 7785 3187 7789
rect 3312 7796 3316 7800
rect 3325 7799 3329 7805
rect 3362 7799 3366 7805
rect 3375 7801 3379 7805
rect 3399 7805 3403 7809
rect 3473 7805 3477 7809
rect 3383 7799 3387 7805
rect 3420 7799 3424 7805
rect 3436 7799 3440 7805
rect 3457 7799 3461 7805
rect 3494 7799 3498 7805
rect 3507 7801 3511 7805
rect 3531 7805 3535 7809
rect 3605 7805 3609 7809
rect 3515 7799 3519 7805
rect 3552 7799 3556 7805
rect 3568 7799 3572 7805
rect 3589 7799 3593 7805
rect 3626 7799 3630 7805
rect 3639 7801 3643 7805
rect 3663 7805 3667 7809
rect 3733 7812 3739 7816
rect 3815 7812 3819 7816
rect 3824 7812 3828 7816
rect 3874 7812 3878 7816
rect 3899 7812 3903 7816
rect 3930 7812 3934 7816
rect 3647 7799 3651 7805
rect 3684 7799 3688 7805
rect 3700 7801 3704 7805
rect 3815 7804 3819 7808
rect 3858 7805 3862 7809
rect 3880 7804 3887 7808
rect 3930 7805 3934 7809
rect 3801 7800 3805 7804
rect 3833 7800 3837 7804
rect 3851 7800 3855 7804
rect 3908 7800 3912 7804
rect 3923 7800 3927 7804
rect 3951 7800 3955 7804
rect 3202 7786 3206 7790
rect 3221 7786 3225 7790
rect 3234 7787 3238 7791
rect 3256 7786 3260 7790
rect 3264 7787 3268 7791
rect 3276 7787 3280 7791
rect 3325 7786 3329 7790
rect 3341 7786 3345 7792
rect 3375 7792 3379 7796
rect 3362 7786 3366 7790
rect 3383 7786 3387 7790
rect 3399 7786 3403 7792
rect 3420 7786 3424 7790
rect 3436 7786 3440 7790
rect 3457 7786 3461 7790
rect 3473 7786 3477 7792
rect 3507 7792 3511 7796
rect 3494 7786 3498 7790
rect 3515 7786 3519 7790
rect 3531 7786 3535 7792
rect 3552 7786 3556 7790
rect 3568 7786 3572 7790
rect 3589 7786 3593 7790
rect 3605 7786 3609 7792
rect 3639 7792 3643 7796
rect 3626 7786 3630 7790
rect 3647 7786 3651 7790
rect 3663 7786 3667 7792
rect 3684 7786 3688 7790
rect 3700 7786 3704 7790
rect 3796 7788 3800 7792
rect 3090 7770 3094 7774
rect 3116 7770 3120 7774
rect 664 7761 668 7765
rect 674 7761 678 7765
rect 684 7761 688 7765
rect 2373 7759 2377 7763
rect 2424 7759 2428 7763
rect 2474 7759 2478 7763
rect 2505 7759 2509 7763
rect 2556 7759 2560 7763
rect 2606 7759 2610 7763
rect 2637 7759 2641 7763
rect 2688 7759 2692 7763
rect 2738 7759 2742 7763
rect 2812 7760 2818 7764
rect 2864 7760 2868 7764
rect 2882 7760 2886 7764
rect 2913 7760 2917 7764
rect 2935 7760 2939 7764
rect 3000 7760 3004 7764
rect 3142 7767 3146 7771
rect 3149 7770 3153 7774
rect 3167 7770 3171 7774
rect 3189 7767 3193 7771
rect 3214 7767 3218 7771
rect 3224 7770 3228 7774
rect 3240 7770 3244 7774
rect 3260 7767 3264 7771
rect 3267 7770 3271 7774
rect 3318 7775 3322 7779
rect 3355 7773 3359 7777
rect 3375 7773 3379 7777
rect 3419 7773 3423 7777
rect 3450 7775 3454 7779
rect 3487 7773 3491 7777
rect 3507 7773 3511 7777
rect 3551 7773 3555 7777
rect 3582 7775 3586 7779
rect 3619 7773 3623 7777
rect 3639 7773 3643 7777
rect 3683 7773 3687 7777
rect 3828 7786 3832 7790
rect 3848 7789 3852 7793
rect 3867 7785 3871 7789
rect 3886 7786 3890 7790
rect 3905 7786 3909 7790
rect 3918 7787 3922 7791
rect 4054 7812 4058 7816
rect 4076 7812 4080 7816
rect 4135 7812 4139 7816
rect 4160 7812 4164 7816
rect 4191 7812 4195 7816
rect 4076 7804 4080 7808
rect 4119 7805 4123 7809
rect 4141 7804 4148 7808
rect 4191 7805 4195 7809
rect 4094 7800 4098 7804
rect 4112 7800 4116 7804
rect 4169 7800 4173 7804
rect 4184 7800 4188 7804
rect 4212 7800 4216 7804
rect 4015 7796 4019 7800
rect 3940 7786 3944 7790
rect 3948 7787 3952 7791
rect 3960 7787 3964 7791
rect 3994 7781 3998 7785
rect 4034 7787 4038 7791
rect 4023 7780 4027 7784
rect 3801 7770 3805 7774
rect 3721 7766 3727 7770
rect 3826 7767 3830 7771
rect 3833 7770 3837 7774
rect 3851 7770 3855 7774
rect 3873 7767 3877 7771
rect 3898 7767 3902 7771
rect 3908 7770 3912 7774
rect 3924 7770 3928 7774
rect 3944 7767 3948 7771
rect 3951 7770 3955 7774
rect 4089 7786 4093 7790
rect 4109 7789 4113 7793
rect 4128 7785 4132 7789
rect 4147 7786 4151 7790
rect 4166 7786 4170 7790
rect 4179 7787 4183 7791
rect 4201 7786 4205 7790
rect 4209 7787 4213 7791
rect 4221 7787 4225 7791
rect 4484 7789 4488 7793
rect 4494 7789 4498 7793
rect 4504 7789 4508 7793
rect 4484 7784 4488 7788
rect 4494 7784 4498 7788
rect 4504 7784 4508 7788
rect 4484 7779 4488 7783
rect 4494 7779 4498 7783
rect 4504 7779 4508 7783
rect 4484 7774 4488 7778
rect 4494 7774 4498 7778
rect 4504 7774 4508 7778
rect 4530 7789 4534 7793
rect 4540 7789 4544 7793
rect 4550 7789 4554 7793
rect 4530 7784 4534 7788
rect 4540 7784 4544 7788
rect 4550 7784 4554 7788
rect 4530 7779 4534 7783
rect 4540 7779 4544 7783
rect 4550 7779 4554 7783
rect 4530 7774 4534 7778
rect 4540 7774 4544 7778
rect 4550 7774 4554 7778
rect 4035 7770 4039 7774
rect 4061 7770 4065 7774
rect 3060 7760 3064 7764
rect 3099 7760 3103 7764
rect 3143 7760 3147 7764
rect 3174 7760 3178 7764
rect 3196 7760 3200 7764
rect 3261 7760 3265 7764
rect 3318 7759 3322 7763
rect 3369 7759 3373 7763
rect 3419 7759 3423 7763
rect 3450 7759 3454 7763
rect 3501 7759 3505 7763
rect 3551 7759 3555 7763
rect 3582 7759 3586 7763
rect 3633 7759 3637 7763
rect 3683 7759 3687 7763
rect 3757 7760 3763 7764
rect 3809 7760 3813 7764
rect 3827 7760 3831 7764
rect 3858 7760 3862 7764
rect 3880 7760 3884 7764
rect 3945 7760 3949 7764
rect 4087 7767 4091 7771
rect 4094 7770 4098 7774
rect 4112 7770 4116 7774
rect 4134 7767 4138 7771
rect 4159 7767 4163 7771
rect 4169 7770 4173 7774
rect 4185 7770 4189 7774
rect 4205 7767 4209 7771
rect 4212 7770 4216 7774
rect 4005 7760 4009 7764
rect 4044 7760 4048 7764
rect 4088 7760 4092 7764
rect 4119 7760 4123 7764
rect 4141 7760 4145 7764
rect 4206 7760 4210 7764
rect 2367 7752 2371 7756
rect 2755 7752 2759 7756
rect 2764 7753 2770 7757
rect 2855 7753 2859 7757
rect 2889 7753 2893 7757
rect 2906 7753 2910 7757
rect 2962 7753 2966 7757
rect 2979 7753 2983 7757
rect 3007 7753 3011 7757
rect 3090 7753 3094 7757
rect 3116 7753 3120 7757
rect 3150 7753 3154 7757
rect 3167 7753 3171 7757
rect 3223 7753 3227 7757
rect 3240 7753 3244 7757
rect 3268 7753 3272 7757
rect 3312 7752 3316 7756
rect 3700 7752 3704 7756
rect 3709 7753 3715 7757
rect 3800 7753 3804 7757
rect 3834 7753 3838 7757
rect 3851 7753 3855 7757
rect 3907 7753 3911 7757
rect 3924 7753 3928 7757
rect 3952 7753 3956 7757
rect 4035 7753 4039 7757
rect 4061 7753 4065 7757
rect 4095 7753 4099 7757
rect 4112 7753 4116 7757
rect 4168 7753 4172 7757
rect 4185 7753 4189 7757
rect 4213 7753 4217 7757
rect 2490 7745 2495 7749
rect 2623 7745 2627 7749
rect 2800 7746 2806 7750
rect 2864 7746 2868 7750
rect 3098 7746 3102 7750
rect 3284 7747 3288 7751
rect 3296 7747 3300 7751
rect 3435 7745 3440 7749
rect 3568 7745 3572 7749
rect 3745 7746 3751 7750
rect 3809 7746 3813 7750
rect 4043 7746 4047 7750
rect 4229 7747 4233 7751
rect 4241 7747 4245 7751
rect 2498 7738 2502 7742
rect 2788 7738 2794 7742
rect 3108 7739 3112 7743
rect 3273 7739 3277 7743
rect 2482 7734 2486 7738
rect 2514 7734 2518 7738
rect 2836 7732 2842 7736
rect 3443 7738 3447 7742
rect 3733 7738 3739 7742
rect 4053 7739 4057 7743
rect 4218 7739 4222 7743
rect 3427 7734 3431 7738
rect 3459 7734 3463 7738
rect 3781 7732 3787 7736
rect 2482 7725 2486 7729
rect 2514 7725 2518 7729
rect 3427 7725 3431 7729
rect 3459 7725 3463 7729
rect 2498 7718 2502 7722
rect 2755 7718 2759 7722
rect 2824 7718 2830 7722
rect 3156 7718 3160 7722
rect 3192 7718 3196 7722
rect 3259 7718 3263 7722
rect 3443 7718 3447 7722
rect 3700 7718 3704 7722
rect 3769 7718 3775 7722
rect 4101 7718 4105 7722
rect 4137 7718 4141 7722
rect 4204 7718 4208 7722
rect 2755 7710 2759 7714
rect 2764 7711 2770 7715
rect 3142 7711 3146 7715
rect 2482 7706 2486 7710
rect 2514 7706 2518 7710
rect 2498 7702 2502 7706
rect 3156 7704 3160 7708
rect 3206 7704 3210 7708
rect 3259 7704 3263 7708
rect 3700 7710 3704 7714
rect 3709 7711 3715 7715
rect 4087 7711 4091 7715
rect 3427 7706 3431 7710
rect 3459 7706 3463 7710
rect 3443 7702 3447 7706
rect 4101 7704 4105 7708
rect 4151 7704 4155 7708
rect 4204 7704 4208 7708
rect 2490 7695 2495 7699
rect 2624 7695 2628 7699
rect 3179 7693 3183 7697
rect 2373 7688 2377 7692
rect 2409 7688 2413 7692
rect 2476 7688 2480 7692
rect 2505 7688 2509 7692
rect 2541 7688 2545 7692
rect 2608 7688 2612 7692
rect 2637 7688 2641 7692
rect 2673 7688 2677 7692
rect 2740 7688 2744 7692
rect 2824 7688 2830 7692
rect 2764 7681 2770 7685
rect 3150 7684 3154 7688
rect 3163 7687 3167 7693
rect 3200 7687 3204 7693
rect 3213 7689 3217 7693
rect 3237 7693 3241 7697
rect 3435 7695 3440 7699
rect 3569 7695 3573 7699
rect 4124 7693 4128 7697
rect 3221 7687 3225 7693
rect 3258 7687 3262 7693
rect 3274 7687 3278 7693
rect 3318 7688 3322 7692
rect 3354 7688 3358 7692
rect 3421 7688 3425 7692
rect 3450 7688 3454 7692
rect 3486 7688 3490 7692
rect 3553 7688 3557 7692
rect 3582 7688 3586 7692
rect 3618 7688 3622 7692
rect 3685 7688 3689 7692
rect 3769 7688 3775 7692
rect 2373 7674 2377 7678
rect 2423 7674 2427 7678
rect 2476 7674 2480 7678
rect 2505 7674 2509 7678
rect 2555 7674 2559 7678
rect 2608 7674 2612 7678
rect 2637 7674 2641 7678
rect 2687 7674 2691 7678
rect 2740 7674 2744 7678
rect 3163 7674 3167 7678
rect 3179 7674 3183 7680
rect 3213 7680 3217 7684
rect 3200 7674 3204 7678
rect 2396 7663 2400 7667
rect 2367 7654 2371 7658
rect 2380 7657 2384 7663
rect 2417 7657 2421 7663
rect 2430 7659 2434 7663
rect 2454 7663 2458 7667
rect 2528 7663 2532 7667
rect 2438 7657 2442 7663
rect 2475 7657 2479 7663
rect 2491 7657 2495 7663
rect 2512 7657 2516 7663
rect 2549 7657 2553 7663
rect 2562 7659 2566 7663
rect 2586 7663 2590 7667
rect 2660 7663 2664 7667
rect 2570 7657 2574 7663
rect 2607 7657 2611 7663
rect 2623 7657 2627 7663
rect 2644 7657 2648 7663
rect 2681 7657 2685 7663
rect 2694 7659 2698 7663
rect 2718 7663 2722 7667
rect 2702 7657 2706 7663
rect 2739 7657 2743 7663
rect 2755 7659 2759 7663
rect 3221 7674 3225 7678
rect 3237 7674 3241 7680
rect 3709 7681 3715 7685
rect 4095 7684 4099 7688
rect 4108 7687 4112 7693
rect 4145 7687 4149 7693
rect 4158 7689 4162 7693
rect 4182 7693 4186 7697
rect 4166 7687 4170 7693
rect 4203 7687 4207 7693
rect 4219 7687 4223 7693
rect 3258 7674 3262 7678
rect 3274 7674 3278 7678
rect 3318 7674 3322 7678
rect 3368 7674 3372 7678
rect 3421 7674 3425 7678
rect 3450 7674 3454 7678
rect 3500 7674 3504 7678
rect 3553 7674 3557 7678
rect 3582 7674 3586 7678
rect 3632 7674 3636 7678
rect 3685 7674 3689 7678
rect 4108 7674 4112 7678
rect 4124 7674 4128 7680
rect 4158 7680 4162 7684
rect 4145 7674 4149 7678
rect 3156 7663 3160 7667
rect 3193 7661 3197 7665
rect 3213 7661 3217 7665
rect 3257 7661 3261 7665
rect 3341 7663 3345 7667
rect 2380 7644 2384 7648
rect 2396 7644 2400 7650
rect 2430 7650 2434 7654
rect 2417 7644 2421 7648
rect 2438 7644 2442 7648
rect 2454 7644 2458 7650
rect 2475 7644 2479 7648
rect 2491 7644 2495 7648
rect 2512 7644 2516 7648
rect 2528 7644 2532 7650
rect 2562 7650 2566 7654
rect 2549 7644 2553 7648
rect 2570 7644 2574 7648
rect 2586 7644 2590 7650
rect 2607 7644 2611 7648
rect 2623 7644 2627 7648
rect 2644 7644 2648 7648
rect 2660 7644 2664 7650
rect 2694 7650 2698 7654
rect 2681 7644 2685 7648
rect 2702 7644 2706 7648
rect 2718 7644 2722 7650
rect 2776 7654 2782 7658
rect 3312 7654 3316 7658
rect 3325 7657 3329 7663
rect 3362 7657 3366 7663
rect 3375 7659 3379 7663
rect 3399 7663 3403 7667
rect 3473 7663 3477 7667
rect 3383 7657 3387 7663
rect 3420 7657 3424 7663
rect 3436 7657 3440 7663
rect 3457 7657 3461 7663
rect 3494 7657 3498 7663
rect 3507 7659 3511 7663
rect 3531 7663 3535 7667
rect 3605 7663 3609 7667
rect 3515 7657 3519 7663
rect 3552 7657 3556 7663
rect 3568 7657 3572 7663
rect 3589 7657 3593 7663
rect 3626 7657 3630 7663
rect 3639 7659 3643 7663
rect 3663 7663 3667 7667
rect 3647 7657 3651 7663
rect 3684 7657 3688 7663
rect 3700 7659 3704 7663
rect 4166 7674 4170 7678
rect 4182 7674 4186 7680
rect 4203 7674 4207 7678
rect 4219 7674 4223 7678
rect 4101 7663 4105 7667
rect 4138 7661 4142 7665
rect 4158 7661 4162 7665
rect 4202 7661 4206 7665
rect 2739 7644 2743 7648
rect 2755 7644 2759 7648
rect 2812 7647 2818 7651
rect 3156 7647 3160 7651
rect 3207 7647 3211 7651
rect 3257 7647 3261 7651
rect 3325 7644 3329 7648
rect 3341 7644 3345 7650
rect 3375 7650 3379 7654
rect 3362 7644 3366 7648
rect 2373 7633 2377 7637
rect 2410 7631 2414 7635
rect 2430 7631 2434 7635
rect 2474 7631 2478 7635
rect 2505 7633 2509 7637
rect 2542 7631 2546 7635
rect 2562 7631 2566 7635
rect 2606 7631 2610 7635
rect 2637 7633 2641 7637
rect 2674 7631 2678 7635
rect 2694 7631 2698 7635
rect 2738 7631 2742 7635
rect 3149 7639 3153 7643
rect 3274 7640 3278 7644
rect 3383 7644 3387 7648
rect 3399 7644 3403 7650
rect 3420 7644 3424 7648
rect 3436 7644 3440 7648
rect 3457 7644 3461 7648
rect 3473 7644 3477 7650
rect 3507 7650 3511 7654
rect 3494 7644 3498 7648
rect 3515 7644 3519 7648
rect 3531 7644 3535 7650
rect 3552 7644 3556 7648
rect 3568 7644 3572 7648
rect 3589 7644 3593 7648
rect 3605 7644 3609 7650
rect 3639 7650 3643 7654
rect 3626 7644 3630 7648
rect 3647 7644 3651 7648
rect 3663 7644 3667 7650
rect 3721 7654 3727 7658
rect 3684 7644 3688 7648
rect 3700 7644 3704 7648
rect 3757 7647 3763 7651
rect 4101 7647 4105 7651
rect 4152 7647 4156 7651
rect 4202 7647 4206 7651
rect 2824 7632 2830 7636
rect 3156 7632 3160 7636
rect 3192 7632 3196 7636
rect 3259 7632 3263 7636
rect 2776 7624 2782 7628
rect 3142 7625 3146 7629
rect 3318 7633 3322 7637
rect 3355 7631 3359 7635
rect 3375 7631 3379 7635
rect 3419 7631 3423 7635
rect 3450 7633 3454 7637
rect 3487 7631 3491 7635
rect 3507 7631 3511 7635
rect 3551 7631 3555 7635
rect 3582 7633 3586 7637
rect 3619 7631 3623 7635
rect 3639 7631 3643 7635
rect 3683 7631 3687 7635
rect 4094 7639 4098 7643
rect 4219 7640 4223 7644
rect 3769 7632 3775 7636
rect 4101 7632 4105 7636
rect 4137 7632 4141 7636
rect 4204 7632 4208 7636
rect 2373 7617 2377 7621
rect 2424 7617 2428 7621
rect 2474 7617 2478 7621
rect 2505 7617 2509 7621
rect 2556 7617 2560 7621
rect 2606 7617 2610 7621
rect 2637 7617 2641 7621
rect 2688 7617 2692 7621
rect 2738 7617 2742 7621
rect 2812 7617 2818 7621
rect 3156 7618 3160 7622
rect 3206 7618 3210 7622
rect 3259 7618 3263 7622
rect 3721 7624 3727 7628
rect 4087 7625 4091 7629
rect 3318 7617 3322 7621
rect 3369 7617 3373 7621
rect 3419 7617 3423 7621
rect 3450 7617 3454 7621
rect 3501 7617 3505 7621
rect 3551 7617 3555 7621
rect 3582 7617 3586 7621
rect 3633 7617 3637 7621
rect 3683 7617 3687 7621
rect 3757 7617 3763 7621
rect 4101 7618 4105 7622
rect 4151 7618 4155 7622
rect 4204 7618 4208 7622
rect 2366 7610 2370 7614
rect 2755 7610 2759 7614
rect 3179 7607 3183 7611
rect 2373 7602 2377 7606
rect 2409 7602 2413 7606
rect 2476 7602 2480 7606
rect 2505 7602 2509 7606
rect 2541 7602 2545 7606
rect 2608 7602 2612 7606
rect 2637 7602 2641 7606
rect 2673 7602 2677 7606
rect 2740 7602 2744 7606
rect 2824 7602 2830 7606
rect 2764 7595 2770 7599
rect 3150 7598 3154 7602
rect 3163 7601 3167 7607
rect 3200 7601 3204 7607
rect 3213 7603 3217 7607
rect 3237 7607 3241 7611
rect 3311 7610 3315 7614
rect 3700 7610 3704 7614
rect 4124 7607 4128 7611
rect 3221 7601 3225 7607
rect 3258 7601 3262 7607
rect 3274 7603 3278 7607
rect 3296 7601 3300 7605
rect 3318 7602 3322 7606
rect 3354 7602 3358 7606
rect 3421 7602 3425 7606
rect 3450 7602 3454 7606
rect 3486 7602 3490 7606
rect 3553 7602 3557 7606
rect 3582 7602 3586 7606
rect 3618 7602 3622 7606
rect 3685 7602 3689 7606
rect 3769 7602 3775 7606
rect 2373 7588 2377 7592
rect 2423 7588 2427 7592
rect 2476 7588 2480 7592
rect 2505 7588 2509 7592
rect 2555 7588 2559 7592
rect 2608 7588 2612 7592
rect 2637 7588 2641 7592
rect 2687 7588 2691 7592
rect 2740 7588 2744 7592
rect 3163 7588 3167 7592
rect 3179 7588 3183 7594
rect 3213 7594 3217 7598
rect 3200 7588 3204 7592
rect 2396 7577 2400 7581
rect 2367 7568 2371 7572
rect 2380 7571 2384 7577
rect 2417 7571 2421 7577
rect 2430 7573 2434 7577
rect 2454 7577 2458 7581
rect 2528 7577 2532 7581
rect 2438 7571 2442 7577
rect 2475 7571 2479 7577
rect 2491 7571 2495 7577
rect 2512 7571 2516 7577
rect 2549 7571 2553 7577
rect 2562 7573 2566 7577
rect 2586 7577 2590 7581
rect 2660 7577 2664 7581
rect 2570 7571 2574 7577
rect 2607 7571 2611 7577
rect 2623 7571 2627 7577
rect 2644 7571 2648 7577
rect 2681 7571 2685 7577
rect 2694 7573 2698 7577
rect 2718 7577 2722 7581
rect 2702 7571 2706 7577
rect 2739 7571 2743 7577
rect 2755 7573 2759 7577
rect 3221 7588 3225 7592
rect 3237 7588 3241 7594
rect 3258 7588 3262 7592
rect 3274 7588 3278 7597
rect 3709 7595 3715 7599
rect 4095 7598 4099 7602
rect 4108 7601 4112 7607
rect 4145 7601 4149 7607
rect 4158 7603 4162 7607
rect 4182 7607 4186 7611
rect 4166 7601 4170 7607
rect 4203 7601 4207 7607
rect 4219 7603 4223 7607
rect 4241 7601 4245 7605
rect 3296 7585 3300 7589
rect 3318 7588 3322 7592
rect 3368 7588 3372 7592
rect 3421 7588 3425 7592
rect 3450 7588 3454 7592
rect 3500 7588 3504 7592
rect 3553 7588 3557 7592
rect 3582 7588 3586 7592
rect 3632 7588 3636 7592
rect 3685 7588 3689 7592
rect 4108 7588 4112 7592
rect 4124 7588 4128 7594
rect 4158 7594 4162 7598
rect 4145 7588 4149 7592
rect 3156 7577 3160 7581
rect 3193 7575 3197 7579
rect 3213 7575 3217 7579
rect 3257 7575 3261 7579
rect 3341 7577 3345 7581
rect 2380 7558 2384 7562
rect 2396 7558 2400 7564
rect 2430 7564 2434 7568
rect 2417 7558 2421 7562
rect 2438 7558 2442 7562
rect 2454 7558 2458 7564
rect 2475 7558 2479 7562
rect 2491 7558 2495 7562
rect 2512 7558 2516 7562
rect 2528 7558 2532 7564
rect 2562 7564 2566 7568
rect 2549 7558 2553 7562
rect 2570 7558 2574 7562
rect 2586 7558 2590 7564
rect 2607 7558 2611 7562
rect 2623 7558 2627 7562
rect 2644 7558 2648 7562
rect 2660 7558 2664 7564
rect 2694 7564 2698 7568
rect 2681 7558 2685 7562
rect 2702 7558 2706 7562
rect 2718 7558 2722 7564
rect 2776 7568 2782 7572
rect 3312 7568 3316 7572
rect 3325 7571 3329 7577
rect 3362 7571 3366 7577
rect 3375 7573 3379 7577
rect 3399 7577 3403 7581
rect 3473 7577 3477 7581
rect 3383 7571 3387 7577
rect 3420 7571 3424 7577
rect 3436 7571 3440 7577
rect 3457 7571 3461 7577
rect 3494 7571 3498 7577
rect 3507 7573 3511 7577
rect 3531 7577 3535 7581
rect 3605 7577 3609 7581
rect 3515 7571 3519 7577
rect 3552 7571 3556 7577
rect 3568 7571 3572 7577
rect 3589 7571 3593 7577
rect 3626 7571 3630 7577
rect 3639 7573 3643 7577
rect 3663 7577 3667 7581
rect 3647 7571 3651 7577
rect 3684 7571 3688 7577
rect 3700 7573 3704 7577
rect 4166 7588 4170 7592
rect 4182 7588 4186 7594
rect 4203 7588 4207 7592
rect 4219 7588 4223 7597
rect 4241 7585 4245 7589
rect 4101 7577 4105 7581
rect 4138 7575 4142 7579
rect 4158 7575 4162 7579
rect 4202 7575 4206 7579
rect 2739 7558 2743 7562
rect 2755 7558 2759 7562
rect 2812 7561 2818 7565
rect 3156 7561 3160 7565
rect 3207 7561 3211 7565
rect 3257 7561 3261 7565
rect 3325 7558 3329 7562
rect 3341 7558 3345 7564
rect 3375 7564 3379 7568
rect 3362 7558 3366 7562
rect 3383 7558 3387 7562
rect 3399 7558 3403 7564
rect 3420 7558 3424 7562
rect 3436 7558 3440 7562
rect 3457 7558 3461 7562
rect 3473 7558 3477 7564
rect 3507 7564 3511 7568
rect 3494 7558 3498 7562
rect 3515 7558 3519 7562
rect 3531 7558 3535 7564
rect 3552 7558 3556 7562
rect 3568 7558 3572 7562
rect 3589 7558 3593 7562
rect 3605 7558 3609 7564
rect 3639 7564 3643 7568
rect 3626 7558 3630 7562
rect 3647 7558 3651 7562
rect 3663 7558 3667 7564
rect 3721 7568 3727 7572
rect 3684 7558 3688 7562
rect 3700 7558 3704 7562
rect 3757 7561 3763 7565
rect 4101 7561 4105 7565
rect 4152 7561 4156 7565
rect 4202 7561 4206 7565
rect 2373 7547 2377 7551
rect 2410 7545 2414 7549
rect 2430 7545 2434 7549
rect 2474 7545 2478 7549
rect 2505 7547 2509 7551
rect 2542 7545 2546 7549
rect 2562 7545 2566 7549
rect 2606 7545 2610 7549
rect 2637 7547 2641 7551
rect 2674 7545 2678 7549
rect 2694 7545 2698 7549
rect 2738 7545 2742 7549
rect 3318 7547 3322 7551
rect 3355 7545 3359 7549
rect 3375 7545 3379 7549
rect 3419 7545 3423 7549
rect 3450 7547 3454 7551
rect 3487 7545 3491 7549
rect 3507 7545 3511 7549
rect 3551 7545 3555 7549
rect 3582 7547 3586 7551
rect 3619 7545 3623 7549
rect 3639 7545 3643 7549
rect 3683 7545 3687 7549
rect 2776 7538 2782 7542
rect 3721 7538 3727 7542
rect 2373 7531 2377 7535
rect 2424 7531 2428 7535
rect 2474 7531 2478 7535
rect 2505 7531 2509 7535
rect 2556 7531 2560 7535
rect 2606 7531 2610 7535
rect 2637 7531 2641 7535
rect 2688 7531 2692 7535
rect 2738 7531 2742 7535
rect 2812 7531 2818 7535
rect 3318 7531 3322 7535
rect 3369 7531 3373 7535
rect 3419 7531 3423 7535
rect 3450 7531 3454 7535
rect 3501 7531 3505 7535
rect 3551 7531 3555 7535
rect 3582 7531 3586 7535
rect 3633 7531 3637 7535
rect 3683 7531 3687 7535
rect 3757 7531 3763 7535
rect 2366 7524 2370 7528
rect 2755 7524 2759 7528
rect 3311 7524 3315 7528
rect 3700 7524 3704 7528
rect 2491 7517 2495 7521
rect 2599 7517 2603 7521
rect 2623 7517 2627 7521
rect 3436 7517 3440 7521
rect 3544 7517 3548 7521
rect 3568 7517 3572 7521
rect 2615 7510 2619 7514
rect 2599 7506 2603 7510
rect 2631 7506 2635 7510
rect 3560 7510 3564 7514
rect 3544 7506 3548 7510
rect 3576 7506 3580 7510
rect 2599 7499 2603 7503
rect 2631 7499 2635 7503
rect 3296 7499 3300 7503
rect 3544 7499 3548 7503
rect 3576 7499 3580 7503
rect 4241 7499 4245 7503
rect 2615 7492 2619 7496
rect 2755 7492 2759 7496
rect 3560 7492 3564 7496
rect 3700 7492 3704 7496
rect 2755 7484 2759 7488
rect 3700 7484 3704 7488
rect 2599 7480 2603 7484
rect 2631 7480 2635 7484
rect 2615 7476 2619 7480
rect 3544 7480 3548 7484
rect 3576 7480 3580 7484
rect 3560 7476 3564 7480
rect 618 7467 622 7471
rect 628 7467 632 7471
rect 638 7467 642 7471
rect 618 7462 622 7466
rect 628 7462 632 7466
rect 638 7462 642 7466
rect 618 7457 622 7461
rect 628 7457 632 7461
rect 638 7457 642 7461
rect 618 7452 622 7456
rect 628 7452 632 7456
rect 638 7452 642 7456
rect 664 7467 668 7471
rect 674 7467 678 7471
rect 684 7467 688 7471
rect 2491 7469 2495 7473
rect 2599 7469 2603 7473
rect 2623 7469 2627 7473
rect 3436 7469 3440 7473
rect 3544 7469 3548 7473
rect 3568 7469 3572 7473
rect 664 7462 668 7466
rect 674 7462 678 7466
rect 684 7462 688 7466
rect 2373 7462 2377 7466
rect 2409 7462 2413 7466
rect 2476 7462 2480 7466
rect 2505 7462 2509 7466
rect 2541 7462 2545 7466
rect 2608 7462 2612 7466
rect 2637 7462 2641 7466
rect 2673 7462 2677 7466
rect 2740 7462 2744 7466
rect 2824 7462 2830 7466
rect 3318 7462 3322 7466
rect 3354 7462 3358 7466
rect 3421 7462 3425 7466
rect 3450 7462 3454 7466
rect 3486 7462 3490 7466
rect 3553 7462 3557 7466
rect 3582 7462 3586 7466
rect 3618 7462 3622 7466
rect 3685 7462 3689 7466
rect 3769 7462 3775 7466
rect 664 7457 668 7461
rect 674 7457 678 7461
rect 684 7457 688 7461
rect 664 7452 668 7456
rect 674 7452 678 7456
rect 684 7452 688 7456
rect 2764 7455 2770 7459
rect 3709 7455 3715 7459
rect 2373 7448 2377 7452
rect 2423 7448 2427 7452
rect 2476 7448 2480 7452
rect 2505 7448 2509 7452
rect 2555 7448 2559 7452
rect 2608 7448 2612 7452
rect 2637 7448 2641 7452
rect 2687 7448 2691 7452
rect 2740 7448 2744 7452
rect 3318 7448 3322 7452
rect 3368 7448 3372 7452
rect 3421 7448 3425 7452
rect 3450 7448 3454 7452
rect 3500 7448 3504 7452
rect 3553 7448 3557 7452
rect 3582 7448 3586 7452
rect 3632 7448 3636 7452
rect 3685 7448 3689 7452
rect 2396 7437 2400 7441
rect 2367 7428 2371 7432
rect 2380 7431 2384 7437
rect 2417 7431 2421 7437
rect 2430 7433 2434 7437
rect 2454 7437 2458 7441
rect 2528 7437 2532 7441
rect 2438 7431 2442 7437
rect 2475 7431 2479 7437
rect 2491 7431 2495 7437
rect 2512 7431 2516 7437
rect 2549 7431 2553 7437
rect 2562 7433 2566 7437
rect 2586 7437 2590 7441
rect 2660 7437 2664 7441
rect 2570 7431 2574 7437
rect 2607 7431 2611 7437
rect 2623 7431 2627 7437
rect 2644 7431 2648 7437
rect 2681 7431 2685 7437
rect 2694 7433 2698 7437
rect 2718 7437 2722 7441
rect 3341 7437 3345 7441
rect 2702 7431 2706 7437
rect 2739 7431 2743 7437
rect 2755 7433 2759 7437
rect 2380 7418 2384 7422
rect 2396 7418 2400 7424
rect 2430 7424 2434 7428
rect 2417 7418 2421 7422
rect 2438 7418 2442 7422
rect 2454 7418 2458 7424
rect 2475 7418 2479 7422
rect 2491 7418 2495 7422
rect 2512 7418 2516 7422
rect 2528 7418 2532 7424
rect 2562 7424 2566 7428
rect 2549 7418 2553 7422
rect 2570 7418 2574 7422
rect 2586 7418 2590 7424
rect 2607 7418 2611 7422
rect 2623 7418 2627 7422
rect 2644 7418 2648 7422
rect 2660 7418 2664 7424
rect 2694 7424 2698 7428
rect 2681 7418 2685 7422
rect 2702 7418 2706 7422
rect 2718 7418 2722 7424
rect 3312 7428 3316 7432
rect 3325 7431 3329 7437
rect 3362 7431 3366 7437
rect 3375 7433 3379 7437
rect 3399 7437 3403 7441
rect 3473 7437 3477 7441
rect 3383 7431 3387 7437
rect 3420 7431 3424 7437
rect 3436 7431 3440 7437
rect 3457 7431 3461 7437
rect 3494 7431 3498 7437
rect 3507 7433 3511 7437
rect 3531 7437 3535 7441
rect 3605 7437 3609 7441
rect 3515 7431 3519 7437
rect 3552 7431 3556 7437
rect 3568 7431 3572 7437
rect 3589 7431 3593 7437
rect 3626 7431 3630 7437
rect 3639 7433 3643 7437
rect 3663 7437 3667 7441
rect 3647 7431 3651 7437
rect 3684 7431 3688 7437
rect 3700 7433 3704 7437
rect 2739 7418 2743 7422
rect 2755 7418 2759 7422
rect 3325 7418 3329 7422
rect 3341 7418 3345 7424
rect 3375 7424 3379 7428
rect 3362 7418 3366 7422
rect 3383 7418 3387 7422
rect 3399 7418 3403 7424
rect 3420 7418 3424 7422
rect 3436 7418 3440 7422
rect 3457 7418 3461 7422
rect 3473 7418 3477 7424
rect 3507 7424 3511 7428
rect 3494 7418 3498 7422
rect 3515 7418 3519 7422
rect 3531 7418 3535 7424
rect 3552 7418 3556 7422
rect 3568 7418 3572 7422
rect 3589 7418 3593 7422
rect 3605 7418 3609 7424
rect 3639 7424 3643 7428
rect 3626 7418 3630 7422
rect 3647 7418 3651 7422
rect 3663 7418 3667 7424
rect 3684 7418 3688 7422
rect 3700 7418 3704 7422
rect 2373 7407 2377 7411
rect 2410 7405 2414 7409
rect 2430 7405 2434 7409
rect 2474 7405 2478 7409
rect 2505 7407 2509 7411
rect 2542 7405 2546 7409
rect 2562 7405 2566 7409
rect 2606 7405 2610 7409
rect 2637 7407 2641 7411
rect 2674 7405 2678 7409
rect 2694 7405 2698 7409
rect 2738 7405 2742 7409
rect 3318 7407 3322 7411
rect 3355 7405 3359 7409
rect 3375 7405 3379 7409
rect 3419 7405 3423 7409
rect 3450 7407 3454 7411
rect 3487 7405 3491 7409
rect 3507 7405 3511 7409
rect 3551 7405 3555 7409
rect 3582 7407 3586 7411
rect 3619 7405 3623 7409
rect 3639 7405 3643 7409
rect 3683 7405 3687 7409
rect 2776 7398 2782 7402
rect 3721 7398 3727 7402
rect 2373 7391 2377 7395
rect 2424 7391 2428 7395
rect 2474 7391 2478 7395
rect 2505 7391 2509 7395
rect 2556 7391 2560 7395
rect 2606 7391 2610 7395
rect 2637 7391 2641 7395
rect 2688 7391 2692 7395
rect 2738 7391 2742 7395
rect 2812 7391 2818 7395
rect 3318 7391 3322 7395
rect 3369 7391 3373 7395
rect 3419 7391 3423 7395
rect 3450 7391 3454 7395
rect 3501 7391 3505 7395
rect 3551 7391 3555 7395
rect 3582 7391 3586 7395
rect 3633 7391 3637 7395
rect 3683 7391 3687 7395
rect 3757 7391 3763 7395
rect 4484 7202 4488 7206
rect 4494 7202 4498 7206
rect 4504 7202 4508 7206
rect 4484 7197 4488 7201
rect 4494 7197 4498 7201
rect 4504 7197 4508 7201
rect 4484 7192 4488 7196
rect 4494 7192 4498 7196
rect 4504 7192 4508 7196
rect 4484 7187 4488 7191
rect 4494 7187 4498 7191
rect 4504 7187 4508 7191
rect 4530 7202 4534 7206
rect 4540 7202 4544 7206
rect 4550 7202 4554 7206
rect 4530 7197 4534 7201
rect 4540 7197 4544 7201
rect 4550 7197 4554 7201
rect 4530 7192 4534 7196
rect 4540 7192 4544 7196
rect 4550 7192 4554 7196
rect 4530 7187 4534 7191
rect 4540 7187 4544 7191
rect 4550 7187 4554 7191
rect 618 7158 622 7162
rect 628 7158 632 7162
rect 638 7158 642 7162
rect 618 7153 622 7157
rect 628 7153 632 7157
rect 638 7153 642 7157
rect 618 7148 622 7152
rect 628 7148 632 7152
rect 638 7148 642 7152
rect 618 7143 622 7147
rect 628 7143 632 7147
rect 638 7143 642 7147
rect 664 7158 668 7162
rect 674 7158 678 7162
rect 684 7158 688 7162
rect 664 7153 668 7157
rect 674 7153 678 7157
rect 684 7153 688 7157
rect 664 7148 668 7152
rect 674 7148 678 7152
rect 684 7148 688 7152
rect 664 7143 668 7147
rect 674 7143 678 7147
rect 684 7143 688 7147
rect 4484 6893 4488 6897
rect 4494 6893 4498 6897
rect 4504 6893 4508 6897
rect 4484 6888 4488 6892
rect 4494 6888 4498 6892
rect 4504 6888 4508 6892
rect 4484 6883 4488 6887
rect 4494 6883 4498 6887
rect 4504 6883 4508 6887
rect 4484 6878 4488 6882
rect 4494 6878 4498 6882
rect 4504 6878 4508 6882
rect 4530 6893 4534 6897
rect 4540 6893 4544 6897
rect 4550 6893 4554 6897
rect 4530 6888 4534 6892
rect 4540 6888 4544 6892
rect 4550 6888 4554 6892
rect 4530 6883 4534 6887
rect 4540 6883 4544 6887
rect 4550 6883 4554 6887
rect 4530 6878 4534 6882
rect 4540 6878 4544 6882
rect 4550 6878 4554 6882
rect 618 6849 622 6853
rect 628 6849 632 6853
rect 638 6849 642 6853
rect 618 6844 622 6848
rect 628 6844 632 6848
rect 638 6844 642 6848
rect 618 6839 622 6843
rect 628 6839 632 6843
rect 638 6839 642 6843
rect 618 6834 622 6838
rect 628 6834 632 6838
rect 638 6834 642 6838
rect 664 6849 668 6853
rect 674 6849 678 6853
rect 684 6849 688 6853
rect 664 6844 668 6848
rect 674 6844 678 6848
rect 684 6844 688 6848
rect 664 6839 668 6843
rect 674 6839 678 6843
rect 684 6839 688 6843
rect 664 6834 668 6838
rect 674 6834 678 6838
rect 684 6834 688 6838
rect 4484 6584 4488 6588
rect 4494 6584 4498 6588
rect 4504 6584 4508 6588
rect 4484 6579 4488 6583
rect 4494 6579 4498 6583
rect 4504 6579 4508 6583
rect 4484 6574 4488 6578
rect 4494 6574 4498 6578
rect 4504 6574 4508 6578
rect 4484 6569 4488 6573
rect 4494 6569 4498 6573
rect 4504 6569 4508 6573
rect 4530 6584 4534 6588
rect 4540 6584 4544 6588
rect 4550 6584 4554 6588
rect 4530 6579 4534 6583
rect 4540 6579 4544 6583
rect 4550 6579 4554 6583
rect 4530 6574 4534 6578
rect 4540 6574 4544 6578
rect 4550 6574 4554 6578
rect 4530 6569 4534 6573
rect 4540 6569 4544 6573
rect 4550 6569 4554 6573
rect 618 6540 622 6544
rect 628 6540 632 6544
rect 638 6540 642 6544
rect 618 6535 622 6539
rect 628 6535 632 6539
rect 638 6535 642 6539
rect 618 6530 622 6534
rect 628 6530 632 6534
rect 638 6530 642 6534
rect 618 6525 622 6529
rect 628 6525 632 6529
rect 638 6525 642 6529
rect 664 6540 668 6544
rect 674 6540 678 6544
rect 684 6540 688 6544
rect 664 6535 668 6539
rect 674 6535 678 6539
rect 684 6535 688 6539
rect 664 6530 668 6534
rect 674 6530 678 6534
rect 684 6530 688 6534
rect 664 6525 668 6529
rect 674 6525 678 6529
rect 684 6525 688 6529
rect 4484 6275 4488 6279
rect 4494 6275 4498 6279
rect 4504 6275 4508 6279
rect 4484 6270 4488 6274
rect 4494 6270 4498 6274
rect 4504 6270 4508 6274
rect 4484 6265 4488 6269
rect 4494 6265 4498 6269
rect 4504 6265 4508 6269
rect 4484 6260 4488 6264
rect 4494 6260 4498 6264
rect 4504 6260 4508 6264
rect 4530 6275 4534 6279
rect 4540 6275 4544 6279
rect 4550 6275 4554 6279
rect 4530 6270 4534 6274
rect 4540 6270 4544 6274
rect 4550 6270 4554 6274
rect 4530 6265 4534 6269
rect 4540 6265 4544 6269
rect 4550 6265 4554 6269
rect 4530 6260 4534 6264
rect 4540 6260 4544 6264
rect 4550 6260 4554 6264
rect 618 6140 622 6144
rect 628 6140 632 6144
rect 638 6140 642 6144
rect 618 6135 622 6139
rect 628 6135 632 6139
rect 638 6135 642 6139
rect 618 6130 622 6134
rect 628 6130 632 6134
rect 638 6130 642 6134
rect 618 6125 622 6129
rect 628 6125 632 6129
rect 638 6125 642 6129
rect 664 6140 668 6144
rect 674 6140 678 6144
rect 684 6140 688 6144
rect 664 6135 668 6139
rect 674 6135 678 6139
rect 684 6135 688 6139
rect 664 6130 668 6134
rect 674 6130 678 6134
rect 684 6130 688 6134
rect 664 6125 668 6129
rect 674 6125 678 6129
rect 684 6125 688 6129
rect 618 6111 622 6115
rect 628 6111 632 6115
rect 638 6111 642 6115
rect 618 6106 622 6110
rect 628 6106 632 6110
rect 638 6106 642 6110
rect 618 6101 622 6105
rect 628 6101 632 6105
rect 638 6101 642 6105
rect 618 6096 622 6100
rect 628 6096 632 6100
rect 638 6096 642 6100
rect 664 6111 668 6115
rect 674 6111 678 6115
rect 684 6111 688 6115
rect 664 6106 668 6110
rect 674 6106 678 6110
rect 684 6106 688 6110
rect 664 6101 668 6105
rect 674 6101 678 6105
rect 684 6101 688 6105
rect 664 6096 668 6100
rect 674 6096 678 6100
rect 684 6096 688 6100
rect 618 6082 622 6086
rect 628 6082 632 6086
rect 638 6082 642 6086
rect 618 6077 622 6081
rect 628 6077 632 6081
rect 638 6077 642 6081
rect 618 6072 622 6076
rect 628 6072 632 6076
rect 638 6072 642 6076
rect 618 6067 622 6071
rect 628 6067 632 6071
rect 638 6067 642 6071
rect 664 6082 668 6086
rect 674 6082 678 6086
rect 684 6082 688 6086
rect 664 6077 668 6081
rect 674 6077 678 6081
rect 684 6077 688 6081
rect 664 6072 668 6076
rect 674 6072 678 6076
rect 684 6072 688 6076
rect 664 6067 668 6071
rect 674 6067 678 6071
rect 684 6067 688 6071
rect 4484 6083 4488 6087
rect 4494 6083 4498 6087
rect 4504 6083 4508 6087
rect 4484 6078 4488 6082
rect 4494 6078 4498 6082
rect 4504 6078 4508 6082
rect 4484 6073 4488 6077
rect 4494 6073 4498 6077
rect 4504 6073 4508 6077
rect 4484 6068 4488 6072
rect 4494 6068 4498 6072
rect 4504 6068 4508 6072
rect 4530 6083 4534 6087
rect 4540 6083 4544 6087
rect 4550 6083 4554 6087
rect 4530 6078 4534 6082
rect 4540 6078 4544 6082
rect 4550 6078 4554 6082
rect 4530 6073 4534 6077
rect 4540 6073 4544 6077
rect 4550 6073 4554 6077
rect 4530 6068 4534 6072
rect 4540 6068 4544 6072
rect 4550 6068 4554 6072
rect 4484 6057 4488 6061
rect 4494 6057 4498 6061
rect 4504 6057 4508 6061
rect 618 6053 622 6057
rect 628 6053 632 6057
rect 638 6053 642 6057
rect 618 6048 622 6052
rect 628 6048 632 6052
rect 638 6048 642 6052
rect 618 6043 622 6047
rect 628 6043 632 6047
rect 638 6043 642 6047
rect 618 6038 622 6042
rect 628 6038 632 6042
rect 638 6038 642 6042
rect 664 6053 668 6057
rect 674 6053 678 6057
rect 684 6053 688 6057
rect 664 6048 668 6052
rect 674 6048 678 6052
rect 684 6048 688 6052
rect 664 6043 668 6047
rect 674 6043 678 6047
rect 684 6043 688 6047
rect 4484 6052 4488 6056
rect 4494 6052 4498 6056
rect 4504 6052 4508 6056
rect 4484 6047 4488 6051
rect 4494 6047 4498 6051
rect 4504 6047 4508 6051
rect 4484 6042 4488 6046
rect 4494 6042 4498 6046
rect 4504 6042 4508 6046
rect 4530 6057 4534 6061
rect 4540 6057 4544 6061
rect 4550 6057 4554 6061
rect 4530 6052 4534 6056
rect 4540 6052 4544 6056
rect 4550 6052 4554 6056
rect 4530 6047 4534 6051
rect 4540 6047 4544 6051
rect 4550 6047 4554 6051
rect 4530 6042 4534 6046
rect 4540 6042 4544 6046
rect 4550 6042 4554 6046
rect 664 6038 668 6042
rect 674 6038 678 6042
rect 684 6038 688 6042
rect 4484 6031 4488 6035
rect 4494 6031 4498 6035
rect 4504 6031 4508 6035
rect 618 6024 622 6028
rect 628 6024 632 6028
rect 638 6024 642 6028
rect 618 6019 622 6023
rect 628 6019 632 6023
rect 638 6019 642 6023
rect 618 6014 622 6018
rect 628 6014 632 6018
rect 638 6014 642 6018
rect 618 6009 622 6013
rect 628 6009 632 6013
rect 638 6009 642 6013
rect 664 6024 668 6028
rect 674 6024 678 6028
rect 684 6024 688 6028
rect 664 6019 668 6023
rect 674 6019 678 6023
rect 684 6019 688 6023
rect 664 6014 668 6018
rect 674 6014 678 6018
rect 684 6014 688 6018
rect 4484 6026 4488 6030
rect 4494 6026 4498 6030
rect 4504 6026 4508 6030
rect 4484 6021 4488 6025
rect 4494 6021 4498 6025
rect 4504 6021 4508 6025
rect 4484 6016 4488 6020
rect 4494 6016 4498 6020
rect 4504 6016 4508 6020
rect 4530 6031 4534 6035
rect 4540 6031 4544 6035
rect 4550 6031 4554 6035
rect 4530 6026 4534 6030
rect 4540 6026 4544 6030
rect 4550 6026 4554 6030
rect 4530 6021 4534 6025
rect 4540 6021 4544 6025
rect 4550 6021 4554 6025
rect 4530 6016 4534 6020
rect 4540 6016 4544 6020
rect 4550 6016 4554 6020
rect 664 6009 668 6013
rect 674 6009 678 6013
rect 684 6009 688 6013
rect 4484 6005 4488 6009
rect 4494 6005 4498 6009
rect 4504 6005 4508 6009
rect 4484 6000 4488 6004
rect 4494 6000 4498 6004
rect 4504 6000 4508 6004
rect 4484 5995 4488 5999
rect 4494 5995 4498 5999
rect 4504 5995 4508 5999
rect 4484 5990 4488 5994
rect 4494 5990 4498 5994
rect 4504 5990 4508 5994
rect 4530 6005 4534 6009
rect 4540 6005 4544 6009
rect 4550 6005 4554 6009
rect 4530 6000 4534 6004
rect 4540 6000 4544 6004
rect 4550 6000 4554 6004
rect 4530 5995 4534 5999
rect 4540 5995 4544 5999
rect 4550 5995 4554 5999
rect 4530 5990 4534 5994
rect 4540 5990 4544 5994
rect 4550 5990 4554 5994
rect 4484 5979 4488 5983
rect 4494 5979 4498 5983
rect 4504 5979 4508 5983
rect 757 5891 761 5895
rect 762 5891 766 5895
rect 767 5891 771 5895
rect 772 5891 776 5895
rect 757 5881 761 5885
rect 762 5881 766 5885
rect 767 5881 771 5885
rect 772 5881 776 5885
rect 757 5871 761 5875
rect 762 5871 766 5875
rect 767 5871 771 5875
rect 772 5871 776 5875
rect 783 5891 787 5895
rect 788 5891 792 5895
rect 793 5891 797 5895
rect 798 5891 802 5895
rect 783 5881 787 5885
rect 788 5881 792 5885
rect 793 5881 797 5885
rect 798 5881 802 5885
rect 783 5871 787 5875
rect 788 5871 792 5875
rect 793 5871 797 5875
rect 798 5871 802 5875
rect 809 5891 813 5895
rect 814 5891 818 5895
rect 819 5891 823 5895
rect 824 5891 828 5895
rect 809 5881 813 5885
rect 814 5881 818 5885
rect 819 5881 823 5885
rect 824 5881 828 5885
rect 809 5871 813 5875
rect 814 5871 818 5875
rect 819 5871 823 5875
rect 824 5871 828 5875
rect 835 5891 839 5895
rect 840 5891 844 5895
rect 845 5891 849 5895
rect 850 5891 854 5895
rect 835 5881 839 5885
rect 840 5881 844 5885
rect 845 5881 849 5885
rect 850 5881 854 5885
rect 835 5871 839 5875
rect 840 5871 844 5875
rect 845 5871 849 5875
rect 850 5871 854 5875
rect 861 5891 865 5895
rect 866 5891 870 5895
rect 871 5891 875 5895
rect 876 5891 880 5895
rect 861 5881 865 5885
rect 866 5881 870 5885
rect 871 5881 875 5885
rect 876 5881 880 5885
rect 861 5871 865 5875
rect 866 5871 870 5875
rect 871 5871 875 5875
rect 876 5871 880 5875
rect 1054 5891 1058 5895
rect 1059 5891 1063 5895
rect 1064 5891 1068 5895
rect 1069 5891 1073 5895
rect 1054 5881 1058 5885
rect 1059 5881 1063 5885
rect 1064 5881 1068 5885
rect 1069 5881 1073 5885
rect 1054 5871 1058 5875
rect 1059 5871 1063 5875
rect 1064 5871 1068 5875
rect 1069 5871 1073 5875
rect 757 5845 761 5849
rect 762 5845 766 5849
rect 767 5845 771 5849
rect 772 5845 776 5849
rect 757 5835 761 5839
rect 762 5835 766 5839
rect 767 5835 771 5839
rect 772 5835 776 5839
rect 757 5825 761 5829
rect 762 5825 766 5829
rect 767 5825 771 5829
rect 772 5825 776 5829
rect 783 5845 787 5849
rect 788 5845 792 5849
rect 793 5845 797 5849
rect 798 5845 802 5849
rect 783 5835 787 5839
rect 788 5835 792 5839
rect 793 5835 797 5839
rect 798 5835 802 5839
rect 783 5825 787 5829
rect 788 5825 792 5829
rect 793 5825 797 5829
rect 798 5825 802 5829
rect 809 5845 813 5849
rect 814 5845 818 5849
rect 819 5845 823 5849
rect 824 5845 828 5849
rect 809 5835 813 5839
rect 814 5835 818 5839
rect 819 5835 823 5839
rect 824 5835 828 5839
rect 809 5825 813 5829
rect 814 5825 818 5829
rect 819 5825 823 5829
rect 824 5825 828 5829
rect 835 5845 839 5849
rect 840 5845 844 5849
rect 845 5845 849 5849
rect 850 5845 854 5849
rect 835 5835 839 5839
rect 840 5835 844 5839
rect 845 5835 849 5839
rect 850 5835 854 5839
rect 835 5825 839 5829
rect 840 5825 844 5829
rect 845 5825 849 5829
rect 850 5825 854 5829
rect 861 5845 865 5849
rect 866 5845 870 5849
rect 871 5845 875 5849
rect 876 5845 880 5849
rect 861 5835 865 5839
rect 866 5835 870 5839
rect 871 5835 875 5839
rect 876 5835 880 5839
rect 861 5825 865 5829
rect 866 5825 870 5829
rect 871 5825 875 5829
rect 876 5825 880 5829
rect 1054 5845 1058 5849
rect 1059 5845 1063 5849
rect 1064 5845 1068 5849
rect 1069 5845 1073 5849
rect 1054 5835 1058 5839
rect 1059 5835 1063 5839
rect 1064 5835 1068 5839
rect 1069 5835 1073 5839
rect 1054 5825 1058 5829
rect 1059 5825 1063 5829
rect 1064 5825 1068 5829
rect 1069 5825 1073 5829
rect 1363 5891 1367 5895
rect 1368 5891 1372 5895
rect 1373 5891 1377 5895
rect 1378 5891 1382 5895
rect 1363 5881 1367 5885
rect 1368 5881 1372 5885
rect 1373 5881 1377 5885
rect 1378 5881 1382 5885
rect 1363 5871 1367 5875
rect 1368 5871 1372 5875
rect 1373 5871 1377 5875
rect 1378 5871 1382 5875
rect 1363 5845 1367 5849
rect 1368 5845 1372 5849
rect 1373 5845 1377 5849
rect 1378 5845 1382 5849
rect 1363 5835 1367 5839
rect 1368 5835 1372 5839
rect 1373 5835 1377 5839
rect 1378 5835 1382 5839
rect 1363 5825 1367 5829
rect 1368 5825 1372 5829
rect 1373 5825 1377 5829
rect 1378 5825 1382 5829
rect 1672 5891 1676 5895
rect 1677 5891 1681 5895
rect 1682 5891 1686 5895
rect 1687 5891 1691 5895
rect 1672 5881 1676 5885
rect 1677 5881 1681 5885
rect 1682 5881 1686 5885
rect 1687 5881 1691 5885
rect 1672 5871 1676 5875
rect 1677 5871 1681 5875
rect 1682 5871 1686 5875
rect 1687 5871 1691 5875
rect 1672 5845 1676 5849
rect 1677 5845 1681 5849
rect 1682 5845 1686 5849
rect 1687 5845 1691 5849
rect 1672 5835 1676 5839
rect 1677 5835 1681 5839
rect 1682 5835 1686 5839
rect 1687 5835 1691 5839
rect 1672 5825 1676 5829
rect 1677 5825 1681 5829
rect 1682 5825 1686 5829
rect 1687 5825 1691 5829
rect 1981 5891 1985 5895
rect 1986 5891 1990 5895
rect 1991 5891 1995 5895
rect 1996 5891 2000 5895
rect 1981 5881 1985 5885
rect 1986 5881 1990 5885
rect 1991 5881 1995 5885
rect 1996 5881 2000 5885
rect 1981 5871 1985 5875
rect 1986 5871 1990 5875
rect 1991 5871 1995 5875
rect 1996 5871 2000 5875
rect 1981 5845 1985 5849
rect 1986 5845 1990 5849
rect 1991 5845 1995 5849
rect 1996 5845 2000 5849
rect 1981 5835 1985 5839
rect 1986 5835 1990 5839
rect 1991 5835 1995 5839
rect 1996 5835 2000 5839
rect 1981 5825 1985 5829
rect 1986 5825 1990 5829
rect 1991 5825 1995 5829
rect 1996 5825 2000 5829
rect 2290 5891 2294 5895
rect 2295 5891 2299 5895
rect 2300 5891 2304 5895
rect 2305 5891 2309 5895
rect 2290 5881 2294 5885
rect 2295 5881 2299 5885
rect 2300 5881 2304 5885
rect 2305 5881 2309 5885
rect 2290 5871 2294 5875
rect 2295 5871 2299 5875
rect 2300 5871 2304 5875
rect 2305 5871 2309 5875
rect 2290 5845 2294 5849
rect 2295 5845 2299 5849
rect 2300 5845 2304 5849
rect 2305 5845 2309 5849
rect 2290 5835 2294 5839
rect 2295 5835 2299 5839
rect 2300 5835 2304 5839
rect 2305 5835 2309 5839
rect 2290 5825 2294 5829
rect 2295 5825 2299 5829
rect 2300 5825 2304 5829
rect 2305 5825 2309 5829
rect 2599 5891 2603 5895
rect 2604 5891 2608 5895
rect 2609 5891 2613 5895
rect 2614 5891 2618 5895
rect 2599 5881 2603 5885
rect 2604 5881 2608 5885
rect 2609 5881 2613 5885
rect 2614 5881 2618 5885
rect 2599 5871 2603 5875
rect 2604 5871 2608 5875
rect 2609 5871 2613 5875
rect 2614 5871 2618 5875
rect 2599 5845 2603 5849
rect 2604 5845 2608 5849
rect 2609 5845 2613 5849
rect 2614 5845 2618 5849
rect 2599 5835 2603 5839
rect 2604 5835 2608 5839
rect 2609 5835 2613 5839
rect 2614 5835 2618 5839
rect 2599 5825 2603 5829
rect 2604 5825 2608 5829
rect 2609 5825 2613 5829
rect 2614 5825 2618 5829
rect 2908 5891 2912 5895
rect 2913 5891 2917 5895
rect 2918 5891 2922 5895
rect 2923 5891 2927 5895
rect 2908 5881 2912 5885
rect 2913 5881 2917 5885
rect 2918 5881 2922 5885
rect 2923 5881 2927 5885
rect 2908 5871 2912 5875
rect 2913 5871 2917 5875
rect 2918 5871 2922 5875
rect 2923 5871 2927 5875
rect 2908 5845 2912 5849
rect 2913 5845 2917 5849
rect 2918 5845 2922 5849
rect 2923 5845 2927 5849
rect 2908 5835 2912 5839
rect 2913 5835 2917 5839
rect 2918 5835 2922 5839
rect 2923 5835 2927 5839
rect 2908 5825 2912 5829
rect 2913 5825 2917 5829
rect 2918 5825 2922 5829
rect 2923 5825 2927 5829
rect 3217 5891 3221 5895
rect 3222 5891 3226 5895
rect 3227 5891 3231 5895
rect 3232 5891 3236 5895
rect 3217 5881 3221 5885
rect 3222 5881 3226 5885
rect 3227 5881 3231 5885
rect 3232 5881 3236 5885
rect 3217 5871 3221 5875
rect 3222 5871 3226 5875
rect 3227 5871 3231 5875
rect 3232 5871 3236 5875
rect 3217 5845 3221 5849
rect 3222 5845 3226 5849
rect 3227 5845 3231 5849
rect 3232 5845 3236 5849
rect 3217 5835 3221 5839
rect 3222 5835 3226 5839
rect 3227 5835 3231 5839
rect 3232 5835 3236 5839
rect 3217 5825 3221 5829
rect 3222 5825 3226 5829
rect 3227 5825 3231 5829
rect 3232 5825 3236 5829
rect 3526 5891 3530 5895
rect 3531 5891 3535 5895
rect 3536 5891 3540 5895
rect 3541 5891 3545 5895
rect 3526 5881 3530 5885
rect 3531 5881 3535 5885
rect 3536 5881 3540 5885
rect 3541 5881 3545 5885
rect 3526 5871 3530 5875
rect 3531 5871 3535 5875
rect 3536 5871 3540 5875
rect 3541 5871 3545 5875
rect 3526 5845 3530 5849
rect 3531 5845 3535 5849
rect 3536 5845 3540 5849
rect 3541 5845 3545 5849
rect 3526 5835 3530 5839
rect 3531 5835 3535 5839
rect 3536 5835 3540 5839
rect 3541 5835 3545 5839
rect 3526 5825 3530 5829
rect 3531 5825 3535 5829
rect 3536 5825 3540 5829
rect 3541 5825 3545 5829
rect 3835 5891 3839 5895
rect 3840 5891 3844 5895
rect 3845 5891 3849 5895
rect 3850 5891 3854 5895
rect 3835 5881 3839 5885
rect 3840 5881 3844 5885
rect 3845 5881 3849 5885
rect 3850 5881 3854 5885
rect 3835 5871 3839 5875
rect 3840 5871 3844 5875
rect 3845 5871 3849 5875
rect 3850 5871 3854 5875
rect 3835 5845 3839 5849
rect 3840 5845 3844 5849
rect 3845 5845 3849 5849
rect 3850 5845 3854 5849
rect 3835 5835 3839 5839
rect 3840 5835 3844 5839
rect 3845 5835 3849 5839
rect 3850 5835 3854 5839
rect 3835 5825 3839 5829
rect 3840 5825 3844 5829
rect 3845 5825 3849 5829
rect 3850 5825 3854 5829
rect 4484 5974 4488 5978
rect 4494 5974 4498 5978
rect 4504 5974 4508 5978
rect 4484 5969 4488 5973
rect 4494 5969 4498 5973
rect 4504 5969 4508 5973
rect 4484 5964 4488 5968
rect 4494 5964 4498 5968
rect 4504 5964 4508 5968
rect 4530 5979 4534 5983
rect 4540 5979 4544 5983
rect 4550 5979 4554 5983
rect 4530 5974 4534 5978
rect 4540 5974 4544 5978
rect 4550 5974 4554 5978
rect 4530 5969 4534 5973
rect 4540 5969 4544 5973
rect 4550 5969 4554 5973
rect 4530 5964 4534 5968
rect 4540 5964 4544 5968
rect 4550 5964 4554 5968
rect 4235 5891 4239 5895
rect 4240 5891 4244 5895
rect 4245 5891 4249 5895
rect 4250 5891 4254 5895
rect 4235 5881 4239 5885
rect 4240 5881 4244 5885
rect 4245 5881 4249 5885
rect 4250 5881 4254 5885
rect 4235 5871 4239 5875
rect 4240 5871 4244 5875
rect 4245 5871 4249 5875
rect 4250 5871 4254 5875
rect 4264 5891 4268 5895
rect 4269 5891 4273 5895
rect 4274 5891 4278 5895
rect 4279 5891 4283 5895
rect 4264 5881 4268 5885
rect 4269 5881 4273 5885
rect 4274 5881 4278 5885
rect 4279 5881 4283 5885
rect 4264 5871 4268 5875
rect 4269 5871 4273 5875
rect 4274 5871 4278 5875
rect 4279 5871 4283 5875
rect 4293 5891 4297 5895
rect 4298 5891 4302 5895
rect 4303 5891 4307 5895
rect 4308 5891 4312 5895
rect 4293 5881 4297 5885
rect 4298 5881 4302 5885
rect 4303 5881 4307 5885
rect 4308 5881 4312 5885
rect 4293 5871 4297 5875
rect 4298 5871 4302 5875
rect 4303 5871 4307 5875
rect 4308 5871 4312 5875
rect 4322 5891 4326 5895
rect 4327 5891 4331 5895
rect 4332 5891 4336 5895
rect 4337 5891 4341 5895
rect 4322 5881 4326 5885
rect 4327 5881 4331 5885
rect 4332 5881 4336 5885
rect 4337 5881 4341 5885
rect 4322 5871 4326 5875
rect 4327 5871 4331 5875
rect 4332 5871 4336 5875
rect 4337 5871 4341 5875
rect 4351 5891 4355 5895
rect 4356 5891 4360 5895
rect 4361 5891 4365 5895
rect 4366 5891 4370 5895
rect 4351 5881 4355 5885
rect 4356 5881 4360 5885
rect 4361 5881 4365 5885
rect 4366 5881 4370 5885
rect 4351 5871 4355 5875
rect 4356 5871 4360 5875
rect 4361 5871 4365 5875
rect 4366 5871 4370 5875
rect 4235 5845 4239 5849
rect 4240 5845 4244 5849
rect 4245 5845 4249 5849
rect 4250 5845 4254 5849
rect 4235 5835 4239 5839
rect 4240 5835 4244 5839
rect 4245 5835 4249 5839
rect 4250 5835 4254 5839
rect 4235 5825 4239 5829
rect 4240 5825 4244 5829
rect 4245 5825 4249 5829
rect 4250 5825 4254 5829
rect 4264 5845 4268 5849
rect 4269 5845 4273 5849
rect 4274 5845 4278 5849
rect 4279 5845 4283 5849
rect 4264 5835 4268 5839
rect 4269 5835 4273 5839
rect 4274 5835 4278 5839
rect 4279 5835 4283 5839
rect 4264 5825 4268 5829
rect 4269 5825 4273 5829
rect 4274 5825 4278 5829
rect 4279 5825 4283 5829
rect 4293 5845 4297 5849
rect 4298 5845 4302 5849
rect 4303 5845 4307 5849
rect 4308 5845 4312 5849
rect 4293 5835 4297 5839
rect 4298 5835 4302 5839
rect 4303 5835 4307 5839
rect 4308 5835 4312 5839
rect 4293 5825 4297 5829
rect 4298 5825 4302 5829
rect 4303 5825 4307 5829
rect 4308 5825 4312 5829
rect 4322 5845 4326 5849
rect 4327 5845 4331 5849
rect 4332 5845 4336 5849
rect 4337 5845 4341 5849
rect 4322 5835 4326 5839
rect 4327 5835 4331 5839
rect 4332 5835 4336 5839
rect 4337 5835 4341 5839
rect 4322 5825 4326 5829
rect 4327 5825 4331 5829
rect 4332 5825 4336 5829
rect 4337 5825 4341 5829
rect 4351 5845 4355 5849
rect 4356 5845 4360 5849
rect 4361 5845 4365 5849
rect 4366 5845 4370 5849
rect 4351 5835 4355 5839
rect 4356 5835 4360 5839
rect 4361 5835 4365 5839
rect 4366 5835 4370 5839
rect 4351 5825 4355 5829
rect 4356 5825 4360 5829
rect 4361 5825 4365 5829
rect 4366 5825 4370 5829
<< metal2 >>
rect 1060 10290 1320 10293
rect 118 9786 1024 10280
rect 1060 10036 1063 10290
rect 1317 10036 1320 10290
rect 1060 10033 1320 10036
rect 1369 10290 1629 10293
rect 1369 10036 1372 10290
rect 1626 10036 1629 10290
rect 1369 10033 1629 10036
rect 1678 10290 1938 10293
rect 1678 10036 1681 10290
rect 1935 10036 1938 10290
rect 1678 10033 1938 10036
rect 1987 10290 2247 10293
rect 1987 10036 1990 10290
rect 2244 10036 2247 10290
rect 1987 10033 2247 10036
rect 2296 10290 2556 10293
rect 2296 10036 2299 10290
rect 2553 10036 2556 10290
rect 2296 10033 2556 10036
rect 2605 10290 2865 10293
rect 2605 10036 2608 10290
rect 2862 10036 2865 10290
rect 2605 10033 2865 10036
rect 2914 10290 3174 10293
rect 2914 10036 2917 10290
rect 3171 10036 3174 10290
rect 2914 10033 3174 10036
rect 3223 10290 3483 10293
rect 3223 10036 3226 10290
rect 3480 10036 3483 10290
rect 3223 10033 3483 10036
rect 3532 10290 3792 10293
rect 3532 10036 3535 10290
rect 3789 10036 3792 10290
rect 3532 10033 3792 10036
rect 3841 10290 4101 10293
rect 3841 10036 3844 10290
rect 4098 10036 4101 10290
rect 3841 10033 4101 10036
rect 1441 10001 1557 10002
rect 1441 9997 1454 10001
rect 1458 9997 1461 10001
rect 1465 9997 1468 10001
rect 1472 9997 1475 10001
rect 1479 9997 1482 10001
rect 1486 9997 1489 10001
rect 1493 9997 1496 10001
rect 1500 9997 1503 10001
rect 1507 9997 1510 10001
rect 1514 9997 1517 10001
rect 1521 9997 1524 10001
rect 1528 9997 1531 10001
rect 1535 9997 1538 10001
rect 1542 9997 1557 10001
rect 1441 9996 1557 9997
rect 1441 9993 1454 9996
rect 1451 9992 1454 9993
rect 1458 9992 1461 9996
rect 1465 9992 1468 9996
rect 1472 9992 1475 9996
rect 1479 9992 1482 9996
rect 1486 9992 1489 9996
rect 1493 9992 1496 9996
rect 1500 9992 1503 9996
rect 1507 9992 1510 9996
rect 1514 9992 1517 9996
rect 1521 9992 1524 9996
rect 1528 9992 1531 9996
rect 1535 9992 1538 9996
rect 1542 9993 1557 9996
rect 1750 10001 1866 10002
rect 1750 9997 1763 10001
rect 1767 9997 1770 10001
rect 1774 9997 1777 10001
rect 1781 9997 1784 10001
rect 1788 9997 1791 10001
rect 1795 9997 1798 10001
rect 1802 9997 1805 10001
rect 1809 9997 1812 10001
rect 1816 9997 1819 10001
rect 1823 9997 1826 10001
rect 1830 9997 1833 10001
rect 1837 9997 1840 10001
rect 1844 9997 1847 10001
rect 1851 9997 1866 10001
rect 1750 9996 1866 9997
rect 1750 9993 1763 9996
rect 1542 9992 1547 9993
rect 1451 9991 1547 9992
rect 1451 9987 1454 9991
rect 1458 9987 1461 9991
rect 1465 9987 1468 9991
rect 1472 9987 1475 9991
rect 1479 9987 1482 9991
rect 1486 9987 1489 9991
rect 1493 9987 1496 9991
rect 1500 9987 1503 9991
rect 1507 9987 1510 9991
rect 1514 9987 1517 9991
rect 1521 9987 1524 9991
rect 1528 9987 1531 9991
rect 1535 9987 1538 9991
rect 1542 9987 1547 9991
rect 1451 9986 1547 9987
rect 1451 9982 1454 9986
rect 1458 9982 1461 9986
rect 1465 9982 1468 9986
rect 1472 9982 1475 9986
rect 1479 9982 1482 9986
rect 1486 9982 1489 9986
rect 1493 9982 1496 9986
rect 1500 9982 1503 9986
rect 1507 9982 1510 9986
rect 1514 9982 1517 9986
rect 1521 9982 1524 9986
rect 1528 9982 1531 9986
rect 1535 9982 1538 9986
rect 1542 9982 1547 9986
rect 1451 9953 1547 9982
rect 1760 9992 1763 9993
rect 1767 9992 1770 9996
rect 1774 9992 1777 9996
rect 1781 9992 1784 9996
rect 1788 9992 1791 9996
rect 1795 9992 1798 9996
rect 1802 9992 1805 9996
rect 1809 9992 1812 9996
rect 1816 9992 1819 9996
rect 1823 9992 1826 9996
rect 1830 9992 1833 9996
rect 1837 9992 1840 9996
rect 1844 9992 1847 9996
rect 1851 9993 1866 9996
rect 2059 10001 2175 10002
rect 2059 9997 2072 10001
rect 2076 9997 2079 10001
rect 2083 9997 2086 10001
rect 2090 9997 2093 10001
rect 2097 9997 2100 10001
rect 2104 9997 2107 10001
rect 2111 9997 2114 10001
rect 2118 9997 2121 10001
rect 2125 9997 2128 10001
rect 2132 9997 2135 10001
rect 2139 9997 2142 10001
rect 2146 9997 2149 10001
rect 2153 9997 2156 10001
rect 2160 9997 2175 10001
rect 2059 9996 2175 9997
rect 2059 9993 2072 9996
rect 1851 9992 1856 9993
rect 1760 9991 1856 9992
rect 1760 9987 1763 9991
rect 1767 9987 1770 9991
rect 1774 9987 1777 9991
rect 1781 9987 1784 9991
rect 1788 9987 1791 9991
rect 1795 9987 1798 9991
rect 1802 9987 1805 9991
rect 1809 9987 1812 9991
rect 1816 9987 1819 9991
rect 1823 9987 1826 9991
rect 1830 9987 1833 9991
rect 1837 9987 1840 9991
rect 1844 9987 1847 9991
rect 1851 9987 1856 9991
rect 1760 9986 1856 9987
rect 1760 9982 1763 9986
rect 1767 9982 1770 9986
rect 1774 9982 1777 9986
rect 1781 9982 1784 9986
rect 1788 9982 1791 9986
rect 1795 9982 1798 9986
rect 1802 9982 1805 9986
rect 1809 9982 1812 9986
rect 1816 9982 1819 9986
rect 1823 9982 1826 9986
rect 1830 9982 1833 9986
rect 1837 9982 1840 9986
rect 1844 9982 1847 9986
rect 1851 9982 1856 9986
rect 1760 9953 1856 9982
rect 2069 9992 2072 9993
rect 2076 9992 2079 9996
rect 2083 9992 2086 9996
rect 2090 9992 2093 9996
rect 2097 9992 2100 9996
rect 2104 9992 2107 9996
rect 2111 9992 2114 9996
rect 2118 9992 2121 9996
rect 2125 9992 2128 9996
rect 2132 9992 2135 9996
rect 2139 9992 2142 9996
rect 2146 9992 2149 9996
rect 2153 9992 2156 9996
rect 2160 9993 2175 9996
rect 2368 10001 2484 10002
rect 2368 9997 2381 10001
rect 2385 9997 2388 10001
rect 2392 9997 2395 10001
rect 2399 9997 2402 10001
rect 2406 9997 2409 10001
rect 2413 9997 2416 10001
rect 2420 9997 2423 10001
rect 2427 9997 2430 10001
rect 2434 9997 2437 10001
rect 2441 9997 2444 10001
rect 2448 9997 2451 10001
rect 2455 9997 2458 10001
rect 2462 9997 2465 10001
rect 2469 9997 2484 10001
rect 2368 9996 2484 9997
rect 2368 9993 2381 9996
rect 2160 9992 2165 9993
rect 2069 9991 2165 9992
rect 2069 9987 2072 9991
rect 2076 9987 2079 9991
rect 2083 9987 2086 9991
rect 2090 9987 2093 9991
rect 2097 9987 2100 9991
rect 2104 9987 2107 9991
rect 2111 9987 2114 9991
rect 2118 9987 2121 9991
rect 2125 9987 2128 9991
rect 2132 9987 2135 9991
rect 2139 9987 2142 9991
rect 2146 9987 2149 9991
rect 2153 9987 2156 9991
rect 2160 9987 2165 9991
rect 2069 9986 2165 9987
rect 2069 9982 2072 9986
rect 2076 9982 2079 9986
rect 2083 9982 2086 9986
rect 2090 9982 2093 9986
rect 2097 9982 2100 9986
rect 2104 9982 2107 9986
rect 2111 9982 2114 9986
rect 2118 9982 2121 9986
rect 2125 9982 2128 9986
rect 2132 9982 2135 9986
rect 2139 9982 2142 9986
rect 2146 9982 2149 9986
rect 2153 9982 2156 9986
rect 2160 9982 2165 9986
rect 2069 9953 2165 9982
rect 2378 9992 2381 9993
rect 2385 9992 2388 9996
rect 2392 9992 2395 9996
rect 2399 9992 2402 9996
rect 2406 9992 2409 9996
rect 2413 9992 2416 9996
rect 2420 9992 2423 9996
rect 2427 9992 2430 9996
rect 2434 9992 2437 9996
rect 2441 9992 2444 9996
rect 2448 9992 2451 9996
rect 2455 9992 2458 9996
rect 2462 9992 2465 9996
rect 2469 9993 2484 9996
rect 2677 10001 2793 10002
rect 2677 9997 2690 10001
rect 2694 9997 2697 10001
rect 2701 9997 2704 10001
rect 2708 9997 2711 10001
rect 2715 9997 2718 10001
rect 2722 9997 2725 10001
rect 2729 9997 2732 10001
rect 2736 9997 2739 10001
rect 2743 9997 2746 10001
rect 2750 9997 2753 10001
rect 2757 9997 2760 10001
rect 2764 9997 2767 10001
rect 2771 9997 2774 10001
rect 2778 9997 2793 10001
rect 2677 9996 2793 9997
rect 2677 9993 2690 9996
rect 2469 9992 2474 9993
rect 2378 9991 2474 9992
rect 2378 9987 2381 9991
rect 2385 9987 2388 9991
rect 2392 9987 2395 9991
rect 2399 9987 2402 9991
rect 2406 9987 2409 9991
rect 2413 9987 2416 9991
rect 2420 9987 2423 9991
rect 2427 9987 2430 9991
rect 2434 9987 2437 9991
rect 2441 9987 2444 9991
rect 2448 9987 2451 9991
rect 2455 9987 2458 9991
rect 2462 9987 2465 9991
rect 2469 9987 2474 9991
rect 2378 9986 2474 9987
rect 2378 9982 2381 9986
rect 2385 9982 2388 9986
rect 2392 9982 2395 9986
rect 2399 9982 2402 9986
rect 2406 9982 2409 9986
rect 2413 9982 2416 9986
rect 2420 9982 2423 9986
rect 2427 9982 2430 9986
rect 2434 9982 2437 9986
rect 2441 9982 2444 9986
rect 2448 9982 2451 9986
rect 2455 9982 2458 9986
rect 2462 9982 2465 9986
rect 2469 9982 2474 9986
rect 2378 9953 2474 9982
rect 2687 9992 2690 9993
rect 2694 9992 2697 9996
rect 2701 9992 2704 9996
rect 2708 9992 2711 9996
rect 2715 9992 2718 9996
rect 2722 9992 2725 9996
rect 2729 9992 2732 9996
rect 2736 9992 2739 9996
rect 2743 9992 2746 9996
rect 2750 9992 2753 9996
rect 2757 9992 2760 9996
rect 2764 9992 2767 9996
rect 2771 9992 2774 9996
rect 2778 9993 2793 9996
rect 2986 10001 3102 10002
rect 2986 9997 2999 10001
rect 3003 9997 3006 10001
rect 3010 9997 3013 10001
rect 3017 9997 3020 10001
rect 3024 9997 3027 10001
rect 3031 9997 3034 10001
rect 3038 9997 3041 10001
rect 3045 9997 3048 10001
rect 3052 9997 3055 10001
rect 3059 9997 3062 10001
rect 3066 9997 3069 10001
rect 3073 9997 3076 10001
rect 3080 9997 3083 10001
rect 3087 9997 3102 10001
rect 2986 9996 3102 9997
rect 2986 9993 2999 9996
rect 2778 9992 2783 9993
rect 2687 9991 2783 9992
rect 2687 9987 2690 9991
rect 2694 9987 2697 9991
rect 2701 9987 2704 9991
rect 2708 9987 2711 9991
rect 2715 9987 2718 9991
rect 2722 9987 2725 9991
rect 2729 9987 2732 9991
rect 2736 9987 2739 9991
rect 2743 9987 2746 9991
rect 2750 9987 2753 9991
rect 2757 9987 2760 9991
rect 2764 9987 2767 9991
rect 2771 9987 2774 9991
rect 2778 9987 2783 9991
rect 2687 9986 2783 9987
rect 2687 9982 2690 9986
rect 2694 9982 2697 9986
rect 2701 9982 2704 9986
rect 2708 9982 2711 9986
rect 2715 9982 2718 9986
rect 2722 9982 2725 9986
rect 2729 9982 2732 9986
rect 2736 9982 2739 9986
rect 2743 9982 2746 9986
rect 2750 9982 2753 9986
rect 2757 9982 2760 9986
rect 2764 9982 2767 9986
rect 2771 9982 2774 9986
rect 2778 9982 2783 9986
rect 2687 9953 2783 9982
rect 2996 9992 2999 9993
rect 3003 9992 3006 9996
rect 3010 9992 3013 9996
rect 3017 9992 3020 9996
rect 3024 9992 3027 9996
rect 3031 9992 3034 9996
rect 3038 9992 3041 9996
rect 3045 9992 3048 9996
rect 3052 9992 3055 9996
rect 3059 9992 3062 9996
rect 3066 9992 3069 9996
rect 3073 9992 3076 9996
rect 3080 9992 3083 9996
rect 3087 9993 3102 9996
rect 3295 10001 3411 10002
rect 3295 9997 3308 10001
rect 3312 9997 3315 10001
rect 3319 9997 3322 10001
rect 3326 9997 3329 10001
rect 3333 9997 3336 10001
rect 3340 9997 3343 10001
rect 3347 9997 3350 10001
rect 3354 9997 3357 10001
rect 3361 9997 3364 10001
rect 3368 9997 3371 10001
rect 3375 9997 3378 10001
rect 3382 9997 3385 10001
rect 3389 9997 3392 10001
rect 3396 9997 3411 10001
rect 3295 9996 3411 9997
rect 3295 9993 3308 9996
rect 3087 9992 3092 9993
rect 2996 9991 3092 9992
rect 2996 9987 2999 9991
rect 3003 9987 3006 9991
rect 3010 9987 3013 9991
rect 3017 9987 3020 9991
rect 3024 9987 3027 9991
rect 3031 9987 3034 9991
rect 3038 9987 3041 9991
rect 3045 9987 3048 9991
rect 3052 9987 3055 9991
rect 3059 9987 3062 9991
rect 3066 9987 3069 9991
rect 3073 9987 3076 9991
rect 3080 9987 3083 9991
rect 3087 9987 3092 9991
rect 2996 9986 3092 9987
rect 2996 9982 2999 9986
rect 3003 9982 3006 9986
rect 3010 9982 3013 9986
rect 3017 9982 3020 9986
rect 3024 9982 3027 9986
rect 3031 9982 3034 9986
rect 3038 9982 3041 9986
rect 3045 9982 3048 9986
rect 3052 9982 3055 9986
rect 3059 9982 3062 9986
rect 3066 9982 3069 9986
rect 3073 9982 3076 9986
rect 3080 9982 3083 9986
rect 3087 9982 3092 9986
rect 2996 9953 3092 9982
rect 3305 9992 3308 9993
rect 3312 9992 3315 9996
rect 3319 9992 3322 9996
rect 3326 9992 3329 9996
rect 3333 9992 3336 9996
rect 3340 9992 3343 9996
rect 3347 9992 3350 9996
rect 3354 9992 3357 9996
rect 3361 9992 3364 9996
rect 3368 9992 3371 9996
rect 3375 9992 3378 9996
rect 3382 9992 3385 9996
rect 3389 9992 3392 9996
rect 3396 9993 3411 9996
rect 3604 10001 3720 10002
rect 3604 9997 3617 10001
rect 3621 9997 3624 10001
rect 3628 9997 3631 10001
rect 3635 9997 3638 10001
rect 3642 9997 3645 10001
rect 3649 9997 3652 10001
rect 3656 9997 3659 10001
rect 3663 9997 3666 10001
rect 3670 9997 3673 10001
rect 3677 9997 3680 10001
rect 3684 9997 3687 10001
rect 3691 9997 3694 10001
rect 3698 9997 3701 10001
rect 3705 9997 3720 10001
rect 3604 9996 3720 9997
rect 3604 9993 3617 9996
rect 3396 9992 3401 9993
rect 3305 9991 3401 9992
rect 3305 9987 3308 9991
rect 3312 9987 3315 9991
rect 3319 9987 3322 9991
rect 3326 9987 3329 9991
rect 3333 9987 3336 9991
rect 3340 9987 3343 9991
rect 3347 9987 3350 9991
rect 3354 9987 3357 9991
rect 3361 9987 3364 9991
rect 3368 9987 3371 9991
rect 3375 9987 3378 9991
rect 3382 9987 3385 9991
rect 3389 9987 3392 9991
rect 3396 9987 3401 9991
rect 3305 9986 3401 9987
rect 3305 9982 3308 9986
rect 3312 9982 3315 9986
rect 3319 9982 3322 9986
rect 3326 9982 3329 9986
rect 3333 9982 3336 9986
rect 3340 9982 3343 9986
rect 3347 9982 3350 9986
rect 3354 9982 3357 9986
rect 3361 9982 3364 9986
rect 3368 9982 3371 9986
rect 3375 9982 3378 9986
rect 3382 9982 3385 9986
rect 3389 9982 3392 9986
rect 3396 9982 3401 9986
rect 3305 9953 3401 9982
rect 3614 9992 3617 9993
rect 3621 9992 3624 9996
rect 3628 9992 3631 9996
rect 3635 9992 3638 9996
rect 3642 9992 3645 9996
rect 3649 9992 3652 9996
rect 3656 9992 3659 9996
rect 3663 9992 3666 9996
rect 3670 9992 3673 9996
rect 3677 9992 3680 9996
rect 3684 9992 3687 9996
rect 3691 9992 3694 9996
rect 3698 9992 3701 9996
rect 3705 9993 3720 9996
rect 3913 10001 4029 10002
rect 3913 9997 3926 10001
rect 3930 9997 3933 10001
rect 3937 9997 3940 10001
rect 3944 9997 3947 10001
rect 3951 9997 3954 10001
rect 3958 9997 3961 10001
rect 3965 9997 3968 10001
rect 3972 9997 3975 10001
rect 3979 9997 3982 10001
rect 3986 9997 3989 10001
rect 3993 9997 3996 10001
rect 4000 9997 4003 10001
rect 4007 9997 4010 10001
rect 4014 9997 4029 10001
rect 3913 9996 4029 9997
rect 3913 9993 3926 9996
rect 3705 9992 3710 9993
rect 3614 9991 3710 9992
rect 3614 9987 3617 9991
rect 3621 9987 3624 9991
rect 3628 9987 3631 9991
rect 3635 9987 3638 9991
rect 3642 9987 3645 9991
rect 3649 9987 3652 9991
rect 3656 9987 3659 9991
rect 3663 9987 3666 9991
rect 3670 9987 3673 9991
rect 3677 9987 3680 9991
rect 3684 9987 3687 9991
rect 3691 9987 3694 9991
rect 3698 9987 3701 9991
rect 3705 9987 3710 9991
rect 3614 9986 3710 9987
rect 3614 9982 3617 9986
rect 3621 9982 3624 9986
rect 3628 9982 3631 9986
rect 3635 9982 3638 9986
rect 3642 9982 3645 9986
rect 3649 9982 3652 9986
rect 3656 9982 3659 9986
rect 3663 9982 3666 9986
rect 3670 9982 3673 9986
rect 3677 9982 3680 9986
rect 3684 9982 3687 9986
rect 3691 9982 3694 9986
rect 3698 9982 3701 9986
rect 3705 9982 3710 9986
rect 3614 9953 3710 9982
rect 3923 9992 3926 9993
rect 3930 9992 3933 9996
rect 3937 9992 3940 9996
rect 3944 9992 3947 9996
rect 3951 9992 3954 9996
rect 3958 9992 3961 9996
rect 3965 9992 3968 9996
rect 3972 9992 3975 9996
rect 3979 9992 3982 9996
rect 3986 9992 3989 9996
rect 3993 9992 3996 9996
rect 4000 9992 4003 9996
rect 4007 9992 4010 9996
rect 4014 9993 4029 9996
rect 4014 9992 4019 9993
rect 3923 9991 4019 9992
rect 3923 9987 3926 9991
rect 3930 9987 3933 9991
rect 3937 9987 3940 9991
rect 3944 9987 3947 9991
rect 3951 9987 3954 9991
rect 3958 9987 3961 9991
rect 3965 9987 3968 9991
rect 3972 9987 3975 9991
rect 3979 9987 3982 9991
rect 3986 9987 3989 9991
rect 3993 9987 3996 9991
rect 4000 9987 4003 9991
rect 4007 9987 4010 9991
rect 4014 9987 4019 9991
rect 3923 9986 4019 9987
rect 3923 9982 3926 9986
rect 3930 9982 3933 9986
rect 3937 9982 3940 9986
rect 3944 9982 3947 9986
rect 3951 9982 3954 9986
rect 3958 9982 3961 9986
rect 3965 9982 3968 9986
rect 3972 9982 3975 9986
rect 3979 9982 3982 9986
rect 3986 9982 3989 9986
rect 3993 9982 3996 9986
rect 4000 9982 4003 9986
rect 4007 9982 4010 9986
rect 4014 9982 4019 9986
rect 3923 9953 4019 9982
rect 1401 9949 1407 9953
rect 1411 9949 1417 9953
rect 1421 9949 1427 9953
rect 1431 9949 1437 9953
rect 1441 9949 1557 9953
rect 1561 9949 1567 9953
rect 1571 9949 1577 9953
rect 1581 9949 1587 9953
rect 1591 9949 1597 9953
rect 1397 9948 1601 9949
rect 1397 9944 1402 9948
rect 1406 9944 1412 9948
rect 1416 9944 1422 9948
rect 1426 9944 1432 9948
rect 1436 9944 1562 9948
rect 1566 9944 1572 9948
rect 1576 9944 1582 9948
rect 1586 9944 1592 9948
rect 1596 9944 1601 9948
rect 1397 9943 1601 9944
rect 1401 9939 1407 9943
rect 1411 9939 1417 9943
rect 1421 9939 1427 9943
rect 1431 9939 1437 9943
rect 1441 9939 1557 9943
rect 1561 9939 1567 9943
rect 1571 9939 1577 9943
rect 1581 9939 1587 9943
rect 1591 9939 1597 9943
rect 1397 9938 1601 9939
rect 1397 9934 1402 9938
rect 1406 9934 1412 9938
rect 1416 9934 1422 9938
rect 1426 9934 1432 9938
rect 1436 9934 1562 9938
rect 1566 9934 1572 9938
rect 1576 9934 1582 9938
rect 1586 9934 1592 9938
rect 1596 9934 1601 9938
rect 1397 9933 1601 9934
rect 1401 9929 1407 9933
rect 1411 9929 1417 9933
rect 1421 9929 1427 9933
rect 1431 9929 1437 9933
rect 1441 9929 1557 9933
rect 1561 9929 1567 9933
rect 1571 9929 1577 9933
rect 1581 9929 1587 9933
rect 1591 9929 1597 9933
rect 1397 9928 1601 9929
rect 1397 9924 1402 9928
rect 1406 9924 1412 9928
rect 1416 9924 1422 9928
rect 1426 9924 1432 9928
rect 1436 9924 1562 9928
rect 1566 9924 1572 9928
rect 1576 9924 1582 9928
rect 1586 9924 1592 9928
rect 1596 9924 1601 9928
rect 1397 9923 1601 9924
rect 1401 9919 1407 9923
rect 1411 9919 1417 9923
rect 1421 9919 1427 9923
rect 1431 9919 1437 9923
rect 1441 9919 1557 9923
rect 1561 9919 1567 9923
rect 1571 9919 1577 9923
rect 1581 9919 1587 9923
rect 1591 9919 1597 9923
rect 1397 9918 1601 9919
rect 1397 9914 1402 9918
rect 1406 9914 1412 9918
rect 1416 9914 1422 9918
rect 1426 9914 1432 9918
rect 1436 9914 1562 9918
rect 1566 9914 1572 9918
rect 1576 9914 1582 9918
rect 1586 9914 1592 9918
rect 1596 9914 1601 9918
rect 1397 9913 1601 9914
rect 1401 9909 1407 9913
rect 1411 9909 1417 9913
rect 1421 9909 1427 9913
rect 1431 9909 1437 9913
rect 1441 9909 1557 9913
rect 1561 9909 1567 9913
rect 1571 9909 1577 9913
rect 1581 9909 1587 9913
rect 1591 9909 1597 9913
rect 1397 9908 1601 9909
rect 1397 9904 1402 9908
rect 1406 9904 1412 9908
rect 1416 9904 1422 9908
rect 1426 9904 1432 9908
rect 1436 9904 1562 9908
rect 1566 9904 1572 9908
rect 1576 9904 1582 9908
rect 1586 9904 1592 9908
rect 1596 9904 1601 9908
rect 1397 9903 1601 9904
rect 1401 9899 1407 9903
rect 1411 9899 1417 9903
rect 1421 9899 1427 9903
rect 1431 9899 1437 9903
rect 1441 9899 1557 9903
rect 1561 9899 1567 9903
rect 1571 9899 1577 9903
rect 1581 9899 1587 9903
rect 1591 9899 1597 9903
rect 1397 9898 1601 9899
rect 1397 9894 1402 9898
rect 1406 9894 1412 9898
rect 1416 9894 1422 9898
rect 1426 9894 1432 9898
rect 1436 9894 1562 9898
rect 1566 9894 1572 9898
rect 1576 9894 1582 9898
rect 1586 9894 1592 9898
rect 1596 9894 1601 9898
rect 1397 9893 1601 9894
rect 1401 9889 1407 9893
rect 1411 9889 1417 9893
rect 1421 9889 1427 9893
rect 1431 9889 1437 9893
rect 1441 9889 1557 9893
rect 1561 9889 1567 9893
rect 1571 9889 1577 9893
rect 1581 9889 1587 9893
rect 1591 9889 1597 9893
rect 1397 9888 1601 9889
rect 1397 9884 1402 9888
rect 1406 9884 1412 9888
rect 1416 9884 1422 9888
rect 1426 9884 1432 9888
rect 1436 9884 1562 9888
rect 1566 9884 1572 9888
rect 1576 9884 1582 9888
rect 1586 9884 1592 9888
rect 1596 9884 1601 9888
rect 1397 9883 1601 9884
rect 1401 9879 1407 9883
rect 1411 9879 1417 9883
rect 1421 9879 1427 9883
rect 1431 9879 1437 9883
rect 1441 9879 1557 9883
rect 1561 9879 1567 9883
rect 1571 9879 1577 9883
rect 1581 9879 1587 9883
rect 1591 9879 1597 9883
rect 1397 9878 1601 9879
rect 1397 9874 1402 9878
rect 1406 9874 1412 9878
rect 1416 9874 1422 9878
rect 1426 9874 1432 9878
rect 1436 9874 1562 9878
rect 1566 9874 1572 9878
rect 1576 9874 1582 9878
rect 1586 9874 1592 9878
rect 1596 9874 1601 9878
rect 1397 9873 1601 9874
rect 1401 9869 1407 9873
rect 1411 9869 1417 9873
rect 1421 9869 1427 9873
rect 1431 9869 1437 9873
rect 1441 9869 1557 9873
rect 1561 9869 1567 9873
rect 1571 9869 1577 9873
rect 1581 9869 1587 9873
rect 1591 9869 1597 9873
rect 1397 9868 1601 9869
rect 1397 9864 1402 9868
rect 1406 9864 1412 9868
rect 1416 9864 1422 9868
rect 1426 9864 1432 9868
rect 1436 9864 1562 9868
rect 1566 9864 1572 9868
rect 1576 9864 1582 9868
rect 1586 9864 1592 9868
rect 1596 9864 1601 9868
rect 1710 9949 1716 9953
rect 1720 9949 1726 9953
rect 1730 9949 1736 9953
rect 1740 9949 1746 9953
rect 1750 9949 1866 9953
rect 1870 9949 1876 9953
rect 1880 9949 1886 9953
rect 1890 9949 1896 9953
rect 1900 9949 1906 9953
rect 1706 9948 1910 9949
rect 1706 9944 1711 9948
rect 1715 9944 1721 9948
rect 1725 9944 1731 9948
rect 1735 9944 1741 9948
rect 1745 9944 1871 9948
rect 1875 9944 1881 9948
rect 1885 9944 1891 9948
rect 1895 9944 1901 9948
rect 1905 9944 1910 9948
rect 1706 9943 1910 9944
rect 1710 9939 1716 9943
rect 1720 9939 1726 9943
rect 1730 9939 1736 9943
rect 1740 9939 1746 9943
rect 1750 9939 1866 9943
rect 1870 9939 1876 9943
rect 1880 9939 1886 9943
rect 1890 9939 1896 9943
rect 1900 9939 1906 9943
rect 1706 9938 1910 9939
rect 1706 9934 1711 9938
rect 1715 9934 1721 9938
rect 1725 9934 1731 9938
rect 1735 9934 1741 9938
rect 1745 9934 1871 9938
rect 1875 9934 1881 9938
rect 1885 9934 1891 9938
rect 1895 9934 1901 9938
rect 1905 9934 1910 9938
rect 1706 9933 1910 9934
rect 1710 9929 1716 9933
rect 1720 9929 1726 9933
rect 1730 9929 1736 9933
rect 1740 9929 1746 9933
rect 1750 9929 1866 9933
rect 1870 9929 1876 9933
rect 1880 9929 1886 9933
rect 1890 9929 1896 9933
rect 1900 9929 1906 9933
rect 1706 9928 1910 9929
rect 1706 9924 1711 9928
rect 1715 9924 1721 9928
rect 1725 9924 1731 9928
rect 1735 9924 1741 9928
rect 1745 9924 1871 9928
rect 1875 9924 1881 9928
rect 1885 9924 1891 9928
rect 1895 9924 1901 9928
rect 1905 9924 1910 9928
rect 1706 9923 1910 9924
rect 1710 9919 1716 9923
rect 1720 9919 1726 9923
rect 1730 9919 1736 9923
rect 1740 9919 1746 9923
rect 1750 9919 1866 9923
rect 1870 9919 1876 9923
rect 1880 9919 1886 9923
rect 1890 9919 1896 9923
rect 1900 9919 1906 9923
rect 1706 9918 1910 9919
rect 1706 9914 1711 9918
rect 1715 9914 1721 9918
rect 1725 9914 1731 9918
rect 1735 9914 1741 9918
rect 1745 9914 1871 9918
rect 1875 9914 1881 9918
rect 1885 9914 1891 9918
rect 1895 9914 1901 9918
rect 1905 9914 1910 9918
rect 1706 9913 1910 9914
rect 1710 9909 1716 9913
rect 1720 9909 1726 9913
rect 1730 9909 1736 9913
rect 1740 9909 1746 9913
rect 1750 9909 1866 9913
rect 1870 9909 1876 9913
rect 1880 9909 1886 9913
rect 1890 9909 1896 9913
rect 1900 9909 1906 9913
rect 1706 9908 1910 9909
rect 1706 9904 1711 9908
rect 1715 9904 1721 9908
rect 1725 9904 1731 9908
rect 1735 9904 1741 9908
rect 1745 9904 1871 9908
rect 1875 9904 1881 9908
rect 1885 9904 1891 9908
rect 1895 9904 1901 9908
rect 1905 9904 1910 9908
rect 1706 9903 1910 9904
rect 1710 9899 1716 9903
rect 1720 9899 1726 9903
rect 1730 9899 1736 9903
rect 1740 9899 1746 9903
rect 1750 9899 1866 9903
rect 1870 9899 1876 9903
rect 1880 9899 1886 9903
rect 1890 9899 1896 9903
rect 1900 9899 1906 9903
rect 1706 9898 1910 9899
rect 1706 9894 1711 9898
rect 1715 9894 1721 9898
rect 1725 9894 1731 9898
rect 1735 9894 1741 9898
rect 1745 9894 1871 9898
rect 1875 9894 1881 9898
rect 1885 9894 1891 9898
rect 1895 9894 1901 9898
rect 1905 9894 1910 9898
rect 1706 9893 1910 9894
rect 1710 9889 1716 9893
rect 1720 9889 1726 9893
rect 1730 9889 1736 9893
rect 1740 9889 1746 9893
rect 1750 9889 1866 9893
rect 1870 9889 1876 9893
rect 1880 9889 1886 9893
rect 1890 9889 1896 9893
rect 1900 9889 1906 9893
rect 1706 9888 1910 9889
rect 1706 9884 1711 9888
rect 1715 9884 1721 9888
rect 1725 9884 1731 9888
rect 1735 9884 1741 9888
rect 1745 9884 1871 9888
rect 1875 9884 1881 9888
rect 1885 9884 1891 9888
rect 1895 9884 1901 9888
rect 1905 9884 1910 9888
rect 1706 9883 1910 9884
rect 1710 9879 1716 9883
rect 1720 9879 1726 9883
rect 1730 9879 1736 9883
rect 1740 9879 1746 9883
rect 1750 9879 1866 9883
rect 1870 9879 1876 9883
rect 1880 9879 1886 9883
rect 1890 9879 1896 9883
rect 1900 9879 1906 9883
rect 1706 9878 1910 9879
rect 1706 9874 1711 9878
rect 1715 9874 1721 9878
rect 1725 9874 1731 9878
rect 1735 9874 1741 9878
rect 1745 9874 1871 9878
rect 1875 9874 1881 9878
rect 1885 9874 1891 9878
rect 1895 9874 1901 9878
rect 1905 9874 1910 9878
rect 1706 9873 1910 9874
rect 1710 9869 1716 9873
rect 1720 9869 1726 9873
rect 1730 9869 1736 9873
rect 1740 9869 1746 9873
rect 1750 9869 1866 9873
rect 1870 9869 1876 9873
rect 1880 9869 1886 9873
rect 1890 9869 1896 9873
rect 1900 9869 1906 9873
rect 1706 9868 1910 9869
rect 1706 9864 1711 9868
rect 1715 9864 1721 9868
rect 1725 9864 1731 9868
rect 1735 9864 1741 9868
rect 1745 9864 1871 9868
rect 1875 9864 1881 9868
rect 1885 9864 1891 9868
rect 1895 9864 1901 9868
rect 1905 9864 1910 9868
rect 2019 9949 2025 9953
rect 2029 9949 2035 9953
rect 2039 9949 2045 9953
rect 2049 9949 2055 9953
rect 2059 9949 2175 9953
rect 2179 9949 2185 9953
rect 2189 9949 2195 9953
rect 2199 9949 2205 9953
rect 2209 9949 2215 9953
rect 2015 9948 2219 9949
rect 2015 9944 2020 9948
rect 2024 9944 2030 9948
rect 2034 9944 2040 9948
rect 2044 9944 2050 9948
rect 2054 9944 2180 9948
rect 2184 9944 2190 9948
rect 2194 9944 2200 9948
rect 2204 9944 2210 9948
rect 2214 9944 2219 9948
rect 2015 9943 2219 9944
rect 2019 9939 2025 9943
rect 2029 9939 2035 9943
rect 2039 9939 2045 9943
rect 2049 9939 2055 9943
rect 2059 9939 2175 9943
rect 2179 9939 2185 9943
rect 2189 9939 2195 9943
rect 2199 9939 2205 9943
rect 2209 9939 2215 9943
rect 2015 9938 2219 9939
rect 2015 9934 2020 9938
rect 2024 9934 2030 9938
rect 2034 9934 2040 9938
rect 2044 9934 2050 9938
rect 2054 9934 2180 9938
rect 2184 9934 2190 9938
rect 2194 9934 2200 9938
rect 2204 9934 2210 9938
rect 2214 9934 2219 9938
rect 2015 9933 2219 9934
rect 2019 9929 2025 9933
rect 2029 9929 2035 9933
rect 2039 9929 2045 9933
rect 2049 9929 2055 9933
rect 2059 9929 2175 9933
rect 2179 9929 2185 9933
rect 2189 9929 2195 9933
rect 2199 9929 2205 9933
rect 2209 9929 2215 9933
rect 2015 9928 2219 9929
rect 2015 9924 2020 9928
rect 2024 9924 2030 9928
rect 2034 9924 2040 9928
rect 2044 9924 2050 9928
rect 2054 9924 2180 9928
rect 2184 9924 2190 9928
rect 2194 9924 2200 9928
rect 2204 9924 2210 9928
rect 2214 9924 2219 9928
rect 2015 9923 2219 9924
rect 2019 9919 2025 9923
rect 2029 9919 2035 9923
rect 2039 9919 2045 9923
rect 2049 9919 2055 9923
rect 2059 9919 2175 9923
rect 2179 9919 2185 9923
rect 2189 9919 2195 9923
rect 2199 9919 2205 9923
rect 2209 9919 2215 9923
rect 2015 9918 2219 9919
rect 2015 9914 2020 9918
rect 2024 9914 2030 9918
rect 2034 9914 2040 9918
rect 2044 9914 2050 9918
rect 2054 9914 2180 9918
rect 2184 9914 2190 9918
rect 2194 9914 2200 9918
rect 2204 9914 2210 9918
rect 2214 9914 2219 9918
rect 2015 9913 2219 9914
rect 2019 9909 2025 9913
rect 2029 9909 2035 9913
rect 2039 9909 2045 9913
rect 2049 9909 2055 9913
rect 2059 9909 2175 9913
rect 2179 9909 2185 9913
rect 2189 9909 2195 9913
rect 2199 9909 2205 9913
rect 2209 9909 2215 9913
rect 2015 9908 2219 9909
rect 2015 9904 2020 9908
rect 2024 9904 2030 9908
rect 2034 9904 2040 9908
rect 2044 9904 2050 9908
rect 2054 9904 2180 9908
rect 2184 9904 2190 9908
rect 2194 9904 2200 9908
rect 2204 9904 2210 9908
rect 2214 9904 2219 9908
rect 2015 9903 2219 9904
rect 2019 9899 2025 9903
rect 2029 9899 2035 9903
rect 2039 9899 2045 9903
rect 2049 9899 2055 9903
rect 2059 9899 2175 9903
rect 2179 9899 2185 9903
rect 2189 9899 2195 9903
rect 2199 9899 2205 9903
rect 2209 9899 2215 9903
rect 2015 9898 2219 9899
rect 2015 9894 2020 9898
rect 2024 9894 2030 9898
rect 2034 9894 2040 9898
rect 2044 9894 2050 9898
rect 2054 9894 2180 9898
rect 2184 9894 2190 9898
rect 2194 9894 2200 9898
rect 2204 9894 2210 9898
rect 2214 9894 2219 9898
rect 2015 9893 2219 9894
rect 2019 9889 2025 9893
rect 2029 9889 2035 9893
rect 2039 9889 2045 9893
rect 2049 9889 2055 9893
rect 2059 9889 2175 9893
rect 2179 9889 2185 9893
rect 2189 9889 2195 9893
rect 2199 9889 2205 9893
rect 2209 9889 2215 9893
rect 2015 9888 2219 9889
rect 2015 9884 2020 9888
rect 2024 9884 2030 9888
rect 2034 9884 2040 9888
rect 2044 9884 2050 9888
rect 2054 9884 2180 9888
rect 2184 9884 2190 9888
rect 2194 9884 2200 9888
rect 2204 9884 2210 9888
rect 2214 9884 2219 9888
rect 2015 9883 2219 9884
rect 2019 9879 2025 9883
rect 2029 9879 2035 9883
rect 2039 9879 2045 9883
rect 2049 9879 2055 9883
rect 2059 9879 2175 9883
rect 2179 9879 2185 9883
rect 2189 9879 2195 9883
rect 2199 9879 2205 9883
rect 2209 9879 2215 9883
rect 2015 9878 2219 9879
rect 2015 9874 2020 9878
rect 2024 9874 2030 9878
rect 2034 9874 2040 9878
rect 2044 9874 2050 9878
rect 2054 9874 2180 9878
rect 2184 9874 2190 9878
rect 2194 9874 2200 9878
rect 2204 9874 2210 9878
rect 2214 9874 2219 9878
rect 2015 9873 2219 9874
rect 2019 9869 2025 9873
rect 2029 9869 2035 9873
rect 2039 9869 2045 9873
rect 2049 9869 2055 9873
rect 2059 9869 2175 9873
rect 2179 9869 2185 9873
rect 2189 9869 2195 9873
rect 2199 9869 2205 9873
rect 2209 9869 2215 9873
rect 2015 9868 2219 9869
rect 2015 9864 2020 9868
rect 2024 9864 2030 9868
rect 2034 9864 2040 9868
rect 2044 9864 2050 9868
rect 2054 9864 2180 9868
rect 2184 9864 2190 9868
rect 2194 9864 2200 9868
rect 2204 9864 2210 9868
rect 2214 9864 2219 9868
rect 2328 9949 2334 9953
rect 2338 9949 2344 9953
rect 2348 9949 2354 9953
rect 2358 9949 2364 9953
rect 2368 9949 2484 9953
rect 2488 9949 2494 9953
rect 2498 9949 2504 9953
rect 2508 9949 2514 9953
rect 2518 9949 2524 9953
rect 2324 9948 2528 9949
rect 2324 9944 2329 9948
rect 2333 9944 2339 9948
rect 2343 9944 2349 9948
rect 2353 9944 2359 9948
rect 2363 9944 2489 9948
rect 2493 9944 2499 9948
rect 2503 9944 2509 9948
rect 2513 9944 2519 9948
rect 2523 9944 2528 9948
rect 2324 9943 2528 9944
rect 2328 9939 2334 9943
rect 2338 9939 2344 9943
rect 2348 9939 2354 9943
rect 2358 9939 2364 9943
rect 2368 9939 2484 9943
rect 2488 9939 2494 9943
rect 2498 9939 2504 9943
rect 2508 9939 2514 9943
rect 2518 9939 2524 9943
rect 2324 9938 2528 9939
rect 2324 9934 2329 9938
rect 2333 9934 2339 9938
rect 2343 9934 2349 9938
rect 2353 9934 2359 9938
rect 2363 9934 2489 9938
rect 2493 9934 2499 9938
rect 2503 9934 2509 9938
rect 2513 9934 2519 9938
rect 2523 9934 2528 9938
rect 2324 9933 2528 9934
rect 2328 9929 2334 9933
rect 2338 9929 2344 9933
rect 2348 9929 2354 9933
rect 2358 9929 2364 9933
rect 2368 9929 2484 9933
rect 2488 9929 2494 9933
rect 2498 9929 2504 9933
rect 2508 9929 2514 9933
rect 2518 9929 2524 9933
rect 2324 9928 2528 9929
rect 2324 9924 2329 9928
rect 2333 9924 2339 9928
rect 2343 9924 2349 9928
rect 2353 9924 2359 9928
rect 2363 9924 2489 9928
rect 2493 9924 2499 9928
rect 2503 9924 2509 9928
rect 2513 9924 2519 9928
rect 2523 9924 2528 9928
rect 2324 9923 2528 9924
rect 2328 9919 2334 9923
rect 2338 9919 2344 9923
rect 2348 9919 2354 9923
rect 2358 9919 2364 9923
rect 2368 9919 2484 9923
rect 2488 9919 2494 9923
rect 2498 9919 2504 9923
rect 2508 9919 2514 9923
rect 2518 9919 2524 9923
rect 2324 9918 2528 9919
rect 2324 9914 2329 9918
rect 2333 9914 2339 9918
rect 2343 9914 2349 9918
rect 2353 9914 2359 9918
rect 2363 9914 2489 9918
rect 2493 9914 2499 9918
rect 2503 9914 2509 9918
rect 2513 9914 2519 9918
rect 2523 9914 2528 9918
rect 2324 9913 2528 9914
rect 2328 9909 2334 9913
rect 2338 9909 2344 9913
rect 2348 9909 2354 9913
rect 2358 9909 2364 9913
rect 2368 9909 2484 9913
rect 2488 9909 2494 9913
rect 2498 9909 2504 9913
rect 2508 9909 2514 9913
rect 2518 9909 2524 9913
rect 2324 9908 2528 9909
rect 2324 9904 2329 9908
rect 2333 9904 2339 9908
rect 2343 9904 2349 9908
rect 2353 9904 2359 9908
rect 2363 9904 2489 9908
rect 2493 9904 2499 9908
rect 2503 9904 2509 9908
rect 2513 9904 2519 9908
rect 2523 9904 2528 9908
rect 2324 9903 2528 9904
rect 2328 9899 2334 9903
rect 2338 9899 2344 9903
rect 2348 9899 2354 9903
rect 2358 9899 2364 9903
rect 2368 9899 2484 9903
rect 2488 9899 2494 9903
rect 2498 9899 2504 9903
rect 2508 9899 2514 9903
rect 2518 9899 2524 9903
rect 2324 9898 2528 9899
rect 2324 9894 2329 9898
rect 2333 9894 2339 9898
rect 2343 9894 2349 9898
rect 2353 9894 2359 9898
rect 2363 9894 2489 9898
rect 2493 9894 2499 9898
rect 2503 9894 2509 9898
rect 2513 9894 2519 9898
rect 2523 9894 2528 9898
rect 2324 9893 2528 9894
rect 2328 9889 2334 9893
rect 2338 9889 2344 9893
rect 2348 9889 2354 9893
rect 2358 9889 2364 9893
rect 2368 9889 2484 9893
rect 2488 9889 2494 9893
rect 2498 9889 2504 9893
rect 2508 9889 2514 9893
rect 2518 9889 2524 9893
rect 2324 9888 2528 9889
rect 2324 9884 2329 9888
rect 2333 9884 2339 9888
rect 2343 9884 2349 9888
rect 2353 9884 2359 9888
rect 2363 9884 2489 9888
rect 2493 9884 2499 9888
rect 2503 9884 2509 9888
rect 2513 9884 2519 9888
rect 2523 9884 2528 9888
rect 2324 9883 2528 9884
rect 2328 9879 2334 9883
rect 2338 9879 2344 9883
rect 2348 9879 2354 9883
rect 2358 9879 2364 9883
rect 2368 9879 2484 9883
rect 2488 9879 2494 9883
rect 2498 9879 2504 9883
rect 2508 9879 2514 9883
rect 2518 9879 2524 9883
rect 2324 9878 2528 9879
rect 2324 9874 2329 9878
rect 2333 9874 2339 9878
rect 2343 9874 2349 9878
rect 2353 9874 2359 9878
rect 2363 9874 2489 9878
rect 2493 9874 2499 9878
rect 2503 9874 2509 9878
rect 2513 9874 2519 9878
rect 2523 9874 2528 9878
rect 2324 9873 2528 9874
rect 2328 9869 2334 9873
rect 2338 9869 2344 9873
rect 2348 9869 2354 9873
rect 2358 9869 2364 9873
rect 2368 9869 2484 9873
rect 2488 9869 2494 9873
rect 2498 9869 2504 9873
rect 2508 9869 2514 9873
rect 2518 9869 2524 9873
rect 2324 9868 2528 9869
rect 2324 9864 2329 9868
rect 2333 9864 2339 9868
rect 2343 9864 2349 9868
rect 2353 9864 2359 9868
rect 2363 9864 2489 9868
rect 2493 9864 2499 9868
rect 2503 9864 2509 9868
rect 2513 9864 2519 9868
rect 2523 9864 2528 9868
rect 2637 9949 2643 9953
rect 2647 9949 2653 9953
rect 2657 9949 2663 9953
rect 2667 9949 2673 9953
rect 2677 9949 2793 9953
rect 2797 9949 2803 9953
rect 2807 9949 2813 9953
rect 2817 9949 2823 9953
rect 2827 9949 2833 9953
rect 2633 9948 2837 9949
rect 2633 9944 2638 9948
rect 2642 9944 2648 9948
rect 2652 9944 2658 9948
rect 2662 9944 2668 9948
rect 2672 9944 2798 9948
rect 2802 9944 2808 9948
rect 2812 9944 2818 9948
rect 2822 9944 2828 9948
rect 2832 9944 2837 9948
rect 2633 9943 2837 9944
rect 2637 9939 2643 9943
rect 2647 9939 2653 9943
rect 2657 9939 2663 9943
rect 2667 9939 2673 9943
rect 2677 9939 2793 9943
rect 2797 9939 2803 9943
rect 2807 9939 2813 9943
rect 2817 9939 2823 9943
rect 2827 9939 2833 9943
rect 2633 9938 2837 9939
rect 2633 9934 2638 9938
rect 2642 9934 2648 9938
rect 2652 9934 2658 9938
rect 2662 9934 2668 9938
rect 2672 9934 2798 9938
rect 2802 9934 2808 9938
rect 2812 9934 2818 9938
rect 2822 9934 2828 9938
rect 2832 9934 2837 9938
rect 2633 9933 2837 9934
rect 2637 9929 2643 9933
rect 2647 9929 2653 9933
rect 2657 9929 2663 9933
rect 2667 9929 2673 9933
rect 2677 9929 2793 9933
rect 2797 9929 2803 9933
rect 2807 9929 2813 9933
rect 2817 9929 2823 9933
rect 2827 9929 2833 9933
rect 2633 9928 2837 9929
rect 2633 9924 2638 9928
rect 2642 9924 2648 9928
rect 2652 9924 2658 9928
rect 2662 9924 2668 9928
rect 2672 9924 2798 9928
rect 2802 9924 2808 9928
rect 2812 9924 2818 9928
rect 2822 9924 2828 9928
rect 2832 9924 2837 9928
rect 2633 9923 2837 9924
rect 2637 9919 2643 9923
rect 2647 9919 2653 9923
rect 2657 9919 2663 9923
rect 2667 9919 2673 9923
rect 2677 9919 2793 9923
rect 2797 9919 2803 9923
rect 2807 9919 2813 9923
rect 2817 9919 2823 9923
rect 2827 9919 2833 9923
rect 2633 9918 2837 9919
rect 2633 9914 2638 9918
rect 2642 9914 2648 9918
rect 2652 9914 2658 9918
rect 2662 9914 2668 9918
rect 2672 9914 2798 9918
rect 2802 9914 2808 9918
rect 2812 9914 2818 9918
rect 2822 9914 2828 9918
rect 2832 9914 2837 9918
rect 2633 9913 2837 9914
rect 2637 9909 2643 9913
rect 2647 9909 2653 9913
rect 2657 9909 2663 9913
rect 2667 9909 2673 9913
rect 2677 9909 2793 9913
rect 2797 9909 2803 9913
rect 2807 9909 2813 9913
rect 2817 9909 2823 9913
rect 2827 9909 2833 9913
rect 2633 9908 2837 9909
rect 2633 9904 2638 9908
rect 2642 9904 2648 9908
rect 2652 9904 2658 9908
rect 2662 9904 2668 9908
rect 2672 9904 2798 9908
rect 2802 9904 2808 9908
rect 2812 9904 2818 9908
rect 2822 9904 2828 9908
rect 2832 9904 2837 9908
rect 2633 9903 2837 9904
rect 2637 9899 2643 9903
rect 2647 9899 2653 9903
rect 2657 9899 2663 9903
rect 2667 9899 2673 9903
rect 2677 9899 2793 9903
rect 2797 9899 2803 9903
rect 2807 9899 2813 9903
rect 2817 9899 2823 9903
rect 2827 9899 2833 9903
rect 2633 9898 2837 9899
rect 2633 9894 2638 9898
rect 2642 9894 2648 9898
rect 2652 9894 2658 9898
rect 2662 9894 2668 9898
rect 2672 9894 2798 9898
rect 2802 9894 2808 9898
rect 2812 9894 2818 9898
rect 2822 9894 2828 9898
rect 2832 9894 2837 9898
rect 2633 9893 2837 9894
rect 2637 9889 2643 9893
rect 2647 9889 2653 9893
rect 2657 9889 2663 9893
rect 2667 9889 2673 9893
rect 2677 9889 2793 9893
rect 2797 9889 2803 9893
rect 2807 9889 2813 9893
rect 2817 9889 2823 9893
rect 2827 9889 2833 9893
rect 2633 9888 2837 9889
rect 2633 9884 2638 9888
rect 2642 9884 2648 9888
rect 2652 9884 2658 9888
rect 2662 9884 2668 9888
rect 2672 9884 2798 9888
rect 2802 9884 2808 9888
rect 2812 9884 2818 9888
rect 2822 9884 2828 9888
rect 2832 9884 2837 9888
rect 2633 9883 2837 9884
rect 2637 9879 2643 9883
rect 2647 9879 2653 9883
rect 2657 9879 2663 9883
rect 2667 9879 2673 9883
rect 2677 9879 2793 9883
rect 2797 9879 2803 9883
rect 2807 9879 2813 9883
rect 2817 9879 2823 9883
rect 2827 9879 2833 9883
rect 2633 9878 2837 9879
rect 2633 9874 2638 9878
rect 2642 9874 2648 9878
rect 2652 9874 2658 9878
rect 2662 9874 2668 9878
rect 2672 9874 2798 9878
rect 2802 9874 2808 9878
rect 2812 9874 2818 9878
rect 2822 9874 2828 9878
rect 2832 9874 2837 9878
rect 2633 9873 2837 9874
rect 2637 9869 2643 9873
rect 2647 9869 2653 9873
rect 2657 9869 2663 9873
rect 2667 9869 2673 9873
rect 2677 9869 2793 9873
rect 2797 9869 2803 9873
rect 2807 9869 2813 9873
rect 2817 9869 2823 9873
rect 2827 9869 2833 9873
rect 2633 9868 2837 9869
rect 2633 9864 2638 9868
rect 2642 9864 2648 9868
rect 2652 9864 2658 9868
rect 2662 9864 2668 9868
rect 2672 9864 2798 9868
rect 2802 9864 2808 9868
rect 2812 9864 2818 9868
rect 2822 9864 2828 9868
rect 2832 9864 2837 9868
rect 2946 9949 2952 9953
rect 2956 9949 2962 9953
rect 2966 9949 2972 9953
rect 2976 9949 2982 9953
rect 2986 9949 3102 9953
rect 3106 9949 3112 9953
rect 3116 9949 3122 9953
rect 3126 9949 3132 9953
rect 3136 9949 3142 9953
rect 2942 9948 3146 9949
rect 2942 9944 2947 9948
rect 2951 9944 2957 9948
rect 2961 9944 2967 9948
rect 2971 9944 2977 9948
rect 2981 9944 3107 9948
rect 3111 9944 3117 9948
rect 3121 9944 3127 9948
rect 3131 9944 3137 9948
rect 3141 9944 3146 9948
rect 2942 9943 3146 9944
rect 2946 9939 2952 9943
rect 2956 9939 2962 9943
rect 2966 9939 2972 9943
rect 2976 9939 2982 9943
rect 2986 9939 3102 9943
rect 3106 9939 3112 9943
rect 3116 9939 3122 9943
rect 3126 9939 3132 9943
rect 3136 9939 3142 9943
rect 2942 9938 3146 9939
rect 2942 9934 2947 9938
rect 2951 9934 2957 9938
rect 2961 9934 2967 9938
rect 2971 9934 2977 9938
rect 2981 9934 3107 9938
rect 3111 9934 3117 9938
rect 3121 9934 3127 9938
rect 3131 9934 3137 9938
rect 3141 9934 3146 9938
rect 2942 9933 3146 9934
rect 2946 9929 2952 9933
rect 2956 9929 2962 9933
rect 2966 9929 2972 9933
rect 2976 9929 2982 9933
rect 2986 9929 3102 9933
rect 3106 9929 3112 9933
rect 3116 9929 3122 9933
rect 3126 9929 3132 9933
rect 3136 9929 3142 9933
rect 2942 9928 3146 9929
rect 2942 9924 2947 9928
rect 2951 9924 2957 9928
rect 2961 9924 2967 9928
rect 2971 9924 2977 9928
rect 2981 9924 3107 9928
rect 3111 9924 3117 9928
rect 3121 9924 3127 9928
rect 3131 9924 3137 9928
rect 3141 9924 3146 9928
rect 2942 9923 3146 9924
rect 2946 9919 2952 9923
rect 2956 9919 2962 9923
rect 2966 9919 2972 9923
rect 2976 9919 2982 9923
rect 2986 9919 3102 9923
rect 3106 9919 3112 9923
rect 3116 9919 3122 9923
rect 3126 9919 3132 9923
rect 3136 9919 3142 9923
rect 2942 9918 3146 9919
rect 2942 9914 2947 9918
rect 2951 9914 2957 9918
rect 2961 9914 2967 9918
rect 2971 9914 2977 9918
rect 2981 9914 3107 9918
rect 3111 9914 3117 9918
rect 3121 9914 3127 9918
rect 3131 9914 3137 9918
rect 3141 9914 3146 9918
rect 2942 9913 3146 9914
rect 2946 9909 2952 9913
rect 2956 9909 2962 9913
rect 2966 9909 2972 9913
rect 2976 9909 2982 9913
rect 2986 9909 3102 9913
rect 3106 9909 3112 9913
rect 3116 9909 3122 9913
rect 3126 9909 3132 9913
rect 3136 9909 3142 9913
rect 2942 9908 3146 9909
rect 2942 9904 2947 9908
rect 2951 9904 2957 9908
rect 2961 9904 2967 9908
rect 2971 9904 2977 9908
rect 2981 9904 3107 9908
rect 3111 9904 3117 9908
rect 3121 9904 3127 9908
rect 3131 9904 3137 9908
rect 3141 9904 3146 9908
rect 2942 9903 3146 9904
rect 2946 9899 2952 9903
rect 2956 9899 2962 9903
rect 2966 9899 2972 9903
rect 2976 9899 2982 9903
rect 2986 9899 3102 9903
rect 3106 9899 3112 9903
rect 3116 9899 3122 9903
rect 3126 9899 3132 9903
rect 3136 9899 3142 9903
rect 2942 9898 3146 9899
rect 2942 9894 2947 9898
rect 2951 9894 2957 9898
rect 2961 9894 2967 9898
rect 2971 9894 2977 9898
rect 2981 9894 3107 9898
rect 3111 9894 3117 9898
rect 3121 9894 3127 9898
rect 3131 9894 3137 9898
rect 3141 9894 3146 9898
rect 2942 9893 3146 9894
rect 2946 9889 2952 9893
rect 2956 9889 2962 9893
rect 2966 9889 2972 9893
rect 2976 9889 2982 9893
rect 2986 9889 3102 9893
rect 3106 9889 3112 9893
rect 3116 9889 3122 9893
rect 3126 9889 3132 9893
rect 3136 9889 3142 9893
rect 2942 9888 3146 9889
rect 2942 9884 2947 9888
rect 2951 9884 2957 9888
rect 2961 9884 2967 9888
rect 2971 9884 2977 9888
rect 2981 9884 3107 9888
rect 3111 9884 3117 9888
rect 3121 9884 3127 9888
rect 3131 9884 3137 9888
rect 3141 9884 3146 9888
rect 2942 9883 3146 9884
rect 2946 9879 2952 9883
rect 2956 9879 2962 9883
rect 2966 9879 2972 9883
rect 2976 9879 2982 9883
rect 2986 9879 3102 9883
rect 3106 9879 3112 9883
rect 3116 9879 3122 9883
rect 3126 9879 3132 9883
rect 3136 9879 3142 9883
rect 2942 9878 3146 9879
rect 2942 9874 2947 9878
rect 2951 9874 2957 9878
rect 2961 9874 2967 9878
rect 2971 9874 2977 9878
rect 2981 9874 3107 9878
rect 3111 9874 3117 9878
rect 3121 9874 3127 9878
rect 3131 9874 3137 9878
rect 3141 9874 3146 9878
rect 2942 9873 3146 9874
rect 2946 9869 2952 9873
rect 2956 9869 2962 9873
rect 2966 9869 2972 9873
rect 2976 9869 2982 9873
rect 2986 9869 3102 9873
rect 3106 9869 3112 9873
rect 3116 9869 3122 9873
rect 3126 9869 3132 9873
rect 3136 9869 3142 9873
rect 2942 9868 3146 9869
rect 2942 9864 2947 9868
rect 2951 9864 2957 9868
rect 2961 9864 2967 9868
rect 2971 9864 2977 9868
rect 2981 9864 3107 9868
rect 3111 9864 3117 9868
rect 3121 9864 3127 9868
rect 3131 9864 3137 9868
rect 3141 9864 3146 9868
rect 3255 9949 3261 9953
rect 3265 9949 3271 9953
rect 3275 9949 3281 9953
rect 3285 9949 3291 9953
rect 3295 9949 3411 9953
rect 3415 9949 3421 9953
rect 3425 9949 3431 9953
rect 3435 9949 3441 9953
rect 3445 9949 3451 9953
rect 3251 9948 3455 9949
rect 3251 9944 3256 9948
rect 3260 9944 3266 9948
rect 3270 9944 3276 9948
rect 3280 9944 3286 9948
rect 3290 9944 3416 9948
rect 3420 9944 3426 9948
rect 3430 9944 3436 9948
rect 3440 9944 3446 9948
rect 3450 9944 3455 9948
rect 3251 9943 3455 9944
rect 3255 9939 3261 9943
rect 3265 9939 3271 9943
rect 3275 9939 3281 9943
rect 3285 9939 3291 9943
rect 3295 9939 3411 9943
rect 3415 9939 3421 9943
rect 3425 9939 3431 9943
rect 3435 9939 3441 9943
rect 3445 9939 3451 9943
rect 3251 9938 3455 9939
rect 3251 9934 3256 9938
rect 3260 9934 3266 9938
rect 3270 9934 3276 9938
rect 3280 9934 3286 9938
rect 3290 9934 3416 9938
rect 3420 9934 3426 9938
rect 3430 9934 3436 9938
rect 3440 9934 3446 9938
rect 3450 9934 3455 9938
rect 3251 9933 3455 9934
rect 3255 9929 3261 9933
rect 3265 9929 3271 9933
rect 3275 9929 3281 9933
rect 3285 9929 3291 9933
rect 3295 9929 3411 9933
rect 3415 9929 3421 9933
rect 3425 9929 3431 9933
rect 3435 9929 3441 9933
rect 3445 9929 3451 9933
rect 3251 9928 3455 9929
rect 3251 9924 3256 9928
rect 3260 9924 3266 9928
rect 3270 9924 3276 9928
rect 3280 9924 3286 9928
rect 3290 9924 3416 9928
rect 3420 9924 3426 9928
rect 3430 9924 3436 9928
rect 3440 9924 3446 9928
rect 3450 9924 3455 9928
rect 3251 9923 3455 9924
rect 3255 9919 3261 9923
rect 3265 9919 3271 9923
rect 3275 9919 3281 9923
rect 3285 9919 3291 9923
rect 3295 9919 3411 9923
rect 3415 9919 3421 9923
rect 3425 9919 3431 9923
rect 3435 9919 3441 9923
rect 3445 9919 3451 9923
rect 3251 9918 3455 9919
rect 3251 9914 3256 9918
rect 3260 9914 3266 9918
rect 3270 9914 3276 9918
rect 3280 9914 3286 9918
rect 3290 9914 3416 9918
rect 3420 9914 3426 9918
rect 3430 9914 3436 9918
rect 3440 9914 3446 9918
rect 3450 9914 3455 9918
rect 3251 9913 3455 9914
rect 3255 9909 3261 9913
rect 3265 9909 3271 9913
rect 3275 9909 3281 9913
rect 3285 9909 3291 9913
rect 3295 9909 3411 9913
rect 3415 9909 3421 9913
rect 3425 9909 3431 9913
rect 3435 9909 3441 9913
rect 3445 9909 3451 9913
rect 3251 9908 3455 9909
rect 3251 9904 3256 9908
rect 3260 9904 3266 9908
rect 3270 9904 3276 9908
rect 3280 9904 3286 9908
rect 3290 9904 3416 9908
rect 3420 9904 3426 9908
rect 3430 9904 3436 9908
rect 3440 9904 3446 9908
rect 3450 9904 3455 9908
rect 3251 9903 3455 9904
rect 3255 9899 3261 9903
rect 3265 9899 3271 9903
rect 3275 9899 3281 9903
rect 3285 9899 3291 9903
rect 3295 9899 3411 9903
rect 3415 9899 3421 9903
rect 3425 9899 3431 9903
rect 3435 9899 3441 9903
rect 3445 9899 3451 9903
rect 3251 9898 3455 9899
rect 3251 9894 3256 9898
rect 3260 9894 3266 9898
rect 3270 9894 3276 9898
rect 3280 9894 3286 9898
rect 3290 9894 3416 9898
rect 3420 9894 3426 9898
rect 3430 9894 3436 9898
rect 3440 9894 3446 9898
rect 3450 9894 3455 9898
rect 3251 9893 3455 9894
rect 3255 9889 3261 9893
rect 3265 9889 3271 9893
rect 3275 9889 3281 9893
rect 3285 9889 3291 9893
rect 3295 9889 3411 9893
rect 3415 9889 3421 9893
rect 3425 9889 3431 9893
rect 3435 9889 3441 9893
rect 3445 9889 3451 9893
rect 3251 9888 3455 9889
rect 3251 9884 3256 9888
rect 3260 9884 3266 9888
rect 3270 9884 3276 9888
rect 3280 9884 3286 9888
rect 3290 9884 3416 9888
rect 3420 9884 3426 9888
rect 3430 9884 3436 9888
rect 3440 9884 3446 9888
rect 3450 9884 3455 9888
rect 3251 9883 3455 9884
rect 3255 9879 3261 9883
rect 3265 9879 3271 9883
rect 3275 9879 3281 9883
rect 3285 9879 3291 9883
rect 3295 9879 3411 9883
rect 3415 9879 3421 9883
rect 3425 9879 3431 9883
rect 3435 9879 3441 9883
rect 3445 9879 3451 9883
rect 3251 9878 3455 9879
rect 3251 9874 3256 9878
rect 3260 9874 3266 9878
rect 3270 9874 3276 9878
rect 3280 9874 3286 9878
rect 3290 9874 3416 9878
rect 3420 9874 3426 9878
rect 3430 9874 3436 9878
rect 3440 9874 3446 9878
rect 3450 9874 3455 9878
rect 3251 9873 3455 9874
rect 3255 9869 3261 9873
rect 3265 9869 3271 9873
rect 3275 9869 3281 9873
rect 3285 9869 3291 9873
rect 3295 9869 3411 9873
rect 3415 9869 3421 9873
rect 3425 9869 3431 9873
rect 3435 9869 3441 9873
rect 3445 9869 3451 9873
rect 3251 9868 3455 9869
rect 3251 9864 3256 9868
rect 3260 9864 3266 9868
rect 3270 9864 3276 9868
rect 3280 9864 3286 9868
rect 3290 9864 3416 9868
rect 3420 9864 3426 9868
rect 3430 9864 3436 9868
rect 3440 9864 3446 9868
rect 3450 9864 3455 9868
rect 3564 9949 3570 9953
rect 3574 9949 3580 9953
rect 3584 9949 3590 9953
rect 3594 9949 3600 9953
rect 3604 9949 3720 9953
rect 3724 9949 3730 9953
rect 3734 9949 3740 9953
rect 3744 9949 3750 9953
rect 3754 9949 3760 9953
rect 3560 9948 3764 9949
rect 3560 9944 3565 9948
rect 3569 9944 3575 9948
rect 3579 9944 3585 9948
rect 3589 9944 3595 9948
rect 3599 9944 3725 9948
rect 3729 9944 3735 9948
rect 3739 9944 3745 9948
rect 3749 9944 3755 9948
rect 3759 9944 3764 9948
rect 3560 9943 3764 9944
rect 3564 9939 3570 9943
rect 3574 9939 3580 9943
rect 3584 9939 3590 9943
rect 3594 9939 3600 9943
rect 3604 9939 3720 9943
rect 3724 9939 3730 9943
rect 3734 9939 3740 9943
rect 3744 9939 3750 9943
rect 3754 9939 3760 9943
rect 3560 9938 3764 9939
rect 3560 9934 3565 9938
rect 3569 9934 3575 9938
rect 3579 9934 3585 9938
rect 3589 9934 3595 9938
rect 3599 9934 3725 9938
rect 3729 9934 3735 9938
rect 3739 9934 3745 9938
rect 3749 9934 3755 9938
rect 3759 9934 3764 9938
rect 3560 9933 3764 9934
rect 3564 9929 3570 9933
rect 3574 9929 3580 9933
rect 3584 9929 3590 9933
rect 3594 9929 3600 9933
rect 3604 9929 3720 9933
rect 3724 9929 3730 9933
rect 3734 9929 3740 9933
rect 3744 9929 3750 9933
rect 3754 9929 3760 9933
rect 3560 9928 3764 9929
rect 3560 9924 3565 9928
rect 3569 9924 3575 9928
rect 3579 9924 3585 9928
rect 3589 9924 3595 9928
rect 3599 9924 3725 9928
rect 3729 9924 3735 9928
rect 3739 9924 3745 9928
rect 3749 9924 3755 9928
rect 3759 9924 3764 9928
rect 3560 9923 3764 9924
rect 3564 9919 3570 9923
rect 3574 9919 3580 9923
rect 3584 9919 3590 9923
rect 3594 9919 3600 9923
rect 3604 9919 3720 9923
rect 3724 9919 3730 9923
rect 3734 9919 3740 9923
rect 3744 9919 3750 9923
rect 3754 9919 3760 9923
rect 3560 9918 3764 9919
rect 3560 9914 3565 9918
rect 3569 9914 3575 9918
rect 3579 9914 3585 9918
rect 3589 9914 3595 9918
rect 3599 9914 3725 9918
rect 3729 9914 3735 9918
rect 3739 9914 3745 9918
rect 3749 9914 3755 9918
rect 3759 9914 3764 9918
rect 3560 9913 3764 9914
rect 3564 9909 3570 9913
rect 3574 9909 3580 9913
rect 3584 9909 3590 9913
rect 3594 9909 3600 9913
rect 3604 9909 3720 9913
rect 3724 9909 3730 9913
rect 3734 9909 3740 9913
rect 3744 9909 3750 9913
rect 3754 9909 3760 9913
rect 3560 9908 3764 9909
rect 3560 9904 3565 9908
rect 3569 9904 3575 9908
rect 3579 9904 3585 9908
rect 3589 9904 3595 9908
rect 3599 9904 3725 9908
rect 3729 9904 3735 9908
rect 3739 9904 3745 9908
rect 3749 9904 3755 9908
rect 3759 9904 3764 9908
rect 3560 9903 3764 9904
rect 3564 9899 3570 9903
rect 3574 9899 3580 9903
rect 3584 9899 3590 9903
rect 3594 9899 3600 9903
rect 3604 9899 3720 9903
rect 3724 9899 3730 9903
rect 3734 9899 3740 9903
rect 3744 9899 3750 9903
rect 3754 9899 3760 9903
rect 3560 9898 3764 9899
rect 3560 9894 3565 9898
rect 3569 9894 3575 9898
rect 3579 9894 3585 9898
rect 3589 9894 3595 9898
rect 3599 9894 3725 9898
rect 3729 9894 3735 9898
rect 3739 9894 3745 9898
rect 3749 9894 3755 9898
rect 3759 9894 3764 9898
rect 3560 9893 3764 9894
rect 3564 9889 3570 9893
rect 3574 9889 3580 9893
rect 3584 9889 3590 9893
rect 3594 9889 3600 9893
rect 3604 9889 3720 9893
rect 3724 9889 3730 9893
rect 3734 9889 3740 9893
rect 3744 9889 3750 9893
rect 3754 9889 3760 9893
rect 3560 9888 3764 9889
rect 3560 9884 3565 9888
rect 3569 9884 3575 9888
rect 3579 9884 3585 9888
rect 3589 9884 3595 9888
rect 3599 9884 3725 9888
rect 3729 9884 3735 9888
rect 3739 9884 3745 9888
rect 3749 9884 3755 9888
rect 3759 9884 3764 9888
rect 3560 9883 3764 9884
rect 3564 9879 3570 9883
rect 3574 9879 3580 9883
rect 3584 9879 3590 9883
rect 3594 9879 3600 9883
rect 3604 9879 3720 9883
rect 3724 9879 3730 9883
rect 3734 9879 3740 9883
rect 3744 9879 3750 9883
rect 3754 9879 3760 9883
rect 3560 9878 3764 9879
rect 3560 9874 3565 9878
rect 3569 9874 3575 9878
rect 3579 9874 3585 9878
rect 3589 9874 3595 9878
rect 3599 9874 3725 9878
rect 3729 9874 3735 9878
rect 3739 9874 3745 9878
rect 3749 9874 3755 9878
rect 3759 9874 3764 9878
rect 3560 9873 3764 9874
rect 3564 9869 3570 9873
rect 3574 9869 3580 9873
rect 3584 9869 3590 9873
rect 3594 9869 3600 9873
rect 3604 9869 3720 9873
rect 3724 9869 3730 9873
rect 3734 9869 3740 9873
rect 3744 9869 3750 9873
rect 3754 9869 3760 9873
rect 3560 9868 3764 9869
rect 3560 9864 3565 9868
rect 3569 9864 3575 9868
rect 3579 9864 3585 9868
rect 3589 9864 3595 9868
rect 3599 9864 3725 9868
rect 3729 9864 3735 9868
rect 3739 9864 3745 9868
rect 3749 9864 3755 9868
rect 3759 9864 3764 9868
rect 3873 9949 3879 9953
rect 3883 9949 3889 9953
rect 3893 9949 3899 9953
rect 3903 9949 3909 9953
rect 3913 9949 4029 9953
rect 4033 9949 4039 9953
rect 4043 9949 4049 9953
rect 4053 9949 4059 9953
rect 4063 9949 4069 9953
rect 3869 9948 4073 9949
rect 3869 9944 3874 9948
rect 3878 9944 3884 9948
rect 3888 9944 3894 9948
rect 3898 9944 3904 9948
rect 3908 9944 4034 9948
rect 4038 9944 4044 9948
rect 4048 9944 4054 9948
rect 4058 9944 4064 9948
rect 4068 9944 4073 9948
rect 3869 9943 4073 9944
rect 3873 9939 3879 9943
rect 3883 9939 3889 9943
rect 3893 9939 3899 9943
rect 3903 9939 3909 9943
rect 3913 9939 4029 9943
rect 4033 9939 4039 9943
rect 4043 9939 4049 9943
rect 4053 9939 4059 9943
rect 4063 9939 4069 9943
rect 3869 9938 4073 9939
rect 3869 9934 3874 9938
rect 3878 9934 3884 9938
rect 3888 9934 3894 9938
rect 3898 9934 3904 9938
rect 3908 9934 4034 9938
rect 4038 9934 4044 9938
rect 4048 9934 4054 9938
rect 4058 9934 4064 9938
rect 4068 9934 4073 9938
rect 3869 9933 4073 9934
rect 3873 9929 3879 9933
rect 3883 9929 3889 9933
rect 3893 9929 3899 9933
rect 3903 9929 3909 9933
rect 3913 9929 4029 9933
rect 4033 9929 4039 9933
rect 4043 9929 4049 9933
rect 4053 9929 4059 9933
rect 4063 9929 4069 9933
rect 3869 9928 4073 9929
rect 3869 9924 3874 9928
rect 3878 9924 3884 9928
rect 3888 9924 3894 9928
rect 3898 9924 3904 9928
rect 3908 9924 4034 9928
rect 4038 9924 4044 9928
rect 4048 9924 4054 9928
rect 4058 9924 4064 9928
rect 4068 9924 4073 9928
rect 3869 9923 4073 9924
rect 3873 9919 3879 9923
rect 3883 9919 3889 9923
rect 3893 9919 3899 9923
rect 3903 9919 3909 9923
rect 3913 9919 4029 9923
rect 4033 9919 4039 9923
rect 4043 9919 4049 9923
rect 4053 9919 4059 9923
rect 4063 9919 4069 9923
rect 3869 9918 4073 9919
rect 3869 9914 3874 9918
rect 3878 9914 3884 9918
rect 3888 9914 3894 9918
rect 3898 9914 3904 9918
rect 3908 9914 4034 9918
rect 4038 9914 4044 9918
rect 4048 9914 4054 9918
rect 4058 9914 4064 9918
rect 4068 9914 4073 9918
rect 3869 9913 4073 9914
rect 3873 9909 3879 9913
rect 3883 9909 3889 9913
rect 3893 9909 3899 9913
rect 3903 9909 3909 9913
rect 3913 9909 4029 9913
rect 4033 9909 4039 9913
rect 4043 9909 4049 9913
rect 4053 9909 4059 9913
rect 4063 9909 4069 9913
rect 3869 9908 4073 9909
rect 3869 9904 3874 9908
rect 3878 9904 3884 9908
rect 3888 9904 3894 9908
rect 3898 9904 3904 9908
rect 3908 9904 4034 9908
rect 4038 9904 4044 9908
rect 4048 9904 4054 9908
rect 4058 9904 4064 9908
rect 4068 9904 4073 9908
rect 3869 9903 4073 9904
rect 3873 9899 3879 9903
rect 3883 9899 3889 9903
rect 3893 9899 3899 9903
rect 3903 9899 3909 9903
rect 3913 9899 4029 9903
rect 4033 9899 4039 9903
rect 4043 9899 4049 9903
rect 4053 9899 4059 9903
rect 4063 9899 4069 9903
rect 3869 9898 4073 9899
rect 3869 9894 3874 9898
rect 3878 9894 3884 9898
rect 3888 9894 3894 9898
rect 3898 9894 3904 9898
rect 3908 9894 4034 9898
rect 4038 9894 4044 9898
rect 4048 9894 4054 9898
rect 4058 9894 4064 9898
rect 4068 9894 4073 9898
rect 3869 9893 4073 9894
rect 3873 9889 3879 9893
rect 3883 9889 3889 9893
rect 3893 9889 3899 9893
rect 3903 9889 3909 9893
rect 3913 9889 4029 9893
rect 4033 9889 4039 9893
rect 4043 9889 4049 9893
rect 4053 9889 4059 9893
rect 4063 9889 4069 9893
rect 3869 9888 4073 9889
rect 3869 9884 3874 9888
rect 3878 9884 3884 9888
rect 3888 9884 3894 9888
rect 3898 9884 3904 9888
rect 3908 9884 4034 9888
rect 4038 9884 4044 9888
rect 4048 9884 4054 9888
rect 4058 9884 4064 9888
rect 4068 9884 4073 9888
rect 3869 9883 4073 9884
rect 3873 9879 3879 9883
rect 3883 9879 3889 9883
rect 3893 9879 3899 9883
rect 3903 9879 3909 9883
rect 3913 9879 4029 9883
rect 4033 9879 4039 9883
rect 4043 9879 4049 9883
rect 4053 9879 4059 9883
rect 4063 9879 4069 9883
rect 3869 9878 4073 9879
rect 3869 9874 3874 9878
rect 3878 9874 3884 9878
rect 3888 9874 3894 9878
rect 3898 9874 3904 9878
rect 3908 9874 4034 9878
rect 4038 9874 4044 9878
rect 4048 9874 4054 9878
rect 4058 9874 4064 9878
rect 4068 9874 4073 9878
rect 3869 9873 4073 9874
rect 3873 9869 3879 9873
rect 3883 9869 3889 9873
rect 3893 9869 3899 9873
rect 3903 9869 3909 9873
rect 3913 9869 4029 9873
rect 4033 9869 4039 9873
rect 4043 9869 4049 9873
rect 4053 9869 4059 9873
rect 4063 9869 4069 9873
rect 3869 9868 4073 9869
rect 3869 9864 3874 9868
rect 3878 9864 3884 9868
rect 3888 9864 3894 9868
rect 3898 9864 3904 9868
rect 3908 9864 4034 9868
rect 4038 9864 4044 9868
rect 4048 9864 4054 9868
rect 4058 9864 4064 9868
rect 4068 9864 4073 9868
rect 1389 9848 1392 9852
rect 1396 9848 1397 9852
rect 1401 9848 1402 9852
rect 1406 9848 1407 9852
rect 1411 9848 1412 9852
rect 1416 9848 1417 9852
rect 1421 9848 1422 9852
rect 1426 9848 1427 9852
rect 1431 9848 1432 9852
rect 1436 9848 1437 9852
rect 1441 9848 1442 9852
rect 1446 9848 1449 9852
rect 1352 9800 1373 9802
rect 1352 9796 1354 9800
rect 1358 9796 1359 9800
rect 1363 9796 1364 9800
rect 1368 9796 1369 9800
rect 1352 9795 1373 9796
rect 1352 9791 1354 9795
rect 1358 9791 1359 9795
rect 1363 9791 1364 9795
rect 1368 9791 1369 9795
rect 1352 9790 1373 9791
rect 1352 9786 1354 9790
rect 1358 9786 1359 9790
rect 1363 9786 1364 9790
rect 1368 9786 1369 9790
rect 118 9348 593 9786
rect 1352 9785 1373 9786
rect 1352 9781 1354 9785
rect 1358 9781 1359 9785
rect 1363 9781 1364 9785
rect 1368 9781 1369 9785
rect 1352 9780 1373 9781
rect 1352 9776 1354 9780
rect 1358 9776 1359 9780
rect 1363 9776 1364 9780
rect 1368 9776 1369 9780
rect 1352 9775 1373 9776
rect 1352 9771 1354 9775
rect 1358 9771 1359 9775
rect 1363 9771 1364 9775
rect 1368 9771 1369 9775
rect 1352 9770 1373 9771
rect 1352 9766 1354 9770
rect 1358 9766 1359 9770
rect 1363 9766 1364 9770
rect 1368 9766 1369 9770
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 802 9761 821 9762
rect 806 9757 807 9761
rect 811 9757 812 9761
rect 816 9757 817 9761
rect 802 9756 821 9757
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 802 9751 821 9752
rect 806 9747 807 9751
rect 811 9747 812 9751
rect 816 9747 817 9751
rect 802 9746 821 9747
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 802 9741 821 9742
rect 806 9737 807 9741
rect 811 9737 812 9741
rect 816 9737 817 9741
rect 802 9736 821 9737
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 831 9761 850 9762
rect 835 9757 836 9761
rect 840 9757 841 9761
rect 845 9757 846 9761
rect 831 9756 850 9757
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 831 9751 850 9752
rect 835 9747 836 9751
rect 840 9747 841 9751
rect 845 9747 846 9751
rect 831 9746 850 9747
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 831 9741 850 9742
rect 835 9737 836 9741
rect 840 9737 841 9741
rect 845 9737 846 9741
rect 831 9736 850 9737
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 860 9761 879 9762
rect 864 9757 865 9761
rect 869 9757 870 9761
rect 874 9757 875 9761
rect 860 9756 879 9757
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 860 9751 879 9752
rect 864 9747 865 9751
rect 869 9747 870 9751
rect 874 9747 875 9751
rect 860 9746 879 9747
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 860 9741 879 9742
rect 864 9737 865 9741
rect 869 9737 870 9741
rect 874 9737 875 9741
rect 860 9736 879 9737
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 889 9761 908 9762
rect 893 9757 894 9761
rect 898 9757 899 9761
rect 903 9757 904 9761
rect 889 9756 908 9757
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 889 9751 908 9752
rect 893 9747 894 9751
rect 898 9747 899 9751
rect 903 9747 904 9751
rect 889 9746 908 9747
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 889 9741 908 9742
rect 893 9737 894 9741
rect 898 9737 899 9741
rect 903 9737 904 9741
rect 889 9736 908 9737
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 918 9761 937 9762
rect 922 9757 923 9761
rect 927 9757 928 9761
rect 932 9757 933 9761
rect 918 9756 937 9757
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 918 9751 937 9752
rect 922 9747 923 9751
rect 927 9747 928 9751
rect 932 9747 933 9751
rect 918 9746 937 9747
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 918 9741 937 9742
rect 922 9737 923 9741
rect 927 9737 928 9741
rect 932 9737 933 9741
rect 918 9736 937 9737
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1319 9761 1338 9762
rect 1323 9757 1324 9761
rect 1328 9757 1329 9761
rect 1333 9757 1334 9761
rect 1319 9756 1338 9757
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1319 9751 1338 9752
rect 1323 9747 1324 9751
rect 1328 9747 1329 9751
rect 1333 9747 1334 9751
rect 1319 9746 1338 9747
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1319 9741 1338 9742
rect 1323 9737 1324 9741
rect 1328 9737 1329 9741
rect 1333 9737 1334 9741
rect 1319 9736 1338 9737
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1352 9765 1373 9766
rect 1352 9761 1354 9765
rect 1358 9761 1359 9765
rect 1363 9761 1364 9765
rect 1368 9761 1369 9765
rect 1352 9760 1373 9761
rect 1352 9756 1354 9760
rect 1358 9756 1359 9760
rect 1363 9756 1364 9760
rect 1368 9756 1369 9760
rect 1352 9755 1373 9756
rect 1352 9751 1354 9755
rect 1358 9751 1359 9755
rect 1363 9751 1364 9755
rect 1368 9751 1369 9755
rect 1352 9750 1373 9751
rect 1352 9746 1354 9750
rect 1358 9746 1359 9750
rect 1363 9746 1364 9750
rect 1368 9746 1369 9750
rect 1352 9745 1373 9746
rect 1352 9741 1354 9745
rect 1358 9741 1359 9745
rect 1363 9741 1364 9745
rect 1368 9741 1369 9745
rect 1352 9740 1373 9741
rect 1352 9736 1354 9740
rect 1358 9736 1359 9740
rect 1363 9736 1364 9740
rect 1368 9736 1369 9740
rect 1352 9734 1373 9736
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 802 9715 821 9716
rect 806 9711 807 9715
rect 811 9711 812 9715
rect 816 9711 817 9715
rect 802 9710 821 9711
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 802 9705 821 9706
rect 806 9701 807 9705
rect 811 9701 812 9705
rect 816 9701 817 9705
rect 802 9700 821 9701
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 802 9695 821 9696
rect 806 9691 807 9695
rect 811 9691 812 9695
rect 816 9691 817 9695
rect 802 9690 821 9691
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 831 9715 850 9716
rect 835 9711 836 9715
rect 840 9711 841 9715
rect 845 9711 846 9715
rect 831 9710 850 9711
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 831 9705 850 9706
rect 835 9701 836 9705
rect 840 9701 841 9705
rect 845 9701 846 9705
rect 831 9700 850 9701
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 831 9695 850 9696
rect 835 9691 836 9695
rect 840 9691 841 9695
rect 845 9691 846 9695
rect 831 9690 850 9691
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 860 9715 879 9716
rect 864 9711 865 9715
rect 869 9711 870 9715
rect 874 9711 875 9715
rect 860 9710 879 9711
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 860 9705 879 9706
rect 864 9701 865 9705
rect 869 9701 870 9705
rect 874 9701 875 9705
rect 860 9700 879 9701
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 860 9695 879 9696
rect 864 9691 865 9695
rect 869 9691 870 9695
rect 874 9691 875 9695
rect 860 9690 879 9691
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 889 9715 908 9716
rect 893 9711 894 9715
rect 898 9711 899 9715
rect 903 9711 904 9715
rect 889 9710 908 9711
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 889 9705 908 9706
rect 893 9701 894 9705
rect 898 9701 899 9705
rect 903 9701 904 9705
rect 889 9700 908 9701
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 889 9695 908 9696
rect 893 9691 894 9695
rect 898 9691 899 9695
rect 903 9691 904 9695
rect 889 9690 908 9691
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 918 9715 937 9716
rect 922 9711 923 9715
rect 927 9711 928 9715
rect 932 9711 933 9715
rect 918 9710 937 9711
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 918 9705 937 9706
rect 922 9701 923 9705
rect 927 9701 928 9705
rect 932 9701 933 9705
rect 918 9700 937 9701
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 918 9695 937 9696
rect 922 9691 923 9695
rect 927 9691 928 9695
rect 932 9691 933 9695
rect 918 9690 937 9691
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1319 9715 1338 9716
rect 1323 9711 1324 9715
rect 1328 9711 1329 9715
rect 1333 9711 1334 9715
rect 1319 9710 1338 9711
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1319 9705 1338 9706
rect 1323 9701 1324 9705
rect 1328 9701 1329 9705
rect 1333 9701 1334 9705
rect 1319 9700 1338 9701
rect 1385 9712 1453 9848
rect 1549 9848 1552 9852
rect 1556 9848 1557 9852
rect 1561 9848 1562 9852
rect 1566 9848 1567 9852
rect 1571 9848 1572 9852
rect 1576 9848 1577 9852
rect 1581 9848 1582 9852
rect 1586 9848 1587 9852
rect 1591 9848 1592 9852
rect 1596 9848 1597 9852
rect 1601 9848 1602 9852
rect 1606 9848 1609 9852
rect 1545 9769 1613 9848
rect 1698 9848 1701 9852
rect 1705 9848 1706 9852
rect 1710 9848 1711 9852
rect 1715 9848 1716 9852
rect 1720 9848 1721 9852
rect 1725 9848 1726 9852
rect 1730 9848 1731 9852
rect 1735 9848 1736 9852
rect 1740 9848 1741 9852
rect 1745 9848 1746 9852
rect 1750 9848 1751 9852
rect 1755 9848 1758 9852
rect 1545 9765 1547 9769
rect 1551 9765 1552 9769
rect 1556 9765 1557 9769
rect 1561 9765 1562 9769
rect 1566 9765 1567 9769
rect 1571 9765 1572 9769
rect 1576 9765 1577 9769
rect 1581 9765 1582 9769
rect 1586 9765 1587 9769
rect 1591 9765 1592 9769
rect 1596 9765 1597 9769
rect 1601 9765 1602 9769
rect 1606 9765 1607 9769
rect 1611 9765 1613 9769
rect 1661 9800 1682 9802
rect 1661 9796 1663 9800
rect 1667 9796 1668 9800
rect 1672 9796 1673 9800
rect 1677 9796 1678 9800
rect 1661 9795 1682 9796
rect 1661 9791 1663 9795
rect 1667 9791 1668 9795
rect 1672 9791 1673 9795
rect 1677 9791 1678 9795
rect 1661 9790 1682 9791
rect 1661 9786 1663 9790
rect 1667 9786 1668 9790
rect 1672 9786 1673 9790
rect 1677 9786 1678 9790
rect 1661 9785 1682 9786
rect 1661 9781 1663 9785
rect 1667 9781 1668 9785
rect 1672 9781 1673 9785
rect 1677 9781 1678 9785
rect 1661 9780 1682 9781
rect 1661 9776 1663 9780
rect 1667 9776 1668 9780
rect 1672 9776 1673 9780
rect 1677 9776 1678 9780
rect 1661 9775 1682 9776
rect 1661 9771 1663 9775
rect 1667 9771 1668 9775
rect 1672 9771 1673 9775
rect 1677 9771 1678 9775
rect 1661 9770 1682 9771
rect 1661 9766 1663 9770
rect 1667 9766 1668 9770
rect 1672 9766 1673 9770
rect 1677 9766 1678 9770
rect 1545 9764 1613 9765
rect 1545 9760 1547 9764
rect 1551 9760 1552 9764
rect 1556 9760 1557 9764
rect 1561 9760 1562 9764
rect 1566 9760 1567 9764
rect 1571 9760 1572 9764
rect 1576 9760 1577 9764
rect 1581 9760 1582 9764
rect 1586 9760 1587 9764
rect 1591 9760 1592 9764
rect 1596 9760 1597 9764
rect 1601 9760 1602 9764
rect 1606 9760 1607 9764
rect 1611 9760 1613 9764
rect 1545 9757 1613 9760
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1628 9761 1647 9762
rect 1632 9757 1633 9761
rect 1637 9757 1638 9761
rect 1642 9757 1643 9761
rect 1628 9756 1647 9757
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1628 9751 1647 9752
rect 1632 9747 1633 9751
rect 1637 9747 1638 9751
rect 1642 9747 1643 9751
rect 1628 9746 1647 9747
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1628 9741 1647 9742
rect 1632 9737 1633 9741
rect 1637 9737 1638 9741
rect 1642 9737 1643 9741
rect 1628 9736 1647 9737
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1661 9765 1682 9766
rect 1661 9761 1663 9765
rect 1667 9761 1668 9765
rect 1672 9761 1673 9765
rect 1677 9761 1678 9765
rect 1661 9760 1682 9761
rect 1661 9756 1663 9760
rect 1667 9756 1668 9760
rect 1672 9756 1673 9760
rect 1677 9756 1678 9760
rect 1661 9755 1682 9756
rect 1661 9751 1663 9755
rect 1667 9751 1668 9755
rect 1672 9751 1673 9755
rect 1677 9751 1678 9755
rect 1661 9750 1682 9751
rect 1661 9746 1663 9750
rect 1667 9746 1668 9750
rect 1672 9746 1673 9750
rect 1677 9746 1678 9750
rect 1661 9745 1682 9746
rect 1661 9741 1663 9745
rect 1667 9741 1668 9745
rect 1672 9741 1673 9745
rect 1677 9741 1678 9745
rect 1661 9740 1682 9741
rect 1661 9736 1663 9740
rect 1667 9736 1668 9740
rect 1672 9736 1673 9740
rect 1677 9736 1678 9740
rect 1661 9734 1682 9736
rect 1573 9718 1574 9722
rect 1578 9718 1579 9722
rect 1583 9718 1584 9722
rect 1588 9718 1589 9722
rect 1593 9718 1594 9722
rect 1598 9718 1599 9722
rect 1603 9718 1604 9722
rect 1608 9718 1609 9722
rect 1613 9718 1614 9722
rect 1618 9718 1619 9722
rect 1623 9718 1625 9722
rect 1569 9717 1625 9718
rect 1385 9708 1387 9712
rect 1391 9708 1392 9712
rect 1396 9708 1397 9712
rect 1401 9708 1402 9712
rect 1406 9708 1407 9712
rect 1411 9708 1412 9712
rect 1416 9708 1417 9712
rect 1421 9708 1422 9712
rect 1426 9708 1427 9712
rect 1431 9708 1432 9712
rect 1436 9708 1437 9712
rect 1441 9708 1442 9712
rect 1446 9708 1447 9712
rect 1451 9708 1453 9712
rect 1385 9707 1453 9708
rect 1385 9703 1387 9707
rect 1391 9703 1392 9707
rect 1396 9703 1397 9707
rect 1401 9703 1402 9707
rect 1406 9703 1407 9707
rect 1411 9703 1412 9707
rect 1416 9703 1417 9707
rect 1421 9703 1422 9707
rect 1426 9703 1427 9707
rect 1431 9703 1432 9707
rect 1436 9703 1437 9707
rect 1441 9703 1442 9707
rect 1446 9703 1447 9707
rect 1451 9703 1453 9707
rect 1385 9700 1453 9703
rect 1488 9711 1489 9715
rect 1493 9711 1494 9715
rect 1498 9711 1499 9715
rect 1503 9711 1504 9715
rect 1488 9710 1508 9711
rect 1488 9706 1489 9710
rect 1493 9706 1494 9710
rect 1498 9706 1499 9710
rect 1503 9706 1504 9710
rect 1488 9705 1508 9706
rect 1488 9701 1489 9705
rect 1493 9701 1494 9705
rect 1498 9701 1499 9705
rect 1503 9701 1504 9705
rect 1573 9713 1574 9717
rect 1578 9713 1579 9717
rect 1583 9713 1584 9717
rect 1588 9713 1589 9717
rect 1593 9713 1594 9717
rect 1598 9713 1599 9717
rect 1603 9713 1604 9717
rect 1608 9713 1609 9717
rect 1613 9713 1614 9717
rect 1618 9713 1619 9717
rect 1623 9713 1625 9717
rect 1569 9712 1625 9713
rect 1573 9708 1574 9712
rect 1578 9708 1579 9712
rect 1583 9708 1584 9712
rect 1588 9708 1589 9712
rect 1593 9708 1594 9712
rect 1598 9708 1599 9712
rect 1603 9708 1604 9712
rect 1608 9708 1609 9712
rect 1613 9708 1614 9712
rect 1618 9708 1619 9712
rect 1623 9708 1625 9712
rect 1569 9707 1625 9708
rect 1573 9703 1574 9707
rect 1578 9703 1579 9707
rect 1583 9703 1584 9707
rect 1588 9703 1589 9707
rect 1593 9703 1594 9707
rect 1598 9703 1599 9707
rect 1603 9703 1604 9707
rect 1608 9703 1609 9707
rect 1613 9703 1614 9707
rect 1618 9703 1619 9707
rect 1623 9703 1625 9707
rect 1569 9701 1625 9703
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1628 9715 1647 9716
rect 1632 9711 1633 9715
rect 1637 9711 1638 9715
rect 1642 9711 1643 9715
rect 1628 9710 1647 9711
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1628 9705 1647 9706
rect 1632 9701 1633 9705
rect 1637 9701 1638 9705
rect 1642 9701 1643 9705
rect 1488 9700 1508 9701
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1319 9695 1338 9696
rect 1323 9691 1324 9695
rect 1328 9691 1329 9695
rect 1333 9691 1334 9695
rect 1319 9690 1338 9691
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1488 9696 1489 9700
rect 1493 9696 1494 9700
rect 1498 9696 1499 9700
rect 1503 9696 1504 9700
rect 1488 9695 1508 9696
rect 1488 9691 1489 9695
rect 1493 9691 1494 9695
rect 1498 9691 1499 9695
rect 1503 9691 1504 9695
rect 1488 9690 1508 9691
rect 1488 9686 1489 9690
rect 1493 9686 1494 9690
rect 1498 9686 1499 9690
rect 1503 9686 1504 9690
rect 1628 9700 1647 9701
rect 1694 9712 1762 9848
rect 1858 9848 1861 9852
rect 1865 9848 1866 9852
rect 1870 9848 1871 9852
rect 1875 9848 1876 9852
rect 1880 9848 1881 9852
rect 1885 9848 1886 9852
rect 1890 9848 1891 9852
rect 1895 9848 1896 9852
rect 1900 9848 1901 9852
rect 1905 9848 1906 9852
rect 1910 9848 1911 9852
rect 1915 9848 1918 9852
rect 1778 9815 1782 9827
rect 1778 9799 1782 9811
rect 1778 9783 1782 9795
rect 1836 9815 1840 9827
rect 1836 9799 1840 9811
rect 1836 9783 1840 9795
rect 1854 9769 1922 9848
rect 2007 9848 2010 9852
rect 2014 9848 2015 9852
rect 2019 9848 2020 9852
rect 2024 9848 2025 9852
rect 2029 9848 2030 9852
rect 2034 9848 2035 9852
rect 2039 9848 2040 9852
rect 2044 9848 2045 9852
rect 2049 9848 2050 9852
rect 2054 9848 2055 9852
rect 2059 9848 2060 9852
rect 2064 9848 2067 9852
rect 1854 9765 1856 9769
rect 1860 9765 1861 9769
rect 1865 9765 1866 9769
rect 1870 9765 1871 9769
rect 1875 9765 1876 9769
rect 1880 9765 1881 9769
rect 1885 9765 1886 9769
rect 1890 9765 1891 9769
rect 1895 9765 1896 9769
rect 1900 9765 1901 9769
rect 1905 9765 1906 9769
rect 1910 9765 1911 9769
rect 1915 9765 1916 9769
rect 1920 9765 1922 9769
rect 1970 9800 1991 9802
rect 1970 9796 1972 9800
rect 1976 9796 1977 9800
rect 1981 9796 1982 9800
rect 1986 9796 1987 9800
rect 1970 9795 1991 9796
rect 1970 9791 1972 9795
rect 1976 9791 1977 9795
rect 1981 9791 1982 9795
rect 1986 9791 1987 9795
rect 1970 9790 1991 9791
rect 1970 9786 1972 9790
rect 1976 9786 1977 9790
rect 1981 9786 1982 9790
rect 1986 9786 1987 9790
rect 1970 9785 1991 9786
rect 1970 9781 1972 9785
rect 1976 9781 1977 9785
rect 1981 9781 1982 9785
rect 1986 9781 1987 9785
rect 1970 9780 1991 9781
rect 1970 9776 1972 9780
rect 1976 9776 1977 9780
rect 1981 9776 1982 9780
rect 1986 9776 1987 9780
rect 1970 9775 1991 9776
rect 1970 9771 1972 9775
rect 1976 9771 1977 9775
rect 1981 9771 1982 9775
rect 1986 9771 1987 9775
rect 1970 9770 1991 9771
rect 1970 9766 1972 9770
rect 1976 9766 1977 9770
rect 1981 9766 1982 9770
rect 1986 9766 1987 9770
rect 1854 9764 1922 9765
rect 1854 9760 1856 9764
rect 1860 9760 1861 9764
rect 1865 9760 1866 9764
rect 1870 9760 1871 9764
rect 1875 9760 1876 9764
rect 1880 9760 1881 9764
rect 1885 9760 1886 9764
rect 1890 9760 1891 9764
rect 1895 9760 1896 9764
rect 1900 9760 1901 9764
rect 1905 9760 1906 9764
rect 1910 9760 1911 9764
rect 1915 9760 1916 9764
rect 1920 9760 1922 9764
rect 1854 9757 1922 9760
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1937 9761 1956 9762
rect 1941 9757 1942 9761
rect 1946 9757 1947 9761
rect 1951 9757 1952 9761
rect 1937 9756 1956 9757
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1937 9751 1956 9752
rect 1941 9747 1942 9751
rect 1946 9747 1947 9751
rect 1951 9747 1952 9751
rect 1937 9746 1956 9747
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1937 9741 1956 9742
rect 1941 9737 1942 9741
rect 1946 9737 1947 9741
rect 1951 9737 1952 9741
rect 1937 9736 1956 9737
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1970 9765 1991 9766
rect 1970 9761 1972 9765
rect 1976 9761 1977 9765
rect 1981 9761 1982 9765
rect 1986 9761 1987 9765
rect 1970 9760 1991 9761
rect 1970 9756 1972 9760
rect 1976 9756 1977 9760
rect 1981 9756 1982 9760
rect 1986 9756 1987 9760
rect 1970 9755 1991 9756
rect 1970 9751 1972 9755
rect 1976 9751 1977 9755
rect 1981 9751 1982 9755
rect 1986 9751 1987 9755
rect 1970 9750 1991 9751
rect 1970 9746 1972 9750
rect 1976 9746 1977 9750
rect 1981 9746 1982 9750
rect 1986 9746 1987 9750
rect 1970 9745 1991 9746
rect 1970 9741 1972 9745
rect 1976 9741 1977 9745
rect 1981 9741 1982 9745
rect 1986 9741 1987 9745
rect 1970 9740 1991 9741
rect 1970 9736 1972 9740
rect 1976 9736 1977 9740
rect 1981 9736 1982 9740
rect 1986 9736 1987 9740
rect 1970 9734 1991 9736
rect 1694 9708 1696 9712
rect 1700 9708 1701 9712
rect 1705 9708 1706 9712
rect 1710 9708 1711 9712
rect 1715 9708 1716 9712
rect 1720 9708 1721 9712
rect 1725 9708 1726 9712
rect 1730 9708 1731 9712
rect 1735 9708 1736 9712
rect 1740 9708 1741 9712
rect 1745 9708 1746 9712
rect 1750 9708 1751 9712
rect 1755 9708 1756 9712
rect 1760 9708 1762 9712
rect 1694 9707 1762 9708
rect 1694 9703 1696 9707
rect 1700 9703 1701 9707
rect 1705 9703 1706 9707
rect 1710 9703 1711 9707
rect 1715 9703 1716 9707
rect 1720 9703 1721 9707
rect 1725 9703 1726 9707
rect 1730 9703 1731 9707
rect 1735 9703 1736 9707
rect 1740 9703 1741 9707
rect 1745 9703 1746 9707
rect 1750 9703 1751 9707
rect 1755 9703 1756 9707
rect 1760 9703 1762 9707
rect 1694 9700 1762 9703
rect 1882 9718 1883 9722
rect 1887 9718 1888 9722
rect 1892 9718 1893 9722
rect 1897 9718 1898 9722
rect 1902 9718 1903 9722
rect 1907 9718 1908 9722
rect 1912 9718 1913 9722
rect 1917 9718 1918 9722
rect 1922 9718 1923 9722
rect 1927 9718 1928 9722
rect 1932 9718 1934 9722
rect 1878 9717 1934 9718
rect 1882 9713 1883 9717
rect 1887 9713 1888 9717
rect 1892 9713 1893 9717
rect 1897 9713 1898 9717
rect 1902 9713 1903 9717
rect 1907 9713 1908 9717
rect 1912 9713 1913 9717
rect 1917 9713 1918 9717
rect 1922 9713 1923 9717
rect 1927 9713 1928 9717
rect 1932 9713 1934 9717
rect 1878 9712 1934 9713
rect 1882 9708 1883 9712
rect 1887 9708 1888 9712
rect 1892 9708 1893 9712
rect 1897 9708 1898 9712
rect 1902 9708 1903 9712
rect 1907 9708 1908 9712
rect 1912 9708 1913 9712
rect 1917 9708 1918 9712
rect 1922 9708 1923 9712
rect 1927 9708 1928 9712
rect 1932 9708 1934 9712
rect 1878 9707 1934 9708
rect 1882 9703 1883 9707
rect 1887 9703 1888 9707
rect 1892 9703 1893 9707
rect 1897 9703 1898 9707
rect 1902 9703 1903 9707
rect 1907 9703 1908 9707
rect 1912 9703 1913 9707
rect 1917 9703 1918 9707
rect 1922 9703 1923 9707
rect 1927 9703 1928 9707
rect 1932 9703 1934 9707
rect 1878 9701 1934 9703
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1937 9715 1956 9716
rect 1941 9711 1942 9715
rect 1946 9711 1947 9715
rect 1951 9711 1952 9715
rect 1937 9710 1956 9711
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1937 9705 1956 9706
rect 1941 9701 1942 9705
rect 1946 9701 1947 9705
rect 1951 9701 1952 9705
rect 1937 9700 1956 9701
rect 2003 9712 2071 9848
rect 2167 9848 2170 9852
rect 2174 9848 2175 9852
rect 2179 9848 2180 9852
rect 2184 9848 2185 9852
rect 2189 9848 2190 9852
rect 2194 9848 2195 9852
rect 2199 9848 2200 9852
rect 2204 9848 2205 9852
rect 2209 9848 2210 9852
rect 2214 9848 2215 9852
rect 2219 9848 2220 9852
rect 2224 9848 2227 9852
rect 2087 9815 2091 9827
rect 2087 9799 2091 9811
rect 2087 9783 2091 9795
rect 2145 9815 2149 9827
rect 2145 9799 2149 9811
rect 2145 9783 2149 9795
rect 2163 9769 2231 9848
rect 2316 9848 2319 9852
rect 2323 9848 2324 9852
rect 2328 9848 2329 9852
rect 2333 9848 2334 9852
rect 2338 9848 2339 9852
rect 2343 9848 2344 9852
rect 2348 9848 2349 9852
rect 2353 9848 2354 9852
rect 2358 9848 2359 9852
rect 2363 9848 2364 9852
rect 2368 9848 2369 9852
rect 2373 9848 2376 9852
rect 2163 9765 2165 9769
rect 2169 9765 2170 9769
rect 2174 9765 2175 9769
rect 2179 9765 2180 9769
rect 2184 9765 2185 9769
rect 2189 9765 2190 9769
rect 2194 9765 2195 9769
rect 2199 9765 2200 9769
rect 2204 9765 2205 9769
rect 2209 9765 2210 9769
rect 2214 9765 2215 9769
rect 2219 9765 2220 9769
rect 2224 9765 2225 9769
rect 2229 9765 2231 9769
rect 2279 9800 2300 9802
rect 2279 9796 2281 9800
rect 2285 9796 2286 9800
rect 2290 9796 2291 9800
rect 2295 9796 2296 9800
rect 2279 9795 2300 9796
rect 2279 9791 2281 9795
rect 2285 9791 2286 9795
rect 2290 9791 2291 9795
rect 2295 9791 2296 9795
rect 2279 9790 2300 9791
rect 2279 9786 2281 9790
rect 2285 9786 2286 9790
rect 2290 9786 2291 9790
rect 2295 9786 2296 9790
rect 2279 9785 2300 9786
rect 2279 9781 2281 9785
rect 2285 9781 2286 9785
rect 2290 9781 2291 9785
rect 2295 9781 2296 9785
rect 2279 9780 2300 9781
rect 2279 9776 2281 9780
rect 2285 9776 2286 9780
rect 2290 9776 2291 9780
rect 2295 9776 2296 9780
rect 2279 9775 2300 9776
rect 2279 9771 2281 9775
rect 2285 9771 2286 9775
rect 2290 9771 2291 9775
rect 2295 9771 2296 9775
rect 2279 9770 2300 9771
rect 2279 9766 2281 9770
rect 2285 9766 2286 9770
rect 2290 9766 2291 9770
rect 2295 9766 2296 9770
rect 2163 9764 2231 9765
rect 2163 9760 2165 9764
rect 2169 9760 2170 9764
rect 2174 9760 2175 9764
rect 2179 9760 2180 9764
rect 2184 9760 2185 9764
rect 2189 9760 2190 9764
rect 2194 9760 2195 9764
rect 2199 9760 2200 9764
rect 2204 9760 2205 9764
rect 2209 9760 2210 9764
rect 2214 9760 2215 9764
rect 2219 9760 2220 9764
rect 2224 9760 2225 9764
rect 2229 9760 2231 9764
rect 2163 9757 2231 9760
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2246 9761 2265 9762
rect 2250 9757 2251 9761
rect 2255 9757 2256 9761
rect 2260 9757 2261 9761
rect 2246 9756 2265 9757
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2246 9751 2265 9752
rect 2250 9747 2251 9751
rect 2255 9747 2256 9751
rect 2260 9747 2261 9751
rect 2246 9746 2265 9747
rect 2003 9708 2005 9712
rect 2009 9708 2010 9712
rect 2014 9708 2015 9712
rect 2019 9708 2020 9712
rect 2024 9708 2025 9712
rect 2029 9708 2030 9712
rect 2034 9708 2035 9712
rect 2039 9708 2040 9712
rect 2044 9708 2045 9712
rect 2049 9708 2050 9712
rect 2054 9708 2055 9712
rect 2059 9708 2060 9712
rect 2064 9708 2065 9712
rect 2069 9708 2071 9712
rect 2003 9707 2071 9708
rect 2003 9703 2005 9707
rect 2009 9703 2010 9707
rect 2014 9703 2015 9707
rect 2019 9703 2020 9707
rect 2024 9703 2025 9707
rect 2029 9703 2030 9707
rect 2034 9703 2035 9707
rect 2039 9703 2040 9707
rect 2044 9703 2045 9707
rect 2049 9703 2050 9707
rect 2054 9703 2055 9707
rect 2059 9703 2060 9707
rect 2064 9703 2065 9707
rect 2069 9703 2071 9707
rect 2003 9700 2071 9703
rect 2166 9741 2174 9743
rect 2166 9736 2167 9741
rect 2172 9736 2174 9741
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1628 9695 1647 9696
rect 1632 9691 1633 9695
rect 1637 9691 1638 9695
rect 1642 9691 1643 9695
rect 1628 9690 1647 9691
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1937 9695 1956 9696
rect 1941 9691 1942 9695
rect 1946 9691 1947 9695
rect 1951 9691 1952 9695
rect 1937 9690 1956 9691
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 1488 9685 1508 9686
rect 1488 9681 1489 9685
rect 1493 9681 1494 9685
rect 1498 9681 1499 9685
rect 1503 9681 1504 9685
rect 1488 9680 1508 9681
rect 1488 9676 1489 9680
rect 1493 9676 1494 9680
rect 1498 9676 1499 9680
rect 1503 9676 1504 9680
rect 1488 9675 1508 9676
rect 1488 9671 1489 9675
rect 1493 9671 1494 9675
rect 1498 9671 1499 9675
rect 1503 9671 1504 9675
rect 1488 9670 1508 9671
rect 1488 9666 1489 9670
rect 1493 9666 1494 9670
rect 1498 9666 1499 9670
rect 1503 9666 1504 9670
rect 1488 9665 1508 9666
rect 1488 9661 1489 9665
rect 1493 9661 1494 9665
rect 1498 9661 1499 9665
rect 1503 9661 1504 9665
rect 1488 9659 1508 9661
rect 2166 9623 2174 9736
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2246 9741 2265 9742
rect 2250 9737 2251 9741
rect 2255 9737 2256 9741
rect 2260 9737 2261 9741
rect 2246 9736 2265 9737
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2279 9765 2300 9766
rect 2279 9761 2281 9765
rect 2285 9761 2286 9765
rect 2290 9761 2291 9765
rect 2295 9761 2296 9765
rect 2279 9760 2300 9761
rect 2279 9756 2281 9760
rect 2285 9756 2286 9760
rect 2290 9756 2291 9760
rect 2295 9756 2296 9760
rect 2279 9755 2300 9756
rect 2279 9751 2281 9755
rect 2285 9751 2286 9755
rect 2290 9751 2291 9755
rect 2295 9751 2296 9755
rect 2279 9750 2300 9751
rect 2279 9746 2281 9750
rect 2285 9746 2286 9750
rect 2290 9746 2291 9750
rect 2295 9746 2296 9750
rect 2279 9745 2300 9746
rect 2279 9741 2281 9745
rect 2285 9741 2286 9745
rect 2290 9741 2291 9745
rect 2295 9741 2296 9745
rect 2279 9740 2300 9741
rect 2279 9736 2281 9740
rect 2285 9736 2286 9740
rect 2290 9736 2291 9740
rect 2295 9736 2296 9740
rect 2279 9734 2300 9736
rect 2191 9718 2192 9722
rect 2196 9718 2197 9722
rect 2201 9718 2202 9722
rect 2206 9718 2207 9722
rect 2211 9718 2212 9722
rect 2216 9718 2217 9722
rect 2221 9718 2222 9722
rect 2226 9718 2227 9722
rect 2231 9718 2232 9722
rect 2236 9718 2237 9722
rect 2241 9718 2243 9722
rect 2187 9717 2243 9718
rect 2191 9713 2192 9717
rect 2196 9713 2197 9717
rect 2201 9713 2202 9717
rect 2206 9713 2207 9717
rect 2211 9713 2212 9717
rect 2216 9713 2217 9717
rect 2221 9713 2222 9717
rect 2226 9713 2227 9717
rect 2231 9713 2232 9717
rect 2236 9713 2237 9717
rect 2241 9713 2243 9717
rect 2187 9712 2243 9713
rect 2191 9708 2192 9712
rect 2196 9708 2197 9712
rect 2201 9708 2202 9712
rect 2206 9708 2207 9712
rect 2211 9708 2212 9712
rect 2216 9708 2217 9712
rect 2221 9708 2222 9712
rect 2226 9708 2227 9712
rect 2231 9708 2232 9712
rect 2236 9708 2237 9712
rect 2241 9708 2243 9712
rect 2187 9707 2243 9708
rect 2191 9703 2192 9707
rect 2196 9703 2197 9707
rect 2201 9703 2202 9707
rect 2206 9703 2207 9707
rect 2211 9703 2212 9707
rect 2216 9703 2217 9707
rect 2221 9703 2222 9707
rect 2226 9703 2227 9707
rect 2231 9703 2232 9707
rect 2236 9703 2237 9707
rect 2241 9703 2243 9707
rect 2187 9701 2243 9703
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2246 9715 2265 9716
rect 2250 9711 2251 9715
rect 2255 9711 2256 9715
rect 2260 9711 2261 9715
rect 2246 9710 2265 9711
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2246 9705 2265 9706
rect 2250 9701 2251 9705
rect 2255 9701 2256 9705
rect 2260 9701 2261 9705
rect 2246 9700 2265 9701
rect 2312 9712 2380 9848
rect 2476 9848 2479 9852
rect 2483 9848 2484 9852
rect 2488 9848 2489 9852
rect 2493 9848 2494 9852
rect 2498 9848 2499 9852
rect 2503 9848 2504 9852
rect 2508 9848 2509 9852
rect 2513 9848 2514 9852
rect 2518 9848 2519 9852
rect 2523 9848 2524 9852
rect 2528 9848 2529 9852
rect 2533 9848 2536 9852
rect 2396 9815 2400 9827
rect 2396 9799 2400 9811
rect 2396 9783 2400 9795
rect 2454 9815 2458 9827
rect 2454 9799 2458 9811
rect 2454 9783 2458 9795
rect 2472 9769 2540 9848
rect 2625 9848 2628 9852
rect 2632 9848 2633 9852
rect 2637 9848 2638 9852
rect 2642 9848 2643 9852
rect 2647 9848 2648 9852
rect 2652 9848 2653 9852
rect 2657 9848 2658 9852
rect 2662 9848 2663 9852
rect 2667 9848 2668 9852
rect 2672 9848 2673 9852
rect 2677 9848 2678 9852
rect 2682 9848 2685 9852
rect 2472 9765 2474 9769
rect 2478 9765 2479 9769
rect 2483 9765 2484 9769
rect 2488 9765 2489 9769
rect 2493 9765 2494 9769
rect 2498 9765 2499 9769
rect 2503 9765 2504 9769
rect 2508 9765 2509 9769
rect 2513 9765 2514 9769
rect 2518 9765 2519 9769
rect 2523 9765 2524 9769
rect 2528 9765 2529 9769
rect 2533 9765 2534 9769
rect 2538 9765 2540 9769
rect 2588 9800 2609 9802
rect 2588 9796 2590 9800
rect 2594 9796 2595 9800
rect 2599 9796 2600 9800
rect 2604 9796 2605 9800
rect 2588 9795 2609 9796
rect 2588 9791 2590 9795
rect 2594 9791 2595 9795
rect 2599 9791 2600 9795
rect 2604 9791 2605 9795
rect 2588 9790 2609 9791
rect 2588 9786 2590 9790
rect 2594 9786 2595 9790
rect 2599 9786 2600 9790
rect 2604 9786 2605 9790
rect 2588 9785 2609 9786
rect 2588 9781 2590 9785
rect 2594 9781 2595 9785
rect 2599 9781 2600 9785
rect 2604 9781 2605 9785
rect 2588 9780 2609 9781
rect 2588 9776 2590 9780
rect 2594 9776 2595 9780
rect 2599 9776 2600 9780
rect 2604 9776 2605 9780
rect 2588 9775 2609 9776
rect 2588 9771 2590 9775
rect 2594 9771 2595 9775
rect 2599 9771 2600 9775
rect 2604 9771 2605 9775
rect 2588 9770 2609 9771
rect 2588 9766 2590 9770
rect 2594 9766 2595 9770
rect 2599 9766 2600 9770
rect 2604 9766 2605 9770
rect 2472 9764 2540 9765
rect 2472 9760 2474 9764
rect 2478 9760 2479 9764
rect 2483 9760 2484 9764
rect 2488 9760 2489 9764
rect 2493 9760 2494 9764
rect 2498 9760 2499 9764
rect 2503 9760 2504 9764
rect 2508 9760 2509 9764
rect 2513 9760 2514 9764
rect 2518 9760 2519 9764
rect 2523 9760 2524 9764
rect 2528 9760 2529 9764
rect 2533 9760 2534 9764
rect 2538 9760 2540 9764
rect 2472 9757 2540 9760
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2555 9761 2574 9762
rect 2559 9757 2560 9761
rect 2564 9757 2565 9761
rect 2569 9757 2570 9761
rect 2555 9756 2574 9757
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2555 9751 2574 9752
rect 2559 9747 2560 9751
rect 2564 9747 2565 9751
rect 2569 9747 2570 9751
rect 2555 9746 2574 9747
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2555 9741 2574 9742
rect 2559 9737 2560 9741
rect 2564 9737 2565 9741
rect 2569 9737 2570 9741
rect 2555 9736 2574 9737
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2588 9765 2609 9766
rect 2588 9761 2590 9765
rect 2594 9761 2595 9765
rect 2599 9761 2600 9765
rect 2604 9761 2605 9765
rect 2588 9760 2609 9761
rect 2588 9756 2590 9760
rect 2594 9756 2595 9760
rect 2599 9756 2600 9760
rect 2604 9756 2605 9760
rect 2588 9755 2609 9756
rect 2588 9751 2590 9755
rect 2594 9751 2595 9755
rect 2599 9751 2600 9755
rect 2604 9751 2605 9755
rect 2588 9750 2609 9751
rect 2588 9746 2590 9750
rect 2594 9746 2595 9750
rect 2599 9746 2600 9750
rect 2604 9746 2605 9750
rect 2588 9745 2609 9746
rect 2588 9741 2590 9745
rect 2594 9741 2595 9745
rect 2599 9741 2600 9745
rect 2604 9741 2605 9745
rect 2588 9740 2609 9741
rect 2588 9736 2590 9740
rect 2594 9736 2595 9740
rect 2599 9736 2600 9740
rect 2604 9736 2605 9740
rect 2588 9734 2609 9736
rect 2312 9708 2314 9712
rect 2318 9708 2319 9712
rect 2323 9708 2324 9712
rect 2328 9708 2329 9712
rect 2333 9708 2334 9712
rect 2338 9708 2339 9712
rect 2343 9708 2344 9712
rect 2348 9708 2349 9712
rect 2353 9708 2354 9712
rect 2358 9708 2359 9712
rect 2363 9708 2364 9712
rect 2368 9708 2369 9712
rect 2373 9708 2374 9712
rect 2378 9708 2380 9712
rect 2312 9707 2380 9708
rect 2312 9703 2314 9707
rect 2318 9703 2319 9707
rect 2323 9703 2324 9707
rect 2328 9703 2329 9707
rect 2333 9703 2334 9707
rect 2338 9703 2339 9707
rect 2343 9703 2344 9707
rect 2348 9703 2349 9707
rect 2353 9703 2354 9707
rect 2358 9703 2359 9707
rect 2363 9703 2364 9707
rect 2368 9703 2369 9707
rect 2373 9703 2374 9707
rect 2378 9703 2380 9707
rect 2312 9700 2380 9703
rect 2500 9718 2501 9722
rect 2505 9718 2506 9722
rect 2510 9718 2511 9722
rect 2515 9718 2516 9722
rect 2520 9718 2521 9722
rect 2525 9718 2526 9722
rect 2530 9718 2531 9722
rect 2535 9718 2536 9722
rect 2540 9718 2541 9722
rect 2545 9718 2546 9722
rect 2550 9718 2552 9722
rect 2496 9717 2552 9718
rect 2500 9713 2501 9717
rect 2505 9713 2506 9717
rect 2510 9713 2511 9717
rect 2515 9713 2516 9717
rect 2520 9713 2521 9717
rect 2525 9713 2526 9717
rect 2530 9713 2531 9717
rect 2535 9713 2536 9717
rect 2540 9713 2541 9717
rect 2545 9713 2546 9717
rect 2550 9713 2552 9717
rect 2496 9712 2552 9713
rect 2500 9708 2501 9712
rect 2505 9708 2506 9712
rect 2510 9708 2511 9712
rect 2515 9708 2516 9712
rect 2520 9708 2521 9712
rect 2525 9708 2526 9712
rect 2530 9708 2531 9712
rect 2535 9708 2536 9712
rect 2540 9708 2541 9712
rect 2545 9708 2546 9712
rect 2550 9708 2552 9712
rect 2496 9707 2552 9708
rect 2500 9703 2501 9707
rect 2505 9703 2506 9707
rect 2510 9703 2511 9707
rect 2515 9703 2516 9707
rect 2520 9703 2521 9707
rect 2525 9703 2526 9707
rect 2530 9703 2531 9707
rect 2535 9703 2536 9707
rect 2540 9703 2541 9707
rect 2545 9703 2546 9707
rect 2550 9703 2552 9707
rect 2496 9701 2552 9703
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2555 9715 2574 9716
rect 2559 9711 2560 9715
rect 2564 9711 2565 9715
rect 2569 9711 2570 9715
rect 2555 9710 2574 9711
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2555 9705 2574 9706
rect 2559 9701 2560 9705
rect 2564 9701 2565 9705
rect 2569 9701 2570 9705
rect 2555 9700 2574 9701
rect 2621 9712 2689 9848
rect 2785 9848 2788 9852
rect 2792 9848 2793 9852
rect 2797 9848 2798 9852
rect 2802 9848 2803 9852
rect 2807 9848 2808 9852
rect 2812 9848 2813 9852
rect 2817 9848 2818 9852
rect 2822 9848 2823 9852
rect 2827 9848 2828 9852
rect 2832 9848 2833 9852
rect 2837 9848 2838 9852
rect 2842 9848 2845 9852
rect 2705 9815 2709 9827
rect 2705 9799 2709 9811
rect 2705 9783 2709 9795
rect 2763 9815 2767 9827
rect 2763 9799 2767 9811
rect 2763 9783 2767 9795
rect 2781 9769 2849 9848
rect 2934 9848 2937 9852
rect 2941 9848 2942 9852
rect 2946 9848 2947 9852
rect 2951 9848 2952 9852
rect 2956 9848 2957 9852
rect 2961 9848 2962 9852
rect 2966 9848 2967 9852
rect 2971 9848 2972 9852
rect 2976 9848 2977 9852
rect 2981 9848 2982 9852
rect 2986 9848 2987 9852
rect 2991 9848 2994 9852
rect 2781 9765 2783 9769
rect 2787 9765 2788 9769
rect 2792 9765 2793 9769
rect 2797 9765 2798 9769
rect 2802 9765 2803 9769
rect 2807 9765 2808 9769
rect 2812 9765 2813 9769
rect 2817 9765 2818 9769
rect 2822 9765 2823 9769
rect 2827 9765 2828 9769
rect 2832 9765 2833 9769
rect 2837 9765 2838 9769
rect 2842 9765 2843 9769
rect 2847 9765 2849 9769
rect 2897 9800 2918 9802
rect 2897 9796 2899 9800
rect 2903 9796 2904 9800
rect 2908 9796 2909 9800
rect 2913 9796 2914 9800
rect 2897 9795 2918 9796
rect 2897 9791 2899 9795
rect 2903 9791 2904 9795
rect 2908 9791 2909 9795
rect 2913 9791 2914 9795
rect 2897 9790 2918 9791
rect 2897 9786 2899 9790
rect 2903 9786 2904 9790
rect 2908 9786 2909 9790
rect 2913 9786 2914 9790
rect 2897 9785 2918 9786
rect 2897 9781 2899 9785
rect 2903 9781 2904 9785
rect 2908 9781 2909 9785
rect 2913 9781 2914 9785
rect 2897 9780 2918 9781
rect 2897 9776 2899 9780
rect 2903 9776 2904 9780
rect 2908 9776 2909 9780
rect 2913 9776 2914 9780
rect 2897 9775 2918 9776
rect 2897 9771 2899 9775
rect 2903 9771 2904 9775
rect 2908 9771 2909 9775
rect 2913 9771 2914 9775
rect 2897 9770 2918 9771
rect 2897 9766 2899 9770
rect 2903 9766 2904 9770
rect 2908 9766 2909 9770
rect 2913 9766 2914 9770
rect 2781 9764 2849 9765
rect 2781 9760 2783 9764
rect 2787 9760 2788 9764
rect 2792 9760 2793 9764
rect 2797 9760 2798 9764
rect 2802 9760 2803 9764
rect 2807 9760 2808 9764
rect 2812 9760 2813 9764
rect 2817 9760 2818 9764
rect 2822 9760 2823 9764
rect 2827 9760 2828 9764
rect 2832 9760 2833 9764
rect 2837 9760 2838 9764
rect 2842 9760 2843 9764
rect 2847 9760 2849 9764
rect 2781 9757 2849 9760
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2864 9761 2883 9762
rect 2868 9757 2869 9761
rect 2873 9757 2874 9761
rect 2878 9757 2879 9761
rect 2864 9756 2883 9757
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2864 9751 2883 9752
rect 2868 9747 2869 9751
rect 2873 9747 2874 9751
rect 2878 9747 2879 9751
rect 2864 9746 2883 9747
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2864 9741 2883 9742
rect 2868 9737 2869 9741
rect 2873 9737 2874 9741
rect 2878 9737 2879 9741
rect 2864 9736 2883 9737
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2897 9765 2918 9766
rect 2897 9761 2899 9765
rect 2903 9761 2904 9765
rect 2908 9761 2909 9765
rect 2913 9761 2914 9765
rect 2897 9760 2918 9761
rect 2897 9756 2899 9760
rect 2903 9756 2904 9760
rect 2908 9756 2909 9760
rect 2913 9756 2914 9760
rect 2897 9755 2918 9756
rect 2897 9751 2899 9755
rect 2903 9751 2904 9755
rect 2908 9751 2909 9755
rect 2913 9751 2914 9755
rect 2897 9750 2918 9751
rect 2897 9746 2899 9750
rect 2903 9746 2904 9750
rect 2908 9746 2909 9750
rect 2913 9746 2914 9750
rect 2897 9745 2918 9746
rect 2897 9741 2899 9745
rect 2903 9741 2904 9745
rect 2908 9741 2909 9745
rect 2913 9741 2914 9745
rect 2897 9740 2918 9741
rect 2897 9736 2899 9740
rect 2903 9736 2904 9740
rect 2908 9736 2909 9740
rect 2913 9736 2914 9740
rect 2897 9734 2918 9736
rect 2621 9708 2623 9712
rect 2627 9708 2628 9712
rect 2632 9708 2633 9712
rect 2637 9708 2638 9712
rect 2642 9708 2643 9712
rect 2647 9708 2648 9712
rect 2652 9708 2653 9712
rect 2657 9708 2658 9712
rect 2662 9708 2663 9712
rect 2667 9708 2668 9712
rect 2672 9708 2673 9712
rect 2677 9708 2678 9712
rect 2682 9708 2683 9712
rect 2687 9708 2689 9712
rect 2621 9707 2689 9708
rect 2621 9703 2623 9707
rect 2627 9703 2628 9707
rect 2632 9703 2633 9707
rect 2637 9703 2638 9707
rect 2642 9703 2643 9707
rect 2647 9703 2648 9707
rect 2652 9703 2653 9707
rect 2657 9703 2658 9707
rect 2662 9703 2663 9707
rect 2667 9703 2668 9707
rect 2672 9703 2673 9707
rect 2677 9703 2678 9707
rect 2682 9703 2683 9707
rect 2687 9703 2689 9707
rect 2621 9700 2689 9703
rect 2809 9718 2810 9722
rect 2814 9718 2815 9722
rect 2819 9718 2820 9722
rect 2824 9718 2825 9722
rect 2829 9718 2830 9722
rect 2834 9718 2835 9722
rect 2839 9718 2840 9722
rect 2844 9718 2845 9722
rect 2849 9718 2850 9722
rect 2854 9718 2855 9722
rect 2859 9718 2861 9722
rect 2805 9717 2861 9718
rect 2809 9713 2810 9717
rect 2814 9713 2815 9717
rect 2819 9713 2820 9717
rect 2824 9713 2825 9717
rect 2829 9713 2830 9717
rect 2834 9713 2835 9717
rect 2839 9713 2840 9717
rect 2844 9713 2845 9717
rect 2849 9713 2850 9717
rect 2854 9713 2855 9717
rect 2859 9713 2861 9717
rect 2805 9712 2861 9713
rect 2809 9708 2810 9712
rect 2814 9708 2815 9712
rect 2819 9708 2820 9712
rect 2824 9708 2825 9712
rect 2829 9708 2830 9712
rect 2834 9708 2835 9712
rect 2839 9708 2840 9712
rect 2844 9708 2845 9712
rect 2849 9708 2850 9712
rect 2854 9708 2855 9712
rect 2859 9708 2861 9712
rect 2805 9707 2861 9708
rect 2809 9703 2810 9707
rect 2814 9703 2815 9707
rect 2819 9703 2820 9707
rect 2824 9703 2825 9707
rect 2829 9703 2830 9707
rect 2834 9703 2835 9707
rect 2839 9703 2840 9707
rect 2844 9703 2845 9707
rect 2849 9703 2850 9707
rect 2854 9703 2855 9707
rect 2859 9703 2861 9707
rect 2805 9701 2861 9703
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2864 9715 2883 9716
rect 2868 9711 2869 9715
rect 2873 9711 2874 9715
rect 2878 9711 2879 9715
rect 2864 9710 2883 9711
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2864 9705 2883 9706
rect 2868 9701 2869 9705
rect 2873 9701 2874 9705
rect 2878 9701 2879 9705
rect 2864 9700 2883 9701
rect 2930 9712 2998 9848
rect 3094 9848 3097 9852
rect 3101 9848 3102 9852
rect 3106 9848 3107 9852
rect 3111 9848 3112 9852
rect 3116 9848 3117 9852
rect 3121 9848 3122 9852
rect 3126 9848 3127 9852
rect 3131 9848 3132 9852
rect 3136 9848 3137 9852
rect 3141 9848 3142 9852
rect 3146 9848 3147 9852
rect 3151 9848 3154 9852
rect 3014 9815 3018 9827
rect 3014 9799 3018 9811
rect 3014 9783 3018 9795
rect 3072 9815 3076 9827
rect 3072 9799 3076 9811
rect 3072 9783 3076 9795
rect 3090 9769 3158 9848
rect 3243 9848 3246 9852
rect 3250 9848 3251 9852
rect 3255 9848 3256 9852
rect 3260 9848 3261 9852
rect 3265 9848 3266 9852
rect 3270 9848 3271 9852
rect 3275 9848 3276 9852
rect 3280 9848 3281 9852
rect 3285 9848 3286 9852
rect 3290 9848 3291 9852
rect 3295 9848 3296 9852
rect 3300 9848 3303 9852
rect 3090 9765 3092 9769
rect 3096 9765 3097 9769
rect 3101 9765 3102 9769
rect 3106 9765 3107 9769
rect 3111 9765 3112 9769
rect 3116 9765 3117 9769
rect 3121 9765 3122 9769
rect 3126 9765 3127 9769
rect 3131 9765 3132 9769
rect 3136 9765 3137 9769
rect 3141 9765 3142 9769
rect 3146 9765 3147 9769
rect 3151 9765 3152 9769
rect 3156 9765 3158 9769
rect 3206 9800 3227 9802
rect 3206 9796 3208 9800
rect 3212 9796 3213 9800
rect 3217 9796 3218 9800
rect 3222 9796 3223 9800
rect 3206 9795 3227 9796
rect 3206 9791 3208 9795
rect 3212 9791 3213 9795
rect 3217 9791 3218 9795
rect 3222 9791 3223 9795
rect 3206 9790 3227 9791
rect 3206 9786 3208 9790
rect 3212 9786 3213 9790
rect 3217 9786 3218 9790
rect 3222 9786 3223 9790
rect 3206 9785 3227 9786
rect 3206 9781 3208 9785
rect 3212 9781 3213 9785
rect 3217 9781 3218 9785
rect 3222 9781 3223 9785
rect 3206 9780 3227 9781
rect 3206 9776 3208 9780
rect 3212 9776 3213 9780
rect 3217 9776 3218 9780
rect 3222 9776 3223 9780
rect 3206 9775 3227 9776
rect 3206 9771 3208 9775
rect 3212 9771 3213 9775
rect 3217 9771 3218 9775
rect 3222 9771 3223 9775
rect 3206 9770 3227 9771
rect 3206 9766 3208 9770
rect 3212 9766 3213 9770
rect 3217 9766 3218 9770
rect 3222 9766 3223 9770
rect 3090 9764 3158 9765
rect 3090 9760 3092 9764
rect 3096 9760 3097 9764
rect 3101 9760 3102 9764
rect 3106 9760 3107 9764
rect 3111 9760 3112 9764
rect 3116 9760 3117 9764
rect 3121 9760 3122 9764
rect 3126 9760 3127 9764
rect 3131 9760 3132 9764
rect 3136 9760 3137 9764
rect 3141 9760 3142 9764
rect 3146 9760 3147 9764
rect 3151 9760 3152 9764
rect 3156 9760 3158 9764
rect 3090 9757 3158 9760
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3173 9761 3192 9762
rect 3177 9757 3178 9761
rect 3182 9757 3183 9761
rect 3187 9757 3188 9761
rect 3173 9756 3192 9757
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3173 9751 3192 9752
rect 3177 9747 3178 9751
rect 3182 9747 3183 9751
rect 3187 9747 3188 9751
rect 3173 9746 3192 9747
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3173 9741 3192 9742
rect 3177 9737 3178 9741
rect 3182 9737 3183 9741
rect 3187 9737 3188 9741
rect 3173 9736 3192 9737
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3206 9765 3227 9766
rect 3206 9761 3208 9765
rect 3212 9761 3213 9765
rect 3217 9761 3218 9765
rect 3222 9761 3223 9765
rect 3206 9760 3227 9761
rect 3206 9756 3208 9760
rect 3212 9756 3213 9760
rect 3217 9756 3218 9760
rect 3222 9756 3223 9760
rect 3206 9755 3227 9756
rect 3206 9751 3208 9755
rect 3212 9751 3213 9755
rect 3217 9751 3218 9755
rect 3222 9751 3223 9755
rect 3206 9750 3227 9751
rect 3206 9746 3208 9750
rect 3212 9746 3213 9750
rect 3217 9746 3218 9750
rect 3222 9746 3223 9750
rect 3206 9745 3227 9746
rect 3206 9741 3208 9745
rect 3212 9741 3213 9745
rect 3217 9741 3218 9745
rect 3222 9741 3223 9745
rect 3206 9740 3227 9741
rect 3206 9736 3208 9740
rect 3212 9736 3213 9740
rect 3217 9736 3218 9740
rect 3222 9736 3223 9740
rect 3206 9734 3227 9736
rect 2930 9708 2932 9712
rect 2936 9708 2937 9712
rect 2941 9708 2942 9712
rect 2946 9708 2947 9712
rect 2951 9708 2952 9712
rect 2956 9708 2957 9712
rect 2961 9708 2962 9712
rect 2966 9708 2967 9712
rect 2971 9708 2972 9712
rect 2976 9708 2977 9712
rect 2981 9708 2982 9712
rect 2986 9708 2987 9712
rect 2991 9708 2992 9712
rect 2996 9708 2998 9712
rect 2930 9707 2998 9708
rect 2930 9703 2932 9707
rect 2936 9703 2937 9707
rect 2941 9703 2942 9707
rect 2946 9703 2947 9707
rect 2951 9703 2952 9707
rect 2956 9703 2957 9707
rect 2961 9703 2962 9707
rect 2966 9703 2967 9707
rect 2971 9703 2972 9707
rect 2976 9703 2977 9707
rect 2981 9703 2982 9707
rect 2986 9703 2987 9707
rect 2991 9703 2992 9707
rect 2996 9703 2998 9707
rect 2930 9700 2998 9703
rect 3118 9718 3119 9722
rect 3123 9718 3124 9722
rect 3128 9718 3129 9722
rect 3133 9718 3134 9722
rect 3138 9718 3139 9722
rect 3143 9718 3144 9722
rect 3148 9718 3149 9722
rect 3153 9718 3154 9722
rect 3158 9718 3159 9722
rect 3163 9718 3164 9722
rect 3168 9718 3170 9722
rect 3114 9717 3170 9718
rect 3118 9713 3119 9717
rect 3123 9713 3124 9717
rect 3128 9713 3129 9717
rect 3133 9713 3134 9717
rect 3138 9713 3139 9717
rect 3143 9713 3144 9717
rect 3148 9713 3149 9717
rect 3153 9713 3154 9717
rect 3158 9713 3159 9717
rect 3163 9713 3164 9717
rect 3168 9713 3170 9717
rect 3114 9712 3170 9713
rect 3118 9708 3119 9712
rect 3123 9708 3124 9712
rect 3128 9708 3129 9712
rect 3133 9708 3134 9712
rect 3138 9708 3139 9712
rect 3143 9708 3144 9712
rect 3148 9708 3149 9712
rect 3153 9708 3154 9712
rect 3158 9708 3159 9712
rect 3163 9708 3164 9712
rect 3168 9708 3170 9712
rect 3114 9707 3170 9708
rect 3118 9703 3119 9707
rect 3123 9703 3124 9707
rect 3128 9703 3129 9707
rect 3133 9703 3134 9707
rect 3138 9703 3139 9707
rect 3143 9703 3144 9707
rect 3148 9703 3149 9707
rect 3153 9703 3154 9707
rect 3158 9703 3159 9707
rect 3163 9703 3164 9707
rect 3168 9703 3170 9707
rect 3114 9701 3170 9703
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3173 9715 3192 9716
rect 3177 9711 3178 9715
rect 3182 9711 3183 9715
rect 3187 9711 3188 9715
rect 3173 9710 3192 9711
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3173 9705 3192 9706
rect 3177 9701 3178 9705
rect 3182 9701 3183 9705
rect 3187 9701 3188 9705
rect 3173 9700 3192 9701
rect 3239 9712 3307 9848
rect 3403 9848 3406 9852
rect 3410 9848 3411 9852
rect 3415 9848 3416 9852
rect 3420 9848 3421 9852
rect 3425 9848 3426 9852
rect 3430 9848 3431 9852
rect 3435 9848 3436 9852
rect 3440 9848 3441 9852
rect 3445 9848 3446 9852
rect 3450 9848 3451 9852
rect 3455 9848 3456 9852
rect 3460 9848 3463 9852
rect 3399 9769 3467 9848
rect 3552 9848 3555 9852
rect 3559 9848 3560 9852
rect 3564 9848 3565 9852
rect 3569 9848 3570 9852
rect 3574 9848 3575 9852
rect 3579 9848 3580 9852
rect 3584 9848 3585 9852
rect 3589 9848 3590 9852
rect 3594 9848 3595 9852
rect 3599 9848 3600 9852
rect 3604 9848 3605 9852
rect 3609 9848 3612 9852
rect 3399 9765 3401 9769
rect 3405 9765 3406 9769
rect 3410 9765 3411 9769
rect 3415 9765 3416 9769
rect 3420 9765 3421 9769
rect 3425 9765 3426 9769
rect 3430 9765 3431 9769
rect 3435 9765 3436 9769
rect 3440 9765 3441 9769
rect 3445 9765 3446 9769
rect 3450 9765 3451 9769
rect 3455 9765 3456 9769
rect 3460 9765 3461 9769
rect 3465 9765 3467 9769
rect 3515 9800 3536 9802
rect 3515 9796 3517 9800
rect 3521 9796 3522 9800
rect 3526 9796 3527 9800
rect 3531 9796 3532 9800
rect 3515 9795 3536 9796
rect 3515 9791 3517 9795
rect 3521 9791 3522 9795
rect 3526 9791 3527 9795
rect 3531 9791 3532 9795
rect 3515 9790 3536 9791
rect 3515 9786 3517 9790
rect 3521 9786 3522 9790
rect 3526 9786 3527 9790
rect 3531 9786 3532 9790
rect 3515 9785 3536 9786
rect 3515 9781 3517 9785
rect 3521 9781 3522 9785
rect 3526 9781 3527 9785
rect 3531 9781 3532 9785
rect 3515 9780 3536 9781
rect 3515 9776 3517 9780
rect 3521 9776 3522 9780
rect 3526 9776 3527 9780
rect 3531 9776 3532 9780
rect 3515 9775 3536 9776
rect 3515 9771 3517 9775
rect 3521 9771 3522 9775
rect 3526 9771 3527 9775
rect 3531 9771 3532 9775
rect 3515 9770 3536 9771
rect 3515 9766 3517 9770
rect 3521 9766 3522 9770
rect 3526 9766 3527 9770
rect 3531 9766 3532 9770
rect 3399 9764 3467 9765
rect 3399 9760 3401 9764
rect 3405 9760 3406 9764
rect 3410 9760 3411 9764
rect 3415 9760 3416 9764
rect 3420 9760 3421 9764
rect 3425 9760 3426 9764
rect 3430 9760 3431 9764
rect 3435 9760 3436 9764
rect 3440 9760 3441 9764
rect 3445 9760 3446 9764
rect 3450 9760 3451 9764
rect 3455 9760 3456 9764
rect 3460 9760 3461 9764
rect 3465 9760 3467 9764
rect 3399 9757 3467 9760
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3482 9761 3501 9762
rect 3486 9757 3487 9761
rect 3491 9757 3492 9761
rect 3496 9757 3497 9761
rect 3482 9756 3501 9757
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3482 9751 3501 9752
rect 3486 9747 3487 9751
rect 3491 9747 3492 9751
rect 3496 9747 3497 9751
rect 3482 9746 3501 9747
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3482 9741 3501 9742
rect 3486 9737 3487 9741
rect 3491 9737 3492 9741
rect 3496 9737 3497 9741
rect 3482 9736 3501 9737
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3515 9765 3536 9766
rect 3515 9761 3517 9765
rect 3521 9761 3522 9765
rect 3526 9761 3527 9765
rect 3531 9761 3532 9765
rect 3515 9760 3536 9761
rect 3515 9756 3517 9760
rect 3521 9756 3522 9760
rect 3526 9756 3527 9760
rect 3531 9756 3532 9760
rect 3515 9755 3536 9756
rect 3515 9751 3517 9755
rect 3521 9751 3522 9755
rect 3526 9751 3527 9755
rect 3531 9751 3532 9755
rect 3515 9750 3536 9751
rect 3515 9746 3517 9750
rect 3521 9746 3522 9750
rect 3526 9746 3527 9750
rect 3531 9746 3532 9750
rect 3515 9745 3536 9746
rect 3515 9741 3517 9745
rect 3521 9741 3522 9745
rect 3526 9741 3527 9745
rect 3531 9741 3532 9745
rect 3515 9740 3536 9741
rect 3515 9736 3517 9740
rect 3521 9736 3522 9740
rect 3526 9736 3527 9740
rect 3531 9736 3532 9740
rect 3515 9734 3536 9736
rect 3427 9718 3428 9722
rect 3432 9718 3433 9722
rect 3437 9718 3438 9722
rect 3442 9718 3443 9722
rect 3447 9718 3448 9722
rect 3452 9718 3453 9722
rect 3457 9718 3458 9722
rect 3462 9718 3463 9722
rect 3467 9718 3468 9722
rect 3472 9718 3473 9722
rect 3477 9718 3479 9722
rect 3423 9717 3479 9718
rect 3239 9708 3241 9712
rect 3245 9708 3246 9712
rect 3250 9708 3251 9712
rect 3255 9708 3256 9712
rect 3260 9708 3261 9712
rect 3265 9708 3266 9712
rect 3270 9708 3271 9712
rect 3275 9708 3276 9712
rect 3280 9708 3281 9712
rect 3285 9708 3286 9712
rect 3290 9708 3291 9712
rect 3295 9708 3296 9712
rect 3300 9708 3301 9712
rect 3305 9708 3307 9712
rect 3239 9707 3307 9708
rect 3239 9703 3241 9707
rect 3245 9703 3246 9707
rect 3250 9703 3251 9707
rect 3255 9703 3256 9707
rect 3260 9703 3261 9707
rect 3265 9703 3266 9707
rect 3270 9703 3271 9707
rect 3275 9703 3276 9707
rect 3280 9703 3281 9707
rect 3285 9703 3286 9707
rect 3290 9703 3291 9707
rect 3295 9703 3296 9707
rect 3300 9703 3301 9707
rect 3305 9703 3307 9707
rect 3239 9700 3307 9703
rect 3342 9711 3343 9715
rect 3347 9711 3348 9715
rect 3352 9711 3353 9715
rect 3357 9711 3358 9715
rect 3342 9710 3362 9711
rect 3342 9706 3343 9710
rect 3347 9706 3348 9710
rect 3352 9706 3353 9710
rect 3357 9706 3358 9710
rect 3342 9705 3362 9706
rect 3342 9701 3343 9705
rect 3347 9701 3348 9705
rect 3352 9701 3353 9705
rect 3357 9701 3358 9705
rect 3427 9713 3428 9717
rect 3432 9713 3433 9717
rect 3437 9713 3438 9717
rect 3442 9713 3443 9717
rect 3447 9713 3448 9717
rect 3452 9713 3453 9717
rect 3457 9713 3458 9717
rect 3462 9713 3463 9717
rect 3467 9713 3468 9717
rect 3472 9713 3473 9717
rect 3477 9713 3479 9717
rect 3423 9712 3479 9713
rect 3427 9708 3428 9712
rect 3432 9708 3433 9712
rect 3437 9708 3438 9712
rect 3442 9708 3443 9712
rect 3447 9708 3448 9712
rect 3452 9708 3453 9712
rect 3457 9708 3458 9712
rect 3462 9708 3463 9712
rect 3467 9708 3468 9712
rect 3472 9708 3473 9712
rect 3477 9708 3479 9712
rect 3423 9707 3479 9708
rect 3427 9703 3428 9707
rect 3432 9703 3433 9707
rect 3437 9703 3438 9707
rect 3442 9703 3443 9707
rect 3447 9703 3448 9707
rect 3452 9703 3453 9707
rect 3457 9703 3458 9707
rect 3462 9703 3463 9707
rect 3467 9703 3468 9707
rect 3472 9703 3473 9707
rect 3477 9703 3479 9707
rect 3423 9701 3479 9703
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3482 9715 3501 9716
rect 3486 9711 3487 9715
rect 3491 9711 3492 9715
rect 3496 9711 3497 9715
rect 3482 9710 3501 9711
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3482 9705 3501 9706
rect 3486 9701 3487 9705
rect 3491 9701 3492 9705
rect 3496 9701 3497 9705
rect 3342 9700 3362 9701
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2246 9695 2265 9696
rect 2250 9691 2251 9695
rect 2255 9691 2256 9695
rect 2260 9691 2261 9695
rect 2246 9690 2265 9691
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2555 9695 2574 9696
rect 2559 9691 2560 9695
rect 2564 9691 2565 9695
rect 2569 9691 2570 9695
rect 2555 9690 2574 9691
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2864 9695 2883 9696
rect 2868 9691 2869 9695
rect 2873 9691 2874 9695
rect 2878 9691 2879 9695
rect 2864 9690 2883 9691
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3173 9695 3192 9696
rect 3177 9691 3178 9695
rect 3182 9691 3183 9695
rect 3187 9691 3188 9695
rect 3173 9690 3192 9691
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3342 9696 3343 9700
rect 3347 9696 3348 9700
rect 3352 9696 3353 9700
rect 3357 9696 3358 9700
rect 3342 9695 3362 9696
rect 3342 9691 3343 9695
rect 3347 9691 3348 9695
rect 3352 9691 3353 9695
rect 3357 9691 3358 9695
rect 3342 9690 3362 9691
rect 3342 9686 3343 9690
rect 3347 9686 3348 9690
rect 3352 9686 3353 9690
rect 3357 9686 3358 9690
rect 3482 9700 3501 9701
rect 3548 9712 3616 9848
rect 3712 9848 3715 9852
rect 3719 9848 3720 9852
rect 3724 9848 3725 9852
rect 3729 9848 3730 9852
rect 3734 9848 3735 9852
rect 3739 9848 3740 9852
rect 3744 9848 3745 9852
rect 3749 9848 3750 9852
rect 3754 9848 3755 9852
rect 3759 9848 3760 9852
rect 3764 9848 3765 9852
rect 3769 9848 3772 9852
rect 3651 9791 3652 9795
rect 3656 9791 3657 9795
rect 3661 9791 3662 9795
rect 3666 9791 3667 9795
rect 3651 9790 3671 9791
rect 3651 9786 3652 9790
rect 3656 9786 3657 9790
rect 3661 9786 3662 9790
rect 3666 9786 3667 9790
rect 3651 9785 3671 9786
rect 3651 9781 3652 9785
rect 3656 9781 3657 9785
rect 3661 9781 3662 9785
rect 3666 9781 3667 9785
rect 3651 9780 3671 9781
rect 3651 9776 3652 9780
rect 3656 9776 3657 9780
rect 3661 9776 3662 9780
rect 3666 9776 3667 9780
rect 3651 9775 3671 9776
rect 3651 9771 3652 9775
rect 3656 9771 3657 9775
rect 3661 9771 3662 9775
rect 3666 9771 3667 9775
rect 3651 9770 3671 9771
rect 3651 9766 3652 9770
rect 3656 9766 3657 9770
rect 3661 9766 3662 9770
rect 3666 9766 3667 9770
rect 3651 9765 3671 9766
rect 3651 9761 3652 9765
rect 3656 9761 3657 9765
rect 3661 9761 3662 9765
rect 3666 9761 3667 9765
rect 3651 9760 3671 9761
rect 3651 9756 3652 9760
rect 3656 9756 3657 9760
rect 3661 9756 3662 9760
rect 3666 9756 3667 9760
rect 3708 9769 3776 9848
rect 3861 9848 3864 9852
rect 3868 9848 3869 9852
rect 3873 9848 3874 9852
rect 3878 9848 3879 9852
rect 3883 9848 3884 9852
rect 3888 9848 3889 9852
rect 3893 9848 3894 9852
rect 3898 9848 3899 9852
rect 3903 9848 3904 9852
rect 3908 9848 3909 9852
rect 3913 9848 3914 9852
rect 3918 9848 3921 9852
rect 3708 9765 3710 9769
rect 3714 9765 3715 9769
rect 3719 9765 3720 9769
rect 3724 9765 3725 9769
rect 3729 9765 3730 9769
rect 3734 9765 3735 9769
rect 3739 9765 3740 9769
rect 3744 9765 3745 9769
rect 3749 9765 3750 9769
rect 3754 9765 3755 9769
rect 3759 9765 3760 9769
rect 3764 9765 3765 9769
rect 3769 9765 3770 9769
rect 3774 9765 3776 9769
rect 3824 9800 3845 9802
rect 3824 9796 3826 9800
rect 3830 9796 3831 9800
rect 3835 9796 3836 9800
rect 3840 9796 3841 9800
rect 3824 9795 3845 9796
rect 3824 9791 3826 9795
rect 3830 9791 3831 9795
rect 3835 9791 3836 9795
rect 3840 9791 3841 9795
rect 3824 9790 3845 9791
rect 3824 9786 3826 9790
rect 3830 9786 3831 9790
rect 3835 9786 3836 9790
rect 3840 9786 3841 9790
rect 3824 9785 3845 9786
rect 3824 9781 3826 9785
rect 3830 9781 3831 9785
rect 3835 9781 3836 9785
rect 3840 9781 3841 9785
rect 3824 9780 3845 9781
rect 3824 9776 3826 9780
rect 3830 9776 3831 9780
rect 3835 9776 3836 9780
rect 3840 9776 3841 9780
rect 3824 9775 3845 9776
rect 3824 9771 3826 9775
rect 3830 9771 3831 9775
rect 3835 9771 3836 9775
rect 3840 9771 3841 9775
rect 3824 9770 3845 9771
rect 3824 9766 3826 9770
rect 3830 9766 3831 9770
rect 3835 9766 3836 9770
rect 3840 9766 3841 9770
rect 3708 9764 3776 9765
rect 3708 9760 3710 9764
rect 3714 9760 3715 9764
rect 3719 9760 3720 9764
rect 3724 9760 3725 9764
rect 3729 9760 3730 9764
rect 3734 9760 3735 9764
rect 3739 9760 3740 9764
rect 3744 9760 3745 9764
rect 3749 9760 3750 9764
rect 3754 9760 3755 9764
rect 3759 9760 3760 9764
rect 3764 9760 3765 9764
rect 3769 9760 3770 9764
rect 3774 9760 3776 9764
rect 3708 9757 3776 9760
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3791 9761 3810 9762
rect 3795 9757 3796 9761
rect 3800 9757 3801 9761
rect 3805 9757 3806 9761
rect 3651 9755 3671 9756
rect 3651 9751 3652 9755
rect 3656 9751 3657 9755
rect 3661 9751 3662 9755
rect 3666 9751 3667 9755
rect 3651 9750 3671 9751
rect 3651 9746 3652 9750
rect 3656 9746 3657 9750
rect 3661 9746 3662 9750
rect 3666 9746 3667 9750
rect 3651 9745 3671 9746
rect 3651 9741 3652 9745
rect 3656 9741 3657 9745
rect 3661 9741 3662 9745
rect 3666 9741 3667 9745
rect 3651 9739 3671 9741
rect 3791 9756 3810 9757
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3791 9751 3810 9752
rect 3795 9747 3796 9751
rect 3800 9747 3801 9751
rect 3805 9747 3806 9751
rect 3791 9746 3810 9747
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3791 9741 3810 9742
rect 3795 9737 3796 9741
rect 3800 9737 3801 9741
rect 3805 9737 3806 9741
rect 3791 9736 3810 9737
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3824 9765 3845 9766
rect 3824 9761 3826 9765
rect 3830 9761 3831 9765
rect 3835 9761 3836 9765
rect 3840 9761 3841 9765
rect 3824 9760 3845 9761
rect 3824 9756 3826 9760
rect 3830 9756 3831 9760
rect 3835 9756 3836 9760
rect 3840 9756 3841 9760
rect 3824 9755 3845 9756
rect 3824 9751 3826 9755
rect 3830 9751 3831 9755
rect 3835 9751 3836 9755
rect 3840 9751 3841 9755
rect 3824 9750 3845 9751
rect 3824 9746 3826 9750
rect 3830 9746 3831 9750
rect 3835 9746 3836 9750
rect 3840 9746 3841 9750
rect 3824 9745 3845 9746
rect 3824 9741 3826 9745
rect 3830 9741 3831 9745
rect 3835 9741 3836 9745
rect 3840 9741 3841 9745
rect 3824 9740 3845 9741
rect 3824 9736 3826 9740
rect 3830 9736 3831 9740
rect 3835 9736 3836 9740
rect 3840 9736 3841 9740
rect 3824 9734 3845 9736
rect 3548 9708 3550 9712
rect 3554 9708 3555 9712
rect 3559 9708 3560 9712
rect 3564 9708 3565 9712
rect 3569 9708 3570 9712
rect 3574 9708 3575 9712
rect 3579 9708 3580 9712
rect 3584 9708 3585 9712
rect 3589 9708 3590 9712
rect 3594 9708 3595 9712
rect 3599 9708 3600 9712
rect 3604 9708 3605 9712
rect 3609 9708 3610 9712
rect 3614 9708 3616 9712
rect 3548 9707 3616 9708
rect 3548 9703 3550 9707
rect 3554 9703 3555 9707
rect 3559 9703 3560 9707
rect 3564 9703 3565 9707
rect 3569 9703 3570 9707
rect 3574 9703 3575 9707
rect 3579 9703 3580 9707
rect 3584 9703 3585 9707
rect 3589 9703 3590 9707
rect 3594 9703 3595 9707
rect 3599 9703 3600 9707
rect 3604 9703 3605 9707
rect 3609 9703 3610 9707
rect 3614 9703 3616 9707
rect 3548 9700 3616 9703
rect 3736 9718 3737 9722
rect 3741 9718 3742 9722
rect 3746 9718 3747 9722
rect 3751 9718 3752 9722
rect 3756 9718 3757 9722
rect 3761 9718 3762 9722
rect 3766 9718 3767 9722
rect 3771 9718 3772 9722
rect 3776 9718 3777 9722
rect 3781 9718 3782 9722
rect 3786 9718 3788 9722
rect 3732 9717 3788 9718
rect 3736 9713 3737 9717
rect 3741 9713 3742 9717
rect 3746 9713 3747 9717
rect 3751 9713 3752 9717
rect 3756 9713 3757 9717
rect 3761 9713 3762 9717
rect 3766 9713 3767 9717
rect 3771 9713 3772 9717
rect 3776 9713 3777 9717
rect 3781 9713 3782 9717
rect 3786 9713 3788 9717
rect 3732 9712 3788 9713
rect 3736 9708 3737 9712
rect 3741 9708 3742 9712
rect 3746 9708 3747 9712
rect 3751 9708 3752 9712
rect 3756 9708 3757 9712
rect 3761 9708 3762 9712
rect 3766 9708 3767 9712
rect 3771 9708 3772 9712
rect 3776 9708 3777 9712
rect 3781 9708 3782 9712
rect 3786 9708 3788 9712
rect 3732 9707 3788 9708
rect 3736 9703 3737 9707
rect 3741 9703 3742 9707
rect 3746 9703 3747 9707
rect 3751 9703 3752 9707
rect 3756 9703 3757 9707
rect 3761 9703 3762 9707
rect 3766 9703 3767 9707
rect 3771 9703 3772 9707
rect 3776 9703 3777 9707
rect 3781 9703 3782 9707
rect 3786 9703 3788 9707
rect 3732 9701 3788 9703
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3791 9715 3810 9716
rect 3795 9711 3796 9715
rect 3800 9711 3801 9715
rect 3805 9711 3806 9715
rect 3791 9710 3810 9711
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3791 9705 3810 9706
rect 3795 9701 3796 9705
rect 3800 9701 3801 9705
rect 3805 9701 3806 9705
rect 3791 9700 3810 9701
rect 3857 9712 3925 9848
rect 4021 9848 4024 9852
rect 4028 9848 4029 9852
rect 4033 9848 4034 9852
rect 4038 9848 4039 9852
rect 4043 9848 4044 9852
rect 4048 9848 4049 9852
rect 4053 9848 4054 9852
rect 4058 9848 4059 9852
rect 4063 9848 4064 9852
rect 4068 9848 4069 9852
rect 4073 9848 4074 9852
rect 4078 9848 4081 9852
rect 3941 9815 3945 9827
rect 3941 9799 3945 9811
rect 3941 9783 3945 9795
rect 3999 9815 4003 9827
rect 3999 9799 4003 9811
rect 3999 9783 4003 9795
rect 4017 9769 4085 9848
rect 4141 9786 5073 10261
rect 4017 9765 4019 9769
rect 4023 9765 4024 9769
rect 4028 9765 4029 9769
rect 4033 9765 4034 9769
rect 4038 9765 4039 9769
rect 4043 9765 4044 9769
rect 4048 9765 4049 9769
rect 4053 9765 4054 9769
rect 4058 9765 4059 9769
rect 4063 9765 4064 9769
rect 4068 9765 4069 9769
rect 4073 9765 4074 9769
rect 4078 9765 4079 9769
rect 4083 9765 4085 9769
rect 4017 9764 4085 9765
rect 4017 9760 4019 9764
rect 4023 9760 4024 9764
rect 4028 9760 4029 9764
rect 4033 9760 4034 9764
rect 4038 9760 4039 9764
rect 4043 9760 4044 9764
rect 4048 9760 4049 9764
rect 4053 9760 4054 9764
rect 4058 9760 4059 9764
rect 4063 9760 4064 9764
rect 4068 9760 4069 9764
rect 4073 9760 4074 9764
rect 4078 9760 4079 9764
rect 4083 9760 4085 9764
rect 4017 9757 4085 9760
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4100 9761 4119 9762
rect 4104 9757 4105 9761
rect 4109 9757 4110 9761
rect 4114 9757 4115 9761
rect 4100 9756 4119 9757
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4100 9751 4119 9752
rect 4104 9747 4105 9751
rect 4109 9747 4110 9751
rect 4114 9747 4115 9751
rect 4100 9746 4119 9747
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4100 9741 4119 9742
rect 4104 9737 4105 9741
rect 4109 9737 4110 9741
rect 4114 9737 4115 9741
rect 4100 9736 4119 9737
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4292 9761 4311 9762
rect 4296 9757 4297 9761
rect 4301 9757 4302 9761
rect 4306 9757 4307 9761
rect 4292 9756 4311 9757
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4292 9751 4311 9752
rect 4296 9747 4297 9751
rect 4301 9747 4302 9751
rect 4306 9747 4307 9751
rect 4292 9746 4311 9747
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4292 9741 4311 9742
rect 4296 9737 4297 9741
rect 4301 9737 4302 9741
rect 4306 9737 4307 9741
rect 4292 9736 4311 9737
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4318 9761 4337 9762
rect 4322 9757 4323 9761
rect 4327 9757 4328 9761
rect 4332 9757 4333 9761
rect 4318 9756 4337 9757
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4318 9751 4337 9752
rect 4322 9747 4323 9751
rect 4327 9747 4328 9751
rect 4332 9747 4333 9751
rect 4318 9746 4337 9747
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4318 9741 4337 9742
rect 4322 9737 4323 9741
rect 4327 9737 4328 9741
rect 4332 9737 4333 9741
rect 4318 9736 4337 9737
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4344 9761 4363 9762
rect 4348 9757 4349 9761
rect 4353 9757 4354 9761
rect 4358 9757 4359 9761
rect 4344 9756 4363 9757
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4344 9751 4363 9752
rect 4348 9747 4349 9751
rect 4353 9747 4354 9751
rect 4358 9747 4359 9751
rect 4344 9746 4363 9747
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4344 9741 4363 9742
rect 4348 9737 4349 9741
rect 4353 9737 4354 9741
rect 4358 9737 4359 9741
rect 4344 9736 4363 9737
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4370 9761 4389 9762
rect 4374 9757 4375 9761
rect 4379 9757 4380 9761
rect 4384 9757 4385 9761
rect 4370 9756 4389 9757
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4370 9751 4389 9752
rect 4374 9747 4375 9751
rect 4379 9747 4380 9751
rect 4384 9747 4385 9751
rect 4370 9746 4389 9747
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4370 9741 4389 9742
rect 4374 9737 4375 9741
rect 4379 9737 4380 9741
rect 4384 9737 4385 9741
rect 4370 9736 4389 9737
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4396 9761 4415 9762
rect 4400 9757 4401 9761
rect 4405 9757 4406 9761
rect 4410 9757 4411 9761
rect 4396 9756 4415 9757
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4396 9751 4415 9752
rect 4400 9747 4401 9751
rect 4405 9747 4406 9751
rect 4410 9747 4411 9751
rect 4396 9746 4415 9747
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4396 9741 4415 9742
rect 4400 9737 4401 9741
rect 4405 9737 4406 9741
rect 4410 9737 4411 9741
rect 4396 9736 4415 9737
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 3857 9708 3859 9712
rect 3863 9708 3864 9712
rect 3868 9708 3869 9712
rect 3873 9708 3874 9712
rect 3878 9708 3879 9712
rect 3883 9708 3884 9712
rect 3888 9708 3889 9712
rect 3893 9708 3894 9712
rect 3898 9708 3899 9712
rect 3903 9708 3904 9712
rect 3908 9708 3909 9712
rect 3913 9708 3914 9712
rect 3918 9708 3919 9712
rect 3923 9708 3925 9712
rect 3857 9707 3925 9708
rect 3857 9703 3859 9707
rect 3863 9703 3864 9707
rect 3868 9703 3869 9707
rect 3873 9703 3874 9707
rect 3878 9703 3879 9707
rect 3883 9703 3884 9707
rect 3888 9703 3889 9707
rect 3893 9703 3894 9707
rect 3898 9703 3899 9707
rect 3903 9703 3904 9707
rect 3908 9703 3909 9707
rect 3913 9703 3914 9707
rect 3918 9703 3919 9707
rect 3923 9703 3925 9707
rect 3857 9700 3925 9703
rect 4045 9718 4046 9722
rect 4050 9718 4051 9722
rect 4055 9718 4056 9722
rect 4060 9718 4061 9722
rect 4065 9718 4066 9722
rect 4070 9718 4071 9722
rect 4075 9718 4076 9722
rect 4080 9718 4081 9722
rect 4085 9718 4086 9722
rect 4090 9718 4091 9722
rect 4095 9718 4097 9722
rect 4041 9717 4097 9718
rect 4045 9713 4046 9717
rect 4050 9713 4051 9717
rect 4055 9713 4056 9717
rect 4060 9713 4061 9717
rect 4065 9713 4066 9717
rect 4070 9713 4071 9717
rect 4075 9713 4076 9717
rect 4080 9713 4081 9717
rect 4085 9713 4086 9717
rect 4090 9713 4091 9717
rect 4095 9713 4097 9717
rect 4041 9712 4097 9713
rect 4045 9708 4046 9712
rect 4050 9708 4051 9712
rect 4055 9708 4056 9712
rect 4060 9708 4061 9712
rect 4065 9708 4066 9712
rect 4070 9708 4071 9712
rect 4075 9708 4076 9712
rect 4080 9708 4081 9712
rect 4085 9708 4086 9712
rect 4090 9708 4091 9712
rect 4095 9708 4097 9712
rect 4041 9707 4097 9708
rect 4045 9703 4046 9707
rect 4050 9703 4051 9707
rect 4055 9703 4056 9707
rect 4060 9703 4061 9707
rect 4065 9703 4066 9707
rect 4070 9703 4071 9707
rect 4075 9703 4076 9707
rect 4080 9703 4081 9707
rect 4085 9703 4086 9707
rect 4090 9703 4091 9707
rect 4095 9703 4097 9707
rect 4041 9701 4097 9703
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4100 9715 4119 9716
rect 4104 9711 4105 9715
rect 4109 9711 4110 9715
rect 4114 9711 4115 9715
rect 4100 9710 4119 9711
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4100 9705 4119 9706
rect 4104 9701 4105 9705
rect 4109 9701 4110 9705
rect 4114 9701 4115 9705
rect 4100 9700 4119 9701
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3482 9695 3501 9696
rect 3486 9691 3487 9695
rect 3491 9691 3492 9695
rect 3496 9691 3497 9695
rect 3482 9690 3501 9691
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3791 9695 3810 9696
rect 3795 9691 3796 9695
rect 3800 9691 3801 9695
rect 3805 9691 3806 9695
rect 3791 9690 3810 9691
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4100 9695 4119 9696
rect 4104 9691 4105 9695
rect 4109 9691 4110 9695
rect 4114 9691 4115 9695
rect 4100 9690 4119 9691
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4292 9715 4311 9716
rect 4296 9711 4297 9715
rect 4301 9711 4302 9715
rect 4306 9711 4307 9715
rect 4292 9710 4311 9711
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4292 9705 4311 9706
rect 4296 9701 4297 9705
rect 4301 9701 4302 9705
rect 4306 9701 4307 9705
rect 4292 9700 4311 9701
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4292 9695 4311 9696
rect 4296 9691 4297 9695
rect 4301 9691 4302 9695
rect 4306 9691 4307 9695
rect 4292 9690 4311 9691
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4318 9715 4337 9716
rect 4322 9711 4323 9715
rect 4327 9711 4328 9715
rect 4332 9711 4333 9715
rect 4318 9710 4337 9711
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4318 9705 4337 9706
rect 4322 9701 4323 9705
rect 4327 9701 4328 9705
rect 4332 9701 4333 9705
rect 4318 9700 4337 9701
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4318 9695 4337 9696
rect 4322 9691 4323 9695
rect 4327 9691 4328 9695
rect 4332 9691 4333 9695
rect 4318 9690 4337 9691
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4344 9715 4363 9716
rect 4348 9711 4349 9715
rect 4353 9711 4354 9715
rect 4358 9711 4359 9715
rect 4344 9710 4363 9711
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4344 9705 4363 9706
rect 4348 9701 4349 9705
rect 4353 9701 4354 9705
rect 4358 9701 4359 9705
rect 4344 9700 4363 9701
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4344 9695 4363 9696
rect 4348 9691 4349 9695
rect 4353 9691 4354 9695
rect 4358 9691 4359 9695
rect 4344 9690 4363 9691
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4370 9715 4389 9716
rect 4374 9711 4375 9715
rect 4379 9711 4380 9715
rect 4384 9711 4385 9715
rect 4370 9710 4389 9711
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4370 9705 4389 9706
rect 4374 9701 4375 9705
rect 4379 9701 4380 9705
rect 4384 9701 4385 9705
rect 4370 9700 4389 9701
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4370 9695 4389 9696
rect 4374 9691 4375 9695
rect 4379 9691 4380 9695
rect 4384 9691 4385 9695
rect 4370 9690 4389 9691
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4396 9715 4415 9716
rect 4400 9711 4401 9715
rect 4405 9711 4406 9715
rect 4410 9711 4411 9715
rect 4396 9710 4415 9711
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4396 9705 4415 9706
rect 4400 9701 4401 9705
rect 4405 9701 4406 9705
rect 4410 9701 4411 9705
rect 4396 9700 4415 9701
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4396 9695 4415 9696
rect 4400 9691 4401 9695
rect 4405 9691 4406 9695
rect 4410 9691 4411 9695
rect 4396 9690 4415 9691
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 3342 9685 3362 9686
rect 3342 9681 3343 9685
rect 3347 9681 3348 9685
rect 3352 9681 3353 9685
rect 3357 9681 3358 9685
rect 3342 9680 3362 9681
rect 3342 9676 3343 9680
rect 3347 9676 3348 9680
rect 3352 9676 3353 9680
rect 3357 9676 3358 9680
rect 3342 9675 3362 9676
rect 3342 9671 3343 9675
rect 3347 9671 3348 9675
rect 3352 9671 3353 9675
rect 3357 9671 3358 9675
rect 3342 9670 3362 9671
rect 3342 9666 3343 9670
rect 3347 9666 3348 9670
rect 3352 9666 3353 9670
rect 3357 9666 3358 9670
rect 3342 9665 3362 9666
rect 3342 9661 3343 9665
rect 3347 9661 3348 9665
rect 3352 9661 3353 9665
rect 3357 9661 3358 9665
rect 3342 9659 3362 9661
rect 617 9618 618 9622
rect 622 9618 623 9622
rect 627 9618 628 9622
rect 632 9618 633 9622
rect 637 9618 638 9622
rect 642 9618 643 9622
rect 613 9617 647 9618
rect 617 9613 618 9617
rect 622 9613 623 9617
rect 627 9613 628 9617
rect 632 9613 633 9617
rect 637 9613 638 9617
rect 642 9613 643 9617
rect 613 9612 647 9613
rect 617 9608 618 9612
rect 622 9608 623 9612
rect 627 9608 628 9612
rect 632 9608 633 9612
rect 637 9608 638 9612
rect 642 9608 643 9612
rect 613 9607 647 9608
rect 617 9603 618 9607
rect 622 9603 623 9607
rect 627 9603 628 9607
rect 632 9603 633 9607
rect 637 9603 638 9607
rect 642 9603 643 9607
rect 663 9618 664 9622
rect 668 9618 669 9622
rect 673 9618 674 9622
rect 678 9618 679 9622
rect 683 9618 684 9622
rect 688 9618 689 9622
rect 659 9617 693 9618
rect 663 9613 664 9617
rect 668 9613 669 9617
rect 673 9613 674 9617
rect 678 9613 679 9617
rect 683 9613 684 9617
rect 688 9613 689 9617
rect 2166 9616 2179 9623
rect 659 9612 693 9613
rect 663 9608 664 9612
rect 668 9608 669 9612
rect 673 9608 674 9612
rect 678 9608 679 9612
rect 683 9608 684 9612
rect 688 9608 689 9612
rect 659 9607 693 9608
rect 663 9603 664 9607
rect 668 9603 669 9607
rect 673 9603 674 9607
rect 678 9603 679 9607
rect 683 9603 684 9607
rect 688 9603 689 9607
rect 617 9592 618 9596
rect 622 9592 623 9596
rect 627 9592 628 9596
rect 632 9592 633 9596
rect 637 9592 638 9596
rect 642 9592 643 9596
rect 613 9591 647 9592
rect 617 9587 618 9591
rect 622 9587 623 9591
rect 627 9587 628 9591
rect 632 9587 633 9591
rect 637 9587 638 9591
rect 642 9587 643 9591
rect 613 9586 647 9587
rect 617 9582 618 9586
rect 622 9582 623 9586
rect 627 9582 628 9586
rect 632 9582 633 9586
rect 637 9582 638 9586
rect 642 9582 643 9586
rect 613 9581 647 9582
rect 617 9577 618 9581
rect 622 9577 623 9581
rect 627 9577 628 9581
rect 632 9577 633 9581
rect 637 9577 638 9581
rect 642 9577 643 9581
rect 663 9592 664 9596
rect 668 9592 669 9596
rect 673 9592 674 9596
rect 678 9592 679 9596
rect 683 9592 684 9596
rect 688 9592 689 9596
rect 659 9591 693 9592
rect 663 9587 664 9591
rect 668 9587 669 9591
rect 673 9587 674 9591
rect 678 9587 679 9591
rect 683 9587 684 9591
rect 688 9587 689 9591
rect 659 9586 693 9587
rect 663 9582 664 9586
rect 668 9582 669 9586
rect 673 9582 674 9586
rect 678 9582 679 9586
rect 683 9582 684 9586
rect 688 9582 689 9586
rect 659 9581 693 9582
rect 663 9577 664 9581
rect 668 9577 669 9581
rect 673 9577 674 9581
rect 678 9577 679 9581
rect 683 9577 684 9581
rect 688 9577 689 9581
rect 2173 9593 2179 9616
rect 2257 9619 2258 9623
rect 2257 9593 2261 9619
rect 2113 9572 2126 9593
rect 617 9566 618 9570
rect 622 9566 623 9570
rect 627 9566 628 9570
rect 632 9566 633 9570
rect 637 9566 638 9570
rect 642 9566 643 9570
rect 613 9565 647 9566
rect 617 9561 618 9565
rect 622 9561 623 9565
rect 627 9561 628 9565
rect 632 9561 633 9565
rect 637 9561 638 9565
rect 642 9561 643 9565
rect 613 9560 647 9561
rect 617 9556 618 9560
rect 622 9556 623 9560
rect 627 9556 628 9560
rect 632 9556 633 9560
rect 637 9556 638 9560
rect 642 9556 643 9560
rect 613 9555 647 9556
rect 617 9551 618 9555
rect 622 9551 623 9555
rect 627 9551 628 9555
rect 632 9551 633 9555
rect 637 9551 638 9555
rect 642 9551 643 9555
rect 663 9566 664 9570
rect 668 9566 669 9570
rect 673 9566 674 9570
rect 678 9566 679 9570
rect 683 9566 684 9570
rect 688 9566 689 9570
rect 659 9565 693 9566
rect 663 9561 664 9565
rect 668 9561 669 9565
rect 673 9561 674 9565
rect 678 9561 679 9565
rect 683 9561 684 9565
rect 688 9561 689 9565
rect 659 9560 693 9561
rect 663 9556 664 9560
rect 668 9556 669 9560
rect 673 9556 674 9560
rect 678 9556 679 9560
rect 683 9556 684 9560
rect 688 9556 689 9560
rect 659 9555 693 9556
rect 663 9551 664 9555
rect 668 9551 669 9555
rect 673 9551 674 9555
rect 678 9551 679 9555
rect 683 9551 684 9555
rect 688 9551 689 9555
rect 2476 9548 2481 9549
rect 617 9540 618 9544
rect 622 9540 623 9544
rect 627 9540 628 9544
rect 632 9540 633 9544
rect 637 9540 638 9544
rect 642 9540 643 9544
rect 613 9539 647 9540
rect 617 9535 618 9539
rect 622 9535 623 9539
rect 627 9535 628 9539
rect 632 9535 633 9539
rect 637 9535 638 9539
rect 642 9535 643 9539
rect 613 9534 647 9535
rect 617 9530 618 9534
rect 622 9530 623 9534
rect 627 9530 628 9534
rect 632 9530 633 9534
rect 637 9530 638 9534
rect 642 9530 643 9534
rect 613 9529 647 9530
rect 617 9525 618 9529
rect 622 9525 623 9529
rect 627 9525 628 9529
rect 632 9525 633 9529
rect 637 9525 638 9529
rect 642 9525 643 9529
rect 663 9540 664 9544
rect 668 9540 669 9544
rect 673 9540 674 9544
rect 678 9540 679 9544
rect 683 9540 684 9544
rect 688 9540 689 9544
rect 659 9539 693 9540
rect 663 9535 664 9539
rect 668 9535 669 9539
rect 673 9535 674 9539
rect 678 9535 679 9539
rect 683 9535 684 9539
rect 688 9535 689 9539
rect 659 9534 693 9535
rect 663 9530 664 9534
rect 668 9530 669 9534
rect 673 9530 674 9534
rect 678 9530 679 9534
rect 683 9530 684 9534
rect 688 9530 689 9534
rect 659 9529 693 9530
rect 663 9525 664 9529
rect 668 9525 669 9529
rect 673 9525 674 9529
rect 678 9525 679 9529
rect 683 9525 684 9529
rect 688 9525 689 9529
rect 617 9514 618 9518
rect 622 9514 623 9518
rect 627 9514 628 9518
rect 632 9514 633 9518
rect 637 9514 638 9518
rect 642 9514 643 9518
rect 613 9513 647 9514
rect 617 9509 618 9513
rect 622 9509 623 9513
rect 627 9509 628 9513
rect 632 9509 633 9513
rect 637 9509 638 9513
rect 642 9509 643 9513
rect 613 9508 647 9509
rect 617 9504 618 9508
rect 622 9504 623 9508
rect 627 9504 628 9508
rect 632 9504 633 9508
rect 637 9504 638 9508
rect 642 9504 643 9508
rect 613 9503 647 9504
rect 617 9499 618 9503
rect 622 9499 623 9503
rect 627 9499 628 9503
rect 632 9499 633 9503
rect 637 9499 638 9503
rect 642 9499 643 9503
rect 663 9514 664 9518
rect 668 9514 669 9518
rect 673 9514 674 9518
rect 678 9514 679 9518
rect 683 9514 684 9518
rect 688 9514 689 9518
rect 659 9513 693 9514
rect 663 9509 664 9513
rect 668 9509 669 9513
rect 673 9509 674 9513
rect 678 9509 679 9513
rect 683 9509 684 9513
rect 688 9509 689 9513
rect 659 9508 693 9509
rect 663 9504 664 9508
rect 668 9504 669 9508
rect 673 9504 674 9508
rect 678 9504 679 9508
rect 683 9504 684 9508
rect 688 9504 689 9508
rect 659 9503 693 9504
rect 663 9499 664 9503
rect 668 9499 669 9503
rect 673 9499 674 9503
rect 678 9499 679 9503
rect 683 9499 684 9503
rect 688 9499 689 9503
rect 617 9321 618 9325
rect 622 9321 623 9325
rect 627 9321 628 9325
rect 632 9321 633 9325
rect 637 9321 638 9325
rect 642 9321 643 9325
rect 613 9320 647 9321
rect 617 9316 618 9320
rect 622 9316 623 9320
rect 627 9316 628 9320
rect 632 9316 633 9320
rect 637 9316 638 9320
rect 642 9316 643 9320
rect 613 9315 647 9316
rect 617 9311 618 9315
rect 622 9311 623 9315
rect 627 9311 628 9315
rect 632 9311 633 9315
rect 637 9311 638 9315
rect 642 9311 643 9315
rect 613 9310 647 9311
rect 86 9304 346 9307
rect 617 9306 618 9310
rect 622 9306 623 9310
rect 627 9306 628 9310
rect 632 9306 633 9310
rect 637 9306 638 9310
rect 642 9306 643 9310
rect 663 9321 664 9325
rect 668 9321 669 9325
rect 673 9321 674 9325
rect 678 9321 679 9325
rect 683 9321 684 9325
rect 688 9321 689 9325
rect 659 9320 693 9321
rect 663 9316 664 9320
rect 668 9316 669 9320
rect 673 9316 674 9320
rect 678 9316 679 9320
rect 683 9316 684 9320
rect 688 9316 689 9320
rect 659 9315 693 9316
rect 663 9311 664 9315
rect 668 9311 669 9315
rect 673 9311 674 9315
rect 678 9311 679 9315
rect 683 9311 684 9315
rect 688 9311 689 9315
rect 659 9310 693 9311
rect 663 9306 664 9310
rect 668 9306 669 9310
rect 673 9306 674 9310
rect 678 9306 679 9310
rect 683 9306 684 9310
rect 688 9306 689 9310
rect 86 9050 89 9304
rect 343 9050 346 9304
rect 86 9047 346 9050
rect 617 9012 618 9016
rect 622 9012 623 9016
rect 627 9012 628 9016
rect 632 9012 633 9016
rect 637 9012 638 9016
rect 642 9012 643 9016
rect 613 9011 647 9012
rect 617 9007 618 9011
rect 622 9007 623 9011
rect 627 9007 628 9011
rect 632 9007 633 9011
rect 637 9007 638 9011
rect 642 9007 643 9011
rect 613 9006 647 9007
rect 617 9002 618 9006
rect 622 9002 623 9006
rect 627 9002 628 9006
rect 632 9002 633 9006
rect 637 9002 638 9006
rect 642 9002 643 9006
rect 613 9001 647 9002
rect 86 8995 346 8998
rect 617 8997 618 9001
rect 622 8997 623 9001
rect 627 8997 628 9001
rect 632 8997 633 9001
rect 637 8997 638 9001
rect 642 8997 643 9001
rect 663 9012 664 9016
rect 668 9012 669 9016
rect 673 9012 674 9016
rect 678 9012 679 9016
rect 683 9012 684 9016
rect 688 9012 689 9016
rect 659 9011 693 9012
rect 663 9007 664 9011
rect 668 9007 669 9011
rect 673 9007 674 9011
rect 678 9007 679 9011
rect 683 9007 684 9011
rect 688 9007 689 9011
rect 659 9006 693 9007
rect 663 9002 664 9006
rect 668 9002 669 9006
rect 673 9002 674 9006
rect 678 9002 679 9006
rect 683 9002 684 9006
rect 688 9002 689 9006
rect 659 9001 693 9002
rect 663 8997 664 9001
rect 668 8997 669 9001
rect 673 8997 674 9001
rect 678 8997 679 9001
rect 683 8997 684 9001
rect 688 8997 689 9001
rect 86 8741 89 8995
rect 343 8741 346 8995
rect 2476 8823 2480 9548
rect 2497 9386 2502 9575
rect 2788 9479 2794 9501
rect 2764 9430 2770 9459
rect 2776 9430 2782 9466
rect 2788 9430 2794 9475
rect 2800 9486 2806 9501
rect 2800 9430 2806 9482
rect 2812 9493 2818 9501
rect 2812 9430 2818 9489
rect 2824 9430 2830 9497
rect 2836 9430 2842 9452
rect 3021 9438 3026 9605
rect 3040 9448 3053 9607
rect 3379 9606 3382 9608
rect 3327 9471 3382 9606
rect 3634 9469 3690 9604
rect 4483 9573 4484 9577
rect 4488 9573 4489 9577
rect 4493 9573 4494 9577
rect 4498 9573 4499 9577
rect 4503 9573 4504 9577
rect 4508 9573 4509 9577
rect 4479 9572 4513 9573
rect 4483 9568 4484 9572
rect 4488 9568 4489 9572
rect 4493 9568 4494 9572
rect 4498 9568 4499 9572
rect 4503 9568 4504 9572
rect 4508 9568 4509 9572
rect 4479 9567 4513 9568
rect 4483 9563 4484 9567
rect 4488 9563 4489 9567
rect 4493 9563 4494 9567
rect 4498 9563 4499 9567
rect 4503 9563 4504 9567
rect 4508 9563 4509 9567
rect 4479 9562 4513 9563
rect 4483 9558 4484 9562
rect 4488 9558 4489 9562
rect 4493 9558 4494 9562
rect 4498 9558 4499 9562
rect 4503 9558 4504 9562
rect 4508 9558 4509 9562
rect 4529 9573 4530 9577
rect 4534 9573 4535 9577
rect 4539 9573 4540 9577
rect 4544 9573 4545 9577
rect 4549 9573 4550 9577
rect 4554 9573 4555 9577
rect 4525 9572 4559 9573
rect 4529 9568 4530 9572
rect 4534 9568 4535 9572
rect 4539 9568 4540 9572
rect 4544 9568 4545 9572
rect 4549 9568 4550 9572
rect 4554 9568 4555 9572
rect 4525 9567 4559 9568
rect 4529 9563 4530 9567
rect 4534 9563 4535 9567
rect 4539 9563 4540 9567
rect 4544 9563 4545 9567
rect 4549 9563 4550 9567
rect 4554 9563 4555 9567
rect 4525 9562 4559 9563
rect 4529 9558 4530 9562
rect 4534 9558 4535 9562
rect 4539 9558 4540 9562
rect 4544 9558 4545 9562
rect 4549 9558 4550 9562
rect 4554 9558 4555 9562
rect 4483 9544 4484 9548
rect 4488 9544 4489 9548
rect 4493 9544 4494 9548
rect 4498 9544 4499 9548
rect 4503 9544 4504 9548
rect 4508 9544 4509 9548
rect 4479 9543 4513 9544
rect 4483 9539 4484 9543
rect 4488 9539 4489 9543
rect 4493 9539 4494 9543
rect 4498 9539 4499 9543
rect 4503 9539 4504 9543
rect 4508 9539 4509 9543
rect 4479 9538 4513 9539
rect 4483 9534 4484 9538
rect 4488 9534 4489 9538
rect 4493 9534 4494 9538
rect 4498 9534 4499 9538
rect 4503 9534 4504 9538
rect 4508 9534 4509 9538
rect 4479 9533 4513 9534
rect 4483 9529 4484 9533
rect 4488 9529 4489 9533
rect 4493 9529 4494 9533
rect 4498 9529 4499 9533
rect 4503 9529 4504 9533
rect 4508 9529 4509 9533
rect 4529 9544 4530 9548
rect 4534 9544 4535 9548
rect 4539 9544 4540 9548
rect 4544 9544 4545 9548
rect 4549 9544 4550 9548
rect 4554 9544 4555 9548
rect 4525 9543 4559 9544
rect 4529 9539 4530 9543
rect 4534 9539 4535 9543
rect 4539 9539 4540 9543
rect 4544 9539 4545 9543
rect 4549 9539 4550 9543
rect 4554 9539 4555 9543
rect 4525 9538 4559 9539
rect 4529 9534 4530 9538
rect 4534 9534 4535 9538
rect 4539 9534 4540 9538
rect 4544 9534 4545 9538
rect 4549 9534 4550 9538
rect 4554 9534 4555 9538
rect 4525 9533 4559 9534
rect 4529 9529 4530 9533
rect 4534 9529 4535 9533
rect 4539 9529 4540 9533
rect 4544 9529 4545 9533
rect 4549 9529 4550 9533
rect 4554 9529 4555 9533
rect 4483 9515 4484 9519
rect 4488 9515 4489 9519
rect 4493 9515 4494 9519
rect 4498 9515 4499 9519
rect 4503 9515 4504 9519
rect 4508 9515 4509 9519
rect 4479 9514 4513 9515
rect 4483 9510 4484 9514
rect 4488 9510 4489 9514
rect 4493 9510 4494 9514
rect 4498 9510 4499 9514
rect 4503 9510 4504 9514
rect 4508 9510 4509 9514
rect 4479 9509 4513 9510
rect 4483 9505 4484 9509
rect 4488 9505 4489 9509
rect 4493 9505 4494 9509
rect 4498 9505 4499 9509
rect 4503 9505 4504 9509
rect 4508 9505 4509 9509
rect 4479 9504 4513 9505
rect 4483 9500 4484 9504
rect 4488 9500 4489 9504
rect 4493 9500 4494 9504
rect 4498 9500 4499 9504
rect 4503 9500 4504 9504
rect 4508 9500 4509 9504
rect 4529 9515 4530 9519
rect 4534 9515 4535 9519
rect 4539 9515 4540 9519
rect 4544 9515 4545 9519
rect 4549 9515 4550 9519
rect 4554 9515 4555 9519
rect 4525 9514 4559 9515
rect 4529 9510 4530 9514
rect 4534 9510 4535 9514
rect 4539 9510 4540 9514
rect 4544 9510 4545 9514
rect 4549 9510 4550 9514
rect 4554 9510 4555 9514
rect 4525 9509 4559 9510
rect 4529 9505 4530 9509
rect 4534 9505 4535 9509
rect 4539 9505 4540 9509
rect 4544 9505 4545 9509
rect 4549 9505 4550 9509
rect 4554 9505 4555 9509
rect 4525 9504 4559 9505
rect 4529 9500 4530 9504
rect 4534 9500 4535 9504
rect 4539 9500 4540 9504
rect 4544 9500 4545 9504
rect 4549 9500 4550 9504
rect 4554 9500 4555 9504
rect 3327 9466 3382 9467
rect 3635 9463 3690 9469
rect 2490 9231 2493 9280
rect 2490 9187 2493 9227
rect 2498 9224 2502 9386
rect 2506 9304 2509 9314
rect 2513 9274 2516 9283
rect 2529 9276 2532 9289
rect 2542 9261 2545 9314
rect 2609 9304 2612 9314
rect 2549 9289 2553 9293
rect 2550 9274 2553 9283
rect 2505 9247 2508 9259
rect 2546 9257 2547 9261
rect 2556 9247 2559 9300
rect 2562 9280 2565 9285
rect 2571 9274 2574 9283
rect 2587 9276 2590 9289
rect 2608 9274 2611 9283
rect 2607 9247 2610 9257
rect 2490 9172 2493 9181
rect 86 8738 346 8741
rect 2351 8711 2355 8819
rect 2374 8802 2377 8812
rect 2381 8772 2384 8781
rect 2397 8774 2400 8787
rect 2410 8759 2413 8812
rect 2477 8802 2480 8812
rect 2417 8787 2421 8791
rect 2418 8772 2421 8781
rect 2373 8745 2376 8757
rect 2414 8755 2415 8759
rect 2424 8745 2427 8798
rect 2430 8778 2433 8783
rect 2439 8772 2442 8781
rect 2455 8774 2458 8787
rect 2476 8772 2479 8781
rect 2492 8772 2495 8781
rect 2475 8745 2478 8755
rect 617 8703 618 8707
rect 622 8703 623 8707
rect 627 8703 628 8707
rect 632 8703 633 8707
rect 637 8703 638 8707
rect 642 8703 643 8707
rect 613 8702 647 8703
rect 617 8698 618 8702
rect 622 8698 623 8702
rect 627 8698 628 8702
rect 632 8698 633 8702
rect 637 8698 638 8702
rect 642 8698 643 8702
rect 613 8697 647 8698
rect 617 8693 618 8697
rect 622 8693 623 8697
rect 627 8693 628 8697
rect 632 8693 633 8697
rect 637 8693 638 8697
rect 642 8693 643 8697
rect 613 8692 647 8693
rect 86 8686 346 8689
rect 617 8688 618 8692
rect 622 8688 623 8692
rect 627 8688 628 8692
rect 632 8688 633 8692
rect 637 8688 638 8692
rect 642 8688 643 8692
rect 663 8703 664 8707
rect 668 8703 669 8707
rect 673 8703 674 8707
rect 678 8703 679 8707
rect 683 8703 684 8707
rect 688 8703 689 8707
rect 659 8702 693 8703
rect 663 8698 664 8702
rect 668 8698 669 8702
rect 673 8698 674 8702
rect 678 8698 679 8702
rect 683 8698 684 8702
rect 688 8698 689 8702
rect 659 8697 693 8698
rect 663 8693 664 8697
rect 668 8693 669 8697
rect 673 8693 674 8697
rect 678 8693 679 8697
rect 683 8693 684 8697
rect 688 8693 689 8697
rect 659 8692 693 8693
rect 663 8688 664 8692
rect 668 8688 669 8692
rect 673 8688 674 8692
rect 678 8688 679 8692
rect 683 8688 684 8692
rect 688 8688 689 8692
rect 86 8432 89 8686
rect 343 8432 346 8686
rect 2367 8640 2370 8734
rect 2492 8731 2495 8768
rect 2498 8724 2502 9220
rect 2615 9233 2619 9367
rect 2764 9344 2770 9391
rect 2764 9311 2770 9340
rect 2624 9281 2627 9283
rect 2624 9274 2627 9277
rect 2624 9240 2627 9270
rect 2764 9267 2770 9307
rect 2505 9202 2508 9212
rect 2506 9172 2509 9181
rect 2527 9174 2530 9187
rect 2543 9172 2546 9181
rect 2552 9178 2555 9183
rect 2507 9145 2510 9155
rect 2558 9145 2561 9198
rect 2564 9187 2568 9191
rect 2564 9172 2567 9181
rect 2572 9159 2575 9212
rect 2608 9202 2611 9212
rect 2585 9174 2588 9187
rect 2601 9172 2604 9181
rect 2570 9155 2571 9159
rect 2609 9145 2612 9157
rect 2506 8802 2509 8812
rect 2513 8772 2516 8781
rect 2529 8774 2532 8787
rect 2542 8759 2545 8812
rect 2609 8802 2612 8812
rect 2549 8787 2553 8791
rect 2550 8772 2553 8781
rect 2505 8745 2508 8757
rect 2546 8755 2547 8759
rect 2556 8745 2559 8798
rect 2562 8778 2565 8783
rect 2571 8772 2574 8781
rect 2587 8774 2590 8787
rect 2608 8772 2611 8781
rect 2607 8745 2610 8755
rect 2482 8711 2486 8715
rect 2482 8692 2486 8707
rect 2498 8704 2502 8720
rect 2514 8719 2518 8724
rect 2514 8711 2518 8715
rect 2514 8692 2518 8707
rect 2498 8688 2502 8689
rect 2514 8684 2518 8688
rect 2374 8660 2377 8670
rect 2381 8630 2384 8639
rect 2397 8632 2400 8645
rect 2410 8617 2413 8670
rect 2477 8660 2480 8670
rect 2417 8645 2421 8649
rect 2418 8630 2421 8639
rect 2373 8603 2376 8615
rect 2414 8613 2415 8617
rect 2424 8603 2427 8656
rect 2492 8645 2495 8677
rect 2430 8636 2433 8641
rect 2439 8630 2442 8639
rect 2455 8632 2458 8645
rect 2476 8630 2479 8639
rect 2492 8630 2495 8639
rect 2475 8603 2478 8613
rect 2367 8554 2370 8592
rect 2374 8574 2377 8584
rect 2381 8544 2384 8553
rect 2397 8546 2400 8559
rect 2410 8531 2413 8584
rect 2477 8574 2480 8584
rect 2417 8559 2421 8563
rect 2418 8544 2421 8553
rect 2373 8517 2376 8529
rect 2414 8527 2415 8531
rect 2424 8517 2427 8570
rect 2430 8550 2433 8555
rect 2439 8544 2442 8553
rect 2455 8546 2458 8559
rect 2476 8544 2479 8553
rect 2492 8544 2495 8553
rect 2475 8517 2478 8527
rect 86 8429 346 8432
rect 2367 8414 2370 8506
rect 2492 8503 2495 8540
rect 2374 8434 2377 8444
rect 2381 8404 2384 8413
rect 2397 8406 2400 8419
rect 617 8394 618 8398
rect 622 8394 623 8398
rect 627 8394 628 8398
rect 632 8394 633 8398
rect 637 8394 638 8398
rect 642 8394 643 8398
rect 613 8393 647 8394
rect 617 8389 618 8393
rect 622 8389 623 8393
rect 627 8389 628 8393
rect 632 8389 633 8393
rect 637 8389 638 8393
rect 642 8389 643 8393
rect 613 8388 647 8389
rect 617 8384 618 8388
rect 622 8384 623 8388
rect 627 8384 628 8388
rect 632 8384 633 8388
rect 637 8384 638 8388
rect 642 8384 643 8388
rect 613 8383 647 8384
rect 86 8377 346 8380
rect 617 8379 618 8383
rect 622 8379 623 8383
rect 627 8379 628 8383
rect 632 8379 633 8383
rect 637 8379 638 8383
rect 642 8379 643 8383
rect 663 8394 664 8398
rect 668 8394 669 8398
rect 673 8394 674 8398
rect 678 8394 679 8398
rect 683 8394 684 8398
rect 688 8394 689 8398
rect 659 8393 693 8394
rect 663 8389 664 8393
rect 668 8389 669 8393
rect 673 8389 674 8393
rect 678 8389 679 8393
rect 683 8389 684 8393
rect 688 8389 689 8393
rect 659 8388 693 8389
rect 663 8384 664 8388
rect 668 8384 669 8388
rect 673 8384 674 8388
rect 678 8384 679 8388
rect 683 8384 684 8388
rect 688 8384 689 8388
rect 659 8383 693 8384
rect 663 8379 664 8383
rect 668 8379 669 8383
rect 673 8379 674 8383
rect 678 8379 679 8383
rect 683 8379 684 8383
rect 688 8379 689 8383
rect 2410 8391 2413 8444
rect 2477 8434 2480 8444
rect 2417 8419 2421 8423
rect 2418 8404 2421 8413
rect 86 8123 89 8377
rect 343 8123 346 8377
rect 2373 8377 2376 8389
rect 2414 8387 2415 8391
rect 2424 8377 2427 8430
rect 2492 8419 2495 8451
rect 2430 8410 2433 8415
rect 2439 8404 2442 8413
rect 2455 8406 2458 8419
rect 2476 8404 2479 8413
rect 2492 8404 2495 8413
rect 2475 8377 2478 8387
rect 2490 8249 2493 8298
rect 2490 8205 2493 8245
rect 2498 8242 2502 8684
rect 2506 8660 2509 8670
rect 2513 8630 2516 8639
rect 2529 8632 2532 8645
rect 2542 8617 2545 8670
rect 2609 8660 2612 8670
rect 2549 8645 2553 8649
rect 2550 8630 2553 8639
rect 2505 8603 2508 8615
rect 2546 8613 2547 8617
rect 2556 8603 2559 8656
rect 2562 8636 2565 8641
rect 2571 8630 2574 8639
rect 2587 8632 2590 8645
rect 2608 8630 2611 8639
rect 2607 8603 2610 8613
rect 2506 8574 2509 8584
rect 2513 8544 2516 8553
rect 2529 8546 2532 8559
rect 2542 8531 2545 8584
rect 2609 8574 2612 8584
rect 2549 8559 2553 8563
rect 2550 8544 2553 8553
rect 2505 8517 2508 8529
rect 2546 8527 2547 8531
rect 2556 8517 2559 8570
rect 2562 8550 2565 8555
rect 2571 8544 2574 8553
rect 2587 8546 2590 8559
rect 2608 8544 2611 8553
rect 2607 8517 2610 8527
rect 2615 8496 2619 9229
rect 2639 9224 2643 9229
rect 2764 9209 2770 9263
rect 2764 9135 2770 9205
rect 2764 9003 2770 9131
rect 2764 8871 2770 8999
rect 2638 8802 2641 8812
rect 2624 8772 2627 8781
rect 2645 8772 2648 8781
rect 2661 8774 2664 8787
rect 2624 8731 2627 8768
rect 2674 8759 2677 8812
rect 2741 8802 2744 8812
rect 2764 8809 2770 8867
rect 2681 8787 2685 8791
rect 2682 8772 2685 8781
rect 2637 8745 2640 8757
rect 2678 8755 2679 8759
rect 2688 8745 2691 8798
rect 2694 8778 2697 8783
rect 2703 8772 2706 8781
rect 2719 8774 2722 8787
rect 2740 8772 2743 8781
rect 2756 8772 2759 8783
rect 2739 8745 2742 8755
rect 2756 8738 2759 8768
rect 2756 8704 2759 8734
rect 2764 8739 2770 8805
rect 2764 8697 2770 8735
rect 2624 8645 2627 8677
rect 2638 8660 2641 8670
rect 2624 8630 2627 8639
rect 2645 8630 2648 8639
rect 2661 8632 2664 8645
rect 2674 8617 2677 8670
rect 2741 8660 2744 8670
rect 2681 8645 2685 8649
rect 2682 8630 2685 8639
rect 2637 8603 2640 8615
rect 2678 8613 2679 8617
rect 2688 8603 2691 8656
rect 2756 8645 2759 8692
rect 2694 8636 2697 8641
rect 2703 8630 2706 8639
rect 2719 8632 2722 8645
rect 2740 8630 2743 8639
rect 2756 8630 2759 8641
rect 2739 8603 2742 8613
rect 2756 8596 2759 8626
rect 2764 8667 2770 8693
rect 2638 8574 2641 8584
rect 2624 8544 2627 8553
rect 2645 8544 2648 8553
rect 2661 8546 2664 8559
rect 2624 8503 2627 8540
rect 2674 8531 2677 8584
rect 2741 8574 2744 8584
rect 2764 8581 2770 8663
rect 2681 8559 2685 8563
rect 2682 8544 2685 8553
rect 2637 8517 2640 8529
rect 2678 8527 2679 8531
rect 2688 8517 2691 8570
rect 2694 8550 2697 8555
rect 2703 8544 2706 8553
rect 2719 8546 2722 8559
rect 2740 8544 2743 8553
rect 2756 8544 2759 8555
rect 2739 8517 2742 8527
rect 2756 8510 2759 8540
rect 2599 8485 2603 8488
rect 2599 8466 2603 8481
rect 2615 8478 2619 8492
rect 2631 8492 2635 8496
rect 2631 8485 2635 8488
rect 2631 8466 2635 8481
rect 2756 8478 2759 8506
rect 2615 8462 2619 8463
rect 2631 8458 2635 8462
rect 2506 8434 2509 8444
rect 2513 8404 2516 8413
rect 2529 8406 2532 8419
rect 2542 8391 2545 8444
rect 2609 8434 2612 8444
rect 2549 8419 2553 8423
rect 2550 8404 2553 8413
rect 2505 8377 2508 8389
rect 2546 8387 2547 8391
rect 2556 8377 2559 8430
rect 2562 8410 2565 8415
rect 2571 8404 2574 8413
rect 2587 8406 2590 8419
rect 2608 8404 2611 8413
rect 2607 8377 2610 8387
rect 2506 8322 2509 8332
rect 2513 8292 2516 8301
rect 2529 8294 2532 8307
rect 2542 8279 2545 8332
rect 2609 8322 2612 8332
rect 2549 8307 2553 8311
rect 2550 8292 2553 8301
rect 2505 8265 2508 8277
rect 2546 8275 2547 8279
rect 2556 8265 2559 8318
rect 2562 8298 2565 8303
rect 2571 8292 2574 8301
rect 2587 8294 2590 8307
rect 2608 8292 2611 8301
rect 2607 8265 2610 8275
rect 2490 8190 2493 8199
rect 86 8120 346 8123
rect 617 8085 618 8089
rect 622 8085 623 8089
rect 627 8085 628 8089
rect 632 8085 633 8089
rect 637 8085 638 8089
rect 642 8085 643 8089
rect 613 8084 647 8085
rect 617 8080 618 8084
rect 622 8080 623 8084
rect 627 8080 628 8084
rect 632 8080 633 8084
rect 637 8080 638 8084
rect 642 8080 643 8084
rect 613 8079 647 8080
rect 617 8075 618 8079
rect 622 8075 623 8079
rect 627 8075 628 8079
rect 632 8075 633 8079
rect 637 8075 638 8079
rect 642 8075 643 8079
rect 613 8074 647 8075
rect 86 8068 346 8071
rect 617 8070 618 8074
rect 622 8070 623 8074
rect 627 8070 628 8074
rect 632 8070 633 8074
rect 637 8070 638 8074
rect 642 8070 643 8074
rect 663 8085 664 8089
rect 668 8085 669 8089
rect 673 8085 674 8089
rect 678 8085 679 8089
rect 683 8085 684 8089
rect 688 8085 689 8089
rect 659 8084 693 8085
rect 663 8080 664 8084
rect 668 8080 669 8084
rect 673 8080 674 8084
rect 678 8080 679 8084
rect 683 8080 684 8084
rect 688 8080 689 8084
rect 659 8079 693 8080
rect 663 8075 664 8079
rect 668 8075 669 8079
rect 673 8075 674 8079
rect 678 8075 679 8079
rect 683 8075 684 8079
rect 688 8075 689 8079
rect 659 8074 693 8075
rect 663 8070 664 8074
rect 668 8070 669 8074
rect 673 8070 674 8074
rect 678 8070 679 8074
rect 683 8070 684 8074
rect 688 8070 689 8074
rect 86 7814 89 8068
rect 343 7814 346 8068
rect 2374 7820 2377 7830
rect 86 7811 346 7814
rect 2381 7790 2384 7799
rect 2397 7792 2400 7805
rect 617 7776 618 7780
rect 622 7776 623 7780
rect 627 7776 628 7780
rect 632 7776 633 7780
rect 637 7776 638 7780
rect 642 7776 643 7780
rect 613 7775 647 7776
rect 617 7771 618 7775
rect 622 7771 623 7775
rect 627 7771 628 7775
rect 632 7771 633 7775
rect 637 7771 638 7775
rect 642 7771 643 7775
rect 613 7770 647 7771
rect 617 7766 618 7770
rect 622 7766 623 7770
rect 627 7766 628 7770
rect 632 7766 633 7770
rect 637 7766 638 7770
rect 642 7766 643 7770
rect 613 7765 647 7766
rect 86 7759 346 7762
rect 617 7761 618 7765
rect 622 7761 623 7765
rect 627 7761 628 7765
rect 632 7761 633 7765
rect 637 7761 638 7765
rect 642 7761 643 7765
rect 663 7776 664 7780
rect 668 7776 669 7780
rect 673 7776 674 7780
rect 678 7776 679 7780
rect 683 7776 684 7780
rect 688 7776 689 7780
rect 659 7775 693 7776
rect 663 7771 664 7775
rect 668 7771 669 7775
rect 673 7771 674 7775
rect 678 7771 679 7775
rect 683 7771 684 7775
rect 688 7771 689 7775
rect 659 7770 693 7771
rect 663 7766 664 7770
rect 668 7766 669 7770
rect 673 7766 674 7770
rect 678 7766 679 7770
rect 683 7766 684 7770
rect 688 7766 689 7770
rect 659 7765 693 7766
rect 663 7761 664 7765
rect 668 7761 669 7765
rect 673 7761 674 7765
rect 678 7761 679 7765
rect 683 7761 684 7765
rect 688 7761 689 7765
rect 2410 7777 2413 7830
rect 2477 7820 2480 7830
rect 2417 7805 2421 7809
rect 2418 7790 2421 7799
rect 2373 7763 2376 7775
rect 2414 7773 2415 7777
rect 2424 7763 2427 7816
rect 2430 7796 2433 7801
rect 2439 7790 2442 7799
rect 2455 7792 2458 7805
rect 2476 7790 2479 7799
rect 2492 7790 2495 7799
rect 2475 7763 2478 7773
rect 86 7505 89 7759
rect 343 7505 346 7759
rect 2367 7658 2370 7752
rect 2492 7749 2495 7786
rect 2498 7742 2502 8238
rect 2615 8251 2619 8458
rect 2624 8419 2627 8451
rect 2638 8434 2641 8444
rect 2624 8404 2627 8413
rect 2645 8404 2648 8413
rect 2661 8406 2664 8419
rect 2674 8391 2677 8444
rect 2741 8434 2744 8444
rect 2681 8419 2685 8423
rect 2682 8404 2685 8413
rect 2637 8377 2640 8389
rect 2678 8387 2679 8391
rect 2688 8377 2691 8430
rect 2756 8419 2759 8466
rect 2694 8410 2697 8415
rect 2703 8404 2706 8413
rect 2719 8406 2722 8419
rect 2740 8404 2743 8413
rect 2756 8411 2759 8415
rect 2764 8441 2770 8577
rect 2756 8404 2759 8407
rect 2739 8377 2742 8387
rect 2764 8362 2770 8437
rect 2764 8329 2770 8358
rect 2624 8299 2627 8301
rect 2624 8292 2627 8295
rect 2624 8258 2627 8288
rect 2764 8285 2770 8325
rect 2505 8220 2508 8230
rect 2506 8190 2509 8199
rect 2527 8192 2530 8205
rect 2543 8190 2546 8199
rect 2552 8196 2555 8201
rect 2507 8163 2510 8173
rect 2558 8163 2561 8216
rect 2564 8205 2568 8209
rect 2564 8190 2567 8199
rect 2572 8177 2575 8230
rect 2608 8220 2611 8230
rect 2585 8192 2588 8205
rect 2601 8190 2604 8199
rect 2570 8173 2571 8177
rect 2609 8163 2612 8175
rect 2506 7820 2509 7830
rect 2513 7790 2516 7799
rect 2529 7792 2532 7805
rect 2542 7777 2545 7830
rect 2609 7820 2612 7830
rect 2549 7805 2553 7809
rect 2550 7790 2553 7799
rect 2505 7763 2508 7775
rect 2546 7773 2547 7777
rect 2556 7763 2559 7816
rect 2562 7796 2565 7801
rect 2571 7790 2574 7799
rect 2587 7792 2590 7805
rect 2608 7790 2611 7799
rect 2607 7763 2610 7773
rect 2482 7729 2486 7734
rect 2482 7710 2486 7725
rect 2498 7722 2502 7738
rect 2514 7738 2518 7742
rect 2514 7729 2518 7734
rect 2514 7710 2518 7725
rect 2498 7706 2502 7707
rect 2514 7702 2518 7706
rect 2374 7678 2377 7688
rect 2381 7648 2384 7657
rect 2397 7650 2400 7663
rect 2410 7635 2413 7688
rect 2477 7678 2480 7688
rect 2417 7663 2421 7667
rect 2418 7648 2421 7657
rect 2373 7621 2376 7633
rect 2414 7631 2415 7635
rect 2424 7621 2427 7674
rect 2492 7663 2495 7695
rect 2430 7654 2433 7659
rect 2439 7648 2442 7657
rect 2455 7650 2458 7663
rect 2476 7648 2479 7657
rect 2492 7648 2495 7657
rect 2475 7621 2478 7631
rect 2367 7572 2370 7610
rect 2374 7592 2377 7602
rect 2381 7562 2384 7571
rect 2397 7564 2400 7577
rect 2410 7549 2413 7602
rect 2477 7592 2480 7602
rect 2417 7577 2421 7581
rect 2418 7562 2421 7571
rect 2373 7535 2376 7547
rect 2414 7545 2415 7549
rect 2424 7535 2427 7588
rect 2430 7568 2433 7573
rect 2439 7562 2442 7571
rect 2455 7564 2458 7577
rect 2476 7562 2479 7571
rect 2492 7562 2495 7571
rect 2475 7535 2478 7545
rect 86 7502 346 7505
rect 617 7467 618 7471
rect 622 7467 623 7471
rect 627 7467 628 7471
rect 632 7467 633 7471
rect 637 7467 638 7471
rect 642 7467 643 7471
rect 613 7466 647 7467
rect 617 7462 618 7466
rect 622 7462 623 7466
rect 627 7462 628 7466
rect 632 7462 633 7466
rect 637 7462 638 7466
rect 642 7462 643 7466
rect 613 7461 647 7462
rect 617 7457 618 7461
rect 622 7457 623 7461
rect 627 7457 628 7461
rect 632 7457 633 7461
rect 637 7457 638 7461
rect 642 7457 643 7461
rect 613 7456 647 7457
rect 86 7450 346 7453
rect 617 7452 618 7456
rect 622 7452 623 7456
rect 627 7452 628 7456
rect 632 7452 633 7456
rect 637 7452 638 7456
rect 642 7452 643 7456
rect 663 7467 664 7471
rect 668 7467 669 7471
rect 673 7467 674 7471
rect 678 7467 679 7471
rect 683 7467 684 7471
rect 688 7467 689 7471
rect 659 7466 693 7467
rect 663 7462 664 7466
rect 668 7462 669 7466
rect 673 7462 674 7466
rect 678 7462 679 7466
rect 683 7462 684 7466
rect 688 7462 689 7466
rect 659 7461 693 7462
rect 663 7457 664 7461
rect 668 7457 669 7461
rect 673 7457 674 7461
rect 678 7457 679 7461
rect 683 7457 684 7461
rect 688 7457 689 7461
rect 659 7456 693 7457
rect 663 7452 664 7456
rect 668 7452 669 7456
rect 673 7452 674 7456
rect 678 7452 679 7456
rect 683 7452 684 7456
rect 688 7452 689 7456
rect 86 7196 89 7450
rect 343 7196 346 7450
rect 2367 7432 2370 7524
rect 2492 7521 2495 7558
rect 2374 7452 2377 7462
rect 2381 7422 2384 7431
rect 2397 7424 2400 7437
rect 2410 7409 2413 7462
rect 2477 7452 2480 7462
rect 2417 7437 2421 7441
rect 2418 7422 2421 7431
rect 2373 7395 2376 7407
rect 2414 7405 2415 7409
rect 2424 7395 2427 7448
rect 2492 7437 2495 7469
rect 2430 7428 2433 7433
rect 2439 7422 2442 7431
rect 2455 7424 2458 7437
rect 2476 7422 2479 7431
rect 2492 7422 2495 7431
rect 2475 7395 2478 7405
rect 2498 7381 2502 7702
rect 2506 7678 2509 7688
rect 2513 7648 2516 7657
rect 2529 7650 2532 7663
rect 2542 7635 2545 7688
rect 2609 7678 2612 7688
rect 2549 7663 2553 7667
rect 2550 7648 2553 7657
rect 2505 7621 2508 7633
rect 2546 7631 2547 7635
rect 2556 7621 2559 7674
rect 2562 7654 2565 7659
rect 2571 7648 2574 7657
rect 2587 7650 2590 7663
rect 2608 7648 2611 7657
rect 2607 7621 2610 7631
rect 2506 7592 2509 7602
rect 2513 7562 2516 7571
rect 2529 7564 2532 7577
rect 2542 7549 2545 7602
rect 2609 7592 2612 7602
rect 2549 7577 2553 7581
rect 2550 7562 2553 7571
rect 2505 7535 2508 7547
rect 2546 7545 2547 7549
rect 2556 7535 2559 7588
rect 2562 7568 2565 7573
rect 2571 7562 2574 7571
rect 2587 7564 2590 7577
rect 2608 7562 2611 7571
rect 2607 7535 2610 7545
rect 2615 7514 2619 8247
rect 2639 8242 2643 8247
rect 2764 8227 2770 8281
rect 2764 8153 2770 8223
rect 2764 8021 2770 8149
rect 2764 7889 2770 8017
rect 2638 7820 2641 7830
rect 2624 7790 2627 7799
rect 2645 7790 2648 7799
rect 2661 7792 2664 7805
rect 2624 7749 2627 7786
rect 2674 7777 2677 7830
rect 2741 7820 2744 7830
rect 2764 7827 2770 7885
rect 2681 7805 2685 7809
rect 2682 7790 2685 7799
rect 2637 7763 2640 7775
rect 2678 7773 2679 7777
rect 2688 7763 2691 7816
rect 2694 7796 2697 7801
rect 2703 7790 2706 7799
rect 2719 7792 2722 7805
rect 2740 7790 2743 7799
rect 2756 7790 2759 7801
rect 2739 7763 2742 7773
rect 2756 7756 2759 7786
rect 2756 7722 2759 7752
rect 2764 7757 2770 7823
rect 2764 7715 2770 7753
rect 2624 7663 2627 7695
rect 2638 7678 2641 7688
rect 2624 7648 2627 7657
rect 2645 7648 2648 7657
rect 2661 7650 2664 7663
rect 2674 7635 2677 7688
rect 2741 7678 2744 7688
rect 2681 7663 2685 7667
rect 2682 7648 2685 7657
rect 2637 7621 2640 7633
rect 2678 7631 2679 7635
rect 2688 7621 2691 7674
rect 2756 7663 2759 7710
rect 2694 7654 2697 7659
rect 2703 7648 2706 7657
rect 2719 7650 2722 7663
rect 2740 7648 2743 7657
rect 2756 7648 2759 7659
rect 2739 7621 2742 7631
rect 2756 7614 2759 7644
rect 2764 7685 2770 7711
rect 2638 7592 2641 7602
rect 2624 7562 2627 7571
rect 2645 7562 2648 7571
rect 2661 7564 2664 7577
rect 2624 7521 2627 7558
rect 2674 7549 2677 7602
rect 2741 7592 2744 7602
rect 2764 7599 2770 7681
rect 2681 7577 2685 7581
rect 2682 7562 2685 7571
rect 2637 7535 2640 7547
rect 2678 7545 2679 7549
rect 2688 7535 2691 7588
rect 2694 7568 2697 7573
rect 2703 7562 2706 7571
rect 2719 7564 2722 7577
rect 2740 7562 2743 7571
rect 2756 7562 2759 7573
rect 2739 7535 2742 7545
rect 2756 7528 2759 7558
rect 2599 7503 2603 7506
rect 2599 7484 2603 7499
rect 2615 7496 2619 7510
rect 2631 7510 2635 7514
rect 2631 7503 2635 7506
rect 2631 7484 2635 7499
rect 2756 7496 2759 7524
rect 2615 7480 2619 7481
rect 2631 7476 2635 7480
rect 2506 7452 2509 7462
rect 2513 7422 2516 7431
rect 2529 7424 2532 7437
rect 2542 7409 2545 7462
rect 2609 7452 2612 7462
rect 2549 7437 2553 7441
rect 2550 7422 2553 7431
rect 2505 7395 2508 7407
rect 2546 7405 2547 7409
rect 2556 7395 2559 7448
rect 2562 7428 2565 7433
rect 2571 7422 2574 7431
rect 2587 7424 2590 7437
rect 2608 7422 2611 7431
rect 2607 7395 2610 7405
rect 2615 7381 2619 7476
rect 2624 7437 2627 7469
rect 2638 7452 2641 7462
rect 2624 7422 2627 7431
rect 2645 7422 2648 7431
rect 2661 7424 2664 7437
rect 2674 7409 2677 7462
rect 2741 7452 2744 7462
rect 2681 7437 2685 7441
rect 2682 7422 2685 7431
rect 2637 7395 2640 7407
rect 2678 7405 2679 7409
rect 2688 7395 2691 7448
rect 2756 7437 2759 7484
rect 2694 7428 2697 7433
rect 2703 7422 2706 7431
rect 2719 7424 2722 7437
rect 2740 7422 2743 7431
rect 2756 7429 2759 7433
rect 2764 7459 2770 7595
rect 2756 7422 2759 7425
rect 2739 7395 2742 7405
rect 2764 7381 2770 7455
rect 2776 9287 2782 9391
rect 2776 9254 2782 9283
rect 2776 9201 2782 9250
rect 2776 9152 2782 9197
rect 2776 9069 2782 9148
rect 2776 8937 2782 9065
rect 2776 8805 2782 8933
rect 2776 8752 2782 8801
rect 2776 8640 2782 8748
rect 2776 8610 2782 8636
rect 2776 8554 2782 8606
rect 2776 8524 2782 8550
rect 2776 8384 2782 8520
rect 2776 8305 2782 8380
rect 2776 8272 2782 8301
rect 2776 8219 2782 8268
rect 2776 8170 2782 8215
rect 2776 8087 2782 8166
rect 2776 7955 2782 8083
rect 2776 7823 2782 7951
rect 2776 7770 2782 7819
rect 2776 7658 2782 7766
rect 2776 7628 2782 7654
rect 2776 7572 2782 7624
rect 2776 7542 2782 7568
rect 2776 7402 2782 7538
rect 2776 7381 2782 7398
rect 2788 9208 2794 9391
rect 2788 9194 2794 9204
rect 2788 9076 2794 9190
rect 2788 9062 2794 9072
rect 2788 8944 2794 9058
rect 2788 8930 2794 8940
rect 2788 8798 2794 8926
rect 2788 8724 2794 8794
rect 2788 8226 2794 8720
rect 2788 8212 2794 8222
rect 2788 8094 2794 8208
rect 2788 8080 2794 8090
rect 2788 7962 2794 8076
rect 2788 7948 2794 7958
rect 2788 7816 2794 7944
rect 2788 7742 2794 7812
rect 2788 7381 2794 7738
rect 2800 9260 2806 9391
rect 2800 9128 2806 9256
rect 2800 9010 2806 9124
rect 2800 8996 2806 9006
rect 2800 8878 2806 8992
rect 2800 8864 2806 8874
rect 2800 8732 2806 8860
rect 2800 8278 2806 8728
rect 2800 8146 2806 8274
rect 2800 8028 2806 8142
rect 2800 8014 2806 8024
rect 2800 7896 2806 8010
rect 2800 7882 2806 7892
rect 2800 7750 2806 7878
rect 2800 7381 2806 7746
rect 2812 9280 2818 9391
rect 2812 9247 2818 9276
rect 2812 9145 2818 9243
rect 2812 8746 2818 9141
rect 2812 8633 2818 8742
rect 2812 8603 2818 8629
rect 2812 8547 2818 8599
rect 2812 8517 2818 8543
rect 2812 8377 2818 8513
rect 2812 8298 2818 8373
rect 2812 8265 2818 8294
rect 2812 8163 2818 8261
rect 2812 7764 2818 8159
rect 2812 7651 2818 7760
rect 2812 7621 2818 7647
rect 2812 7565 2818 7617
rect 2812 7535 2818 7561
rect 2812 7395 2818 7531
rect 2812 7381 2818 7391
rect 2824 9351 2830 9391
rect 2824 9318 2830 9347
rect 2824 9216 2830 9314
rect 2824 8816 2830 9212
rect 2824 8704 2830 8812
rect 2824 8674 2830 8700
rect 2824 8618 2830 8670
rect 2824 8588 2830 8614
rect 2824 8448 2830 8584
rect 2824 8369 2830 8444
rect 2824 8336 2830 8365
rect 2824 8234 2830 8332
rect 2824 7834 2830 8230
rect 2824 7722 2830 7830
rect 2824 7692 2830 7718
rect 2824 7636 2830 7688
rect 2824 7606 2830 7632
rect 2824 7466 2830 7602
rect 2824 7381 2830 7462
rect 2836 8718 2842 9391
rect 2858 9337 2861 9347
rect 2847 9317 2851 9318
rect 2865 9307 2868 9316
rect 2881 9309 2884 9322
rect 2894 9294 2897 9347
rect 2961 9337 2964 9347
rect 2990 9337 2993 9347
rect 2901 9322 2905 9326
rect 2902 9307 2905 9316
rect 2857 9280 2860 9292
rect 2898 9290 2899 9294
rect 2908 9280 2911 9333
rect 2914 9313 2917 9318
rect 2923 9307 2926 9316
rect 2939 9309 2942 9322
rect 2960 9307 2963 9316
rect 2976 9316 2979 9318
rect 2976 9313 2983 9316
rect 2976 9307 2979 9313
rect 2997 9307 3000 9316
rect 3013 9309 3016 9322
rect 2959 9280 2962 9290
rect 2976 9273 2979 9303
rect 3026 9294 3029 9347
rect 3093 9337 3096 9347
rect 3122 9337 3125 9347
rect 3033 9322 3037 9326
rect 3034 9307 3037 9316
rect 2989 9280 2992 9292
rect 3030 9290 3031 9294
rect 3040 9280 3043 9333
rect 3046 9313 3049 9318
rect 3055 9307 3058 9316
rect 3071 9309 3074 9322
rect 3092 9307 3095 9316
rect 3108 9316 3111 9318
rect 3108 9313 3115 9316
rect 3108 9307 3111 9313
rect 3129 9307 3132 9316
rect 3145 9309 3148 9322
rect 3091 9280 3094 9290
rect 2976 9270 3028 9273
rect 2856 9250 2859 9263
rect 2882 9253 2885 9256
rect 2889 9250 2892 9263
rect 2906 9250 2909 9263
rect 2856 9201 2859 9216
rect 2870 9208 2873 9212
rect 2888 9201 2891 9216
rect 2907 9201 2910 9216
rect 2913 9215 2916 9256
rect 2929 9208 2932 9249
rect 2935 9216 2938 9256
rect 2954 9208 2957 9249
rect 2963 9250 2966 9263
rect 2979 9250 2982 9263
rect 3000 9253 3003 9256
rect 3007 9250 3010 9263
rect 3025 9259 3028 9270
rect 3108 9267 3111 9303
rect 3158 9294 3161 9347
rect 3225 9337 3228 9347
rect 3254 9337 3257 9347
rect 3165 9322 3169 9326
rect 3166 9307 3169 9316
rect 3121 9280 3124 9292
rect 3162 9290 3163 9294
rect 3172 9280 3175 9333
rect 3178 9313 3181 9318
rect 3187 9307 3190 9316
rect 3203 9309 3206 9322
rect 3224 9307 3227 9316
rect 3240 9316 3243 9318
rect 3240 9313 3247 9316
rect 3240 9307 3243 9313
rect 3261 9307 3264 9316
rect 3277 9309 3280 9322
rect 3223 9280 3226 9290
rect 3240 9273 3243 9295
rect 3290 9294 3293 9347
rect 3357 9337 3360 9347
rect 3297 9322 3301 9326
rect 3298 9307 3301 9316
rect 3253 9280 3256 9292
rect 3294 9290 3295 9294
rect 3304 9280 3307 9333
rect 3310 9313 3313 9318
rect 3319 9307 3322 9316
rect 3335 9309 3338 9322
rect 3356 9307 3359 9316
rect 3372 9316 3375 9318
rect 3372 9313 3376 9316
rect 3372 9307 3375 9313
rect 3372 9299 3375 9303
rect 3355 9280 3358 9290
rect 3106 9262 3111 9267
rect 3168 9269 3243 9273
rect 3025 9256 3070 9259
rect 3025 9246 3028 9256
rect 3043 9243 3063 9246
rect 3060 9224 3063 9243
rect 2963 9201 2966 9216
rect 2978 9201 2981 9216
rect 2985 9208 2989 9211
rect 3006 9201 3009 9216
rect 2856 9182 2859 9197
rect 2870 9186 2873 9190
rect 2888 9182 2891 9197
rect 2907 9182 2910 9197
rect 2856 9135 2859 9148
rect 2882 9142 2885 9145
rect 2856 9118 2859 9131
rect 2866 9128 2870 9138
rect 2889 9135 2892 9148
rect 2906 9135 2909 9148
rect 2913 9142 2916 9183
rect 2929 9149 2932 9190
rect 2935 9142 2938 9182
rect 2954 9149 2957 9190
rect 2963 9182 2966 9197
rect 2978 9182 2981 9197
rect 2985 9187 2989 9190
rect 3006 9182 3009 9197
rect 2963 9135 2966 9148
rect 2882 9121 2885 9124
rect 2889 9118 2892 9131
rect 2906 9118 2909 9131
rect 2856 9069 2859 9084
rect 2870 9076 2873 9080
rect 2888 9069 2891 9084
rect 2907 9069 2910 9084
rect 2913 9083 2916 9124
rect 2929 9076 2932 9117
rect 2935 9084 2938 9124
rect 2954 9076 2957 9117
rect 2963 9118 2966 9131
rect 2979 9135 2982 9148
rect 3000 9142 3003 9145
rect 3007 9135 3010 9148
rect 3060 9148 3063 9220
rect 3071 9184 3074 9256
rect 3106 9259 3109 9262
rect 3106 9256 3151 9259
rect 3106 9246 3109 9256
rect 2979 9118 2982 9131
rect 3000 9121 3003 9124
rect 3007 9118 3010 9131
rect 3060 9114 3063 9144
rect 3071 9128 3074 9180
rect 3078 9168 3082 9234
rect 3066 9124 3070 9127
rect 3059 9111 3063 9114
rect 3060 9092 3063 9111
rect 2963 9069 2966 9084
rect 2978 9069 2981 9084
rect 2985 9076 2989 9079
rect 3006 9069 3009 9084
rect 2856 9050 2859 9065
rect 2870 9054 2873 9058
rect 2888 9050 2891 9065
rect 2907 9050 2910 9065
rect 2856 9003 2859 9016
rect 2882 9010 2885 9013
rect 2856 8986 2859 8999
rect 2889 9003 2892 9016
rect 2906 9003 2909 9016
rect 2913 9010 2916 9051
rect 2929 9017 2932 9058
rect 2935 9010 2938 9050
rect 2954 9017 2957 9058
rect 2963 9050 2966 9065
rect 2978 9050 2981 9065
rect 2985 9055 2989 9058
rect 3006 9050 3009 9065
rect 2963 9003 2966 9016
rect 2882 8989 2885 8992
rect 2889 8986 2892 8999
rect 2906 8986 2909 8999
rect 2856 8937 2859 8952
rect 2870 8944 2873 8948
rect 2888 8937 2891 8952
rect 2907 8937 2910 8952
rect 2913 8951 2916 8992
rect 2929 8944 2932 8985
rect 2935 8952 2938 8992
rect 2954 8944 2957 8985
rect 2963 8986 2966 8999
rect 2979 9003 2982 9016
rect 3000 9010 3003 9013
rect 3007 9003 3010 9016
rect 3060 9017 3063 9088
rect 3071 9053 3074 9124
rect 2979 8986 2982 8999
rect 3000 8989 3003 8992
rect 3007 8986 3010 8999
rect 3060 8960 3063 9013
rect 3071 8996 3074 9049
rect 3078 9037 3082 9102
rect 3066 8992 3070 8995
rect 3109 8995 3112 9246
rect 3124 9243 3144 9246
rect 3141 9224 3144 9243
rect 3141 9148 3144 9220
rect 3152 9184 3155 9256
rect 3159 9168 3163 9234
rect 3168 9135 3171 9269
rect 3372 9266 3375 9295
rect 3196 9263 3303 9266
rect 3130 9131 3171 9135
rect 3130 9127 3133 9131
rect 3130 9124 3175 9127
rect 3130 9114 3133 9124
rect 3148 9111 3168 9114
rect 3130 9109 3133 9110
rect 3165 9092 3168 9111
rect 3165 9017 3168 9088
rect 3176 9053 3179 9124
rect 3183 9037 3187 9102
rect 2963 8937 2966 8952
rect 2978 8937 2981 8952
rect 2985 8944 2989 8947
rect 3006 8937 3009 8952
rect 2856 8918 2859 8933
rect 2870 8922 2873 8926
rect 2888 8918 2891 8933
rect 2907 8918 2910 8933
rect 2856 8871 2859 8884
rect 2882 8878 2885 8881
rect 2856 8854 2859 8867
rect 2889 8871 2892 8884
rect 2906 8871 2909 8884
rect 2913 8878 2916 8919
rect 2929 8885 2932 8926
rect 2935 8878 2938 8918
rect 2954 8885 2957 8926
rect 2963 8918 2966 8933
rect 2978 8918 2981 8933
rect 2985 8923 2989 8926
rect 3006 8918 3009 8933
rect 2963 8871 2966 8884
rect 2882 8857 2885 8860
rect 2889 8854 2892 8867
rect 2906 8854 2909 8867
rect 2856 8805 2859 8820
rect 2870 8812 2873 8816
rect 2856 8786 2859 8801
rect 2879 8798 2883 8808
rect 2888 8805 2891 8820
rect 2907 8805 2910 8820
rect 2913 8819 2916 8860
rect 2929 8812 2932 8853
rect 2935 8820 2938 8860
rect 2954 8812 2957 8853
rect 2963 8854 2966 8867
rect 2979 8871 2982 8884
rect 3000 8878 3003 8881
rect 3007 8871 3010 8884
rect 3060 8882 3063 8956
rect 3071 8918 3074 8992
rect 3106 8992 3151 8995
rect 3106 8982 3109 8992
rect 3124 8979 3144 8982
rect 2979 8854 2982 8867
rect 3000 8857 3003 8860
rect 3007 8854 3010 8867
rect 3060 8828 3063 8878
rect 3071 8864 3074 8914
rect 3078 8902 3082 8970
rect 3141 8960 3144 8979
rect 3141 8882 3144 8956
rect 3152 8918 3155 8992
rect 3196 8995 3199 9263
rect 3307 9263 3375 9266
rect 3411 9258 3416 9434
rect 3315 9018 3328 9250
rect 3423 9245 3427 9444
rect 3709 9384 3715 9460
rect 3709 9344 3715 9380
rect 3361 9124 3365 9241
rect 3435 9231 3438 9280
rect 3435 9187 3438 9227
rect 3443 9224 3447 9333
rect 3451 9304 3454 9314
rect 3458 9274 3461 9283
rect 3474 9276 3477 9289
rect 3487 9261 3490 9314
rect 3554 9304 3557 9314
rect 3494 9289 3498 9293
rect 3495 9274 3498 9283
rect 3450 9247 3453 9259
rect 3491 9257 3492 9261
rect 3501 9247 3504 9300
rect 3507 9280 3510 9285
rect 3516 9274 3519 9283
rect 3532 9276 3535 9289
rect 3553 9274 3556 9283
rect 3552 9247 3555 9257
rect 3435 9172 3438 9181
rect 3443 9140 3447 9220
rect 3560 9233 3564 9333
rect 3709 9311 3715 9340
rect 3569 9281 3572 9283
rect 3569 9274 3572 9277
rect 3569 9240 3572 9270
rect 3709 9267 3715 9307
rect 3450 9202 3453 9212
rect 3451 9172 3454 9181
rect 3472 9174 3475 9187
rect 3488 9172 3491 9181
rect 3497 9178 3500 9183
rect 3452 9145 3455 9155
rect 3503 9145 3506 9198
rect 3509 9187 3513 9191
rect 3509 9172 3512 9181
rect 3517 9159 3520 9212
rect 3553 9202 3556 9212
rect 3530 9174 3533 9187
rect 3546 9172 3549 9181
rect 3515 9155 3516 9159
rect 3554 9145 3557 9157
rect 3560 9141 3564 9229
rect 3584 9224 3588 9229
rect 3709 9209 3715 9263
rect 3709 9135 3715 9205
rect 3361 9098 3364 9120
rect 3361 9095 3406 9098
rect 3361 9085 3364 9095
rect 3339 9081 3360 9085
rect 3379 9082 3399 9085
rect 3315 9004 3330 9018
rect 3315 9000 3326 9004
rect 3196 8992 3241 8995
rect 3196 8982 3199 8992
rect 3214 8979 3234 8982
rect 3159 8902 3163 8970
rect 3231 8960 3234 8979
rect 3231 8882 3234 8956
rect 3242 8918 3245 8992
rect 3249 8902 3253 8970
rect 3066 8860 3070 8863
rect 2963 8805 2966 8820
rect 2978 8805 2981 8820
rect 2985 8812 2989 8815
rect 3006 8805 3009 8820
rect 2870 8790 2873 8794
rect 2888 8786 2891 8801
rect 2907 8786 2910 8801
rect 2856 8739 2859 8752
rect 2882 8746 2885 8749
rect 2864 8732 2868 8742
rect 2889 8739 2892 8752
rect 2906 8739 2909 8752
rect 2913 8746 2916 8787
rect 2929 8753 2932 8794
rect 2935 8746 2938 8786
rect 2954 8753 2957 8794
rect 2963 8786 2966 8801
rect 2978 8786 2981 8801
rect 2985 8791 2989 8794
rect 3006 8786 3009 8801
rect 2963 8739 2966 8752
rect 2979 8739 2982 8752
rect 3000 8746 3003 8749
rect 3007 8739 3010 8752
rect 3060 8746 3063 8824
rect 3071 8782 3074 8860
rect 3078 8766 3082 8838
rect 3090 8739 3094 8752
rect 3099 8732 3102 8742
rect 3109 8725 3112 8794
rect 3131 8790 3134 8794
rect 3149 8786 3152 8801
rect 3168 8786 3171 8801
rect 3116 8739 3120 8752
rect 3143 8746 3146 8749
rect 3150 8739 3153 8752
rect 3167 8739 3170 8752
rect 3174 8746 3177 8787
rect 3190 8753 3193 8794
rect 3196 8746 3199 8786
rect 3215 8753 3218 8794
rect 3224 8786 3227 8801
rect 3239 8786 3242 8801
rect 3246 8791 3250 8794
rect 3267 8786 3270 8801
rect 3224 8739 3227 8752
rect 3240 8739 3243 8752
rect 3261 8746 3264 8749
rect 3268 8739 3271 8752
rect 3284 8733 3288 8969
rect 3326 8874 3330 9000
rect 3339 8955 3342 9081
rect 3361 9076 3364 9081
rect 3361 9073 3383 9076
rect 3396 9063 3399 9082
rect 3396 8983 3399 9059
rect 3407 9019 3410 9095
rect 3414 9003 3418 9073
rect 3593 9012 3597 9053
rect 3660 9026 3665 9065
rect 3361 8965 3406 8968
rect 3361 8955 3364 8965
rect 3379 8952 3399 8955
rect 3339 8946 3342 8951
rect 3339 8943 3383 8946
rect 3396 8933 3399 8952
rect 3326 8870 3328 8874
rect 3396 8853 3399 8929
rect 3407 8889 3410 8965
rect 3414 8873 3418 8943
rect 3488 8886 3492 8923
rect 3660 8896 3665 9022
rect 3660 8833 3665 8892
rect 3668 9037 3672 9102
rect 3668 8976 3672 9033
rect 3668 8846 3672 8972
rect 3668 8833 3672 8842
rect 3676 9021 3680 9065
rect 3676 8833 3680 9017
rect 3709 9037 3715 9131
rect 3709 9003 3715 9033
rect 3709 8871 3715 8999
rect 3443 8824 3447 8825
rect 3560 8823 3564 8824
rect 3319 8802 3322 8812
rect 3326 8772 3329 8781
rect 3342 8774 3345 8787
rect 3355 8759 3358 8812
rect 3422 8802 3425 8812
rect 3362 8787 3366 8791
rect 3363 8772 3366 8781
rect 3318 8745 3321 8757
rect 3359 8755 3360 8759
rect 3369 8745 3372 8798
rect 3375 8778 3378 8783
rect 3384 8772 3387 8781
rect 3400 8774 3403 8787
rect 3421 8772 3424 8781
rect 3437 8772 3440 8781
rect 3420 8745 3423 8755
rect 3277 8721 3278 8724
rect 2836 7736 2842 8714
rect 3142 8611 3146 8693
rect 3157 8690 3160 8700
rect 3164 8660 3167 8669
rect 3180 8662 3183 8675
rect 3193 8647 3196 8700
rect 3260 8690 3263 8700
rect 3200 8675 3204 8679
rect 3201 8660 3204 8669
rect 3156 8633 3159 8645
rect 3197 8643 3198 8647
rect 3207 8633 3210 8686
rect 3275 8675 3278 8721
rect 3213 8666 3216 8671
rect 3222 8660 3225 8669
rect 3238 8662 3241 8675
rect 3259 8660 3262 8669
rect 3275 8660 3278 8669
rect 3258 8633 3261 8643
rect 3275 8626 3278 8656
rect 3150 8584 3153 8621
rect 3157 8604 3160 8614
rect 3164 8574 3167 8583
rect 3180 8576 3183 8589
rect 3193 8561 3196 8614
rect 3260 8604 3263 8614
rect 3200 8589 3204 8593
rect 3201 8574 3204 8583
rect 3156 8547 3159 8559
rect 3197 8557 3198 8561
rect 3207 8547 3210 8600
rect 3213 8580 3216 8585
rect 3222 8574 3225 8583
rect 3238 8576 3241 8589
rect 3259 8574 3262 8583
rect 3275 8584 3278 8585
rect 3296 8587 3300 8729
rect 3312 8640 3315 8734
rect 3437 8731 3440 8768
rect 3443 8724 3447 8819
rect 3451 8802 3454 8812
rect 3458 8772 3461 8781
rect 3474 8774 3477 8787
rect 3487 8759 3490 8812
rect 3554 8802 3557 8812
rect 3494 8787 3498 8791
rect 3495 8772 3498 8781
rect 3450 8745 3453 8757
rect 3491 8755 3492 8759
rect 3501 8745 3504 8798
rect 3507 8778 3510 8783
rect 3516 8772 3519 8781
rect 3532 8774 3535 8787
rect 3553 8772 3556 8781
rect 3552 8745 3555 8755
rect 3427 8711 3431 8715
rect 3427 8692 3431 8707
rect 3443 8704 3447 8720
rect 3459 8719 3463 8724
rect 3459 8711 3463 8715
rect 3459 8692 3463 8707
rect 3443 8688 3447 8689
rect 3459 8684 3463 8688
rect 3319 8660 3322 8670
rect 3326 8630 3329 8639
rect 3342 8632 3345 8645
rect 3355 8617 3358 8670
rect 3422 8660 3425 8670
rect 3362 8645 3366 8649
rect 3363 8630 3366 8639
rect 3318 8603 3321 8615
rect 3359 8613 3360 8617
rect 3369 8603 3372 8656
rect 3437 8645 3440 8677
rect 3375 8636 3378 8641
rect 3384 8630 3387 8639
rect 3400 8632 3403 8645
rect 3421 8630 3424 8639
rect 3437 8630 3440 8639
rect 3420 8603 3423 8613
rect 3275 8579 3278 8580
rect 3258 8547 3261 8557
rect 3296 8485 3300 8567
rect 3312 8554 3315 8592
rect 3319 8574 3322 8584
rect 3326 8544 3329 8553
rect 3342 8546 3345 8559
rect 3355 8531 3358 8584
rect 3422 8574 3425 8584
rect 3362 8559 3366 8563
rect 3363 8544 3366 8553
rect 3318 8517 3321 8529
rect 3359 8527 3360 8531
rect 3369 8517 3372 8570
rect 3375 8550 3378 8555
rect 3384 8544 3387 8553
rect 3400 8546 3403 8559
rect 3421 8544 3424 8553
rect 3437 8544 3440 8553
rect 3420 8517 3423 8527
rect 3312 8414 3315 8506
rect 3437 8503 3440 8540
rect 3319 8434 3322 8444
rect 3326 8404 3329 8413
rect 3342 8406 3345 8419
rect 3355 8391 3358 8444
rect 3422 8434 3425 8444
rect 3362 8419 3366 8423
rect 3363 8404 3366 8413
rect 3318 8377 3321 8389
rect 3359 8387 3360 8391
rect 3369 8377 3372 8430
rect 3437 8419 3440 8451
rect 3375 8410 3378 8415
rect 3384 8404 3387 8413
rect 3400 8406 3403 8419
rect 3421 8404 3424 8413
rect 3437 8404 3440 8413
rect 3420 8377 3423 8387
rect 2858 8355 2861 8365
rect 2865 8325 2868 8334
rect 2881 8327 2884 8340
rect 2894 8312 2897 8365
rect 2961 8355 2964 8365
rect 2990 8355 2993 8365
rect 2901 8340 2905 8344
rect 2902 8325 2905 8334
rect 2857 8298 2860 8310
rect 2898 8308 2899 8312
rect 2908 8298 2911 8351
rect 2914 8331 2917 8336
rect 2923 8325 2926 8334
rect 2939 8327 2942 8340
rect 2960 8325 2963 8334
rect 2976 8334 2979 8336
rect 2976 8331 2983 8334
rect 2976 8325 2979 8331
rect 2997 8325 3000 8334
rect 3013 8327 3016 8340
rect 2959 8298 2962 8308
rect 2976 8291 2979 8321
rect 3026 8312 3029 8365
rect 3093 8355 3096 8365
rect 3122 8355 3125 8365
rect 3033 8340 3037 8344
rect 3034 8325 3037 8334
rect 2989 8298 2992 8310
rect 3030 8308 3031 8312
rect 3040 8298 3043 8351
rect 3046 8331 3049 8336
rect 3055 8325 3058 8334
rect 3071 8327 3074 8340
rect 3092 8325 3095 8334
rect 3108 8334 3111 8336
rect 3108 8331 3115 8334
rect 3108 8325 3111 8331
rect 3129 8325 3132 8334
rect 3145 8327 3148 8340
rect 3091 8298 3094 8308
rect 2976 8288 3028 8291
rect 2856 8268 2859 8281
rect 2882 8271 2885 8274
rect 2889 8268 2892 8281
rect 2906 8268 2909 8281
rect 2856 8219 2859 8234
rect 2870 8226 2873 8230
rect 2888 8219 2891 8234
rect 2907 8219 2910 8234
rect 2913 8233 2916 8274
rect 2929 8226 2932 8267
rect 2935 8234 2938 8274
rect 2954 8226 2957 8267
rect 2963 8268 2966 8281
rect 2979 8268 2982 8281
rect 3000 8271 3003 8274
rect 3007 8268 3010 8281
rect 3025 8277 3028 8288
rect 3108 8285 3111 8321
rect 3158 8312 3161 8365
rect 3225 8355 3228 8365
rect 3254 8355 3257 8365
rect 3165 8340 3169 8344
rect 3166 8325 3169 8334
rect 3121 8298 3124 8310
rect 3162 8308 3163 8312
rect 3172 8298 3175 8351
rect 3178 8331 3181 8336
rect 3187 8325 3190 8334
rect 3203 8327 3206 8340
rect 3224 8325 3227 8334
rect 3240 8334 3243 8336
rect 3240 8331 3247 8334
rect 3240 8325 3243 8331
rect 3261 8325 3264 8334
rect 3277 8327 3280 8340
rect 3223 8298 3226 8308
rect 3240 8291 3243 8313
rect 3290 8312 3293 8365
rect 3357 8355 3360 8365
rect 3297 8340 3301 8344
rect 3298 8325 3301 8334
rect 3253 8298 3256 8310
rect 3294 8308 3295 8312
rect 3304 8298 3307 8351
rect 3310 8331 3313 8336
rect 3319 8325 3322 8334
rect 3335 8327 3338 8340
rect 3356 8325 3359 8334
rect 3372 8334 3375 8336
rect 3372 8331 3376 8334
rect 3372 8325 3375 8331
rect 3372 8317 3375 8321
rect 3355 8298 3358 8308
rect 3106 8280 3111 8285
rect 3168 8287 3243 8291
rect 3025 8274 3070 8277
rect 3025 8264 3028 8274
rect 3043 8261 3063 8264
rect 3060 8242 3063 8261
rect 2963 8219 2966 8234
rect 2978 8219 2981 8234
rect 2985 8226 2989 8229
rect 3006 8219 3009 8234
rect 2856 8200 2859 8215
rect 2870 8204 2873 8208
rect 2888 8200 2891 8215
rect 2907 8200 2910 8215
rect 2856 8153 2859 8166
rect 2882 8160 2885 8163
rect 2856 8136 2859 8149
rect 2866 8146 2870 8156
rect 2889 8153 2892 8166
rect 2906 8153 2909 8166
rect 2913 8160 2916 8201
rect 2929 8167 2932 8208
rect 2935 8160 2938 8200
rect 2954 8167 2957 8208
rect 2963 8200 2966 8215
rect 2978 8200 2981 8215
rect 2985 8205 2989 8208
rect 3006 8200 3009 8215
rect 2963 8153 2966 8166
rect 2882 8139 2885 8142
rect 2889 8136 2892 8149
rect 2906 8136 2909 8149
rect 2856 8087 2859 8102
rect 2870 8094 2873 8098
rect 2888 8087 2891 8102
rect 2907 8087 2910 8102
rect 2913 8101 2916 8142
rect 2929 8094 2932 8135
rect 2935 8102 2938 8142
rect 2954 8094 2957 8135
rect 2963 8136 2966 8149
rect 2979 8153 2982 8166
rect 3000 8160 3003 8163
rect 3007 8153 3010 8166
rect 3060 8166 3063 8238
rect 3071 8202 3074 8274
rect 3106 8277 3109 8280
rect 3106 8274 3151 8277
rect 3106 8264 3109 8274
rect 2979 8136 2982 8149
rect 3000 8139 3003 8142
rect 3007 8136 3010 8149
rect 3060 8132 3063 8162
rect 3071 8146 3074 8198
rect 3078 8186 3082 8252
rect 3066 8142 3070 8145
rect 3059 8129 3063 8132
rect 3060 8110 3063 8129
rect 2963 8087 2966 8102
rect 2978 8087 2981 8102
rect 2985 8094 2989 8097
rect 3006 8087 3009 8102
rect 2856 8068 2859 8083
rect 2870 8072 2873 8076
rect 2888 8068 2891 8083
rect 2907 8068 2910 8083
rect 2856 8021 2859 8034
rect 2882 8028 2885 8031
rect 2856 8004 2859 8017
rect 2889 8021 2892 8034
rect 2906 8021 2909 8034
rect 2913 8028 2916 8069
rect 2929 8035 2932 8076
rect 2935 8028 2938 8068
rect 2954 8035 2957 8076
rect 2963 8068 2966 8083
rect 2978 8068 2981 8083
rect 2985 8073 2989 8076
rect 3006 8068 3009 8083
rect 2963 8021 2966 8034
rect 2882 8007 2885 8010
rect 2889 8004 2892 8017
rect 2906 8004 2909 8017
rect 2856 7955 2859 7970
rect 2870 7962 2873 7966
rect 2888 7955 2891 7970
rect 2907 7955 2910 7970
rect 2913 7969 2916 8010
rect 2929 7962 2932 8003
rect 2935 7970 2938 8010
rect 2954 7962 2957 8003
rect 2963 8004 2966 8017
rect 2979 8021 2982 8034
rect 3000 8028 3003 8031
rect 3007 8021 3010 8034
rect 3060 8035 3063 8106
rect 3071 8071 3074 8142
rect 2979 8004 2982 8017
rect 3000 8007 3003 8010
rect 3007 8004 3010 8017
rect 3060 7978 3063 8031
rect 3071 8014 3074 8067
rect 3078 8055 3082 8120
rect 3066 8010 3070 8013
rect 3109 8013 3112 8264
rect 3124 8261 3144 8264
rect 3141 8242 3144 8261
rect 3141 8166 3144 8238
rect 3152 8202 3155 8274
rect 3159 8186 3163 8252
rect 3168 8153 3171 8287
rect 3372 8284 3375 8313
rect 3196 8281 3303 8284
rect 3130 8149 3171 8153
rect 3130 8145 3133 8149
rect 3130 8142 3175 8145
rect 3130 8132 3133 8142
rect 3148 8129 3168 8132
rect 3130 8127 3133 8128
rect 3165 8110 3168 8129
rect 3165 8035 3168 8106
rect 3176 8071 3179 8142
rect 3183 8055 3187 8120
rect 2963 7955 2966 7970
rect 2978 7955 2981 7970
rect 2985 7962 2989 7965
rect 3006 7955 3009 7970
rect 2856 7936 2859 7951
rect 2870 7940 2873 7944
rect 2888 7936 2891 7951
rect 2907 7936 2910 7951
rect 2856 7889 2859 7902
rect 2882 7896 2885 7899
rect 2856 7872 2859 7885
rect 2889 7889 2892 7902
rect 2906 7889 2909 7902
rect 2913 7896 2916 7937
rect 2929 7903 2932 7944
rect 2935 7896 2938 7936
rect 2954 7903 2957 7944
rect 2963 7936 2966 7951
rect 2978 7936 2981 7951
rect 2985 7941 2989 7944
rect 3006 7936 3009 7951
rect 2963 7889 2966 7902
rect 2882 7875 2885 7878
rect 2889 7872 2892 7885
rect 2906 7872 2909 7885
rect 2856 7823 2859 7838
rect 2870 7830 2873 7834
rect 2856 7804 2859 7819
rect 2879 7816 2883 7826
rect 2888 7823 2891 7838
rect 2907 7823 2910 7838
rect 2913 7837 2916 7878
rect 2929 7830 2932 7871
rect 2935 7838 2938 7878
rect 2954 7830 2957 7871
rect 2963 7872 2966 7885
rect 2979 7889 2982 7902
rect 3000 7896 3003 7899
rect 3007 7889 3010 7902
rect 3060 7900 3063 7974
rect 3071 7936 3074 8010
rect 3106 8010 3151 8013
rect 3106 8000 3109 8010
rect 3124 7997 3144 8000
rect 2979 7872 2982 7885
rect 3000 7875 3003 7878
rect 3007 7872 3010 7885
rect 3060 7846 3063 7896
rect 3071 7882 3074 7932
rect 3078 7920 3082 7988
rect 3141 7978 3144 7997
rect 3141 7900 3144 7974
rect 3152 7936 3155 8010
rect 3196 8013 3199 8281
rect 3307 8281 3375 8284
rect 3435 8249 3438 8298
rect 3435 8205 3438 8245
rect 3443 8242 3447 8684
rect 3451 8660 3454 8670
rect 3458 8630 3461 8639
rect 3474 8632 3477 8645
rect 3487 8617 3490 8670
rect 3554 8660 3557 8670
rect 3494 8645 3498 8649
rect 3495 8630 3498 8639
rect 3450 8603 3453 8615
rect 3491 8613 3492 8617
rect 3501 8603 3504 8656
rect 3507 8636 3510 8641
rect 3516 8630 3519 8639
rect 3532 8632 3535 8645
rect 3553 8630 3556 8639
rect 3552 8603 3555 8613
rect 3451 8574 3454 8584
rect 3458 8544 3461 8553
rect 3474 8546 3477 8559
rect 3487 8531 3490 8584
rect 3554 8574 3557 8584
rect 3494 8559 3498 8563
rect 3495 8544 3498 8553
rect 3450 8517 3453 8529
rect 3491 8527 3492 8531
rect 3501 8517 3504 8570
rect 3507 8550 3510 8555
rect 3516 8544 3519 8553
rect 3532 8546 3535 8559
rect 3553 8544 3556 8553
rect 3552 8517 3555 8527
rect 3560 8496 3564 8818
rect 3583 8802 3586 8812
rect 3569 8772 3572 8781
rect 3590 8772 3593 8781
rect 3606 8774 3609 8787
rect 3569 8731 3572 8768
rect 3619 8759 3622 8812
rect 3686 8802 3689 8812
rect 3709 8809 3715 8867
rect 3626 8787 3630 8791
rect 3627 8772 3630 8781
rect 3582 8745 3585 8757
rect 3623 8755 3624 8759
rect 3633 8745 3636 8798
rect 3639 8778 3642 8783
rect 3648 8772 3651 8781
rect 3664 8774 3667 8787
rect 3685 8772 3688 8781
rect 3701 8772 3704 8783
rect 3684 8745 3687 8755
rect 3701 8738 3704 8768
rect 3701 8704 3704 8734
rect 3709 8739 3715 8805
rect 3709 8697 3715 8735
rect 3569 8645 3572 8677
rect 3583 8660 3586 8670
rect 3569 8630 3572 8639
rect 3590 8630 3593 8639
rect 3606 8632 3609 8645
rect 3619 8617 3622 8670
rect 3686 8660 3689 8670
rect 3626 8645 3630 8649
rect 3627 8630 3630 8639
rect 3582 8603 3585 8615
rect 3623 8613 3624 8617
rect 3633 8603 3636 8656
rect 3701 8645 3704 8692
rect 3639 8636 3642 8641
rect 3648 8630 3651 8639
rect 3664 8632 3667 8645
rect 3685 8630 3688 8639
rect 3701 8630 3704 8641
rect 3684 8603 3687 8613
rect 3701 8596 3704 8626
rect 3709 8667 3715 8693
rect 3583 8574 3586 8584
rect 3569 8544 3572 8553
rect 3590 8544 3593 8553
rect 3606 8546 3609 8559
rect 3569 8503 3572 8540
rect 3619 8531 3622 8584
rect 3686 8574 3689 8584
rect 3709 8581 3715 8663
rect 3626 8559 3630 8563
rect 3627 8544 3630 8553
rect 3582 8517 3585 8529
rect 3623 8527 3624 8531
rect 3633 8517 3636 8570
rect 3639 8550 3642 8555
rect 3648 8544 3651 8553
rect 3664 8546 3667 8559
rect 3685 8544 3688 8553
rect 3701 8544 3704 8555
rect 3684 8517 3687 8527
rect 3701 8510 3704 8540
rect 3544 8485 3548 8488
rect 3544 8466 3548 8481
rect 3560 8478 3564 8492
rect 3576 8492 3580 8496
rect 3576 8485 3580 8488
rect 3576 8466 3580 8481
rect 3701 8478 3704 8506
rect 3560 8462 3564 8463
rect 3576 8458 3580 8462
rect 3451 8434 3454 8444
rect 3458 8404 3461 8413
rect 3474 8406 3477 8419
rect 3487 8391 3490 8444
rect 3554 8434 3557 8444
rect 3494 8419 3498 8423
rect 3495 8404 3498 8413
rect 3450 8377 3453 8389
rect 3491 8387 3492 8391
rect 3501 8377 3504 8430
rect 3507 8410 3510 8415
rect 3516 8404 3519 8413
rect 3532 8406 3535 8419
rect 3553 8404 3556 8413
rect 3552 8377 3555 8387
rect 3451 8322 3454 8332
rect 3458 8292 3461 8301
rect 3474 8294 3477 8307
rect 3487 8279 3490 8332
rect 3554 8322 3557 8332
rect 3494 8307 3498 8311
rect 3495 8292 3498 8301
rect 3450 8265 3453 8277
rect 3491 8275 3492 8279
rect 3501 8265 3504 8318
rect 3507 8298 3510 8303
rect 3516 8292 3519 8301
rect 3532 8294 3535 8307
rect 3553 8292 3556 8301
rect 3552 8265 3555 8275
rect 3435 8190 3438 8199
rect 3196 8010 3241 8013
rect 3196 8000 3199 8010
rect 3214 7997 3234 8000
rect 3159 7920 3163 7988
rect 3231 7978 3234 7997
rect 3231 7900 3234 7974
rect 3242 7936 3245 8010
rect 3249 7920 3253 7988
rect 3066 7878 3070 7881
rect 2963 7823 2966 7838
rect 2978 7823 2981 7838
rect 2985 7830 2989 7833
rect 3006 7823 3009 7838
rect 2870 7808 2873 7812
rect 2888 7804 2891 7819
rect 2907 7804 2910 7819
rect 2856 7757 2859 7770
rect 2882 7764 2885 7767
rect 2864 7750 2868 7760
rect 2889 7757 2892 7770
rect 2906 7757 2909 7770
rect 2913 7764 2916 7805
rect 2929 7771 2932 7812
rect 2935 7764 2938 7804
rect 2954 7771 2957 7812
rect 2963 7804 2966 7819
rect 2978 7804 2981 7819
rect 2985 7809 2989 7812
rect 3006 7804 3009 7819
rect 2963 7757 2966 7770
rect 2979 7757 2982 7770
rect 3000 7764 3003 7767
rect 3007 7757 3010 7770
rect 3060 7764 3063 7842
rect 3071 7800 3074 7878
rect 3078 7784 3082 7856
rect 3090 7757 3094 7770
rect 3099 7750 3102 7760
rect 3109 7743 3112 7812
rect 3131 7808 3134 7812
rect 3149 7804 3152 7819
rect 3168 7804 3171 7819
rect 3116 7757 3120 7770
rect 3143 7764 3146 7767
rect 3150 7757 3153 7770
rect 3167 7757 3170 7770
rect 3174 7764 3177 7805
rect 3190 7771 3193 7812
rect 3196 7764 3199 7804
rect 3215 7771 3218 7812
rect 3224 7804 3227 7819
rect 3239 7804 3242 7819
rect 3246 7809 3250 7812
rect 3267 7804 3270 7819
rect 3224 7757 3227 7770
rect 3240 7757 3243 7770
rect 3261 7764 3264 7767
rect 3268 7757 3271 7770
rect 3284 7751 3288 7987
rect 3319 7820 3322 7830
rect 3326 7790 3329 7799
rect 3342 7792 3345 7805
rect 3355 7777 3358 7830
rect 3422 7820 3425 7830
rect 3362 7805 3366 7809
rect 3363 7790 3366 7799
rect 3318 7763 3321 7775
rect 3359 7773 3360 7777
rect 3369 7763 3372 7816
rect 3375 7796 3378 7801
rect 3384 7790 3387 7799
rect 3400 7792 3403 7805
rect 3421 7790 3424 7799
rect 3437 7790 3440 7799
rect 3420 7763 3423 7773
rect 3277 7739 3278 7742
rect 2836 7381 2842 7732
rect 3142 7629 3146 7711
rect 3157 7708 3160 7718
rect 3164 7678 3167 7687
rect 3180 7680 3183 7693
rect 3193 7665 3196 7718
rect 3260 7708 3263 7718
rect 3200 7693 3204 7697
rect 3201 7678 3204 7687
rect 3156 7651 3159 7663
rect 3197 7661 3198 7665
rect 3207 7651 3210 7704
rect 3275 7693 3278 7739
rect 3213 7684 3216 7689
rect 3222 7678 3225 7687
rect 3238 7680 3241 7693
rect 3259 7678 3262 7687
rect 3275 7678 3278 7687
rect 3258 7651 3261 7661
rect 3275 7644 3278 7674
rect 3150 7602 3153 7639
rect 3157 7622 3160 7632
rect 3164 7592 3167 7601
rect 3180 7594 3183 7607
rect 3193 7579 3196 7632
rect 3260 7622 3263 7632
rect 3200 7607 3204 7611
rect 3201 7592 3204 7601
rect 3156 7565 3159 7577
rect 3197 7575 3198 7579
rect 3207 7565 3210 7618
rect 3213 7598 3216 7603
rect 3222 7592 3225 7601
rect 3238 7594 3241 7607
rect 3259 7592 3262 7601
rect 3275 7602 3278 7603
rect 3296 7605 3300 7747
rect 3312 7658 3315 7752
rect 3437 7749 3440 7786
rect 3443 7742 3447 8238
rect 3560 8251 3564 8458
rect 3569 8419 3572 8451
rect 3583 8434 3586 8444
rect 3569 8404 3572 8413
rect 3590 8404 3593 8413
rect 3606 8406 3609 8419
rect 3619 8391 3622 8444
rect 3686 8434 3689 8444
rect 3626 8419 3630 8423
rect 3627 8404 3630 8413
rect 3582 8377 3585 8389
rect 3623 8387 3624 8391
rect 3633 8377 3636 8430
rect 3701 8419 3704 8466
rect 3639 8410 3642 8415
rect 3648 8404 3651 8413
rect 3664 8406 3667 8419
rect 3685 8404 3688 8413
rect 3701 8411 3704 8415
rect 3709 8441 3715 8577
rect 3701 8404 3704 8407
rect 3684 8377 3687 8387
rect 3709 8362 3715 8437
rect 3709 8329 3715 8358
rect 3569 8300 3572 8301
rect 3569 8295 3573 8296
rect 3569 8292 3572 8295
rect 3569 8258 3572 8288
rect 3709 8285 3715 8325
rect 3450 8220 3453 8230
rect 3451 8190 3454 8199
rect 3472 8192 3475 8205
rect 3488 8190 3491 8199
rect 3497 8196 3500 8201
rect 3452 8163 3455 8173
rect 3503 8163 3506 8216
rect 3509 8205 3513 8209
rect 3509 8190 3512 8199
rect 3517 8177 3520 8230
rect 3553 8220 3556 8230
rect 3530 8192 3533 8205
rect 3546 8190 3549 8199
rect 3515 8173 3516 8177
rect 3554 8163 3557 8175
rect 3451 7820 3454 7830
rect 3458 7790 3461 7799
rect 3474 7792 3477 7805
rect 3487 7777 3490 7830
rect 3554 7820 3557 7830
rect 3494 7805 3498 7809
rect 3495 7790 3498 7799
rect 3450 7763 3453 7775
rect 3491 7773 3492 7777
rect 3501 7763 3504 7816
rect 3507 7796 3510 7801
rect 3516 7790 3519 7799
rect 3532 7792 3535 7805
rect 3553 7790 3556 7799
rect 3552 7763 3555 7773
rect 3427 7729 3431 7734
rect 3427 7710 3431 7725
rect 3443 7722 3447 7738
rect 3459 7738 3463 7742
rect 3459 7729 3463 7734
rect 3459 7710 3463 7725
rect 3443 7706 3447 7707
rect 3459 7702 3463 7706
rect 3319 7678 3322 7688
rect 3326 7648 3329 7657
rect 3342 7650 3345 7663
rect 3355 7635 3358 7688
rect 3422 7678 3425 7688
rect 3362 7663 3366 7667
rect 3363 7648 3366 7657
rect 3318 7621 3321 7633
rect 3359 7631 3360 7635
rect 3369 7621 3372 7674
rect 3437 7663 3440 7695
rect 3375 7654 3378 7659
rect 3384 7648 3387 7657
rect 3400 7650 3403 7663
rect 3421 7648 3424 7657
rect 3437 7648 3440 7657
rect 3420 7621 3423 7631
rect 3275 7597 3278 7598
rect 3258 7565 3261 7575
rect 3296 7503 3300 7585
rect 3312 7572 3315 7610
rect 3319 7592 3322 7602
rect 3326 7562 3329 7571
rect 3342 7564 3345 7577
rect 3355 7549 3358 7602
rect 3422 7592 3425 7602
rect 3362 7577 3366 7581
rect 3363 7562 3366 7571
rect 3318 7535 3321 7547
rect 3359 7545 3360 7549
rect 3369 7535 3372 7588
rect 3375 7568 3378 7573
rect 3384 7562 3387 7571
rect 3400 7564 3403 7577
rect 3421 7562 3424 7571
rect 3437 7562 3440 7571
rect 3420 7535 3423 7545
rect 3312 7432 3315 7524
rect 3437 7521 3440 7558
rect 3319 7452 3322 7462
rect 3326 7422 3329 7431
rect 3342 7424 3345 7437
rect 3355 7409 3358 7462
rect 3422 7452 3425 7462
rect 3362 7437 3366 7441
rect 3363 7422 3366 7431
rect 3318 7395 3321 7407
rect 3359 7405 3360 7409
rect 3369 7395 3372 7448
rect 3437 7437 3440 7469
rect 3375 7428 3378 7433
rect 3384 7422 3387 7431
rect 3400 7424 3403 7437
rect 3421 7422 3424 7431
rect 3437 7422 3440 7431
rect 3420 7395 3423 7405
rect 3443 7381 3447 7702
rect 3451 7678 3454 7688
rect 3458 7648 3461 7657
rect 3474 7650 3477 7663
rect 3487 7635 3490 7688
rect 3554 7678 3557 7688
rect 3494 7663 3498 7667
rect 3495 7648 3498 7657
rect 3450 7621 3453 7633
rect 3491 7631 3492 7635
rect 3501 7621 3504 7674
rect 3507 7654 3510 7659
rect 3516 7648 3519 7657
rect 3532 7650 3535 7663
rect 3553 7648 3556 7657
rect 3552 7621 3555 7631
rect 3451 7592 3454 7602
rect 3458 7562 3461 7571
rect 3474 7564 3477 7577
rect 3487 7549 3490 7602
rect 3554 7592 3557 7602
rect 3494 7577 3498 7581
rect 3495 7562 3498 7571
rect 3450 7535 3453 7547
rect 3491 7545 3492 7549
rect 3501 7535 3504 7588
rect 3507 7568 3510 7573
rect 3516 7562 3519 7571
rect 3532 7564 3535 7577
rect 3553 7562 3556 7571
rect 3552 7535 3555 7545
rect 3560 7514 3564 8247
rect 3584 8242 3588 8247
rect 3709 8227 3715 8281
rect 3709 8153 3715 8223
rect 3709 8021 3715 8149
rect 3709 7889 3715 8017
rect 3583 7820 3586 7830
rect 3569 7790 3572 7799
rect 3590 7790 3593 7799
rect 3606 7792 3609 7805
rect 3569 7749 3572 7786
rect 3619 7777 3622 7830
rect 3686 7820 3689 7830
rect 3709 7827 3715 7885
rect 3626 7805 3630 7809
rect 3627 7790 3630 7799
rect 3582 7763 3585 7775
rect 3623 7773 3624 7777
rect 3633 7763 3636 7816
rect 3639 7796 3642 7801
rect 3648 7790 3651 7799
rect 3664 7792 3667 7805
rect 3685 7790 3688 7799
rect 3701 7790 3704 7801
rect 3684 7763 3687 7773
rect 3701 7756 3704 7786
rect 3701 7722 3704 7752
rect 3709 7757 3715 7823
rect 3709 7715 3715 7753
rect 3569 7663 3572 7695
rect 3583 7678 3586 7688
rect 3569 7648 3572 7657
rect 3590 7648 3593 7657
rect 3606 7650 3609 7663
rect 3619 7635 3622 7688
rect 3686 7678 3689 7688
rect 3626 7663 3630 7667
rect 3627 7648 3630 7657
rect 3582 7621 3585 7633
rect 3623 7631 3624 7635
rect 3633 7621 3636 7674
rect 3701 7663 3704 7710
rect 3639 7654 3642 7659
rect 3648 7648 3651 7657
rect 3664 7650 3667 7663
rect 3685 7648 3688 7657
rect 3701 7648 3704 7659
rect 3684 7621 3687 7631
rect 3701 7614 3704 7644
rect 3709 7685 3715 7711
rect 3583 7592 3586 7602
rect 3569 7562 3572 7571
rect 3590 7562 3593 7571
rect 3606 7564 3609 7577
rect 3569 7521 3572 7558
rect 3619 7549 3622 7602
rect 3686 7592 3689 7602
rect 3709 7599 3715 7681
rect 3626 7577 3630 7581
rect 3627 7562 3630 7571
rect 3582 7535 3585 7547
rect 3623 7545 3624 7549
rect 3633 7535 3636 7588
rect 3639 7568 3642 7573
rect 3648 7562 3651 7571
rect 3664 7564 3667 7577
rect 3685 7562 3688 7571
rect 3701 7562 3704 7573
rect 3684 7535 3687 7545
rect 3701 7528 3704 7558
rect 3544 7503 3548 7506
rect 3544 7484 3548 7499
rect 3560 7496 3564 7510
rect 3576 7510 3580 7514
rect 3576 7503 3580 7506
rect 3576 7484 3580 7499
rect 3701 7496 3704 7524
rect 3560 7480 3564 7481
rect 3576 7476 3580 7480
rect 3451 7452 3454 7462
rect 3458 7422 3461 7431
rect 3474 7424 3477 7437
rect 3487 7409 3490 7462
rect 3554 7452 3557 7462
rect 3494 7437 3498 7441
rect 3495 7422 3498 7431
rect 3450 7395 3453 7407
rect 3491 7405 3492 7409
rect 3501 7395 3504 7448
rect 3507 7428 3510 7433
rect 3516 7422 3519 7431
rect 3532 7424 3535 7437
rect 3553 7422 3556 7431
rect 3552 7395 3555 7405
rect 3560 7381 3564 7476
rect 3569 7437 3572 7469
rect 3583 7452 3586 7462
rect 3569 7422 3572 7431
rect 3590 7422 3593 7431
rect 3606 7424 3609 7437
rect 3619 7409 3622 7462
rect 3686 7452 3689 7462
rect 3626 7437 3630 7441
rect 3627 7422 3630 7431
rect 3582 7395 3585 7407
rect 3623 7405 3624 7409
rect 3633 7395 3636 7448
rect 3701 7437 3704 7484
rect 3639 7428 3642 7433
rect 3648 7422 3651 7431
rect 3664 7424 3667 7437
rect 3685 7422 3688 7431
rect 3701 7429 3704 7433
rect 3709 7459 3715 7595
rect 3701 7422 3704 7425
rect 3684 7395 3687 7405
rect 3709 7381 3715 7455
rect 3721 9392 3727 9467
rect 3721 9287 3727 9388
rect 3721 9254 3727 9283
rect 3721 9201 3727 9250
rect 3721 9152 3727 9197
rect 3721 9069 3727 9148
rect 3721 9030 3727 9065
rect 3721 8937 3727 9026
rect 3721 8805 3727 8933
rect 3721 8752 3727 8801
rect 3721 8640 3727 8748
rect 3721 8610 3727 8636
rect 3721 8554 3727 8606
rect 3721 8524 3727 8550
rect 3721 8384 3727 8520
rect 3721 8305 3727 8380
rect 3721 8272 3727 8301
rect 3721 8219 3727 8268
rect 3721 8170 3727 8215
rect 3721 8087 3727 8166
rect 3721 7955 3727 8083
rect 3721 7823 3727 7951
rect 3721 7770 3727 7819
rect 3721 7658 3727 7766
rect 3721 7628 3727 7654
rect 3721 7572 3727 7624
rect 3721 7542 3727 7568
rect 3721 7402 3727 7538
rect 3721 7381 3727 7398
rect 3733 9400 3739 9475
rect 3733 9208 3739 9396
rect 3733 9194 3739 9204
rect 3733 9076 3739 9190
rect 3733 9062 3739 9072
rect 3733 9012 3739 9058
rect 3733 8944 3739 9008
rect 3733 8930 3739 8940
rect 3733 8798 3739 8926
rect 3733 8724 3739 8794
rect 3733 8226 3739 8720
rect 3733 8212 3739 8222
rect 3733 8094 3739 8208
rect 3733 8080 3739 8090
rect 3733 7962 3739 8076
rect 3733 7948 3739 7958
rect 3733 7816 3739 7944
rect 3733 7742 3739 7812
rect 3733 7381 3739 7738
rect 3745 9408 3751 9482
rect 3745 9260 3751 9404
rect 3745 9128 3751 9256
rect 3745 9049 3751 9124
rect 3745 9010 3751 9045
rect 3745 8996 3751 9006
rect 3745 8878 3751 8992
rect 3745 8864 3751 8874
rect 3745 8732 3751 8860
rect 3745 8278 3751 8728
rect 3745 8146 3751 8274
rect 3745 8028 3751 8142
rect 3745 8014 3751 8024
rect 3745 7896 3751 8010
rect 3745 7882 3751 7892
rect 3745 7750 3751 7878
rect 3745 7381 3751 7746
rect 3757 9416 3763 9489
rect 3757 9280 3763 9412
rect 3757 9247 3763 9276
rect 3757 9145 3763 9243
rect 3757 8886 3763 9141
rect 3757 8746 3763 8882
rect 3757 8633 3763 8742
rect 3757 8603 3763 8629
rect 3757 8547 3763 8599
rect 3757 8517 3763 8543
rect 3757 8377 3763 8513
rect 3757 8298 3763 8373
rect 3757 8265 3763 8294
rect 3757 8163 3763 8261
rect 3757 7764 3763 8159
rect 3757 7651 3763 7760
rect 3757 7621 3763 7647
rect 3757 7565 3763 7617
rect 3757 7535 3763 7561
rect 3757 7395 3763 7531
rect 3757 7381 3763 7391
rect 3769 9351 3775 9497
rect 4483 9486 4484 9490
rect 4488 9486 4489 9490
rect 4493 9486 4494 9490
rect 4498 9486 4499 9490
rect 4503 9486 4504 9490
rect 4508 9486 4509 9490
rect 4479 9485 4513 9486
rect 4483 9481 4484 9485
rect 4488 9481 4489 9485
rect 4493 9481 4494 9485
rect 4498 9481 4499 9485
rect 4503 9481 4504 9485
rect 4508 9481 4509 9485
rect 4479 9480 4513 9481
rect 4483 9476 4484 9480
rect 4488 9476 4489 9480
rect 4493 9476 4494 9480
rect 4498 9476 4499 9480
rect 4503 9476 4504 9480
rect 4508 9476 4509 9480
rect 4479 9475 4513 9476
rect 4483 9471 4484 9475
rect 4488 9471 4489 9475
rect 4493 9471 4494 9475
rect 4498 9471 4499 9475
rect 4503 9471 4504 9475
rect 4508 9471 4509 9475
rect 4529 9486 4530 9490
rect 4534 9486 4535 9490
rect 4539 9486 4540 9490
rect 4544 9486 4545 9490
rect 4549 9486 4550 9490
rect 4554 9486 4555 9490
rect 4525 9485 4559 9486
rect 4529 9481 4530 9485
rect 4534 9481 4535 9485
rect 4539 9481 4540 9485
rect 4544 9481 4545 9485
rect 4549 9481 4550 9485
rect 4554 9481 4555 9485
rect 4525 9480 4559 9481
rect 4529 9476 4530 9480
rect 4534 9476 4535 9480
rect 4539 9476 4540 9480
rect 4544 9476 4545 9480
rect 4549 9476 4550 9480
rect 4554 9476 4555 9480
rect 4525 9475 4559 9476
rect 4529 9471 4530 9475
rect 4534 9471 4535 9475
rect 4539 9471 4540 9475
rect 4544 9471 4545 9475
rect 4549 9471 4550 9475
rect 4554 9471 4555 9475
rect 4483 9457 4484 9461
rect 4488 9457 4489 9461
rect 4493 9457 4494 9461
rect 4498 9457 4499 9461
rect 4503 9457 4504 9461
rect 4508 9457 4509 9461
rect 4479 9456 4513 9457
rect 3769 9318 3775 9347
rect 3769 9216 3775 9314
rect 3769 8916 3775 9212
rect 3769 8816 3775 8912
rect 3769 8704 3775 8812
rect 3769 8674 3775 8700
rect 3769 8618 3775 8670
rect 3769 8588 3775 8614
rect 3769 8448 3775 8584
rect 3769 8369 3775 8444
rect 3769 8336 3775 8365
rect 3769 8234 3775 8332
rect 3769 7834 3775 8230
rect 3769 7722 3775 7830
rect 3769 7692 3775 7718
rect 3769 7636 3775 7688
rect 3769 7606 3775 7632
rect 3769 7466 3775 7602
rect 3769 7381 3775 7462
rect 3781 9021 3787 9452
rect 4483 9452 4484 9456
rect 4488 9452 4489 9456
rect 4493 9452 4494 9456
rect 4498 9452 4499 9456
rect 4503 9452 4504 9456
rect 4508 9452 4509 9456
rect 4479 9451 4513 9452
rect 4483 9447 4484 9451
rect 4488 9447 4489 9451
rect 4493 9447 4494 9451
rect 4498 9447 4499 9451
rect 4503 9447 4504 9451
rect 4508 9447 4509 9451
rect 4479 9446 4513 9447
rect 4483 9442 4484 9446
rect 4488 9442 4489 9446
rect 4493 9442 4494 9446
rect 4498 9442 4499 9446
rect 4503 9442 4504 9446
rect 4508 9442 4509 9446
rect 4529 9457 4530 9461
rect 4534 9457 4535 9461
rect 4539 9457 4540 9461
rect 4544 9457 4545 9461
rect 4549 9457 4550 9461
rect 4554 9457 4555 9461
rect 4525 9456 4559 9457
rect 4529 9452 4530 9456
rect 4534 9452 4535 9456
rect 4539 9452 4540 9456
rect 4544 9452 4545 9456
rect 4549 9452 4550 9456
rect 4554 9452 4555 9456
rect 4525 9451 4559 9452
rect 4529 9447 4530 9451
rect 4534 9447 4535 9451
rect 4539 9447 4540 9451
rect 4544 9447 4545 9451
rect 4549 9447 4550 9451
rect 4554 9447 4555 9451
rect 4525 9446 4559 9447
rect 4529 9442 4530 9446
rect 4534 9442 4535 9446
rect 4539 9442 4540 9446
rect 4544 9442 4545 9446
rect 4549 9442 4550 9446
rect 4554 9442 4555 9446
rect 4579 9355 5073 9786
rect 3803 9337 3806 9347
rect 3810 9307 3813 9316
rect 3826 9309 3829 9322
rect 3839 9294 3842 9347
rect 3906 9337 3909 9347
rect 3935 9337 3938 9347
rect 3846 9322 3850 9326
rect 3847 9307 3850 9316
rect 3802 9280 3805 9292
rect 3843 9290 3844 9294
rect 3853 9280 3856 9333
rect 3859 9313 3862 9318
rect 3868 9307 3871 9316
rect 3884 9309 3887 9322
rect 3905 9307 3908 9316
rect 3921 9316 3924 9318
rect 3921 9313 3928 9316
rect 3921 9307 3924 9313
rect 3942 9307 3945 9316
rect 3958 9309 3961 9322
rect 3904 9280 3907 9290
rect 3921 9273 3924 9303
rect 3971 9294 3974 9347
rect 4038 9337 4041 9347
rect 4067 9337 4070 9347
rect 3978 9322 3982 9326
rect 3979 9307 3982 9316
rect 3934 9280 3937 9292
rect 3975 9290 3976 9294
rect 3985 9280 3988 9333
rect 3991 9313 3994 9318
rect 4000 9307 4003 9316
rect 4016 9309 4019 9322
rect 4037 9307 4040 9316
rect 4053 9316 4056 9318
rect 4053 9313 4060 9316
rect 4053 9307 4056 9313
rect 4074 9307 4077 9316
rect 4090 9309 4093 9322
rect 4036 9280 4039 9290
rect 3921 9270 3973 9273
rect 3801 9250 3804 9263
rect 3827 9253 3830 9256
rect 3834 9250 3837 9263
rect 3851 9250 3854 9263
rect 3801 9201 3804 9216
rect 3815 9208 3818 9212
rect 3833 9201 3836 9216
rect 3852 9201 3855 9216
rect 3858 9215 3861 9256
rect 3874 9208 3877 9249
rect 3880 9216 3883 9256
rect 3899 9208 3902 9249
rect 3908 9250 3911 9263
rect 3924 9250 3927 9263
rect 3945 9253 3948 9256
rect 3952 9250 3955 9263
rect 3970 9259 3973 9270
rect 4053 9267 4056 9303
rect 4103 9294 4106 9347
rect 4170 9337 4173 9347
rect 4199 9337 4202 9347
rect 4110 9322 4114 9326
rect 4111 9307 4114 9316
rect 4066 9280 4069 9292
rect 4107 9290 4108 9294
rect 4117 9280 4120 9333
rect 4123 9313 4126 9318
rect 4132 9307 4135 9316
rect 4148 9309 4151 9322
rect 4169 9307 4172 9316
rect 4185 9316 4188 9318
rect 4185 9313 4192 9316
rect 4185 9307 4188 9313
rect 4206 9307 4209 9316
rect 4222 9309 4225 9322
rect 4168 9280 4171 9290
rect 4185 9273 4188 9295
rect 4235 9294 4238 9347
rect 4302 9337 4305 9347
rect 4242 9322 4246 9326
rect 4243 9307 4246 9316
rect 4198 9280 4201 9292
rect 4239 9290 4240 9294
rect 4249 9280 4252 9333
rect 4255 9313 4258 9318
rect 4264 9307 4267 9316
rect 4280 9309 4283 9322
rect 4301 9307 4304 9316
rect 4317 9316 4320 9318
rect 4826 9316 5086 9319
rect 4317 9313 4321 9316
rect 4317 9307 4320 9313
rect 4317 9299 4320 9303
rect 4300 9280 4303 9290
rect 4051 9262 4056 9267
rect 4113 9269 4188 9273
rect 3970 9256 4015 9259
rect 3970 9246 3973 9256
rect 3988 9243 4008 9246
rect 4005 9224 4008 9243
rect 3908 9201 3911 9216
rect 3923 9201 3926 9216
rect 3930 9208 3934 9211
rect 3951 9201 3954 9216
rect 3801 9182 3804 9197
rect 3815 9186 3818 9190
rect 3833 9182 3836 9197
rect 3852 9182 3855 9197
rect 3801 9135 3804 9148
rect 3827 9142 3830 9145
rect 3801 9118 3804 9131
rect 3811 9128 3815 9138
rect 3834 9135 3837 9148
rect 3851 9135 3854 9148
rect 3858 9142 3861 9183
rect 3874 9149 3877 9190
rect 3880 9142 3883 9182
rect 3899 9149 3902 9190
rect 3908 9182 3911 9197
rect 3923 9182 3926 9197
rect 3930 9187 3934 9190
rect 3951 9182 3954 9197
rect 3908 9135 3911 9148
rect 3827 9121 3830 9124
rect 3834 9118 3837 9131
rect 3851 9118 3854 9131
rect 3801 9069 3804 9084
rect 3815 9076 3818 9080
rect 3833 9069 3836 9084
rect 3852 9069 3855 9084
rect 3858 9083 3861 9124
rect 3874 9076 3877 9117
rect 3880 9084 3883 9124
rect 3899 9076 3902 9117
rect 3908 9118 3911 9131
rect 3924 9135 3927 9148
rect 3945 9142 3948 9145
rect 3952 9135 3955 9148
rect 4005 9148 4008 9220
rect 4016 9184 4019 9256
rect 4051 9259 4054 9262
rect 4051 9256 4096 9259
rect 4051 9246 4054 9256
rect 3924 9118 3927 9131
rect 3945 9121 3948 9124
rect 3952 9118 3955 9131
rect 4005 9114 4008 9144
rect 4016 9128 4019 9180
rect 4023 9168 4027 9234
rect 4011 9124 4015 9127
rect 4004 9111 4008 9114
rect 4005 9092 4008 9111
rect 3908 9069 3911 9084
rect 3923 9069 3926 9084
rect 3930 9076 3934 9079
rect 3951 9069 3954 9084
rect 3801 9050 3804 9065
rect 3815 9054 3818 9058
rect 3833 9050 3836 9065
rect 3852 9050 3855 9065
rect 3781 8718 3787 9017
rect 3801 9003 3804 9016
rect 3827 9010 3830 9013
rect 3801 8986 3804 8999
rect 3834 9003 3837 9016
rect 3851 9003 3854 9016
rect 3858 9010 3861 9051
rect 3874 9017 3877 9058
rect 3880 9010 3883 9050
rect 3899 9017 3902 9058
rect 3908 9050 3911 9065
rect 3923 9050 3926 9065
rect 3930 9055 3934 9058
rect 3951 9050 3954 9065
rect 3908 9003 3911 9016
rect 3827 8989 3830 8992
rect 3834 8986 3837 8999
rect 3851 8986 3854 8999
rect 3801 8937 3804 8952
rect 3815 8944 3818 8948
rect 3833 8937 3836 8952
rect 3852 8937 3855 8952
rect 3858 8951 3861 8992
rect 3874 8944 3877 8985
rect 3880 8952 3883 8992
rect 3899 8944 3902 8985
rect 3908 8986 3911 8999
rect 3924 9003 3927 9016
rect 3945 9010 3948 9013
rect 3952 9003 3955 9016
rect 4005 9017 4008 9088
rect 4016 9053 4019 9124
rect 3924 8986 3927 8999
rect 3945 8989 3948 8992
rect 3952 8986 3955 8999
rect 4005 8960 4008 9013
rect 4016 8996 4019 9049
rect 4023 9037 4027 9102
rect 4011 8992 4015 8995
rect 4054 8995 4057 9246
rect 4069 9243 4089 9246
rect 4086 9224 4089 9243
rect 4086 9148 4089 9220
rect 4097 9184 4100 9256
rect 4104 9168 4108 9234
rect 4113 9135 4116 9269
rect 4317 9266 4320 9295
rect 4141 9263 4248 9266
rect 4075 9131 4116 9135
rect 4075 9127 4078 9131
rect 4075 9124 4120 9127
rect 4075 9114 4078 9124
rect 4093 9111 4113 9114
rect 4075 9109 4078 9110
rect 4110 9092 4113 9111
rect 4110 9017 4113 9088
rect 4121 9053 4124 9124
rect 4128 9037 4132 9102
rect 3908 8937 3911 8952
rect 3923 8937 3926 8952
rect 3930 8944 3934 8947
rect 3951 8937 3954 8952
rect 3801 8918 3804 8933
rect 3815 8922 3818 8926
rect 3833 8918 3836 8933
rect 3852 8918 3855 8933
rect 3801 8871 3804 8884
rect 3827 8878 3830 8881
rect 3801 8854 3804 8867
rect 3834 8871 3837 8884
rect 3851 8871 3854 8884
rect 3858 8878 3861 8919
rect 3874 8885 3877 8926
rect 3880 8878 3883 8918
rect 3899 8885 3902 8926
rect 3908 8918 3911 8933
rect 3923 8918 3926 8933
rect 3930 8923 3934 8926
rect 3951 8918 3954 8933
rect 3908 8871 3911 8884
rect 3827 8857 3830 8860
rect 3834 8854 3837 8867
rect 3851 8854 3854 8867
rect 3801 8805 3804 8820
rect 3815 8812 3818 8816
rect 3801 8786 3804 8801
rect 3824 8798 3828 8808
rect 3833 8805 3836 8820
rect 3852 8805 3855 8820
rect 3858 8819 3861 8860
rect 3874 8812 3877 8853
rect 3880 8820 3883 8860
rect 3899 8812 3902 8853
rect 3908 8854 3911 8867
rect 3924 8871 3927 8884
rect 3945 8878 3948 8881
rect 3952 8871 3955 8884
rect 4005 8882 4008 8956
rect 4016 8918 4019 8992
rect 4051 8992 4096 8995
rect 4051 8982 4054 8992
rect 4069 8979 4089 8982
rect 3924 8854 3927 8867
rect 3945 8857 3948 8860
rect 3952 8854 3955 8867
rect 4005 8828 4008 8878
rect 4016 8864 4019 8914
rect 4023 8902 4027 8970
rect 4086 8960 4089 8979
rect 4086 8882 4089 8956
rect 4097 8918 4100 8992
rect 4141 8995 4144 9263
rect 4252 9263 4320 9266
rect 4826 9062 4829 9316
rect 5083 9062 5086 9316
rect 4483 9056 4484 9060
rect 4488 9056 4489 9060
rect 4493 9056 4494 9060
rect 4498 9056 4499 9060
rect 4503 9056 4504 9060
rect 4508 9056 4509 9060
rect 4479 9055 4513 9056
rect 4483 9051 4484 9055
rect 4488 9051 4489 9055
rect 4493 9051 4494 9055
rect 4498 9051 4499 9055
rect 4503 9051 4504 9055
rect 4508 9051 4509 9055
rect 4479 9050 4513 9051
rect 4483 9046 4484 9050
rect 4488 9046 4489 9050
rect 4493 9046 4494 9050
rect 4498 9046 4499 9050
rect 4503 9046 4504 9050
rect 4508 9046 4509 9050
rect 4479 9045 4513 9046
rect 4483 9041 4484 9045
rect 4488 9041 4489 9045
rect 4493 9041 4494 9045
rect 4498 9041 4499 9045
rect 4503 9041 4504 9045
rect 4508 9041 4509 9045
rect 4529 9056 4530 9060
rect 4534 9056 4535 9060
rect 4539 9056 4540 9060
rect 4544 9056 4545 9060
rect 4549 9056 4550 9060
rect 4554 9056 4555 9060
rect 4826 9059 5086 9062
rect 4525 9055 4559 9056
rect 4529 9051 4530 9055
rect 4534 9051 4535 9055
rect 4539 9051 4540 9055
rect 4544 9051 4545 9055
rect 4549 9051 4550 9055
rect 4554 9051 4555 9055
rect 4525 9050 4559 9051
rect 4529 9046 4530 9050
rect 4534 9046 4535 9050
rect 4539 9046 4540 9050
rect 4544 9046 4545 9050
rect 4549 9046 4550 9050
rect 4554 9046 4555 9050
rect 4525 9045 4559 9046
rect 4529 9041 4530 9045
rect 4534 9041 4535 9045
rect 4539 9041 4540 9045
rect 4544 9041 4545 9045
rect 4549 9041 4550 9045
rect 4554 9041 4555 9045
rect 4826 9007 5086 9010
rect 4141 8992 4186 8995
rect 4141 8982 4144 8992
rect 4159 8979 4179 8982
rect 4104 8902 4108 8970
rect 4176 8960 4179 8979
rect 4176 8882 4179 8956
rect 4187 8918 4190 8992
rect 4194 8902 4198 8970
rect 4011 8860 4015 8863
rect 3908 8805 3911 8820
rect 3923 8805 3926 8820
rect 3930 8812 3934 8815
rect 3951 8805 3954 8820
rect 3815 8790 3818 8794
rect 3833 8786 3836 8801
rect 3852 8786 3855 8801
rect 3801 8739 3804 8752
rect 3827 8746 3830 8749
rect 3809 8732 3813 8742
rect 3834 8739 3837 8752
rect 3851 8739 3854 8752
rect 3858 8746 3861 8787
rect 3874 8753 3877 8794
rect 3880 8746 3883 8786
rect 3899 8753 3902 8794
rect 3908 8786 3911 8801
rect 3923 8786 3926 8801
rect 3930 8791 3934 8794
rect 3951 8786 3954 8801
rect 3908 8739 3911 8752
rect 3924 8739 3927 8752
rect 3945 8746 3948 8749
rect 3952 8739 3955 8752
rect 4005 8746 4008 8824
rect 4016 8782 4019 8860
rect 4023 8766 4027 8838
rect 4035 8739 4039 8752
rect 4044 8732 4047 8742
rect 4054 8725 4057 8794
rect 4076 8790 4079 8794
rect 4094 8786 4097 8801
rect 4113 8786 4116 8801
rect 4061 8739 4065 8752
rect 4088 8746 4091 8749
rect 4095 8739 4098 8752
rect 4112 8739 4115 8752
rect 4119 8746 4122 8787
rect 4135 8753 4138 8794
rect 4141 8746 4144 8786
rect 4160 8753 4163 8794
rect 4169 8786 4172 8801
rect 4184 8786 4187 8801
rect 4191 8791 4195 8794
rect 4212 8786 4215 8801
rect 4169 8739 4172 8752
rect 4185 8739 4188 8752
rect 4206 8746 4209 8749
rect 4213 8739 4216 8752
rect 4229 8733 4233 8969
rect 4826 8753 4829 9007
rect 5083 8753 5086 9007
rect 4483 8747 4484 8751
rect 4488 8747 4489 8751
rect 4493 8747 4494 8751
rect 4498 8747 4499 8751
rect 4503 8747 4504 8751
rect 4508 8747 4509 8751
rect 4479 8746 4513 8747
rect 4483 8742 4484 8746
rect 4488 8742 4489 8746
rect 4493 8742 4494 8746
rect 4498 8742 4499 8746
rect 4503 8742 4504 8746
rect 4508 8742 4509 8746
rect 4479 8741 4513 8742
rect 4483 8737 4484 8741
rect 4488 8737 4489 8741
rect 4493 8737 4494 8741
rect 4498 8737 4499 8741
rect 4503 8737 4504 8741
rect 4508 8737 4509 8741
rect 4479 8736 4513 8737
rect 4483 8732 4484 8736
rect 4488 8732 4489 8736
rect 4493 8732 4494 8736
rect 4498 8732 4499 8736
rect 4503 8732 4504 8736
rect 4508 8732 4509 8736
rect 4529 8747 4530 8751
rect 4534 8747 4535 8751
rect 4539 8747 4540 8751
rect 4544 8747 4545 8751
rect 4549 8747 4550 8751
rect 4554 8747 4555 8751
rect 4826 8750 5086 8753
rect 4525 8746 4559 8747
rect 4529 8742 4530 8746
rect 4534 8742 4535 8746
rect 4539 8742 4540 8746
rect 4544 8742 4545 8746
rect 4549 8742 4550 8746
rect 4554 8742 4555 8746
rect 4525 8741 4559 8742
rect 4529 8737 4530 8741
rect 4534 8737 4535 8741
rect 4539 8737 4540 8741
rect 4544 8737 4545 8741
rect 4549 8737 4550 8741
rect 4554 8737 4555 8741
rect 4525 8736 4559 8737
rect 4529 8732 4530 8736
rect 4534 8732 4535 8736
rect 4539 8732 4540 8736
rect 4544 8732 4545 8736
rect 4549 8732 4550 8736
rect 4554 8732 4555 8736
rect 4222 8721 4223 8724
rect 3781 7736 3787 8714
rect 4087 8611 4091 8693
rect 4102 8690 4105 8700
rect 4109 8660 4112 8669
rect 4125 8662 4128 8675
rect 4138 8647 4141 8700
rect 4205 8690 4208 8700
rect 4145 8675 4149 8679
rect 4146 8660 4149 8669
rect 4101 8633 4104 8645
rect 4142 8643 4143 8647
rect 4152 8633 4155 8686
rect 4220 8675 4223 8721
rect 4158 8666 4161 8671
rect 4167 8660 4170 8669
rect 4183 8662 4186 8675
rect 4204 8660 4207 8669
rect 4220 8660 4223 8669
rect 4203 8633 4206 8643
rect 4220 8626 4223 8656
rect 4095 8584 4098 8621
rect 4102 8604 4105 8614
rect 4109 8574 4112 8583
rect 4125 8576 4128 8589
rect 4138 8561 4141 8614
rect 4205 8604 4208 8614
rect 4145 8589 4149 8593
rect 4146 8574 4149 8583
rect 4101 8547 4104 8559
rect 4142 8557 4143 8561
rect 4152 8547 4155 8600
rect 4158 8580 4161 8585
rect 4167 8574 4170 8583
rect 4183 8576 4186 8589
rect 4204 8574 4207 8583
rect 4220 8584 4223 8585
rect 4241 8587 4245 8729
rect 4826 8698 5086 8701
rect 4220 8579 4223 8580
rect 4203 8547 4206 8557
rect 4241 8485 4245 8567
rect 4826 8444 4829 8698
rect 5083 8444 5086 8698
rect 4483 8438 4484 8442
rect 4488 8438 4489 8442
rect 4493 8438 4494 8442
rect 4498 8438 4499 8442
rect 4503 8438 4504 8442
rect 4508 8438 4509 8442
rect 4479 8437 4513 8438
rect 4483 8433 4484 8437
rect 4488 8433 4489 8437
rect 4493 8433 4494 8437
rect 4498 8433 4499 8437
rect 4503 8433 4504 8437
rect 4508 8433 4509 8437
rect 4479 8432 4513 8433
rect 4483 8428 4484 8432
rect 4488 8428 4489 8432
rect 4493 8428 4494 8432
rect 4498 8428 4499 8432
rect 4503 8428 4504 8432
rect 4508 8428 4509 8432
rect 4479 8427 4513 8428
rect 4483 8423 4484 8427
rect 4488 8423 4489 8427
rect 4493 8423 4494 8427
rect 4498 8423 4499 8427
rect 4503 8423 4504 8427
rect 4508 8423 4509 8427
rect 4529 8438 4530 8442
rect 4534 8438 4535 8442
rect 4539 8438 4540 8442
rect 4544 8438 4545 8442
rect 4549 8438 4550 8442
rect 4554 8438 4555 8442
rect 4826 8441 5086 8444
rect 4525 8437 4559 8438
rect 4529 8433 4530 8437
rect 4534 8433 4535 8437
rect 4539 8433 4540 8437
rect 4544 8433 4545 8437
rect 4549 8433 4550 8437
rect 4554 8433 4555 8437
rect 4525 8432 4559 8433
rect 4529 8428 4530 8432
rect 4534 8428 4535 8432
rect 4539 8428 4540 8432
rect 4544 8428 4545 8432
rect 4549 8428 4550 8432
rect 4554 8428 4555 8432
rect 4525 8427 4559 8428
rect 4529 8423 4530 8427
rect 4534 8423 4535 8427
rect 4539 8423 4540 8427
rect 4544 8423 4545 8427
rect 4549 8423 4550 8427
rect 4554 8423 4555 8427
rect 4826 8389 5086 8392
rect 3803 8355 3806 8365
rect 3810 8325 3813 8334
rect 3826 8327 3829 8340
rect 3839 8312 3842 8365
rect 3906 8355 3909 8365
rect 3935 8355 3938 8365
rect 3846 8340 3850 8344
rect 3847 8325 3850 8334
rect 3802 8298 3805 8310
rect 3843 8308 3844 8312
rect 3853 8298 3856 8351
rect 3859 8331 3862 8336
rect 3868 8325 3871 8334
rect 3884 8327 3887 8340
rect 3905 8325 3908 8334
rect 3921 8334 3924 8336
rect 3921 8331 3928 8334
rect 3921 8325 3924 8331
rect 3942 8325 3945 8334
rect 3958 8327 3961 8340
rect 3904 8298 3907 8308
rect 3921 8291 3924 8321
rect 3971 8312 3974 8365
rect 4038 8355 4041 8365
rect 4067 8355 4070 8365
rect 3978 8340 3982 8344
rect 3979 8325 3982 8334
rect 3934 8298 3937 8310
rect 3975 8308 3976 8312
rect 3985 8298 3988 8351
rect 3991 8331 3994 8336
rect 4000 8325 4003 8334
rect 4016 8327 4019 8340
rect 4037 8325 4040 8334
rect 4053 8334 4056 8336
rect 4053 8331 4060 8334
rect 4053 8325 4056 8331
rect 4074 8325 4077 8334
rect 4090 8327 4093 8340
rect 4036 8298 4039 8308
rect 3921 8288 3973 8291
rect 3801 8268 3804 8281
rect 3827 8271 3830 8274
rect 3834 8268 3837 8281
rect 3851 8268 3854 8281
rect 3801 8219 3804 8234
rect 3815 8226 3818 8230
rect 3833 8219 3836 8234
rect 3852 8219 3855 8234
rect 3858 8233 3861 8274
rect 3874 8226 3877 8267
rect 3880 8234 3883 8274
rect 3899 8226 3902 8267
rect 3908 8268 3911 8281
rect 3924 8268 3927 8281
rect 3945 8271 3948 8274
rect 3952 8268 3955 8281
rect 3970 8277 3973 8288
rect 4053 8285 4056 8321
rect 4103 8312 4106 8365
rect 4170 8355 4173 8365
rect 4199 8355 4202 8365
rect 4110 8340 4114 8344
rect 4111 8325 4114 8334
rect 4066 8298 4069 8310
rect 4107 8308 4108 8312
rect 4117 8298 4120 8351
rect 4123 8331 4126 8336
rect 4132 8325 4135 8334
rect 4148 8327 4151 8340
rect 4169 8325 4172 8334
rect 4185 8334 4188 8336
rect 4185 8331 4192 8334
rect 4185 8325 4188 8331
rect 4206 8325 4209 8334
rect 4222 8327 4225 8340
rect 4168 8298 4171 8308
rect 4185 8291 4188 8313
rect 4235 8312 4238 8365
rect 4302 8355 4305 8365
rect 4242 8340 4246 8344
rect 4243 8325 4246 8334
rect 4198 8298 4201 8310
rect 4239 8308 4240 8312
rect 4249 8298 4252 8351
rect 4255 8331 4258 8336
rect 4264 8325 4267 8334
rect 4280 8327 4283 8340
rect 4301 8325 4304 8334
rect 4317 8334 4320 8336
rect 4317 8331 4321 8334
rect 4317 8325 4320 8331
rect 4317 8317 4320 8321
rect 4300 8298 4303 8308
rect 4051 8280 4056 8285
rect 4113 8287 4188 8291
rect 3970 8274 4015 8277
rect 3970 8264 3973 8274
rect 3988 8261 4008 8264
rect 4005 8242 4008 8261
rect 3908 8219 3911 8234
rect 3923 8219 3926 8234
rect 3930 8226 3934 8229
rect 3951 8219 3954 8234
rect 3801 8200 3804 8215
rect 3815 8204 3818 8208
rect 3833 8200 3836 8215
rect 3852 8200 3855 8215
rect 3801 8153 3804 8166
rect 3827 8160 3830 8163
rect 3801 8136 3804 8149
rect 3811 8146 3815 8156
rect 3834 8153 3837 8166
rect 3851 8153 3854 8166
rect 3858 8160 3861 8201
rect 3874 8167 3877 8208
rect 3880 8160 3883 8200
rect 3899 8167 3902 8208
rect 3908 8200 3911 8215
rect 3923 8200 3926 8215
rect 3930 8205 3934 8208
rect 3951 8200 3954 8215
rect 3908 8153 3911 8166
rect 3827 8139 3830 8142
rect 3834 8136 3837 8149
rect 3851 8136 3854 8149
rect 3801 8087 3804 8102
rect 3815 8094 3818 8098
rect 3833 8087 3836 8102
rect 3852 8087 3855 8102
rect 3858 8101 3861 8142
rect 3874 8094 3877 8135
rect 3880 8102 3883 8142
rect 3899 8094 3902 8135
rect 3908 8136 3911 8149
rect 3924 8153 3927 8166
rect 3945 8160 3948 8163
rect 3952 8153 3955 8166
rect 4005 8166 4008 8238
rect 4016 8202 4019 8274
rect 4051 8277 4054 8280
rect 4051 8274 4096 8277
rect 4051 8264 4054 8274
rect 3924 8136 3927 8149
rect 3945 8139 3948 8142
rect 3952 8136 3955 8149
rect 4005 8132 4008 8162
rect 4016 8146 4019 8198
rect 4023 8186 4027 8252
rect 4011 8142 4015 8145
rect 4004 8129 4008 8132
rect 4005 8110 4008 8129
rect 3908 8087 3911 8102
rect 3923 8087 3926 8102
rect 3930 8094 3934 8097
rect 3951 8087 3954 8102
rect 3801 8068 3804 8083
rect 3815 8072 3818 8076
rect 3833 8068 3836 8083
rect 3852 8068 3855 8083
rect 3801 8021 3804 8034
rect 3827 8028 3830 8031
rect 3801 8004 3804 8017
rect 3834 8021 3837 8034
rect 3851 8021 3854 8034
rect 3858 8028 3861 8069
rect 3874 8035 3877 8076
rect 3880 8028 3883 8068
rect 3899 8035 3902 8076
rect 3908 8068 3911 8083
rect 3923 8068 3926 8083
rect 3930 8073 3934 8076
rect 3951 8068 3954 8083
rect 3908 8021 3911 8034
rect 3827 8007 3830 8010
rect 3834 8004 3837 8017
rect 3851 8004 3854 8017
rect 3801 7955 3804 7970
rect 3815 7962 3818 7966
rect 3833 7955 3836 7970
rect 3852 7955 3855 7970
rect 3858 7969 3861 8010
rect 3874 7962 3877 8003
rect 3880 7970 3883 8010
rect 3899 7962 3902 8003
rect 3908 8004 3911 8017
rect 3924 8021 3927 8034
rect 3945 8028 3948 8031
rect 3952 8021 3955 8034
rect 4005 8035 4008 8106
rect 4016 8071 4019 8142
rect 3924 8004 3927 8017
rect 3945 8007 3948 8010
rect 3952 8004 3955 8017
rect 4005 7978 4008 8031
rect 4016 8014 4019 8067
rect 4023 8055 4027 8120
rect 4011 8010 4015 8013
rect 4054 8013 4057 8264
rect 4069 8261 4089 8264
rect 4086 8242 4089 8261
rect 4086 8166 4089 8238
rect 4097 8202 4100 8274
rect 4104 8186 4108 8252
rect 4113 8153 4116 8287
rect 4317 8284 4320 8313
rect 4141 8281 4248 8284
rect 4075 8149 4116 8153
rect 4075 8145 4078 8149
rect 4075 8142 4120 8145
rect 4075 8132 4078 8142
rect 4093 8129 4113 8132
rect 4075 8127 4078 8128
rect 4110 8110 4113 8129
rect 4110 8035 4113 8106
rect 4121 8071 4124 8142
rect 4128 8055 4132 8120
rect 3908 7955 3911 7970
rect 3923 7955 3926 7970
rect 3930 7962 3934 7965
rect 3951 7955 3954 7970
rect 3801 7936 3804 7951
rect 3815 7940 3818 7944
rect 3833 7936 3836 7951
rect 3852 7936 3855 7951
rect 3801 7889 3804 7902
rect 3827 7896 3830 7899
rect 3801 7872 3804 7885
rect 3834 7889 3837 7902
rect 3851 7889 3854 7902
rect 3858 7896 3861 7937
rect 3874 7903 3877 7944
rect 3880 7896 3883 7936
rect 3899 7903 3902 7944
rect 3908 7936 3911 7951
rect 3923 7936 3926 7951
rect 3930 7941 3934 7944
rect 3951 7936 3954 7951
rect 3908 7889 3911 7902
rect 3827 7875 3830 7878
rect 3834 7872 3837 7885
rect 3851 7872 3854 7885
rect 3801 7823 3804 7838
rect 3815 7830 3818 7834
rect 3801 7804 3804 7819
rect 3824 7816 3828 7826
rect 3833 7823 3836 7838
rect 3852 7823 3855 7838
rect 3858 7837 3861 7878
rect 3874 7830 3877 7871
rect 3880 7838 3883 7878
rect 3899 7830 3902 7871
rect 3908 7872 3911 7885
rect 3924 7889 3927 7902
rect 3945 7896 3948 7899
rect 3952 7889 3955 7902
rect 4005 7900 4008 7974
rect 4016 7936 4019 8010
rect 4051 8010 4096 8013
rect 4051 8000 4054 8010
rect 4069 7997 4089 8000
rect 3924 7872 3927 7885
rect 3945 7875 3948 7878
rect 3952 7872 3955 7885
rect 4005 7846 4008 7896
rect 4016 7882 4019 7932
rect 4023 7920 4027 7988
rect 4086 7978 4089 7997
rect 4086 7900 4089 7974
rect 4097 7936 4100 8010
rect 4141 8013 4144 8281
rect 4252 8281 4320 8284
rect 4826 8135 4829 8389
rect 5083 8135 5086 8389
rect 4483 8129 4484 8133
rect 4488 8129 4489 8133
rect 4493 8129 4494 8133
rect 4498 8129 4499 8133
rect 4503 8129 4504 8133
rect 4508 8129 4509 8133
rect 4479 8128 4513 8129
rect 4483 8124 4484 8128
rect 4488 8124 4489 8128
rect 4493 8124 4494 8128
rect 4498 8124 4499 8128
rect 4503 8124 4504 8128
rect 4508 8124 4509 8128
rect 4479 8123 4513 8124
rect 4483 8119 4484 8123
rect 4488 8119 4489 8123
rect 4493 8119 4494 8123
rect 4498 8119 4499 8123
rect 4503 8119 4504 8123
rect 4508 8119 4509 8123
rect 4479 8118 4513 8119
rect 4483 8114 4484 8118
rect 4488 8114 4489 8118
rect 4493 8114 4494 8118
rect 4498 8114 4499 8118
rect 4503 8114 4504 8118
rect 4508 8114 4509 8118
rect 4529 8129 4530 8133
rect 4534 8129 4535 8133
rect 4539 8129 4540 8133
rect 4544 8129 4545 8133
rect 4549 8129 4550 8133
rect 4554 8129 4555 8133
rect 4826 8132 5086 8135
rect 4525 8128 4559 8129
rect 4529 8124 4530 8128
rect 4534 8124 4535 8128
rect 4539 8124 4540 8128
rect 4544 8124 4545 8128
rect 4549 8124 4550 8128
rect 4554 8124 4555 8128
rect 4525 8123 4559 8124
rect 4529 8119 4530 8123
rect 4534 8119 4535 8123
rect 4539 8119 4540 8123
rect 4544 8119 4545 8123
rect 4549 8119 4550 8123
rect 4554 8119 4555 8123
rect 4525 8118 4559 8119
rect 4529 8114 4530 8118
rect 4534 8114 4535 8118
rect 4539 8114 4540 8118
rect 4544 8114 4545 8118
rect 4549 8114 4550 8118
rect 4554 8114 4555 8118
rect 4483 8098 4484 8102
rect 4488 8098 4489 8102
rect 4493 8098 4494 8102
rect 4498 8098 4499 8102
rect 4503 8098 4504 8102
rect 4508 8098 4509 8102
rect 4479 8097 4513 8098
rect 4483 8093 4484 8097
rect 4488 8093 4489 8097
rect 4493 8093 4494 8097
rect 4498 8093 4499 8097
rect 4503 8093 4504 8097
rect 4508 8093 4509 8097
rect 4479 8092 4513 8093
rect 4483 8088 4484 8092
rect 4488 8088 4489 8092
rect 4493 8088 4494 8092
rect 4498 8088 4499 8092
rect 4503 8088 4504 8092
rect 4508 8088 4509 8092
rect 4479 8087 4513 8088
rect 4483 8083 4484 8087
rect 4488 8083 4489 8087
rect 4493 8083 4494 8087
rect 4498 8083 4499 8087
rect 4503 8083 4504 8087
rect 4508 8083 4509 8087
rect 4529 8098 4530 8102
rect 4534 8098 4535 8102
rect 4539 8098 4540 8102
rect 4544 8098 4545 8102
rect 4549 8098 4550 8102
rect 4554 8098 4555 8102
rect 4525 8097 4559 8098
rect 4529 8093 4530 8097
rect 4534 8093 4535 8097
rect 4539 8093 4540 8097
rect 4544 8093 4545 8097
rect 4549 8093 4550 8097
rect 4554 8093 4555 8097
rect 4525 8092 4559 8093
rect 4529 8088 4530 8092
rect 4534 8088 4535 8092
rect 4539 8088 4540 8092
rect 4544 8088 4545 8092
rect 4549 8088 4550 8092
rect 4554 8088 4555 8092
rect 4525 8087 4559 8088
rect 4529 8083 4530 8087
rect 4534 8083 4535 8087
rect 4539 8083 4540 8087
rect 4544 8083 4545 8087
rect 4549 8083 4550 8087
rect 4554 8083 4555 8087
rect 4826 8081 5086 8084
rect 4494 8078 4515 8080
rect 4494 8074 4496 8078
rect 4500 8074 4501 8078
rect 4505 8074 4506 8078
rect 4510 8074 4511 8078
rect 4494 8073 4515 8074
rect 4494 8069 4496 8073
rect 4500 8069 4501 8073
rect 4505 8069 4506 8073
rect 4510 8069 4511 8073
rect 4494 8068 4515 8069
rect 4494 8064 4496 8068
rect 4500 8064 4501 8068
rect 4505 8064 4506 8068
rect 4510 8064 4511 8068
rect 4494 8063 4515 8064
rect 4494 8059 4496 8063
rect 4500 8059 4501 8063
rect 4505 8059 4506 8063
rect 4510 8059 4511 8063
rect 4494 8058 4515 8059
rect 4494 8054 4496 8058
rect 4500 8054 4501 8058
rect 4505 8054 4506 8058
rect 4510 8054 4511 8058
rect 4494 8053 4515 8054
rect 4494 8049 4496 8053
rect 4500 8049 4501 8053
rect 4505 8049 4506 8053
rect 4510 8049 4511 8053
rect 4494 8048 4515 8049
rect 4494 8044 4496 8048
rect 4500 8044 4501 8048
rect 4505 8044 4506 8048
rect 4510 8044 4511 8048
rect 4494 8043 4515 8044
rect 4494 8039 4496 8043
rect 4500 8039 4501 8043
rect 4505 8039 4506 8043
rect 4510 8039 4511 8043
rect 4494 8038 4515 8039
rect 4494 8034 4496 8038
rect 4500 8034 4501 8038
rect 4505 8034 4506 8038
rect 4510 8034 4511 8038
rect 4494 8033 4515 8034
rect 4494 8029 4496 8033
rect 4500 8029 4501 8033
rect 4505 8029 4506 8033
rect 4510 8029 4511 8033
rect 4494 8028 4515 8029
rect 4494 8024 4496 8028
rect 4500 8024 4501 8028
rect 4505 8024 4506 8028
rect 4510 8024 4511 8028
rect 4141 8010 4186 8013
rect 4141 8000 4144 8010
rect 4159 7997 4179 8000
rect 4104 7920 4108 7988
rect 4176 7978 4179 7997
rect 4176 7900 4179 7974
rect 4187 7936 4190 8010
rect 4194 7920 4198 7988
rect 4011 7878 4015 7881
rect 3908 7823 3911 7838
rect 3923 7823 3926 7838
rect 3930 7830 3934 7833
rect 3951 7823 3954 7838
rect 3815 7808 3818 7812
rect 3833 7804 3836 7819
rect 3852 7804 3855 7819
rect 3801 7757 3804 7770
rect 3827 7764 3830 7767
rect 3809 7750 3813 7760
rect 3834 7757 3837 7770
rect 3851 7757 3854 7770
rect 3858 7764 3861 7805
rect 3874 7771 3877 7812
rect 3880 7764 3883 7804
rect 3899 7771 3902 7812
rect 3908 7804 3911 7819
rect 3923 7804 3926 7819
rect 3930 7809 3934 7812
rect 3951 7804 3954 7819
rect 3908 7757 3911 7770
rect 3924 7757 3927 7770
rect 3945 7764 3948 7767
rect 3952 7757 3955 7770
rect 4005 7764 4008 7842
rect 4016 7800 4019 7878
rect 4023 7784 4027 7856
rect 4035 7757 4039 7770
rect 4044 7750 4047 7760
rect 4054 7743 4057 7812
rect 4076 7808 4079 7812
rect 4094 7804 4097 7819
rect 4113 7804 4116 7819
rect 4061 7757 4065 7770
rect 4088 7764 4091 7767
rect 4095 7757 4098 7770
rect 4112 7757 4115 7770
rect 4119 7764 4122 7805
rect 4135 7771 4138 7812
rect 4141 7764 4144 7804
rect 4160 7771 4163 7812
rect 4169 7804 4172 7819
rect 4184 7804 4187 7819
rect 4191 7809 4195 7812
rect 4212 7804 4215 7819
rect 4169 7757 4172 7770
rect 4185 7757 4188 7770
rect 4206 7764 4209 7767
rect 4213 7757 4216 7770
rect 4229 7751 4233 7987
rect 4377 7963 4386 7987
rect 4578 7982 4590 7986
rect 4594 7982 4606 7986
rect 4610 7982 4622 7986
rect 4626 7982 4645 7986
rect 4649 7982 4661 7986
rect 4665 7982 4688 7986
rect 4692 7982 4704 7986
rect 4708 7982 4729 7986
rect 4733 7982 4745 7986
rect 4657 7963 4717 7965
rect 4657 7954 4659 7963
rect 4667 7954 4703 7963
rect 4711 7954 4717 7963
rect 4657 7952 4717 7954
rect 4578 7924 4590 7928
rect 4594 7924 4606 7928
rect 4610 7924 4622 7928
rect 4626 7924 4645 7928
rect 4649 7924 4661 7928
rect 4665 7924 4688 7928
rect 4692 7924 4704 7928
rect 4708 7924 4729 7928
rect 4733 7924 4745 7928
rect 4527 7824 4529 7828
rect 4533 7824 4534 7828
rect 4538 7824 4539 7828
rect 4543 7824 4544 7828
rect 4548 7824 4549 7828
rect 4553 7824 4554 7828
rect 4558 7824 4559 7828
rect 4563 7824 4564 7828
rect 4568 7824 4569 7828
rect 4573 7824 4574 7828
rect 4578 7824 4579 7828
rect 4583 7824 4584 7828
rect 4588 7824 4589 7828
rect 4593 7824 4595 7828
rect 4826 7827 4829 8081
rect 5083 7827 5086 8081
rect 4826 7824 5086 7827
rect 4527 7823 4595 7824
rect 4527 7819 4529 7823
rect 4533 7819 4534 7823
rect 4538 7819 4539 7823
rect 4543 7819 4544 7823
rect 4548 7819 4549 7823
rect 4553 7819 4554 7823
rect 4558 7819 4559 7823
rect 4563 7819 4564 7823
rect 4568 7819 4569 7823
rect 4573 7819 4574 7823
rect 4578 7819 4579 7823
rect 4583 7819 4584 7823
rect 4588 7819 4589 7823
rect 4593 7819 4595 7823
rect 4527 7818 4595 7819
rect 4527 7814 4529 7818
rect 4533 7814 4534 7818
rect 4538 7814 4539 7818
rect 4543 7814 4544 7818
rect 4548 7814 4549 7818
rect 4553 7814 4554 7818
rect 4558 7814 4559 7818
rect 4563 7814 4564 7818
rect 4568 7814 4569 7818
rect 4573 7814 4574 7818
rect 4578 7814 4579 7818
rect 4583 7814 4584 7818
rect 4588 7814 4589 7818
rect 4593 7814 4595 7818
rect 4527 7813 4595 7814
rect 4527 7809 4529 7813
rect 4533 7809 4534 7813
rect 4538 7809 4539 7813
rect 4543 7809 4544 7813
rect 4548 7809 4549 7813
rect 4553 7809 4554 7813
rect 4558 7809 4559 7813
rect 4563 7809 4564 7813
rect 4568 7809 4569 7813
rect 4573 7809 4574 7813
rect 4578 7809 4579 7813
rect 4583 7809 4584 7813
rect 4588 7809 4589 7813
rect 4593 7809 4595 7813
rect 4527 7807 4595 7809
rect 4483 7789 4484 7793
rect 4488 7789 4489 7793
rect 4493 7789 4494 7793
rect 4498 7789 4499 7793
rect 4503 7789 4504 7793
rect 4508 7789 4509 7793
rect 4479 7788 4513 7789
rect 4483 7784 4484 7788
rect 4488 7784 4489 7788
rect 4493 7784 4494 7788
rect 4498 7784 4499 7788
rect 4503 7784 4504 7788
rect 4508 7784 4509 7788
rect 4479 7783 4513 7784
rect 4483 7779 4484 7783
rect 4488 7779 4489 7783
rect 4493 7779 4494 7783
rect 4498 7779 4499 7783
rect 4503 7779 4504 7783
rect 4508 7779 4509 7783
rect 4479 7778 4513 7779
rect 4483 7774 4484 7778
rect 4488 7774 4489 7778
rect 4493 7774 4494 7778
rect 4498 7774 4499 7778
rect 4503 7774 4504 7778
rect 4508 7774 4509 7778
rect 4529 7789 4530 7793
rect 4534 7789 4535 7793
rect 4539 7789 4540 7793
rect 4544 7789 4545 7793
rect 4549 7789 4550 7793
rect 4554 7789 4555 7793
rect 4525 7788 4559 7789
rect 4529 7784 4530 7788
rect 4534 7784 4535 7788
rect 4539 7784 4540 7788
rect 4544 7784 4545 7788
rect 4549 7784 4550 7788
rect 4554 7784 4555 7788
rect 4525 7783 4559 7784
rect 4529 7779 4530 7783
rect 4534 7779 4535 7783
rect 4539 7779 4540 7783
rect 4544 7779 4545 7783
rect 4549 7779 4550 7783
rect 4554 7779 4555 7783
rect 4525 7778 4559 7779
rect 4529 7774 4530 7778
rect 4534 7774 4535 7778
rect 4539 7774 4540 7778
rect 4544 7774 4545 7778
rect 4549 7774 4550 7778
rect 4554 7774 4555 7778
rect 4826 7772 5086 7775
rect 4222 7739 4223 7742
rect 3781 7381 3787 7732
rect 4087 7629 4091 7711
rect 4102 7708 4105 7718
rect 4109 7678 4112 7687
rect 4125 7680 4128 7693
rect 4138 7665 4141 7718
rect 4205 7708 4208 7718
rect 4145 7693 4149 7697
rect 4146 7678 4149 7687
rect 4101 7651 4104 7663
rect 4142 7661 4143 7665
rect 4152 7651 4155 7704
rect 4220 7693 4223 7739
rect 4158 7684 4161 7689
rect 4167 7678 4170 7687
rect 4183 7680 4186 7693
rect 4204 7678 4207 7687
rect 4220 7678 4223 7687
rect 4203 7651 4206 7661
rect 4220 7644 4223 7674
rect 4095 7602 4098 7639
rect 4102 7622 4105 7632
rect 4109 7592 4112 7601
rect 4125 7594 4128 7607
rect 4138 7579 4141 7632
rect 4205 7622 4208 7632
rect 4145 7607 4149 7611
rect 4146 7592 4149 7601
rect 4101 7565 4104 7577
rect 4142 7575 4143 7579
rect 4152 7565 4155 7618
rect 4158 7598 4161 7603
rect 4167 7592 4170 7601
rect 4183 7594 4186 7607
rect 4204 7592 4207 7601
rect 4220 7602 4223 7603
rect 4241 7605 4245 7747
rect 4220 7597 4223 7598
rect 4203 7565 4206 7575
rect 4241 7503 4245 7585
rect 4826 7518 4829 7772
rect 5083 7518 5086 7772
rect 4826 7515 5086 7518
rect 4826 7462 5086 7465
rect 4826 7208 4829 7462
rect 5083 7208 5086 7462
rect 86 7193 346 7196
rect 4483 7202 4484 7206
rect 4488 7202 4489 7206
rect 4493 7202 4494 7206
rect 4498 7202 4499 7206
rect 4503 7202 4504 7206
rect 4508 7202 4509 7206
rect 4479 7201 4513 7202
rect 4483 7197 4484 7201
rect 4488 7197 4489 7201
rect 4493 7197 4494 7201
rect 4498 7197 4499 7201
rect 4503 7197 4504 7201
rect 4508 7197 4509 7201
rect 4479 7196 4513 7197
rect 4483 7192 4484 7196
rect 4488 7192 4489 7196
rect 4493 7192 4494 7196
rect 4498 7192 4499 7196
rect 4503 7192 4504 7196
rect 4508 7192 4509 7196
rect 4479 7191 4513 7192
rect 4483 7187 4484 7191
rect 4488 7187 4489 7191
rect 4493 7187 4494 7191
rect 4498 7187 4499 7191
rect 4503 7187 4504 7191
rect 4508 7187 4509 7191
rect 4529 7202 4530 7206
rect 4534 7202 4535 7206
rect 4539 7202 4540 7206
rect 4544 7202 4545 7206
rect 4549 7202 4550 7206
rect 4554 7202 4555 7206
rect 4826 7205 5086 7208
rect 4525 7201 4559 7202
rect 4529 7197 4530 7201
rect 4534 7197 4535 7201
rect 4539 7197 4540 7201
rect 4544 7197 4545 7201
rect 4549 7197 4550 7201
rect 4554 7197 4555 7201
rect 4525 7196 4559 7197
rect 4529 7192 4530 7196
rect 4534 7192 4535 7196
rect 4539 7192 4540 7196
rect 4544 7192 4545 7196
rect 4549 7192 4550 7196
rect 4554 7192 4555 7196
rect 4525 7191 4559 7192
rect 4529 7187 4530 7191
rect 4534 7187 4535 7191
rect 4539 7187 4540 7191
rect 4544 7187 4545 7191
rect 4549 7187 4550 7191
rect 4554 7187 4555 7191
rect 617 7158 618 7162
rect 622 7158 623 7162
rect 627 7158 628 7162
rect 632 7158 633 7162
rect 637 7158 638 7162
rect 642 7158 643 7162
rect 613 7157 647 7158
rect 617 7153 618 7157
rect 622 7153 623 7157
rect 627 7153 628 7157
rect 632 7153 633 7157
rect 637 7153 638 7157
rect 642 7153 643 7157
rect 613 7152 647 7153
rect 617 7148 618 7152
rect 622 7148 623 7152
rect 627 7148 628 7152
rect 632 7148 633 7152
rect 637 7148 638 7152
rect 642 7148 643 7152
rect 613 7147 647 7148
rect 86 7141 346 7144
rect 617 7143 618 7147
rect 622 7143 623 7147
rect 627 7143 628 7147
rect 632 7143 633 7147
rect 637 7143 638 7147
rect 642 7143 643 7147
rect 663 7158 664 7162
rect 668 7158 669 7162
rect 673 7158 674 7162
rect 678 7158 679 7162
rect 683 7158 684 7162
rect 688 7158 689 7162
rect 659 7157 693 7158
rect 663 7153 664 7157
rect 668 7153 669 7157
rect 673 7153 674 7157
rect 678 7153 679 7157
rect 683 7153 684 7157
rect 688 7153 689 7157
rect 659 7152 693 7153
rect 663 7148 664 7152
rect 668 7148 669 7152
rect 673 7148 674 7152
rect 678 7148 679 7152
rect 683 7148 684 7152
rect 688 7148 689 7152
rect 659 7147 693 7148
rect 663 7143 664 7147
rect 668 7143 669 7147
rect 673 7143 674 7147
rect 678 7143 679 7147
rect 683 7143 684 7147
rect 688 7143 689 7147
rect 4826 7153 5086 7156
rect 86 6887 89 7141
rect 343 6887 346 7141
rect 4826 6899 4829 7153
rect 5083 6899 5086 7153
rect 86 6884 346 6887
rect 4483 6893 4484 6897
rect 4488 6893 4489 6897
rect 4493 6893 4494 6897
rect 4498 6893 4499 6897
rect 4503 6893 4504 6897
rect 4508 6893 4509 6897
rect 4479 6892 4513 6893
rect 4483 6888 4484 6892
rect 4488 6888 4489 6892
rect 4493 6888 4494 6892
rect 4498 6888 4499 6892
rect 4503 6888 4504 6892
rect 4508 6888 4509 6892
rect 4479 6887 4513 6888
rect 4483 6883 4484 6887
rect 4488 6883 4489 6887
rect 4493 6883 4494 6887
rect 4498 6883 4499 6887
rect 4503 6883 4504 6887
rect 4508 6883 4509 6887
rect 4479 6882 4513 6883
rect 4483 6878 4484 6882
rect 4488 6878 4489 6882
rect 4493 6878 4494 6882
rect 4498 6878 4499 6882
rect 4503 6878 4504 6882
rect 4508 6878 4509 6882
rect 4529 6893 4530 6897
rect 4534 6893 4535 6897
rect 4539 6893 4540 6897
rect 4544 6893 4545 6897
rect 4549 6893 4550 6897
rect 4554 6893 4555 6897
rect 4826 6896 5086 6899
rect 4525 6892 4559 6893
rect 4529 6888 4530 6892
rect 4534 6888 4535 6892
rect 4539 6888 4540 6892
rect 4544 6888 4545 6892
rect 4549 6888 4550 6892
rect 4554 6888 4555 6892
rect 4525 6887 4559 6888
rect 4529 6883 4530 6887
rect 4534 6883 4535 6887
rect 4539 6883 4540 6887
rect 4544 6883 4545 6887
rect 4549 6883 4550 6887
rect 4554 6883 4555 6887
rect 4525 6882 4559 6883
rect 4529 6878 4530 6882
rect 4534 6878 4535 6882
rect 4539 6878 4540 6882
rect 4544 6878 4545 6882
rect 4549 6878 4550 6882
rect 4554 6878 4555 6882
rect 617 6849 618 6853
rect 622 6849 623 6853
rect 627 6849 628 6853
rect 632 6849 633 6853
rect 637 6849 638 6853
rect 642 6849 643 6853
rect 613 6848 647 6849
rect 617 6844 618 6848
rect 622 6844 623 6848
rect 627 6844 628 6848
rect 632 6844 633 6848
rect 637 6844 638 6848
rect 642 6844 643 6848
rect 613 6843 647 6844
rect 617 6839 618 6843
rect 622 6839 623 6843
rect 627 6839 628 6843
rect 632 6839 633 6843
rect 637 6839 638 6843
rect 642 6839 643 6843
rect 613 6838 647 6839
rect 86 6832 346 6835
rect 617 6834 618 6838
rect 622 6834 623 6838
rect 627 6834 628 6838
rect 632 6834 633 6838
rect 637 6834 638 6838
rect 642 6834 643 6838
rect 663 6849 664 6853
rect 668 6849 669 6853
rect 673 6849 674 6853
rect 678 6849 679 6853
rect 683 6849 684 6853
rect 688 6849 689 6853
rect 659 6848 693 6849
rect 663 6844 664 6848
rect 668 6844 669 6848
rect 673 6844 674 6848
rect 678 6844 679 6848
rect 683 6844 684 6848
rect 688 6844 689 6848
rect 659 6843 693 6844
rect 663 6839 664 6843
rect 668 6839 669 6843
rect 673 6839 674 6843
rect 678 6839 679 6843
rect 683 6839 684 6843
rect 688 6839 689 6843
rect 659 6838 693 6839
rect 663 6834 664 6838
rect 668 6834 669 6838
rect 673 6834 674 6838
rect 678 6834 679 6838
rect 683 6834 684 6838
rect 688 6834 689 6838
rect 4826 6844 5086 6847
rect 86 6578 89 6832
rect 343 6578 346 6832
rect 4826 6590 4829 6844
rect 5083 6590 5086 6844
rect 86 6575 346 6578
rect 4483 6584 4484 6588
rect 4488 6584 4489 6588
rect 4493 6584 4494 6588
rect 4498 6584 4499 6588
rect 4503 6584 4504 6588
rect 4508 6584 4509 6588
rect 4479 6583 4513 6584
rect 4483 6579 4484 6583
rect 4488 6579 4489 6583
rect 4493 6579 4494 6583
rect 4498 6579 4499 6583
rect 4503 6579 4504 6583
rect 4508 6579 4509 6583
rect 4479 6578 4513 6579
rect 4483 6574 4484 6578
rect 4488 6574 4489 6578
rect 4493 6574 4494 6578
rect 4498 6574 4499 6578
rect 4503 6574 4504 6578
rect 4508 6574 4509 6578
rect 4479 6573 4513 6574
rect 4483 6569 4484 6573
rect 4488 6569 4489 6573
rect 4493 6569 4494 6573
rect 4498 6569 4499 6573
rect 4503 6569 4504 6573
rect 4508 6569 4509 6573
rect 4529 6584 4530 6588
rect 4534 6584 4535 6588
rect 4539 6584 4540 6588
rect 4544 6584 4545 6588
rect 4549 6584 4550 6588
rect 4554 6584 4555 6588
rect 4826 6587 5086 6590
rect 4525 6583 4559 6584
rect 4529 6579 4530 6583
rect 4534 6579 4535 6583
rect 4539 6579 4540 6583
rect 4544 6579 4545 6583
rect 4549 6579 4550 6583
rect 4554 6579 4555 6583
rect 4525 6578 4559 6579
rect 4529 6574 4530 6578
rect 4534 6574 4535 6578
rect 4539 6574 4540 6578
rect 4544 6574 4545 6578
rect 4549 6574 4550 6578
rect 4554 6574 4555 6578
rect 4525 6573 4559 6574
rect 4529 6569 4530 6573
rect 4534 6569 4535 6573
rect 4539 6569 4540 6573
rect 4544 6569 4545 6573
rect 4549 6569 4550 6573
rect 4554 6569 4555 6573
rect 617 6540 618 6544
rect 622 6540 623 6544
rect 627 6540 628 6544
rect 632 6540 633 6544
rect 637 6540 638 6544
rect 642 6540 643 6544
rect 613 6539 647 6540
rect 617 6535 618 6539
rect 622 6535 623 6539
rect 627 6535 628 6539
rect 632 6535 633 6539
rect 637 6535 638 6539
rect 642 6535 643 6539
rect 613 6534 647 6535
rect 617 6530 618 6534
rect 622 6530 623 6534
rect 627 6530 628 6534
rect 632 6530 633 6534
rect 637 6530 638 6534
rect 642 6530 643 6534
rect 613 6529 647 6530
rect 86 6523 346 6526
rect 617 6525 618 6529
rect 622 6525 623 6529
rect 627 6525 628 6529
rect 632 6525 633 6529
rect 637 6525 638 6529
rect 642 6525 643 6529
rect 663 6540 664 6544
rect 668 6540 669 6544
rect 673 6540 674 6544
rect 678 6540 679 6544
rect 683 6540 684 6544
rect 688 6540 689 6544
rect 659 6539 693 6540
rect 663 6535 664 6539
rect 668 6535 669 6539
rect 673 6535 674 6539
rect 678 6535 679 6539
rect 683 6535 684 6539
rect 688 6535 689 6539
rect 659 6534 693 6535
rect 663 6530 664 6534
rect 668 6530 669 6534
rect 673 6530 674 6534
rect 678 6530 679 6534
rect 683 6530 684 6534
rect 688 6530 689 6534
rect 659 6529 693 6530
rect 663 6525 664 6529
rect 668 6525 669 6529
rect 673 6525 674 6529
rect 678 6525 679 6529
rect 683 6525 684 6529
rect 688 6525 689 6529
rect 4826 6535 5086 6538
rect 86 6269 89 6523
rect 343 6269 346 6523
rect 4826 6281 4829 6535
rect 5083 6281 5086 6535
rect 86 6266 346 6269
rect 4483 6275 4484 6279
rect 4488 6275 4489 6279
rect 4493 6275 4494 6279
rect 4498 6275 4499 6279
rect 4503 6275 4504 6279
rect 4508 6275 4509 6279
rect 4479 6274 4513 6275
rect 4483 6270 4484 6274
rect 4488 6270 4489 6274
rect 4493 6270 4494 6274
rect 4498 6270 4499 6274
rect 4503 6270 4504 6274
rect 4508 6270 4509 6274
rect 4479 6269 4513 6270
rect 4483 6265 4484 6269
rect 4488 6265 4489 6269
rect 4493 6265 4494 6269
rect 4498 6265 4499 6269
rect 4503 6265 4504 6269
rect 4508 6265 4509 6269
rect 4479 6264 4513 6265
rect 4483 6260 4484 6264
rect 4488 6260 4489 6264
rect 4493 6260 4494 6264
rect 4498 6260 4499 6264
rect 4503 6260 4504 6264
rect 4508 6260 4509 6264
rect 4529 6275 4530 6279
rect 4534 6275 4535 6279
rect 4539 6275 4540 6279
rect 4544 6275 4545 6279
rect 4549 6275 4550 6279
rect 4554 6275 4555 6279
rect 4826 6278 5086 6281
rect 4525 6274 4559 6275
rect 4529 6270 4530 6274
rect 4534 6270 4535 6274
rect 4539 6270 4540 6274
rect 4544 6270 4545 6274
rect 4549 6270 4550 6274
rect 4554 6270 4555 6274
rect 4525 6269 4559 6270
rect 4529 6265 4530 6269
rect 4534 6265 4535 6269
rect 4539 6265 4540 6269
rect 4544 6265 4545 6269
rect 4549 6265 4550 6269
rect 4554 6265 4555 6269
rect 4525 6264 4559 6265
rect 4529 6260 4530 6264
rect 4534 6260 4535 6264
rect 4539 6260 4540 6264
rect 4544 6260 4545 6264
rect 4549 6260 4550 6264
rect 4554 6260 4555 6264
rect 99 5800 593 6231
rect 617 6140 618 6144
rect 622 6140 623 6144
rect 627 6140 628 6144
rect 632 6140 633 6144
rect 637 6140 638 6144
rect 642 6140 643 6144
rect 613 6139 647 6140
rect 617 6135 618 6139
rect 622 6135 623 6139
rect 627 6135 628 6139
rect 632 6135 633 6139
rect 637 6135 638 6139
rect 642 6135 643 6139
rect 613 6134 647 6135
rect 617 6130 618 6134
rect 622 6130 623 6134
rect 627 6130 628 6134
rect 632 6130 633 6134
rect 637 6130 638 6134
rect 642 6130 643 6134
rect 613 6129 647 6130
rect 617 6125 618 6129
rect 622 6125 623 6129
rect 627 6125 628 6129
rect 632 6125 633 6129
rect 637 6125 638 6129
rect 642 6125 643 6129
rect 663 6140 664 6144
rect 668 6140 669 6144
rect 673 6140 674 6144
rect 678 6140 679 6144
rect 683 6140 684 6144
rect 688 6140 689 6144
rect 659 6139 693 6140
rect 663 6135 664 6139
rect 668 6135 669 6139
rect 673 6135 674 6139
rect 678 6135 679 6139
rect 683 6135 684 6139
rect 688 6135 689 6139
rect 659 6134 693 6135
rect 663 6130 664 6134
rect 668 6130 669 6134
rect 673 6130 674 6134
rect 678 6130 679 6134
rect 683 6130 684 6134
rect 688 6130 689 6134
rect 659 6129 693 6130
rect 663 6125 664 6129
rect 668 6125 669 6129
rect 673 6125 674 6129
rect 678 6125 679 6129
rect 683 6125 684 6129
rect 688 6125 689 6129
rect 617 6111 618 6115
rect 622 6111 623 6115
rect 627 6111 628 6115
rect 632 6111 633 6115
rect 637 6111 638 6115
rect 642 6111 643 6115
rect 613 6110 647 6111
rect 617 6106 618 6110
rect 622 6106 623 6110
rect 627 6106 628 6110
rect 632 6106 633 6110
rect 637 6106 638 6110
rect 642 6106 643 6110
rect 613 6105 647 6106
rect 617 6101 618 6105
rect 622 6101 623 6105
rect 627 6101 628 6105
rect 632 6101 633 6105
rect 637 6101 638 6105
rect 642 6101 643 6105
rect 613 6100 647 6101
rect 617 6096 618 6100
rect 622 6096 623 6100
rect 627 6096 628 6100
rect 632 6096 633 6100
rect 637 6096 638 6100
rect 642 6096 643 6100
rect 663 6111 664 6115
rect 668 6111 669 6115
rect 673 6111 674 6115
rect 678 6111 679 6115
rect 683 6111 684 6115
rect 688 6111 689 6115
rect 659 6110 693 6111
rect 663 6106 664 6110
rect 668 6106 669 6110
rect 673 6106 674 6110
rect 678 6106 679 6110
rect 683 6106 684 6110
rect 688 6106 689 6110
rect 659 6105 693 6106
rect 663 6101 664 6105
rect 668 6101 669 6105
rect 673 6101 674 6105
rect 678 6101 679 6105
rect 683 6101 684 6105
rect 688 6101 689 6105
rect 659 6100 693 6101
rect 663 6096 664 6100
rect 668 6096 669 6100
rect 673 6096 674 6100
rect 678 6096 679 6100
rect 683 6096 684 6100
rect 688 6096 689 6100
rect 617 6082 618 6086
rect 622 6082 623 6086
rect 627 6082 628 6086
rect 632 6082 633 6086
rect 637 6082 638 6086
rect 642 6082 643 6086
rect 613 6081 647 6082
rect 617 6077 618 6081
rect 622 6077 623 6081
rect 627 6077 628 6081
rect 632 6077 633 6081
rect 637 6077 638 6081
rect 642 6077 643 6081
rect 613 6076 647 6077
rect 617 6072 618 6076
rect 622 6072 623 6076
rect 627 6072 628 6076
rect 632 6072 633 6076
rect 637 6072 638 6076
rect 642 6072 643 6076
rect 613 6071 647 6072
rect 617 6067 618 6071
rect 622 6067 623 6071
rect 627 6067 628 6071
rect 632 6067 633 6071
rect 637 6067 638 6071
rect 642 6067 643 6071
rect 663 6082 664 6086
rect 668 6082 669 6086
rect 673 6082 674 6086
rect 678 6082 679 6086
rect 683 6082 684 6086
rect 688 6082 689 6086
rect 659 6081 693 6082
rect 663 6077 664 6081
rect 668 6077 669 6081
rect 673 6077 674 6081
rect 678 6077 679 6081
rect 683 6077 684 6081
rect 688 6077 689 6081
rect 659 6076 693 6077
rect 663 6072 664 6076
rect 668 6072 669 6076
rect 673 6072 674 6076
rect 678 6072 679 6076
rect 683 6072 684 6076
rect 688 6072 689 6076
rect 659 6071 693 6072
rect 663 6067 664 6071
rect 668 6067 669 6071
rect 673 6067 674 6071
rect 678 6067 679 6071
rect 683 6067 684 6071
rect 688 6067 689 6071
rect 4483 6083 4484 6087
rect 4488 6083 4489 6087
rect 4493 6083 4494 6087
rect 4498 6083 4499 6087
rect 4503 6083 4504 6087
rect 4508 6083 4509 6087
rect 4479 6082 4513 6083
rect 4483 6078 4484 6082
rect 4488 6078 4489 6082
rect 4493 6078 4494 6082
rect 4498 6078 4499 6082
rect 4503 6078 4504 6082
rect 4508 6078 4509 6082
rect 4479 6077 4513 6078
rect 4483 6073 4484 6077
rect 4488 6073 4489 6077
rect 4493 6073 4494 6077
rect 4498 6073 4499 6077
rect 4503 6073 4504 6077
rect 4508 6073 4509 6077
rect 4479 6072 4513 6073
rect 4483 6068 4484 6072
rect 4488 6068 4489 6072
rect 4493 6068 4494 6072
rect 4498 6068 4499 6072
rect 4503 6068 4504 6072
rect 4508 6068 4509 6072
rect 4529 6083 4530 6087
rect 4534 6083 4535 6087
rect 4539 6083 4540 6087
rect 4544 6083 4545 6087
rect 4549 6083 4550 6087
rect 4554 6083 4555 6087
rect 4525 6082 4559 6083
rect 4529 6078 4530 6082
rect 4534 6078 4535 6082
rect 4539 6078 4540 6082
rect 4544 6078 4545 6082
rect 4549 6078 4550 6082
rect 4554 6078 4555 6082
rect 4525 6077 4559 6078
rect 4529 6073 4530 6077
rect 4534 6073 4535 6077
rect 4539 6073 4540 6077
rect 4544 6073 4545 6077
rect 4549 6073 4550 6077
rect 4554 6073 4555 6077
rect 4525 6072 4559 6073
rect 4529 6068 4530 6072
rect 4534 6068 4535 6072
rect 4539 6068 4540 6072
rect 4544 6068 4545 6072
rect 4549 6068 4550 6072
rect 4554 6068 4555 6072
rect 4483 6057 4484 6061
rect 4488 6057 4489 6061
rect 4493 6057 4494 6061
rect 4498 6057 4499 6061
rect 4503 6057 4504 6061
rect 4508 6057 4509 6061
rect 617 6053 618 6057
rect 622 6053 623 6057
rect 627 6053 628 6057
rect 632 6053 633 6057
rect 637 6053 638 6057
rect 642 6053 643 6057
rect 613 6052 647 6053
rect 617 6048 618 6052
rect 622 6048 623 6052
rect 627 6048 628 6052
rect 632 6048 633 6052
rect 637 6048 638 6052
rect 642 6048 643 6052
rect 613 6047 647 6048
rect 617 6043 618 6047
rect 622 6043 623 6047
rect 627 6043 628 6047
rect 632 6043 633 6047
rect 637 6043 638 6047
rect 642 6043 643 6047
rect 613 6042 647 6043
rect 617 6038 618 6042
rect 622 6038 623 6042
rect 627 6038 628 6042
rect 632 6038 633 6042
rect 637 6038 638 6042
rect 642 6038 643 6042
rect 663 6053 664 6057
rect 668 6053 669 6057
rect 673 6053 674 6057
rect 678 6053 679 6057
rect 683 6053 684 6057
rect 688 6053 689 6057
rect 659 6052 693 6053
rect 663 6048 664 6052
rect 668 6048 669 6052
rect 673 6048 674 6052
rect 678 6048 679 6052
rect 683 6048 684 6052
rect 688 6048 689 6052
rect 659 6047 693 6048
rect 663 6043 664 6047
rect 668 6043 669 6047
rect 673 6043 674 6047
rect 678 6043 679 6047
rect 683 6043 684 6047
rect 688 6043 689 6047
rect 659 6042 693 6043
rect 4479 6056 4513 6057
rect 4483 6052 4484 6056
rect 4488 6052 4489 6056
rect 4493 6052 4494 6056
rect 4498 6052 4499 6056
rect 4503 6052 4504 6056
rect 4508 6052 4509 6056
rect 4479 6051 4513 6052
rect 4483 6047 4484 6051
rect 4488 6047 4489 6051
rect 4493 6047 4494 6051
rect 4498 6047 4499 6051
rect 4503 6047 4504 6051
rect 4508 6047 4509 6051
rect 4479 6046 4513 6047
rect 4483 6042 4484 6046
rect 4488 6042 4489 6046
rect 4493 6042 4494 6046
rect 4498 6042 4499 6046
rect 4503 6042 4504 6046
rect 4508 6042 4509 6046
rect 4529 6057 4530 6061
rect 4534 6057 4535 6061
rect 4539 6057 4540 6061
rect 4544 6057 4545 6061
rect 4549 6057 4550 6061
rect 4554 6057 4555 6061
rect 4525 6056 4559 6057
rect 4529 6052 4530 6056
rect 4534 6052 4535 6056
rect 4539 6052 4540 6056
rect 4544 6052 4545 6056
rect 4549 6052 4550 6056
rect 4554 6052 4555 6056
rect 4525 6051 4559 6052
rect 4529 6047 4530 6051
rect 4534 6047 4535 6051
rect 4539 6047 4540 6051
rect 4544 6047 4545 6051
rect 4549 6047 4550 6051
rect 4554 6047 4555 6051
rect 4525 6046 4559 6047
rect 4529 6042 4530 6046
rect 4534 6042 4535 6046
rect 4539 6042 4540 6046
rect 4544 6042 4545 6046
rect 4549 6042 4550 6046
rect 4554 6042 4555 6046
rect 663 6038 664 6042
rect 668 6038 669 6042
rect 673 6038 674 6042
rect 678 6038 679 6042
rect 683 6038 684 6042
rect 688 6038 689 6042
rect 4483 6031 4484 6035
rect 4488 6031 4489 6035
rect 4493 6031 4494 6035
rect 4498 6031 4499 6035
rect 4503 6031 4504 6035
rect 4508 6031 4509 6035
rect 4479 6030 4513 6031
rect 617 6024 618 6028
rect 622 6024 623 6028
rect 627 6024 628 6028
rect 632 6024 633 6028
rect 637 6024 638 6028
rect 642 6024 643 6028
rect 613 6023 647 6024
rect 617 6019 618 6023
rect 622 6019 623 6023
rect 627 6019 628 6023
rect 632 6019 633 6023
rect 637 6019 638 6023
rect 642 6019 643 6023
rect 613 6018 647 6019
rect 617 6014 618 6018
rect 622 6014 623 6018
rect 627 6014 628 6018
rect 632 6014 633 6018
rect 637 6014 638 6018
rect 642 6014 643 6018
rect 613 6013 647 6014
rect 617 6009 618 6013
rect 622 6009 623 6013
rect 627 6009 628 6013
rect 632 6009 633 6013
rect 637 6009 638 6013
rect 642 6009 643 6013
rect 663 6024 664 6028
rect 668 6024 669 6028
rect 673 6024 674 6028
rect 678 6024 679 6028
rect 683 6024 684 6028
rect 688 6024 689 6028
rect 659 6023 693 6024
rect 663 6019 664 6023
rect 668 6019 669 6023
rect 673 6019 674 6023
rect 678 6019 679 6023
rect 683 6019 684 6023
rect 688 6019 689 6023
rect 659 6018 693 6019
rect 663 6014 664 6018
rect 668 6014 669 6018
rect 673 6014 674 6018
rect 678 6014 679 6018
rect 683 6014 684 6018
rect 688 6014 689 6018
rect 4483 6026 4484 6030
rect 4488 6026 4489 6030
rect 4493 6026 4494 6030
rect 4498 6026 4499 6030
rect 4503 6026 4504 6030
rect 4508 6026 4509 6030
rect 4479 6025 4513 6026
rect 4483 6021 4484 6025
rect 4488 6021 4489 6025
rect 4493 6021 4494 6025
rect 4498 6021 4499 6025
rect 4503 6021 4504 6025
rect 4508 6021 4509 6025
rect 4479 6020 4513 6021
rect 4483 6016 4484 6020
rect 4488 6016 4489 6020
rect 4493 6016 4494 6020
rect 4498 6016 4499 6020
rect 4503 6016 4504 6020
rect 4508 6016 4509 6020
rect 4529 6031 4530 6035
rect 4534 6031 4535 6035
rect 4539 6031 4540 6035
rect 4544 6031 4545 6035
rect 4549 6031 4550 6035
rect 4554 6031 4555 6035
rect 4525 6030 4559 6031
rect 4529 6026 4530 6030
rect 4534 6026 4535 6030
rect 4539 6026 4540 6030
rect 4544 6026 4545 6030
rect 4549 6026 4550 6030
rect 4554 6026 4555 6030
rect 4525 6025 4559 6026
rect 4529 6021 4530 6025
rect 4534 6021 4535 6025
rect 4539 6021 4540 6025
rect 4544 6021 4545 6025
rect 4549 6021 4550 6025
rect 4554 6021 4555 6025
rect 4525 6020 4559 6021
rect 4529 6016 4530 6020
rect 4534 6016 4535 6020
rect 4539 6016 4540 6020
rect 4544 6016 4545 6020
rect 4549 6016 4550 6020
rect 4554 6016 4555 6020
rect 659 6013 693 6014
rect 663 6009 664 6013
rect 668 6009 669 6013
rect 673 6009 674 6013
rect 678 6009 679 6013
rect 683 6009 684 6013
rect 688 6009 689 6013
rect 4483 6005 4484 6009
rect 4488 6005 4489 6009
rect 4493 6005 4494 6009
rect 4498 6005 4499 6009
rect 4503 6005 4504 6009
rect 4508 6005 4509 6009
rect 4479 6004 4513 6005
rect 4483 6000 4484 6004
rect 4488 6000 4489 6004
rect 4493 6000 4494 6004
rect 4498 6000 4499 6004
rect 4503 6000 4504 6004
rect 4508 6000 4509 6004
rect 4479 5999 4513 6000
rect 4483 5995 4484 5999
rect 4488 5995 4489 5999
rect 4493 5995 4494 5999
rect 4498 5995 4499 5999
rect 4503 5995 4504 5999
rect 4508 5995 4509 5999
rect 4479 5994 4513 5995
rect 4483 5990 4484 5994
rect 4488 5990 4489 5994
rect 4493 5990 4494 5994
rect 4498 5990 4499 5994
rect 4503 5990 4504 5994
rect 4508 5990 4509 5994
rect 4529 6005 4530 6009
rect 4534 6005 4535 6009
rect 4539 6005 4540 6009
rect 4544 6005 4545 6009
rect 4549 6005 4550 6009
rect 4554 6005 4555 6009
rect 4525 6004 4559 6005
rect 4529 6000 4530 6004
rect 4534 6000 4535 6004
rect 4539 6000 4540 6004
rect 4544 6000 4545 6004
rect 4549 6000 4550 6004
rect 4554 6000 4555 6004
rect 4525 5999 4559 6000
rect 4529 5995 4530 5999
rect 4534 5995 4535 5999
rect 4539 5995 4540 5999
rect 4544 5995 4545 5999
rect 4549 5995 4550 5999
rect 4554 5995 4555 5999
rect 4525 5994 4559 5995
rect 4529 5990 4530 5994
rect 4534 5990 4535 5994
rect 4539 5990 4540 5994
rect 4544 5990 4545 5994
rect 4549 5990 4550 5994
rect 4554 5990 4555 5994
rect 4483 5979 4484 5983
rect 4488 5979 4489 5983
rect 4493 5979 4494 5983
rect 4498 5979 4499 5983
rect 4503 5979 4504 5983
rect 4508 5979 4509 5983
rect 4479 5978 4513 5979
rect 4483 5974 4484 5978
rect 4488 5974 4489 5978
rect 4493 5974 4494 5978
rect 4498 5974 4499 5978
rect 4503 5974 4504 5978
rect 4508 5974 4509 5978
rect 4479 5973 4513 5974
rect 4483 5969 4484 5973
rect 4488 5969 4489 5973
rect 4493 5969 4494 5973
rect 4498 5969 4499 5973
rect 4503 5969 4504 5973
rect 4508 5969 4509 5973
rect 4479 5968 4513 5969
rect 4483 5964 4484 5968
rect 4488 5964 4489 5968
rect 4493 5964 4494 5968
rect 4498 5964 4499 5968
rect 4503 5964 4504 5968
rect 4508 5964 4509 5968
rect 4529 5979 4530 5983
rect 4534 5979 4535 5983
rect 4539 5979 4540 5983
rect 4544 5979 4545 5983
rect 4549 5979 4550 5983
rect 4554 5979 4555 5983
rect 4525 5978 4559 5979
rect 4529 5974 4530 5978
rect 4534 5974 4535 5978
rect 4539 5974 4540 5978
rect 4544 5974 4545 5978
rect 4549 5974 4550 5978
rect 4554 5974 4555 5978
rect 4525 5973 4559 5974
rect 4529 5969 4530 5973
rect 4534 5969 4535 5973
rect 4539 5969 4540 5973
rect 4544 5969 4545 5973
rect 4549 5969 4550 5973
rect 4554 5969 4555 5973
rect 4525 5968 4559 5969
rect 4529 5964 4530 5968
rect 4534 5964 4535 5968
rect 4539 5964 4540 5968
rect 4544 5964 4545 5968
rect 4549 5964 4550 5968
rect 4554 5964 4555 5968
rect 761 5896 762 5900
rect 766 5896 767 5900
rect 771 5896 772 5900
rect 757 5895 776 5896
rect 761 5891 762 5895
rect 766 5891 767 5895
rect 771 5891 772 5895
rect 757 5890 776 5891
rect 761 5886 762 5890
rect 766 5886 767 5890
rect 771 5886 772 5890
rect 757 5885 776 5886
rect 761 5881 762 5885
rect 766 5881 767 5885
rect 771 5881 772 5885
rect 757 5880 776 5881
rect 761 5876 762 5880
rect 766 5876 767 5880
rect 771 5876 772 5880
rect 757 5875 776 5876
rect 761 5871 762 5875
rect 766 5871 767 5875
rect 771 5871 772 5875
rect 757 5870 776 5871
rect 761 5866 762 5870
rect 766 5866 767 5870
rect 771 5866 772 5870
rect 787 5896 788 5900
rect 792 5896 793 5900
rect 797 5896 798 5900
rect 783 5895 802 5896
rect 787 5891 788 5895
rect 792 5891 793 5895
rect 797 5891 798 5895
rect 783 5890 802 5891
rect 787 5886 788 5890
rect 792 5886 793 5890
rect 797 5886 798 5890
rect 783 5885 802 5886
rect 787 5881 788 5885
rect 792 5881 793 5885
rect 797 5881 798 5885
rect 783 5880 802 5881
rect 787 5876 788 5880
rect 792 5876 793 5880
rect 797 5876 798 5880
rect 783 5875 802 5876
rect 787 5871 788 5875
rect 792 5871 793 5875
rect 797 5871 798 5875
rect 783 5870 802 5871
rect 787 5866 788 5870
rect 792 5866 793 5870
rect 797 5866 798 5870
rect 813 5896 814 5900
rect 818 5896 819 5900
rect 823 5896 824 5900
rect 809 5895 828 5896
rect 813 5891 814 5895
rect 818 5891 819 5895
rect 823 5891 824 5895
rect 809 5890 828 5891
rect 813 5886 814 5890
rect 818 5886 819 5890
rect 823 5886 824 5890
rect 809 5885 828 5886
rect 813 5881 814 5885
rect 818 5881 819 5885
rect 823 5881 824 5885
rect 809 5880 828 5881
rect 813 5876 814 5880
rect 818 5876 819 5880
rect 823 5876 824 5880
rect 809 5875 828 5876
rect 813 5871 814 5875
rect 818 5871 819 5875
rect 823 5871 824 5875
rect 809 5870 828 5871
rect 813 5866 814 5870
rect 818 5866 819 5870
rect 823 5866 824 5870
rect 839 5896 840 5900
rect 844 5896 845 5900
rect 849 5896 850 5900
rect 835 5895 854 5896
rect 839 5891 840 5895
rect 844 5891 845 5895
rect 849 5891 850 5895
rect 835 5890 854 5891
rect 839 5886 840 5890
rect 844 5886 845 5890
rect 849 5886 850 5890
rect 835 5885 854 5886
rect 839 5881 840 5885
rect 844 5881 845 5885
rect 849 5881 850 5885
rect 835 5880 854 5881
rect 839 5876 840 5880
rect 844 5876 845 5880
rect 849 5876 850 5880
rect 835 5875 854 5876
rect 839 5871 840 5875
rect 844 5871 845 5875
rect 849 5871 850 5875
rect 835 5870 854 5871
rect 839 5866 840 5870
rect 844 5866 845 5870
rect 849 5866 850 5870
rect 865 5896 866 5900
rect 870 5896 871 5900
rect 875 5896 876 5900
rect 861 5895 880 5896
rect 865 5891 866 5895
rect 870 5891 871 5895
rect 875 5891 876 5895
rect 861 5890 880 5891
rect 865 5886 866 5890
rect 870 5886 871 5890
rect 875 5886 876 5890
rect 861 5885 880 5886
rect 865 5881 866 5885
rect 870 5881 871 5885
rect 875 5881 876 5885
rect 861 5880 880 5881
rect 865 5876 866 5880
rect 870 5876 871 5880
rect 875 5876 876 5880
rect 861 5875 880 5876
rect 865 5871 866 5875
rect 870 5871 871 5875
rect 875 5871 876 5875
rect 861 5870 880 5871
rect 865 5866 866 5870
rect 870 5866 871 5870
rect 875 5866 876 5870
rect 1058 5896 1059 5900
rect 1063 5896 1064 5900
rect 1068 5896 1069 5900
rect 1054 5895 1073 5896
rect 1058 5891 1059 5895
rect 1063 5891 1064 5895
rect 1068 5891 1069 5895
rect 1054 5890 1073 5891
rect 1058 5886 1059 5890
rect 1063 5886 1064 5890
rect 1068 5886 1069 5890
rect 1054 5885 1073 5886
rect 1058 5881 1059 5885
rect 1063 5881 1064 5885
rect 1068 5881 1069 5885
rect 1054 5880 1073 5881
rect 1058 5876 1059 5880
rect 1063 5876 1064 5880
rect 1068 5876 1069 5880
rect 1054 5875 1073 5876
rect 1058 5871 1059 5875
rect 1063 5871 1064 5875
rect 1068 5871 1069 5875
rect 1054 5870 1073 5871
rect 1058 5866 1059 5870
rect 1063 5866 1064 5870
rect 1068 5866 1069 5870
rect 1367 5896 1368 5900
rect 1372 5896 1373 5900
rect 1377 5896 1378 5900
rect 1363 5895 1382 5896
rect 1367 5891 1368 5895
rect 1372 5891 1373 5895
rect 1377 5891 1378 5895
rect 1363 5890 1382 5891
rect 1367 5886 1368 5890
rect 1372 5886 1373 5890
rect 1377 5886 1378 5890
rect 1363 5885 1382 5886
rect 1367 5881 1368 5885
rect 1372 5881 1373 5885
rect 1377 5881 1378 5885
rect 1363 5880 1382 5881
rect 1367 5876 1368 5880
rect 1372 5876 1373 5880
rect 1377 5876 1378 5880
rect 1363 5875 1382 5876
rect 1367 5871 1368 5875
rect 1372 5871 1373 5875
rect 1377 5871 1378 5875
rect 1363 5870 1382 5871
rect 1367 5866 1368 5870
rect 1372 5866 1373 5870
rect 1377 5866 1378 5870
rect 1676 5896 1677 5900
rect 1681 5896 1682 5900
rect 1686 5896 1687 5900
rect 1672 5895 1691 5896
rect 1676 5891 1677 5895
rect 1681 5891 1682 5895
rect 1686 5891 1687 5895
rect 1672 5890 1691 5891
rect 1676 5886 1677 5890
rect 1681 5886 1682 5890
rect 1686 5886 1687 5890
rect 1672 5885 1691 5886
rect 1676 5881 1677 5885
rect 1681 5881 1682 5885
rect 1686 5881 1687 5885
rect 1672 5880 1691 5881
rect 1676 5876 1677 5880
rect 1681 5876 1682 5880
rect 1686 5876 1687 5880
rect 1672 5875 1691 5876
rect 1676 5871 1677 5875
rect 1681 5871 1682 5875
rect 1686 5871 1687 5875
rect 1672 5870 1691 5871
rect 1676 5866 1677 5870
rect 1681 5866 1682 5870
rect 1686 5866 1687 5870
rect 1985 5896 1986 5900
rect 1990 5896 1991 5900
rect 1995 5896 1996 5900
rect 1981 5895 2000 5896
rect 1985 5891 1986 5895
rect 1990 5891 1991 5895
rect 1995 5891 1996 5895
rect 1981 5890 2000 5891
rect 1985 5886 1986 5890
rect 1990 5886 1991 5890
rect 1995 5886 1996 5890
rect 1981 5885 2000 5886
rect 1985 5881 1986 5885
rect 1990 5881 1991 5885
rect 1995 5881 1996 5885
rect 1981 5880 2000 5881
rect 1985 5876 1986 5880
rect 1990 5876 1991 5880
rect 1995 5876 1996 5880
rect 1981 5875 2000 5876
rect 1985 5871 1986 5875
rect 1990 5871 1991 5875
rect 1995 5871 1996 5875
rect 1981 5870 2000 5871
rect 1985 5866 1986 5870
rect 1990 5866 1991 5870
rect 1995 5866 1996 5870
rect 2294 5896 2295 5900
rect 2299 5896 2300 5900
rect 2304 5896 2305 5900
rect 2290 5895 2309 5896
rect 2294 5891 2295 5895
rect 2299 5891 2300 5895
rect 2304 5891 2305 5895
rect 2290 5890 2309 5891
rect 2294 5886 2295 5890
rect 2299 5886 2300 5890
rect 2304 5886 2305 5890
rect 2290 5885 2309 5886
rect 2294 5881 2295 5885
rect 2299 5881 2300 5885
rect 2304 5881 2305 5885
rect 2290 5880 2309 5881
rect 2294 5876 2295 5880
rect 2299 5876 2300 5880
rect 2304 5876 2305 5880
rect 2290 5875 2309 5876
rect 2294 5871 2295 5875
rect 2299 5871 2300 5875
rect 2304 5871 2305 5875
rect 2290 5870 2309 5871
rect 2294 5866 2295 5870
rect 2299 5866 2300 5870
rect 2304 5866 2305 5870
rect 2603 5896 2604 5900
rect 2608 5896 2609 5900
rect 2613 5896 2614 5900
rect 2599 5895 2618 5896
rect 2603 5891 2604 5895
rect 2608 5891 2609 5895
rect 2613 5891 2614 5895
rect 2599 5890 2618 5891
rect 2603 5886 2604 5890
rect 2608 5886 2609 5890
rect 2613 5886 2614 5890
rect 2599 5885 2618 5886
rect 2603 5881 2604 5885
rect 2608 5881 2609 5885
rect 2613 5881 2614 5885
rect 2599 5880 2618 5881
rect 2603 5876 2604 5880
rect 2608 5876 2609 5880
rect 2613 5876 2614 5880
rect 2599 5875 2618 5876
rect 2603 5871 2604 5875
rect 2608 5871 2609 5875
rect 2613 5871 2614 5875
rect 2599 5870 2618 5871
rect 2603 5866 2604 5870
rect 2608 5866 2609 5870
rect 2613 5866 2614 5870
rect 2912 5896 2913 5900
rect 2917 5896 2918 5900
rect 2922 5896 2923 5900
rect 2908 5895 2927 5896
rect 2912 5891 2913 5895
rect 2917 5891 2918 5895
rect 2922 5891 2923 5895
rect 2908 5890 2927 5891
rect 2912 5886 2913 5890
rect 2917 5886 2918 5890
rect 2922 5886 2923 5890
rect 2908 5885 2927 5886
rect 2912 5881 2913 5885
rect 2917 5881 2918 5885
rect 2922 5881 2923 5885
rect 2908 5880 2927 5881
rect 2912 5876 2913 5880
rect 2917 5876 2918 5880
rect 2922 5876 2923 5880
rect 2908 5875 2927 5876
rect 2912 5871 2913 5875
rect 2917 5871 2918 5875
rect 2922 5871 2923 5875
rect 2908 5870 2927 5871
rect 2912 5866 2913 5870
rect 2917 5866 2918 5870
rect 2922 5866 2923 5870
rect 3221 5896 3222 5900
rect 3226 5896 3227 5900
rect 3231 5896 3232 5900
rect 3217 5895 3236 5896
rect 3221 5891 3222 5895
rect 3226 5891 3227 5895
rect 3231 5891 3232 5895
rect 3217 5890 3236 5891
rect 3221 5886 3222 5890
rect 3226 5886 3227 5890
rect 3231 5886 3232 5890
rect 3217 5885 3236 5886
rect 3221 5881 3222 5885
rect 3226 5881 3227 5885
rect 3231 5881 3232 5885
rect 3217 5880 3236 5881
rect 3221 5876 3222 5880
rect 3226 5876 3227 5880
rect 3231 5876 3232 5880
rect 3217 5875 3236 5876
rect 3221 5871 3222 5875
rect 3226 5871 3227 5875
rect 3231 5871 3232 5875
rect 3217 5870 3236 5871
rect 3221 5866 3222 5870
rect 3226 5866 3227 5870
rect 3231 5866 3232 5870
rect 3530 5896 3531 5900
rect 3535 5896 3536 5900
rect 3540 5896 3541 5900
rect 3526 5895 3545 5896
rect 3530 5891 3531 5895
rect 3535 5891 3536 5895
rect 3540 5891 3541 5895
rect 3526 5890 3545 5891
rect 3530 5886 3531 5890
rect 3535 5886 3536 5890
rect 3540 5886 3541 5890
rect 3526 5885 3545 5886
rect 3530 5881 3531 5885
rect 3535 5881 3536 5885
rect 3540 5881 3541 5885
rect 3526 5880 3545 5881
rect 3530 5876 3531 5880
rect 3535 5876 3536 5880
rect 3540 5876 3541 5880
rect 3526 5875 3545 5876
rect 3530 5871 3531 5875
rect 3535 5871 3536 5875
rect 3540 5871 3541 5875
rect 3526 5870 3545 5871
rect 3530 5866 3531 5870
rect 3535 5866 3536 5870
rect 3540 5866 3541 5870
rect 3839 5896 3840 5900
rect 3844 5896 3845 5900
rect 3849 5896 3850 5900
rect 3835 5895 3854 5896
rect 3839 5891 3840 5895
rect 3844 5891 3845 5895
rect 3849 5891 3850 5895
rect 3835 5890 3854 5891
rect 3839 5886 3840 5890
rect 3844 5886 3845 5890
rect 3849 5886 3850 5890
rect 3835 5885 3854 5886
rect 3839 5881 3840 5885
rect 3844 5881 3845 5885
rect 3849 5881 3850 5885
rect 3835 5880 3854 5881
rect 3839 5876 3840 5880
rect 3844 5876 3845 5880
rect 3849 5876 3850 5880
rect 3835 5875 3854 5876
rect 3839 5871 3840 5875
rect 3844 5871 3845 5875
rect 3849 5871 3850 5875
rect 3835 5870 3854 5871
rect 3839 5866 3840 5870
rect 3844 5866 3845 5870
rect 3849 5866 3850 5870
rect 4239 5896 4240 5900
rect 4244 5896 4245 5900
rect 4249 5896 4250 5900
rect 4235 5895 4254 5896
rect 4239 5891 4240 5895
rect 4244 5891 4245 5895
rect 4249 5891 4250 5895
rect 4235 5890 4254 5891
rect 4239 5886 4240 5890
rect 4244 5886 4245 5890
rect 4249 5886 4250 5890
rect 4235 5885 4254 5886
rect 4239 5881 4240 5885
rect 4244 5881 4245 5885
rect 4249 5881 4250 5885
rect 4235 5880 4254 5881
rect 4239 5876 4240 5880
rect 4244 5876 4245 5880
rect 4249 5876 4250 5880
rect 4235 5875 4254 5876
rect 4239 5871 4240 5875
rect 4244 5871 4245 5875
rect 4249 5871 4250 5875
rect 4235 5870 4254 5871
rect 4239 5866 4240 5870
rect 4244 5866 4245 5870
rect 4249 5866 4250 5870
rect 4268 5896 4269 5900
rect 4273 5896 4274 5900
rect 4278 5896 4279 5900
rect 4264 5895 4283 5896
rect 4268 5891 4269 5895
rect 4273 5891 4274 5895
rect 4278 5891 4279 5895
rect 4264 5890 4283 5891
rect 4268 5886 4269 5890
rect 4273 5886 4274 5890
rect 4278 5886 4279 5890
rect 4264 5885 4283 5886
rect 4268 5881 4269 5885
rect 4273 5881 4274 5885
rect 4278 5881 4279 5885
rect 4264 5880 4283 5881
rect 4268 5876 4269 5880
rect 4273 5876 4274 5880
rect 4278 5876 4279 5880
rect 4264 5875 4283 5876
rect 4268 5871 4269 5875
rect 4273 5871 4274 5875
rect 4278 5871 4279 5875
rect 4264 5870 4283 5871
rect 4268 5866 4269 5870
rect 4273 5866 4274 5870
rect 4278 5866 4279 5870
rect 4297 5896 4298 5900
rect 4302 5896 4303 5900
rect 4307 5896 4308 5900
rect 4293 5895 4312 5896
rect 4297 5891 4298 5895
rect 4302 5891 4303 5895
rect 4307 5891 4308 5895
rect 4293 5890 4312 5891
rect 4297 5886 4298 5890
rect 4302 5886 4303 5890
rect 4307 5886 4308 5890
rect 4293 5885 4312 5886
rect 4297 5881 4298 5885
rect 4302 5881 4303 5885
rect 4307 5881 4308 5885
rect 4293 5880 4312 5881
rect 4297 5876 4298 5880
rect 4302 5876 4303 5880
rect 4307 5876 4308 5880
rect 4293 5875 4312 5876
rect 4297 5871 4298 5875
rect 4302 5871 4303 5875
rect 4307 5871 4308 5875
rect 4293 5870 4312 5871
rect 4297 5866 4298 5870
rect 4302 5866 4303 5870
rect 4307 5866 4308 5870
rect 4326 5896 4327 5900
rect 4331 5896 4332 5900
rect 4336 5896 4337 5900
rect 4322 5895 4341 5896
rect 4326 5891 4327 5895
rect 4331 5891 4332 5895
rect 4336 5891 4337 5895
rect 4322 5890 4341 5891
rect 4326 5886 4327 5890
rect 4331 5886 4332 5890
rect 4336 5886 4337 5890
rect 4322 5885 4341 5886
rect 4326 5881 4327 5885
rect 4331 5881 4332 5885
rect 4336 5881 4337 5885
rect 4322 5880 4341 5881
rect 4326 5876 4327 5880
rect 4331 5876 4332 5880
rect 4336 5876 4337 5880
rect 4322 5875 4341 5876
rect 4326 5871 4327 5875
rect 4331 5871 4332 5875
rect 4336 5871 4337 5875
rect 4322 5870 4341 5871
rect 4326 5866 4327 5870
rect 4331 5866 4332 5870
rect 4336 5866 4337 5870
rect 4355 5896 4356 5900
rect 4360 5896 4361 5900
rect 4365 5896 4366 5900
rect 4351 5895 4370 5896
rect 4355 5891 4356 5895
rect 4360 5891 4361 5895
rect 4365 5891 4366 5895
rect 4351 5890 4370 5891
rect 4355 5886 4356 5890
rect 4360 5886 4361 5890
rect 4365 5886 4366 5890
rect 4351 5885 4370 5886
rect 4355 5881 4356 5885
rect 4360 5881 4361 5885
rect 4365 5881 4366 5885
rect 4351 5880 4370 5881
rect 4355 5876 4356 5880
rect 4360 5876 4361 5880
rect 4365 5876 4366 5880
rect 4351 5875 4370 5876
rect 4355 5871 4356 5875
rect 4360 5871 4361 5875
rect 4365 5871 4366 5875
rect 4351 5870 4370 5871
rect 4355 5866 4356 5870
rect 4360 5866 4361 5870
rect 4365 5866 4366 5870
rect 761 5850 762 5854
rect 766 5850 767 5854
rect 771 5850 772 5854
rect 757 5849 776 5850
rect 761 5845 762 5849
rect 766 5845 767 5849
rect 771 5845 772 5849
rect 757 5844 776 5845
rect 761 5840 762 5844
rect 766 5840 767 5844
rect 771 5840 772 5844
rect 757 5839 776 5840
rect 761 5835 762 5839
rect 766 5835 767 5839
rect 771 5835 772 5839
rect 757 5834 776 5835
rect 761 5830 762 5834
rect 766 5830 767 5834
rect 771 5830 772 5834
rect 757 5829 776 5830
rect 761 5825 762 5829
rect 766 5825 767 5829
rect 771 5825 772 5829
rect 757 5824 776 5825
rect 761 5820 762 5824
rect 766 5820 767 5824
rect 771 5820 772 5824
rect 787 5850 788 5854
rect 792 5850 793 5854
rect 797 5850 798 5854
rect 783 5849 802 5850
rect 787 5845 788 5849
rect 792 5845 793 5849
rect 797 5845 798 5849
rect 783 5844 802 5845
rect 787 5840 788 5844
rect 792 5840 793 5844
rect 797 5840 798 5844
rect 783 5839 802 5840
rect 787 5835 788 5839
rect 792 5835 793 5839
rect 797 5835 798 5839
rect 783 5834 802 5835
rect 787 5830 788 5834
rect 792 5830 793 5834
rect 797 5830 798 5834
rect 783 5829 802 5830
rect 787 5825 788 5829
rect 792 5825 793 5829
rect 797 5825 798 5829
rect 783 5824 802 5825
rect 787 5820 788 5824
rect 792 5820 793 5824
rect 797 5820 798 5824
rect 813 5850 814 5854
rect 818 5850 819 5854
rect 823 5850 824 5854
rect 809 5849 828 5850
rect 813 5845 814 5849
rect 818 5845 819 5849
rect 823 5845 824 5849
rect 809 5844 828 5845
rect 813 5840 814 5844
rect 818 5840 819 5844
rect 823 5840 824 5844
rect 809 5839 828 5840
rect 813 5835 814 5839
rect 818 5835 819 5839
rect 823 5835 824 5839
rect 809 5834 828 5835
rect 813 5830 814 5834
rect 818 5830 819 5834
rect 823 5830 824 5834
rect 809 5829 828 5830
rect 813 5825 814 5829
rect 818 5825 819 5829
rect 823 5825 824 5829
rect 809 5824 828 5825
rect 813 5820 814 5824
rect 818 5820 819 5824
rect 823 5820 824 5824
rect 839 5850 840 5854
rect 844 5850 845 5854
rect 849 5850 850 5854
rect 835 5849 854 5850
rect 839 5845 840 5849
rect 844 5845 845 5849
rect 849 5845 850 5849
rect 835 5844 854 5845
rect 839 5840 840 5844
rect 844 5840 845 5844
rect 849 5840 850 5844
rect 835 5839 854 5840
rect 839 5835 840 5839
rect 844 5835 845 5839
rect 849 5835 850 5839
rect 835 5834 854 5835
rect 839 5830 840 5834
rect 844 5830 845 5834
rect 849 5830 850 5834
rect 835 5829 854 5830
rect 839 5825 840 5829
rect 844 5825 845 5829
rect 849 5825 850 5829
rect 835 5824 854 5825
rect 839 5820 840 5824
rect 844 5820 845 5824
rect 849 5820 850 5824
rect 865 5850 866 5854
rect 870 5850 871 5854
rect 875 5850 876 5854
rect 861 5849 880 5850
rect 865 5845 866 5849
rect 870 5845 871 5849
rect 875 5845 876 5849
rect 861 5844 880 5845
rect 865 5840 866 5844
rect 870 5840 871 5844
rect 875 5840 876 5844
rect 861 5839 880 5840
rect 865 5835 866 5839
rect 870 5835 871 5839
rect 875 5835 876 5839
rect 861 5834 880 5835
rect 865 5830 866 5834
rect 870 5830 871 5834
rect 875 5830 876 5834
rect 861 5829 880 5830
rect 865 5825 866 5829
rect 870 5825 871 5829
rect 875 5825 876 5829
rect 861 5824 880 5825
rect 865 5820 866 5824
rect 870 5820 871 5824
rect 875 5820 876 5824
rect 1058 5850 1059 5854
rect 1063 5850 1064 5854
rect 1068 5850 1069 5854
rect 1054 5849 1073 5850
rect 1058 5845 1059 5849
rect 1063 5845 1064 5849
rect 1068 5845 1069 5849
rect 1054 5844 1073 5845
rect 1058 5840 1059 5844
rect 1063 5840 1064 5844
rect 1068 5840 1069 5844
rect 1054 5839 1073 5840
rect 1058 5835 1059 5839
rect 1063 5835 1064 5839
rect 1068 5835 1069 5839
rect 1054 5834 1073 5835
rect 1058 5830 1059 5834
rect 1063 5830 1064 5834
rect 1068 5830 1069 5834
rect 1054 5829 1073 5830
rect 1058 5825 1059 5829
rect 1063 5825 1064 5829
rect 1068 5825 1069 5829
rect 1054 5824 1073 5825
rect 1058 5820 1059 5824
rect 1063 5820 1064 5824
rect 1068 5820 1069 5824
rect 1367 5850 1368 5854
rect 1372 5850 1373 5854
rect 1377 5850 1378 5854
rect 1363 5849 1382 5850
rect 1367 5845 1368 5849
rect 1372 5845 1373 5849
rect 1377 5845 1378 5849
rect 1363 5844 1382 5845
rect 1367 5840 1368 5844
rect 1372 5840 1373 5844
rect 1377 5840 1378 5844
rect 1363 5839 1382 5840
rect 1367 5835 1368 5839
rect 1372 5835 1373 5839
rect 1377 5835 1378 5839
rect 1363 5834 1382 5835
rect 1367 5830 1368 5834
rect 1372 5830 1373 5834
rect 1377 5830 1378 5834
rect 1363 5829 1382 5830
rect 1367 5825 1368 5829
rect 1372 5825 1373 5829
rect 1377 5825 1378 5829
rect 1363 5824 1382 5825
rect 1367 5820 1368 5824
rect 1372 5820 1373 5824
rect 1377 5820 1378 5824
rect 1676 5850 1677 5854
rect 1681 5850 1682 5854
rect 1686 5850 1687 5854
rect 1672 5849 1691 5850
rect 1676 5845 1677 5849
rect 1681 5845 1682 5849
rect 1686 5845 1687 5849
rect 1672 5844 1691 5845
rect 1676 5840 1677 5844
rect 1681 5840 1682 5844
rect 1686 5840 1687 5844
rect 1672 5839 1691 5840
rect 1676 5835 1677 5839
rect 1681 5835 1682 5839
rect 1686 5835 1687 5839
rect 1672 5834 1691 5835
rect 1676 5830 1677 5834
rect 1681 5830 1682 5834
rect 1686 5830 1687 5834
rect 1672 5829 1691 5830
rect 1676 5825 1677 5829
rect 1681 5825 1682 5829
rect 1686 5825 1687 5829
rect 1672 5824 1691 5825
rect 1676 5820 1677 5824
rect 1681 5820 1682 5824
rect 1686 5820 1687 5824
rect 1985 5850 1986 5854
rect 1990 5850 1991 5854
rect 1995 5850 1996 5854
rect 1981 5849 2000 5850
rect 1985 5845 1986 5849
rect 1990 5845 1991 5849
rect 1995 5845 1996 5849
rect 1981 5844 2000 5845
rect 1985 5840 1986 5844
rect 1990 5840 1991 5844
rect 1995 5840 1996 5844
rect 1981 5839 2000 5840
rect 1985 5835 1986 5839
rect 1990 5835 1991 5839
rect 1995 5835 1996 5839
rect 1981 5834 2000 5835
rect 1985 5830 1986 5834
rect 1990 5830 1991 5834
rect 1995 5830 1996 5834
rect 1981 5829 2000 5830
rect 1985 5825 1986 5829
rect 1990 5825 1991 5829
rect 1995 5825 1996 5829
rect 1981 5824 2000 5825
rect 1985 5820 1986 5824
rect 1990 5820 1991 5824
rect 1995 5820 1996 5824
rect 2294 5850 2295 5854
rect 2299 5850 2300 5854
rect 2304 5850 2305 5854
rect 2290 5849 2309 5850
rect 2294 5845 2295 5849
rect 2299 5845 2300 5849
rect 2304 5845 2305 5849
rect 2290 5844 2309 5845
rect 2294 5840 2295 5844
rect 2299 5840 2300 5844
rect 2304 5840 2305 5844
rect 2290 5839 2309 5840
rect 2294 5835 2295 5839
rect 2299 5835 2300 5839
rect 2304 5835 2305 5839
rect 2290 5834 2309 5835
rect 2294 5830 2295 5834
rect 2299 5830 2300 5834
rect 2304 5830 2305 5834
rect 2290 5829 2309 5830
rect 2294 5825 2295 5829
rect 2299 5825 2300 5829
rect 2304 5825 2305 5829
rect 2290 5824 2309 5825
rect 2294 5820 2295 5824
rect 2299 5820 2300 5824
rect 2304 5820 2305 5824
rect 2603 5850 2604 5854
rect 2608 5850 2609 5854
rect 2613 5850 2614 5854
rect 2599 5849 2618 5850
rect 2603 5845 2604 5849
rect 2608 5845 2609 5849
rect 2613 5845 2614 5849
rect 2599 5844 2618 5845
rect 2603 5840 2604 5844
rect 2608 5840 2609 5844
rect 2613 5840 2614 5844
rect 2599 5839 2618 5840
rect 2603 5835 2604 5839
rect 2608 5835 2609 5839
rect 2613 5835 2614 5839
rect 2599 5834 2618 5835
rect 2603 5830 2604 5834
rect 2608 5830 2609 5834
rect 2613 5830 2614 5834
rect 2599 5829 2618 5830
rect 2603 5825 2604 5829
rect 2608 5825 2609 5829
rect 2613 5825 2614 5829
rect 2599 5824 2618 5825
rect 2603 5820 2604 5824
rect 2608 5820 2609 5824
rect 2613 5820 2614 5824
rect 2912 5850 2913 5854
rect 2917 5850 2918 5854
rect 2922 5850 2923 5854
rect 2908 5849 2927 5850
rect 2912 5845 2913 5849
rect 2917 5845 2918 5849
rect 2922 5845 2923 5849
rect 2908 5844 2927 5845
rect 2912 5840 2913 5844
rect 2917 5840 2918 5844
rect 2922 5840 2923 5844
rect 2908 5839 2927 5840
rect 2912 5835 2913 5839
rect 2917 5835 2918 5839
rect 2922 5835 2923 5839
rect 2908 5834 2927 5835
rect 2912 5830 2913 5834
rect 2917 5830 2918 5834
rect 2922 5830 2923 5834
rect 2908 5829 2927 5830
rect 2912 5825 2913 5829
rect 2917 5825 2918 5829
rect 2922 5825 2923 5829
rect 2908 5824 2927 5825
rect 2912 5820 2913 5824
rect 2917 5820 2918 5824
rect 2922 5820 2923 5824
rect 3221 5850 3222 5854
rect 3226 5850 3227 5854
rect 3231 5850 3232 5854
rect 3217 5849 3236 5850
rect 3221 5845 3222 5849
rect 3226 5845 3227 5849
rect 3231 5845 3232 5849
rect 3217 5844 3236 5845
rect 3221 5840 3222 5844
rect 3226 5840 3227 5844
rect 3231 5840 3232 5844
rect 3217 5839 3236 5840
rect 3221 5835 3222 5839
rect 3226 5835 3227 5839
rect 3231 5835 3232 5839
rect 3217 5834 3236 5835
rect 3221 5830 3222 5834
rect 3226 5830 3227 5834
rect 3231 5830 3232 5834
rect 3217 5829 3236 5830
rect 3221 5825 3222 5829
rect 3226 5825 3227 5829
rect 3231 5825 3232 5829
rect 3217 5824 3236 5825
rect 3221 5820 3222 5824
rect 3226 5820 3227 5824
rect 3231 5820 3232 5824
rect 3530 5850 3531 5854
rect 3535 5850 3536 5854
rect 3540 5850 3541 5854
rect 3526 5849 3545 5850
rect 3530 5845 3531 5849
rect 3535 5845 3536 5849
rect 3540 5845 3541 5849
rect 3526 5844 3545 5845
rect 3530 5840 3531 5844
rect 3535 5840 3536 5844
rect 3540 5840 3541 5844
rect 3526 5839 3545 5840
rect 3530 5835 3531 5839
rect 3535 5835 3536 5839
rect 3540 5835 3541 5839
rect 3526 5834 3545 5835
rect 3530 5830 3531 5834
rect 3535 5830 3536 5834
rect 3540 5830 3541 5834
rect 3526 5829 3545 5830
rect 3530 5825 3531 5829
rect 3535 5825 3536 5829
rect 3540 5825 3541 5829
rect 3526 5824 3545 5825
rect 3530 5820 3531 5824
rect 3535 5820 3536 5824
rect 3540 5820 3541 5824
rect 3839 5850 3840 5854
rect 3844 5850 3845 5854
rect 3849 5850 3850 5854
rect 3835 5849 3854 5850
rect 3839 5845 3840 5849
rect 3844 5845 3845 5849
rect 3849 5845 3850 5849
rect 3835 5844 3854 5845
rect 3839 5840 3840 5844
rect 3844 5840 3845 5844
rect 3849 5840 3850 5844
rect 3835 5839 3854 5840
rect 3839 5835 3840 5839
rect 3844 5835 3845 5839
rect 3849 5835 3850 5839
rect 3835 5834 3854 5835
rect 3839 5830 3840 5834
rect 3844 5830 3845 5834
rect 3849 5830 3850 5834
rect 3835 5829 3854 5830
rect 3839 5825 3840 5829
rect 3844 5825 3845 5829
rect 3849 5825 3850 5829
rect 3835 5824 3854 5825
rect 3839 5820 3840 5824
rect 3844 5820 3845 5824
rect 3849 5820 3850 5824
rect 4239 5850 4240 5854
rect 4244 5850 4245 5854
rect 4249 5850 4250 5854
rect 4235 5849 4254 5850
rect 4239 5845 4240 5849
rect 4244 5845 4245 5849
rect 4249 5845 4250 5849
rect 4235 5844 4254 5845
rect 4239 5840 4240 5844
rect 4244 5840 4245 5844
rect 4249 5840 4250 5844
rect 4235 5839 4254 5840
rect 4239 5835 4240 5839
rect 4244 5835 4245 5839
rect 4249 5835 4250 5839
rect 4235 5834 4254 5835
rect 4239 5830 4240 5834
rect 4244 5830 4245 5834
rect 4249 5830 4250 5834
rect 4235 5829 4254 5830
rect 4239 5825 4240 5829
rect 4244 5825 4245 5829
rect 4249 5825 4250 5829
rect 4235 5824 4254 5825
rect 4239 5820 4240 5824
rect 4244 5820 4245 5824
rect 4249 5820 4250 5824
rect 4268 5850 4269 5854
rect 4273 5850 4274 5854
rect 4278 5850 4279 5854
rect 4264 5849 4283 5850
rect 4268 5845 4269 5849
rect 4273 5845 4274 5849
rect 4278 5845 4279 5849
rect 4264 5844 4283 5845
rect 4268 5840 4269 5844
rect 4273 5840 4274 5844
rect 4278 5840 4279 5844
rect 4264 5839 4283 5840
rect 4268 5835 4269 5839
rect 4273 5835 4274 5839
rect 4278 5835 4279 5839
rect 4264 5834 4283 5835
rect 4268 5830 4269 5834
rect 4273 5830 4274 5834
rect 4278 5830 4279 5834
rect 4264 5829 4283 5830
rect 4268 5825 4269 5829
rect 4273 5825 4274 5829
rect 4278 5825 4279 5829
rect 4264 5824 4283 5825
rect 4268 5820 4269 5824
rect 4273 5820 4274 5824
rect 4278 5820 4279 5824
rect 4297 5850 4298 5854
rect 4302 5850 4303 5854
rect 4307 5850 4308 5854
rect 4293 5849 4312 5850
rect 4297 5845 4298 5849
rect 4302 5845 4303 5849
rect 4307 5845 4308 5849
rect 4293 5844 4312 5845
rect 4297 5840 4298 5844
rect 4302 5840 4303 5844
rect 4307 5840 4308 5844
rect 4293 5839 4312 5840
rect 4297 5835 4298 5839
rect 4302 5835 4303 5839
rect 4307 5835 4308 5839
rect 4293 5834 4312 5835
rect 4297 5830 4298 5834
rect 4302 5830 4303 5834
rect 4307 5830 4308 5834
rect 4293 5829 4312 5830
rect 4297 5825 4298 5829
rect 4302 5825 4303 5829
rect 4307 5825 4308 5829
rect 4293 5824 4312 5825
rect 4297 5820 4298 5824
rect 4302 5820 4303 5824
rect 4307 5820 4308 5824
rect 4326 5850 4327 5854
rect 4331 5850 4332 5854
rect 4336 5850 4337 5854
rect 4322 5849 4341 5850
rect 4326 5845 4327 5849
rect 4331 5845 4332 5849
rect 4336 5845 4337 5849
rect 4322 5844 4341 5845
rect 4326 5840 4327 5844
rect 4331 5840 4332 5844
rect 4336 5840 4337 5844
rect 4322 5839 4341 5840
rect 4326 5835 4327 5839
rect 4331 5835 4332 5839
rect 4336 5835 4337 5839
rect 4322 5834 4341 5835
rect 4326 5830 4327 5834
rect 4331 5830 4332 5834
rect 4336 5830 4337 5834
rect 4322 5829 4341 5830
rect 4326 5825 4327 5829
rect 4331 5825 4332 5829
rect 4336 5825 4337 5829
rect 4322 5824 4341 5825
rect 4326 5820 4327 5824
rect 4331 5820 4332 5824
rect 4336 5820 4337 5824
rect 4355 5850 4356 5854
rect 4360 5850 4361 5854
rect 4365 5850 4366 5854
rect 4351 5849 4370 5850
rect 4355 5845 4356 5849
rect 4360 5845 4361 5849
rect 4365 5845 4366 5849
rect 4351 5844 4370 5845
rect 4355 5840 4356 5844
rect 4360 5840 4361 5844
rect 4365 5840 4366 5844
rect 4351 5839 4370 5840
rect 4355 5835 4356 5839
rect 4360 5835 4361 5839
rect 4365 5835 4366 5839
rect 4351 5834 4370 5835
rect 4355 5830 4356 5834
rect 4360 5830 4361 5834
rect 4365 5830 4366 5834
rect 4351 5829 4370 5830
rect 4355 5825 4356 5829
rect 4360 5825 4361 5829
rect 4365 5825 4366 5829
rect 4351 5824 4370 5825
rect 4355 5820 4356 5824
rect 4360 5820 4361 5824
rect 4365 5820 4366 5824
rect 4579 5800 5054 6238
rect 99 5325 1031 5800
rect 1072 5550 1332 5553
rect 1072 5296 1075 5550
rect 1329 5296 1332 5550
rect 1072 5293 1332 5296
rect 1381 5550 1641 5553
rect 1381 5296 1384 5550
rect 1638 5296 1641 5550
rect 1381 5293 1641 5296
rect 1690 5550 1950 5553
rect 1690 5296 1693 5550
rect 1947 5296 1950 5550
rect 1690 5293 1950 5296
rect 1999 5550 2259 5553
rect 1999 5296 2002 5550
rect 2256 5296 2259 5550
rect 1999 5293 2259 5296
rect 2308 5550 2568 5553
rect 2308 5296 2311 5550
rect 2565 5296 2568 5550
rect 2308 5293 2568 5296
rect 2617 5550 2877 5553
rect 2617 5296 2620 5550
rect 2874 5296 2877 5550
rect 2617 5293 2877 5296
rect 2926 5550 3186 5553
rect 2926 5296 2929 5550
rect 3183 5296 3186 5550
rect 2926 5293 3186 5296
rect 3235 5550 3495 5553
rect 3235 5296 3238 5550
rect 3492 5296 3495 5550
rect 3235 5293 3495 5296
rect 3544 5550 3804 5553
rect 3544 5296 3547 5550
rect 3801 5296 3804 5550
rect 3544 5293 3804 5296
rect 3853 5550 4113 5553
rect 3853 5296 3856 5550
rect 4110 5296 4113 5550
rect 4148 5306 5054 5800
rect 3853 5293 4113 5296
<< m3contact >>
rect 1354 9796 1358 9800
rect 1359 9796 1363 9800
rect 1354 9791 1358 9795
rect 1359 9791 1363 9795
rect 1354 9786 1358 9790
rect 1359 9786 1363 9790
rect 1354 9781 1358 9785
rect 1359 9781 1363 9785
rect 1354 9776 1358 9780
rect 1359 9776 1363 9780
rect 1354 9771 1358 9775
rect 1359 9771 1363 9775
rect 1354 9766 1358 9770
rect 1359 9766 1363 9770
rect 802 9762 806 9766
rect 807 9762 811 9766
rect 812 9762 816 9766
rect 817 9762 821 9766
rect 802 9752 806 9756
rect 807 9752 811 9756
rect 812 9752 816 9756
rect 817 9752 821 9756
rect 802 9742 806 9746
rect 807 9742 811 9746
rect 812 9742 816 9746
rect 817 9742 821 9746
rect 802 9732 806 9736
rect 807 9732 811 9736
rect 812 9732 816 9736
rect 817 9732 821 9736
rect 831 9762 835 9766
rect 836 9762 840 9766
rect 841 9762 845 9766
rect 846 9762 850 9766
rect 831 9752 835 9756
rect 836 9752 840 9756
rect 841 9752 845 9756
rect 846 9752 850 9756
rect 831 9742 835 9746
rect 836 9742 840 9746
rect 841 9742 845 9746
rect 846 9742 850 9746
rect 831 9732 835 9736
rect 836 9732 840 9736
rect 841 9732 845 9736
rect 846 9732 850 9736
rect 860 9762 864 9766
rect 865 9762 869 9766
rect 870 9762 874 9766
rect 875 9762 879 9766
rect 860 9752 864 9756
rect 865 9752 869 9756
rect 870 9752 874 9756
rect 875 9752 879 9756
rect 860 9742 864 9746
rect 865 9742 869 9746
rect 870 9742 874 9746
rect 875 9742 879 9746
rect 860 9732 864 9736
rect 865 9732 869 9736
rect 870 9732 874 9736
rect 875 9732 879 9736
rect 889 9762 893 9766
rect 894 9762 898 9766
rect 899 9762 903 9766
rect 904 9762 908 9766
rect 889 9752 893 9756
rect 894 9752 898 9756
rect 899 9752 903 9756
rect 904 9752 908 9756
rect 889 9742 893 9746
rect 894 9742 898 9746
rect 899 9742 903 9746
rect 904 9742 908 9746
rect 889 9732 893 9736
rect 894 9732 898 9736
rect 899 9732 903 9736
rect 904 9732 908 9736
rect 918 9762 922 9766
rect 923 9762 927 9766
rect 928 9762 932 9766
rect 933 9762 937 9766
rect 918 9752 922 9756
rect 923 9752 927 9756
rect 928 9752 932 9756
rect 933 9752 937 9756
rect 918 9742 922 9746
rect 923 9742 927 9746
rect 928 9742 932 9746
rect 933 9742 937 9746
rect 918 9732 922 9736
rect 923 9732 927 9736
rect 928 9732 932 9736
rect 933 9732 937 9736
rect 1319 9762 1323 9766
rect 1324 9762 1328 9766
rect 1329 9762 1333 9766
rect 1334 9762 1338 9766
rect 1319 9752 1323 9756
rect 1324 9752 1328 9756
rect 1329 9752 1333 9756
rect 1334 9752 1338 9756
rect 1319 9742 1323 9746
rect 1324 9742 1328 9746
rect 1329 9742 1333 9746
rect 1334 9742 1338 9746
rect 1319 9732 1323 9736
rect 1324 9732 1328 9736
rect 1329 9732 1333 9736
rect 1334 9732 1338 9736
rect 1354 9761 1358 9765
rect 1359 9761 1363 9765
rect 1354 9756 1358 9760
rect 1359 9756 1363 9760
rect 1354 9751 1358 9755
rect 1359 9751 1363 9755
rect 1354 9746 1358 9750
rect 1359 9746 1363 9750
rect 1354 9741 1358 9745
rect 1359 9741 1363 9745
rect 1354 9736 1358 9740
rect 1359 9736 1363 9740
rect 802 9716 806 9720
rect 807 9716 811 9720
rect 812 9716 816 9720
rect 817 9716 821 9720
rect 802 9706 806 9710
rect 807 9706 811 9710
rect 812 9706 816 9710
rect 817 9706 821 9710
rect 802 9696 806 9700
rect 807 9696 811 9700
rect 812 9696 816 9700
rect 817 9696 821 9700
rect 802 9686 806 9690
rect 807 9686 811 9690
rect 812 9686 816 9690
rect 817 9686 821 9690
rect 831 9716 835 9720
rect 836 9716 840 9720
rect 841 9716 845 9720
rect 846 9716 850 9720
rect 831 9706 835 9710
rect 836 9706 840 9710
rect 841 9706 845 9710
rect 846 9706 850 9710
rect 831 9696 835 9700
rect 836 9696 840 9700
rect 841 9696 845 9700
rect 846 9696 850 9700
rect 831 9686 835 9690
rect 836 9686 840 9690
rect 841 9686 845 9690
rect 846 9686 850 9690
rect 860 9716 864 9720
rect 865 9716 869 9720
rect 870 9716 874 9720
rect 875 9716 879 9720
rect 860 9706 864 9710
rect 865 9706 869 9710
rect 870 9706 874 9710
rect 875 9706 879 9710
rect 860 9696 864 9700
rect 865 9696 869 9700
rect 870 9696 874 9700
rect 875 9696 879 9700
rect 860 9686 864 9690
rect 865 9686 869 9690
rect 870 9686 874 9690
rect 875 9686 879 9690
rect 889 9716 893 9720
rect 894 9716 898 9720
rect 899 9716 903 9720
rect 904 9716 908 9720
rect 889 9706 893 9710
rect 894 9706 898 9710
rect 899 9706 903 9710
rect 904 9706 908 9710
rect 889 9696 893 9700
rect 894 9696 898 9700
rect 899 9696 903 9700
rect 904 9696 908 9700
rect 889 9686 893 9690
rect 894 9686 898 9690
rect 899 9686 903 9690
rect 904 9686 908 9690
rect 918 9716 922 9720
rect 923 9716 927 9720
rect 928 9716 932 9720
rect 933 9716 937 9720
rect 918 9706 922 9710
rect 923 9706 927 9710
rect 928 9706 932 9710
rect 933 9706 937 9710
rect 918 9696 922 9700
rect 923 9696 927 9700
rect 928 9696 932 9700
rect 933 9696 937 9700
rect 918 9686 922 9690
rect 923 9686 927 9690
rect 928 9686 932 9690
rect 933 9686 937 9690
rect 1319 9716 1323 9720
rect 1324 9716 1328 9720
rect 1329 9716 1333 9720
rect 1334 9716 1338 9720
rect 1319 9706 1323 9710
rect 1324 9706 1328 9710
rect 1329 9706 1333 9710
rect 1334 9706 1338 9710
rect 1547 9765 1551 9769
rect 1552 9765 1556 9769
rect 1557 9765 1561 9769
rect 1562 9765 1566 9769
rect 1567 9765 1571 9769
rect 1572 9765 1576 9769
rect 1577 9765 1581 9769
rect 1582 9765 1586 9769
rect 1587 9765 1591 9769
rect 1592 9765 1596 9769
rect 1597 9765 1601 9769
rect 1602 9765 1606 9769
rect 1607 9765 1611 9769
rect 1663 9796 1667 9800
rect 1668 9796 1672 9800
rect 1663 9791 1667 9795
rect 1668 9791 1672 9795
rect 1663 9786 1667 9790
rect 1668 9786 1672 9790
rect 1663 9781 1667 9785
rect 1668 9781 1672 9785
rect 1663 9776 1667 9780
rect 1668 9776 1672 9780
rect 1663 9771 1667 9775
rect 1668 9771 1672 9775
rect 1663 9766 1667 9770
rect 1668 9766 1672 9770
rect 1547 9760 1551 9764
rect 1552 9760 1556 9764
rect 1557 9760 1561 9764
rect 1562 9760 1566 9764
rect 1567 9760 1571 9764
rect 1572 9760 1576 9764
rect 1577 9760 1581 9764
rect 1582 9760 1586 9764
rect 1587 9760 1591 9764
rect 1592 9760 1596 9764
rect 1597 9760 1601 9764
rect 1602 9760 1606 9764
rect 1607 9760 1611 9764
rect 1628 9762 1632 9766
rect 1633 9762 1637 9766
rect 1638 9762 1642 9766
rect 1643 9762 1647 9766
rect 1628 9752 1632 9756
rect 1633 9752 1637 9756
rect 1638 9752 1642 9756
rect 1643 9752 1647 9756
rect 1628 9742 1632 9746
rect 1633 9742 1637 9746
rect 1638 9742 1642 9746
rect 1643 9742 1647 9746
rect 1628 9732 1632 9736
rect 1633 9732 1637 9736
rect 1638 9732 1642 9736
rect 1643 9732 1647 9736
rect 1663 9761 1667 9765
rect 1668 9761 1672 9765
rect 1663 9756 1667 9760
rect 1668 9756 1672 9760
rect 1663 9751 1667 9755
rect 1668 9751 1672 9755
rect 1663 9746 1667 9750
rect 1668 9746 1672 9750
rect 1663 9741 1667 9745
rect 1668 9741 1672 9745
rect 1663 9736 1667 9740
rect 1668 9736 1672 9740
rect 1387 9708 1391 9712
rect 1392 9708 1396 9712
rect 1397 9708 1401 9712
rect 1402 9708 1406 9712
rect 1407 9708 1411 9712
rect 1412 9708 1416 9712
rect 1417 9708 1421 9712
rect 1422 9708 1426 9712
rect 1427 9708 1431 9712
rect 1432 9708 1436 9712
rect 1437 9708 1441 9712
rect 1442 9708 1446 9712
rect 1447 9708 1451 9712
rect 1387 9703 1391 9707
rect 1392 9703 1396 9707
rect 1397 9703 1401 9707
rect 1402 9703 1406 9707
rect 1407 9703 1411 9707
rect 1412 9703 1416 9707
rect 1417 9703 1421 9707
rect 1422 9703 1426 9707
rect 1427 9703 1431 9707
rect 1432 9703 1436 9707
rect 1437 9703 1441 9707
rect 1442 9703 1446 9707
rect 1447 9703 1451 9707
rect 1489 9711 1493 9715
rect 1494 9711 1498 9715
rect 1489 9706 1493 9710
rect 1494 9706 1498 9710
rect 1489 9701 1493 9705
rect 1494 9701 1498 9705
rect 1569 9708 1573 9712
rect 1574 9708 1578 9712
rect 1579 9708 1583 9712
rect 1584 9708 1588 9712
rect 1589 9708 1593 9712
rect 1594 9708 1598 9712
rect 1599 9708 1603 9712
rect 1604 9708 1608 9712
rect 1609 9708 1613 9712
rect 1614 9708 1618 9712
rect 1619 9708 1623 9712
rect 1569 9703 1573 9707
rect 1574 9703 1578 9707
rect 1579 9703 1583 9707
rect 1584 9703 1588 9707
rect 1589 9703 1593 9707
rect 1594 9703 1598 9707
rect 1599 9703 1603 9707
rect 1604 9703 1608 9707
rect 1609 9703 1613 9707
rect 1614 9703 1618 9707
rect 1619 9703 1623 9707
rect 1628 9716 1632 9720
rect 1633 9716 1637 9720
rect 1638 9716 1642 9720
rect 1643 9716 1647 9720
rect 1628 9706 1632 9710
rect 1633 9706 1637 9710
rect 1638 9706 1642 9710
rect 1643 9706 1647 9710
rect 1319 9696 1323 9700
rect 1324 9696 1328 9700
rect 1329 9696 1333 9700
rect 1334 9696 1338 9700
rect 1319 9686 1323 9690
rect 1324 9686 1328 9690
rect 1329 9686 1333 9690
rect 1334 9686 1338 9690
rect 1489 9696 1493 9700
rect 1494 9696 1498 9700
rect 1489 9691 1493 9695
rect 1494 9691 1498 9695
rect 1489 9686 1493 9690
rect 1494 9686 1498 9690
rect 1856 9765 1860 9769
rect 1861 9765 1865 9769
rect 1866 9765 1870 9769
rect 1871 9765 1875 9769
rect 1876 9765 1880 9769
rect 1881 9765 1885 9769
rect 1886 9765 1890 9769
rect 1891 9765 1895 9769
rect 1896 9765 1900 9769
rect 1901 9765 1905 9769
rect 1906 9765 1910 9769
rect 1911 9765 1915 9769
rect 1916 9765 1920 9769
rect 1972 9796 1976 9800
rect 1977 9796 1981 9800
rect 1972 9791 1976 9795
rect 1977 9791 1981 9795
rect 1972 9786 1976 9790
rect 1977 9786 1981 9790
rect 1972 9781 1976 9785
rect 1977 9781 1981 9785
rect 1972 9776 1976 9780
rect 1977 9776 1981 9780
rect 1972 9771 1976 9775
rect 1977 9771 1981 9775
rect 1972 9766 1976 9770
rect 1977 9766 1981 9770
rect 1856 9760 1860 9764
rect 1861 9760 1865 9764
rect 1866 9760 1870 9764
rect 1871 9760 1875 9764
rect 1876 9760 1880 9764
rect 1881 9760 1885 9764
rect 1886 9760 1890 9764
rect 1891 9760 1895 9764
rect 1896 9760 1900 9764
rect 1901 9760 1905 9764
rect 1906 9760 1910 9764
rect 1911 9760 1915 9764
rect 1916 9760 1920 9764
rect 1937 9762 1941 9766
rect 1942 9762 1946 9766
rect 1947 9762 1951 9766
rect 1952 9762 1956 9766
rect 1937 9752 1941 9756
rect 1942 9752 1946 9756
rect 1947 9752 1951 9756
rect 1952 9752 1956 9756
rect 1937 9742 1941 9746
rect 1942 9742 1946 9746
rect 1947 9742 1951 9746
rect 1952 9742 1956 9746
rect 1937 9732 1941 9736
rect 1942 9732 1946 9736
rect 1947 9732 1951 9736
rect 1952 9732 1956 9736
rect 1972 9761 1976 9765
rect 1977 9761 1981 9765
rect 1972 9756 1976 9760
rect 1977 9756 1981 9760
rect 1972 9751 1976 9755
rect 1977 9751 1981 9755
rect 1972 9746 1976 9750
rect 1977 9746 1981 9750
rect 1972 9741 1976 9745
rect 1977 9741 1981 9745
rect 1972 9736 1976 9740
rect 1977 9736 1981 9740
rect 1696 9708 1700 9712
rect 1701 9708 1705 9712
rect 1706 9708 1710 9712
rect 1711 9708 1715 9712
rect 1716 9708 1720 9712
rect 1721 9708 1725 9712
rect 1726 9708 1730 9712
rect 1731 9708 1735 9712
rect 1736 9708 1740 9712
rect 1741 9708 1745 9712
rect 1746 9708 1750 9712
rect 1751 9708 1755 9712
rect 1756 9708 1760 9712
rect 1696 9703 1700 9707
rect 1701 9703 1705 9707
rect 1706 9703 1710 9707
rect 1711 9703 1715 9707
rect 1716 9703 1720 9707
rect 1721 9703 1725 9707
rect 1726 9703 1730 9707
rect 1731 9703 1735 9707
rect 1736 9703 1740 9707
rect 1741 9703 1745 9707
rect 1746 9703 1750 9707
rect 1751 9703 1755 9707
rect 1756 9703 1760 9707
rect 1878 9708 1882 9712
rect 1883 9708 1887 9712
rect 1888 9708 1892 9712
rect 1893 9708 1897 9712
rect 1898 9708 1902 9712
rect 1903 9708 1907 9712
rect 1908 9708 1912 9712
rect 1913 9708 1917 9712
rect 1918 9708 1922 9712
rect 1923 9708 1927 9712
rect 1928 9708 1932 9712
rect 1878 9703 1882 9707
rect 1883 9703 1887 9707
rect 1888 9703 1892 9707
rect 1893 9703 1897 9707
rect 1898 9703 1902 9707
rect 1903 9703 1907 9707
rect 1908 9703 1912 9707
rect 1913 9703 1917 9707
rect 1918 9703 1922 9707
rect 1923 9703 1927 9707
rect 1928 9703 1932 9707
rect 1937 9716 1941 9720
rect 1942 9716 1946 9720
rect 1947 9716 1951 9720
rect 1952 9716 1956 9720
rect 1937 9706 1941 9710
rect 1942 9706 1946 9710
rect 1947 9706 1951 9710
rect 1952 9706 1956 9710
rect 2165 9765 2169 9769
rect 2170 9765 2174 9769
rect 2175 9765 2179 9769
rect 2180 9765 2184 9769
rect 2185 9765 2189 9769
rect 2190 9765 2194 9769
rect 2195 9765 2199 9769
rect 2200 9765 2204 9769
rect 2205 9765 2209 9769
rect 2210 9765 2214 9769
rect 2215 9765 2219 9769
rect 2220 9765 2224 9769
rect 2225 9765 2229 9769
rect 2281 9796 2285 9800
rect 2286 9796 2290 9800
rect 2281 9791 2285 9795
rect 2286 9791 2290 9795
rect 2281 9786 2285 9790
rect 2286 9786 2290 9790
rect 2281 9781 2285 9785
rect 2286 9781 2290 9785
rect 2281 9776 2285 9780
rect 2286 9776 2290 9780
rect 2281 9771 2285 9775
rect 2286 9771 2290 9775
rect 2281 9766 2285 9770
rect 2286 9766 2290 9770
rect 2165 9760 2169 9764
rect 2170 9760 2174 9764
rect 2175 9760 2179 9764
rect 2180 9760 2184 9764
rect 2185 9760 2189 9764
rect 2190 9760 2194 9764
rect 2195 9760 2199 9764
rect 2200 9760 2204 9764
rect 2205 9760 2209 9764
rect 2210 9760 2214 9764
rect 2215 9760 2219 9764
rect 2220 9760 2224 9764
rect 2225 9760 2229 9764
rect 2246 9762 2250 9766
rect 2251 9762 2255 9766
rect 2256 9762 2260 9766
rect 2261 9762 2265 9766
rect 2246 9752 2250 9756
rect 2251 9752 2255 9756
rect 2256 9752 2260 9756
rect 2261 9752 2265 9756
rect 2005 9708 2009 9712
rect 2010 9708 2014 9712
rect 2015 9708 2019 9712
rect 2020 9708 2024 9712
rect 2025 9708 2029 9712
rect 2030 9708 2034 9712
rect 2035 9708 2039 9712
rect 2040 9708 2044 9712
rect 2045 9708 2049 9712
rect 2050 9708 2054 9712
rect 2055 9708 2059 9712
rect 2060 9708 2064 9712
rect 2065 9708 2069 9712
rect 2005 9703 2009 9707
rect 2010 9703 2014 9707
rect 2015 9703 2019 9707
rect 2020 9703 2024 9707
rect 2025 9703 2029 9707
rect 2030 9703 2034 9707
rect 2035 9703 2039 9707
rect 2040 9703 2044 9707
rect 2045 9703 2049 9707
rect 2050 9703 2054 9707
rect 2055 9703 2059 9707
rect 2060 9703 2064 9707
rect 2065 9703 2069 9707
rect 2167 9736 2172 9741
rect 1628 9696 1632 9700
rect 1633 9696 1637 9700
rect 1638 9696 1642 9700
rect 1643 9696 1647 9700
rect 1628 9686 1632 9690
rect 1633 9686 1637 9690
rect 1638 9686 1642 9690
rect 1643 9686 1647 9690
rect 1937 9696 1941 9700
rect 1942 9696 1946 9700
rect 1947 9696 1951 9700
rect 1952 9696 1956 9700
rect 1937 9686 1941 9690
rect 1942 9686 1946 9690
rect 1947 9686 1951 9690
rect 1952 9686 1956 9690
rect 1489 9681 1493 9685
rect 1494 9681 1498 9685
rect 1489 9676 1493 9680
rect 1494 9676 1498 9680
rect 1489 9671 1493 9675
rect 1494 9671 1498 9675
rect 1489 9666 1493 9670
rect 1494 9666 1498 9670
rect 1489 9661 1493 9665
rect 1494 9661 1498 9665
rect 2246 9742 2250 9746
rect 2251 9742 2255 9746
rect 2256 9742 2260 9746
rect 2261 9742 2265 9746
rect 2246 9732 2250 9736
rect 2251 9732 2255 9736
rect 2256 9732 2260 9736
rect 2261 9732 2265 9736
rect 2281 9761 2285 9765
rect 2286 9761 2290 9765
rect 2281 9756 2285 9760
rect 2286 9756 2290 9760
rect 2281 9751 2285 9755
rect 2286 9751 2290 9755
rect 2281 9746 2285 9750
rect 2286 9746 2290 9750
rect 2281 9741 2285 9745
rect 2286 9741 2290 9745
rect 2281 9736 2285 9740
rect 2286 9736 2290 9740
rect 2187 9708 2191 9712
rect 2192 9708 2196 9712
rect 2197 9708 2201 9712
rect 2202 9708 2206 9712
rect 2207 9708 2211 9712
rect 2212 9708 2216 9712
rect 2217 9708 2221 9712
rect 2222 9708 2226 9712
rect 2227 9708 2231 9712
rect 2232 9708 2236 9712
rect 2237 9708 2241 9712
rect 2187 9703 2191 9707
rect 2192 9703 2196 9707
rect 2197 9703 2201 9707
rect 2202 9703 2206 9707
rect 2207 9703 2211 9707
rect 2212 9703 2216 9707
rect 2217 9703 2221 9707
rect 2222 9703 2226 9707
rect 2227 9703 2231 9707
rect 2232 9703 2236 9707
rect 2237 9703 2241 9707
rect 2246 9716 2250 9720
rect 2251 9716 2255 9720
rect 2256 9716 2260 9720
rect 2261 9716 2265 9720
rect 2246 9706 2250 9710
rect 2251 9706 2255 9710
rect 2256 9706 2260 9710
rect 2261 9706 2265 9710
rect 2474 9765 2478 9769
rect 2479 9765 2483 9769
rect 2484 9765 2488 9769
rect 2489 9765 2493 9769
rect 2494 9765 2498 9769
rect 2499 9765 2503 9769
rect 2504 9765 2508 9769
rect 2509 9765 2513 9769
rect 2514 9765 2518 9769
rect 2519 9765 2523 9769
rect 2524 9765 2528 9769
rect 2529 9765 2533 9769
rect 2534 9765 2538 9769
rect 2590 9796 2594 9800
rect 2595 9796 2599 9800
rect 2590 9791 2594 9795
rect 2595 9791 2599 9795
rect 2590 9786 2594 9790
rect 2595 9786 2599 9790
rect 2590 9781 2594 9785
rect 2595 9781 2599 9785
rect 2590 9776 2594 9780
rect 2595 9776 2599 9780
rect 2590 9771 2594 9775
rect 2595 9771 2599 9775
rect 2590 9766 2594 9770
rect 2595 9766 2599 9770
rect 2474 9760 2478 9764
rect 2479 9760 2483 9764
rect 2484 9760 2488 9764
rect 2489 9760 2493 9764
rect 2494 9760 2498 9764
rect 2499 9760 2503 9764
rect 2504 9760 2508 9764
rect 2509 9760 2513 9764
rect 2514 9760 2518 9764
rect 2519 9760 2523 9764
rect 2524 9760 2528 9764
rect 2529 9760 2533 9764
rect 2534 9760 2538 9764
rect 2555 9762 2559 9766
rect 2560 9762 2564 9766
rect 2565 9762 2569 9766
rect 2570 9762 2574 9766
rect 2555 9752 2559 9756
rect 2560 9752 2564 9756
rect 2565 9752 2569 9756
rect 2570 9752 2574 9756
rect 2555 9742 2559 9746
rect 2560 9742 2564 9746
rect 2565 9742 2569 9746
rect 2570 9742 2574 9746
rect 2555 9732 2559 9736
rect 2560 9732 2564 9736
rect 2565 9732 2569 9736
rect 2570 9732 2574 9736
rect 2590 9761 2594 9765
rect 2595 9761 2599 9765
rect 2590 9756 2594 9760
rect 2595 9756 2599 9760
rect 2590 9751 2594 9755
rect 2595 9751 2599 9755
rect 2590 9746 2594 9750
rect 2595 9746 2599 9750
rect 2590 9741 2594 9745
rect 2595 9741 2599 9745
rect 2590 9736 2594 9740
rect 2595 9736 2599 9740
rect 2314 9708 2318 9712
rect 2319 9708 2323 9712
rect 2324 9708 2328 9712
rect 2329 9708 2333 9712
rect 2334 9708 2338 9712
rect 2339 9708 2343 9712
rect 2344 9708 2348 9712
rect 2349 9708 2353 9712
rect 2354 9708 2358 9712
rect 2359 9708 2363 9712
rect 2364 9708 2368 9712
rect 2369 9708 2373 9712
rect 2374 9708 2378 9712
rect 2314 9703 2318 9707
rect 2319 9703 2323 9707
rect 2324 9703 2328 9707
rect 2329 9703 2333 9707
rect 2334 9703 2338 9707
rect 2339 9703 2343 9707
rect 2344 9703 2348 9707
rect 2349 9703 2353 9707
rect 2354 9703 2358 9707
rect 2359 9703 2363 9707
rect 2364 9703 2368 9707
rect 2369 9703 2373 9707
rect 2374 9703 2378 9707
rect 2496 9708 2500 9712
rect 2501 9708 2505 9712
rect 2506 9708 2510 9712
rect 2511 9708 2515 9712
rect 2516 9708 2520 9712
rect 2521 9708 2525 9712
rect 2526 9708 2530 9712
rect 2531 9708 2535 9712
rect 2536 9708 2540 9712
rect 2541 9708 2545 9712
rect 2546 9708 2550 9712
rect 2496 9703 2500 9707
rect 2501 9703 2505 9707
rect 2506 9703 2510 9707
rect 2511 9703 2515 9707
rect 2516 9703 2520 9707
rect 2521 9703 2525 9707
rect 2526 9703 2530 9707
rect 2531 9703 2535 9707
rect 2536 9703 2540 9707
rect 2541 9703 2545 9707
rect 2546 9703 2550 9707
rect 2555 9716 2559 9720
rect 2560 9716 2564 9720
rect 2565 9716 2569 9720
rect 2570 9716 2574 9720
rect 2555 9706 2559 9710
rect 2560 9706 2564 9710
rect 2565 9706 2569 9710
rect 2570 9706 2574 9710
rect 2783 9765 2787 9769
rect 2788 9765 2792 9769
rect 2793 9765 2797 9769
rect 2798 9765 2802 9769
rect 2803 9765 2807 9769
rect 2808 9765 2812 9769
rect 2813 9765 2817 9769
rect 2818 9765 2822 9769
rect 2823 9765 2827 9769
rect 2828 9765 2832 9769
rect 2833 9765 2837 9769
rect 2838 9765 2842 9769
rect 2843 9765 2847 9769
rect 2899 9796 2903 9800
rect 2904 9796 2908 9800
rect 2899 9791 2903 9795
rect 2904 9791 2908 9795
rect 2899 9786 2903 9790
rect 2904 9786 2908 9790
rect 2899 9781 2903 9785
rect 2904 9781 2908 9785
rect 2899 9776 2903 9780
rect 2904 9776 2908 9780
rect 2899 9771 2903 9775
rect 2904 9771 2908 9775
rect 2899 9766 2903 9770
rect 2904 9766 2908 9770
rect 2783 9760 2787 9764
rect 2788 9760 2792 9764
rect 2793 9760 2797 9764
rect 2798 9760 2802 9764
rect 2803 9760 2807 9764
rect 2808 9760 2812 9764
rect 2813 9760 2817 9764
rect 2818 9760 2822 9764
rect 2823 9760 2827 9764
rect 2828 9760 2832 9764
rect 2833 9760 2837 9764
rect 2838 9760 2842 9764
rect 2843 9760 2847 9764
rect 2864 9762 2868 9766
rect 2869 9762 2873 9766
rect 2874 9762 2878 9766
rect 2879 9762 2883 9766
rect 2864 9752 2868 9756
rect 2869 9752 2873 9756
rect 2874 9752 2878 9756
rect 2879 9752 2883 9756
rect 2864 9742 2868 9746
rect 2869 9742 2873 9746
rect 2874 9742 2878 9746
rect 2879 9742 2883 9746
rect 2864 9732 2868 9736
rect 2869 9732 2873 9736
rect 2874 9732 2878 9736
rect 2879 9732 2883 9736
rect 2899 9761 2903 9765
rect 2904 9761 2908 9765
rect 2899 9756 2903 9760
rect 2904 9756 2908 9760
rect 2899 9751 2903 9755
rect 2904 9751 2908 9755
rect 2899 9746 2903 9750
rect 2904 9746 2908 9750
rect 2899 9741 2903 9745
rect 2904 9741 2908 9745
rect 2899 9736 2903 9740
rect 2904 9736 2908 9740
rect 2623 9708 2627 9712
rect 2628 9708 2632 9712
rect 2633 9708 2637 9712
rect 2638 9708 2642 9712
rect 2643 9708 2647 9712
rect 2648 9708 2652 9712
rect 2653 9708 2657 9712
rect 2658 9708 2662 9712
rect 2663 9708 2667 9712
rect 2668 9708 2672 9712
rect 2673 9708 2677 9712
rect 2678 9708 2682 9712
rect 2683 9708 2687 9712
rect 2623 9703 2627 9707
rect 2628 9703 2632 9707
rect 2633 9703 2637 9707
rect 2638 9703 2642 9707
rect 2643 9703 2647 9707
rect 2648 9703 2652 9707
rect 2653 9703 2657 9707
rect 2658 9703 2662 9707
rect 2663 9703 2667 9707
rect 2668 9703 2672 9707
rect 2673 9703 2677 9707
rect 2678 9703 2682 9707
rect 2683 9703 2687 9707
rect 2805 9708 2809 9712
rect 2810 9708 2814 9712
rect 2815 9708 2819 9712
rect 2820 9708 2824 9712
rect 2825 9708 2829 9712
rect 2830 9708 2834 9712
rect 2835 9708 2839 9712
rect 2840 9708 2844 9712
rect 2845 9708 2849 9712
rect 2850 9708 2854 9712
rect 2855 9708 2859 9712
rect 2805 9703 2809 9707
rect 2810 9703 2814 9707
rect 2815 9703 2819 9707
rect 2820 9703 2824 9707
rect 2825 9703 2829 9707
rect 2830 9703 2834 9707
rect 2835 9703 2839 9707
rect 2840 9703 2844 9707
rect 2845 9703 2849 9707
rect 2850 9703 2854 9707
rect 2855 9703 2859 9707
rect 2864 9716 2868 9720
rect 2869 9716 2873 9720
rect 2874 9716 2878 9720
rect 2879 9716 2883 9720
rect 2864 9706 2868 9710
rect 2869 9706 2873 9710
rect 2874 9706 2878 9710
rect 2879 9706 2883 9710
rect 3092 9765 3096 9769
rect 3097 9765 3101 9769
rect 3102 9765 3106 9769
rect 3107 9765 3111 9769
rect 3112 9765 3116 9769
rect 3117 9765 3121 9769
rect 3122 9765 3126 9769
rect 3127 9765 3131 9769
rect 3132 9765 3136 9769
rect 3137 9765 3141 9769
rect 3142 9765 3146 9769
rect 3147 9765 3151 9769
rect 3152 9765 3156 9769
rect 3208 9796 3212 9800
rect 3213 9796 3217 9800
rect 3208 9791 3212 9795
rect 3213 9791 3217 9795
rect 3208 9786 3212 9790
rect 3213 9786 3217 9790
rect 3208 9781 3212 9785
rect 3213 9781 3217 9785
rect 3208 9776 3212 9780
rect 3213 9776 3217 9780
rect 3208 9771 3212 9775
rect 3213 9771 3217 9775
rect 3208 9766 3212 9770
rect 3213 9766 3217 9770
rect 3092 9760 3096 9764
rect 3097 9760 3101 9764
rect 3102 9760 3106 9764
rect 3107 9760 3111 9764
rect 3112 9760 3116 9764
rect 3117 9760 3121 9764
rect 3122 9760 3126 9764
rect 3127 9760 3131 9764
rect 3132 9760 3136 9764
rect 3137 9760 3141 9764
rect 3142 9760 3146 9764
rect 3147 9760 3151 9764
rect 3152 9760 3156 9764
rect 3173 9762 3177 9766
rect 3178 9762 3182 9766
rect 3183 9762 3187 9766
rect 3188 9762 3192 9766
rect 3173 9752 3177 9756
rect 3178 9752 3182 9756
rect 3183 9752 3187 9756
rect 3188 9752 3192 9756
rect 3173 9742 3177 9746
rect 3178 9742 3182 9746
rect 3183 9742 3187 9746
rect 3188 9742 3192 9746
rect 3173 9732 3177 9736
rect 3178 9732 3182 9736
rect 3183 9732 3187 9736
rect 3188 9732 3192 9736
rect 3208 9761 3212 9765
rect 3213 9761 3217 9765
rect 3208 9756 3212 9760
rect 3213 9756 3217 9760
rect 3208 9751 3212 9755
rect 3213 9751 3217 9755
rect 3208 9746 3212 9750
rect 3213 9746 3217 9750
rect 3208 9741 3212 9745
rect 3213 9741 3217 9745
rect 3208 9736 3212 9740
rect 3213 9736 3217 9740
rect 2932 9708 2936 9712
rect 2937 9708 2941 9712
rect 2942 9708 2946 9712
rect 2947 9708 2951 9712
rect 2952 9708 2956 9712
rect 2957 9708 2961 9712
rect 2962 9708 2966 9712
rect 2967 9708 2971 9712
rect 2972 9708 2976 9712
rect 2977 9708 2981 9712
rect 2982 9708 2986 9712
rect 2987 9708 2991 9712
rect 2992 9708 2996 9712
rect 2932 9703 2936 9707
rect 2937 9703 2941 9707
rect 2942 9703 2946 9707
rect 2947 9703 2951 9707
rect 2952 9703 2956 9707
rect 2957 9703 2961 9707
rect 2962 9703 2966 9707
rect 2967 9703 2971 9707
rect 2972 9703 2976 9707
rect 2977 9703 2981 9707
rect 2982 9703 2986 9707
rect 2987 9703 2991 9707
rect 2992 9703 2996 9707
rect 3114 9708 3118 9712
rect 3119 9708 3123 9712
rect 3124 9708 3128 9712
rect 3129 9708 3133 9712
rect 3134 9708 3138 9712
rect 3139 9708 3143 9712
rect 3144 9708 3148 9712
rect 3149 9708 3153 9712
rect 3154 9708 3158 9712
rect 3159 9708 3163 9712
rect 3164 9708 3168 9712
rect 3114 9703 3118 9707
rect 3119 9703 3123 9707
rect 3124 9703 3128 9707
rect 3129 9703 3133 9707
rect 3134 9703 3138 9707
rect 3139 9703 3143 9707
rect 3144 9703 3148 9707
rect 3149 9703 3153 9707
rect 3154 9703 3158 9707
rect 3159 9703 3163 9707
rect 3164 9703 3168 9707
rect 3173 9716 3177 9720
rect 3178 9716 3182 9720
rect 3183 9716 3187 9720
rect 3188 9716 3192 9720
rect 3173 9706 3177 9710
rect 3178 9706 3182 9710
rect 3183 9706 3187 9710
rect 3188 9706 3192 9710
rect 3401 9765 3405 9769
rect 3406 9765 3410 9769
rect 3411 9765 3415 9769
rect 3416 9765 3420 9769
rect 3421 9765 3425 9769
rect 3426 9765 3430 9769
rect 3431 9765 3435 9769
rect 3436 9765 3440 9769
rect 3441 9765 3445 9769
rect 3446 9765 3450 9769
rect 3451 9765 3455 9769
rect 3456 9765 3460 9769
rect 3461 9765 3465 9769
rect 3517 9796 3521 9800
rect 3522 9796 3526 9800
rect 3517 9791 3521 9795
rect 3522 9791 3526 9795
rect 3517 9786 3521 9790
rect 3522 9786 3526 9790
rect 3517 9781 3521 9785
rect 3522 9781 3526 9785
rect 3517 9776 3521 9780
rect 3522 9776 3526 9780
rect 3517 9771 3521 9775
rect 3522 9771 3526 9775
rect 3517 9766 3521 9770
rect 3522 9766 3526 9770
rect 3401 9760 3405 9764
rect 3406 9760 3410 9764
rect 3411 9760 3415 9764
rect 3416 9760 3420 9764
rect 3421 9760 3425 9764
rect 3426 9760 3430 9764
rect 3431 9760 3435 9764
rect 3436 9760 3440 9764
rect 3441 9760 3445 9764
rect 3446 9760 3450 9764
rect 3451 9760 3455 9764
rect 3456 9760 3460 9764
rect 3461 9760 3465 9764
rect 3482 9762 3486 9766
rect 3487 9762 3491 9766
rect 3492 9762 3496 9766
rect 3497 9762 3501 9766
rect 3482 9752 3486 9756
rect 3487 9752 3491 9756
rect 3492 9752 3496 9756
rect 3497 9752 3501 9756
rect 3482 9742 3486 9746
rect 3487 9742 3491 9746
rect 3492 9742 3496 9746
rect 3497 9742 3501 9746
rect 3482 9732 3486 9736
rect 3487 9732 3491 9736
rect 3492 9732 3496 9736
rect 3497 9732 3501 9736
rect 3517 9761 3521 9765
rect 3522 9761 3526 9765
rect 3517 9756 3521 9760
rect 3522 9756 3526 9760
rect 3517 9751 3521 9755
rect 3522 9751 3526 9755
rect 3517 9746 3521 9750
rect 3522 9746 3526 9750
rect 3517 9741 3521 9745
rect 3522 9741 3526 9745
rect 3517 9736 3521 9740
rect 3522 9736 3526 9740
rect 3241 9708 3245 9712
rect 3246 9708 3250 9712
rect 3251 9708 3255 9712
rect 3256 9708 3260 9712
rect 3261 9708 3265 9712
rect 3266 9708 3270 9712
rect 3271 9708 3275 9712
rect 3276 9708 3280 9712
rect 3281 9708 3285 9712
rect 3286 9708 3290 9712
rect 3291 9708 3295 9712
rect 3296 9708 3300 9712
rect 3301 9708 3305 9712
rect 3241 9703 3245 9707
rect 3246 9703 3250 9707
rect 3251 9703 3255 9707
rect 3256 9703 3260 9707
rect 3261 9703 3265 9707
rect 3266 9703 3270 9707
rect 3271 9703 3275 9707
rect 3276 9703 3280 9707
rect 3281 9703 3285 9707
rect 3286 9703 3290 9707
rect 3291 9703 3295 9707
rect 3296 9703 3300 9707
rect 3301 9703 3305 9707
rect 3343 9711 3347 9715
rect 3348 9711 3352 9715
rect 3343 9706 3347 9710
rect 3348 9706 3352 9710
rect 3343 9701 3347 9705
rect 3348 9701 3352 9705
rect 3423 9708 3427 9712
rect 3428 9708 3432 9712
rect 3433 9708 3437 9712
rect 3438 9708 3442 9712
rect 3443 9708 3447 9712
rect 3448 9708 3452 9712
rect 3453 9708 3457 9712
rect 3458 9708 3462 9712
rect 3463 9708 3467 9712
rect 3468 9708 3472 9712
rect 3473 9708 3477 9712
rect 3423 9703 3427 9707
rect 3428 9703 3432 9707
rect 3433 9703 3437 9707
rect 3438 9703 3442 9707
rect 3443 9703 3447 9707
rect 3448 9703 3452 9707
rect 3453 9703 3457 9707
rect 3458 9703 3462 9707
rect 3463 9703 3467 9707
rect 3468 9703 3472 9707
rect 3473 9703 3477 9707
rect 3482 9716 3486 9720
rect 3487 9716 3491 9720
rect 3492 9716 3496 9720
rect 3497 9716 3501 9720
rect 3482 9706 3486 9710
rect 3487 9706 3491 9710
rect 3492 9706 3496 9710
rect 3497 9706 3501 9710
rect 2246 9696 2250 9700
rect 2251 9696 2255 9700
rect 2256 9696 2260 9700
rect 2261 9696 2265 9700
rect 2246 9686 2250 9690
rect 2251 9686 2255 9690
rect 2256 9686 2260 9690
rect 2261 9686 2265 9690
rect 2555 9696 2559 9700
rect 2560 9696 2564 9700
rect 2565 9696 2569 9700
rect 2570 9696 2574 9700
rect 2555 9686 2559 9690
rect 2560 9686 2564 9690
rect 2565 9686 2569 9690
rect 2570 9686 2574 9690
rect 2864 9696 2868 9700
rect 2869 9696 2873 9700
rect 2874 9696 2878 9700
rect 2879 9696 2883 9700
rect 2864 9686 2868 9690
rect 2869 9686 2873 9690
rect 2874 9686 2878 9690
rect 2879 9686 2883 9690
rect 3173 9696 3177 9700
rect 3178 9696 3182 9700
rect 3183 9696 3187 9700
rect 3188 9696 3192 9700
rect 3173 9686 3177 9690
rect 3178 9686 3182 9690
rect 3183 9686 3187 9690
rect 3188 9686 3192 9690
rect 3343 9696 3347 9700
rect 3348 9696 3352 9700
rect 3343 9691 3347 9695
rect 3348 9691 3352 9695
rect 3343 9686 3347 9690
rect 3348 9686 3352 9690
rect 3652 9791 3656 9795
rect 3657 9791 3661 9795
rect 3652 9786 3656 9790
rect 3657 9786 3661 9790
rect 3652 9781 3656 9785
rect 3657 9781 3661 9785
rect 3652 9776 3656 9780
rect 3657 9776 3661 9780
rect 3652 9771 3656 9775
rect 3657 9771 3661 9775
rect 3652 9766 3656 9770
rect 3657 9766 3661 9770
rect 3652 9761 3656 9765
rect 3657 9761 3661 9765
rect 3652 9756 3656 9760
rect 3657 9756 3661 9760
rect 3710 9765 3714 9769
rect 3715 9765 3719 9769
rect 3720 9765 3724 9769
rect 3725 9765 3729 9769
rect 3730 9765 3734 9769
rect 3735 9765 3739 9769
rect 3740 9765 3744 9769
rect 3745 9765 3749 9769
rect 3750 9765 3754 9769
rect 3755 9765 3759 9769
rect 3760 9765 3764 9769
rect 3765 9765 3769 9769
rect 3770 9765 3774 9769
rect 3826 9796 3830 9800
rect 3831 9796 3835 9800
rect 3826 9791 3830 9795
rect 3831 9791 3835 9795
rect 3826 9786 3830 9790
rect 3831 9786 3835 9790
rect 3826 9781 3830 9785
rect 3831 9781 3835 9785
rect 3826 9776 3830 9780
rect 3831 9776 3835 9780
rect 3826 9771 3830 9775
rect 3831 9771 3835 9775
rect 3826 9766 3830 9770
rect 3831 9766 3835 9770
rect 3710 9760 3714 9764
rect 3715 9760 3719 9764
rect 3720 9760 3724 9764
rect 3725 9760 3729 9764
rect 3730 9760 3734 9764
rect 3735 9760 3739 9764
rect 3740 9760 3744 9764
rect 3745 9760 3749 9764
rect 3750 9760 3754 9764
rect 3755 9760 3759 9764
rect 3760 9760 3764 9764
rect 3765 9760 3769 9764
rect 3770 9760 3774 9764
rect 3791 9762 3795 9766
rect 3796 9762 3800 9766
rect 3801 9762 3805 9766
rect 3806 9762 3810 9766
rect 3652 9751 3656 9755
rect 3657 9751 3661 9755
rect 3652 9746 3656 9750
rect 3657 9746 3661 9750
rect 3652 9741 3656 9745
rect 3657 9741 3661 9745
rect 3791 9752 3795 9756
rect 3796 9752 3800 9756
rect 3801 9752 3805 9756
rect 3806 9752 3810 9756
rect 3791 9742 3795 9746
rect 3796 9742 3800 9746
rect 3801 9742 3805 9746
rect 3806 9742 3810 9746
rect 3791 9732 3795 9736
rect 3796 9732 3800 9736
rect 3801 9732 3805 9736
rect 3806 9732 3810 9736
rect 3826 9761 3830 9765
rect 3831 9761 3835 9765
rect 3826 9756 3830 9760
rect 3831 9756 3835 9760
rect 3826 9751 3830 9755
rect 3831 9751 3835 9755
rect 3826 9746 3830 9750
rect 3831 9746 3835 9750
rect 3826 9741 3830 9745
rect 3831 9741 3835 9745
rect 3826 9736 3830 9740
rect 3831 9736 3835 9740
rect 3550 9708 3554 9712
rect 3555 9708 3559 9712
rect 3560 9708 3564 9712
rect 3565 9708 3569 9712
rect 3570 9708 3574 9712
rect 3575 9708 3579 9712
rect 3580 9708 3584 9712
rect 3585 9708 3589 9712
rect 3590 9708 3594 9712
rect 3595 9708 3599 9712
rect 3600 9708 3604 9712
rect 3605 9708 3609 9712
rect 3610 9708 3614 9712
rect 3550 9703 3554 9707
rect 3555 9703 3559 9707
rect 3560 9703 3564 9707
rect 3565 9703 3569 9707
rect 3570 9703 3574 9707
rect 3575 9703 3579 9707
rect 3580 9703 3584 9707
rect 3585 9703 3589 9707
rect 3590 9703 3594 9707
rect 3595 9703 3599 9707
rect 3600 9703 3604 9707
rect 3605 9703 3609 9707
rect 3610 9703 3614 9707
rect 3732 9708 3736 9712
rect 3737 9708 3741 9712
rect 3742 9708 3746 9712
rect 3747 9708 3751 9712
rect 3752 9708 3756 9712
rect 3757 9708 3761 9712
rect 3762 9708 3766 9712
rect 3767 9708 3771 9712
rect 3772 9708 3776 9712
rect 3777 9708 3781 9712
rect 3782 9708 3786 9712
rect 3732 9703 3736 9707
rect 3737 9703 3741 9707
rect 3742 9703 3746 9707
rect 3747 9703 3751 9707
rect 3752 9703 3756 9707
rect 3757 9703 3761 9707
rect 3762 9703 3766 9707
rect 3767 9703 3771 9707
rect 3772 9703 3776 9707
rect 3777 9703 3781 9707
rect 3782 9703 3786 9707
rect 3791 9716 3795 9720
rect 3796 9716 3800 9720
rect 3801 9716 3805 9720
rect 3806 9716 3810 9720
rect 3791 9706 3795 9710
rect 3796 9706 3800 9710
rect 3801 9706 3805 9710
rect 3806 9706 3810 9710
rect 4019 9765 4023 9769
rect 4024 9765 4028 9769
rect 4029 9765 4033 9769
rect 4034 9765 4038 9769
rect 4039 9765 4043 9769
rect 4044 9765 4048 9769
rect 4049 9765 4053 9769
rect 4054 9765 4058 9769
rect 4059 9765 4063 9769
rect 4064 9765 4068 9769
rect 4069 9765 4073 9769
rect 4074 9765 4078 9769
rect 4079 9765 4083 9769
rect 4019 9760 4023 9764
rect 4024 9760 4028 9764
rect 4029 9760 4033 9764
rect 4034 9760 4038 9764
rect 4039 9760 4043 9764
rect 4044 9760 4048 9764
rect 4049 9760 4053 9764
rect 4054 9760 4058 9764
rect 4059 9760 4063 9764
rect 4064 9760 4068 9764
rect 4069 9760 4073 9764
rect 4074 9760 4078 9764
rect 4079 9760 4083 9764
rect 4100 9762 4104 9766
rect 4105 9762 4109 9766
rect 4110 9762 4114 9766
rect 4115 9762 4119 9766
rect 4100 9752 4104 9756
rect 4105 9752 4109 9756
rect 4110 9752 4114 9756
rect 4115 9752 4119 9756
rect 4100 9742 4104 9746
rect 4105 9742 4109 9746
rect 4110 9742 4114 9746
rect 4115 9742 4119 9746
rect 4100 9732 4104 9736
rect 4105 9732 4109 9736
rect 4110 9732 4114 9736
rect 4115 9732 4119 9736
rect 4292 9762 4296 9766
rect 4297 9762 4301 9766
rect 4302 9762 4306 9766
rect 4307 9762 4311 9766
rect 4292 9752 4296 9756
rect 4297 9752 4301 9756
rect 4302 9752 4306 9756
rect 4307 9752 4311 9756
rect 4292 9742 4296 9746
rect 4297 9742 4301 9746
rect 4302 9742 4306 9746
rect 4307 9742 4311 9746
rect 4292 9732 4296 9736
rect 4297 9732 4301 9736
rect 4302 9732 4306 9736
rect 4307 9732 4311 9736
rect 4318 9762 4322 9766
rect 4323 9762 4327 9766
rect 4328 9762 4332 9766
rect 4333 9762 4337 9766
rect 4318 9752 4322 9756
rect 4323 9752 4327 9756
rect 4328 9752 4332 9756
rect 4333 9752 4337 9756
rect 4318 9742 4322 9746
rect 4323 9742 4327 9746
rect 4328 9742 4332 9746
rect 4333 9742 4337 9746
rect 4318 9732 4322 9736
rect 4323 9732 4327 9736
rect 4328 9732 4332 9736
rect 4333 9732 4337 9736
rect 4344 9762 4348 9766
rect 4349 9762 4353 9766
rect 4354 9762 4358 9766
rect 4359 9762 4363 9766
rect 4344 9752 4348 9756
rect 4349 9752 4353 9756
rect 4354 9752 4358 9756
rect 4359 9752 4363 9756
rect 4344 9742 4348 9746
rect 4349 9742 4353 9746
rect 4354 9742 4358 9746
rect 4359 9742 4363 9746
rect 4344 9732 4348 9736
rect 4349 9732 4353 9736
rect 4354 9732 4358 9736
rect 4359 9732 4363 9736
rect 4370 9762 4374 9766
rect 4375 9762 4379 9766
rect 4380 9762 4384 9766
rect 4385 9762 4389 9766
rect 4370 9752 4374 9756
rect 4375 9752 4379 9756
rect 4380 9752 4384 9756
rect 4385 9752 4389 9756
rect 4370 9742 4374 9746
rect 4375 9742 4379 9746
rect 4380 9742 4384 9746
rect 4385 9742 4389 9746
rect 4370 9732 4374 9736
rect 4375 9732 4379 9736
rect 4380 9732 4384 9736
rect 4385 9732 4389 9736
rect 4396 9762 4400 9766
rect 4401 9762 4405 9766
rect 4406 9762 4410 9766
rect 4411 9762 4415 9766
rect 4396 9752 4400 9756
rect 4401 9752 4405 9756
rect 4406 9752 4410 9756
rect 4411 9752 4415 9756
rect 4396 9742 4400 9746
rect 4401 9742 4405 9746
rect 4406 9742 4410 9746
rect 4411 9742 4415 9746
rect 4396 9732 4400 9736
rect 4401 9732 4405 9736
rect 4406 9732 4410 9736
rect 4411 9732 4415 9736
rect 3859 9708 3863 9712
rect 3864 9708 3868 9712
rect 3869 9708 3873 9712
rect 3874 9708 3878 9712
rect 3879 9708 3883 9712
rect 3884 9708 3888 9712
rect 3889 9708 3893 9712
rect 3894 9708 3898 9712
rect 3899 9708 3903 9712
rect 3904 9708 3908 9712
rect 3909 9708 3913 9712
rect 3914 9708 3918 9712
rect 3919 9708 3923 9712
rect 3859 9703 3863 9707
rect 3864 9703 3868 9707
rect 3869 9703 3873 9707
rect 3874 9703 3878 9707
rect 3879 9703 3883 9707
rect 3884 9703 3888 9707
rect 3889 9703 3893 9707
rect 3894 9703 3898 9707
rect 3899 9703 3903 9707
rect 3904 9703 3908 9707
rect 3909 9703 3913 9707
rect 3914 9703 3918 9707
rect 3919 9703 3923 9707
rect 4041 9708 4045 9712
rect 4046 9708 4050 9712
rect 4051 9708 4055 9712
rect 4056 9708 4060 9712
rect 4061 9708 4065 9712
rect 4066 9708 4070 9712
rect 4071 9708 4075 9712
rect 4076 9708 4080 9712
rect 4081 9708 4085 9712
rect 4086 9708 4090 9712
rect 4091 9708 4095 9712
rect 4041 9703 4045 9707
rect 4046 9703 4050 9707
rect 4051 9703 4055 9707
rect 4056 9703 4060 9707
rect 4061 9703 4065 9707
rect 4066 9703 4070 9707
rect 4071 9703 4075 9707
rect 4076 9703 4080 9707
rect 4081 9703 4085 9707
rect 4086 9703 4090 9707
rect 4091 9703 4095 9707
rect 4100 9716 4104 9720
rect 4105 9716 4109 9720
rect 4110 9716 4114 9720
rect 4115 9716 4119 9720
rect 4100 9706 4104 9710
rect 4105 9706 4109 9710
rect 4110 9706 4114 9710
rect 4115 9706 4119 9710
rect 3482 9696 3486 9700
rect 3487 9696 3491 9700
rect 3492 9696 3496 9700
rect 3497 9696 3501 9700
rect 3482 9686 3486 9690
rect 3487 9686 3491 9690
rect 3492 9686 3496 9690
rect 3497 9686 3501 9690
rect 3791 9696 3795 9700
rect 3796 9696 3800 9700
rect 3801 9696 3805 9700
rect 3806 9696 3810 9700
rect 3791 9686 3795 9690
rect 3796 9686 3800 9690
rect 3801 9686 3805 9690
rect 3806 9686 3810 9690
rect 4100 9696 4104 9700
rect 4105 9696 4109 9700
rect 4110 9696 4114 9700
rect 4115 9696 4119 9700
rect 4100 9686 4104 9690
rect 4105 9686 4109 9690
rect 4110 9686 4114 9690
rect 4115 9686 4119 9690
rect 4292 9716 4296 9720
rect 4297 9716 4301 9720
rect 4302 9716 4306 9720
rect 4307 9716 4311 9720
rect 4292 9706 4296 9710
rect 4297 9706 4301 9710
rect 4302 9706 4306 9710
rect 4307 9706 4311 9710
rect 4292 9696 4296 9700
rect 4297 9696 4301 9700
rect 4302 9696 4306 9700
rect 4307 9696 4311 9700
rect 4292 9686 4296 9690
rect 4297 9686 4301 9690
rect 4302 9686 4306 9690
rect 4307 9686 4311 9690
rect 4318 9716 4322 9720
rect 4323 9716 4327 9720
rect 4328 9716 4332 9720
rect 4333 9716 4337 9720
rect 4318 9706 4322 9710
rect 4323 9706 4327 9710
rect 4328 9706 4332 9710
rect 4333 9706 4337 9710
rect 4318 9696 4322 9700
rect 4323 9696 4327 9700
rect 4328 9696 4332 9700
rect 4333 9696 4337 9700
rect 4318 9686 4322 9690
rect 4323 9686 4327 9690
rect 4328 9686 4332 9690
rect 4333 9686 4337 9690
rect 4344 9716 4348 9720
rect 4349 9716 4353 9720
rect 4354 9716 4358 9720
rect 4359 9716 4363 9720
rect 4344 9706 4348 9710
rect 4349 9706 4353 9710
rect 4354 9706 4358 9710
rect 4359 9706 4363 9710
rect 4344 9696 4348 9700
rect 4349 9696 4353 9700
rect 4354 9696 4358 9700
rect 4359 9696 4363 9700
rect 4344 9686 4348 9690
rect 4349 9686 4353 9690
rect 4354 9686 4358 9690
rect 4359 9686 4363 9690
rect 4370 9716 4374 9720
rect 4375 9716 4379 9720
rect 4380 9716 4384 9720
rect 4385 9716 4389 9720
rect 4370 9706 4374 9710
rect 4375 9706 4379 9710
rect 4380 9706 4384 9710
rect 4385 9706 4389 9710
rect 4370 9696 4374 9700
rect 4375 9696 4379 9700
rect 4380 9696 4384 9700
rect 4385 9696 4389 9700
rect 4370 9686 4374 9690
rect 4375 9686 4379 9690
rect 4380 9686 4384 9690
rect 4385 9686 4389 9690
rect 4396 9716 4400 9720
rect 4401 9716 4405 9720
rect 4406 9716 4410 9720
rect 4411 9716 4415 9720
rect 4396 9706 4400 9710
rect 4401 9706 4405 9710
rect 4406 9706 4410 9710
rect 4411 9706 4415 9710
rect 4396 9696 4400 9700
rect 4401 9696 4405 9700
rect 4406 9696 4410 9700
rect 4411 9696 4415 9700
rect 4396 9686 4400 9690
rect 4401 9686 4405 9690
rect 4406 9686 4410 9690
rect 4411 9686 4415 9690
rect 3343 9681 3347 9685
rect 3348 9681 3352 9685
rect 3343 9676 3347 9680
rect 3348 9676 3352 9680
rect 3343 9671 3347 9675
rect 3348 9671 3352 9675
rect 3343 9666 3347 9670
rect 3348 9666 3352 9670
rect 3343 9661 3347 9665
rect 3348 9661 3352 9665
rect 613 9618 617 9622
rect 623 9618 627 9622
rect 633 9618 637 9622
rect 643 9618 647 9622
rect 613 9613 617 9617
rect 623 9613 627 9617
rect 633 9613 637 9617
rect 643 9613 647 9617
rect 613 9608 617 9612
rect 623 9608 627 9612
rect 633 9608 637 9612
rect 643 9608 647 9612
rect 613 9603 617 9607
rect 623 9603 627 9607
rect 633 9603 637 9607
rect 643 9603 647 9607
rect 659 9618 663 9622
rect 669 9618 673 9622
rect 679 9618 683 9622
rect 689 9618 693 9622
rect 659 9613 663 9617
rect 669 9613 673 9617
rect 679 9613 683 9617
rect 689 9613 693 9617
rect 659 9608 663 9612
rect 669 9608 673 9612
rect 679 9608 683 9612
rect 689 9608 693 9612
rect 659 9603 663 9607
rect 669 9603 673 9607
rect 679 9603 683 9607
rect 689 9603 693 9607
rect 613 9592 617 9596
rect 623 9592 627 9596
rect 633 9592 637 9596
rect 643 9592 647 9596
rect 613 9587 617 9591
rect 623 9587 627 9591
rect 633 9587 637 9591
rect 643 9587 647 9591
rect 613 9582 617 9586
rect 623 9582 627 9586
rect 633 9582 637 9586
rect 643 9582 647 9586
rect 613 9577 617 9581
rect 623 9577 627 9581
rect 633 9577 637 9581
rect 643 9577 647 9581
rect 659 9592 663 9596
rect 669 9592 673 9596
rect 679 9592 683 9596
rect 689 9592 693 9596
rect 659 9587 663 9591
rect 669 9587 673 9591
rect 679 9587 683 9591
rect 689 9587 693 9591
rect 659 9582 663 9586
rect 669 9582 673 9586
rect 679 9582 683 9586
rect 689 9582 693 9586
rect 659 9577 663 9581
rect 669 9577 673 9581
rect 679 9577 683 9581
rect 689 9577 693 9581
rect 2258 9619 2262 9623
rect 613 9566 617 9570
rect 623 9566 627 9570
rect 633 9566 637 9570
rect 643 9566 647 9570
rect 613 9561 617 9565
rect 623 9561 627 9565
rect 633 9561 637 9565
rect 643 9561 647 9565
rect 613 9556 617 9560
rect 623 9556 627 9560
rect 633 9556 637 9560
rect 643 9556 647 9560
rect 613 9551 617 9555
rect 623 9551 627 9555
rect 633 9551 637 9555
rect 643 9551 647 9555
rect 659 9566 663 9570
rect 669 9566 673 9570
rect 679 9566 683 9570
rect 689 9566 693 9570
rect 659 9561 663 9565
rect 669 9561 673 9565
rect 679 9561 683 9565
rect 689 9561 693 9565
rect 659 9556 663 9560
rect 669 9556 673 9560
rect 679 9556 683 9560
rect 689 9556 693 9560
rect 659 9551 663 9555
rect 669 9551 673 9555
rect 679 9551 683 9555
rect 689 9551 693 9555
rect 613 9540 617 9544
rect 623 9540 627 9544
rect 633 9540 637 9544
rect 643 9540 647 9544
rect 613 9535 617 9539
rect 623 9535 627 9539
rect 633 9535 637 9539
rect 643 9535 647 9539
rect 613 9530 617 9534
rect 623 9530 627 9534
rect 633 9530 637 9534
rect 643 9530 647 9534
rect 613 9525 617 9529
rect 623 9525 627 9529
rect 633 9525 637 9529
rect 643 9525 647 9529
rect 659 9540 663 9544
rect 669 9540 673 9544
rect 679 9540 683 9544
rect 689 9540 693 9544
rect 659 9535 663 9539
rect 669 9535 673 9539
rect 679 9535 683 9539
rect 689 9535 693 9539
rect 659 9530 663 9534
rect 669 9530 673 9534
rect 679 9530 683 9534
rect 689 9530 693 9534
rect 659 9525 663 9529
rect 669 9525 673 9529
rect 679 9525 683 9529
rect 689 9525 693 9529
rect 613 9514 617 9518
rect 623 9514 627 9518
rect 633 9514 637 9518
rect 643 9514 647 9518
rect 613 9509 617 9513
rect 623 9509 627 9513
rect 633 9509 637 9513
rect 643 9509 647 9513
rect 613 9504 617 9508
rect 623 9504 627 9508
rect 633 9504 637 9508
rect 643 9504 647 9508
rect 613 9499 617 9503
rect 623 9499 627 9503
rect 633 9499 637 9503
rect 643 9499 647 9503
rect 659 9514 663 9518
rect 669 9514 673 9518
rect 679 9514 683 9518
rect 689 9514 693 9518
rect 659 9509 663 9513
rect 669 9509 673 9513
rect 679 9509 683 9513
rect 689 9509 693 9513
rect 659 9504 663 9508
rect 669 9504 673 9508
rect 679 9504 683 9508
rect 689 9504 693 9508
rect 659 9499 663 9503
rect 669 9499 673 9503
rect 679 9499 683 9503
rect 689 9499 693 9503
rect 613 9321 617 9325
rect 623 9321 627 9325
rect 633 9321 637 9325
rect 643 9321 647 9325
rect 613 9316 617 9320
rect 623 9316 627 9320
rect 633 9316 637 9320
rect 643 9316 647 9320
rect 613 9311 617 9315
rect 623 9311 627 9315
rect 633 9311 637 9315
rect 643 9311 647 9315
rect 613 9306 617 9310
rect 623 9306 627 9310
rect 633 9306 637 9310
rect 643 9306 647 9310
rect 659 9321 663 9325
rect 669 9321 673 9325
rect 679 9321 683 9325
rect 689 9321 693 9325
rect 659 9316 663 9320
rect 669 9316 673 9320
rect 679 9316 683 9320
rect 689 9316 693 9320
rect 659 9311 663 9315
rect 669 9311 673 9315
rect 679 9311 683 9315
rect 689 9311 693 9315
rect 659 9306 663 9310
rect 669 9306 673 9310
rect 679 9306 683 9310
rect 689 9306 693 9310
rect 613 9012 617 9016
rect 623 9012 627 9016
rect 633 9012 637 9016
rect 643 9012 647 9016
rect 613 9007 617 9011
rect 623 9007 627 9011
rect 633 9007 637 9011
rect 643 9007 647 9011
rect 613 9002 617 9006
rect 623 9002 627 9006
rect 633 9002 637 9006
rect 643 9002 647 9006
rect 613 8997 617 9001
rect 623 8997 627 9001
rect 633 8997 637 9001
rect 643 8997 647 9001
rect 659 9012 663 9016
rect 669 9012 673 9016
rect 679 9012 683 9016
rect 689 9012 693 9016
rect 659 9007 663 9011
rect 669 9007 673 9011
rect 679 9007 683 9011
rect 689 9007 693 9011
rect 659 9002 663 9006
rect 669 9002 673 9006
rect 679 9002 683 9006
rect 689 9002 693 9006
rect 659 8997 663 9001
rect 669 8997 673 9001
rect 679 8997 683 9001
rect 689 8997 693 9001
rect 4479 9573 4483 9577
rect 4489 9573 4493 9577
rect 4499 9573 4503 9577
rect 4509 9573 4513 9577
rect 4479 9568 4483 9572
rect 4489 9568 4493 9572
rect 4499 9568 4503 9572
rect 4509 9568 4513 9572
rect 4479 9563 4483 9567
rect 4489 9563 4493 9567
rect 4499 9563 4503 9567
rect 4509 9563 4513 9567
rect 4479 9558 4483 9562
rect 4489 9558 4493 9562
rect 4499 9558 4503 9562
rect 4509 9558 4513 9562
rect 4525 9573 4529 9577
rect 4535 9573 4539 9577
rect 4545 9573 4549 9577
rect 4555 9573 4559 9577
rect 4525 9568 4529 9572
rect 4535 9568 4539 9572
rect 4545 9568 4549 9572
rect 4555 9568 4559 9572
rect 4525 9563 4529 9567
rect 4535 9563 4539 9567
rect 4545 9563 4549 9567
rect 4555 9563 4559 9567
rect 4525 9558 4529 9562
rect 4535 9558 4539 9562
rect 4545 9558 4549 9562
rect 4555 9558 4559 9562
rect 4479 9544 4483 9548
rect 4489 9544 4493 9548
rect 4499 9544 4503 9548
rect 4509 9544 4513 9548
rect 4479 9539 4483 9543
rect 4489 9539 4493 9543
rect 4499 9539 4503 9543
rect 4509 9539 4513 9543
rect 4479 9534 4483 9538
rect 4489 9534 4493 9538
rect 4499 9534 4503 9538
rect 4509 9534 4513 9538
rect 4479 9529 4483 9533
rect 4489 9529 4493 9533
rect 4499 9529 4503 9533
rect 4509 9529 4513 9533
rect 4525 9544 4529 9548
rect 4535 9544 4539 9548
rect 4545 9544 4549 9548
rect 4555 9544 4559 9548
rect 4525 9539 4529 9543
rect 4535 9539 4539 9543
rect 4545 9539 4549 9543
rect 4555 9539 4559 9543
rect 4525 9534 4529 9538
rect 4535 9534 4539 9538
rect 4545 9534 4549 9538
rect 4555 9534 4559 9538
rect 4525 9529 4529 9533
rect 4535 9529 4539 9533
rect 4545 9529 4549 9533
rect 4555 9529 4559 9533
rect 4479 9515 4483 9519
rect 4489 9515 4493 9519
rect 4499 9515 4503 9519
rect 4509 9515 4513 9519
rect 4479 9510 4483 9514
rect 4489 9510 4493 9514
rect 4499 9510 4503 9514
rect 4509 9510 4513 9514
rect 4479 9505 4483 9509
rect 4489 9505 4493 9509
rect 4499 9505 4503 9509
rect 4509 9505 4513 9509
rect 4479 9500 4483 9504
rect 4489 9500 4493 9504
rect 4499 9500 4503 9504
rect 4509 9500 4513 9504
rect 4525 9515 4529 9519
rect 4535 9515 4539 9519
rect 4545 9515 4549 9519
rect 4555 9515 4559 9519
rect 4525 9510 4529 9514
rect 4535 9510 4539 9514
rect 4545 9510 4549 9514
rect 4555 9510 4559 9514
rect 4525 9505 4529 9509
rect 4535 9505 4539 9509
rect 4545 9505 4549 9509
rect 4555 9505 4559 9509
rect 4525 9500 4529 9504
rect 4535 9500 4539 9504
rect 4545 9500 4549 9504
rect 4555 9500 4559 9504
rect 2367 8774 2371 8778
rect 613 8703 617 8707
rect 623 8703 627 8707
rect 633 8703 637 8707
rect 643 8703 647 8707
rect 613 8698 617 8702
rect 623 8698 627 8702
rect 633 8698 637 8702
rect 643 8698 647 8702
rect 613 8693 617 8697
rect 623 8693 627 8697
rect 633 8693 637 8697
rect 643 8693 647 8697
rect 613 8688 617 8692
rect 623 8688 627 8692
rect 633 8688 637 8692
rect 643 8688 647 8692
rect 659 8703 663 8707
rect 669 8703 673 8707
rect 679 8703 683 8707
rect 689 8703 693 8707
rect 659 8698 663 8702
rect 669 8698 673 8702
rect 679 8698 683 8702
rect 689 8698 693 8702
rect 659 8693 663 8697
rect 669 8693 673 8697
rect 679 8693 683 8697
rect 689 8693 693 8697
rect 659 8688 663 8692
rect 669 8688 673 8692
rect 679 8688 683 8692
rect 689 8688 693 8692
rect 2624 9277 2628 9281
rect 613 8394 617 8398
rect 623 8394 627 8398
rect 633 8394 637 8398
rect 643 8394 647 8398
rect 613 8389 617 8393
rect 623 8389 627 8393
rect 633 8389 637 8393
rect 643 8389 647 8393
rect 613 8384 617 8388
rect 623 8384 627 8388
rect 633 8384 637 8388
rect 643 8384 647 8388
rect 613 8379 617 8383
rect 623 8379 627 8383
rect 633 8379 637 8383
rect 643 8379 647 8383
rect 659 8394 663 8398
rect 669 8394 673 8398
rect 679 8394 683 8398
rect 689 8394 693 8398
rect 659 8389 663 8393
rect 669 8389 673 8393
rect 679 8389 683 8393
rect 689 8389 693 8393
rect 659 8384 663 8388
rect 669 8384 673 8388
rect 679 8384 683 8388
rect 689 8384 693 8388
rect 659 8379 663 8383
rect 669 8379 673 8383
rect 679 8379 683 8383
rect 689 8379 693 8383
rect 2623 9174 2627 9178
rect 613 8085 617 8089
rect 623 8085 627 8089
rect 633 8085 637 8089
rect 643 8085 647 8089
rect 613 8080 617 8084
rect 623 8080 627 8084
rect 633 8080 637 8084
rect 643 8080 647 8084
rect 613 8075 617 8079
rect 623 8075 627 8079
rect 633 8075 637 8079
rect 643 8075 647 8079
rect 613 8070 617 8074
rect 623 8070 627 8074
rect 633 8070 637 8074
rect 643 8070 647 8074
rect 659 8085 663 8089
rect 669 8085 673 8089
rect 679 8085 683 8089
rect 689 8085 693 8089
rect 659 8080 663 8084
rect 669 8080 673 8084
rect 679 8080 683 8084
rect 689 8080 693 8084
rect 659 8075 663 8079
rect 669 8075 673 8079
rect 679 8075 683 8079
rect 689 8075 693 8079
rect 659 8070 663 8074
rect 669 8070 673 8074
rect 679 8070 683 8074
rect 689 8070 693 8074
rect 2367 7792 2371 7796
rect 613 7776 617 7780
rect 623 7776 627 7780
rect 633 7776 637 7780
rect 643 7776 647 7780
rect 613 7771 617 7775
rect 623 7771 627 7775
rect 633 7771 637 7775
rect 643 7771 647 7775
rect 613 7766 617 7770
rect 623 7766 627 7770
rect 633 7766 637 7770
rect 643 7766 647 7770
rect 613 7761 617 7765
rect 623 7761 627 7765
rect 633 7761 637 7765
rect 643 7761 647 7765
rect 659 7776 663 7780
rect 669 7776 673 7780
rect 679 7776 683 7780
rect 689 7776 693 7780
rect 659 7771 663 7775
rect 669 7771 673 7775
rect 679 7771 683 7775
rect 689 7771 693 7775
rect 659 7766 663 7770
rect 669 7766 673 7770
rect 679 7766 683 7770
rect 689 7766 693 7770
rect 659 7761 663 7765
rect 669 7761 673 7765
rect 679 7761 683 7765
rect 689 7761 693 7765
rect 2756 8407 2760 8411
rect 2624 8295 2628 8299
rect 613 7467 617 7471
rect 623 7467 627 7471
rect 633 7467 637 7471
rect 643 7467 647 7471
rect 613 7462 617 7466
rect 623 7462 627 7466
rect 633 7462 637 7466
rect 643 7462 647 7466
rect 613 7457 617 7461
rect 623 7457 627 7461
rect 633 7457 637 7461
rect 643 7457 647 7461
rect 613 7452 617 7456
rect 623 7452 627 7456
rect 633 7452 637 7456
rect 643 7452 647 7456
rect 659 7467 663 7471
rect 669 7467 673 7471
rect 679 7467 683 7471
rect 689 7467 693 7471
rect 659 7462 663 7466
rect 669 7462 673 7466
rect 679 7462 683 7466
rect 689 7462 693 7466
rect 659 7457 663 7461
rect 669 7457 673 7461
rect 679 7457 683 7461
rect 689 7457 693 7461
rect 659 7452 663 7456
rect 669 7452 673 7456
rect 679 7452 683 7456
rect 689 7452 693 7456
rect 2623 8192 2627 8196
rect 2756 7425 2760 7429
rect 2847 9313 2851 9317
rect 2887 9230 2892 9235
rect 2898 9226 2903 9231
rect 2921 9235 2926 9240
rect 2945 9230 2950 9235
rect 2960 9234 2965 9240
rect 2990 9230 2995 9235
rect 3019 9229 3024 9234
rect 2974 9224 2979 9229
rect 3003 9224 3007 9229
rect 3045 9223 3050 9228
rect 2851 9170 2856 9175
rect 2887 9163 2892 9168
rect 2898 9167 2903 9172
rect 2921 9158 2926 9163
rect 2945 9163 2950 9168
rect 2974 9169 2979 9174
rect 3003 9169 3007 9174
rect 2960 9158 2965 9164
rect 2990 9163 2995 9168
rect 3019 9164 3024 9169
rect 3045 9164 3050 9169
rect 2850 9101 2855 9106
rect 2887 9098 2892 9103
rect 2898 9094 2903 9099
rect 2921 9103 2926 9108
rect 2945 9098 2950 9103
rect 3101 9229 3106 9234
rect 2960 9102 2965 9108
rect 2990 9098 2995 9103
rect 3019 9097 3024 9102
rect 2974 9092 2979 9097
rect 3003 9092 3007 9097
rect 3045 9091 3050 9096
rect 2851 9038 2856 9043
rect 2887 9031 2892 9036
rect 2898 9035 2903 9040
rect 2921 9026 2926 9031
rect 2945 9031 2950 9036
rect 2974 9037 2979 9042
rect 3003 9037 3007 9042
rect 2960 9026 2965 9032
rect 2990 9031 2995 9036
rect 3019 9032 3024 9037
rect 3044 9033 3049 9038
rect 2850 8969 2855 8974
rect 2887 8966 2892 8971
rect 2898 8962 2903 8967
rect 2921 8971 2926 8976
rect 2945 8966 2950 8971
rect 2960 8970 2965 8976
rect 2990 8966 2995 8971
rect 3019 8965 3024 8970
rect 2974 8960 2979 8965
rect 3003 8960 3007 8965
rect 3045 8959 3050 8964
rect 3101 9105 3106 9110
rect 3126 9223 3131 9228
rect 3125 9164 3130 9169
rect 3186 9229 3191 9234
rect 3150 9091 3155 9096
rect 3150 9033 3155 9038
rect 2851 8906 2856 8911
rect 2887 8899 2892 8904
rect 2898 8903 2903 8908
rect 2921 8894 2926 8899
rect 2945 8899 2950 8904
rect 2974 8905 2979 8910
rect 3003 8905 3007 8910
rect 2960 8894 2965 8900
rect 2990 8899 2995 8904
rect 3019 8900 3024 8905
rect 3045 8898 3050 8903
rect 2850 8837 2855 8842
rect 2887 8834 2892 8839
rect 2898 8830 2903 8835
rect 2921 8839 2926 8844
rect 2945 8834 2950 8839
rect 2960 8838 2965 8844
rect 2990 8834 2995 8839
rect 3019 8833 3024 8838
rect 2974 8828 2979 8833
rect 3003 8828 3007 8833
rect 3045 8827 3050 8832
rect 3101 8965 3106 8970
rect 3126 8959 3131 8964
rect 3125 8898 3130 8903
rect 3303 9262 3307 9266
rect 3208 9102 3213 9107
rect 3569 9277 3573 9281
rect 3568 9174 3572 9178
rect 3443 9135 3448 9140
rect 3560 9136 3565 9141
rect 3183 8974 3188 8979
rect 3217 8967 3222 8972
rect 3214 8894 3219 8899
rect 2851 8774 2856 8779
rect 2887 8767 2892 8772
rect 2898 8771 2903 8776
rect 2921 8762 2926 8767
rect 2945 8767 2950 8772
rect 2974 8773 2979 8778
rect 3003 8773 3007 8778
rect 2960 8762 2965 8768
rect 2990 8767 2995 8772
rect 3019 8768 3024 8773
rect 3044 8762 3049 8767
rect 3101 8841 3106 8846
rect 3089 8773 3094 8778
rect 3148 8767 3153 8772
rect 3159 8771 3164 8776
rect 3182 8762 3187 8767
rect 3206 8767 3211 8772
rect 3235 8773 3240 8778
rect 3264 8773 3268 8778
rect 3221 8762 3226 8768
rect 3251 8767 3256 8772
rect 3276 8773 3281 8778
rect 3443 8819 3448 8824
rect 3312 8774 3316 8778
rect 3150 8662 3154 8666
rect 3560 8818 3565 8823
rect 3275 8580 3279 8584
rect 2847 8331 2851 8335
rect 2849 8251 2854 8256
rect 2887 8248 2892 8253
rect 2898 8244 2903 8249
rect 2921 8253 2926 8258
rect 2945 8248 2950 8253
rect 2960 8252 2965 8258
rect 2990 8248 2995 8253
rect 3019 8247 3024 8252
rect 2974 8242 2979 8247
rect 3003 8242 3007 8247
rect 3045 8241 3050 8246
rect 2851 8188 2856 8193
rect 2887 8181 2892 8186
rect 2898 8185 2903 8190
rect 2921 8176 2926 8181
rect 2945 8181 2950 8186
rect 2974 8187 2979 8192
rect 3003 8187 3007 8192
rect 2960 8176 2965 8182
rect 2990 8181 2995 8186
rect 3019 8182 3024 8187
rect 3045 8182 3050 8187
rect 2850 8119 2855 8124
rect 2887 8116 2892 8121
rect 2898 8112 2903 8117
rect 2921 8121 2926 8126
rect 2945 8116 2950 8121
rect 3101 8247 3106 8252
rect 2960 8120 2965 8126
rect 2990 8116 2995 8121
rect 3019 8115 3024 8120
rect 2974 8110 2979 8115
rect 3003 8110 3007 8115
rect 3045 8109 3050 8114
rect 2851 8056 2856 8061
rect 2887 8049 2892 8054
rect 2898 8053 2903 8058
rect 2921 8044 2926 8049
rect 2945 8049 2950 8054
rect 2974 8055 2979 8060
rect 3003 8055 3007 8060
rect 2960 8044 2965 8050
rect 2990 8049 2995 8054
rect 3019 8050 3024 8055
rect 3044 8051 3049 8056
rect 2850 7987 2855 7992
rect 2887 7984 2892 7989
rect 2898 7980 2903 7985
rect 2921 7989 2926 7994
rect 2945 7984 2950 7989
rect 2960 7988 2965 7994
rect 2990 7984 2995 7989
rect 3019 7983 3024 7988
rect 2974 7978 2979 7983
rect 3003 7978 3007 7983
rect 3045 7977 3050 7982
rect 3101 8123 3106 8128
rect 3126 8241 3131 8246
rect 3125 8182 3130 8187
rect 3186 8247 3191 8252
rect 3150 8109 3155 8114
rect 3150 8051 3155 8056
rect 2851 7924 2856 7929
rect 2887 7917 2892 7922
rect 2898 7921 2903 7926
rect 2921 7912 2926 7917
rect 2945 7917 2950 7922
rect 2974 7923 2979 7928
rect 3003 7923 3007 7928
rect 2960 7912 2965 7918
rect 2990 7917 2995 7922
rect 3019 7918 3024 7923
rect 3045 7916 3050 7921
rect 2850 7855 2855 7860
rect 2887 7852 2892 7857
rect 2898 7848 2903 7853
rect 2921 7857 2926 7862
rect 2945 7852 2950 7857
rect 2960 7856 2965 7862
rect 2990 7852 2995 7857
rect 3019 7851 3024 7856
rect 2974 7846 2979 7851
rect 3003 7846 3007 7851
rect 3045 7845 3050 7850
rect 3101 7983 3106 7988
rect 3126 7977 3131 7982
rect 3125 7916 3130 7921
rect 3303 8280 3307 8284
rect 3208 8120 3213 8125
rect 3183 7992 3188 7997
rect 3217 7985 3222 7990
rect 3214 7912 3219 7917
rect 2851 7792 2856 7797
rect 2887 7785 2892 7790
rect 2898 7789 2903 7794
rect 2921 7780 2926 7785
rect 2945 7785 2950 7790
rect 2974 7791 2979 7796
rect 3003 7791 3007 7796
rect 2960 7780 2965 7786
rect 2990 7785 2995 7790
rect 3019 7786 3024 7791
rect 3044 7780 3049 7785
rect 3101 7859 3106 7864
rect 3089 7791 3094 7796
rect 3148 7785 3153 7790
rect 3159 7789 3164 7794
rect 3182 7780 3187 7785
rect 3206 7785 3211 7790
rect 3235 7791 3240 7796
rect 3264 7791 3268 7796
rect 3221 7780 3226 7786
rect 3251 7785 3256 7790
rect 3276 7791 3281 7796
rect 3312 7792 3316 7796
rect 3150 7680 3154 7684
rect 3701 8407 3705 8411
rect 3569 8296 3573 8300
rect 3275 7598 3279 7602
rect 3568 8192 3572 8196
rect 3701 7425 3705 7429
rect 4479 9486 4483 9490
rect 4489 9486 4493 9490
rect 4499 9486 4503 9490
rect 4509 9486 4513 9490
rect 4479 9481 4483 9485
rect 4489 9481 4493 9485
rect 4499 9481 4503 9485
rect 4509 9481 4513 9485
rect 4479 9476 4483 9480
rect 4489 9476 4493 9480
rect 4499 9476 4503 9480
rect 4509 9476 4513 9480
rect 4479 9471 4483 9475
rect 4489 9471 4493 9475
rect 4499 9471 4503 9475
rect 4509 9471 4513 9475
rect 4525 9486 4529 9490
rect 4535 9486 4539 9490
rect 4545 9486 4549 9490
rect 4555 9486 4559 9490
rect 4525 9481 4529 9485
rect 4535 9481 4539 9485
rect 4545 9481 4549 9485
rect 4555 9481 4559 9485
rect 4525 9476 4529 9480
rect 4535 9476 4539 9480
rect 4545 9476 4549 9480
rect 4555 9476 4559 9480
rect 4525 9471 4529 9475
rect 4535 9471 4539 9475
rect 4545 9471 4549 9475
rect 4555 9471 4559 9475
rect 4479 9457 4483 9461
rect 4489 9457 4493 9461
rect 4499 9457 4503 9461
rect 4509 9457 4513 9461
rect 4479 9452 4483 9456
rect 4489 9452 4493 9456
rect 4499 9452 4503 9456
rect 4509 9452 4513 9456
rect 4479 9447 4483 9451
rect 4489 9447 4493 9451
rect 4499 9447 4503 9451
rect 4509 9447 4513 9451
rect 4479 9442 4483 9446
rect 4489 9442 4493 9446
rect 4499 9442 4503 9446
rect 4509 9442 4513 9446
rect 4525 9457 4529 9461
rect 4535 9457 4539 9461
rect 4545 9457 4549 9461
rect 4555 9457 4559 9461
rect 4525 9452 4529 9456
rect 4535 9452 4539 9456
rect 4545 9452 4549 9456
rect 4555 9452 4559 9456
rect 4525 9447 4529 9451
rect 4535 9447 4539 9451
rect 4545 9447 4549 9451
rect 4555 9447 4559 9451
rect 4525 9442 4529 9446
rect 4535 9442 4539 9446
rect 4545 9442 4549 9446
rect 4555 9442 4559 9446
rect 3792 9313 3796 9317
rect 3793 9233 3798 9238
rect 3832 9230 3837 9235
rect 3843 9226 3848 9231
rect 3866 9235 3871 9240
rect 3890 9230 3895 9235
rect 3905 9234 3910 9240
rect 3935 9230 3940 9235
rect 3964 9229 3969 9234
rect 3919 9224 3924 9229
rect 3948 9224 3952 9229
rect 3990 9223 3995 9228
rect 3796 9170 3801 9175
rect 3832 9163 3837 9168
rect 3843 9167 3848 9172
rect 3866 9158 3871 9163
rect 3890 9163 3895 9168
rect 3919 9169 3924 9174
rect 3948 9169 3952 9174
rect 3905 9158 3910 9164
rect 3935 9163 3940 9168
rect 3964 9164 3969 9169
rect 3990 9164 3995 9169
rect 3795 9101 3800 9106
rect 3832 9098 3837 9103
rect 3843 9094 3848 9099
rect 3866 9103 3871 9108
rect 3890 9098 3895 9103
rect 4046 9229 4051 9234
rect 3905 9102 3910 9108
rect 3935 9098 3940 9103
rect 3964 9097 3969 9102
rect 3919 9092 3924 9097
rect 3948 9092 3952 9097
rect 3990 9091 3995 9096
rect 3796 9038 3801 9043
rect 3832 9031 3837 9036
rect 3843 9035 3848 9040
rect 3866 9026 3871 9031
rect 3890 9031 3895 9036
rect 3919 9037 3924 9042
rect 3948 9037 3952 9042
rect 3905 9026 3910 9032
rect 3935 9031 3940 9036
rect 3964 9032 3969 9037
rect 3989 9033 3994 9038
rect 3795 8969 3800 8974
rect 3832 8966 3837 8971
rect 3843 8962 3848 8967
rect 3866 8971 3871 8976
rect 3890 8966 3895 8971
rect 3905 8970 3910 8976
rect 3935 8966 3940 8971
rect 3964 8965 3969 8970
rect 3919 8960 3924 8965
rect 3948 8960 3952 8965
rect 3990 8959 3995 8964
rect 4046 9105 4051 9110
rect 4071 9223 4076 9228
rect 4070 9164 4075 9169
rect 4131 9229 4136 9234
rect 4095 9091 4100 9096
rect 4095 9033 4100 9038
rect 3796 8906 3801 8911
rect 3832 8899 3837 8904
rect 3843 8903 3848 8908
rect 3866 8894 3871 8899
rect 3890 8899 3895 8904
rect 3919 8905 3924 8910
rect 3948 8905 3952 8910
rect 3905 8894 3910 8900
rect 3935 8899 3940 8904
rect 3964 8900 3969 8905
rect 3990 8898 3995 8903
rect 3795 8837 3800 8842
rect 3832 8834 3837 8839
rect 3843 8830 3848 8835
rect 3866 8839 3871 8844
rect 3890 8834 3895 8839
rect 3905 8838 3910 8844
rect 3935 8834 3940 8839
rect 3964 8833 3969 8838
rect 3919 8828 3924 8833
rect 3948 8828 3952 8833
rect 3990 8827 3995 8832
rect 4046 8965 4051 8970
rect 4071 8959 4076 8964
rect 4070 8898 4075 8903
rect 4248 9262 4252 9266
rect 4153 9102 4158 9107
rect 4479 9056 4483 9060
rect 4489 9056 4493 9060
rect 4499 9056 4503 9060
rect 4509 9056 4513 9060
rect 4479 9051 4483 9055
rect 4489 9051 4493 9055
rect 4499 9051 4503 9055
rect 4509 9051 4513 9055
rect 4479 9046 4483 9050
rect 4489 9046 4493 9050
rect 4499 9046 4503 9050
rect 4509 9046 4513 9050
rect 4479 9041 4483 9045
rect 4489 9041 4493 9045
rect 4499 9041 4503 9045
rect 4509 9041 4513 9045
rect 4525 9056 4529 9060
rect 4535 9056 4539 9060
rect 4545 9056 4549 9060
rect 4555 9056 4559 9060
rect 4525 9051 4529 9055
rect 4535 9051 4539 9055
rect 4545 9051 4549 9055
rect 4555 9051 4559 9055
rect 4525 9046 4529 9050
rect 4535 9046 4539 9050
rect 4545 9046 4549 9050
rect 4555 9046 4559 9050
rect 4525 9041 4529 9045
rect 4535 9041 4539 9045
rect 4545 9041 4549 9045
rect 4555 9041 4559 9045
rect 4128 8974 4133 8979
rect 4162 8967 4167 8972
rect 4159 8894 4164 8899
rect 3796 8774 3801 8779
rect 3832 8767 3837 8772
rect 3843 8771 3848 8776
rect 3866 8762 3871 8767
rect 3890 8767 3895 8772
rect 3919 8773 3924 8778
rect 3948 8773 3952 8778
rect 3905 8762 3910 8768
rect 3935 8767 3940 8772
rect 3964 8768 3969 8773
rect 3989 8762 3994 8767
rect 4046 8841 4051 8846
rect 4034 8773 4039 8778
rect 4093 8767 4098 8772
rect 4104 8771 4109 8776
rect 4127 8762 4132 8767
rect 4151 8767 4156 8772
rect 4180 8773 4185 8778
rect 4209 8773 4213 8778
rect 4166 8762 4171 8768
rect 4196 8767 4201 8772
rect 4221 8773 4226 8778
rect 4479 8747 4483 8751
rect 4489 8747 4493 8751
rect 4499 8747 4503 8751
rect 4509 8747 4513 8751
rect 4479 8742 4483 8746
rect 4489 8742 4493 8746
rect 4499 8742 4503 8746
rect 4509 8742 4513 8746
rect 4479 8737 4483 8741
rect 4489 8737 4493 8741
rect 4499 8737 4503 8741
rect 4509 8737 4513 8741
rect 4479 8732 4483 8736
rect 4489 8732 4493 8736
rect 4499 8732 4503 8736
rect 4509 8732 4513 8736
rect 4525 8747 4529 8751
rect 4535 8747 4539 8751
rect 4545 8747 4549 8751
rect 4555 8747 4559 8751
rect 4525 8742 4529 8746
rect 4535 8742 4539 8746
rect 4545 8742 4549 8746
rect 4555 8742 4559 8746
rect 4525 8737 4529 8741
rect 4535 8737 4539 8741
rect 4545 8737 4549 8741
rect 4555 8737 4559 8741
rect 4525 8732 4529 8736
rect 4535 8732 4539 8736
rect 4545 8732 4549 8736
rect 4555 8732 4559 8736
rect 4095 8662 4099 8666
rect 4220 8580 4224 8584
rect 4479 8438 4483 8442
rect 4489 8438 4493 8442
rect 4499 8438 4503 8442
rect 4509 8438 4513 8442
rect 4479 8433 4483 8437
rect 4489 8433 4493 8437
rect 4499 8433 4503 8437
rect 4509 8433 4513 8437
rect 4479 8428 4483 8432
rect 4489 8428 4493 8432
rect 4499 8428 4503 8432
rect 4509 8428 4513 8432
rect 4479 8423 4483 8427
rect 4489 8423 4493 8427
rect 4499 8423 4503 8427
rect 4509 8423 4513 8427
rect 4525 8438 4529 8442
rect 4535 8438 4539 8442
rect 4545 8438 4549 8442
rect 4555 8438 4559 8442
rect 4525 8433 4529 8437
rect 4535 8433 4539 8437
rect 4545 8433 4549 8437
rect 4555 8433 4559 8437
rect 4525 8428 4529 8432
rect 4535 8428 4539 8432
rect 4545 8428 4549 8432
rect 4555 8428 4559 8432
rect 4525 8423 4529 8427
rect 4535 8423 4539 8427
rect 4545 8423 4549 8427
rect 4555 8423 4559 8427
rect 3792 8331 3796 8335
rect 3794 8251 3799 8256
rect 3832 8248 3837 8253
rect 3843 8244 3848 8249
rect 3866 8253 3871 8258
rect 3890 8248 3895 8253
rect 3905 8252 3910 8258
rect 3935 8248 3940 8253
rect 3964 8247 3969 8252
rect 3919 8242 3924 8247
rect 3948 8242 3952 8247
rect 3990 8241 3995 8246
rect 3796 8188 3801 8193
rect 3832 8181 3837 8186
rect 3843 8185 3848 8190
rect 3866 8176 3871 8181
rect 3890 8181 3895 8186
rect 3919 8187 3924 8192
rect 3948 8187 3952 8192
rect 3905 8176 3910 8182
rect 3935 8181 3940 8186
rect 3964 8182 3969 8187
rect 3990 8182 3995 8187
rect 3795 8119 3800 8124
rect 3832 8116 3837 8121
rect 3843 8112 3848 8117
rect 3866 8121 3871 8126
rect 3890 8116 3895 8121
rect 4046 8247 4051 8252
rect 3905 8120 3910 8126
rect 3935 8116 3940 8121
rect 3964 8115 3969 8120
rect 3919 8110 3924 8115
rect 3948 8110 3952 8115
rect 3990 8109 3995 8114
rect 3796 8056 3801 8061
rect 3832 8049 3837 8054
rect 3843 8053 3848 8058
rect 3866 8044 3871 8049
rect 3890 8049 3895 8054
rect 3919 8055 3924 8060
rect 3948 8055 3952 8060
rect 3905 8044 3910 8050
rect 3935 8049 3940 8054
rect 3964 8050 3969 8055
rect 3989 8051 3994 8056
rect 3795 7987 3800 7992
rect 3832 7984 3837 7989
rect 3843 7980 3848 7985
rect 3866 7989 3871 7994
rect 3890 7984 3895 7989
rect 3905 7988 3910 7994
rect 3935 7984 3940 7989
rect 3964 7983 3969 7988
rect 3919 7978 3924 7983
rect 3948 7978 3952 7983
rect 3990 7977 3995 7982
rect 4046 8123 4051 8128
rect 4071 8241 4076 8246
rect 4070 8182 4075 8187
rect 4131 8247 4136 8252
rect 4095 8109 4100 8114
rect 4095 8051 4100 8056
rect 3796 7924 3801 7929
rect 3832 7917 3837 7922
rect 3843 7921 3848 7926
rect 3866 7912 3871 7917
rect 3890 7917 3895 7922
rect 3919 7923 3924 7928
rect 3948 7923 3952 7928
rect 3905 7912 3910 7918
rect 3935 7917 3940 7922
rect 3964 7918 3969 7923
rect 3990 7916 3995 7921
rect 3795 7855 3800 7860
rect 3832 7852 3837 7857
rect 3843 7848 3848 7853
rect 3866 7857 3871 7862
rect 3890 7852 3895 7857
rect 3905 7856 3910 7862
rect 3935 7852 3940 7857
rect 3964 7851 3969 7856
rect 3919 7846 3924 7851
rect 3948 7846 3952 7851
rect 3990 7845 3995 7850
rect 4046 7983 4051 7988
rect 4071 7977 4076 7982
rect 4070 7916 4075 7921
rect 4248 8280 4252 8284
rect 4479 8129 4483 8133
rect 4489 8129 4493 8133
rect 4499 8129 4503 8133
rect 4509 8129 4513 8133
rect 4153 8120 4158 8125
rect 4479 8124 4483 8128
rect 4489 8124 4493 8128
rect 4499 8124 4503 8128
rect 4509 8124 4513 8128
rect 4479 8119 4483 8123
rect 4489 8119 4493 8123
rect 4499 8119 4503 8123
rect 4509 8119 4513 8123
rect 4479 8114 4483 8118
rect 4489 8114 4493 8118
rect 4499 8114 4503 8118
rect 4509 8114 4513 8118
rect 4525 8129 4529 8133
rect 4535 8129 4539 8133
rect 4545 8129 4549 8133
rect 4555 8129 4559 8133
rect 4525 8124 4529 8128
rect 4535 8124 4539 8128
rect 4545 8124 4549 8128
rect 4555 8124 4559 8128
rect 4525 8119 4529 8123
rect 4535 8119 4539 8123
rect 4545 8119 4549 8123
rect 4555 8119 4559 8123
rect 4525 8114 4529 8118
rect 4535 8114 4539 8118
rect 4545 8114 4549 8118
rect 4555 8114 4559 8118
rect 4479 8098 4483 8102
rect 4489 8098 4493 8102
rect 4499 8098 4503 8102
rect 4509 8098 4513 8102
rect 4479 8093 4483 8097
rect 4489 8093 4493 8097
rect 4499 8093 4503 8097
rect 4509 8093 4513 8097
rect 4479 8088 4483 8092
rect 4489 8088 4493 8092
rect 4499 8088 4503 8092
rect 4509 8088 4513 8092
rect 4479 8083 4483 8087
rect 4489 8083 4493 8087
rect 4499 8083 4503 8087
rect 4509 8083 4513 8087
rect 4525 8098 4529 8102
rect 4535 8098 4539 8102
rect 4545 8098 4549 8102
rect 4555 8098 4559 8102
rect 4525 8093 4529 8097
rect 4535 8093 4539 8097
rect 4545 8093 4549 8097
rect 4555 8093 4559 8097
rect 4525 8088 4529 8092
rect 4535 8088 4539 8092
rect 4545 8088 4549 8092
rect 4555 8088 4559 8092
rect 4525 8083 4529 8087
rect 4535 8083 4539 8087
rect 4545 8083 4549 8087
rect 4555 8083 4559 8087
rect 4496 8074 4500 8078
rect 4501 8074 4505 8078
rect 4496 8069 4500 8073
rect 4501 8069 4505 8073
rect 4496 8064 4500 8068
rect 4501 8064 4505 8068
rect 4496 8059 4500 8063
rect 4501 8059 4505 8063
rect 4496 8054 4500 8058
rect 4501 8054 4505 8058
rect 4496 8049 4500 8053
rect 4501 8049 4505 8053
rect 4496 8044 4500 8048
rect 4501 8044 4505 8048
rect 4496 8039 4500 8043
rect 4501 8039 4505 8043
rect 4496 8034 4500 8038
rect 4501 8034 4505 8038
rect 4496 8029 4500 8033
rect 4501 8029 4505 8033
rect 4496 8024 4500 8028
rect 4501 8024 4505 8028
rect 4128 7992 4133 7997
rect 4162 7985 4167 7990
rect 4159 7912 4164 7917
rect 3796 7792 3801 7797
rect 3832 7785 3837 7790
rect 3843 7789 3848 7794
rect 3866 7780 3871 7785
rect 3890 7785 3895 7790
rect 3919 7791 3924 7796
rect 3948 7791 3952 7796
rect 3905 7780 3910 7786
rect 3935 7785 3940 7790
rect 3964 7786 3969 7791
rect 3989 7780 3994 7785
rect 4046 7859 4051 7864
rect 4034 7791 4039 7796
rect 4093 7785 4098 7790
rect 4104 7789 4109 7794
rect 4127 7780 4132 7785
rect 4151 7785 4156 7790
rect 4180 7791 4185 7796
rect 4209 7791 4213 7796
rect 4166 7780 4171 7786
rect 4196 7785 4201 7790
rect 4221 7791 4226 7796
rect 4529 7814 4533 7818
rect 4534 7814 4538 7818
rect 4539 7814 4543 7818
rect 4544 7814 4548 7818
rect 4549 7814 4553 7818
rect 4554 7814 4558 7818
rect 4559 7814 4563 7818
rect 4564 7814 4568 7818
rect 4569 7814 4573 7818
rect 4574 7814 4578 7818
rect 4579 7814 4583 7818
rect 4584 7814 4588 7818
rect 4589 7814 4593 7818
rect 4529 7809 4533 7813
rect 4534 7809 4538 7813
rect 4539 7809 4543 7813
rect 4544 7809 4548 7813
rect 4549 7809 4553 7813
rect 4554 7809 4558 7813
rect 4559 7809 4563 7813
rect 4564 7809 4568 7813
rect 4569 7809 4573 7813
rect 4574 7809 4578 7813
rect 4579 7809 4583 7813
rect 4584 7809 4588 7813
rect 4589 7809 4593 7813
rect 4479 7789 4483 7793
rect 4489 7789 4493 7793
rect 4499 7789 4503 7793
rect 4509 7789 4513 7793
rect 4479 7784 4483 7788
rect 4489 7784 4493 7788
rect 4499 7784 4503 7788
rect 4509 7784 4513 7788
rect 4479 7779 4483 7783
rect 4489 7779 4493 7783
rect 4499 7779 4503 7783
rect 4509 7779 4513 7783
rect 4479 7774 4483 7778
rect 4489 7774 4493 7778
rect 4499 7774 4503 7778
rect 4509 7774 4513 7778
rect 4525 7789 4529 7793
rect 4535 7789 4539 7793
rect 4545 7789 4549 7793
rect 4555 7789 4559 7793
rect 4525 7784 4529 7788
rect 4535 7784 4539 7788
rect 4545 7784 4549 7788
rect 4555 7784 4559 7788
rect 4525 7779 4529 7783
rect 4535 7779 4539 7783
rect 4545 7779 4549 7783
rect 4555 7779 4559 7783
rect 4525 7774 4529 7778
rect 4535 7774 4539 7778
rect 4545 7774 4549 7778
rect 4555 7774 4559 7778
rect 4095 7680 4099 7684
rect 4220 7598 4224 7602
rect 4479 7202 4483 7206
rect 4489 7202 4493 7206
rect 4499 7202 4503 7206
rect 4509 7202 4513 7206
rect 4479 7197 4483 7201
rect 4489 7197 4493 7201
rect 4499 7197 4503 7201
rect 4509 7197 4513 7201
rect 4479 7192 4483 7196
rect 4489 7192 4493 7196
rect 4499 7192 4503 7196
rect 4509 7192 4513 7196
rect 4479 7187 4483 7191
rect 4489 7187 4493 7191
rect 4499 7187 4503 7191
rect 4509 7187 4513 7191
rect 4525 7202 4529 7206
rect 4535 7202 4539 7206
rect 4545 7202 4549 7206
rect 4555 7202 4559 7206
rect 4525 7197 4529 7201
rect 4535 7197 4539 7201
rect 4545 7197 4549 7201
rect 4555 7197 4559 7201
rect 4525 7192 4529 7196
rect 4535 7192 4539 7196
rect 4545 7192 4549 7196
rect 4555 7192 4559 7196
rect 4525 7187 4529 7191
rect 4535 7187 4539 7191
rect 4545 7187 4549 7191
rect 4555 7187 4559 7191
rect 613 7158 617 7162
rect 623 7158 627 7162
rect 633 7158 637 7162
rect 643 7158 647 7162
rect 613 7153 617 7157
rect 623 7153 627 7157
rect 633 7153 637 7157
rect 643 7153 647 7157
rect 613 7148 617 7152
rect 623 7148 627 7152
rect 633 7148 637 7152
rect 643 7148 647 7152
rect 613 7143 617 7147
rect 623 7143 627 7147
rect 633 7143 637 7147
rect 643 7143 647 7147
rect 659 7158 663 7162
rect 669 7158 673 7162
rect 679 7158 683 7162
rect 689 7158 693 7162
rect 659 7153 663 7157
rect 669 7153 673 7157
rect 679 7153 683 7157
rect 689 7153 693 7157
rect 659 7148 663 7152
rect 669 7148 673 7152
rect 679 7148 683 7152
rect 689 7148 693 7152
rect 659 7143 663 7147
rect 669 7143 673 7147
rect 679 7143 683 7147
rect 689 7143 693 7147
rect 4479 6893 4483 6897
rect 4489 6893 4493 6897
rect 4499 6893 4503 6897
rect 4509 6893 4513 6897
rect 4479 6888 4483 6892
rect 4489 6888 4493 6892
rect 4499 6888 4503 6892
rect 4509 6888 4513 6892
rect 4479 6883 4483 6887
rect 4489 6883 4493 6887
rect 4499 6883 4503 6887
rect 4509 6883 4513 6887
rect 4479 6878 4483 6882
rect 4489 6878 4493 6882
rect 4499 6878 4503 6882
rect 4509 6878 4513 6882
rect 4525 6893 4529 6897
rect 4535 6893 4539 6897
rect 4545 6893 4549 6897
rect 4555 6893 4559 6897
rect 4525 6888 4529 6892
rect 4535 6888 4539 6892
rect 4545 6888 4549 6892
rect 4555 6888 4559 6892
rect 4525 6883 4529 6887
rect 4535 6883 4539 6887
rect 4545 6883 4549 6887
rect 4555 6883 4559 6887
rect 4525 6878 4529 6882
rect 4535 6878 4539 6882
rect 4545 6878 4549 6882
rect 4555 6878 4559 6882
rect 613 6849 617 6853
rect 623 6849 627 6853
rect 633 6849 637 6853
rect 643 6849 647 6853
rect 613 6844 617 6848
rect 623 6844 627 6848
rect 633 6844 637 6848
rect 643 6844 647 6848
rect 613 6839 617 6843
rect 623 6839 627 6843
rect 633 6839 637 6843
rect 643 6839 647 6843
rect 613 6834 617 6838
rect 623 6834 627 6838
rect 633 6834 637 6838
rect 643 6834 647 6838
rect 659 6849 663 6853
rect 669 6849 673 6853
rect 679 6849 683 6853
rect 689 6849 693 6853
rect 659 6844 663 6848
rect 669 6844 673 6848
rect 679 6844 683 6848
rect 689 6844 693 6848
rect 659 6839 663 6843
rect 669 6839 673 6843
rect 679 6839 683 6843
rect 689 6839 693 6843
rect 659 6834 663 6838
rect 669 6834 673 6838
rect 679 6834 683 6838
rect 689 6834 693 6838
rect 4479 6584 4483 6588
rect 4489 6584 4493 6588
rect 4499 6584 4503 6588
rect 4509 6584 4513 6588
rect 4479 6579 4483 6583
rect 4489 6579 4493 6583
rect 4499 6579 4503 6583
rect 4509 6579 4513 6583
rect 4479 6574 4483 6578
rect 4489 6574 4493 6578
rect 4499 6574 4503 6578
rect 4509 6574 4513 6578
rect 4479 6569 4483 6573
rect 4489 6569 4493 6573
rect 4499 6569 4503 6573
rect 4509 6569 4513 6573
rect 4525 6584 4529 6588
rect 4535 6584 4539 6588
rect 4545 6584 4549 6588
rect 4555 6584 4559 6588
rect 4525 6579 4529 6583
rect 4535 6579 4539 6583
rect 4545 6579 4549 6583
rect 4555 6579 4559 6583
rect 4525 6574 4529 6578
rect 4535 6574 4539 6578
rect 4545 6574 4549 6578
rect 4555 6574 4559 6578
rect 4525 6569 4529 6573
rect 4535 6569 4539 6573
rect 4545 6569 4549 6573
rect 4555 6569 4559 6573
rect 613 6540 617 6544
rect 623 6540 627 6544
rect 633 6540 637 6544
rect 643 6540 647 6544
rect 613 6535 617 6539
rect 623 6535 627 6539
rect 633 6535 637 6539
rect 643 6535 647 6539
rect 613 6530 617 6534
rect 623 6530 627 6534
rect 633 6530 637 6534
rect 643 6530 647 6534
rect 613 6525 617 6529
rect 623 6525 627 6529
rect 633 6525 637 6529
rect 643 6525 647 6529
rect 659 6540 663 6544
rect 669 6540 673 6544
rect 679 6540 683 6544
rect 689 6540 693 6544
rect 659 6535 663 6539
rect 669 6535 673 6539
rect 679 6535 683 6539
rect 689 6535 693 6539
rect 659 6530 663 6534
rect 669 6530 673 6534
rect 679 6530 683 6534
rect 689 6530 693 6534
rect 659 6525 663 6529
rect 669 6525 673 6529
rect 679 6525 683 6529
rect 689 6525 693 6529
rect 4479 6275 4483 6279
rect 4489 6275 4493 6279
rect 4499 6275 4503 6279
rect 4509 6275 4513 6279
rect 4479 6270 4483 6274
rect 4489 6270 4493 6274
rect 4499 6270 4503 6274
rect 4509 6270 4513 6274
rect 4479 6265 4483 6269
rect 4489 6265 4493 6269
rect 4499 6265 4503 6269
rect 4509 6265 4513 6269
rect 4479 6260 4483 6264
rect 4489 6260 4493 6264
rect 4499 6260 4503 6264
rect 4509 6260 4513 6264
rect 4525 6275 4529 6279
rect 4535 6275 4539 6279
rect 4545 6275 4549 6279
rect 4555 6275 4559 6279
rect 4525 6270 4529 6274
rect 4535 6270 4539 6274
rect 4545 6270 4549 6274
rect 4555 6270 4559 6274
rect 4525 6265 4529 6269
rect 4535 6265 4539 6269
rect 4545 6265 4549 6269
rect 4555 6265 4559 6269
rect 4525 6260 4529 6264
rect 4535 6260 4539 6264
rect 4545 6260 4549 6264
rect 4555 6260 4559 6264
rect 613 6140 617 6144
rect 623 6140 627 6144
rect 633 6140 637 6144
rect 643 6140 647 6144
rect 613 6135 617 6139
rect 623 6135 627 6139
rect 633 6135 637 6139
rect 643 6135 647 6139
rect 613 6130 617 6134
rect 623 6130 627 6134
rect 633 6130 637 6134
rect 643 6130 647 6134
rect 613 6125 617 6129
rect 623 6125 627 6129
rect 633 6125 637 6129
rect 643 6125 647 6129
rect 659 6140 663 6144
rect 669 6140 673 6144
rect 679 6140 683 6144
rect 689 6140 693 6144
rect 659 6135 663 6139
rect 669 6135 673 6139
rect 679 6135 683 6139
rect 689 6135 693 6139
rect 659 6130 663 6134
rect 669 6130 673 6134
rect 679 6130 683 6134
rect 689 6130 693 6134
rect 659 6125 663 6129
rect 669 6125 673 6129
rect 679 6125 683 6129
rect 689 6125 693 6129
rect 613 6111 617 6115
rect 623 6111 627 6115
rect 633 6111 637 6115
rect 643 6111 647 6115
rect 613 6106 617 6110
rect 623 6106 627 6110
rect 633 6106 637 6110
rect 643 6106 647 6110
rect 613 6101 617 6105
rect 623 6101 627 6105
rect 633 6101 637 6105
rect 643 6101 647 6105
rect 613 6096 617 6100
rect 623 6096 627 6100
rect 633 6096 637 6100
rect 643 6096 647 6100
rect 659 6111 663 6115
rect 669 6111 673 6115
rect 679 6111 683 6115
rect 689 6111 693 6115
rect 659 6106 663 6110
rect 669 6106 673 6110
rect 679 6106 683 6110
rect 689 6106 693 6110
rect 659 6101 663 6105
rect 669 6101 673 6105
rect 679 6101 683 6105
rect 689 6101 693 6105
rect 659 6096 663 6100
rect 669 6096 673 6100
rect 679 6096 683 6100
rect 689 6096 693 6100
rect 613 6082 617 6086
rect 623 6082 627 6086
rect 633 6082 637 6086
rect 643 6082 647 6086
rect 613 6077 617 6081
rect 623 6077 627 6081
rect 633 6077 637 6081
rect 643 6077 647 6081
rect 613 6072 617 6076
rect 623 6072 627 6076
rect 633 6072 637 6076
rect 643 6072 647 6076
rect 613 6067 617 6071
rect 623 6067 627 6071
rect 633 6067 637 6071
rect 643 6067 647 6071
rect 659 6082 663 6086
rect 669 6082 673 6086
rect 679 6082 683 6086
rect 689 6082 693 6086
rect 659 6077 663 6081
rect 669 6077 673 6081
rect 679 6077 683 6081
rect 689 6077 693 6081
rect 659 6072 663 6076
rect 669 6072 673 6076
rect 679 6072 683 6076
rect 689 6072 693 6076
rect 659 6067 663 6071
rect 669 6067 673 6071
rect 679 6067 683 6071
rect 689 6067 693 6071
rect 4479 6083 4483 6087
rect 4489 6083 4493 6087
rect 4499 6083 4503 6087
rect 4509 6083 4513 6087
rect 4479 6078 4483 6082
rect 4489 6078 4493 6082
rect 4499 6078 4503 6082
rect 4509 6078 4513 6082
rect 4479 6073 4483 6077
rect 4489 6073 4493 6077
rect 4499 6073 4503 6077
rect 4509 6073 4513 6077
rect 4479 6068 4483 6072
rect 4489 6068 4493 6072
rect 4499 6068 4503 6072
rect 4509 6068 4513 6072
rect 4525 6083 4529 6087
rect 4535 6083 4539 6087
rect 4545 6083 4549 6087
rect 4555 6083 4559 6087
rect 4525 6078 4529 6082
rect 4535 6078 4539 6082
rect 4545 6078 4549 6082
rect 4555 6078 4559 6082
rect 4525 6073 4529 6077
rect 4535 6073 4539 6077
rect 4545 6073 4549 6077
rect 4555 6073 4559 6077
rect 4525 6068 4529 6072
rect 4535 6068 4539 6072
rect 4545 6068 4549 6072
rect 4555 6068 4559 6072
rect 4479 6057 4483 6061
rect 4489 6057 4493 6061
rect 4499 6057 4503 6061
rect 4509 6057 4513 6061
rect 613 6053 617 6057
rect 623 6053 627 6057
rect 633 6053 637 6057
rect 643 6053 647 6057
rect 613 6048 617 6052
rect 623 6048 627 6052
rect 633 6048 637 6052
rect 643 6048 647 6052
rect 613 6043 617 6047
rect 623 6043 627 6047
rect 633 6043 637 6047
rect 643 6043 647 6047
rect 613 6038 617 6042
rect 623 6038 627 6042
rect 633 6038 637 6042
rect 643 6038 647 6042
rect 659 6053 663 6057
rect 669 6053 673 6057
rect 679 6053 683 6057
rect 689 6053 693 6057
rect 659 6048 663 6052
rect 669 6048 673 6052
rect 679 6048 683 6052
rect 689 6048 693 6052
rect 659 6043 663 6047
rect 669 6043 673 6047
rect 679 6043 683 6047
rect 689 6043 693 6047
rect 4479 6052 4483 6056
rect 4489 6052 4493 6056
rect 4499 6052 4503 6056
rect 4509 6052 4513 6056
rect 4479 6047 4483 6051
rect 4489 6047 4493 6051
rect 4499 6047 4503 6051
rect 4509 6047 4513 6051
rect 4479 6042 4483 6046
rect 4489 6042 4493 6046
rect 4499 6042 4503 6046
rect 4509 6042 4513 6046
rect 4525 6057 4529 6061
rect 4535 6057 4539 6061
rect 4545 6057 4549 6061
rect 4555 6057 4559 6061
rect 4525 6052 4529 6056
rect 4535 6052 4539 6056
rect 4545 6052 4549 6056
rect 4555 6052 4559 6056
rect 4525 6047 4529 6051
rect 4535 6047 4539 6051
rect 4545 6047 4549 6051
rect 4555 6047 4559 6051
rect 4525 6042 4529 6046
rect 4535 6042 4539 6046
rect 4545 6042 4549 6046
rect 4555 6042 4559 6046
rect 659 6038 663 6042
rect 669 6038 673 6042
rect 679 6038 683 6042
rect 689 6038 693 6042
rect 4479 6031 4483 6035
rect 4489 6031 4493 6035
rect 4499 6031 4503 6035
rect 4509 6031 4513 6035
rect 613 6024 617 6028
rect 623 6024 627 6028
rect 633 6024 637 6028
rect 643 6024 647 6028
rect 613 6019 617 6023
rect 623 6019 627 6023
rect 633 6019 637 6023
rect 643 6019 647 6023
rect 613 6014 617 6018
rect 623 6014 627 6018
rect 633 6014 637 6018
rect 643 6014 647 6018
rect 613 6009 617 6013
rect 623 6009 627 6013
rect 633 6009 637 6013
rect 643 6009 647 6013
rect 659 6024 663 6028
rect 669 6024 673 6028
rect 679 6024 683 6028
rect 689 6024 693 6028
rect 659 6019 663 6023
rect 669 6019 673 6023
rect 679 6019 683 6023
rect 689 6019 693 6023
rect 659 6014 663 6018
rect 669 6014 673 6018
rect 679 6014 683 6018
rect 689 6014 693 6018
rect 4479 6026 4483 6030
rect 4489 6026 4493 6030
rect 4499 6026 4503 6030
rect 4509 6026 4513 6030
rect 4479 6021 4483 6025
rect 4489 6021 4493 6025
rect 4499 6021 4503 6025
rect 4509 6021 4513 6025
rect 4479 6016 4483 6020
rect 4489 6016 4493 6020
rect 4499 6016 4503 6020
rect 4509 6016 4513 6020
rect 4525 6031 4529 6035
rect 4535 6031 4539 6035
rect 4545 6031 4549 6035
rect 4555 6031 4559 6035
rect 4525 6026 4529 6030
rect 4535 6026 4539 6030
rect 4545 6026 4549 6030
rect 4555 6026 4559 6030
rect 4525 6021 4529 6025
rect 4535 6021 4539 6025
rect 4545 6021 4549 6025
rect 4555 6021 4559 6025
rect 4525 6016 4529 6020
rect 4535 6016 4539 6020
rect 4545 6016 4549 6020
rect 4555 6016 4559 6020
rect 659 6009 663 6013
rect 669 6009 673 6013
rect 679 6009 683 6013
rect 689 6009 693 6013
rect 4479 6005 4483 6009
rect 4489 6005 4493 6009
rect 4499 6005 4503 6009
rect 4509 6005 4513 6009
rect 4479 6000 4483 6004
rect 4489 6000 4493 6004
rect 4499 6000 4503 6004
rect 4509 6000 4513 6004
rect 4479 5995 4483 5999
rect 4489 5995 4493 5999
rect 4499 5995 4503 5999
rect 4509 5995 4513 5999
rect 4479 5990 4483 5994
rect 4489 5990 4493 5994
rect 4499 5990 4503 5994
rect 4509 5990 4513 5994
rect 4525 6005 4529 6009
rect 4535 6005 4539 6009
rect 4545 6005 4549 6009
rect 4555 6005 4559 6009
rect 4525 6000 4529 6004
rect 4535 6000 4539 6004
rect 4545 6000 4549 6004
rect 4555 6000 4559 6004
rect 4525 5995 4529 5999
rect 4535 5995 4539 5999
rect 4545 5995 4549 5999
rect 4555 5995 4559 5999
rect 4525 5990 4529 5994
rect 4535 5990 4539 5994
rect 4545 5990 4549 5994
rect 4555 5990 4559 5994
rect 4479 5979 4483 5983
rect 4489 5979 4493 5983
rect 4499 5979 4503 5983
rect 4509 5979 4513 5983
rect 4479 5974 4483 5978
rect 4489 5974 4493 5978
rect 4499 5974 4503 5978
rect 4509 5974 4513 5978
rect 4479 5969 4483 5973
rect 4489 5969 4493 5973
rect 4499 5969 4503 5973
rect 4509 5969 4513 5973
rect 4479 5964 4483 5968
rect 4489 5964 4493 5968
rect 4499 5964 4503 5968
rect 4509 5964 4513 5968
rect 4525 5979 4529 5983
rect 4535 5979 4539 5983
rect 4545 5979 4549 5983
rect 4555 5979 4559 5983
rect 4525 5974 4529 5978
rect 4535 5974 4539 5978
rect 4545 5974 4549 5978
rect 4555 5974 4559 5978
rect 4525 5969 4529 5973
rect 4535 5969 4539 5973
rect 4545 5969 4549 5973
rect 4555 5969 4559 5973
rect 4525 5964 4529 5968
rect 4535 5964 4539 5968
rect 4545 5964 4549 5968
rect 4555 5964 4559 5968
rect 757 5896 761 5900
rect 762 5896 766 5900
rect 767 5896 771 5900
rect 772 5896 776 5900
rect 757 5886 761 5890
rect 762 5886 766 5890
rect 767 5886 771 5890
rect 772 5886 776 5890
rect 757 5876 761 5880
rect 762 5876 766 5880
rect 767 5876 771 5880
rect 772 5876 776 5880
rect 757 5866 761 5870
rect 762 5866 766 5870
rect 767 5866 771 5870
rect 772 5866 776 5870
rect 783 5896 787 5900
rect 788 5896 792 5900
rect 793 5896 797 5900
rect 798 5896 802 5900
rect 783 5886 787 5890
rect 788 5886 792 5890
rect 793 5886 797 5890
rect 798 5886 802 5890
rect 783 5876 787 5880
rect 788 5876 792 5880
rect 793 5876 797 5880
rect 798 5876 802 5880
rect 783 5866 787 5870
rect 788 5866 792 5870
rect 793 5866 797 5870
rect 798 5866 802 5870
rect 809 5896 813 5900
rect 814 5896 818 5900
rect 819 5896 823 5900
rect 824 5896 828 5900
rect 809 5886 813 5890
rect 814 5886 818 5890
rect 819 5886 823 5890
rect 824 5886 828 5890
rect 809 5876 813 5880
rect 814 5876 818 5880
rect 819 5876 823 5880
rect 824 5876 828 5880
rect 809 5866 813 5870
rect 814 5866 818 5870
rect 819 5866 823 5870
rect 824 5866 828 5870
rect 835 5896 839 5900
rect 840 5896 844 5900
rect 845 5896 849 5900
rect 850 5896 854 5900
rect 835 5886 839 5890
rect 840 5886 844 5890
rect 845 5886 849 5890
rect 850 5886 854 5890
rect 835 5876 839 5880
rect 840 5876 844 5880
rect 845 5876 849 5880
rect 850 5876 854 5880
rect 835 5866 839 5870
rect 840 5866 844 5870
rect 845 5866 849 5870
rect 850 5866 854 5870
rect 861 5896 865 5900
rect 866 5896 870 5900
rect 871 5896 875 5900
rect 876 5896 880 5900
rect 861 5886 865 5890
rect 866 5886 870 5890
rect 871 5886 875 5890
rect 876 5886 880 5890
rect 861 5876 865 5880
rect 866 5876 870 5880
rect 871 5876 875 5880
rect 876 5876 880 5880
rect 861 5866 865 5870
rect 866 5866 870 5870
rect 871 5866 875 5870
rect 876 5866 880 5870
rect 1054 5896 1058 5900
rect 1059 5896 1063 5900
rect 1064 5896 1068 5900
rect 1069 5896 1073 5900
rect 1054 5886 1058 5890
rect 1059 5886 1063 5890
rect 1064 5886 1068 5890
rect 1069 5886 1073 5890
rect 1054 5876 1058 5880
rect 1059 5876 1063 5880
rect 1064 5876 1068 5880
rect 1069 5876 1073 5880
rect 1054 5866 1058 5870
rect 1059 5866 1063 5870
rect 1064 5866 1068 5870
rect 1069 5866 1073 5870
rect 1363 5896 1367 5900
rect 1368 5896 1372 5900
rect 1373 5896 1377 5900
rect 1378 5896 1382 5900
rect 1363 5886 1367 5890
rect 1368 5886 1372 5890
rect 1373 5886 1377 5890
rect 1378 5886 1382 5890
rect 1363 5876 1367 5880
rect 1368 5876 1372 5880
rect 1373 5876 1377 5880
rect 1378 5876 1382 5880
rect 1363 5866 1367 5870
rect 1368 5866 1372 5870
rect 1373 5866 1377 5870
rect 1378 5866 1382 5870
rect 1672 5896 1676 5900
rect 1677 5896 1681 5900
rect 1682 5896 1686 5900
rect 1687 5896 1691 5900
rect 1672 5886 1676 5890
rect 1677 5886 1681 5890
rect 1682 5886 1686 5890
rect 1687 5886 1691 5890
rect 1672 5876 1676 5880
rect 1677 5876 1681 5880
rect 1682 5876 1686 5880
rect 1687 5876 1691 5880
rect 1672 5866 1676 5870
rect 1677 5866 1681 5870
rect 1682 5866 1686 5870
rect 1687 5866 1691 5870
rect 1981 5896 1985 5900
rect 1986 5896 1990 5900
rect 1991 5896 1995 5900
rect 1996 5896 2000 5900
rect 1981 5886 1985 5890
rect 1986 5886 1990 5890
rect 1991 5886 1995 5890
rect 1996 5886 2000 5890
rect 1981 5876 1985 5880
rect 1986 5876 1990 5880
rect 1991 5876 1995 5880
rect 1996 5876 2000 5880
rect 1981 5866 1985 5870
rect 1986 5866 1990 5870
rect 1991 5866 1995 5870
rect 1996 5866 2000 5870
rect 2290 5896 2294 5900
rect 2295 5896 2299 5900
rect 2300 5896 2304 5900
rect 2305 5896 2309 5900
rect 2290 5886 2294 5890
rect 2295 5886 2299 5890
rect 2300 5886 2304 5890
rect 2305 5886 2309 5890
rect 2290 5876 2294 5880
rect 2295 5876 2299 5880
rect 2300 5876 2304 5880
rect 2305 5876 2309 5880
rect 2290 5866 2294 5870
rect 2295 5866 2299 5870
rect 2300 5866 2304 5870
rect 2305 5866 2309 5870
rect 2599 5896 2603 5900
rect 2604 5896 2608 5900
rect 2609 5896 2613 5900
rect 2614 5896 2618 5900
rect 2599 5886 2603 5890
rect 2604 5886 2608 5890
rect 2609 5886 2613 5890
rect 2614 5886 2618 5890
rect 2599 5876 2603 5880
rect 2604 5876 2608 5880
rect 2609 5876 2613 5880
rect 2614 5876 2618 5880
rect 2599 5866 2603 5870
rect 2604 5866 2608 5870
rect 2609 5866 2613 5870
rect 2614 5866 2618 5870
rect 2908 5896 2912 5900
rect 2913 5896 2917 5900
rect 2918 5896 2922 5900
rect 2923 5896 2927 5900
rect 2908 5886 2912 5890
rect 2913 5886 2917 5890
rect 2918 5886 2922 5890
rect 2923 5886 2927 5890
rect 2908 5876 2912 5880
rect 2913 5876 2917 5880
rect 2918 5876 2922 5880
rect 2923 5876 2927 5880
rect 2908 5866 2912 5870
rect 2913 5866 2917 5870
rect 2918 5866 2922 5870
rect 2923 5866 2927 5870
rect 3217 5896 3221 5900
rect 3222 5896 3226 5900
rect 3227 5896 3231 5900
rect 3232 5896 3236 5900
rect 3217 5886 3221 5890
rect 3222 5886 3226 5890
rect 3227 5886 3231 5890
rect 3232 5886 3236 5890
rect 3217 5876 3221 5880
rect 3222 5876 3226 5880
rect 3227 5876 3231 5880
rect 3232 5876 3236 5880
rect 3217 5866 3221 5870
rect 3222 5866 3226 5870
rect 3227 5866 3231 5870
rect 3232 5866 3236 5870
rect 3526 5896 3530 5900
rect 3531 5896 3535 5900
rect 3536 5896 3540 5900
rect 3541 5896 3545 5900
rect 3526 5886 3530 5890
rect 3531 5886 3535 5890
rect 3536 5886 3540 5890
rect 3541 5886 3545 5890
rect 3526 5876 3530 5880
rect 3531 5876 3535 5880
rect 3536 5876 3540 5880
rect 3541 5876 3545 5880
rect 3526 5866 3530 5870
rect 3531 5866 3535 5870
rect 3536 5866 3540 5870
rect 3541 5866 3545 5870
rect 3835 5896 3839 5900
rect 3840 5896 3844 5900
rect 3845 5896 3849 5900
rect 3850 5896 3854 5900
rect 3835 5886 3839 5890
rect 3840 5886 3844 5890
rect 3845 5886 3849 5890
rect 3850 5886 3854 5890
rect 3835 5876 3839 5880
rect 3840 5876 3844 5880
rect 3845 5876 3849 5880
rect 3850 5876 3854 5880
rect 3835 5866 3839 5870
rect 3840 5866 3844 5870
rect 3845 5866 3849 5870
rect 3850 5866 3854 5870
rect 4235 5896 4239 5900
rect 4240 5896 4244 5900
rect 4245 5896 4249 5900
rect 4250 5896 4254 5900
rect 4235 5886 4239 5890
rect 4240 5886 4244 5890
rect 4245 5886 4249 5890
rect 4250 5886 4254 5890
rect 4235 5876 4239 5880
rect 4240 5876 4244 5880
rect 4245 5876 4249 5880
rect 4250 5876 4254 5880
rect 4235 5866 4239 5870
rect 4240 5866 4244 5870
rect 4245 5866 4249 5870
rect 4250 5866 4254 5870
rect 4264 5896 4268 5900
rect 4269 5896 4273 5900
rect 4274 5896 4278 5900
rect 4279 5896 4283 5900
rect 4264 5886 4268 5890
rect 4269 5886 4273 5890
rect 4274 5886 4278 5890
rect 4279 5886 4283 5890
rect 4264 5876 4268 5880
rect 4269 5876 4273 5880
rect 4274 5876 4278 5880
rect 4279 5876 4283 5880
rect 4264 5866 4268 5870
rect 4269 5866 4273 5870
rect 4274 5866 4278 5870
rect 4279 5866 4283 5870
rect 4293 5896 4297 5900
rect 4298 5896 4302 5900
rect 4303 5896 4307 5900
rect 4308 5896 4312 5900
rect 4293 5886 4297 5890
rect 4298 5886 4302 5890
rect 4303 5886 4307 5890
rect 4308 5886 4312 5890
rect 4293 5876 4297 5880
rect 4298 5876 4302 5880
rect 4303 5876 4307 5880
rect 4308 5876 4312 5880
rect 4293 5866 4297 5870
rect 4298 5866 4302 5870
rect 4303 5866 4307 5870
rect 4308 5866 4312 5870
rect 4322 5896 4326 5900
rect 4327 5896 4331 5900
rect 4332 5896 4336 5900
rect 4337 5896 4341 5900
rect 4322 5886 4326 5890
rect 4327 5886 4331 5890
rect 4332 5886 4336 5890
rect 4337 5886 4341 5890
rect 4322 5876 4326 5880
rect 4327 5876 4331 5880
rect 4332 5876 4336 5880
rect 4337 5876 4341 5880
rect 4322 5866 4326 5870
rect 4327 5866 4331 5870
rect 4332 5866 4336 5870
rect 4337 5866 4341 5870
rect 4351 5896 4355 5900
rect 4356 5896 4360 5900
rect 4361 5896 4365 5900
rect 4366 5896 4370 5900
rect 4351 5886 4355 5890
rect 4356 5886 4360 5890
rect 4361 5886 4365 5890
rect 4366 5886 4370 5890
rect 4351 5876 4355 5880
rect 4356 5876 4360 5880
rect 4361 5876 4365 5880
rect 4366 5876 4370 5880
rect 4351 5866 4355 5870
rect 4356 5866 4360 5870
rect 4361 5866 4365 5870
rect 4366 5866 4370 5870
rect 757 5850 761 5854
rect 762 5850 766 5854
rect 767 5850 771 5854
rect 772 5850 776 5854
rect 757 5840 761 5844
rect 762 5840 766 5844
rect 767 5840 771 5844
rect 772 5840 776 5844
rect 757 5830 761 5834
rect 762 5830 766 5834
rect 767 5830 771 5834
rect 772 5830 776 5834
rect 757 5820 761 5824
rect 762 5820 766 5824
rect 767 5820 771 5824
rect 772 5820 776 5824
rect 783 5850 787 5854
rect 788 5850 792 5854
rect 793 5850 797 5854
rect 798 5850 802 5854
rect 783 5840 787 5844
rect 788 5840 792 5844
rect 793 5840 797 5844
rect 798 5840 802 5844
rect 783 5830 787 5834
rect 788 5830 792 5834
rect 793 5830 797 5834
rect 798 5830 802 5834
rect 783 5820 787 5824
rect 788 5820 792 5824
rect 793 5820 797 5824
rect 798 5820 802 5824
rect 809 5850 813 5854
rect 814 5850 818 5854
rect 819 5850 823 5854
rect 824 5850 828 5854
rect 809 5840 813 5844
rect 814 5840 818 5844
rect 819 5840 823 5844
rect 824 5840 828 5844
rect 809 5830 813 5834
rect 814 5830 818 5834
rect 819 5830 823 5834
rect 824 5830 828 5834
rect 809 5820 813 5824
rect 814 5820 818 5824
rect 819 5820 823 5824
rect 824 5820 828 5824
rect 835 5850 839 5854
rect 840 5850 844 5854
rect 845 5850 849 5854
rect 850 5850 854 5854
rect 835 5840 839 5844
rect 840 5840 844 5844
rect 845 5840 849 5844
rect 850 5840 854 5844
rect 835 5830 839 5834
rect 840 5830 844 5834
rect 845 5830 849 5834
rect 850 5830 854 5834
rect 835 5820 839 5824
rect 840 5820 844 5824
rect 845 5820 849 5824
rect 850 5820 854 5824
rect 861 5850 865 5854
rect 866 5850 870 5854
rect 871 5850 875 5854
rect 876 5850 880 5854
rect 861 5840 865 5844
rect 866 5840 870 5844
rect 871 5840 875 5844
rect 876 5840 880 5844
rect 861 5830 865 5834
rect 866 5830 870 5834
rect 871 5830 875 5834
rect 876 5830 880 5834
rect 861 5820 865 5824
rect 866 5820 870 5824
rect 871 5820 875 5824
rect 876 5820 880 5824
rect 1054 5850 1058 5854
rect 1059 5850 1063 5854
rect 1064 5850 1068 5854
rect 1069 5850 1073 5854
rect 1054 5840 1058 5844
rect 1059 5840 1063 5844
rect 1064 5840 1068 5844
rect 1069 5840 1073 5844
rect 1054 5830 1058 5834
rect 1059 5830 1063 5834
rect 1064 5830 1068 5834
rect 1069 5830 1073 5834
rect 1054 5820 1058 5824
rect 1059 5820 1063 5824
rect 1064 5820 1068 5824
rect 1069 5820 1073 5824
rect 1363 5850 1367 5854
rect 1368 5850 1372 5854
rect 1373 5850 1377 5854
rect 1378 5850 1382 5854
rect 1363 5840 1367 5844
rect 1368 5840 1372 5844
rect 1373 5840 1377 5844
rect 1378 5840 1382 5844
rect 1363 5830 1367 5834
rect 1368 5830 1372 5834
rect 1373 5830 1377 5834
rect 1378 5830 1382 5834
rect 1363 5820 1367 5824
rect 1368 5820 1372 5824
rect 1373 5820 1377 5824
rect 1378 5820 1382 5824
rect 1672 5850 1676 5854
rect 1677 5850 1681 5854
rect 1682 5850 1686 5854
rect 1687 5850 1691 5854
rect 1672 5840 1676 5844
rect 1677 5840 1681 5844
rect 1682 5840 1686 5844
rect 1687 5840 1691 5844
rect 1672 5830 1676 5834
rect 1677 5830 1681 5834
rect 1682 5830 1686 5834
rect 1687 5830 1691 5834
rect 1672 5820 1676 5824
rect 1677 5820 1681 5824
rect 1682 5820 1686 5824
rect 1687 5820 1691 5824
rect 1981 5850 1985 5854
rect 1986 5850 1990 5854
rect 1991 5850 1995 5854
rect 1996 5850 2000 5854
rect 1981 5840 1985 5844
rect 1986 5840 1990 5844
rect 1991 5840 1995 5844
rect 1996 5840 2000 5844
rect 1981 5830 1985 5834
rect 1986 5830 1990 5834
rect 1991 5830 1995 5834
rect 1996 5830 2000 5834
rect 1981 5820 1985 5824
rect 1986 5820 1990 5824
rect 1991 5820 1995 5824
rect 1996 5820 2000 5824
rect 2290 5850 2294 5854
rect 2295 5850 2299 5854
rect 2300 5850 2304 5854
rect 2305 5850 2309 5854
rect 2290 5840 2294 5844
rect 2295 5840 2299 5844
rect 2300 5840 2304 5844
rect 2305 5840 2309 5844
rect 2290 5830 2294 5834
rect 2295 5830 2299 5834
rect 2300 5830 2304 5834
rect 2305 5830 2309 5834
rect 2290 5820 2294 5824
rect 2295 5820 2299 5824
rect 2300 5820 2304 5824
rect 2305 5820 2309 5824
rect 2599 5850 2603 5854
rect 2604 5850 2608 5854
rect 2609 5850 2613 5854
rect 2614 5850 2618 5854
rect 2599 5840 2603 5844
rect 2604 5840 2608 5844
rect 2609 5840 2613 5844
rect 2614 5840 2618 5844
rect 2599 5830 2603 5834
rect 2604 5830 2608 5834
rect 2609 5830 2613 5834
rect 2614 5830 2618 5834
rect 2599 5820 2603 5824
rect 2604 5820 2608 5824
rect 2609 5820 2613 5824
rect 2614 5820 2618 5824
rect 2908 5850 2912 5854
rect 2913 5850 2917 5854
rect 2918 5850 2922 5854
rect 2923 5850 2927 5854
rect 2908 5840 2912 5844
rect 2913 5840 2917 5844
rect 2918 5840 2922 5844
rect 2923 5840 2927 5844
rect 2908 5830 2912 5834
rect 2913 5830 2917 5834
rect 2918 5830 2922 5834
rect 2923 5830 2927 5834
rect 2908 5820 2912 5824
rect 2913 5820 2917 5824
rect 2918 5820 2922 5824
rect 2923 5820 2927 5824
rect 3217 5850 3221 5854
rect 3222 5850 3226 5854
rect 3227 5850 3231 5854
rect 3232 5850 3236 5854
rect 3217 5840 3221 5844
rect 3222 5840 3226 5844
rect 3227 5840 3231 5844
rect 3232 5840 3236 5844
rect 3217 5830 3221 5834
rect 3222 5830 3226 5834
rect 3227 5830 3231 5834
rect 3232 5830 3236 5834
rect 3217 5820 3221 5824
rect 3222 5820 3226 5824
rect 3227 5820 3231 5824
rect 3232 5820 3236 5824
rect 3526 5850 3530 5854
rect 3531 5850 3535 5854
rect 3536 5850 3540 5854
rect 3541 5850 3545 5854
rect 3526 5840 3530 5844
rect 3531 5840 3535 5844
rect 3536 5840 3540 5844
rect 3541 5840 3545 5844
rect 3526 5830 3530 5834
rect 3531 5830 3535 5834
rect 3536 5830 3540 5834
rect 3541 5830 3545 5834
rect 3526 5820 3530 5824
rect 3531 5820 3535 5824
rect 3536 5820 3540 5824
rect 3541 5820 3545 5824
rect 3835 5850 3839 5854
rect 3840 5850 3844 5854
rect 3845 5850 3849 5854
rect 3850 5850 3854 5854
rect 3835 5840 3839 5844
rect 3840 5840 3844 5844
rect 3845 5840 3849 5844
rect 3850 5840 3854 5844
rect 3835 5830 3839 5834
rect 3840 5830 3844 5834
rect 3845 5830 3849 5834
rect 3850 5830 3854 5834
rect 3835 5820 3839 5824
rect 3840 5820 3844 5824
rect 3845 5820 3849 5824
rect 3850 5820 3854 5824
rect 4235 5850 4239 5854
rect 4240 5850 4244 5854
rect 4245 5850 4249 5854
rect 4250 5850 4254 5854
rect 4235 5840 4239 5844
rect 4240 5840 4244 5844
rect 4245 5840 4249 5844
rect 4250 5840 4254 5844
rect 4235 5830 4239 5834
rect 4240 5830 4244 5834
rect 4245 5830 4249 5834
rect 4250 5830 4254 5834
rect 4235 5820 4239 5824
rect 4240 5820 4244 5824
rect 4245 5820 4249 5824
rect 4250 5820 4254 5824
rect 4264 5850 4268 5854
rect 4269 5850 4273 5854
rect 4274 5850 4278 5854
rect 4279 5850 4283 5854
rect 4264 5840 4268 5844
rect 4269 5840 4273 5844
rect 4274 5840 4278 5844
rect 4279 5840 4283 5844
rect 4264 5830 4268 5834
rect 4269 5830 4273 5834
rect 4274 5830 4278 5834
rect 4279 5830 4283 5834
rect 4264 5820 4268 5824
rect 4269 5820 4273 5824
rect 4274 5820 4278 5824
rect 4279 5820 4283 5824
rect 4293 5850 4297 5854
rect 4298 5850 4302 5854
rect 4303 5850 4307 5854
rect 4308 5850 4312 5854
rect 4293 5840 4297 5844
rect 4298 5840 4302 5844
rect 4303 5840 4307 5844
rect 4308 5840 4312 5844
rect 4293 5830 4297 5834
rect 4298 5830 4302 5834
rect 4303 5830 4307 5834
rect 4308 5830 4312 5834
rect 4293 5820 4297 5824
rect 4298 5820 4302 5824
rect 4303 5820 4307 5824
rect 4308 5820 4312 5824
rect 4322 5850 4326 5854
rect 4327 5850 4331 5854
rect 4332 5850 4336 5854
rect 4337 5850 4341 5854
rect 4322 5840 4326 5844
rect 4327 5840 4331 5844
rect 4332 5840 4336 5844
rect 4337 5840 4341 5844
rect 4322 5830 4326 5834
rect 4327 5830 4331 5834
rect 4332 5830 4336 5834
rect 4337 5830 4341 5834
rect 4322 5820 4326 5824
rect 4327 5820 4331 5824
rect 4332 5820 4336 5824
rect 4337 5820 4341 5824
rect 4351 5850 4355 5854
rect 4356 5850 4360 5854
rect 4361 5850 4365 5854
rect 4366 5850 4370 5854
rect 4351 5840 4355 5844
rect 4356 5840 4360 5844
rect 4361 5840 4365 5844
rect 4366 5840 4370 5844
rect 4351 5830 4355 5834
rect 4356 5830 4360 5834
rect 4361 5830 4365 5834
rect 4366 5830 4370 5834
rect 4351 5820 4355 5824
rect 4356 5820 4360 5824
rect 4361 5820 4365 5824
rect 4366 5820 4370 5824
<< metal3 >>
rect 570 9800 4602 9809
rect 570 9796 1354 9800
rect 1358 9796 1359 9800
rect 1363 9796 1663 9800
rect 1667 9796 1668 9800
rect 1672 9796 1972 9800
rect 1976 9796 1977 9800
rect 1981 9796 2281 9800
rect 2285 9796 2286 9800
rect 2290 9796 2590 9800
rect 2594 9796 2595 9800
rect 2599 9796 2899 9800
rect 2903 9796 2904 9800
rect 2908 9796 3208 9800
rect 3212 9796 3213 9800
rect 3217 9796 3517 9800
rect 3521 9796 3522 9800
rect 3526 9796 3826 9800
rect 3830 9796 3831 9800
rect 3835 9796 4602 9800
rect 570 9795 4602 9796
rect 570 9791 1354 9795
rect 1358 9791 1359 9795
rect 1363 9791 1663 9795
rect 1667 9791 1668 9795
rect 1672 9791 1972 9795
rect 1976 9791 1977 9795
rect 1981 9791 2281 9795
rect 2285 9791 2286 9795
rect 2290 9791 2590 9795
rect 2594 9791 2595 9795
rect 2599 9791 2899 9795
rect 2903 9791 2904 9795
rect 2908 9791 3208 9795
rect 3212 9791 3213 9795
rect 3217 9791 3517 9795
rect 3521 9791 3522 9795
rect 3526 9791 3652 9795
rect 3656 9791 3657 9795
rect 3661 9791 3826 9795
rect 3830 9791 3831 9795
rect 3835 9791 4602 9795
rect 570 9790 4602 9791
rect 570 9786 1354 9790
rect 1358 9786 1359 9790
rect 1363 9786 1663 9790
rect 1667 9786 1668 9790
rect 1672 9786 1972 9790
rect 1976 9786 1977 9790
rect 1981 9786 2281 9790
rect 2285 9786 2286 9790
rect 2290 9786 2590 9790
rect 2594 9786 2595 9790
rect 2599 9786 2899 9790
rect 2903 9786 2904 9790
rect 2908 9786 3208 9790
rect 3212 9786 3213 9790
rect 3217 9786 3517 9790
rect 3521 9786 3522 9790
rect 3526 9786 3652 9790
rect 3656 9786 3657 9790
rect 3661 9786 3826 9790
rect 3830 9786 3831 9790
rect 3835 9786 4602 9790
rect 570 9785 4602 9786
rect 570 9781 1354 9785
rect 1358 9781 1359 9785
rect 1363 9781 1663 9785
rect 1667 9781 1668 9785
rect 1672 9781 1972 9785
rect 1976 9781 1977 9785
rect 1981 9781 2281 9785
rect 2285 9781 2286 9785
rect 2290 9781 2590 9785
rect 2594 9781 2595 9785
rect 2599 9781 2899 9785
rect 2903 9781 2904 9785
rect 2908 9781 3208 9785
rect 3212 9781 3213 9785
rect 3217 9781 3517 9785
rect 3521 9781 3522 9785
rect 3526 9781 3652 9785
rect 3656 9781 3657 9785
rect 3661 9781 3826 9785
rect 3830 9781 3831 9785
rect 3835 9781 4602 9785
rect 570 9780 4602 9781
rect 570 9776 1354 9780
rect 1358 9776 1359 9780
rect 1363 9776 1663 9780
rect 1667 9776 1668 9780
rect 1672 9776 1972 9780
rect 1976 9776 1977 9780
rect 1981 9776 2281 9780
rect 2285 9776 2286 9780
rect 2290 9776 2590 9780
rect 2594 9776 2595 9780
rect 2599 9776 2899 9780
rect 2903 9776 2904 9780
rect 2908 9776 3208 9780
rect 3212 9776 3213 9780
rect 3217 9776 3517 9780
rect 3521 9776 3522 9780
rect 3526 9776 3652 9780
rect 3656 9776 3657 9780
rect 3661 9776 3826 9780
rect 3830 9776 3831 9780
rect 3835 9776 4602 9780
rect 570 9775 4602 9776
rect 570 9771 1354 9775
rect 1358 9771 1359 9775
rect 1363 9771 1663 9775
rect 1667 9771 1668 9775
rect 1672 9771 1972 9775
rect 1976 9771 1977 9775
rect 1981 9771 2281 9775
rect 2285 9771 2286 9775
rect 2290 9771 2590 9775
rect 2594 9771 2595 9775
rect 2599 9771 2899 9775
rect 2903 9771 2904 9775
rect 2908 9771 3208 9775
rect 3212 9771 3213 9775
rect 3217 9771 3517 9775
rect 3521 9771 3522 9775
rect 3526 9771 3652 9775
rect 3656 9771 3657 9775
rect 3661 9771 3826 9775
rect 3830 9771 3831 9775
rect 3835 9771 4602 9775
rect 570 9770 4602 9771
rect 570 9766 1354 9770
rect 1358 9766 1359 9770
rect 1363 9769 1663 9770
rect 1363 9766 1547 9769
rect 570 9762 802 9766
rect 806 9762 807 9766
rect 811 9762 812 9766
rect 816 9762 817 9766
rect 821 9762 831 9766
rect 835 9762 836 9766
rect 840 9762 841 9766
rect 845 9762 846 9766
rect 850 9762 860 9766
rect 864 9762 865 9766
rect 869 9762 870 9766
rect 874 9762 875 9766
rect 879 9762 889 9766
rect 893 9762 894 9766
rect 898 9762 899 9766
rect 903 9762 904 9766
rect 908 9762 918 9766
rect 922 9762 923 9766
rect 927 9762 928 9766
rect 932 9762 933 9766
rect 937 9762 1319 9766
rect 1323 9762 1324 9766
rect 1328 9762 1329 9766
rect 1333 9762 1334 9766
rect 1338 9765 1547 9766
rect 1551 9765 1552 9769
rect 1556 9765 1557 9769
rect 1561 9765 1562 9769
rect 1566 9765 1567 9769
rect 1571 9765 1572 9769
rect 1576 9765 1577 9769
rect 1581 9765 1582 9769
rect 1586 9765 1587 9769
rect 1591 9765 1592 9769
rect 1596 9765 1597 9769
rect 1601 9765 1602 9769
rect 1606 9765 1607 9769
rect 1611 9766 1663 9769
rect 1667 9766 1668 9770
rect 1672 9769 1972 9770
rect 1672 9766 1856 9769
rect 1611 9765 1628 9766
rect 1338 9762 1354 9765
rect 570 9761 1354 9762
rect 1358 9761 1359 9765
rect 1363 9764 1628 9765
rect 1363 9761 1547 9764
rect 570 9760 1547 9761
rect 1551 9760 1552 9764
rect 1556 9760 1557 9764
rect 1561 9760 1562 9764
rect 1566 9760 1567 9764
rect 1571 9760 1572 9764
rect 1576 9760 1577 9764
rect 1581 9760 1582 9764
rect 1586 9760 1587 9764
rect 1591 9760 1592 9764
rect 1596 9760 1597 9764
rect 1601 9760 1602 9764
rect 1606 9760 1607 9764
rect 1611 9762 1628 9764
rect 1632 9762 1633 9766
rect 1637 9762 1638 9766
rect 1642 9762 1643 9766
rect 1647 9765 1856 9766
rect 1860 9765 1861 9769
rect 1865 9765 1866 9769
rect 1870 9765 1871 9769
rect 1875 9765 1876 9769
rect 1880 9765 1881 9769
rect 1885 9765 1886 9769
rect 1890 9765 1891 9769
rect 1895 9765 1896 9769
rect 1900 9765 1901 9769
rect 1905 9765 1906 9769
rect 1910 9765 1911 9769
rect 1915 9765 1916 9769
rect 1920 9766 1972 9769
rect 1976 9766 1977 9770
rect 1981 9769 2281 9770
rect 1981 9766 2165 9769
rect 1920 9765 1937 9766
rect 1647 9762 1663 9765
rect 1611 9761 1663 9762
rect 1667 9761 1668 9765
rect 1672 9764 1937 9765
rect 1672 9761 1856 9764
rect 1611 9760 1856 9761
rect 1860 9760 1861 9764
rect 1865 9760 1866 9764
rect 1870 9760 1871 9764
rect 1875 9760 1876 9764
rect 1880 9760 1881 9764
rect 1885 9760 1886 9764
rect 1890 9760 1891 9764
rect 1895 9760 1896 9764
rect 1900 9760 1901 9764
rect 1905 9760 1906 9764
rect 1910 9760 1911 9764
rect 1915 9760 1916 9764
rect 1920 9762 1937 9764
rect 1941 9762 1942 9766
rect 1946 9762 1947 9766
rect 1951 9762 1952 9766
rect 1956 9765 2165 9766
rect 2169 9765 2170 9769
rect 2174 9765 2175 9769
rect 2179 9765 2180 9769
rect 2184 9765 2185 9769
rect 2189 9765 2190 9769
rect 2194 9765 2195 9769
rect 2199 9765 2200 9769
rect 2204 9765 2205 9769
rect 2209 9765 2210 9769
rect 2214 9765 2215 9769
rect 2219 9765 2220 9769
rect 2224 9765 2225 9769
rect 2229 9766 2281 9769
rect 2285 9766 2286 9770
rect 2290 9769 2590 9770
rect 2290 9766 2474 9769
rect 2229 9765 2246 9766
rect 1956 9762 1972 9765
rect 1920 9761 1972 9762
rect 1976 9761 1977 9765
rect 1981 9764 2246 9765
rect 1981 9761 2165 9764
rect 1920 9760 2165 9761
rect 2169 9760 2170 9764
rect 2174 9760 2175 9764
rect 2179 9760 2180 9764
rect 2184 9760 2185 9764
rect 2189 9760 2190 9764
rect 2194 9760 2195 9764
rect 2199 9760 2200 9764
rect 2204 9760 2205 9764
rect 2209 9760 2210 9764
rect 2214 9760 2215 9764
rect 2219 9760 2220 9764
rect 2224 9760 2225 9764
rect 2229 9762 2246 9764
rect 2250 9762 2251 9766
rect 2255 9762 2256 9766
rect 2260 9762 2261 9766
rect 2265 9765 2474 9766
rect 2478 9765 2479 9769
rect 2483 9765 2484 9769
rect 2488 9765 2489 9769
rect 2493 9765 2494 9769
rect 2498 9765 2499 9769
rect 2503 9765 2504 9769
rect 2508 9765 2509 9769
rect 2513 9765 2514 9769
rect 2518 9765 2519 9769
rect 2523 9765 2524 9769
rect 2528 9765 2529 9769
rect 2533 9765 2534 9769
rect 2538 9766 2590 9769
rect 2594 9766 2595 9770
rect 2599 9769 2899 9770
rect 2599 9766 2783 9769
rect 2538 9765 2555 9766
rect 2265 9762 2281 9765
rect 2229 9761 2281 9762
rect 2285 9761 2286 9765
rect 2290 9764 2555 9765
rect 2290 9761 2474 9764
rect 2229 9760 2474 9761
rect 2478 9760 2479 9764
rect 2483 9760 2484 9764
rect 2488 9760 2489 9764
rect 2493 9760 2494 9764
rect 2498 9760 2499 9764
rect 2503 9760 2504 9764
rect 2508 9760 2509 9764
rect 2513 9760 2514 9764
rect 2518 9760 2519 9764
rect 2523 9760 2524 9764
rect 2528 9760 2529 9764
rect 2533 9760 2534 9764
rect 2538 9762 2555 9764
rect 2559 9762 2560 9766
rect 2564 9762 2565 9766
rect 2569 9762 2570 9766
rect 2574 9765 2783 9766
rect 2787 9765 2788 9769
rect 2792 9765 2793 9769
rect 2797 9765 2798 9769
rect 2802 9765 2803 9769
rect 2807 9765 2808 9769
rect 2812 9765 2813 9769
rect 2817 9765 2818 9769
rect 2822 9765 2823 9769
rect 2827 9765 2828 9769
rect 2832 9765 2833 9769
rect 2837 9765 2838 9769
rect 2842 9765 2843 9769
rect 2847 9766 2899 9769
rect 2903 9766 2904 9770
rect 2908 9769 3208 9770
rect 2908 9766 3092 9769
rect 2847 9765 2864 9766
rect 2574 9762 2590 9765
rect 2538 9761 2590 9762
rect 2594 9761 2595 9765
rect 2599 9764 2864 9765
rect 2599 9761 2783 9764
rect 2538 9760 2783 9761
rect 2787 9760 2788 9764
rect 2792 9760 2793 9764
rect 2797 9760 2798 9764
rect 2802 9760 2803 9764
rect 2807 9760 2808 9764
rect 2812 9760 2813 9764
rect 2817 9760 2818 9764
rect 2822 9760 2823 9764
rect 2827 9760 2828 9764
rect 2832 9760 2833 9764
rect 2837 9760 2838 9764
rect 2842 9760 2843 9764
rect 2847 9762 2864 9764
rect 2868 9762 2869 9766
rect 2873 9762 2874 9766
rect 2878 9762 2879 9766
rect 2883 9765 3092 9766
rect 3096 9765 3097 9769
rect 3101 9765 3102 9769
rect 3106 9765 3107 9769
rect 3111 9765 3112 9769
rect 3116 9765 3117 9769
rect 3121 9765 3122 9769
rect 3126 9765 3127 9769
rect 3131 9765 3132 9769
rect 3136 9765 3137 9769
rect 3141 9765 3142 9769
rect 3146 9765 3147 9769
rect 3151 9765 3152 9769
rect 3156 9766 3208 9769
rect 3212 9766 3213 9770
rect 3217 9769 3517 9770
rect 3217 9766 3401 9769
rect 3156 9765 3173 9766
rect 2883 9762 2899 9765
rect 2847 9761 2899 9762
rect 2903 9761 2904 9765
rect 2908 9764 3173 9765
rect 2908 9761 3092 9764
rect 2847 9760 3092 9761
rect 3096 9760 3097 9764
rect 3101 9760 3102 9764
rect 3106 9760 3107 9764
rect 3111 9760 3112 9764
rect 3116 9760 3117 9764
rect 3121 9760 3122 9764
rect 3126 9760 3127 9764
rect 3131 9760 3132 9764
rect 3136 9760 3137 9764
rect 3141 9760 3142 9764
rect 3146 9760 3147 9764
rect 3151 9760 3152 9764
rect 3156 9762 3173 9764
rect 3177 9762 3178 9766
rect 3182 9762 3183 9766
rect 3187 9762 3188 9766
rect 3192 9765 3401 9766
rect 3405 9765 3406 9769
rect 3410 9765 3411 9769
rect 3415 9765 3416 9769
rect 3420 9765 3421 9769
rect 3425 9765 3426 9769
rect 3430 9765 3431 9769
rect 3435 9765 3436 9769
rect 3440 9765 3441 9769
rect 3445 9765 3446 9769
rect 3450 9765 3451 9769
rect 3455 9765 3456 9769
rect 3460 9765 3461 9769
rect 3465 9766 3517 9769
rect 3521 9766 3522 9770
rect 3526 9766 3652 9770
rect 3656 9766 3657 9770
rect 3661 9769 3826 9770
rect 3661 9766 3710 9769
rect 3465 9765 3482 9766
rect 3192 9762 3208 9765
rect 3156 9761 3208 9762
rect 3212 9761 3213 9765
rect 3217 9764 3482 9765
rect 3217 9761 3401 9764
rect 3156 9760 3401 9761
rect 3405 9760 3406 9764
rect 3410 9760 3411 9764
rect 3415 9760 3416 9764
rect 3420 9760 3421 9764
rect 3425 9760 3426 9764
rect 3430 9760 3431 9764
rect 3435 9760 3436 9764
rect 3440 9760 3441 9764
rect 3445 9760 3446 9764
rect 3450 9760 3451 9764
rect 3455 9760 3456 9764
rect 3460 9760 3461 9764
rect 3465 9762 3482 9764
rect 3486 9762 3487 9766
rect 3491 9762 3492 9766
rect 3496 9762 3497 9766
rect 3501 9765 3710 9766
rect 3714 9765 3715 9769
rect 3719 9765 3720 9769
rect 3724 9765 3725 9769
rect 3729 9765 3730 9769
rect 3734 9765 3735 9769
rect 3739 9765 3740 9769
rect 3744 9765 3745 9769
rect 3749 9765 3750 9769
rect 3754 9765 3755 9769
rect 3759 9765 3760 9769
rect 3764 9765 3765 9769
rect 3769 9765 3770 9769
rect 3774 9766 3826 9769
rect 3830 9766 3831 9770
rect 3835 9769 4602 9770
rect 3835 9766 4019 9769
rect 3774 9765 3791 9766
rect 3501 9762 3517 9765
rect 3465 9761 3517 9762
rect 3521 9761 3522 9765
rect 3526 9761 3652 9765
rect 3656 9761 3657 9765
rect 3661 9764 3791 9765
rect 3661 9761 3710 9764
rect 3465 9760 3710 9761
rect 3714 9760 3715 9764
rect 3719 9760 3720 9764
rect 3724 9760 3725 9764
rect 3729 9760 3730 9764
rect 3734 9760 3735 9764
rect 3739 9760 3740 9764
rect 3744 9760 3745 9764
rect 3749 9760 3750 9764
rect 3754 9760 3755 9764
rect 3759 9760 3760 9764
rect 3764 9760 3765 9764
rect 3769 9760 3770 9764
rect 3774 9762 3791 9764
rect 3795 9762 3796 9766
rect 3800 9762 3801 9766
rect 3805 9762 3806 9766
rect 3810 9765 4019 9766
rect 4023 9765 4024 9769
rect 4028 9765 4029 9769
rect 4033 9765 4034 9769
rect 4038 9765 4039 9769
rect 4043 9765 4044 9769
rect 4048 9765 4049 9769
rect 4053 9765 4054 9769
rect 4058 9765 4059 9769
rect 4063 9765 4064 9769
rect 4068 9765 4069 9769
rect 4073 9765 4074 9769
rect 4078 9765 4079 9769
rect 4083 9766 4602 9769
rect 4083 9765 4100 9766
rect 3810 9762 3826 9765
rect 3774 9761 3826 9762
rect 3830 9761 3831 9765
rect 3835 9764 4100 9765
rect 3835 9761 4019 9764
rect 3774 9760 4019 9761
rect 4023 9760 4024 9764
rect 4028 9760 4029 9764
rect 4033 9760 4034 9764
rect 4038 9760 4039 9764
rect 4043 9760 4044 9764
rect 4048 9760 4049 9764
rect 4053 9760 4054 9764
rect 4058 9760 4059 9764
rect 4063 9760 4064 9764
rect 4068 9760 4069 9764
rect 4073 9760 4074 9764
rect 4078 9760 4079 9764
rect 4083 9762 4100 9764
rect 4104 9762 4105 9766
rect 4109 9762 4110 9766
rect 4114 9762 4115 9766
rect 4119 9762 4292 9766
rect 4296 9762 4297 9766
rect 4301 9762 4302 9766
rect 4306 9762 4307 9766
rect 4311 9762 4318 9766
rect 4322 9762 4323 9766
rect 4327 9762 4328 9766
rect 4332 9762 4333 9766
rect 4337 9762 4344 9766
rect 4348 9762 4349 9766
rect 4353 9762 4354 9766
rect 4358 9762 4359 9766
rect 4363 9762 4370 9766
rect 4374 9762 4375 9766
rect 4379 9762 4380 9766
rect 4384 9762 4385 9766
rect 4389 9762 4396 9766
rect 4400 9762 4401 9766
rect 4405 9762 4406 9766
rect 4410 9762 4411 9766
rect 4415 9762 4602 9766
rect 4083 9760 4602 9762
rect 570 9756 1354 9760
rect 1358 9756 1359 9760
rect 1363 9756 1663 9760
rect 1667 9756 1668 9760
rect 1672 9756 1972 9760
rect 1976 9756 1977 9760
rect 1981 9756 2281 9760
rect 2285 9756 2286 9760
rect 2290 9756 2590 9760
rect 2594 9756 2595 9760
rect 2599 9756 2899 9760
rect 2903 9756 2904 9760
rect 2908 9756 3208 9760
rect 3212 9756 3213 9760
rect 3217 9756 3517 9760
rect 3521 9756 3522 9760
rect 3526 9756 3652 9760
rect 3656 9756 3657 9760
rect 3661 9756 3826 9760
rect 3830 9756 3831 9760
rect 3835 9756 4602 9760
rect 570 9752 802 9756
rect 806 9752 807 9756
rect 811 9752 812 9756
rect 816 9752 817 9756
rect 821 9752 831 9756
rect 835 9752 836 9756
rect 840 9752 841 9756
rect 845 9752 846 9756
rect 850 9752 860 9756
rect 864 9752 865 9756
rect 869 9752 870 9756
rect 874 9752 875 9756
rect 879 9752 889 9756
rect 893 9752 894 9756
rect 898 9752 899 9756
rect 903 9752 904 9756
rect 908 9752 918 9756
rect 922 9752 923 9756
rect 927 9752 928 9756
rect 932 9752 933 9756
rect 937 9752 1319 9756
rect 1323 9752 1324 9756
rect 1328 9752 1329 9756
rect 1333 9752 1334 9756
rect 1338 9755 1628 9756
rect 1338 9752 1354 9755
rect 570 9751 1354 9752
rect 1358 9751 1359 9755
rect 1363 9752 1628 9755
rect 1632 9752 1633 9756
rect 1637 9752 1638 9756
rect 1642 9752 1643 9756
rect 1647 9755 1937 9756
rect 1647 9752 1663 9755
rect 1363 9751 1663 9752
rect 1667 9751 1668 9755
rect 1672 9752 1937 9755
rect 1941 9752 1942 9756
rect 1946 9752 1947 9756
rect 1951 9752 1952 9756
rect 1956 9755 2246 9756
rect 1956 9752 1972 9755
rect 1672 9751 1972 9752
rect 1976 9751 1977 9755
rect 1981 9752 2246 9755
rect 2250 9752 2251 9756
rect 2255 9752 2256 9756
rect 2260 9752 2261 9756
rect 2265 9755 2555 9756
rect 2265 9752 2281 9755
rect 1981 9751 2281 9752
rect 2285 9751 2286 9755
rect 2290 9752 2555 9755
rect 2559 9752 2560 9756
rect 2564 9752 2565 9756
rect 2569 9752 2570 9756
rect 2574 9755 2864 9756
rect 2574 9752 2590 9755
rect 2290 9751 2590 9752
rect 2594 9751 2595 9755
rect 2599 9752 2864 9755
rect 2868 9752 2869 9756
rect 2873 9752 2874 9756
rect 2878 9752 2879 9756
rect 2883 9755 3173 9756
rect 2883 9752 2899 9755
rect 2599 9751 2899 9752
rect 2903 9751 2904 9755
rect 2908 9752 3173 9755
rect 3177 9752 3178 9756
rect 3182 9752 3183 9756
rect 3187 9752 3188 9756
rect 3192 9755 3482 9756
rect 3192 9752 3208 9755
rect 2908 9751 3208 9752
rect 3212 9751 3213 9755
rect 3217 9752 3482 9755
rect 3486 9752 3487 9756
rect 3491 9752 3492 9756
rect 3496 9752 3497 9756
rect 3501 9755 3791 9756
rect 3501 9752 3517 9755
rect 3217 9751 3517 9752
rect 3521 9751 3522 9755
rect 3526 9751 3652 9755
rect 3656 9751 3657 9755
rect 3661 9752 3791 9755
rect 3795 9752 3796 9756
rect 3800 9752 3801 9756
rect 3805 9752 3806 9756
rect 3810 9755 4100 9756
rect 3810 9752 3826 9755
rect 3661 9751 3826 9752
rect 3830 9751 3831 9755
rect 3835 9752 4100 9755
rect 4104 9752 4105 9756
rect 4109 9752 4110 9756
rect 4114 9752 4115 9756
rect 4119 9752 4292 9756
rect 4296 9752 4297 9756
rect 4301 9752 4302 9756
rect 4306 9752 4307 9756
rect 4311 9752 4318 9756
rect 4322 9752 4323 9756
rect 4327 9752 4328 9756
rect 4332 9752 4333 9756
rect 4337 9752 4344 9756
rect 4348 9752 4349 9756
rect 4353 9752 4354 9756
rect 4358 9752 4359 9756
rect 4363 9752 4370 9756
rect 4374 9752 4375 9756
rect 4379 9752 4380 9756
rect 4384 9752 4385 9756
rect 4389 9752 4396 9756
rect 4400 9752 4401 9756
rect 4405 9752 4406 9756
rect 4410 9752 4411 9756
rect 4415 9752 4602 9756
rect 3835 9751 4602 9752
rect 570 9750 4602 9751
rect 570 9746 1354 9750
rect 1358 9746 1359 9750
rect 1363 9746 1663 9750
rect 1667 9746 1668 9750
rect 1672 9746 1972 9750
rect 1976 9746 1977 9750
rect 1981 9746 2281 9750
rect 2285 9746 2286 9750
rect 2290 9746 2590 9750
rect 2594 9746 2595 9750
rect 2599 9746 2899 9750
rect 2903 9746 2904 9750
rect 2908 9746 3208 9750
rect 3212 9746 3213 9750
rect 3217 9746 3517 9750
rect 3521 9746 3522 9750
rect 3526 9746 3652 9750
rect 3656 9746 3657 9750
rect 3661 9746 3826 9750
rect 3830 9746 3831 9750
rect 3835 9746 4602 9750
rect 570 9742 802 9746
rect 806 9742 807 9746
rect 811 9742 812 9746
rect 816 9742 817 9746
rect 821 9742 831 9746
rect 835 9742 836 9746
rect 840 9742 841 9746
rect 845 9742 846 9746
rect 850 9742 860 9746
rect 864 9742 865 9746
rect 869 9742 870 9746
rect 874 9742 875 9746
rect 879 9742 889 9746
rect 893 9742 894 9746
rect 898 9742 899 9746
rect 903 9742 904 9746
rect 908 9742 918 9746
rect 922 9742 923 9746
rect 927 9742 928 9746
rect 932 9742 933 9746
rect 937 9742 1319 9746
rect 1323 9742 1324 9746
rect 1328 9742 1329 9746
rect 1333 9742 1334 9746
rect 1338 9745 1628 9746
rect 1338 9742 1354 9745
rect 570 9741 1354 9742
rect 1358 9741 1359 9745
rect 1363 9742 1628 9745
rect 1632 9742 1633 9746
rect 1637 9742 1638 9746
rect 1642 9742 1643 9746
rect 1647 9745 1937 9746
rect 1647 9742 1663 9745
rect 1363 9741 1663 9742
rect 1667 9741 1668 9745
rect 1672 9742 1937 9745
rect 1941 9742 1942 9746
rect 1946 9742 1947 9746
rect 1951 9742 1952 9746
rect 1956 9745 2246 9746
rect 1956 9742 1972 9745
rect 1672 9741 1972 9742
rect 1976 9741 1977 9745
rect 1981 9742 2246 9745
rect 2250 9742 2251 9746
rect 2255 9742 2256 9746
rect 2260 9742 2261 9746
rect 2265 9745 2555 9746
rect 2265 9742 2281 9745
rect 1981 9741 2281 9742
rect 2285 9741 2286 9745
rect 2290 9742 2555 9745
rect 2559 9742 2560 9746
rect 2564 9742 2565 9746
rect 2569 9742 2570 9746
rect 2574 9745 2864 9746
rect 2574 9742 2590 9745
rect 2290 9741 2590 9742
rect 2594 9741 2595 9745
rect 2599 9742 2864 9745
rect 2868 9742 2869 9746
rect 2873 9742 2874 9746
rect 2878 9742 2879 9746
rect 2883 9745 3173 9746
rect 2883 9742 2899 9745
rect 2599 9741 2899 9742
rect 2903 9741 2904 9745
rect 2908 9742 3173 9745
rect 3177 9742 3178 9746
rect 3182 9742 3183 9746
rect 3187 9742 3188 9746
rect 3192 9745 3482 9746
rect 3192 9742 3208 9745
rect 2908 9741 3208 9742
rect 3212 9741 3213 9745
rect 3217 9742 3482 9745
rect 3486 9742 3487 9746
rect 3491 9742 3492 9746
rect 3496 9742 3497 9746
rect 3501 9745 3791 9746
rect 3501 9742 3517 9745
rect 3217 9741 3517 9742
rect 3521 9741 3522 9745
rect 3526 9741 3652 9745
rect 3656 9741 3657 9745
rect 3661 9742 3791 9745
rect 3795 9742 3796 9746
rect 3800 9742 3801 9746
rect 3805 9742 3806 9746
rect 3810 9745 4100 9746
rect 3810 9742 3826 9745
rect 3661 9741 3826 9742
rect 3830 9741 3831 9745
rect 3835 9742 4100 9745
rect 4104 9742 4105 9746
rect 4109 9742 4110 9746
rect 4114 9742 4115 9746
rect 4119 9742 4292 9746
rect 4296 9742 4297 9746
rect 4301 9742 4302 9746
rect 4306 9742 4307 9746
rect 4311 9742 4318 9746
rect 4322 9742 4323 9746
rect 4327 9742 4328 9746
rect 4332 9742 4333 9746
rect 4337 9742 4344 9746
rect 4348 9742 4349 9746
rect 4353 9742 4354 9746
rect 4358 9742 4359 9746
rect 4363 9742 4370 9746
rect 4374 9742 4375 9746
rect 4379 9742 4380 9746
rect 4384 9742 4385 9746
rect 4389 9742 4396 9746
rect 4400 9742 4401 9746
rect 4405 9742 4406 9746
rect 4410 9742 4411 9746
rect 4415 9742 4602 9746
rect 3835 9741 4602 9742
rect 570 9740 2167 9741
rect 570 9736 1354 9740
rect 1358 9736 1359 9740
rect 1363 9736 1663 9740
rect 1667 9736 1668 9740
rect 1672 9736 1972 9740
rect 1976 9736 1977 9740
rect 1981 9736 2167 9740
rect 2172 9740 4602 9741
rect 2172 9736 2281 9740
rect 2285 9736 2286 9740
rect 2290 9736 2590 9740
rect 2594 9736 2595 9740
rect 2599 9736 2899 9740
rect 2903 9736 2904 9740
rect 2908 9736 3208 9740
rect 3212 9736 3213 9740
rect 3217 9736 3517 9740
rect 3521 9736 3522 9740
rect 3526 9736 3826 9740
rect 3830 9736 3831 9740
rect 3835 9736 4602 9740
rect 570 9732 802 9736
rect 806 9732 807 9736
rect 811 9732 812 9736
rect 816 9732 817 9736
rect 821 9732 831 9736
rect 835 9732 836 9736
rect 840 9732 841 9736
rect 845 9732 846 9736
rect 850 9732 860 9736
rect 864 9732 865 9736
rect 869 9732 870 9736
rect 874 9732 875 9736
rect 879 9732 889 9736
rect 893 9732 894 9736
rect 898 9732 899 9736
rect 903 9732 904 9736
rect 908 9732 918 9736
rect 922 9732 923 9736
rect 927 9732 928 9736
rect 932 9732 933 9736
rect 937 9732 1319 9736
rect 1323 9732 1324 9736
rect 1328 9732 1329 9736
rect 1333 9732 1334 9736
rect 1338 9732 1628 9736
rect 1632 9732 1633 9736
rect 1637 9732 1638 9736
rect 1642 9732 1643 9736
rect 1647 9732 1937 9736
rect 1941 9732 1942 9736
rect 1946 9732 1947 9736
rect 1951 9732 1952 9736
rect 1956 9732 2246 9736
rect 2250 9732 2251 9736
rect 2255 9732 2256 9736
rect 2260 9732 2261 9736
rect 2265 9732 2555 9736
rect 2559 9732 2560 9736
rect 2564 9732 2565 9736
rect 2569 9732 2570 9736
rect 2574 9732 2864 9736
rect 2868 9732 2869 9736
rect 2873 9732 2874 9736
rect 2878 9732 2879 9736
rect 2883 9732 3173 9736
rect 3177 9732 3178 9736
rect 3182 9732 3183 9736
rect 3187 9732 3188 9736
rect 3192 9732 3482 9736
rect 3486 9732 3487 9736
rect 3491 9732 3492 9736
rect 3496 9732 3497 9736
rect 3501 9732 3791 9736
rect 3795 9732 3796 9736
rect 3800 9732 3801 9736
rect 3805 9732 3806 9736
rect 3810 9732 4100 9736
rect 4104 9732 4105 9736
rect 4109 9732 4110 9736
rect 4114 9732 4115 9736
rect 4119 9732 4292 9736
rect 4296 9732 4297 9736
rect 4301 9732 4302 9736
rect 4306 9732 4307 9736
rect 4311 9732 4318 9736
rect 4322 9732 4323 9736
rect 4327 9732 4328 9736
rect 4332 9732 4333 9736
rect 4337 9732 4344 9736
rect 4348 9732 4349 9736
rect 4353 9732 4354 9736
rect 4358 9732 4359 9736
rect 4363 9732 4370 9736
rect 4374 9732 4375 9736
rect 4379 9732 4380 9736
rect 4384 9732 4385 9736
rect 4389 9732 4396 9736
rect 4400 9732 4401 9736
rect 4405 9732 4406 9736
rect 4410 9732 4411 9736
rect 4415 9732 4602 9736
rect 570 9729 4602 9732
rect 570 9622 650 9729
rect 570 9618 613 9622
rect 617 9618 623 9622
rect 627 9618 633 9622
rect 637 9618 643 9622
rect 647 9618 650 9622
rect 570 9617 650 9618
rect 570 9613 613 9617
rect 617 9613 623 9617
rect 627 9613 633 9617
rect 637 9613 643 9617
rect 647 9613 650 9617
rect 570 9612 650 9613
rect 570 9608 613 9612
rect 617 9608 623 9612
rect 627 9608 633 9612
rect 637 9608 643 9612
rect 647 9608 650 9612
rect 570 9607 650 9608
rect 570 9603 613 9607
rect 617 9603 623 9607
rect 627 9603 633 9607
rect 637 9603 643 9607
rect 647 9603 650 9607
rect 570 9596 650 9603
rect 570 9592 613 9596
rect 617 9592 623 9596
rect 627 9592 633 9596
rect 637 9592 643 9596
rect 647 9592 650 9596
rect 570 9591 650 9592
rect 570 9587 613 9591
rect 617 9587 623 9591
rect 627 9587 633 9591
rect 637 9587 643 9591
rect 647 9587 650 9591
rect 570 9586 650 9587
rect 570 9582 613 9586
rect 617 9582 623 9586
rect 627 9582 633 9586
rect 637 9582 643 9586
rect 647 9582 650 9586
rect 570 9581 650 9582
rect 570 9577 613 9581
rect 617 9577 623 9581
rect 627 9577 633 9581
rect 637 9577 643 9581
rect 647 9577 650 9581
rect 570 9570 650 9577
rect 570 9566 613 9570
rect 617 9566 623 9570
rect 627 9566 633 9570
rect 637 9566 643 9570
rect 647 9566 650 9570
rect 570 9565 650 9566
rect 570 9561 613 9565
rect 617 9561 623 9565
rect 627 9561 633 9565
rect 637 9561 643 9565
rect 647 9561 650 9565
rect 570 9560 650 9561
rect 570 9556 613 9560
rect 617 9556 623 9560
rect 627 9556 633 9560
rect 637 9556 643 9560
rect 647 9556 650 9560
rect 570 9555 650 9556
rect 570 9551 613 9555
rect 617 9551 623 9555
rect 627 9551 633 9555
rect 637 9551 643 9555
rect 647 9551 650 9555
rect 570 9544 650 9551
rect 570 9540 613 9544
rect 617 9540 623 9544
rect 627 9540 633 9544
rect 637 9540 643 9544
rect 647 9540 650 9544
rect 570 9539 650 9540
rect 570 9535 613 9539
rect 617 9535 623 9539
rect 627 9535 633 9539
rect 637 9535 643 9539
rect 647 9535 650 9539
rect 570 9534 650 9535
rect 570 9530 613 9534
rect 617 9530 623 9534
rect 627 9530 633 9534
rect 637 9530 643 9534
rect 647 9530 650 9534
rect 570 9529 650 9530
rect 570 9525 613 9529
rect 617 9525 623 9529
rect 627 9525 633 9529
rect 637 9525 643 9529
rect 647 9525 650 9529
rect 570 9518 650 9525
rect 570 9514 613 9518
rect 617 9514 623 9518
rect 627 9514 633 9518
rect 637 9514 643 9518
rect 647 9514 650 9518
rect 570 9513 650 9514
rect 570 9509 613 9513
rect 617 9509 623 9513
rect 627 9509 633 9513
rect 637 9509 643 9513
rect 647 9509 650 9513
rect 570 9508 650 9509
rect 570 9504 613 9508
rect 617 9504 623 9508
rect 627 9504 633 9508
rect 637 9504 643 9508
rect 647 9504 650 9508
rect 570 9503 650 9504
rect 570 9499 613 9503
rect 617 9499 623 9503
rect 627 9499 633 9503
rect 637 9499 643 9503
rect 647 9499 650 9503
rect 570 9325 650 9499
rect 570 9321 613 9325
rect 617 9321 623 9325
rect 627 9321 633 9325
rect 637 9321 643 9325
rect 647 9321 650 9325
rect 570 9320 650 9321
rect 570 9316 613 9320
rect 617 9316 623 9320
rect 627 9316 633 9320
rect 637 9316 643 9320
rect 647 9316 650 9320
rect 570 9315 650 9316
rect 570 9311 613 9315
rect 617 9311 623 9315
rect 627 9311 633 9315
rect 637 9311 643 9315
rect 647 9311 650 9315
rect 570 9310 650 9311
rect 570 9306 613 9310
rect 617 9306 623 9310
rect 627 9306 633 9310
rect 637 9306 643 9310
rect 647 9306 650 9310
rect 570 9016 650 9306
rect 570 9012 613 9016
rect 617 9012 623 9016
rect 627 9012 633 9016
rect 637 9012 643 9016
rect 647 9012 650 9016
rect 570 9011 650 9012
rect 570 9007 613 9011
rect 617 9007 623 9011
rect 627 9007 633 9011
rect 637 9007 643 9011
rect 647 9007 650 9011
rect 570 9006 650 9007
rect 570 9002 613 9006
rect 617 9002 623 9006
rect 627 9002 633 9006
rect 637 9002 643 9006
rect 647 9002 650 9006
rect 570 9001 650 9002
rect 570 8997 613 9001
rect 617 8997 623 9001
rect 627 8997 633 9001
rect 637 8997 643 9001
rect 647 8997 650 9001
rect 570 8707 650 8997
rect 570 8703 613 8707
rect 617 8703 623 8707
rect 627 8703 633 8707
rect 637 8703 643 8707
rect 647 8703 650 8707
rect 570 8702 650 8703
rect 570 8698 613 8702
rect 617 8698 623 8702
rect 627 8698 633 8702
rect 637 8698 643 8702
rect 647 8698 650 8702
rect 570 8697 650 8698
rect 570 8693 613 8697
rect 617 8693 623 8697
rect 627 8693 633 8697
rect 637 8693 643 8697
rect 647 8693 650 8697
rect 570 8692 650 8693
rect 570 8688 613 8692
rect 617 8688 623 8692
rect 627 8688 633 8692
rect 637 8688 643 8692
rect 647 8688 650 8692
rect 570 8398 650 8688
rect 570 8394 613 8398
rect 617 8394 623 8398
rect 627 8394 633 8398
rect 637 8394 643 8398
rect 647 8394 650 8398
rect 570 8393 650 8394
rect 570 8389 613 8393
rect 617 8389 623 8393
rect 627 8389 633 8393
rect 637 8389 643 8393
rect 647 8389 650 8393
rect 570 8388 650 8389
rect 570 8384 613 8388
rect 617 8384 623 8388
rect 627 8384 633 8388
rect 637 8384 643 8388
rect 647 8384 650 8388
rect 570 8383 650 8384
rect 570 8379 613 8383
rect 617 8379 623 8383
rect 627 8379 633 8383
rect 637 8379 643 8383
rect 647 8379 650 8383
rect 570 8089 650 8379
rect 570 8085 613 8089
rect 617 8085 623 8089
rect 627 8085 633 8089
rect 637 8085 643 8089
rect 647 8085 650 8089
rect 570 8084 650 8085
rect 570 8080 613 8084
rect 617 8080 623 8084
rect 627 8080 633 8084
rect 637 8080 643 8084
rect 647 8080 650 8084
rect 570 8079 650 8080
rect 570 8075 613 8079
rect 617 8075 623 8079
rect 627 8075 633 8079
rect 637 8075 643 8079
rect 647 8075 650 8079
rect 570 8074 650 8075
rect 570 8070 613 8074
rect 617 8070 623 8074
rect 627 8070 633 8074
rect 637 8070 643 8074
rect 647 8070 650 8074
rect 570 7780 650 8070
rect 570 7776 613 7780
rect 617 7776 623 7780
rect 627 7776 633 7780
rect 637 7776 643 7780
rect 647 7776 650 7780
rect 570 7775 650 7776
rect 570 7771 613 7775
rect 617 7771 623 7775
rect 627 7771 633 7775
rect 637 7771 643 7775
rect 647 7771 650 7775
rect 570 7770 650 7771
rect 570 7766 613 7770
rect 617 7766 623 7770
rect 627 7766 633 7770
rect 637 7766 643 7770
rect 647 7766 650 7770
rect 570 7765 650 7766
rect 570 7761 613 7765
rect 617 7761 623 7765
rect 627 7761 633 7765
rect 637 7761 643 7765
rect 647 7761 650 7765
rect 570 7471 650 7761
rect 570 7467 613 7471
rect 617 7467 623 7471
rect 627 7467 633 7471
rect 637 7467 643 7471
rect 647 7467 650 7471
rect 570 7466 650 7467
rect 570 7462 613 7466
rect 617 7462 623 7466
rect 627 7462 633 7466
rect 637 7462 643 7466
rect 647 7462 650 7466
rect 570 7461 650 7462
rect 570 7457 613 7461
rect 617 7457 623 7461
rect 627 7457 633 7461
rect 637 7457 643 7461
rect 647 7457 650 7461
rect 570 7456 650 7457
rect 570 7452 613 7456
rect 617 7452 623 7456
rect 627 7452 633 7456
rect 637 7452 643 7456
rect 647 7452 650 7456
rect 570 7162 650 7452
rect 570 7158 613 7162
rect 617 7158 623 7162
rect 627 7158 633 7162
rect 637 7158 643 7162
rect 647 7158 650 7162
rect 570 7157 650 7158
rect 570 7153 613 7157
rect 617 7153 623 7157
rect 627 7153 633 7157
rect 637 7153 643 7157
rect 647 7153 650 7157
rect 570 7152 650 7153
rect 570 7148 613 7152
rect 617 7148 623 7152
rect 627 7148 633 7152
rect 637 7148 643 7152
rect 647 7148 650 7152
rect 570 7147 650 7148
rect 570 7143 613 7147
rect 617 7143 623 7147
rect 627 7143 633 7147
rect 637 7143 643 7147
rect 647 7143 650 7147
rect 570 6853 650 7143
rect 570 6849 613 6853
rect 617 6849 623 6853
rect 627 6849 633 6853
rect 637 6849 643 6853
rect 647 6849 650 6853
rect 570 6848 650 6849
rect 570 6844 613 6848
rect 617 6844 623 6848
rect 627 6844 633 6848
rect 637 6844 643 6848
rect 647 6844 650 6848
rect 570 6843 650 6844
rect 570 6839 613 6843
rect 617 6839 623 6843
rect 627 6839 633 6843
rect 637 6839 643 6843
rect 647 6839 650 6843
rect 570 6838 650 6839
rect 570 6834 613 6838
rect 617 6834 623 6838
rect 627 6834 633 6838
rect 637 6834 643 6838
rect 647 6834 650 6838
rect 570 6544 650 6834
rect 570 6540 613 6544
rect 617 6540 623 6544
rect 627 6540 633 6544
rect 637 6540 643 6544
rect 647 6540 650 6544
rect 570 6539 650 6540
rect 570 6535 613 6539
rect 617 6535 623 6539
rect 627 6535 633 6539
rect 637 6535 643 6539
rect 647 6535 650 6539
rect 570 6534 650 6535
rect 570 6530 613 6534
rect 617 6530 623 6534
rect 627 6530 633 6534
rect 637 6530 643 6534
rect 647 6530 650 6534
rect 570 6529 650 6530
rect 570 6525 613 6529
rect 617 6525 623 6529
rect 627 6525 633 6529
rect 637 6525 643 6529
rect 647 6525 650 6529
rect 570 6144 650 6525
rect 570 6140 613 6144
rect 617 6140 623 6144
rect 627 6140 633 6144
rect 637 6140 643 6144
rect 647 6140 650 6144
rect 570 6139 650 6140
rect 570 6135 613 6139
rect 617 6135 623 6139
rect 627 6135 633 6139
rect 637 6135 643 6139
rect 647 6135 650 6139
rect 570 6134 650 6135
rect 570 6130 613 6134
rect 617 6130 623 6134
rect 627 6130 633 6134
rect 637 6130 643 6134
rect 647 6130 650 6134
rect 570 6129 650 6130
rect 570 6125 613 6129
rect 617 6125 623 6129
rect 627 6125 633 6129
rect 637 6125 643 6129
rect 647 6125 650 6129
rect 570 6115 650 6125
rect 570 6111 613 6115
rect 617 6111 623 6115
rect 627 6111 633 6115
rect 637 6111 643 6115
rect 647 6111 650 6115
rect 570 6110 650 6111
rect 570 6106 613 6110
rect 617 6106 623 6110
rect 627 6106 633 6110
rect 637 6106 643 6110
rect 647 6106 650 6110
rect 570 6105 650 6106
rect 570 6101 613 6105
rect 617 6101 623 6105
rect 627 6101 633 6105
rect 637 6101 643 6105
rect 647 6101 650 6105
rect 570 6100 650 6101
rect 570 6096 613 6100
rect 617 6096 623 6100
rect 627 6096 633 6100
rect 637 6096 643 6100
rect 647 6096 650 6100
rect 570 6086 650 6096
rect 570 6082 613 6086
rect 617 6082 623 6086
rect 627 6082 633 6086
rect 637 6082 643 6086
rect 647 6082 650 6086
rect 570 6081 650 6082
rect 570 6077 613 6081
rect 617 6077 623 6081
rect 627 6077 633 6081
rect 637 6077 643 6081
rect 647 6077 650 6081
rect 570 6076 650 6077
rect 570 6072 613 6076
rect 617 6072 623 6076
rect 627 6072 633 6076
rect 637 6072 643 6076
rect 647 6072 650 6076
rect 570 6071 650 6072
rect 570 6067 613 6071
rect 617 6067 623 6071
rect 627 6067 633 6071
rect 637 6067 643 6071
rect 647 6067 650 6071
rect 570 6057 650 6067
rect 570 6053 613 6057
rect 617 6053 623 6057
rect 627 6053 633 6057
rect 637 6053 643 6057
rect 647 6053 650 6057
rect 570 6052 650 6053
rect 570 6048 613 6052
rect 617 6048 623 6052
rect 627 6048 633 6052
rect 637 6048 643 6052
rect 647 6048 650 6052
rect 570 6047 650 6048
rect 570 6043 613 6047
rect 617 6043 623 6047
rect 627 6043 633 6047
rect 637 6043 643 6047
rect 647 6043 650 6047
rect 570 6042 650 6043
rect 570 6038 613 6042
rect 617 6038 623 6042
rect 627 6038 633 6042
rect 637 6038 643 6042
rect 647 6038 650 6042
rect 570 6028 650 6038
rect 570 6024 613 6028
rect 617 6024 623 6028
rect 627 6024 633 6028
rect 637 6024 643 6028
rect 647 6024 650 6028
rect 570 6023 650 6024
rect 570 6019 613 6023
rect 617 6019 623 6023
rect 627 6019 633 6023
rect 637 6019 643 6023
rect 647 6019 650 6023
rect 570 6018 650 6019
rect 570 6014 613 6018
rect 617 6014 623 6018
rect 627 6014 633 6018
rect 637 6014 643 6018
rect 647 6014 650 6018
rect 570 6013 650 6014
rect 570 6009 613 6013
rect 617 6009 623 6013
rect 627 6009 633 6013
rect 637 6009 643 6013
rect 647 6009 650 6013
rect 570 5857 650 6009
rect 654 9720 4518 9725
rect 654 9716 802 9720
rect 806 9716 807 9720
rect 811 9716 812 9720
rect 816 9716 817 9720
rect 821 9716 831 9720
rect 835 9716 836 9720
rect 840 9716 841 9720
rect 845 9716 846 9720
rect 850 9716 860 9720
rect 864 9716 865 9720
rect 869 9716 870 9720
rect 874 9716 875 9720
rect 879 9716 889 9720
rect 893 9716 894 9720
rect 898 9716 899 9720
rect 903 9716 904 9720
rect 908 9716 918 9720
rect 922 9716 923 9720
rect 927 9716 928 9720
rect 932 9716 933 9720
rect 937 9716 1319 9720
rect 1323 9716 1324 9720
rect 1328 9716 1329 9720
rect 1333 9716 1334 9720
rect 1338 9716 1628 9720
rect 1632 9716 1633 9720
rect 1637 9716 1638 9720
rect 1642 9716 1643 9720
rect 1647 9716 1937 9720
rect 1941 9716 1942 9720
rect 1946 9716 1947 9720
rect 1951 9716 1952 9720
rect 1956 9716 2246 9720
rect 2250 9716 2251 9720
rect 2255 9716 2256 9720
rect 2260 9716 2261 9720
rect 2265 9716 2555 9720
rect 2559 9716 2560 9720
rect 2564 9716 2565 9720
rect 2569 9716 2570 9720
rect 2574 9716 2864 9720
rect 2868 9716 2869 9720
rect 2873 9716 2874 9720
rect 2878 9716 2879 9720
rect 2883 9716 3173 9720
rect 3177 9716 3178 9720
rect 3182 9716 3183 9720
rect 3187 9716 3188 9720
rect 3192 9716 3482 9720
rect 3486 9716 3487 9720
rect 3491 9716 3492 9720
rect 3496 9716 3497 9720
rect 3501 9716 3791 9720
rect 3795 9716 3796 9720
rect 3800 9716 3801 9720
rect 3805 9716 3806 9720
rect 3810 9716 4100 9720
rect 4104 9716 4105 9720
rect 4109 9716 4110 9720
rect 4114 9716 4115 9720
rect 4119 9716 4292 9720
rect 4296 9716 4297 9720
rect 4301 9716 4302 9720
rect 4306 9716 4307 9720
rect 4311 9716 4318 9720
rect 4322 9716 4323 9720
rect 4327 9716 4328 9720
rect 4332 9716 4333 9720
rect 4337 9716 4344 9720
rect 4348 9716 4349 9720
rect 4353 9716 4354 9720
rect 4358 9716 4359 9720
rect 4363 9716 4370 9720
rect 4374 9716 4375 9720
rect 4379 9716 4380 9720
rect 4384 9716 4385 9720
rect 4389 9716 4396 9720
rect 4400 9716 4401 9720
rect 4405 9716 4406 9720
rect 4410 9716 4411 9720
rect 4415 9716 4518 9720
rect 654 9715 4518 9716
rect 654 9712 1489 9715
rect 654 9710 1387 9712
rect 654 9706 802 9710
rect 806 9706 807 9710
rect 811 9706 812 9710
rect 816 9706 817 9710
rect 821 9706 831 9710
rect 835 9706 836 9710
rect 840 9706 841 9710
rect 845 9706 846 9710
rect 850 9706 860 9710
rect 864 9706 865 9710
rect 869 9706 870 9710
rect 874 9706 875 9710
rect 879 9706 889 9710
rect 893 9706 894 9710
rect 898 9706 899 9710
rect 903 9706 904 9710
rect 908 9706 918 9710
rect 922 9706 923 9710
rect 927 9706 928 9710
rect 932 9706 933 9710
rect 937 9706 1319 9710
rect 1323 9706 1324 9710
rect 1328 9706 1329 9710
rect 1333 9706 1334 9710
rect 1338 9708 1387 9710
rect 1391 9708 1392 9712
rect 1396 9708 1397 9712
rect 1401 9708 1402 9712
rect 1406 9708 1407 9712
rect 1411 9708 1412 9712
rect 1416 9708 1417 9712
rect 1421 9708 1422 9712
rect 1426 9708 1427 9712
rect 1431 9708 1432 9712
rect 1436 9708 1437 9712
rect 1441 9708 1442 9712
rect 1446 9708 1447 9712
rect 1451 9711 1489 9712
rect 1493 9711 1494 9715
rect 1498 9712 3343 9715
rect 1498 9711 1569 9712
rect 1451 9710 1569 9711
rect 1451 9708 1489 9710
rect 1338 9707 1489 9708
rect 1338 9706 1387 9707
rect 654 9703 1387 9706
rect 1391 9703 1392 9707
rect 1396 9703 1397 9707
rect 1401 9703 1402 9707
rect 1406 9703 1407 9707
rect 1411 9703 1412 9707
rect 1416 9703 1417 9707
rect 1421 9703 1422 9707
rect 1426 9703 1427 9707
rect 1431 9703 1432 9707
rect 1436 9703 1437 9707
rect 1441 9703 1442 9707
rect 1446 9703 1447 9707
rect 1451 9706 1489 9707
rect 1493 9706 1494 9710
rect 1498 9708 1569 9710
rect 1573 9708 1574 9712
rect 1578 9708 1579 9712
rect 1583 9708 1584 9712
rect 1588 9708 1589 9712
rect 1593 9708 1594 9712
rect 1598 9708 1599 9712
rect 1603 9708 1604 9712
rect 1608 9708 1609 9712
rect 1613 9708 1614 9712
rect 1618 9708 1619 9712
rect 1623 9710 1696 9712
rect 1623 9708 1628 9710
rect 1498 9707 1628 9708
rect 1498 9706 1569 9707
rect 1451 9705 1569 9706
rect 1451 9703 1489 9705
rect 654 9701 1489 9703
rect 1493 9701 1494 9705
rect 1498 9703 1569 9705
rect 1573 9703 1574 9707
rect 1578 9703 1579 9707
rect 1583 9703 1584 9707
rect 1588 9703 1589 9707
rect 1593 9703 1594 9707
rect 1598 9703 1599 9707
rect 1603 9703 1604 9707
rect 1608 9703 1609 9707
rect 1613 9703 1614 9707
rect 1618 9703 1619 9707
rect 1623 9706 1628 9707
rect 1632 9706 1633 9710
rect 1637 9706 1638 9710
rect 1642 9706 1643 9710
rect 1647 9708 1696 9710
rect 1700 9708 1701 9712
rect 1705 9708 1706 9712
rect 1710 9708 1711 9712
rect 1715 9708 1716 9712
rect 1720 9708 1721 9712
rect 1725 9708 1726 9712
rect 1730 9708 1731 9712
rect 1735 9708 1736 9712
rect 1740 9708 1741 9712
rect 1745 9708 1746 9712
rect 1750 9708 1751 9712
rect 1755 9708 1756 9712
rect 1760 9708 1878 9712
rect 1882 9708 1883 9712
rect 1887 9708 1888 9712
rect 1892 9708 1893 9712
rect 1897 9708 1898 9712
rect 1902 9708 1903 9712
rect 1907 9708 1908 9712
rect 1912 9708 1913 9712
rect 1917 9708 1918 9712
rect 1922 9708 1923 9712
rect 1927 9708 1928 9712
rect 1932 9710 2005 9712
rect 1932 9708 1937 9710
rect 1647 9707 1937 9708
rect 1647 9706 1696 9707
rect 1623 9703 1696 9706
rect 1700 9703 1701 9707
rect 1705 9703 1706 9707
rect 1710 9703 1711 9707
rect 1715 9703 1716 9707
rect 1720 9703 1721 9707
rect 1725 9703 1726 9707
rect 1730 9703 1731 9707
rect 1735 9703 1736 9707
rect 1740 9703 1741 9707
rect 1745 9703 1746 9707
rect 1750 9703 1751 9707
rect 1755 9703 1756 9707
rect 1760 9703 1878 9707
rect 1882 9703 1883 9707
rect 1887 9703 1888 9707
rect 1892 9703 1893 9707
rect 1897 9703 1898 9707
rect 1902 9703 1903 9707
rect 1907 9703 1908 9707
rect 1912 9703 1913 9707
rect 1917 9703 1918 9707
rect 1922 9703 1923 9707
rect 1927 9703 1928 9707
rect 1932 9706 1937 9707
rect 1941 9706 1942 9710
rect 1946 9706 1947 9710
rect 1951 9706 1952 9710
rect 1956 9708 2005 9710
rect 2009 9708 2010 9712
rect 2014 9708 2015 9712
rect 2019 9708 2020 9712
rect 2024 9708 2025 9712
rect 2029 9708 2030 9712
rect 2034 9708 2035 9712
rect 2039 9708 2040 9712
rect 2044 9708 2045 9712
rect 2049 9708 2050 9712
rect 2054 9708 2055 9712
rect 2059 9708 2060 9712
rect 2064 9708 2065 9712
rect 2069 9708 2187 9712
rect 2191 9708 2192 9712
rect 2196 9708 2197 9712
rect 2201 9708 2202 9712
rect 2206 9708 2207 9712
rect 2211 9708 2212 9712
rect 2216 9708 2217 9712
rect 2221 9708 2222 9712
rect 2226 9708 2227 9712
rect 2231 9708 2232 9712
rect 2236 9708 2237 9712
rect 2241 9710 2314 9712
rect 2241 9708 2246 9710
rect 1956 9707 2246 9708
rect 1956 9706 2005 9707
rect 1932 9703 2005 9706
rect 2009 9703 2010 9707
rect 2014 9703 2015 9707
rect 2019 9703 2020 9707
rect 2024 9703 2025 9707
rect 2029 9703 2030 9707
rect 2034 9703 2035 9707
rect 2039 9703 2040 9707
rect 2044 9703 2045 9707
rect 2049 9703 2050 9707
rect 2054 9703 2055 9707
rect 2059 9703 2060 9707
rect 2064 9703 2065 9707
rect 2069 9703 2187 9707
rect 2191 9703 2192 9707
rect 2196 9703 2197 9707
rect 2201 9703 2202 9707
rect 2206 9703 2207 9707
rect 2211 9703 2212 9707
rect 2216 9703 2217 9707
rect 2221 9703 2222 9707
rect 2226 9703 2227 9707
rect 2231 9703 2232 9707
rect 2236 9703 2237 9707
rect 2241 9706 2246 9707
rect 2250 9706 2251 9710
rect 2255 9706 2256 9710
rect 2260 9706 2261 9710
rect 2265 9708 2314 9710
rect 2318 9708 2319 9712
rect 2323 9708 2324 9712
rect 2328 9708 2329 9712
rect 2333 9708 2334 9712
rect 2338 9708 2339 9712
rect 2343 9708 2344 9712
rect 2348 9708 2349 9712
rect 2353 9708 2354 9712
rect 2358 9708 2359 9712
rect 2363 9708 2364 9712
rect 2368 9708 2369 9712
rect 2373 9708 2374 9712
rect 2378 9708 2496 9712
rect 2500 9708 2501 9712
rect 2505 9708 2506 9712
rect 2510 9708 2511 9712
rect 2515 9708 2516 9712
rect 2520 9708 2521 9712
rect 2525 9708 2526 9712
rect 2530 9708 2531 9712
rect 2535 9708 2536 9712
rect 2540 9708 2541 9712
rect 2545 9708 2546 9712
rect 2550 9710 2623 9712
rect 2550 9708 2555 9710
rect 2265 9707 2555 9708
rect 2265 9706 2314 9707
rect 2241 9703 2314 9706
rect 2318 9703 2319 9707
rect 2323 9703 2324 9707
rect 2328 9703 2329 9707
rect 2333 9703 2334 9707
rect 2338 9703 2339 9707
rect 2343 9703 2344 9707
rect 2348 9703 2349 9707
rect 2353 9703 2354 9707
rect 2358 9703 2359 9707
rect 2363 9703 2364 9707
rect 2368 9703 2369 9707
rect 2373 9703 2374 9707
rect 2378 9703 2496 9707
rect 2500 9703 2501 9707
rect 2505 9703 2506 9707
rect 2510 9703 2511 9707
rect 2515 9703 2516 9707
rect 2520 9703 2521 9707
rect 2525 9703 2526 9707
rect 2530 9703 2531 9707
rect 2535 9703 2536 9707
rect 2540 9703 2541 9707
rect 2545 9703 2546 9707
rect 2550 9706 2555 9707
rect 2559 9706 2560 9710
rect 2564 9706 2565 9710
rect 2569 9706 2570 9710
rect 2574 9708 2623 9710
rect 2627 9708 2628 9712
rect 2632 9708 2633 9712
rect 2637 9708 2638 9712
rect 2642 9708 2643 9712
rect 2647 9708 2648 9712
rect 2652 9708 2653 9712
rect 2657 9708 2658 9712
rect 2662 9708 2663 9712
rect 2667 9708 2668 9712
rect 2672 9708 2673 9712
rect 2677 9708 2678 9712
rect 2682 9708 2683 9712
rect 2687 9708 2805 9712
rect 2809 9708 2810 9712
rect 2814 9708 2815 9712
rect 2819 9708 2820 9712
rect 2824 9708 2825 9712
rect 2829 9708 2830 9712
rect 2834 9708 2835 9712
rect 2839 9708 2840 9712
rect 2844 9708 2845 9712
rect 2849 9708 2850 9712
rect 2854 9708 2855 9712
rect 2859 9710 2932 9712
rect 2859 9708 2864 9710
rect 2574 9707 2864 9708
rect 2574 9706 2623 9707
rect 2550 9703 2623 9706
rect 2627 9703 2628 9707
rect 2632 9703 2633 9707
rect 2637 9703 2638 9707
rect 2642 9703 2643 9707
rect 2647 9703 2648 9707
rect 2652 9703 2653 9707
rect 2657 9703 2658 9707
rect 2662 9703 2663 9707
rect 2667 9703 2668 9707
rect 2672 9703 2673 9707
rect 2677 9703 2678 9707
rect 2682 9703 2683 9707
rect 2687 9703 2805 9707
rect 2809 9703 2810 9707
rect 2814 9703 2815 9707
rect 2819 9703 2820 9707
rect 2824 9703 2825 9707
rect 2829 9703 2830 9707
rect 2834 9703 2835 9707
rect 2839 9703 2840 9707
rect 2844 9703 2845 9707
rect 2849 9703 2850 9707
rect 2854 9703 2855 9707
rect 2859 9706 2864 9707
rect 2868 9706 2869 9710
rect 2873 9706 2874 9710
rect 2878 9706 2879 9710
rect 2883 9708 2932 9710
rect 2936 9708 2937 9712
rect 2941 9708 2942 9712
rect 2946 9708 2947 9712
rect 2951 9708 2952 9712
rect 2956 9708 2957 9712
rect 2961 9708 2962 9712
rect 2966 9708 2967 9712
rect 2971 9708 2972 9712
rect 2976 9708 2977 9712
rect 2981 9708 2982 9712
rect 2986 9708 2987 9712
rect 2991 9708 2992 9712
rect 2996 9708 3114 9712
rect 3118 9708 3119 9712
rect 3123 9708 3124 9712
rect 3128 9708 3129 9712
rect 3133 9708 3134 9712
rect 3138 9708 3139 9712
rect 3143 9708 3144 9712
rect 3148 9708 3149 9712
rect 3153 9708 3154 9712
rect 3158 9708 3159 9712
rect 3163 9708 3164 9712
rect 3168 9710 3241 9712
rect 3168 9708 3173 9710
rect 2883 9707 3173 9708
rect 2883 9706 2932 9707
rect 2859 9703 2932 9706
rect 2936 9703 2937 9707
rect 2941 9703 2942 9707
rect 2946 9703 2947 9707
rect 2951 9703 2952 9707
rect 2956 9703 2957 9707
rect 2961 9703 2962 9707
rect 2966 9703 2967 9707
rect 2971 9703 2972 9707
rect 2976 9703 2977 9707
rect 2981 9703 2982 9707
rect 2986 9703 2987 9707
rect 2991 9703 2992 9707
rect 2996 9703 3114 9707
rect 3118 9703 3119 9707
rect 3123 9703 3124 9707
rect 3128 9703 3129 9707
rect 3133 9703 3134 9707
rect 3138 9703 3139 9707
rect 3143 9703 3144 9707
rect 3148 9703 3149 9707
rect 3153 9703 3154 9707
rect 3158 9703 3159 9707
rect 3163 9703 3164 9707
rect 3168 9706 3173 9707
rect 3177 9706 3178 9710
rect 3182 9706 3183 9710
rect 3187 9706 3188 9710
rect 3192 9708 3241 9710
rect 3245 9708 3246 9712
rect 3250 9708 3251 9712
rect 3255 9708 3256 9712
rect 3260 9708 3261 9712
rect 3265 9708 3266 9712
rect 3270 9708 3271 9712
rect 3275 9708 3276 9712
rect 3280 9708 3281 9712
rect 3285 9708 3286 9712
rect 3290 9708 3291 9712
rect 3295 9708 3296 9712
rect 3300 9708 3301 9712
rect 3305 9711 3343 9712
rect 3347 9711 3348 9715
rect 3352 9712 4518 9715
rect 3352 9711 3423 9712
rect 3305 9710 3423 9711
rect 3305 9708 3343 9710
rect 3192 9707 3343 9708
rect 3192 9706 3241 9707
rect 3168 9703 3241 9706
rect 3245 9703 3246 9707
rect 3250 9703 3251 9707
rect 3255 9703 3256 9707
rect 3260 9703 3261 9707
rect 3265 9703 3266 9707
rect 3270 9703 3271 9707
rect 3275 9703 3276 9707
rect 3280 9703 3281 9707
rect 3285 9703 3286 9707
rect 3290 9703 3291 9707
rect 3295 9703 3296 9707
rect 3300 9703 3301 9707
rect 3305 9706 3343 9707
rect 3347 9706 3348 9710
rect 3352 9708 3423 9710
rect 3427 9708 3428 9712
rect 3432 9708 3433 9712
rect 3437 9708 3438 9712
rect 3442 9708 3443 9712
rect 3447 9708 3448 9712
rect 3452 9708 3453 9712
rect 3457 9708 3458 9712
rect 3462 9708 3463 9712
rect 3467 9708 3468 9712
rect 3472 9708 3473 9712
rect 3477 9710 3550 9712
rect 3477 9708 3482 9710
rect 3352 9707 3482 9708
rect 3352 9706 3423 9707
rect 3305 9705 3423 9706
rect 3305 9703 3343 9705
rect 1498 9701 3343 9703
rect 3347 9701 3348 9705
rect 3352 9703 3423 9705
rect 3427 9703 3428 9707
rect 3432 9703 3433 9707
rect 3437 9703 3438 9707
rect 3442 9703 3443 9707
rect 3447 9703 3448 9707
rect 3452 9703 3453 9707
rect 3457 9703 3458 9707
rect 3462 9703 3463 9707
rect 3467 9703 3468 9707
rect 3472 9703 3473 9707
rect 3477 9706 3482 9707
rect 3486 9706 3487 9710
rect 3491 9706 3492 9710
rect 3496 9706 3497 9710
rect 3501 9708 3550 9710
rect 3554 9708 3555 9712
rect 3559 9708 3560 9712
rect 3564 9708 3565 9712
rect 3569 9708 3570 9712
rect 3574 9708 3575 9712
rect 3579 9708 3580 9712
rect 3584 9708 3585 9712
rect 3589 9708 3590 9712
rect 3594 9708 3595 9712
rect 3599 9708 3600 9712
rect 3604 9708 3605 9712
rect 3609 9708 3610 9712
rect 3614 9708 3732 9712
rect 3736 9708 3737 9712
rect 3741 9708 3742 9712
rect 3746 9708 3747 9712
rect 3751 9708 3752 9712
rect 3756 9708 3757 9712
rect 3761 9708 3762 9712
rect 3766 9708 3767 9712
rect 3771 9708 3772 9712
rect 3776 9708 3777 9712
rect 3781 9708 3782 9712
rect 3786 9710 3859 9712
rect 3786 9708 3791 9710
rect 3501 9707 3791 9708
rect 3501 9706 3550 9707
rect 3477 9703 3550 9706
rect 3554 9703 3555 9707
rect 3559 9703 3560 9707
rect 3564 9703 3565 9707
rect 3569 9703 3570 9707
rect 3574 9703 3575 9707
rect 3579 9703 3580 9707
rect 3584 9703 3585 9707
rect 3589 9703 3590 9707
rect 3594 9703 3595 9707
rect 3599 9703 3600 9707
rect 3604 9703 3605 9707
rect 3609 9703 3610 9707
rect 3614 9703 3732 9707
rect 3736 9703 3737 9707
rect 3741 9703 3742 9707
rect 3746 9703 3747 9707
rect 3751 9703 3752 9707
rect 3756 9703 3757 9707
rect 3761 9703 3762 9707
rect 3766 9703 3767 9707
rect 3771 9703 3772 9707
rect 3776 9703 3777 9707
rect 3781 9703 3782 9707
rect 3786 9706 3791 9707
rect 3795 9706 3796 9710
rect 3800 9706 3801 9710
rect 3805 9706 3806 9710
rect 3810 9708 3859 9710
rect 3863 9708 3864 9712
rect 3868 9708 3869 9712
rect 3873 9708 3874 9712
rect 3878 9708 3879 9712
rect 3883 9708 3884 9712
rect 3888 9708 3889 9712
rect 3893 9708 3894 9712
rect 3898 9708 3899 9712
rect 3903 9708 3904 9712
rect 3908 9708 3909 9712
rect 3913 9708 3914 9712
rect 3918 9708 3919 9712
rect 3923 9708 4041 9712
rect 4045 9708 4046 9712
rect 4050 9708 4051 9712
rect 4055 9708 4056 9712
rect 4060 9708 4061 9712
rect 4065 9708 4066 9712
rect 4070 9708 4071 9712
rect 4075 9708 4076 9712
rect 4080 9708 4081 9712
rect 4085 9708 4086 9712
rect 4090 9708 4091 9712
rect 4095 9710 4518 9712
rect 4095 9708 4100 9710
rect 3810 9707 4100 9708
rect 3810 9706 3859 9707
rect 3786 9703 3859 9706
rect 3863 9703 3864 9707
rect 3868 9703 3869 9707
rect 3873 9703 3874 9707
rect 3878 9703 3879 9707
rect 3883 9703 3884 9707
rect 3888 9703 3889 9707
rect 3893 9703 3894 9707
rect 3898 9703 3899 9707
rect 3903 9703 3904 9707
rect 3908 9703 3909 9707
rect 3913 9703 3914 9707
rect 3918 9703 3919 9707
rect 3923 9703 4041 9707
rect 4045 9703 4046 9707
rect 4050 9703 4051 9707
rect 4055 9703 4056 9707
rect 4060 9703 4061 9707
rect 4065 9703 4066 9707
rect 4070 9703 4071 9707
rect 4075 9703 4076 9707
rect 4080 9703 4081 9707
rect 4085 9703 4086 9707
rect 4090 9703 4091 9707
rect 4095 9706 4100 9707
rect 4104 9706 4105 9710
rect 4109 9706 4110 9710
rect 4114 9706 4115 9710
rect 4119 9706 4292 9710
rect 4296 9706 4297 9710
rect 4301 9706 4302 9710
rect 4306 9706 4307 9710
rect 4311 9706 4318 9710
rect 4322 9706 4323 9710
rect 4327 9706 4328 9710
rect 4332 9706 4333 9710
rect 4337 9706 4344 9710
rect 4348 9706 4349 9710
rect 4353 9706 4354 9710
rect 4358 9706 4359 9710
rect 4363 9706 4370 9710
rect 4374 9706 4375 9710
rect 4379 9706 4380 9710
rect 4384 9706 4385 9710
rect 4389 9706 4396 9710
rect 4400 9706 4401 9710
rect 4405 9706 4406 9710
rect 4410 9706 4411 9710
rect 4415 9706 4518 9710
rect 4095 9703 4518 9706
rect 3352 9701 4518 9703
rect 654 9700 4518 9701
rect 654 9696 802 9700
rect 806 9696 807 9700
rect 811 9696 812 9700
rect 816 9696 817 9700
rect 821 9696 831 9700
rect 835 9696 836 9700
rect 840 9696 841 9700
rect 845 9696 846 9700
rect 850 9696 860 9700
rect 864 9696 865 9700
rect 869 9696 870 9700
rect 874 9696 875 9700
rect 879 9696 889 9700
rect 893 9696 894 9700
rect 898 9696 899 9700
rect 903 9696 904 9700
rect 908 9696 918 9700
rect 922 9696 923 9700
rect 927 9696 928 9700
rect 932 9696 933 9700
rect 937 9696 1319 9700
rect 1323 9696 1324 9700
rect 1328 9696 1329 9700
rect 1333 9696 1334 9700
rect 1338 9696 1489 9700
rect 1493 9696 1494 9700
rect 1498 9696 1628 9700
rect 1632 9696 1633 9700
rect 1637 9696 1638 9700
rect 1642 9696 1643 9700
rect 1647 9696 1937 9700
rect 1941 9696 1942 9700
rect 1946 9696 1947 9700
rect 1951 9696 1952 9700
rect 1956 9696 2246 9700
rect 2250 9696 2251 9700
rect 2255 9696 2256 9700
rect 2260 9696 2261 9700
rect 2265 9696 2555 9700
rect 2559 9696 2560 9700
rect 2564 9696 2565 9700
rect 2569 9696 2570 9700
rect 2574 9696 2864 9700
rect 2868 9696 2869 9700
rect 2873 9696 2874 9700
rect 2878 9696 2879 9700
rect 2883 9696 3173 9700
rect 3177 9696 3178 9700
rect 3182 9696 3183 9700
rect 3187 9696 3188 9700
rect 3192 9696 3343 9700
rect 3347 9696 3348 9700
rect 3352 9696 3482 9700
rect 3486 9696 3487 9700
rect 3491 9696 3492 9700
rect 3496 9696 3497 9700
rect 3501 9696 3791 9700
rect 3795 9696 3796 9700
rect 3800 9696 3801 9700
rect 3805 9696 3806 9700
rect 3810 9696 4100 9700
rect 4104 9696 4105 9700
rect 4109 9696 4110 9700
rect 4114 9696 4115 9700
rect 4119 9696 4292 9700
rect 4296 9696 4297 9700
rect 4301 9696 4302 9700
rect 4306 9696 4307 9700
rect 4311 9696 4318 9700
rect 4322 9696 4323 9700
rect 4327 9696 4328 9700
rect 4332 9696 4333 9700
rect 4337 9696 4344 9700
rect 4348 9696 4349 9700
rect 4353 9696 4354 9700
rect 4358 9696 4359 9700
rect 4363 9696 4370 9700
rect 4374 9696 4375 9700
rect 4379 9696 4380 9700
rect 4384 9696 4385 9700
rect 4389 9696 4396 9700
rect 4400 9696 4401 9700
rect 4405 9696 4406 9700
rect 4410 9696 4411 9700
rect 4415 9696 4518 9700
rect 654 9695 4518 9696
rect 654 9691 1489 9695
rect 1493 9691 1494 9695
rect 1498 9691 3343 9695
rect 3347 9691 3348 9695
rect 3352 9691 4518 9695
rect 654 9690 4518 9691
rect 654 9686 802 9690
rect 806 9686 807 9690
rect 811 9686 812 9690
rect 816 9686 817 9690
rect 821 9686 831 9690
rect 835 9686 836 9690
rect 840 9686 841 9690
rect 845 9686 846 9690
rect 850 9686 860 9690
rect 864 9686 865 9690
rect 869 9686 870 9690
rect 874 9686 875 9690
rect 879 9686 889 9690
rect 893 9686 894 9690
rect 898 9686 899 9690
rect 903 9686 904 9690
rect 908 9686 918 9690
rect 922 9686 923 9690
rect 927 9686 928 9690
rect 932 9686 933 9690
rect 937 9686 1319 9690
rect 1323 9686 1324 9690
rect 1328 9686 1329 9690
rect 1333 9686 1334 9690
rect 1338 9686 1489 9690
rect 1493 9686 1494 9690
rect 1498 9686 1628 9690
rect 1632 9686 1633 9690
rect 1637 9686 1638 9690
rect 1642 9686 1643 9690
rect 1647 9686 1937 9690
rect 1941 9686 1942 9690
rect 1946 9686 1947 9690
rect 1951 9686 1952 9690
rect 1956 9686 2246 9690
rect 2250 9686 2251 9690
rect 2255 9686 2256 9690
rect 2260 9686 2261 9690
rect 2265 9686 2555 9690
rect 2559 9686 2560 9690
rect 2564 9686 2565 9690
rect 2569 9686 2570 9690
rect 2574 9686 2864 9690
rect 2868 9686 2869 9690
rect 2873 9686 2874 9690
rect 2878 9686 2879 9690
rect 2883 9686 3173 9690
rect 3177 9686 3178 9690
rect 3182 9686 3183 9690
rect 3187 9686 3188 9690
rect 3192 9686 3343 9690
rect 3347 9686 3348 9690
rect 3352 9686 3482 9690
rect 3486 9686 3487 9690
rect 3491 9686 3492 9690
rect 3496 9686 3497 9690
rect 3501 9686 3791 9690
rect 3795 9686 3796 9690
rect 3800 9686 3801 9690
rect 3805 9686 3806 9690
rect 3810 9686 4100 9690
rect 4104 9686 4105 9690
rect 4109 9686 4110 9690
rect 4114 9686 4115 9690
rect 4119 9686 4292 9690
rect 4296 9686 4297 9690
rect 4301 9686 4302 9690
rect 4306 9686 4307 9690
rect 4311 9686 4318 9690
rect 4322 9686 4323 9690
rect 4327 9686 4328 9690
rect 4332 9686 4333 9690
rect 4337 9686 4344 9690
rect 4348 9686 4349 9690
rect 4353 9686 4354 9690
rect 4358 9686 4359 9690
rect 4363 9686 4370 9690
rect 4374 9686 4375 9690
rect 4379 9686 4380 9690
rect 4384 9686 4385 9690
rect 4389 9686 4396 9690
rect 4400 9686 4401 9690
rect 4405 9686 4406 9690
rect 4410 9686 4411 9690
rect 4415 9686 4518 9690
rect 654 9685 4518 9686
rect 654 9681 1489 9685
rect 1493 9681 1494 9685
rect 1498 9681 3343 9685
rect 3347 9681 3348 9685
rect 3352 9681 4518 9685
rect 654 9680 4518 9681
rect 654 9676 1489 9680
rect 1493 9676 1494 9680
rect 1498 9676 3343 9680
rect 3347 9676 3348 9680
rect 3352 9676 4518 9680
rect 654 9675 4518 9676
rect 654 9671 1489 9675
rect 1493 9671 1494 9675
rect 1498 9671 3343 9675
rect 3347 9671 3348 9675
rect 3352 9671 4518 9675
rect 654 9670 4518 9671
rect 654 9666 1489 9670
rect 1493 9666 1494 9670
rect 1498 9666 3343 9670
rect 3347 9666 3348 9670
rect 3352 9666 4518 9670
rect 654 9665 4518 9666
rect 654 9661 1489 9665
rect 1493 9661 1494 9665
rect 1498 9661 3343 9665
rect 3347 9661 3348 9665
rect 3352 9661 4518 9665
rect 654 9623 4518 9661
rect 654 9622 2258 9623
rect 654 9618 659 9622
rect 663 9618 669 9622
rect 673 9618 679 9622
rect 683 9618 689 9622
rect 693 9619 2258 9622
rect 2262 9619 4518 9623
rect 693 9618 4518 9619
rect 654 9617 4518 9618
rect 654 9613 659 9617
rect 663 9613 669 9617
rect 673 9613 679 9617
rect 683 9613 689 9617
rect 693 9613 4518 9617
rect 654 9612 4518 9613
rect 654 9608 659 9612
rect 663 9608 669 9612
rect 673 9608 679 9612
rect 683 9608 689 9612
rect 693 9610 4518 9612
rect 693 9608 769 9610
rect 654 9607 769 9608
rect 654 9603 659 9607
rect 663 9603 669 9607
rect 673 9603 679 9607
rect 683 9603 689 9607
rect 693 9603 769 9607
rect 654 9596 769 9603
rect 654 9592 659 9596
rect 663 9592 669 9596
rect 673 9592 679 9596
rect 683 9592 689 9596
rect 693 9592 769 9596
rect 654 9591 769 9592
rect 654 9587 659 9591
rect 663 9587 669 9591
rect 673 9587 679 9591
rect 683 9587 689 9591
rect 693 9587 769 9591
rect 654 9586 769 9587
rect 654 9582 659 9586
rect 663 9582 669 9586
rect 673 9582 679 9586
rect 683 9582 689 9586
rect 693 9582 769 9586
rect 654 9581 769 9582
rect 654 9577 659 9581
rect 663 9577 669 9581
rect 673 9577 679 9581
rect 683 9577 689 9581
rect 693 9577 769 9581
rect 654 9570 769 9577
rect 654 9566 659 9570
rect 663 9566 669 9570
rect 673 9566 679 9570
rect 683 9566 689 9570
rect 693 9566 769 9570
rect 654 9565 769 9566
rect 654 9561 659 9565
rect 663 9561 669 9565
rect 673 9561 679 9565
rect 683 9561 689 9565
rect 693 9561 769 9565
rect 654 9560 769 9561
rect 654 9556 659 9560
rect 663 9556 669 9560
rect 673 9556 679 9560
rect 683 9556 689 9560
rect 693 9556 769 9560
rect 654 9555 769 9556
rect 654 9551 659 9555
rect 663 9551 669 9555
rect 673 9551 679 9555
rect 683 9551 689 9555
rect 693 9551 769 9555
rect 654 9544 769 9551
rect 654 9540 659 9544
rect 663 9540 669 9544
rect 673 9540 679 9544
rect 683 9540 689 9544
rect 693 9540 769 9544
rect 654 9539 769 9540
rect 654 9535 659 9539
rect 663 9535 669 9539
rect 673 9535 679 9539
rect 683 9535 689 9539
rect 693 9535 769 9539
rect 654 9534 769 9535
rect 654 9530 659 9534
rect 663 9530 669 9534
rect 673 9530 679 9534
rect 683 9530 689 9534
rect 693 9530 769 9534
rect 654 9529 769 9530
rect 654 9525 659 9529
rect 663 9525 669 9529
rect 673 9525 679 9529
rect 683 9525 689 9529
rect 693 9525 769 9529
rect 654 9518 769 9525
rect 654 9514 659 9518
rect 663 9514 669 9518
rect 673 9514 679 9518
rect 683 9514 689 9518
rect 693 9514 769 9518
rect 654 9513 769 9514
rect 654 9509 659 9513
rect 663 9509 669 9513
rect 673 9509 679 9513
rect 683 9509 689 9513
rect 693 9509 769 9513
rect 654 9508 769 9509
rect 654 9504 659 9508
rect 663 9504 669 9508
rect 673 9504 679 9508
rect 683 9504 689 9508
rect 693 9504 769 9508
rect 654 9503 769 9504
rect 654 9499 659 9503
rect 663 9499 669 9503
rect 673 9499 679 9503
rect 683 9499 689 9503
rect 693 9499 769 9503
rect 654 9325 769 9499
rect 654 9321 659 9325
rect 663 9321 669 9325
rect 673 9321 679 9325
rect 683 9321 689 9325
rect 693 9321 769 9325
rect 654 9320 769 9321
rect 654 9316 659 9320
rect 663 9316 669 9320
rect 673 9316 679 9320
rect 683 9316 689 9320
rect 693 9316 769 9320
rect 4403 9577 4518 9610
rect 4403 9573 4479 9577
rect 4483 9573 4489 9577
rect 4493 9573 4499 9577
rect 4503 9573 4509 9577
rect 4513 9573 4518 9577
rect 4403 9572 4518 9573
rect 4403 9568 4479 9572
rect 4483 9568 4489 9572
rect 4493 9568 4499 9572
rect 4503 9568 4509 9572
rect 4513 9568 4518 9572
rect 4403 9567 4518 9568
rect 4403 9563 4479 9567
rect 4483 9563 4489 9567
rect 4493 9563 4499 9567
rect 4503 9563 4509 9567
rect 4513 9563 4518 9567
rect 4403 9562 4518 9563
rect 4403 9558 4479 9562
rect 4483 9558 4489 9562
rect 4493 9558 4499 9562
rect 4503 9558 4509 9562
rect 4513 9558 4518 9562
rect 4403 9548 4518 9558
rect 4403 9544 4479 9548
rect 4483 9544 4489 9548
rect 4493 9544 4499 9548
rect 4503 9544 4509 9548
rect 4513 9544 4518 9548
rect 4403 9543 4518 9544
rect 4403 9539 4479 9543
rect 4483 9539 4489 9543
rect 4493 9539 4499 9543
rect 4503 9539 4509 9543
rect 4513 9539 4518 9543
rect 4403 9538 4518 9539
rect 4403 9534 4479 9538
rect 4483 9534 4489 9538
rect 4493 9534 4499 9538
rect 4503 9534 4509 9538
rect 4513 9534 4518 9538
rect 4403 9533 4518 9534
rect 4403 9529 4479 9533
rect 4483 9529 4489 9533
rect 4493 9529 4499 9533
rect 4503 9529 4509 9533
rect 4513 9529 4518 9533
rect 4403 9519 4518 9529
rect 4403 9515 4479 9519
rect 4483 9515 4489 9519
rect 4493 9515 4499 9519
rect 4503 9515 4509 9519
rect 4513 9515 4518 9519
rect 4403 9514 4518 9515
rect 4403 9510 4479 9514
rect 4483 9510 4489 9514
rect 4493 9510 4499 9514
rect 4503 9510 4509 9514
rect 4513 9510 4518 9514
rect 4403 9509 4518 9510
rect 4403 9505 4479 9509
rect 4483 9505 4489 9509
rect 4493 9505 4499 9509
rect 4503 9505 4509 9509
rect 4513 9505 4518 9509
rect 4403 9504 4518 9505
rect 4403 9500 4479 9504
rect 4483 9500 4489 9504
rect 4493 9500 4499 9504
rect 4503 9500 4509 9504
rect 4513 9500 4518 9504
rect 4403 9490 4518 9500
rect 4403 9486 4479 9490
rect 4483 9486 4489 9490
rect 4493 9486 4499 9490
rect 4503 9486 4509 9490
rect 4513 9486 4518 9490
rect 4403 9485 4518 9486
rect 4403 9481 4479 9485
rect 4483 9481 4489 9485
rect 4493 9481 4499 9485
rect 4503 9481 4509 9485
rect 4513 9481 4518 9485
rect 4403 9480 4518 9481
rect 4403 9476 4479 9480
rect 4483 9476 4489 9480
rect 4493 9476 4499 9480
rect 4503 9476 4509 9480
rect 4513 9476 4518 9480
rect 4403 9475 4518 9476
rect 4403 9471 4479 9475
rect 4483 9471 4489 9475
rect 4493 9471 4499 9475
rect 4503 9471 4509 9475
rect 4513 9471 4518 9475
rect 4403 9461 4518 9471
rect 4403 9457 4479 9461
rect 4483 9457 4489 9461
rect 4493 9457 4499 9461
rect 4503 9457 4509 9461
rect 4513 9457 4518 9461
rect 4403 9456 4518 9457
rect 4403 9452 4479 9456
rect 4483 9452 4489 9456
rect 4493 9452 4499 9456
rect 4503 9452 4509 9456
rect 4513 9452 4518 9456
rect 4403 9451 4518 9452
rect 4403 9447 4479 9451
rect 4483 9447 4489 9451
rect 4493 9447 4499 9451
rect 4503 9447 4509 9451
rect 4513 9447 4518 9451
rect 4403 9446 4518 9447
rect 4403 9442 4479 9446
rect 4483 9442 4489 9446
rect 4493 9442 4499 9446
rect 4503 9442 4509 9446
rect 4513 9442 4518 9446
rect 654 9315 769 9316
rect 654 9311 659 9315
rect 663 9311 669 9315
rect 673 9311 679 9315
rect 683 9311 689 9315
rect 693 9311 769 9315
rect 654 9310 769 9311
rect 654 9306 659 9310
rect 663 9306 669 9310
rect 673 9306 679 9310
rect 683 9306 689 9310
rect 693 9306 769 9310
rect 654 9016 769 9306
rect 2846 9317 2852 9318
rect 2846 9313 2847 9317
rect 2851 9313 2852 9317
rect 2846 9312 2852 9313
rect 3791 9317 3797 9318
rect 3791 9313 3792 9317
rect 3796 9313 3797 9317
rect 3791 9312 3797 9313
rect 2846 9282 2851 9312
rect 3791 9282 3796 9312
rect 2623 9281 2851 9282
rect 2623 9277 2624 9281
rect 2628 9277 2851 9281
rect 3568 9281 3796 9282
rect 3568 9277 3569 9281
rect 3573 9277 3796 9281
rect 2623 9276 2629 9277
rect 3568 9276 3574 9277
rect 3302 9266 3308 9267
rect 3302 9262 3303 9266
rect 3307 9262 3308 9266
rect 3302 9261 3308 9262
rect 4247 9266 4253 9267
rect 4247 9262 4248 9266
rect 4252 9262 4253 9266
rect 4247 9261 4253 9262
rect 2887 9240 2927 9241
rect 2887 9236 2921 9240
rect 2886 9235 2893 9236
rect 2886 9230 2887 9235
rect 2892 9230 2893 9235
rect 2920 9235 2921 9236
rect 2926 9235 2927 9240
rect 2959 9240 2995 9245
rect 2920 9234 2927 9235
rect 2944 9235 2951 9236
rect 2886 9229 2893 9230
rect 2897 9231 2904 9232
rect 2897 9226 2898 9231
rect 2903 9226 2904 9231
rect 2944 9230 2945 9235
rect 2950 9230 2951 9235
rect 2959 9234 2960 9240
rect 2965 9239 2995 9240
rect 2965 9234 2966 9239
rect 2990 9236 2995 9239
rect 2959 9233 2966 9234
rect 2989 9235 2996 9236
rect 2989 9230 2990 9235
rect 2995 9230 2996 9235
rect 3018 9234 3025 9235
rect 2944 9229 2951 9230
rect 2973 9229 2980 9230
rect 2989 9229 2996 9230
rect 3002 9229 3008 9230
rect 2945 9226 2950 9229
rect 2897 9221 2950 9226
rect 2973 9224 2974 9229
rect 2979 9224 2980 9229
rect 3002 9224 3003 9229
rect 3007 9224 3008 9229
rect 2973 9223 3008 9224
rect 2974 9219 3008 9223
rect 3018 9229 3019 9234
rect 3024 9229 3025 9234
rect 3100 9234 3107 9235
rect 3100 9229 3101 9234
rect 3106 9229 3107 9234
rect 3185 9234 3192 9235
rect 3185 9229 3186 9234
rect 3191 9229 3192 9234
rect 3018 9228 3025 9229
rect 3044 9228 3051 9229
rect 3100 9228 3107 9229
rect 3125 9228 3132 9229
rect 3185 9228 3192 9229
rect 3018 9223 3045 9228
rect 3050 9223 3051 9228
rect 3101 9223 3126 9228
rect 3131 9223 3132 9228
rect 3018 9202 3023 9223
rect 3044 9222 3051 9223
rect 3125 9222 3132 9223
rect 3182 9223 3191 9228
rect 2851 9196 3023 9202
rect 2622 9178 2628 9179
rect 2622 9174 2623 9178
rect 2627 9174 2760 9178
rect 2851 9176 2856 9196
rect 2622 9173 2760 9174
rect 654 9012 659 9016
rect 663 9012 669 9016
rect 673 9012 679 9016
rect 683 9012 689 9016
rect 693 9012 769 9016
rect 654 9011 769 9012
rect 654 9007 659 9011
rect 663 9007 669 9011
rect 673 9007 679 9011
rect 683 9007 689 9011
rect 693 9007 769 9011
rect 654 9006 769 9007
rect 654 9002 659 9006
rect 663 9002 669 9006
rect 673 9002 679 9006
rect 683 9002 689 9006
rect 693 9002 769 9006
rect 654 9001 769 9002
rect 654 8997 659 9001
rect 663 8997 669 9001
rect 673 8997 679 9001
rect 683 8997 689 9001
rect 693 8997 769 9001
rect 654 8707 769 8997
rect 2366 8778 2372 8779
rect 2366 8774 2367 8778
rect 2371 8774 2372 8778
rect 2366 8773 2372 8774
rect 654 8703 659 8707
rect 663 8703 669 8707
rect 673 8703 679 8707
rect 683 8703 689 8707
rect 693 8703 769 8707
rect 654 8702 769 8703
rect 654 8698 659 8702
rect 663 8698 669 8702
rect 673 8698 679 8702
rect 683 8698 689 8702
rect 693 8698 769 8702
rect 654 8697 769 8698
rect 654 8693 659 8697
rect 663 8693 669 8697
rect 673 8693 679 8697
rect 683 8693 689 8697
rect 693 8693 769 8697
rect 654 8692 769 8693
rect 654 8688 659 8692
rect 663 8688 669 8692
rect 673 8688 679 8692
rect 683 8688 689 8692
rect 693 8688 769 8692
rect 654 8398 769 8688
rect 2755 8412 2760 9173
rect 2850 9175 2857 9176
rect 2850 9170 2851 9175
rect 2856 9170 2857 9175
rect 2850 9169 2857 9170
rect 2897 9172 2950 9177
rect 2974 9175 3008 9179
rect 2886 9168 2893 9169
rect 2886 9163 2887 9168
rect 2892 9163 2893 9168
rect 2897 9167 2898 9172
rect 2903 9167 2904 9172
rect 2945 9169 2950 9172
rect 2973 9174 3008 9175
rect 2973 9169 2974 9174
rect 2979 9169 2980 9174
rect 3002 9169 3003 9174
rect 3007 9169 3008 9174
rect 2897 9166 2904 9167
rect 2944 9168 2951 9169
rect 2973 9168 2980 9169
rect 2989 9168 2996 9169
rect 3002 9168 3008 9169
rect 3018 9169 3025 9170
rect 3044 9169 3051 9170
rect 3124 9169 3131 9170
rect 2886 9162 2893 9163
rect 2920 9163 2927 9164
rect 2920 9162 2921 9163
rect 2887 9158 2921 9162
rect 2926 9158 2927 9163
rect 2944 9163 2945 9168
rect 2950 9163 2951 9168
rect 2944 9162 2951 9163
rect 2959 9164 2966 9165
rect 2887 9157 2927 9158
rect 2959 9158 2960 9164
rect 2965 9159 2966 9164
rect 2989 9163 2990 9168
rect 2995 9163 2996 9168
rect 3018 9164 3019 9169
rect 3024 9164 3045 9169
rect 3050 9164 3051 9169
rect 3018 9163 3025 9164
rect 3044 9163 3051 9164
rect 3101 9164 3125 9169
rect 3130 9164 3131 9169
rect 2989 9162 2996 9163
rect 2990 9159 2995 9162
rect 2965 9158 2995 9159
rect 2959 9153 2995 9158
rect 3019 9136 3024 9163
rect 2850 9130 3024 9136
rect 2850 9107 2855 9130
rect 2887 9108 2927 9109
rect 2849 9106 2856 9107
rect 2849 9101 2850 9106
rect 2855 9101 2856 9106
rect 2887 9104 2921 9108
rect 2849 9100 2856 9101
rect 2886 9103 2893 9104
rect 2886 9098 2887 9103
rect 2892 9098 2893 9103
rect 2920 9103 2921 9104
rect 2926 9103 2927 9108
rect 2959 9108 2995 9113
rect 3101 9111 3106 9164
rect 3124 9163 3131 9164
rect 3182 9135 3187 9223
rect 3144 9130 3187 9135
rect 2920 9102 2927 9103
rect 2944 9103 2951 9104
rect 2886 9097 2893 9098
rect 2897 9099 2904 9100
rect 2897 9094 2898 9099
rect 2903 9094 2904 9099
rect 2944 9098 2945 9103
rect 2950 9098 2951 9103
rect 2959 9102 2960 9108
rect 2965 9107 2995 9108
rect 2965 9102 2966 9107
rect 2990 9104 2995 9107
rect 3100 9110 3107 9111
rect 3100 9105 3101 9110
rect 3106 9105 3107 9110
rect 3100 9104 3107 9105
rect 2959 9101 2966 9102
rect 2989 9103 2996 9104
rect 2989 9098 2990 9103
rect 2995 9098 2996 9103
rect 3018 9102 3025 9103
rect 2944 9097 2951 9098
rect 2973 9097 2980 9098
rect 2989 9097 2996 9098
rect 3002 9097 3008 9098
rect 2945 9094 2950 9097
rect 2897 9089 2950 9094
rect 2973 9092 2974 9097
rect 2979 9092 2980 9097
rect 3002 9092 3003 9097
rect 3007 9092 3008 9097
rect 2973 9091 3008 9092
rect 2974 9087 3008 9091
rect 3018 9097 3019 9102
rect 3024 9097 3025 9102
rect 3144 9097 3149 9130
rect 3207 9107 3214 9108
rect 3207 9102 3208 9107
rect 3213 9102 3214 9107
rect 3207 9101 3214 9102
rect 3018 9096 3025 9097
rect 3044 9096 3051 9097
rect 3018 9091 3045 9096
rect 3050 9091 3051 9096
rect 3144 9096 3156 9097
rect 3144 9091 3150 9096
rect 3155 9091 3156 9096
rect 3018 9070 3023 9091
rect 3044 9090 3051 9091
rect 3149 9090 3156 9091
rect 2851 9064 3023 9070
rect 2851 9044 2856 9064
rect 2850 9043 2857 9044
rect 2850 9038 2851 9043
rect 2856 9038 2857 9043
rect 2850 9037 2857 9038
rect 2897 9040 2950 9045
rect 2974 9043 3008 9047
rect 2886 9036 2893 9037
rect 2886 9031 2887 9036
rect 2892 9031 2893 9036
rect 2897 9035 2898 9040
rect 2903 9035 2904 9040
rect 2945 9037 2950 9040
rect 2973 9042 3008 9043
rect 2973 9037 2974 9042
rect 2979 9037 2980 9042
rect 3002 9037 3003 9042
rect 3007 9037 3008 9042
rect 3043 9038 3050 9039
rect 3149 9038 3156 9039
rect 2897 9034 2904 9035
rect 2944 9036 2951 9037
rect 2973 9036 2980 9037
rect 2989 9036 2996 9037
rect 3002 9036 3008 9037
rect 3018 9037 3044 9038
rect 2886 9030 2893 9031
rect 2920 9031 2927 9032
rect 2920 9030 2921 9031
rect 2887 9026 2921 9030
rect 2926 9026 2927 9031
rect 2944 9031 2945 9036
rect 2950 9031 2951 9036
rect 2944 9030 2951 9031
rect 2959 9032 2966 9033
rect 2887 9025 2927 9026
rect 2959 9026 2960 9032
rect 2965 9027 2966 9032
rect 2989 9031 2990 9036
rect 2995 9031 2996 9036
rect 2989 9030 2996 9031
rect 3018 9032 3019 9037
rect 3024 9033 3044 9037
rect 3049 9033 3050 9038
rect 3024 9032 3025 9033
rect 3043 9032 3050 9033
rect 3145 9033 3150 9038
rect 3155 9033 3156 9038
rect 3145 9032 3156 9033
rect 3018 9031 3025 9032
rect 2990 9027 2995 9030
rect 2965 9026 2995 9027
rect 2959 9021 2995 9026
rect 3018 9004 3023 9031
rect 2850 8998 3023 9004
rect 3145 9004 3150 9032
rect 3145 8999 3188 9004
rect 2850 8975 2855 8998
rect 2887 8976 2927 8977
rect 2849 8974 2856 8975
rect 2849 8969 2850 8974
rect 2855 8969 2856 8974
rect 2887 8972 2921 8976
rect 2849 8968 2856 8969
rect 2886 8971 2893 8972
rect 2886 8966 2887 8971
rect 2892 8966 2893 8971
rect 2920 8971 2921 8972
rect 2926 8971 2927 8976
rect 2959 8976 2995 8981
rect 3183 8980 3188 8999
rect 2920 8970 2927 8971
rect 2944 8971 2951 8972
rect 2886 8965 2893 8966
rect 2897 8967 2904 8968
rect 2897 8962 2898 8967
rect 2903 8962 2904 8967
rect 2944 8966 2945 8971
rect 2950 8966 2951 8971
rect 2959 8970 2960 8976
rect 2965 8975 2995 8976
rect 2965 8970 2966 8975
rect 2990 8972 2995 8975
rect 3182 8979 3189 8980
rect 3182 8974 3183 8979
rect 3188 8974 3189 8979
rect 3182 8973 3189 8974
rect 3208 8972 3213 9101
rect 3216 8972 3223 8973
rect 2959 8969 2966 8970
rect 2989 8971 2996 8972
rect 2989 8966 2990 8971
rect 2995 8966 2996 8971
rect 3018 8970 3025 8971
rect 2944 8965 2951 8966
rect 2973 8965 2980 8966
rect 2989 8965 2996 8966
rect 3002 8965 3008 8966
rect 2945 8962 2950 8965
rect 2897 8957 2950 8962
rect 2973 8960 2974 8965
rect 2979 8960 2980 8965
rect 3002 8960 3003 8965
rect 3007 8960 3008 8965
rect 2973 8959 3008 8960
rect 2974 8955 3008 8959
rect 3018 8965 3019 8970
rect 3024 8965 3025 8970
rect 3100 8970 3107 8971
rect 3100 8965 3101 8970
rect 3106 8965 3107 8970
rect 3196 8967 3217 8972
rect 3222 8967 3223 8972
rect 3196 8966 3208 8967
rect 3216 8966 3223 8967
rect 3018 8964 3025 8965
rect 3044 8964 3051 8965
rect 3100 8964 3107 8965
rect 3125 8964 3132 8965
rect 3018 8959 3045 8964
rect 3050 8959 3051 8964
rect 3101 8959 3126 8964
rect 3131 8959 3132 8964
rect 3018 8938 3023 8959
rect 3044 8958 3051 8959
rect 3125 8958 3132 8959
rect 3196 8958 3201 8966
rect 2851 8932 3023 8938
rect 3163 8937 3201 8958
rect 2851 8912 2856 8932
rect 2850 8911 2857 8912
rect 2850 8906 2851 8911
rect 2856 8906 2857 8911
rect 2850 8905 2857 8906
rect 2897 8908 2950 8913
rect 2974 8911 3008 8915
rect 2886 8904 2893 8905
rect 2886 8899 2887 8904
rect 2892 8899 2893 8904
rect 2897 8903 2898 8908
rect 2903 8903 2904 8908
rect 2945 8905 2950 8908
rect 2973 8910 3008 8911
rect 2973 8905 2974 8910
rect 2979 8905 2980 8910
rect 3002 8905 3003 8910
rect 3007 8905 3008 8910
rect 2897 8902 2904 8903
rect 2944 8904 2951 8905
rect 2973 8904 2980 8905
rect 2989 8904 2996 8905
rect 3002 8904 3008 8905
rect 3018 8905 3025 8906
rect 2886 8898 2893 8899
rect 2920 8899 2927 8900
rect 2920 8898 2921 8899
rect 2887 8894 2921 8898
rect 2926 8894 2927 8899
rect 2944 8899 2945 8904
rect 2950 8899 2951 8904
rect 2944 8898 2951 8899
rect 2959 8900 2966 8901
rect 2887 8893 2927 8894
rect 2959 8894 2960 8900
rect 2965 8895 2966 8900
rect 2989 8899 2990 8904
rect 2995 8899 2996 8904
rect 3018 8900 3019 8905
rect 3024 8903 3025 8905
rect 3044 8903 3051 8904
rect 3124 8903 3131 8904
rect 3024 8900 3045 8903
rect 3018 8899 3045 8900
rect 2989 8898 2996 8899
rect 3019 8898 3045 8899
rect 3050 8898 3051 8903
rect 2990 8895 2995 8898
rect 2965 8894 2995 8895
rect 2959 8889 2995 8894
rect 3019 8872 3024 8898
rect 3044 8897 3051 8898
rect 3101 8898 3125 8903
rect 3130 8898 3131 8903
rect 2850 8866 3024 8872
rect 2850 8843 2855 8866
rect 2887 8844 2927 8845
rect 2849 8842 2856 8843
rect 2849 8837 2850 8842
rect 2855 8837 2856 8842
rect 2887 8840 2921 8844
rect 2849 8836 2856 8837
rect 2886 8839 2893 8840
rect 2886 8834 2887 8839
rect 2892 8834 2893 8839
rect 2920 8839 2921 8840
rect 2926 8839 2927 8844
rect 2959 8844 2995 8849
rect 3101 8847 3106 8898
rect 3124 8897 3131 8898
rect 2920 8838 2927 8839
rect 2944 8839 2951 8840
rect 2886 8833 2893 8834
rect 2897 8835 2904 8836
rect 2897 8830 2898 8835
rect 2903 8830 2904 8835
rect 2944 8834 2945 8839
rect 2950 8834 2951 8839
rect 2959 8838 2960 8844
rect 2965 8843 2995 8844
rect 2965 8838 2966 8843
rect 2990 8840 2995 8843
rect 3100 8846 3107 8847
rect 3100 8841 3101 8846
rect 3106 8841 3107 8846
rect 3100 8840 3107 8841
rect 2959 8837 2966 8838
rect 2989 8839 2996 8840
rect 2989 8834 2990 8839
rect 2995 8834 2996 8839
rect 3018 8838 3025 8839
rect 2944 8833 2951 8834
rect 2973 8833 2980 8834
rect 2989 8833 2996 8834
rect 3002 8833 3008 8834
rect 2945 8830 2950 8833
rect 2897 8825 2950 8830
rect 2973 8828 2974 8833
rect 2979 8828 2980 8833
rect 3002 8828 3003 8833
rect 3007 8828 3008 8833
rect 2973 8827 3008 8828
rect 2974 8823 3008 8827
rect 3018 8833 3019 8838
rect 3024 8833 3025 8838
rect 3018 8832 3025 8833
rect 3044 8832 3051 8833
rect 3018 8827 3045 8832
rect 3050 8827 3051 8832
rect 3163 8828 3168 8937
rect 3213 8899 3220 8900
rect 3213 8894 3214 8899
rect 3219 8894 3220 8899
rect 3213 8893 3220 8894
rect 3120 8827 3168 8828
rect 3018 8806 3023 8827
rect 3044 8826 3051 8827
rect 2851 8800 3023 8806
rect 3089 8822 3168 8827
rect 3214 8831 3219 8893
rect 3214 8825 3281 8831
rect 2851 8780 2856 8800
rect 2850 8779 2857 8780
rect 2850 8774 2851 8779
rect 2856 8774 2857 8779
rect 2850 8773 2857 8774
rect 2897 8776 2950 8781
rect 2974 8779 3008 8783
rect 3089 8779 3094 8822
rect 2886 8772 2893 8773
rect 2886 8767 2887 8772
rect 2892 8767 2893 8772
rect 2897 8771 2898 8776
rect 2903 8771 2904 8776
rect 2945 8773 2950 8776
rect 2973 8778 3008 8779
rect 2973 8773 2974 8778
rect 2979 8773 2980 8778
rect 3002 8773 3003 8778
rect 3007 8773 3008 8778
rect 3088 8778 3095 8779
rect 2897 8770 2904 8771
rect 2944 8772 2951 8773
rect 2973 8772 2980 8773
rect 2989 8772 2996 8773
rect 3002 8772 3008 8773
rect 3018 8773 3025 8774
rect 2886 8766 2893 8767
rect 2920 8767 2927 8768
rect 2920 8766 2921 8767
rect 2887 8762 2921 8766
rect 2926 8762 2927 8767
rect 2944 8767 2945 8772
rect 2950 8767 2951 8772
rect 2944 8766 2951 8767
rect 2959 8768 2966 8769
rect 2887 8761 2927 8762
rect 2959 8762 2960 8768
rect 2965 8763 2966 8768
rect 2989 8767 2990 8772
rect 2995 8767 2996 8772
rect 3018 8768 3019 8773
rect 3024 8768 3025 8773
rect 3088 8773 3089 8778
rect 3094 8773 3095 8778
rect 3158 8776 3211 8781
rect 3235 8779 3269 8783
rect 3276 8779 3281 8825
rect 3088 8772 3095 8773
rect 3147 8772 3154 8773
rect 3018 8767 3025 8768
rect 3043 8767 3050 8768
rect 2989 8766 2996 8767
rect 2990 8763 2995 8766
rect 2965 8762 2995 8763
rect 2959 8757 2995 8762
rect 3020 8762 3044 8767
rect 3049 8762 3050 8767
rect 3147 8767 3148 8772
rect 3153 8767 3154 8772
rect 3158 8771 3159 8776
rect 3164 8771 3165 8776
rect 3206 8773 3211 8776
rect 3234 8778 3269 8779
rect 3234 8773 3235 8778
rect 3240 8773 3241 8778
rect 3263 8773 3264 8778
rect 3268 8773 3269 8778
rect 3158 8770 3165 8771
rect 3205 8772 3212 8773
rect 3234 8772 3241 8773
rect 3250 8772 3257 8773
rect 3263 8772 3269 8773
rect 3275 8778 3282 8779
rect 3275 8773 3276 8778
rect 3281 8773 3282 8778
rect 3275 8772 3282 8773
rect 3147 8766 3154 8767
rect 3181 8767 3188 8768
rect 3181 8766 3182 8767
rect 2755 8411 2761 8412
rect 2755 8407 2756 8411
rect 2760 8407 2761 8411
rect 2755 8406 2761 8407
rect 654 8394 659 8398
rect 663 8394 669 8398
rect 673 8394 679 8398
rect 683 8394 689 8398
rect 693 8394 769 8398
rect 654 8393 769 8394
rect 654 8389 659 8393
rect 663 8389 669 8393
rect 673 8389 679 8393
rect 683 8389 689 8393
rect 693 8389 769 8393
rect 654 8388 769 8389
rect 3020 8394 3025 8762
rect 3043 8761 3050 8762
rect 3148 8762 3182 8766
rect 3187 8762 3188 8767
rect 3205 8767 3206 8772
rect 3211 8767 3212 8772
rect 3205 8766 3212 8767
rect 3220 8768 3227 8769
rect 3148 8761 3188 8762
rect 3220 8762 3221 8768
rect 3226 8763 3227 8768
rect 3250 8767 3251 8772
rect 3256 8767 3257 8772
rect 3250 8766 3257 8767
rect 3251 8763 3256 8766
rect 3226 8762 3256 8763
rect 3220 8757 3256 8762
rect 3303 8734 3308 9261
rect 3832 9240 3872 9241
rect 3792 9238 3799 9239
rect 3770 9233 3793 9238
rect 3798 9233 3799 9238
rect 3832 9236 3866 9240
rect 3567 9178 3573 9179
rect 3567 9174 3568 9178
rect 3572 9174 3705 9178
rect 3567 9173 3705 9174
rect 3559 9141 3566 9142
rect 3442 9140 3449 9141
rect 3442 9135 3443 9140
rect 3448 9135 3449 9140
rect 3559 9136 3560 9141
rect 3565 9136 3566 9141
rect 3559 9135 3566 9136
rect 3442 9134 3449 9135
rect 3443 8825 3448 9134
rect 3442 8824 3449 8825
rect 3560 8824 3565 9135
rect 3442 8819 3443 8824
rect 3448 8819 3449 8824
rect 3442 8818 3449 8819
rect 3559 8823 3566 8824
rect 3559 8818 3560 8823
rect 3565 8818 3566 8823
rect 3559 8817 3566 8818
rect 3311 8778 3317 8779
rect 3311 8774 3312 8778
rect 3316 8774 3317 8778
rect 3311 8773 3317 8774
rect 3150 8729 3308 8734
rect 3150 8667 3155 8729
rect 3149 8666 3155 8667
rect 3149 8662 3150 8666
rect 3154 8662 3155 8666
rect 3149 8661 3155 8662
rect 3312 8604 3317 8773
rect 3275 8599 3317 8604
rect 3275 8585 3280 8599
rect 3274 8584 3280 8585
rect 3274 8580 3275 8584
rect 3279 8580 3280 8584
rect 3274 8579 3280 8580
rect 3700 8412 3705 9173
rect 3700 8411 3706 8412
rect 3700 8407 3701 8411
rect 3705 8407 3706 8411
rect 3700 8406 3706 8407
rect 3770 8394 3775 9233
rect 3792 9232 3799 9233
rect 3831 9235 3838 9236
rect 3831 9230 3832 9235
rect 3837 9230 3838 9235
rect 3865 9235 3866 9236
rect 3871 9235 3872 9240
rect 3904 9240 3940 9245
rect 3865 9234 3872 9235
rect 3889 9235 3896 9236
rect 3831 9229 3838 9230
rect 3842 9231 3849 9232
rect 3842 9226 3843 9231
rect 3848 9226 3849 9231
rect 3889 9230 3890 9235
rect 3895 9230 3896 9235
rect 3904 9234 3905 9240
rect 3910 9239 3940 9240
rect 3910 9234 3911 9239
rect 3935 9236 3940 9239
rect 3904 9233 3911 9234
rect 3934 9235 3941 9236
rect 3934 9230 3935 9235
rect 3940 9230 3941 9235
rect 3963 9234 3970 9235
rect 3889 9229 3896 9230
rect 3918 9229 3925 9230
rect 3934 9229 3941 9230
rect 3947 9229 3953 9230
rect 3890 9226 3895 9229
rect 3842 9221 3895 9226
rect 3918 9224 3919 9229
rect 3924 9224 3925 9229
rect 3947 9224 3948 9229
rect 3952 9224 3953 9229
rect 3918 9223 3953 9224
rect 3919 9219 3953 9223
rect 3963 9229 3964 9234
rect 3969 9229 3970 9234
rect 4045 9234 4052 9235
rect 4045 9229 4046 9234
rect 4051 9229 4052 9234
rect 4130 9234 4137 9235
rect 4130 9229 4131 9234
rect 4136 9229 4137 9234
rect 3963 9228 3970 9229
rect 3989 9228 3996 9229
rect 4045 9228 4052 9229
rect 4070 9228 4077 9229
rect 4130 9228 4137 9229
rect 3963 9223 3990 9228
rect 3995 9223 3996 9228
rect 4046 9223 4071 9228
rect 4076 9223 4077 9228
rect 3963 9202 3968 9223
rect 3989 9222 3996 9223
rect 4070 9222 4077 9223
rect 4127 9223 4136 9228
rect 3796 9196 3968 9202
rect 3796 9176 3801 9196
rect 3795 9175 3802 9176
rect 3795 9170 3796 9175
rect 3801 9170 3802 9175
rect 3795 9169 3802 9170
rect 3842 9172 3895 9177
rect 3919 9175 3953 9179
rect 3831 9168 3838 9169
rect 3831 9163 3832 9168
rect 3837 9163 3838 9168
rect 3842 9167 3843 9172
rect 3848 9167 3849 9172
rect 3890 9169 3895 9172
rect 3918 9174 3953 9175
rect 3918 9169 3919 9174
rect 3924 9169 3925 9174
rect 3947 9169 3948 9174
rect 3952 9169 3953 9174
rect 3842 9166 3849 9167
rect 3889 9168 3896 9169
rect 3918 9168 3925 9169
rect 3934 9168 3941 9169
rect 3947 9168 3953 9169
rect 3963 9169 3970 9170
rect 3989 9169 3996 9170
rect 4069 9169 4076 9170
rect 3831 9162 3838 9163
rect 3865 9163 3872 9164
rect 3865 9162 3866 9163
rect 3832 9158 3866 9162
rect 3871 9158 3872 9163
rect 3889 9163 3890 9168
rect 3895 9163 3896 9168
rect 3889 9162 3896 9163
rect 3904 9164 3911 9165
rect 3832 9157 3872 9158
rect 3904 9158 3905 9164
rect 3910 9159 3911 9164
rect 3934 9163 3935 9168
rect 3940 9163 3941 9168
rect 3963 9164 3964 9169
rect 3969 9164 3990 9169
rect 3995 9164 3996 9169
rect 3963 9163 3970 9164
rect 3989 9163 3996 9164
rect 4046 9164 4070 9169
rect 4075 9164 4076 9169
rect 3934 9162 3941 9163
rect 3935 9159 3940 9162
rect 3910 9158 3940 9159
rect 3904 9153 3940 9158
rect 3964 9136 3969 9163
rect 3795 9130 3969 9136
rect 3795 9107 3800 9130
rect 3832 9108 3872 9109
rect 3794 9106 3801 9107
rect 3794 9101 3795 9106
rect 3800 9101 3801 9106
rect 3832 9104 3866 9108
rect 3794 9100 3801 9101
rect 3831 9103 3838 9104
rect 3831 9098 3832 9103
rect 3837 9098 3838 9103
rect 3865 9103 3866 9104
rect 3871 9103 3872 9108
rect 3904 9108 3940 9113
rect 4046 9111 4051 9164
rect 4069 9163 4076 9164
rect 4127 9135 4132 9223
rect 4089 9130 4132 9135
rect 3865 9102 3872 9103
rect 3889 9103 3896 9104
rect 3831 9097 3838 9098
rect 3842 9099 3849 9100
rect 3842 9094 3843 9099
rect 3848 9094 3849 9099
rect 3889 9098 3890 9103
rect 3895 9098 3896 9103
rect 3904 9102 3905 9108
rect 3910 9107 3940 9108
rect 3910 9102 3911 9107
rect 3935 9104 3940 9107
rect 4045 9110 4052 9111
rect 4045 9105 4046 9110
rect 4051 9105 4052 9110
rect 4045 9104 4052 9105
rect 3904 9101 3911 9102
rect 3934 9103 3941 9104
rect 3934 9098 3935 9103
rect 3940 9098 3941 9103
rect 3963 9102 3970 9103
rect 3889 9097 3896 9098
rect 3918 9097 3925 9098
rect 3934 9097 3941 9098
rect 3947 9097 3953 9098
rect 3890 9094 3895 9097
rect 3842 9089 3895 9094
rect 3918 9092 3919 9097
rect 3924 9092 3925 9097
rect 3947 9092 3948 9097
rect 3952 9092 3953 9097
rect 3918 9091 3953 9092
rect 3919 9087 3953 9091
rect 3963 9097 3964 9102
rect 3969 9097 3970 9102
rect 4089 9097 4094 9130
rect 4152 9107 4159 9108
rect 4152 9102 4153 9107
rect 4158 9102 4159 9107
rect 4152 9101 4159 9102
rect 3963 9096 3970 9097
rect 3989 9096 3996 9097
rect 3963 9091 3990 9096
rect 3995 9091 3996 9096
rect 4089 9096 4101 9097
rect 4089 9091 4095 9096
rect 4100 9091 4101 9096
rect 3963 9070 3968 9091
rect 3989 9090 3996 9091
rect 4094 9090 4101 9091
rect 3796 9064 3968 9070
rect 3796 9044 3801 9064
rect 3795 9043 3802 9044
rect 3795 9038 3796 9043
rect 3801 9038 3802 9043
rect 3795 9037 3802 9038
rect 3842 9040 3895 9045
rect 3919 9043 3953 9047
rect 3831 9036 3838 9037
rect 3831 9031 3832 9036
rect 3837 9031 3838 9036
rect 3842 9035 3843 9040
rect 3848 9035 3849 9040
rect 3890 9037 3895 9040
rect 3918 9042 3953 9043
rect 3918 9037 3919 9042
rect 3924 9037 3925 9042
rect 3947 9037 3948 9042
rect 3952 9037 3953 9042
rect 3988 9038 3995 9039
rect 4094 9038 4101 9039
rect 3842 9034 3849 9035
rect 3889 9036 3896 9037
rect 3918 9036 3925 9037
rect 3934 9036 3941 9037
rect 3947 9036 3953 9037
rect 3963 9037 3989 9038
rect 3831 9030 3838 9031
rect 3865 9031 3872 9032
rect 3865 9030 3866 9031
rect 3832 9026 3866 9030
rect 3871 9026 3872 9031
rect 3889 9031 3890 9036
rect 3895 9031 3896 9036
rect 3889 9030 3896 9031
rect 3904 9032 3911 9033
rect 3832 9025 3872 9026
rect 3904 9026 3905 9032
rect 3910 9027 3911 9032
rect 3934 9031 3935 9036
rect 3940 9031 3941 9036
rect 3934 9030 3941 9031
rect 3963 9032 3964 9037
rect 3969 9033 3989 9037
rect 3994 9033 3995 9038
rect 3969 9032 3970 9033
rect 3988 9032 3995 9033
rect 4090 9033 4095 9038
rect 4100 9033 4101 9038
rect 4090 9032 4101 9033
rect 3963 9031 3970 9032
rect 3935 9027 3940 9030
rect 3910 9026 3940 9027
rect 3904 9021 3940 9026
rect 3963 9004 3968 9031
rect 3795 8998 3968 9004
rect 4090 9004 4095 9032
rect 4090 8999 4133 9004
rect 3795 8975 3800 8998
rect 3832 8976 3872 8977
rect 3794 8974 3801 8975
rect 3794 8969 3795 8974
rect 3800 8969 3801 8974
rect 3832 8972 3866 8976
rect 3794 8968 3801 8969
rect 3831 8971 3838 8972
rect 3831 8966 3832 8971
rect 3837 8966 3838 8971
rect 3865 8971 3866 8972
rect 3871 8971 3872 8976
rect 3904 8976 3940 8981
rect 4128 8980 4133 8999
rect 3865 8970 3872 8971
rect 3889 8971 3896 8972
rect 3831 8965 3838 8966
rect 3842 8967 3849 8968
rect 3842 8962 3843 8967
rect 3848 8962 3849 8967
rect 3889 8966 3890 8971
rect 3895 8966 3896 8971
rect 3904 8970 3905 8976
rect 3910 8975 3940 8976
rect 3910 8970 3911 8975
rect 3935 8972 3940 8975
rect 4127 8979 4134 8980
rect 4127 8974 4128 8979
rect 4133 8974 4134 8979
rect 4127 8973 4134 8974
rect 4153 8972 4158 9101
rect 4161 8972 4168 8973
rect 3904 8969 3911 8970
rect 3934 8971 3941 8972
rect 3934 8966 3935 8971
rect 3940 8966 3941 8971
rect 3963 8970 3970 8971
rect 3889 8965 3896 8966
rect 3918 8965 3925 8966
rect 3934 8965 3941 8966
rect 3947 8965 3953 8966
rect 3890 8962 3895 8965
rect 3842 8957 3895 8962
rect 3918 8960 3919 8965
rect 3924 8960 3925 8965
rect 3947 8960 3948 8965
rect 3952 8960 3953 8965
rect 3918 8959 3953 8960
rect 3919 8955 3953 8959
rect 3963 8965 3964 8970
rect 3969 8965 3970 8970
rect 4045 8970 4052 8971
rect 4045 8965 4046 8970
rect 4051 8965 4052 8970
rect 4141 8967 4162 8972
rect 4167 8967 4168 8972
rect 4141 8966 4153 8967
rect 4161 8966 4168 8967
rect 3963 8964 3970 8965
rect 3989 8964 3996 8965
rect 4045 8964 4052 8965
rect 4070 8964 4077 8965
rect 3963 8959 3990 8964
rect 3995 8959 3996 8964
rect 4046 8959 4071 8964
rect 4076 8959 4077 8964
rect 3963 8938 3968 8959
rect 3989 8958 3996 8959
rect 4070 8958 4077 8959
rect 4141 8958 4146 8966
rect 3796 8932 3968 8938
rect 4108 8937 4146 8958
rect 3796 8912 3801 8932
rect 3795 8911 3802 8912
rect 3795 8906 3796 8911
rect 3801 8906 3802 8911
rect 3795 8905 3802 8906
rect 3842 8908 3895 8913
rect 3919 8911 3953 8915
rect 3831 8904 3838 8905
rect 3831 8899 3832 8904
rect 3837 8899 3838 8904
rect 3842 8903 3843 8908
rect 3848 8903 3849 8908
rect 3890 8905 3895 8908
rect 3918 8910 3953 8911
rect 3918 8905 3919 8910
rect 3924 8905 3925 8910
rect 3947 8905 3948 8910
rect 3952 8905 3953 8910
rect 3842 8902 3849 8903
rect 3889 8904 3896 8905
rect 3918 8904 3925 8905
rect 3934 8904 3941 8905
rect 3947 8904 3953 8905
rect 3963 8905 3970 8906
rect 3831 8898 3838 8899
rect 3865 8899 3872 8900
rect 3865 8898 3866 8899
rect 3832 8894 3866 8898
rect 3871 8894 3872 8899
rect 3889 8899 3890 8904
rect 3895 8899 3896 8904
rect 3889 8898 3896 8899
rect 3904 8900 3911 8901
rect 3832 8893 3872 8894
rect 3904 8894 3905 8900
rect 3910 8895 3911 8900
rect 3934 8899 3935 8904
rect 3940 8899 3941 8904
rect 3963 8900 3964 8905
rect 3969 8903 3970 8905
rect 3989 8903 3996 8904
rect 4069 8903 4076 8904
rect 3969 8900 3990 8903
rect 3963 8899 3990 8900
rect 3934 8898 3941 8899
rect 3964 8898 3990 8899
rect 3995 8898 3996 8903
rect 3935 8895 3940 8898
rect 3910 8894 3940 8895
rect 3904 8889 3940 8894
rect 3964 8872 3969 8898
rect 3989 8897 3996 8898
rect 4046 8898 4070 8903
rect 4075 8898 4076 8903
rect 3795 8866 3969 8872
rect 3795 8843 3800 8866
rect 3832 8844 3872 8845
rect 3794 8842 3801 8843
rect 3794 8837 3795 8842
rect 3800 8837 3801 8842
rect 3832 8840 3866 8844
rect 3794 8836 3801 8837
rect 3831 8839 3838 8840
rect 3831 8834 3832 8839
rect 3837 8834 3838 8839
rect 3865 8839 3866 8840
rect 3871 8839 3872 8844
rect 3904 8844 3940 8849
rect 4046 8847 4051 8898
rect 4069 8897 4076 8898
rect 3865 8838 3872 8839
rect 3889 8839 3896 8840
rect 3831 8833 3838 8834
rect 3842 8835 3849 8836
rect 3842 8830 3843 8835
rect 3848 8830 3849 8835
rect 3889 8834 3890 8839
rect 3895 8834 3896 8839
rect 3904 8838 3905 8844
rect 3910 8843 3940 8844
rect 3910 8838 3911 8843
rect 3935 8840 3940 8843
rect 4045 8846 4052 8847
rect 4045 8841 4046 8846
rect 4051 8841 4052 8846
rect 4045 8840 4052 8841
rect 3904 8837 3911 8838
rect 3934 8839 3941 8840
rect 3934 8834 3935 8839
rect 3940 8834 3941 8839
rect 3963 8838 3970 8839
rect 3889 8833 3896 8834
rect 3918 8833 3925 8834
rect 3934 8833 3941 8834
rect 3947 8833 3953 8834
rect 3890 8830 3895 8833
rect 3842 8825 3895 8830
rect 3918 8828 3919 8833
rect 3924 8828 3925 8833
rect 3947 8828 3948 8833
rect 3952 8828 3953 8833
rect 3918 8827 3953 8828
rect 3919 8823 3953 8827
rect 3963 8833 3964 8838
rect 3969 8833 3970 8838
rect 3963 8832 3970 8833
rect 3989 8832 3996 8833
rect 3963 8827 3990 8832
rect 3995 8827 3996 8832
rect 4108 8828 4113 8937
rect 4158 8899 4165 8900
rect 4158 8894 4159 8899
rect 4164 8894 4165 8899
rect 4158 8893 4165 8894
rect 4065 8827 4113 8828
rect 3963 8806 3968 8827
rect 3989 8826 3996 8827
rect 3796 8800 3968 8806
rect 4034 8822 4113 8827
rect 4159 8831 4164 8893
rect 4159 8825 4226 8831
rect 3796 8780 3801 8800
rect 3795 8779 3802 8780
rect 3795 8774 3796 8779
rect 3801 8774 3802 8779
rect 3795 8773 3802 8774
rect 3842 8776 3895 8781
rect 3919 8779 3953 8783
rect 4034 8779 4039 8822
rect 3831 8772 3838 8773
rect 3831 8767 3832 8772
rect 3837 8767 3838 8772
rect 3842 8771 3843 8776
rect 3848 8771 3849 8776
rect 3890 8773 3895 8776
rect 3918 8778 3953 8779
rect 3918 8773 3919 8778
rect 3924 8773 3925 8778
rect 3947 8773 3948 8778
rect 3952 8773 3953 8778
rect 4033 8778 4040 8779
rect 3842 8770 3849 8771
rect 3889 8772 3896 8773
rect 3918 8772 3925 8773
rect 3934 8772 3941 8773
rect 3947 8772 3953 8773
rect 3963 8773 3970 8774
rect 3831 8766 3838 8767
rect 3865 8767 3872 8768
rect 3865 8766 3866 8767
rect 3832 8762 3866 8766
rect 3871 8762 3872 8767
rect 3889 8767 3890 8772
rect 3895 8767 3896 8772
rect 3889 8766 3896 8767
rect 3904 8768 3911 8769
rect 3832 8761 3872 8762
rect 3904 8762 3905 8768
rect 3910 8763 3911 8768
rect 3934 8767 3935 8772
rect 3940 8767 3941 8772
rect 3963 8768 3964 8773
rect 3969 8768 3970 8773
rect 4033 8773 4034 8778
rect 4039 8773 4040 8778
rect 4103 8776 4156 8781
rect 4180 8779 4214 8783
rect 4221 8779 4226 8825
rect 4033 8772 4040 8773
rect 4092 8772 4099 8773
rect 3963 8767 3970 8768
rect 3988 8767 3995 8768
rect 3934 8766 3941 8767
rect 3935 8763 3940 8766
rect 3910 8762 3940 8763
rect 3904 8757 3940 8762
rect 3965 8762 3989 8767
rect 3994 8762 3995 8767
rect 4092 8767 4093 8772
rect 4098 8767 4099 8772
rect 4103 8771 4104 8776
rect 4109 8771 4110 8776
rect 4151 8773 4156 8776
rect 4179 8778 4214 8779
rect 4179 8773 4180 8778
rect 4185 8773 4186 8778
rect 4208 8773 4209 8778
rect 4213 8773 4214 8778
rect 4103 8770 4110 8771
rect 4150 8772 4157 8773
rect 4179 8772 4186 8773
rect 4195 8772 4202 8773
rect 4208 8772 4214 8773
rect 4220 8778 4227 8779
rect 4220 8773 4221 8778
rect 4226 8773 4227 8778
rect 4220 8772 4227 8773
rect 4092 8766 4099 8767
rect 4126 8767 4133 8768
rect 4126 8766 4127 8767
rect 3965 8631 3970 8762
rect 3988 8761 3995 8762
rect 4093 8762 4127 8766
rect 4132 8762 4133 8767
rect 4150 8767 4151 8772
rect 4156 8767 4157 8772
rect 4150 8766 4157 8767
rect 4165 8768 4172 8769
rect 4093 8761 4133 8762
rect 4165 8762 4166 8768
rect 4171 8763 4172 8768
rect 4195 8767 4196 8772
rect 4201 8767 4202 8772
rect 4195 8766 4202 8767
rect 4196 8763 4201 8766
rect 4171 8762 4201 8763
rect 4165 8757 4201 8762
rect 4248 8734 4253 9261
rect 4095 8729 4253 8734
rect 4403 9060 4518 9442
rect 4403 9056 4479 9060
rect 4483 9056 4489 9060
rect 4493 9056 4499 9060
rect 4503 9056 4509 9060
rect 4513 9056 4518 9060
rect 4403 9055 4518 9056
rect 4403 9051 4479 9055
rect 4483 9051 4489 9055
rect 4493 9051 4499 9055
rect 4503 9051 4509 9055
rect 4513 9051 4518 9055
rect 4403 9050 4518 9051
rect 4403 9046 4479 9050
rect 4483 9046 4489 9050
rect 4493 9046 4499 9050
rect 4503 9046 4509 9050
rect 4513 9046 4518 9050
rect 4403 9045 4518 9046
rect 4403 9041 4479 9045
rect 4483 9041 4489 9045
rect 4493 9041 4499 9045
rect 4503 9041 4509 9045
rect 4513 9041 4518 9045
rect 4403 8751 4518 9041
rect 4403 8747 4479 8751
rect 4483 8747 4489 8751
rect 4493 8747 4499 8751
rect 4503 8747 4509 8751
rect 4513 8747 4518 8751
rect 4403 8746 4518 8747
rect 4403 8742 4479 8746
rect 4483 8742 4489 8746
rect 4493 8742 4499 8746
rect 4503 8742 4509 8746
rect 4513 8742 4518 8746
rect 4403 8741 4518 8742
rect 4403 8737 4479 8741
rect 4483 8737 4489 8741
rect 4493 8737 4499 8741
rect 4503 8737 4509 8741
rect 4513 8737 4518 8741
rect 4403 8736 4518 8737
rect 4403 8732 4479 8736
rect 4483 8732 4489 8736
rect 4493 8732 4499 8736
rect 4503 8732 4509 8736
rect 4513 8732 4518 8736
rect 4095 8667 4100 8729
rect 4094 8666 4100 8667
rect 4094 8662 4095 8666
rect 4099 8662 4100 8666
rect 4094 8661 4100 8662
rect 3965 8625 4276 8631
rect 4219 8584 4225 8585
rect 4219 8580 4220 8584
rect 4224 8580 4225 8584
rect 4219 8579 4225 8580
rect 3020 8388 3775 8394
rect 654 8384 659 8388
rect 663 8384 669 8388
rect 673 8384 679 8388
rect 683 8384 689 8388
rect 693 8384 769 8388
rect 654 8383 769 8384
rect 654 8379 659 8383
rect 663 8379 669 8383
rect 673 8379 679 8383
rect 683 8379 689 8383
rect 693 8379 769 8383
rect 654 8089 769 8379
rect 4220 8375 4225 8579
rect 654 8085 659 8089
rect 663 8085 669 8089
rect 673 8085 679 8089
rect 683 8085 689 8089
rect 693 8085 769 8089
rect 654 8084 769 8085
rect 654 8080 659 8084
rect 663 8080 669 8084
rect 673 8080 679 8084
rect 683 8080 689 8084
rect 693 8080 769 8084
rect 654 8079 769 8080
rect 654 8075 659 8079
rect 663 8075 669 8079
rect 673 8075 679 8079
rect 683 8075 689 8079
rect 693 8075 769 8079
rect 654 8074 769 8075
rect 654 8070 659 8074
rect 663 8070 669 8074
rect 673 8070 679 8074
rect 683 8070 689 8074
rect 693 8070 769 8074
rect 654 7780 769 8070
rect 2367 8370 4225 8375
rect 2367 7797 2372 8370
rect 2761 8335 2852 8336
rect 2761 8331 2847 8335
rect 2851 8331 2852 8335
rect 2762 8300 2767 8331
rect 2846 8330 2852 8331
rect 3791 8335 3797 8336
rect 3791 8331 3792 8335
rect 3796 8331 3797 8335
rect 3791 8330 3797 8331
rect 2623 8299 2767 8300
rect 2623 8295 2624 8299
rect 2628 8295 2767 8299
rect 3568 8300 3574 8301
rect 3791 8300 3796 8330
rect 2623 8294 2629 8295
rect 2849 8292 3329 8297
rect 3568 8296 3569 8300
rect 3573 8296 3796 8300
rect 4271 8297 4276 8625
rect 3568 8295 3796 8296
rect 3934 8292 4276 8297
rect 4403 8442 4518 8732
rect 4403 8438 4479 8442
rect 4483 8438 4489 8442
rect 4493 8438 4499 8442
rect 4503 8438 4509 8442
rect 4513 8438 4518 8442
rect 4403 8437 4518 8438
rect 4403 8433 4479 8437
rect 4483 8433 4489 8437
rect 4493 8433 4499 8437
rect 4503 8433 4509 8437
rect 4513 8433 4518 8437
rect 4403 8432 4518 8433
rect 4403 8428 4479 8432
rect 4483 8428 4489 8432
rect 4493 8428 4499 8432
rect 4503 8428 4509 8432
rect 4513 8428 4518 8432
rect 4403 8427 4518 8428
rect 4403 8423 4479 8427
rect 4483 8423 4489 8427
rect 4493 8423 4499 8427
rect 4503 8423 4509 8427
rect 4513 8423 4518 8427
rect 2849 8257 2854 8292
rect 3324 8287 3962 8292
rect 3302 8284 3308 8285
rect 3302 8280 3303 8284
rect 3307 8280 3308 8284
rect 3302 8279 3308 8280
rect 4247 8284 4253 8285
rect 4247 8280 4248 8284
rect 4252 8280 4253 8284
rect 4247 8279 4253 8280
rect 2887 8258 2927 8259
rect 2848 8256 2855 8257
rect 2848 8251 2849 8256
rect 2854 8251 2855 8256
rect 2887 8254 2921 8258
rect 2848 8250 2855 8251
rect 2886 8253 2893 8254
rect 2886 8248 2887 8253
rect 2892 8248 2893 8253
rect 2920 8253 2921 8254
rect 2926 8253 2927 8258
rect 2959 8258 2995 8263
rect 2920 8252 2927 8253
rect 2944 8253 2951 8254
rect 2886 8247 2893 8248
rect 2897 8249 2904 8250
rect 2897 8244 2898 8249
rect 2903 8244 2904 8249
rect 2944 8248 2945 8253
rect 2950 8248 2951 8253
rect 2959 8252 2960 8258
rect 2965 8257 2995 8258
rect 2965 8252 2966 8257
rect 2990 8254 2995 8257
rect 2959 8251 2966 8252
rect 2989 8253 2996 8254
rect 2989 8248 2990 8253
rect 2995 8248 2996 8253
rect 3018 8252 3025 8253
rect 2944 8247 2951 8248
rect 2973 8247 2980 8248
rect 2989 8247 2996 8248
rect 3002 8247 3008 8248
rect 2945 8244 2950 8247
rect 2897 8239 2950 8244
rect 2973 8242 2974 8247
rect 2979 8242 2980 8247
rect 3002 8242 3003 8247
rect 3007 8242 3008 8247
rect 2973 8241 3008 8242
rect 2974 8237 3008 8241
rect 3018 8247 3019 8252
rect 3024 8247 3025 8252
rect 3100 8252 3107 8253
rect 3100 8247 3101 8252
rect 3106 8247 3107 8252
rect 3185 8252 3192 8253
rect 3185 8247 3186 8252
rect 3191 8247 3192 8252
rect 3018 8246 3025 8247
rect 3044 8246 3051 8247
rect 3100 8246 3107 8247
rect 3125 8246 3132 8247
rect 3185 8246 3192 8247
rect 3018 8241 3045 8246
rect 3050 8241 3051 8246
rect 3101 8241 3126 8246
rect 3131 8241 3132 8246
rect 3018 8220 3023 8241
rect 3044 8240 3051 8241
rect 3125 8240 3132 8241
rect 3182 8241 3191 8246
rect 2851 8214 3023 8220
rect 2622 8196 2628 8197
rect 2622 8192 2623 8196
rect 2627 8192 2760 8196
rect 2851 8194 2856 8214
rect 2622 8191 2760 8192
rect 2366 7796 2372 7797
rect 2366 7792 2367 7796
rect 2371 7792 2372 7796
rect 2366 7791 2372 7792
rect 654 7776 659 7780
rect 663 7776 669 7780
rect 673 7776 679 7780
rect 683 7776 689 7780
rect 693 7776 769 7780
rect 654 7775 769 7776
rect 654 7771 659 7775
rect 663 7771 669 7775
rect 673 7771 679 7775
rect 683 7771 689 7775
rect 693 7771 769 7775
rect 654 7770 769 7771
rect 654 7766 659 7770
rect 663 7766 669 7770
rect 673 7766 679 7770
rect 683 7766 689 7770
rect 693 7766 769 7770
rect 654 7765 769 7766
rect 654 7761 659 7765
rect 663 7761 669 7765
rect 673 7761 679 7765
rect 683 7761 689 7765
rect 693 7761 769 7765
rect 654 7471 769 7761
rect 654 7467 659 7471
rect 663 7467 669 7471
rect 673 7467 679 7471
rect 683 7467 689 7471
rect 693 7467 769 7471
rect 654 7466 769 7467
rect 654 7462 659 7466
rect 663 7462 669 7466
rect 673 7462 679 7466
rect 683 7462 689 7466
rect 693 7462 769 7466
rect 654 7461 769 7462
rect 654 7457 659 7461
rect 663 7457 669 7461
rect 673 7457 679 7461
rect 683 7457 689 7461
rect 693 7457 769 7461
rect 654 7456 769 7457
rect 654 7452 659 7456
rect 663 7452 669 7456
rect 673 7452 679 7456
rect 683 7452 689 7456
rect 693 7452 769 7456
rect 654 7162 769 7452
rect 2755 7430 2760 8191
rect 2850 8193 2857 8194
rect 2850 8188 2851 8193
rect 2856 8188 2857 8193
rect 2850 8187 2857 8188
rect 2897 8190 2950 8195
rect 2974 8193 3008 8197
rect 2886 8186 2893 8187
rect 2886 8181 2887 8186
rect 2892 8181 2893 8186
rect 2897 8185 2898 8190
rect 2903 8185 2904 8190
rect 2945 8187 2950 8190
rect 2973 8192 3008 8193
rect 2973 8187 2974 8192
rect 2979 8187 2980 8192
rect 3002 8187 3003 8192
rect 3007 8187 3008 8192
rect 2897 8184 2904 8185
rect 2944 8186 2951 8187
rect 2973 8186 2980 8187
rect 2989 8186 2996 8187
rect 3002 8186 3008 8187
rect 3018 8187 3025 8188
rect 3044 8187 3051 8188
rect 3124 8187 3131 8188
rect 2886 8180 2893 8181
rect 2920 8181 2927 8182
rect 2920 8180 2921 8181
rect 2887 8176 2921 8180
rect 2926 8176 2927 8181
rect 2944 8181 2945 8186
rect 2950 8181 2951 8186
rect 2944 8180 2951 8181
rect 2959 8182 2966 8183
rect 2887 8175 2927 8176
rect 2959 8176 2960 8182
rect 2965 8177 2966 8182
rect 2989 8181 2990 8186
rect 2995 8181 2996 8186
rect 3018 8182 3019 8187
rect 3024 8182 3045 8187
rect 3050 8182 3051 8187
rect 3018 8181 3025 8182
rect 3044 8181 3051 8182
rect 3101 8182 3125 8187
rect 3130 8182 3131 8187
rect 2989 8180 2996 8181
rect 2990 8177 2995 8180
rect 2965 8176 2995 8177
rect 2959 8171 2995 8176
rect 3019 8154 3024 8181
rect 2850 8148 3024 8154
rect 2850 8125 2855 8148
rect 2887 8126 2927 8127
rect 2849 8124 2856 8125
rect 2849 8119 2850 8124
rect 2855 8119 2856 8124
rect 2887 8122 2921 8126
rect 2849 8118 2856 8119
rect 2886 8121 2893 8122
rect 2886 8116 2887 8121
rect 2892 8116 2893 8121
rect 2920 8121 2921 8122
rect 2926 8121 2927 8126
rect 2959 8126 2995 8131
rect 3101 8129 3106 8182
rect 3124 8181 3131 8182
rect 3182 8153 3187 8241
rect 3144 8148 3187 8153
rect 2920 8120 2927 8121
rect 2944 8121 2951 8122
rect 2886 8115 2893 8116
rect 2897 8117 2904 8118
rect 2897 8112 2898 8117
rect 2903 8112 2904 8117
rect 2944 8116 2945 8121
rect 2950 8116 2951 8121
rect 2959 8120 2960 8126
rect 2965 8125 2995 8126
rect 2965 8120 2966 8125
rect 2990 8122 2995 8125
rect 3100 8128 3107 8129
rect 3100 8123 3101 8128
rect 3106 8123 3107 8128
rect 3100 8122 3107 8123
rect 2959 8119 2966 8120
rect 2989 8121 2996 8122
rect 2989 8116 2990 8121
rect 2995 8116 2996 8121
rect 3018 8120 3025 8121
rect 2944 8115 2951 8116
rect 2973 8115 2980 8116
rect 2989 8115 2996 8116
rect 3002 8115 3008 8116
rect 2945 8112 2950 8115
rect 2897 8107 2950 8112
rect 2973 8110 2974 8115
rect 2979 8110 2980 8115
rect 3002 8110 3003 8115
rect 3007 8110 3008 8115
rect 2973 8109 3008 8110
rect 2974 8105 3008 8109
rect 3018 8115 3019 8120
rect 3024 8115 3025 8120
rect 3144 8115 3149 8148
rect 3207 8125 3214 8126
rect 3207 8120 3208 8125
rect 3213 8120 3214 8125
rect 3207 8119 3214 8120
rect 3018 8114 3025 8115
rect 3044 8114 3051 8115
rect 3018 8109 3045 8114
rect 3050 8109 3051 8114
rect 3144 8114 3156 8115
rect 3144 8109 3150 8114
rect 3155 8109 3156 8114
rect 3018 8088 3023 8109
rect 3044 8108 3051 8109
rect 3149 8108 3156 8109
rect 2851 8082 3023 8088
rect 2851 8062 2856 8082
rect 2850 8061 2857 8062
rect 2850 8056 2851 8061
rect 2856 8056 2857 8061
rect 2850 8055 2857 8056
rect 2897 8058 2950 8063
rect 2974 8061 3008 8065
rect 2886 8054 2893 8055
rect 2886 8049 2887 8054
rect 2892 8049 2893 8054
rect 2897 8053 2898 8058
rect 2903 8053 2904 8058
rect 2945 8055 2950 8058
rect 2973 8060 3008 8061
rect 2973 8055 2974 8060
rect 2979 8055 2980 8060
rect 3002 8055 3003 8060
rect 3007 8055 3008 8060
rect 3043 8056 3050 8057
rect 3149 8056 3156 8057
rect 2897 8052 2904 8053
rect 2944 8054 2951 8055
rect 2973 8054 2980 8055
rect 2989 8054 2996 8055
rect 3002 8054 3008 8055
rect 3018 8055 3044 8056
rect 2886 8048 2893 8049
rect 2920 8049 2927 8050
rect 2920 8048 2921 8049
rect 2887 8044 2921 8048
rect 2926 8044 2927 8049
rect 2944 8049 2945 8054
rect 2950 8049 2951 8054
rect 2944 8048 2951 8049
rect 2959 8050 2966 8051
rect 2887 8043 2927 8044
rect 2959 8044 2960 8050
rect 2965 8045 2966 8050
rect 2989 8049 2990 8054
rect 2995 8049 2996 8054
rect 2989 8048 2996 8049
rect 3018 8050 3019 8055
rect 3024 8051 3044 8055
rect 3049 8051 3050 8056
rect 3024 8050 3025 8051
rect 3043 8050 3050 8051
rect 3145 8051 3150 8056
rect 3155 8051 3156 8056
rect 3145 8050 3156 8051
rect 3018 8049 3025 8050
rect 2990 8045 2995 8048
rect 2965 8044 2995 8045
rect 2959 8039 2995 8044
rect 3018 8022 3023 8049
rect 2850 8016 3023 8022
rect 3145 8022 3150 8050
rect 3145 8017 3188 8022
rect 2850 7993 2855 8016
rect 2887 7994 2927 7995
rect 2849 7992 2856 7993
rect 2849 7987 2850 7992
rect 2855 7987 2856 7992
rect 2887 7990 2921 7994
rect 2849 7986 2856 7987
rect 2886 7989 2893 7990
rect 2886 7984 2887 7989
rect 2892 7984 2893 7989
rect 2920 7989 2921 7990
rect 2926 7989 2927 7994
rect 2959 7994 2995 7999
rect 3183 7998 3188 8017
rect 2920 7988 2927 7989
rect 2944 7989 2951 7990
rect 2886 7983 2893 7984
rect 2897 7985 2904 7986
rect 2897 7980 2898 7985
rect 2903 7980 2904 7985
rect 2944 7984 2945 7989
rect 2950 7984 2951 7989
rect 2959 7988 2960 7994
rect 2965 7993 2995 7994
rect 2965 7988 2966 7993
rect 2990 7990 2995 7993
rect 3182 7997 3189 7998
rect 3182 7992 3183 7997
rect 3188 7992 3189 7997
rect 3182 7991 3189 7992
rect 3208 7990 3213 8119
rect 3216 7990 3223 7991
rect 2959 7987 2966 7988
rect 2989 7989 2996 7990
rect 2989 7984 2990 7989
rect 2995 7984 2996 7989
rect 3018 7988 3025 7989
rect 2944 7983 2951 7984
rect 2973 7983 2980 7984
rect 2989 7983 2996 7984
rect 3002 7983 3008 7984
rect 2945 7980 2950 7983
rect 2897 7975 2950 7980
rect 2973 7978 2974 7983
rect 2979 7978 2980 7983
rect 3002 7978 3003 7983
rect 3007 7978 3008 7983
rect 2973 7977 3008 7978
rect 2974 7973 3008 7977
rect 3018 7983 3019 7988
rect 3024 7983 3025 7988
rect 3100 7988 3107 7989
rect 3100 7983 3101 7988
rect 3106 7983 3107 7988
rect 3196 7985 3217 7990
rect 3222 7985 3223 7990
rect 3196 7984 3208 7985
rect 3216 7984 3223 7985
rect 3018 7982 3025 7983
rect 3044 7982 3051 7983
rect 3100 7982 3107 7983
rect 3125 7982 3132 7983
rect 3018 7977 3045 7982
rect 3050 7977 3051 7982
rect 3101 7977 3126 7982
rect 3131 7977 3132 7982
rect 3018 7956 3023 7977
rect 3044 7976 3051 7977
rect 3125 7976 3132 7977
rect 3196 7976 3201 7984
rect 2851 7950 3023 7956
rect 3163 7955 3201 7976
rect 2851 7930 2856 7950
rect 2850 7929 2857 7930
rect 2850 7924 2851 7929
rect 2856 7924 2857 7929
rect 2850 7923 2857 7924
rect 2897 7926 2950 7931
rect 2974 7929 3008 7933
rect 2886 7922 2893 7923
rect 2886 7917 2887 7922
rect 2892 7917 2893 7922
rect 2897 7921 2898 7926
rect 2903 7921 2904 7926
rect 2945 7923 2950 7926
rect 2973 7928 3008 7929
rect 2973 7923 2974 7928
rect 2979 7923 2980 7928
rect 3002 7923 3003 7928
rect 3007 7923 3008 7928
rect 2897 7920 2904 7921
rect 2944 7922 2951 7923
rect 2973 7922 2980 7923
rect 2989 7922 2996 7923
rect 3002 7922 3008 7923
rect 3018 7923 3025 7924
rect 2886 7916 2893 7917
rect 2920 7917 2927 7918
rect 2920 7916 2921 7917
rect 2887 7912 2921 7916
rect 2926 7912 2927 7917
rect 2944 7917 2945 7922
rect 2950 7917 2951 7922
rect 2944 7916 2951 7917
rect 2959 7918 2966 7919
rect 2887 7911 2927 7912
rect 2959 7912 2960 7918
rect 2965 7913 2966 7918
rect 2989 7917 2990 7922
rect 2995 7917 2996 7922
rect 3018 7918 3019 7923
rect 3024 7921 3025 7923
rect 3044 7921 3051 7922
rect 3124 7921 3131 7922
rect 3024 7918 3045 7921
rect 3018 7917 3045 7918
rect 2989 7916 2996 7917
rect 3019 7916 3045 7917
rect 3050 7916 3051 7921
rect 2990 7913 2995 7916
rect 2965 7912 2995 7913
rect 2959 7907 2995 7912
rect 3019 7890 3024 7916
rect 3044 7915 3051 7916
rect 3101 7916 3125 7921
rect 3130 7916 3131 7921
rect 2850 7884 3024 7890
rect 2850 7861 2855 7884
rect 2887 7862 2927 7863
rect 2849 7860 2856 7861
rect 2849 7855 2850 7860
rect 2855 7855 2856 7860
rect 2887 7858 2921 7862
rect 2849 7854 2856 7855
rect 2886 7857 2893 7858
rect 2886 7852 2887 7857
rect 2892 7852 2893 7857
rect 2920 7857 2921 7858
rect 2926 7857 2927 7862
rect 2959 7862 2995 7867
rect 3101 7865 3106 7916
rect 3124 7915 3131 7916
rect 2920 7856 2927 7857
rect 2944 7857 2951 7858
rect 2886 7851 2893 7852
rect 2897 7853 2904 7854
rect 2897 7848 2898 7853
rect 2903 7848 2904 7853
rect 2944 7852 2945 7857
rect 2950 7852 2951 7857
rect 2959 7856 2960 7862
rect 2965 7861 2995 7862
rect 2965 7856 2966 7861
rect 2990 7858 2995 7861
rect 3100 7864 3107 7865
rect 3100 7859 3101 7864
rect 3106 7859 3107 7864
rect 3100 7858 3107 7859
rect 2959 7855 2966 7856
rect 2989 7857 2996 7858
rect 2989 7852 2990 7857
rect 2995 7852 2996 7857
rect 3018 7856 3025 7857
rect 2944 7851 2951 7852
rect 2973 7851 2980 7852
rect 2989 7851 2996 7852
rect 3002 7851 3008 7852
rect 2945 7848 2950 7851
rect 2897 7843 2950 7848
rect 2973 7846 2974 7851
rect 2979 7846 2980 7851
rect 3002 7846 3003 7851
rect 3007 7846 3008 7851
rect 2973 7845 3008 7846
rect 2974 7841 3008 7845
rect 3018 7851 3019 7856
rect 3024 7851 3025 7856
rect 3018 7850 3025 7851
rect 3044 7850 3051 7851
rect 3018 7845 3045 7850
rect 3050 7845 3051 7850
rect 3163 7846 3168 7955
rect 3213 7917 3220 7918
rect 3213 7912 3214 7917
rect 3219 7912 3220 7917
rect 3213 7911 3220 7912
rect 3120 7845 3168 7846
rect 3018 7824 3023 7845
rect 3044 7844 3051 7845
rect 2851 7818 3023 7824
rect 3089 7840 3168 7845
rect 3214 7849 3219 7911
rect 3214 7843 3281 7849
rect 2851 7798 2856 7818
rect 2850 7797 2857 7798
rect 2850 7792 2851 7797
rect 2856 7792 2857 7797
rect 2850 7791 2857 7792
rect 2897 7794 2950 7799
rect 2974 7797 3008 7801
rect 3089 7797 3094 7840
rect 2886 7790 2893 7791
rect 2886 7785 2887 7790
rect 2892 7785 2893 7790
rect 2897 7789 2898 7794
rect 2903 7789 2904 7794
rect 2945 7791 2950 7794
rect 2973 7796 3008 7797
rect 2973 7791 2974 7796
rect 2979 7791 2980 7796
rect 3002 7791 3003 7796
rect 3007 7791 3008 7796
rect 3088 7796 3095 7797
rect 2897 7788 2904 7789
rect 2944 7790 2951 7791
rect 2973 7790 2980 7791
rect 2989 7790 2996 7791
rect 3002 7790 3008 7791
rect 3018 7791 3025 7792
rect 2886 7784 2893 7785
rect 2920 7785 2927 7786
rect 2920 7784 2921 7785
rect 2887 7780 2921 7784
rect 2926 7780 2927 7785
rect 2944 7785 2945 7790
rect 2950 7785 2951 7790
rect 2944 7784 2951 7785
rect 2959 7786 2966 7787
rect 2887 7779 2927 7780
rect 2959 7780 2960 7786
rect 2965 7781 2966 7786
rect 2989 7785 2990 7790
rect 2995 7785 2996 7790
rect 3018 7786 3019 7791
rect 3024 7786 3025 7791
rect 3088 7791 3089 7796
rect 3094 7791 3095 7796
rect 3158 7794 3211 7799
rect 3235 7797 3269 7801
rect 3276 7797 3281 7843
rect 3088 7790 3095 7791
rect 3147 7790 3154 7791
rect 3018 7785 3025 7786
rect 3043 7785 3050 7786
rect 2989 7784 2996 7785
rect 2990 7781 2995 7784
rect 2965 7780 2995 7781
rect 2959 7775 2995 7780
rect 3020 7780 3044 7785
rect 3049 7780 3050 7785
rect 3147 7785 3148 7790
rect 3153 7785 3154 7790
rect 3158 7789 3159 7794
rect 3164 7789 3165 7794
rect 3206 7791 3211 7794
rect 3234 7796 3269 7797
rect 3234 7791 3235 7796
rect 3240 7791 3241 7796
rect 3263 7791 3264 7796
rect 3268 7791 3269 7796
rect 3158 7788 3165 7789
rect 3205 7790 3212 7791
rect 3234 7790 3241 7791
rect 3250 7790 3257 7791
rect 3263 7790 3269 7791
rect 3275 7796 3282 7797
rect 3275 7791 3276 7796
rect 3281 7791 3282 7796
rect 3275 7790 3282 7791
rect 3147 7784 3154 7785
rect 3181 7785 3188 7786
rect 3181 7784 3182 7785
rect 2755 7429 2761 7430
rect 2755 7425 2756 7429
rect 2760 7425 2761 7429
rect 2755 7424 2761 7425
rect 3020 7427 3025 7780
rect 3043 7779 3050 7780
rect 3148 7780 3182 7784
rect 3187 7780 3188 7785
rect 3205 7785 3206 7790
rect 3211 7785 3212 7790
rect 3205 7784 3212 7785
rect 3220 7786 3227 7787
rect 3148 7779 3188 7780
rect 3220 7780 3221 7786
rect 3226 7781 3227 7786
rect 3250 7785 3251 7790
rect 3256 7785 3257 7790
rect 3250 7784 3257 7785
rect 3251 7781 3256 7784
rect 3226 7780 3256 7781
rect 3220 7775 3256 7780
rect 3303 7752 3308 8279
rect 3832 8258 3872 8259
rect 3793 8256 3800 8257
rect 3770 8251 3794 8256
rect 3799 8251 3800 8256
rect 3832 8254 3866 8258
rect 3567 8196 3573 8197
rect 3567 8192 3568 8196
rect 3572 8192 3705 8196
rect 3567 8191 3705 8192
rect 3311 7796 3317 7797
rect 3311 7792 3312 7796
rect 3316 7792 3317 7796
rect 3311 7791 3317 7792
rect 3150 7747 3308 7752
rect 3150 7685 3155 7747
rect 3149 7684 3155 7685
rect 3149 7680 3150 7684
rect 3154 7680 3155 7684
rect 3149 7679 3155 7680
rect 3312 7622 3317 7791
rect 3275 7617 3317 7622
rect 3275 7603 3280 7617
rect 3274 7602 3280 7603
rect 3274 7598 3275 7602
rect 3279 7598 3280 7602
rect 3274 7597 3280 7598
rect 3700 7430 3705 8191
rect 3700 7429 3706 7430
rect 3020 7422 3065 7427
rect 3700 7425 3701 7429
rect 3705 7425 3706 7429
rect 3700 7424 3706 7425
rect 3770 7418 3775 8251
rect 3793 8250 3800 8251
rect 3831 8253 3838 8254
rect 3831 8248 3832 8253
rect 3837 8248 3838 8253
rect 3865 8253 3866 8254
rect 3871 8253 3872 8258
rect 3904 8258 3940 8263
rect 3865 8252 3872 8253
rect 3889 8253 3896 8254
rect 3831 8247 3838 8248
rect 3842 8249 3849 8250
rect 3842 8244 3843 8249
rect 3848 8244 3849 8249
rect 3889 8248 3890 8253
rect 3895 8248 3896 8253
rect 3904 8252 3905 8258
rect 3910 8257 3940 8258
rect 3910 8252 3911 8257
rect 3935 8254 3940 8257
rect 3904 8251 3911 8252
rect 3934 8253 3941 8254
rect 3934 8248 3935 8253
rect 3940 8248 3941 8253
rect 3963 8252 3970 8253
rect 3889 8247 3896 8248
rect 3918 8247 3925 8248
rect 3934 8247 3941 8248
rect 3947 8247 3953 8248
rect 3890 8244 3895 8247
rect 3842 8239 3895 8244
rect 3918 8242 3919 8247
rect 3924 8242 3925 8247
rect 3947 8242 3948 8247
rect 3952 8242 3953 8247
rect 3918 8241 3953 8242
rect 3919 8237 3953 8241
rect 3963 8247 3964 8252
rect 3969 8247 3970 8252
rect 4045 8252 4052 8253
rect 4045 8247 4046 8252
rect 4051 8247 4052 8252
rect 4130 8252 4137 8253
rect 4130 8247 4131 8252
rect 4136 8247 4137 8252
rect 3963 8246 3970 8247
rect 3989 8246 3996 8247
rect 4045 8246 4052 8247
rect 4070 8246 4077 8247
rect 4130 8246 4137 8247
rect 3963 8241 3990 8246
rect 3995 8241 3996 8246
rect 4046 8241 4071 8246
rect 4076 8241 4077 8246
rect 3963 8220 3968 8241
rect 3989 8240 3996 8241
rect 4070 8240 4077 8241
rect 4127 8241 4136 8246
rect 3796 8214 3968 8220
rect 3796 8194 3801 8214
rect 3795 8193 3802 8194
rect 3795 8188 3796 8193
rect 3801 8188 3802 8193
rect 3795 8187 3802 8188
rect 3842 8190 3895 8195
rect 3919 8193 3953 8197
rect 3831 8186 3838 8187
rect 3831 8181 3832 8186
rect 3837 8181 3838 8186
rect 3842 8185 3843 8190
rect 3848 8185 3849 8190
rect 3890 8187 3895 8190
rect 3918 8192 3953 8193
rect 3918 8187 3919 8192
rect 3924 8187 3925 8192
rect 3947 8187 3948 8192
rect 3952 8187 3953 8192
rect 3842 8184 3849 8185
rect 3889 8186 3896 8187
rect 3918 8186 3925 8187
rect 3934 8186 3941 8187
rect 3947 8186 3953 8187
rect 3963 8187 3970 8188
rect 3989 8187 3996 8188
rect 4069 8187 4076 8188
rect 3831 8180 3838 8181
rect 3865 8181 3872 8182
rect 3865 8180 3866 8181
rect 3832 8176 3866 8180
rect 3871 8176 3872 8181
rect 3889 8181 3890 8186
rect 3895 8181 3896 8186
rect 3889 8180 3896 8181
rect 3904 8182 3911 8183
rect 3832 8175 3872 8176
rect 3904 8176 3905 8182
rect 3910 8177 3911 8182
rect 3934 8181 3935 8186
rect 3940 8181 3941 8186
rect 3963 8182 3964 8187
rect 3969 8182 3990 8187
rect 3995 8182 3996 8187
rect 3963 8181 3970 8182
rect 3989 8181 3996 8182
rect 4046 8182 4070 8187
rect 4075 8182 4076 8187
rect 3934 8180 3941 8181
rect 3935 8177 3940 8180
rect 3910 8176 3940 8177
rect 3904 8171 3940 8176
rect 3964 8154 3969 8181
rect 3795 8148 3969 8154
rect 3795 8125 3800 8148
rect 3832 8126 3872 8127
rect 3794 8124 3801 8125
rect 3794 8119 3795 8124
rect 3800 8119 3801 8124
rect 3832 8122 3866 8126
rect 3794 8118 3801 8119
rect 3831 8121 3838 8122
rect 3831 8116 3832 8121
rect 3837 8116 3838 8121
rect 3865 8121 3866 8122
rect 3871 8121 3872 8126
rect 3904 8126 3940 8131
rect 4046 8129 4051 8182
rect 4069 8181 4076 8182
rect 4127 8153 4132 8241
rect 4089 8148 4132 8153
rect 3865 8120 3872 8121
rect 3889 8121 3896 8122
rect 3831 8115 3838 8116
rect 3842 8117 3849 8118
rect 3842 8112 3843 8117
rect 3848 8112 3849 8117
rect 3889 8116 3890 8121
rect 3895 8116 3896 8121
rect 3904 8120 3905 8126
rect 3910 8125 3940 8126
rect 3910 8120 3911 8125
rect 3935 8122 3940 8125
rect 4045 8128 4052 8129
rect 4045 8123 4046 8128
rect 4051 8123 4052 8128
rect 4045 8122 4052 8123
rect 3904 8119 3911 8120
rect 3934 8121 3941 8122
rect 3934 8116 3935 8121
rect 3940 8116 3941 8121
rect 3963 8120 3970 8121
rect 3889 8115 3896 8116
rect 3918 8115 3925 8116
rect 3934 8115 3941 8116
rect 3947 8115 3953 8116
rect 3890 8112 3895 8115
rect 3842 8107 3895 8112
rect 3918 8110 3919 8115
rect 3924 8110 3925 8115
rect 3947 8110 3948 8115
rect 3952 8110 3953 8115
rect 3918 8109 3953 8110
rect 3919 8105 3953 8109
rect 3963 8115 3964 8120
rect 3969 8115 3970 8120
rect 4089 8115 4094 8148
rect 4152 8125 4159 8126
rect 4152 8120 4153 8125
rect 4158 8120 4159 8125
rect 4152 8119 4159 8120
rect 3963 8114 3970 8115
rect 3989 8114 3996 8115
rect 3963 8109 3990 8114
rect 3995 8109 3996 8114
rect 4089 8114 4101 8115
rect 4089 8109 4095 8114
rect 4100 8109 4101 8114
rect 3963 8088 3968 8109
rect 3989 8108 3996 8109
rect 4094 8108 4101 8109
rect 3796 8082 3968 8088
rect 3796 8062 3801 8082
rect 3795 8061 3802 8062
rect 3795 8056 3796 8061
rect 3801 8056 3802 8061
rect 3795 8055 3802 8056
rect 3842 8058 3895 8063
rect 3919 8061 3953 8065
rect 3831 8054 3838 8055
rect 3831 8049 3832 8054
rect 3837 8049 3838 8054
rect 3842 8053 3843 8058
rect 3848 8053 3849 8058
rect 3890 8055 3895 8058
rect 3918 8060 3953 8061
rect 3918 8055 3919 8060
rect 3924 8055 3925 8060
rect 3947 8055 3948 8060
rect 3952 8055 3953 8060
rect 3988 8056 3995 8057
rect 4094 8056 4101 8057
rect 3842 8052 3849 8053
rect 3889 8054 3896 8055
rect 3918 8054 3925 8055
rect 3934 8054 3941 8055
rect 3947 8054 3953 8055
rect 3963 8055 3989 8056
rect 3831 8048 3838 8049
rect 3865 8049 3872 8050
rect 3865 8048 3866 8049
rect 3832 8044 3866 8048
rect 3871 8044 3872 8049
rect 3889 8049 3890 8054
rect 3895 8049 3896 8054
rect 3889 8048 3896 8049
rect 3904 8050 3911 8051
rect 3832 8043 3872 8044
rect 3904 8044 3905 8050
rect 3910 8045 3911 8050
rect 3934 8049 3935 8054
rect 3940 8049 3941 8054
rect 3934 8048 3941 8049
rect 3963 8050 3964 8055
rect 3969 8051 3989 8055
rect 3994 8051 3995 8056
rect 3969 8050 3970 8051
rect 3988 8050 3995 8051
rect 4090 8051 4095 8056
rect 4100 8051 4101 8056
rect 4090 8050 4101 8051
rect 3963 8049 3970 8050
rect 3935 8045 3940 8048
rect 3910 8044 3940 8045
rect 3904 8039 3940 8044
rect 3963 8022 3968 8049
rect 3795 8016 3968 8022
rect 4090 8022 4095 8050
rect 4090 8017 4133 8022
rect 3795 7993 3800 8016
rect 3832 7994 3872 7995
rect 3794 7992 3801 7993
rect 3794 7987 3795 7992
rect 3800 7987 3801 7992
rect 3832 7990 3866 7994
rect 3794 7986 3801 7987
rect 3831 7989 3838 7990
rect 3831 7984 3832 7989
rect 3837 7984 3838 7989
rect 3865 7989 3866 7990
rect 3871 7989 3872 7994
rect 3904 7994 3940 7999
rect 4128 7998 4133 8017
rect 3865 7988 3872 7989
rect 3889 7989 3896 7990
rect 3831 7983 3838 7984
rect 3842 7985 3849 7986
rect 3842 7980 3843 7985
rect 3848 7980 3849 7985
rect 3889 7984 3890 7989
rect 3895 7984 3896 7989
rect 3904 7988 3905 7994
rect 3910 7993 3940 7994
rect 3910 7988 3911 7993
rect 3935 7990 3940 7993
rect 4127 7997 4134 7998
rect 4127 7992 4128 7997
rect 4133 7992 4134 7997
rect 4127 7991 4134 7992
rect 4153 7990 4158 8119
rect 4161 7990 4168 7991
rect 3904 7987 3911 7988
rect 3934 7989 3941 7990
rect 3934 7984 3935 7989
rect 3940 7984 3941 7989
rect 3963 7988 3970 7989
rect 3889 7983 3896 7984
rect 3918 7983 3925 7984
rect 3934 7983 3941 7984
rect 3947 7983 3953 7984
rect 3890 7980 3895 7983
rect 3842 7975 3895 7980
rect 3918 7978 3919 7983
rect 3924 7978 3925 7983
rect 3947 7978 3948 7983
rect 3952 7978 3953 7983
rect 3918 7977 3953 7978
rect 3919 7973 3953 7977
rect 3963 7983 3964 7988
rect 3969 7983 3970 7988
rect 4045 7988 4052 7989
rect 4045 7983 4046 7988
rect 4051 7983 4052 7988
rect 4141 7985 4162 7990
rect 4167 7985 4168 7990
rect 4141 7984 4153 7985
rect 4161 7984 4168 7985
rect 3963 7982 3970 7983
rect 3989 7982 3996 7983
rect 4045 7982 4052 7983
rect 4070 7982 4077 7983
rect 3963 7977 3990 7982
rect 3995 7977 3996 7982
rect 4046 7977 4071 7982
rect 4076 7977 4077 7982
rect 3963 7956 3968 7977
rect 3989 7976 3996 7977
rect 4070 7976 4077 7977
rect 4141 7976 4146 7984
rect 3796 7950 3968 7956
rect 4108 7955 4146 7976
rect 3796 7930 3801 7950
rect 3795 7929 3802 7930
rect 3795 7924 3796 7929
rect 3801 7924 3802 7929
rect 3795 7923 3802 7924
rect 3842 7926 3895 7931
rect 3919 7929 3953 7933
rect 3831 7922 3838 7923
rect 3831 7917 3832 7922
rect 3837 7917 3838 7922
rect 3842 7921 3843 7926
rect 3848 7921 3849 7926
rect 3890 7923 3895 7926
rect 3918 7928 3953 7929
rect 3918 7923 3919 7928
rect 3924 7923 3925 7928
rect 3947 7923 3948 7928
rect 3952 7923 3953 7928
rect 3842 7920 3849 7921
rect 3889 7922 3896 7923
rect 3918 7922 3925 7923
rect 3934 7922 3941 7923
rect 3947 7922 3953 7923
rect 3963 7923 3970 7924
rect 3831 7916 3838 7917
rect 3865 7917 3872 7918
rect 3865 7916 3866 7917
rect 3832 7912 3866 7916
rect 3871 7912 3872 7917
rect 3889 7917 3890 7922
rect 3895 7917 3896 7922
rect 3889 7916 3896 7917
rect 3904 7918 3911 7919
rect 3832 7911 3872 7912
rect 3904 7912 3905 7918
rect 3910 7913 3911 7918
rect 3934 7917 3935 7922
rect 3940 7917 3941 7922
rect 3963 7918 3964 7923
rect 3969 7921 3970 7923
rect 3989 7921 3996 7922
rect 4069 7921 4076 7922
rect 3969 7918 3990 7921
rect 3963 7917 3990 7918
rect 3934 7916 3941 7917
rect 3964 7916 3990 7917
rect 3995 7916 3996 7921
rect 3935 7913 3940 7916
rect 3910 7912 3940 7913
rect 3904 7907 3940 7912
rect 3964 7890 3969 7916
rect 3989 7915 3996 7916
rect 4046 7916 4070 7921
rect 4075 7916 4076 7921
rect 3795 7884 3969 7890
rect 3795 7861 3800 7884
rect 3832 7862 3872 7863
rect 3794 7860 3801 7861
rect 3794 7855 3795 7860
rect 3800 7855 3801 7860
rect 3832 7858 3866 7862
rect 3794 7854 3801 7855
rect 3831 7857 3838 7858
rect 3831 7852 3832 7857
rect 3837 7852 3838 7857
rect 3865 7857 3866 7858
rect 3871 7857 3872 7862
rect 3904 7862 3940 7867
rect 4046 7865 4051 7916
rect 4069 7915 4076 7916
rect 3865 7856 3872 7857
rect 3889 7857 3896 7858
rect 3831 7851 3838 7852
rect 3842 7853 3849 7854
rect 3842 7848 3843 7853
rect 3848 7848 3849 7853
rect 3889 7852 3890 7857
rect 3895 7852 3896 7857
rect 3904 7856 3905 7862
rect 3910 7861 3940 7862
rect 3910 7856 3911 7861
rect 3935 7858 3940 7861
rect 4045 7864 4052 7865
rect 4045 7859 4046 7864
rect 4051 7859 4052 7864
rect 4045 7858 4052 7859
rect 3904 7855 3911 7856
rect 3934 7857 3941 7858
rect 3934 7852 3935 7857
rect 3940 7852 3941 7857
rect 3963 7856 3970 7857
rect 3889 7851 3896 7852
rect 3918 7851 3925 7852
rect 3934 7851 3941 7852
rect 3947 7851 3953 7852
rect 3890 7848 3895 7851
rect 3842 7843 3895 7848
rect 3918 7846 3919 7851
rect 3924 7846 3925 7851
rect 3947 7846 3948 7851
rect 3952 7846 3953 7851
rect 3918 7845 3953 7846
rect 3919 7841 3953 7845
rect 3963 7851 3964 7856
rect 3969 7851 3970 7856
rect 3963 7850 3970 7851
rect 3989 7850 3996 7851
rect 3963 7845 3990 7850
rect 3995 7845 3996 7850
rect 4108 7846 4113 7955
rect 4158 7917 4165 7918
rect 4158 7912 4159 7917
rect 4164 7912 4165 7917
rect 4158 7911 4165 7912
rect 4065 7845 4113 7846
rect 3963 7824 3968 7845
rect 3989 7844 3996 7845
rect 3796 7818 3968 7824
rect 4034 7840 4113 7845
rect 4159 7849 4164 7911
rect 4159 7843 4226 7849
rect 3796 7798 3801 7818
rect 3795 7797 3802 7798
rect 3795 7792 3796 7797
rect 3801 7792 3802 7797
rect 3795 7791 3802 7792
rect 3842 7794 3895 7799
rect 3919 7797 3953 7801
rect 4034 7797 4039 7840
rect 3831 7790 3838 7791
rect 3831 7785 3832 7790
rect 3837 7785 3838 7790
rect 3842 7789 3843 7794
rect 3848 7789 3849 7794
rect 3890 7791 3895 7794
rect 3918 7796 3953 7797
rect 3918 7791 3919 7796
rect 3924 7791 3925 7796
rect 3947 7791 3948 7796
rect 3952 7791 3953 7796
rect 4033 7796 4040 7797
rect 3842 7788 3849 7789
rect 3889 7790 3896 7791
rect 3918 7790 3925 7791
rect 3934 7790 3941 7791
rect 3947 7790 3953 7791
rect 3963 7791 3970 7792
rect 3831 7784 3838 7785
rect 3865 7785 3872 7786
rect 3865 7784 3866 7785
rect 3832 7780 3866 7784
rect 3871 7780 3872 7785
rect 3889 7785 3890 7790
rect 3895 7785 3896 7790
rect 3889 7784 3896 7785
rect 3904 7786 3911 7787
rect 3832 7779 3872 7780
rect 3904 7780 3905 7786
rect 3910 7781 3911 7786
rect 3934 7785 3935 7790
rect 3940 7785 3941 7790
rect 3963 7786 3964 7791
rect 3969 7786 3970 7791
rect 4033 7791 4034 7796
rect 4039 7791 4040 7796
rect 4103 7794 4156 7799
rect 4180 7797 4214 7801
rect 4221 7797 4226 7843
rect 4033 7790 4040 7791
rect 4092 7790 4099 7791
rect 3963 7785 3970 7786
rect 3988 7785 3995 7786
rect 3934 7784 3941 7785
rect 3935 7781 3940 7784
rect 3910 7780 3940 7781
rect 3965 7780 3989 7785
rect 3994 7780 3995 7785
rect 4092 7785 4093 7790
rect 4098 7785 4099 7790
rect 4103 7789 4104 7794
rect 4109 7789 4110 7794
rect 4151 7791 4156 7794
rect 4179 7796 4214 7797
rect 4179 7791 4180 7796
rect 4185 7791 4186 7796
rect 4208 7791 4209 7796
rect 4213 7791 4214 7796
rect 4103 7788 4110 7789
rect 4150 7790 4157 7791
rect 4179 7790 4186 7791
rect 4195 7790 4202 7791
rect 4208 7790 4214 7791
rect 4220 7796 4227 7797
rect 4220 7791 4221 7796
rect 4226 7791 4227 7796
rect 4220 7790 4227 7791
rect 4092 7784 4099 7785
rect 4126 7785 4133 7786
rect 4126 7784 4127 7785
rect 3904 7775 3940 7780
rect 3988 7779 3995 7780
rect 4093 7780 4127 7784
rect 4132 7780 4133 7785
rect 4150 7785 4151 7790
rect 4156 7785 4157 7790
rect 4150 7784 4157 7785
rect 4165 7786 4172 7787
rect 4093 7779 4133 7780
rect 4165 7780 4166 7786
rect 4171 7781 4172 7786
rect 4195 7785 4196 7790
rect 4201 7785 4202 7790
rect 4195 7784 4202 7785
rect 4196 7781 4201 7784
rect 4171 7780 4201 7781
rect 4165 7775 4201 7780
rect 4248 7752 4253 8279
rect 4403 8133 4518 8423
rect 4403 8129 4479 8133
rect 4483 8129 4489 8133
rect 4493 8129 4499 8133
rect 4503 8129 4509 8133
rect 4513 8129 4518 8133
rect 4403 8128 4518 8129
rect 4403 8124 4479 8128
rect 4483 8124 4489 8128
rect 4493 8124 4499 8128
rect 4503 8124 4509 8128
rect 4513 8124 4518 8128
rect 4403 8123 4518 8124
rect 4403 8119 4479 8123
rect 4483 8119 4489 8123
rect 4493 8119 4499 8123
rect 4503 8119 4509 8123
rect 4513 8119 4518 8123
rect 4403 8118 4518 8119
rect 4403 8114 4479 8118
rect 4483 8114 4489 8118
rect 4493 8114 4499 8118
rect 4503 8114 4509 8118
rect 4513 8114 4518 8118
rect 4403 8102 4518 8114
rect 4403 8098 4479 8102
rect 4483 8098 4489 8102
rect 4493 8098 4499 8102
rect 4503 8098 4509 8102
rect 4513 8098 4518 8102
rect 4403 8097 4518 8098
rect 4403 8093 4479 8097
rect 4483 8093 4489 8097
rect 4493 8093 4499 8097
rect 4503 8093 4509 8097
rect 4513 8093 4518 8097
rect 4403 8092 4518 8093
rect 4403 8088 4479 8092
rect 4483 8088 4489 8092
rect 4493 8088 4499 8092
rect 4503 8088 4509 8092
rect 4513 8088 4518 8092
rect 4403 8087 4518 8088
rect 4403 8083 4479 8087
rect 4483 8083 4489 8087
rect 4493 8083 4499 8087
rect 4503 8083 4509 8087
rect 4513 8083 4518 8087
rect 4403 8078 4518 8083
rect 4403 8074 4496 8078
rect 4500 8074 4501 8078
rect 4505 8074 4518 8078
rect 4403 8073 4518 8074
rect 4403 8069 4496 8073
rect 4500 8069 4501 8073
rect 4505 8069 4518 8073
rect 4403 8068 4518 8069
rect 4403 8064 4496 8068
rect 4500 8064 4501 8068
rect 4505 8064 4518 8068
rect 4403 8063 4518 8064
rect 4403 8059 4496 8063
rect 4500 8059 4501 8063
rect 4505 8059 4518 8063
rect 4403 8058 4518 8059
rect 4403 8054 4496 8058
rect 4500 8054 4501 8058
rect 4505 8054 4518 8058
rect 4403 8053 4518 8054
rect 4403 8049 4496 8053
rect 4500 8049 4501 8053
rect 4505 8049 4518 8053
rect 4403 8048 4518 8049
rect 4403 8044 4496 8048
rect 4500 8044 4501 8048
rect 4505 8044 4518 8048
rect 4403 8043 4518 8044
rect 4403 8039 4496 8043
rect 4500 8039 4501 8043
rect 4505 8039 4518 8043
rect 4403 8038 4518 8039
rect 4403 8034 4496 8038
rect 4500 8034 4501 8038
rect 4505 8034 4518 8038
rect 4403 8033 4518 8034
rect 4403 8029 4496 8033
rect 4500 8029 4501 8033
rect 4505 8029 4518 8033
rect 4403 8028 4518 8029
rect 4403 8024 4496 8028
rect 4500 8024 4501 8028
rect 4505 8024 4518 8028
rect 4095 7747 4253 7752
rect 4266 7796 4322 7801
rect 4095 7685 4100 7747
rect 4094 7684 4100 7685
rect 4094 7680 4095 7684
rect 4099 7680 4100 7684
rect 4094 7679 4100 7680
rect 4266 7622 4271 7796
rect 4220 7617 4271 7622
rect 4403 7793 4518 8024
rect 4403 7789 4479 7793
rect 4483 7789 4489 7793
rect 4493 7789 4499 7793
rect 4503 7789 4509 7793
rect 4513 7789 4518 7793
rect 4403 7788 4518 7789
rect 4403 7784 4479 7788
rect 4483 7784 4489 7788
rect 4493 7784 4499 7788
rect 4503 7784 4509 7788
rect 4513 7784 4518 7788
rect 4403 7783 4518 7784
rect 4403 7779 4479 7783
rect 4483 7779 4489 7783
rect 4493 7779 4499 7783
rect 4503 7779 4509 7783
rect 4513 7779 4518 7783
rect 4403 7778 4518 7779
rect 4403 7774 4479 7778
rect 4483 7774 4489 7778
rect 4493 7774 4499 7778
rect 4503 7774 4509 7778
rect 4513 7774 4518 7778
rect 4220 7603 4225 7617
rect 4219 7602 4225 7603
rect 4219 7598 4220 7602
rect 4224 7598 4225 7602
rect 4219 7597 4225 7598
rect 3020 7413 3775 7418
rect 654 7158 659 7162
rect 663 7158 669 7162
rect 673 7158 679 7162
rect 683 7158 689 7162
rect 693 7158 769 7162
rect 654 7157 769 7158
rect 654 7153 659 7157
rect 663 7153 669 7157
rect 673 7153 679 7157
rect 683 7153 689 7157
rect 693 7153 769 7157
rect 654 7152 769 7153
rect 654 7148 659 7152
rect 663 7148 669 7152
rect 673 7148 679 7152
rect 683 7148 689 7152
rect 693 7148 769 7152
rect 654 7147 769 7148
rect 654 7143 659 7147
rect 663 7143 669 7147
rect 673 7143 679 7147
rect 683 7143 689 7147
rect 693 7143 769 7147
rect 654 6853 769 7143
rect 654 6849 659 6853
rect 663 6849 669 6853
rect 673 6849 679 6853
rect 683 6849 689 6853
rect 693 6849 769 6853
rect 654 6848 769 6849
rect 654 6844 659 6848
rect 663 6844 669 6848
rect 673 6844 679 6848
rect 683 6844 689 6848
rect 693 6844 769 6848
rect 654 6843 769 6844
rect 654 6839 659 6843
rect 663 6839 669 6843
rect 673 6839 679 6843
rect 683 6839 689 6843
rect 693 6839 769 6843
rect 654 6838 769 6839
rect 654 6834 659 6838
rect 663 6834 669 6838
rect 673 6834 679 6838
rect 683 6834 689 6838
rect 693 6834 769 6838
rect 654 6544 769 6834
rect 654 6540 659 6544
rect 663 6540 669 6544
rect 673 6540 679 6544
rect 683 6540 689 6544
rect 693 6540 769 6544
rect 654 6539 769 6540
rect 654 6535 659 6539
rect 663 6535 669 6539
rect 673 6535 679 6539
rect 683 6535 689 6539
rect 693 6535 769 6539
rect 654 6534 769 6535
rect 654 6530 659 6534
rect 663 6530 669 6534
rect 673 6530 679 6534
rect 683 6530 689 6534
rect 693 6530 769 6534
rect 654 6529 769 6530
rect 654 6525 659 6529
rect 663 6525 669 6529
rect 673 6525 679 6529
rect 683 6525 689 6529
rect 693 6525 769 6529
rect 654 6144 769 6525
rect 654 6140 659 6144
rect 663 6140 669 6144
rect 673 6140 679 6144
rect 683 6140 689 6144
rect 693 6140 769 6144
rect 654 6139 769 6140
rect 654 6135 659 6139
rect 663 6135 669 6139
rect 673 6135 679 6139
rect 683 6135 689 6139
rect 693 6135 769 6139
rect 654 6134 769 6135
rect 654 6130 659 6134
rect 663 6130 669 6134
rect 673 6130 679 6134
rect 683 6130 689 6134
rect 693 6130 769 6134
rect 654 6129 769 6130
rect 654 6125 659 6129
rect 663 6125 669 6129
rect 673 6125 679 6129
rect 683 6125 689 6129
rect 693 6125 769 6129
rect 654 6115 769 6125
rect 654 6111 659 6115
rect 663 6111 669 6115
rect 673 6111 679 6115
rect 683 6111 689 6115
rect 693 6111 769 6115
rect 654 6110 769 6111
rect 654 6106 659 6110
rect 663 6106 669 6110
rect 673 6106 679 6110
rect 683 6106 689 6110
rect 693 6106 769 6110
rect 654 6105 769 6106
rect 654 6101 659 6105
rect 663 6101 669 6105
rect 673 6101 679 6105
rect 683 6101 689 6105
rect 693 6101 769 6105
rect 654 6100 769 6101
rect 654 6096 659 6100
rect 663 6096 669 6100
rect 673 6096 679 6100
rect 683 6096 689 6100
rect 693 6096 769 6100
rect 654 6086 769 6096
rect 654 6082 659 6086
rect 663 6082 669 6086
rect 673 6082 679 6086
rect 683 6082 689 6086
rect 693 6082 769 6086
rect 654 6081 769 6082
rect 654 6077 659 6081
rect 663 6077 669 6081
rect 673 6077 679 6081
rect 683 6077 689 6081
rect 693 6077 769 6081
rect 654 6076 769 6077
rect 654 6072 659 6076
rect 663 6072 669 6076
rect 673 6072 679 6076
rect 683 6072 689 6076
rect 693 6072 769 6076
rect 654 6071 769 6072
rect 654 6067 659 6071
rect 663 6067 669 6071
rect 673 6067 679 6071
rect 683 6067 689 6071
rect 693 6067 769 6071
rect 654 6057 769 6067
rect 654 6053 659 6057
rect 663 6053 669 6057
rect 673 6053 679 6057
rect 683 6053 689 6057
rect 693 6053 769 6057
rect 654 6052 769 6053
rect 654 6048 659 6052
rect 663 6048 669 6052
rect 673 6048 679 6052
rect 683 6048 689 6052
rect 693 6048 769 6052
rect 654 6047 769 6048
rect 654 6043 659 6047
rect 663 6043 669 6047
rect 673 6043 679 6047
rect 683 6043 689 6047
rect 693 6043 769 6047
rect 654 6042 769 6043
rect 654 6038 659 6042
rect 663 6038 669 6042
rect 673 6038 679 6042
rect 683 6038 689 6042
rect 693 6038 769 6042
rect 654 6028 769 6038
rect 654 6024 659 6028
rect 663 6024 669 6028
rect 673 6024 679 6028
rect 683 6024 689 6028
rect 693 6024 769 6028
rect 654 6023 769 6024
rect 654 6019 659 6023
rect 663 6019 669 6023
rect 673 6019 679 6023
rect 683 6019 689 6023
rect 693 6019 769 6023
rect 654 6018 769 6019
rect 654 6014 659 6018
rect 663 6014 669 6018
rect 673 6014 679 6018
rect 683 6014 689 6018
rect 693 6014 769 6018
rect 654 6013 769 6014
rect 654 6009 659 6013
rect 663 6009 669 6013
rect 673 6009 679 6013
rect 683 6009 689 6013
rect 693 6009 769 6013
rect 654 5976 769 6009
rect 4403 7206 4518 7774
rect 4403 7202 4479 7206
rect 4483 7202 4489 7206
rect 4493 7202 4499 7206
rect 4503 7202 4509 7206
rect 4513 7202 4518 7206
rect 4403 7201 4518 7202
rect 4403 7197 4479 7201
rect 4483 7197 4489 7201
rect 4493 7197 4499 7201
rect 4503 7197 4509 7201
rect 4513 7197 4518 7201
rect 4403 7196 4518 7197
rect 4403 7192 4479 7196
rect 4483 7192 4489 7196
rect 4493 7192 4499 7196
rect 4503 7192 4509 7196
rect 4513 7192 4518 7196
rect 4403 7191 4518 7192
rect 4403 7187 4479 7191
rect 4483 7187 4489 7191
rect 4493 7187 4499 7191
rect 4503 7187 4509 7191
rect 4513 7187 4518 7191
rect 4403 6897 4518 7187
rect 4403 6893 4479 6897
rect 4483 6893 4489 6897
rect 4493 6893 4499 6897
rect 4503 6893 4509 6897
rect 4513 6893 4518 6897
rect 4403 6892 4518 6893
rect 4403 6888 4479 6892
rect 4483 6888 4489 6892
rect 4493 6888 4499 6892
rect 4503 6888 4509 6892
rect 4513 6888 4518 6892
rect 4403 6887 4518 6888
rect 4403 6883 4479 6887
rect 4483 6883 4489 6887
rect 4493 6883 4499 6887
rect 4503 6883 4509 6887
rect 4513 6883 4518 6887
rect 4403 6882 4518 6883
rect 4403 6878 4479 6882
rect 4483 6878 4489 6882
rect 4493 6878 4499 6882
rect 4503 6878 4509 6882
rect 4513 6878 4518 6882
rect 4403 6588 4518 6878
rect 4403 6584 4479 6588
rect 4483 6584 4489 6588
rect 4493 6584 4499 6588
rect 4503 6584 4509 6588
rect 4513 6584 4518 6588
rect 4403 6583 4518 6584
rect 4403 6579 4479 6583
rect 4483 6579 4489 6583
rect 4493 6579 4499 6583
rect 4503 6579 4509 6583
rect 4513 6579 4518 6583
rect 4403 6578 4518 6579
rect 4403 6574 4479 6578
rect 4483 6574 4489 6578
rect 4493 6574 4499 6578
rect 4503 6574 4509 6578
rect 4513 6574 4518 6578
rect 4403 6573 4518 6574
rect 4403 6569 4479 6573
rect 4483 6569 4489 6573
rect 4493 6569 4499 6573
rect 4503 6569 4509 6573
rect 4513 6569 4518 6573
rect 4403 6279 4518 6569
rect 4403 6275 4479 6279
rect 4483 6275 4489 6279
rect 4493 6275 4499 6279
rect 4503 6275 4509 6279
rect 4513 6275 4518 6279
rect 4403 6274 4518 6275
rect 4403 6270 4479 6274
rect 4483 6270 4489 6274
rect 4493 6270 4499 6274
rect 4503 6270 4509 6274
rect 4513 6270 4518 6274
rect 4403 6269 4518 6270
rect 4403 6265 4479 6269
rect 4483 6265 4489 6269
rect 4493 6265 4499 6269
rect 4503 6265 4509 6269
rect 4513 6265 4518 6269
rect 4403 6264 4518 6265
rect 4403 6260 4479 6264
rect 4483 6260 4489 6264
rect 4493 6260 4499 6264
rect 4503 6260 4509 6264
rect 4513 6260 4518 6264
rect 4403 6087 4518 6260
rect 4403 6083 4479 6087
rect 4483 6083 4489 6087
rect 4493 6083 4499 6087
rect 4503 6083 4509 6087
rect 4513 6083 4518 6087
rect 4403 6082 4518 6083
rect 4403 6078 4479 6082
rect 4483 6078 4489 6082
rect 4493 6078 4499 6082
rect 4503 6078 4509 6082
rect 4513 6078 4518 6082
rect 4403 6077 4518 6078
rect 4403 6073 4479 6077
rect 4483 6073 4489 6077
rect 4493 6073 4499 6077
rect 4503 6073 4509 6077
rect 4513 6073 4518 6077
rect 4403 6072 4518 6073
rect 4403 6068 4479 6072
rect 4483 6068 4489 6072
rect 4493 6068 4499 6072
rect 4503 6068 4509 6072
rect 4513 6068 4518 6072
rect 4403 6061 4518 6068
rect 4403 6057 4479 6061
rect 4483 6057 4489 6061
rect 4493 6057 4499 6061
rect 4503 6057 4509 6061
rect 4513 6057 4518 6061
rect 4403 6056 4518 6057
rect 4403 6052 4479 6056
rect 4483 6052 4489 6056
rect 4493 6052 4499 6056
rect 4503 6052 4509 6056
rect 4513 6052 4518 6056
rect 4403 6051 4518 6052
rect 4403 6047 4479 6051
rect 4483 6047 4489 6051
rect 4493 6047 4499 6051
rect 4503 6047 4509 6051
rect 4513 6047 4518 6051
rect 4403 6046 4518 6047
rect 4403 6042 4479 6046
rect 4483 6042 4489 6046
rect 4493 6042 4499 6046
rect 4503 6042 4509 6046
rect 4513 6042 4518 6046
rect 4403 6035 4518 6042
rect 4403 6031 4479 6035
rect 4483 6031 4489 6035
rect 4493 6031 4499 6035
rect 4503 6031 4509 6035
rect 4513 6031 4518 6035
rect 4403 6030 4518 6031
rect 4403 6026 4479 6030
rect 4483 6026 4489 6030
rect 4493 6026 4499 6030
rect 4503 6026 4509 6030
rect 4513 6026 4518 6030
rect 4403 6025 4518 6026
rect 4403 6021 4479 6025
rect 4483 6021 4489 6025
rect 4493 6021 4499 6025
rect 4503 6021 4509 6025
rect 4513 6021 4518 6025
rect 4403 6020 4518 6021
rect 4403 6016 4479 6020
rect 4483 6016 4489 6020
rect 4493 6016 4499 6020
rect 4503 6016 4509 6020
rect 4513 6016 4518 6020
rect 4403 6009 4518 6016
rect 4403 6005 4479 6009
rect 4483 6005 4489 6009
rect 4493 6005 4499 6009
rect 4503 6005 4509 6009
rect 4513 6005 4518 6009
rect 4403 6004 4518 6005
rect 4403 6000 4479 6004
rect 4483 6000 4489 6004
rect 4493 6000 4499 6004
rect 4503 6000 4509 6004
rect 4513 6000 4518 6004
rect 4403 5999 4518 6000
rect 4403 5995 4479 5999
rect 4483 5995 4489 5999
rect 4493 5995 4499 5999
rect 4503 5995 4509 5999
rect 4513 5995 4518 5999
rect 4403 5994 4518 5995
rect 4403 5990 4479 5994
rect 4483 5990 4489 5994
rect 4493 5990 4499 5994
rect 4503 5990 4509 5994
rect 4513 5990 4518 5994
rect 4403 5983 4518 5990
rect 4403 5979 4479 5983
rect 4483 5979 4489 5983
rect 4493 5979 4499 5983
rect 4503 5979 4509 5983
rect 4513 5979 4518 5983
rect 4403 5978 4518 5979
rect 4403 5976 4479 5978
rect 654 5974 4479 5976
rect 4483 5974 4489 5978
rect 4493 5974 4499 5978
rect 4503 5974 4509 5978
rect 4513 5974 4518 5978
rect 654 5973 4518 5974
rect 654 5969 4479 5973
rect 4483 5969 4489 5973
rect 4493 5969 4499 5973
rect 4503 5969 4509 5973
rect 4513 5969 4518 5973
rect 654 5968 4518 5969
rect 654 5964 4479 5968
rect 4483 5964 4489 5968
rect 4493 5964 4499 5968
rect 4503 5964 4509 5968
rect 4513 5964 4518 5968
rect 654 5900 4518 5964
rect 654 5896 757 5900
rect 761 5896 762 5900
rect 766 5896 767 5900
rect 771 5896 772 5900
rect 776 5896 783 5900
rect 787 5896 788 5900
rect 792 5896 793 5900
rect 797 5896 798 5900
rect 802 5896 809 5900
rect 813 5896 814 5900
rect 818 5896 819 5900
rect 823 5896 824 5900
rect 828 5896 835 5900
rect 839 5896 840 5900
rect 844 5896 845 5900
rect 849 5896 850 5900
rect 854 5896 861 5900
rect 865 5896 866 5900
rect 870 5896 871 5900
rect 875 5896 876 5900
rect 880 5896 1054 5900
rect 1058 5896 1059 5900
rect 1063 5896 1064 5900
rect 1068 5896 1069 5900
rect 1073 5896 1363 5900
rect 1367 5896 1368 5900
rect 1372 5896 1373 5900
rect 1377 5896 1378 5900
rect 1382 5896 1672 5900
rect 1676 5896 1677 5900
rect 1681 5896 1682 5900
rect 1686 5896 1687 5900
rect 1691 5896 1981 5900
rect 1985 5896 1986 5900
rect 1990 5896 1991 5900
rect 1995 5896 1996 5900
rect 2000 5896 2290 5900
rect 2294 5896 2295 5900
rect 2299 5896 2300 5900
rect 2304 5896 2305 5900
rect 2309 5896 2599 5900
rect 2603 5896 2604 5900
rect 2608 5896 2609 5900
rect 2613 5896 2614 5900
rect 2618 5896 2908 5900
rect 2912 5896 2913 5900
rect 2917 5896 2918 5900
rect 2922 5896 2923 5900
rect 2927 5896 3217 5900
rect 3221 5896 3222 5900
rect 3226 5896 3227 5900
rect 3231 5896 3232 5900
rect 3236 5896 3526 5900
rect 3530 5896 3531 5900
rect 3535 5896 3536 5900
rect 3540 5896 3541 5900
rect 3545 5896 3835 5900
rect 3839 5896 3840 5900
rect 3844 5896 3845 5900
rect 3849 5896 3850 5900
rect 3854 5896 4235 5900
rect 4239 5896 4240 5900
rect 4244 5896 4245 5900
rect 4249 5896 4250 5900
rect 4254 5896 4264 5900
rect 4268 5896 4269 5900
rect 4273 5896 4274 5900
rect 4278 5896 4279 5900
rect 4283 5896 4293 5900
rect 4297 5896 4298 5900
rect 4302 5896 4303 5900
rect 4307 5896 4308 5900
rect 4312 5896 4322 5900
rect 4326 5896 4327 5900
rect 4331 5896 4332 5900
rect 4336 5896 4337 5900
rect 4341 5896 4351 5900
rect 4355 5896 4356 5900
rect 4360 5896 4361 5900
rect 4365 5896 4366 5900
rect 4370 5896 4518 5900
rect 654 5890 4518 5896
rect 654 5886 757 5890
rect 761 5886 762 5890
rect 766 5886 767 5890
rect 771 5886 772 5890
rect 776 5886 783 5890
rect 787 5886 788 5890
rect 792 5886 793 5890
rect 797 5886 798 5890
rect 802 5886 809 5890
rect 813 5886 814 5890
rect 818 5886 819 5890
rect 823 5886 824 5890
rect 828 5886 835 5890
rect 839 5886 840 5890
rect 844 5886 845 5890
rect 849 5886 850 5890
rect 854 5886 861 5890
rect 865 5886 866 5890
rect 870 5886 871 5890
rect 875 5886 876 5890
rect 880 5886 1054 5890
rect 1058 5886 1059 5890
rect 1063 5886 1064 5890
rect 1068 5886 1069 5890
rect 1073 5886 1363 5890
rect 1367 5886 1368 5890
rect 1372 5886 1373 5890
rect 1377 5886 1378 5890
rect 1382 5886 1672 5890
rect 1676 5886 1677 5890
rect 1681 5886 1682 5890
rect 1686 5886 1687 5890
rect 1691 5886 1981 5890
rect 1985 5886 1986 5890
rect 1990 5886 1991 5890
rect 1995 5886 1996 5890
rect 2000 5886 2290 5890
rect 2294 5886 2295 5890
rect 2299 5886 2300 5890
rect 2304 5886 2305 5890
rect 2309 5886 2599 5890
rect 2603 5886 2604 5890
rect 2608 5886 2609 5890
rect 2613 5886 2614 5890
rect 2618 5886 2908 5890
rect 2912 5886 2913 5890
rect 2917 5886 2918 5890
rect 2922 5886 2923 5890
rect 2927 5886 3217 5890
rect 3221 5886 3222 5890
rect 3226 5886 3227 5890
rect 3231 5886 3232 5890
rect 3236 5886 3526 5890
rect 3530 5886 3531 5890
rect 3535 5886 3536 5890
rect 3540 5886 3541 5890
rect 3545 5886 3835 5890
rect 3839 5886 3840 5890
rect 3844 5886 3845 5890
rect 3849 5886 3850 5890
rect 3854 5886 4235 5890
rect 4239 5886 4240 5890
rect 4244 5886 4245 5890
rect 4249 5886 4250 5890
rect 4254 5886 4264 5890
rect 4268 5886 4269 5890
rect 4273 5886 4274 5890
rect 4278 5886 4279 5890
rect 4283 5886 4293 5890
rect 4297 5886 4298 5890
rect 4302 5886 4303 5890
rect 4307 5886 4308 5890
rect 4312 5886 4322 5890
rect 4326 5886 4327 5890
rect 4331 5886 4332 5890
rect 4336 5886 4337 5890
rect 4341 5886 4351 5890
rect 4355 5886 4356 5890
rect 4360 5886 4361 5890
rect 4365 5886 4366 5890
rect 4370 5886 4518 5890
rect 654 5880 4518 5886
rect 654 5876 757 5880
rect 761 5876 762 5880
rect 766 5876 767 5880
rect 771 5876 772 5880
rect 776 5876 783 5880
rect 787 5876 788 5880
rect 792 5876 793 5880
rect 797 5876 798 5880
rect 802 5876 809 5880
rect 813 5876 814 5880
rect 818 5876 819 5880
rect 823 5876 824 5880
rect 828 5876 835 5880
rect 839 5876 840 5880
rect 844 5876 845 5880
rect 849 5876 850 5880
rect 854 5876 861 5880
rect 865 5876 866 5880
rect 870 5876 871 5880
rect 875 5876 876 5880
rect 880 5876 1054 5880
rect 1058 5876 1059 5880
rect 1063 5876 1064 5880
rect 1068 5876 1069 5880
rect 1073 5876 1363 5880
rect 1367 5876 1368 5880
rect 1372 5876 1373 5880
rect 1377 5876 1378 5880
rect 1382 5876 1672 5880
rect 1676 5876 1677 5880
rect 1681 5876 1682 5880
rect 1686 5876 1687 5880
rect 1691 5876 1981 5880
rect 1985 5876 1986 5880
rect 1990 5876 1991 5880
rect 1995 5876 1996 5880
rect 2000 5876 2290 5880
rect 2294 5876 2295 5880
rect 2299 5876 2300 5880
rect 2304 5876 2305 5880
rect 2309 5876 2599 5880
rect 2603 5876 2604 5880
rect 2608 5876 2609 5880
rect 2613 5876 2614 5880
rect 2618 5876 2908 5880
rect 2912 5876 2913 5880
rect 2917 5876 2918 5880
rect 2922 5876 2923 5880
rect 2927 5876 3217 5880
rect 3221 5876 3222 5880
rect 3226 5876 3227 5880
rect 3231 5876 3232 5880
rect 3236 5876 3526 5880
rect 3530 5876 3531 5880
rect 3535 5876 3536 5880
rect 3540 5876 3541 5880
rect 3545 5876 3835 5880
rect 3839 5876 3840 5880
rect 3844 5876 3845 5880
rect 3849 5876 3850 5880
rect 3854 5876 4235 5880
rect 4239 5876 4240 5880
rect 4244 5876 4245 5880
rect 4249 5876 4250 5880
rect 4254 5876 4264 5880
rect 4268 5876 4269 5880
rect 4273 5876 4274 5880
rect 4278 5876 4279 5880
rect 4283 5876 4293 5880
rect 4297 5876 4298 5880
rect 4302 5876 4303 5880
rect 4307 5876 4308 5880
rect 4312 5876 4322 5880
rect 4326 5876 4327 5880
rect 4331 5876 4332 5880
rect 4336 5876 4337 5880
rect 4341 5876 4351 5880
rect 4355 5876 4356 5880
rect 4360 5876 4361 5880
rect 4365 5876 4366 5880
rect 4370 5876 4518 5880
rect 654 5870 4518 5876
rect 654 5866 757 5870
rect 761 5866 762 5870
rect 766 5866 767 5870
rect 771 5866 772 5870
rect 776 5866 783 5870
rect 787 5866 788 5870
rect 792 5866 793 5870
rect 797 5866 798 5870
rect 802 5866 809 5870
rect 813 5866 814 5870
rect 818 5866 819 5870
rect 823 5866 824 5870
rect 828 5866 835 5870
rect 839 5866 840 5870
rect 844 5866 845 5870
rect 849 5866 850 5870
rect 854 5866 861 5870
rect 865 5866 866 5870
rect 870 5866 871 5870
rect 875 5866 876 5870
rect 880 5866 1054 5870
rect 1058 5866 1059 5870
rect 1063 5866 1064 5870
rect 1068 5866 1069 5870
rect 1073 5866 1363 5870
rect 1367 5866 1368 5870
rect 1372 5866 1373 5870
rect 1377 5866 1378 5870
rect 1382 5866 1672 5870
rect 1676 5866 1677 5870
rect 1681 5866 1682 5870
rect 1686 5866 1687 5870
rect 1691 5866 1981 5870
rect 1985 5866 1986 5870
rect 1990 5866 1991 5870
rect 1995 5866 1996 5870
rect 2000 5866 2290 5870
rect 2294 5866 2295 5870
rect 2299 5866 2300 5870
rect 2304 5866 2305 5870
rect 2309 5866 2599 5870
rect 2603 5866 2604 5870
rect 2608 5866 2609 5870
rect 2613 5866 2614 5870
rect 2618 5866 2908 5870
rect 2912 5866 2913 5870
rect 2917 5866 2918 5870
rect 2922 5866 2923 5870
rect 2927 5866 3217 5870
rect 3221 5866 3222 5870
rect 3226 5866 3227 5870
rect 3231 5866 3232 5870
rect 3236 5866 3526 5870
rect 3530 5866 3531 5870
rect 3535 5866 3536 5870
rect 3540 5866 3541 5870
rect 3545 5866 3835 5870
rect 3839 5866 3840 5870
rect 3844 5866 3845 5870
rect 3849 5866 3850 5870
rect 3854 5866 4235 5870
rect 4239 5866 4240 5870
rect 4244 5866 4245 5870
rect 4249 5866 4250 5870
rect 4254 5866 4264 5870
rect 4268 5866 4269 5870
rect 4273 5866 4274 5870
rect 4278 5866 4279 5870
rect 4283 5866 4293 5870
rect 4297 5866 4298 5870
rect 4302 5866 4303 5870
rect 4307 5866 4308 5870
rect 4312 5866 4322 5870
rect 4326 5866 4327 5870
rect 4331 5866 4332 5870
rect 4336 5866 4337 5870
rect 4341 5866 4351 5870
rect 4355 5866 4356 5870
rect 4360 5866 4361 5870
rect 4365 5866 4366 5870
rect 4370 5866 4518 5870
rect 654 5861 4518 5866
rect 4522 9577 4602 9729
rect 4522 9573 4525 9577
rect 4529 9573 4535 9577
rect 4539 9573 4545 9577
rect 4549 9573 4555 9577
rect 4559 9573 4602 9577
rect 4522 9572 4602 9573
rect 4522 9568 4525 9572
rect 4529 9568 4535 9572
rect 4539 9568 4545 9572
rect 4549 9568 4555 9572
rect 4559 9568 4602 9572
rect 4522 9567 4602 9568
rect 4522 9563 4525 9567
rect 4529 9563 4535 9567
rect 4539 9563 4545 9567
rect 4549 9563 4555 9567
rect 4559 9563 4602 9567
rect 4522 9562 4602 9563
rect 4522 9558 4525 9562
rect 4529 9558 4535 9562
rect 4539 9558 4545 9562
rect 4549 9558 4555 9562
rect 4559 9558 4602 9562
rect 4522 9548 4602 9558
rect 4522 9544 4525 9548
rect 4529 9544 4535 9548
rect 4539 9544 4545 9548
rect 4549 9544 4555 9548
rect 4559 9544 4602 9548
rect 4522 9543 4602 9544
rect 4522 9539 4525 9543
rect 4529 9539 4535 9543
rect 4539 9539 4545 9543
rect 4549 9539 4555 9543
rect 4559 9539 4602 9543
rect 4522 9538 4602 9539
rect 4522 9534 4525 9538
rect 4529 9534 4535 9538
rect 4539 9534 4545 9538
rect 4549 9534 4555 9538
rect 4559 9534 4602 9538
rect 4522 9533 4602 9534
rect 4522 9529 4525 9533
rect 4529 9529 4535 9533
rect 4539 9529 4545 9533
rect 4549 9529 4555 9533
rect 4559 9529 4602 9533
rect 4522 9519 4602 9529
rect 4522 9515 4525 9519
rect 4529 9515 4535 9519
rect 4539 9515 4545 9519
rect 4549 9515 4555 9519
rect 4559 9515 4602 9519
rect 4522 9514 4602 9515
rect 4522 9510 4525 9514
rect 4529 9510 4535 9514
rect 4539 9510 4545 9514
rect 4549 9510 4555 9514
rect 4559 9510 4602 9514
rect 4522 9509 4602 9510
rect 4522 9505 4525 9509
rect 4529 9505 4535 9509
rect 4539 9505 4545 9509
rect 4549 9505 4555 9509
rect 4559 9505 4602 9509
rect 4522 9504 4602 9505
rect 4522 9500 4525 9504
rect 4529 9500 4535 9504
rect 4539 9500 4545 9504
rect 4549 9500 4555 9504
rect 4559 9500 4602 9504
rect 4522 9490 4602 9500
rect 4522 9486 4525 9490
rect 4529 9486 4535 9490
rect 4539 9486 4545 9490
rect 4549 9486 4555 9490
rect 4559 9486 4602 9490
rect 4522 9485 4602 9486
rect 4522 9481 4525 9485
rect 4529 9481 4535 9485
rect 4539 9481 4545 9485
rect 4549 9481 4555 9485
rect 4559 9481 4602 9485
rect 4522 9480 4602 9481
rect 4522 9476 4525 9480
rect 4529 9476 4535 9480
rect 4539 9476 4545 9480
rect 4549 9476 4555 9480
rect 4559 9476 4602 9480
rect 4522 9475 4602 9476
rect 4522 9471 4525 9475
rect 4529 9471 4535 9475
rect 4539 9471 4545 9475
rect 4549 9471 4555 9475
rect 4559 9471 4602 9475
rect 4522 9461 4602 9471
rect 4522 9457 4525 9461
rect 4529 9457 4535 9461
rect 4539 9457 4545 9461
rect 4549 9457 4555 9461
rect 4559 9457 4602 9461
rect 4522 9456 4602 9457
rect 4522 9452 4525 9456
rect 4529 9452 4535 9456
rect 4539 9452 4545 9456
rect 4549 9452 4555 9456
rect 4559 9452 4602 9456
rect 4522 9451 4602 9452
rect 4522 9447 4525 9451
rect 4529 9447 4535 9451
rect 4539 9447 4545 9451
rect 4549 9447 4555 9451
rect 4559 9447 4602 9451
rect 4522 9446 4602 9447
rect 4522 9442 4525 9446
rect 4529 9442 4535 9446
rect 4539 9442 4545 9446
rect 4549 9442 4555 9446
rect 4559 9442 4602 9446
rect 4522 9060 4602 9442
rect 4522 9056 4525 9060
rect 4529 9056 4535 9060
rect 4539 9056 4545 9060
rect 4549 9056 4555 9060
rect 4559 9056 4602 9060
rect 4522 9055 4602 9056
rect 4522 9051 4525 9055
rect 4529 9051 4535 9055
rect 4539 9051 4545 9055
rect 4549 9051 4555 9055
rect 4559 9051 4602 9055
rect 4522 9050 4602 9051
rect 4522 9046 4525 9050
rect 4529 9046 4535 9050
rect 4539 9046 4545 9050
rect 4549 9046 4555 9050
rect 4559 9046 4602 9050
rect 4522 9045 4602 9046
rect 4522 9041 4525 9045
rect 4529 9041 4535 9045
rect 4539 9041 4545 9045
rect 4549 9041 4555 9045
rect 4559 9041 4602 9045
rect 4522 8751 4602 9041
rect 4522 8747 4525 8751
rect 4529 8747 4535 8751
rect 4539 8747 4545 8751
rect 4549 8747 4555 8751
rect 4559 8747 4602 8751
rect 4522 8746 4602 8747
rect 4522 8742 4525 8746
rect 4529 8742 4535 8746
rect 4539 8742 4545 8746
rect 4549 8742 4555 8746
rect 4559 8742 4602 8746
rect 4522 8741 4602 8742
rect 4522 8737 4525 8741
rect 4529 8737 4535 8741
rect 4539 8737 4545 8741
rect 4549 8737 4555 8741
rect 4559 8737 4602 8741
rect 4522 8736 4602 8737
rect 4522 8732 4525 8736
rect 4529 8732 4535 8736
rect 4539 8732 4545 8736
rect 4549 8732 4555 8736
rect 4559 8732 4602 8736
rect 4522 8442 4602 8732
rect 4522 8438 4525 8442
rect 4529 8438 4535 8442
rect 4539 8438 4545 8442
rect 4549 8438 4555 8442
rect 4559 8438 4602 8442
rect 4522 8437 4602 8438
rect 4522 8433 4525 8437
rect 4529 8433 4535 8437
rect 4539 8433 4545 8437
rect 4549 8433 4555 8437
rect 4559 8433 4602 8437
rect 4522 8432 4602 8433
rect 4522 8428 4525 8432
rect 4529 8428 4535 8432
rect 4539 8428 4545 8432
rect 4549 8428 4555 8432
rect 4559 8428 4602 8432
rect 4522 8427 4602 8428
rect 4522 8423 4525 8427
rect 4529 8423 4535 8427
rect 4539 8423 4545 8427
rect 4549 8423 4555 8427
rect 4559 8423 4602 8427
rect 4522 8133 4602 8423
rect 4522 8129 4525 8133
rect 4529 8129 4535 8133
rect 4539 8129 4545 8133
rect 4549 8129 4555 8133
rect 4559 8129 4602 8133
rect 4522 8128 4602 8129
rect 4522 8124 4525 8128
rect 4529 8124 4535 8128
rect 4539 8124 4545 8128
rect 4549 8124 4555 8128
rect 4559 8124 4602 8128
rect 4522 8123 4602 8124
rect 4522 8119 4525 8123
rect 4529 8119 4535 8123
rect 4539 8119 4545 8123
rect 4549 8119 4555 8123
rect 4559 8119 4602 8123
rect 4522 8118 4602 8119
rect 4522 8114 4525 8118
rect 4529 8114 4535 8118
rect 4539 8114 4545 8118
rect 4549 8114 4555 8118
rect 4559 8114 4602 8118
rect 4522 8102 4602 8114
rect 4522 8098 4525 8102
rect 4529 8098 4535 8102
rect 4539 8098 4545 8102
rect 4549 8098 4555 8102
rect 4559 8098 4602 8102
rect 4522 8097 4602 8098
rect 4522 8093 4525 8097
rect 4529 8093 4535 8097
rect 4539 8093 4545 8097
rect 4549 8093 4555 8097
rect 4559 8093 4602 8097
rect 4522 8092 4602 8093
rect 4522 8088 4525 8092
rect 4529 8088 4535 8092
rect 4539 8088 4545 8092
rect 4549 8088 4555 8092
rect 4559 8088 4602 8092
rect 4522 8087 4602 8088
rect 4522 8083 4525 8087
rect 4529 8083 4535 8087
rect 4539 8083 4545 8087
rect 4549 8083 4555 8087
rect 4559 8083 4602 8087
rect 4522 7818 4602 8083
rect 4522 7814 4529 7818
rect 4533 7814 4534 7818
rect 4538 7814 4539 7818
rect 4543 7814 4544 7818
rect 4548 7814 4549 7818
rect 4553 7814 4554 7818
rect 4558 7814 4559 7818
rect 4563 7814 4564 7818
rect 4568 7814 4569 7818
rect 4573 7814 4574 7818
rect 4578 7814 4579 7818
rect 4583 7814 4584 7818
rect 4588 7814 4589 7818
rect 4593 7814 4602 7818
rect 4522 7813 4602 7814
rect 4522 7809 4529 7813
rect 4533 7809 4534 7813
rect 4538 7809 4539 7813
rect 4543 7809 4544 7813
rect 4548 7809 4549 7813
rect 4553 7809 4554 7813
rect 4558 7809 4559 7813
rect 4563 7809 4564 7813
rect 4568 7809 4569 7813
rect 4573 7809 4574 7813
rect 4578 7809 4579 7813
rect 4583 7809 4584 7813
rect 4588 7809 4589 7813
rect 4593 7809 4602 7813
rect 4522 7793 4602 7809
rect 4522 7789 4525 7793
rect 4529 7789 4535 7793
rect 4539 7789 4545 7793
rect 4549 7789 4555 7793
rect 4559 7789 4602 7793
rect 4522 7788 4602 7789
rect 4522 7784 4525 7788
rect 4529 7784 4535 7788
rect 4539 7784 4545 7788
rect 4549 7784 4555 7788
rect 4559 7784 4602 7788
rect 4522 7783 4602 7784
rect 4522 7779 4525 7783
rect 4529 7779 4535 7783
rect 4539 7779 4545 7783
rect 4549 7779 4555 7783
rect 4559 7779 4602 7783
rect 4522 7778 4602 7779
rect 4522 7774 4525 7778
rect 4529 7774 4535 7778
rect 4539 7774 4545 7778
rect 4549 7774 4555 7778
rect 4559 7774 4602 7778
rect 4522 7206 4602 7774
rect 4522 7202 4525 7206
rect 4529 7202 4535 7206
rect 4539 7202 4545 7206
rect 4549 7202 4555 7206
rect 4559 7202 4602 7206
rect 4522 7201 4602 7202
rect 4522 7197 4525 7201
rect 4529 7197 4535 7201
rect 4539 7197 4545 7201
rect 4549 7197 4555 7201
rect 4559 7197 4602 7201
rect 4522 7196 4602 7197
rect 4522 7192 4525 7196
rect 4529 7192 4535 7196
rect 4539 7192 4545 7196
rect 4549 7192 4555 7196
rect 4559 7192 4602 7196
rect 4522 7191 4602 7192
rect 4522 7187 4525 7191
rect 4529 7187 4535 7191
rect 4539 7187 4545 7191
rect 4549 7187 4555 7191
rect 4559 7187 4602 7191
rect 4522 6897 4602 7187
rect 4522 6893 4525 6897
rect 4529 6893 4535 6897
rect 4539 6893 4545 6897
rect 4549 6893 4555 6897
rect 4559 6893 4602 6897
rect 4522 6892 4602 6893
rect 4522 6888 4525 6892
rect 4529 6888 4535 6892
rect 4539 6888 4545 6892
rect 4549 6888 4555 6892
rect 4559 6888 4602 6892
rect 4522 6887 4602 6888
rect 4522 6883 4525 6887
rect 4529 6883 4535 6887
rect 4539 6883 4545 6887
rect 4549 6883 4555 6887
rect 4559 6883 4602 6887
rect 4522 6882 4602 6883
rect 4522 6878 4525 6882
rect 4529 6878 4535 6882
rect 4539 6878 4545 6882
rect 4549 6878 4555 6882
rect 4559 6878 4602 6882
rect 4522 6588 4602 6878
rect 4522 6584 4525 6588
rect 4529 6584 4535 6588
rect 4539 6584 4545 6588
rect 4549 6584 4555 6588
rect 4559 6584 4602 6588
rect 4522 6583 4602 6584
rect 4522 6579 4525 6583
rect 4529 6579 4535 6583
rect 4539 6579 4545 6583
rect 4549 6579 4555 6583
rect 4559 6579 4602 6583
rect 4522 6578 4602 6579
rect 4522 6574 4525 6578
rect 4529 6574 4535 6578
rect 4539 6574 4545 6578
rect 4549 6574 4555 6578
rect 4559 6574 4602 6578
rect 4522 6573 4602 6574
rect 4522 6569 4525 6573
rect 4529 6569 4535 6573
rect 4539 6569 4545 6573
rect 4549 6569 4555 6573
rect 4559 6569 4602 6573
rect 4522 6279 4602 6569
rect 4522 6275 4525 6279
rect 4529 6275 4535 6279
rect 4539 6275 4545 6279
rect 4549 6275 4555 6279
rect 4559 6275 4602 6279
rect 4522 6274 4602 6275
rect 4522 6270 4525 6274
rect 4529 6270 4535 6274
rect 4539 6270 4545 6274
rect 4549 6270 4555 6274
rect 4559 6270 4602 6274
rect 4522 6269 4602 6270
rect 4522 6265 4525 6269
rect 4529 6265 4535 6269
rect 4539 6265 4545 6269
rect 4549 6265 4555 6269
rect 4559 6265 4602 6269
rect 4522 6264 4602 6265
rect 4522 6260 4525 6264
rect 4529 6260 4535 6264
rect 4539 6260 4545 6264
rect 4549 6260 4555 6264
rect 4559 6260 4602 6264
rect 4522 6087 4602 6260
rect 4522 6083 4525 6087
rect 4529 6083 4535 6087
rect 4539 6083 4545 6087
rect 4549 6083 4555 6087
rect 4559 6083 4602 6087
rect 4522 6082 4602 6083
rect 4522 6078 4525 6082
rect 4529 6078 4535 6082
rect 4539 6078 4545 6082
rect 4549 6078 4555 6082
rect 4559 6078 4602 6082
rect 4522 6077 4602 6078
rect 4522 6073 4525 6077
rect 4529 6073 4535 6077
rect 4539 6073 4545 6077
rect 4549 6073 4555 6077
rect 4559 6073 4602 6077
rect 4522 6072 4602 6073
rect 4522 6068 4525 6072
rect 4529 6068 4535 6072
rect 4539 6068 4545 6072
rect 4549 6068 4555 6072
rect 4559 6068 4602 6072
rect 4522 6061 4602 6068
rect 4522 6057 4525 6061
rect 4529 6057 4535 6061
rect 4539 6057 4545 6061
rect 4549 6057 4555 6061
rect 4559 6057 4602 6061
rect 4522 6056 4602 6057
rect 4522 6052 4525 6056
rect 4529 6052 4535 6056
rect 4539 6052 4545 6056
rect 4549 6052 4555 6056
rect 4559 6052 4602 6056
rect 4522 6051 4602 6052
rect 4522 6047 4525 6051
rect 4529 6047 4535 6051
rect 4539 6047 4545 6051
rect 4549 6047 4555 6051
rect 4559 6047 4602 6051
rect 4522 6046 4602 6047
rect 4522 6042 4525 6046
rect 4529 6042 4535 6046
rect 4539 6042 4545 6046
rect 4549 6042 4555 6046
rect 4559 6042 4602 6046
rect 4522 6035 4602 6042
rect 4522 6031 4525 6035
rect 4529 6031 4535 6035
rect 4539 6031 4545 6035
rect 4549 6031 4555 6035
rect 4559 6031 4602 6035
rect 4522 6030 4602 6031
rect 4522 6026 4525 6030
rect 4529 6026 4535 6030
rect 4539 6026 4545 6030
rect 4549 6026 4555 6030
rect 4559 6026 4602 6030
rect 4522 6025 4602 6026
rect 4522 6021 4525 6025
rect 4529 6021 4535 6025
rect 4539 6021 4545 6025
rect 4549 6021 4555 6025
rect 4559 6021 4602 6025
rect 4522 6020 4602 6021
rect 4522 6016 4525 6020
rect 4529 6016 4535 6020
rect 4539 6016 4545 6020
rect 4549 6016 4555 6020
rect 4559 6016 4602 6020
rect 4522 6009 4602 6016
rect 4522 6005 4525 6009
rect 4529 6005 4535 6009
rect 4539 6005 4545 6009
rect 4549 6005 4555 6009
rect 4559 6005 4602 6009
rect 4522 6004 4602 6005
rect 4522 6000 4525 6004
rect 4529 6000 4535 6004
rect 4539 6000 4545 6004
rect 4549 6000 4555 6004
rect 4559 6000 4602 6004
rect 4522 5999 4602 6000
rect 4522 5995 4525 5999
rect 4529 5995 4535 5999
rect 4539 5995 4545 5999
rect 4549 5995 4555 5999
rect 4559 5995 4602 5999
rect 4522 5994 4602 5995
rect 4522 5990 4525 5994
rect 4529 5990 4535 5994
rect 4539 5990 4545 5994
rect 4549 5990 4555 5994
rect 4559 5990 4602 5994
rect 4522 5983 4602 5990
rect 4522 5979 4525 5983
rect 4529 5979 4535 5983
rect 4539 5979 4545 5983
rect 4549 5979 4555 5983
rect 4559 5979 4602 5983
rect 4522 5978 4602 5979
rect 4522 5974 4525 5978
rect 4529 5974 4535 5978
rect 4539 5974 4545 5978
rect 4549 5974 4555 5978
rect 4559 5974 4602 5978
rect 4522 5973 4602 5974
rect 4522 5969 4525 5973
rect 4529 5969 4535 5973
rect 4539 5969 4545 5973
rect 4549 5969 4555 5973
rect 4559 5969 4602 5973
rect 4522 5968 4602 5969
rect 4522 5964 4525 5968
rect 4529 5964 4535 5968
rect 4539 5964 4545 5968
rect 4549 5964 4555 5968
rect 4559 5964 4602 5968
rect 4522 5857 4602 5964
rect 570 5854 4602 5857
rect 570 5850 757 5854
rect 761 5850 762 5854
rect 766 5850 767 5854
rect 771 5850 772 5854
rect 776 5850 783 5854
rect 787 5850 788 5854
rect 792 5850 793 5854
rect 797 5850 798 5854
rect 802 5850 809 5854
rect 813 5850 814 5854
rect 818 5850 819 5854
rect 823 5850 824 5854
rect 828 5850 835 5854
rect 839 5850 840 5854
rect 844 5850 845 5854
rect 849 5850 850 5854
rect 854 5850 861 5854
rect 865 5850 866 5854
rect 870 5850 871 5854
rect 875 5850 876 5854
rect 880 5850 1054 5854
rect 1058 5850 1059 5854
rect 1063 5850 1064 5854
rect 1068 5850 1069 5854
rect 1073 5850 1363 5854
rect 1367 5850 1368 5854
rect 1372 5850 1373 5854
rect 1377 5850 1378 5854
rect 1382 5850 1672 5854
rect 1676 5850 1677 5854
rect 1681 5850 1682 5854
rect 1686 5850 1687 5854
rect 1691 5850 1981 5854
rect 1985 5850 1986 5854
rect 1990 5850 1991 5854
rect 1995 5850 1996 5854
rect 2000 5850 2290 5854
rect 2294 5850 2295 5854
rect 2299 5850 2300 5854
rect 2304 5850 2305 5854
rect 2309 5850 2599 5854
rect 2603 5850 2604 5854
rect 2608 5850 2609 5854
rect 2613 5850 2614 5854
rect 2618 5850 2908 5854
rect 2912 5850 2913 5854
rect 2917 5850 2918 5854
rect 2922 5850 2923 5854
rect 2927 5850 3217 5854
rect 3221 5850 3222 5854
rect 3226 5850 3227 5854
rect 3231 5850 3232 5854
rect 3236 5850 3526 5854
rect 3530 5850 3531 5854
rect 3535 5850 3536 5854
rect 3540 5850 3541 5854
rect 3545 5850 3835 5854
rect 3839 5850 3840 5854
rect 3844 5850 3845 5854
rect 3849 5850 3850 5854
rect 3854 5850 4235 5854
rect 4239 5850 4240 5854
rect 4244 5850 4245 5854
rect 4249 5850 4250 5854
rect 4254 5850 4264 5854
rect 4268 5850 4269 5854
rect 4273 5850 4274 5854
rect 4278 5850 4279 5854
rect 4283 5850 4293 5854
rect 4297 5850 4298 5854
rect 4302 5850 4303 5854
rect 4307 5850 4308 5854
rect 4312 5850 4322 5854
rect 4326 5850 4327 5854
rect 4331 5850 4332 5854
rect 4336 5850 4337 5854
rect 4341 5850 4351 5854
rect 4355 5850 4356 5854
rect 4360 5850 4361 5854
rect 4365 5850 4366 5854
rect 4370 5850 4602 5854
rect 570 5844 4602 5850
rect 570 5840 757 5844
rect 761 5840 762 5844
rect 766 5840 767 5844
rect 771 5840 772 5844
rect 776 5840 783 5844
rect 787 5840 788 5844
rect 792 5840 793 5844
rect 797 5840 798 5844
rect 802 5840 809 5844
rect 813 5840 814 5844
rect 818 5840 819 5844
rect 823 5840 824 5844
rect 828 5840 835 5844
rect 839 5840 840 5844
rect 844 5840 845 5844
rect 849 5840 850 5844
rect 854 5840 861 5844
rect 865 5840 866 5844
rect 870 5840 871 5844
rect 875 5840 876 5844
rect 880 5840 1054 5844
rect 1058 5840 1059 5844
rect 1063 5840 1064 5844
rect 1068 5840 1069 5844
rect 1073 5840 1363 5844
rect 1367 5840 1368 5844
rect 1372 5840 1373 5844
rect 1377 5840 1378 5844
rect 1382 5840 1672 5844
rect 1676 5840 1677 5844
rect 1681 5840 1682 5844
rect 1686 5840 1687 5844
rect 1691 5840 1981 5844
rect 1985 5840 1986 5844
rect 1990 5840 1991 5844
rect 1995 5840 1996 5844
rect 2000 5840 2290 5844
rect 2294 5840 2295 5844
rect 2299 5840 2300 5844
rect 2304 5840 2305 5844
rect 2309 5840 2599 5844
rect 2603 5840 2604 5844
rect 2608 5840 2609 5844
rect 2613 5840 2614 5844
rect 2618 5840 2908 5844
rect 2912 5840 2913 5844
rect 2917 5840 2918 5844
rect 2922 5840 2923 5844
rect 2927 5840 3217 5844
rect 3221 5840 3222 5844
rect 3226 5840 3227 5844
rect 3231 5840 3232 5844
rect 3236 5840 3526 5844
rect 3530 5840 3531 5844
rect 3535 5840 3536 5844
rect 3540 5840 3541 5844
rect 3545 5840 3835 5844
rect 3839 5840 3840 5844
rect 3844 5840 3845 5844
rect 3849 5840 3850 5844
rect 3854 5840 4235 5844
rect 4239 5840 4240 5844
rect 4244 5840 4245 5844
rect 4249 5840 4250 5844
rect 4254 5840 4264 5844
rect 4268 5840 4269 5844
rect 4273 5840 4274 5844
rect 4278 5840 4279 5844
rect 4283 5840 4293 5844
rect 4297 5840 4298 5844
rect 4302 5840 4303 5844
rect 4307 5840 4308 5844
rect 4312 5840 4322 5844
rect 4326 5840 4327 5844
rect 4331 5840 4332 5844
rect 4336 5840 4337 5844
rect 4341 5840 4351 5844
rect 4355 5840 4356 5844
rect 4360 5840 4361 5844
rect 4365 5840 4366 5844
rect 4370 5840 4602 5844
rect 570 5834 4602 5840
rect 570 5830 757 5834
rect 761 5830 762 5834
rect 766 5830 767 5834
rect 771 5830 772 5834
rect 776 5830 783 5834
rect 787 5830 788 5834
rect 792 5830 793 5834
rect 797 5830 798 5834
rect 802 5830 809 5834
rect 813 5830 814 5834
rect 818 5830 819 5834
rect 823 5830 824 5834
rect 828 5830 835 5834
rect 839 5830 840 5834
rect 844 5830 845 5834
rect 849 5830 850 5834
rect 854 5830 861 5834
rect 865 5830 866 5834
rect 870 5830 871 5834
rect 875 5830 876 5834
rect 880 5830 1054 5834
rect 1058 5830 1059 5834
rect 1063 5830 1064 5834
rect 1068 5830 1069 5834
rect 1073 5830 1363 5834
rect 1367 5830 1368 5834
rect 1372 5830 1373 5834
rect 1377 5830 1378 5834
rect 1382 5830 1672 5834
rect 1676 5830 1677 5834
rect 1681 5830 1682 5834
rect 1686 5830 1687 5834
rect 1691 5830 1981 5834
rect 1985 5830 1986 5834
rect 1990 5830 1991 5834
rect 1995 5830 1996 5834
rect 2000 5830 2290 5834
rect 2294 5830 2295 5834
rect 2299 5830 2300 5834
rect 2304 5830 2305 5834
rect 2309 5830 2599 5834
rect 2603 5830 2604 5834
rect 2608 5830 2609 5834
rect 2613 5830 2614 5834
rect 2618 5830 2908 5834
rect 2912 5830 2913 5834
rect 2917 5830 2918 5834
rect 2922 5830 2923 5834
rect 2927 5830 3217 5834
rect 3221 5830 3222 5834
rect 3226 5830 3227 5834
rect 3231 5830 3232 5834
rect 3236 5830 3526 5834
rect 3530 5830 3531 5834
rect 3535 5830 3536 5834
rect 3540 5830 3541 5834
rect 3545 5830 3835 5834
rect 3839 5830 3840 5834
rect 3844 5830 3845 5834
rect 3849 5830 3850 5834
rect 3854 5830 4235 5834
rect 4239 5830 4240 5834
rect 4244 5830 4245 5834
rect 4249 5830 4250 5834
rect 4254 5830 4264 5834
rect 4268 5830 4269 5834
rect 4273 5830 4274 5834
rect 4278 5830 4279 5834
rect 4283 5830 4293 5834
rect 4297 5830 4298 5834
rect 4302 5830 4303 5834
rect 4307 5830 4308 5834
rect 4312 5830 4322 5834
rect 4326 5830 4327 5834
rect 4331 5830 4332 5834
rect 4336 5830 4337 5834
rect 4341 5830 4351 5834
rect 4355 5830 4356 5834
rect 4360 5830 4361 5834
rect 4365 5830 4366 5834
rect 4370 5830 4602 5834
rect 570 5824 4602 5830
rect 570 5820 757 5824
rect 761 5820 762 5824
rect 766 5820 767 5824
rect 771 5820 772 5824
rect 776 5820 783 5824
rect 787 5820 788 5824
rect 792 5820 793 5824
rect 797 5820 798 5824
rect 802 5820 809 5824
rect 813 5820 814 5824
rect 818 5820 819 5824
rect 823 5820 824 5824
rect 828 5820 835 5824
rect 839 5820 840 5824
rect 844 5820 845 5824
rect 849 5820 850 5824
rect 854 5820 861 5824
rect 865 5820 866 5824
rect 870 5820 871 5824
rect 875 5820 876 5824
rect 880 5820 1054 5824
rect 1058 5820 1059 5824
rect 1063 5820 1064 5824
rect 1068 5820 1069 5824
rect 1073 5820 1363 5824
rect 1367 5820 1368 5824
rect 1372 5820 1373 5824
rect 1377 5820 1378 5824
rect 1382 5820 1672 5824
rect 1676 5820 1677 5824
rect 1681 5820 1682 5824
rect 1686 5820 1687 5824
rect 1691 5820 1981 5824
rect 1985 5820 1986 5824
rect 1990 5820 1991 5824
rect 1995 5820 1996 5824
rect 2000 5820 2290 5824
rect 2294 5820 2295 5824
rect 2299 5820 2300 5824
rect 2304 5820 2305 5824
rect 2309 5820 2599 5824
rect 2603 5820 2604 5824
rect 2608 5820 2609 5824
rect 2613 5820 2614 5824
rect 2618 5820 2908 5824
rect 2912 5820 2913 5824
rect 2917 5820 2918 5824
rect 2922 5820 2923 5824
rect 2927 5820 3217 5824
rect 3221 5820 3222 5824
rect 3226 5820 3227 5824
rect 3231 5820 3232 5824
rect 3236 5820 3526 5824
rect 3530 5820 3531 5824
rect 3535 5820 3536 5824
rect 3540 5820 3541 5824
rect 3545 5820 3835 5824
rect 3839 5820 3840 5824
rect 3844 5820 3845 5824
rect 3849 5820 3850 5824
rect 3854 5820 4235 5824
rect 4239 5820 4240 5824
rect 4244 5820 4245 5824
rect 4249 5820 4250 5824
rect 4254 5820 4264 5824
rect 4268 5820 4269 5824
rect 4273 5820 4274 5824
rect 4278 5820 4279 5824
rect 4283 5820 4293 5824
rect 4297 5820 4298 5824
rect 4302 5820 4303 5824
rect 4307 5820 4308 5824
rect 4312 5820 4322 5824
rect 4326 5820 4327 5824
rect 4331 5820 4332 5824
rect 4336 5820 4337 5824
rect 4341 5820 4351 5824
rect 4355 5820 4356 5824
rect 4360 5820 4361 5824
rect 4365 5820 4366 5824
rect 4370 5820 4602 5824
rect 570 5777 4602 5820
<< pad >>
rect 1063 10036 1317 10290
rect 1372 10036 1626 10290
rect 1681 10036 1935 10290
rect 1990 10036 2244 10290
rect 2299 10036 2553 10290
rect 2608 10036 2862 10290
rect 2917 10036 3171 10290
rect 3226 10036 3480 10290
rect 3535 10036 3789 10290
rect 3844 10036 4098 10290
rect 89 9050 343 9304
rect 89 8741 343 8995
rect 89 8432 343 8686
rect 89 8123 343 8377
rect 89 7814 343 8068
rect 89 7505 343 7759
rect 89 7196 343 7450
rect 89 6887 343 7141
rect 89 6578 343 6832
rect 89 6269 343 6523
rect 4829 9062 5083 9316
rect 4829 8753 5083 9007
rect 4829 8444 5083 8698
rect 4829 8135 5083 8389
rect 4829 7827 5083 8081
rect 4829 7518 5083 7772
rect 4829 7208 5083 7462
rect 4829 6899 5083 7153
rect 4829 6590 5083 6844
rect 4829 6281 5083 6535
rect 1075 5296 1329 5550
rect 1384 5296 1638 5550
rect 1693 5296 1947 5550
rect 2002 5296 2256 5550
rect 2311 5296 2565 5550
rect 2620 5296 2874 5550
rect 2929 5296 3183 5550
rect 3238 5296 3492 5550
rect 3547 5296 3801 5550
rect 3856 5296 4110 5550
<< labels >>
rlabel metal3 4125 5872 4125 5872 5 GND!
rlabel metal3 4124 5846 4124 5846 5 Vdd!
rlabel metal1 3982 5720 3982 5720 5 Raw
rlabel metal3 4507 6242 4507 6242 3 GND!
rlabel metal3 4533 6241 4533 6241 3 Vdd!
rlabel metal3 4433 5872 4433 5872 5 GND!
rlabel metal3 4432 5846 4432 5846 5 Vdd!
rlabel metal3 3816 5872 3816 5872 5 GND!
rlabel metal3 3815 5846 3815 5846 5 Vdd!
rlabel metal1 3673 5720 3673 5720 5 Raw
rlabel metal3 3507 5872 3507 5872 5 GND!
rlabel metal3 3506 5846 3506 5846 5 Vdd!
rlabel metal1 3364 5720 3364 5720 5 Raw
rlabel metal3 3198 5872 3198 5872 5 GND!
rlabel metal3 3197 5846 3197 5846 5 Vdd!
rlabel metal1 3055 5720 3055 5720 5 Raw
rlabel metal3 2889 5872 2889 5872 5 GND!
rlabel metal3 2888 5846 2888 5846 5 Vdd!
rlabel metal1 2746 5720 2746 5720 5 Raw
rlabel metal3 2580 5872 2580 5872 5 GND!
rlabel metal3 2579 5846 2579 5846 5 Vdd!
rlabel metal1 2437 5720 2437 5720 5 Raw
rlabel metal3 2271 5872 2271 5872 5 GND!
rlabel metal3 2270 5846 2270 5846 5 Vdd!
rlabel metal1 2128 5720 2128 5720 5 Raw
rlabel metal3 1962 5872 1962 5872 5 GND!
rlabel metal3 1961 5846 1961 5846 5 Vdd!
rlabel metal1 1819 5720 1819 5720 5 Raw
rlabel metal3 1653 5872 1653 5872 5 GND!
rlabel metal3 1652 5846 1652 5846 5 Vdd!
rlabel metal1 1510 5720 1510 5720 5 Raw
rlabel metal3 1344 5872 1344 5872 5 GND!
rlabel metal3 1343 5846 1343 5846 5 Vdd!
rlabel metal1 1201 5720 1201 5720 5 Raw
rlabel metal3 1035 5872 1035 5872 5 GND!
rlabel metal3 1034 5846 1034 5846 5 Vdd!
rlabel metal3 665 5946 665 5946 7 GND!
rlabel metal3 639 5947 639 5947 7 Vdd!
rlabel metal3 665 6254 665 6254 7 GND!
rlabel metal3 639 6255 639 6255 7 Vdd!
rlabel metal1 513 6397 513 6397 7 Raw
rlabel metal3 4507 6550 4507 6550 3 GND!
rlabel metal3 4533 6549 4533 6549 3 Vdd!
rlabel metal1 4659 6407 4659 6407 3 Raw
rlabel metal3 4507 6859 4507 6859 3 GND!
rlabel metal3 4533 6858 4533 6858 3 Vdd!
rlabel metal1 4659 6716 4659 6716 3 Raw
rlabel metal3 4507 7168 4507 7168 3 GND!
rlabel metal3 4533 7167 4533 7167 3 Vdd!
rlabel metal1 4659 7025 4659 7025 3 Raw
rlabel metal3 4507 7477 4507 7477 3 GND!
rlabel metal3 4533 7476 4533 7476 3 Vdd!
rlabel metal1 4659 7334 4659 7334 3 Raw
rlabel metal3 4507 7503 4507 7503 3 GND!
rlabel metal3 4533 7504 4533 7504 3 Vdd!
rlabel metal1 4659 7646 4659 7646 3 Raw
rlabel metal3 4507 7812 4507 7812 3 GND!
rlabel metal3 4533 7813 4533 7813 3 Vdd!
rlabel metal1 4781 7954 4781 7954 3 RawOut
rlabel polycontact 4595 7962 4595 7962 3 _out
rlabel metal1 4441 7956 4441 7956 3 out
rlabel metal3 4532 7814 4532 7814 3 Vdd!
rlabel metal3 4507 8404 4507 8404 3 GND!
rlabel metal3 4533 8403 4533 8403 3 Vdd!
rlabel metal1 4659 8261 4659 8261 3 Raw
rlabel metal3 4507 8713 4507 8713 3 GND!
rlabel metal3 4533 8712 4533 8712 3 Vdd!
rlabel metal1 4659 8570 4659 8570 3 Raw
rlabel metal3 4507 9022 4507 9022 3 GND!
rlabel metal3 4533 9021 4533 9021 3 Vdd!
rlabel metal1 4659 8879 4659 8879 3 Raw
rlabel metal3 4507 9331 4507 9331 3 GND!
rlabel metal3 4533 9330 4533 9330 3 Vdd!
rlabel metal1 4659 9188 4659 9188 3 Raw
rlabel metal3 665 6563 665 6563 7 GND!
rlabel metal3 639 6564 639 6564 7 Vdd!
rlabel metal1 513 6706 513 6706 7 Raw
rlabel metal3 665 6872 665 6872 7 GND!
rlabel metal3 639 6873 639 6873 7 Vdd!
rlabel metal1 513 7015 513 7015 7 Raw
rlabel metal3 665 7181 665 7181 7 GND!
rlabel metal3 639 7182 639 7182 7 Vdd!
rlabel metal1 513 7324 513 7324 7 Raw
rlabel metal3 665 7490 665 7490 7 GND!
rlabel metal3 639 7491 639 7491 7 Vdd!
rlabel metal1 513 7633 513 7633 7 Raw
rlabel metal3 665 7799 665 7799 7 GND!
rlabel metal3 639 7800 639 7800 7 Vdd!
rlabel metal1 513 7942 513 7942 7 Raw
rlabel metal3 665 8108 665 8108 7 GND!
rlabel metal3 639 8109 639 8109 7 Vdd!
rlabel metal1 513 8251 513 8251 7 Raw
rlabel metal3 665 8417 665 8417 7 GND!
rlabel metal3 639 8418 639 8418 7 Vdd!
rlabel metal1 513 8560 513 8560 7 Raw
rlabel metal3 665 8726 665 8726 7 GND!
rlabel metal3 639 8727 639 8727 7 Vdd!
rlabel metal1 513 8869 513 8869 7 Raw
rlabel metal3 665 9035 665 9035 7 GND!
rlabel metal3 639 9036 639 9036 7 Vdd!
rlabel metal1 513 9178 513 9178 7 Raw
rlabel metal3 665 9344 665 9344 7 GND!
rlabel metal3 639 9345 639 9345 7 Vdd!
rlabel metal3 739 9714 739 9714 1 GND!
rlabel metal3 740 9740 740 9740 1 Vdd!
rlabel metal3 4137 9714 4137 9714 1 GND!
rlabel metal3 4138 9740 4138 9740 1 Vdd!
rlabel metal3 4507 9640 4507 9640 3 GND!
rlabel metal3 4533 9639 4533 9639 3 Vdd!
rlabel metal3 3829 9714 3829 9714 1 GND!
rlabel metal3 3830 9740 3830 9740 1 Vdd!
rlabel metal1 3964 9821 3964 9821 1 _RawIn
rlabel metal1 3970 9776 3970 9776 1 in
rlabel metal1 3971 9854 3971 9854 1 RawIn
rlabel metal3 3831 9739 3831 9739 1 Vdd!
rlabel metal3 3520 9714 3520 9714 1 GND!
rlabel metal3 3521 9740 3521 9740 1 Vdd!
rlabel m3contact 3524 9743 3524 9743 1 Vdd!0
rlabel metal3 3522 9739 3522 9739 1 Vdd!_uq0
rlabel metal1 3660 9855 3660 9855 1 Vdd!
rlabel metal3 3211 9714 3211 9714 1 GND!
rlabel metal3 3212 9740 3212 9740 1 Vdd!
rlabel metal1 3351 9855 3351 9855 1 GND!
rlabel metal3 3213 9739 3213 9739 1 Vdd!
rlabel metal3 2902 9714 2902 9714 1 GND!
rlabel metal3 2903 9740 2903 9740 1 Vdd!
rlabel metal1 3037 9821 3037 9821 1 _RawIn
rlabel metal1 3043 9776 3043 9776 1 in
rlabel metal1 3044 9854 3044 9854 1 RawIn
rlabel metal3 2904 9739 2904 9739 1 Vdd!
rlabel metal3 2593 9714 2593 9714 1 GND!
rlabel metal3 2594 9740 2594 9740 1 Vdd!
rlabel metal1 2728 9821 2728 9821 1 _RawIn
rlabel metal1 2734 9776 2734 9776 1 in
rlabel metal1 2735 9854 2735 9854 1 RawIn
rlabel metal3 2595 9739 2595 9739 1 Vdd!
rlabel metal3 2284 9714 2284 9714 1 GND!
rlabel metal3 2285 9740 2285 9740 1 Vdd!
rlabel metal1 2419 9821 2419 9821 1 _RawIn
rlabel metal1 2425 9776 2425 9776 1 in
rlabel metal1 2426 9854 2426 9854 1 RawIn
rlabel metal3 2286 9739 2286 9739 1 Vdd!
rlabel metal3 1975 9714 1975 9714 1 GND!
rlabel metal3 1976 9740 1976 9740 1 Vdd!
rlabel metal1 2110 9821 2110 9821 1 _RawIn
rlabel metal1 2116 9776 2116 9776 1 in
rlabel metal1 2117 9854 2117 9854 1 RawIn
rlabel metal3 1977 9739 1977 9739 1 Vdd!
rlabel metal3 1666 9714 1666 9714 1 GND!
rlabel metal3 1667 9740 1667 9740 1 Vdd!
rlabel metal1 1801 9821 1801 9821 1 _RawIn
rlabel metal1 1807 9776 1807 9776 1 in
rlabel metal1 1808 9854 1808 9854 1 RawIn
rlabel metal3 1668 9739 1668 9739 1 Vdd!
rlabel metal3 1357 9714 1357 9714 1 GND!
rlabel metal3 1358 9740 1358 9740 1 Vdd!
rlabel metal1 1497 9855 1497 9855 1 GND!
rlabel metal3 1359 9739 1359 9739 1 Vdd!
rlabel metal3 1048 9714 1048 9714 1 GND!
rlabel metal3 1049 9740 1049 9740 1 Vdd!
rlabel metal1 1191 9866 1191 9866 1 Raw
rlabel space 1998 10058 2232 10296 1 PROGRAM
rlabel pad 2309 10051 2543 10289 1 DATA
rlabel pad 2620 10045 2854 10283 1 clk
rlabel pad 3848 10042 4082 10280 1 RESET_b
rlabel space 2913 10037 3173 10297 1 MODE
rlabel space 3224 10034 3484 10294 1 GND!
rlabel space 3531 10034 3791 10294 1 Vdd!
rlabel space 4826 7826 5086 8086 1 OUT
rlabel metal2 3781 9351 3787 9355 1 reset_b
rlabel polysilicon 4247 7595 4247 7595 1 CB4
rlabel metal1 4095 7632 4098 7636 4 clk
rlabel metal1 4097 7561 4100 7565 2 ~clk
rlabel metal1 4096 7568 4099 7572 1 GND!
rlabel metal1 4095 7625 4098 7629 1 Vdd!
rlabel metal1 4095 7711 4098 7715 1 Vdd!
rlabel metal1 4096 7654 4099 7658 1 GND!
rlabel metal1 4097 7647 4100 7651 2 ~clk
rlabel metal1 4095 7718 4098 7722 4 clk
rlabel metal1 4095 8700 4098 8704 4 clk
rlabel metal1 4097 8629 4100 8633 2 ~clk
rlabel metal1 4096 8636 4099 8640 1 GND!
rlabel metal1 4095 8693 4098 8697 1 Vdd!
rlabel metal1 4095 8607 4098 8611 1 Vdd!
rlabel metal1 4096 8550 4099 8554 1 GND!
rlabel metal1 4097 8543 4100 8547 2 ~clk
rlabel metal1 4095 8614 4098 8618 4 clk
rlabel polysilicon 4235 7741 4235 7741 1 CB3
rlabel metal1 3928 8358 3931 8362 1 Vdd!
rlabel metal1 4050 7760 4053 7764 1 clk
rlabel metal1 4047 7812 4051 7816 1 ~clk
rlabel metal1 4046 7819 4050 7823 1 GND!
rlabel metal1 4057 7753 4061 7757 1 Vdd!
rlabel metal2 4113 8285 4116 8291 1 select2
rlabel metal2 4053 8285 4056 8292 1 select1
rlabel metal2 3970 8286 3973 8291 1 select0
rlabel m3contact 3793 8331 3796 8334 3 ctrl_reg
rlabel metal1 4192 8358 4195 8362 1 Vdd!
rlabel metal1 4193 8301 4196 8305 1 GND!
rlabel metal1 4194 8294 4197 8298 2 ~clk
rlabel metal1 4192 8365 4195 8369 4 clk
rlabel metal1 4060 8365 4063 8369 4 clk
rlabel metal1 4062 8294 4065 8298 2 ~clk
rlabel metal1 4061 8301 4064 8305 1 GND!
rlabel metal1 4060 8358 4063 8362 1 Vdd!
rlabel metal1 3928 8365 3931 8369 4 clk
rlabel metal1 3930 8294 3933 8298 2 ~clk
rlabel metal1 3929 8301 3932 8305 1 GND!
rlabel metal1 3796 8365 3799 8369 4 clk
rlabel metal1 3798 8294 3801 8298 2 ~clk
rlabel metal1 3797 8301 3800 8305 1 GND!
rlabel metal1 3796 8358 3799 8362 1 Vdd!
rlabel metal2 4141 8276 4144 8281 1 select_out
rlabel metal1 4078 8215 4081 8219 1 GND!
rlabel metal1 3997 8215 4000 8219 1 GND!
rlabel metal1 4077 8281 4081 8285 1 Vdd!
rlabel metal1 3996 8281 4000 8285 1 Vdd!
rlabel metal1 4146 8120 4149 8123 7 Y
rlabel metal1 4077 8149 4081 8153 1 Vdd!
rlabel metal1 3996 8149 4000 8153 1 Vdd!
rlabel metal1 4102 8083 4105 8087 1 GND!
rlabel metal1 3997 8083 4000 8087 1 GND!
rlabel metal1 4077 8017 4081 8021 1 Vdd!
rlabel metal1 3996 8017 4000 8021 1 Vdd!
rlabel metal1 4167 8017 4171 8021 1 Vdd!
rlabel metal1 3997 7951 4000 7955 1 GND!
rlabel metal1 4078 7951 4081 7955 1 GND!
rlabel metal1 4168 7951 4171 7955 1 GND!
rlabel metal1 3996 7885 4000 7889 1 Vdd!
rlabel metal1 4077 7885 4081 7889 1 Vdd!
rlabel metal1 4167 7885 4171 7889 1 Vdd!
rlabel metal1 3997 7819 4000 7823 1 GND!
rlabel metal1 3996 7753 4000 7757 1 Vdd!
rlabel polysilicon 4040 7783 4042 7786 5 D
rlabel polysilicon 4058 7792 4060 7795 5 reset
rlabel metal1 3794 8010 3798 8014 3 clk
rlabel metal1 3794 8017 3798 8021 3 Vdd!
rlabel metal1 3794 7958 3798 7962 3 ~clk
rlabel metal1 3794 7892 3798 7896 3 clk
rlabel metal1 3794 7944 3798 7948 3 ~clk
rlabel metal1 3794 7951 3798 7955 3 GND!
rlabel metal1 3794 7878 3798 7882 3 clk
rlabel metal1 3794 7885 3798 7889 3 Vdd!
rlabel metal1 3794 7826 3798 7830 3 ~clk
rlabel metal1 3794 7753 3798 7757 3 Vdd!
rlabel metal1 3794 7812 3798 7816 3 ~clk
rlabel metal1 3794 7819 3798 7823 3 GND!
rlabel metal1 3794 8083 3798 8087 3 GND!
rlabel metal1 3794 8076 3798 8080 3 ~clk
rlabel metal1 3794 8024 3798 8028 3 clk
rlabel metal1 3794 8090 3798 8094 3 ~clk
rlabel metal1 3794 8149 3798 8153 3 Vdd!
rlabel metal1 3794 8142 3798 8146 3 clk
rlabel metal1 3794 8215 3798 8219 3 GND!
rlabel metal1 3794 8208 3798 8212 3 ~clk
rlabel metal1 3794 8222 3798 8226 3 ~clk
rlabel metal1 3794 8281 3798 8285 3 Vdd!
rlabel metal1 3794 8274 3798 8278 3 clk
rlabel metal1 3794 9256 3798 9260 3 clk
rlabel metal1 3794 9263 3798 9267 3 Vdd!
rlabel metal1 3794 9204 3798 9208 3 ~clk
rlabel metal1 3794 9190 3798 9194 3 ~clk
rlabel metal1 3794 9197 3798 9201 3 GND!
rlabel metal1 3794 9124 3798 9128 3 clk
rlabel metal1 3794 9131 3798 9135 3 Vdd!
rlabel metal1 3794 9072 3798 9076 3 ~clk
rlabel metal1 3794 9006 3798 9010 3 clk
rlabel metal1 3794 9058 3798 9062 3 ~clk
rlabel metal1 3794 9065 3798 9069 3 GND!
rlabel metal1 3794 8801 3798 8805 3 GND!
rlabel metal1 3794 8794 3798 8798 3 ~clk
rlabel metal1 3794 8735 3798 8739 3 Vdd!
rlabel metal1 3794 8808 3798 8812 3 ~clk
rlabel metal1 3794 8867 3798 8871 3 Vdd!
rlabel metal1 3794 8860 3798 8864 3 clk
rlabel metal1 3794 8933 3798 8937 3 GND!
rlabel metal1 3794 8926 3798 8930 3 ~clk
rlabel metal1 3794 8874 3798 8878 3 clk
rlabel metal1 3794 8940 3798 8944 3 ~clk
rlabel metal1 3794 8999 3798 9003 3 Vdd!
rlabel metal1 3794 8992 3798 8996 3 clk
rlabel polysilicon 4058 8774 4060 8777 5 reset
rlabel metal1 3996 8735 4000 8739 1 Vdd!
rlabel metal1 3997 8801 4000 8805 1 GND!
rlabel metal1 4167 8867 4171 8871 1 Vdd!
rlabel metal1 4077 8867 4081 8871 1 Vdd!
rlabel metal1 3996 8867 4000 8871 1 Vdd!
rlabel metal1 4168 8933 4171 8937 1 GND!
rlabel metal1 4078 8933 4081 8937 1 GND!
rlabel metal1 3997 8933 4000 8937 1 GND!
rlabel metal1 4167 8999 4171 9003 1 Vdd!
rlabel metal1 3996 8999 4000 9003 1 Vdd!
rlabel metal1 4077 8999 4081 9003 1 Vdd!
rlabel metal1 3997 9065 4000 9069 1 GND!
rlabel metal1 4102 9065 4105 9069 1 GND!
rlabel metal1 3996 9131 4000 9135 1 Vdd!
rlabel metal1 4077 9131 4081 9135 1 Vdd!
rlabel metal1 4146 9102 4149 9105 7 Y
rlabel metal1 3996 9263 4000 9267 1 Vdd!
rlabel metal1 4077 9263 4081 9267 1 Vdd!
rlabel metal1 3997 9197 4000 9201 1 GND!
rlabel metal1 4078 9197 4081 9201 1 GND!
rlabel metal2 4141 9258 4144 9263 1 select_out
rlabel metal1 3796 9340 3799 9344 1 Vdd!
rlabel metal1 3797 9283 3800 9287 1 GND!
rlabel metal1 3798 9276 3801 9280 2 ~clk
rlabel metal1 3796 9347 3799 9351 4 clk
rlabel metal1 3929 9283 3932 9287 1 GND!
rlabel metal1 3930 9276 3933 9280 2 ~clk
rlabel metal1 3928 9347 3931 9351 4 clk
rlabel metal1 4060 9340 4063 9344 1 Vdd!
rlabel metal1 4061 9283 4064 9287 1 GND!
rlabel metal1 4062 9276 4065 9280 2 ~clk
rlabel metal1 4060 9347 4063 9351 4 clk
rlabel metal1 4192 9347 4195 9351 4 clk
rlabel metal1 4194 9276 4197 9280 2 ~clk
rlabel metal1 4193 9283 4196 9287 1 GND!
rlabel metal1 4192 9340 4195 9344 1 Vdd!
rlabel m3contact 3793 9313 3796 9316 3 ctrl_reg
rlabel metal2 3970 9268 3973 9273 1 select0
rlabel metal2 4053 9267 4056 9274 1 select1
rlabel metal2 4113 9267 4116 9273 1 select2
rlabel metal1 4057 8735 4061 8739 1 Vdd!
rlabel metal1 4046 8801 4050 8805 1 GND!
rlabel metal1 4047 8794 4051 8798 1 ~clk
rlabel metal1 4050 8742 4053 8746 1 clk
rlabel metal1 3928 9340 3931 9344 1 Vdd!
rlabel metal1 4226 8972 4226 8972 1 out
rlabel metal2 3772 8373 3772 8373 5 p_clk
rlabel metal2 3772 9355 3772 9355 5 p_clk
rlabel metal1 3163 7711 3166 7715 1 Vdd!
rlabel metal1 3312 7455 3315 7459 1 Vdd!
rlabel metal1 3313 7398 3316 7402 1 GND!
rlabel metal1 3314 7391 3317 7395 2 ~clk
rlabel metal1 3312 7462 3315 7466 4 clk
rlabel metal1 3444 7455 3447 7459 1 Vdd!
rlabel metal1 3445 7398 3448 7402 1 GND!
rlabel metal1 3446 7391 3449 7395 2 ~clk
rlabel metal1 3444 7462 3447 7466 4 clk
rlabel metal1 3576 7455 3579 7459 1 Vdd!
rlabel metal1 3577 7398 3580 7402 1 GND!
rlabel metal1 3578 7391 3581 7395 2 ~clk
rlabel metal1 3576 7462 3579 7466 4 clk
rlabel metal1 3312 7595 3315 7599 1 Vdd!
rlabel metal1 3313 7538 3316 7542 1 GND!
rlabel metal1 3314 7531 3317 7535 2 ~clk
rlabel metal1 3312 7602 3315 7606 4 clk
rlabel metal1 3444 7595 3447 7599 1 Vdd!
rlabel metal1 3445 7538 3448 7542 1 GND!
rlabel metal1 3446 7531 3449 7535 2 ~clk
rlabel metal1 3444 7602 3447 7606 4 clk
rlabel metal1 3576 7595 3579 7599 1 Vdd!
rlabel metal1 3577 7538 3580 7542 1 GND!
rlabel metal1 3578 7531 3581 7535 2 ~clk
rlabel metal1 3576 7602 3579 7606 4 clk
rlabel metal1 3576 7688 3579 7692 4 clk
rlabel metal1 3578 7617 3581 7621 2 ~clk
rlabel metal1 3577 7624 3580 7628 1 GND!
rlabel metal1 3576 7681 3579 7685 1 Vdd!
rlabel metal1 3444 7688 3447 7692 4 clk
rlabel metal1 3446 7617 3449 7621 2 ~clk
rlabel metal1 3445 7624 3448 7628 1 GND!
rlabel metal1 3444 7681 3447 7685 1 Vdd!
rlabel metal1 3312 7688 3315 7692 4 clk
rlabel metal1 3314 7617 3317 7621 2 ~clk
rlabel metal1 3313 7624 3316 7628 1 GND!
rlabel metal1 3312 7681 3315 7685 1 Vdd!
rlabel metal1 3150 7632 3153 7636 4 clk
rlabel metal1 3152 7561 3155 7565 2 ~clk
rlabel metal1 3151 7568 3154 7572 1 GND!
rlabel metal1 3150 7625 3153 7629 1 Vdd!
rlabel metal1 3151 7654 3154 7658 1 GND!
rlabel metal1 3152 7647 3155 7651 2 ~clk
rlabel metal1 3150 7718 3153 7722 4 clk
rlabel metal1 2367 7455 2370 7459 1 Vdd!
rlabel metal1 2368 7398 2371 7402 1 GND!
rlabel metal1 2369 7391 2372 7395 2 ~clk
rlabel metal1 2367 7462 2370 7466 4 clk
rlabel metal1 2499 7455 2502 7459 1 Vdd!
rlabel metal1 2500 7398 2503 7402 1 GND!
rlabel metal1 2501 7391 2504 7395 2 ~clk
rlabel metal1 2499 7462 2502 7466 4 clk
rlabel metal1 2631 7455 2634 7459 1 Vdd!
rlabel metal1 2632 7398 2635 7402 1 GND!
rlabel metal1 2633 7391 2636 7395 2 ~clk
rlabel metal1 2631 7462 2634 7466 4 clk
rlabel metal1 2367 7595 2370 7599 1 Vdd!
rlabel metal1 2368 7538 2371 7542 1 GND!
rlabel metal1 2369 7531 2372 7535 2 ~clk
rlabel metal1 2367 7602 2370 7606 4 clk
rlabel metal1 2499 7595 2502 7599 1 Vdd!
rlabel metal1 2500 7538 2503 7542 1 GND!
rlabel metal1 2501 7531 2504 7535 2 ~clk
rlabel metal1 2499 7602 2502 7606 4 clk
rlabel metal1 2631 7595 2634 7599 1 Vdd!
rlabel metal1 2632 7538 2635 7542 1 GND!
rlabel metal1 2633 7531 2636 7535 2 ~clk
rlabel metal1 2631 7602 2634 7606 4 clk
rlabel metal1 2631 7688 2634 7692 4 clk
rlabel metal1 2633 7617 2636 7621 2 ~clk
rlabel metal1 2632 7624 2635 7628 1 GND!
rlabel metal1 2631 7681 2634 7685 1 Vdd!
rlabel metal1 2499 7688 2502 7692 4 clk
rlabel metal1 2501 7617 2504 7621 2 ~clk
rlabel metal1 2500 7624 2503 7628 1 GND!
rlabel metal1 2499 7681 2502 7685 1 Vdd!
rlabel metal1 2367 7688 2370 7692 4 clk
rlabel metal1 2369 7617 2372 7621 2 ~clk
rlabel metal1 2368 7624 2371 7628 1 GND!
rlabel metal1 2367 7681 2370 7685 1 Vdd!
rlabel metal1 3150 8700 3153 8704 4 clk
rlabel metal1 3152 8629 3155 8633 2 ~clk
rlabel metal1 3151 8636 3154 8640 1 GND!
rlabel metal1 3150 8693 3153 8697 1 Vdd!
rlabel metal1 3150 8607 3153 8611 1 Vdd!
rlabel metal1 3151 8550 3154 8554 1 GND!
rlabel metal1 3152 8543 3155 8547 2 ~clk
rlabel metal1 3150 8614 3153 8618 4 clk
rlabel polysilicon 3302 8577 3302 8577 1 CB4
rlabel metal1 3312 8663 3315 8667 1 Vdd!
rlabel metal1 3313 8606 3316 8610 1 GND!
rlabel metal1 3314 8599 3317 8603 2 ~clk
rlabel metal1 3312 8670 3315 8674 4 clk
rlabel metal1 3444 8663 3447 8667 1 Vdd!
rlabel metal1 3445 8606 3448 8610 1 GND!
rlabel metal1 3446 8599 3449 8603 2 ~clk
rlabel metal1 3444 8670 3447 8674 4 clk
rlabel metal1 3576 8663 3579 8667 1 Vdd!
rlabel metal1 3577 8606 3580 8610 1 GND!
rlabel metal1 3578 8599 3581 8603 2 ~clk
rlabel metal1 3576 8670 3579 8674 4 clk
rlabel metal1 3576 8584 3579 8588 4 clk
rlabel metal1 3578 8513 3581 8517 2 ~clk
rlabel metal1 3577 8520 3580 8524 1 GND!
rlabel metal1 3576 8577 3579 8581 1 Vdd!
rlabel metal1 3444 8584 3447 8588 4 clk
rlabel metal1 3446 8513 3449 8517 2 ~clk
rlabel metal1 3445 8520 3448 8524 1 GND!
rlabel metal1 3444 8577 3447 8581 1 Vdd!
rlabel metal1 3312 8584 3315 8588 4 clk
rlabel metal1 3314 8513 3317 8517 2 ~clk
rlabel metal1 3313 8520 3316 8524 1 GND!
rlabel metal1 3312 8577 3315 8581 1 Vdd!
rlabel metal1 3576 8444 3579 8448 4 clk
rlabel metal1 3578 8373 3581 8377 2 ~clk
rlabel metal1 3577 8380 3580 8384 1 GND!
rlabel metal1 3576 8437 3579 8441 1 Vdd!
rlabel metal1 3444 8444 3447 8448 4 clk
rlabel metal1 3446 8373 3449 8377 2 ~clk
rlabel metal1 3445 8380 3448 8384 1 GND!
rlabel metal1 3444 8437 3447 8441 1 Vdd!
rlabel metal1 3312 8444 3315 8448 4 clk
rlabel metal1 3314 8373 3317 8377 2 ~clk
rlabel metal1 3313 8380 3316 8384 1 GND!
rlabel metal1 3312 8437 3315 8441 1 Vdd!
rlabel metal2 3723 8374 3723 8374 1 GND!
rlabel metal2 3711 8374 3711 8374 1 Vdd!
rlabel polysilicon 3457 8244 3457 8244 1 CB1
rlabel metal1 3560 8230 3563 8234 6 clk
rlabel metal1 3558 8159 3561 8163 8 ~clk
rlabel metal1 3559 8166 3562 8170 1 GND!
rlabel metal1 3560 8223 3563 8227 1 Vdd!
rlabel polysilicon 3574 8252 3574 8252 1 CB2
rlabel metal1 3444 8332 3447 8336 4 clk
rlabel metal1 3446 8261 3449 8265 2 ~clk
rlabel metal1 3445 8268 3448 8272 1 GND!
rlabel metal1 3444 8325 3447 8329 1 Vdd!
rlabel metal2 3736 8373 3736 8373 4 f_clk_b
rlabel metal2 3748 8372 3748 8372 5 f_clk
rlabel metal2 3760 8373 3760 8373 5 p_clk_b
rlabel metal1 3576 7830 3579 7834 4 clk
rlabel metal1 3578 7759 3581 7763 2 ~clk
rlabel metal1 3577 7766 3580 7770 1 GND!
rlabel metal1 3576 7823 3579 7827 1 Vdd!
rlabel metal1 3444 7830 3447 7834 4 clk
rlabel metal1 3446 7759 3449 7763 2 ~clk
rlabel metal1 3445 7766 3448 7770 1 GND!
rlabel metal1 3444 7823 3447 7827 1 Vdd!
rlabel metal1 3312 7830 3315 7834 4 clk
rlabel metal1 3314 7759 3317 7763 2 ~clk
rlabel metal1 3313 7766 3316 7770 1 GND!
rlabel metal1 3312 7823 3315 7827 1 Vdd!
rlabel metal1 2983 8358 2986 8362 1 Vdd!
rlabel metal1 3105 7760 3108 7764 1 clk
rlabel metal1 3102 7812 3106 7816 1 ~clk
rlabel metal1 3101 7819 3105 7823 1 GND!
rlabel metal1 3112 7753 3116 7757 1 Vdd!
rlabel metal2 3168 8285 3171 8291 1 select2
rlabel metal2 3108 8285 3111 8292 1 select1
rlabel metal2 3025 8286 3028 8291 1 select0
rlabel metal1 3247 8358 3250 8362 1 Vdd!
rlabel metal1 3248 8301 3251 8305 1 GND!
rlabel metal1 3249 8294 3252 8298 2 ~clk
rlabel metal1 3247 8365 3250 8369 4 clk
rlabel metal1 3115 8365 3118 8369 4 clk
rlabel metal1 3117 8294 3120 8298 2 ~clk
rlabel metal1 3116 8301 3119 8305 1 GND!
rlabel metal1 3115 8358 3118 8362 1 Vdd!
rlabel metal1 2983 8365 2986 8369 4 clk
rlabel metal1 2985 8294 2988 8298 2 ~clk
rlabel metal1 2984 8301 2987 8305 1 GND!
rlabel metal1 2851 8365 2854 8369 4 clk
rlabel metal1 2853 8294 2856 8298 2 ~clk
rlabel metal1 2852 8301 2855 8305 1 GND!
rlabel metal1 2851 8358 2854 8362 1 Vdd!
rlabel metal2 3196 8276 3199 8281 1 select_out
rlabel metal1 3133 8215 3136 8219 1 GND!
rlabel metal1 3052 8215 3055 8219 1 GND!
rlabel metal1 3132 8281 3136 8285 1 Vdd!
rlabel metal1 3051 8281 3055 8285 1 Vdd!
rlabel metal1 3201 8120 3204 8123 7 Y
rlabel metal1 3132 8149 3136 8153 1 Vdd!
rlabel metal1 3051 8149 3055 8153 1 Vdd!
rlabel metal1 3157 8083 3160 8087 1 GND!
rlabel metal1 3052 8083 3055 8087 1 GND!
rlabel metal1 3132 8017 3136 8021 1 Vdd!
rlabel metal1 3051 8017 3055 8021 1 Vdd!
rlabel metal1 3222 8017 3226 8021 1 Vdd!
rlabel metal1 3052 7951 3055 7955 1 GND!
rlabel metal1 3133 7951 3136 7955 1 GND!
rlabel metal1 3223 7951 3226 7955 1 GND!
rlabel metal1 3051 7885 3055 7889 1 Vdd!
rlabel metal1 3132 7885 3136 7889 1 Vdd!
rlabel metal1 3222 7885 3226 7889 1 Vdd!
rlabel metal1 3052 7819 3055 7823 1 GND!
rlabel metal1 3051 7753 3055 7757 1 Vdd!
rlabel polysilicon 3095 7783 3097 7786 5 D
rlabel polysilicon 3113 7792 3115 7795 5 reset
rlabel metal1 2849 8010 2853 8014 3 clk
rlabel metal1 2849 8017 2853 8021 3 Vdd!
rlabel metal1 2849 7958 2853 7962 3 ~clk
rlabel metal1 2849 7892 2853 7896 3 clk
rlabel metal1 2849 7944 2853 7948 3 ~clk
rlabel metal1 2849 7951 2853 7955 3 GND!
rlabel metal1 2849 7878 2853 7882 3 clk
rlabel metal1 2849 7885 2853 7889 3 Vdd!
rlabel metal1 2849 7826 2853 7830 3 ~clk
rlabel metal1 2849 7753 2853 7757 3 Vdd!
rlabel metal1 2849 7812 2853 7816 3 ~clk
rlabel metal1 2849 7819 2853 7823 3 GND!
rlabel metal1 2849 8083 2853 8087 3 GND!
rlabel metal1 2849 8076 2853 8080 3 ~clk
rlabel metal1 2849 8024 2853 8028 3 clk
rlabel metal1 2849 8090 2853 8094 3 ~clk
rlabel metal1 2849 8149 2853 8153 3 Vdd!
rlabel metal1 2849 8142 2853 8146 3 clk
rlabel metal1 2849 8215 2853 8219 3 GND!
rlabel metal1 2849 8208 2853 8212 3 ~clk
rlabel metal1 2849 8222 2853 8226 3 ~clk
rlabel metal1 2849 8281 2853 8285 3 Vdd!
rlabel metal1 2849 8274 2853 8278 3 clk
rlabel metal2 3184 8112 3184 8112 2 Core
rlabel metal1 2367 8663 2370 8667 1 Vdd!
rlabel metal1 2368 8606 2371 8610 1 GND!
rlabel metal1 2369 8599 2372 8603 2 ~clk
rlabel metal1 2367 8670 2370 8674 4 clk
rlabel metal1 2499 8663 2502 8667 1 Vdd!
rlabel metal1 2500 8606 2503 8610 1 GND!
rlabel metal1 2501 8599 2504 8603 2 ~clk
rlabel metal1 2499 8670 2502 8674 4 clk
rlabel metal1 2631 8663 2634 8667 1 Vdd!
rlabel metal1 2632 8606 2635 8610 1 GND!
rlabel metal1 2633 8599 2636 8603 2 ~clk
rlabel metal1 2631 8670 2634 8674 4 clk
rlabel metal1 2631 8584 2634 8588 4 clk
rlabel metal1 2633 8513 2636 8517 2 ~clk
rlabel metal1 2632 8520 2635 8524 1 GND!
rlabel metal1 2631 8577 2634 8581 1 Vdd!
rlabel metal1 2499 8584 2502 8588 4 clk
rlabel metal1 2501 8513 2504 8517 2 ~clk
rlabel metal1 2500 8520 2503 8524 1 GND!
rlabel metal1 2499 8577 2502 8581 1 Vdd!
rlabel metal1 2367 8584 2370 8588 4 clk
rlabel metal1 2369 8513 2372 8517 2 ~clk
rlabel metal1 2368 8520 2371 8524 1 GND!
rlabel metal1 2367 8577 2370 8581 1 Vdd!
rlabel metal1 2631 8444 2634 8448 4 clk
rlabel metal1 2633 8373 2636 8377 2 ~clk
rlabel metal1 2632 8380 2635 8384 1 GND!
rlabel metal1 2631 8437 2634 8441 1 Vdd!
rlabel metal1 2499 8444 2502 8448 4 clk
rlabel metal1 2501 8373 2504 8377 2 ~clk
rlabel metal1 2500 8380 2503 8384 1 GND!
rlabel metal1 2499 8437 2502 8441 1 Vdd!
rlabel metal1 2367 8444 2370 8448 4 clk
rlabel metal1 2369 8373 2372 8377 2 ~clk
rlabel metal1 2368 8380 2371 8384 1 GND!
rlabel metal1 2367 8437 2370 8441 1 Vdd!
rlabel metal2 2778 8374 2778 8374 1 GND!
rlabel metal2 2766 8374 2766 8374 1 Vdd!
rlabel metal1 2615 8230 2618 8234 6 clk
rlabel metal1 2613 8159 2616 8163 8 ~clk
rlabel metal1 2614 8166 2617 8170 1 GND!
rlabel metal1 2615 8223 2618 8227 1 Vdd!
rlabel polysilicon 2629 8252 2629 8252 1 CB2
rlabel metal1 2499 8332 2502 8336 4 clk
rlabel metal1 2501 8261 2504 8265 2 ~clk
rlabel metal1 2500 8268 2503 8272 1 GND!
rlabel metal1 2499 8325 2502 8329 1 Vdd!
rlabel metal2 2791 8373 2791 8373 4 f_clk_b
rlabel metal2 2803 8372 2803 8372 5 f_clk
rlabel metal2 2827 8373 2827 8373 5 p_clk
rlabel metal2 2815 8373 2815 8373 5 p_clk_b
rlabel metal1 2631 7830 2634 7834 4 clk
rlabel metal1 2633 7759 2636 7763 2 ~clk
rlabel metal1 2632 7766 2635 7770 1 GND!
rlabel metal1 2631 7823 2634 7827 1 Vdd!
rlabel metal1 2499 7830 2502 7834 4 clk
rlabel metal1 2501 7759 2504 7763 2 ~clk
rlabel metal1 2500 7766 2503 7770 1 GND!
rlabel metal1 2499 7823 2502 7827 1 Vdd!
rlabel metal1 2369 7759 2372 7763 2 ~clk
rlabel metal1 2368 7766 2371 7770 1 GND!
rlabel metal1 2849 9256 2853 9260 3 clk
rlabel metal1 2849 9263 2853 9267 3 Vdd!
rlabel metal1 2849 9204 2853 9208 3 ~clk
rlabel metal1 2849 9190 2853 9194 3 ~clk
rlabel metal1 2849 9197 2853 9201 3 GND!
rlabel metal1 2849 9124 2853 9128 3 clk
rlabel metal1 2849 9131 2853 9135 3 Vdd!
rlabel metal1 2849 9072 2853 9076 3 ~clk
rlabel metal1 2849 9006 2853 9010 3 clk
rlabel metal1 2849 9058 2853 9062 3 ~clk
rlabel metal1 2849 9065 2853 9069 3 GND!
rlabel metal1 2849 8801 2853 8805 3 GND!
rlabel metal1 2849 8794 2853 8798 3 ~clk
rlabel metal1 2849 8735 2853 8739 3 Vdd!
rlabel metal1 2849 8808 2853 8812 3 ~clk
rlabel metal1 2849 8867 2853 8871 3 Vdd!
rlabel metal1 2849 8860 2853 8864 3 clk
rlabel metal1 2849 8933 2853 8937 3 GND!
rlabel metal1 2849 8926 2853 8930 3 ~clk
rlabel metal1 2849 8874 2853 8878 3 clk
rlabel metal1 2849 8940 2853 8944 3 ~clk
rlabel metal1 2849 8999 2853 9003 3 Vdd!
rlabel metal1 2849 8992 2853 8996 3 clk
rlabel polysilicon 3113 8774 3115 8777 5 reset
rlabel polysilicon 3095 8765 3097 8768 5 D
rlabel metal1 3051 8735 3055 8739 1 Vdd!
rlabel metal1 3052 8801 3055 8805 1 GND!
rlabel metal1 3222 8867 3226 8871 1 Vdd!
rlabel metal1 3132 8867 3136 8871 1 Vdd!
rlabel metal1 3051 8867 3055 8871 1 Vdd!
rlabel metal1 3223 8933 3226 8937 1 GND!
rlabel metal1 3133 8933 3136 8937 1 GND!
rlabel metal1 3052 8933 3055 8937 1 GND!
rlabel metal1 3222 8999 3226 9003 1 Vdd!
rlabel metal1 3051 8999 3055 9003 1 Vdd!
rlabel metal1 3132 8999 3136 9003 1 Vdd!
rlabel metal1 3052 9065 3055 9069 1 GND!
rlabel metal1 3157 9065 3160 9069 1 GND!
rlabel metal1 3051 9131 3055 9135 1 Vdd!
rlabel metal1 3132 9131 3136 9135 1 Vdd!
rlabel metal1 3201 9102 3204 9105 7 Y
rlabel metal1 3051 9263 3055 9267 1 Vdd!
rlabel metal1 3132 9263 3136 9267 1 Vdd!
rlabel metal1 3052 9197 3055 9201 1 GND!
rlabel metal1 3133 9197 3136 9201 1 GND!
rlabel metal2 3196 9258 3199 9263 1 select_out
rlabel metal1 2851 9340 2854 9344 1 Vdd!
rlabel metal1 2852 9283 2855 9287 1 GND!
rlabel metal1 2853 9276 2856 9280 2 ~clk
rlabel metal1 2851 9347 2854 9351 4 clk
rlabel metal1 2984 9283 2987 9287 1 GND!
rlabel metal1 2985 9276 2988 9280 2 ~clk
rlabel metal1 2983 9347 2986 9351 4 clk
rlabel metal1 3115 9340 3118 9344 1 Vdd!
rlabel metal1 3116 9283 3119 9287 1 GND!
rlabel metal1 3117 9276 3120 9280 2 ~clk
rlabel metal1 3115 9347 3118 9351 4 clk
rlabel metal1 3247 9347 3250 9351 4 clk
rlabel metal1 3249 9276 3252 9280 2 ~clk
rlabel metal1 3248 9283 3251 9287 1 GND!
rlabel metal1 3247 9340 3250 9344 1 Vdd!
rlabel m3contact 2848 9313 2851 9316 3 ctrl_reg
rlabel metal2 3025 9268 3028 9273 1 select0
rlabel metal2 3108 9267 3111 9274 1 select1
rlabel metal2 3168 9267 3171 9273 1 select2
rlabel metal1 3112 8735 3116 8739 1 Vdd!
rlabel metal1 3101 8801 3105 8805 1 GND!
rlabel metal1 3102 8794 3106 8798 1 ~clk
rlabel metal1 3105 8742 3108 8746 1 clk
rlabel metal1 2983 9340 2986 9344 1 Vdd!
rlabel polysilicon 3290 8723 3290 8723 1 CB3
rlabel metal1 3312 8805 3315 8809 1 Vdd!
rlabel metal1 3313 8748 3316 8752 1 GND!
rlabel metal1 3314 8741 3317 8745 2 ~clk
rlabel metal1 3312 8812 3315 8816 4 clk
rlabel metal1 3444 8805 3447 8809 1 Vdd!
rlabel metal1 3445 8748 3448 8752 1 GND!
rlabel metal1 3446 8741 3449 8745 2 ~clk
rlabel metal1 3444 8812 3447 8816 4 clk
rlabel metal1 3576 8805 3579 8809 1 Vdd!
rlabel metal1 3577 8748 3580 8752 1 GND!
rlabel metal1 3578 8741 3581 8745 2 ~clk
rlabel metal1 3576 8812 3579 8816 4 clk
rlabel metal2 3760 9355 3760 9355 5 p_clk_b
rlabel metal2 3748 9354 3748 9354 5 f_clk
rlabel metal2 3736 9355 3736 9355 4 f_clk_b
rlabel metal1 3444 9307 3447 9311 1 Vdd!
rlabel metal1 3445 9250 3448 9254 1 GND!
rlabel metal1 3446 9243 3449 9247 2 ~clk
rlabel metal1 3444 9314 3447 9318 4 clk
rlabel polysilicon 3574 9234 3574 9234 1 CB2
rlabel metal1 3560 9205 3563 9209 1 Vdd!
rlabel metal1 3559 9148 3562 9152 1 GND!
rlabel metal1 3558 9141 3561 9145 8 ~clk
rlabel metal1 3560 9212 3563 9216 6 clk
rlabel metal1 3565 9180 3565 9180 1 D
rlabel polysilicon 3457 9226 3457 9226 1 CB1
rlabel metal2 3711 9356 3711 9356 1 Vdd!
rlabel metal2 3723 9356 3723 9356 1 GND!
rlabel metal1 2367 8805 2370 8809 1 Vdd!
rlabel metal1 2368 8748 2371 8752 1 GND!
rlabel metal1 2369 8741 2372 8745 2 ~clk
rlabel metal1 2367 8812 2370 8816 4 clk
rlabel metal1 2499 8805 2502 8809 1 Vdd!
rlabel metal1 2500 8748 2503 8752 1 GND!
rlabel metal1 2501 8741 2504 8745 2 ~clk
rlabel metal1 2499 8812 2502 8816 4 clk
rlabel metal1 2631 8805 2634 8809 1 Vdd!
rlabel metal1 2632 8748 2635 8752 1 GND!
rlabel metal1 2633 8741 2636 8745 2 ~clk
rlabel metal1 2631 8812 2634 8816 4 clk
rlabel metal2 2815 9355 2815 9355 5 p_clk_b
rlabel metal2 2827 9355 2827 9355 5 p_clk
rlabel metal2 2803 9354 2803 9354 5 f_clk
rlabel metal2 2791 9355 2791 9355 4 f_clk_b
rlabel metal1 2499 9307 2502 9311 1 Vdd!
rlabel metal1 2500 9250 2503 9254 1 GND!
rlabel metal1 2501 9243 2504 9247 2 ~clk
rlabel metal1 2499 9314 2502 9318 4 clk
rlabel metal1 2615 9205 2618 9209 1 Vdd!
rlabel metal1 2614 9148 2617 9152 1 GND!
rlabel metal1 2613 9141 2616 9145 8 ~clk
rlabel metal1 2615 9212 2618 9216 6 clk
rlabel metal2 2766 9356 2766 9356 1 Vdd!
rlabel metal2 2778 9356 2778 9356 1 GND!
rlabel metal1 3387 9102 3391 9106 1 Vdd!
rlabel metal1 3337 8951 3338 8954 3 enable
rlabel metal1 3387 8972 3391 8976 1 Vdd!
rlabel metal1 3386 9000 3390 9003 1 clk
rlabel metal1 3388 9022 3391 9026 1 GND!
rlabel metal1 3386 8870 3390 8873 1 clk
rlabel metal1 3387 8842 3391 8846 1 Vdd!
rlabel metal1 3388 8892 3391 8896 1 GND!
rlabel metal2 3676 9011 3680 9028 1 reset_b
rlabel metal2 3668 9011 3672 9028 1 Vdd!
rlabel metal2 3660 9001 3664 9018 1 GND!
rlabel metal2 3315 9121 3328 9134 1 clk
rlabel metal2 3040 9597 3053 9610 1 mode
rlabel metal1 3037 10155 3037 10155 1 p4
rlabel metal1 2723 10161 2723 10161 1 p3
rlabel metal1 3657 10154 3658 10154 1 p7
rlabel metal1 1503 10176 1505 10177 1 p6
rlabel metal1 3353 10155 3353 10155 1 p5
rlabel metal1 2426 10158 2426 10158 1 p2
rlabel metal1 2117 10166 2117 10166 1 p1
rlabel metal1 1802 10150 1806 10150 1 p0
<< end >>
