magic
tech scmos
timestamp 1608296550
<< ntransistor >>
rect 573 1706 575 1710
rect 578 1706 580 1710
rect 594 1706 596 1710
rect 610 1706 612 1710
rect 615 1706 617 1710
rect 636 1706 638 1710
rect 652 1706 654 1710
rect 668 1706 670 1710
rect 673 1706 675 1710
rect 689 1706 691 1710
rect 705 1706 707 1710
rect 710 1706 712 1710
rect 726 1706 728 1710
rect 742 1706 744 1710
rect 747 1706 749 1710
rect 768 1706 770 1710
rect 784 1706 786 1710
rect 800 1706 802 1710
rect 805 1706 807 1710
rect 821 1706 823 1710
rect 837 1706 839 1710
rect 842 1706 844 1710
rect 858 1706 860 1710
rect 874 1706 876 1710
rect 879 1706 881 1710
rect 900 1706 902 1710
rect 916 1706 918 1710
rect 932 1706 934 1710
rect 937 1706 939 1710
rect 953 1706 955 1710
rect 969 1706 971 1710
rect 974 1706 976 1710
rect 990 1706 992 1710
rect 1006 1706 1008 1710
rect 1011 1706 1013 1710
rect 1032 1706 1034 1710
rect 1048 1706 1050 1710
rect 1064 1706 1066 1710
rect 1069 1706 1071 1710
rect 1085 1706 1087 1710
rect 1506 1706 1508 1710
rect 1511 1706 1513 1710
rect 1527 1706 1529 1710
rect 1543 1706 1545 1710
rect 1548 1706 1550 1710
rect 1569 1706 1571 1710
rect 1585 1706 1587 1710
rect 1601 1706 1603 1710
rect 1606 1706 1608 1710
rect 1622 1706 1624 1710
rect 1638 1706 1640 1710
rect 1643 1706 1645 1710
rect 1659 1706 1661 1710
rect 1675 1706 1677 1710
rect 1680 1706 1682 1710
rect 1701 1706 1703 1710
rect 1717 1706 1719 1710
rect 1733 1706 1735 1710
rect 1738 1706 1740 1710
rect 1754 1706 1756 1710
rect 1770 1706 1772 1710
rect 1775 1706 1777 1710
rect 1791 1706 1793 1710
rect 1807 1706 1809 1710
rect 1812 1706 1814 1710
rect 1833 1706 1835 1710
rect 1849 1706 1851 1710
rect 1865 1706 1867 1710
rect 1870 1706 1872 1710
rect 1886 1706 1888 1710
rect 1902 1706 1904 1710
rect 1907 1706 1909 1710
rect 1923 1706 1925 1710
rect 1939 1706 1941 1710
rect 1944 1706 1946 1710
rect 1965 1706 1967 1710
rect 1981 1706 1983 1710
rect 1997 1706 1999 1710
rect 2002 1706 2004 1710
rect 2018 1706 2020 1710
rect 233 1673 235 1677
rect 238 1673 240 1677
rect 254 1673 256 1677
rect 270 1673 272 1677
rect 275 1673 277 1677
rect 296 1673 298 1677
rect 312 1673 314 1677
rect 328 1673 330 1677
rect 333 1673 335 1677
rect 349 1673 351 1677
rect 1166 1673 1168 1677
rect 1171 1673 1173 1677
rect 1187 1673 1189 1677
rect 1203 1673 1205 1677
rect 1208 1673 1210 1677
rect 1229 1673 1231 1677
rect 1245 1673 1247 1677
rect 1261 1673 1263 1677
rect 1266 1673 1268 1677
rect 1282 1673 1284 1677
rect 357 1636 359 1640
rect 752 1640 754 1644
rect 778 1636 780 1640
rect 783 1636 785 1640
rect 833 1640 835 1644
rect 859 1636 861 1640
rect 864 1636 866 1640
rect 806 1632 808 1636
rect 240 1627 242 1631
rect 578 1627 580 1631
rect 594 1627 596 1631
rect 610 1627 612 1631
rect 633 1627 635 1631
rect 638 1627 640 1631
rect 664 1627 666 1631
rect 685 1627 687 1631
rect 705 1627 707 1631
rect 710 1627 712 1631
rect 728 1627 730 1631
rect 887 1632 889 1636
rect 1290 1636 1292 1640
rect 1685 1640 1687 1644
rect 1711 1636 1713 1640
rect 1716 1636 1718 1640
rect 1766 1640 1768 1644
rect 1792 1636 1794 1640
rect 1797 1636 1799 1640
rect 1739 1632 1741 1636
rect 1173 1627 1175 1631
rect 1511 1627 1513 1631
rect 1527 1627 1529 1631
rect 1543 1627 1545 1631
rect 1566 1627 1568 1631
rect 1571 1627 1573 1631
rect 1597 1627 1599 1631
rect 1618 1627 1620 1631
rect 1638 1627 1640 1631
rect 1643 1627 1645 1631
rect 1661 1627 1663 1631
rect 1820 1632 1822 1636
rect 578 1581 580 1585
rect 594 1581 596 1585
rect 610 1581 612 1585
rect 633 1581 635 1585
rect 638 1581 640 1585
rect 664 1581 666 1585
rect 685 1581 687 1585
rect 705 1581 707 1585
rect 710 1581 712 1585
rect 728 1581 730 1585
rect 224 1571 226 1575
rect 240 1571 242 1575
rect 245 1571 247 1575
rect 261 1571 263 1575
rect 277 1571 279 1575
rect 298 1571 300 1575
rect 303 1571 305 1575
rect 319 1571 321 1575
rect 335 1571 337 1575
rect 340 1571 342 1575
rect 778 1580 780 1584
rect 783 1580 785 1584
rect 859 1580 861 1584
rect 864 1580 866 1584
rect 1511 1581 1513 1585
rect 1527 1581 1529 1585
rect 1543 1581 1545 1585
rect 1566 1581 1568 1585
rect 1571 1581 1573 1585
rect 1597 1581 1599 1585
rect 1618 1581 1620 1585
rect 1638 1581 1640 1585
rect 1643 1581 1645 1585
rect 1661 1581 1663 1585
rect 1157 1571 1159 1575
rect 1173 1571 1175 1575
rect 1178 1571 1180 1575
rect 1194 1571 1196 1575
rect 1210 1571 1212 1575
rect 1231 1571 1233 1575
rect 1236 1571 1238 1575
rect 1252 1571 1254 1575
rect 1268 1571 1270 1575
rect 1273 1571 1275 1575
rect 1711 1580 1713 1584
rect 1716 1580 1718 1584
rect 1792 1580 1794 1584
rect 1797 1580 1799 1584
rect 778 1504 780 1508
rect 783 1504 785 1508
rect 857 1508 859 1512
rect 883 1504 885 1508
rect 888 1504 890 1508
rect 806 1500 808 1504
rect 578 1495 580 1499
rect 594 1495 596 1499
rect 610 1495 612 1499
rect 633 1495 635 1499
rect 638 1495 640 1499
rect 664 1495 666 1499
rect 685 1495 687 1499
rect 705 1495 707 1499
rect 710 1495 712 1499
rect 728 1495 730 1499
rect 911 1500 913 1504
rect 1711 1504 1713 1508
rect 1716 1504 1718 1508
rect 1790 1508 1792 1512
rect 1816 1504 1818 1508
rect 1821 1504 1823 1508
rect 1739 1500 1741 1504
rect 1511 1495 1513 1499
rect 1527 1495 1529 1499
rect 1543 1495 1545 1499
rect 1566 1495 1568 1499
rect 1571 1495 1573 1499
rect 1597 1495 1599 1499
rect 1618 1495 1620 1499
rect 1638 1495 1640 1499
rect 1643 1495 1645 1499
rect 1661 1495 1663 1499
rect 1844 1500 1846 1504
rect 578 1449 580 1453
rect 594 1449 596 1453
rect 610 1449 612 1453
rect 633 1449 635 1453
rect 638 1449 640 1453
rect 664 1449 666 1453
rect 685 1449 687 1453
rect 705 1449 707 1453
rect 710 1449 712 1453
rect 728 1449 730 1453
rect 778 1449 780 1453
rect 783 1449 785 1453
rect 883 1449 885 1453
rect 888 1449 890 1453
rect 1511 1449 1513 1453
rect 1527 1449 1529 1453
rect 1543 1449 1545 1453
rect 1566 1449 1568 1453
rect 1571 1449 1573 1453
rect 1597 1449 1599 1453
rect 1618 1449 1620 1453
rect 1638 1449 1640 1453
rect 1643 1449 1645 1453
rect 1661 1449 1663 1453
rect 1711 1449 1713 1453
rect 1716 1449 1718 1453
rect 1816 1449 1818 1453
rect 1821 1449 1823 1453
rect 778 1372 780 1376
rect 783 1372 785 1376
rect 833 1376 835 1380
rect 859 1372 861 1376
rect 864 1372 866 1376
rect 923 1376 925 1380
rect 949 1372 951 1376
rect 954 1372 956 1376
rect 806 1368 808 1372
rect 578 1363 580 1367
rect 594 1363 596 1367
rect 610 1363 612 1367
rect 633 1363 635 1367
rect 638 1363 640 1367
rect 664 1363 666 1367
rect 685 1363 687 1367
rect 705 1363 707 1367
rect 710 1363 712 1367
rect 728 1363 730 1367
rect 887 1368 889 1372
rect 977 1368 979 1372
rect 1711 1372 1713 1376
rect 1716 1372 1718 1376
rect 1766 1376 1768 1380
rect 1792 1372 1794 1376
rect 1797 1372 1799 1376
rect 1856 1376 1858 1380
rect 1882 1372 1884 1376
rect 1887 1372 1889 1376
rect 1739 1368 1741 1372
rect 1511 1363 1513 1367
rect 1527 1363 1529 1367
rect 1543 1363 1545 1367
rect 1566 1363 1568 1367
rect 1571 1363 1573 1367
rect 1597 1363 1599 1367
rect 1618 1363 1620 1367
rect 1638 1363 1640 1367
rect 1643 1363 1645 1367
rect 1661 1363 1663 1367
rect 1820 1368 1822 1372
rect 1910 1368 1912 1372
rect 578 1317 580 1321
rect 594 1317 596 1321
rect 610 1317 612 1321
rect 633 1317 635 1321
rect 638 1317 640 1321
rect 664 1317 666 1321
rect 685 1317 687 1321
rect 705 1317 707 1321
rect 710 1317 712 1321
rect 728 1317 730 1321
rect 778 1314 780 1318
rect 783 1314 785 1318
rect 859 1314 861 1318
rect 864 1314 866 1318
rect 949 1314 951 1318
rect 954 1314 956 1318
rect 1511 1317 1513 1321
rect 1527 1317 1529 1321
rect 1543 1317 1545 1321
rect 1566 1317 1568 1321
rect 1571 1317 1573 1321
rect 1597 1317 1599 1321
rect 1618 1317 1620 1321
rect 1638 1317 1640 1321
rect 1643 1317 1645 1321
rect 1661 1317 1663 1321
rect 1711 1314 1713 1318
rect 1716 1314 1718 1318
rect 1792 1314 1794 1318
rect 1797 1314 1799 1318
rect 1882 1314 1884 1318
rect 1887 1314 1889 1318
rect 778 1240 780 1244
rect 783 1240 785 1244
rect 806 1236 808 1240
rect 578 1231 580 1235
rect 594 1231 596 1235
rect 610 1231 612 1235
rect 633 1231 635 1235
rect 638 1231 640 1235
rect 664 1231 666 1235
rect 685 1231 687 1235
rect 705 1231 707 1235
rect 710 1231 712 1235
rect 728 1231 730 1235
rect 1711 1240 1713 1244
rect 1716 1240 1718 1244
rect 1739 1236 1741 1240
rect 1511 1231 1513 1235
rect 1527 1231 1529 1235
rect 1543 1231 1545 1235
rect 1566 1231 1568 1235
rect 1571 1231 1573 1235
rect 1597 1231 1599 1235
rect 1618 1231 1620 1235
rect 1638 1231 1640 1235
rect 1643 1231 1645 1235
rect 1661 1231 1663 1235
rect 578 1185 580 1189
rect 594 1185 596 1189
rect 610 1185 612 1189
rect 633 1185 635 1189
rect 638 1185 640 1189
rect 664 1185 666 1189
rect 685 1185 687 1189
rect 705 1185 707 1189
rect 710 1185 712 1189
rect 728 1185 730 1189
rect 812 1185 814 1189
rect 830 1185 832 1189
rect 855 1185 857 1189
rect 871 1185 873 1189
rect 894 1185 896 1189
rect 899 1185 901 1189
rect 925 1185 927 1189
rect 946 1185 948 1189
rect 966 1185 968 1189
rect 971 1185 973 1189
rect 989 1185 991 1189
rect 101 1171 103 1175
rect 106 1171 108 1175
rect 122 1171 124 1175
rect 138 1171 140 1175
rect 143 1171 145 1175
rect 164 1171 166 1175
rect 180 1171 182 1175
rect 196 1171 198 1175
rect 201 1171 203 1175
rect 217 1171 219 1175
rect 233 1171 235 1175
rect 238 1171 240 1175
rect 254 1171 256 1175
rect 270 1171 272 1175
rect 275 1171 277 1175
rect 296 1171 298 1175
rect 312 1171 314 1175
rect 328 1171 330 1175
rect 333 1171 335 1175
rect 349 1171 351 1175
rect 365 1171 367 1175
rect 370 1171 372 1175
rect 386 1171 388 1175
rect 402 1171 404 1175
rect 407 1171 409 1175
rect 428 1171 430 1175
rect 444 1171 446 1175
rect 460 1171 462 1175
rect 465 1171 467 1175
rect 481 1171 483 1175
rect 778 1178 780 1182
rect 783 1178 785 1182
rect 1511 1185 1513 1189
rect 1527 1185 1529 1189
rect 1543 1185 1545 1189
rect 1566 1185 1568 1189
rect 1571 1185 1573 1189
rect 1597 1185 1599 1189
rect 1618 1185 1620 1189
rect 1638 1185 1640 1189
rect 1643 1185 1645 1189
rect 1661 1185 1663 1189
rect 1745 1185 1747 1189
rect 1763 1185 1765 1189
rect 1788 1185 1790 1189
rect 1804 1185 1806 1189
rect 1827 1185 1829 1189
rect 1832 1185 1834 1189
rect 1858 1185 1860 1189
rect 1879 1185 1881 1189
rect 1899 1185 1901 1189
rect 1904 1185 1906 1189
rect 1922 1185 1924 1189
rect 1034 1171 1036 1175
rect 1039 1171 1041 1175
rect 1055 1171 1057 1175
rect 1071 1171 1073 1175
rect 1076 1171 1078 1175
rect 1097 1171 1099 1175
rect 1113 1171 1115 1175
rect 1129 1171 1131 1175
rect 1134 1171 1136 1175
rect 1150 1171 1152 1175
rect 1166 1171 1168 1175
rect 1171 1171 1173 1175
rect 1187 1171 1189 1175
rect 1203 1171 1205 1175
rect 1208 1171 1210 1175
rect 1229 1171 1231 1175
rect 1245 1171 1247 1175
rect 1261 1171 1263 1175
rect 1266 1171 1268 1175
rect 1282 1171 1284 1175
rect 1298 1171 1300 1175
rect 1303 1171 1305 1175
rect 1319 1171 1321 1175
rect 1335 1171 1337 1175
rect 1340 1171 1342 1175
rect 1361 1171 1363 1175
rect 1377 1171 1379 1175
rect 1393 1171 1395 1175
rect 1398 1171 1400 1175
rect 1414 1171 1416 1175
rect 1711 1178 1713 1182
rect 1716 1178 1718 1182
rect 216 1127 218 1131
rect 240 1127 242 1131
rect 1001 1129 1005 1131
rect 1149 1127 1151 1131
rect 1173 1127 1175 1131
rect 1934 1129 1938 1131
rect 236 1116 238 1120
rect 1169 1116 1171 1120
rect 227 1102 231 1104
rect 1160 1102 1164 1104
rect 216 1093 218 1097
rect 240 1093 242 1097
rect 1149 1093 1151 1097
rect 1173 1093 1175 1097
rect 872 1061 874 1065
rect 877 1061 879 1065
rect 893 1061 895 1065
rect 909 1061 911 1065
rect 914 1061 916 1065
rect 935 1061 937 1065
rect 951 1061 953 1065
rect 967 1061 969 1065
rect 972 1061 974 1065
rect 988 1061 990 1065
rect 1805 1061 1807 1065
rect 1810 1061 1812 1065
rect 1826 1061 1828 1065
rect 1842 1061 1844 1065
rect 1847 1061 1849 1065
rect 1868 1061 1870 1065
rect 1884 1061 1886 1065
rect 1900 1061 1902 1065
rect 1905 1061 1907 1065
rect 1921 1061 1923 1065
rect 101 1031 103 1035
rect 106 1031 108 1035
rect 122 1031 124 1035
rect 138 1031 140 1035
rect 143 1031 145 1035
rect 164 1031 166 1035
rect 180 1031 182 1035
rect 196 1031 198 1035
rect 201 1031 203 1035
rect 217 1031 219 1035
rect 233 1031 235 1035
rect 238 1031 240 1035
rect 254 1031 256 1035
rect 270 1031 272 1035
rect 275 1031 277 1035
rect 296 1031 298 1035
rect 312 1031 314 1035
rect 328 1031 330 1035
rect 333 1031 335 1035
rect 349 1031 351 1035
rect 365 1031 367 1035
rect 370 1031 372 1035
rect 386 1031 388 1035
rect 402 1031 404 1035
rect 407 1031 409 1035
rect 428 1031 430 1035
rect 444 1031 446 1035
rect 460 1031 462 1035
rect 465 1031 467 1035
rect 481 1031 483 1035
rect 1034 1031 1036 1035
rect 1039 1031 1041 1035
rect 1055 1031 1057 1035
rect 1071 1031 1073 1035
rect 1076 1031 1078 1035
rect 1097 1031 1099 1035
rect 1113 1031 1115 1035
rect 1129 1031 1131 1035
rect 1134 1031 1136 1035
rect 1150 1031 1152 1035
rect 1166 1031 1168 1035
rect 1171 1031 1173 1035
rect 1187 1031 1189 1035
rect 1203 1031 1205 1035
rect 1208 1031 1210 1035
rect 1229 1031 1231 1035
rect 1245 1031 1247 1035
rect 1261 1031 1263 1035
rect 1266 1031 1268 1035
rect 1282 1031 1284 1035
rect 1298 1031 1300 1035
rect 1303 1031 1305 1035
rect 1319 1031 1321 1035
rect 1335 1031 1337 1035
rect 1340 1031 1342 1035
rect 1361 1031 1363 1035
rect 1377 1031 1379 1035
rect 1393 1031 1395 1035
rect 1398 1031 1400 1035
rect 1414 1031 1416 1035
rect 1013 985 1017 987
rect 1946 985 1950 987
rect 872 975 874 979
rect 877 975 879 979
rect 893 975 895 979
rect 909 975 911 979
rect 914 975 916 979
rect 935 975 937 979
rect 951 975 953 979
rect 967 975 969 979
rect 972 975 974 979
rect 988 975 990 979
rect 1805 975 1807 979
rect 1810 975 1812 979
rect 1826 975 1828 979
rect 1842 975 1844 979
rect 1847 975 1849 979
rect 1868 975 1870 979
rect 1884 975 1886 979
rect 1900 975 1902 979
rect 1905 975 1907 979
rect 1921 975 1923 979
rect 101 945 103 949
rect 106 945 108 949
rect 122 945 124 949
rect 138 945 140 949
rect 143 945 145 949
rect 164 945 166 949
rect 180 945 182 949
rect 196 945 198 949
rect 201 945 203 949
rect 217 945 219 949
rect 233 945 235 949
rect 238 945 240 949
rect 254 945 256 949
rect 270 945 272 949
rect 275 945 277 949
rect 296 945 298 949
rect 312 945 314 949
rect 328 945 330 949
rect 333 945 335 949
rect 349 945 351 949
rect 365 945 367 949
rect 370 945 372 949
rect 386 945 388 949
rect 402 945 404 949
rect 407 945 409 949
rect 428 945 430 949
rect 444 945 446 949
rect 460 945 462 949
rect 465 945 467 949
rect 481 945 483 949
rect 1034 945 1036 949
rect 1039 945 1041 949
rect 1055 945 1057 949
rect 1071 945 1073 949
rect 1076 945 1078 949
rect 1097 945 1099 949
rect 1113 945 1115 949
rect 1129 945 1131 949
rect 1134 945 1136 949
rect 1150 945 1152 949
rect 1166 945 1168 949
rect 1171 945 1173 949
rect 1187 945 1189 949
rect 1203 945 1205 949
rect 1208 945 1210 949
rect 1229 945 1231 949
rect 1245 945 1247 949
rect 1261 945 1263 949
rect 1266 945 1268 949
rect 1282 945 1284 949
rect 1298 945 1300 949
rect 1303 945 1305 949
rect 1319 945 1321 949
rect 1335 945 1337 949
rect 1340 945 1342 949
rect 1361 945 1363 949
rect 1377 945 1379 949
rect 1393 945 1395 949
rect 1398 945 1400 949
rect 1414 945 1416 949
rect 333 901 335 905
rect 357 901 359 905
rect 1266 901 1268 905
rect 1290 901 1292 905
rect 353 890 355 894
rect 1286 890 1288 894
rect 344 876 348 878
rect 1277 876 1281 878
rect 333 867 335 871
rect 357 867 359 871
rect 1266 867 1268 871
rect 1290 867 1292 871
rect 101 805 103 809
rect 106 805 108 809
rect 122 805 124 809
rect 138 805 140 809
rect 143 805 145 809
rect 164 805 166 809
rect 180 805 182 809
rect 196 805 198 809
rect 201 805 203 809
rect 217 805 219 809
rect 233 805 235 809
rect 238 805 240 809
rect 254 805 256 809
rect 270 805 272 809
rect 275 805 277 809
rect 296 805 298 809
rect 312 805 314 809
rect 328 805 330 809
rect 333 805 335 809
rect 349 805 351 809
rect 365 805 367 809
rect 370 805 372 809
rect 386 805 388 809
rect 402 805 404 809
rect 407 805 409 809
rect 428 805 430 809
rect 444 805 446 809
rect 460 805 462 809
rect 465 805 467 809
rect 481 805 483 809
rect 1034 805 1036 809
rect 1039 805 1041 809
rect 1055 805 1057 809
rect 1071 805 1073 809
rect 1076 805 1078 809
rect 1097 805 1099 809
rect 1113 805 1115 809
rect 1129 805 1131 809
rect 1134 805 1136 809
rect 1150 805 1152 809
rect 1166 805 1168 809
rect 1171 805 1173 809
rect 1187 805 1189 809
rect 1203 805 1205 809
rect 1208 805 1210 809
rect 1229 805 1231 809
rect 1245 805 1247 809
rect 1261 805 1263 809
rect 1266 805 1268 809
rect 1282 805 1284 809
rect 1298 805 1300 809
rect 1303 805 1305 809
rect 1319 805 1321 809
rect 1335 805 1337 809
rect 1340 805 1342 809
rect 1361 805 1363 809
rect 1377 805 1379 809
rect 1393 805 1395 809
rect 1398 805 1400 809
rect 1414 805 1416 809
rect 573 726 575 730
rect 578 726 580 730
rect 594 726 596 730
rect 610 726 612 730
rect 615 726 617 730
rect 636 726 638 730
rect 652 726 654 730
rect 668 726 670 730
rect 673 726 675 730
rect 689 726 691 730
rect 705 726 707 730
rect 710 726 712 730
rect 726 726 728 730
rect 742 726 744 730
rect 747 726 749 730
rect 768 726 770 730
rect 784 726 786 730
rect 800 726 802 730
rect 805 726 807 730
rect 821 726 823 730
rect 837 726 839 730
rect 842 726 844 730
rect 858 726 860 730
rect 874 726 876 730
rect 879 726 881 730
rect 900 726 902 730
rect 916 726 918 730
rect 932 726 934 730
rect 937 726 939 730
rect 953 726 955 730
rect 969 726 971 730
rect 974 726 976 730
rect 990 726 992 730
rect 1006 726 1008 730
rect 1011 726 1013 730
rect 1032 726 1034 730
rect 1048 726 1050 730
rect 1064 726 1066 730
rect 1069 726 1071 730
rect 1085 726 1087 730
rect 1506 726 1508 730
rect 1511 726 1513 730
rect 1527 726 1529 730
rect 1543 726 1545 730
rect 1548 726 1550 730
rect 1569 726 1571 730
rect 1585 726 1587 730
rect 1601 726 1603 730
rect 1606 726 1608 730
rect 1622 726 1624 730
rect 1638 726 1640 730
rect 1643 726 1645 730
rect 1659 726 1661 730
rect 1675 726 1677 730
rect 1680 726 1682 730
rect 1701 726 1703 730
rect 1717 726 1719 730
rect 1733 726 1735 730
rect 1738 726 1740 730
rect 1754 726 1756 730
rect 1770 726 1772 730
rect 1775 726 1777 730
rect 1791 726 1793 730
rect 1807 726 1809 730
rect 1812 726 1814 730
rect 1833 726 1835 730
rect 1849 726 1851 730
rect 1865 726 1867 730
rect 1870 726 1872 730
rect 1886 726 1888 730
rect 1902 726 1904 730
rect 1907 726 1909 730
rect 1923 726 1925 730
rect 1939 726 1941 730
rect 1944 726 1946 730
rect 1965 726 1967 730
rect 1981 726 1983 730
rect 1997 726 1999 730
rect 2002 726 2004 730
rect 2018 726 2020 730
rect 233 693 235 697
rect 238 693 240 697
rect 254 693 256 697
rect 270 693 272 697
rect 275 693 277 697
rect 296 693 298 697
rect 312 693 314 697
rect 328 693 330 697
rect 333 693 335 697
rect 349 693 351 697
rect 1166 693 1168 697
rect 1171 693 1173 697
rect 1187 693 1189 697
rect 1203 693 1205 697
rect 1208 693 1210 697
rect 1229 693 1231 697
rect 1245 693 1247 697
rect 1261 693 1263 697
rect 1266 693 1268 697
rect 1282 693 1284 697
rect 357 656 359 660
rect 752 660 754 664
rect 778 656 780 660
rect 783 656 785 660
rect 833 660 835 664
rect 859 656 861 660
rect 864 656 866 660
rect 806 652 808 656
rect 240 647 242 651
rect 578 647 580 651
rect 594 647 596 651
rect 610 647 612 651
rect 633 647 635 651
rect 638 647 640 651
rect 664 647 666 651
rect 685 647 687 651
rect 705 647 707 651
rect 710 647 712 651
rect 728 647 730 651
rect 887 652 889 656
rect 1290 656 1292 660
rect 1685 660 1687 664
rect 1711 656 1713 660
rect 1716 656 1718 660
rect 1766 660 1768 664
rect 1792 656 1794 660
rect 1797 656 1799 660
rect 1739 652 1741 656
rect 1173 647 1175 651
rect 1511 647 1513 651
rect 1527 647 1529 651
rect 1543 647 1545 651
rect 1566 647 1568 651
rect 1571 647 1573 651
rect 1597 647 1599 651
rect 1618 647 1620 651
rect 1638 647 1640 651
rect 1643 647 1645 651
rect 1661 647 1663 651
rect 1820 652 1822 656
rect 578 601 580 605
rect 594 601 596 605
rect 610 601 612 605
rect 633 601 635 605
rect 638 601 640 605
rect 664 601 666 605
rect 685 601 687 605
rect 705 601 707 605
rect 710 601 712 605
rect 728 601 730 605
rect 224 591 226 595
rect 240 591 242 595
rect 245 591 247 595
rect 261 591 263 595
rect 277 591 279 595
rect 298 591 300 595
rect 303 591 305 595
rect 319 591 321 595
rect 335 591 337 595
rect 340 591 342 595
rect 778 600 780 604
rect 783 600 785 604
rect 859 600 861 604
rect 864 600 866 604
rect 1511 601 1513 605
rect 1527 601 1529 605
rect 1543 601 1545 605
rect 1566 601 1568 605
rect 1571 601 1573 605
rect 1597 601 1599 605
rect 1618 601 1620 605
rect 1638 601 1640 605
rect 1643 601 1645 605
rect 1661 601 1663 605
rect 1157 591 1159 595
rect 1173 591 1175 595
rect 1178 591 1180 595
rect 1194 591 1196 595
rect 1210 591 1212 595
rect 1231 591 1233 595
rect 1236 591 1238 595
rect 1252 591 1254 595
rect 1268 591 1270 595
rect 1273 591 1275 595
rect 1711 600 1713 604
rect 1716 600 1718 604
rect 1792 600 1794 604
rect 1797 600 1799 604
rect 778 524 780 528
rect 783 524 785 528
rect 857 528 859 532
rect 883 524 885 528
rect 888 524 890 528
rect 806 520 808 524
rect 578 515 580 519
rect 594 515 596 519
rect 610 515 612 519
rect 633 515 635 519
rect 638 515 640 519
rect 664 515 666 519
rect 685 515 687 519
rect 705 515 707 519
rect 710 515 712 519
rect 728 515 730 519
rect 911 520 913 524
rect 1711 524 1713 528
rect 1716 524 1718 528
rect 1790 528 1792 532
rect 1816 524 1818 528
rect 1821 524 1823 528
rect 1739 520 1741 524
rect 1511 515 1513 519
rect 1527 515 1529 519
rect 1543 515 1545 519
rect 1566 515 1568 519
rect 1571 515 1573 519
rect 1597 515 1599 519
rect 1618 515 1620 519
rect 1638 515 1640 519
rect 1643 515 1645 519
rect 1661 515 1663 519
rect 1844 520 1846 524
rect 578 469 580 473
rect 594 469 596 473
rect 610 469 612 473
rect 633 469 635 473
rect 638 469 640 473
rect 664 469 666 473
rect 685 469 687 473
rect 705 469 707 473
rect 710 469 712 473
rect 728 469 730 473
rect 778 469 780 473
rect 783 469 785 473
rect 883 469 885 473
rect 888 469 890 473
rect 1511 469 1513 473
rect 1527 469 1529 473
rect 1543 469 1545 473
rect 1566 469 1568 473
rect 1571 469 1573 473
rect 1597 469 1599 473
rect 1618 469 1620 473
rect 1638 469 1640 473
rect 1643 469 1645 473
rect 1661 469 1663 473
rect 1711 469 1713 473
rect 1716 469 1718 473
rect 1816 469 1818 473
rect 1821 469 1823 473
rect 778 392 780 396
rect 783 392 785 396
rect 833 396 835 400
rect 859 392 861 396
rect 864 392 866 396
rect 923 396 925 400
rect 949 392 951 396
rect 954 392 956 396
rect 806 388 808 392
rect 578 383 580 387
rect 594 383 596 387
rect 610 383 612 387
rect 633 383 635 387
rect 638 383 640 387
rect 664 383 666 387
rect 685 383 687 387
rect 705 383 707 387
rect 710 383 712 387
rect 728 383 730 387
rect 887 388 889 392
rect 977 388 979 392
rect 1711 392 1713 396
rect 1716 392 1718 396
rect 1766 396 1768 400
rect 1792 392 1794 396
rect 1797 392 1799 396
rect 1856 396 1858 400
rect 1882 392 1884 396
rect 1887 392 1889 396
rect 1739 388 1741 392
rect 1511 383 1513 387
rect 1527 383 1529 387
rect 1543 383 1545 387
rect 1566 383 1568 387
rect 1571 383 1573 387
rect 1597 383 1599 387
rect 1618 383 1620 387
rect 1638 383 1640 387
rect 1643 383 1645 387
rect 1661 383 1663 387
rect 1820 388 1822 392
rect 1910 388 1912 392
rect 578 337 580 341
rect 594 337 596 341
rect 610 337 612 341
rect 633 337 635 341
rect 638 337 640 341
rect 664 337 666 341
rect 685 337 687 341
rect 705 337 707 341
rect 710 337 712 341
rect 728 337 730 341
rect 778 334 780 338
rect 783 334 785 338
rect 859 334 861 338
rect 864 334 866 338
rect 949 334 951 338
rect 954 334 956 338
rect 1511 337 1513 341
rect 1527 337 1529 341
rect 1543 337 1545 341
rect 1566 337 1568 341
rect 1571 337 1573 341
rect 1597 337 1599 341
rect 1618 337 1620 341
rect 1638 337 1640 341
rect 1643 337 1645 341
rect 1661 337 1663 341
rect 1711 334 1713 338
rect 1716 334 1718 338
rect 1792 334 1794 338
rect 1797 334 1799 338
rect 1882 334 1884 338
rect 1887 334 1889 338
rect 778 260 780 264
rect 783 260 785 264
rect 806 256 808 260
rect 578 251 580 255
rect 594 251 596 255
rect 610 251 612 255
rect 633 251 635 255
rect 638 251 640 255
rect 664 251 666 255
rect 685 251 687 255
rect 705 251 707 255
rect 710 251 712 255
rect 728 251 730 255
rect 1711 260 1713 264
rect 1716 260 1718 264
rect 1739 256 1741 260
rect 1511 251 1513 255
rect 1527 251 1529 255
rect 1543 251 1545 255
rect 1566 251 1568 255
rect 1571 251 1573 255
rect 1597 251 1599 255
rect 1618 251 1620 255
rect 1638 251 1640 255
rect 1643 251 1645 255
rect 1661 251 1663 255
rect 578 205 580 209
rect 594 205 596 209
rect 610 205 612 209
rect 633 205 635 209
rect 638 205 640 209
rect 664 205 666 209
rect 685 205 687 209
rect 705 205 707 209
rect 710 205 712 209
rect 728 205 730 209
rect 812 205 814 209
rect 830 205 832 209
rect 855 205 857 209
rect 871 205 873 209
rect 894 205 896 209
rect 899 205 901 209
rect 925 205 927 209
rect 946 205 948 209
rect 966 205 968 209
rect 971 205 973 209
rect 989 205 991 209
rect 101 191 103 195
rect 106 191 108 195
rect 122 191 124 195
rect 138 191 140 195
rect 143 191 145 195
rect 164 191 166 195
rect 180 191 182 195
rect 196 191 198 195
rect 201 191 203 195
rect 217 191 219 195
rect 233 191 235 195
rect 238 191 240 195
rect 254 191 256 195
rect 270 191 272 195
rect 275 191 277 195
rect 296 191 298 195
rect 312 191 314 195
rect 328 191 330 195
rect 333 191 335 195
rect 349 191 351 195
rect 365 191 367 195
rect 370 191 372 195
rect 386 191 388 195
rect 402 191 404 195
rect 407 191 409 195
rect 428 191 430 195
rect 444 191 446 195
rect 460 191 462 195
rect 465 191 467 195
rect 481 191 483 195
rect 778 198 780 202
rect 783 198 785 202
rect 1511 205 1513 209
rect 1527 205 1529 209
rect 1543 205 1545 209
rect 1566 205 1568 209
rect 1571 205 1573 209
rect 1597 205 1599 209
rect 1618 205 1620 209
rect 1638 205 1640 209
rect 1643 205 1645 209
rect 1661 205 1663 209
rect 1745 205 1747 209
rect 1763 205 1765 209
rect 1788 205 1790 209
rect 1804 205 1806 209
rect 1827 205 1829 209
rect 1832 205 1834 209
rect 1858 205 1860 209
rect 1879 205 1881 209
rect 1899 205 1901 209
rect 1904 205 1906 209
rect 1922 205 1924 209
rect 1034 191 1036 195
rect 1039 191 1041 195
rect 1055 191 1057 195
rect 1071 191 1073 195
rect 1076 191 1078 195
rect 1097 191 1099 195
rect 1113 191 1115 195
rect 1129 191 1131 195
rect 1134 191 1136 195
rect 1150 191 1152 195
rect 1166 191 1168 195
rect 1171 191 1173 195
rect 1187 191 1189 195
rect 1203 191 1205 195
rect 1208 191 1210 195
rect 1229 191 1231 195
rect 1245 191 1247 195
rect 1261 191 1263 195
rect 1266 191 1268 195
rect 1282 191 1284 195
rect 1298 191 1300 195
rect 1303 191 1305 195
rect 1319 191 1321 195
rect 1335 191 1337 195
rect 1340 191 1342 195
rect 1361 191 1363 195
rect 1377 191 1379 195
rect 1393 191 1395 195
rect 1398 191 1400 195
rect 1414 191 1416 195
rect 1711 198 1713 202
rect 1716 198 1718 202
rect 216 147 218 151
rect 240 147 242 151
rect 1001 149 1005 151
rect 1149 147 1151 151
rect 1173 147 1175 151
rect 1934 149 1938 151
rect 236 136 238 140
rect 1169 136 1171 140
rect 227 122 231 124
rect 1160 122 1164 124
rect 216 113 218 117
rect 240 113 242 117
rect 1149 113 1151 117
rect 1173 113 1175 117
rect 872 81 874 85
rect 877 81 879 85
rect 893 81 895 85
rect 909 81 911 85
rect 914 81 916 85
rect 935 81 937 85
rect 951 81 953 85
rect 967 81 969 85
rect 972 81 974 85
rect 988 81 990 85
rect 1805 81 1807 85
rect 1810 81 1812 85
rect 1826 81 1828 85
rect 1842 81 1844 85
rect 1847 81 1849 85
rect 1868 81 1870 85
rect 1884 81 1886 85
rect 1900 81 1902 85
rect 1905 81 1907 85
rect 1921 81 1923 85
rect 101 51 103 55
rect 106 51 108 55
rect 122 51 124 55
rect 138 51 140 55
rect 143 51 145 55
rect 164 51 166 55
rect 180 51 182 55
rect 196 51 198 55
rect 201 51 203 55
rect 217 51 219 55
rect 233 51 235 55
rect 238 51 240 55
rect 254 51 256 55
rect 270 51 272 55
rect 275 51 277 55
rect 296 51 298 55
rect 312 51 314 55
rect 328 51 330 55
rect 333 51 335 55
rect 349 51 351 55
rect 365 51 367 55
rect 370 51 372 55
rect 386 51 388 55
rect 402 51 404 55
rect 407 51 409 55
rect 428 51 430 55
rect 444 51 446 55
rect 460 51 462 55
rect 465 51 467 55
rect 481 51 483 55
rect 1034 51 1036 55
rect 1039 51 1041 55
rect 1055 51 1057 55
rect 1071 51 1073 55
rect 1076 51 1078 55
rect 1097 51 1099 55
rect 1113 51 1115 55
rect 1129 51 1131 55
rect 1134 51 1136 55
rect 1150 51 1152 55
rect 1166 51 1168 55
rect 1171 51 1173 55
rect 1187 51 1189 55
rect 1203 51 1205 55
rect 1208 51 1210 55
rect 1229 51 1231 55
rect 1245 51 1247 55
rect 1261 51 1263 55
rect 1266 51 1268 55
rect 1282 51 1284 55
rect 1298 51 1300 55
rect 1303 51 1305 55
rect 1319 51 1321 55
rect 1335 51 1337 55
rect 1340 51 1342 55
rect 1361 51 1363 55
rect 1377 51 1379 55
rect 1393 51 1395 55
rect 1398 51 1400 55
rect 1414 51 1416 55
rect 1013 5 1017 7
rect 1946 5 1950 7
rect 872 -5 874 -1
rect 877 -5 879 -1
rect 893 -5 895 -1
rect 909 -5 911 -1
rect 914 -5 916 -1
rect 935 -5 937 -1
rect 951 -5 953 -1
rect 967 -5 969 -1
rect 972 -5 974 -1
rect 988 -5 990 -1
rect 1805 -5 1807 -1
rect 1810 -5 1812 -1
rect 1826 -5 1828 -1
rect 1842 -5 1844 -1
rect 1847 -5 1849 -1
rect 1868 -5 1870 -1
rect 1884 -5 1886 -1
rect 1900 -5 1902 -1
rect 1905 -5 1907 -1
rect 1921 -5 1923 -1
rect 101 -35 103 -31
rect 106 -35 108 -31
rect 122 -35 124 -31
rect 138 -35 140 -31
rect 143 -35 145 -31
rect 164 -35 166 -31
rect 180 -35 182 -31
rect 196 -35 198 -31
rect 201 -35 203 -31
rect 217 -35 219 -31
rect 233 -35 235 -31
rect 238 -35 240 -31
rect 254 -35 256 -31
rect 270 -35 272 -31
rect 275 -35 277 -31
rect 296 -35 298 -31
rect 312 -35 314 -31
rect 328 -35 330 -31
rect 333 -35 335 -31
rect 349 -35 351 -31
rect 365 -35 367 -31
rect 370 -35 372 -31
rect 386 -35 388 -31
rect 402 -35 404 -31
rect 407 -35 409 -31
rect 428 -35 430 -31
rect 444 -35 446 -31
rect 460 -35 462 -31
rect 465 -35 467 -31
rect 481 -35 483 -31
rect 1034 -35 1036 -31
rect 1039 -35 1041 -31
rect 1055 -35 1057 -31
rect 1071 -35 1073 -31
rect 1076 -35 1078 -31
rect 1097 -35 1099 -31
rect 1113 -35 1115 -31
rect 1129 -35 1131 -31
rect 1134 -35 1136 -31
rect 1150 -35 1152 -31
rect 1166 -35 1168 -31
rect 1171 -35 1173 -31
rect 1187 -35 1189 -31
rect 1203 -35 1205 -31
rect 1208 -35 1210 -31
rect 1229 -35 1231 -31
rect 1245 -35 1247 -31
rect 1261 -35 1263 -31
rect 1266 -35 1268 -31
rect 1282 -35 1284 -31
rect 1298 -35 1300 -31
rect 1303 -35 1305 -31
rect 1319 -35 1321 -31
rect 1335 -35 1337 -31
rect 1340 -35 1342 -31
rect 1361 -35 1363 -31
rect 1377 -35 1379 -31
rect 1393 -35 1395 -31
rect 1398 -35 1400 -31
rect 1414 -35 1416 -31
rect 333 -79 335 -75
rect 357 -79 359 -75
rect 1266 -79 1268 -75
rect 1290 -79 1292 -75
rect 353 -90 355 -86
rect 1286 -90 1288 -86
rect 344 -104 348 -102
rect 1277 -104 1281 -102
rect 333 -113 335 -109
rect 357 -113 359 -109
rect 1266 -113 1268 -109
rect 1290 -113 1292 -109
rect 101 -175 103 -171
rect 106 -175 108 -171
rect 122 -175 124 -171
rect 138 -175 140 -171
rect 143 -175 145 -171
rect 164 -175 166 -171
rect 180 -175 182 -171
rect 196 -175 198 -171
rect 201 -175 203 -171
rect 217 -175 219 -171
rect 233 -175 235 -171
rect 238 -175 240 -171
rect 254 -175 256 -171
rect 270 -175 272 -171
rect 275 -175 277 -171
rect 296 -175 298 -171
rect 312 -175 314 -171
rect 328 -175 330 -171
rect 333 -175 335 -171
rect 349 -175 351 -171
rect 365 -175 367 -171
rect 370 -175 372 -171
rect 386 -175 388 -171
rect 402 -175 404 -171
rect 407 -175 409 -171
rect 428 -175 430 -171
rect 444 -175 446 -171
rect 460 -175 462 -171
rect 465 -175 467 -171
rect 481 -175 483 -171
rect 1034 -175 1036 -171
rect 1039 -175 1041 -171
rect 1055 -175 1057 -171
rect 1071 -175 1073 -171
rect 1076 -175 1078 -171
rect 1097 -175 1099 -171
rect 1113 -175 1115 -171
rect 1129 -175 1131 -171
rect 1134 -175 1136 -171
rect 1150 -175 1152 -171
rect 1166 -175 1168 -171
rect 1171 -175 1173 -171
rect 1187 -175 1189 -171
rect 1203 -175 1205 -171
rect 1208 -175 1210 -171
rect 1229 -175 1231 -171
rect 1245 -175 1247 -171
rect 1261 -175 1263 -171
rect 1266 -175 1268 -171
rect 1282 -175 1284 -171
rect 1298 -175 1300 -171
rect 1303 -175 1305 -171
rect 1319 -175 1321 -171
rect 1335 -175 1337 -171
rect 1340 -175 1342 -171
rect 1361 -175 1363 -171
rect 1377 -175 1379 -171
rect 1393 -175 1395 -171
rect 1398 -175 1400 -171
rect 1414 -175 1416 -171
<< ptransistor >>
rect 573 1729 575 1737
rect 578 1729 580 1737
rect 594 1729 596 1737
rect 610 1729 612 1737
rect 615 1729 617 1737
rect 636 1729 638 1737
rect 652 1729 654 1737
rect 668 1729 670 1737
rect 673 1729 675 1737
rect 689 1729 691 1737
rect 705 1729 707 1737
rect 710 1729 712 1737
rect 726 1729 728 1737
rect 742 1729 744 1737
rect 747 1729 749 1737
rect 768 1729 770 1737
rect 784 1729 786 1737
rect 800 1729 802 1737
rect 805 1729 807 1737
rect 821 1729 823 1737
rect 837 1729 839 1737
rect 842 1729 844 1737
rect 858 1729 860 1737
rect 874 1729 876 1737
rect 879 1729 881 1737
rect 900 1729 902 1737
rect 916 1729 918 1737
rect 932 1729 934 1737
rect 937 1729 939 1737
rect 953 1729 955 1737
rect 969 1729 971 1737
rect 974 1729 976 1737
rect 990 1729 992 1737
rect 1006 1729 1008 1737
rect 1011 1729 1013 1737
rect 1032 1729 1034 1737
rect 1048 1729 1050 1737
rect 1064 1729 1066 1737
rect 1069 1729 1071 1737
rect 1085 1729 1087 1737
rect 1506 1729 1508 1737
rect 1511 1729 1513 1737
rect 1527 1729 1529 1737
rect 1543 1729 1545 1737
rect 1548 1729 1550 1737
rect 1569 1729 1571 1737
rect 1585 1729 1587 1737
rect 1601 1729 1603 1737
rect 1606 1729 1608 1737
rect 1622 1729 1624 1737
rect 1638 1729 1640 1737
rect 1643 1729 1645 1737
rect 1659 1729 1661 1737
rect 1675 1729 1677 1737
rect 1680 1729 1682 1737
rect 1701 1729 1703 1737
rect 1717 1729 1719 1737
rect 1733 1729 1735 1737
rect 1738 1729 1740 1737
rect 1754 1729 1756 1737
rect 1770 1729 1772 1737
rect 1775 1729 1777 1737
rect 1791 1729 1793 1737
rect 1807 1729 1809 1737
rect 1812 1729 1814 1737
rect 1833 1729 1835 1737
rect 1849 1729 1851 1737
rect 1865 1729 1867 1737
rect 1870 1729 1872 1737
rect 1886 1729 1888 1737
rect 1902 1729 1904 1737
rect 1907 1729 1909 1737
rect 1923 1729 1925 1737
rect 1939 1729 1941 1737
rect 1944 1729 1946 1737
rect 1965 1729 1967 1737
rect 1981 1729 1983 1737
rect 1997 1729 1999 1737
rect 2002 1729 2004 1737
rect 2018 1729 2020 1737
rect 233 1696 235 1704
rect 238 1696 240 1704
rect 254 1696 256 1704
rect 270 1696 272 1704
rect 275 1696 277 1704
rect 296 1696 298 1704
rect 312 1696 314 1704
rect 328 1696 330 1704
rect 333 1696 335 1704
rect 349 1696 351 1704
rect 1166 1696 1168 1704
rect 1171 1696 1173 1704
rect 1187 1696 1189 1704
rect 1203 1696 1205 1704
rect 1208 1696 1210 1704
rect 1229 1696 1231 1704
rect 1245 1696 1247 1704
rect 1261 1696 1263 1704
rect 1266 1696 1268 1704
rect 1282 1696 1284 1704
rect 752 1658 754 1666
rect 578 1645 580 1653
rect 594 1645 596 1653
rect 610 1645 612 1653
rect 633 1645 635 1653
rect 638 1645 640 1653
rect 664 1645 666 1653
rect 685 1645 687 1653
rect 705 1645 707 1653
rect 710 1645 712 1653
rect 728 1645 730 1653
rect 778 1652 780 1660
rect 783 1652 785 1660
rect 806 1658 808 1666
rect 833 1658 835 1666
rect 859 1652 861 1660
rect 864 1652 866 1660
rect 887 1658 889 1666
rect 1685 1658 1687 1666
rect 1511 1645 1513 1653
rect 1527 1645 1529 1653
rect 1543 1645 1545 1653
rect 1566 1645 1568 1653
rect 1571 1645 1573 1653
rect 1597 1645 1599 1653
rect 1618 1645 1620 1653
rect 1638 1645 1640 1653
rect 1643 1645 1645 1653
rect 1661 1645 1663 1653
rect 1711 1652 1713 1660
rect 1716 1652 1718 1660
rect 1739 1658 1741 1666
rect 1766 1658 1768 1666
rect 1792 1652 1794 1660
rect 1797 1652 1799 1660
rect 1820 1658 1822 1666
rect 224 1594 226 1602
rect 240 1594 242 1602
rect 245 1594 247 1602
rect 261 1594 263 1602
rect 277 1594 279 1602
rect 298 1594 300 1602
rect 303 1594 305 1602
rect 319 1594 321 1602
rect 335 1594 337 1602
rect 340 1594 342 1602
rect 1157 1594 1159 1602
rect 1173 1594 1175 1602
rect 1178 1594 1180 1602
rect 1194 1594 1196 1602
rect 1210 1594 1212 1602
rect 1231 1594 1233 1602
rect 1236 1594 1238 1602
rect 1252 1594 1254 1602
rect 1268 1594 1270 1602
rect 1273 1594 1275 1602
rect 578 1559 580 1567
rect 594 1559 596 1567
rect 610 1559 612 1567
rect 633 1559 635 1567
rect 638 1559 640 1567
rect 664 1559 666 1567
rect 685 1559 687 1567
rect 705 1559 707 1567
rect 710 1559 712 1567
rect 728 1559 730 1567
rect 778 1560 780 1568
rect 783 1560 785 1568
rect 859 1560 861 1568
rect 864 1560 866 1568
rect 1511 1559 1513 1567
rect 1527 1559 1529 1567
rect 1543 1559 1545 1567
rect 1566 1559 1568 1567
rect 1571 1559 1573 1567
rect 1597 1559 1599 1567
rect 1618 1559 1620 1567
rect 1638 1559 1640 1567
rect 1643 1559 1645 1567
rect 1661 1559 1663 1567
rect 1711 1560 1713 1568
rect 1716 1560 1718 1568
rect 1792 1560 1794 1568
rect 1797 1560 1799 1568
rect 578 1513 580 1521
rect 594 1513 596 1521
rect 610 1513 612 1521
rect 633 1513 635 1521
rect 638 1513 640 1521
rect 664 1513 666 1521
rect 685 1513 687 1521
rect 705 1513 707 1521
rect 710 1513 712 1521
rect 728 1513 730 1521
rect 778 1520 780 1528
rect 783 1520 785 1528
rect 806 1526 808 1534
rect 857 1526 859 1534
rect 883 1520 885 1528
rect 888 1520 890 1528
rect 911 1526 913 1534
rect 1511 1513 1513 1521
rect 1527 1513 1529 1521
rect 1543 1513 1545 1521
rect 1566 1513 1568 1521
rect 1571 1513 1573 1521
rect 1597 1513 1599 1521
rect 1618 1513 1620 1521
rect 1638 1513 1640 1521
rect 1643 1513 1645 1521
rect 1661 1513 1663 1521
rect 1711 1520 1713 1528
rect 1716 1520 1718 1528
rect 1739 1526 1741 1534
rect 1790 1526 1792 1534
rect 1816 1520 1818 1528
rect 1821 1520 1823 1528
rect 1844 1526 1846 1534
rect 578 1427 580 1435
rect 594 1427 596 1435
rect 610 1427 612 1435
rect 633 1427 635 1435
rect 638 1427 640 1435
rect 664 1427 666 1435
rect 685 1427 687 1435
rect 705 1427 707 1435
rect 710 1427 712 1435
rect 728 1427 730 1435
rect 778 1429 780 1437
rect 783 1429 785 1437
rect 883 1429 885 1437
rect 888 1429 890 1437
rect 1511 1427 1513 1435
rect 1527 1427 1529 1435
rect 1543 1427 1545 1435
rect 1566 1427 1568 1435
rect 1571 1427 1573 1435
rect 1597 1427 1599 1435
rect 1618 1427 1620 1435
rect 1638 1427 1640 1435
rect 1643 1427 1645 1435
rect 1661 1427 1663 1435
rect 1711 1429 1713 1437
rect 1716 1429 1718 1437
rect 1816 1429 1818 1437
rect 1821 1429 1823 1437
rect 578 1381 580 1389
rect 594 1381 596 1389
rect 610 1381 612 1389
rect 633 1381 635 1389
rect 638 1381 640 1389
rect 664 1381 666 1389
rect 685 1381 687 1389
rect 705 1381 707 1389
rect 710 1381 712 1389
rect 728 1381 730 1389
rect 778 1388 780 1396
rect 783 1388 785 1396
rect 806 1394 808 1402
rect 833 1394 835 1402
rect 859 1388 861 1396
rect 864 1388 866 1396
rect 887 1394 889 1402
rect 923 1394 925 1402
rect 949 1388 951 1396
rect 954 1388 956 1396
rect 977 1394 979 1402
rect 1511 1381 1513 1389
rect 1527 1381 1529 1389
rect 1543 1381 1545 1389
rect 1566 1381 1568 1389
rect 1571 1381 1573 1389
rect 1597 1381 1599 1389
rect 1618 1381 1620 1389
rect 1638 1381 1640 1389
rect 1643 1381 1645 1389
rect 1661 1381 1663 1389
rect 1711 1388 1713 1396
rect 1716 1388 1718 1396
rect 1739 1394 1741 1402
rect 1766 1394 1768 1402
rect 1792 1388 1794 1396
rect 1797 1388 1799 1396
rect 1820 1394 1822 1402
rect 1856 1394 1858 1402
rect 1882 1388 1884 1396
rect 1887 1388 1889 1396
rect 1910 1394 1912 1402
rect 578 1295 580 1303
rect 594 1295 596 1303
rect 610 1295 612 1303
rect 633 1295 635 1303
rect 638 1295 640 1303
rect 664 1295 666 1303
rect 685 1295 687 1303
rect 705 1295 707 1303
rect 710 1295 712 1303
rect 728 1295 730 1303
rect 778 1294 780 1302
rect 783 1294 785 1302
rect 859 1294 861 1302
rect 864 1294 866 1302
rect 949 1294 951 1302
rect 954 1294 956 1302
rect 1511 1295 1513 1303
rect 1527 1295 1529 1303
rect 1543 1295 1545 1303
rect 1566 1295 1568 1303
rect 1571 1295 1573 1303
rect 1597 1295 1599 1303
rect 1618 1295 1620 1303
rect 1638 1295 1640 1303
rect 1643 1295 1645 1303
rect 1661 1295 1663 1303
rect 1711 1294 1713 1302
rect 1716 1294 1718 1302
rect 1792 1294 1794 1302
rect 1797 1294 1799 1302
rect 1882 1294 1884 1302
rect 1887 1294 1889 1302
rect 578 1249 580 1257
rect 594 1249 596 1257
rect 610 1249 612 1257
rect 633 1249 635 1257
rect 638 1249 640 1257
rect 664 1249 666 1257
rect 685 1249 687 1257
rect 705 1249 707 1257
rect 710 1249 712 1257
rect 728 1249 730 1257
rect 778 1256 780 1264
rect 783 1256 785 1264
rect 806 1262 808 1270
rect 1511 1249 1513 1257
rect 1527 1249 1529 1257
rect 1543 1249 1545 1257
rect 1566 1249 1568 1257
rect 1571 1249 1573 1257
rect 1597 1249 1599 1257
rect 1618 1249 1620 1257
rect 1638 1249 1640 1257
rect 1643 1249 1645 1257
rect 1661 1249 1663 1257
rect 1711 1256 1713 1264
rect 1716 1256 1718 1264
rect 1739 1262 1741 1270
rect 101 1194 103 1202
rect 106 1194 108 1202
rect 122 1194 124 1202
rect 138 1194 140 1202
rect 143 1194 145 1202
rect 164 1194 166 1202
rect 180 1194 182 1202
rect 196 1194 198 1202
rect 201 1194 203 1202
rect 217 1194 219 1202
rect 233 1194 235 1202
rect 238 1194 240 1202
rect 254 1194 256 1202
rect 270 1194 272 1202
rect 275 1194 277 1202
rect 296 1194 298 1202
rect 312 1194 314 1202
rect 328 1194 330 1202
rect 333 1194 335 1202
rect 349 1194 351 1202
rect 365 1194 367 1202
rect 370 1194 372 1202
rect 386 1194 388 1202
rect 402 1194 404 1202
rect 407 1194 409 1202
rect 428 1194 430 1202
rect 444 1194 446 1202
rect 460 1194 462 1202
rect 465 1194 467 1202
rect 481 1194 483 1202
rect 1034 1194 1036 1202
rect 1039 1194 1041 1202
rect 1055 1194 1057 1202
rect 1071 1194 1073 1202
rect 1076 1194 1078 1202
rect 1097 1194 1099 1202
rect 1113 1194 1115 1202
rect 1129 1194 1131 1202
rect 1134 1194 1136 1202
rect 1150 1194 1152 1202
rect 1166 1194 1168 1202
rect 1171 1194 1173 1202
rect 1187 1194 1189 1202
rect 1203 1194 1205 1202
rect 1208 1194 1210 1202
rect 1229 1194 1231 1202
rect 1245 1194 1247 1202
rect 1261 1194 1263 1202
rect 1266 1194 1268 1202
rect 1282 1194 1284 1202
rect 1298 1194 1300 1202
rect 1303 1194 1305 1202
rect 1319 1194 1321 1202
rect 1335 1194 1337 1202
rect 1340 1194 1342 1202
rect 1361 1194 1363 1202
rect 1377 1194 1379 1202
rect 1393 1194 1395 1202
rect 1398 1194 1400 1202
rect 1414 1194 1416 1202
rect 578 1163 580 1171
rect 594 1163 596 1171
rect 610 1163 612 1171
rect 633 1163 635 1171
rect 638 1163 640 1171
rect 664 1163 666 1171
rect 685 1163 687 1171
rect 705 1163 707 1171
rect 710 1163 712 1171
rect 728 1163 730 1171
rect 778 1158 780 1166
rect 783 1158 785 1166
rect 812 1163 814 1171
rect 830 1163 832 1171
rect 855 1163 857 1171
rect 871 1163 873 1171
rect 894 1163 896 1171
rect 899 1163 901 1171
rect 925 1163 927 1171
rect 946 1163 948 1171
rect 966 1163 968 1171
rect 971 1163 973 1171
rect 989 1163 991 1171
rect 1511 1163 1513 1171
rect 1527 1163 1529 1171
rect 1543 1163 1545 1171
rect 1566 1163 1568 1171
rect 1571 1163 1573 1171
rect 1597 1163 1599 1171
rect 1618 1163 1620 1171
rect 1638 1163 1640 1171
rect 1643 1163 1645 1171
rect 1661 1163 1663 1171
rect 1711 1158 1713 1166
rect 1716 1158 1718 1166
rect 1745 1163 1747 1171
rect 1763 1163 1765 1171
rect 1788 1163 1790 1171
rect 1804 1163 1806 1171
rect 1827 1163 1829 1171
rect 1832 1163 1834 1171
rect 1858 1163 1860 1171
rect 1879 1163 1881 1171
rect 1899 1163 1901 1171
rect 1904 1163 1906 1171
rect 1922 1163 1924 1171
rect 872 1084 874 1092
rect 877 1084 879 1092
rect 893 1084 895 1092
rect 909 1084 911 1092
rect 914 1084 916 1092
rect 935 1084 937 1092
rect 951 1084 953 1092
rect 967 1084 969 1092
rect 972 1084 974 1092
rect 988 1084 990 1092
rect 1805 1084 1807 1092
rect 1810 1084 1812 1092
rect 1826 1084 1828 1092
rect 1842 1084 1844 1092
rect 1847 1084 1849 1092
rect 1868 1084 1870 1092
rect 1884 1084 1886 1092
rect 1900 1084 1902 1092
rect 1905 1084 1907 1092
rect 1921 1084 1923 1092
rect 101 1054 103 1062
rect 106 1054 108 1062
rect 122 1054 124 1062
rect 138 1054 140 1062
rect 143 1054 145 1062
rect 164 1054 166 1062
rect 180 1054 182 1062
rect 196 1054 198 1062
rect 201 1054 203 1062
rect 217 1054 219 1062
rect 233 1054 235 1062
rect 238 1054 240 1062
rect 254 1054 256 1062
rect 270 1054 272 1062
rect 275 1054 277 1062
rect 296 1054 298 1062
rect 312 1054 314 1062
rect 328 1054 330 1062
rect 333 1054 335 1062
rect 349 1054 351 1062
rect 365 1054 367 1062
rect 370 1054 372 1062
rect 386 1054 388 1062
rect 402 1054 404 1062
rect 407 1054 409 1062
rect 428 1054 430 1062
rect 444 1054 446 1062
rect 460 1054 462 1062
rect 465 1054 467 1062
rect 481 1054 483 1062
rect 1034 1054 1036 1062
rect 1039 1054 1041 1062
rect 1055 1054 1057 1062
rect 1071 1054 1073 1062
rect 1076 1054 1078 1062
rect 1097 1054 1099 1062
rect 1113 1054 1115 1062
rect 1129 1054 1131 1062
rect 1134 1054 1136 1062
rect 1150 1054 1152 1062
rect 1166 1054 1168 1062
rect 1171 1054 1173 1062
rect 1187 1054 1189 1062
rect 1203 1054 1205 1062
rect 1208 1054 1210 1062
rect 1229 1054 1231 1062
rect 1245 1054 1247 1062
rect 1261 1054 1263 1062
rect 1266 1054 1268 1062
rect 1282 1054 1284 1062
rect 1298 1054 1300 1062
rect 1303 1054 1305 1062
rect 1319 1054 1321 1062
rect 1335 1054 1337 1062
rect 1340 1054 1342 1062
rect 1361 1054 1363 1062
rect 1377 1054 1379 1062
rect 1393 1054 1395 1062
rect 1398 1054 1400 1062
rect 1414 1054 1416 1062
rect 872 998 874 1006
rect 877 998 879 1006
rect 893 998 895 1006
rect 909 998 911 1006
rect 914 998 916 1006
rect 935 998 937 1006
rect 951 998 953 1006
rect 967 998 969 1006
rect 972 998 974 1006
rect 988 998 990 1006
rect 1805 998 1807 1006
rect 1810 998 1812 1006
rect 1826 998 1828 1006
rect 1842 998 1844 1006
rect 1847 998 1849 1006
rect 1868 998 1870 1006
rect 1884 998 1886 1006
rect 1900 998 1902 1006
rect 1905 998 1907 1006
rect 1921 998 1923 1006
rect 101 968 103 976
rect 106 968 108 976
rect 122 968 124 976
rect 138 968 140 976
rect 143 968 145 976
rect 164 968 166 976
rect 180 968 182 976
rect 196 968 198 976
rect 201 968 203 976
rect 217 968 219 976
rect 233 968 235 976
rect 238 968 240 976
rect 254 968 256 976
rect 270 968 272 976
rect 275 968 277 976
rect 296 968 298 976
rect 312 968 314 976
rect 328 968 330 976
rect 333 968 335 976
rect 349 968 351 976
rect 365 968 367 976
rect 370 968 372 976
rect 386 968 388 976
rect 402 968 404 976
rect 407 968 409 976
rect 428 968 430 976
rect 444 968 446 976
rect 460 968 462 976
rect 465 968 467 976
rect 481 968 483 976
rect 1034 968 1036 976
rect 1039 968 1041 976
rect 1055 968 1057 976
rect 1071 968 1073 976
rect 1076 968 1078 976
rect 1097 968 1099 976
rect 1113 968 1115 976
rect 1129 968 1131 976
rect 1134 968 1136 976
rect 1150 968 1152 976
rect 1166 968 1168 976
rect 1171 968 1173 976
rect 1187 968 1189 976
rect 1203 968 1205 976
rect 1208 968 1210 976
rect 1229 968 1231 976
rect 1245 968 1247 976
rect 1261 968 1263 976
rect 1266 968 1268 976
rect 1282 968 1284 976
rect 1298 968 1300 976
rect 1303 968 1305 976
rect 1319 968 1321 976
rect 1335 968 1337 976
rect 1340 968 1342 976
rect 1361 968 1363 976
rect 1377 968 1379 976
rect 1393 968 1395 976
rect 1398 968 1400 976
rect 1414 968 1416 976
rect 101 828 103 836
rect 106 828 108 836
rect 122 828 124 836
rect 138 828 140 836
rect 143 828 145 836
rect 164 828 166 836
rect 180 828 182 836
rect 196 828 198 836
rect 201 828 203 836
rect 217 828 219 836
rect 233 828 235 836
rect 238 828 240 836
rect 254 828 256 836
rect 270 828 272 836
rect 275 828 277 836
rect 296 828 298 836
rect 312 828 314 836
rect 328 828 330 836
rect 333 828 335 836
rect 349 828 351 836
rect 365 828 367 836
rect 370 828 372 836
rect 386 828 388 836
rect 402 828 404 836
rect 407 828 409 836
rect 428 828 430 836
rect 444 828 446 836
rect 460 828 462 836
rect 465 828 467 836
rect 481 828 483 836
rect 1034 828 1036 836
rect 1039 828 1041 836
rect 1055 828 1057 836
rect 1071 828 1073 836
rect 1076 828 1078 836
rect 1097 828 1099 836
rect 1113 828 1115 836
rect 1129 828 1131 836
rect 1134 828 1136 836
rect 1150 828 1152 836
rect 1166 828 1168 836
rect 1171 828 1173 836
rect 1187 828 1189 836
rect 1203 828 1205 836
rect 1208 828 1210 836
rect 1229 828 1231 836
rect 1245 828 1247 836
rect 1261 828 1263 836
rect 1266 828 1268 836
rect 1282 828 1284 836
rect 1298 828 1300 836
rect 1303 828 1305 836
rect 1319 828 1321 836
rect 1335 828 1337 836
rect 1340 828 1342 836
rect 1361 828 1363 836
rect 1377 828 1379 836
rect 1393 828 1395 836
rect 1398 828 1400 836
rect 1414 828 1416 836
rect 573 749 575 757
rect 578 749 580 757
rect 594 749 596 757
rect 610 749 612 757
rect 615 749 617 757
rect 636 749 638 757
rect 652 749 654 757
rect 668 749 670 757
rect 673 749 675 757
rect 689 749 691 757
rect 705 749 707 757
rect 710 749 712 757
rect 726 749 728 757
rect 742 749 744 757
rect 747 749 749 757
rect 768 749 770 757
rect 784 749 786 757
rect 800 749 802 757
rect 805 749 807 757
rect 821 749 823 757
rect 837 749 839 757
rect 842 749 844 757
rect 858 749 860 757
rect 874 749 876 757
rect 879 749 881 757
rect 900 749 902 757
rect 916 749 918 757
rect 932 749 934 757
rect 937 749 939 757
rect 953 749 955 757
rect 969 749 971 757
rect 974 749 976 757
rect 990 749 992 757
rect 1006 749 1008 757
rect 1011 749 1013 757
rect 1032 749 1034 757
rect 1048 749 1050 757
rect 1064 749 1066 757
rect 1069 749 1071 757
rect 1085 749 1087 757
rect 1506 749 1508 757
rect 1511 749 1513 757
rect 1527 749 1529 757
rect 1543 749 1545 757
rect 1548 749 1550 757
rect 1569 749 1571 757
rect 1585 749 1587 757
rect 1601 749 1603 757
rect 1606 749 1608 757
rect 1622 749 1624 757
rect 1638 749 1640 757
rect 1643 749 1645 757
rect 1659 749 1661 757
rect 1675 749 1677 757
rect 1680 749 1682 757
rect 1701 749 1703 757
rect 1717 749 1719 757
rect 1733 749 1735 757
rect 1738 749 1740 757
rect 1754 749 1756 757
rect 1770 749 1772 757
rect 1775 749 1777 757
rect 1791 749 1793 757
rect 1807 749 1809 757
rect 1812 749 1814 757
rect 1833 749 1835 757
rect 1849 749 1851 757
rect 1865 749 1867 757
rect 1870 749 1872 757
rect 1886 749 1888 757
rect 1902 749 1904 757
rect 1907 749 1909 757
rect 1923 749 1925 757
rect 1939 749 1941 757
rect 1944 749 1946 757
rect 1965 749 1967 757
rect 1981 749 1983 757
rect 1997 749 1999 757
rect 2002 749 2004 757
rect 2018 749 2020 757
rect 233 716 235 724
rect 238 716 240 724
rect 254 716 256 724
rect 270 716 272 724
rect 275 716 277 724
rect 296 716 298 724
rect 312 716 314 724
rect 328 716 330 724
rect 333 716 335 724
rect 349 716 351 724
rect 1166 716 1168 724
rect 1171 716 1173 724
rect 1187 716 1189 724
rect 1203 716 1205 724
rect 1208 716 1210 724
rect 1229 716 1231 724
rect 1245 716 1247 724
rect 1261 716 1263 724
rect 1266 716 1268 724
rect 1282 716 1284 724
rect 752 678 754 686
rect 578 665 580 673
rect 594 665 596 673
rect 610 665 612 673
rect 633 665 635 673
rect 638 665 640 673
rect 664 665 666 673
rect 685 665 687 673
rect 705 665 707 673
rect 710 665 712 673
rect 728 665 730 673
rect 778 672 780 680
rect 783 672 785 680
rect 806 678 808 686
rect 833 678 835 686
rect 859 672 861 680
rect 864 672 866 680
rect 887 678 889 686
rect 1685 678 1687 686
rect 1511 665 1513 673
rect 1527 665 1529 673
rect 1543 665 1545 673
rect 1566 665 1568 673
rect 1571 665 1573 673
rect 1597 665 1599 673
rect 1618 665 1620 673
rect 1638 665 1640 673
rect 1643 665 1645 673
rect 1661 665 1663 673
rect 1711 672 1713 680
rect 1716 672 1718 680
rect 1739 678 1741 686
rect 1766 678 1768 686
rect 1792 672 1794 680
rect 1797 672 1799 680
rect 1820 678 1822 686
rect 224 614 226 622
rect 240 614 242 622
rect 245 614 247 622
rect 261 614 263 622
rect 277 614 279 622
rect 298 614 300 622
rect 303 614 305 622
rect 319 614 321 622
rect 335 614 337 622
rect 340 614 342 622
rect 1157 614 1159 622
rect 1173 614 1175 622
rect 1178 614 1180 622
rect 1194 614 1196 622
rect 1210 614 1212 622
rect 1231 614 1233 622
rect 1236 614 1238 622
rect 1252 614 1254 622
rect 1268 614 1270 622
rect 1273 614 1275 622
rect 578 579 580 587
rect 594 579 596 587
rect 610 579 612 587
rect 633 579 635 587
rect 638 579 640 587
rect 664 579 666 587
rect 685 579 687 587
rect 705 579 707 587
rect 710 579 712 587
rect 728 579 730 587
rect 778 580 780 588
rect 783 580 785 588
rect 859 580 861 588
rect 864 580 866 588
rect 1511 579 1513 587
rect 1527 579 1529 587
rect 1543 579 1545 587
rect 1566 579 1568 587
rect 1571 579 1573 587
rect 1597 579 1599 587
rect 1618 579 1620 587
rect 1638 579 1640 587
rect 1643 579 1645 587
rect 1661 579 1663 587
rect 1711 580 1713 588
rect 1716 580 1718 588
rect 1792 580 1794 588
rect 1797 580 1799 588
rect 578 533 580 541
rect 594 533 596 541
rect 610 533 612 541
rect 633 533 635 541
rect 638 533 640 541
rect 664 533 666 541
rect 685 533 687 541
rect 705 533 707 541
rect 710 533 712 541
rect 728 533 730 541
rect 778 540 780 548
rect 783 540 785 548
rect 806 546 808 554
rect 857 546 859 554
rect 883 540 885 548
rect 888 540 890 548
rect 911 546 913 554
rect 1511 533 1513 541
rect 1527 533 1529 541
rect 1543 533 1545 541
rect 1566 533 1568 541
rect 1571 533 1573 541
rect 1597 533 1599 541
rect 1618 533 1620 541
rect 1638 533 1640 541
rect 1643 533 1645 541
rect 1661 533 1663 541
rect 1711 540 1713 548
rect 1716 540 1718 548
rect 1739 546 1741 554
rect 1790 546 1792 554
rect 1816 540 1818 548
rect 1821 540 1823 548
rect 1844 546 1846 554
rect 578 447 580 455
rect 594 447 596 455
rect 610 447 612 455
rect 633 447 635 455
rect 638 447 640 455
rect 664 447 666 455
rect 685 447 687 455
rect 705 447 707 455
rect 710 447 712 455
rect 728 447 730 455
rect 778 449 780 457
rect 783 449 785 457
rect 883 449 885 457
rect 888 449 890 457
rect 1511 447 1513 455
rect 1527 447 1529 455
rect 1543 447 1545 455
rect 1566 447 1568 455
rect 1571 447 1573 455
rect 1597 447 1599 455
rect 1618 447 1620 455
rect 1638 447 1640 455
rect 1643 447 1645 455
rect 1661 447 1663 455
rect 1711 449 1713 457
rect 1716 449 1718 457
rect 1816 449 1818 457
rect 1821 449 1823 457
rect 578 401 580 409
rect 594 401 596 409
rect 610 401 612 409
rect 633 401 635 409
rect 638 401 640 409
rect 664 401 666 409
rect 685 401 687 409
rect 705 401 707 409
rect 710 401 712 409
rect 728 401 730 409
rect 778 408 780 416
rect 783 408 785 416
rect 806 414 808 422
rect 833 414 835 422
rect 859 408 861 416
rect 864 408 866 416
rect 887 414 889 422
rect 923 414 925 422
rect 949 408 951 416
rect 954 408 956 416
rect 977 414 979 422
rect 1511 401 1513 409
rect 1527 401 1529 409
rect 1543 401 1545 409
rect 1566 401 1568 409
rect 1571 401 1573 409
rect 1597 401 1599 409
rect 1618 401 1620 409
rect 1638 401 1640 409
rect 1643 401 1645 409
rect 1661 401 1663 409
rect 1711 408 1713 416
rect 1716 408 1718 416
rect 1739 414 1741 422
rect 1766 414 1768 422
rect 1792 408 1794 416
rect 1797 408 1799 416
rect 1820 414 1822 422
rect 1856 414 1858 422
rect 1882 408 1884 416
rect 1887 408 1889 416
rect 1910 414 1912 422
rect 578 315 580 323
rect 594 315 596 323
rect 610 315 612 323
rect 633 315 635 323
rect 638 315 640 323
rect 664 315 666 323
rect 685 315 687 323
rect 705 315 707 323
rect 710 315 712 323
rect 728 315 730 323
rect 778 314 780 322
rect 783 314 785 322
rect 859 314 861 322
rect 864 314 866 322
rect 949 314 951 322
rect 954 314 956 322
rect 1511 315 1513 323
rect 1527 315 1529 323
rect 1543 315 1545 323
rect 1566 315 1568 323
rect 1571 315 1573 323
rect 1597 315 1599 323
rect 1618 315 1620 323
rect 1638 315 1640 323
rect 1643 315 1645 323
rect 1661 315 1663 323
rect 1711 314 1713 322
rect 1716 314 1718 322
rect 1792 314 1794 322
rect 1797 314 1799 322
rect 1882 314 1884 322
rect 1887 314 1889 322
rect 578 269 580 277
rect 594 269 596 277
rect 610 269 612 277
rect 633 269 635 277
rect 638 269 640 277
rect 664 269 666 277
rect 685 269 687 277
rect 705 269 707 277
rect 710 269 712 277
rect 728 269 730 277
rect 778 276 780 284
rect 783 276 785 284
rect 806 282 808 290
rect 1511 269 1513 277
rect 1527 269 1529 277
rect 1543 269 1545 277
rect 1566 269 1568 277
rect 1571 269 1573 277
rect 1597 269 1599 277
rect 1618 269 1620 277
rect 1638 269 1640 277
rect 1643 269 1645 277
rect 1661 269 1663 277
rect 1711 276 1713 284
rect 1716 276 1718 284
rect 1739 282 1741 290
rect 101 214 103 222
rect 106 214 108 222
rect 122 214 124 222
rect 138 214 140 222
rect 143 214 145 222
rect 164 214 166 222
rect 180 214 182 222
rect 196 214 198 222
rect 201 214 203 222
rect 217 214 219 222
rect 233 214 235 222
rect 238 214 240 222
rect 254 214 256 222
rect 270 214 272 222
rect 275 214 277 222
rect 296 214 298 222
rect 312 214 314 222
rect 328 214 330 222
rect 333 214 335 222
rect 349 214 351 222
rect 365 214 367 222
rect 370 214 372 222
rect 386 214 388 222
rect 402 214 404 222
rect 407 214 409 222
rect 428 214 430 222
rect 444 214 446 222
rect 460 214 462 222
rect 465 214 467 222
rect 481 214 483 222
rect 1034 214 1036 222
rect 1039 214 1041 222
rect 1055 214 1057 222
rect 1071 214 1073 222
rect 1076 214 1078 222
rect 1097 214 1099 222
rect 1113 214 1115 222
rect 1129 214 1131 222
rect 1134 214 1136 222
rect 1150 214 1152 222
rect 1166 214 1168 222
rect 1171 214 1173 222
rect 1187 214 1189 222
rect 1203 214 1205 222
rect 1208 214 1210 222
rect 1229 214 1231 222
rect 1245 214 1247 222
rect 1261 214 1263 222
rect 1266 214 1268 222
rect 1282 214 1284 222
rect 1298 214 1300 222
rect 1303 214 1305 222
rect 1319 214 1321 222
rect 1335 214 1337 222
rect 1340 214 1342 222
rect 1361 214 1363 222
rect 1377 214 1379 222
rect 1393 214 1395 222
rect 1398 214 1400 222
rect 1414 214 1416 222
rect 578 183 580 191
rect 594 183 596 191
rect 610 183 612 191
rect 633 183 635 191
rect 638 183 640 191
rect 664 183 666 191
rect 685 183 687 191
rect 705 183 707 191
rect 710 183 712 191
rect 728 183 730 191
rect 778 178 780 186
rect 783 178 785 186
rect 812 183 814 191
rect 830 183 832 191
rect 855 183 857 191
rect 871 183 873 191
rect 894 183 896 191
rect 899 183 901 191
rect 925 183 927 191
rect 946 183 948 191
rect 966 183 968 191
rect 971 183 973 191
rect 989 183 991 191
rect 1511 183 1513 191
rect 1527 183 1529 191
rect 1543 183 1545 191
rect 1566 183 1568 191
rect 1571 183 1573 191
rect 1597 183 1599 191
rect 1618 183 1620 191
rect 1638 183 1640 191
rect 1643 183 1645 191
rect 1661 183 1663 191
rect 1711 178 1713 186
rect 1716 178 1718 186
rect 1745 183 1747 191
rect 1763 183 1765 191
rect 1788 183 1790 191
rect 1804 183 1806 191
rect 1827 183 1829 191
rect 1832 183 1834 191
rect 1858 183 1860 191
rect 1879 183 1881 191
rect 1899 183 1901 191
rect 1904 183 1906 191
rect 1922 183 1924 191
rect 872 104 874 112
rect 877 104 879 112
rect 893 104 895 112
rect 909 104 911 112
rect 914 104 916 112
rect 935 104 937 112
rect 951 104 953 112
rect 967 104 969 112
rect 972 104 974 112
rect 988 104 990 112
rect 1805 104 1807 112
rect 1810 104 1812 112
rect 1826 104 1828 112
rect 1842 104 1844 112
rect 1847 104 1849 112
rect 1868 104 1870 112
rect 1884 104 1886 112
rect 1900 104 1902 112
rect 1905 104 1907 112
rect 1921 104 1923 112
rect 101 74 103 82
rect 106 74 108 82
rect 122 74 124 82
rect 138 74 140 82
rect 143 74 145 82
rect 164 74 166 82
rect 180 74 182 82
rect 196 74 198 82
rect 201 74 203 82
rect 217 74 219 82
rect 233 74 235 82
rect 238 74 240 82
rect 254 74 256 82
rect 270 74 272 82
rect 275 74 277 82
rect 296 74 298 82
rect 312 74 314 82
rect 328 74 330 82
rect 333 74 335 82
rect 349 74 351 82
rect 365 74 367 82
rect 370 74 372 82
rect 386 74 388 82
rect 402 74 404 82
rect 407 74 409 82
rect 428 74 430 82
rect 444 74 446 82
rect 460 74 462 82
rect 465 74 467 82
rect 481 74 483 82
rect 1034 74 1036 82
rect 1039 74 1041 82
rect 1055 74 1057 82
rect 1071 74 1073 82
rect 1076 74 1078 82
rect 1097 74 1099 82
rect 1113 74 1115 82
rect 1129 74 1131 82
rect 1134 74 1136 82
rect 1150 74 1152 82
rect 1166 74 1168 82
rect 1171 74 1173 82
rect 1187 74 1189 82
rect 1203 74 1205 82
rect 1208 74 1210 82
rect 1229 74 1231 82
rect 1245 74 1247 82
rect 1261 74 1263 82
rect 1266 74 1268 82
rect 1282 74 1284 82
rect 1298 74 1300 82
rect 1303 74 1305 82
rect 1319 74 1321 82
rect 1335 74 1337 82
rect 1340 74 1342 82
rect 1361 74 1363 82
rect 1377 74 1379 82
rect 1393 74 1395 82
rect 1398 74 1400 82
rect 1414 74 1416 82
rect 872 18 874 26
rect 877 18 879 26
rect 893 18 895 26
rect 909 18 911 26
rect 914 18 916 26
rect 935 18 937 26
rect 951 18 953 26
rect 967 18 969 26
rect 972 18 974 26
rect 988 18 990 26
rect 1805 18 1807 26
rect 1810 18 1812 26
rect 1826 18 1828 26
rect 1842 18 1844 26
rect 1847 18 1849 26
rect 1868 18 1870 26
rect 1884 18 1886 26
rect 1900 18 1902 26
rect 1905 18 1907 26
rect 1921 18 1923 26
rect 101 -12 103 -4
rect 106 -12 108 -4
rect 122 -12 124 -4
rect 138 -12 140 -4
rect 143 -12 145 -4
rect 164 -12 166 -4
rect 180 -12 182 -4
rect 196 -12 198 -4
rect 201 -12 203 -4
rect 217 -12 219 -4
rect 233 -12 235 -4
rect 238 -12 240 -4
rect 254 -12 256 -4
rect 270 -12 272 -4
rect 275 -12 277 -4
rect 296 -12 298 -4
rect 312 -12 314 -4
rect 328 -12 330 -4
rect 333 -12 335 -4
rect 349 -12 351 -4
rect 365 -12 367 -4
rect 370 -12 372 -4
rect 386 -12 388 -4
rect 402 -12 404 -4
rect 407 -12 409 -4
rect 428 -12 430 -4
rect 444 -12 446 -4
rect 460 -12 462 -4
rect 465 -12 467 -4
rect 481 -12 483 -4
rect 1034 -12 1036 -4
rect 1039 -12 1041 -4
rect 1055 -12 1057 -4
rect 1071 -12 1073 -4
rect 1076 -12 1078 -4
rect 1097 -12 1099 -4
rect 1113 -12 1115 -4
rect 1129 -12 1131 -4
rect 1134 -12 1136 -4
rect 1150 -12 1152 -4
rect 1166 -12 1168 -4
rect 1171 -12 1173 -4
rect 1187 -12 1189 -4
rect 1203 -12 1205 -4
rect 1208 -12 1210 -4
rect 1229 -12 1231 -4
rect 1245 -12 1247 -4
rect 1261 -12 1263 -4
rect 1266 -12 1268 -4
rect 1282 -12 1284 -4
rect 1298 -12 1300 -4
rect 1303 -12 1305 -4
rect 1319 -12 1321 -4
rect 1335 -12 1337 -4
rect 1340 -12 1342 -4
rect 1361 -12 1363 -4
rect 1377 -12 1379 -4
rect 1393 -12 1395 -4
rect 1398 -12 1400 -4
rect 1414 -12 1416 -4
rect 101 -152 103 -144
rect 106 -152 108 -144
rect 122 -152 124 -144
rect 138 -152 140 -144
rect 143 -152 145 -144
rect 164 -152 166 -144
rect 180 -152 182 -144
rect 196 -152 198 -144
rect 201 -152 203 -144
rect 217 -152 219 -144
rect 233 -152 235 -144
rect 238 -152 240 -144
rect 254 -152 256 -144
rect 270 -152 272 -144
rect 275 -152 277 -144
rect 296 -152 298 -144
rect 312 -152 314 -144
rect 328 -152 330 -144
rect 333 -152 335 -144
rect 349 -152 351 -144
rect 365 -152 367 -144
rect 370 -152 372 -144
rect 386 -152 388 -144
rect 402 -152 404 -144
rect 407 -152 409 -144
rect 428 -152 430 -144
rect 444 -152 446 -144
rect 460 -152 462 -144
rect 465 -152 467 -144
rect 481 -152 483 -144
rect 1034 -152 1036 -144
rect 1039 -152 1041 -144
rect 1055 -152 1057 -144
rect 1071 -152 1073 -144
rect 1076 -152 1078 -144
rect 1097 -152 1099 -144
rect 1113 -152 1115 -144
rect 1129 -152 1131 -144
rect 1134 -152 1136 -144
rect 1150 -152 1152 -144
rect 1166 -152 1168 -144
rect 1171 -152 1173 -144
rect 1187 -152 1189 -144
rect 1203 -152 1205 -144
rect 1208 -152 1210 -144
rect 1229 -152 1231 -144
rect 1245 -152 1247 -144
rect 1261 -152 1263 -144
rect 1266 -152 1268 -144
rect 1282 -152 1284 -144
rect 1298 -152 1300 -144
rect 1303 -152 1305 -144
rect 1319 -152 1321 -144
rect 1335 -152 1337 -144
rect 1340 -152 1342 -144
rect 1361 -152 1363 -144
rect 1377 -152 1379 -144
rect 1393 -152 1395 -144
rect 1398 -152 1400 -144
rect 1414 -152 1416 -144
<< ndiffusion >>
rect 572 1706 573 1710
rect 575 1706 578 1710
rect 580 1706 581 1710
rect 593 1706 594 1710
rect 596 1706 597 1710
rect 609 1706 610 1710
rect 612 1706 615 1710
rect 617 1706 618 1710
rect 635 1706 636 1710
rect 638 1706 639 1710
rect 651 1706 652 1710
rect 654 1706 655 1710
rect 667 1706 668 1710
rect 670 1706 673 1710
rect 675 1706 676 1710
rect 688 1706 689 1710
rect 691 1706 692 1710
rect 704 1706 705 1710
rect 707 1706 710 1710
rect 712 1706 713 1710
rect 725 1706 726 1710
rect 728 1706 729 1710
rect 741 1706 742 1710
rect 744 1706 747 1710
rect 749 1706 750 1710
rect 767 1706 768 1710
rect 770 1706 771 1710
rect 783 1706 784 1710
rect 786 1706 787 1710
rect 799 1706 800 1710
rect 802 1706 805 1710
rect 807 1706 808 1710
rect 820 1706 821 1710
rect 823 1706 824 1710
rect 836 1706 837 1710
rect 839 1706 842 1710
rect 844 1706 845 1710
rect 857 1706 858 1710
rect 860 1706 861 1710
rect 873 1706 874 1710
rect 876 1706 879 1710
rect 881 1706 882 1710
rect 899 1706 900 1710
rect 902 1706 903 1710
rect 915 1706 916 1710
rect 918 1706 919 1710
rect 931 1706 932 1710
rect 934 1706 937 1710
rect 939 1706 940 1710
rect 952 1706 953 1710
rect 955 1706 956 1710
rect 968 1706 969 1710
rect 971 1706 974 1710
rect 976 1706 977 1710
rect 989 1706 990 1710
rect 992 1706 993 1710
rect 1005 1706 1006 1710
rect 1008 1706 1011 1710
rect 1013 1706 1014 1710
rect 1031 1706 1032 1710
rect 1034 1706 1035 1710
rect 1047 1706 1048 1710
rect 1050 1706 1051 1710
rect 1063 1706 1064 1710
rect 1066 1706 1069 1710
rect 1071 1706 1072 1710
rect 1084 1706 1085 1710
rect 1087 1706 1088 1710
rect 1505 1706 1506 1710
rect 1508 1706 1511 1710
rect 1513 1706 1514 1710
rect 1526 1706 1527 1710
rect 1529 1706 1530 1710
rect 1542 1706 1543 1710
rect 1545 1706 1548 1710
rect 1550 1706 1551 1710
rect 1568 1706 1569 1710
rect 1571 1706 1572 1710
rect 1584 1706 1585 1710
rect 1587 1706 1588 1710
rect 1600 1706 1601 1710
rect 1603 1706 1606 1710
rect 1608 1706 1609 1710
rect 1621 1706 1622 1710
rect 1624 1706 1625 1710
rect 1637 1706 1638 1710
rect 1640 1706 1643 1710
rect 1645 1706 1646 1710
rect 1658 1706 1659 1710
rect 1661 1706 1662 1710
rect 1674 1706 1675 1710
rect 1677 1706 1680 1710
rect 1682 1706 1683 1710
rect 1700 1706 1701 1710
rect 1703 1706 1704 1710
rect 1716 1706 1717 1710
rect 1719 1706 1720 1710
rect 1732 1706 1733 1710
rect 1735 1706 1738 1710
rect 1740 1706 1741 1710
rect 1753 1706 1754 1710
rect 1756 1706 1757 1710
rect 1769 1706 1770 1710
rect 1772 1706 1775 1710
rect 1777 1706 1778 1710
rect 1790 1706 1791 1710
rect 1793 1706 1794 1710
rect 1806 1706 1807 1710
rect 1809 1706 1812 1710
rect 1814 1706 1815 1710
rect 1832 1706 1833 1710
rect 1835 1706 1836 1710
rect 1848 1706 1849 1710
rect 1851 1706 1852 1710
rect 1864 1706 1865 1710
rect 1867 1706 1870 1710
rect 1872 1706 1873 1710
rect 1885 1706 1886 1710
rect 1888 1706 1889 1710
rect 1901 1706 1902 1710
rect 1904 1706 1907 1710
rect 1909 1706 1910 1710
rect 1922 1706 1923 1710
rect 1925 1706 1926 1710
rect 1938 1706 1939 1710
rect 1941 1706 1944 1710
rect 1946 1706 1947 1710
rect 1964 1706 1965 1710
rect 1967 1706 1968 1710
rect 1980 1706 1981 1710
rect 1983 1706 1984 1710
rect 1996 1706 1997 1710
rect 1999 1706 2002 1710
rect 2004 1706 2005 1710
rect 2017 1706 2018 1710
rect 2020 1706 2021 1710
rect 232 1673 233 1677
rect 235 1673 238 1677
rect 240 1673 241 1677
rect 253 1673 254 1677
rect 256 1673 257 1677
rect 269 1673 270 1677
rect 272 1673 275 1677
rect 277 1673 278 1677
rect 295 1673 296 1677
rect 298 1673 299 1677
rect 311 1673 312 1677
rect 314 1673 315 1677
rect 327 1673 328 1677
rect 330 1673 333 1677
rect 335 1673 336 1677
rect 348 1673 349 1677
rect 351 1673 352 1677
rect 1165 1673 1166 1677
rect 1168 1673 1171 1677
rect 1173 1673 1174 1677
rect 1186 1673 1187 1677
rect 1189 1673 1190 1677
rect 1202 1673 1203 1677
rect 1205 1673 1208 1677
rect 1210 1673 1211 1677
rect 1228 1673 1229 1677
rect 1231 1673 1232 1677
rect 1244 1673 1245 1677
rect 1247 1673 1248 1677
rect 1260 1673 1261 1677
rect 1263 1673 1266 1677
rect 1268 1673 1269 1677
rect 1281 1673 1282 1677
rect 1284 1673 1285 1677
rect 356 1636 357 1640
rect 359 1636 360 1640
rect 751 1640 752 1644
rect 754 1640 755 1644
rect 775 1636 778 1640
rect 780 1636 783 1640
rect 785 1636 786 1640
rect 832 1640 833 1644
rect 835 1640 836 1644
rect 856 1636 859 1640
rect 861 1636 864 1640
rect 866 1636 867 1640
rect 805 1632 806 1636
rect 808 1632 809 1636
rect 239 1627 240 1631
rect 242 1627 243 1631
rect 577 1627 578 1631
rect 580 1627 581 1631
rect 593 1627 594 1631
rect 596 1627 597 1631
rect 609 1627 610 1631
rect 612 1627 613 1631
rect 628 1627 633 1631
rect 635 1627 638 1631
rect 640 1627 641 1631
rect 662 1627 664 1631
rect 666 1627 667 1631
rect 684 1627 685 1631
rect 687 1627 688 1631
rect 700 1627 705 1631
rect 707 1627 710 1631
rect 712 1627 713 1631
rect 727 1627 728 1631
rect 730 1627 731 1631
rect 886 1632 887 1636
rect 889 1632 890 1636
rect 1289 1636 1290 1640
rect 1292 1636 1293 1640
rect 1684 1640 1685 1644
rect 1687 1640 1688 1644
rect 1708 1636 1711 1640
rect 1713 1636 1716 1640
rect 1718 1636 1719 1640
rect 1765 1640 1766 1644
rect 1768 1640 1769 1644
rect 1789 1636 1792 1640
rect 1794 1636 1797 1640
rect 1799 1636 1800 1640
rect 1738 1632 1739 1636
rect 1741 1632 1742 1636
rect 1172 1627 1173 1631
rect 1175 1627 1176 1631
rect 1510 1627 1511 1631
rect 1513 1627 1514 1631
rect 1526 1627 1527 1631
rect 1529 1627 1530 1631
rect 1542 1627 1543 1631
rect 1545 1627 1546 1631
rect 1561 1627 1566 1631
rect 1568 1627 1571 1631
rect 1573 1627 1574 1631
rect 1595 1627 1597 1631
rect 1599 1627 1600 1631
rect 1617 1627 1618 1631
rect 1620 1627 1621 1631
rect 1633 1627 1638 1631
rect 1640 1627 1643 1631
rect 1645 1627 1646 1631
rect 1660 1627 1661 1631
rect 1663 1627 1664 1631
rect 1819 1632 1820 1636
rect 1822 1632 1823 1636
rect 577 1581 578 1585
rect 580 1581 581 1585
rect 593 1581 594 1585
rect 596 1581 597 1585
rect 609 1581 610 1585
rect 612 1581 613 1585
rect 628 1581 633 1585
rect 635 1581 638 1585
rect 640 1581 641 1585
rect 662 1581 664 1585
rect 666 1581 667 1585
rect 684 1581 685 1585
rect 687 1581 688 1585
rect 700 1581 705 1585
rect 707 1581 710 1585
rect 712 1581 713 1585
rect 727 1581 728 1585
rect 730 1581 731 1585
rect 223 1571 224 1575
rect 226 1571 227 1575
rect 239 1571 240 1575
rect 242 1571 245 1575
rect 247 1571 248 1575
rect 260 1571 261 1575
rect 263 1571 264 1575
rect 276 1571 277 1575
rect 279 1571 280 1575
rect 297 1571 298 1575
rect 300 1571 303 1575
rect 305 1571 306 1575
rect 318 1571 319 1575
rect 321 1571 322 1575
rect 334 1571 335 1575
rect 337 1571 340 1575
rect 342 1571 343 1575
rect 775 1580 778 1584
rect 780 1580 783 1584
rect 785 1580 786 1584
rect 856 1580 859 1584
rect 861 1580 864 1584
rect 866 1580 867 1584
rect 1510 1581 1511 1585
rect 1513 1581 1514 1585
rect 1526 1581 1527 1585
rect 1529 1581 1530 1585
rect 1542 1581 1543 1585
rect 1545 1581 1546 1585
rect 1561 1581 1566 1585
rect 1568 1581 1571 1585
rect 1573 1581 1574 1585
rect 1595 1581 1597 1585
rect 1599 1581 1600 1585
rect 1617 1581 1618 1585
rect 1620 1581 1621 1585
rect 1633 1581 1638 1585
rect 1640 1581 1643 1585
rect 1645 1581 1646 1585
rect 1660 1581 1661 1585
rect 1663 1581 1664 1585
rect 1156 1571 1157 1575
rect 1159 1571 1160 1575
rect 1172 1571 1173 1575
rect 1175 1571 1178 1575
rect 1180 1571 1181 1575
rect 1193 1571 1194 1575
rect 1196 1571 1197 1575
rect 1209 1571 1210 1575
rect 1212 1571 1213 1575
rect 1230 1571 1231 1575
rect 1233 1571 1236 1575
rect 1238 1571 1239 1575
rect 1251 1571 1252 1575
rect 1254 1571 1255 1575
rect 1267 1571 1268 1575
rect 1270 1571 1273 1575
rect 1275 1571 1276 1575
rect 1708 1580 1711 1584
rect 1713 1580 1716 1584
rect 1718 1580 1719 1584
rect 1789 1580 1792 1584
rect 1794 1580 1797 1584
rect 1799 1580 1800 1584
rect 775 1504 778 1508
rect 780 1504 783 1508
rect 785 1504 786 1508
rect 856 1508 857 1512
rect 859 1508 860 1512
rect 880 1504 883 1508
rect 885 1504 888 1508
rect 890 1504 891 1508
rect 805 1500 806 1504
rect 808 1500 809 1504
rect 577 1495 578 1499
rect 580 1495 581 1499
rect 593 1495 594 1499
rect 596 1495 597 1499
rect 609 1495 610 1499
rect 612 1495 613 1499
rect 628 1495 633 1499
rect 635 1495 638 1499
rect 640 1495 641 1499
rect 662 1495 664 1499
rect 666 1495 667 1499
rect 684 1495 685 1499
rect 687 1495 688 1499
rect 700 1495 705 1499
rect 707 1495 710 1499
rect 712 1495 713 1499
rect 727 1495 728 1499
rect 730 1495 731 1499
rect 910 1500 911 1504
rect 913 1500 914 1504
rect 1708 1504 1711 1508
rect 1713 1504 1716 1508
rect 1718 1504 1719 1508
rect 1789 1508 1790 1512
rect 1792 1508 1793 1512
rect 1813 1504 1816 1508
rect 1818 1504 1821 1508
rect 1823 1504 1824 1508
rect 1738 1500 1739 1504
rect 1741 1500 1742 1504
rect 1510 1495 1511 1499
rect 1513 1495 1514 1499
rect 1526 1495 1527 1499
rect 1529 1495 1530 1499
rect 1542 1495 1543 1499
rect 1545 1495 1546 1499
rect 1561 1495 1566 1499
rect 1568 1495 1571 1499
rect 1573 1495 1574 1499
rect 1595 1495 1597 1499
rect 1599 1495 1600 1499
rect 1617 1495 1618 1499
rect 1620 1495 1621 1499
rect 1633 1495 1638 1499
rect 1640 1495 1643 1499
rect 1645 1495 1646 1499
rect 1660 1495 1661 1499
rect 1663 1495 1664 1499
rect 1843 1500 1844 1504
rect 1846 1500 1847 1504
rect 577 1449 578 1453
rect 580 1449 581 1453
rect 593 1449 594 1453
rect 596 1449 597 1453
rect 609 1449 610 1453
rect 612 1449 613 1453
rect 628 1449 633 1453
rect 635 1449 638 1453
rect 640 1449 641 1453
rect 662 1449 664 1453
rect 666 1449 667 1453
rect 684 1449 685 1453
rect 687 1449 688 1453
rect 700 1449 705 1453
rect 707 1449 710 1453
rect 712 1449 713 1453
rect 727 1449 728 1453
rect 730 1449 731 1453
rect 775 1449 778 1453
rect 780 1449 783 1453
rect 785 1449 786 1453
rect 880 1449 883 1453
rect 885 1449 888 1453
rect 890 1449 891 1453
rect 1510 1449 1511 1453
rect 1513 1449 1514 1453
rect 1526 1449 1527 1453
rect 1529 1449 1530 1453
rect 1542 1449 1543 1453
rect 1545 1449 1546 1453
rect 1561 1449 1566 1453
rect 1568 1449 1571 1453
rect 1573 1449 1574 1453
rect 1595 1449 1597 1453
rect 1599 1449 1600 1453
rect 1617 1449 1618 1453
rect 1620 1449 1621 1453
rect 1633 1449 1638 1453
rect 1640 1449 1643 1453
rect 1645 1449 1646 1453
rect 1660 1449 1661 1453
rect 1663 1449 1664 1453
rect 1708 1449 1711 1453
rect 1713 1449 1716 1453
rect 1718 1449 1719 1453
rect 1813 1449 1816 1453
rect 1818 1449 1821 1453
rect 1823 1449 1824 1453
rect 775 1372 778 1376
rect 780 1372 783 1376
rect 785 1372 786 1376
rect 832 1376 833 1380
rect 835 1376 836 1380
rect 856 1372 859 1376
rect 861 1372 864 1376
rect 866 1372 867 1376
rect 922 1376 923 1380
rect 925 1376 926 1380
rect 946 1372 949 1376
rect 951 1372 954 1376
rect 956 1372 957 1376
rect 805 1368 806 1372
rect 808 1368 809 1372
rect 577 1363 578 1367
rect 580 1363 581 1367
rect 593 1363 594 1367
rect 596 1363 597 1367
rect 609 1363 610 1367
rect 612 1363 613 1367
rect 628 1363 633 1367
rect 635 1363 638 1367
rect 640 1363 641 1367
rect 662 1363 664 1367
rect 666 1363 667 1367
rect 684 1363 685 1367
rect 687 1363 688 1367
rect 700 1363 705 1367
rect 707 1363 710 1367
rect 712 1363 713 1367
rect 727 1363 728 1367
rect 730 1363 731 1367
rect 886 1368 887 1372
rect 889 1368 890 1372
rect 976 1368 977 1372
rect 979 1368 980 1372
rect 1708 1372 1711 1376
rect 1713 1372 1716 1376
rect 1718 1372 1719 1376
rect 1765 1376 1766 1380
rect 1768 1376 1769 1380
rect 1789 1372 1792 1376
rect 1794 1372 1797 1376
rect 1799 1372 1800 1376
rect 1855 1376 1856 1380
rect 1858 1376 1859 1380
rect 1879 1372 1882 1376
rect 1884 1372 1887 1376
rect 1889 1372 1890 1376
rect 1738 1368 1739 1372
rect 1741 1368 1742 1372
rect 1510 1363 1511 1367
rect 1513 1363 1514 1367
rect 1526 1363 1527 1367
rect 1529 1363 1530 1367
rect 1542 1363 1543 1367
rect 1545 1363 1546 1367
rect 1561 1363 1566 1367
rect 1568 1363 1571 1367
rect 1573 1363 1574 1367
rect 1595 1363 1597 1367
rect 1599 1363 1600 1367
rect 1617 1363 1618 1367
rect 1620 1363 1621 1367
rect 1633 1363 1638 1367
rect 1640 1363 1643 1367
rect 1645 1363 1646 1367
rect 1660 1363 1661 1367
rect 1663 1363 1664 1367
rect 1819 1368 1820 1372
rect 1822 1368 1823 1372
rect 1909 1368 1910 1372
rect 1912 1368 1913 1372
rect 577 1317 578 1321
rect 580 1317 581 1321
rect 593 1317 594 1321
rect 596 1317 597 1321
rect 609 1317 610 1321
rect 612 1317 613 1321
rect 628 1317 633 1321
rect 635 1317 638 1321
rect 640 1317 641 1321
rect 662 1317 664 1321
rect 666 1317 667 1321
rect 684 1317 685 1321
rect 687 1317 688 1321
rect 700 1317 705 1321
rect 707 1317 710 1321
rect 712 1317 713 1321
rect 727 1317 728 1321
rect 730 1317 731 1321
rect 775 1314 778 1318
rect 780 1314 783 1318
rect 785 1314 786 1318
rect 856 1314 859 1318
rect 861 1314 864 1318
rect 866 1314 867 1318
rect 946 1314 949 1318
rect 951 1314 954 1318
rect 956 1314 957 1318
rect 1510 1317 1511 1321
rect 1513 1317 1514 1321
rect 1526 1317 1527 1321
rect 1529 1317 1530 1321
rect 1542 1317 1543 1321
rect 1545 1317 1546 1321
rect 1561 1317 1566 1321
rect 1568 1317 1571 1321
rect 1573 1317 1574 1321
rect 1595 1317 1597 1321
rect 1599 1317 1600 1321
rect 1617 1317 1618 1321
rect 1620 1317 1621 1321
rect 1633 1317 1638 1321
rect 1640 1317 1643 1321
rect 1645 1317 1646 1321
rect 1660 1317 1661 1321
rect 1663 1317 1664 1321
rect 1708 1314 1711 1318
rect 1713 1314 1716 1318
rect 1718 1314 1719 1318
rect 1789 1314 1792 1318
rect 1794 1314 1797 1318
rect 1799 1314 1800 1318
rect 1879 1314 1882 1318
rect 1884 1314 1887 1318
rect 1889 1314 1890 1318
rect 775 1240 778 1244
rect 780 1240 783 1244
rect 785 1240 786 1244
rect 805 1236 806 1240
rect 808 1236 809 1240
rect 577 1231 578 1235
rect 580 1231 581 1235
rect 593 1231 594 1235
rect 596 1231 597 1235
rect 609 1231 610 1235
rect 612 1231 613 1235
rect 628 1231 633 1235
rect 635 1231 638 1235
rect 640 1231 641 1235
rect 662 1231 664 1235
rect 666 1231 667 1235
rect 684 1231 685 1235
rect 687 1231 688 1235
rect 700 1231 705 1235
rect 707 1231 710 1235
rect 712 1231 713 1235
rect 727 1231 728 1235
rect 730 1231 731 1235
rect 1708 1240 1711 1244
rect 1713 1240 1716 1244
rect 1718 1240 1719 1244
rect 1738 1236 1739 1240
rect 1741 1236 1742 1240
rect 1510 1231 1511 1235
rect 1513 1231 1514 1235
rect 1526 1231 1527 1235
rect 1529 1231 1530 1235
rect 1542 1231 1543 1235
rect 1545 1231 1546 1235
rect 1561 1231 1566 1235
rect 1568 1231 1571 1235
rect 1573 1231 1574 1235
rect 1595 1231 1597 1235
rect 1599 1231 1600 1235
rect 1617 1231 1618 1235
rect 1620 1231 1621 1235
rect 1633 1231 1638 1235
rect 1640 1231 1643 1235
rect 1645 1231 1646 1235
rect 1660 1231 1661 1235
rect 1663 1231 1664 1235
rect 577 1185 578 1189
rect 580 1185 581 1189
rect 593 1185 594 1189
rect 596 1185 597 1189
rect 609 1185 610 1189
rect 612 1185 613 1189
rect 628 1185 633 1189
rect 635 1185 638 1189
rect 640 1185 641 1189
rect 662 1185 664 1189
rect 666 1185 667 1189
rect 684 1185 685 1189
rect 687 1185 688 1189
rect 700 1185 705 1189
rect 707 1185 710 1189
rect 712 1185 713 1189
rect 727 1185 728 1189
rect 730 1185 731 1189
rect 811 1185 812 1189
rect 814 1185 815 1189
rect 819 1185 825 1189
rect 829 1185 830 1189
rect 832 1185 833 1189
rect 854 1185 855 1189
rect 857 1185 858 1189
rect 870 1185 871 1189
rect 873 1185 874 1189
rect 889 1185 894 1189
rect 896 1185 899 1189
rect 901 1185 902 1189
rect 923 1185 925 1189
rect 927 1185 928 1189
rect 945 1185 946 1189
rect 948 1185 949 1189
rect 961 1185 966 1189
rect 968 1185 971 1189
rect 973 1185 974 1189
rect 988 1185 989 1189
rect 991 1185 992 1189
rect 100 1171 101 1175
rect 103 1171 106 1175
rect 108 1171 109 1175
rect 121 1171 122 1175
rect 124 1171 125 1175
rect 137 1171 138 1175
rect 140 1171 143 1175
rect 145 1171 146 1175
rect 163 1171 164 1175
rect 166 1171 167 1175
rect 179 1171 180 1175
rect 182 1171 183 1175
rect 195 1171 196 1175
rect 198 1171 201 1175
rect 203 1171 204 1175
rect 216 1171 217 1175
rect 219 1171 220 1175
rect 232 1171 233 1175
rect 235 1171 238 1175
rect 240 1171 241 1175
rect 253 1171 254 1175
rect 256 1171 257 1175
rect 269 1171 270 1175
rect 272 1171 275 1175
rect 277 1171 278 1175
rect 295 1171 296 1175
rect 298 1171 299 1175
rect 311 1171 312 1175
rect 314 1171 315 1175
rect 327 1171 328 1175
rect 330 1171 333 1175
rect 335 1171 336 1175
rect 348 1171 349 1175
rect 351 1171 352 1175
rect 364 1171 365 1175
rect 367 1171 370 1175
rect 372 1171 373 1175
rect 385 1171 386 1175
rect 388 1171 389 1175
rect 401 1171 402 1175
rect 404 1171 407 1175
rect 409 1171 410 1175
rect 427 1171 428 1175
rect 430 1171 431 1175
rect 443 1171 444 1175
rect 446 1171 447 1175
rect 459 1171 460 1175
rect 462 1171 465 1175
rect 467 1171 468 1175
rect 480 1171 481 1175
rect 483 1171 484 1175
rect 775 1178 778 1182
rect 780 1178 783 1182
rect 785 1178 786 1182
rect 1510 1185 1511 1189
rect 1513 1185 1514 1189
rect 1526 1185 1527 1189
rect 1529 1185 1530 1189
rect 1542 1185 1543 1189
rect 1545 1185 1546 1189
rect 1561 1185 1566 1189
rect 1568 1185 1571 1189
rect 1573 1185 1574 1189
rect 1595 1185 1597 1189
rect 1599 1185 1600 1189
rect 1617 1185 1618 1189
rect 1620 1185 1621 1189
rect 1633 1185 1638 1189
rect 1640 1185 1643 1189
rect 1645 1185 1646 1189
rect 1660 1185 1661 1189
rect 1663 1185 1664 1189
rect 1744 1185 1745 1189
rect 1747 1185 1748 1189
rect 1752 1185 1758 1189
rect 1762 1185 1763 1189
rect 1765 1185 1766 1189
rect 1787 1185 1788 1189
rect 1790 1185 1791 1189
rect 1803 1185 1804 1189
rect 1806 1185 1807 1189
rect 1822 1185 1827 1189
rect 1829 1185 1832 1189
rect 1834 1185 1835 1189
rect 1856 1185 1858 1189
rect 1860 1185 1861 1189
rect 1878 1185 1879 1189
rect 1881 1185 1882 1189
rect 1894 1185 1899 1189
rect 1901 1185 1904 1189
rect 1906 1185 1907 1189
rect 1921 1185 1922 1189
rect 1924 1185 1925 1189
rect 1033 1171 1034 1175
rect 1036 1171 1039 1175
rect 1041 1171 1042 1175
rect 1054 1171 1055 1175
rect 1057 1171 1058 1175
rect 1070 1171 1071 1175
rect 1073 1171 1076 1175
rect 1078 1171 1079 1175
rect 1096 1171 1097 1175
rect 1099 1171 1100 1175
rect 1112 1171 1113 1175
rect 1115 1171 1116 1175
rect 1128 1171 1129 1175
rect 1131 1171 1134 1175
rect 1136 1171 1137 1175
rect 1149 1171 1150 1175
rect 1152 1171 1153 1175
rect 1165 1171 1166 1175
rect 1168 1171 1171 1175
rect 1173 1171 1174 1175
rect 1186 1171 1187 1175
rect 1189 1171 1190 1175
rect 1202 1171 1203 1175
rect 1205 1171 1208 1175
rect 1210 1171 1211 1175
rect 1228 1171 1229 1175
rect 1231 1171 1232 1175
rect 1244 1171 1245 1175
rect 1247 1171 1248 1175
rect 1260 1171 1261 1175
rect 1263 1171 1266 1175
rect 1268 1171 1269 1175
rect 1281 1171 1282 1175
rect 1284 1171 1285 1175
rect 1297 1171 1298 1175
rect 1300 1171 1303 1175
rect 1305 1171 1306 1175
rect 1318 1171 1319 1175
rect 1321 1171 1322 1175
rect 1334 1171 1335 1175
rect 1337 1171 1340 1175
rect 1342 1171 1343 1175
rect 1360 1171 1361 1175
rect 1363 1171 1364 1175
rect 1376 1171 1377 1175
rect 1379 1171 1380 1175
rect 1392 1171 1393 1175
rect 1395 1171 1398 1175
rect 1400 1171 1401 1175
rect 1413 1171 1414 1175
rect 1416 1171 1417 1175
rect 1708 1178 1711 1182
rect 1713 1178 1716 1182
rect 1718 1178 1719 1182
rect 215 1127 216 1131
rect 218 1127 219 1131
rect 239 1127 240 1131
rect 242 1127 243 1131
rect 1001 1131 1005 1132
rect 1001 1128 1005 1129
rect 1148 1127 1149 1131
rect 1151 1127 1152 1131
rect 1172 1127 1173 1131
rect 1175 1127 1176 1131
rect 1934 1131 1938 1132
rect 1934 1128 1938 1129
rect 235 1116 236 1120
rect 238 1116 239 1120
rect 1168 1116 1169 1120
rect 1171 1116 1172 1120
rect 227 1104 231 1105
rect 227 1101 231 1102
rect 1160 1104 1164 1105
rect 1160 1101 1164 1102
rect 215 1093 216 1097
rect 218 1093 219 1097
rect 239 1093 240 1097
rect 242 1093 243 1097
rect 1148 1093 1149 1097
rect 1151 1093 1152 1097
rect 1172 1093 1173 1097
rect 1175 1093 1176 1097
rect 871 1061 872 1065
rect 874 1061 877 1065
rect 879 1061 880 1065
rect 892 1061 893 1065
rect 895 1061 896 1065
rect 908 1061 909 1065
rect 911 1061 914 1065
rect 916 1061 917 1065
rect 934 1061 935 1065
rect 937 1061 938 1065
rect 950 1061 951 1065
rect 953 1061 954 1065
rect 966 1061 967 1065
rect 969 1061 972 1065
rect 974 1061 975 1065
rect 987 1061 988 1065
rect 990 1061 991 1065
rect 1804 1061 1805 1065
rect 1807 1061 1810 1065
rect 1812 1061 1813 1065
rect 1825 1061 1826 1065
rect 1828 1061 1829 1065
rect 1841 1061 1842 1065
rect 1844 1061 1847 1065
rect 1849 1061 1850 1065
rect 1867 1061 1868 1065
rect 1870 1061 1871 1065
rect 1883 1061 1884 1065
rect 1886 1061 1887 1065
rect 1899 1061 1900 1065
rect 1902 1061 1905 1065
rect 1907 1061 1908 1065
rect 1920 1061 1921 1065
rect 1923 1061 1924 1065
rect 100 1031 101 1035
rect 103 1031 106 1035
rect 108 1031 109 1035
rect 121 1031 122 1035
rect 124 1031 125 1035
rect 137 1031 138 1035
rect 140 1031 143 1035
rect 145 1031 146 1035
rect 163 1031 164 1035
rect 166 1031 167 1035
rect 179 1031 180 1035
rect 182 1031 183 1035
rect 195 1031 196 1035
rect 198 1031 201 1035
rect 203 1031 204 1035
rect 216 1031 217 1035
rect 219 1031 220 1035
rect 232 1031 233 1035
rect 235 1031 238 1035
rect 240 1031 241 1035
rect 253 1031 254 1035
rect 256 1031 257 1035
rect 269 1031 270 1035
rect 272 1031 275 1035
rect 277 1031 278 1035
rect 295 1031 296 1035
rect 298 1031 299 1035
rect 311 1031 312 1035
rect 314 1031 315 1035
rect 327 1031 328 1035
rect 330 1031 333 1035
rect 335 1031 336 1035
rect 348 1031 349 1035
rect 351 1031 352 1035
rect 364 1031 365 1035
rect 367 1031 370 1035
rect 372 1031 373 1035
rect 385 1031 386 1035
rect 388 1031 389 1035
rect 401 1031 402 1035
rect 404 1031 407 1035
rect 409 1031 410 1035
rect 427 1031 428 1035
rect 430 1031 431 1035
rect 443 1031 444 1035
rect 446 1031 447 1035
rect 459 1031 460 1035
rect 462 1031 465 1035
rect 467 1031 468 1035
rect 480 1031 481 1035
rect 483 1031 484 1035
rect 1033 1031 1034 1035
rect 1036 1031 1039 1035
rect 1041 1031 1042 1035
rect 1054 1031 1055 1035
rect 1057 1031 1058 1035
rect 1070 1031 1071 1035
rect 1073 1031 1076 1035
rect 1078 1031 1079 1035
rect 1096 1031 1097 1035
rect 1099 1031 1100 1035
rect 1112 1031 1113 1035
rect 1115 1031 1116 1035
rect 1128 1031 1129 1035
rect 1131 1031 1134 1035
rect 1136 1031 1137 1035
rect 1149 1031 1150 1035
rect 1152 1031 1153 1035
rect 1165 1031 1166 1035
rect 1168 1031 1171 1035
rect 1173 1031 1174 1035
rect 1186 1031 1187 1035
rect 1189 1031 1190 1035
rect 1202 1031 1203 1035
rect 1205 1031 1208 1035
rect 1210 1031 1211 1035
rect 1228 1031 1229 1035
rect 1231 1031 1232 1035
rect 1244 1031 1245 1035
rect 1247 1031 1248 1035
rect 1260 1031 1261 1035
rect 1263 1031 1266 1035
rect 1268 1031 1269 1035
rect 1281 1031 1282 1035
rect 1284 1031 1285 1035
rect 1297 1031 1298 1035
rect 1300 1031 1303 1035
rect 1305 1031 1306 1035
rect 1318 1031 1319 1035
rect 1321 1031 1322 1035
rect 1334 1031 1335 1035
rect 1337 1031 1340 1035
rect 1342 1031 1343 1035
rect 1360 1031 1361 1035
rect 1363 1031 1364 1035
rect 1376 1031 1377 1035
rect 1379 1031 1380 1035
rect 1392 1031 1393 1035
rect 1395 1031 1398 1035
rect 1400 1031 1401 1035
rect 1413 1031 1414 1035
rect 1416 1031 1417 1035
rect 1013 987 1017 988
rect 1013 984 1017 985
rect 1946 987 1950 988
rect 1946 984 1950 985
rect 871 975 872 979
rect 874 975 877 979
rect 879 975 880 979
rect 892 975 893 979
rect 895 975 896 979
rect 908 975 909 979
rect 911 975 914 979
rect 916 975 917 979
rect 934 975 935 979
rect 937 975 938 979
rect 950 975 951 979
rect 953 975 954 979
rect 966 975 967 979
rect 969 975 972 979
rect 974 975 975 979
rect 987 975 988 979
rect 990 975 991 979
rect 1804 975 1805 979
rect 1807 975 1810 979
rect 1812 975 1813 979
rect 1825 975 1826 979
rect 1828 975 1829 979
rect 1841 975 1842 979
rect 1844 975 1847 979
rect 1849 975 1850 979
rect 1867 975 1868 979
rect 1870 975 1871 979
rect 1883 975 1884 979
rect 1886 975 1887 979
rect 1899 975 1900 979
rect 1902 975 1905 979
rect 1907 975 1908 979
rect 1920 975 1921 979
rect 1923 975 1924 979
rect 100 945 101 949
rect 103 945 106 949
rect 108 945 109 949
rect 121 945 122 949
rect 124 945 125 949
rect 137 945 138 949
rect 140 945 143 949
rect 145 945 146 949
rect 163 945 164 949
rect 166 945 167 949
rect 179 945 180 949
rect 182 945 183 949
rect 195 945 196 949
rect 198 945 201 949
rect 203 945 204 949
rect 216 945 217 949
rect 219 945 220 949
rect 232 945 233 949
rect 235 945 238 949
rect 240 945 241 949
rect 253 945 254 949
rect 256 945 257 949
rect 269 945 270 949
rect 272 945 275 949
rect 277 945 278 949
rect 295 945 296 949
rect 298 945 299 949
rect 311 945 312 949
rect 314 945 315 949
rect 327 945 328 949
rect 330 945 333 949
rect 335 945 336 949
rect 348 945 349 949
rect 351 945 352 949
rect 364 945 365 949
rect 367 945 370 949
rect 372 945 373 949
rect 385 945 386 949
rect 388 945 389 949
rect 401 945 402 949
rect 404 945 407 949
rect 409 945 410 949
rect 427 945 428 949
rect 430 945 431 949
rect 443 945 444 949
rect 446 945 447 949
rect 459 945 460 949
rect 462 945 465 949
rect 467 945 468 949
rect 480 945 481 949
rect 483 945 484 949
rect 1033 945 1034 949
rect 1036 945 1039 949
rect 1041 945 1042 949
rect 1054 945 1055 949
rect 1057 945 1058 949
rect 1070 945 1071 949
rect 1073 945 1076 949
rect 1078 945 1079 949
rect 1096 945 1097 949
rect 1099 945 1100 949
rect 1112 945 1113 949
rect 1115 945 1116 949
rect 1128 945 1129 949
rect 1131 945 1134 949
rect 1136 945 1137 949
rect 1149 945 1150 949
rect 1152 945 1153 949
rect 1165 945 1166 949
rect 1168 945 1171 949
rect 1173 945 1174 949
rect 1186 945 1187 949
rect 1189 945 1190 949
rect 1202 945 1203 949
rect 1205 945 1208 949
rect 1210 945 1211 949
rect 1228 945 1229 949
rect 1231 945 1232 949
rect 1244 945 1245 949
rect 1247 945 1248 949
rect 1260 945 1261 949
rect 1263 945 1266 949
rect 1268 945 1269 949
rect 1281 945 1282 949
rect 1284 945 1285 949
rect 1297 945 1298 949
rect 1300 945 1303 949
rect 1305 945 1306 949
rect 1318 945 1319 949
rect 1321 945 1322 949
rect 1334 945 1335 949
rect 1337 945 1340 949
rect 1342 945 1343 949
rect 1360 945 1361 949
rect 1363 945 1364 949
rect 1376 945 1377 949
rect 1379 945 1380 949
rect 1392 945 1393 949
rect 1395 945 1398 949
rect 1400 945 1401 949
rect 1413 945 1414 949
rect 1416 945 1417 949
rect 332 901 333 905
rect 335 901 336 905
rect 356 901 357 905
rect 359 901 360 905
rect 1265 901 1266 905
rect 1268 901 1269 905
rect 1289 901 1290 905
rect 1292 901 1293 905
rect 352 890 353 894
rect 355 890 356 894
rect 1285 890 1286 894
rect 1288 890 1289 894
rect 344 878 348 879
rect 344 875 348 876
rect 1277 878 1281 879
rect 1277 875 1281 876
rect 332 867 333 871
rect 335 867 336 871
rect 356 867 357 871
rect 359 867 360 871
rect 1265 867 1266 871
rect 1268 867 1269 871
rect 1289 867 1290 871
rect 1292 867 1293 871
rect 100 805 101 809
rect 103 805 106 809
rect 108 805 109 809
rect 121 805 122 809
rect 124 805 125 809
rect 137 805 138 809
rect 140 805 143 809
rect 145 805 146 809
rect 163 805 164 809
rect 166 805 167 809
rect 179 805 180 809
rect 182 805 183 809
rect 195 805 196 809
rect 198 805 201 809
rect 203 805 204 809
rect 216 805 217 809
rect 219 805 220 809
rect 232 805 233 809
rect 235 805 238 809
rect 240 805 241 809
rect 253 805 254 809
rect 256 805 257 809
rect 269 805 270 809
rect 272 805 275 809
rect 277 805 278 809
rect 295 805 296 809
rect 298 805 299 809
rect 311 805 312 809
rect 314 805 315 809
rect 327 805 328 809
rect 330 805 333 809
rect 335 805 336 809
rect 348 805 349 809
rect 351 805 352 809
rect 364 805 365 809
rect 367 805 370 809
rect 372 805 373 809
rect 385 805 386 809
rect 388 805 389 809
rect 401 805 402 809
rect 404 805 407 809
rect 409 805 410 809
rect 427 805 428 809
rect 430 805 431 809
rect 443 805 444 809
rect 446 805 447 809
rect 459 805 460 809
rect 462 805 465 809
rect 467 805 468 809
rect 480 805 481 809
rect 483 805 484 809
rect 1033 805 1034 809
rect 1036 805 1039 809
rect 1041 805 1042 809
rect 1054 805 1055 809
rect 1057 805 1058 809
rect 1070 805 1071 809
rect 1073 805 1076 809
rect 1078 805 1079 809
rect 1096 805 1097 809
rect 1099 805 1100 809
rect 1112 805 1113 809
rect 1115 805 1116 809
rect 1128 805 1129 809
rect 1131 805 1134 809
rect 1136 805 1137 809
rect 1149 805 1150 809
rect 1152 805 1153 809
rect 1165 805 1166 809
rect 1168 805 1171 809
rect 1173 805 1174 809
rect 1186 805 1187 809
rect 1189 805 1190 809
rect 1202 805 1203 809
rect 1205 805 1208 809
rect 1210 805 1211 809
rect 1228 805 1229 809
rect 1231 805 1232 809
rect 1244 805 1245 809
rect 1247 805 1248 809
rect 1260 805 1261 809
rect 1263 805 1266 809
rect 1268 805 1269 809
rect 1281 805 1282 809
rect 1284 805 1285 809
rect 1297 805 1298 809
rect 1300 805 1303 809
rect 1305 805 1306 809
rect 1318 805 1319 809
rect 1321 805 1322 809
rect 1334 805 1335 809
rect 1337 805 1340 809
rect 1342 805 1343 809
rect 1360 805 1361 809
rect 1363 805 1364 809
rect 1376 805 1377 809
rect 1379 805 1380 809
rect 1392 805 1393 809
rect 1395 805 1398 809
rect 1400 805 1401 809
rect 1413 805 1414 809
rect 1416 805 1417 809
rect 572 726 573 730
rect 575 726 578 730
rect 580 726 581 730
rect 593 726 594 730
rect 596 726 597 730
rect 609 726 610 730
rect 612 726 615 730
rect 617 726 618 730
rect 635 726 636 730
rect 638 726 639 730
rect 651 726 652 730
rect 654 726 655 730
rect 667 726 668 730
rect 670 726 673 730
rect 675 726 676 730
rect 688 726 689 730
rect 691 726 692 730
rect 704 726 705 730
rect 707 726 710 730
rect 712 726 713 730
rect 725 726 726 730
rect 728 726 729 730
rect 741 726 742 730
rect 744 726 747 730
rect 749 726 750 730
rect 767 726 768 730
rect 770 726 771 730
rect 783 726 784 730
rect 786 726 787 730
rect 799 726 800 730
rect 802 726 805 730
rect 807 726 808 730
rect 820 726 821 730
rect 823 726 824 730
rect 836 726 837 730
rect 839 726 842 730
rect 844 726 845 730
rect 857 726 858 730
rect 860 726 861 730
rect 873 726 874 730
rect 876 726 879 730
rect 881 726 882 730
rect 899 726 900 730
rect 902 726 903 730
rect 915 726 916 730
rect 918 726 919 730
rect 931 726 932 730
rect 934 726 937 730
rect 939 726 940 730
rect 952 726 953 730
rect 955 726 956 730
rect 968 726 969 730
rect 971 726 974 730
rect 976 726 977 730
rect 989 726 990 730
rect 992 726 993 730
rect 1005 726 1006 730
rect 1008 726 1011 730
rect 1013 726 1014 730
rect 1031 726 1032 730
rect 1034 726 1035 730
rect 1047 726 1048 730
rect 1050 726 1051 730
rect 1063 726 1064 730
rect 1066 726 1069 730
rect 1071 726 1072 730
rect 1084 726 1085 730
rect 1087 726 1088 730
rect 1505 726 1506 730
rect 1508 726 1511 730
rect 1513 726 1514 730
rect 1526 726 1527 730
rect 1529 726 1530 730
rect 1542 726 1543 730
rect 1545 726 1548 730
rect 1550 726 1551 730
rect 1568 726 1569 730
rect 1571 726 1572 730
rect 1584 726 1585 730
rect 1587 726 1588 730
rect 1600 726 1601 730
rect 1603 726 1606 730
rect 1608 726 1609 730
rect 1621 726 1622 730
rect 1624 726 1625 730
rect 1637 726 1638 730
rect 1640 726 1643 730
rect 1645 726 1646 730
rect 1658 726 1659 730
rect 1661 726 1662 730
rect 1674 726 1675 730
rect 1677 726 1680 730
rect 1682 726 1683 730
rect 1700 726 1701 730
rect 1703 726 1704 730
rect 1716 726 1717 730
rect 1719 726 1720 730
rect 1732 726 1733 730
rect 1735 726 1738 730
rect 1740 726 1741 730
rect 1753 726 1754 730
rect 1756 726 1757 730
rect 1769 726 1770 730
rect 1772 726 1775 730
rect 1777 726 1778 730
rect 1790 726 1791 730
rect 1793 726 1794 730
rect 1806 726 1807 730
rect 1809 726 1812 730
rect 1814 726 1815 730
rect 1832 726 1833 730
rect 1835 726 1836 730
rect 1848 726 1849 730
rect 1851 726 1852 730
rect 1864 726 1865 730
rect 1867 726 1870 730
rect 1872 726 1873 730
rect 1885 726 1886 730
rect 1888 726 1889 730
rect 1901 726 1902 730
rect 1904 726 1907 730
rect 1909 726 1910 730
rect 1922 726 1923 730
rect 1925 726 1926 730
rect 1938 726 1939 730
rect 1941 726 1944 730
rect 1946 726 1947 730
rect 1964 726 1965 730
rect 1967 726 1968 730
rect 1980 726 1981 730
rect 1983 726 1984 730
rect 1996 726 1997 730
rect 1999 726 2002 730
rect 2004 726 2005 730
rect 2017 726 2018 730
rect 2020 726 2021 730
rect 232 693 233 697
rect 235 693 238 697
rect 240 693 241 697
rect 253 693 254 697
rect 256 693 257 697
rect 269 693 270 697
rect 272 693 275 697
rect 277 693 278 697
rect 295 693 296 697
rect 298 693 299 697
rect 311 693 312 697
rect 314 693 315 697
rect 327 693 328 697
rect 330 693 333 697
rect 335 693 336 697
rect 348 693 349 697
rect 351 693 352 697
rect 1165 693 1166 697
rect 1168 693 1171 697
rect 1173 693 1174 697
rect 1186 693 1187 697
rect 1189 693 1190 697
rect 1202 693 1203 697
rect 1205 693 1208 697
rect 1210 693 1211 697
rect 1228 693 1229 697
rect 1231 693 1232 697
rect 1244 693 1245 697
rect 1247 693 1248 697
rect 1260 693 1261 697
rect 1263 693 1266 697
rect 1268 693 1269 697
rect 1281 693 1282 697
rect 1284 693 1285 697
rect 356 656 357 660
rect 359 656 360 660
rect 751 660 752 664
rect 754 660 755 664
rect 775 656 778 660
rect 780 656 783 660
rect 785 656 786 660
rect 832 660 833 664
rect 835 660 836 664
rect 856 656 859 660
rect 861 656 864 660
rect 866 656 867 660
rect 805 652 806 656
rect 808 652 809 656
rect 239 647 240 651
rect 242 647 243 651
rect 577 647 578 651
rect 580 647 581 651
rect 593 647 594 651
rect 596 647 597 651
rect 609 647 610 651
rect 612 647 613 651
rect 628 647 633 651
rect 635 647 638 651
rect 640 647 641 651
rect 662 647 664 651
rect 666 647 667 651
rect 684 647 685 651
rect 687 647 688 651
rect 700 647 705 651
rect 707 647 710 651
rect 712 647 713 651
rect 727 647 728 651
rect 730 647 731 651
rect 886 652 887 656
rect 889 652 890 656
rect 1289 656 1290 660
rect 1292 656 1293 660
rect 1684 660 1685 664
rect 1687 660 1688 664
rect 1708 656 1711 660
rect 1713 656 1716 660
rect 1718 656 1719 660
rect 1765 660 1766 664
rect 1768 660 1769 664
rect 1789 656 1792 660
rect 1794 656 1797 660
rect 1799 656 1800 660
rect 1738 652 1739 656
rect 1741 652 1742 656
rect 1172 647 1173 651
rect 1175 647 1176 651
rect 1510 647 1511 651
rect 1513 647 1514 651
rect 1526 647 1527 651
rect 1529 647 1530 651
rect 1542 647 1543 651
rect 1545 647 1546 651
rect 1561 647 1566 651
rect 1568 647 1571 651
rect 1573 647 1574 651
rect 1595 647 1597 651
rect 1599 647 1600 651
rect 1617 647 1618 651
rect 1620 647 1621 651
rect 1633 647 1638 651
rect 1640 647 1643 651
rect 1645 647 1646 651
rect 1660 647 1661 651
rect 1663 647 1664 651
rect 1819 652 1820 656
rect 1822 652 1823 656
rect 577 601 578 605
rect 580 601 581 605
rect 593 601 594 605
rect 596 601 597 605
rect 609 601 610 605
rect 612 601 613 605
rect 628 601 633 605
rect 635 601 638 605
rect 640 601 641 605
rect 662 601 664 605
rect 666 601 667 605
rect 684 601 685 605
rect 687 601 688 605
rect 700 601 705 605
rect 707 601 710 605
rect 712 601 713 605
rect 727 601 728 605
rect 730 601 731 605
rect 223 591 224 595
rect 226 591 227 595
rect 239 591 240 595
rect 242 591 245 595
rect 247 591 248 595
rect 260 591 261 595
rect 263 591 264 595
rect 276 591 277 595
rect 279 591 280 595
rect 297 591 298 595
rect 300 591 303 595
rect 305 591 306 595
rect 318 591 319 595
rect 321 591 322 595
rect 334 591 335 595
rect 337 591 340 595
rect 342 591 343 595
rect 775 600 778 604
rect 780 600 783 604
rect 785 600 786 604
rect 856 600 859 604
rect 861 600 864 604
rect 866 600 867 604
rect 1510 601 1511 605
rect 1513 601 1514 605
rect 1526 601 1527 605
rect 1529 601 1530 605
rect 1542 601 1543 605
rect 1545 601 1546 605
rect 1561 601 1566 605
rect 1568 601 1571 605
rect 1573 601 1574 605
rect 1595 601 1597 605
rect 1599 601 1600 605
rect 1617 601 1618 605
rect 1620 601 1621 605
rect 1633 601 1638 605
rect 1640 601 1643 605
rect 1645 601 1646 605
rect 1660 601 1661 605
rect 1663 601 1664 605
rect 1156 591 1157 595
rect 1159 591 1160 595
rect 1172 591 1173 595
rect 1175 591 1178 595
rect 1180 591 1181 595
rect 1193 591 1194 595
rect 1196 591 1197 595
rect 1209 591 1210 595
rect 1212 591 1213 595
rect 1230 591 1231 595
rect 1233 591 1236 595
rect 1238 591 1239 595
rect 1251 591 1252 595
rect 1254 591 1255 595
rect 1267 591 1268 595
rect 1270 591 1273 595
rect 1275 591 1276 595
rect 1708 600 1711 604
rect 1713 600 1716 604
rect 1718 600 1719 604
rect 1789 600 1792 604
rect 1794 600 1797 604
rect 1799 600 1800 604
rect 775 524 778 528
rect 780 524 783 528
rect 785 524 786 528
rect 856 528 857 532
rect 859 528 860 532
rect 880 524 883 528
rect 885 524 888 528
rect 890 524 891 528
rect 805 520 806 524
rect 808 520 809 524
rect 577 515 578 519
rect 580 515 581 519
rect 593 515 594 519
rect 596 515 597 519
rect 609 515 610 519
rect 612 515 613 519
rect 628 515 633 519
rect 635 515 638 519
rect 640 515 641 519
rect 662 515 664 519
rect 666 515 667 519
rect 684 515 685 519
rect 687 515 688 519
rect 700 515 705 519
rect 707 515 710 519
rect 712 515 713 519
rect 727 515 728 519
rect 730 515 731 519
rect 910 520 911 524
rect 913 520 914 524
rect 1708 524 1711 528
rect 1713 524 1716 528
rect 1718 524 1719 528
rect 1789 528 1790 532
rect 1792 528 1793 532
rect 1813 524 1816 528
rect 1818 524 1821 528
rect 1823 524 1824 528
rect 1738 520 1739 524
rect 1741 520 1742 524
rect 1510 515 1511 519
rect 1513 515 1514 519
rect 1526 515 1527 519
rect 1529 515 1530 519
rect 1542 515 1543 519
rect 1545 515 1546 519
rect 1561 515 1566 519
rect 1568 515 1571 519
rect 1573 515 1574 519
rect 1595 515 1597 519
rect 1599 515 1600 519
rect 1617 515 1618 519
rect 1620 515 1621 519
rect 1633 515 1638 519
rect 1640 515 1643 519
rect 1645 515 1646 519
rect 1660 515 1661 519
rect 1663 515 1664 519
rect 1843 520 1844 524
rect 1846 520 1847 524
rect 577 469 578 473
rect 580 469 581 473
rect 593 469 594 473
rect 596 469 597 473
rect 609 469 610 473
rect 612 469 613 473
rect 628 469 633 473
rect 635 469 638 473
rect 640 469 641 473
rect 662 469 664 473
rect 666 469 667 473
rect 684 469 685 473
rect 687 469 688 473
rect 700 469 705 473
rect 707 469 710 473
rect 712 469 713 473
rect 727 469 728 473
rect 730 469 731 473
rect 775 469 778 473
rect 780 469 783 473
rect 785 469 786 473
rect 880 469 883 473
rect 885 469 888 473
rect 890 469 891 473
rect 1510 469 1511 473
rect 1513 469 1514 473
rect 1526 469 1527 473
rect 1529 469 1530 473
rect 1542 469 1543 473
rect 1545 469 1546 473
rect 1561 469 1566 473
rect 1568 469 1571 473
rect 1573 469 1574 473
rect 1595 469 1597 473
rect 1599 469 1600 473
rect 1617 469 1618 473
rect 1620 469 1621 473
rect 1633 469 1638 473
rect 1640 469 1643 473
rect 1645 469 1646 473
rect 1660 469 1661 473
rect 1663 469 1664 473
rect 1708 469 1711 473
rect 1713 469 1716 473
rect 1718 469 1719 473
rect 1813 469 1816 473
rect 1818 469 1821 473
rect 1823 469 1824 473
rect 775 392 778 396
rect 780 392 783 396
rect 785 392 786 396
rect 832 396 833 400
rect 835 396 836 400
rect 856 392 859 396
rect 861 392 864 396
rect 866 392 867 396
rect 922 396 923 400
rect 925 396 926 400
rect 946 392 949 396
rect 951 392 954 396
rect 956 392 957 396
rect 805 388 806 392
rect 808 388 809 392
rect 577 383 578 387
rect 580 383 581 387
rect 593 383 594 387
rect 596 383 597 387
rect 609 383 610 387
rect 612 383 613 387
rect 628 383 633 387
rect 635 383 638 387
rect 640 383 641 387
rect 662 383 664 387
rect 666 383 667 387
rect 684 383 685 387
rect 687 383 688 387
rect 700 383 705 387
rect 707 383 710 387
rect 712 383 713 387
rect 727 383 728 387
rect 730 383 731 387
rect 886 388 887 392
rect 889 388 890 392
rect 976 388 977 392
rect 979 388 980 392
rect 1708 392 1711 396
rect 1713 392 1716 396
rect 1718 392 1719 396
rect 1765 396 1766 400
rect 1768 396 1769 400
rect 1789 392 1792 396
rect 1794 392 1797 396
rect 1799 392 1800 396
rect 1855 396 1856 400
rect 1858 396 1859 400
rect 1879 392 1882 396
rect 1884 392 1887 396
rect 1889 392 1890 396
rect 1738 388 1739 392
rect 1741 388 1742 392
rect 1510 383 1511 387
rect 1513 383 1514 387
rect 1526 383 1527 387
rect 1529 383 1530 387
rect 1542 383 1543 387
rect 1545 383 1546 387
rect 1561 383 1566 387
rect 1568 383 1571 387
rect 1573 383 1574 387
rect 1595 383 1597 387
rect 1599 383 1600 387
rect 1617 383 1618 387
rect 1620 383 1621 387
rect 1633 383 1638 387
rect 1640 383 1643 387
rect 1645 383 1646 387
rect 1660 383 1661 387
rect 1663 383 1664 387
rect 1819 388 1820 392
rect 1822 388 1823 392
rect 1909 388 1910 392
rect 1912 388 1913 392
rect 577 337 578 341
rect 580 337 581 341
rect 593 337 594 341
rect 596 337 597 341
rect 609 337 610 341
rect 612 337 613 341
rect 628 337 633 341
rect 635 337 638 341
rect 640 337 641 341
rect 662 337 664 341
rect 666 337 667 341
rect 684 337 685 341
rect 687 337 688 341
rect 700 337 705 341
rect 707 337 710 341
rect 712 337 713 341
rect 727 337 728 341
rect 730 337 731 341
rect 775 334 778 338
rect 780 334 783 338
rect 785 334 786 338
rect 856 334 859 338
rect 861 334 864 338
rect 866 334 867 338
rect 946 334 949 338
rect 951 334 954 338
rect 956 334 957 338
rect 1510 337 1511 341
rect 1513 337 1514 341
rect 1526 337 1527 341
rect 1529 337 1530 341
rect 1542 337 1543 341
rect 1545 337 1546 341
rect 1561 337 1566 341
rect 1568 337 1571 341
rect 1573 337 1574 341
rect 1595 337 1597 341
rect 1599 337 1600 341
rect 1617 337 1618 341
rect 1620 337 1621 341
rect 1633 337 1638 341
rect 1640 337 1643 341
rect 1645 337 1646 341
rect 1660 337 1661 341
rect 1663 337 1664 341
rect 1708 334 1711 338
rect 1713 334 1716 338
rect 1718 334 1719 338
rect 1789 334 1792 338
rect 1794 334 1797 338
rect 1799 334 1800 338
rect 1879 334 1882 338
rect 1884 334 1887 338
rect 1889 334 1890 338
rect 775 260 778 264
rect 780 260 783 264
rect 785 260 786 264
rect 805 256 806 260
rect 808 256 809 260
rect 577 251 578 255
rect 580 251 581 255
rect 593 251 594 255
rect 596 251 597 255
rect 609 251 610 255
rect 612 251 613 255
rect 628 251 633 255
rect 635 251 638 255
rect 640 251 641 255
rect 662 251 664 255
rect 666 251 667 255
rect 684 251 685 255
rect 687 251 688 255
rect 700 251 705 255
rect 707 251 710 255
rect 712 251 713 255
rect 727 251 728 255
rect 730 251 731 255
rect 1708 260 1711 264
rect 1713 260 1716 264
rect 1718 260 1719 264
rect 1738 256 1739 260
rect 1741 256 1742 260
rect 1510 251 1511 255
rect 1513 251 1514 255
rect 1526 251 1527 255
rect 1529 251 1530 255
rect 1542 251 1543 255
rect 1545 251 1546 255
rect 1561 251 1566 255
rect 1568 251 1571 255
rect 1573 251 1574 255
rect 1595 251 1597 255
rect 1599 251 1600 255
rect 1617 251 1618 255
rect 1620 251 1621 255
rect 1633 251 1638 255
rect 1640 251 1643 255
rect 1645 251 1646 255
rect 1660 251 1661 255
rect 1663 251 1664 255
rect 577 205 578 209
rect 580 205 581 209
rect 593 205 594 209
rect 596 205 597 209
rect 609 205 610 209
rect 612 205 613 209
rect 628 205 633 209
rect 635 205 638 209
rect 640 205 641 209
rect 662 205 664 209
rect 666 205 667 209
rect 684 205 685 209
rect 687 205 688 209
rect 700 205 705 209
rect 707 205 710 209
rect 712 205 713 209
rect 727 205 728 209
rect 730 205 731 209
rect 811 205 812 209
rect 814 205 815 209
rect 819 205 825 209
rect 829 205 830 209
rect 832 205 833 209
rect 854 205 855 209
rect 857 205 858 209
rect 870 205 871 209
rect 873 205 874 209
rect 889 205 894 209
rect 896 205 899 209
rect 901 205 902 209
rect 923 205 925 209
rect 927 205 928 209
rect 945 205 946 209
rect 948 205 949 209
rect 961 205 966 209
rect 968 205 971 209
rect 973 205 974 209
rect 988 205 989 209
rect 991 205 992 209
rect 100 191 101 195
rect 103 191 106 195
rect 108 191 109 195
rect 121 191 122 195
rect 124 191 125 195
rect 137 191 138 195
rect 140 191 143 195
rect 145 191 146 195
rect 163 191 164 195
rect 166 191 167 195
rect 179 191 180 195
rect 182 191 183 195
rect 195 191 196 195
rect 198 191 201 195
rect 203 191 204 195
rect 216 191 217 195
rect 219 191 220 195
rect 232 191 233 195
rect 235 191 238 195
rect 240 191 241 195
rect 253 191 254 195
rect 256 191 257 195
rect 269 191 270 195
rect 272 191 275 195
rect 277 191 278 195
rect 295 191 296 195
rect 298 191 299 195
rect 311 191 312 195
rect 314 191 315 195
rect 327 191 328 195
rect 330 191 333 195
rect 335 191 336 195
rect 348 191 349 195
rect 351 191 352 195
rect 364 191 365 195
rect 367 191 370 195
rect 372 191 373 195
rect 385 191 386 195
rect 388 191 389 195
rect 401 191 402 195
rect 404 191 407 195
rect 409 191 410 195
rect 427 191 428 195
rect 430 191 431 195
rect 443 191 444 195
rect 446 191 447 195
rect 459 191 460 195
rect 462 191 465 195
rect 467 191 468 195
rect 480 191 481 195
rect 483 191 484 195
rect 775 198 778 202
rect 780 198 783 202
rect 785 198 786 202
rect 1510 205 1511 209
rect 1513 205 1514 209
rect 1526 205 1527 209
rect 1529 205 1530 209
rect 1542 205 1543 209
rect 1545 205 1546 209
rect 1561 205 1566 209
rect 1568 205 1571 209
rect 1573 205 1574 209
rect 1595 205 1597 209
rect 1599 205 1600 209
rect 1617 205 1618 209
rect 1620 205 1621 209
rect 1633 205 1638 209
rect 1640 205 1643 209
rect 1645 205 1646 209
rect 1660 205 1661 209
rect 1663 205 1664 209
rect 1744 205 1745 209
rect 1747 205 1748 209
rect 1752 205 1758 209
rect 1762 205 1763 209
rect 1765 205 1766 209
rect 1787 205 1788 209
rect 1790 205 1791 209
rect 1803 205 1804 209
rect 1806 205 1807 209
rect 1822 205 1827 209
rect 1829 205 1832 209
rect 1834 205 1835 209
rect 1856 205 1858 209
rect 1860 205 1861 209
rect 1878 205 1879 209
rect 1881 205 1882 209
rect 1894 205 1899 209
rect 1901 205 1904 209
rect 1906 205 1907 209
rect 1921 205 1922 209
rect 1924 205 1925 209
rect 1033 191 1034 195
rect 1036 191 1039 195
rect 1041 191 1042 195
rect 1054 191 1055 195
rect 1057 191 1058 195
rect 1070 191 1071 195
rect 1073 191 1076 195
rect 1078 191 1079 195
rect 1096 191 1097 195
rect 1099 191 1100 195
rect 1112 191 1113 195
rect 1115 191 1116 195
rect 1128 191 1129 195
rect 1131 191 1134 195
rect 1136 191 1137 195
rect 1149 191 1150 195
rect 1152 191 1153 195
rect 1165 191 1166 195
rect 1168 191 1171 195
rect 1173 191 1174 195
rect 1186 191 1187 195
rect 1189 191 1190 195
rect 1202 191 1203 195
rect 1205 191 1208 195
rect 1210 191 1211 195
rect 1228 191 1229 195
rect 1231 191 1232 195
rect 1244 191 1245 195
rect 1247 191 1248 195
rect 1260 191 1261 195
rect 1263 191 1266 195
rect 1268 191 1269 195
rect 1281 191 1282 195
rect 1284 191 1285 195
rect 1297 191 1298 195
rect 1300 191 1303 195
rect 1305 191 1306 195
rect 1318 191 1319 195
rect 1321 191 1322 195
rect 1334 191 1335 195
rect 1337 191 1340 195
rect 1342 191 1343 195
rect 1360 191 1361 195
rect 1363 191 1364 195
rect 1376 191 1377 195
rect 1379 191 1380 195
rect 1392 191 1393 195
rect 1395 191 1398 195
rect 1400 191 1401 195
rect 1413 191 1414 195
rect 1416 191 1417 195
rect 1708 198 1711 202
rect 1713 198 1716 202
rect 1718 198 1719 202
rect 215 147 216 151
rect 218 147 219 151
rect 239 147 240 151
rect 242 147 243 151
rect 1001 151 1005 152
rect 1001 148 1005 149
rect 1148 147 1149 151
rect 1151 147 1152 151
rect 1172 147 1173 151
rect 1175 147 1176 151
rect 1934 151 1938 152
rect 1934 148 1938 149
rect 235 136 236 140
rect 238 136 239 140
rect 1168 136 1169 140
rect 1171 136 1172 140
rect 227 124 231 125
rect 227 121 231 122
rect 1160 124 1164 125
rect 1160 121 1164 122
rect 215 113 216 117
rect 218 113 219 117
rect 239 113 240 117
rect 242 113 243 117
rect 1148 113 1149 117
rect 1151 113 1152 117
rect 1172 113 1173 117
rect 1175 113 1176 117
rect 871 81 872 85
rect 874 81 877 85
rect 879 81 880 85
rect 892 81 893 85
rect 895 81 896 85
rect 908 81 909 85
rect 911 81 914 85
rect 916 81 917 85
rect 934 81 935 85
rect 937 81 938 85
rect 950 81 951 85
rect 953 81 954 85
rect 966 81 967 85
rect 969 81 972 85
rect 974 81 975 85
rect 987 81 988 85
rect 990 81 991 85
rect 1804 81 1805 85
rect 1807 81 1810 85
rect 1812 81 1813 85
rect 1825 81 1826 85
rect 1828 81 1829 85
rect 1841 81 1842 85
rect 1844 81 1847 85
rect 1849 81 1850 85
rect 1867 81 1868 85
rect 1870 81 1871 85
rect 1883 81 1884 85
rect 1886 81 1887 85
rect 1899 81 1900 85
rect 1902 81 1905 85
rect 1907 81 1908 85
rect 1920 81 1921 85
rect 1923 81 1924 85
rect 100 51 101 55
rect 103 51 106 55
rect 108 51 109 55
rect 121 51 122 55
rect 124 51 125 55
rect 137 51 138 55
rect 140 51 143 55
rect 145 51 146 55
rect 163 51 164 55
rect 166 51 167 55
rect 179 51 180 55
rect 182 51 183 55
rect 195 51 196 55
rect 198 51 201 55
rect 203 51 204 55
rect 216 51 217 55
rect 219 51 220 55
rect 232 51 233 55
rect 235 51 238 55
rect 240 51 241 55
rect 253 51 254 55
rect 256 51 257 55
rect 269 51 270 55
rect 272 51 275 55
rect 277 51 278 55
rect 295 51 296 55
rect 298 51 299 55
rect 311 51 312 55
rect 314 51 315 55
rect 327 51 328 55
rect 330 51 333 55
rect 335 51 336 55
rect 348 51 349 55
rect 351 51 352 55
rect 364 51 365 55
rect 367 51 370 55
rect 372 51 373 55
rect 385 51 386 55
rect 388 51 389 55
rect 401 51 402 55
rect 404 51 407 55
rect 409 51 410 55
rect 427 51 428 55
rect 430 51 431 55
rect 443 51 444 55
rect 446 51 447 55
rect 459 51 460 55
rect 462 51 465 55
rect 467 51 468 55
rect 480 51 481 55
rect 483 51 484 55
rect 1033 51 1034 55
rect 1036 51 1039 55
rect 1041 51 1042 55
rect 1054 51 1055 55
rect 1057 51 1058 55
rect 1070 51 1071 55
rect 1073 51 1076 55
rect 1078 51 1079 55
rect 1096 51 1097 55
rect 1099 51 1100 55
rect 1112 51 1113 55
rect 1115 51 1116 55
rect 1128 51 1129 55
rect 1131 51 1134 55
rect 1136 51 1137 55
rect 1149 51 1150 55
rect 1152 51 1153 55
rect 1165 51 1166 55
rect 1168 51 1171 55
rect 1173 51 1174 55
rect 1186 51 1187 55
rect 1189 51 1190 55
rect 1202 51 1203 55
rect 1205 51 1208 55
rect 1210 51 1211 55
rect 1228 51 1229 55
rect 1231 51 1232 55
rect 1244 51 1245 55
rect 1247 51 1248 55
rect 1260 51 1261 55
rect 1263 51 1266 55
rect 1268 51 1269 55
rect 1281 51 1282 55
rect 1284 51 1285 55
rect 1297 51 1298 55
rect 1300 51 1303 55
rect 1305 51 1306 55
rect 1318 51 1319 55
rect 1321 51 1322 55
rect 1334 51 1335 55
rect 1337 51 1340 55
rect 1342 51 1343 55
rect 1360 51 1361 55
rect 1363 51 1364 55
rect 1376 51 1377 55
rect 1379 51 1380 55
rect 1392 51 1393 55
rect 1395 51 1398 55
rect 1400 51 1401 55
rect 1413 51 1414 55
rect 1416 51 1417 55
rect 1013 7 1017 8
rect 1013 4 1017 5
rect 1946 7 1950 8
rect 1946 4 1950 5
rect 871 -5 872 -1
rect 874 -5 877 -1
rect 879 -5 880 -1
rect 892 -5 893 -1
rect 895 -5 896 -1
rect 908 -5 909 -1
rect 911 -5 914 -1
rect 916 -5 917 -1
rect 934 -5 935 -1
rect 937 -5 938 -1
rect 950 -5 951 -1
rect 953 -5 954 -1
rect 966 -5 967 -1
rect 969 -5 972 -1
rect 974 -5 975 -1
rect 987 -5 988 -1
rect 990 -5 991 -1
rect 1804 -5 1805 -1
rect 1807 -5 1810 -1
rect 1812 -5 1813 -1
rect 1825 -5 1826 -1
rect 1828 -5 1829 -1
rect 1841 -5 1842 -1
rect 1844 -5 1847 -1
rect 1849 -5 1850 -1
rect 1867 -5 1868 -1
rect 1870 -5 1871 -1
rect 1883 -5 1884 -1
rect 1886 -5 1887 -1
rect 1899 -5 1900 -1
rect 1902 -5 1905 -1
rect 1907 -5 1908 -1
rect 1920 -5 1921 -1
rect 1923 -5 1924 -1
rect 100 -35 101 -31
rect 103 -35 106 -31
rect 108 -35 109 -31
rect 121 -35 122 -31
rect 124 -35 125 -31
rect 137 -35 138 -31
rect 140 -35 143 -31
rect 145 -35 146 -31
rect 163 -35 164 -31
rect 166 -35 167 -31
rect 179 -35 180 -31
rect 182 -35 183 -31
rect 195 -35 196 -31
rect 198 -35 201 -31
rect 203 -35 204 -31
rect 216 -35 217 -31
rect 219 -35 220 -31
rect 232 -35 233 -31
rect 235 -35 238 -31
rect 240 -35 241 -31
rect 253 -35 254 -31
rect 256 -35 257 -31
rect 269 -35 270 -31
rect 272 -35 275 -31
rect 277 -35 278 -31
rect 295 -35 296 -31
rect 298 -35 299 -31
rect 311 -35 312 -31
rect 314 -35 315 -31
rect 327 -35 328 -31
rect 330 -35 333 -31
rect 335 -35 336 -31
rect 348 -35 349 -31
rect 351 -35 352 -31
rect 364 -35 365 -31
rect 367 -35 370 -31
rect 372 -35 373 -31
rect 385 -35 386 -31
rect 388 -35 389 -31
rect 401 -35 402 -31
rect 404 -35 407 -31
rect 409 -35 410 -31
rect 427 -35 428 -31
rect 430 -35 431 -31
rect 443 -35 444 -31
rect 446 -35 447 -31
rect 459 -35 460 -31
rect 462 -35 465 -31
rect 467 -35 468 -31
rect 480 -35 481 -31
rect 483 -35 484 -31
rect 1033 -35 1034 -31
rect 1036 -35 1039 -31
rect 1041 -35 1042 -31
rect 1054 -35 1055 -31
rect 1057 -35 1058 -31
rect 1070 -35 1071 -31
rect 1073 -35 1076 -31
rect 1078 -35 1079 -31
rect 1096 -35 1097 -31
rect 1099 -35 1100 -31
rect 1112 -35 1113 -31
rect 1115 -35 1116 -31
rect 1128 -35 1129 -31
rect 1131 -35 1134 -31
rect 1136 -35 1137 -31
rect 1149 -35 1150 -31
rect 1152 -35 1153 -31
rect 1165 -35 1166 -31
rect 1168 -35 1171 -31
rect 1173 -35 1174 -31
rect 1186 -35 1187 -31
rect 1189 -35 1190 -31
rect 1202 -35 1203 -31
rect 1205 -35 1208 -31
rect 1210 -35 1211 -31
rect 1228 -35 1229 -31
rect 1231 -35 1232 -31
rect 1244 -35 1245 -31
rect 1247 -35 1248 -31
rect 1260 -35 1261 -31
rect 1263 -35 1266 -31
rect 1268 -35 1269 -31
rect 1281 -35 1282 -31
rect 1284 -35 1285 -31
rect 1297 -35 1298 -31
rect 1300 -35 1303 -31
rect 1305 -35 1306 -31
rect 1318 -35 1319 -31
rect 1321 -35 1322 -31
rect 1334 -35 1335 -31
rect 1337 -35 1340 -31
rect 1342 -35 1343 -31
rect 1360 -35 1361 -31
rect 1363 -35 1364 -31
rect 1376 -35 1377 -31
rect 1379 -35 1380 -31
rect 1392 -35 1393 -31
rect 1395 -35 1398 -31
rect 1400 -35 1401 -31
rect 1413 -35 1414 -31
rect 1416 -35 1417 -31
rect 332 -79 333 -75
rect 335 -79 336 -75
rect 356 -79 357 -75
rect 359 -79 360 -75
rect 1265 -79 1266 -75
rect 1268 -79 1269 -75
rect 1289 -79 1290 -75
rect 1292 -79 1293 -75
rect 352 -90 353 -86
rect 355 -90 356 -86
rect 1285 -90 1286 -86
rect 1288 -90 1289 -86
rect 344 -102 348 -101
rect 344 -105 348 -104
rect 1277 -102 1281 -101
rect 1277 -105 1281 -104
rect 332 -113 333 -109
rect 335 -113 336 -109
rect 356 -113 357 -109
rect 359 -113 360 -109
rect 1265 -113 1266 -109
rect 1268 -113 1269 -109
rect 1289 -113 1290 -109
rect 1292 -113 1293 -109
rect 100 -175 101 -171
rect 103 -175 106 -171
rect 108 -175 109 -171
rect 121 -175 122 -171
rect 124 -175 125 -171
rect 137 -175 138 -171
rect 140 -175 143 -171
rect 145 -175 146 -171
rect 163 -175 164 -171
rect 166 -175 167 -171
rect 179 -175 180 -171
rect 182 -175 183 -171
rect 195 -175 196 -171
rect 198 -175 201 -171
rect 203 -175 204 -171
rect 216 -175 217 -171
rect 219 -175 220 -171
rect 232 -175 233 -171
rect 235 -175 238 -171
rect 240 -175 241 -171
rect 253 -175 254 -171
rect 256 -175 257 -171
rect 269 -175 270 -171
rect 272 -175 275 -171
rect 277 -175 278 -171
rect 295 -175 296 -171
rect 298 -175 299 -171
rect 311 -175 312 -171
rect 314 -175 315 -171
rect 327 -175 328 -171
rect 330 -175 333 -171
rect 335 -175 336 -171
rect 348 -175 349 -171
rect 351 -175 352 -171
rect 364 -175 365 -171
rect 367 -175 370 -171
rect 372 -175 373 -171
rect 385 -175 386 -171
rect 388 -175 389 -171
rect 401 -175 402 -171
rect 404 -175 407 -171
rect 409 -175 410 -171
rect 427 -175 428 -171
rect 430 -175 431 -171
rect 443 -175 444 -171
rect 446 -175 447 -171
rect 459 -175 460 -171
rect 462 -175 465 -171
rect 467 -175 468 -171
rect 480 -175 481 -171
rect 483 -175 484 -171
rect 1033 -175 1034 -171
rect 1036 -175 1039 -171
rect 1041 -175 1042 -171
rect 1054 -175 1055 -171
rect 1057 -175 1058 -171
rect 1070 -175 1071 -171
rect 1073 -175 1076 -171
rect 1078 -175 1079 -171
rect 1096 -175 1097 -171
rect 1099 -175 1100 -171
rect 1112 -175 1113 -171
rect 1115 -175 1116 -171
rect 1128 -175 1129 -171
rect 1131 -175 1134 -171
rect 1136 -175 1137 -171
rect 1149 -175 1150 -171
rect 1152 -175 1153 -171
rect 1165 -175 1166 -171
rect 1168 -175 1171 -171
rect 1173 -175 1174 -171
rect 1186 -175 1187 -171
rect 1189 -175 1190 -171
rect 1202 -175 1203 -171
rect 1205 -175 1208 -171
rect 1210 -175 1211 -171
rect 1228 -175 1229 -171
rect 1231 -175 1232 -171
rect 1244 -175 1245 -171
rect 1247 -175 1248 -171
rect 1260 -175 1261 -171
rect 1263 -175 1266 -171
rect 1268 -175 1269 -171
rect 1281 -175 1282 -171
rect 1284 -175 1285 -171
rect 1297 -175 1298 -171
rect 1300 -175 1303 -171
rect 1305 -175 1306 -171
rect 1318 -175 1319 -171
rect 1321 -175 1322 -171
rect 1334 -175 1335 -171
rect 1337 -175 1340 -171
rect 1342 -175 1343 -171
rect 1360 -175 1361 -171
rect 1363 -175 1364 -171
rect 1376 -175 1377 -171
rect 1379 -175 1380 -171
rect 1392 -175 1393 -171
rect 1395 -175 1398 -171
rect 1400 -175 1401 -171
rect 1413 -175 1414 -171
rect 1416 -175 1417 -171
<< pdiffusion >>
rect 572 1729 573 1737
rect 575 1729 578 1737
rect 580 1729 581 1737
rect 593 1729 594 1737
rect 596 1733 597 1737
rect 596 1729 601 1733
rect 609 1729 610 1737
rect 612 1729 615 1737
rect 617 1729 618 1737
rect 635 1729 636 1737
rect 638 1729 639 1737
rect 651 1729 652 1737
rect 654 1733 655 1737
rect 654 1729 659 1733
rect 667 1729 668 1737
rect 670 1729 673 1737
rect 675 1729 676 1737
rect 688 1729 689 1737
rect 691 1729 692 1737
rect 704 1729 705 1737
rect 707 1729 710 1737
rect 712 1729 713 1737
rect 725 1729 726 1737
rect 728 1733 729 1737
rect 728 1729 733 1733
rect 741 1729 742 1737
rect 744 1729 747 1737
rect 749 1729 750 1737
rect 767 1729 768 1737
rect 770 1729 771 1737
rect 783 1729 784 1737
rect 786 1733 787 1737
rect 786 1729 791 1733
rect 799 1729 800 1737
rect 802 1729 805 1737
rect 807 1729 808 1737
rect 820 1729 821 1737
rect 823 1729 824 1737
rect 836 1729 837 1737
rect 839 1729 842 1737
rect 844 1729 845 1737
rect 857 1729 858 1737
rect 860 1733 861 1737
rect 860 1729 865 1733
rect 873 1729 874 1737
rect 876 1729 879 1737
rect 881 1729 882 1737
rect 899 1729 900 1737
rect 902 1729 903 1737
rect 915 1729 916 1737
rect 918 1733 919 1737
rect 918 1729 923 1733
rect 931 1729 932 1737
rect 934 1729 937 1737
rect 939 1729 940 1737
rect 952 1729 953 1737
rect 955 1729 956 1737
rect 968 1729 969 1737
rect 971 1729 974 1737
rect 976 1729 977 1737
rect 989 1729 990 1737
rect 992 1733 993 1737
rect 992 1729 997 1733
rect 1005 1729 1006 1737
rect 1008 1729 1011 1737
rect 1013 1729 1014 1737
rect 1031 1729 1032 1737
rect 1034 1729 1035 1737
rect 1047 1729 1048 1737
rect 1050 1733 1051 1737
rect 1050 1729 1055 1733
rect 1063 1729 1064 1737
rect 1066 1729 1069 1737
rect 1071 1729 1072 1737
rect 1084 1729 1085 1737
rect 1087 1729 1088 1737
rect 1505 1729 1506 1737
rect 1508 1729 1511 1737
rect 1513 1729 1514 1737
rect 1526 1729 1527 1737
rect 1529 1733 1530 1737
rect 1529 1729 1534 1733
rect 1542 1729 1543 1737
rect 1545 1729 1548 1737
rect 1550 1729 1551 1737
rect 1568 1729 1569 1737
rect 1571 1729 1572 1737
rect 1584 1729 1585 1737
rect 1587 1733 1588 1737
rect 1587 1729 1592 1733
rect 1600 1729 1601 1737
rect 1603 1729 1606 1737
rect 1608 1729 1609 1737
rect 1621 1729 1622 1737
rect 1624 1729 1625 1737
rect 1637 1729 1638 1737
rect 1640 1729 1643 1737
rect 1645 1729 1646 1737
rect 1658 1729 1659 1737
rect 1661 1733 1662 1737
rect 1661 1729 1666 1733
rect 1674 1729 1675 1737
rect 1677 1729 1680 1737
rect 1682 1729 1683 1737
rect 1700 1729 1701 1737
rect 1703 1729 1704 1737
rect 1716 1729 1717 1737
rect 1719 1733 1720 1737
rect 1719 1729 1724 1733
rect 1732 1729 1733 1737
rect 1735 1729 1738 1737
rect 1740 1729 1741 1737
rect 1753 1729 1754 1737
rect 1756 1729 1757 1737
rect 1769 1729 1770 1737
rect 1772 1729 1775 1737
rect 1777 1729 1778 1737
rect 1790 1729 1791 1737
rect 1793 1733 1794 1737
rect 1793 1729 1798 1733
rect 1806 1729 1807 1737
rect 1809 1729 1812 1737
rect 1814 1729 1815 1737
rect 1832 1729 1833 1737
rect 1835 1729 1836 1737
rect 1848 1729 1849 1737
rect 1851 1733 1852 1737
rect 1851 1729 1856 1733
rect 1864 1729 1865 1737
rect 1867 1729 1870 1737
rect 1872 1729 1873 1737
rect 1885 1729 1886 1737
rect 1888 1729 1889 1737
rect 1901 1729 1902 1737
rect 1904 1729 1907 1737
rect 1909 1729 1910 1737
rect 1922 1729 1923 1737
rect 1925 1733 1926 1737
rect 1925 1729 1930 1733
rect 1938 1729 1939 1737
rect 1941 1729 1944 1737
rect 1946 1729 1947 1737
rect 1964 1729 1965 1737
rect 1967 1729 1968 1737
rect 1980 1729 1981 1737
rect 1983 1733 1984 1737
rect 1983 1729 1988 1733
rect 1996 1729 1997 1737
rect 1999 1729 2002 1737
rect 2004 1729 2005 1737
rect 2017 1729 2018 1737
rect 2020 1729 2021 1737
rect 232 1696 233 1704
rect 235 1696 238 1704
rect 240 1696 241 1704
rect 253 1696 254 1704
rect 256 1700 257 1704
rect 256 1696 261 1700
rect 269 1696 270 1704
rect 272 1696 275 1704
rect 277 1696 278 1704
rect 295 1696 296 1704
rect 298 1696 299 1704
rect 311 1696 312 1704
rect 314 1700 315 1704
rect 314 1696 319 1700
rect 327 1696 328 1704
rect 330 1696 333 1704
rect 335 1696 336 1704
rect 348 1696 349 1704
rect 351 1696 352 1704
rect 1165 1696 1166 1704
rect 1168 1696 1171 1704
rect 1173 1696 1174 1704
rect 1186 1696 1187 1704
rect 1189 1700 1190 1704
rect 1189 1696 1194 1700
rect 1202 1696 1203 1704
rect 1205 1696 1208 1704
rect 1210 1696 1211 1704
rect 1228 1696 1229 1704
rect 1231 1696 1232 1704
rect 1244 1696 1245 1704
rect 1247 1700 1248 1704
rect 1247 1696 1252 1700
rect 1260 1696 1261 1704
rect 1263 1696 1266 1704
rect 1268 1696 1269 1704
rect 1281 1696 1282 1704
rect 1284 1696 1285 1704
rect 751 1658 752 1666
rect 754 1658 755 1666
rect 577 1645 578 1653
rect 580 1645 581 1653
rect 593 1645 594 1653
rect 596 1645 597 1653
rect 609 1645 610 1653
rect 612 1645 613 1653
rect 628 1645 633 1653
rect 635 1645 638 1653
rect 640 1645 641 1653
rect 662 1645 664 1653
rect 666 1645 667 1653
rect 684 1645 685 1653
rect 687 1645 688 1653
rect 700 1645 705 1653
rect 707 1645 710 1653
rect 712 1645 713 1653
rect 727 1645 728 1653
rect 730 1645 731 1653
rect 775 1652 778 1660
rect 780 1652 783 1660
rect 785 1652 786 1660
rect 805 1658 806 1666
rect 808 1658 809 1666
rect 832 1658 833 1666
rect 835 1658 836 1666
rect 856 1652 859 1660
rect 861 1652 864 1660
rect 866 1652 867 1660
rect 886 1658 887 1666
rect 889 1658 890 1666
rect 1684 1658 1685 1666
rect 1687 1658 1688 1666
rect 1510 1645 1511 1653
rect 1513 1645 1514 1653
rect 1526 1645 1527 1653
rect 1529 1645 1530 1653
rect 1542 1645 1543 1653
rect 1545 1645 1546 1653
rect 1561 1645 1566 1653
rect 1568 1645 1571 1653
rect 1573 1645 1574 1653
rect 1595 1645 1597 1653
rect 1599 1645 1600 1653
rect 1617 1645 1618 1653
rect 1620 1645 1621 1653
rect 1633 1645 1638 1653
rect 1640 1645 1643 1653
rect 1645 1645 1646 1653
rect 1660 1645 1661 1653
rect 1663 1645 1664 1653
rect 1708 1652 1711 1660
rect 1713 1652 1716 1660
rect 1718 1652 1719 1660
rect 1738 1658 1739 1666
rect 1741 1658 1742 1666
rect 1765 1658 1766 1666
rect 1768 1658 1769 1666
rect 1789 1652 1792 1660
rect 1794 1652 1797 1660
rect 1799 1652 1800 1660
rect 1819 1658 1820 1666
rect 1822 1658 1823 1666
rect 223 1594 224 1602
rect 226 1594 227 1602
rect 239 1594 240 1602
rect 242 1594 245 1602
rect 247 1594 248 1602
rect 260 1598 261 1602
rect 256 1594 261 1598
rect 263 1594 264 1602
rect 276 1594 277 1602
rect 279 1594 280 1602
rect 297 1594 298 1602
rect 300 1594 303 1602
rect 305 1594 306 1602
rect 318 1598 319 1602
rect 314 1594 319 1598
rect 321 1594 322 1602
rect 334 1594 335 1602
rect 337 1594 340 1602
rect 342 1594 343 1602
rect 1156 1594 1157 1602
rect 1159 1594 1160 1602
rect 1172 1594 1173 1602
rect 1175 1594 1178 1602
rect 1180 1594 1181 1602
rect 1193 1598 1194 1602
rect 1189 1594 1194 1598
rect 1196 1594 1197 1602
rect 1209 1594 1210 1602
rect 1212 1594 1213 1602
rect 1230 1594 1231 1602
rect 1233 1594 1236 1602
rect 1238 1594 1239 1602
rect 1251 1598 1252 1602
rect 1247 1594 1252 1598
rect 1254 1594 1255 1602
rect 1267 1594 1268 1602
rect 1270 1594 1273 1602
rect 1275 1594 1276 1602
rect 577 1559 578 1567
rect 580 1559 581 1567
rect 593 1559 594 1567
rect 596 1559 597 1567
rect 609 1559 610 1567
rect 612 1559 613 1567
rect 628 1559 633 1567
rect 635 1559 638 1567
rect 640 1559 641 1567
rect 662 1559 664 1567
rect 666 1559 667 1567
rect 684 1559 685 1567
rect 687 1559 688 1567
rect 700 1559 705 1567
rect 707 1559 710 1567
rect 712 1559 713 1567
rect 727 1559 728 1567
rect 730 1559 731 1567
rect 775 1560 778 1568
rect 780 1560 783 1568
rect 785 1560 786 1568
rect 856 1560 859 1568
rect 861 1560 864 1568
rect 866 1560 867 1568
rect 1510 1559 1511 1567
rect 1513 1559 1514 1567
rect 1526 1559 1527 1567
rect 1529 1559 1530 1567
rect 1542 1559 1543 1567
rect 1545 1559 1546 1567
rect 1561 1559 1566 1567
rect 1568 1559 1571 1567
rect 1573 1559 1574 1567
rect 1595 1559 1597 1567
rect 1599 1559 1600 1567
rect 1617 1559 1618 1567
rect 1620 1559 1621 1567
rect 1633 1559 1638 1567
rect 1640 1559 1643 1567
rect 1645 1559 1646 1567
rect 1660 1559 1661 1567
rect 1663 1559 1664 1567
rect 1708 1560 1711 1568
rect 1713 1560 1716 1568
rect 1718 1560 1719 1568
rect 1789 1560 1792 1568
rect 1794 1560 1797 1568
rect 1799 1560 1800 1568
rect 577 1513 578 1521
rect 580 1513 581 1521
rect 593 1513 594 1521
rect 596 1513 597 1521
rect 609 1513 610 1521
rect 612 1513 613 1521
rect 628 1513 633 1521
rect 635 1513 638 1521
rect 640 1513 641 1521
rect 662 1513 664 1521
rect 666 1513 667 1521
rect 684 1513 685 1521
rect 687 1513 688 1521
rect 700 1513 705 1521
rect 707 1513 710 1521
rect 712 1513 713 1521
rect 727 1513 728 1521
rect 730 1513 731 1521
rect 775 1520 778 1528
rect 780 1520 783 1528
rect 785 1520 786 1528
rect 805 1526 806 1534
rect 808 1526 809 1534
rect 856 1526 857 1534
rect 859 1526 860 1534
rect 880 1520 883 1528
rect 885 1520 888 1528
rect 890 1520 891 1528
rect 910 1526 911 1534
rect 913 1526 914 1534
rect 1510 1513 1511 1521
rect 1513 1513 1514 1521
rect 1526 1513 1527 1521
rect 1529 1513 1530 1521
rect 1542 1513 1543 1521
rect 1545 1513 1546 1521
rect 1561 1513 1566 1521
rect 1568 1513 1571 1521
rect 1573 1513 1574 1521
rect 1595 1513 1597 1521
rect 1599 1513 1600 1521
rect 1617 1513 1618 1521
rect 1620 1513 1621 1521
rect 1633 1513 1638 1521
rect 1640 1513 1643 1521
rect 1645 1513 1646 1521
rect 1660 1513 1661 1521
rect 1663 1513 1664 1521
rect 1708 1520 1711 1528
rect 1713 1520 1716 1528
rect 1718 1520 1719 1528
rect 1738 1526 1739 1534
rect 1741 1526 1742 1534
rect 1789 1526 1790 1534
rect 1792 1526 1793 1534
rect 1813 1520 1816 1528
rect 1818 1520 1821 1528
rect 1823 1520 1824 1528
rect 1843 1526 1844 1534
rect 1846 1526 1847 1534
rect 577 1427 578 1435
rect 580 1427 581 1435
rect 593 1427 594 1435
rect 596 1427 597 1435
rect 609 1427 610 1435
rect 612 1427 613 1435
rect 628 1427 633 1435
rect 635 1427 638 1435
rect 640 1427 641 1435
rect 662 1427 664 1435
rect 666 1427 667 1435
rect 684 1427 685 1435
rect 687 1427 688 1435
rect 700 1427 705 1435
rect 707 1427 710 1435
rect 712 1427 713 1435
rect 727 1427 728 1435
rect 730 1427 731 1435
rect 775 1429 778 1437
rect 780 1429 783 1437
rect 785 1429 786 1437
rect 880 1429 883 1437
rect 885 1429 888 1437
rect 890 1429 891 1437
rect 1510 1427 1511 1435
rect 1513 1427 1514 1435
rect 1526 1427 1527 1435
rect 1529 1427 1530 1435
rect 1542 1427 1543 1435
rect 1545 1427 1546 1435
rect 1561 1427 1566 1435
rect 1568 1427 1571 1435
rect 1573 1427 1574 1435
rect 1595 1427 1597 1435
rect 1599 1427 1600 1435
rect 1617 1427 1618 1435
rect 1620 1427 1621 1435
rect 1633 1427 1638 1435
rect 1640 1427 1643 1435
rect 1645 1427 1646 1435
rect 1660 1427 1661 1435
rect 1663 1427 1664 1435
rect 1708 1429 1711 1437
rect 1713 1429 1716 1437
rect 1718 1429 1719 1437
rect 1813 1429 1816 1437
rect 1818 1429 1821 1437
rect 1823 1429 1824 1437
rect 577 1381 578 1389
rect 580 1381 581 1389
rect 593 1381 594 1389
rect 596 1381 597 1389
rect 609 1381 610 1389
rect 612 1381 613 1389
rect 628 1381 633 1389
rect 635 1381 638 1389
rect 640 1381 641 1389
rect 662 1381 664 1389
rect 666 1381 667 1389
rect 684 1381 685 1389
rect 687 1381 688 1389
rect 700 1381 705 1389
rect 707 1381 710 1389
rect 712 1381 713 1389
rect 727 1381 728 1389
rect 730 1381 731 1389
rect 775 1388 778 1396
rect 780 1388 783 1396
rect 785 1388 786 1396
rect 805 1394 806 1402
rect 808 1394 809 1402
rect 832 1394 833 1402
rect 835 1394 836 1402
rect 856 1388 859 1396
rect 861 1388 864 1396
rect 866 1388 867 1396
rect 886 1394 887 1402
rect 889 1394 890 1402
rect 922 1394 923 1402
rect 925 1394 926 1402
rect 946 1388 949 1396
rect 951 1388 954 1396
rect 956 1388 957 1396
rect 976 1394 977 1402
rect 979 1394 980 1402
rect 1510 1381 1511 1389
rect 1513 1381 1514 1389
rect 1526 1381 1527 1389
rect 1529 1381 1530 1389
rect 1542 1381 1543 1389
rect 1545 1381 1546 1389
rect 1561 1381 1566 1389
rect 1568 1381 1571 1389
rect 1573 1381 1574 1389
rect 1595 1381 1597 1389
rect 1599 1381 1600 1389
rect 1617 1381 1618 1389
rect 1620 1381 1621 1389
rect 1633 1381 1638 1389
rect 1640 1381 1643 1389
rect 1645 1381 1646 1389
rect 1660 1381 1661 1389
rect 1663 1381 1664 1389
rect 1708 1388 1711 1396
rect 1713 1388 1716 1396
rect 1718 1388 1719 1396
rect 1738 1394 1739 1402
rect 1741 1394 1742 1402
rect 1765 1394 1766 1402
rect 1768 1394 1769 1402
rect 1789 1388 1792 1396
rect 1794 1388 1797 1396
rect 1799 1388 1800 1396
rect 1819 1394 1820 1402
rect 1822 1394 1823 1402
rect 1855 1394 1856 1402
rect 1858 1394 1859 1402
rect 1879 1388 1882 1396
rect 1884 1388 1887 1396
rect 1889 1388 1890 1396
rect 1909 1394 1910 1402
rect 1912 1394 1913 1402
rect 577 1295 578 1303
rect 580 1295 581 1303
rect 593 1295 594 1303
rect 596 1295 597 1303
rect 609 1295 610 1303
rect 612 1295 613 1303
rect 628 1295 633 1303
rect 635 1295 638 1303
rect 640 1295 641 1303
rect 662 1295 664 1303
rect 666 1295 667 1303
rect 684 1295 685 1303
rect 687 1295 688 1303
rect 700 1295 705 1303
rect 707 1295 710 1303
rect 712 1295 713 1303
rect 727 1295 728 1303
rect 730 1295 731 1303
rect 775 1294 778 1302
rect 780 1294 783 1302
rect 785 1294 786 1302
rect 856 1294 859 1302
rect 861 1294 864 1302
rect 866 1294 867 1302
rect 946 1294 949 1302
rect 951 1294 954 1302
rect 956 1294 957 1302
rect 1510 1295 1511 1303
rect 1513 1295 1514 1303
rect 1526 1295 1527 1303
rect 1529 1295 1530 1303
rect 1542 1295 1543 1303
rect 1545 1295 1546 1303
rect 1561 1295 1566 1303
rect 1568 1295 1571 1303
rect 1573 1295 1574 1303
rect 1595 1295 1597 1303
rect 1599 1295 1600 1303
rect 1617 1295 1618 1303
rect 1620 1295 1621 1303
rect 1633 1295 1638 1303
rect 1640 1295 1643 1303
rect 1645 1295 1646 1303
rect 1660 1295 1661 1303
rect 1663 1295 1664 1303
rect 1708 1294 1711 1302
rect 1713 1294 1716 1302
rect 1718 1294 1719 1302
rect 1789 1294 1792 1302
rect 1794 1294 1797 1302
rect 1799 1294 1800 1302
rect 1879 1294 1882 1302
rect 1884 1294 1887 1302
rect 1889 1294 1890 1302
rect 577 1249 578 1257
rect 580 1249 581 1257
rect 593 1249 594 1257
rect 596 1249 597 1257
rect 609 1249 610 1257
rect 612 1249 613 1257
rect 628 1249 633 1257
rect 635 1249 638 1257
rect 640 1249 641 1257
rect 662 1249 664 1257
rect 666 1249 667 1257
rect 684 1249 685 1257
rect 687 1249 688 1257
rect 700 1249 705 1257
rect 707 1249 710 1257
rect 712 1249 713 1257
rect 727 1249 728 1257
rect 730 1249 731 1257
rect 775 1256 778 1264
rect 780 1256 783 1264
rect 785 1256 786 1264
rect 805 1262 806 1270
rect 808 1262 809 1270
rect 1510 1249 1511 1257
rect 1513 1249 1514 1257
rect 1526 1249 1527 1257
rect 1529 1249 1530 1257
rect 1542 1249 1543 1257
rect 1545 1249 1546 1257
rect 1561 1249 1566 1257
rect 1568 1249 1571 1257
rect 1573 1249 1574 1257
rect 1595 1249 1597 1257
rect 1599 1249 1600 1257
rect 1617 1249 1618 1257
rect 1620 1249 1621 1257
rect 1633 1249 1638 1257
rect 1640 1249 1643 1257
rect 1645 1249 1646 1257
rect 1660 1249 1661 1257
rect 1663 1249 1664 1257
rect 1708 1256 1711 1264
rect 1713 1256 1716 1264
rect 1718 1256 1719 1264
rect 1738 1262 1739 1270
rect 1741 1262 1742 1270
rect 100 1194 101 1202
rect 103 1194 106 1202
rect 108 1194 109 1202
rect 121 1194 122 1202
rect 124 1198 125 1202
rect 124 1194 129 1198
rect 137 1194 138 1202
rect 140 1194 143 1202
rect 145 1194 146 1202
rect 163 1194 164 1202
rect 166 1194 167 1202
rect 179 1194 180 1202
rect 182 1198 183 1202
rect 182 1194 187 1198
rect 195 1194 196 1202
rect 198 1194 201 1202
rect 203 1194 204 1202
rect 216 1194 217 1202
rect 219 1194 220 1202
rect 232 1194 233 1202
rect 235 1194 238 1202
rect 240 1194 241 1202
rect 253 1194 254 1202
rect 256 1198 257 1202
rect 256 1194 261 1198
rect 269 1194 270 1202
rect 272 1194 275 1202
rect 277 1194 278 1202
rect 295 1194 296 1202
rect 298 1194 299 1202
rect 311 1194 312 1202
rect 314 1198 315 1202
rect 314 1194 319 1198
rect 327 1194 328 1202
rect 330 1194 333 1202
rect 335 1194 336 1202
rect 348 1194 349 1202
rect 351 1194 352 1202
rect 364 1194 365 1202
rect 367 1194 370 1202
rect 372 1194 373 1202
rect 385 1194 386 1202
rect 388 1198 389 1202
rect 388 1194 393 1198
rect 401 1194 402 1202
rect 404 1194 407 1202
rect 409 1194 410 1202
rect 427 1194 428 1202
rect 430 1194 431 1202
rect 443 1194 444 1202
rect 446 1198 447 1202
rect 446 1194 451 1198
rect 459 1194 460 1202
rect 462 1194 465 1202
rect 467 1194 468 1202
rect 480 1194 481 1202
rect 483 1194 484 1202
rect 1033 1194 1034 1202
rect 1036 1194 1039 1202
rect 1041 1194 1042 1202
rect 1054 1194 1055 1202
rect 1057 1198 1058 1202
rect 1057 1194 1062 1198
rect 1070 1194 1071 1202
rect 1073 1194 1076 1202
rect 1078 1194 1079 1202
rect 1096 1194 1097 1202
rect 1099 1194 1100 1202
rect 1112 1194 1113 1202
rect 1115 1198 1116 1202
rect 1115 1194 1120 1198
rect 1128 1194 1129 1202
rect 1131 1194 1134 1202
rect 1136 1194 1137 1202
rect 1149 1194 1150 1202
rect 1152 1194 1153 1202
rect 1165 1194 1166 1202
rect 1168 1194 1171 1202
rect 1173 1194 1174 1202
rect 1186 1194 1187 1202
rect 1189 1198 1190 1202
rect 1189 1194 1194 1198
rect 1202 1194 1203 1202
rect 1205 1194 1208 1202
rect 1210 1194 1211 1202
rect 1228 1194 1229 1202
rect 1231 1194 1232 1202
rect 1244 1194 1245 1202
rect 1247 1198 1248 1202
rect 1247 1194 1252 1198
rect 1260 1194 1261 1202
rect 1263 1194 1266 1202
rect 1268 1194 1269 1202
rect 1281 1194 1282 1202
rect 1284 1194 1285 1202
rect 1297 1194 1298 1202
rect 1300 1194 1303 1202
rect 1305 1194 1306 1202
rect 1318 1194 1319 1202
rect 1321 1198 1322 1202
rect 1321 1194 1326 1198
rect 1334 1194 1335 1202
rect 1337 1194 1340 1202
rect 1342 1194 1343 1202
rect 1360 1194 1361 1202
rect 1363 1194 1364 1202
rect 1376 1194 1377 1202
rect 1379 1198 1380 1202
rect 1379 1194 1384 1198
rect 1392 1194 1393 1202
rect 1395 1194 1398 1202
rect 1400 1194 1401 1202
rect 1413 1194 1414 1202
rect 1416 1194 1417 1202
rect 577 1163 578 1171
rect 580 1163 581 1171
rect 593 1163 594 1171
rect 596 1163 597 1171
rect 609 1163 610 1171
rect 612 1163 613 1171
rect 628 1163 633 1171
rect 635 1163 638 1171
rect 640 1163 641 1171
rect 662 1163 664 1171
rect 666 1163 667 1171
rect 684 1163 685 1171
rect 687 1163 688 1171
rect 700 1163 705 1171
rect 707 1163 710 1171
rect 712 1163 713 1171
rect 727 1163 728 1171
rect 730 1163 731 1171
rect 775 1158 778 1166
rect 780 1158 783 1166
rect 785 1158 786 1166
rect 811 1163 812 1171
rect 814 1163 815 1171
rect 819 1163 825 1171
rect 829 1163 830 1171
rect 832 1163 833 1171
rect 854 1163 855 1171
rect 857 1163 858 1171
rect 870 1163 871 1171
rect 873 1163 874 1171
rect 889 1163 894 1171
rect 896 1163 899 1171
rect 901 1163 902 1171
rect 923 1163 925 1171
rect 927 1163 928 1171
rect 945 1163 946 1171
rect 948 1163 949 1171
rect 961 1163 966 1171
rect 968 1163 971 1171
rect 973 1163 974 1171
rect 988 1163 989 1171
rect 991 1163 992 1171
rect 1510 1163 1511 1171
rect 1513 1163 1514 1171
rect 1526 1163 1527 1171
rect 1529 1163 1530 1171
rect 1542 1163 1543 1171
rect 1545 1163 1546 1171
rect 1561 1163 1566 1171
rect 1568 1163 1571 1171
rect 1573 1163 1574 1171
rect 1595 1163 1597 1171
rect 1599 1163 1600 1171
rect 1617 1163 1618 1171
rect 1620 1163 1621 1171
rect 1633 1163 1638 1171
rect 1640 1163 1643 1171
rect 1645 1163 1646 1171
rect 1660 1163 1661 1171
rect 1663 1163 1664 1171
rect 1708 1158 1711 1166
rect 1713 1158 1716 1166
rect 1718 1158 1719 1166
rect 1744 1163 1745 1171
rect 1747 1163 1748 1171
rect 1752 1163 1758 1171
rect 1762 1163 1763 1171
rect 1765 1163 1766 1171
rect 1787 1163 1788 1171
rect 1790 1163 1791 1171
rect 1803 1163 1804 1171
rect 1806 1163 1807 1171
rect 1822 1163 1827 1171
rect 1829 1163 1832 1171
rect 1834 1163 1835 1171
rect 1856 1163 1858 1171
rect 1860 1163 1861 1171
rect 1878 1163 1879 1171
rect 1881 1163 1882 1171
rect 1894 1163 1899 1171
rect 1901 1163 1904 1171
rect 1906 1163 1907 1171
rect 1921 1163 1922 1171
rect 1924 1163 1925 1171
rect 871 1084 872 1092
rect 874 1084 877 1092
rect 879 1084 880 1092
rect 892 1084 893 1092
rect 895 1088 896 1092
rect 895 1084 900 1088
rect 908 1084 909 1092
rect 911 1084 914 1092
rect 916 1084 917 1092
rect 934 1084 935 1092
rect 937 1084 938 1092
rect 950 1084 951 1092
rect 953 1088 954 1092
rect 953 1084 958 1088
rect 966 1084 967 1092
rect 969 1084 972 1092
rect 974 1084 975 1092
rect 987 1084 988 1092
rect 990 1084 991 1092
rect 1804 1084 1805 1092
rect 1807 1084 1810 1092
rect 1812 1084 1813 1092
rect 1825 1084 1826 1092
rect 1828 1088 1829 1092
rect 1828 1084 1833 1088
rect 1841 1084 1842 1092
rect 1844 1084 1847 1092
rect 1849 1084 1850 1092
rect 1867 1084 1868 1092
rect 1870 1084 1871 1092
rect 1883 1084 1884 1092
rect 1886 1088 1887 1092
rect 1886 1084 1891 1088
rect 1899 1084 1900 1092
rect 1902 1084 1905 1092
rect 1907 1084 1908 1092
rect 1920 1084 1921 1092
rect 1923 1084 1924 1092
rect 100 1054 101 1062
rect 103 1054 106 1062
rect 108 1054 109 1062
rect 121 1054 122 1062
rect 124 1058 125 1062
rect 124 1054 129 1058
rect 137 1054 138 1062
rect 140 1054 143 1062
rect 145 1054 146 1062
rect 163 1054 164 1062
rect 166 1054 167 1062
rect 179 1054 180 1062
rect 182 1058 183 1062
rect 182 1054 187 1058
rect 195 1054 196 1062
rect 198 1054 201 1062
rect 203 1054 204 1062
rect 216 1054 217 1062
rect 219 1054 220 1062
rect 232 1054 233 1062
rect 235 1054 238 1062
rect 240 1054 241 1062
rect 253 1054 254 1062
rect 256 1058 257 1062
rect 256 1054 261 1058
rect 269 1054 270 1062
rect 272 1054 275 1062
rect 277 1054 278 1062
rect 295 1054 296 1062
rect 298 1054 299 1062
rect 311 1054 312 1062
rect 314 1058 315 1062
rect 314 1054 319 1058
rect 327 1054 328 1062
rect 330 1054 333 1062
rect 335 1054 336 1062
rect 348 1054 349 1062
rect 351 1054 352 1062
rect 364 1054 365 1062
rect 367 1054 370 1062
rect 372 1054 373 1062
rect 385 1054 386 1062
rect 388 1058 389 1062
rect 388 1054 393 1058
rect 401 1054 402 1062
rect 404 1054 407 1062
rect 409 1054 410 1062
rect 427 1054 428 1062
rect 430 1054 431 1062
rect 443 1054 444 1062
rect 446 1058 447 1062
rect 446 1054 451 1058
rect 459 1054 460 1062
rect 462 1054 465 1062
rect 467 1054 468 1062
rect 480 1054 481 1062
rect 483 1054 484 1062
rect 1033 1054 1034 1062
rect 1036 1054 1039 1062
rect 1041 1054 1042 1062
rect 1054 1054 1055 1062
rect 1057 1058 1058 1062
rect 1057 1054 1062 1058
rect 1070 1054 1071 1062
rect 1073 1054 1076 1062
rect 1078 1054 1079 1062
rect 1096 1054 1097 1062
rect 1099 1054 1100 1062
rect 1112 1054 1113 1062
rect 1115 1058 1116 1062
rect 1115 1054 1120 1058
rect 1128 1054 1129 1062
rect 1131 1054 1134 1062
rect 1136 1054 1137 1062
rect 1149 1054 1150 1062
rect 1152 1054 1153 1062
rect 1165 1054 1166 1062
rect 1168 1054 1171 1062
rect 1173 1054 1174 1062
rect 1186 1054 1187 1062
rect 1189 1058 1190 1062
rect 1189 1054 1194 1058
rect 1202 1054 1203 1062
rect 1205 1054 1208 1062
rect 1210 1054 1211 1062
rect 1228 1054 1229 1062
rect 1231 1054 1232 1062
rect 1244 1054 1245 1062
rect 1247 1058 1248 1062
rect 1247 1054 1252 1058
rect 1260 1054 1261 1062
rect 1263 1054 1266 1062
rect 1268 1054 1269 1062
rect 1281 1054 1282 1062
rect 1284 1054 1285 1062
rect 1297 1054 1298 1062
rect 1300 1054 1303 1062
rect 1305 1054 1306 1062
rect 1318 1054 1319 1062
rect 1321 1058 1322 1062
rect 1321 1054 1326 1058
rect 1334 1054 1335 1062
rect 1337 1054 1340 1062
rect 1342 1054 1343 1062
rect 1360 1054 1361 1062
rect 1363 1054 1364 1062
rect 1376 1054 1377 1062
rect 1379 1058 1380 1062
rect 1379 1054 1384 1058
rect 1392 1054 1393 1062
rect 1395 1054 1398 1062
rect 1400 1054 1401 1062
rect 1413 1054 1414 1062
rect 1416 1054 1417 1062
rect 871 998 872 1006
rect 874 998 877 1006
rect 879 998 880 1006
rect 892 998 893 1006
rect 895 1002 896 1006
rect 895 998 900 1002
rect 908 998 909 1006
rect 911 998 914 1006
rect 916 998 917 1006
rect 934 998 935 1006
rect 937 998 938 1006
rect 950 998 951 1006
rect 953 1002 954 1006
rect 953 998 958 1002
rect 966 998 967 1006
rect 969 998 972 1006
rect 974 998 975 1006
rect 987 998 988 1006
rect 990 998 991 1006
rect 1804 998 1805 1006
rect 1807 998 1810 1006
rect 1812 998 1813 1006
rect 1825 998 1826 1006
rect 1828 1002 1829 1006
rect 1828 998 1833 1002
rect 1841 998 1842 1006
rect 1844 998 1847 1006
rect 1849 998 1850 1006
rect 1867 998 1868 1006
rect 1870 998 1871 1006
rect 1883 998 1884 1006
rect 1886 1002 1887 1006
rect 1886 998 1891 1002
rect 1899 998 1900 1006
rect 1902 998 1905 1006
rect 1907 998 1908 1006
rect 1920 998 1921 1006
rect 1923 998 1924 1006
rect 100 968 101 976
rect 103 968 106 976
rect 108 968 109 976
rect 121 968 122 976
rect 124 972 125 976
rect 124 968 129 972
rect 137 968 138 976
rect 140 968 143 976
rect 145 968 146 976
rect 163 968 164 976
rect 166 968 167 976
rect 179 968 180 976
rect 182 972 183 976
rect 182 968 187 972
rect 195 968 196 976
rect 198 968 201 976
rect 203 968 204 976
rect 216 968 217 976
rect 219 968 220 976
rect 232 968 233 976
rect 235 968 238 976
rect 240 968 241 976
rect 253 968 254 976
rect 256 972 257 976
rect 256 968 261 972
rect 269 968 270 976
rect 272 968 275 976
rect 277 968 278 976
rect 295 968 296 976
rect 298 968 299 976
rect 311 968 312 976
rect 314 972 315 976
rect 314 968 319 972
rect 327 968 328 976
rect 330 968 333 976
rect 335 968 336 976
rect 348 968 349 976
rect 351 968 352 976
rect 364 968 365 976
rect 367 968 370 976
rect 372 968 373 976
rect 385 968 386 976
rect 388 972 389 976
rect 388 968 393 972
rect 401 968 402 976
rect 404 968 407 976
rect 409 968 410 976
rect 427 968 428 976
rect 430 968 431 976
rect 443 968 444 976
rect 446 972 447 976
rect 446 968 451 972
rect 459 968 460 976
rect 462 968 465 976
rect 467 968 468 976
rect 480 968 481 976
rect 483 968 484 976
rect 1033 968 1034 976
rect 1036 968 1039 976
rect 1041 968 1042 976
rect 1054 968 1055 976
rect 1057 972 1058 976
rect 1057 968 1062 972
rect 1070 968 1071 976
rect 1073 968 1076 976
rect 1078 968 1079 976
rect 1096 968 1097 976
rect 1099 968 1100 976
rect 1112 968 1113 976
rect 1115 972 1116 976
rect 1115 968 1120 972
rect 1128 968 1129 976
rect 1131 968 1134 976
rect 1136 968 1137 976
rect 1149 968 1150 976
rect 1152 968 1153 976
rect 1165 968 1166 976
rect 1168 968 1171 976
rect 1173 968 1174 976
rect 1186 968 1187 976
rect 1189 972 1190 976
rect 1189 968 1194 972
rect 1202 968 1203 976
rect 1205 968 1208 976
rect 1210 968 1211 976
rect 1228 968 1229 976
rect 1231 968 1232 976
rect 1244 968 1245 976
rect 1247 972 1248 976
rect 1247 968 1252 972
rect 1260 968 1261 976
rect 1263 968 1266 976
rect 1268 968 1269 976
rect 1281 968 1282 976
rect 1284 968 1285 976
rect 1297 968 1298 976
rect 1300 968 1303 976
rect 1305 968 1306 976
rect 1318 968 1319 976
rect 1321 972 1322 976
rect 1321 968 1326 972
rect 1334 968 1335 976
rect 1337 968 1340 976
rect 1342 968 1343 976
rect 1360 968 1361 976
rect 1363 968 1364 976
rect 1376 968 1377 976
rect 1379 972 1380 976
rect 1379 968 1384 972
rect 1392 968 1393 976
rect 1395 968 1398 976
rect 1400 968 1401 976
rect 1413 968 1414 976
rect 1416 968 1417 976
rect 100 828 101 836
rect 103 828 106 836
rect 108 828 109 836
rect 121 828 122 836
rect 124 832 125 836
rect 124 828 129 832
rect 137 828 138 836
rect 140 828 143 836
rect 145 828 146 836
rect 163 828 164 836
rect 166 828 167 836
rect 179 828 180 836
rect 182 832 183 836
rect 182 828 187 832
rect 195 828 196 836
rect 198 828 201 836
rect 203 828 204 836
rect 216 828 217 836
rect 219 828 220 836
rect 232 828 233 836
rect 235 828 238 836
rect 240 828 241 836
rect 253 828 254 836
rect 256 832 257 836
rect 256 828 261 832
rect 269 828 270 836
rect 272 828 275 836
rect 277 828 278 836
rect 295 828 296 836
rect 298 828 299 836
rect 311 828 312 836
rect 314 832 315 836
rect 314 828 319 832
rect 327 828 328 836
rect 330 828 333 836
rect 335 828 336 836
rect 348 828 349 836
rect 351 828 352 836
rect 364 828 365 836
rect 367 828 370 836
rect 372 828 373 836
rect 385 828 386 836
rect 388 832 389 836
rect 388 828 393 832
rect 401 828 402 836
rect 404 828 407 836
rect 409 828 410 836
rect 427 828 428 836
rect 430 828 431 836
rect 443 828 444 836
rect 446 832 447 836
rect 446 828 451 832
rect 459 828 460 836
rect 462 828 465 836
rect 467 828 468 836
rect 480 828 481 836
rect 483 828 484 836
rect 1033 828 1034 836
rect 1036 828 1039 836
rect 1041 828 1042 836
rect 1054 828 1055 836
rect 1057 832 1058 836
rect 1057 828 1062 832
rect 1070 828 1071 836
rect 1073 828 1076 836
rect 1078 828 1079 836
rect 1096 828 1097 836
rect 1099 828 1100 836
rect 1112 828 1113 836
rect 1115 832 1116 836
rect 1115 828 1120 832
rect 1128 828 1129 836
rect 1131 828 1134 836
rect 1136 828 1137 836
rect 1149 828 1150 836
rect 1152 828 1153 836
rect 1165 828 1166 836
rect 1168 828 1171 836
rect 1173 828 1174 836
rect 1186 828 1187 836
rect 1189 832 1190 836
rect 1189 828 1194 832
rect 1202 828 1203 836
rect 1205 828 1208 836
rect 1210 828 1211 836
rect 1228 828 1229 836
rect 1231 828 1232 836
rect 1244 828 1245 836
rect 1247 832 1248 836
rect 1247 828 1252 832
rect 1260 828 1261 836
rect 1263 828 1266 836
rect 1268 828 1269 836
rect 1281 828 1282 836
rect 1284 828 1285 836
rect 1297 828 1298 836
rect 1300 828 1303 836
rect 1305 828 1306 836
rect 1318 828 1319 836
rect 1321 832 1322 836
rect 1321 828 1326 832
rect 1334 828 1335 836
rect 1337 828 1340 836
rect 1342 828 1343 836
rect 1360 828 1361 836
rect 1363 828 1364 836
rect 1376 828 1377 836
rect 1379 832 1380 836
rect 1379 828 1384 832
rect 1392 828 1393 836
rect 1395 828 1398 836
rect 1400 828 1401 836
rect 1413 828 1414 836
rect 1416 828 1417 836
rect 572 749 573 757
rect 575 749 578 757
rect 580 749 581 757
rect 593 749 594 757
rect 596 753 597 757
rect 596 749 601 753
rect 609 749 610 757
rect 612 749 615 757
rect 617 749 618 757
rect 635 749 636 757
rect 638 749 639 757
rect 651 749 652 757
rect 654 753 655 757
rect 654 749 659 753
rect 667 749 668 757
rect 670 749 673 757
rect 675 749 676 757
rect 688 749 689 757
rect 691 749 692 757
rect 704 749 705 757
rect 707 749 710 757
rect 712 749 713 757
rect 725 749 726 757
rect 728 753 729 757
rect 728 749 733 753
rect 741 749 742 757
rect 744 749 747 757
rect 749 749 750 757
rect 767 749 768 757
rect 770 749 771 757
rect 783 749 784 757
rect 786 753 787 757
rect 786 749 791 753
rect 799 749 800 757
rect 802 749 805 757
rect 807 749 808 757
rect 820 749 821 757
rect 823 749 824 757
rect 836 749 837 757
rect 839 749 842 757
rect 844 749 845 757
rect 857 749 858 757
rect 860 753 861 757
rect 860 749 865 753
rect 873 749 874 757
rect 876 749 879 757
rect 881 749 882 757
rect 899 749 900 757
rect 902 749 903 757
rect 915 749 916 757
rect 918 753 919 757
rect 918 749 923 753
rect 931 749 932 757
rect 934 749 937 757
rect 939 749 940 757
rect 952 749 953 757
rect 955 749 956 757
rect 968 749 969 757
rect 971 749 974 757
rect 976 749 977 757
rect 989 749 990 757
rect 992 753 993 757
rect 992 749 997 753
rect 1005 749 1006 757
rect 1008 749 1011 757
rect 1013 749 1014 757
rect 1031 749 1032 757
rect 1034 749 1035 757
rect 1047 749 1048 757
rect 1050 753 1051 757
rect 1050 749 1055 753
rect 1063 749 1064 757
rect 1066 749 1069 757
rect 1071 749 1072 757
rect 1084 749 1085 757
rect 1087 749 1088 757
rect 1505 749 1506 757
rect 1508 749 1511 757
rect 1513 749 1514 757
rect 1526 749 1527 757
rect 1529 753 1530 757
rect 1529 749 1534 753
rect 1542 749 1543 757
rect 1545 749 1548 757
rect 1550 749 1551 757
rect 1568 749 1569 757
rect 1571 749 1572 757
rect 1584 749 1585 757
rect 1587 753 1588 757
rect 1587 749 1592 753
rect 1600 749 1601 757
rect 1603 749 1606 757
rect 1608 749 1609 757
rect 1621 749 1622 757
rect 1624 749 1625 757
rect 1637 749 1638 757
rect 1640 749 1643 757
rect 1645 749 1646 757
rect 1658 749 1659 757
rect 1661 753 1662 757
rect 1661 749 1666 753
rect 1674 749 1675 757
rect 1677 749 1680 757
rect 1682 749 1683 757
rect 1700 749 1701 757
rect 1703 749 1704 757
rect 1716 749 1717 757
rect 1719 753 1720 757
rect 1719 749 1724 753
rect 1732 749 1733 757
rect 1735 749 1738 757
rect 1740 749 1741 757
rect 1753 749 1754 757
rect 1756 749 1757 757
rect 1769 749 1770 757
rect 1772 749 1775 757
rect 1777 749 1778 757
rect 1790 749 1791 757
rect 1793 753 1794 757
rect 1793 749 1798 753
rect 1806 749 1807 757
rect 1809 749 1812 757
rect 1814 749 1815 757
rect 1832 749 1833 757
rect 1835 749 1836 757
rect 1848 749 1849 757
rect 1851 753 1852 757
rect 1851 749 1856 753
rect 1864 749 1865 757
rect 1867 749 1870 757
rect 1872 749 1873 757
rect 1885 749 1886 757
rect 1888 749 1889 757
rect 1901 749 1902 757
rect 1904 749 1907 757
rect 1909 749 1910 757
rect 1922 749 1923 757
rect 1925 753 1926 757
rect 1925 749 1930 753
rect 1938 749 1939 757
rect 1941 749 1944 757
rect 1946 749 1947 757
rect 1964 749 1965 757
rect 1967 749 1968 757
rect 1980 749 1981 757
rect 1983 753 1984 757
rect 1983 749 1988 753
rect 1996 749 1997 757
rect 1999 749 2002 757
rect 2004 749 2005 757
rect 2017 749 2018 757
rect 2020 749 2021 757
rect 232 716 233 724
rect 235 716 238 724
rect 240 716 241 724
rect 253 716 254 724
rect 256 720 257 724
rect 256 716 261 720
rect 269 716 270 724
rect 272 716 275 724
rect 277 716 278 724
rect 295 716 296 724
rect 298 716 299 724
rect 311 716 312 724
rect 314 720 315 724
rect 314 716 319 720
rect 327 716 328 724
rect 330 716 333 724
rect 335 716 336 724
rect 348 716 349 724
rect 351 716 352 724
rect 1165 716 1166 724
rect 1168 716 1171 724
rect 1173 716 1174 724
rect 1186 716 1187 724
rect 1189 720 1190 724
rect 1189 716 1194 720
rect 1202 716 1203 724
rect 1205 716 1208 724
rect 1210 716 1211 724
rect 1228 716 1229 724
rect 1231 716 1232 724
rect 1244 716 1245 724
rect 1247 720 1248 724
rect 1247 716 1252 720
rect 1260 716 1261 724
rect 1263 716 1266 724
rect 1268 716 1269 724
rect 1281 716 1282 724
rect 1284 716 1285 724
rect 751 678 752 686
rect 754 678 755 686
rect 577 665 578 673
rect 580 665 581 673
rect 593 665 594 673
rect 596 665 597 673
rect 609 665 610 673
rect 612 665 613 673
rect 628 665 633 673
rect 635 665 638 673
rect 640 665 641 673
rect 662 665 664 673
rect 666 665 667 673
rect 684 665 685 673
rect 687 665 688 673
rect 700 665 705 673
rect 707 665 710 673
rect 712 665 713 673
rect 727 665 728 673
rect 730 665 731 673
rect 775 672 778 680
rect 780 672 783 680
rect 785 672 786 680
rect 805 678 806 686
rect 808 678 809 686
rect 832 678 833 686
rect 835 678 836 686
rect 856 672 859 680
rect 861 672 864 680
rect 866 672 867 680
rect 886 678 887 686
rect 889 678 890 686
rect 1684 678 1685 686
rect 1687 678 1688 686
rect 1510 665 1511 673
rect 1513 665 1514 673
rect 1526 665 1527 673
rect 1529 665 1530 673
rect 1542 665 1543 673
rect 1545 665 1546 673
rect 1561 665 1566 673
rect 1568 665 1571 673
rect 1573 665 1574 673
rect 1595 665 1597 673
rect 1599 665 1600 673
rect 1617 665 1618 673
rect 1620 665 1621 673
rect 1633 665 1638 673
rect 1640 665 1643 673
rect 1645 665 1646 673
rect 1660 665 1661 673
rect 1663 665 1664 673
rect 1708 672 1711 680
rect 1713 672 1716 680
rect 1718 672 1719 680
rect 1738 678 1739 686
rect 1741 678 1742 686
rect 1765 678 1766 686
rect 1768 678 1769 686
rect 1789 672 1792 680
rect 1794 672 1797 680
rect 1799 672 1800 680
rect 1819 678 1820 686
rect 1822 678 1823 686
rect 223 614 224 622
rect 226 614 227 622
rect 239 614 240 622
rect 242 614 245 622
rect 247 614 248 622
rect 260 618 261 622
rect 256 614 261 618
rect 263 614 264 622
rect 276 614 277 622
rect 279 614 280 622
rect 297 614 298 622
rect 300 614 303 622
rect 305 614 306 622
rect 318 618 319 622
rect 314 614 319 618
rect 321 614 322 622
rect 334 614 335 622
rect 337 614 340 622
rect 342 614 343 622
rect 1156 614 1157 622
rect 1159 614 1160 622
rect 1172 614 1173 622
rect 1175 614 1178 622
rect 1180 614 1181 622
rect 1193 618 1194 622
rect 1189 614 1194 618
rect 1196 614 1197 622
rect 1209 614 1210 622
rect 1212 614 1213 622
rect 1230 614 1231 622
rect 1233 614 1236 622
rect 1238 614 1239 622
rect 1251 618 1252 622
rect 1247 614 1252 618
rect 1254 614 1255 622
rect 1267 614 1268 622
rect 1270 614 1273 622
rect 1275 614 1276 622
rect 577 579 578 587
rect 580 579 581 587
rect 593 579 594 587
rect 596 579 597 587
rect 609 579 610 587
rect 612 579 613 587
rect 628 579 633 587
rect 635 579 638 587
rect 640 579 641 587
rect 662 579 664 587
rect 666 579 667 587
rect 684 579 685 587
rect 687 579 688 587
rect 700 579 705 587
rect 707 579 710 587
rect 712 579 713 587
rect 727 579 728 587
rect 730 579 731 587
rect 775 580 778 588
rect 780 580 783 588
rect 785 580 786 588
rect 856 580 859 588
rect 861 580 864 588
rect 866 580 867 588
rect 1510 579 1511 587
rect 1513 579 1514 587
rect 1526 579 1527 587
rect 1529 579 1530 587
rect 1542 579 1543 587
rect 1545 579 1546 587
rect 1561 579 1566 587
rect 1568 579 1571 587
rect 1573 579 1574 587
rect 1595 579 1597 587
rect 1599 579 1600 587
rect 1617 579 1618 587
rect 1620 579 1621 587
rect 1633 579 1638 587
rect 1640 579 1643 587
rect 1645 579 1646 587
rect 1660 579 1661 587
rect 1663 579 1664 587
rect 1708 580 1711 588
rect 1713 580 1716 588
rect 1718 580 1719 588
rect 1789 580 1792 588
rect 1794 580 1797 588
rect 1799 580 1800 588
rect 577 533 578 541
rect 580 533 581 541
rect 593 533 594 541
rect 596 533 597 541
rect 609 533 610 541
rect 612 533 613 541
rect 628 533 633 541
rect 635 533 638 541
rect 640 533 641 541
rect 662 533 664 541
rect 666 533 667 541
rect 684 533 685 541
rect 687 533 688 541
rect 700 533 705 541
rect 707 533 710 541
rect 712 533 713 541
rect 727 533 728 541
rect 730 533 731 541
rect 775 540 778 548
rect 780 540 783 548
rect 785 540 786 548
rect 805 546 806 554
rect 808 546 809 554
rect 856 546 857 554
rect 859 546 860 554
rect 880 540 883 548
rect 885 540 888 548
rect 890 540 891 548
rect 910 546 911 554
rect 913 546 914 554
rect 1510 533 1511 541
rect 1513 533 1514 541
rect 1526 533 1527 541
rect 1529 533 1530 541
rect 1542 533 1543 541
rect 1545 533 1546 541
rect 1561 533 1566 541
rect 1568 533 1571 541
rect 1573 533 1574 541
rect 1595 533 1597 541
rect 1599 533 1600 541
rect 1617 533 1618 541
rect 1620 533 1621 541
rect 1633 533 1638 541
rect 1640 533 1643 541
rect 1645 533 1646 541
rect 1660 533 1661 541
rect 1663 533 1664 541
rect 1708 540 1711 548
rect 1713 540 1716 548
rect 1718 540 1719 548
rect 1738 546 1739 554
rect 1741 546 1742 554
rect 1789 546 1790 554
rect 1792 546 1793 554
rect 1813 540 1816 548
rect 1818 540 1821 548
rect 1823 540 1824 548
rect 1843 546 1844 554
rect 1846 546 1847 554
rect 577 447 578 455
rect 580 447 581 455
rect 593 447 594 455
rect 596 447 597 455
rect 609 447 610 455
rect 612 447 613 455
rect 628 447 633 455
rect 635 447 638 455
rect 640 447 641 455
rect 662 447 664 455
rect 666 447 667 455
rect 684 447 685 455
rect 687 447 688 455
rect 700 447 705 455
rect 707 447 710 455
rect 712 447 713 455
rect 727 447 728 455
rect 730 447 731 455
rect 775 449 778 457
rect 780 449 783 457
rect 785 449 786 457
rect 880 449 883 457
rect 885 449 888 457
rect 890 449 891 457
rect 1510 447 1511 455
rect 1513 447 1514 455
rect 1526 447 1527 455
rect 1529 447 1530 455
rect 1542 447 1543 455
rect 1545 447 1546 455
rect 1561 447 1566 455
rect 1568 447 1571 455
rect 1573 447 1574 455
rect 1595 447 1597 455
rect 1599 447 1600 455
rect 1617 447 1618 455
rect 1620 447 1621 455
rect 1633 447 1638 455
rect 1640 447 1643 455
rect 1645 447 1646 455
rect 1660 447 1661 455
rect 1663 447 1664 455
rect 1708 449 1711 457
rect 1713 449 1716 457
rect 1718 449 1719 457
rect 1813 449 1816 457
rect 1818 449 1821 457
rect 1823 449 1824 457
rect 577 401 578 409
rect 580 401 581 409
rect 593 401 594 409
rect 596 401 597 409
rect 609 401 610 409
rect 612 401 613 409
rect 628 401 633 409
rect 635 401 638 409
rect 640 401 641 409
rect 662 401 664 409
rect 666 401 667 409
rect 684 401 685 409
rect 687 401 688 409
rect 700 401 705 409
rect 707 401 710 409
rect 712 401 713 409
rect 727 401 728 409
rect 730 401 731 409
rect 775 408 778 416
rect 780 408 783 416
rect 785 408 786 416
rect 805 414 806 422
rect 808 414 809 422
rect 832 414 833 422
rect 835 414 836 422
rect 856 408 859 416
rect 861 408 864 416
rect 866 408 867 416
rect 886 414 887 422
rect 889 414 890 422
rect 922 414 923 422
rect 925 414 926 422
rect 946 408 949 416
rect 951 408 954 416
rect 956 408 957 416
rect 976 414 977 422
rect 979 414 980 422
rect 1510 401 1511 409
rect 1513 401 1514 409
rect 1526 401 1527 409
rect 1529 401 1530 409
rect 1542 401 1543 409
rect 1545 401 1546 409
rect 1561 401 1566 409
rect 1568 401 1571 409
rect 1573 401 1574 409
rect 1595 401 1597 409
rect 1599 401 1600 409
rect 1617 401 1618 409
rect 1620 401 1621 409
rect 1633 401 1638 409
rect 1640 401 1643 409
rect 1645 401 1646 409
rect 1660 401 1661 409
rect 1663 401 1664 409
rect 1708 408 1711 416
rect 1713 408 1716 416
rect 1718 408 1719 416
rect 1738 414 1739 422
rect 1741 414 1742 422
rect 1765 414 1766 422
rect 1768 414 1769 422
rect 1789 408 1792 416
rect 1794 408 1797 416
rect 1799 408 1800 416
rect 1819 414 1820 422
rect 1822 414 1823 422
rect 1855 414 1856 422
rect 1858 414 1859 422
rect 1879 408 1882 416
rect 1884 408 1887 416
rect 1889 408 1890 416
rect 1909 414 1910 422
rect 1912 414 1913 422
rect 577 315 578 323
rect 580 315 581 323
rect 593 315 594 323
rect 596 315 597 323
rect 609 315 610 323
rect 612 315 613 323
rect 628 315 633 323
rect 635 315 638 323
rect 640 315 641 323
rect 662 315 664 323
rect 666 315 667 323
rect 684 315 685 323
rect 687 315 688 323
rect 700 315 705 323
rect 707 315 710 323
rect 712 315 713 323
rect 727 315 728 323
rect 730 315 731 323
rect 775 314 778 322
rect 780 314 783 322
rect 785 314 786 322
rect 856 314 859 322
rect 861 314 864 322
rect 866 314 867 322
rect 946 314 949 322
rect 951 314 954 322
rect 956 314 957 322
rect 1510 315 1511 323
rect 1513 315 1514 323
rect 1526 315 1527 323
rect 1529 315 1530 323
rect 1542 315 1543 323
rect 1545 315 1546 323
rect 1561 315 1566 323
rect 1568 315 1571 323
rect 1573 315 1574 323
rect 1595 315 1597 323
rect 1599 315 1600 323
rect 1617 315 1618 323
rect 1620 315 1621 323
rect 1633 315 1638 323
rect 1640 315 1643 323
rect 1645 315 1646 323
rect 1660 315 1661 323
rect 1663 315 1664 323
rect 1708 314 1711 322
rect 1713 314 1716 322
rect 1718 314 1719 322
rect 1789 314 1792 322
rect 1794 314 1797 322
rect 1799 314 1800 322
rect 1879 314 1882 322
rect 1884 314 1887 322
rect 1889 314 1890 322
rect 577 269 578 277
rect 580 269 581 277
rect 593 269 594 277
rect 596 269 597 277
rect 609 269 610 277
rect 612 269 613 277
rect 628 269 633 277
rect 635 269 638 277
rect 640 269 641 277
rect 662 269 664 277
rect 666 269 667 277
rect 684 269 685 277
rect 687 269 688 277
rect 700 269 705 277
rect 707 269 710 277
rect 712 269 713 277
rect 727 269 728 277
rect 730 269 731 277
rect 775 276 778 284
rect 780 276 783 284
rect 785 276 786 284
rect 805 282 806 290
rect 808 282 809 290
rect 1510 269 1511 277
rect 1513 269 1514 277
rect 1526 269 1527 277
rect 1529 269 1530 277
rect 1542 269 1543 277
rect 1545 269 1546 277
rect 1561 269 1566 277
rect 1568 269 1571 277
rect 1573 269 1574 277
rect 1595 269 1597 277
rect 1599 269 1600 277
rect 1617 269 1618 277
rect 1620 269 1621 277
rect 1633 269 1638 277
rect 1640 269 1643 277
rect 1645 269 1646 277
rect 1660 269 1661 277
rect 1663 269 1664 277
rect 1708 276 1711 284
rect 1713 276 1716 284
rect 1718 276 1719 284
rect 1738 282 1739 290
rect 1741 282 1742 290
rect 100 214 101 222
rect 103 214 106 222
rect 108 214 109 222
rect 121 214 122 222
rect 124 218 125 222
rect 124 214 129 218
rect 137 214 138 222
rect 140 214 143 222
rect 145 214 146 222
rect 163 214 164 222
rect 166 214 167 222
rect 179 214 180 222
rect 182 218 183 222
rect 182 214 187 218
rect 195 214 196 222
rect 198 214 201 222
rect 203 214 204 222
rect 216 214 217 222
rect 219 214 220 222
rect 232 214 233 222
rect 235 214 238 222
rect 240 214 241 222
rect 253 214 254 222
rect 256 218 257 222
rect 256 214 261 218
rect 269 214 270 222
rect 272 214 275 222
rect 277 214 278 222
rect 295 214 296 222
rect 298 214 299 222
rect 311 214 312 222
rect 314 218 315 222
rect 314 214 319 218
rect 327 214 328 222
rect 330 214 333 222
rect 335 214 336 222
rect 348 214 349 222
rect 351 214 352 222
rect 364 214 365 222
rect 367 214 370 222
rect 372 214 373 222
rect 385 214 386 222
rect 388 218 389 222
rect 388 214 393 218
rect 401 214 402 222
rect 404 214 407 222
rect 409 214 410 222
rect 427 214 428 222
rect 430 214 431 222
rect 443 214 444 222
rect 446 218 447 222
rect 446 214 451 218
rect 459 214 460 222
rect 462 214 465 222
rect 467 214 468 222
rect 480 214 481 222
rect 483 214 484 222
rect 1033 214 1034 222
rect 1036 214 1039 222
rect 1041 214 1042 222
rect 1054 214 1055 222
rect 1057 218 1058 222
rect 1057 214 1062 218
rect 1070 214 1071 222
rect 1073 214 1076 222
rect 1078 214 1079 222
rect 1096 214 1097 222
rect 1099 214 1100 222
rect 1112 214 1113 222
rect 1115 218 1116 222
rect 1115 214 1120 218
rect 1128 214 1129 222
rect 1131 214 1134 222
rect 1136 214 1137 222
rect 1149 214 1150 222
rect 1152 214 1153 222
rect 1165 214 1166 222
rect 1168 214 1171 222
rect 1173 214 1174 222
rect 1186 214 1187 222
rect 1189 218 1190 222
rect 1189 214 1194 218
rect 1202 214 1203 222
rect 1205 214 1208 222
rect 1210 214 1211 222
rect 1228 214 1229 222
rect 1231 214 1232 222
rect 1244 214 1245 222
rect 1247 218 1248 222
rect 1247 214 1252 218
rect 1260 214 1261 222
rect 1263 214 1266 222
rect 1268 214 1269 222
rect 1281 214 1282 222
rect 1284 214 1285 222
rect 1297 214 1298 222
rect 1300 214 1303 222
rect 1305 214 1306 222
rect 1318 214 1319 222
rect 1321 218 1322 222
rect 1321 214 1326 218
rect 1334 214 1335 222
rect 1337 214 1340 222
rect 1342 214 1343 222
rect 1360 214 1361 222
rect 1363 214 1364 222
rect 1376 214 1377 222
rect 1379 218 1380 222
rect 1379 214 1384 218
rect 1392 214 1393 222
rect 1395 214 1398 222
rect 1400 214 1401 222
rect 1413 214 1414 222
rect 1416 214 1417 222
rect 577 183 578 191
rect 580 183 581 191
rect 593 183 594 191
rect 596 183 597 191
rect 609 183 610 191
rect 612 183 613 191
rect 628 183 633 191
rect 635 183 638 191
rect 640 183 641 191
rect 662 183 664 191
rect 666 183 667 191
rect 684 183 685 191
rect 687 183 688 191
rect 700 183 705 191
rect 707 183 710 191
rect 712 183 713 191
rect 727 183 728 191
rect 730 183 731 191
rect 775 178 778 186
rect 780 178 783 186
rect 785 178 786 186
rect 811 183 812 191
rect 814 183 815 191
rect 819 183 825 191
rect 829 183 830 191
rect 832 183 833 191
rect 854 183 855 191
rect 857 183 858 191
rect 870 183 871 191
rect 873 183 874 191
rect 889 183 894 191
rect 896 183 899 191
rect 901 183 902 191
rect 923 183 925 191
rect 927 183 928 191
rect 945 183 946 191
rect 948 183 949 191
rect 961 183 966 191
rect 968 183 971 191
rect 973 183 974 191
rect 988 183 989 191
rect 991 183 992 191
rect 1510 183 1511 191
rect 1513 183 1514 191
rect 1526 183 1527 191
rect 1529 183 1530 191
rect 1542 183 1543 191
rect 1545 183 1546 191
rect 1561 183 1566 191
rect 1568 183 1571 191
rect 1573 183 1574 191
rect 1595 183 1597 191
rect 1599 183 1600 191
rect 1617 183 1618 191
rect 1620 183 1621 191
rect 1633 183 1638 191
rect 1640 183 1643 191
rect 1645 183 1646 191
rect 1660 183 1661 191
rect 1663 183 1664 191
rect 1708 178 1711 186
rect 1713 178 1716 186
rect 1718 178 1719 186
rect 1744 183 1745 191
rect 1747 183 1748 191
rect 1752 183 1758 191
rect 1762 183 1763 191
rect 1765 183 1766 191
rect 1787 183 1788 191
rect 1790 183 1791 191
rect 1803 183 1804 191
rect 1806 183 1807 191
rect 1822 183 1827 191
rect 1829 183 1832 191
rect 1834 183 1835 191
rect 1856 183 1858 191
rect 1860 183 1861 191
rect 1878 183 1879 191
rect 1881 183 1882 191
rect 1894 183 1899 191
rect 1901 183 1904 191
rect 1906 183 1907 191
rect 1921 183 1922 191
rect 1924 183 1925 191
rect 871 104 872 112
rect 874 104 877 112
rect 879 104 880 112
rect 892 104 893 112
rect 895 108 896 112
rect 895 104 900 108
rect 908 104 909 112
rect 911 104 914 112
rect 916 104 917 112
rect 934 104 935 112
rect 937 104 938 112
rect 950 104 951 112
rect 953 108 954 112
rect 953 104 958 108
rect 966 104 967 112
rect 969 104 972 112
rect 974 104 975 112
rect 987 104 988 112
rect 990 104 991 112
rect 1804 104 1805 112
rect 1807 104 1810 112
rect 1812 104 1813 112
rect 1825 104 1826 112
rect 1828 108 1829 112
rect 1828 104 1833 108
rect 1841 104 1842 112
rect 1844 104 1847 112
rect 1849 104 1850 112
rect 1867 104 1868 112
rect 1870 104 1871 112
rect 1883 104 1884 112
rect 1886 108 1887 112
rect 1886 104 1891 108
rect 1899 104 1900 112
rect 1902 104 1905 112
rect 1907 104 1908 112
rect 1920 104 1921 112
rect 1923 104 1924 112
rect 100 74 101 82
rect 103 74 106 82
rect 108 74 109 82
rect 121 74 122 82
rect 124 78 125 82
rect 124 74 129 78
rect 137 74 138 82
rect 140 74 143 82
rect 145 74 146 82
rect 163 74 164 82
rect 166 74 167 82
rect 179 74 180 82
rect 182 78 183 82
rect 182 74 187 78
rect 195 74 196 82
rect 198 74 201 82
rect 203 74 204 82
rect 216 74 217 82
rect 219 74 220 82
rect 232 74 233 82
rect 235 74 238 82
rect 240 74 241 82
rect 253 74 254 82
rect 256 78 257 82
rect 256 74 261 78
rect 269 74 270 82
rect 272 74 275 82
rect 277 74 278 82
rect 295 74 296 82
rect 298 74 299 82
rect 311 74 312 82
rect 314 78 315 82
rect 314 74 319 78
rect 327 74 328 82
rect 330 74 333 82
rect 335 74 336 82
rect 348 74 349 82
rect 351 74 352 82
rect 364 74 365 82
rect 367 74 370 82
rect 372 74 373 82
rect 385 74 386 82
rect 388 78 389 82
rect 388 74 393 78
rect 401 74 402 82
rect 404 74 407 82
rect 409 74 410 82
rect 427 74 428 82
rect 430 74 431 82
rect 443 74 444 82
rect 446 78 447 82
rect 446 74 451 78
rect 459 74 460 82
rect 462 74 465 82
rect 467 74 468 82
rect 480 74 481 82
rect 483 74 484 82
rect 1033 74 1034 82
rect 1036 74 1039 82
rect 1041 74 1042 82
rect 1054 74 1055 82
rect 1057 78 1058 82
rect 1057 74 1062 78
rect 1070 74 1071 82
rect 1073 74 1076 82
rect 1078 74 1079 82
rect 1096 74 1097 82
rect 1099 74 1100 82
rect 1112 74 1113 82
rect 1115 78 1116 82
rect 1115 74 1120 78
rect 1128 74 1129 82
rect 1131 74 1134 82
rect 1136 74 1137 82
rect 1149 74 1150 82
rect 1152 74 1153 82
rect 1165 74 1166 82
rect 1168 74 1171 82
rect 1173 74 1174 82
rect 1186 74 1187 82
rect 1189 78 1190 82
rect 1189 74 1194 78
rect 1202 74 1203 82
rect 1205 74 1208 82
rect 1210 74 1211 82
rect 1228 74 1229 82
rect 1231 74 1232 82
rect 1244 74 1245 82
rect 1247 78 1248 82
rect 1247 74 1252 78
rect 1260 74 1261 82
rect 1263 74 1266 82
rect 1268 74 1269 82
rect 1281 74 1282 82
rect 1284 74 1285 82
rect 1297 74 1298 82
rect 1300 74 1303 82
rect 1305 74 1306 82
rect 1318 74 1319 82
rect 1321 78 1322 82
rect 1321 74 1326 78
rect 1334 74 1335 82
rect 1337 74 1340 82
rect 1342 74 1343 82
rect 1360 74 1361 82
rect 1363 74 1364 82
rect 1376 74 1377 82
rect 1379 78 1380 82
rect 1379 74 1384 78
rect 1392 74 1393 82
rect 1395 74 1398 82
rect 1400 74 1401 82
rect 1413 74 1414 82
rect 1416 74 1417 82
rect 871 18 872 26
rect 874 18 877 26
rect 879 18 880 26
rect 892 18 893 26
rect 895 22 896 26
rect 895 18 900 22
rect 908 18 909 26
rect 911 18 914 26
rect 916 18 917 26
rect 934 18 935 26
rect 937 18 938 26
rect 950 18 951 26
rect 953 22 954 26
rect 953 18 958 22
rect 966 18 967 26
rect 969 18 972 26
rect 974 18 975 26
rect 987 18 988 26
rect 990 18 991 26
rect 1804 18 1805 26
rect 1807 18 1810 26
rect 1812 18 1813 26
rect 1825 18 1826 26
rect 1828 22 1829 26
rect 1828 18 1833 22
rect 1841 18 1842 26
rect 1844 18 1847 26
rect 1849 18 1850 26
rect 1867 18 1868 26
rect 1870 18 1871 26
rect 1883 18 1884 26
rect 1886 22 1887 26
rect 1886 18 1891 22
rect 1899 18 1900 26
rect 1902 18 1905 26
rect 1907 18 1908 26
rect 1920 18 1921 26
rect 1923 18 1924 26
rect 100 -12 101 -4
rect 103 -12 106 -4
rect 108 -12 109 -4
rect 121 -12 122 -4
rect 124 -8 125 -4
rect 124 -12 129 -8
rect 137 -12 138 -4
rect 140 -12 143 -4
rect 145 -12 146 -4
rect 163 -12 164 -4
rect 166 -12 167 -4
rect 179 -12 180 -4
rect 182 -8 183 -4
rect 182 -12 187 -8
rect 195 -12 196 -4
rect 198 -12 201 -4
rect 203 -12 204 -4
rect 216 -12 217 -4
rect 219 -12 220 -4
rect 232 -12 233 -4
rect 235 -12 238 -4
rect 240 -12 241 -4
rect 253 -12 254 -4
rect 256 -8 257 -4
rect 256 -12 261 -8
rect 269 -12 270 -4
rect 272 -12 275 -4
rect 277 -12 278 -4
rect 295 -12 296 -4
rect 298 -12 299 -4
rect 311 -12 312 -4
rect 314 -8 315 -4
rect 314 -12 319 -8
rect 327 -12 328 -4
rect 330 -12 333 -4
rect 335 -12 336 -4
rect 348 -12 349 -4
rect 351 -12 352 -4
rect 364 -12 365 -4
rect 367 -12 370 -4
rect 372 -12 373 -4
rect 385 -12 386 -4
rect 388 -8 389 -4
rect 388 -12 393 -8
rect 401 -12 402 -4
rect 404 -12 407 -4
rect 409 -12 410 -4
rect 427 -12 428 -4
rect 430 -12 431 -4
rect 443 -12 444 -4
rect 446 -8 447 -4
rect 446 -12 451 -8
rect 459 -12 460 -4
rect 462 -12 465 -4
rect 467 -12 468 -4
rect 480 -12 481 -4
rect 483 -12 484 -4
rect 1033 -12 1034 -4
rect 1036 -12 1039 -4
rect 1041 -12 1042 -4
rect 1054 -12 1055 -4
rect 1057 -8 1058 -4
rect 1057 -12 1062 -8
rect 1070 -12 1071 -4
rect 1073 -12 1076 -4
rect 1078 -12 1079 -4
rect 1096 -12 1097 -4
rect 1099 -12 1100 -4
rect 1112 -12 1113 -4
rect 1115 -8 1116 -4
rect 1115 -12 1120 -8
rect 1128 -12 1129 -4
rect 1131 -12 1134 -4
rect 1136 -12 1137 -4
rect 1149 -12 1150 -4
rect 1152 -12 1153 -4
rect 1165 -12 1166 -4
rect 1168 -12 1171 -4
rect 1173 -12 1174 -4
rect 1186 -12 1187 -4
rect 1189 -8 1190 -4
rect 1189 -12 1194 -8
rect 1202 -12 1203 -4
rect 1205 -12 1208 -4
rect 1210 -12 1211 -4
rect 1228 -12 1229 -4
rect 1231 -12 1232 -4
rect 1244 -12 1245 -4
rect 1247 -8 1248 -4
rect 1247 -12 1252 -8
rect 1260 -12 1261 -4
rect 1263 -12 1266 -4
rect 1268 -12 1269 -4
rect 1281 -12 1282 -4
rect 1284 -12 1285 -4
rect 1297 -12 1298 -4
rect 1300 -12 1303 -4
rect 1305 -12 1306 -4
rect 1318 -12 1319 -4
rect 1321 -8 1322 -4
rect 1321 -12 1326 -8
rect 1334 -12 1335 -4
rect 1337 -12 1340 -4
rect 1342 -12 1343 -4
rect 1360 -12 1361 -4
rect 1363 -12 1364 -4
rect 1376 -12 1377 -4
rect 1379 -8 1380 -4
rect 1379 -12 1384 -8
rect 1392 -12 1393 -4
rect 1395 -12 1398 -4
rect 1400 -12 1401 -4
rect 1413 -12 1414 -4
rect 1416 -12 1417 -4
rect 100 -152 101 -144
rect 103 -152 106 -144
rect 108 -152 109 -144
rect 121 -152 122 -144
rect 124 -148 125 -144
rect 124 -152 129 -148
rect 137 -152 138 -144
rect 140 -152 143 -144
rect 145 -152 146 -144
rect 163 -152 164 -144
rect 166 -152 167 -144
rect 179 -152 180 -144
rect 182 -148 183 -144
rect 182 -152 187 -148
rect 195 -152 196 -144
rect 198 -152 201 -144
rect 203 -152 204 -144
rect 216 -152 217 -144
rect 219 -152 220 -144
rect 232 -152 233 -144
rect 235 -152 238 -144
rect 240 -152 241 -144
rect 253 -152 254 -144
rect 256 -148 257 -144
rect 256 -152 261 -148
rect 269 -152 270 -144
rect 272 -152 275 -144
rect 277 -152 278 -144
rect 295 -152 296 -144
rect 298 -152 299 -144
rect 311 -152 312 -144
rect 314 -148 315 -144
rect 314 -152 319 -148
rect 327 -152 328 -144
rect 330 -152 333 -144
rect 335 -152 336 -144
rect 348 -152 349 -144
rect 351 -152 352 -144
rect 364 -152 365 -144
rect 367 -152 370 -144
rect 372 -152 373 -144
rect 385 -152 386 -144
rect 388 -148 389 -144
rect 388 -152 393 -148
rect 401 -152 402 -144
rect 404 -152 407 -144
rect 409 -152 410 -144
rect 427 -152 428 -144
rect 430 -152 431 -144
rect 443 -152 444 -144
rect 446 -148 447 -144
rect 446 -152 451 -148
rect 459 -152 460 -144
rect 462 -152 465 -144
rect 467 -152 468 -144
rect 480 -152 481 -144
rect 483 -152 484 -144
rect 1033 -152 1034 -144
rect 1036 -152 1039 -144
rect 1041 -152 1042 -144
rect 1054 -152 1055 -144
rect 1057 -148 1058 -144
rect 1057 -152 1062 -148
rect 1070 -152 1071 -144
rect 1073 -152 1076 -144
rect 1078 -152 1079 -144
rect 1096 -152 1097 -144
rect 1099 -152 1100 -144
rect 1112 -152 1113 -144
rect 1115 -148 1116 -144
rect 1115 -152 1120 -148
rect 1128 -152 1129 -144
rect 1131 -152 1134 -144
rect 1136 -152 1137 -144
rect 1149 -152 1150 -144
rect 1152 -152 1153 -144
rect 1165 -152 1166 -144
rect 1168 -152 1171 -144
rect 1173 -152 1174 -144
rect 1186 -152 1187 -144
rect 1189 -148 1190 -144
rect 1189 -152 1194 -148
rect 1202 -152 1203 -144
rect 1205 -152 1208 -144
rect 1210 -152 1211 -144
rect 1228 -152 1229 -144
rect 1231 -152 1232 -144
rect 1244 -152 1245 -144
rect 1247 -148 1248 -144
rect 1247 -152 1252 -148
rect 1260 -152 1261 -144
rect 1263 -152 1266 -144
rect 1268 -152 1269 -144
rect 1281 -152 1282 -144
rect 1284 -152 1285 -144
rect 1297 -152 1298 -144
rect 1300 -152 1303 -144
rect 1305 -152 1306 -144
rect 1318 -152 1319 -144
rect 1321 -148 1322 -144
rect 1321 -152 1326 -148
rect 1334 -152 1335 -144
rect 1337 -152 1340 -144
rect 1342 -152 1343 -144
rect 1360 -152 1361 -144
rect 1363 -152 1364 -144
rect 1376 -152 1377 -144
rect 1379 -148 1380 -144
rect 1379 -152 1384 -148
rect 1392 -152 1393 -144
rect 1395 -152 1398 -144
rect 1400 -152 1401 -144
rect 1413 -152 1414 -144
rect 1416 -152 1417 -144
<< ndcontact >>
rect 568 1706 572 1710
rect 581 1706 585 1710
rect 589 1706 593 1710
rect 597 1706 601 1710
rect 605 1706 609 1710
rect 618 1706 622 1710
rect 631 1706 635 1710
rect 639 1706 643 1710
rect 647 1706 651 1710
rect 655 1706 659 1710
rect 663 1706 667 1710
rect 676 1706 680 1710
rect 684 1706 688 1710
rect 692 1706 696 1710
rect 700 1706 704 1710
rect 713 1706 717 1710
rect 721 1706 725 1710
rect 729 1706 733 1710
rect 737 1706 741 1710
rect 750 1706 754 1710
rect 763 1706 767 1710
rect 771 1706 775 1710
rect 779 1706 783 1710
rect 787 1706 791 1710
rect 795 1706 799 1710
rect 808 1706 812 1710
rect 816 1706 820 1710
rect 824 1706 828 1710
rect 832 1706 836 1710
rect 845 1706 849 1710
rect 853 1706 857 1710
rect 861 1706 865 1710
rect 869 1706 873 1710
rect 882 1706 886 1710
rect 895 1706 899 1710
rect 903 1706 907 1710
rect 911 1706 915 1710
rect 919 1706 923 1710
rect 927 1706 931 1710
rect 940 1706 944 1710
rect 948 1706 952 1710
rect 956 1706 960 1710
rect 964 1706 968 1710
rect 977 1706 981 1710
rect 985 1706 989 1710
rect 993 1706 997 1710
rect 1001 1706 1005 1710
rect 1014 1706 1018 1710
rect 1027 1706 1031 1710
rect 1035 1706 1039 1710
rect 1043 1706 1047 1710
rect 1051 1706 1055 1710
rect 1059 1706 1063 1710
rect 1072 1706 1076 1710
rect 1080 1706 1084 1710
rect 1088 1706 1092 1710
rect 1501 1706 1505 1710
rect 1514 1706 1518 1710
rect 1522 1706 1526 1710
rect 1530 1706 1534 1710
rect 1538 1706 1542 1710
rect 1551 1706 1555 1710
rect 1564 1706 1568 1710
rect 1572 1706 1576 1710
rect 1580 1706 1584 1710
rect 1588 1706 1592 1710
rect 1596 1706 1600 1710
rect 1609 1706 1613 1710
rect 1617 1706 1621 1710
rect 1625 1706 1629 1710
rect 1633 1706 1637 1710
rect 1646 1706 1650 1710
rect 1654 1706 1658 1710
rect 1662 1706 1666 1710
rect 1670 1706 1674 1710
rect 1683 1706 1687 1710
rect 1696 1706 1700 1710
rect 1704 1706 1708 1710
rect 1712 1706 1716 1710
rect 1720 1706 1724 1710
rect 1728 1706 1732 1710
rect 1741 1706 1745 1710
rect 1749 1706 1753 1710
rect 1757 1706 1761 1710
rect 1765 1706 1769 1710
rect 1778 1706 1782 1710
rect 1786 1706 1790 1710
rect 1794 1706 1798 1710
rect 1802 1706 1806 1710
rect 1815 1706 1819 1710
rect 1828 1706 1832 1710
rect 1836 1706 1840 1710
rect 1844 1706 1848 1710
rect 1852 1706 1856 1710
rect 1860 1706 1864 1710
rect 1873 1706 1877 1710
rect 1881 1706 1885 1710
rect 1889 1706 1893 1710
rect 1897 1706 1901 1710
rect 1910 1706 1914 1710
rect 1918 1706 1922 1710
rect 1926 1706 1930 1710
rect 1934 1706 1938 1710
rect 1947 1706 1951 1710
rect 1960 1706 1964 1710
rect 1968 1706 1972 1710
rect 1976 1706 1980 1710
rect 1984 1706 1988 1710
rect 1992 1706 1996 1710
rect 2005 1706 2009 1710
rect 2013 1706 2017 1710
rect 2021 1706 2025 1710
rect 228 1673 232 1677
rect 241 1673 245 1677
rect 249 1673 253 1677
rect 257 1673 261 1677
rect 265 1673 269 1677
rect 278 1673 282 1677
rect 291 1673 295 1677
rect 299 1673 303 1677
rect 307 1673 311 1677
rect 315 1673 319 1677
rect 323 1673 327 1677
rect 336 1673 340 1677
rect 344 1673 348 1677
rect 352 1673 356 1677
rect 1161 1673 1165 1677
rect 1174 1673 1178 1677
rect 1182 1673 1186 1677
rect 1190 1673 1194 1677
rect 1198 1673 1202 1677
rect 1211 1673 1215 1677
rect 1224 1673 1228 1677
rect 1232 1673 1236 1677
rect 1240 1673 1244 1677
rect 1248 1673 1252 1677
rect 1256 1673 1260 1677
rect 1269 1673 1273 1677
rect 1277 1673 1281 1677
rect 1285 1673 1289 1677
rect 352 1636 356 1640
rect 360 1636 364 1640
rect 747 1640 751 1644
rect 755 1640 759 1644
rect 771 1636 775 1640
rect 786 1636 790 1640
rect 828 1640 832 1644
rect 836 1640 840 1644
rect 852 1636 856 1640
rect 867 1636 871 1640
rect 801 1632 805 1636
rect 809 1632 813 1636
rect 235 1627 239 1631
rect 243 1627 247 1631
rect 573 1627 577 1631
rect 581 1627 585 1631
rect 589 1627 593 1631
rect 597 1627 601 1631
rect 605 1627 609 1631
rect 613 1627 617 1631
rect 624 1627 628 1631
rect 641 1627 645 1631
rect 658 1627 662 1631
rect 667 1627 671 1631
rect 680 1627 684 1631
rect 688 1627 692 1631
rect 696 1627 700 1631
rect 713 1627 717 1631
rect 723 1627 727 1631
rect 731 1627 735 1631
rect 882 1632 886 1636
rect 890 1632 894 1636
rect 1285 1636 1289 1640
rect 1293 1636 1297 1640
rect 1680 1640 1684 1644
rect 1688 1640 1692 1644
rect 1704 1636 1708 1640
rect 1719 1636 1723 1640
rect 1761 1640 1765 1644
rect 1769 1640 1773 1644
rect 1785 1636 1789 1640
rect 1800 1636 1804 1640
rect 1734 1632 1738 1636
rect 1742 1632 1746 1636
rect 1168 1627 1172 1631
rect 1176 1627 1180 1631
rect 1506 1627 1510 1631
rect 1514 1627 1518 1631
rect 1522 1627 1526 1631
rect 1530 1627 1534 1631
rect 1538 1627 1542 1631
rect 1546 1627 1550 1631
rect 1557 1627 1561 1631
rect 1574 1627 1578 1631
rect 1591 1627 1595 1631
rect 1600 1627 1604 1631
rect 1613 1627 1617 1631
rect 1621 1627 1625 1631
rect 1629 1627 1633 1631
rect 1646 1627 1650 1631
rect 1656 1627 1660 1631
rect 1664 1627 1668 1631
rect 1815 1632 1819 1636
rect 1823 1632 1827 1636
rect 573 1581 577 1585
rect 581 1581 585 1585
rect 589 1581 593 1585
rect 597 1581 601 1585
rect 605 1581 609 1585
rect 613 1581 617 1585
rect 624 1581 628 1585
rect 641 1581 645 1585
rect 658 1581 662 1585
rect 667 1581 671 1585
rect 680 1581 684 1585
rect 688 1581 692 1585
rect 696 1581 700 1585
rect 713 1581 717 1585
rect 723 1581 727 1585
rect 731 1581 735 1585
rect 219 1571 223 1575
rect 227 1571 231 1575
rect 235 1571 239 1575
rect 248 1571 252 1575
rect 256 1571 260 1575
rect 264 1571 268 1575
rect 272 1571 276 1575
rect 280 1571 284 1575
rect 293 1571 297 1575
rect 306 1571 310 1575
rect 314 1571 318 1575
rect 322 1571 326 1575
rect 330 1571 334 1575
rect 343 1571 347 1575
rect 771 1580 775 1584
rect 786 1580 790 1584
rect 852 1580 856 1584
rect 867 1580 871 1584
rect 1506 1581 1510 1585
rect 1514 1581 1518 1585
rect 1522 1581 1526 1585
rect 1530 1581 1534 1585
rect 1538 1581 1542 1585
rect 1546 1581 1550 1585
rect 1557 1581 1561 1585
rect 1574 1581 1578 1585
rect 1591 1581 1595 1585
rect 1600 1581 1604 1585
rect 1613 1581 1617 1585
rect 1621 1581 1625 1585
rect 1629 1581 1633 1585
rect 1646 1581 1650 1585
rect 1656 1581 1660 1585
rect 1664 1581 1668 1585
rect 1152 1571 1156 1575
rect 1160 1571 1164 1575
rect 1168 1571 1172 1575
rect 1181 1571 1185 1575
rect 1189 1571 1193 1575
rect 1197 1571 1201 1575
rect 1205 1571 1209 1575
rect 1213 1571 1217 1575
rect 1226 1571 1230 1575
rect 1239 1571 1243 1575
rect 1247 1571 1251 1575
rect 1255 1571 1259 1575
rect 1263 1571 1267 1575
rect 1276 1571 1280 1575
rect 1704 1580 1708 1584
rect 1719 1580 1723 1584
rect 1785 1580 1789 1584
rect 1800 1580 1804 1584
rect 771 1504 775 1508
rect 786 1504 790 1508
rect 852 1508 856 1512
rect 860 1508 864 1512
rect 876 1504 880 1508
rect 891 1504 895 1508
rect 801 1500 805 1504
rect 809 1500 813 1504
rect 573 1495 577 1499
rect 581 1495 585 1499
rect 589 1495 593 1499
rect 597 1495 601 1499
rect 605 1495 609 1499
rect 613 1495 617 1499
rect 624 1495 628 1499
rect 641 1495 645 1499
rect 658 1495 662 1499
rect 667 1495 671 1499
rect 680 1495 684 1499
rect 688 1495 692 1499
rect 696 1495 700 1499
rect 713 1495 717 1499
rect 723 1495 727 1499
rect 731 1495 735 1499
rect 906 1500 910 1504
rect 914 1500 918 1504
rect 1704 1504 1708 1508
rect 1719 1504 1723 1508
rect 1785 1508 1789 1512
rect 1793 1508 1797 1512
rect 1809 1504 1813 1508
rect 1824 1504 1828 1508
rect 1734 1500 1738 1504
rect 1742 1500 1746 1504
rect 1506 1495 1510 1499
rect 1514 1495 1518 1499
rect 1522 1495 1526 1499
rect 1530 1495 1534 1499
rect 1538 1495 1542 1499
rect 1546 1495 1550 1499
rect 1557 1495 1561 1499
rect 1574 1495 1578 1499
rect 1591 1495 1595 1499
rect 1600 1495 1604 1499
rect 1613 1495 1617 1499
rect 1621 1495 1625 1499
rect 1629 1495 1633 1499
rect 1646 1495 1650 1499
rect 1656 1495 1660 1499
rect 1664 1495 1668 1499
rect 1839 1500 1843 1504
rect 1847 1500 1851 1504
rect 573 1449 577 1453
rect 581 1449 585 1453
rect 589 1449 593 1453
rect 597 1449 601 1453
rect 605 1449 609 1453
rect 613 1449 617 1453
rect 624 1449 628 1453
rect 641 1449 645 1453
rect 658 1449 662 1453
rect 667 1449 671 1453
rect 680 1449 684 1453
rect 688 1449 692 1453
rect 696 1449 700 1453
rect 713 1449 717 1453
rect 723 1449 727 1453
rect 731 1449 735 1453
rect 771 1449 775 1453
rect 786 1449 790 1453
rect 876 1449 880 1453
rect 891 1449 895 1453
rect 1506 1449 1510 1453
rect 1514 1449 1518 1453
rect 1522 1449 1526 1453
rect 1530 1449 1534 1453
rect 1538 1449 1542 1453
rect 1546 1449 1550 1453
rect 1557 1449 1561 1453
rect 1574 1449 1578 1453
rect 1591 1449 1595 1453
rect 1600 1449 1604 1453
rect 1613 1449 1617 1453
rect 1621 1449 1625 1453
rect 1629 1449 1633 1453
rect 1646 1449 1650 1453
rect 1656 1449 1660 1453
rect 1664 1449 1668 1453
rect 1704 1449 1708 1453
rect 1719 1449 1723 1453
rect 1809 1449 1813 1453
rect 1824 1449 1828 1453
rect 771 1372 775 1376
rect 786 1372 790 1376
rect 828 1376 832 1380
rect 836 1376 840 1380
rect 852 1372 856 1376
rect 867 1372 871 1376
rect 918 1376 922 1380
rect 926 1376 930 1380
rect 942 1372 946 1376
rect 957 1372 961 1376
rect 801 1368 805 1372
rect 809 1368 813 1372
rect 573 1363 577 1367
rect 581 1363 585 1367
rect 589 1363 593 1367
rect 597 1363 601 1367
rect 605 1363 609 1367
rect 613 1363 617 1367
rect 624 1363 628 1367
rect 641 1363 645 1367
rect 658 1363 662 1367
rect 667 1363 671 1367
rect 680 1363 684 1367
rect 688 1363 692 1367
rect 696 1363 700 1367
rect 713 1363 717 1367
rect 723 1363 727 1367
rect 731 1363 735 1367
rect 882 1368 886 1372
rect 890 1368 894 1372
rect 972 1368 976 1372
rect 980 1368 984 1372
rect 1704 1372 1708 1376
rect 1719 1372 1723 1376
rect 1761 1376 1765 1380
rect 1769 1376 1773 1380
rect 1785 1372 1789 1376
rect 1800 1372 1804 1376
rect 1851 1376 1855 1380
rect 1859 1376 1863 1380
rect 1875 1372 1879 1376
rect 1890 1372 1894 1376
rect 1734 1368 1738 1372
rect 1742 1368 1746 1372
rect 1506 1363 1510 1367
rect 1514 1363 1518 1367
rect 1522 1363 1526 1367
rect 1530 1363 1534 1367
rect 1538 1363 1542 1367
rect 1546 1363 1550 1367
rect 1557 1363 1561 1367
rect 1574 1363 1578 1367
rect 1591 1363 1595 1367
rect 1600 1363 1604 1367
rect 1613 1363 1617 1367
rect 1621 1363 1625 1367
rect 1629 1363 1633 1367
rect 1646 1363 1650 1367
rect 1656 1363 1660 1367
rect 1664 1363 1668 1367
rect 1815 1368 1819 1372
rect 1823 1368 1827 1372
rect 1905 1368 1909 1372
rect 1913 1368 1917 1372
rect 573 1317 577 1321
rect 581 1317 585 1321
rect 589 1317 593 1321
rect 597 1317 601 1321
rect 605 1317 609 1321
rect 613 1317 617 1321
rect 624 1317 628 1321
rect 641 1317 645 1321
rect 658 1317 662 1321
rect 667 1317 671 1321
rect 680 1317 684 1321
rect 688 1317 692 1321
rect 696 1317 700 1321
rect 713 1317 717 1321
rect 723 1317 727 1321
rect 731 1317 735 1321
rect 771 1314 775 1318
rect 786 1314 790 1318
rect 852 1314 856 1318
rect 867 1314 871 1318
rect 942 1314 946 1318
rect 957 1314 961 1318
rect 1506 1317 1510 1321
rect 1514 1317 1518 1321
rect 1522 1317 1526 1321
rect 1530 1317 1534 1321
rect 1538 1317 1542 1321
rect 1546 1317 1550 1321
rect 1557 1317 1561 1321
rect 1574 1317 1578 1321
rect 1591 1317 1595 1321
rect 1600 1317 1604 1321
rect 1613 1317 1617 1321
rect 1621 1317 1625 1321
rect 1629 1317 1633 1321
rect 1646 1317 1650 1321
rect 1656 1317 1660 1321
rect 1664 1317 1668 1321
rect 1704 1314 1708 1318
rect 1719 1314 1723 1318
rect 1785 1314 1789 1318
rect 1800 1314 1804 1318
rect 1875 1314 1879 1318
rect 1890 1314 1894 1318
rect 771 1240 775 1244
rect 786 1240 790 1244
rect 801 1236 805 1240
rect 809 1236 813 1240
rect 573 1231 577 1235
rect 581 1231 585 1235
rect 589 1231 593 1235
rect 597 1231 601 1235
rect 605 1231 609 1235
rect 613 1231 617 1235
rect 624 1231 628 1235
rect 641 1231 645 1235
rect 658 1231 662 1235
rect 667 1231 671 1235
rect 680 1231 684 1235
rect 688 1231 692 1235
rect 696 1231 700 1235
rect 713 1231 717 1235
rect 723 1231 727 1235
rect 731 1231 735 1235
rect 1704 1240 1708 1244
rect 1719 1240 1723 1244
rect 1734 1236 1738 1240
rect 1742 1236 1746 1240
rect 1506 1231 1510 1235
rect 1514 1231 1518 1235
rect 1522 1231 1526 1235
rect 1530 1231 1534 1235
rect 1538 1231 1542 1235
rect 1546 1231 1550 1235
rect 1557 1231 1561 1235
rect 1574 1231 1578 1235
rect 1591 1231 1595 1235
rect 1600 1231 1604 1235
rect 1613 1231 1617 1235
rect 1621 1231 1625 1235
rect 1629 1231 1633 1235
rect 1646 1231 1650 1235
rect 1656 1231 1660 1235
rect 1664 1231 1668 1235
rect 573 1185 577 1189
rect 581 1185 585 1189
rect 589 1185 593 1189
rect 597 1185 601 1189
rect 605 1185 609 1189
rect 613 1185 617 1189
rect 624 1185 628 1189
rect 641 1185 645 1189
rect 658 1185 662 1189
rect 667 1185 671 1189
rect 680 1185 684 1189
rect 688 1185 692 1189
rect 696 1185 700 1189
rect 713 1185 717 1189
rect 723 1185 727 1189
rect 731 1185 735 1189
rect 807 1185 811 1189
rect 815 1185 819 1189
rect 825 1185 829 1189
rect 833 1185 837 1189
rect 842 1185 846 1189
rect 850 1185 854 1189
rect 858 1185 862 1189
rect 866 1185 870 1189
rect 874 1185 878 1189
rect 885 1185 889 1189
rect 902 1185 906 1189
rect 919 1185 923 1189
rect 928 1185 932 1189
rect 941 1185 945 1189
rect 949 1185 953 1189
rect 957 1185 961 1189
rect 974 1185 978 1189
rect 984 1185 988 1189
rect 992 1185 996 1189
rect 96 1171 100 1175
rect 109 1171 113 1175
rect 117 1171 121 1175
rect 125 1171 129 1175
rect 133 1171 137 1175
rect 146 1171 150 1175
rect 159 1171 163 1175
rect 167 1171 171 1175
rect 175 1171 179 1175
rect 183 1171 187 1175
rect 191 1171 195 1175
rect 204 1171 208 1175
rect 212 1171 216 1175
rect 220 1171 224 1175
rect 228 1171 232 1175
rect 241 1171 245 1175
rect 249 1171 253 1175
rect 257 1171 261 1175
rect 265 1171 269 1175
rect 278 1171 282 1175
rect 291 1171 295 1175
rect 299 1171 303 1175
rect 307 1171 311 1175
rect 315 1171 319 1175
rect 323 1171 327 1175
rect 336 1171 340 1175
rect 344 1171 348 1175
rect 352 1171 356 1175
rect 360 1171 364 1175
rect 373 1171 377 1175
rect 381 1171 385 1175
rect 389 1171 393 1175
rect 397 1171 401 1175
rect 410 1171 414 1175
rect 423 1171 427 1175
rect 431 1171 435 1175
rect 439 1171 443 1175
rect 447 1171 451 1175
rect 455 1171 459 1175
rect 468 1171 472 1175
rect 476 1171 480 1175
rect 484 1171 488 1175
rect 771 1178 775 1182
rect 786 1178 790 1182
rect 1506 1185 1510 1189
rect 1514 1185 1518 1189
rect 1522 1185 1526 1189
rect 1530 1185 1534 1189
rect 1538 1185 1542 1189
rect 1546 1185 1550 1189
rect 1557 1185 1561 1189
rect 1574 1185 1578 1189
rect 1591 1185 1595 1189
rect 1600 1185 1604 1189
rect 1613 1185 1617 1189
rect 1621 1185 1625 1189
rect 1629 1185 1633 1189
rect 1646 1185 1650 1189
rect 1656 1185 1660 1189
rect 1664 1185 1668 1189
rect 1740 1185 1744 1189
rect 1748 1185 1752 1189
rect 1758 1185 1762 1189
rect 1766 1185 1770 1189
rect 1775 1185 1779 1189
rect 1783 1185 1787 1189
rect 1791 1185 1795 1189
rect 1799 1185 1803 1189
rect 1807 1185 1811 1189
rect 1818 1185 1822 1189
rect 1835 1185 1839 1189
rect 1852 1185 1856 1189
rect 1861 1185 1865 1189
rect 1874 1185 1878 1189
rect 1882 1185 1886 1189
rect 1890 1185 1894 1189
rect 1907 1185 1911 1189
rect 1917 1185 1921 1189
rect 1925 1185 1929 1189
rect 1029 1171 1033 1175
rect 1042 1171 1046 1175
rect 1050 1171 1054 1175
rect 1058 1171 1062 1175
rect 1066 1171 1070 1175
rect 1079 1171 1083 1175
rect 1092 1171 1096 1175
rect 1100 1171 1104 1175
rect 1108 1171 1112 1175
rect 1116 1171 1120 1175
rect 1124 1171 1128 1175
rect 1137 1171 1141 1175
rect 1145 1171 1149 1175
rect 1153 1171 1157 1175
rect 1161 1171 1165 1175
rect 1174 1171 1178 1175
rect 1182 1171 1186 1175
rect 1190 1171 1194 1175
rect 1198 1171 1202 1175
rect 1211 1171 1215 1175
rect 1224 1171 1228 1175
rect 1232 1171 1236 1175
rect 1240 1171 1244 1175
rect 1248 1171 1252 1175
rect 1256 1171 1260 1175
rect 1269 1171 1273 1175
rect 1277 1171 1281 1175
rect 1285 1171 1289 1175
rect 1293 1171 1297 1175
rect 1306 1171 1310 1175
rect 1314 1171 1318 1175
rect 1322 1171 1326 1175
rect 1330 1171 1334 1175
rect 1343 1171 1347 1175
rect 1356 1171 1360 1175
rect 1364 1171 1368 1175
rect 1372 1171 1376 1175
rect 1380 1171 1384 1175
rect 1388 1171 1392 1175
rect 1401 1171 1405 1175
rect 1409 1171 1413 1175
rect 1417 1171 1421 1175
rect 1704 1178 1708 1182
rect 1719 1178 1723 1182
rect 1001 1132 1005 1136
rect 211 1127 215 1131
rect 219 1127 223 1131
rect 235 1127 239 1131
rect 243 1127 247 1131
rect 1934 1132 1938 1136
rect 1001 1124 1005 1128
rect 1144 1127 1148 1131
rect 1152 1127 1156 1131
rect 1168 1127 1172 1131
rect 1176 1127 1180 1131
rect 1934 1124 1938 1128
rect 231 1116 235 1120
rect 239 1116 243 1120
rect 1164 1116 1168 1120
rect 1172 1116 1176 1120
rect 227 1105 231 1109
rect 1160 1105 1164 1109
rect 227 1097 231 1101
rect 211 1093 215 1097
rect 219 1093 223 1097
rect 235 1093 239 1097
rect 243 1093 247 1097
rect 1160 1097 1164 1101
rect 1144 1093 1148 1097
rect 1152 1093 1156 1097
rect 1168 1093 1172 1097
rect 1176 1093 1180 1097
rect 867 1061 871 1065
rect 880 1061 884 1065
rect 888 1061 892 1065
rect 896 1061 900 1065
rect 904 1061 908 1065
rect 917 1061 921 1065
rect 930 1061 934 1065
rect 938 1061 942 1065
rect 946 1061 950 1065
rect 954 1061 958 1065
rect 962 1061 966 1065
rect 975 1061 979 1065
rect 983 1061 987 1065
rect 991 1061 995 1065
rect 1800 1061 1804 1065
rect 1813 1061 1817 1065
rect 1821 1061 1825 1065
rect 1829 1061 1833 1065
rect 1837 1061 1841 1065
rect 1850 1061 1854 1065
rect 1863 1061 1867 1065
rect 1871 1061 1875 1065
rect 1879 1061 1883 1065
rect 1887 1061 1891 1065
rect 1895 1061 1899 1065
rect 1908 1061 1912 1065
rect 1916 1061 1920 1065
rect 1924 1061 1928 1065
rect 96 1031 100 1035
rect 109 1031 113 1035
rect 117 1031 121 1035
rect 125 1031 129 1035
rect 133 1031 137 1035
rect 146 1031 150 1035
rect 159 1031 163 1035
rect 167 1031 171 1035
rect 175 1031 179 1035
rect 183 1031 187 1035
rect 191 1031 195 1035
rect 204 1031 208 1035
rect 212 1031 216 1035
rect 220 1031 224 1035
rect 228 1031 232 1035
rect 241 1031 245 1035
rect 249 1031 253 1035
rect 257 1031 261 1035
rect 265 1031 269 1035
rect 278 1031 282 1035
rect 291 1031 295 1035
rect 299 1031 303 1035
rect 307 1031 311 1035
rect 315 1031 319 1035
rect 323 1031 327 1035
rect 336 1031 340 1035
rect 344 1031 348 1035
rect 352 1031 356 1035
rect 360 1031 364 1035
rect 373 1031 377 1035
rect 381 1031 385 1035
rect 389 1031 393 1035
rect 397 1031 401 1035
rect 410 1031 414 1035
rect 423 1031 427 1035
rect 431 1031 435 1035
rect 439 1031 443 1035
rect 447 1031 451 1035
rect 455 1031 459 1035
rect 468 1031 472 1035
rect 476 1031 480 1035
rect 484 1031 488 1035
rect 1029 1031 1033 1035
rect 1042 1031 1046 1035
rect 1050 1031 1054 1035
rect 1058 1031 1062 1035
rect 1066 1031 1070 1035
rect 1079 1031 1083 1035
rect 1092 1031 1096 1035
rect 1100 1031 1104 1035
rect 1108 1031 1112 1035
rect 1116 1031 1120 1035
rect 1124 1031 1128 1035
rect 1137 1031 1141 1035
rect 1145 1031 1149 1035
rect 1153 1031 1157 1035
rect 1161 1031 1165 1035
rect 1174 1031 1178 1035
rect 1182 1031 1186 1035
rect 1190 1031 1194 1035
rect 1198 1031 1202 1035
rect 1211 1031 1215 1035
rect 1224 1031 1228 1035
rect 1232 1031 1236 1035
rect 1240 1031 1244 1035
rect 1248 1031 1252 1035
rect 1256 1031 1260 1035
rect 1269 1031 1273 1035
rect 1277 1031 1281 1035
rect 1285 1031 1289 1035
rect 1293 1031 1297 1035
rect 1306 1031 1310 1035
rect 1314 1031 1318 1035
rect 1322 1031 1326 1035
rect 1330 1031 1334 1035
rect 1343 1031 1347 1035
rect 1356 1031 1360 1035
rect 1364 1031 1368 1035
rect 1372 1031 1376 1035
rect 1380 1031 1384 1035
rect 1388 1031 1392 1035
rect 1401 1031 1405 1035
rect 1409 1031 1413 1035
rect 1417 1031 1421 1035
rect 1013 988 1017 992
rect 1013 980 1017 984
rect 1946 988 1950 992
rect 1946 980 1950 984
rect 867 975 871 979
rect 880 975 884 979
rect 888 975 892 979
rect 896 975 900 979
rect 904 975 908 979
rect 917 975 921 979
rect 930 975 934 979
rect 938 975 942 979
rect 946 975 950 979
rect 954 975 958 979
rect 962 975 966 979
rect 975 975 979 979
rect 983 975 987 979
rect 991 975 995 979
rect 1800 975 1804 979
rect 1813 975 1817 979
rect 1821 975 1825 979
rect 1829 975 1833 979
rect 1837 975 1841 979
rect 1850 975 1854 979
rect 1863 975 1867 979
rect 1871 975 1875 979
rect 1879 975 1883 979
rect 1887 975 1891 979
rect 1895 975 1899 979
rect 1908 975 1912 979
rect 1916 975 1920 979
rect 1924 975 1928 979
rect 96 945 100 949
rect 109 945 113 949
rect 117 945 121 949
rect 125 945 129 949
rect 133 945 137 949
rect 146 945 150 949
rect 159 945 163 949
rect 167 945 171 949
rect 175 945 179 949
rect 183 945 187 949
rect 191 945 195 949
rect 204 945 208 949
rect 212 945 216 949
rect 220 945 224 949
rect 228 945 232 949
rect 241 945 245 949
rect 249 945 253 949
rect 257 945 261 949
rect 265 945 269 949
rect 278 945 282 949
rect 291 945 295 949
rect 299 945 303 949
rect 307 945 311 949
rect 315 945 319 949
rect 323 945 327 949
rect 336 945 340 949
rect 344 945 348 949
rect 352 945 356 949
rect 360 945 364 949
rect 373 945 377 949
rect 381 945 385 949
rect 389 945 393 949
rect 397 945 401 949
rect 410 945 414 949
rect 423 945 427 949
rect 431 945 435 949
rect 439 945 443 949
rect 447 945 451 949
rect 455 945 459 949
rect 468 945 472 949
rect 476 945 480 949
rect 484 945 488 949
rect 1029 945 1033 949
rect 1042 945 1046 949
rect 1050 945 1054 949
rect 1058 945 1062 949
rect 1066 945 1070 949
rect 1079 945 1083 949
rect 1092 945 1096 949
rect 1100 945 1104 949
rect 1108 945 1112 949
rect 1116 945 1120 949
rect 1124 945 1128 949
rect 1137 945 1141 949
rect 1145 945 1149 949
rect 1153 945 1157 949
rect 1161 945 1165 949
rect 1174 945 1178 949
rect 1182 945 1186 949
rect 1190 945 1194 949
rect 1198 945 1202 949
rect 1211 945 1215 949
rect 1224 945 1228 949
rect 1232 945 1236 949
rect 1240 945 1244 949
rect 1248 945 1252 949
rect 1256 945 1260 949
rect 1269 945 1273 949
rect 1277 945 1281 949
rect 1285 945 1289 949
rect 1293 945 1297 949
rect 1306 945 1310 949
rect 1314 945 1318 949
rect 1322 945 1326 949
rect 1330 945 1334 949
rect 1343 945 1347 949
rect 1356 945 1360 949
rect 1364 945 1368 949
rect 1372 945 1376 949
rect 1380 945 1384 949
rect 1388 945 1392 949
rect 1401 945 1405 949
rect 1409 945 1413 949
rect 1417 945 1421 949
rect 328 901 332 905
rect 336 901 340 905
rect 352 901 356 905
rect 360 901 364 905
rect 1261 901 1265 905
rect 1269 901 1273 905
rect 1285 901 1289 905
rect 1293 901 1297 905
rect 348 890 352 894
rect 356 890 360 894
rect 1281 890 1285 894
rect 1289 890 1293 894
rect 344 879 348 883
rect 1277 879 1281 883
rect 344 871 348 875
rect 1277 871 1281 875
rect 328 867 332 871
rect 336 867 340 871
rect 352 867 356 871
rect 360 867 364 871
rect 1261 867 1265 871
rect 1269 867 1273 871
rect 1285 867 1289 871
rect 1293 867 1297 871
rect 96 805 100 809
rect 109 805 113 809
rect 117 805 121 809
rect 125 805 129 809
rect 133 805 137 809
rect 146 805 150 809
rect 159 805 163 809
rect 167 805 171 809
rect 175 805 179 809
rect 183 805 187 809
rect 191 805 195 809
rect 204 805 208 809
rect 212 805 216 809
rect 220 805 224 809
rect 228 805 232 809
rect 241 805 245 809
rect 249 805 253 809
rect 257 805 261 809
rect 265 805 269 809
rect 278 805 282 809
rect 291 805 295 809
rect 299 805 303 809
rect 307 805 311 809
rect 315 805 319 809
rect 323 805 327 809
rect 336 805 340 809
rect 344 805 348 809
rect 352 805 356 809
rect 360 805 364 809
rect 373 805 377 809
rect 381 805 385 809
rect 389 805 393 809
rect 397 805 401 809
rect 410 805 414 809
rect 423 805 427 809
rect 431 805 435 809
rect 439 805 443 809
rect 447 805 451 809
rect 455 805 459 809
rect 468 805 472 809
rect 476 805 480 809
rect 484 805 488 809
rect 1029 805 1033 809
rect 1042 805 1046 809
rect 1050 805 1054 809
rect 1058 805 1062 809
rect 1066 805 1070 809
rect 1079 805 1083 809
rect 1092 805 1096 809
rect 1100 805 1104 809
rect 1108 805 1112 809
rect 1116 805 1120 809
rect 1124 805 1128 809
rect 1137 805 1141 809
rect 1145 805 1149 809
rect 1153 805 1157 809
rect 1161 805 1165 809
rect 1174 805 1178 809
rect 1182 805 1186 809
rect 1190 805 1194 809
rect 1198 805 1202 809
rect 1211 805 1215 809
rect 1224 805 1228 809
rect 1232 805 1236 809
rect 1240 805 1244 809
rect 1248 805 1252 809
rect 1256 805 1260 809
rect 1269 805 1273 809
rect 1277 805 1281 809
rect 1285 805 1289 809
rect 1293 805 1297 809
rect 1306 805 1310 809
rect 1314 805 1318 809
rect 1322 805 1326 809
rect 1330 805 1334 809
rect 1343 805 1347 809
rect 1356 805 1360 809
rect 1364 805 1368 809
rect 1372 805 1376 809
rect 1380 805 1384 809
rect 1388 805 1392 809
rect 1401 805 1405 809
rect 1409 805 1413 809
rect 1417 805 1421 809
rect 568 726 572 730
rect 581 726 585 730
rect 589 726 593 730
rect 597 726 601 730
rect 605 726 609 730
rect 618 726 622 730
rect 631 726 635 730
rect 639 726 643 730
rect 647 726 651 730
rect 655 726 659 730
rect 663 726 667 730
rect 676 726 680 730
rect 684 726 688 730
rect 692 726 696 730
rect 700 726 704 730
rect 713 726 717 730
rect 721 726 725 730
rect 729 726 733 730
rect 737 726 741 730
rect 750 726 754 730
rect 763 726 767 730
rect 771 726 775 730
rect 779 726 783 730
rect 787 726 791 730
rect 795 726 799 730
rect 808 726 812 730
rect 816 726 820 730
rect 824 726 828 730
rect 832 726 836 730
rect 845 726 849 730
rect 853 726 857 730
rect 861 726 865 730
rect 869 726 873 730
rect 882 726 886 730
rect 895 726 899 730
rect 903 726 907 730
rect 911 726 915 730
rect 919 726 923 730
rect 927 726 931 730
rect 940 726 944 730
rect 948 726 952 730
rect 956 726 960 730
rect 964 726 968 730
rect 977 726 981 730
rect 985 726 989 730
rect 993 726 997 730
rect 1001 726 1005 730
rect 1014 726 1018 730
rect 1027 726 1031 730
rect 1035 726 1039 730
rect 1043 726 1047 730
rect 1051 726 1055 730
rect 1059 726 1063 730
rect 1072 726 1076 730
rect 1080 726 1084 730
rect 1088 726 1092 730
rect 1501 726 1505 730
rect 1514 726 1518 730
rect 1522 726 1526 730
rect 1530 726 1534 730
rect 1538 726 1542 730
rect 1551 726 1555 730
rect 1564 726 1568 730
rect 1572 726 1576 730
rect 1580 726 1584 730
rect 1588 726 1592 730
rect 1596 726 1600 730
rect 1609 726 1613 730
rect 1617 726 1621 730
rect 1625 726 1629 730
rect 1633 726 1637 730
rect 1646 726 1650 730
rect 1654 726 1658 730
rect 1662 726 1666 730
rect 1670 726 1674 730
rect 1683 726 1687 730
rect 1696 726 1700 730
rect 1704 726 1708 730
rect 1712 726 1716 730
rect 1720 726 1724 730
rect 1728 726 1732 730
rect 1741 726 1745 730
rect 1749 726 1753 730
rect 1757 726 1761 730
rect 1765 726 1769 730
rect 1778 726 1782 730
rect 1786 726 1790 730
rect 1794 726 1798 730
rect 1802 726 1806 730
rect 1815 726 1819 730
rect 1828 726 1832 730
rect 1836 726 1840 730
rect 1844 726 1848 730
rect 1852 726 1856 730
rect 1860 726 1864 730
rect 1873 726 1877 730
rect 1881 726 1885 730
rect 1889 726 1893 730
rect 1897 726 1901 730
rect 1910 726 1914 730
rect 1918 726 1922 730
rect 1926 726 1930 730
rect 1934 726 1938 730
rect 1947 726 1951 730
rect 1960 726 1964 730
rect 1968 726 1972 730
rect 1976 726 1980 730
rect 1984 726 1988 730
rect 1992 726 1996 730
rect 2005 726 2009 730
rect 2013 726 2017 730
rect 2021 726 2025 730
rect 228 693 232 697
rect 241 693 245 697
rect 249 693 253 697
rect 257 693 261 697
rect 265 693 269 697
rect 278 693 282 697
rect 291 693 295 697
rect 299 693 303 697
rect 307 693 311 697
rect 315 693 319 697
rect 323 693 327 697
rect 336 693 340 697
rect 344 693 348 697
rect 352 693 356 697
rect 1161 693 1165 697
rect 1174 693 1178 697
rect 1182 693 1186 697
rect 1190 693 1194 697
rect 1198 693 1202 697
rect 1211 693 1215 697
rect 1224 693 1228 697
rect 1232 693 1236 697
rect 1240 693 1244 697
rect 1248 693 1252 697
rect 1256 693 1260 697
rect 1269 693 1273 697
rect 1277 693 1281 697
rect 1285 693 1289 697
rect 352 656 356 660
rect 360 656 364 660
rect 747 660 751 664
rect 755 660 759 664
rect 771 656 775 660
rect 786 656 790 660
rect 828 660 832 664
rect 836 660 840 664
rect 852 656 856 660
rect 867 656 871 660
rect 801 652 805 656
rect 809 652 813 656
rect 235 647 239 651
rect 243 647 247 651
rect 573 647 577 651
rect 581 647 585 651
rect 589 647 593 651
rect 597 647 601 651
rect 605 647 609 651
rect 613 647 617 651
rect 624 647 628 651
rect 641 647 645 651
rect 658 647 662 651
rect 667 647 671 651
rect 680 647 684 651
rect 688 647 692 651
rect 696 647 700 651
rect 713 647 717 651
rect 723 647 727 651
rect 731 647 735 651
rect 882 652 886 656
rect 890 652 894 656
rect 1285 656 1289 660
rect 1293 656 1297 660
rect 1680 660 1684 664
rect 1688 660 1692 664
rect 1704 656 1708 660
rect 1719 656 1723 660
rect 1761 660 1765 664
rect 1769 660 1773 664
rect 1785 656 1789 660
rect 1800 656 1804 660
rect 1734 652 1738 656
rect 1742 652 1746 656
rect 1168 647 1172 651
rect 1176 647 1180 651
rect 1506 647 1510 651
rect 1514 647 1518 651
rect 1522 647 1526 651
rect 1530 647 1534 651
rect 1538 647 1542 651
rect 1546 647 1550 651
rect 1557 647 1561 651
rect 1574 647 1578 651
rect 1591 647 1595 651
rect 1600 647 1604 651
rect 1613 647 1617 651
rect 1621 647 1625 651
rect 1629 647 1633 651
rect 1646 647 1650 651
rect 1656 647 1660 651
rect 1664 647 1668 651
rect 1815 652 1819 656
rect 1823 652 1827 656
rect 573 601 577 605
rect 581 601 585 605
rect 589 601 593 605
rect 597 601 601 605
rect 605 601 609 605
rect 613 601 617 605
rect 624 601 628 605
rect 641 601 645 605
rect 658 601 662 605
rect 667 601 671 605
rect 680 601 684 605
rect 688 601 692 605
rect 696 601 700 605
rect 713 601 717 605
rect 723 601 727 605
rect 731 601 735 605
rect 219 591 223 595
rect 227 591 231 595
rect 235 591 239 595
rect 248 591 252 595
rect 256 591 260 595
rect 264 591 268 595
rect 272 591 276 595
rect 280 591 284 595
rect 293 591 297 595
rect 306 591 310 595
rect 314 591 318 595
rect 322 591 326 595
rect 330 591 334 595
rect 343 591 347 595
rect 771 600 775 604
rect 786 600 790 604
rect 852 600 856 604
rect 867 600 871 604
rect 1506 601 1510 605
rect 1514 601 1518 605
rect 1522 601 1526 605
rect 1530 601 1534 605
rect 1538 601 1542 605
rect 1546 601 1550 605
rect 1557 601 1561 605
rect 1574 601 1578 605
rect 1591 601 1595 605
rect 1600 601 1604 605
rect 1613 601 1617 605
rect 1621 601 1625 605
rect 1629 601 1633 605
rect 1646 601 1650 605
rect 1656 601 1660 605
rect 1664 601 1668 605
rect 1152 591 1156 595
rect 1160 591 1164 595
rect 1168 591 1172 595
rect 1181 591 1185 595
rect 1189 591 1193 595
rect 1197 591 1201 595
rect 1205 591 1209 595
rect 1213 591 1217 595
rect 1226 591 1230 595
rect 1239 591 1243 595
rect 1247 591 1251 595
rect 1255 591 1259 595
rect 1263 591 1267 595
rect 1276 591 1280 595
rect 1704 600 1708 604
rect 1719 600 1723 604
rect 1785 600 1789 604
rect 1800 600 1804 604
rect 771 524 775 528
rect 786 524 790 528
rect 852 528 856 532
rect 860 528 864 532
rect 876 524 880 528
rect 891 524 895 528
rect 801 520 805 524
rect 809 520 813 524
rect 573 515 577 519
rect 581 515 585 519
rect 589 515 593 519
rect 597 515 601 519
rect 605 515 609 519
rect 613 515 617 519
rect 624 515 628 519
rect 641 515 645 519
rect 658 515 662 519
rect 667 515 671 519
rect 680 515 684 519
rect 688 515 692 519
rect 696 515 700 519
rect 713 515 717 519
rect 723 515 727 519
rect 731 515 735 519
rect 906 520 910 524
rect 914 520 918 524
rect 1704 524 1708 528
rect 1719 524 1723 528
rect 1785 528 1789 532
rect 1793 528 1797 532
rect 1809 524 1813 528
rect 1824 524 1828 528
rect 1734 520 1738 524
rect 1742 520 1746 524
rect 1506 515 1510 519
rect 1514 515 1518 519
rect 1522 515 1526 519
rect 1530 515 1534 519
rect 1538 515 1542 519
rect 1546 515 1550 519
rect 1557 515 1561 519
rect 1574 515 1578 519
rect 1591 515 1595 519
rect 1600 515 1604 519
rect 1613 515 1617 519
rect 1621 515 1625 519
rect 1629 515 1633 519
rect 1646 515 1650 519
rect 1656 515 1660 519
rect 1664 515 1668 519
rect 1839 520 1843 524
rect 1847 520 1851 524
rect 573 469 577 473
rect 581 469 585 473
rect 589 469 593 473
rect 597 469 601 473
rect 605 469 609 473
rect 613 469 617 473
rect 624 469 628 473
rect 641 469 645 473
rect 658 469 662 473
rect 667 469 671 473
rect 680 469 684 473
rect 688 469 692 473
rect 696 469 700 473
rect 713 469 717 473
rect 723 469 727 473
rect 731 469 735 473
rect 771 469 775 473
rect 786 469 790 473
rect 876 469 880 473
rect 891 469 895 473
rect 1506 469 1510 473
rect 1514 469 1518 473
rect 1522 469 1526 473
rect 1530 469 1534 473
rect 1538 469 1542 473
rect 1546 469 1550 473
rect 1557 469 1561 473
rect 1574 469 1578 473
rect 1591 469 1595 473
rect 1600 469 1604 473
rect 1613 469 1617 473
rect 1621 469 1625 473
rect 1629 469 1633 473
rect 1646 469 1650 473
rect 1656 469 1660 473
rect 1664 469 1668 473
rect 1704 469 1708 473
rect 1719 469 1723 473
rect 1809 469 1813 473
rect 1824 469 1828 473
rect 771 392 775 396
rect 786 392 790 396
rect 828 396 832 400
rect 836 396 840 400
rect 852 392 856 396
rect 867 392 871 396
rect 918 396 922 400
rect 926 396 930 400
rect 942 392 946 396
rect 957 392 961 396
rect 801 388 805 392
rect 809 388 813 392
rect 573 383 577 387
rect 581 383 585 387
rect 589 383 593 387
rect 597 383 601 387
rect 605 383 609 387
rect 613 383 617 387
rect 624 383 628 387
rect 641 383 645 387
rect 658 383 662 387
rect 667 383 671 387
rect 680 383 684 387
rect 688 383 692 387
rect 696 383 700 387
rect 713 383 717 387
rect 723 383 727 387
rect 731 383 735 387
rect 882 388 886 392
rect 890 388 894 392
rect 972 388 976 392
rect 980 388 984 392
rect 1704 392 1708 396
rect 1719 392 1723 396
rect 1761 396 1765 400
rect 1769 396 1773 400
rect 1785 392 1789 396
rect 1800 392 1804 396
rect 1851 396 1855 400
rect 1859 396 1863 400
rect 1875 392 1879 396
rect 1890 392 1894 396
rect 1734 388 1738 392
rect 1742 388 1746 392
rect 1506 383 1510 387
rect 1514 383 1518 387
rect 1522 383 1526 387
rect 1530 383 1534 387
rect 1538 383 1542 387
rect 1546 383 1550 387
rect 1557 383 1561 387
rect 1574 383 1578 387
rect 1591 383 1595 387
rect 1600 383 1604 387
rect 1613 383 1617 387
rect 1621 383 1625 387
rect 1629 383 1633 387
rect 1646 383 1650 387
rect 1656 383 1660 387
rect 1664 383 1668 387
rect 1815 388 1819 392
rect 1823 388 1827 392
rect 1905 388 1909 392
rect 1913 388 1917 392
rect 573 337 577 341
rect 581 337 585 341
rect 589 337 593 341
rect 597 337 601 341
rect 605 337 609 341
rect 613 337 617 341
rect 624 337 628 341
rect 641 337 645 341
rect 658 337 662 341
rect 667 337 671 341
rect 680 337 684 341
rect 688 337 692 341
rect 696 337 700 341
rect 713 337 717 341
rect 723 337 727 341
rect 731 337 735 341
rect 771 334 775 338
rect 786 334 790 338
rect 852 334 856 338
rect 867 334 871 338
rect 942 334 946 338
rect 957 334 961 338
rect 1506 337 1510 341
rect 1514 337 1518 341
rect 1522 337 1526 341
rect 1530 337 1534 341
rect 1538 337 1542 341
rect 1546 337 1550 341
rect 1557 337 1561 341
rect 1574 337 1578 341
rect 1591 337 1595 341
rect 1600 337 1604 341
rect 1613 337 1617 341
rect 1621 337 1625 341
rect 1629 337 1633 341
rect 1646 337 1650 341
rect 1656 337 1660 341
rect 1664 337 1668 341
rect 1704 334 1708 338
rect 1719 334 1723 338
rect 1785 334 1789 338
rect 1800 334 1804 338
rect 1875 334 1879 338
rect 1890 334 1894 338
rect 771 260 775 264
rect 786 260 790 264
rect 801 256 805 260
rect 809 256 813 260
rect 573 251 577 255
rect 581 251 585 255
rect 589 251 593 255
rect 597 251 601 255
rect 605 251 609 255
rect 613 251 617 255
rect 624 251 628 255
rect 641 251 645 255
rect 658 251 662 255
rect 667 251 671 255
rect 680 251 684 255
rect 688 251 692 255
rect 696 251 700 255
rect 713 251 717 255
rect 723 251 727 255
rect 731 251 735 255
rect 1704 260 1708 264
rect 1719 260 1723 264
rect 1734 256 1738 260
rect 1742 256 1746 260
rect 1506 251 1510 255
rect 1514 251 1518 255
rect 1522 251 1526 255
rect 1530 251 1534 255
rect 1538 251 1542 255
rect 1546 251 1550 255
rect 1557 251 1561 255
rect 1574 251 1578 255
rect 1591 251 1595 255
rect 1600 251 1604 255
rect 1613 251 1617 255
rect 1621 251 1625 255
rect 1629 251 1633 255
rect 1646 251 1650 255
rect 1656 251 1660 255
rect 1664 251 1668 255
rect 573 205 577 209
rect 581 205 585 209
rect 589 205 593 209
rect 597 205 601 209
rect 605 205 609 209
rect 613 205 617 209
rect 624 205 628 209
rect 641 205 645 209
rect 658 205 662 209
rect 667 205 671 209
rect 680 205 684 209
rect 688 205 692 209
rect 696 205 700 209
rect 713 205 717 209
rect 723 205 727 209
rect 731 205 735 209
rect 807 205 811 209
rect 815 205 819 209
rect 825 205 829 209
rect 833 205 837 209
rect 842 205 846 209
rect 850 205 854 209
rect 858 205 862 209
rect 866 205 870 209
rect 874 205 878 209
rect 885 205 889 209
rect 902 205 906 209
rect 919 205 923 209
rect 928 205 932 209
rect 941 205 945 209
rect 949 205 953 209
rect 957 205 961 209
rect 974 205 978 209
rect 984 205 988 209
rect 992 205 996 209
rect 96 191 100 195
rect 109 191 113 195
rect 117 191 121 195
rect 125 191 129 195
rect 133 191 137 195
rect 146 191 150 195
rect 159 191 163 195
rect 167 191 171 195
rect 175 191 179 195
rect 183 191 187 195
rect 191 191 195 195
rect 204 191 208 195
rect 212 191 216 195
rect 220 191 224 195
rect 228 191 232 195
rect 241 191 245 195
rect 249 191 253 195
rect 257 191 261 195
rect 265 191 269 195
rect 278 191 282 195
rect 291 191 295 195
rect 299 191 303 195
rect 307 191 311 195
rect 315 191 319 195
rect 323 191 327 195
rect 336 191 340 195
rect 344 191 348 195
rect 352 191 356 195
rect 360 191 364 195
rect 373 191 377 195
rect 381 191 385 195
rect 389 191 393 195
rect 397 191 401 195
rect 410 191 414 195
rect 423 191 427 195
rect 431 191 435 195
rect 439 191 443 195
rect 447 191 451 195
rect 455 191 459 195
rect 468 191 472 195
rect 476 191 480 195
rect 484 191 488 195
rect 771 198 775 202
rect 786 198 790 202
rect 1506 205 1510 209
rect 1514 205 1518 209
rect 1522 205 1526 209
rect 1530 205 1534 209
rect 1538 205 1542 209
rect 1546 205 1550 209
rect 1557 205 1561 209
rect 1574 205 1578 209
rect 1591 205 1595 209
rect 1600 205 1604 209
rect 1613 205 1617 209
rect 1621 205 1625 209
rect 1629 205 1633 209
rect 1646 205 1650 209
rect 1656 205 1660 209
rect 1664 205 1668 209
rect 1740 205 1744 209
rect 1748 205 1752 209
rect 1758 205 1762 209
rect 1766 205 1770 209
rect 1775 205 1779 209
rect 1783 205 1787 209
rect 1791 205 1795 209
rect 1799 205 1803 209
rect 1807 205 1811 209
rect 1818 205 1822 209
rect 1835 205 1839 209
rect 1852 205 1856 209
rect 1861 205 1865 209
rect 1874 205 1878 209
rect 1882 205 1886 209
rect 1890 205 1894 209
rect 1907 205 1911 209
rect 1917 205 1921 209
rect 1925 205 1929 209
rect 1029 191 1033 195
rect 1042 191 1046 195
rect 1050 191 1054 195
rect 1058 191 1062 195
rect 1066 191 1070 195
rect 1079 191 1083 195
rect 1092 191 1096 195
rect 1100 191 1104 195
rect 1108 191 1112 195
rect 1116 191 1120 195
rect 1124 191 1128 195
rect 1137 191 1141 195
rect 1145 191 1149 195
rect 1153 191 1157 195
rect 1161 191 1165 195
rect 1174 191 1178 195
rect 1182 191 1186 195
rect 1190 191 1194 195
rect 1198 191 1202 195
rect 1211 191 1215 195
rect 1224 191 1228 195
rect 1232 191 1236 195
rect 1240 191 1244 195
rect 1248 191 1252 195
rect 1256 191 1260 195
rect 1269 191 1273 195
rect 1277 191 1281 195
rect 1285 191 1289 195
rect 1293 191 1297 195
rect 1306 191 1310 195
rect 1314 191 1318 195
rect 1322 191 1326 195
rect 1330 191 1334 195
rect 1343 191 1347 195
rect 1356 191 1360 195
rect 1364 191 1368 195
rect 1372 191 1376 195
rect 1380 191 1384 195
rect 1388 191 1392 195
rect 1401 191 1405 195
rect 1409 191 1413 195
rect 1417 191 1421 195
rect 1704 198 1708 202
rect 1719 198 1723 202
rect 1001 152 1005 156
rect 211 147 215 151
rect 219 147 223 151
rect 235 147 239 151
rect 243 147 247 151
rect 1934 152 1938 156
rect 1001 144 1005 148
rect 1144 147 1148 151
rect 1152 147 1156 151
rect 1168 147 1172 151
rect 1176 147 1180 151
rect 1934 144 1938 148
rect 231 136 235 140
rect 239 136 243 140
rect 1164 136 1168 140
rect 1172 136 1176 140
rect 227 125 231 129
rect 1160 125 1164 129
rect 227 117 231 121
rect 211 113 215 117
rect 219 113 223 117
rect 235 113 239 117
rect 243 113 247 117
rect 1160 117 1164 121
rect 1144 113 1148 117
rect 1152 113 1156 117
rect 1168 113 1172 117
rect 1176 113 1180 117
rect 867 81 871 85
rect 880 81 884 85
rect 888 81 892 85
rect 896 81 900 85
rect 904 81 908 85
rect 917 81 921 85
rect 930 81 934 85
rect 938 81 942 85
rect 946 81 950 85
rect 954 81 958 85
rect 962 81 966 85
rect 975 81 979 85
rect 983 81 987 85
rect 991 81 995 85
rect 1800 81 1804 85
rect 1813 81 1817 85
rect 1821 81 1825 85
rect 1829 81 1833 85
rect 1837 81 1841 85
rect 1850 81 1854 85
rect 1863 81 1867 85
rect 1871 81 1875 85
rect 1879 81 1883 85
rect 1887 81 1891 85
rect 1895 81 1899 85
rect 1908 81 1912 85
rect 1916 81 1920 85
rect 1924 81 1928 85
rect 96 51 100 55
rect 109 51 113 55
rect 117 51 121 55
rect 125 51 129 55
rect 133 51 137 55
rect 146 51 150 55
rect 159 51 163 55
rect 167 51 171 55
rect 175 51 179 55
rect 183 51 187 55
rect 191 51 195 55
rect 204 51 208 55
rect 212 51 216 55
rect 220 51 224 55
rect 228 51 232 55
rect 241 51 245 55
rect 249 51 253 55
rect 257 51 261 55
rect 265 51 269 55
rect 278 51 282 55
rect 291 51 295 55
rect 299 51 303 55
rect 307 51 311 55
rect 315 51 319 55
rect 323 51 327 55
rect 336 51 340 55
rect 344 51 348 55
rect 352 51 356 55
rect 360 51 364 55
rect 373 51 377 55
rect 381 51 385 55
rect 389 51 393 55
rect 397 51 401 55
rect 410 51 414 55
rect 423 51 427 55
rect 431 51 435 55
rect 439 51 443 55
rect 447 51 451 55
rect 455 51 459 55
rect 468 51 472 55
rect 476 51 480 55
rect 484 51 488 55
rect 1029 51 1033 55
rect 1042 51 1046 55
rect 1050 51 1054 55
rect 1058 51 1062 55
rect 1066 51 1070 55
rect 1079 51 1083 55
rect 1092 51 1096 55
rect 1100 51 1104 55
rect 1108 51 1112 55
rect 1116 51 1120 55
rect 1124 51 1128 55
rect 1137 51 1141 55
rect 1145 51 1149 55
rect 1153 51 1157 55
rect 1161 51 1165 55
rect 1174 51 1178 55
rect 1182 51 1186 55
rect 1190 51 1194 55
rect 1198 51 1202 55
rect 1211 51 1215 55
rect 1224 51 1228 55
rect 1232 51 1236 55
rect 1240 51 1244 55
rect 1248 51 1252 55
rect 1256 51 1260 55
rect 1269 51 1273 55
rect 1277 51 1281 55
rect 1285 51 1289 55
rect 1293 51 1297 55
rect 1306 51 1310 55
rect 1314 51 1318 55
rect 1322 51 1326 55
rect 1330 51 1334 55
rect 1343 51 1347 55
rect 1356 51 1360 55
rect 1364 51 1368 55
rect 1372 51 1376 55
rect 1380 51 1384 55
rect 1388 51 1392 55
rect 1401 51 1405 55
rect 1409 51 1413 55
rect 1417 51 1421 55
rect 1013 8 1017 12
rect 1013 0 1017 4
rect 1946 8 1950 12
rect 1946 0 1950 4
rect 867 -5 871 -1
rect 880 -5 884 -1
rect 888 -5 892 -1
rect 896 -5 900 -1
rect 904 -5 908 -1
rect 917 -5 921 -1
rect 930 -5 934 -1
rect 938 -5 942 -1
rect 946 -5 950 -1
rect 954 -5 958 -1
rect 962 -5 966 -1
rect 975 -5 979 -1
rect 983 -5 987 -1
rect 991 -5 995 -1
rect 1800 -5 1804 -1
rect 1813 -5 1817 -1
rect 1821 -5 1825 -1
rect 1829 -5 1833 -1
rect 1837 -5 1841 -1
rect 1850 -5 1854 -1
rect 1863 -5 1867 -1
rect 1871 -5 1875 -1
rect 1879 -5 1883 -1
rect 1887 -5 1891 -1
rect 1895 -5 1899 -1
rect 1908 -5 1912 -1
rect 1916 -5 1920 -1
rect 1924 -5 1928 -1
rect 96 -35 100 -31
rect 109 -35 113 -31
rect 117 -35 121 -31
rect 125 -35 129 -31
rect 133 -35 137 -31
rect 146 -35 150 -31
rect 159 -35 163 -31
rect 167 -35 171 -31
rect 175 -35 179 -31
rect 183 -35 187 -31
rect 191 -35 195 -31
rect 204 -35 208 -31
rect 212 -35 216 -31
rect 220 -35 224 -31
rect 228 -35 232 -31
rect 241 -35 245 -31
rect 249 -35 253 -31
rect 257 -35 261 -31
rect 265 -35 269 -31
rect 278 -35 282 -31
rect 291 -35 295 -31
rect 299 -35 303 -31
rect 307 -35 311 -31
rect 315 -35 319 -31
rect 323 -35 327 -31
rect 336 -35 340 -31
rect 344 -35 348 -31
rect 352 -35 356 -31
rect 360 -35 364 -31
rect 373 -35 377 -31
rect 381 -35 385 -31
rect 389 -35 393 -31
rect 397 -35 401 -31
rect 410 -35 414 -31
rect 423 -35 427 -31
rect 431 -35 435 -31
rect 439 -35 443 -31
rect 447 -35 451 -31
rect 455 -35 459 -31
rect 468 -35 472 -31
rect 476 -35 480 -31
rect 484 -35 488 -31
rect 1029 -35 1033 -31
rect 1042 -35 1046 -31
rect 1050 -35 1054 -31
rect 1058 -35 1062 -31
rect 1066 -35 1070 -31
rect 1079 -35 1083 -31
rect 1092 -35 1096 -31
rect 1100 -35 1104 -31
rect 1108 -35 1112 -31
rect 1116 -35 1120 -31
rect 1124 -35 1128 -31
rect 1137 -35 1141 -31
rect 1145 -35 1149 -31
rect 1153 -35 1157 -31
rect 1161 -35 1165 -31
rect 1174 -35 1178 -31
rect 1182 -35 1186 -31
rect 1190 -35 1194 -31
rect 1198 -35 1202 -31
rect 1211 -35 1215 -31
rect 1224 -35 1228 -31
rect 1232 -35 1236 -31
rect 1240 -35 1244 -31
rect 1248 -35 1252 -31
rect 1256 -35 1260 -31
rect 1269 -35 1273 -31
rect 1277 -35 1281 -31
rect 1285 -35 1289 -31
rect 1293 -35 1297 -31
rect 1306 -35 1310 -31
rect 1314 -35 1318 -31
rect 1322 -35 1326 -31
rect 1330 -35 1334 -31
rect 1343 -35 1347 -31
rect 1356 -35 1360 -31
rect 1364 -35 1368 -31
rect 1372 -35 1376 -31
rect 1380 -35 1384 -31
rect 1388 -35 1392 -31
rect 1401 -35 1405 -31
rect 1409 -35 1413 -31
rect 1417 -35 1421 -31
rect 328 -79 332 -75
rect 336 -79 340 -75
rect 352 -79 356 -75
rect 360 -79 364 -75
rect 1261 -79 1265 -75
rect 1269 -79 1273 -75
rect 1285 -79 1289 -75
rect 1293 -79 1297 -75
rect 348 -90 352 -86
rect 356 -90 360 -86
rect 1281 -90 1285 -86
rect 1289 -90 1293 -86
rect 344 -101 348 -97
rect 1277 -101 1281 -97
rect 344 -109 348 -105
rect 1277 -109 1281 -105
rect 328 -113 332 -109
rect 336 -113 340 -109
rect 352 -113 356 -109
rect 360 -113 364 -109
rect 1261 -113 1265 -109
rect 1269 -113 1273 -109
rect 1285 -113 1289 -109
rect 1293 -113 1297 -109
rect 96 -175 100 -171
rect 109 -175 113 -171
rect 117 -175 121 -171
rect 125 -175 129 -171
rect 133 -175 137 -171
rect 146 -175 150 -171
rect 159 -175 163 -171
rect 167 -175 171 -171
rect 175 -175 179 -171
rect 183 -175 187 -171
rect 191 -175 195 -171
rect 204 -175 208 -171
rect 212 -175 216 -171
rect 220 -175 224 -171
rect 228 -175 232 -171
rect 241 -175 245 -171
rect 249 -175 253 -171
rect 257 -175 261 -171
rect 265 -175 269 -171
rect 278 -175 282 -171
rect 291 -175 295 -171
rect 299 -175 303 -171
rect 307 -175 311 -171
rect 315 -175 319 -171
rect 323 -175 327 -171
rect 336 -175 340 -171
rect 344 -175 348 -171
rect 352 -175 356 -171
rect 360 -175 364 -171
rect 373 -175 377 -171
rect 381 -175 385 -171
rect 389 -175 393 -171
rect 397 -175 401 -171
rect 410 -175 414 -171
rect 423 -175 427 -171
rect 431 -175 435 -171
rect 439 -175 443 -171
rect 447 -175 451 -171
rect 455 -175 459 -171
rect 468 -175 472 -171
rect 476 -175 480 -171
rect 484 -175 488 -171
rect 1029 -175 1033 -171
rect 1042 -175 1046 -171
rect 1050 -175 1054 -171
rect 1058 -175 1062 -171
rect 1066 -175 1070 -171
rect 1079 -175 1083 -171
rect 1092 -175 1096 -171
rect 1100 -175 1104 -171
rect 1108 -175 1112 -171
rect 1116 -175 1120 -171
rect 1124 -175 1128 -171
rect 1137 -175 1141 -171
rect 1145 -175 1149 -171
rect 1153 -175 1157 -171
rect 1161 -175 1165 -171
rect 1174 -175 1178 -171
rect 1182 -175 1186 -171
rect 1190 -175 1194 -171
rect 1198 -175 1202 -171
rect 1211 -175 1215 -171
rect 1224 -175 1228 -171
rect 1232 -175 1236 -171
rect 1240 -175 1244 -171
rect 1248 -175 1252 -171
rect 1256 -175 1260 -171
rect 1269 -175 1273 -171
rect 1277 -175 1281 -171
rect 1285 -175 1289 -171
rect 1293 -175 1297 -171
rect 1306 -175 1310 -171
rect 1314 -175 1318 -171
rect 1322 -175 1326 -171
rect 1330 -175 1334 -171
rect 1343 -175 1347 -171
rect 1356 -175 1360 -171
rect 1364 -175 1368 -171
rect 1372 -175 1376 -171
rect 1380 -175 1384 -171
rect 1388 -175 1392 -171
rect 1401 -175 1405 -171
rect 1409 -175 1413 -171
rect 1417 -175 1421 -171
<< pdcontact >>
rect 568 1729 572 1737
rect 581 1729 585 1737
rect 589 1729 593 1737
rect 597 1733 601 1737
rect 605 1729 609 1737
rect 618 1729 622 1737
rect 631 1729 635 1737
rect 639 1729 643 1737
rect 647 1729 651 1737
rect 655 1733 659 1737
rect 663 1729 667 1737
rect 676 1729 680 1737
rect 684 1729 688 1737
rect 692 1729 696 1737
rect 700 1729 704 1737
rect 713 1729 717 1737
rect 721 1729 725 1737
rect 729 1733 733 1737
rect 737 1729 741 1737
rect 750 1729 754 1737
rect 763 1729 767 1737
rect 771 1729 775 1737
rect 779 1729 783 1737
rect 787 1733 791 1737
rect 795 1729 799 1737
rect 808 1729 812 1737
rect 816 1729 820 1737
rect 824 1729 828 1737
rect 832 1729 836 1737
rect 845 1729 849 1737
rect 853 1729 857 1737
rect 861 1733 865 1737
rect 869 1729 873 1737
rect 882 1729 886 1737
rect 895 1729 899 1737
rect 903 1729 907 1737
rect 911 1729 915 1737
rect 919 1733 923 1737
rect 927 1729 931 1737
rect 940 1729 944 1737
rect 948 1729 952 1737
rect 956 1729 960 1737
rect 964 1729 968 1737
rect 977 1729 981 1737
rect 985 1729 989 1737
rect 993 1733 997 1737
rect 1001 1729 1005 1737
rect 1014 1729 1018 1737
rect 1027 1729 1031 1737
rect 1035 1729 1039 1737
rect 1043 1729 1047 1737
rect 1051 1733 1055 1737
rect 1059 1729 1063 1737
rect 1072 1729 1076 1737
rect 1080 1729 1084 1737
rect 1088 1729 1092 1737
rect 1501 1729 1505 1737
rect 1514 1729 1518 1737
rect 1522 1729 1526 1737
rect 1530 1733 1534 1737
rect 1538 1729 1542 1737
rect 1551 1729 1555 1737
rect 1564 1729 1568 1737
rect 1572 1729 1576 1737
rect 1580 1729 1584 1737
rect 1588 1733 1592 1737
rect 1596 1729 1600 1737
rect 1609 1729 1613 1737
rect 1617 1729 1621 1737
rect 1625 1729 1629 1737
rect 1633 1729 1637 1737
rect 1646 1729 1650 1737
rect 1654 1729 1658 1737
rect 1662 1733 1666 1737
rect 1670 1729 1674 1737
rect 1683 1729 1687 1737
rect 1696 1729 1700 1737
rect 1704 1729 1708 1737
rect 1712 1729 1716 1737
rect 1720 1733 1724 1737
rect 1728 1729 1732 1737
rect 1741 1729 1745 1737
rect 1749 1729 1753 1737
rect 1757 1729 1761 1737
rect 1765 1729 1769 1737
rect 1778 1729 1782 1737
rect 1786 1729 1790 1737
rect 1794 1733 1798 1737
rect 1802 1729 1806 1737
rect 1815 1729 1819 1737
rect 1828 1729 1832 1737
rect 1836 1729 1840 1737
rect 1844 1729 1848 1737
rect 1852 1733 1856 1737
rect 1860 1729 1864 1737
rect 1873 1729 1877 1737
rect 1881 1729 1885 1737
rect 1889 1729 1893 1737
rect 1897 1729 1901 1737
rect 1910 1729 1914 1737
rect 1918 1729 1922 1737
rect 1926 1733 1930 1737
rect 1934 1729 1938 1737
rect 1947 1729 1951 1737
rect 1960 1729 1964 1737
rect 1968 1729 1972 1737
rect 1976 1729 1980 1737
rect 1984 1733 1988 1737
rect 1992 1729 1996 1737
rect 2005 1729 2009 1737
rect 2013 1729 2017 1737
rect 2021 1729 2025 1737
rect 228 1696 232 1704
rect 241 1696 245 1704
rect 249 1696 253 1704
rect 257 1700 261 1704
rect 265 1696 269 1704
rect 278 1696 282 1704
rect 291 1696 295 1704
rect 299 1696 303 1704
rect 307 1696 311 1704
rect 315 1700 319 1704
rect 323 1696 327 1704
rect 336 1696 340 1704
rect 344 1696 348 1704
rect 352 1696 356 1704
rect 1161 1696 1165 1704
rect 1174 1696 1178 1704
rect 1182 1696 1186 1704
rect 1190 1700 1194 1704
rect 1198 1696 1202 1704
rect 1211 1696 1215 1704
rect 1224 1696 1228 1704
rect 1232 1696 1236 1704
rect 1240 1696 1244 1704
rect 1248 1700 1252 1704
rect 1256 1696 1260 1704
rect 1269 1696 1273 1704
rect 1277 1696 1281 1704
rect 1285 1696 1289 1704
rect 747 1658 751 1666
rect 755 1658 759 1666
rect 573 1645 577 1653
rect 581 1645 585 1653
rect 589 1645 593 1653
rect 597 1645 601 1653
rect 605 1645 609 1653
rect 613 1645 617 1653
rect 624 1645 628 1653
rect 641 1645 645 1653
rect 658 1645 662 1653
rect 667 1645 671 1653
rect 680 1645 684 1653
rect 688 1645 692 1653
rect 696 1645 700 1653
rect 713 1645 717 1653
rect 723 1645 727 1653
rect 731 1645 735 1653
rect 771 1652 775 1660
rect 786 1652 790 1660
rect 801 1658 805 1666
rect 809 1658 813 1666
rect 828 1658 832 1666
rect 836 1658 840 1666
rect 852 1652 856 1660
rect 867 1652 871 1660
rect 882 1658 886 1666
rect 890 1658 894 1666
rect 1680 1658 1684 1666
rect 1688 1658 1692 1666
rect 1506 1645 1510 1653
rect 1514 1645 1518 1653
rect 1522 1645 1526 1653
rect 1530 1645 1534 1653
rect 1538 1645 1542 1653
rect 1546 1645 1550 1653
rect 1557 1645 1561 1653
rect 1574 1645 1578 1653
rect 1591 1645 1595 1653
rect 1600 1645 1604 1653
rect 1613 1645 1617 1653
rect 1621 1645 1625 1653
rect 1629 1645 1633 1653
rect 1646 1645 1650 1653
rect 1656 1645 1660 1653
rect 1664 1645 1668 1653
rect 1704 1652 1708 1660
rect 1719 1652 1723 1660
rect 1734 1658 1738 1666
rect 1742 1658 1746 1666
rect 1761 1658 1765 1666
rect 1769 1658 1773 1666
rect 1785 1652 1789 1660
rect 1800 1652 1804 1660
rect 1815 1658 1819 1666
rect 1823 1658 1827 1666
rect 219 1594 223 1602
rect 227 1594 231 1602
rect 235 1594 239 1602
rect 248 1594 252 1602
rect 256 1598 260 1602
rect 264 1594 268 1602
rect 272 1594 276 1602
rect 280 1594 284 1602
rect 293 1594 297 1602
rect 306 1594 310 1602
rect 314 1598 318 1602
rect 322 1594 326 1602
rect 330 1594 334 1602
rect 343 1594 347 1602
rect 1152 1594 1156 1602
rect 1160 1594 1164 1602
rect 1168 1594 1172 1602
rect 1181 1594 1185 1602
rect 1189 1598 1193 1602
rect 1197 1594 1201 1602
rect 1205 1594 1209 1602
rect 1213 1594 1217 1602
rect 1226 1594 1230 1602
rect 1239 1594 1243 1602
rect 1247 1598 1251 1602
rect 1255 1594 1259 1602
rect 1263 1594 1267 1602
rect 1276 1594 1280 1602
rect 573 1559 577 1567
rect 581 1559 585 1567
rect 589 1559 593 1567
rect 597 1559 601 1567
rect 605 1559 609 1567
rect 613 1559 617 1567
rect 624 1559 628 1567
rect 641 1559 645 1567
rect 658 1559 662 1567
rect 667 1559 671 1567
rect 680 1559 684 1567
rect 688 1559 692 1567
rect 696 1559 700 1567
rect 713 1559 717 1567
rect 723 1559 727 1567
rect 731 1559 735 1567
rect 771 1560 775 1568
rect 786 1560 790 1568
rect 852 1560 856 1568
rect 867 1560 871 1568
rect 1506 1559 1510 1567
rect 1514 1559 1518 1567
rect 1522 1559 1526 1567
rect 1530 1559 1534 1567
rect 1538 1559 1542 1567
rect 1546 1559 1550 1567
rect 1557 1559 1561 1567
rect 1574 1559 1578 1567
rect 1591 1559 1595 1567
rect 1600 1559 1604 1567
rect 1613 1559 1617 1567
rect 1621 1559 1625 1567
rect 1629 1559 1633 1567
rect 1646 1559 1650 1567
rect 1656 1559 1660 1567
rect 1664 1559 1668 1567
rect 1704 1560 1708 1568
rect 1719 1560 1723 1568
rect 1785 1560 1789 1568
rect 1800 1560 1804 1568
rect 573 1513 577 1521
rect 581 1513 585 1521
rect 589 1513 593 1521
rect 597 1513 601 1521
rect 605 1513 609 1521
rect 613 1513 617 1521
rect 624 1513 628 1521
rect 641 1513 645 1521
rect 658 1513 662 1521
rect 667 1513 671 1521
rect 680 1513 684 1521
rect 688 1513 692 1521
rect 696 1513 700 1521
rect 713 1513 717 1521
rect 723 1513 727 1521
rect 731 1513 735 1521
rect 771 1520 775 1528
rect 786 1520 790 1528
rect 801 1526 805 1534
rect 809 1526 813 1534
rect 852 1526 856 1534
rect 860 1526 864 1534
rect 876 1520 880 1528
rect 891 1520 895 1528
rect 906 1526 910 1534
rect 914 1526 918 1534
rect 1506 1513 1510 1521
rect 1514 1513 1518 1521
rect 1522 1513 1526 1521
rect 1530 1513 1534 1521
rect 1538 1513 1542 1521
rect 1546 1513 1550 1521
rect 1557 1513 1561 1521
rect 1574 1513 1578 1521
rect 1591 1513 1595 1521
rect 1600 1513 1604 1521
rect 1613 1513 1617 1521
rect 1621 1513 1625 1521
rect 1629 1513 1633 1521
rect 1646 1513 1650 1521
rect 1656 1513 1660 1521
rect 1664 1513 1668 1521
rect 1704 1520 1708 1528
rect 1719 1520 1723 1528
rect 1734 1526 1738 1534
rect 1742 1526 1746 1534
rect 1785 1526 1789 1534
rect 1793 1526 1797 1534
rect 1809 1520 1813 1528
rect 1824 1520 1828 1528
rect 1839 1526 1843 1534
rect 1847 1526 1851 1534
rect 573 1427 577 1435
rect 581 1427 585 1435
rect 589 1427 593 1435
rect 597 1427 601 1435
rect 605 1427 609 1435
rect 613 1427 617 1435
rect 624 1427 628 1435
rect 641 1427 645 1435
rect 658 1427 662 1435
rect 667 1427 671 1435
rect 680 1427 684 1435
rect 688 1427 692 1435
rect 696 1427 700 1435
rect 713 1427 717 1435
rect 723 1427 727 1435
rect 731 1427 735 1435
rect 771 1429 775 1437
rect 786 1429 790 1437
rect 876 1429 880 1437
rect 891 1429 895 1437
rect 1506 1427 1510 1435
rect 1514 1427 1518 1435
rect 1522 1427 1526 1435
rect 1530 1427 1534 1435
rect 1538 1427 1542 1435
rect 1546 1427 1550 1435
rect 1557 1427 1561 1435
rect 1574 1427 1578 1435
rect 1591 1427 1595 1435
rect 1600 1427 1604 1435
rect 1613 1427 1617 1435
rect 1621 1427 1625 1435
rect 1629 1427 1633 1435
rect 1646 1427 1650 1435
rect 1656 1427 1660 1435
rect 1664 1427 1668 1435
rect 1704 1429 1708 1437
rect 1719 1429 1723 1437
rect 1809 1429 1813 1437
rect 1824 1429 1828 1437
rect 573 1381 577 1389
rect 581 1381 585 1389
rect 589 1381 593 1389
rect 597 1381 601 1389
rect 605 1381 609 1389
rect 613 1381 617 1389
rect 624 1381 628 1389
rect 641 1381 645 1389
rect 658 1381 662 1389
rect 667 1381 671 1389
rect 680 1381 684 1389
rect 688 1381 692 1389
rect 696 1381 700 1389
rect 713 1381 717 1389
rect 723 1381 727 1389
rect 731 1381 735 1389
rect 771 1388 775 1396
rect 786 1388 790 1396
rect 801 1394 805 1402
rect 809 1394 813 1402
rect 828 1394 832 1402
rect 836 1394 840 1402
rect 852 1388 856 1396
rect 867 1388 871 1396
rect 882 1394 886 1402
rect 890 1394 894 1402
rect 918 1394 922 1402
rect 926 1394 930 1402
rect 942 1388 946 1396
rect 957 1388 961 1396
rect 972 1394 976 1402
rect 980 1394 984 1402
rect 1506 1381 1510 1389
rect 1514 1381 1518 1389
rect 1522 1381 1526 1389
rect 1530 1381 1534 1389
rect 1538 1381 1542 1389
rect 1546 1381 1550 1389
rect 1557 1381 1561 1389
rect 1574 1381 1578 1389
rect 1591 1381 1595 1389
rect 1600 1381 1604 1389
rect 1613 1381 1617 1389
rect 1621 1381 1625 1389
rect 1629 1381 1633 1389
rect 1646 1381 1650 1389
rect 1656 1381 1660 1389
rect 1664 1381 1668 1389
rect 1704 1388 1708 1396
rect 1719 1388 1723 1396
rect 1734 1394 1738 1402
rect 1742 1394 1746 1402
rect 1761 1394 1765 1402
rect 1769 1394 1773 1402
rect 1785 1388 1789 1396
rect 1800 1388 1804 1396
rect 1815 1394 1819 1402
rect 1823 1394 1827 1402
rect 1851 1394 1855 1402
rect 1859 1394 1863 1402
rect 1875 1388 1879 1396
rect 1890 1388 1894 1396
rect 1905 1394 1909 1402
rect 1913 1394 1917 1402
rect 573 1295 577 1303
rect 581 1295 585 1303
rect 589 1295 593 1303
rect 597 1295 601 1303
rect 605 1295 609 1303
rect 613 1295 617 1303
rect 624 1295 628 1303
rect 641 1295 645 1303
rect 658 1295 662 1303
rect 667 1295 671 1303
rect 680 1295 684 1303
rect 688 1295 692 1303
rect 696 1295 700 1303
rect 713 1295 717 1303
rect 723 1295 727 1303
rect 731 1295 735 1303
rect 771 1294 775 1302
rect 786 1294 790 1302
rect 852 1294 856 1302
rect 867 1294 871 1302
rect 942 1294 946 1302
rect 957 1294 961 1302
rect 1506 1295 1510 1303
rect 1514 1295 1518 1303
rect 1522 1295 1526 1303
rect 1530 1295 1534 1303
rect 1538 1295 1542 1303
rect 1546 1295 1550 1303
rect 1557 1295 1561 1303
rect 1574 1295 1578 1303
rect 1591 1295 1595 1303
rect 1600 1295 1604 1303
rect 1613 1295 1617 1303
rect 1621 1295 1625 1303
rect 1629 1295 1633 1303
rect 1646 1295 1650 1303
rect 1656 1295 1660 1303
rect 1664 1295 1668 1303
rect 1704 1294 1708 1302
rect 1719 1294 1723 1302
rect 1785 1294 1789 1302
rect 1800 1294 1804 1302
rect 1875 1294 1879 1302
rect 1890 1294 1894 1302
rect 573 1249 577 1257
rect 581 1249 585 1257
rect 589 1249 593 1257
rect 597 1249 601 1257
rect 605 1249 609 1257
rect 613 1249 617 1257
rect 624 1249 628 1257
rect 641 1249 645 1257
rect 658 1249 662 1257
rect 667 1249 671 1257
rect 680 1249 684 1257
rect 688 1249 692 1257
rect 696 1249 700 1257
rect 713 1249 717 1257
rect 723 1249 727 1257
rect 731 1249 735 1257
rect 771 1256 775 1264
rect 786 1256 790 1264
rect 801 1262 805 1270
rect 809 1262 813 1270
rect 1506 1249 1510 1257
rect 1514 1249 1518 1257
rect 1522 1249 1526 1257
rect 1530 1249 1534 1257
rect 1538 1249 1542 1257
rect 1546 1249 1550 1257
rect 1557 1249 1561 1257
rect 1574 1249 1578 1257
rect 1591 1249 1595 1257
rect 1600 1249 1604 1257
rect 1613 1249 1617 1257
rect 1621 1249 1625 1257
rect 1629 1249 1633 1257
rect 1646 1249 1650 1257
rect 1656 1249 1660 1257
rect 1664 1249 1668 1257
rect 1704 1256 1708 1264
rect 1719 1256 1723 1264
rect 1734 1262 1738 1270
rect 1742 1262 1746 1270
rect 96 1194 100 1202
rect 109 1194 113 1202
rect 117 1194 121 1202
rect 125 1198 129 1202
rect 133 1194 137 1202
rect 146 1194 150 1202
rect 159 1194 163 1202
rect 167 1194 171 1202
rect 175 1194 179 1202
rect 183 1198 187 1202
rect 191 1194 195 1202
rect 204 1194 208 1202
rect 212 1194 216 1202
rect 220 1194 224 1202
rect 228 1194 232 1202
rect 241 1194 245 1202
rect 249 1194 253 1202
rect 257 1198 261 1202
rect 265 1194 269 1202
rect 278 1194 282 1202
rect 291 1194 295 1202
rect 299 1194 303 1202
rect 307 1194 311 1202
rect 315 1198 319 1202
rect 323 1194 327 1202
rect 336 1194 340 1202
rect 344 1194 348 1202
rect 352 1194 356 1202
rect 360 1194 364 1202
rect 373 1194 377 1202
rect 381 1194 385 1202
rect 389 1198 393 1202
rect 397 1194 401 1202
rect 410 1194 414 1202
rect 423 1194 427 1202
rect 431 1194 435 1202
rect 439 1194 443 1202
rect 447 1198 451 1202
rect 455 1194 459 1202
rect 468 1194 472 1202
rect 476 1194 480 1202
rect 484 1194 488 1202
rect 1029 1194 1033 1202
rect 1042 1194 1046 1202
rect 1050 1194 1054 1202
rect 1058 1198 1062 1202
rect 1066 1194 1070 1202
rect 1079 1194 1083 1202
rect 1092 1194 1096 1202
rect 1100 1194 1104 1202
rect 1108 1194 1112 1202
rect 1116 1198 1120 1202
rect 1124 1194 1128 1202
rect 1137 1194 1141 1202
rect 1145 1194 1149 1202
rect 1153 1194 1157 1202
rect 1161 1194 1165 1202
rect 1174 1194 1178 1202
rect 1182 1194 1186 1202
rect 1190 1198 1194 1202
rect 1198 1194 1202 1202
rect 1211 1194 1215 1202
rect 1224 1194 1228 1202
rect 1232 1194 1236 1202
rect 1240 1194 1244 1202
rect 1248 1198 1252 1202
rect 1256 1194 1260 1202
rect 1269 1194 1273 1202
rect 1277 1194 1281 1202
rect 1285 1194 1289 1202
rect 1293 1194 1297 1202
rect 1306 1194 1310 1202
rect 1314 1194 1318 1202
rect 1322 1198 1326 1202
rect 1330 1194 1334 1202
rect 1343 1194 1347 1202
rect 1356 1194 1360 1202
rect 1364 1194 1368 1202
rect 1372 1194 1376 1202
rect 1380 1198 1384 1202
rect 1388 1194 1392 1202
rect 1401 1194 1405 1202
rect 1409 1194 1413 1202
rect 1417 1194 1421 1202
rect 573 1163 577 1171
rect 581 1163 585 1171
rect 589 1163 593 1171
rect 597 1163 601 1171
rect 605 1163 609 1171
rect 613 1163 617 1171
rect 624 1163 628 1171
rect 641 1163 645 1171
rect 658 1163 662 1171
rect 667 1163 671 1171
rect 680 1163 684 1171
rect 688 1163 692 1171
rect 696 1163 700 1171
rect 713 1163 717 1171
rect 723 1163 727 1171
rect 731 1163 735 1171
rect 771 1158 775 1166
rect 786 1158 790 1166
rect 807 1163 811 1171
rect 815 1163 819 1171
rect 825 1163 829 1171
rect 833 1163 837 1171
rect 842 1163 846 1171
rect 850 1163 854 1171
rect 858 1163 862 1171
rect 866 1163 870 1171
rect 874 1163 878 1171
rect 885 1163 889 1171
rect 902 1163 906 1171
rect 919 1163 923 1171
rect 928 1163 932 1171
rect 941 1163 945 1171
rect 949 1163 953 1171
rect 957 1163 961 1171
rect 974 1163 978 1171
rect 984 1163 988 1171
rect 992 1163 996 1171
rect 1506 1163 1510 1171
rect 1514 1163 1518 1171
rect 1522 1163 1526 1171
rect 1530 1163 1534 1171
rect 1538 1163 1542 1171
rect 1546 1163 1550 1171
rect 1557 1163 1561 1171
rect 1574 1163 1578 1171
rect 1591 1163 1595 1171
rect 1600 1163 1604 1171
rect 1613 1163 1617 1171
rect 1621 1163 1625 1171
rect 1629 1163 1633 1171
rect 1646 1163 1650 1171
rect 1656 1163 1660 1171
rect 1664 1163 1668 1171
rect 1704 1158 1708 1166
rect 1719 1158 1723 1166
rect 1740 1163 1744 1171
rect 1748 1163 1752 1171
rect 1758 1163 1762 1171
rect 1766 1163 1770 1171
rect 1775 1163 1779 1171
rect 1783 1163 1787 1171
rect 1791 1163 1795 1171
rect 1799 1163 1803 1171
rect 1807 1163 1811 1171
rect 1818 1163 1822 1171
rect 1835 1163 1839 1171
rect 1852 1163 1856 1171
rect 1861 1163 1865 1171
rect 1874 1163 1878 1171
rect 1882 1163 1886 1171
rect 1890 1163 1894 1171
rect 1907 1163 1911 1171
rect 1917 1163 1921 1171
rect 1925 1163 1929 1171
rect 867 1084 871 1092
rect 880 1084 884 1092
rect 888 1084 892 1092
rect 896 1088 900 1092
rect 904 1084 908 1092
rect 917 1084 921 1092
rect 930 1084 934 1092
rect 938 1084 942 1092
rect 946 1084 950 1092
rect 954 1088 958 1092
rect 962 1084 966 1092
rect 975 1084 979 1092
rect 983 1084 987 1092
rect 991 1084 995 1092
rect 1800 1084 1804 1092
rect 1813 1084 1817 1092
rect 1821 1084 1825 1092
rect 1829 1088 1833 1092
rect 1837 1084 1841 1092
rect 1850 1084 1854 1092
rect 1863 1084 1867 1092
rect 1871 1084 1875 1092
rect 1879 1084 1883 1092
rect 1887 1088 1891 1092
rect 1895 1084 1899 1092
rect 1908 1084 1912 1092
rect 1916 1084 1920 1092
rect 1924 1084 1928 1092
rect 96 1054 100 1062
rect 109 1054 113 1062
rect 117 1054 121 1062
rect 125 1058 129 1062
rect 133 1054 137 1062
rect 146 1054 150 1062
rect 159 1054 163 1062
rect 167 1054 171 1062
rect 175 1054 179 1062
rect 183 1058 187 1062
rect 191 1054 195 1062
rect 204 1054 208 1062
rect 212 1054 216 1062
rect 220 1054 224 1062
rect 228 1054 232 1062
rect 241 1054 245 1062
rect 249 1054 253 1062
rect 257 1058 261 1062
rect 265 1054 269 1062
rect 278 1054 282 1062
rect 291 1054 295 1062
rect 299 1054 303 1062
rect 307 1054 311 1062
rect 315 1058 319 1062
rect 323 1054 327 1062
rect 336 1054 340 1062
rect 344 1054 348 1062
rect 352 1054 356 1062
rect 360 1054 364 1062
rect 373 1054 377 1062
rect 381 1054 385 1062
rect 389 1058 393 1062
rect 397 1054 401 1062
rect 410 1054 414 1062
rect 423 1054 427 1062
rect 431 1054 435 1062
rect 439 1054 443 1062
rect 447 1058 451 1062
rect 455 1054 459 1062
rect 468 1054 472 1062
rect 476 1054 480 1062
rect 484 1054 488 1062
rect 1029 1054 1033 1062
rect 1042 1054 1046 1062
rect 1050 1054 1054 1062
rect 1058 1058 1062 1062
rect 1066 1054 1070 1062
rect 1079 1054 1083 1062
rect 1092 1054 1096 1062
rect 1100 1054 1104 1062
rect 1108 1054 1112 1062
rect 1116 1058 1120 1062
rect 1124 1054 1128 1062
rect 1137 1054 1141 1062
rect 1145 1054 1149 1062
rect 1153 1054 1157 1062
rect 1161 1054 1165 1062
rect 1174 1054 1178 1062
rect 1182 1054 1186 1062
rect 1190 1058 1194 1062
rect 1198 1054 1202 1062
rect 1211 1054 1215 1062
rect 1224 1054 1228 1062
rect 1232 1054 1236 1062
rect 1240 1054 1244 1062
rect 1248 1058 1252 1062
rect 1256 1054 1260 1062
rect 1269 1054 1273 1062
rect 1277 1054 1281 1062
rect 1285 1054 1289 1062
rect 1293 1054 1297 1062
rect 1306 1054 1310 1062
rect 1314 1054 1318 1062
rect 1322 1058 1326 1062
rect 1330 1054 1334 1062
rect 1343 1054 1347 1062
rect 1356 1054 1360 1062
rect 1364 1054 1368 1062
rect 1372 1054 1376 1062
rect 1380 1058 1384 1062
rect 1388 1054 1392 1062
rect 1401 1054 1405 1062
rect 1409 1054 1413 1062
rect 1417 1054 1421 1062
rect 867 998 871 1006
rect 880 998 884 1006
rect 888 998 892 1006
rect 896 1002 900 1006
rect 904 998 908 1006
rect 917 998 921 1006
rect 930 998 934 1006
rect 938 998 942 1006
rect 946 998 950 1006
rect 954 1002 958 1006
rect 962 998 966 1006
rect 975 998 979 1006
rect 983 998 987 1006
rect 991 998 995 1006
rect 1800 998 1804 1006
rect 1813 998 1817 1006
rect 1821 998 1825 1006
rect 1829 1002 1833 1006
rect 1837 998 1841 1006
rect 1850 998 1854 1006
rect 1863 998 1867 1006
rect 1871 998 1875 1006
rect 1879 998 1883 1006
rect 1887 1002 1891 1006
rect 1895 998 1899 1006
rect 1908 998 1912 1006
rect 1916 998 1920 1006
rect 1924 998 1928 1006
rect 96 968 100 976
rect 109 968 113 976
rect 117 968 121 976
rect 125 972 129 976
rect 133 968 137 976
rect 146 968 150 976
rect 159 968 163 976
rect 167 968 171 976
rect 175 968 179 976
rect 183 972 187 976
rect 191 968 195 976
rect 204 968 208 976
rect 212 968 216 976
rect 220 968 224 976
rect 228 968 232 976
rect 241 968 245 976
rect 249 968 253 976
rect 257 972 261 976
rect 265 968 269 976
rect 278 968 282 976
rect 291 968 295 976
rect 299 968 303 976
rect 307 968 311 976
rect 315 972 319 976
rect 323 968 327 976
rect 336 968 340 976
rect 344 968 348 976
rect 352 968 356 976
rect 360 968 364 976
rect 373 968 377 976
rect 381 968 385 976
rect 389 972 393 976
rect 397 968 401 976
rect 410 968 414 976
rect 423 968 427 976
rect 431 968 435 976
rect 439 968 443 976
rect 447 972 451 976
rect 455 968 459 976
rect 468 968 472 976
rect 476 968 480 976
rect 484 968 488 976
rect 1029 968 1033 976
rect 1042 968 1046 976
rect 1050 968 1054 976
rect 1058 972 1062 976
rect 1066 968 1070 976
rect 1079 968 1083 976
rect 1092 968 1096 976
rect 1100 968 1104 976
rect 1108 968 1112 976
rect 1116 972 1120 976
rect 1124 968 1128 976
rect 1137 968 1141 976
rect 1145 968 1149 976
rect 1153 968 1157 976
rect 1161 968 1165 976
rect 1174 968 1178 976
rect 1182 968 1186 976
rect 1190 972 1194 976
rect 1198 968 1202 976
rect 1211 968 1215 976
rect 1224 968 1228 976
rect 1232 968 1236 976
rect 1240 968 1244 976
rect 1248 972 1252 976
rect 1256 968 1260 976
rect 1269 968 1273 976
rect 1277 968 1281 976
rect 1285 968 1289 976
rect 1293 968 1297 976
rect 1306 968 1310 976
rect 1314 968 1318 976
rect 1322 972 1326 976
rect 1330 968 1334 976
rect 1343 968 1347 976
rect 1356 968 1360 976
rect 1364 968 1368 976
rect 1372 968 1376 976
rect 1380 972 1384 976
rect 1388 968 1392 976
rect 1401 968 1405 976
rect 1409 968 1413 976
rect 1417 968 1421 976
rect 96 828 100 836
rect 109 828 113 836
rect 117 828 121 836
rect 125 832 129 836
rect 133 828 137 836
rect 146 828 150 836
rect 159 828 163 836
rect 167 828 171 836
rect 175 828 179 836
rect 183 832 187 836
rect 191 828 195 836
rect 204 828 208 836
rect 212 828 216 836
rect 220 828 224 836
rect 228 828 232 836
rect 241 828 245 836
rect 249 828 253 836
rect 257 832 261 836
rect 265 828 269 836
rect 278 828 282 836
rect 291 828 295 836
rect 299 828 303 836
rect 307 828 311 836
rect 315 832 319 836
rect 323 828 327 836
rect 336 828 340 836
rect 344 828 348 836
rect 352 828 356 836
rect 360 828 364 836
rect 373 828 377 836
rect 381 828 385 836
rect 389 832 393 836
rect 397 828 401 836
rect 410 828 414 836
rect 423 828 427 836
rect 431 828 435 836
rect 439 828 443 836
rect 447 832 451 836
rect 455 828 459 836
rect 468 828 472 836
rect 476 828 480 836
rect 484 828 488 836
rect 1029 828 1033 836
rect 1042 828 1046 836
rect 1050 828 1054 836
rect 1058 832 1062 836
rect 1066 828 1070 836
rect 1079 828 1083 836
rect 1092 828 1096 836
rect 1100 828 1104 836
rect 1108 828 1112 836
rect 1116 832 1120 836
rect 1124 828 1128 836
rect 1137 828 1141 836
rect 1145 828 1149 836
rect 1153 828 1157 836
rect 1161 828 1165 836
rect 1174 828 1178 836
rect 1182 828 1186 836
rect 1190 832 1194 836
rect 1198 828 1202 836
rect 1211 828 1215 836
rect 1224 828 1228 836
rect 1232 828 1236 836
rect 1240 828 1244 836
rect 1248 832 1252 836
rect 1256 828 1260 836
rect 1269 828 1273 836
rect 1277 828 1281 836
rect 1285 828 1289 836
rect 1293 828 1297 836
rect 1306 828 1310 836
rect 1314 828 1318 836
rect 1322 832 1326 836
rect 1330 828 1334 836
rect 1343 828 1347 836
rect 1356 828 1360 836
rect 1364 828 1368 836
rect 1372 828 1376 836
rect 1380 832 1384 836
rect 1388 828 1392 836
rect 1401 828 1405 836
rect 1409 828 1413 836
rect 1417 828 1421 836
rect 568 749 572 757
rect 581 749 585 757
rect 589 749 593 757
rect 597 753 601 757
rect 605 749 609 757
rect 618 749 622 757
rect 631 749 635 757
rect 639 749 643 757
rect 647 749 651 757
rect 655 753 659 757
rect 663 749 667 757
rect 676 749 680 757
rect 684 749 688 757
rect 692 749 696 757
rect 700 749 704 757
rect 713 749 717 757
rect 721 749 725 757
rect 729 753 733 757
rect 737 749 741 757
rect 750 749 754 757
rect 763 749 767 757
rect 771 749 775 757
rect 779 749 783 757
rect 787 753 791 757
rect 795 749 799 757
rect 808 749 812 757
rect 816 749 820 757
rect 824 749 828 757
rect 832 749 836 757
rect 845 749 849 757
rect 853 749 857 757
rect 861 753 865 757
rect 869 749 873 757
rect 882 749 886 757
rect 895 749 899 757
rect 903 749 907 757
rect 911 749 915 757
rect 919 753 923 757
rect 927 749 931 757
rect 940 749 944 757
rect 948 749 952 757
rect 956 749 960 757
rect 964 749 968 757
rect 977 749 981 757
rect 985 749 989 757
rect 993 753 997 757
rect 1001 749 1005 757
rect 1014 749 1018 757
rect 1027 749 1031 757
rect 1035 749 1039 757
rect 1043 749 1047 757
rect 1051 753 1055 757
rect 1059 749 1063 757
rect 1072 749 1076 757
rect 1080 749 1084 757
rect 1088 749 1092 757
rect 1501 749 1505 757
rect 1514 749 1518 757
rect 1522 749 1526 757
rect 1530 753 1534 757
rect 1538 749 1542 757
rect 1551 749 1555 757
rect 1564 749 1568 757
rect 1572 749 1576 757
rect 1580 749 1584 757
rect 1588 753 1592 757
rect 1596 749 1600 757
rect 1609 749 1613 757
rect 1617 749 1621 757
rect 1625 749 1629 757
rect 1633 749 1637 757
rect 1646 749 1650 757
rect 1654 749 1658 757
rect 1662 753 1666 757
rect 1670 749 1674 757
rect 1683 749 1687 757
rect 1696 749 1700 757
rect 1704 749 1708 757
rect 1712 749 1716 757
rect 1720 753 1724 757
rect 1728 749 1732 757
rect 1741 749 1745 757
rect 1749 749 1753 757
rect 1757 749 1761 757
rect 1765 749 1769 757
rect 1778 749 1782 757
rect 1786 749 1790 757
rect 1794 753 1798 757
rect 1802 749 1806 757
rect 1815 749 1819 757
rect 1828 749 1832 757
rect 1836 749 1840 757
rect 1844 749 1848 757
rect 1852 753 1856 757
rect 1860 749 1864 757
rect 1873 749 1877 757
rect 1881 749 1885 757
rect 1889 749 1893 757
rect 1897 749 1901 757
rect 1910 749 1914 757
rect 1918 749 1922 757
rect 1926 753 1930 757
rect 1934 749 1938 757
rect 1947 749 1951 757
rect 1960 749 1964 757
rect 1968 749 1972 757
rect 1976 749 1980 757
rect 1984 753 1988 757
rect 1992 749 1996 757
rect 2005 749 2009 757
rect 2013 749 2017 757
rect 2021 749 2025 757
rect 228 716 232 724
rect 241 716 245 724
rect 249 716 253 724
rect 257 720 261 724
rect 265 716 269 724
rect 278 716 282 724
rect 291 716 295 724
rect 299 716 303 724
rect 307 716 311 724
rect 315 720 319 724
rect 323 716 327 724
rect 336 716 340 724
rect 344 716 348 724
rect 352 716 356 724
rect 1161 716 1165 724
rect 1174 716 1178 724
rect 1182 716 1186 724
rect 1190 720 1194 724
rect 1198 716 1202 724
rect 1211 716 1215 724
rect 1224 716 1228 724
rect 1232 716 1236 724
rect 1240 716 1244 724
rect 1248 720 1252 724
rect 1256 716 1260 724
rect 1269 716 1273 724
rect 1277 716 1281 724
rect 1285 716 1289 724
rect 747 678 751 686
rect 755 678 759 686
rect 573 665 577 673
rect 581 665 585 673
rect 589 665 593 673
rect 597 665 601 673
rect 605 665 609 673
rect 613 665 617 673
rect 624 665 628 673
rect 641 665 645 673
rect 658 665 662 673
rect 667 665 671 673
rect 680 665 684 673
rect 688 665 692 673
rect 696 665 700 673
rect 713 665 717 673
rect 723 665 727 673
rect 731 665 735 673
rect 771 672 775 680
rect 786 672 790 680
rect 801 678 805 686
rect 809 678 813 686
rect 828 678 832 686
rect 836 678 840 686
rect 852 672 856 680
rect 867 672 871 680
rect 882 678 886 686
rect 890 678 894 686
rect 1680 678 1684 686
rect 1688 678 1692 686
rect 1506 665 1510 673
rect 1514 665 1518 673
rect 1522 665 1526 673
rect 1530 665 1534 673
rect 1538 665 1542 673
rect 1546 665 1550 673
rect 1557 665 1561 673
rect 1574 665 1578 673
rect 1591 665 1595 673
rect 1600 665 1604 673
rect 1613 665 1617 673
rect 1621 665 1625 673
rect 1629 665 1633 673
rect 1646 665 1650 673
rect 1656 665 1660 673
rect 1664 665 1668 673
rect 1704 672 1708 680
rect 1719 672 1723 680
rect 1734 678 1738 686
rect 1742 678 1746 686
rect 1761 678 1765 686
rect 1769 678 1773 686
rect 1785 672 1789 680
rect 1800 672 1804 680
rect 1815 678 1819 686
rect 1823 678 1827 686
rect 219 614 223 622
rect 227 614 231 622
rect 235 614 239 622
rect 248 614 252 622
rect 256 618 260 622
rect 264 614 268 622
rect 272 614 276 622
rect 280 614 284 622
rect 293 614 297 622
rect 306 614 310 622
rect 314 618 318 622
rect 322 614 326 622
rect 330 614 334 622
rect 343 614 347 622
rect 1152 614 1156 622
rect 1160 614 1164 622
rect 1168 614 1172 622
rect 1181 614 1185 622
rect 1189 618 1193 622
rect 1197 614 1201 622
rect 1205 614 1209 622
rect 1213 614 1217 622
rect 1226 614 1230 622
rect 1239 614 1243 622
rect 1247 618 1251 622
rect 1255 614 1259 622
rect 1263 614 1267 622
rect 1276 614 1280 622
rect 573 579 577 587
rect 581 579 585 587
rect 589 579 593 587
rect 597 579 601 587
rect 605 579 609 587
rect 613 579 617 587
rect 624 579 628 587
rect 641 579 645 587
rect 658 579 662 587
rect 667 579 671 587
rect 680 579 684 587
rect 688 579 692 587
rect 696 579 700 587
rect 713 579 717 587
rect 723 579 727 587
rect 731 579 735 587
rect 771 580 775 588
rect 786 580 790 588
rect 852 580 856 588
rect 867 580 871 588
rect 1506 579 1510 587
rect 1514 579 1518 587
rect 1522 579 1526 587
rect 1530 579 1534 587
rect 1538 579 1542 587
rect 1546 579 1550 587
rect 1557 579 1561 587
rect 1574 579 1578 587
rect 1591 579 1595 587
rect 1600 579 1604 587
rect 1613 579 1617 587
rect 1621 579 1625 587
rect 1629 579 1633 587
rect 1646 579 1650 587
rect 1656 579 1660 587
rect 1664 579 1668 587
rect 1704 580 1708 588
rect 1719 580 1723 588
rect 1785 580 1789 588
rect 1800 580 1804 588
rect 573 533 577 541
rect 581 533 585 541
rect 589 533 593 541
rect 597 533 601 541
rect 605 533 609 541
rect 613 533 617 541
rect 624 533 628 541
rect 641 533 645 541
rect 658 533 662 541
rect 667 533 671 541
rect 680 533 684 541
rect 688 533 692 541
rect 696 533 700 541
rect 713 533 717 541
rect 723 533 727 541
rect 731 533 735 541
rect 771 540 775 548
rect 786 540 790 548
rect 801 546 805 554
rect 809 546 813 554
rect 852 546 856 554
rect 860 546 864 554
rect 876 540 880 548
rect 891 540 895 548
rect 906 546 910 554
rect 914 546 918 554
rect 1506 533 1510 541
rect 1514 533 1518 541
rect 1522 533 1526 541
rect 1530 533 1534 541
rect 1538 533 1542 541
rect 1546 533 1550 541
rect 1557 533 1561 541
rect 1574 533 1578 541
rect 1591 533 1595 541
rect 1600 533 1604 541
rect 1613 533 1617 541
rect 1621 533 1625 541
rect 1629 533 1633 541
rect 1646 533 1650 541
rect 1656 533 1660 541
rect 1664 533 1668 541
rect 1704 540 1708 548
rect 1719 540 1723 548
rect 1734 546 1738 554
rect 1742 546 1746 554
rect 1785 546 1789 554
rect 1793 546 1797 554
rect 1809 540 1813 548
rect 1824 540 1828 548
rect 1839 546 1843 554
rect 1847 546 1851 554
rect 573 447 577 455
rect 581 447 585 455
rect 589 447 593 455
rect 597 447 601 455
rect 605 447 609 455
rect 613 447 617 455
rect 624 447 628 455
rect 641 447 645 455
rect 658 447 662 455
rect 667 447 671 455
rect 680 447 684 455
rect 688 447 692 455
rect 696 447 700 455
rect 713 447 717 455
rect 723 447 727 455
rect 731 447 735 455
rect 771 449 775 457
rect 786 449 790 457
rect 876 449 880 457
rect 891 449 895 457
rect 1506 447 1510 455
rect 1514 447 1518 455
rect 1522 447 1526 455
rect 1530 447 1534 455
rect 1538 447 1542 455
rect 1546 447 1550 455
rect 1557 447 1561 455
rect 1574 447 1578 455
rect 1591 447 1595 455
rect 1600 447 1604 455
rect 1613 447 1617 455
rect 1621 447 1625 455
rect 1629 447 1633 455
rect 1646 447 1650 455
rect 1656 447 1660 455
rect 1664 447 1668 455
rect 1704 449 1708 457
rect 1719 449 1723 457
rect 1809 449 1813 457
rect 1824 449 1828 457
rect 573 401 577 409
rect 581 401 585 409
rect 589 401 593 409
rect 597 401 601 409
rect 605 401 609 409
rect 613 401 617 409
rect 624 401 628 409
rect 641 401 645 409
rect 658 401 662 409
rect 667 401 671 409
rect 680 401 684 409
rect 688 401 692 409
rect 696 401 700 409
rect 713 401 717 409
rect 723 401 727 409
rect 731 401 735 409
rect 771 408 775 416
rect 786 408 790 416
rect 801 414 805 422
rect 809 414 813 422
rect 828 414 832 422
rect 836 414 840 422
rect 852 408 856 416
rect 867 408 871 416
rect 882 414 886 422
rect 890 414 894 422
rect 918 414 922 422
rect 926 414 930 422
rect 942 408 946 416
rect 957 408 961 416
rect 972 414 976 422
rect 980 414 984 422
rect 1506 401 1510 409
rect 1514 401 1518 409
rect 1522 401 1526 409
rect 1530 401 1534 409
rect 1538 401 1542 409
rect 1546 401 1550 409
rect 1557 401 1561 409
rect 1574 401 1578 409
rect 1591 401 1595 409
rect 1600 401 1604 409
rect 1613 401 1617 409
rect 1621 401 1625 409
rect 1629 401 1633 409
rect 1646 401 1650 409
rect 1656 401 1660 409
rect 1664 401 1668 409
rect 1704 408 1708 416
rect 1719 408 1723 416
rect 1734 414 1738 422
rect 1742 414 1746 422
rect 1761 414 1765 422
rect 1769 414 1773 422
rect 1785 408 1789 416
rect 1800 408 1804 416
rect 1815 414 1819 422
rect 1823 414 1827 422
rect 1851 414 1855 422
rect 1859 414 1863 422
rect 1875 408 1879 416
rect 1890 408 1894 416
rect 1905 414 1909 422
rect 1913 414 1917 422
rect 573 315 577 323
rect 581 315 585 323
rect 589 315 593 323
rect 597 315 601 323
rect 605 315 609 323
rect 613 315 617 323
rect 624 315 628 323
rect 641 315 645 323
rect 658 315 662 323
rect 667 315 671 323
rect 680 315 684 323
rect 688 315 692 323
rect 696 315 700 323
rect 713 315 717 323
rect 723 315 727 323
rect 731 315 735 323
rect 771 314 775 322
rect 786 314 790 322
rect 852 314 856 322
rect 867 314 871 322
rect 942 314 946 322
rect 957 314 961 322
rect 1506 315 1510 323
rect 1514 315 1518 323
rect 1522 315 1526 323
rect 1530 315 1534 323
rect 1538 315 1542 323
rect 1546 315 1550 323
rect 1557 315 1561 323
rect 1574 315 1578 323
rect 1591 315 1595 323
rect 1600 315 1604 323
rect 1613 315 1617 323
rect 1621 315 1625 323
rect 1629 315 1633 323
rect 1646 315 1650 323
rect 1656 315 1660 323
rect 1664 315 1668 323
rect 1704 314 1708 322
rect 1719 314 1723 322
rect 1785 314 1789 322
rect 1800 314 1804 322
rect 1875 314 1879 322
rect 1890 314 1894 322
rect 573 269 577 277
rect 581 269 585 277
rect 589 269 593 277
rect 597 269 601 277
rect 605 269 609 277
rect 613 269 617 277
rect 624 269 628 277
rect 641 269 645 277
rect 658 269 662 277
rect 667 269 671 277
rect 680 269 684 277
rect 688 269 692 277
rect 696 269 700 277
rect 713 269 717 277
rect 723 269 727 277
rect 731 269 735 277
rect 771 276 775 284
rect 786 276 790 284
rect 801 282 805 290
rect 809 282 813 290
rect 1506 269 1510 277
rect 1514 269 1518 277
rect 1522 269 1526 277
rect 1530 269 1534 277
rect 1538 269 1542 277
rect 1546 269 1550 277
rect 1557 269 1561 277
rect 1574 269 1578 277
rect 1591 269 1595 277
rect 1600 269 1604 277
rect 1613 269 1617 277
rect 1621 269 1625 277
rect 1629 269 1633 277
rect 1646 269 1650 277
rect 1656 269 1660 277
rect 1664 269 1668 277
rect 1704 276 1708 284
rect 1719 276 1723 284
rect 1734 282 1738 290
rect 1742 282 1746 290
rect 96 214 100 222
rect 109 214 113 222
rect 117 214 121 222
rect 125 218 129 222
rect 133 214 137 222
rect 146 214 150 222
rect 159 214 163 222
rect 167 214 171 222
rect 175 214 179 222
rect 183 218 187 222
rect 191 214 195 222
rect 204 214 208 222
rect 212 214 216 222
rect 220 214 224 222
rect 228 214 232 222
rect 241 214 245 222
rect 249 214 253 222
rect 257 218 261 222
rect 265 214 269 222
rect 278 214 282 222
rect 291 214 295 222
rect 299 214 303 222
rect 307 214 311 222
rect 315 218 319 222
rect 323 214 327 222
rect 336 214 340 222
rect 344 214 348 222
rect 352 214 356 222
rect 360 214 364 222
rect 373 214 377 222
rect 381 214 385 222
rect 389 218 393 222
rect 397 214 401 222
rect 410 214 414 222
rect 423 214 427 222
rect 431 214 435 222
rect 439 214 443 222
rect 447 218 451 222
rect 455 214 459 222
rect 468 214 472 222
rect 476 214 480 222
rect 484 214 488 222
rect 1029 214 1033 222
rect 1042 214 1046 222
rect 1050 214 1054 222
rect 1058 218 1062 222
rect 1066 214 1070 222
rect 1079 214 1083 222
rect 1092 214 1096 222
rect 1100 214 1104 222
rect 1108 214 1112 222
rect 1116 218 1120 222
rect 1124 214 1128 222
rect 1137 214 1141 222
rect 1145 214 1149 222
rect 1153 214 1157 222
rect 1161 214 1165 222
rect 1174 214 1178 222
rect 1182 214 1186 222
rect 1190 218 1194 222
rect 1198 214 1202 222
rect 1211 214 1215 222
rect 1224 214 1228 222
rect 1232 214 1236 222
rect 1240 214 1244 222
rect 1248 218 1252 222
rect 1256 214 1260 222
rect 1269 214 1273 222
rect 1277 214 1281 222
rect 1285 214 1289 222
rect 1293 214 1297 222
rect 1306 214 1310 222
rect 1314 214 1318 222
rect 1322 218 1326 222
rect 1330 214 1334 222
rect 1343 214 1347 222
rect 1356 214 1360 222
rect 1364 214 1368 222
rect 1372 214 1376 222
rect 1380 218 1384 222
rect 1388 214 1392 222
rect 1401 214 1405 222
rect 1409 214 1413 222
rect 1417 214 1421 222
rect 573 183 577 191
rect 581 183 585 191
rect 589 183 593 191
rect 597 183 601 191
rect 605 183 609 191
rect 613 183 617 191
rect 624 183 628 191
rect 641 183 645 191
rect 658 183 662 191
rect 667 183 671 191
rect 680 183 684 191
rect 688 183 692 191
rect 696 183 700 191
rect 713 183 717 191
rect 723 183 727 191
rect 731 183 735 191
rect 771 178 775 186
rect 786 178 790 186
rect 807 183 811 191
rect 815 183 819 191
rect 825 183 829 191
rect 833 183 837 191
rect 842 183 846 191
rect 850 183 854 191
rect 858 183 862 191
rect 866 183 870 191
rect 874 183 878 191
rect 885 183 889 191
rect 902 183 906 191
rect 919 183 923 191
rect 928 183 932 191
rect 941 183 945 191
rect 949 183 953 191
rect 957 183 961 191
rect 974 183 978 191
rect 984 183 988 191
rect 992 183 996 191
rect 1506 183 1510 191
rect 1514 183 1518 191
rect 1522 183 1526 191
rect 1530 183 1534 191
rect 1538 183 1542 191
rect 1546 183 1550 191
rect 1557 183 1561 191
rect 1574 183 1578 191
rect 1591 183 1595 191
rect 1600 183 1604 191
rect 1613 183 1617 191
rect 1621 183 1625 191
rect 1629 183 1633 191
rect 1646 183 1650 191
rect 1656 183 1660 191
rect 1664 183 1668 191
rect 1704 178 1708 186
rect 1719 178 1723 186
rect 1740 183 1744 191
rect 1748 183 1752 191
rect 1758 183 1762 191
rect 1766 183 1770 191
rect 1775 183 1779 191
rect 1783 183 1787 191
rect 1791 183 1795 191
rect 1799 183 1803 191
rect 1807 183 1811 191
rect 1818 183 1822 191
rect 1835 183 1839 191
rect 1852 183 1856 191
rect 1861 183 1865 191
rect 1874 183 1878 191
rect 1882 183 1886 191
rect 1890 183 1894 191
rect 1907 183 1911 191
rect 1917 183 1921 191
rect 1925 183 1929 191
rect 867 104 871 112
rect 880 104 884 112
rect 888 104 892 112
rect 896 108 900 112
rect 904 104 908 112
rect 917 104 921 112
rect 930 104 934 112
rect 938 104 942 112
rect 946 104 950 112
rect 954 108 958 112
rect 962 104 966 112
rect 975 104 979 112
rect 983 104 987 112
rect 991 104 995 112
rect 1800 104 1804 112
rect 1813 104 1817 112
rect 1821 104 1825 112
rect 1829 108 1833 112
rect 1837 104 1841 112
rect 1850 104 1854 112
rect 1863 104 1867 112
rect 1871 104 1875 112
rect 1879 104 1883 112
rect 1887 108 1891 112
rect 1895 104 1899 112
rect 1908 104 1912 112
rect 1916 104 1920 112
rect 1924 104 1928 112
rect 96 74 100 82
rect 109 74 113 82
rect 117 74 121 82
rect 125 78 129 82
rect 133 74 137 82
rect 146 74 150 82
rect 159 74 163 82
rect 167 74 171 82
rect 175 74 179 82
rect 183 78 187 82
rect 191 74 195 82
rect 204 74 208 82
rect 212 74 216 82
rect 220 74 224 82
rect 228 74 232 82
rect 241 74 245 82
rect 249 74 253 82
rect 257 78 261 82
rect 265 74 269 82
rect 278 74 282 82
rect 291 74 295 82
rect 299 74 303 82
rect 307 74 311 82
rect 315 78 319 82
rect 323 74 327 82
rect 336 74 340 82
rect 344 74 348 82
rect 352 74 356 82
rect 360 74 364 82
rect 373 74 377 82
rect 381 74 385 82
rect 389 78 393 82
rect 397 74 401 82
rect 410 74 414 82
rect 423 74 427 82
rect 431 74 435 82
rect 439 74 443 82
rect 447 78 451 82
rect 455 74 459 82
rect 468 74 472 82
rect 476 74 480 82
rect 484 74 488 82
rect 1029 74 1033 82
rect 1042 74 1046 82
rect 1050 74 1054 82
rect 1058 78 1062 82
rect 1066 74 1070 82
rect 1079 74 1083 82
rect 1092 74 1096 82
rect 1100 74 1104 82
rect 1108 74 1112 82
rect 1116 78 1120 82
rect 1124 74 1128 82
rect 1137 74 1141 82
rect 1145 74 1149 82
rect 1153 74 1157 82
rect 1161 74 1165 82
rect 1174 74 1178 82
rect 1182 74 1186 82
rect 1190 78 1194 82
rect 1198 74 1202 82
rect 1211 74 1215 82
rect 1224 74 1228 82
rect 1232 74 1236 82
rect 1240 74 1244 82
rect 1248 78 1252 82
rect 1256 74 1260 82
rect 1269 74 1273 82
rect 1277 74 1281 82
rect 1285 74 1289 82
rect 1293 74 1297 82
rect 1306 74 1310 82
rect 1314 74 1318 82
rect 1322 78 1326 82
rect 1330 74 1334 82
rect 1343 74 1347 82
rect 1356 74 1360 82
rect 1364 74 1368 82
rect 1372 74 1376 82
rect 1380 78 1384 82
rect 1388 74 1392 82
rect 1401 74 1405 82
rect 1409 74 1413 82
rect 1417 74 1421 82
rect 867 18 871 26
rect 880 18 884 26
rect 888 18 892 26
rect 896 22 900 26
rect 904 18 908 26
rect 917 18 921 26
rect 930 18 934 26
rect 938 18 942 26
rect 946 18 950 26
rect 954 22 958 26
rect 962 18 966 26
rect 975 18 979 26
rect 983 18 987 26
rect 991 18 995 26
rect 1800 18 1804 26
rect 1813 18 1817 26
rect 1821 18 1825 26
rect 1829 22 1833 26
rect 1837 18 1841 26
rect 1850 18 1854 26
rect 1863 18 1867 26
rect 1871 18 1875 26
rect 1879 18 1883 26
rect 1887 22 1891 26
rect 1895 18 1899 26
rect 1908 18 1912 26
rect 1916 18 1920 26
rect 1924 18 1928 26
rect 96 -12 100 -4
rect 109 -12 113 -4
rect 117 -12 121 -4
rect 125 -8 129 -4
rect 133 -12 137 -4
rect 146 -12 150 -4
rect 159 -12 163 -4
rect 167 -12 171 -4
rect 175 -12 179 -4
rect 183 -8 187 -4
rect 191 -12 195 -4
rect 204 -12 208 -4
rect 212 -12 216 -4
rect 220 -12 224 -4
rect 228 -12 232 -4
rect 241 -12 245 -4
rect 249 -12 253 -4
rect 257 -8 261 -4
rect 265 -12 269 -4
rect 278 -12 282 -4
rect 291 -12 295 -4
rect 299 -12 303 -4
rect 307 -12 311 -4
rect 315 -8 319 -4
rect 323 -12 327 -4
rect 336 -12 340 -4
rect 344 -12 348 -4
rect 352 -12 356 -4
rect 360 -12 364 -4
rect 373 -12 377 -4
rect 381 -12 385 -4
rect 389 -8 393 -4
rect 397 -12 401 -4
rect 410 -12 414 -4
rect 423 -12 427 -4
rect 431 -12 435 -4
rect 439 -12 443 -4
rect 447 -8 451 -4
rect 455 -12 459 -4
rect 468 -12 472 -4
rect 476 -12 480 -4
rect 484 -12 488 -4
rect 1029 -12 1033 -4
rect 1042 -12 1046 -4
rect 1050 -12 1054 -4
rect 1058 -8 1062 -4
rect 1066 -12 1070 -4
rect 1079 -12 1083 -4
rect 1092 -12 1096 -4
rect 1100 -12 1104 -4
rect 1108 -12 1112 -4
rect 1116 -8 1120 -4
rect 1124 -12 1128 -4
rect 1137 -12 1141 -4
rect 1145 -12 1149 -4
rect 1153 -12 1157 -4
rect 1161 -12 1165 -4
rect 1174 -12 1178 -4
rect 1182 -12 1186 -4
rect 1190 -8 1194 -4
rect 1198 -12 1202 -4
rect 1211 -12 1215 -4
rect 1224 -12 1228 -4
rect 1232 -12 1236 -4
rect 1240 -12 1244 -4
rect 1248 -8 1252 -4
rect 1256 -12 1260 -4
rect 1269 -12 1273 -4
rect 1277 -12 1281 -4
rect 1285 -12 1289 -4
rect 1293 -12 1297 -4
rect 1306 -12 1310 -4
rect 1314 -12 1318 -4
rect 1322 -8 1326 -4
rect 1330 -12 1334 -4
rect 1343 -12 1347 -4
rect 1356 -12 1360 -4
rect 1364 -12 1368 -4
rect 1372 -12 1376 -4
rect 1380 -8 1384 -4
rect 1388 -12 1392 -4
rect 1401 -12 1405 -4
rect 1409 -12 1413 -4
rect 1417 -12 1421 -4
rect 96 -152 100 -144
rect 109 -152 113 -144
rect 117 -152 121 -144
rect 125 -148 129 -144
rect 133 -152 137 -144
rect 146 -152 150 -144
rect 159 -152 163 -144
rect 167 -152 171 -144
rect 175 -152 179 -144
rect 183 -148 187 -144
rect 191 -152 195 -144
rect 204 -152 208 -144
rect 212 -152 216 -144
rect 220 -152 224 -144
rect 228 -152 232 -144
rect 241 -152 245 -144
rect 249 -152 253 -144
rect 257 -148 261 -144
rect 265 -152 269 -144
rect 278 -152 282 -144
rect 291 -152 295 -144
rect 299 -152 303 -144
rect 307 -152 311 -144
rect 315 -148 319 -144
rect 323 -152 327 -144
rect 336 -152 340 -144
rect 344 -152 348 -144
rect 352 -152 356 -144
rect 360 -152 364 -144
rect 373 -152 377 -144
rect 381 -152 385 -144
rect 389 -148 393 -144
rect 397 -152 401 -144
rect 410 -152 414 -144
rect 423 -152 427 -144
rect 431 -152 435 -144
rect 439 -152 443 -144
rect 447 -148 451 -144
rect 455 -152 459 -144
rect 468 -152 472 -144
rect 476 -152 480 -144
rect 484 -152 488 -144
rect 1029 -152 1033 -144
rect 1042 -152 1046 -144
rect 1050 -152 1054 -144
rect 1058 -148 1062 -144
rect 1066 -152 1070 -144
rect 1079 -152 1083 -144
rect 1092 -152 1096 -144
rect 1100 -152 1104 -144
rect 1108 -152 1112 -144
rect 1116 -148 1120 -144
rect 1124 -152 1128 -144
rect 1137 -152 1141 -144
rect 1145 -152 1149 -144
rect 1153 -152 1157 -144
rect 1161 -152 1165 -144
rect 1174 -152 1178 -144
rect 1182 -152 1186 -144
rect 1190 -148 1194 -144
rect 1198 -152 1202 -144
rect 1211 -152 1215 -144
rect 1224 -152 1228 -144
rect 1232 -152 1236 -144
rect 1240 -152 1244 -144
rect 1248 -148 1252 -144
rect 1256 -152 1260 -144
rect 1269 -152 1273 -144
rect 1277 -152 1281 -144
rect 1285 -152 1289 -144
rect 1293 -152 1297 -144
rect 1306 -152 1310 -144
rect 1314 -152 1318 -144
rect 1322 -148 1326 -144
rect 1330 -152 1334 -144
rect 1343 -152 1347 -144
rect 1356 -152 1360 -144
rect 1364 -152 1368 -144
rect 1372 -152 1376 -144
rect 1380 -148 1384 -144
rect 1388 -152 1392 -144
rect 1401 -152 1405 -144
rect 1409 -152 1413 -144
rect 1417 -152 1421 -144
<< psubstratepcontact >>
rect 598 1690 602 1694
rect 626 1690 630 1694
rect 656 1690 660 1694
rect 730 1690 734 1694
rect 758 1690 762 1694
rect 788 1690 792 1694
rect 862 1690 866 1694
rect 890 1690 894 1694
rect 920 1690 924 1694
rect 994 1690 998 1694
rect 1022 1690 1026 1694
rect 1052 1690 1056 1694
rect 1531 1690 1535 1694
rect 1559 1690 1563 1694
rect 1589 1690 1593 1694
rect 1663 1690 1667 1694
rect 1691 1690 1695 1694
rect 1721 1690 1725 1694
rect 1795 1690 1799 1694
rect 1823 1690 1827 1694
rect 1853 1690 1857 1694
rect 1927 1690 1931 1694
rect 1955 1690 1959 1694
rect 1985 1690 1989 1694
rect 258 1657 262 1661
rect 286 1657 290 1661
rect 316 1657 320 1661
rect 1191 1657 1195 1661
rect 1219 1657 1223 1661
rect 1249 1657 1253 1661
rect 579 1604 583 1608
rect 614 1604 618 1608
rect 740 1604 744 1608
rect 764 1604 768 1608
rect 818 1604 825 1608
rect 845 1604 849 1608
rect 899 1604 903 1608
rect 1512 1604 1516 1608
rect 1547 1604 1551 1608
rect 1673 1604 1677 1608
rect 1697 1604 1701 1608
rect 1751 1604 1758 1608
rect 1778 1604 1782 1608
rect 1832 1604 1836 1608
rect 255 1555 259 1559
rect 285 1555 289 1559
rect 313 1555 317 1559
rect 1188 1555 1192 1559
rect 1218 1555 1222 1559
rect 1246 1555 1250 1559
rect 579 1472 583 1476
rect 614 1472 618 1476
rect 740 1472 744 1476
rect 764 1472 768 1476
rect 818 1472 822 1476
rect 845 1472 849 1476
rect 869 1472 873 1476
rect 1512 1472 1516 1476
rect 1547 1472 1551 1476
rect 1673 1472 1677 1476
rect 1697 1472 1701 1476
rect 1751 1472 1755 1476
rect 1778 1472 1782 1476
rect 1802 1472 1806 1476
rect 579 1340 583 1344
rect 614 1340 618 1344
rect 740 1340 744 1344
rect 764 1340 768 1344
rect 818 1340 825 1344
rect 845 1340 849 1344
rect 899 1340 903 1344
rect 935 1340 939 1344
rect 989 1340 993 1344
rect 1512 1340 1516 1344
rect 1547 1340 1551 1344
rect 1673 1340 1677 1344
rect 1697 1340 1701 1344
rect 1751 1340 1758 1344
rect 1778 1340 1782 1344
rect 1832 1340 1836 1344
rect 1868 1340 1872 1344
rect 1922 1340 1926 1344
rect 579 1208 583 1212
rect 614 1208 618 1212
rect 740 1208 744 1212
rect 764 1208 768 1212
rect 875 1208 879 1212
rect 1512 1208 1516 1212
rect 1547 1208 1551 1212
rect 1673 1208 1677 1212
rect 1697 1208 1701 1212
rect 1808 1208 1812 1212
rect 126 1155 130 1159
rect 154 1155 158 1159
rect 184 1155 188 1159
rect 258 1155 262 1159
rect 286 1155 290 1159
rect 316 1155 320 1159
rect 390 1155 394 1159
rect 418 1155 422 1159
rect 448 1155 452 1159
rect 1059 1155 1063 1159
rect 1087 1155 1091 1159
rect 1117 1155 1121 1159
rect 1191 1155 1195 1159
rect 1219 1155 1223 1159
rect 1249 1155 1253 1159
rect 1323 1155 1327 1159
rect 1351 1155 1355 1159
rect 1381 1155 1385 1159
rect 897 1045 901 1049
rect 925 1045 929 1049
rect 955 1045 959 1049
rect 1830 1045 1834 1049
rect 1858 1045 1862 1049
rect 1888 1045 1892 1049
rect 126 1015 130 1019
rect 154 1015 158 1019
rect 184 1015 188 1019
rect 258 1015 262 1019
rect 286 1015 290 1019
rect 316 1015 320 1019
rect 390 1015 394 1019
rect 418 1015 422 1019
rect 448 1015 452 1019
rect 1059 1015 1063 1019
rect 1087 1015 1091 1019
rect 1117 1015 1121 1019
rect 1191 1015 1195 1019
rect 1219 1015 1223 1019
rect 1249 1015 1253 1019
rect 1323 1015 1327 1019
rect 1351 1015 1355 1019
rect 1381 1015 1385 1019
rect 897 959 901 963
rect 925 959 929 963
rect 955 959 959 963
rect 1830 959 1834 963
rect 1858 959 1862 963
rect 1888 959 1892 963
rect 126 929 130 933
rect 154 929 158 933
rect 184 929 188 933
rect 258 929 262 933
rect 286 929 290 933
rect 316 929 320 933
rect 390 929 394 933
rect 418 929 422 933
rect 448 929 452 933
rect 1059 929 1063 933
rect 1087 929 1091 933
rect 1117 929 1121 933
rect 1191 929 1195 933
rect 1219 929 1223 933
rect 1249 929 1253 933
rect 1323 929 1327 933
rect 1351 929 1355 933
rect 1381 929 1385 933
rect 126 789 130 793
rect 154 789 158 793
rect 184 789 188 793
rect 258 789 262 793
rect 286 789 290 793
rect 316 789 320 793
rect 390 789 394 793
rect 418 789 422 793
rect 448 789 452 793
rect 1059 789 1063 793
rect 1087 789 1091 793
rect 1117 789 1121 793
rect 1191 789 1195 793
rect 1219 789 1223 793
rect 1249 789 1253 793
rect 1323 789 1327 793
rect 1351 789 1355 793
rect 1381 789 1385 793
rect 598 710 602 714
rect 626 710 630 714
rect 656 710 660 714
rect 730 710 734 714
rect 758 710 762 714
rect 788 710 792 714
rect 862 710 866 714
rect 890 710 894 714
rect 920 710 924 714
rect 994 710 998 714
rect 1022 710 1026 714
rect 1052 710 1056 714
rect 1531 710 1535 714
rect 1559 710 1563 714
rect 1589 710 1593 714
rect 1663 710 1667 714
rect 1691 710 1695 714
rect 1721 710 1725 714
rect 1795 710 1799 714
rect 1823 710 1827 714
rect 1853 710 1857 714
rect 1927 710 1931 714
rect 1955 710 1959 714
rect 1985 710 1989 714
rect 258 677 262 681
rect 286 677 290 681
rect 316 677 320 681
rect 1191 677 1195 681
rect 1219 677 1223 681
rect 1249 677 1253 681
rect 579 624 583 628
rect 614 624 618 628
rect 740 624 744 628
rect 764 624 768 628
rect 818 624 825 628
rect 845 624 849 628
rect 899 624 903 628
rect 1512 624 1516 628
rect 1547 624 1551 628
rect 1673 624 1677 628
rect 1697 624 1701 628
rect 1751 624 1758 628
rect 1778 624 1782 628
rect 1832 624 1836 628
rect 255 575 259 579
rect 285 575 289 579
rect 313 575 317 579
rect 1188 575 1192 579
rect 1218 575 1222 579
rect 1246 575 1250 579
rect 579 492 583 496
rect 614 492 618 496
rect 740 492 744 496
rect 764 492 768 496
rect 818 492 822 496
rect 845 492 849 496
rect 869 492 873 496
rect 1512 492 1516 496
rect 1547 492 1551 496
rect 1673 492 1677 496
rect 1697 492 1701 496
rect 1751 492 1755 496
rect 1778 492 1782 496
rect 1802 492 1806 496
rect 579 360 583 364
rect 614 360 618 364
rect 740 360 744 364
rect 764 360 768 364
rect 818 360 825 364
rect 845 360 849 364
rect 899 360 903 364
rect 935 360 939 364
rect 989 360 993 364
rect 1512 360 1516 364
rect 1547 360 1551 364
rect 1673 360 1677 364
rect 1697 360 1701 364
rect 1751 360 1758 364
rect 1778 360 1782 364
rect 1832 360 1836 364
rect 1868 360 1872 364
rect 1922 360 1926 364
rect 579 228 583 232
rect 614 228 618 232
rect 740 228 744 232
rect 764 228 768 232
rect 875 228 879 232
rect 1512 228 1516 232
rect 1547 228 1551 232
rect 1673 228 1677 232
rect 1697 228 1701 232
rect 1808 228 1812 232
rect 126 175 130 179
rect 154 175 158 179
rect 184 175 188 179
rect 258 175 262 179
rect 286 175 290 179
rect 316 175 320 179
rect 390 175 394 179
rect 418 175 422 179
rect 448 175 452 179
rect 1059 175 1063 179
rect 1087 175 1091 179
rect 1117 175 1121 179
rect 1191 175 1195 179
rect 1219 175 1223 179
rect 1249 175 1253 179
rect 1323 175 1327 179
rect 1351 175 1355 179
rect 1381 175 1385 179
rect 897 65 901 69
rect 925 65 929 69
rect 955 65 959 69
rect 1830 65 1834 69
rect 1858 65 1862 69
rect 1888 65 1892 69
rect 126 35 130 39
rect 154 35 158 39
rect 184 35 188 39
rect 258 35 262 39
rect 286 35 290 39
rect 316 35 320 39
rect 390 35 394 39
rect 418 35 422 39
rect 448 35 452 39
rect 1059 35 1063 39
rect 1087 35 1091 39
rect 1117 35 1121 39
rect 1191 35 1195 39
rect 1219 35 1223 39
rect 1249 35 1253 39
rect 1323 35 1327 39
rect 1351 35 1355 39
rect 1381 35 1385 39
rect 897 -21 901 -17
rect 925 -21 929 -17
rect 955 -21 959 -17
rect 1830 -21 1834 -17
rect 1858 -21 1862 -17
rect 1888 -21 1892 -17
rect 126 -51 130 -47
rect 154 -51 158 -47
rect 184 -51 188 -47
rect 258 -51 262 -47
rect 286 -51 290 -47
rect 316 -51 320 -47
rect 390 -51 394 -47
rect 418 -51 422 -47
rect 448 -51 452 -47
rect 1059 -51 1063 -47
rect 1087 -51 1091 -47
rect 1117 -51 1121 -47
rect 1191 -51 1195 -47
rect 1219 -51 1223 -47
rect 1249 -51 1253 -47
rect 1323 -51 1327 -47
rect 1351 -51 1355 -47
rect 1381 -51 1385 -47
rect 126 -191 130 -187
rect 154 -191 158 -187
rect 184 -191 188 -187
rect 258 -191 262 -187
rect 286 -191 290 -187
rect 316 -191 320 -187
rect 390 -191 394 -187
rect 418 -191 422 -187
rect 448 -191 452 -187
rect 1059 -191 1063 -187
rect 1087 -191 1091 -187
rect 1117 -191 1121 -187
rect 1191 -191 1195 -187
rect 1219 -191 1223 -187
rect 1249 -191 1253 -187
rect 1323 -191 1327 -187
rect 1351 -191 1355 -187
rect 1381 -191 1385 -187
<< nsubstratencontact >>
rect 598 1747 602 1751
rect 626 1747 630 1751
rect 656 1747 660 1751
rect 693 1747 697 1751
rect 730 1747 734 1751
rect 758 1747 762 1751
rect 788 1747 792 1751
rect 825 1747 829 1751
rect 862 1747 866 1751
rect 890 1747 894 1751
rect 920 1747 924 1751
rect 957 1747 961 1751
rect 994 1747 998 1751
rect 1022 1747 1026 1751
rect 1052 1747 1056 1751
rect 1089 1747 1093 1751
rect 1531 1747 1535 1751
rect 1559 1747 1563 1751
rect 1589 1747 1593 1751
rect 1626 1747 1630 1751
rect 1663 1747 1667 1751
rect 1691 1747 1695 1751
rect 1721 1747 1725 1751
rect 1758 1747 1762 1751
rect 1795 1747 1799 1751
rect 1823 1747 1827 1751
rect 1853 1747 1857 1751
rect 1890 1747 1894 1751
rect 1927 1747 1931 1751
rect 1955 1747 1959 1751
rect 1985 1747 1989 1751
rect 2022 1747 2026 1751
rect 258 1714 262 1718
rect 286 1714 290 1718
rect 316 1714 320 1718
rect 353 1714 357 1718
rect 1191 1714 1195 1718
rect 1219 1714 1223 1718
rect 1249 1714 1253 1718
rect 1286 1714 1290 1718
rect 588 1670 592 1674
rect 617 1670 621 1674
rect 642 1670 646 1674
rect 684 1670 688 1674
rect 740 1670 744 1674
rect 764 1670 768 1674
rect 818 1670 822 1674
rect 845 1670 849 1674
rect 899 1670 903 1674
rect 1521 1670 1525 1674
rect 1550 1670 1554 1674
rect 1575 1670 1579 1674
rect 1617 1670 1621 1674
rect 1673 1670 1677 1674
rect 1697 1670 1701 1674
rect 1751 1670 1755 1674
rect 1778 1670 1782 1674
rect 1832 1670 1836 1674
rect 218 1612 222 1616
rect 255 1612 259 1616
rect 285 1612 289 1616
rect 313 1612 317 1616
rect 1151 1612 1155 1616
rect 1188 1612 1192 1616
rect 1218 1612 1222 1616
rect 1246 1612 1250 1616
rect 588 1538 592 1542
rect 617 1538 621 1542
rect 642 1538 646 1542
rect 684 1538 688 1542
rect 740 1538 744 1542
rect 764 1538 768 1542
rect 818 1538 822 1542
rect 845 1538 849 1542
rect 907 1538 911 1542
rect 1521 1538 1525 1542
rect 1550 1538 1554 1542
rect 1575 1538 1579 1542
rect 1617 1538 1621 1542
rect 1673 1538 1677 1542
rect 1697 1538 1701 1542
rect 1751 1538 1755 1542
rect 1778 1538 1782 1542
rect 1840 1538 1844 1542
rect 588 1406 592 1410
rect 617 1406 621 1410
rect 642 1406 646 1410
rect 684 1406 688 1410
rect 740 1406 744 1410
rect 764 1406 768 1410
rect 818 1406 822 1410
rect 845 1406 849 1410
rect 899 1406 903 1410
rect 907 1406 911 1410
rect 935 1406 939 1410
rect 989 1406 993 1410
rect 1521 1406 1525 1410
rect 1550 1406 1554 1410
rect 1575 1406 1579 1410
rect 1617 1406 1621 1410
rect 1673 1406 1677 1410
rect 1697 1406 1701 1410
rect 1751 1406 1755 1410
rect 1778 1406 1782 1410
rect 1832 1406 1836 1410
rect 1840 1406 1844 1410
rect 1868 1406 1872 1410
rect 1922 1406 1926 1410
rect 588 1274 592 1278
rect 617 1274 621 1278
rect 642 1274 646 1278
rect 684 1274 688 1278
rect 740 1274 744 1278
rect 764 1274 768 1278
rect 818 1274 822 1278
rect 845 1274 849 1278
rect 935 1274 939 1278
rect 1521 1274 1525 1278
rect 1550 1274 1554 1278
rect 1575 1274 1579 1278
rect 1617 1274 1621 1278
rect 1673 1274 1677 1278
rect 1697 1274 1701 1278
rect 1751 1274 1755 1278
rect 1778 1274 1782 1278
rect 1868 1274 1872 1278
rect 126 1212 130 1216
rect 154 1212 158 1216
rect 184 1212 188 1216
rect 221 1212 225 1216
rect 258 1212 262 1216
rect 286 1212 290 1216
rect 316 1212 320 1216
rect 353 1212 357 1216
rect 390 1212 394 1216
rect 418 1212 422 1216
rect 448 1212 452 1216
rect 485 1212 489 1216
rect 1059 1212 1063 1216
rect 1087 1212 1091 1216
rect 1117 1212 1121 1216
rect 1154 1212 1158 1216
rect 1191 1212 1195 1216
rect 1219 1212 1223 1216
rect 1249 1212 1253 1216
rect 1286 1212 1290 1216
rect 1323 1212 1327 1216
rect 1351 1212 1355 1216
rect 1381 1212 1385 1216
rect 1418 1212 1422 1216
rect 588 1142 592 1146
rect 617 1142 621 1146
rect 642 1142 646 1146
rect 684 1142 688 1146
rect 764 1142 768 1146
rect 818 1142 822 1146
rect 849 1142 853 1146
rect 878 1142 882 1146
rect 903 1142 907 1146
rect 945 1142 949 1146
rect 1521 1142 1525 1146
rect 1550 1142 1554 1146
rect 1575 1142 1579 1146
rect 1617 1142 1621 1146
rect 1697 1142 1701 1146
rect 1751 1142 1755 1146
rect 1782 1142 1786 1146
rect 1811 1142 1815 1146
rect 1836 1142 1840 1146
rect 1878 1142 1882 1146
rect 897 1102 901 1106
rect 925 1102 929 1106
rect 955 1102 959 1106
rect 992 1102 996 1106
rect 1830 1102 1834 1106
rect 1858 1102 1862 1106
rect 1888 1102 1892 1106
rect 1925 1102 1929 1106
rect 126 1072 130 1076
rect 154 1072 158 1076
rect 184 1072 188 1076
rect 221 1072 225 1076
rect 258 1072 262 1076
rect 286 1072 290 1076
rect 316 1072 320 1076
rect 353 1072 357 1076
rect 390 1072 394 1076
rect 418 1072 422 1076
rect 448 1072 452 1076
rect 485 1072 489 1076
rect 1059 1072 1063 1076
rect 1087 1072 1091 1076
rect 1117 1072 1121 1076
rect 1154 1072 1158 1076
rect 1191 1072 1195 1076
rect 1219 1072 1223 1076
rect 1249 1072 1253 1076
rect 1286 1072 1290 1076
rect 1323 1072 1327 1076
rect 1351 1072 1355 1076
rect 1381 1072 1385 1076
rect 1418 1072 1422 1076
rect 897 1016 901 1020
rect 925 1016 929 1020
rect 955 1016 959 1020
rect 992 1016 996 1020
rect 1830 1016 1834 1020
rect 1858 1016 1862 1020
rect 1888 1016 1892 1020
rect 1925 1016 1929 1020
rect 126 986 130 990
rect 154 986 158 990
rect 184 986 188 990
rect 221 986 225 990
rect 258 986 262 990
rect 286 986 290 990
rect 316 986 320 990
rect 353 986 357 990
rect 390 986 394 990
rect 418 986 422 990
rect 448 986 452 990
rect 485 986 489 990
rect 1059 986 1063 990
rect 1087 986 1091 990
rect 1117 986 1121 990
rect 1154 986 1158 990
rect 1191 986 1195 990
rect 1219 986 1223 990
rect 1249 986 1253 990
rect 1286 986 1290 990
rect 1323 986 1327 990
rect 1351 986 1355 990
rect 1381 986 1385 990
rect 1418 986 1422 990
rect 126 846 130 850
rect 154 846 158 850
rect 184 846 188 850
rect 221 846 225 850
rect 258 846 262 850
rect 286 846 290 850
rect 316 846 320 850
rect 353 846 357 850
rect 390 846 394 850
rect 418 846 422 850
rect 448 846 452 850
rect 485 846 489 850
rect 1059 846 1063 850
rect 1087 846 1091 850
rect 1117 846 1121 850
rect 1154 846 1158 850
rect 1191 846 1195 850
rect 1219 846 1223 850
rect 1249 846 1253 850
rect 1286 846 1290 850
rect 1323 846 1327 850
rect 1351 846 1355 850
rect 1381 846 1385 850
rect 1418 846 1422 850
rect 598 767 602 771
rect 626 767 630 771
rect 656 767 660 771
rect 693 767 697 771
rect 730 767 734 771
rect 758 767 762 771
rect 788 767 792 771
rect 825 767 829 771
rect 862 767 866 771
rect 890 767 894 771
rect 920 767 924 771
rect 957 767 961 771
rect 994 767 998 771
rect 1022 767 1026 771
rect 1052 767 1056 771
rect 1089 767 1093 771
rect 1531 767 1535 771
rect 1559 767 1563 771
rect 1589 767 1593 771
rect 1626 767 1630 771
rect 1663 767 1667 771
rect 1691 767 1695 771
rect 1721 767 1725 771
rect 1758 767 1762 771
rect 1795 767 1799 771
rect 1823 767 1827 771
rect 1853 767 1857 771
rect 1890 767 1894 771
rect 1927 767 1931 771
rect 1955 767 1959 771
rect 1985 767 1989 771
rect 2022 767 2026 771
rect 258 734 262 738
rect 286 734 290 738
rect 316 734 320 738
rect 353 734 357 738
rect 1191 734 1195 738
rect 1219 734 1223 738
rect 1249 734 1253 738
rect 1286 734 1290 738
rect 588 690 592 694
rect 617 690 621 694
rect 642 690 646 694
rect 684 690 688 694
rect 740 690 744 694
rect 764 690 768 694
rect 818 690 822 694
rect 845 690 849 694
rect 899 690 903 694
rect 1521 690 1525 694
rect 1550 690 1554 694
rect 1575 690 1579 694
rect 1617 690 1621 694
rect 1673 690 1677 694
rect 1697 690 1701 694
rect 1751 690 1755 694
rect 1778 690 1782 694
rect 1832 690 1836 694
rect 218 632 222 636
rect 255 632 259 636
rect 285 632 289 636
rect 313 632 317 636
rect 1151 632 1155 636
rect 1188 632 1192 636
rect 1218 632 1222 636
rect 1246 632 1250 636
rect 588 558 592 562
rect 617 558 621 562
rect 642 558 646 562
rect 684 558 688 562
rect 740 558 744 562
rect 764 558 768 562
rect 818 558 822 562
rect 845 558 849 562
rect 907 558 911 562
rect 1521 558 1525 562
rect 1550 558 1554 562
rect 1575 558 1579 562
rect 1617 558 1621 562
rect 1673 558 1677 562
rect 1697 558 1701 562
rect 1751 558 1755 562
rect 1778 558 1782 562
rect 1840 558 1844 562
rect 588 426 592 430
rect 617 426 621 430
rect 642 426 646 430
rect 684 426 688 430
rect 740 426 744 430
rect 764 426 768 430
rect 818 426 822 430
rect 845 426 849 430
rect 899 426 903 430
rect 907 426 911 430
rect 935 426 939 430
rect 989 426 993 430
rect 1521 426 1525 430
rect 1550 426 1554 430
rect 1575 426 1579 430
rect 1617 426 1621 430
rect 1673 426 1677 430
rect 1697 426 1701 430
rect 1751 426 1755 430
rect 1778 426 1782 430
rect 1832 426 1836 430
rect 1840 426 1844 430
rect 1868 426 1872 430
rect 1922 426 1926 430
rect 588 294 592 298
rect 617 294 621 298
rect 642 294 646 298
rect 684 294 688 298
rect 740 294 744 298
rect 764 294 768 298
rect 818 294 822 298
rect 845 294 849 298
rect 935 294 939 298
rect 1521 294 1525 298
rect 1550 294 1554 298
rect 1575 294 1579 298
rect 1617 294 1621 298
rect 1673 294 1677 298
rect 1697 294 1701 298
rect 1751 294 1755 298
rect 1778 294 1782 298
rect 1868 294 1872 298
rect 126 232 130 236
rect 154 232 158 236
rect 184 232 188 236
rect 221 232 225 236
rect 258 232 262 236
rect 286 232 290 236
rect 316 232 320 236
rect 353 232 357 236
rect 390 232 394 236
rect 418 232 422 236
rect 448 232 452 236
rect 485 232 489 236
rect 1059 232 1063 236
rect 1087 232 1091 236
rect 1117 232 1121 236
rect 1154 232 1158 236
rect 1191 232 1195 236
rect 1219 232 1223 236
rect 1249 232 1253 236
rect 1286 232 1290 236
rect 1323 232 1327 236
rect 1351 232 1355 236
rect 1381 232 1385 236
rect 1418 232 1422 236
rect 588 162 592 166
rect 617 162 621 166
rect 642 162 646 166
rect 684 162 688 166
rect 764 162 768 166
rect 818 162 822 166
rect 849 162 853 166
rect 878 162 882 166
rect 903 162 907 166
rect 945 162 949 166
rect 1521 162 1525 166
rect 1550 162 1554 166
rect 1575 162 1579 166
rect 1617 162 1621 166
rect 1697 162 1701 166
rect 1751 162 1755 166
rect 1782 162 1786 166
rect 1811 162 1815 166
rect 1836 162 1840 166
rect 1878 162 1882 166
rect 897 122 901 126
rect 925 122 929 126
rect 955 122 959 126
rect 992 122 996 126
rect 1830 122 1834 126
rect 1858 122 1862 126
rect 1888 122 1892 126
rect 1925 122 1929 126
rect 126 92 130 96
rect 154 92 158 96
rect 184 92 188 96
rect 221 92 225 96
rect 258 92 262 96
rect 286 92 290 96
rect 316 92 320 96
rect 353 92 357 96
rect 390 92 394 96
rect 418 92 422 96
rect 448 92 452 96
rect 485 92 489 96
rect 1059 92 1063 96
rect 1087 92 1091 96
rect 1117 92 1121 96
rect 1154 92 1158 96
rect 1191 92 1195 96
rect 1219 92 1223 96
rect 1249 92 1253 96
rect 1286 92 1290 96
rect 1323 92 1327 96
rect 1351 92 1355 96
rect 1381 92 1385 96
rect 1418 92 1422 96
rect 897 36 901 40
rect 925 36 929 40
rect 955 36 959 40
rect 992 36 996 40
rect 1830 36 1834 40
rect 1858 36 1862 40
rect 1888 36 1892 40
rect 1925 36 1929 40
rect 126 6 130 10
rect 154 6 158 10
rect 184 6 188 10
rect 221 6 225 10
rect 258 6 262 10
rect 286 6 290 10
rect 316 6 320 10
rect 353 6 357 10
rect 390 6 394 10
rect 418 6 422 10
rect 448 6 452 10
rect 485 6 489 10
rect 1059 6 1063 10
rect 1087 6 1091 10
rect 1117 6 1121 10
rect 1154 6 1158 10
rect 1191 6 1195 10
rect 1219 6 1223 10
rect 1249 6 1253 10
rect 1286 6 1290 10
rect 1323 6 1327 10
rect 1351 6 1355 10
rect 1381 6 1385 10
rect 1418 6 1422 10
rect 126 -134 130 -130
rect 154 -134 158 -130
rect 184 -134 188 -130
rect 221 -134 225 -130
rect 258 -134 262 -130
rect 286 -134 290 -130
rect 316 -134 320 -130
rect 353 -134 357 -130
rect 390 -134 394 -130
rect 418 -134 422 -130
rect 448 -134 452 -130
rect 485 -134 489 -130
rect 1059 -134 1063 -130
rect 1087 -134 1091 -130
rect 1117 -134 1121 -130
rect 1154 -134 1158 -130
rect 1191 -134 1195 -130
rect 1219 -134 1223 -130
rect 1249 -134 1253 -130
rect 1286 -134 1290 -130
rect 1323 -134 1327 -130
rect 1351 -134 1355 -130
rect 1381 -134 1385 -130
rect 1418 -134 1422 -130
<< polysilicon >>
rect 573 1737 575 1739
rect 578 1737 580 1740
rect 594 1737 596 1739
rect 610 1737 612 1739
rect 615 1737 617 1740
rect 636 1737 638 1740
rect 652 1737 654 1740
rect 668 1737 670 1739
rect 673 1737 675 1740
rect 689 1737 691 1739
rect 705 1737 707 1739
rect 710 1737 712 1740
rect 726 1737 728 1739
rect 742 1737 744 1739
rect 747 1737 749 1740
rect 768 1737 770 1740
rect 784 1737 786 1740
rect 800 1737 802 1739
rect 805 1737 807 1740
rect 821 1737 823 1739
rect 837 1737 839 1739
rect 842 1737 844 1740
rect 858 1737 860 1739
rect 874 1737 876 1739
rect 879 1737 881 1740
rect 900 1737 902 1740
rect 916 1737 918 1740
rect 932 1737 934 1739
rect 937 1737 939 1740
rect 953 1737 955 1739
rect 969 1737 971 1739
rect 974 1737 976 1740
rect 990 1737 992 1739
rect 1006 1737 1008 1739
rect 1011 1737 1013 1740
rect 1032 1737 1034 1740
rect 1048 1737 1050 1740
rect 1064 1737 1066 1739
rect 1069 1737 1071 1740
rect 1085 1737 1087 1739
rect 1506 1737 1508 1739
rect 1511 1737 1513 1740
rect 1527 1737 1529 1739
rect 1543 1737 1545 1739
rect 1548 1737 1550 1740
rect 1569 1737 1571 1740
rect 1585 1737 1587 1740
rect 1601 1737 1603 1739
rect 1606 1737 1608 1740
rect 1622 1737 1624 1739
rect 1638 1737 1640 1739
rect 1643 1737 1645 1740
rect 1659 1737 1661 1739
rect 1675 1737 1677 1739
rect 1680 1737 1682 1740
rect 1701 1737 1703 1740
rect 1717 1737 1719 1740
rect 1733 1737 1735 1739
rect 1738 1737 1740 1740
rect 1754 1737 1756 1739
rect 1770 1737 1772 1739
rect 1775 1737 1777 1740
rect 1791 1737 1793 1739
rect 1807 1737 1809 1739
rect 1812 1737 1814 1740
rect 1833 1737 1835 1740
rect 1849 1737 1851 1740
rect 1865 1737 1867 1739
rect 1870 1737 1872 1740
rect 1886 1737 1888 1739
rect 1902 1737 1904 1739
rect 1907 1737 1909 1740
rect 1923 1737 1925 1739
rect 1939 1737 1941 1739
rect 1944 1737 1946 1740
rect 1965 1737 1967 1740
rect 1981 1737 1983 1740
rect 1997 1737 1999 1739
rect 2002 1737 2004 1740
rect 2018 1737 2020 1739
rect 573 1724 575 1729
rect 578 1727 580 1729
rect 573 1710 575 1720
rect 578 1710 580 1717
rect 594 1710 596 1729
rect 610 1720 612 1729
rect 615 1727 617 1729
rect 636 1727 638 1729
rect 652 1726 654 1729
rect 610 1710 612 1713
rect 615 1710 617 1712
rect 636 1710 638 1712
rect 652 1710 654 1722
rect 668 1720 670 1729
rect 673 1727 675 1729
rect 689 1721 691 1729
rect 705 1724 707 1729
rect 710 1727 712 1729
rect 668 1710 670 1713
rect 673 1710 675 1712
rect 689 1710 691 1717
rect 705 1710 707 1720
rect 710 1710 712 1717
rect 726 1710 728 1729
rect 742 1720 744 1729
rect 747 1727 749 1729
rect 768 1727 770 1729
rect 784 1726 786 1729
rect 742 1710 744 1713
rect 747 1710 749 1712
rect 768 1710 770 1712
rect 784 1710 786 1722
rect 800 1720 802 1729
rect 805 1727 807 1729
rect 821 1721 823 1729
rect 837 1724 839 1729
rect 842 1727 844 1729
rect 800 1710 802 1713
rect 805 1710 807 1712
rect 821 1710 823 1717
rect 837 1710 839 1720
rect 842 1710 844 1717
rect 858 1710 860 1729
rect 874 1720 876 1729
rect 879 1727 881 1729
rect 900 1727 902 1729
rect 916 1726 918 1729
rect 874 1710 876 1713
rect 879 1710 881 1712
rect 900 1710 902 1712
rect 916 1710 918 1722
rect 932 1720 934 1729
rect 937 1727 939 1729
rect 953 1721 955 1729
rect 969 1724 971 1729
rect 974 1727 976 1729
rect 932 1710 934 1713
rect 937 1710 939 1712
rect 953 1710 955 1717
rect 969 1710 971 1720
rect 974 1710 976 1717
rect 990 1710 992 1729
rect 1006 1720 1008 1729
rect 1011 1727 1013 1729
rect 1032 1727 1034 1729
rect 1048 1726 1050 1729
rect 1006 1710 1008 1713
rect 1011 1710 1013 1712
rect 1032 1710 1034 1712
rect 1048 1710 1050 1722
rect 1064 1720 1066 1729
rect 1069 1727 1071 1729
rect 1085 1721 1087 1729
rect 1506 1724 1508 1729
rect 1511 1727 1513 1729
rect 1064 1710 1066 1713
rect 1069 1710 1071 1712
rect 1085 1710 1087 1717
rect 233 1704 235 1706
rect 238 1704 240 1707
rect 254 1704 256 1706
rect 270 1704 272 1706
rect 275 1704 277 1707
rect 296 1704 298 1707
rect 312 1704 314 1707
rect 328 1704 330 1706
rect 333 1704 335 1707
rect 1506 1710 1508 1720
rect 1511 1710 1513 1717
rect 1527 1710 1529 1729
rect 1543 1720 1545 1729
rect 1548 1727 1550 1729
rect 1569 1727 1571 1729
rect 1585 1726 1587 1729
rect 1543 1710 1545 1713
rect 1548 1710 1550 1712
rect 1569 1710 1571 1712
rect 1585 1710 1587 1722
rect 1601 1720 1603 1729
rect 1606 1727 1608 1729
rect 1622 1721 1624 1729
rect 1638 1724 1640 1729
rect 1643 1727 1645 1729
rect 1601 1710 1603 1713
rect 1606 1710 1608 1712
rect 1622 1710 1624 1717
rect 1638 1710 1640 1720
rect 1643 1710 1645 1717
rect 1659 1710 1661 1729
rect 1675 1720 1677 1729
rect 1680 1727 1682 1729
rect 1701 1727 1703 1729
rect 1717 1726 1719 1729
rect 1675 1710 1677 1713
rect 1680 1710 1682 1712
rect 1701 1710 1703 1712
rect 1717 1710 1719 1722
rect 1733 1720 1735 1729
rect 1738 1727 1740 1729
rect 1754 1721 1756 1729
rect 1770 1724 1772 1729
rect 1775 1727 1777 1729
rect 1733 1710 1735 1713
rect 1738 1710 1740 1712
rect 1754 1710 1756 1717
rect 1770 1710 1772 1720
rect 1775 1710 1777 1717
rect 1791 1710 1793 1729
rect 1807 1720 1809 1729
rect 1812 1727 1814 1729
rect 1833 1727 1835 1729
rect 1849 1726 1851 1729
rect 1807 1710 1809 1713
rect 1812 1710 1814 1712
rect 1833 1710 1835 1712
rect 1849 1710 1851 1722
rect 1865 1720 1867 1729
rect 1870 1727 1872 1729
rect 1886 1721 1888 1729
rect 1902 1724 1904 1729
rect 1907 1727 1909 1729
rect 1865 1710 1867 1713
rect 1870 1710 1872 1712
rect 1886 1710 1888 1717
rect 1902 1710 1904 1720
rect 1907 1710 1909 1717
rect 1923 1710 1925 1729
rect 1939 1720 1941 1729
rect 1944 1727 1946 1729
rect 1965 1727 1967 1729
rect 1981 1726 1983 1729
rect 1939 1710 1941 1713
rect 1944 1710 1946 1712
rect 1965 1710 1967 1712
rect 1981 1710 1983 1722
rect 1997 1720 1999 1729
rect 2002 1727 2004 1729
rect 2018 1721 2020 1729
rect 1997 1710 1999 1713
rect 2002 1710 2004 1712
rect 2018 1710 2020 1717
rect 349 1704 351 1706
rect 573 1704 575 1706
rect 578 1703 580 1706
rect 594 1704 596 1706
rect 610 1704 612 1706
rect 615 1701 617 1706
rect 636 1701 638 1706
rect 652 1704 654 1706
rect 668 1704 670 1706
rect 673 1701 675 1706
rect 689 1704 691 1706
rect 705 1704 707 1706
rect 710 1703 712 1706
rect 726 1704 728 1706
rect 742 1704 744 1706
rect 747 1701 749 1706
rect 768 1701 770 1706
rect 784 1704 786 1706
rect 800 1704 802 1706
rect 805 1701 807 1706
rect 821 1704 823 1706
rect 837 1704 839 1706
rect 842 1703 844 1706
rect 858 1704 860 1706
rect 874 1704 876 1706
rect 879 1701 881 1706
rect 900 1701 902 1706
rect 916 1704 918 1706
rect 932 1704 934 1706
rect 937 1701 939 1706
rect 953 1704 955 1706
rect 969 1704 971 1706
rect 974 1703 976 1706
rect 990 1704 992 1706
rect 1006 1704 1008 1706
rect 1011 1701 1013 1706
rect 1032 1701 1034 1706
rect 1048 1704 1050 1706
rect 1064 1704 1066 1706
rect 1069 1701 1071 1706
rect 1085 1704 1087 1706
rect 1166 1704 1168 1706
rect 1171 1704 1173 1707
rect 1187 1704 1189 1706
rect 1203 1704 1205 1706
rect 1208 1704 1210 1707
rect 1229 1704 1231 1707
rect 1245 1704 1247 1707
rect 1261 1704 1263 1706
rect 1266 1704 1268 1707
rect 1282 1704 1284 1706
rect 1506 1704 1508 1706
rect 1511 1703 1513 1706
rect 1527 1704 1529 1706
rect 1543 1704 1545 1706
rect 1548 1701 1550 1706
rect 1569 1701 1571 1706
rect 1585 1704 1587 1706
rect 1601 1704 1603 1706
rect 1606 1701 1608 1706
rect 1622 1704 1624 1706
rect 1638 1704 1640 1706
rect 1643 1703 1645 1706
rect 1659 1704 1661 1706
rect 1675 1704 1677 1706
rect 1680 1701 1682 1706
rect 1701 1701 1703 1706
rect 1717 1704 1719 1706
rect 1733 1704 1735 1706
rect 1738 1701 1740 1706
rect 1754 1704 1756 1706
rect 1770 1704 1772 1706
rect 1775 1703 1777 1706
rect 1791 1704 1793 1706
rect 1807 1704 1809 1706
rect 1812 1701 1814 1706
rect 1833 1701 1835 1706
rect 1849 1704 1851 1706
rect 1865 1704 1867 1706
rect 1870 1701 1872 1706
rect 1886 1704 1888 1706
rect 1902 1704 1904 1706
rect 1907 1703 1909 1706
rect 1923 1704 1925 1706
rect 1939 1704 1941 1706
rect 1944 1701 1946 1706
rect 1965 1701 1967 1706
rect 1981 1704 1983 1706
rect 1997 1704 1999 1706
rect 2002 1701 2004 1706
rect 2018 1704 2020 1706
rect 233 1691 235 1696
rect 238 1694 240 1696
rect 233 1677 235 1687
rect 238 1677 240 1684
rect 254 1677 256 1696
rect 270 1687 272 1696
rect 275 1694 277 1696
rect 296 1694 298 1696
rect 312 1693 314 1696
rect 270 1677 272 1680
rect 275 1677 277 1679
rect 296 1677 298 1679
rect 312 1677 314 1689
rect 328 1687 330 1696
rect 333 1694 335 1696
rect 328 1677 330 1680
rect 333 1677 335 1679
rect 349 1677 351 1696
rect 1166 1691 1168 1696
rect 1171 1694 1173 1696
rect 1166 1677 1168 1687
rect 1171 1677 1173 1684
rect 1187 1677 1189 1696
rect 1203 1687 1205 1696
rect 1208 1694 1210 1696
rect 1229 1694 1231 1696
rect 1245 1693 1247 1696
rect 1203 1677 1205 1680
rect 1208 1677 1210 1679
rect 1229 1677 1231 1679
rect 1245 1677 1247 1689
rect 1261 1687 1263 1696
rect 1266 1694 1268 1696
rect 1261 1677 1263 1680
rect 1266 1677 1268 1679
rect 1282 1677 1284 1696
rect 233 1671 235 1673
rect 238 1670 240 1673
rect 254 1671 256 1673
rect 270 1671 272 1673
rect 275 1668 277 1673
rect 296 1668 298 1673
rect 312 1671 314 1673
rect 328 1671 330 1673
rect 333 1668 335 1673
rect 349 1671 351 1673
rect 1166 1671 1168 1673
rect 1171 1670 1173 1673
rect 1187 1671 1189 1673
rect 1203 1671 1205 1673
rect 752 1666 754 1668
rect 594 1660 596 1663
rect 638 1660 640 1663
rect 664 1660 666 1663
rect 710 1660 712 1663
rect 664 1656 665 1660
rect 778 1660 780 1664
rect 806 1666 808 1668
rect 833 1666 835 1668
rect 783 1660 785 1663
rect 578 1653 580 1655
rect 594 1653 596 1656
rect 610 1653 612 1655
rect 633 1653 635 1655
rect 638 1653 640 1656
rect 664 1653 666 1656
rect 685 1653 687 1656
rect 705 1653 707 1655
rect 710 1653 712 1656
rect 728 1653 730 1655
rect 357 1640 359 1643
rect 357 1634 359 1636
rect 240 1631 242 1634
rect 578 1631 580 1645
rect 594 1643 596 1645
rect 594 1631 596 1633
rect 610 1631 612 1645
rect 633 1640 635 1645
rect 638 1643 640 1645
rect 664 1643 666 1645
rect 629 1636 635 1640
rect 633 1631 635 1636
rect 638 1631 640 1633
rect 664 1631 666 1633
rect 685 1631 687 1645
rect 705 1640 707 1645
rect 710 1643 712 1645
rect 701 1636 707 1640
rect 705 1631 707 1636
rect 710 1631 712 1633
rect 728 1631 730 1645
rect 752 1644 754 1658
rect 859 1660 861 1664
rect 887 1666 889 1668
rect 1208 1668 1210 1673
rect 1229 1668 1231 1673
rect 1245 1671 1247 1673
rect 1261 1671 1263 1673
rect 1266 1668 1268 1673
rect 1282 1671 1284 1673
rect 864 1660 866 1663
rect 778 1649 780 1652
rect 783 1650 785 1652
rect 779 1645 780 1649
rect 778 1640 780 1645
rect 783 1640 785 1642
rect 752 1638 754 1640
rect 806 1636 808 1658
rect 833 1644 835 1658
rect 1685 1666 1687 1668
rect 859 1649 861 1652
rect 864 1650 866 1652
rect 860 1645 861 1649
rect 859 1640 861 1645
rect 864 1640 866 1642
rect 833 1638 835 1640
rect 887 1636 889 1658
rect 1527 1660 1529 1663
rect 1571 1660 1573 1663
rect 1597 1660 1599 1663
rect 1643 1660 1645 1663
rect 1597 1656 1598 1660
rect 1711 1660 1713 1664
rect 1739 1666 1741 1668
rect 1766 1666 1768 1668
rect 1716 1660 1718 1663
rect 1511 1653 1513 1655
rect 1527 1653 1529 1656
rect 1543 1653 1545 1655
rect 1566 1653 1568 1655
rect 1571 1653 1573 1656
rect 1597 1653 1599 1656
rect 1618 1653 1620 1656
rect 1638 1653 1640 1655
rect 1643 1653 1645 1656
rect 1661 1653 1663 1655
rect 1290 1640 1292 1643
rect 778 1634 780 1636
rect 783 1631 785 1636
rect 859 1634 861 1636
rect 806 1630 808 1632
rect 864 1631 866 1636
rect 1290 1634 1292 1636
rect 887 1630 889 1632
rect 1173 1631 1175 1634
rect 1511 1631 1513 1645
rect 1527 1643 1529 1645
rect 1527 1631 1529 1633
rect 1543 1631 1545 1645
rect 1566 1640 1568 1645
rect 1571 1643 1573 1645
rect 1597 1643 1599 1645
rect 1562 1636 1568 1640
rect 1566 1631 1568 1636
rect 1571 1631 1573 1633
rect 1597 1631 1599 1633
rect 1618 1631 1620 1645
rect 1638 1640 1640 1645
rect 1643 1643 1645 1645
rect 1634 1636 1640 1640
rect 1638 1631 1640 1636
rect 1643 1631 1645 1633
rect 1661 1631 1663 1645
rect 1685 1644 1687 1658
rect 1792 1660 1794 1664
rect 1820 1666 1822 1668
rect 1797 1660 1799 1663
rect 1711 1649 1713 1652
rect 1716 1650 1718 1652
rect 1712 1645 1713 1649
rect 1711 1640 1713 1645
rect 1716 1640 1718 1642
rect 1685 1638 1687 1640
rect 1739 1636 1741 1658
rect 1766 1644 1768 1658
rect 1792 1649 1794 1652
rect 1797 1650 1799 1652
rect 1793 1645 1794 1649
rect 1792 1640 1794 1645
rect 1797 1640 1799 1642
rect 1766 1638 1768 1640
rect 1820 1636 1822 1658
rect 1711 1634 1713 1636
rect 1716 1631 1718 1636
rect 1792 1634 1794 1636
rect 1739 1630 1741 1632
rect 1797 1631 1799 1636
rect 1820 1630 1822 1632
rect 240 1625 242 1627
rect 578 1625 580 1627
rect 594 1623 596 1627
rect 610 1625 612 1627
rect 633 1625 635 1627
rect 595 1619 596 1623
rect 638 1622 640 1627
rect 664 1623 666 1627
rect 685 1625 687 1627
rect 705 1625 707 1627
rect 594 1616 596 1619
rect 639 1618 640 1622
rect 665 1619 666 1623
rect 710 1622 712 1627
rect 728 1625 730 1627
rect 1173 1625 1175 1627
rect 1511 1625 1513 1627
rect 1527 1623 1529 1627
rect 1543 1625 1545 1627
rect 1566 1625 1568 1627
rect 638 1616 640 1618
rect 664 1615 666 1619
rect 711 1618 712 1622
rect 1528 1619 1529 1623
rect 1571 1622 1573 1627
rect 1597 1623 1599 1627
rect 1618 1625 1620 1627
rect 1638 1625 1640 1627
rect 710 1616 712 1618
rect 1527 1616 1529 1619
rect 1572 1618 1573 1622
rect 1598 1619 1599 1623
rect 1643 1622 1645 1627
rect 1661 1625 1663 1627
rect 1571 1616 1573 1618
rect 1597 1615 1599 1619
rect 1644 1618 1645 1622
rect 1643 1616 1645 1618
rect 224 1602 226 1604
rect 240 1602 242 1605
rect 245 1602 247 1604
rect 261 1602 263 1605
rect 277 1602 279 1605
rect 298 1602 300 1605
rect 303 1602 305 1604
rect 319 1602 321 1604
rect 335 1602 337 1605
rect 340 1602 342 1604
rect 1157 1602 1159 1604
rect 1173 1602 1175 1605
rect 1178 1602 1180 1604
rect 1194 1602 1196 1605
rect 1210 1602 1212 1605
rect 1231 1602 1233 1605
rect 1236 1602 1238 1604
rect 1252 1602 1254 1604
rect 1268 1602 1270 1605
rect 1273 1602 1275 1604
rect 224 1575 226 1594
rect 240 1592 242 1594
rect 245 1585 247 1594
rect 261 1591 263 1594
rect 277 1592 279 1594
rect 298 1592 300 1594
rect 240 1575 242 1577
rect 245 1575 247 1578
rect 261 1575 263 1587
rect 303 1585 305 1594
rect 277 1575 279 1577
rect 298 1575 300 1577
rect 303 1575 305 1578
rect 319 1575 321 1594
rect 335 1592 337 1594
rect 340 1589 342 1594
rect 594 1593 596 1596
rect 638 1594 640 1596
rect 595 1589 596 1593
rect 639 1590 640 1594
rect 664 1593 666 1597
rect 710 1594 712 1596
rect 578 1585 580 1587
rect 594 1585 596 1589
rect 610 1585 612 1587
rect 633 1585 635 1587
rect 638 1585 640 1590
rect 665 1589 666 1593
rect 711 1590 712 1594
rect 664 1585 666 1589
rect 685 1585 687 1587
rect 705 1585 707 1587
rect 710 1585 712 1590
rect 728 1585 730 1587
rect 335 1575 337 1582
rect 340 1575 342 1585
rect 778 1584 780 1587
rect 783 1584 785 1587
rect 859 1584 861 1587
rect 864 1584 866 1587
rect 224 1569 226 1571
rect 240 1566 242 1571
rect 245 1569 247 1571
rect 261 1569 263 1571
rect 277 1566 279 1571
rect 298 1566 300 1571
rect 303 1569 305 1571
rect 319 1569 321 1571
rect 335 1568 337 1571
rect 340 1569 342 1571
rect 578 1567 580 1581
rect 594 1579 596 1581
rect 594 1567 596 1569
rect 610 1567 612 1581
rect 633 1576 635 1581
rect 638 1579 640 1581
rect 664 1579 666 1581
rect 629 1572 635 1576
rect 633 1567 635 1572
rect 638 1567 640 1569
rect 664 1567 666 1569
rect 685 1567 687 1581
rect 705 1576 707 1581
rect 710 1579 712 1581
rect 701 1572 707 1576
rect 705 1567 707 1572
rect 710 1567 712 1569
rect 728 1567 730 1581
rect 778 1568 780 1580
rect 783 1578 785 1580
rect 783 1568 785 1570
rect 859 1568 861 1580
rect 864 1578 866 1580
rect 1157 1575 1159 1594
rect 1173 1592 1175 1594
rect 1178 1585 1180 1594
rect 1194 1591 1196 1594
rect 1210 1592 1212 1594
rect 1231 1592 1233 1594
rect 1173 1575 1175 1577
rect 1178 1575 1180 1578
rect 1194 1575 1196 1587
rect 1236 1585 1238 1594
rect 1210 1575 1212 1577
rect 1231 1575 1233 1577
rect 1236 1575 1238 1578
rect 1252 1575 1254 1594
rect 1268 1592 1270 1594
rect 1273 1589 1275 1594
rect 1527 1593 1529 1596
rect 1571 1594 1573 1596
rect 1528 1589 1529 1593
rect 1572 1590 1573 1594
rect 1597 1593 1599 1597
rect 1643 1594 1645 1596
rect 1511 1585 1513 1587
rect 1527 1585 1529 1589
rect 1543 1585 1545 1587
rect 1566 1585 1568 1587
rect 1571 1585 1573 1590
rect 1598 1589 1599 1593
rect 1644 1590 1645 1594
rect 1597 1585 1599 1589
rect 1618 1585 1620 1587
rect 1638 1585 1640 1587
rect 1643 1585 1645 1590
rect 1661 1585 1663 1587
rect 1268 1575 1270 1582
rect 1273 1575 1275 1585
rect 1711 1584 1713 1587
rect 1716 1584 1718 1587
rect 1792 1584 1794 1587
rect 1797 1584 1799 1587
rect 864 1568 866 1570
rect 1157 1569 1159 1571
rect 1173 1566 1175 1571
rect 1178 1569 1180 1571
rect 1194 1569 1196 1571
rect 1210 1566 1212 1571
rect 1231 1566 1233 1571
rect 1236 1569 1238 1571
rect 1252 1569 1254 1571
rect 1268 1568 1270 1571
rect 1273 1569 1275 1571
rect 1511 1567 1513 1581
rect 1527 1579 1529 1581
rect 1527 1567 1529 1569
rect 1543 1567 1545 1581
rect 1566 1576 1568 1581
rect 1571 1579 1573 1581
rect 1597 1579 1599 1581
rect 1562 1572 1568 1576
rect 1566 1567 1568 1572
rect 1571 1567 1573 1569
rect 1597 1567 1599 1569
rect 1618 1567 1620 1581
rect 1638 1576 1640 1581
rect 1643 1579 1645 1581
rect 1634 1572 1640 1576
rect 1638 1567 1640 1572
rect 1643 1567 1645 1569
rect 1661 1567 1663 1581
rect 1711 1568 1713 1580
rect 1716 1578 1718 1580
rect 1716 1568 1718 1570
rect 1792 1568 1794 1580
rect 1797 1578 1799 1580
rect 1797 1568 1799 1570
rect 578 1557 580 1559
rect 594 1556 596 1559
rect 610 1557 612 1559
rect 633 1557 635 1559
rect 638 1556 640 1559
rect 664 1556 666 1559
rect 685 1556 687 1559
rect 705 1557 707 1559
rect 710 1556 712 1559
rect 728 1557 730 1559
rect 778 1558 780 1560
rect 664 1552 665 1556
rect 783 1555 785 1560
rect 859 1558 861 1560
rect 864 1555 866 1560
rect 1511 1557 1513 1559
rect 1527 1556 1529 1559
rect 1543 1557 1545 1559
rect 1566 1557 1568 1559
rect 1571 1556 1573 1559
rect 1597 1556 1599 1559
rect 1618 1556 1620 1559
rect 1638 1557 1640 1559
rect 1643 1556 1645 1559
rect 1661 1557 1663 1559
rect 1711 1558 1713 1560
rect 594 1549 596 1552
rect 638 1549 640 1552
rect 664 1549 666 1552
rect 710 1549 712 1552
rect 1597 1552 1598 1556
rect 1716 1555 1718 1560
rect 1792 1558 1794 1560
rect 1797 1555 1799 1560
rect 1527 1549 1529 1552
rect 1571 1549 1573 1552
rect 1597 1549 1599 1552
rect 1643 1549 1645 1552
rect 594 1528 596 1531
rect 638 1528 640 1531
rect 664 1528 666 1531
rect 710 1528 712 1531
rect 778 1528 780 1532
rect 806 1534 808 1536
rect 857 1534 859 1536
rect 783 1528 785 1531
rect 664 1524 665 1528
rect 578 1521 580 1523
rect 594 1521 596 1524
rect 610 1521 612 1523
rect 633 1521 635 1523
rect 638 1521 640 1524
rect 664 1521 666 1524
rect 685 1521 687 1524
rect 705 1521 707 1523
rect 710 1521 712 1524
rect 728 1521 730 1523
rect 883 1528 885 1532
rect 911 1534 913 1536
rect 888 1528 890 1531
rect 778 1517 780 1520
rect 783 1518 785 1520
rect 779 1513 780 1517
rect 578 1499 580 1513
rect 594 1511 596 1513
rect 594 1499 596 1501
rect 610 1499 612 1513
rect 633 1508 635 1513
rect 638 1511 640 1513
rect 664 1511 666 1513
rect 629 1504 635 1508
rect 633 1499 635 1504
rect 638 1499 640 1501
rect 664 1499 666 1501
rect 685 1499 687 1513
rect 705 1508 707 1513
rect 710 1511 712 1513
rect 701 1504 707 1508
rect 705 1499 707 1504
rect 710 1499 712 1501
rect 728 1499 730 1513
rect 778 1508 780 1513
rect 783 1508 785 1510
rect 806 1504 808 1526
rect 857 1512 859 1526
rect 1527 1528 1529 1531
rect 1571 1528 1573 1531
rect 1597 1528 1599 1531
rect 1643 1528 1645 1531
rect 1711 1528 1713 1532
rect 1739 1534 1741 1536
rect 1790 1534 1792 1536
rect 1716 1528 1718 1531
rect 883 1517 885 1520
rect 888 1518 890 1520
rect 884 1513 885 1517
rect 883 1508 885 1513
rect 888 1508 890 1510
rect 857 1506 859 1508
rect 911 1504 913 1526
rect 1597 1524 1598 1528
rect 1511 1521 1513 1523
rect 1527 1521 1529 1524
rect 1543 1521 1545 1523
rect 1566 1521 1568 1523
rect 1571 1521 1573 1524
rect 1597 1521 1599 1524
rect 1618 1521 1620 1524
rect 1638 1521 1640 1523
rect 1643 1521 1645 1524
rect 1661 1521 1663 1523
rect 1816 1528 1818 1532
rect 1844 1534 1846 1536
rect 1821 1528 1823 1531
rect 1711 1517 1713 1520
rect 1716 1518 1718 1520
rect 1712 1513 1713 1517
rect 778 1502 780 1504
rect 783 1499 785 1504
rect 883 1502 885 1504
rect 806 1498 808 1500
rect 888 1499 890 1504
rect 911 1498 913 1500
rect 1511 1499 1513 1513
rect 1527 1511 1529 1513
rect 1527 1499 1529 1501
rect 1543 1499 1545 1513
rect 1566 1508 1568 1513
rect 1571 1511 1573 1513
rect 1597 1511 1599 1513
rect 1562 1504 1568 1508
rect 1566 1499 1568 1504
rect 1571 1499 1573 1501
rect 1597 1499 1599 1501
rect 1618 1499 1620 1513
rect 1638 1508 1640 1513
rect 1643 1511 1645 1513
rect 1634 1504 1640 1508
rect 1638 1499 1640 1504
rect 1643 1499 1645 1501
rect 1661 1499 1663 1513
rect 1711 1508 1713 1513
rect 1716 1508 1718 1510
rect 1739 1504 1741 1526
rect 1790 1512 1792 1526
rect 1816 1517 1818 1520
rect 1821 1518 1823 1520
rect 1817 1513 1818 1517
rect 1816 1508 1818 1513
rect 1821 1508 1823 1510
rect 1790 1506 1792 1508
rect 1844 1504 1846 1526
rect 1711 1502 1713 1504
rect 1716 1499 1718 1504
rect 1816 1502 1818 1504
rect 1739 1498 1741 1500
rect 1821 1499 1823 1504
rect 1844 1498 1846 1500
rect 578 1493 580 1495
rect 594 1491 596 1495
rect 610 1493 612 1495
rect 633 1493 635 1495
rect 595 1487 596 1491
rect 638 1490 640 1495
rect 664 1491 666 1495
rect 685 1493 687 1495
rect 705 1493 707 1495
rect 594 1484 596 1487
rect 639 1486 640 1490
rect 665 1487 666 1491
rect 710 1490 712 1495
rect 728 1493 730 1495
rect 1511 1493 1513 1495
rect 1527 1491 1529 1495
rect 1543 1493 1545 1495
rect 1566 1493 1568 1495
rect 638 1484 640 1486
rect 664 1483 666 1487
rect 711 1486 712 1490
rect 1528 1487 1529 1491
rect 1571 1490 1573 1495
rect 1597 1491 1599 1495
rect 1618 1493 1620 1495
rect 1638 1493 1640 1495
rect 710 1484 712 1486
rect 1527 1484 1529 1487
rect 1572 1486 1573 1490
rect 1598 1487 1599 1491
rect 1643 1490 1645 1495
rect 1661 1493 1663 1495
rect 1571 1484 1573 1486
rect 1597 1483 1599 1487
rect 1644 1486 1645 1490
rect 1643 1484 1645 1486
rect 594 1461 596 1464
rect 638 1462 640 1464
rect 595 1457 596 1461
rect 639 1458 640 1462
rect 664 1461 666 1465
rect 710 1462 712 1464
rect 578 1453 580 1455
rect 594 1453 596 1457
rect 610 1453 612 1455
rect 633 1453 635 1455
rect 638 1453 640 1458
rect 665 1457 666 1461
rect 711 1458 712 1462
rect 1527 1461 1529 1464
rect 1571 1462 1573 1464
rect 664 1453 666 1457
rect 685 1453 687 1455
rect 705 1453 707 1455
rect 710 1453 712 1458
rect 1528 1457 1529 1461
rect 1572 1458 1573 1462
rect 1597 1461 1599 1465
rect 1643 1462 1645 1464
rect 728 1453 730 1455
rect 778 1453 780 1456
rect 783 1453 785 1456
rect 883 1453 885 1456
rect 888 1453 890 1456
rect 1511 1453 1513 1455
rect 1527 1453 1529 1457
rect 1543 1453 1545 1455
rect 1566 1453 1568 1455
rect 1571 1453 1573 1458
rect 1598 1457 1599 1461
rect 1644 1458 1645 1462
rect 1597 1453 1599 1457
rect 1618 1453 1620 1455
rect 1638 1453 1640 1455
rect 1643 1453 1645 1458
rect 1661 1453 1663 1455
rect 1711 1453 1713 1456
rect 1716 1453 1718 1456
rect 1816 1453 1818 1456
rect 1821 1453 1823 1456
rect 578 1435 580 1449
rect 594 1447 596 1449
rect 594 1435 596 1437
rect 610 1435 612 1449
rect 633 1444 635 1449
rect 638 1447 640 1449
rect 664 1447 666 1449
rect 629 1440 635 1444
rect 633 1435 635 1440
rect 638 1435 640 1437
rect 664 1435 666 1437
rect 685 1435 687 1449
rect 705 1444 707 1449
rect 710 1447 712 1449
rect 701 1440 707 1444
rect 705 1435 707 1440
rect 710 1435 712 1437
rect 728 1435 730 1449
rect 778 1437 780 1449
rect 783 1447 785 1449
rect 783 1437 785 1439
rect 883 1437 885 1449
rect 888 1447 890 1449
rect 888 1437 890 1439
rect 1511 1435 1513 1449
rect 1527 1447 1529 1449
rect 1527 1435 1529 1437
rect 1543 1435 1545 1449
rect 1566 1444 1568 1449
rect 1571 1447 1573 1449
rect 1597 1447 1599 1449
rect 1562 1440 1568 1444
rect 1566 1435 1568 1440
rect 1571 1435 1573 1437
rect 1597 1435 1599 1437
rect 1618 1435 1620 1449
rect 1638 1444 1640 1449
rect 1643 1447 1645 1449
rect 1634 1440 1640 1444
rect 1638 1435 1640 1440
rect 1643 1435 1645 1437
rect 1661 1435 1663 1449
rect 1711 1437 1713 1449
rect 1716 1447 1718 1449
rect 1716 1437 1718 1439
rect 1816 1437 1818 1449
rect 1821 1447 1823 1449
rect 1821 1437 1823 1439
rect 778 1427 780 1429
rect 578 1425 580 1427
rect 594 1424 596 1427
rect 610 1425 612 1427
rect 633 1425 635 1427
rect 638 1424 640 1427
rect 664 1424 666 1427
rect 685 1424 687 1427
rect 705 1425 707 1427
rect 710 1424 712 1427
rect 728 1425 730 1427
rect 783 1424 785 1429
rect 883 1427 885 1429
rect 888 1424 890 1429
rect 1711 1427 1713 1429
rect 1511 1425 1513 1427
rect 664 1420 665 1424
rect 1527 1424 1529 1427
rect 1543 1425 1545 1427
rect 1566 1425 1568 1427
rect 1571 1424 1573 1427
rect 1597 1424 1599 1427
rect 1618 1424 1620 1427
rect 1638 1425 1640 1427
rect 1643 1424 1645 1427
rect 1661 1425 1663 1427
rect 1716 1424 1718 1429
rect 1816 1427 1818 1429
rect 1821 1424 1823 1429
rect 1597 1420 1598 1424
rect 594 1417 596 1420
rect 638 1417 640 1420
rect 664 1417 666 1420
rect 710 1417 712 1420
rect 1527 1417 1529 1420
rect 1571 1417 1573 1420
rect 1597 1417 1599 1420
rect 1643 1417 1645 1420
rect 594 1396 596 1399
rect 638 1396 640 1399
rect 664 1396 666 1399
rect 710 1396 712 1399
rect 778 1396 780 1400
rect 806 1402 808 1404
rect 833 1402 835 1404
rect 783 1396 785 1399
rect 664 1392 665 1396
rect 578 1389 580 1391
rect 594 1389 596 1392
rect 610 1389 612 1391
rect 633 1389 635 1391
rect 638 1389 640 1392
rect 664 1389 666 1392
rect 685 1389 687 1392
rect 705 1389 707 1391
rect 710 1389 712 1392
rect 728 1389 730 1391
rect 859 1396 861 1400
rect 887 1402 889 1404
rect 923 1402 925 1404
rect 864 1396 866 1399
rect 778 1385 780 1388
rect 783 1386 785 1388
rect 779 1381 780 1385
rect 578 1367 580 1381
rect 594 1379 596 1381
rect 594 1367 596 1369
rect 610 1367 612 1381
rect 633 1376 635 1381
rect 638 1379 640 1381
rect 664 1379 666 1381
rect 629 1372 635 1376
rect 633 1367 635 1372
rect 638 1367 640 1369
rect 664 1367 666 1369
rect 685 1367 687 1381
rect 705 1376 707 1381
rect 710 1379 712 1381
rect 701 1372 707 1376
rect 705 1367 707 1372
rect 710 1367 712 1369
rect 728 1367 730 1381
rect 778 1376 780 1381
rect 783 1376 785 1378
rect 806 1372 808 1394
rect 833 1380 835 1394
rect 949 1396 951 1400
rect 977 1402 979 1404
rect 954 1396 956 1399
rect 859 1385 861 1388
rect 864 1386 866 1388
rect 860 1381 861 1385
rect 859 1376 861 1381
rect 864 1376 866 1378
rect 833 1374 835 1376
rect 887 1372 889 1394
rect 923 1380 925 1394
rect 1527 1396 1529 1399
rect 1571 1396 1573 1399
rect 1597 1396 1599 1399
rect 1643 1396 1645 1399
rect 1711 1396 1713 1400
rect 1739 1402 1741 1404
rect 1766 1402 1768 1404
rect 1716 1396 1718 1399
rect 949 1385 951 1388
rect 954 1386 956 1388
rect 950 1381 951 1385
rect 949 1376 951 1381
rect 954 1376 956 1378
rect 923 1374 925 1376
rect 977 1372 979 1394
rect 1597 1392 1598 1396
rect 1511 1389 1513 1391
rect 1527 1389 1529 1392
rect 1543 1389 1545 1391
rect 1566 1389 1568 1391
rect 1571 1389 1573 1392
rect 1597 1389 1599 1392
rect 1618 1389 1620 1392
rect 1638 1389 1640 1391
rect 1643 1389 1645 1392
rect 1661 1389 1663 1391
rect 1792 1396 1794 1400
rect 1820 1402 1822 1404
rect 1856 1402 1858 1404
rect 1797 1396 1799 1399
rect 1711 1385 1713 1388
rect 1716 1386 1718 1388
rect 1712 1381 1713 1385
rect 778 1370 780 1372
rect 783 1367 785 1372
rect 859 1370 861 1372
rect 806 1366 808 1368
rect 864 1367 866 1372
rect 949 1370 951 1372
rect 887 1366 889 1368
rect 954 1367 956 1372
rect 977 1366 979 1368
rect 1511 1367 1513 1381
rect 1527 1379 1529 1381
rect 1527 1367 1529 1369
rect 1543 1367 1545 1381
rect 1566 1376 1568 1381
rect 1571 1379 1573 1381
rect 1597 1379 1599 1381
rect 1562 1372 1568 1376
rect 1566 1367 1568 1372
rect 1571 1367 1573 1369
rect 1597 1367 1599 1369
rect 1618 1367 1620 1381
rect 1638 1376 1640 1381
rect 1643 1379 1645 1381
rect 1634 1372 1640 1376
rect 1638 1367 1640 1372
rect 1643 1367 1645 1369
rect 1661 1367 1663 1381
rect 1711 1376 1713 1381
rect 1716 1376 1718 1378
rect 1739 1372 1741 1394
rect 1766 1380 1768 1394
rect 1882 1396 1884 1400
rect 1910 1402 1912 1404
rect 1887 1396 1889 1399
rect 1792 1385 1794 1388
rect 1797 1386 1799 1388
rect 1793 1381 1794 1385
rect 1792 1376 1794 1381
rect 1797 1376 1799 1378
rect 1766 1374 1768 1376
rect 1820 1372 1822 1394
rect 1856 1380 1858 1394
rect 1882 1385 1884 1388
rect 1887 1386 1889 1388
rect 1883 1381 1884 1385
rect 1882 1376 1884 1381
rect 1887 1376 1889 1378
rect 1856 1374 1858 1376
rect 1910 1372 1912 1394
rect 1711 1370 1713 1372
rect 1716 1367 1718 1372
rect 1792 1370 1794 1372
rect 1739 1366 1741 1368
rect 1797 1367 1799 1372
rect 1882 1370 1884 1372
rect 1820 1366 1822 1368
rect 1887 1367 1889 1372
rect 1910 1366 1912 1368
rect 578 1361 580 1363
rect 594 1359 596 1363
rect 610 1361 612 1363
rect 633 1361 635 1363
rect 595 1355 596 1359
rect 638 1358 640 1363
rect 664 1359 666 1363
rect 685 1361 687 1363
rect 705 1361 707 1363
rect 594 1352 596 1355
rect 639 1354 640 1358
rect 665 1355 666 1359
rect 710 1358 712 1363
rect 728 1361 730 1363
rect 1511 1361 1513 1363
rect 1527 1359 1529 1363
rect 1543 1361 1545 1363
rect 1566 1361 1568 1363
rect 638 1352 640 1354
rect 664 1351 666 1355
rect 711 1354 712 1358
rect 1528 1355 1529 1359
rect 1571 1358 1573 1363
rect 1597 1359 1599 1363
rect 1618 1361 1620 1363
rect 1638 1361 1640 1363
rect 710 1352 712 1354
rect 1527 1352 1529 1355
rect 1572 1354 1573 1358
rect 1598 1355 1599 1359
rect 1643 1358 1645 1363
rect 1661 1361 1663 1363
rect 1571 1352 1573 1354
rect 1597 1351 1599 1355
rect 1644 1354 1645 1358
rect 1643 1352 1645 1354
rect 594 1329 596 1332
rect 638 1330 640 1332
rect 595 1325 596 1329
rect 639 1326 640 1330
rect 664 1329 666 1333
rect 710 1330 712 1332
rect 578 1321 580 1323
rect 594 1321 596 1325
rect 610 1321 612 1323
rect 633 1321 635 1323
rect 638 1321 640 1326
rect 665 1325 666 1329
rect 711 1326 712 1330
rect 1527 1329 1529 1332
rect 1571 1330 1573 1332
rect 664 1321 666 1325
rect 685 1321 687 1323
rect 705 1321 707 1323
rect 710 1321 712 1326
rect 1528 1325 1529 1329
rect 1572 1326 1573 1330
rect 1597 1329 1599 1333
rect 1643 1330 1645 1332
rect 728 1321 730 1323
rect 1511 1321 1513 1323
rect 1527 1321 1529 1325
rect 1543 1321 1545 1323
rect 1566 1321 1568 1323
rect 1571 1321 1573 1326
rect 1598 1325 1599 1329
rect 1644 1326 1645 1330
rect 1597 1321 1599 1325
rect 1618 1321 1620 1323
rect 1638 1321 1640 1323
rect 1643 1321 1645 1326
rect 1661 1321 1663 1323
rect 778 1318 780 1321
rect 783 1318 785 1321
rect 859 1318 861 1321
rect 864 1318 866 1321
rect 949 1318 951 1321
rect 954 1318 956 1321
rect 578 1303 580 1317
rect 594 1315 596 1317
rect 594 1303 596 1305
rect 610 1303 612 1317
rect 633 1312 635 1317
rect 638 1315 640 1317
rect 664 1315 666 1317
rect 629 1308 635 1312
rect 633 1303 635 1308
rect 638 1303 640 1305
rect 664 1303 666 1305
rect 685 1303 687 1317
rect 705 1312 707 1317
rect 710 1315 712 1317
rect 701 1308 707 1312
rect 705 1303 707 1308
rect 710 1303 712 1305
rect 728 1303 730 1317
rect 1711 1318 1713 1321
rect 1716 1318 1718 1321
rect 1792 1318 1794 1321
rect 1797 1318 1799 1321
rect 1882 1318 1884 1321
rect 1887 1318 1889 1321
rect 778 1302 780 1314
rect 783 1312 785 1314
rect 783 1302 785 1304
rect 859 1302 861 1314
rect 864 1312 866 1314
rect 864 1302 866 1304
rect 949 1302 951 1314
rect 954 1312 956 1314
rect 954 1302 956 1304
rect 1511 1303 1513 1317
rect 1527 1315 1529 1317
rect 1527 1303 1529 1305
rect 1543 1303 1545 1317
rect 1566 1312 1568 1317
rect 1571 1315 1573 1317
rect 1597 1315 1599 1317
rect 1562 1308 1568 1312
rect 1566 1303 1568 1308
rect 1571 1303 1573 1305
rect 1597 1303 1599 1305
rect 1618 1303 1620 1317
rect 1638 1312 1640 1317
rect 1643 1315 1645 1317
rect 1634 1308 1640 1312
rect 1638 1303 1640 1308
rect 1643 1303 1645 1305
rect 1661 1303 1663 1317
rect 578 1293 580 1295
rect 594 1292 596 1295
rect 610 1293 612 1295
rect 633 1293 635 1295
rect 638 1292 640 1295
rect 664 1292 666 1295
rect 685 1292 687 1295
rect 705 1293 707 1295
rect 710 1292 712 1295
rect 728 1293 730 1295
rect 1711 1302 1713 1314
rect 1716 1312 1718 1314
rect 1716 1302 1718 1304
rect 1792 1302 1794 1314
rect 1797 1312 1799 1314
rect 1797 1302 1799 1304
rect 1882 1302 1884 1314
rect 1887 1312 1889 1314
rect 1887 1302 1889 1304
rect 778 1292 780 1294
rect 664 1288 665 1292
rect 783 1289 785 1294
rect 859 1292 861 1294
rect 864 1289 866 1294
rect 949 1292 951 1294
rect 954 1289 956 1294
rect 1511 1293 1513 1295
rect 594 1285 596 1288
rect 638 1285 640 1288
rect 664 1285 666 1288
rect 710 1285 712 1288
rect 1527 1292 1529 1295
rect 1543 1293 1545 1295
rect 1566 1293 1568 1295
rect 1571 1292 1573 1295
rect 1597 1292 1599 1295
rect 1618 1292 1620 1295
rect 1638 1293 1640 1295
rect 1643 1292 1645 1295
rect 1661 1293 1663 1295
rect 1711 1292 1713 1294
rect 1597 1288 1598 1292
rect 1716 1289 1718 1294
rect 1792 1292 1794 1294
rect 1797 1289 1799 1294
rect 1882 1292 1884 1294
rect 1887 1289 1889 1294
rect 1527 1285 1529 1288
rect 1571 1285 1573 1288
rect 1597 1285 1599 1288
rect 1643 1285 1645 1288
rect 594 1264 596 1267
rect 638 1264 640 1267
rect 664 1264 666 1267
rect 710 1264 712 1267
rect 778 1264 780 1268
rect 806 1270 808 1272
rect 783 1264 785 1267
rect 664 1260 665 1264
rect 578 1257 580 1259
rect 594 1257 596 1260
rect 610 1257 612 1259
rect 633 1257 635 1259
rect 638 1257 640 1260
rect 664 1257 666 1260
rect 685 1257 687 1260
rect 705 1257 707 1259
rect 710 1257 712 1260
rect 728 1257 730 1259
rect 1527 1264 1529 1267
rect 1571 1264 1573 1267
rect 1597 1264 1599 1267
rect 1643 1264 1645 1267
rect 1711 1264 1713 1268
rect 1739 1270 1741 1272
rect 1716 1264 1718 1267
rect 778 1253 780 1256
rect 783 1254 785 1256
rect 779 1249 780 1253
rect 578 1235 580 1249
rect 594 1247 596 1249
rect 594 1235 596 1237
rect 610 1235 612 1249
rect 633 1244 635 1249
rect 638 1247 640 1249
rect 664 1247 666 1249
rect 629 1240 635 1244
rect 633 1235 635 1240
rect 638 1235 640 1237
rect 664 1235 666 1237
rect 685 1235 687 1249
rect 705 1244 707 1249
rect 710 1247 712 1249
rect 701 1240 707 1244
rect 705 1235 707 1240
rect 710 1235 712 1237
rect 728 1235 730 1249
rect 778 1244 780 1249
rect 783 1244 785 1246
rect 806 1240 808 1262
rect 1597 1260 1598 1264
rect 1511 1257 1513 1259
rect 1527 1257 1529 1260
rect 1543 1257 1545 1259
rect 1566 1257 1568 1259
rect 1571 1257 1573 1260
rect 1597 1257 1599 1260
rect 1618 1257 1620 1260
rect 1638 1257 1640 1259
rect 1643 1257 1645 1260
rect 1661 1257 1663 1259
rect 1711 1253 1713 1256
rect 1716 1254 1718 1256
rect 1712 1249 1713 1253
rect 778 1238 780 1240
rect 783 1235 785 1240
rect 806 1234 808 1236
rect 1511 1235 1513 1249
rect 1527 1247 1529 1249
rect 1527 1235 1529 1237
rect 1543 1235 1545 1249
rect 1566 1244 1568 1249
rect 1571 1247 1573 1249
rect 1597 1247 1599 1249
rect 1562 1240 1568 1244
rect 1566 1235 1568 1240
rect 1571 1235 1573 1237
rect 1597 1235 1599 1237
rect 1618 1235 1620 1249
rect 1638 1244 1640 1249
rect 1643 1247 1645 1249
rect 1634 1240 1640 1244
rect 1638 1235 1640 1240
rect 1643 1235 1645 1237
rect 1661 1235 1663 1249
rect 1711 1244 1713 1249
rect 1716 1244 1718 1246
rect 1739 1240 1741 1262
rect 1711 1238 1713 1240
rect 1716 1235 1718 1240
rect 1739 1234 1741 1236
rect 578 1229 580 1231
rect 594 1227 596 1231
rect 610 1229 612 1231
rect 633 1229 635 1231
rect 595 1223 596 1227
rect 638 1226 640 1231
rect 664 1227 666 1231
rect 685 1229 687 1231
rect 705 1229 707 1231
rect 594 1220 596 1223
rect 639 1222 640 1226
rect 665 1223 666 1227
rect 710 1226 712 1231
rect 728 1229 730 1231
rect 1511 1229 1513 1231
rect 1527 1227 1529 1231
rect 1543 1229 1545 1231
rect 1566 1229 1568 1231
rect 638 1220 640 1222
rect 664 1219 666 1223
rect 711 1222 712 1226
rect 1528 1223 1529 1227
rect 1571 1226 1573 1231
rect 1597 1227 1599 1231
rect 1618 1229 1620 1231
rect 1638 1229 1640 1231
rect 710 1220 712 1222
rect 1527 1220 1529 1223
rect 1572 1222 1573 1226
rect 1598 1223 1599 1227
rect 1643 1226 1645 1231
rect 1661 1229 1663 1231
rect 1571 1220 1573 1222
rect 1597 1219 1599 1223
rect 1644 1222 1645 1226
rect 1643 1220 1645 1222
rect 101 1202 103 1204
rect 106 1202 108 1205
rect 122 1202 124 1204
rect 138 1202 140 1204
rect 143 1202 145 1205
rect 164 1202 166 1205
rect 180 1202 182 1205
rect 196 1202 198 1204
rect 201 1202 203 1205
rect 217 1202 219 1204
rect 233 1202 235 1204
rect 238 1202 240 1205
rect 254 1202 256 1204
rect 270 1202 272 1204
rect 275 1202 277 1205
rect 296 1202 298 1205
rect 312 1202 314 1205
rect 328 1202 330 1204
rect 333 1202 335 1205
rect 349 1202 351 1204
rect 365 1202 367 1204
rect 370 1202 372 1205
rect 386 1202 388 1204
rect 402 1202 404 1204
rect 407 1202 409 1205
rect 428 1202 430 1205
rect 444 1202 446 1205
rect 460 1202 462 1204
rect 465 1202 467 1205
rect 481 1202 483 1204
rect 1034 1202 1036 1204
rect 1039 1202 1041 1205
rect 1055 1202 1057 1204
rect 1071 1202 1073 1204
rect 1076 1202 1078 1205
rect 1097 1202 1099 1205
rect 1113 1202 1115 1205
rect 1129 1202 1131 1204
rect 1134 1202 1136 1205
rect 1150 1202 1152 1204
rect 1166 1202 1168 1204
rect 1171 1202 1173 1205
rect 1187 1202 1189 1204
rect 1203 1202 1205 1204
rect 1208 1202 1210 1205
rect 1229 1202 1231 1205
rect 1245 1202 1247 1205
rect 1261 1202 1263 1204
rect 1266 1202 1268 1205
rect 1282 1202 1284 1204
rect 1298 1202 1300 1204
rect 1303 1202 1305 1205
rect 1319 1202 1321 1204
rect 1335 1202 1337 1204
rect 1340 1202 1342 1205
rect 1361 1202 1363 1205
rect 1377 1202 1379 1205
rect 1393 1202 1395 1204
rect 1398 1202 1400 1205
rect 1414 1202 1416 1204
rect 594 1197 596 1200
rect 638 1198 640 1200
rect 101 1189 103 1194
rect 106 1192 108 1194
rect 101 1175 103 1185
rect 106 1175 108 1182
rect 122 1175 124 1194
rect 138 1185 140 1194
rect 143 1192 145 1194
rect 164 1192 166 1194
rect 180 1191 182 1194
rect 138 1175 140 1178
rect 143 1175 145 1177
rect 164 1175 166 1177
rect 180 1175 182 1187
rect 196 1185 198 1194
rect 201 1192 203 1194
rect 196 1175 198 1178
rect 201 1175 203 1177
rect 217 1175 219 1194
rect 233 1191 235 1194
rect 238 1192 240 1194
rect 233 1175 235 1187
rect 238 1175 240 1182
rect 254 1175 256 1194
rect 270 1185 272 1194
rect 275 1192 277 1194
rect 296 1192 298 1194
rect 312 1191 314 1194
rect 270 1175 272 1178
rect 275 1175 277 1177
rect 296 1175 298 1177
rect 312 1175 314 1187
rect 328 1185 330 1194
rect 333 1192 335 1194
rect 328 1175 330 1178
rect 333 1175 335 1177
rect 349 1175 351 1194
rect 365 1191 367 1194
rect 370 1192 372 1194
rect 365 1175 367 1187
rect 370 1175 372 1182
rect 386 1175 388 1194
rect 402 1185 404 1194
rect 407 1192 409 1194
rect 428 1192 430 1194
rect 444 1191 446 1194
rect 402 1175 404 1178
rect 407 1175 409 1177
rect 428 1175 430 1177
rect 444 1175 446 1187
rect 460 1185 462 1194
rect 465 1192 467 1194
rect 481 1186 483 1194
rect 595 1193 596 1197
rect 639 1194 640 1198
rect 664 1197 666 1201
rect 710 1198 712 1200
rect 578 1189 580 1191
rect 594 1189 596 1193
rect 610 1189 612 1191
rect 633 1189 635 1191
rect 638 1189 640 1194
rect 665 1193 666 1197
rect 711 1194 712 1198
rect 855 1197 857 1200
rect 899 1198 901 1200
rect 664 1189 666 1193
rect 685 1189 687 1191
rect 705 1189 707 1191
rect 710 1189 712 1194
rect 856 1193 857 1197
rect 900 1194 901 1198
rect 925 1197 927 1201
rect 971 1198 973 1200
rect 728 1189 730 1191
rect 812 1189 814 1192
rect 830 1189 832 1192
rect 855 1189 857 1193
rect 871 1189 873 1191
rect 894 1189 896 1191
rect 899 1189 901 1194
rect 926 1193 927 1197
rect 972 1194 973 1198
rect 1527 1197 1529 1200
rect 1571 1198 1573 1200
rect 925 1189 927 1193
rect 946 1189 948 1191
rect 966 1189 968 1191
rect 971 1189 973 1194
rect 989 1189 991 1191
rect 1034 1189 1036 1194
rect 1039 1192 1041 1194
rect 460 1175 462 1178
rect 465 1175 467 1177
rect 481 1175 483 1182
rect 578 1171 580 1185
rect 594 1183 596 1185
rect 594 1171 596 1173
rect 610 1171 612 1185
rect 633 1180 635 1185
rect 638 1183 640 1185
rect 664 1183 666 1185
rect 629 1176 635 1180
rect 633 1171 635 1176
rect 638 1171 640 1173
rect 664 1171 666 1173
rect 685 1171 687 1185
rect 705 1180 707 1185
rect 710 1183 712 1185
rect 701 1176 707 1180
rect 705 1171 707 1176
rect 710 1171 712 1173
rect 728 1171 730 1185
rect 778 1182 780 1185
rect 783 1182 785 1185
rect 812 1180 814 1185
rect 101 1169 103 1171
rect 106 1168 108 1171
rect 122 1169 124 1171
rect 138 1169 140 1171
rect 143 1166 145 1171
rect 164 1166 166 1171
rect 180 1169 182 1171
rect 196 1169 198 1171
rect 201 1166 203 1171
rect 217 1169 219 1171
rect 233 1169 235 1171
rect 238 1168 240 1171
rect 254 1169 256 1171
rect 270 1169 272 1171
rect 275 1166 277 1171
rect 296 1166 298 1171
rect 312 1169 314 1171
rect 328 1169 330 1171
rect 333 1166 335 1171
rect 349 1169 351 1171
rect 365 1169 367 1171
rect 370 1168 372 1171
rect 386 1169 388 1171
rect 402 1169 404 1171
rect 407 1166 409 1171
rect 428 1166 430 1171
rect 444 1169 446 1171
rect 460 1169 462 1171
rect 465 1166 467 1171
rect 481 1169 483 1171
rect 778 1166 780 1178
rect 783 1176 785 1178
rect 812 1171 814 1176
rect 830 1171 832 1185
rect 855 1183 857 1185
rect 855 1171 857 1173
rect 871 1171 873 1185
rect 894 1180 896 1185
rect 899 1183 901 1185
rect 925 1183 927 1185
rect 890 1176 896 1180
rect 894 1171 896 1176
rect 899 1171 901 1173
rect 925 1171 927 1173
rect 946 1171 948 1185
rect 966 1180 968 1185
rect 971 1183 973 1185
rect 962 1176 968 1180
rect 966 1171 968 1176
rect 971 1171 973 1173
rect 989 1171 991 1185
rect 1034 1175 1036 1185
rect 1039 1175 1041 1182
rect 1055 1175 1057 1194
rect 1071 1185 1073 1194
rect 1076 1192 1078 1194
rect 1097 1192 1099 1194
rect 1113 1191 1115 1194
rect 1071 1175 1073 1178
rect 1076 1175 1078 1177
rect 1097 1175 1099 1177
rect 1113 1175 1115 1187
rect 1129 1185 1131 1194
rect 1134 1192 1136 1194
rect 1129 1175 1131 1178
rect 1134 1175 1136 1177
rect 1150 1175 1152 1194
rect 1166 1191 1168 1194
rect 1171 1192 1173 1194
rect 1166 1175 1168 1187
rect 1171 1175 1173 1182
rect 1187 1175 1189 1194
rect 1203 1185 1205 1194
rect 1208 1192 1210 1194
rect 1229 1192 1231 1194
rect 1245 1191 1247 1194
rect 1203 1175 1205 1178
rect 1208 1175 1210 1177
rect 1229 1175 1231 1177
rect 1245 1175 1247 1187
rect 1261 1185 1263 1194
rect 1266 1192 1268 1194
rect 1261 1175 1263 1178
rect 1266 1175 1268 1177
rect 1282 1175 1284 1194
rect 1298 1191 1300 1194
rect 1303 1192 1305 1194
rect 1298 1175 1300 1187
rect 1303 1175 1305 1182
rect 1319 1175 1321 1194
rect 1335 1185 1337 1194
rect 1340 1192 1342 1194
rect 1361 1192 1363 1194
rect 1377 1191 1379 1194
rect 1335 1175 1337 1178
rect 1340 1175 1342 1177
rect 1361 1175 1363 1177
rect 1377 1175 1379 1187
rect 1393 1185 1395 1194
rect 1398 1192 1400 1194
rect 1414 1186 1416 1194
rect 1528 1193 1529 1197
rect 1572 1194 1573 1198
rect 1597 1197 1599 1201
rect 1643 1198 1645 1200
rect 1511 1189 1513 1191
rect 1527 1189 1529 1193
rect 1543 1189 1545 1191
rect 1566 1189 1568 1191
rect 1571 1189 1573 1194
rect 1598 1193 1599 1197
rect 1644 1194 1645 1198
rect 1788 1197 1790 1200
rect 1832 1198 1834 1200
rect 1597 1189 1599 1193
rect 1618 1189 1620 1191
rect 1638 1189 1640 1191
rect 1643 1189 1645 1194
rect 1789 1193 1790 1197
rect 1833 1194 1834 1198
rect 1858 1197 1860 1201
rect 1904 1198 1906 1200
rect 1661 1189 1663 1191
rect 1745 1189 1747 1192
rect 1763 1189 1765 1192
rect 1788 1189 1790 1193
rect 1804 1189 1806 1191
rect 1827 1189 1829 1191
rect 1832 1189 1834 1194
rect 1859 1193 1860 1197
rect 1905 1194 1906 1198
rect 1858 1189 1860 1193
rect 1879 1189 1881 1191
rect 1899 1189 1901 1191
rect 1904 1189 1906 1194
rect 1922 1189 1924 1191
rect 1393 1175 1395 1178
rect 1398 1175 1400 1177
rect 1414 1175 1416 1182
rect 1511 1171 1513 1185
rect 1527 1183 1529 1185
rect 1527 1171 1529 1173
rect 1543 1171 1545 1185
rect 1566 1180 1568 1185
rect 1571 1183 1573 1185
rect 1597 1183 1599 1185
rect 1562 1176 1568 1180
rect 1566 1171 1568 1176
rect 1571 1171 1573 1173
rect 1597 1171 1599 1173
rect 1618 1171 1620 1185
rect 1638 1180 1640 1185
rect 1643 1183 1645 1185
rect 1634 1176 1640 1180
rect 1638 1171 1640 1176
rect 1643 1171 1645 1173
rect 1661 1171 1663 1185
rect 1711 1182 1713 1185
rect 1716 1182 1718 1185
rect 1745 1180 1747 1185
rect 783 1166 785 1168
rect 578 1161 580 1163
rect 594 1160 596 1163
rect 610 1161 612 1163
rect 633 1161 635 1163
rect 638 1160 640 1163
rect 664 1160 666 1163
rect 685 1160 687 1163
rect 705 1161 707 1163
rect 710 1160 712 1163
rect 728 1161 730 1163
rect 664 1156 665 1160
rect 1034 1169 1036 1171
rect 1039 1168 1041 1171
rect 1055 1169 1057 1171
rect 1071 1169 1073 1171
rect 1076 1166 1078 1171
rect 1097 1166 1099 1171
rect 1113 1169 1115 1171
rect 1129 1169 1131 1171
rect 1134 1166 1136 1171
rect 1150 1169 1152 1171
rect 1166 1169 1168 1171
rect 812 1160 814 1163
rect 830 1160 832 1163
rect 855 1160 857 1163
rect 871 1161 873 1163
rect 894 1161 896 1163
rect 899 1160 901 1163
rect 925 1160 927 1163
rect 946 1160 948 1163
rect 966 1161 968 1163
rect 971 1160 973 1163
rect 989 1161 991 1163
rect 1171 1168 1173 1171
rect 1187 1169 1189 1171
rect 1203 1169 1205 1171
rect 1208 1166 1210 1171
rect 1229 1166 1231 1171
rect 1245 1169 1247 1171
rect 1261 1169 1263 1171
rect 1266 1166 1268 1171
rect 1282 1169 1284 1171
rect 1298 1169 1300 1171
rect 1303 1168 1305 1171
rect 1319 1169 1321 1171
rect 1335 1169 1337 1171
rect 1340 1166 1342 1171
rect 1361 1166 1363 1171
rect 1377 1169 1379 1171
rect 1393 1169 1395 1171
rect 1398 1166 1400 1171
rect 1414 1169 1416 1171
rect 1711 1166 1713 1178
rect 1716 1176 1718 1178
rect 1745 1171 1747 1176
rect 1763 1171 1765 1185
rect 1788 1183 1790 1185
rect 1788 1171 1790 1173
rect 1804 1171 1806 1185
rect 1827 1180 1829 1185
rect 1832 1183 1834 1185
rect 1858 1183 1860 1185
rect 1823 1176 1829 1180
rect 1827 1171 1829 1176
rect 1832 1171 1834 1173
rect 1858 1171 1860 1173
rect 1879 1171 1881 1185
rect 1899 1180 1901 1185
rect 1904 1183 1906 1185
rect 1895 1176 1901 1180
rect 1899 1171 1901 1176
rect 1904 1171 1906 1173
rect 1922 1171 1924 1185
rect 1716 1166 1718 1168
rect 1511 1161 1513 1163
rect 1527 1160 1529 1163
rect 1543 1161 1545 1163
rect 1566 1161 1568 1163
rect 1571 1160 1573 1163
rect 1597 1160 1599 1163
rect 1618 1160 1620 1163
rect 1638 1161 1640 1163
rect 1643 1160 1645 1163
rect 1661 1161 1663 1163
rect 778 1156 780 1158
rect 594 1153 596 1156
rect 638 1153 640 1156
rect 664 1153 666 1156
rect 710 1153 712 1156
rect 783 1153 785 1158
rect 925 1156 926 1160
rect 855 1153 857 1156
rect 899 1153 901 1156
rect 925 1153 927 1156
rect 971 1153 973 1156
rect 1597 1156 1598 1160
rect 1745 1160 1747 1163
rect 1763 1160 1765 1163
rect 1788 1160 1790 1163
rect 1804 1161 1806 1163
rect 1827 1161 1829 1163
rect 1832 1160 1834 1163
rect 1858 1160 1860 1163
rect 1879 1160 1881 1163
rect 1899 1161 1901 1163
rect 1904 1160 1906 1163
rect 1922 1161 1924 1163
rect 1711 1156 1713 1158
rect 1527 1153 1529 1156
rect 1571 1153 1573 1156
rect 1597 1153 1599 1156
rect 1643 1153 1645 1156
rect 1716 1153 1718 1158
rect 1858 1156 1859 1160
rect 1788 1153 1790 1156
rect 1832 1153 1834 1156
rect 1858 1153 1860 1156
rect 1904 1153 1906 1156
rect 216 1131 218 1134
rect 240 1131 242 1134
rect 1149 1131 1151 1134
rect 1173 1131 1175 1134
rect 998 1129 1001 1131
rect 1005 1129 1008 1131
rect 216 1125 218 1127
rect 240 1125 242 1127
rect 1931 1129 1934 1131
rect 1938 1129 1941 1131
rect 1149 1125 1151 1127
rect 1173 1125 1175 1127
rect 236 1120 238 1122
rect 1169 1120 1171 1122
rect 236 1113 238 1116
rect 1169 1113 1171 1116
rect 225 1102 227 1104
rect 231 1102 250 1104
rect 1158 1102 1160 1104
rect 1164 1102 1183 1104
rect 216 1097 218 1099
rect 240 1097 242 1099
rect 1149 1097 1151 1099
rect 1173 1097 1175 1099
rect 216 1090 218 1093
rect 240 1090 242 1093
rect 872 1092 874 1094
rect 877 1092 879 1095
rect 893 1092 895 1094
rect 909 1092 911 1094
rect 914 1092 916 1095
rect 935 1092 937 1095
rect 951 1092 953 1095
rect 967 1092 969 1094
rect 972 1092 974 1095
rect 988 1092 990 1094
rect 1149 1090 1151 1093
rect 1173 1090 1175 1093
rect 1805 1092 1807 1094
rect 1810 1092 1812 1095
rect 1826 1092 1828 1094
rect 1842 1092 1844 1094
rect 1847 1092 1849 1095
rect 1868 1092 1870 1095
rect 1884 1092 1886 1095
rect 1900 1092 1902 1094
rect 1905 1092 1907 1095
rect 1921 1092 1923 1094
rect 872 1079 874 1084
rect 877 1082 879 1084
rect 872 1065 874 1075
rect 877 1065 879 1072
rect 893 1065 895 1084
rect 909 1075 911 1084
rect 914 1082 916 1084
rect 935 1082 937 1084
rect 951 1081 953 1084
rect 909 1065 911 1068
rect 914 1065 916 1067
rect 935 1065 937 1067
rect 951 1065 953 1077
rect 967 1075 969 1084
rect 972 1082 974 1084
rect 967 1065 969 1068
rect 972 1065 974 1067
rect 988 1065 990 1084
rect 1805 1079 1807 1084
rect 1810 1082 1812 1084
rect 1805 1065 1807 1075
rect 1810 1065 1812 1072
rect 1826 1065 1828 1084
rect 1842 1075 1844 1084
rect 1847 1082 1849 1084
rect 1868 1082 1870 1084
rect 1884 1081 1886 1084
rect 1842 1065 1844 1068
rect 1847 1065 1849 1067
rect 1868 1065 1870 1067
rect 1884 1065 1886 1077
rect 1900 1075 1902 1084
rect 1905 1082 1907 1084
rect 1900 1065 1902 1068
rect 1905 1065 1907 1067
rect 1921 1065 1923 1084
rect 101 1062 103 1064
rect 106 1062 108 1065
rect 122 1062 124 1064
rect 138 1062 140 1064
rect 143 1062 145 1065
rect 164 1062 166 1065
rect 180 1062 182 1065
rect 196 1062 198 1064
rect 201 1062 203 1065
rect 217 1062 219 1064
rect 233 1062 235 1064
rect 238 1062 240 1065
rect 254 1062 256 1064
rect 270 1062 272 1064
rect 275 1062 277 1065
rect 296 1062 298 1065
rect 312 1062 314 1065
rect 328 1062 330 1064
rect 333 1062 335 1065
rect 349 1062 351 1064
rect 365 1062 367 1064
rect 370 1062 372 1065
rect 386 1062 388 1064
rect 402 1062 404 1064
rect 407 1062 409 1065
rect 428 1062 430 1065
rect 444 1062 446 1065
rect 460 1062 462 1064
rect 465 1062 467 1065
rect 481 1062 483 1064
rect 1034 1062 1036 1064
rect 1039 1062 1041 1065
rect 1055 1062 1057 1064
rect 1071 1062 1073 1064
rect 1076 1062 1078 1065
rect 1097 1062 1099 1065
rect 1113 1062 1115 1065
rect 1129 1062 1131 1064
rect 1134 1062 1136 1065
rect 1150 1062 1152 1064
rect 1166 1062 1168 1064
rect 1171 1062 1173 1065
rect 1187 1062 1189 1064
rect 1203 1062 1205 1064
rect 1208 1062 1210 1065
rect 1229 1062 1231 1065
rect 1245 1062 1247 1065
rect 1261 1062 1263 1064
rect 1266 1062 1268 1065
rect 1282 1062 1284 1064
rect 1298 1062 1300 1064
rect 1303 1062 1305 1065
rect 1319 1062 1321 1064
rect 1335 1062 1337 1064
rect 1340 1062 1342 1065
rect 1361 1062 1363 1065
rect 1377 1062 1379 1065
rect 1393 1062 1395 1064
rect 1398 1062 1400 1065
rect 1414 1062 1416 1064
rect 872 1059 874 1061
rect 877 1058 879 1061
rect 893 1059 895 1061
rect 909 1059 911 1061
rect 914 1056 916 1061
rect 935 1056 937 1061
rect 951 1059 953 1061
rect 967 1059 969 1061
rect 972 1056 974 1061
rect 988 1059 990 1061
rect 101 1049 103 1054
rect 106 1052 108 1054
rect 101 1035 103 1045
rect 106 1035 108 1042
rect 122 1035 124 1054
rect 138 1045 140 1054
rect 143 1052 145 1054
rect 164 1052 166 1054
rect 180 1051 182 1054
rect 138 1035 140 1038
rect 143 1035 145 1037
rect 164 1035 166 1037
rect 180 1035 182 1047
rect 196 1045 198 1054
rect 201 1052 203 1054
rect 196 1035 198 1038
rect 201 1035 203 1037
rect 217 1035 219 1054
rect 233 1051 235 1054
rect 238 1052 240 1054
rect 233 1035 235 1047
rect 238 1035 240 1042
rect 254 1035 256 1054
rect 270 1045 272 1054
rect 275 1052 277 1054
rect 296 1052 298 1054
rect 312 1051 314 1054
rect 270 1035 272 1038
rect 275 1035 277 1037
rect 296 1035 298 1037
rect 312 1035 314 1047
rect 328 1045 330 1054
rect 333 1052 335 1054
rect 328 1035 330 1038
rect 333 1035 335 1037
rect 349 1035 351 1054
rect 365 1051 367 1054
rect 370 1052 372 1054
rect 365 1035 367 1047
rect 370 1035 372 1042
rect 386 1035 388 1054
rect 402 1045 404 1054
rect 407 1052 409 1054
rect 428 1052 430 1054
rect 444 1051 446 1054
rect 402 1035 404 1038
rect 407 1035 409 1037
rect 428 1035 430 1037
rect 444 1035 446 1047
rect 460 1045 462 1054
rect 465 1052 467 1054
rect 481 1046 483 1054
rect 1805 1059 1807 1061
rect 1810 1058 1812 1061
rect 1826 1059 1828 1061
rect 1842 1059 1844 1061
rect 1847 1056 1849 1061
rect 1868 1056 1870 1061
rect 1884 1059 1886 1061
rect 1900 1059 1902 1061
rect 1905 1056 1907 1061
rect 1921 1059 1923 1061
rect 1034 1049 1036 1054
rect 1039 1052 1041 1054
rect 460 1035 462 1038
rect 465 1035 467 1037
rect 481 1035 483 1042
rect 1034 1035 1036 1045
rect 1039 1035 1041 1042
rect 1055 1035 1057 1054
rect 1071 1045 1073 1054
rect 1076 1052 1078 1054
rect 1097 1052 1099 1054
rect 1113 1051 1115 1054
rect 1071 1035 1073 1038
rect 1076 1035 1078 1037
rect 1097 1035 1099 1037
rect 1113 1035 1115 1047
rect 1129 1045 1131 1054
rect 1134 1052 1136 1054
rect 1129 1035 1131 1038
rect 1134 1035 1136 1037
rect 1150 1035 1152 1054
rect 1166 1051 1168 1054
rect 1171 1052 1173 1054
rect 1166 1035 1168 1047
rect 1171 1035 1173 1042
rect 1187 1035 1189 1054
rect 1203 1045 1205 1054
rect 1208 1052 1210 1054
rect 1229 1052 1231 1054
rect 1245 1051 1247 1054
rect 1203 1035 1205 1038
rect 1208 1035 1210 1037
rect 1229 1035 1231 1037
rect 1245 1035 1247 1047
rect 1261 1045 1263 1054
rect 1266 1052 1268 1054
rect 1261 1035 1263 1038
rect 1266 1035 1268 1037
rect 1282 1035 1284 1054
rect 1298 1051 1300 1054
rect 1303 1052 1305 1054
rect 1298 1035 1300 1047
rect 1303 1035 1305 1042
rect 1319 1035 1321 1054
rect 1335 1045 1337 1054
rect 1340 1052 1342 1054
rect 1361 1052 1363 1054
rect 1377 1051 1379 1054
rect 1335 1035 1337 1038
rect 1340 1035 1342 1037
rect 1361 1035 1363 1037
rect 1377 1035 1379 1047
rect 1393 1045 1395 1054
rect 1398 1052 1400 1054
rect 1414 1046 1416 1054
rect 1393 1035 1395 1038
rect 1398 1035 1400 1037
rect 1414 1035 1416 1042
rect 101 1029 103 1031
rect 106 1028 108 1031
rect 122 1029 124 1031
rect 138 1029 140 1031
rect 143 1026 145 1031
rect 164 1026 166 1031
rect 180 1029 182 1031
rect 196 1029 198 1031
rect 201 1026 203 1031
rect 217 1029 219 1031
rect 233 1029 235 1031
rect 238 1028 240 1031
rect 254 1029 256 1031
rect 270 1029 272 1031
rect 275 1026 277 1031
rect 296 1026 298 1031
rect 312 1029 314 1031
rect 328 1029 330 1031
rect 333 1026 335 1031
rect 349 1029 351 1031
rect 365 1029 367 1031
rect 370 1028 372 1031
rect 386 1029 388 1031
rect 402 1029 404 1031
rect 407 1026 409 1031
rect 428 1026 430 1031
rect 444 1029 446 1031
rect 460 1029 462 1031
rect 465 1026 467 1031
rect 481 1029 483 1031
rect 1034 1029 1036 1031
rect 1039 1028 1041 1031
rect 1055 1029 1057 1031
rect 1071 1029 1073 1031
rect 1076 1026 1078 1031
rect 1097 1026 1099 1031
rect 1113 1029 1115 1031
rect 1129 1029 1131 1031
rect 1134 1026 1136 1031
rect 1150 1029 1152 1031
rect 1166 1029 1168 1031
rect 1171 1028 1173 1031
rect 1187 1029 1189 1031
rect 1203 1029 1205 1031
rect 1208 1026 1210 1031
rect 1229 1026 1231 1031
rect 1245 1029 1247 1031
rect 1261 1029 1263 1031
rect 1266 1026 1268 1031
rect 1282 1029 1284 1031
rect 1298 1029 1300 1031
rect 1303 1028 1305 1031
rect 1319 1029 1321 1031
rect 1335 1029 1337 1031
rect 1340 1026 1342 1031
rect 1361 1026 1363 1031
rect 1377 1029 1379 1031
rect 1393 1029 1395 1031
rect 1398 1026 1400 1031
rect 1414 1029 1416 1031
rect 872 1006 874 1008
rect 877 1006 879 1009
rect 893 1006 895 1008
rect 909 1006 911 1008
rect 914 1006 916 1009
rect 935 1006 937 1009
rect 951 1006 953 1009
rect 967 1006 969 1008
rect 972 1006 974 1009
rect 988 1006 990 1008
rect 1805 1006 1807 1008
rect 1810 1006 1812 1009
rect 1826 1006 1828 1008
rect 1842 1006 1844 1008
rect 1847 1006 1849 1009
rect 1868 1006 1870 1009
rect 1884 1006 1886 1009
rect 1900 1006 1902 1008
rect 1905 1006 1907 1009
rect 1921 1006 1923 1008
rect 872 993 874 998
rect 877 996 879 998
rect 872 979 874 989
rect 877 979 879 986
rect 893 979 895 998
rect 909 989 911 998
rect 914 996 916 998
rect 935 996 937 998
rect 951 995 953 998
rect 909 979 911 982
rect 914 979 916 981
rect 935 979 937 981
rect 951 979 953 991
rect 967 989 969 998
rect 972 996 974 998
rect 967 979 969 982
rect 972 979 974 981
rect 988 979 990 998
rect 1805 993 1807 998
rect 1810 996 1812 998
rect 1010 985 1013 987
rect 1017 985 1020 987
rect 1805 979 1807 989
rect 1810 979 1812 986
rect 1826 979 1828 998
rect 1842 989 1844 998
rect 1847 996 1849 998
rect 1868 996 1870 998
rect 1884 995 1886 998
rect 1842 979 1844 982
rect 1847 979 1849 981
rect 1868 979 1870 981
rect 1884 979 1886 991
rect 1900 989 1902 998
rect 1905 996 1907 998
rect 1900 979 1902 982
rect 1905 979 1907 981
rect 1921 979 1923 998
rect 1943 985 1946 987
rect 1950 985 1953 987
rect 101 976 103 978
rect 106 976 108 979
rect 122 976 124 978
rect 138 976 140 978
rect 143 976 145 979
rect 164 976 166 979
rect 180 976 182 979
rect 196 976 198 978
rect 201 976 203 979
rect 217 976 219 978
rect 233 976 235 978
rect 238 976 240 979
rect 254 976 256 978
rect 270 976 272 978
rect 275 976 277 979
rect 296 976 298 979
rect 312 976 314 979
rect 328 976 330 978
rect 333 976 335 979
rect 349 976 351 978
rect 365 976 367 978
rect 370 976 372 979
rect 386 976 388 978
rect 402 976 404 978
rect 407 976 409 979
rect 428 976 430 979
rect 444 976 446 979
rect 460 976 462 978
rect 465 976 467 979
rect 481 976 483 978
rect 1034 976 1036 978
rect 1039 976 1041 979
rect 1055 976 1057 978
rect 1071 976 1073 978
rect 1076 976 1078 979
rect 1097 976 1099 979
rect 1113 976 1115 979
rect 1129 976 1131 978
rect 1134 976 1136 979
rect 1150 976 1152 978
rect 1166 976 1168 978
rect 1171 976 1173 979
rect 1187 976 1189 978
rect 1203 976 1205 978
rect 1208 976 1210 979
rect 1229 976 1231 979
rect 1245 976 1247 979
rect 1261 976 1263 978
rect 1266 976 1268 979
rect 1282 976 1284 978
rect 1298 976 1300 978
rect 1303 976 1305 979
rect 1319 976 1321 978
rect 1335 976 1337 978
rect 1340 976 1342 979
rect 1361 976 1363 979
rect 1377 976 1379 979
rect 1393 976 1395 978
rect 1398 976 1400 979
rect 1414 976 1416 978
rect 872 973 874 975
rect 877 972 879 975
rect 893 973 895 975
rect 909 973 911 975
rect 914 970 916 975
rect 935 970 937 975
rect 951 973 953 975
rect 967 973 969 975
rect 972 970 974 975
rect 988 973 990 975
rect 101 963 103 968
rect 106 966 108 968
rect 101 949 103 959
rect 106 949 108 956
rect 122 949 124 968
rect 138 959 140 968
rect 143 966 145 968
rect 164 966 166 968
rect 180 965 182 968
rect 138 949 140 952
rect 143 949 145 951
rect 164 949 166 951
rect 180 949 182 961
rect 196 959 198 968
rect 201 966 203 968
rect 196 949 198 952
rect 201 949 203 951
rect 217 949 219 968
rect 233 965 235 968
rect 238 966 240 968
rect 233 949 235 961
rect 238 949 240 956
rect 254 949 256 968
rect 270 959 272 968
rect 275 966 277 968
rect 296 966 298 968
rect 312 965 314 968
rect 270 949 272 952
rect 275 949 277 951
rect 296 949 298 951
rect 312 949 314 961
rect 328 959 330 968
rect 333 966 335 968
rect 328 949 330 952
rect 333 949 335 951
rect 349 949 351 968
rect 365 965 367 968
rect 370 966 372 968
rect 365 949 367 961
rect 370 949 372 956
rect 386 949 388 968
rect 402 959 404 968
rect 407 966 409 968
rect 428 966 430 968
rect 444 965 446 968
rect 402 949 404 952
rect 407 949 409 951
rect 428 949 430 951
rect 444 949 446 961
rect 460 959 462 968
rect 465 966 467 968
rect 481 960 483 968
rect 1805 973 1807 975
rect 1810 972 1812 975
rect 1826 973 1828 975
rect 1842 973 1844 975
rect 1847 970 1849 975
rect 1868 970 1870 975
rect 1884 973 1886 975
rect 1900 973 1902 975
rect 1905 970 1907 975
rect 1921 973 1923 975
rect 1034 963 1036 968
rect 1039 966 1041 968
rect 460 949 462 952
rect 465 949 467 951
rect 481 949 483 956
rect 1034 949 1036 959
rect 1039 949 1041 956
rect 1055 949 1057 968
rect 1071 959 1073 968
rect 1076 966 1078 968
rect 1097 966 1099 968
rect 1113 965 1115 968
rect 1071 949 1073 952
rect 1076 949 1078 951
rect 1097 949 1099 951
rect 1113 949 1115 961
rect 1129 959 1131 968
rect 1134 966 1136 968
rect 1129 949 1131 952
rect 1134 949 1136 951
rect 1150 949 1152 968
rect 1166 965 1168 968
rect 1171 966 1173 968
rect 1166 949 1168 961
rect 1171 949 1173 956
rect 1187 949 1189 968
rect 1203 959 1205 968
rect 1208 966 1210 968
rect 1229 966 1231 968
rect 1245 965 1247 968
rect 1203 949 1205 952
rect 1208 949 1210 951
rect 1229 949 1231 951
rect 1245 949 1247 961
rect 1261 959 1263 968
rect 1266 966 1268 968
rect 1261 949 1263 952
rect 1266 949 1268 951
rect 1282 949 1284 968
rect 1298 965 1300 968
rect 1303 966 1305 968
rect 1298 949 1300 961
rect 1303 949 1305 956
rect 1319 949 1321 968
rect 1335 959 1337 968
rect 1340 966 1342 968
rect 1361 966 1363 968
rect 1377 965 1379 968
rect 1335 949 1337 952
rect 1340 949 1342 951
rect 1361 949 1363 951
rect 1377 949 1379 961
rect 1393 959 1395 968
rect 1398 966 1400 968
rect 1414 960 1416 968
rect 1393 949 1395 952
rect 1398 949 1400 951
rect 1414 949 1416 956
rect 101 943 103 945
rect 106 942 108 945
rect 122 943 124 945
rect 138 943 140 945
rect 143 940 145 945
rect 164 940 166 945
rect 180 943 182 945
rect 196 943 198 945
rect 201 940 203 945
rect 217 943 219 945
rect 233 943 235 945
rect 238 942 240 945
rect 254 943 256 945
rect 270 943 272 945
rect 275 940 277 945
rect 296 940 298 945
rect 312 943 314 945
rect 328 943 330 945
rect 333 940 335 945
rect 349 943 351 945
rect 365 943 367 945
rect 370 942 372 945
rect 386 943 388 945
rect 402 943 404 945
rect 407 940 409 945
rect 428 940 430 945
rect 444 943 446 945
rect 460 943 462 945
rect 465 940 467 945
rect 481 943 483 945
rect 1034 943 1036 945
rect 1039 942 1041 945
rect 1055 943 1057 945
rect 1071 943 1073 945
rect 1076 940 1078 945
rect 1097 940 1099 945
rect 1113 943 1115 945
rect 1129 943 1131 945
rect 1134 940 1136 945
rect 1150 943 1152 945
rect 1166 943 1168 945
rect 1171 942 1173 945
rect 1187 943 1189 945
rect 1203 943 1205 945
rect 1208 940 1210 945
rect 1229 940 1231 945
rect 1245 943 1247 945
rect 1261 943 1263 945
rect 1266 940 1268 945
rect 1282 943 1284 945
rect 1298 943 1300 945
rect 1303 942 1305 945
rect 1319 943 1321 945
rect 1335 943 1337 945
rect 1340 940 1342 945
rect 1361 940 1363 945
rect 1377 943 1379 945
rect 1393 943 1395 945
rect 1398 940 1400 945
rect 1414 943 1416 945
rect 333 905 335 908
rect 357 905 359 908
rect 1266 905 1268 908
rect 1290 905 1292 908
rect 333 899 335 901
rect 357 899 359 901
rect 1266 899 1268 901
rect 1290 899 1292 901
rect 353 894 355 896
rect 1286 894 1288 896
rect 353 887 355 890
rect 1286 887 1288 890
rect 342 876 344 878
rect 348 876 367 878
rect 1275 876 1277 878
rect 1281 876 1300 878
rect 333 871 335 873
rect 357 871 359 873
rect 1266 871 1268 873
rect 1290 871 1292 873
rect 333 864 335 867
rect 357 864 359 867
rect 1266 864 1268 867
rect 1290 864 1292 867
rect 101 836 103 838
rect 106 836 108 839
rect 122 836 124 838
rect 138 836 140 838
rect 143 836 145 839
rect 164 836 166 839
rect 180 836 182 839
rect 196 836 198 838
rect 201 836 203 839
rect 217 836 219 838
rect 233 836 235 838
rect 238 836 240 839
rect 254 836 256 838
rect 270 836 272 838
rect 275 836 277 839
rect 296 836 298 839
rect 312 836 314 839
rect 328 836 330 838
rect 333 836 335 839
rect 349 836 351 838
rect 365 836 367 838
rect 370 836 372 839
rect 386 836 388 838
rect 402 836 404 838
rect 407 836 409 839
rect 428 836 430 839
rect 444 836 446 839
rect 460 836 462 838
rect 465 836 467 839
rect 481 836 483 838
rect 1034 836 1036 838
rect 1039 836 1041 839
rect 1055 836 1057 838
rect 1071 836 1073 838
rect 1076 836 1078 839
rect 1097 836 1099 839
rect 1113 836 1115 839
rect 1129 836 1131 838
rect 1134 836 1136 839
rect 1150 836 1152 838
rect 1166 836 1168 838
rect 1171 836 1173 839
rect 1187 836 1189 838
rect 1203 836 1205 838
rect 1208 836 1210 839
rect 1229 836 1231 839
rect 1245 836 1247 839
rect 1261 836 1263 838
rect 1266 836 1268 839
rect 1282 836 1284 838
rect 1298 836 1300 838
rect 1303 836 1305 839
rect 1319 836 1321 838
rect 1335 836 1337 838
rect 1340 836 1342 839
rect 1361 836 1363 839
rect 1377 836 1379 839
rect 1393 836 1395 838
rect 1398 836 1400 839
rect 1414 836 1416 838
rect 101 823 103 828
rect 106 826 108 828
rect 101 809 103 819
rect 106 809 108 816
rect 122 809 124 828
rect 138 819 140 828
rect 143 826 145 828
rect 164 826 166 828
rect 180 825 182 828
rect 138 809 140 812
rect 143 809 145 811
rect 164 809 166 811
rect 180 809 182 821
rect 196 819 198 828
rect 201 826 203 828
rect 196 809 198 812
rect 201 809 203 811
rect 217 809 219 828
rect 233 825 235 828
rect 238 826 240 828
rect 233 809 235 821
rect 238 809 240 816
rect 254 809 256 828
rect 270 819 272 828
rect 275 826 277 828
rect 296 826 298 828
rect 312 825 314 828
rect 270 809 272 812
rect 275 809 277 811
rect 296 809 298 811
rect 312 809 314 821
rect 328 819 330 828
rect 333 826 335 828
rect 328 809 330 812
rect 333 809 335 811
rect 349 809 351 828
rect 365 825 367 828
rect 370 826 372 828
rect 365 809 367 821
rect 370 809 372 816
rect 386 809 388 828
rect 402 819 404 828
rect 407 826 409 828
rect 428 826 430 828
rect 444 825 446 828
rect 402 809 404 812
rect 407 809 409 811
rect 428 809 430 811
rect 444 809 446 821
rect 460 819 462 828
rect 465 826 467 828
rect 481 820 483 828
rect 1034 823 1036 828
rect 1039 826 1041 828
rect 460 809 462 812
rect 465 809 467 811
rect 481 809 483 816
rect 1034 809 1036 819
rect 1039 809 1041 816
rect 1055 809 1057 828
rect 1071 819 1073 828
rect 1076 826 1078 828
rect 1097 826 1099 828
rect 1113 825 1115 828
rect 1071 809 1073 812
rect 1076 809 1078 811
rect 1097 809 1099 811
rect 1113 809 1115 821
rect 1129 819 1131 828
rect 1134 826 1136 828
rect 1129 809 1131 812
rect 1134 809 1136 811
rect 1150 809 1152 828
rect 1166 825 1168 828
rect 1171 826 1173 828
rect 1166 809 1168 821
rect 1171 809 1173 816
rect 1187 809 1189 828
rect 1203 819 1205 828
rect 1208 826 1210 828
rect 1229 826 1231 828
rect 1245 825 1247 828
rect 1203 809 1205 812
rect 1208 809 1210 811
rect 1229 809 1231 811
rect 1245 809 1247 821
rect 1261 819 1263 828
rect 1266 826 1268 828
rect 1261 809 1263 812
rect 1266 809 1268 811
rect 1282 809 1284 828
rect 1298 825 1300 828
rect 1303 826 1305 828
rect 1298 809 1300 821
rect 1303 809 1305 816
rect 1319 809 1321 828
rect 1335 819 1337 828
rect 1340 826 1342 828
rect 1361 826 1363 828
rect 1377 825 1379 828
rect 1335 809 1337 812
rect 1340 809 1342 811
rect 1361 809 1363 811
rect 1377 809 1379 821
rect 1393 819 1395 828
rect 1398 826 1400 828
rect 1414 820 1416 828
rect 1393 809 1395 812
rect 1398 809 1400 811
rect 1414 809 1416 816
rect 101 803 103 805
rect 106 802 108 805
rect 122 803 124 805
rect 138 803 140 805
rect 143 800 145 805
rect 164 800 166 805
rect 180 803 182 805
rect 196 803 198 805
rect 201 800 203 805
rect 217 803 219 805
rect 233 803 235 805
rect 238 802 240 805
rect 254 803 256 805
rect 270 803 272 805
rect 275 800 277 805
rect 296 800 298 805
rect 312 803 314 805
rect 328 803 330 805
rect 333 800 335 805
rect 349 803 351 805
rect 365 803 367 805
rect 370 802 372 805
rect 386 803 388 805
rect 402 803 404 805
rect 407 800 409 805
rect 428 800 430 805
rect 444 803 446 805
rect 460 803 462 805
rect 465 800 467 805
rect 481 803 483 805
rect 1034 803 1036 805
rect 1039 802 1041 805
rect 1055 803 1057 805
rect 1071 803 1073 805
rect 1076 800 1078 805
rect 1097 800 1099 805
rect 1113 803 1115 805
rect 1129 803 1131 805
rect 1134 800 1136 805
rect 1150 803 1152 805
rect 1166 803 1168 805
rect 1171 802 1173 805
rect 1187 803 1189 805
rect 1203 803 1205 805
rect 1208 800 1210 805
rect 1229 800 1231 805
rect 1245 803 1247 805
rect 1261 803 1263 805
rect 1266 800 1268 805
rect 1282 803 1284 805
rect 1298 803 1300 805
rect 1303 802 1305 805
rect 1319 803 1321 805
rect 1335 803 1337 805
rect 1340 800 1342 805
rect 1361 800 1363 805
rect 1377 803 1379 805
rect 1393 803 1395 805
rect 1398 800 1400 805
rect 1414 803 1416 805
rect 573 757 575 759
rect 578 757 580 760
rect 594 757 596 759
rect 610 757 612 759
rect 615 757 617 760
rect 636 757 638 760
rect 652 757 654 760
rect 668 757 670 759
rect 673 757 675 760
rect 689 757 691 759
rect 705 757 707 759
rect 710 757 712 760
rect 726 757 728 759
rect 742 757 744 759
rect 747 757 749 760
rect 768 757 770 760
rect 784 757 786 760
rect 800 757 802 759
rect 805 757 807 760
rect 821 757 823 759
rect 837 757 839 759
rect 842 757 844 760
rect 858 757 860 759
rect 874 757 876 759
rect 879 757 881 760
rect 900 757 902 760
rect 916 757 918 760
rect 932 757 934 759
rect 937 757 939 760
rect 953 757 955 759
rect 969 757 971 759
rect 974 757 976 760
rect 990 757 992 759
rect 1006 757 1008 759
rect 1011 757 1013 760
rect 1032 757 1034 760
rect 1048 757 1050 760
rect 1064 757 1066 759
rect 1069 757 1071 760
rect 1085 757 1087 759
rect 1506 757 1508 759
rect 1511 757 1513 760
rect 1527 757 1529 759
rect 1543 757 1545 759
rect 1548 757 1550 760
rect 1569 757 1571 760
rect 1585 757 1587 760
rect 1601 757 1603 759
rect 1606 757 1608 760
rect 1622 757 1624 759
rect 1638 757 1640 759
rect 1643 757 1645 760
rect 1659 757 1661 759
rect 1675 757 1677 759
rect 1680 757 1682 760
rect 1701 757 1703 760
rect 1717 757 1719 760
rect 1733 757 1735 759
rect 1738 757 1740 760
rect 1754 757 1756 759
rect 1770 757 1772 759
rect 1775 757 1777 760
rect 1791 757 1793 759
rect 1807 757 1809 759
rect 1812 757 1814 760
rect 1833 757 1835 760
rect 1849 757 1851 760
rect 1865 757 1867 759
rect 1870 757 1872 760
rect 1886 757 1888 759
rect 1902 757 1904 759
rect 1907 757 1909 760
rect 1923 757 1925 759
rect 1939 757 1941 759
rect 1944 757 1946 760
rect 1965 757 1967 760
rect 1981 757 1983 760
rect 1997 757 1999 759
rect 2002 757 2004 760
rect 2018 757 2020 759
rect 573 744 575 749
rect 578 747 580 749
rect 573 730 575 740
rect 578 730 580 737
rect 594 730 596 749
rect 610 740 612 749
rect 615 747 617 749
rect 636 747 638 749
rect 652 746 654 749
rect 610 730 612 733
rect 615 730 617 732
rect 636 730 638 732
rect 652 730 654 742
rect 668 740 670 749
rect 673 747 675 749
rect 689 741 691 749
rect 705 744 707 749
rect 710 747 712 749
rect 668 730 670 733
rect 673 730 675 732
rect 689 730 691 737
rect 705 730 707 740
rect 710 730 712 737
rect 726 730 728 749
rect 742 740 744 749
rect 747 747 749 749
rect 768 747 770 749
rect 784 746 786 749
rect 742 730 744 733
rect 747 730 749 732
rect 768 730 770 732
rect 784 730 786 742
rect 800 740 802 749
rect 805 747 807 749
rect 821 741 823 749
rect 837 744 839 749
rect 842 747 844 749
rect 800 730 802 733
rect 805 730 807 732
rect 821 730 823 737
rect 837 730 839 740
rect 842 730 844 737
rect 858 730 860 749
rect 874 740 876 749
rect 879 747 881 749
rect 900 747 902 749
rect 916 746 918 749
rect 874 730 876 733
rect 879 730 881 732
rect 900 730 902 732
rect 916 730 918 742
rect 932 740 934 749
rect 937 747 939 749
rect 953 741 955 749
rect 969 744 971 749
rect 974 747 976 749
rect 932 730 934 733
rect 937 730 939 732
rect 953 730 955 737
rect 969 730 971 740
rect 974 730 976 737
rect 990 730 992 749
rect 1006 740 1008 749
rect 1011 747 1013 749
rect 1032 747 1034 749
rect 1048 746 1050 749
rect 1006 730 1008 733
rect 1011 730 1013 732
rect 1032 730 1034 732
rect 1048 730 1050 742
rect 1064 740 1066 749
rect 1069 747 1071 749
rect 1085 741 1087 749
rect 1506 744 1508 749
rect 1511 747 1513 749
rect 1064 730 1066 733
rect 1069 730 1071 732
rect 1085 730 1087 737
rect 233 724 235 726
rect 238 724 240 727
rect 254 724 256 726
rect 270 724 272 726
rect 275 724 277 727
rect 296 724 298 727
rect 312 724 314 727
rect 328 724 330 726
rect 333 724 335 727
rect 1506 730 1508 740
rect 1511 730 1513 737
rect 1527 730 1529 749
rect 1543 740 1545 749
rect 1548 747 1550 749
rect 1569 747 1571 749
rect 1585 746 1587 749
rect 1543 730 1545 733
rect 1548 730 1550 732
rect 1569 730 1571 732
rect 1585 730 1587 742
rect 1601 740 1603 749
rect 1606 747 1608 749
rect 1622 741 1624 749
rect 1638 744 1640 749
rect 1643 747 1645 749
rect 1601 730 1603 733
rect 1606 730 1608 732
rect 1622 730 1624 737
rect 1638 730 1640 740
rect 1643 730 1645 737
rect 1659 730 1661 749
rect 1675 740 1677 749
rect 1680 747 1682 749
rect 1701 747 1703 749
rect 1717 746 1719 749
rect 1675 730 1677 733
rect 1680 730 1682 732
rect 1701 730 1703 732
rect 1717 730 1719 742
rect 1733 740 1735 749
rect 1738 747 1740 749
rect 1754 741 1756 749
rect 1770 744 1772 749
rect 1775 747 1777 749
rect 1733 730 1735 733
rect 1738 730 1740 732
rect 1754 730 1756 737
rect 1770 730 1772 740
rect 1775 730 1777 737
rect 1791 730 1793 749
rect 1807 740 1809 749
rect 1812 747 1814 749
rect 1833 747 1835 749
rect 1849 746 1851 749
rect 1807 730 1809 733
rect 1812 730 1814 732
rect 1833 730 1835 732
rect 1849 730 1851 742
rect 1865 740 1867 749
rect 1870 747 1872 749
rect 1886 741 1888 749
rect 1902 744 1904 749
rect 1907 747 1909 749
rect 1865 730 1867 733
rect 1870 730 1872 732
rect 1886 730 1888 737
rect 1902 730 1904 740
rect 1907 730 1909 737
rect 1923 730 1925 749
rect 1939 740 1941 749
rect 1944 747 1946 749
rect 1965 747 1967 749
rect 1981 746 1983 749
rect 1939 730 1941 733
rect 1944 730 1946 732
rect 1965 730 1967 732
rect 1981 730 1983 742
rect 1997 740 1999 749
rect 2002 747 2004 749
rect 2018 741 2020 749
rect 1997 730 1999 733
rect 2002 730 2004 732
rect 2018 730 2020 737
rect 349 724 351 726
rect 573 724 575 726
rect 578 723 580 726
rect 594 724 596 726
rect 610 724 612 726
rect 615 721 617 726
rect 636 721 638 726
rect 652 724 654 726
rect 668 724 670 726
rect 673 721 675 726
rect 689 724 691 726
rect 705 724 707 726
rect 710 723 712 726
rect 726 724 728 726
rect 742 724 744 726
rect 747 721 749 726
rect 768 721 770 726
rect 784 724 786 726
rect 800 724 802 726
rect 805 721 807 726
rect 821 724 823 726
rect 837 724 839 726
rect 842 723 844 726
rect 858 724 860 726
rect 874 724 876 726
rect 879 721 881 726
rect 900 721 902 726
rect 916 724 918 726
rect 932 724 934 726
rect 937 721 939 726
rect 953 724 955 726
rect 969 724 971 726
rect 974 723 976 726
rect 990 724 992 726
rect 1006 724 1008 726
rect 1011 721 1013 726
rect 1032 721 1034 726
rect 1048 724 1050 726
rect 1064 724 1066 726
rect 1069 721 1071 726
rect 1085 724 1087 726
rect 1166 724 1168 726
rect 1171 724 1173 727
rect 1187 724 1189 726
rect 1203 724 1205 726
rect 1208 724 1210 727
rect 1229 724 1231 727
rect 1245 724 1247 727
rect 1261 724 1263 726
rect 1266 724 1268 727
rect 1282 724 1284 726
rect 1506 724 1508 726
rect 1511 723 1513 726
rect 1527 724 1529 726
rect 1543 724 1545 726
rect 1548 721 1550 726
rect 1569 721 1571 726
rect 1585 724 1587 726
rect 1601 724 1603 726
rect 1606 721 1608 726
rect 1622 724 1624 726
rect 1638 724 1640 726
rect 1643 723 1645 726
rect 1659 724 1661 726
rect 1675 724 1677 726
rect 1680 721 1682 726
rect 1701 721 1703 726
rect 1717 724 1719 726
rect 1733 724 1735 726
rect 1738 721 1740 726
rect 1754 724 1756 726
rect 1770 724 1772 726
rect 1775 723 1777 726
rect 1791 724 1793 726
rect 1807 724 1809 726
rect 1812 721 1814 726
rect 1833 721 1835 726
rect 1849 724 1851 726
rect 1865 724 1867 726
rect 1870 721 1872 726
rect 1886 724 1888 726
rect 1902 724 1904 726
rect 1907 723 1909 726
rect 1923 724 1925 726
rect 1939 724 1941 726
rect 1944 721 1946 726
rect 1965 721 1967 726
rect 1981 724 1983 726
rect 1997 724 1999 726
rect 2002 721 2004 726
rect 2018 724 2020 726
rect 233 711 235 716
rect 238 714 240 716
rect 233 697 235 707
rect 238 697 240 704
rect 254 697 256 716
rect 270 707 272 716
rect 275 714 277 716
rect 296 714 298 716
rect 312 713 314 716
rect 270 697 272 700
rect 275 697 277 699
rect 296 697 298 699
rect 312 697 314 709
rect 328 707 330 716
rect 333 714 335 716
rect 328 697 330 700
rect 333 697 335 699
rect 349 697 351 716
rect 1166 711 1168 716
rect 1171 714 1173 716
rect 1166 697 1168 707
rect 1171 697 1173 704
rect 1187 697 1189 716
rect 1203 707 1205 716
rect 1208 714 1210 716
rect 1229 714 1231 716
rect 1245 713 1247 716
rect 1203 697 1205 700
rect 1208 697 1210 699
rect 1229 697 1231 699
rect 1245 697 1247 709
rect 1261 707 1263 716
rect 1266 714 1268 716
rect 1261 697 1263 700
rect 1266 697 1268 699
rect 1282 697 1284 716
rect 233 691 235 693
rect 238 690 240 693
rect 254 691 256 693
rect 270 691 272 693
rect 275 688 277 693
rect 296 688 298 693
rect 312 691 314 693
rect 328 691 330 693
rect 333 688 335 693
rect 349 691 351 693
rect 1166 691 1168 693
rect 1171 690 1173 693
rect 1187 691 1189 693
rect 1203 691 1205 693
rect 752 686 754 688
rect 594 680 596 683
rect 638 680 640 683
rect 664 680 666 683
rect 710 680 712 683
rect 664 676 665 680
rect 778 680 780 684
rect 806 686 808 688
rect 833 686 835 688
rect 783 680 785 683
rect 578 673 580 675
rect 594 673 596 676
rect 610 673 612 675
rect 633 673 635 675
rect 638 673 640 676
rect 664 673 666 676
rect 685 673 687 676
rect 705 673 707 675
rect 710 673 712 676
rect 728 673 730 675
rect 357 660 359 663
rect 357 654 359 656
rect 240 651 242 654
rect 578 651 580 665
rect 594 663 596 665
rect 594 651 596 653
rect 610 651 612 665
rect 633 660 635 665
rect 638 663 640 665
rect 664 663 666 665
rect 629 656 635 660
rect 633 651 635 656
rect 638 651 640 653
rect 664 651 666 653
rect 685 651 687 665
rect 705 660 707 665
rect 710 663 712 665
rect 701 656 707 660
rect 705 651 707 656
rect 710 651 712 653
rect 728 651 730 665
rect 752 664 754 678
rect 859 680 861 684
rect 887 686 889 688
rect 1208 688 1210 693
rect 1229 688 1231 693
rect 1245 691 1247 693
rect 1261 691 1263 693
rect 1266 688 1268 693
rect 1282 691 1284 693
rect 864 680 866 683
rect 778 669 780 672
rect 783 670 785 672
rect 779 665 780 669
rect 778 660 780 665
rect 783 660 785 662
rect 752 658 754 660
rect 806 656 808 678
rect 833 664 835 678
rect 1685 686 1687 688
rect 859 669 861 672
rect 864 670 866 672
rect 860 665 861 669
rect 859 660 861 665
rect 864 660 866 662
rect 833 658 835 660
rect 887 656 889 678
rect 1527 680 1529 683
rect 1571 680 1573 683
rect 1597 680 1599 683
rect 1643 680 1645 683
rect 1597 676 1598 680
rect 1711 680 1713 684
rect 1739 686 1741 688
rect 1766 686 1768 688
rect 1716 680 1718 683
rect 1511 673 1513 675
rect 1527 673 1529 676
rect 1543 673 1545 675
rect 1566 673 1568 675
rect 1571 673 1573 676
rect 1597 673 1599 676
rect 1618 673 1620 676
rect 1638 673 1640 675
rect 1643 673 1645 676
rect 1661 673 1663 675
rect 1290 660 1292 663
rect 778 654 780 656
rect 783 651 785 656
rect 859 654 861 656
rect 806 650 808 652
rect 864 651 866 656
rect 1290 654 1292 656
rect 887 650 889 652
rect 1173 651 1175 654
rect 1511 651 1513 665
rect 1527 663 1529 665
rect 1527 651 1529 653
rect 1543 651 1545 665
rect 1566 660 1568 665
rect 1571 663 1573 665
rect 1597 663 1599 665
rect 1562 656 1568 660
rect 1566 651 1568 656
rect 1571 651 1573 653
rect 1597 651 1599 653
rect 1618 651 1620 665
rect 1638 660 1640 665
rect 1643 663 1645 665
rect 1634 656 1640 660
rect 1638 651 1640 656
rect 1643 651 1645 653
rect 1661 651 1663 665
rect 1685 664 1687 678
rect 1792 680 1794 684
rect 1820 686 1822 688
rect 1797 680 1799 683
rect 1711 669 1713 672
rect 1716 670 1718 672
rect 1712 665 1713 669
rect 1711 660 1713 665
rect 1716 660 1718 662
rect 1685 658 1687 660
rect 1739 656 1741 678
rect 1766 664 1768 678
rect 1792 669 1794 672
rect 1797 670 1799 672
rect 1793 665 1794 669
rect 1792 660 1794 665
rect 1797 660 1799 662
rect 1766 658 1768 660
rect 1820 656 1822 678
rect 1711 654 1713 656
rect 1716 651 1718 656
rect 1792 654 1794 656
rect 1739 650 1741 652
rect 1797 651 1799 656
rect 1820 650 1822 652
rect 240 645 242 647
rect 578 645 580 647
rect 594 643 596 647
rect 610 645 612 647
rect 633 645 635 647
rect 595 639 596 643
rect 638 642 640 647
rect 664 643 666 647
rect 685 645 687 647
rect 705 645 707 647
rect 594 636 596 639
rect 639 638 640 642
rect 665 639 666 643
rect 710 642 712 647
rect 728 645 730 647
rect 1173 645 1175 647
rect 1511 645 1513 647
rect 1527 643 1529 647
rect 1543 645 1545 647
rect 1566 645 1568 647
rect 638 636 640 638
rect 664 635 666 639
rect 711 638 712 642
rect 1528 639 1529 643
rect 1571 642 1573 647
rect 1597 643 1599 647
rect 1618 645 1620 647
rect 1638 645 1640 647
rect 710 636 712 638
rect 1527 636 1529 639
rect 1572 638 1573 642
rect 1598 639 1599 643
rect 1643 642 1645 647
rect 1661 645 1663 647
rect 1571 636 1573 638
rect 1597 635 1599 639
rect 1644 638 1645 642
rect 1643 636 1645 638
rect 224 622 226 624
rect 240 622 242 625
rect 245 622 247 624
rect 261 622 263 625
rect 277 622 279 625
rect 298 622 300 625
rect 303 622 305 624
rect 319 622 321 624
rect 335 622 337 625
rect 340 622 342 624
rect 1157 622 1159 624
rect 1173 622 1175 625
rect 1178 622 1180 624
rect 1194 622 1196 625
rect 1210 622 1212 625
rect 1231 622 1233 625
rect 1236 622 1238 624
rect 1252 622 1254 624
rect 1268 622 1270 625
rect 1273 622 1275 624
rect 224 595 226 614
rect 240 612 242 614
rect 245 605 247 614
rect 261 611 263 614
rect 277 612 279 614
rect 298 612 300 614
rect 240 595 242 597
rect 245 595 247 598
rect 261 595 263 607
rect 303 605 305 614
rect 277 595 279 597
rect 298 595 300 597
rect 303 595 305 598
rect 319 595 321 614
rect 335 612 337 614
rect 340 609 342 614
rect 594 613 596 616
rect 638 614 640 616
rect 595 609 596 613
rect 639 610 640 614
rect 664 613 666 617
rect 710 614 712 616
rect 578 605 580 607
rect 594 605 596 609
rect 610 605 612 607
rect 633 605 635 607
rect 638 605 640 610
rect 665 609 666 613
rect 711 610 712 614
rect 664 605 666 609
rect 685 605 687 607
rect 705 605 707 607
rect 710 605 712 610
rect 728 605 730 607
rect 335 595 337 602
rect 340 595 342 605
rect 778 604 780 607
rect 783 604 785 607
rect 859 604 861 607
rect 864 604 866 607
rect 224 589 226 591
rect 240 586 242 591
rect 245 589 247 591
rect 261 589 263 591
rect 277 586 279 591
rect 298 586 300 591
rect 303 589 305 591
rect 319 589 321 591
rect 335 588 337 591
rect 340 589 342 591
rect 578 587 580 601
rect 594 599 596 601
rect 594 587 596 589
rect 610 587 612 601
rect 633 596 635 601
rect 638 599 640 601
rect 664 599 666 601
rect 629 592 635 596
rect 633 587 635 592
rect 638 587 640 589
rect 664 587 666 589
rect 685 587 687 601
rect 705 596 707 601
rect 710 599 712 601
rect 701 592 707 596
rect 705 587 707 592
rect 710 587 712 589
rect 728 587 730 601
rect 778 588 780 600
rect 783 598 785 600
rect 783 588 785 590
rect 859 588 861 600
rect 864 598 866 600
rect 1157 595 1159 614
rect 1173 612 1175 614
rect 1178 605 1180 614
rect 1194 611 1196 614
rect 1210 612 1212 614
rect 1231 612 1233 614
rect 1173 595 1175 597
rect 1178 595 1180 598
rect 1194 595 1196 607
rect 1236 605 1238 614
rect 1210 595 1212 597
rect 1231 595 1233 597
rect 1236 595 1238 598
rect 1252 595 1254 614
rect 1268 612 1270 614
rect 1273 609 1275 614
rect 1527 613 1529 616
rect 1571 614 1573 616
rect 1528 609 1529 613
rect 1572 610 1573 614
rect 1597 613 1599 617
rect 1643 614 1645 616
rect 1511 605 1513 607
rect 1527 605 1529 609
rect 1543 605 1545 607
rect 1566 605 1568 607
rect 1571 605 1573 610
rect 1598 609 1599 613
rect 1644 610 1645 614
rect 1597 605 1599 609
rect 1618 605 1620 607
rect 1638 605 1640 607
rect 1643 605 1645 610
rect 1661 605 1663 607
rect 1268 595 1270 602
rect 1273 595 1275 605
rect 1711 604 1713 607
rect 1716 604 1718 607
rect 1792 604 1794 607
rect 1797 604 1799 607
rect 864 588 866 590
rect 1157 589 1159 591
rect 1173 586 1175 591
rect 1178 589 1180 591
rect 1194 589 1196 591
rect 1210 586 1212 591
rect 1231 586 1233 591
rect 1236 589 1238 591
rect 1252 589 1254 591
rect 1268 588 1270 591
rect 1273 589 1275 591
rect 1511 587 1513 601
rect 1527 599 1529 601
rect 1527 587 1529 589
rect 1543 587 1545 601
rect 1566 596 1568 601
rect 1571 599 1573 601
rect 1597 599 1599 601
rect 1562 592 1568 596
rect 1566 587 1568 592
rect 1571 587 1573 589
rect 1597 587 1599 589
rect 1618 587 1620 601
rect 1638 596 1640 601
rect 1643 599 1645 601
rect 1634 592 1640 596
rect 1638 587 1640 592
rect 1643 587 1645 589
rect 1661 587 1663 601
rect 1711 588 1713 600
rect 1716 598 1718 600
rect 1716 588 1718 590
rect 1792 588 1794 600
rect 1797 598 1799 600
rect 1797 588 1799 590
rect 578 577 580 579
rect 594 576 596 579
rect 610 577 612 579
rect 633 577 635 579
rect 638 576 640 579
rect 664 576 666 579
rect 685 576 687 579
rect 705 577 707 579
rect 710 576 712 579
rect 728 577 730 579
rect 778 578 780 580
rect 664 572 665 576
rect 783 575 785 580
rect 859 578 861 580
rect 864 575 866 580
rect 1511 577 1513 579
rect 1527 576 1529 579
rect 1543 577 1545 579
rect 1566 577 1568 579
rect 1571 576 1573 579
rect 1597 576 1599 579
rect 1618 576 1620 579
rect 1638 577 1640 579
rect 1643 576 1645 579
rect 1661 577 1663 579
rect 1711 578 1713 580
rect 594 569 596 572
rect 638 569 640 572
rect 664 569 666 572
rect 710 569 712 572
rect 1597 572 1598 576
rect 1716 575 1718 580
rect 1792 578 1794 580
rect 1797 575 1799 580
rect 1527 569 1529 572
rect 1571 569 1573 572
rect 1597 569 1599 572
rect 1643 569 1645 572
rect 594 548 596 551
rect 638 548 640 551
rect 664 548 666 551
rect 710 548 712 551
rect 778 548 780 552
rect 806 554 808 556
rect 857 554 859 556
rect 783 548 785 551
rect 664 544 665 548
rect 578 541 580 543
rect 594 541 596 544
rect 610 541 612 543
rect 633 541 635 543
rect 638 541 640 544
rect 664 541 666 544
rect 685 541 687 544
rect 705 541 707 543
rect 710 541 712 544
rect 728 541 730 543
rect 883 548 885 552
rect 911 554 913 556
rect 888 548 890 551
rect 778 537 780 540
rect 783 538 785 540
rect 779 533 780 537
rect 578 519 580 533
rect 594 531 596 533
rect 594 519 596 521
rect 610 519 612 533
rect 633 528 635 533
rect 638 531 640 533
rect 664 531 666 533
rect 629 524 635 528
rect 633 519 635 524
rect 638 519 640 521
rect 664 519 666 521
rect 685 519 687 533
rect 705 528 707 533
rect 710 531 712 533
rect 701 524 707 528
rect 705 519 707 524
rect 710 519 712 521
rect 728 519 730 533
rect 778 528 780 533
rect 783 528 785 530
rect 806 524 808 546
rect 857 532 859 546
rect 1527 548 1529 551
rect 1571 548 1573 551
rect 1597 548 1599 551
rect 1643 548 1645 551
rect 1711 548 1713 552
rect 1739 554 1741 556
rect 1790 554 1792 556
rect 1716 548 1718 551
rect 883 537 885 540
rect 888 538 890 540
rect 884 533 885 537
rect 883 528 885 533
rect 888 528 890 530
rect 857 526 859 528
rect 911 524 913 546
rect 1597 544 1598 548
rect 1511 541 1513 543
rect 1527 541 1529 544
rect 1543 541 1545 543
rect 1566 541 1568 543
rect 1571 541 1573 544
rect 1597 541 1599 544
rect 1618 541 1620 544
rect 1638 541 1640 543
rect 1643 541 1645 544
rect 1661 541 1663 543
rect 1816 548 1818 552
rect 1844 554 1846 556
rect 1821 548 1823 551
rect 1711 537 1713 540
rect 1716 538 1718 540
rect 1712 533 1713 537
rect 778 522 780 524
rect 783 519 785 524
rect 883 522 885 524
rect 806 518 808 520
rect 888 519 890 524
rect 911 518 913 520
rect 1511 519 1513 533
rect 1527 531 1529 533
rect 1527 519 1529 521
rect 1543 519 1545 533
rect 1566 528 1568 533
rect 1571 531 1573 533
rect 1597 531 1599 533
rect 1562 524 1568 528
rect 1566 519 1568 524
rect 1571 519 1573 521
rect 1597 519 1599 521
rect 1618 519 1620 533
rect 1638 528 1640 533
rect 1643 531 1645 533
rect 1634 524 1640 528
rect 1638 519 1640 524
rect 1643 519 1645 521
rect 1661 519 1663 533
rect 1711 528 1713 533
rect 1716 528 1718 530
rect 1739 524 1741 546
rect 1790 532 1792 546
rect 1816 537 1818 540
rect 1821 538 1823 540
rect 1817 533 1818 537
rect 1816 528 1818 533
rect 1821 528 1823 530
rect 1790 526 1792 528
rect 1844 524 1846 546
rect 1711 522 1713 524
rect 1716 519 1718 524
rect 1816 522 1818 524
rect 1739 518 1741 520
rect 1821 519 1823 524
rect 1844 518 1846 520
rect 578 513 580 515
rect 594 511 596 515
rect 610 513 612 515
rect 633 513 635 515
rect 595 507 596 511
rect 638 510 640 515
rect 664 511 666 515
rect 685 513 687 515
rect 705 513 707 515
rect 594 504 596 507
rect 639 506 640 510
rect 665 507 666 511
rect 710 510 712 515
rect 728 513 730 515
rect 1511 513 1513 515
rect 1527 511 1529 515
rect 1543 513 1545 515
rect 1566 513 1568 515
rect 638 504 640 506
rect 664 503 666 507
rect 711 506 712 510
rect 1528 507 1529 511
rect 1571 510 1573 515
rect 1597 511 1599 515
rect 1618 513 1620 515
rect 1638 513 1640 515
rect 710 504 712 506
rect 1527 504 1529 507
rect 1572 506 1573 510
rect 1598 507 1599 511
rect 1643 510 1645 515
rect 1661 513 1663 515
rect 1571 504 1573 506
rect 1597 503 1599 507
rect 1644 506 1645 510
rect 1643 504 1645 506
rect 594 481 596 484
rect 638 482 640 484
rect 595 477 596 481
rect 639 478 640 482
rect 664 481 666 485
rect 710 482 712 484
rect 578 473 580 475
rect 594 473 596 477
rect 610 473 612 475
rect 633 473 635 475
rect 638 473 640 478
rect 665 477 666 481
rect 711 478 712 482
rect 1527 481 1529 484
rect 1571 482 1573 484
rect 664 473 666 477
rect 685 473 687 475
rect 705 473 707 475
rect 710 473 712 478
rect 1528 477 1529 481
rect 1572 478 1573 482
rect 1597 481 1599 485
rect 1643 482 1645 484
rect 728 473 730 475
rect 778 473 780 476
rect 783 473 785 476
rect 883 473 885 476
rect 888 473 890 476
rect 1511 473 1513 475
rect 1527 473 1529 477
rect 1543 473 1545 475
rect 1566 473 1568 475
rect 1571 473 1573 478
rect 1598 477 1599 481
rect 1644 478 1645 482
rect 1597 473 1599 477
rect 1618 473 1620 475
rect 1638 473 1640 475
rect 1643 473 1645 478
rect 1661 473 1663 475
rect 1711 473 1713 476
rect 1716 473 1718 476
rect 1816 473 1818 476
rect 1821 473 1823 476
rect 578 455 580 469
rect 594 467 596 469
rect 594 455 596 457
rect 610 455 612 469
rect 633 464 635 469
rect 638 467 640 469
rect 664 467 666 469
rect 629 460 635 464
rect 633 455 635 460
rect 638 455 640 457
rect 664 455 666 457
rect 685 455 687 469
rect 705 464 707 469
rect 710 467 712 469
rect 701 460 707 464
rect 705 455 707 460
rect 710 455 712 457
rect 728 455 730 469
rect 778 457 780 469
rect 783 467 785 469
rect 783 457 785 459
rect 883 457 885 469
rect 888 467 890 469
rect 888 457 890 459
rect 1511 455 1513 469
rect 1527 467 1529 469
rect 1527 455 1529 457
rect 1543 455 1545 469
rect 1566 464 1568 469
rect 1571 467 1573 469
rect 1597 467 1599 469
rect 1562 460 1568 464
rect 1566 455 1568 460
rect 1571 455 1573 457
rect 1597 455 1599 457
rect 1618 455 1620 469
rect 1638 464 1640 469
rect 1643 467 1645 469
rect 1634 460 1640 464
rect 1638 455 1640 460
rect 1643 455 1645 457
rect 1661 455 1663 469
rect 1711 457 1713 469
rect 1716 467 1718 469
rect 1716 457 1718 459
rect 1816 457 1818 469
rect 1821 467 1823 469
rect 1821 457 1823 459
rect 778 447 780 449
rect 578 445 580 447
rect 594 444 596 447
rect 610 445 612 447
rect 633 445 635 447
rect 638 444 640 447
rect 664 444 666 447
rect 685 444 687 447
rect 705 445 707 447
rect 710 444 712 447
rect 728 445 730 447
rect 783 444 785 449
rect 883 447 885 449
rect 888 444 890 449
rect 1711 447 1713 449
rect 1511 445 1513 447
rect 664 440 665 444
rect 1527 444 1529 447
rect 1543 445 1545 447
rect 1566 445 1568 447
rect 1571 444 1573 447
rect 1597 444 1599 447
rect 1618 444 1620 447
rect 1638 445 1640 447
rect 1643 444 1645 447
rect 1661 445 1663 447
rect 1716 444 1718 449
rect 1816 447 1818 449
rect 1821 444 1823 449
rect 1597 440 1598 444
rect 594 437 596 440
rect 638 437 640 440
rect 664 437 666 440
rect 710 437 712 440
rect 1527 437 1529 440
rect 1571 437 1573 440
rect 1597 437 1599 440
rect 1643 437 1645 440
rect 594 416 596 419
rect 638 416 640 419
rect 664 416 666 419
rect 710 416 712 419
rect 778 416 780 420
rect 806 422 808 424
rect 833 422 835 424
rect 783 416 785 419
rect 664 412 665 416
rect 578 409 580 411
rect 594 409 596 412
rect 610 409 612 411
rect 633 409 635 411
rect 638 409 640 412
rect 664 409 666 412
rect 685 409 687 412
rect 705 409 707 411
rect 710 409 712 412
rect 728 409 730 411
rect 859 416 861 420
rect 887 422 889 424
rect 923 422 925 424
rect 864 416 866 419
rect 778 405 780 408
rect 783 406 785 408
rect 779 401 780 405
rect 578 387 580 401
rect 594 399 596 401
rect 594 387 596 389
rect 610 387 612 401
rect 633 396 635 401
rect 638 399 640 401
rect 664 399 666 401
rect 629 392 635 396
rect 633 387 635 392
rect 638 387 640 389
rect 664 387 666 389
rect 685 387 687 401
rect 705 396 707 401
rect 710 399 712 401
rect 701 392 707 396
rect 705 387 707 392
rect 710 387 712 389
rect 728 387 730 401
rect 778 396 780 401
rect 783 396 785 398
rect 806 392 808 414
rect 833 400 835 414
rect 949 416 951 420
rect 977 422 979 424
rect 954 416 956 419
rect 859 405 861 408
rect 864 406 866 408
rect 860 401 861 405
rect 859 396 861 401
rect 864 396 866 398
rect 833 394 835 396
rect 887 392 889 414
rect 923 400 925 414
rect 1527 416 1529 419
rect 1571 416 1573 419
rect 1597 416 1599 419
rect 1643 416 1645 419
rect 1711 416 1713 420
rect 1739 422 1741 424
rect 1766 422 1768 424
rect 1716 416 1718 419
rect 949 405 951 408
rect 954 406 956 408
rect 950 401 951 405
rect 949 396 951 401
rect 954 396 956 398
rect 923 394 925 396
rect 977 392 979 414
rect 1597 412 1598 416
rect 1511 409 1513 411
rect 1527 409 1529 412
rect 1543 409 1545 411
rect 1566 409 1568 411
rect 1571 409 1573 412
rect 1597 409 1599 412
rect 1618 409 1620 412
rect 1638 409 1640 411
rect 1643 409 1645 412
rect 1661 409 1663 411
rect 1792 416 1794 420
rect 1820 422 1822 424
rect 1856 422 1858 424
rect 1797 416 1799 419
rect 1711 405 1713 408
rect 1716 406 1718 408
rect 1712 401 1713 405
rect 778 390 780 392
rect 783 387 785 392
rect 859 390 861 392
rect 806 386 808 388
rect 864 387 866 392
rect 949 390 951 392
rect 887 386 889 388
rect 954 387 956 392
rect 977 386 979 388
rect 1511 387 1513 401
rect 1527 399 1529 401
rect 1527 387 1529 389
rect 1543 387 1545 401
rect 1566 396 1568 401
rect 1571 399 1573 401
rect 1597 399 1599 401
rect 1562 392 1568 396
rect 1566 387 1568 392
rect 1571 387 1573 389
rect 1597 387 1599 389
rect 1618 387 1620 401
rect 1638 396 1640 401
rect 1643 399 1645 401
rect 1634 392 1640 396
rect 1638 387 1640 392
rect 1643 387 1645 389
rect 1661 387 1663 401
rect 1711 396 1713 401
rect 1716 396 1718 398
rect 1739 392 1741 414
rect 1766 400 1768 414
rect 1882 416 1884 420
rect 1910 422 1912 424
rect 1887 416 1889 419
rect 1792 405 1794 408
rect 1797 406 1799 408
rect 1793 401 1794 405
rect 1792 396 1794 401
rect 1797 396 1799 398
rect 1766 394 1768 396
rect 1820 392 1822 414
rect 1856 400 1858 414
rect 1882 405 1884 408
rect 1887 406 1889 408
rect 1883 401 1884 405
rect 1882 396 1884 401
rect 1887 396 1889 398
rect 1856 394 1858 396
rect 1910 392 1912 414
rect 1711 390 1713 392
rect 1716 387 1718 392
rect 1792 390 1794 392
rect 1739 386 1741 388
rect 1797 387 1799 392
rect 1882 390 1884 392
rect 1820 386 1822 388
rect 1887 387 1889 392
rect 1910 386 1912 388
rect 578 381 580 383
rect 594 379 596 383
rect 610 381 612 383
rect 633 381 635 383
rect 595 375 596 379
rect 638 378 640 383
rect 664 379 666 383
rect 685 381 687 383
rect 705 381 707 383
rect 594 372 596 375
rect 639 374 640 378
rect 665 375 666 379
rect 710 378 712 383
rect 728 381 730 383
rect 1511 381 1513 383
rect 1527 379 1529 383
rect 1543 381 1545 383
rect 1566 381 1568 383
rect 638 372 640 374
rect 664 371 666 375
rect 711 374 712 378
rect 1528 375 1529 379
rect 1571 378 1573 383
rect 1597 379 1599 383
rect 1618 381 1620 383
rect 1638 381 1640 383
rect 710 372 712 374
rect 1527 372 1529 375
rect 1572 374 1573 378
rect 1598 375 1599 379
rect 1643 378 1645 383
rect 1661 381 1663 383
rect 1571 372 1573 374
rect 1597 371 1599 375
rect 1644 374 1645 378
rect 1643 372 1645 374
rect 594 349 596 352
rect 638 350 640 352
rect 595 345 596 349
rect 639 346 640 350
rect 664 349 666 353
rect 710 350 712 352
rect 578 341 580 343
rect 594 341 596 345
rect 610 341 612 343
rect 633 341 635 343
rect 638 341 640 346
rect 665 345 666 349
rect 711 346 712 350
rect 1527 349 1529 352
rect 1571 350 1573 352
rect 664 341 666 345
rect 685 341 687 343
rect 705 341 707 343
rect 710 341 712 346
rect 1528 345 1529 349
rect 1572 346 1573 350
rect 1597 349 1599 353
rect 1643 350 1645 352
rect 728 341 730 343
rect 1511 341 1513 343
rect 1527 341 1529 345
rect 1543 341 1545 343
rect 1566 341 1568 343
rect 1571 341 1573 346
rect 1598 345 1599 349
rect 1644 346 1645 350
rect 1597 341 1599 345
rect 1618 341 1620 343
rect 1638 341 1640 343
rect 1643 341 1645 346
rect 1661 341 1663 343
rect 778 338 780 341
rect 783 338 785 341
rect 859 338 861 341
rect 864 338 866 341
rect 949 338 951 341
rect 954 338 956 341
rect 578 323 580 337
rect 594 335 596 337
rect 594 323 596 325
rect 610 323 612 337
rect 633 332 635 337
rect 638 335 640 337
rect 664 335 666 337
rect 629 328 635 332
rect 633 323 635 328
rect 638 323 640 325
rect 664 323 666 325
rect 685 323 687 337
rect 705 332 707 337
rect 710 335 712 337
rect 701 328 707 332
rect 705 323 707 328
rect 710 323 712 325
rect 728 323 730 337
rect 1711 338 1713 341
rect 1716 338 1718 341
rect 1792 338 1794 341
rect 1797 338 1799 341
rect 1882 338 1884 341
rect 1887 338 1889 341
rect 778 322 780 334
rect 783 332 785 334
rect 783 322 785 324
rect 859 322 861 334
rect 864 332 866 334
rect 864 322 866 324
rect 949 322 951 334
rect 954 332 956 334
rect 954 322 956 324
rect 1511 323 1513 337
rect 1527 335 1529 337
rect 1527 323 1529 325
rect 1543 323 1545 337
rect 1566 332 1568 337
rect 1571 335 1573 337
rect 1597 335 1599 337
rect 1562 328 1568 332
rect 1566 323 1568 328
rect 1571 323 1573 325
rect 1597 323 1599 325
rect 1618 323 1620 337
rect 1638 332 1640 337
rect 1643 335 1645 337
rect 1634 328 1640 332
rect 1638 323 1640 328
rect 1643 323 1645 325
rect 1661 323 1663 337
rect 578 313 580 315
rect 594 312 596 315
rect 610 313 612 315
rect 633 313 635 315
rect 638 312 640 315
rect 664 312 666 315
rect 685 312 687 315
rect 705 313 707 315
rect 710 312 712 315
rect 728 313 730 315
rect 1711 322 1713 334
rect 1716 332 1718 334
rect 1716 322 1718 324
rect 1792 322 1794 334
rect 1797 332 1799 334
rect 1797 322 1799 324
rect 1882 322 1884 334
rect 1887 332 1889 334
rect 1887 322 1889 324
rect 778 312 780 314
rect 664 308 665 312
rect 783 309 785 314
rect 859 312 861 314
rect 864 309 866 314
rect 949 312 951 314
rect 954 309 956 314
rect 1511 313 1513 315
rect 594 305 596 308
rect 638 305 640 308
rect 664 305 666 308
rect 710 305 712 308
rect 1527 312 1529 315
rect 1543 313 1545 315
rect 1566 313 1568 315
rect 1571 312 1573 315
rect 1597 312 1599 315
rect 1618 312 1620 315
rect 1638 313 1640 315
rect 1643 312 1645 315
rect 1661 313 1663 315
rect 1711 312 1713 314
rect 1597 308 1598 312
rect 1716 309 1718 314
rect 1792 312 1794 314
rect 1797 309 1799 314
rect 1882 312 1884 314
rect 1887 309 1889 314
rect 1527 305 1529 308
rect 1571 305 1573 308
rect 1597 305 1599 308
rect 1643 305 1645 308
rect 594 284 596 287
rect 638 284 640 287
rect 664 284 666 287
rect 710 284 712 287
rect 778 284 780 288
rect 806 290 808 292
rect 783 284 785 287
rect 664 280 665 284
rect 578 277 580 279
rect 594 277 596 280
rect 610 277 612 279
rect 633 277 635 279
rect 638 277 640 280
rect 664 277 666 280
rect 685 277 687 280
rect 705 277 707 279
rect 710 277 712 280
rect 728 277 730 279
rect 1527 284 1529 287
rect 1571 284 1573 287
rect 1597 284 1599 287
rect 1643 284 1645 287
rect 1711 284 1713 288
rect 1739 290 1741 292
rect 1716 284 1718 287
rect 778 273 780 276
rect 783 274 785 276
rect 779 269 780 273
rect 578 255 580 269
rect 594 267 596 269
rect 594 255 596 257
rect 610 255 612 269
rect 633 264 635 269
rect 638 267 640 269
rect 664 267 666 269
rect 629 260 635 264
rect 633 255 635 260
rect 638 255 640 257
rect 664 255 666 257
rect 685 255 687 269
rect 705 264 707 269
rect 710 267 712 269
rect 701 260 707 264
rect 705 255 707 260
rect 710 255 712 257
rect 728 255 730 269
rect 778 264 780 269
rect 783 264 785 266
rect 806 260 808 282
rect 1597 280 1598 284
rect 1511 277 1513 279
rect 1527 277 1529 280
rect 1543 277 1545 279
rect 1566 277 1568 279
rect 1571 277 1573 280
rect 1597 277 1599 280
rect 1618 277 1620 280
rect 1638 277 1640 279
rect 1643 277 1645 280
rect 1661 277 1663 279
rect 1711 273 1713 276
rect 1716 274 1718 276
rect 1712 269 1713 273
rect 778 258 780 260
rect 783 255 785 260
rect 806 254 808 256
rect 1511 255 1513 269
rect 1527 267 1529 269
rect 1527 255 1529 257
rect 1543 255 1545 269
rect 1566 264 1568 269
rect 1571 267 1573 269
rect 1597 267 1599 269
rect 1562 260 1568 264
rect 1566 255 1568 260
rect 1571 255 1573 257
rect 1597 255 1599 257
rect 1618 255 1620 269
rect 1638 264 1640 269
rect 1643 267 1645 269
rect 1634 260 1640 264
rect 1638 255 1640 260
rect 1643 255 1645 257
rect 1661 255 1663 269
rect 1711 264 1713 269
rect 1716 264 1718 266
rect 1739 260 1741 282
rect 1711 258 1713 260
rect 1716 255 1718 260
rect 1739 254 1741 256
rect 578 249 580 251
rect 594 247 596 251
rect 610 249 612 251
rect 633 249 635 251
rect 595 243 596 247
rect 638 246 640 251
rect 664 247 666 251
rect 685 249 687 251
rect 705 249 707 251
rect 594 240 596 243
rect 639 242 640 246
rect 665 243 666 247
rect 710 246 712 251
rect 728 249 730 251
rect 1511 249 1513 251
rect 1527 247 1529 251
rect 1543 249 1545 251
rect 1566 249 1568 251
rect 638 240 640 242
rect 664 239 666 243
rect 711 242 712 246
rect 1528 243 1529 247
rect 1571 246 1573 251
rect 1597 247 1599 251
rect 1618 249 1620 251
rect 1638 249 1640 251
rect 710 240 712 242
rect 1527 240 1529 243
rect 1572 242 1573 246
rect 1598 243 1599 247
rect 1643 246 1645 251
rect 1661 249 1663 251
rect 1571 240 1573 242
rect 1597 239 1599 243
rect 1644 242 1645 246
rect 1643 240 1645 242
rect 101 222 103 224
rect 106 222 108 225
rect 122 222 124 224
rect 138 222 140 224
rect 143 222 145 225
rect 164 222 166 225
rect 180 222 182 225
rect 196 222 198 224
rect 201 222 203 225
rect 217 222 219 224
rect 233 222 235 224
rect 238 222 240 225
rect 254 222 256 224
rect 270 222 272 224
rect 275 222 277 225
rect 296 222 298 225
rect 312 222 314 225
rect 328 222 330 224
rect 333 222 335 225
rect 349 222 351 224
rect 365 222 367 224
rect 370 222 372 225
rect 386 222 388 224
rect 402 222 404 224
rect 407 222 409 225
rect 428 222 430 225
rect 444 222 446 225
rect 460 222 462 224
rect 465 222 467 225
rect 481 222 483 224
rect 1034 222 1036 224
rect 1039 222 1041 225
rect 1055 222 1057 224
rect 1071 222 1073 224
rect 1076 222 1078 225
rect 1097 222 1099 225
rect 1113 222 1115 225
rect 1129 222 1131 224
rect 1134 222 1136 225
rect 1150 222 1152 224
rect 1166 222 1168 224
rect 1171 222 1173 225
rect 1187 222 1189 224
rect 1203 222 1205 224
rect 1208 222 1210 225
rect 1229 222 1231 225
rect 1245 222 1247 225
rect 1261 222 1263 224
rect 1266 222 1268 225
rect 1282 222 1284 224
rect 1298 222 1300 224
rect 1303 222 1305 225
rect 1319 222 1321 224
rect 1335 222 1337 224
rect 1340 222 1342 225
rect 1361 222 1363 225
rect 1377 222 1379 225
rect 1393 222 1395 224
rect 1398 222 1400 225
rect 1414 222 1416 224
rect 594 217 596 220
rect 638 218 640 220
rect 101 209 103 214
rect 106 212 108 214
rect 101 195 103 205
rect 106 195 108 202
rect 122 195 124 214
rect 138 205 140 214
rect 143 212 145 214
rect 164 212 166 214
rect 180 211 182 214
rect 138 195 140 198
rect 143 195 145 197
rect 164 195 166 197
rect 180 195 182 207
rect 196 205 198 214
rect 201 212 203 214
rect 196 195 198 198
rect 201 195 203 197
rect 217 195 219 214
rect 233 211 235 214
rect 238 212 240 214
rect 233 195 235 207
rect 238 195 240 202
rect 254 195 256 214
rect 270 205 272 214
rect 275 212 277 214
rect 296 212 298 214
rect 312 211 314 214
rect 270 195 272 198
rect 275 195 277 197
rect 296 195 298 197
rect 312 195 314 207
rect 328 205 330 214
rect 333 212 335 214
rect 328 195 330 198
rect 333 195 335 197
rect 349 195 351 214
rect 365 211 367 214
rect 370 212 372 214
rect 365 195 367 207
rect 370 195 372 202
rect 386 195 388 214
rect 402 205 404 214
rect 407 212 409 214
rect 428 212 430 214
rect 444 211 446 214
rect 402 195 404 198
rect 407 195 409 197
rect 428 195 430 197
rect 444 195 446 207
rect 460 205 462 214
rect 465 212 467 214
rect 481 206 483 214
rect 595 213 596 217
rect 639 214 640 218
rect 664 217 666 221
rect 710 218 712 220
rect 578 209 580 211
rect 594 209 596 213
rect 610 209 612 211
rect 633 209 635 211
rect 638 209 640 214
rect 665 213 666 217
rect 711 214 712 218
rect 855 217 857 220
rect 899 218 901 220
rect 664 209 666 213
rect 685 209 687 211
rect 705 209 707 211
rect 710 209 712 214
rect 856 213 857 217
rect 900 214 901 218
rect 925 217 927 221
rect 971 218 973 220
rect 728 209 730 211
rect 812 209 814 212
rect 830 209 832 212
rect 855 209 857 213
rect 871 209 873 211
rect 894 209 896 211
rect 899 209 901 214
rect 926 213 927 217
rect 972 214 973 218
rect 1527 217 1529 220
rect 1571 218 1573 220
rect 925 209 927 213
rect 946 209 948 211
rect 966 209 968 211
rect 971 209 973 214
rect 989 209 991 211
rect 1034 209 1036 214
rect 1039 212 1041 214
rect 460 195 462 198
rect 465 195 467 197
rect 481 195 483 202
rect 578 191 580 205
rect 594 203 596 205
rect 594 191 596 193
rect 610 191 612 205
rect 633 200 635 205
rect 638 203 640 205
rect 664 203 666 205
rect 629 196 635 200
rect 633 191 635 196
rect 638 191 640 193
rect 664 191 666 193
rect 685 191 687 205
rect 705 200 707 205
rect 710 203 712 205
rect 701 196 707 200
rect 705 191 707 196
rect 710 191 712 193
rect 728 191 730 205
rect 778 202 780 205
rect 783 202 785 205
rect 812 200 814 205
rect 101 189 103 191
rect 106 188 108 191
rect 122 189 124 191
rect 138 189 140 191
rect 143 186 145 191
rect 164 186 166 191
rect 180 189 182 191
rect 196 189 198 191
rect 201 186 203 191
rect 217 189 219 191
rect 233 189 235 191
rect 238 188 240 191
rect 254 189 256 191
rect 270 189 272 191
rect 275 186 277 191
rect 296 186 298 191
rect 312 189 314 191
rect 328 189 330 191
rect 333 186 335 191
rect 349 189 351 191
rect 365 189 367 191
rect 370 188 372 191
rect 386 189 388 191
rect 402 189 404 191
rect 407 186 409 191
rect 428 186 430 191
rect 444 189 446 191
rect 460 189 462 191
rect 465 186 467 191
rect 481 189 483 191
rect 778 186 780 198
rect 783 196 785 198
rect 812 191 814 196
rect 830 191 832 205
rect 855 203 857 205
rect 855 191 857 193
rect 871 191 873 205
rect 894 200 896 205
rect 899 203 901 205
rect 925 203 927 205
rect 890 196 896 200
rect 894 191 896 196
rect 899 191 901 193
rect 925 191 927 193
rect 946 191 948 205
rect 966 200 968 205
rect 971 203 973 205
rect 962 196 968 200
rect 966 191 968 196
rect 971 191 973 193
rect 989 191 991 205
rect 1034 195 1036 205
rect 1039 195 1041 202
rect 1055 195 1057 214
rect 1071 205 1073 214
rect 1076 212 1078 214
rect 1097 212 1099 214
rect 1113 211 1115 214
rect 1071 195 1073 198
rect 1076 195 1078 197
rect 1097 195 1099 197
rect 1113 195 1115 207
rect 1129 205 1131 214
rect 1134 212 1136 214
rect 1129 195 1131 198
rect 1134 195 1136 197
rect 1150 195 1152 214
rect 1166 211 1168 214
rect 1171 212 1173 214
rect 1166 195 1168 207
rect 1171 195 1173 202
rect 1187 195 1189 214
rect 1203 205 1205 214
rect 1208 212 1210 214
rect 1229 212 1231 214
rect 1245 211 1247 214
rect 1203 195 1205 198
rect 1208 195 1210 197
rect 1229 195 1231 197
rect 1245 195 1247 207
rect 1261 205 1263 214
rect 1266 212 1268 214
rect 1261 195 1263 198
rect 1266 195 1268 197
rect 1282 195 1284 214
rect 1298 211 1300 214
rect 1303 212 1305 214
rect 1298 195 1300 207
rect 1303 195 1305 202
rect 1319 195 1321 214
rect 1335 205 1337 214
rect 1340 212 1342 214
rect 1361 212 1363 214
rect 1377 211 1379 214
rect 1335 195 1337 198
rect 1340 195 1342 197
rect 1361 195 1363 197
rect 1377 195 1379 207
rect 1393 205 1395 214
rect 1398 212 1400 214
rect 1414 206 1416 214
rect 1528 213 1529 217
rect 1572 214 1573 218
rect 1597 217 1599 221
rect 1643 218 1645 220
rect 1511 209 1513 211
rect 1527 209 1529 213
rect 1543 209 1545 211
rect 1566 209 1568 211
rect 1571 209 1573 214
rect 1598 213 1599 217
rect 1644 214 1645 218
rect 1788 217 1790 220
rect 1832 218 1834 220
rect 1597 209 1599 213
rect 1618 209 1620 211
rect 1638 209 1640 211
rect 1643 209 1645 214
rect 1789 213 1790 217
rect 1833 214 1834 218
rect 1858 217 1860 221
rect 1904 218 1906 220
rect 1661 209 1663 211
rect 1745 209 1747 212
rect 1763 209 1765 212
rect 1788 209 1790 213
rect 1804 209 1806 211
rect 1827 209 1829 211
rect 1832 209 1834 214
rect 1859 213 1860 217
rect 1905 214 1906 218
rect 1858 209 1860 213
rect 1879 209 1881 211
rect 1899 209 1901 211
rect 1904 209 1906 214
rect 1922 209 1924 211
rect 1393 195 1395 198
rect 1398 195 1400 197
rect 1414 195 1416 202
rect 1511 191 1513 205
rect 1527 203 1529 205
rect 1527 191 1529 193
rect 1543 191 1545 205
rect 1566 200 1568 205
rect 1571 203 1573 205
rect 1597 203 1599 205
rect 1562 196 1568 200
rect 1566 191 1568 196
rect 1571 191 1573 193
rect 1597 191 1599 193
rect 1618 191 1620 205
rect 1638 200 1640 205
rect 1643 203 1645 205
rect 1634 196 1640 200
rect 1638 191 1640 196
rect 1643 191 1645 193
rect 1661 191 1663 205
rect 1711 202 1713 205
rect 1716 202 1718 205
rect 1745 200 1747 205
rect 783 186 785 188
rect 578 181 580 183
rect 594 180 596 183
rect 610 181 612 183
rect 633 181 635 183
rect 638 180 640 183
rect 664 180 666 183
rect 685 180 687 183
rect 705 181 707 183
rect 710 180 712 183
rect 728 181 730 183
rect 664 176 665 180
rect 1034 189 1036 191
rect 1039 188 1041 191
rect 1055 189 1057 191
rect 1071 189 1073 191
rect 1076 186 1078 191
rect 1097 186 1099 191
rect 1113 189 1115 191
rect 1129 189 1131 191
rect 1134 186 1136 191
rect 1150 189 1152 191
rect 1166 189 1168 191
rect 812 180 814 183
rect 830 180 832 183
rect 855 180 857 183
rect 871 181 873 183
rect 894 181 896 183
rect 899 180 901 183
rect 925 180 927 183
rect 946 180 948 183
rect 966 181 968 183
rect 971 180 973 183
rect 989 181 991 183
rect 1171 188 1173 191
rect 1187 189 1189 191
rect 1203 189 1205 191
rect 1208 186 1210 191
rect 1229 186 1231 191
rect 1245 189 1247 191
rect 1261 189 1263 191
rect 1266 186 1268 191
rect 1282 189 1284 191
rect 1298 189 1300 191
rect 1303 188 1305 191
rect 1319 189 1321 191
rect 1335 189 1337 191
rect 1340 186 1342 191
rect 1361 186 1363 191
rect 1377 189 1379 191
rect 1393 189 1395 191
rect 1398 186 1400 191
rect 1414 189 1416 191
rect 1711 186 1713 198
rect 1716 196 1718 198
rect 1745 191 1747 196
rect 1763 191 1765 205
rect 1788 203 1790 205
rect 1788 191 1790 193
rect 1804 191 1806 205
rect 1827 200 1829 205
rect 1832 203 1834 205
rect 1858 203 1860 205
rect 1823 196 1829 200
rect 1827 191 1829 196
rect 1832 191 1834 193
rect 1858 191 1860 193
rect 1879 191 1881 205
rect 1899 200 1901 205
rect 1904 203 1906 205
rect 1895 196 1901 200
rect 1899 191 1901 196
rect 1904 191 1906 193
rect 1922 191 1924 205
rect 1716 186 1718 188
rect 1511 181 1513 183
rect 1527 180 1529 183
rect 1543 181 1545 183
rect 1566 181 1568 183
rect 1571 180 1573 183
rect 1597 180 1599 183
rect 1618 180 1620 183
rect 1638 181 1640 183
rect 1643 180 1645 183
rect 1661 181 1663 183
rect 778 176 780 178
rect 594 173 596 176
rect 638 173 640 176
rect 664 173 666 176
rect 710 173 712 176
rect 783 173 785 178
rect 925 176 926 180
rect 855 173 857 176
rect 899 173 901 176
rect 925 173 927 176
rect 971 173 973 176
rect 1597 176 1598 180
rect 1745 180 1747 183
rect 1763 180 1765 183
rect 1788 180 1790 183
rect 1804 181 1806 183
rect 1827 181 1829 183
rect 1832 180 1834 183
rect 1858 180 1860 183
rect 1879 180 1881 183
rect 1899 181 1901 183
rect 1904 180 1906 183
rect 1922 181 1924 183
rect 1711 176 1713 178
rect 1527 173 1529 176
rect 1571 173 1573 176
rect 1597 173 1599 176
rect 1643 173 1645 176
rect 1716 173 1718 178
rect 1858 176 1859 180
rect 1788 173 1790 176
rect 1832 173 1834 176
rect 1858 173 1860 176
rect 1904 173 1906 176
rect 216 151 218 154
rect 240 151 242 154
rect 1149 151 1151 154
rect 1173 151 1175 154
rect 998 149 1001 151
rect 1005 149 1008 151
rect 216 145 218 147
rect 240 145 242 147
rect 1931 149 1934 151
rect 1938 149 1941 151
rect 1149 145 1151 147
rect 1173 145 1175 147
rect 236 140 238 142
rect 1169 140 1171 142
rect 236 133 238 136
rect 1169 133 1171 136
rect 225 122 227 124
rect 231 122 250 124
rect 1158 122 1160 124
rect 1164 122 1183 124
rect 216 117 218 119
rect 240 117 242 119
rect 1149 117 1151 119
rect 1173 117 1175 119
rect 216 110 218 113
rect 240 110 242 113
rect 872 112 874 114
rect 877 112 879 115
rect 893 112 895 114
rect 909 112 911 114
rect 914 112 916 115
rect 935 112 937 115
rect 951 112 953 115
rect 967 112 969 114
rect 972 112 974 115
rect 988 112 990 114
rect 1149 110 1151 113
rect 1173 110 1175 113
rect 1805 112 1807 114
rect 1810 112 1812 115
rect 1826 112 1828 114
rect 1842 112 1844 114
rect 1847 112 1849 115
rect 1868 112 1870 115
rect 1884 112 1886 115
rect 1900 112 1902 114
rect 1905 112 1907 115
rect 1921 112 1923 114
rect 872 99 874 104
rect 877 102 879 104
rect 872 85 874 95
rect 877 85 879 92
rect 893 85 895 104
rect 909 95 911 104
rect 914 102 916 104
rect 935 102 937 104
rect 951 101 953 104
rect 909 85 911 88
rect 914 85 916 87
rect 935 85 937 87
rect 951 85 953 97
rect 967 95 969 104
rect 972 102 974 104
rect 967 85 969 88
rect 972 85 974 87
rect 988 85 990 104
rect 1805 99 1807 104
rect 1810 102 1812 104
rect 1805 85 1807 95
rect 1810 85 1812 92
rect 1826 85 1828 104
rect 1842 95 1844 104
rect 1847 102 1849 104
rect 1868 102 1870 104
rect 1884 101 1886 104
rect 1842 85 1844 88
rect 1847 85 1849 87
rect 1868 85 1870 87
rect 1884 85 1886 97
rect 1900 95 1902 104
rect 1905 102 1907 104
rect 1900 85 1902 88
rect 1905 85 1907 87
rect 1921 85 1923 104
rect 101 82 103 84
rect 106 82 108 85
rect 122 82 124 84
rect 138 82 140 84
rect 143 82 145 85
rect 164 82 166 85
rect 180 82 182 85
rect 196 82 198 84
rect 201 82 203 85
rect 217 82 219 84
rect 233 82 235 84
rect 238 82 240 85
rect 254 82 256 84
rect 270 82 272 84
rect 275 82 277 85
rect 296 82 298 85
rect 312 82 314 85
rect 328 82 330 84
rect 333 82 335 85
rect 349 82 351 84
rect 365 82 367 84
rect 370 82 372 85
rect 386 82 388 84
rect 402 82 404 84
rect 407 82 409 85
rect 428 82 430 85
rect 444 82 446 85
rect 460 82 462 84
rect 465 82 467 85
rect 481 82 483 84
rect 1034 82 1036 84
rect 1039 82 1041 85
rect 1055 82 1057 84
rect 1071 82 1073 84
rect 1076 82 1078 85
rect 1097 82 1099 85
rect 1113 82 1115 85
rect 1129 82 1131 84
rect 1134 82 1136 85
rect 1150 82 1152 84
rect 1166 82 1168 84
rect 1171 82 1173 85
rect 1187 82 1189 84
rect 1203 82 1205 84
rect 1208 82 1210 85
rect 1229 82 1231 85
rect 1245 82 1247 85
rect 1261 82 1263 84
rect 1266 82 1268 85
rect 1282 82 1284 84
rect 1298 82 1300 84
rect 1303 82 1305 85
rect 1319 82 1321 84
rect 1335 82 1337 84
rect 1340 82 1342 85
rect 1361 82 1363 85
rect 1377 82 1379 85
rect 1393 82 1395 84
rect 1398 82 1400 85
rect 1414 82 1416 84
rect 872 79 874 81
rect 877 78 879 81
rect 893 79 895 81
rect 909 79 911 81
rect 914 76 916 81
rect 935 76 937 81
rect 951 79 953 81
rect 967 79 969 81
rect 972 76 974 81
rect 988 79 990 81
rect 101 69 103 74
rect 106 72 108 74
rect 101 55 103 65
rect 106 55 108 62
rect 122 55 124 74
rect 138 65 140 74
rect 143 72 145 74
rect 164 72 166 74
rect 180 71 182 74
rect 138 55 140 58
rect 143 55 145 57
rect 164 55 166 57
rect 180 55 182 67
rect 196 65 198 74
rect 201 72 203 74
rect 196 55 198 58
rect 201 55 203 57
rect 217 55 219 74
rect 233 71 235 74
rect 238 72 240 74
rect 233 55 235 67
rect 238 55 240 62
rect 254 55 256 74
rect 270 65 272 74
rect 275 72 277 74
rect 296 72 298 74
rect 312 71 314 74
rect 270 55 272 58
rect 275 55 277 57
rect 296 55 298 57
rect 312 55 314 67
rect 328 65 330 74
rect 333 72 335 74
rect 328 55 330 58
rect 333 55 335 57
rect 349 55 351 74
rect 365 71 367 74
rect 370 72 372 74
rect 365 55 367 67
rect 370 55 372 62
rect 386 55 388 74
rect 402 65 404 74
rect 407 72 409 74
rect 428 72 430 74
rect 444 71 446 74
rect 402 55 404 58
rect 407 55 409 57
rect 428 55 430 57
rect 444 55 446 67
rect 460 65 462 74
rect 465 72 467 74
rect 481 66 483 74
rect 1805 79 1807 81
rect 1810 78 1812 81
rect 1826 79 1828 81
rect 1842 79 1844 81
rect 1847 76 1849 81
rect 1868 76 1870 81
rect 1884 79 1886 81
rect 1900 79 1902 81
rect 1905 76 1907 81
rect 1921 79 1923 81
rect 1034 69 1036 74
rect 1039 72 1041 74
rect 460 55 462 58
rect 465 55 467 57
rect 481 55 483 62
rect 1034 55 1036 65
rect 1039 55 1041 62
rect 1055 55 1057 74
rect 1071 65 1073 74
rect 1076 72 1078 74
rect 1097 72 1099 74
rect 1113 71 1115 74
rect 1071 55 1073 58
rect 1076 55 1078 57
rect 1097 55 1099 57
rect 1113 55 1115 67
rect 1129 65 1131 74
rect 1134 72 1136 74
rect 1129 55 1131 58
rect 1134 55 1136 57
rect 1150 55 1152 74
rect 1166 71 1168 74
rect 1171 72 1173 74
rect 1166 55 1168 67
rect 1171 55 1173 62
rect 1187 55 1189 74
rect 1203 65 1205 74
rect 1208 72 1210 74
rect 1229 72 1231 74
rect 1245 71 1247 74
rect 1203 55 1205 58
rect 1208 55 1210 57
rect 1229 55 1231 57
rect 1245 55 1247 67
rect 1261 65 1263 74
rect 1266 72 1268 74
rect 1261 55 1263 58
rect 1266 55 1268 57
rect 1282 55 1284 74
rect 1298 71 1300 74
rect 1303 72 1305 74
rect 1298 55 1300 67
rect 1303 55 1305 62
rect 1319 55 1321 74
rect 1335 65 1337 74
rect 1340 72 1342 74
rect 1361 72 1363 74
rect 1377 71 1379 74
rect 1335 55 1337 58
rect 1340 55 1342 57
rect 1361 55 1363 57
rect 1377 55 1379 67
rect 1393 65 1395 74
rect 1398 72 1400 74
rect 1414 66 1416 74
rect 1393 55 1395 58
rect 1398 55 1400 57
rect 1414 55 1416 62
rect 101 49 103 51
rect 106 48 108 51
rect 122 49 124 51
rect 138 49 140 51
rect 143 46 145 51
rect 164 46 166 51
rect 180 49 182 51
rect 196 49 198 51
rect 201 46 203 51
rect 217 49 219 51
rect 233 49 235 51
rect 238 48 240 51
rect 254 49 256 51
rect 270 49 272 51
rect 275 46 277 51
rect 296 46 298 51
rect 312 49 314 51
rect 328 49 330 51
rect 333 46 335 51
rect 349 49 351 51
rect 365 49 367 51
rect 370 48 372 51
rect 386 49 388 51
rect 402 49 404 51
rect 407 46 409 51
rect 428 46 430 51
rect 444 49 446 51
rect 460 49 462 51
rect 465 46 467 51
rect 481 49 483 51
rect 1034 49 1036 51
rect 1039 48 1041 51
rect 1055 49 1057 51
rect 1071 49 1073 51
rect 1076 46 1078 51
rect 1097 46 1099 51
rect 1113 49 1115 51
rect 1129 49 1131 51
rect 1134 46 1136 51
rect 1150 49 1152 51
rect 1166 49 1168 51
rect 1171 48 1173 51
rect 1187 49 1189 51
rect 1203 49 1205 51
rect 1208 46 1210 51
rect 1229 46 1231 51
rect 1245 49 1247 51
rect 1261 49 1263 51
rect 1266 46 1268 51
rect 1282 49 1284 51
rect 1298 49 1300 51
rect 1303 48 1305 51
rect 1319 49 1321 51
rect 1335 49 1337 51
rect 1340 46 1342 51
rect 1361 46 1363 51
rect 1377 49 1379 51
rect 1393 49 1395 51
rect 1398 46 1400 51
rect 1414 49 1416 51
rect 872 26 874 28
rect 877 26 879 29
rect 893 26 895 28
rect 909 26 911 28
rect 914 26 916 29
rect 935 26 937 29
rect 951 26 953 29
rect 967 26 969 28
rect 972 26 974 29
rect 988 26 990 28
rect 1805 26 1807 28
rect 1810 26 1812 29
rect 1826 26 1828 28
rect 1842 26 1844 28
rect 1847 26 1849 29
rect 1868 26 1870 29
rect 1884 26 1886 29
rect 1900 26 1902 28
rect 1905 26 1907 29
rect 1921 26 1923 28
rect 872 13 874 18
rect 877 16 879 18
rect 872 -1 874 9
rect 877 -1 879 6
rect 893 -1 895 18
rect 909 9 911 18
rect 914 16 916 18
rect 935 16 937 18
rect 951 15 953 18
rect 909 -1 911 2
rect 914 -1 916 1
rect 935 -1 937 1
rect 951 -1 953 11
rect 967 9 969 18
rect 972 16 974 18
rect 967 -1 969 2
rect 972 -1 974 1
rect 988 -1 990 18
rect 1805 13 1807 18
rect 1810 16 1812 18
rect 1010 5 1013 7
rect 1017 5 1020 7
rect 1805 -1 1807 9
rect 1810 -1 1812 6
rect 1826 -1 1828 18
rect 1842 9 1844 18
rect 1847 16 1849 18
rect 1868 16 1870 18
rect 1884 15 1886 18
rect 1842 -1 1844 2
rect 1847 -1 1849 1
rect 1868 -1 1870 1
rect 1884 -1 1886 11
rect 1900 9 1902 18
rect 1905 16 1907 18
rect 1900 -1 1902 2
rect 1905 -1 1907 1
rect 1921 -1 1923 18
rect 1943 5 1946 7
rect 1950 5 1953 7
rect 101 -4 103 -2
rect 106 -4 108 -1
rect 122 -4 124 -2
rect 138 -4 140 -2
rect 143 -4 145 -1
rect 164 -4 166 -1
rect 180 -4 182 -1
rect 196 -4 198 -2
rect 201 -4 203 -1
rect 217 -4 219 -2
rect 233 -4 235 -2
rect 238 -4 240 -1
rect 254 -4 256 -2
rect 270 -4 272 -2
rect 275 -4 277 -1
rect 296 -4 298 -1
rect 312 -4 314 -1
rect 328 -4 330 -2
rect 333 -4 335 -1
rect 349 -4 351 -2
rect 365 -4 367 -2
rect 370 -4 372 -1
rect 386 -4 388 -2
rect 402 -4 404 -2
rect 407 -4 409 -1
rect 428 -4 430 -1
rect 444 -4 446 -1
rect 460 -4 462 -2
rect 465 -4 467 -1
rect 481 -4 483 -2
rect 1034 -4 1036 -2
rect 1039 -4 1041 -1
rect 1055 -4 1057 -2
rect 1071 -4 1073 -2
rect 1076 -4 1078 -1
rect 1097 -4 1099 -1
rect 1113 -4 1115 -1
rect 1129 -4 1131 -2
rect 1134 -4 1136 -1
rect 1150 -4 1152 -2
rect 1166 -4 1168 -2
rect 1171 -4 1173 -1
rect 1187 -4 1189 -2
rect 1203 -4 1205 -2
rect 1208 -4 1210 -1
rect 1229 -4 1231 -1
rect 1245 -4 1247 -1
rect 1261 -4 1263 -2
rect 1266 -4 1268 -1
rect 1282 -4 1284 -2
rect 1298 -4 1300 -2
rect 1303 -4 1305 -1
rect 1319 -4 1321 -2
rect 1335 -4 1337 -2
rect 1340 -4 1342 -1
rect 1361 -4 1363 -1
rect 1377 -4 1379 -1
rect 1393 -4 1395 -2
rect 1398 -4 1400 -1
rect 1414 -4 1416 -2
rect 872 -7 874 -5
rect 877 -8 879 -5
rect 893 -7 895 -5
rect 909 -7 911 -5
rect 914 -10 916 -5
rect 935 -10 937 -5
rect 951 -7 953 -5
rect 967 -7 969 -5
rect 972 -10 974 -5
rect 988 -7 990 -5
rect 101 -17 103 -12
rect 106 -14 108 -12
rect 101 -31 103 -21
rect 106 -31 108 -24
rect 122 -31 124 -12
rect 138 -21 140 -12
rect 143 -14 145 -12
rect 164 -14 166 -12
rect 180 -15 182 -12
rect 138 -31 140 -28
rect 143 -31 145 -29
rect 164 -31 166 -29
rect 180 -31 182 -19
rect 196 -21 198 -12
rect 201 -14 203 -12
rect 196 -31 198 -28
rect 201 -31 203 -29
rect 217 -31 219 -12
rect 233 -15 235 -12
rect 238 -14 240 -12
rect 233 -31 235 -19
rect 238 -31 240 -24
rect 254 -31 256 -12
rect 270 -21 272 -12
rect 275 -14 277 -12
rect 296 -14 298 -12
rect 312 -15 314 -12
rect 270 -31 272 -28
rect 275 -31 277 -29
rect 296 -31 298 -29
rect 312 -31 314 -19
rect 328 -21 330 -12
rect 333 -14 335 -12
rect 328 -31 330 -28
rect 333 -31 335 -29
rect 349 -31 351 -12
rect 365 -15 367 -12
rect 370 -14 372 -12
rect 365 -31 367 -19
rect 370 -31 372 -24
rect 386 -31 388 -12
rect 402 -21 404 -12
rect 407 -14 409 -12
rect 428 -14 430 -12
rect 444 -15 446 -12
rect 402 -31 404 -28
rect 407 -31 409 -29
rect 428 -31 430 -29
rect 444 -31 446 -19
rect 460 -21 462 -12
rect 465 -14 467 -12
rect 481 -20 483 -12
rect 1805 -7 1807 -5
rect 1810 -8 1812 -5
rect 1826 -7 1828 -5
rect 1842 -7 1844 -5
rect 1847 -10 1849 -5
rect 1868 -10 1870 -5
rect 1884 -7 1886 -5
rect 1900 -7 1902 -5
rect 1905 -10 1907 -5
rect 1921 -7 1923 -5
rect 1034 -17 1036 -12
rect 1039 -14 1041 -12
rect 460 -31 462 -28
rect 465 -31 467 -29
rect 481 -31 483 -24
rect 1034 -31 1036 -21
rect 1039 -31 1041 -24
rect 1055 -31 1057 -12
rect 1071 -21 1073 -12
rect 1076 -14 1078 -12
rect 1097 -14 1099 -12
rect 1113 -15 1115 -12
rect 1071 -31 1073 -28
rect 1076 -31 1078 -29
rect 1097 -31 1099 -29
rect 1113 -31 1115 -19
rect 1129 -21 1131 -12
rect 1134 -14 1136 -12
rect 1129 -31 1131 -28
rect 1134 -31 1136 -29
rect 1150 -31 1152 -12
rect 1166 -15 1168 -12
rect 1171 -14 1173 -12
rect 1166 -31 1168 -19
rect 1171 -31 1173 -24
rect 1187 -31 1189 -12
rect 1203 -21 1205 -12
rect 1208 -14 1210 -12
rect 1229 -14 1231 -12
rect 1245 -15 1247 -12
rect 1203 -31 1205 -28
rect 1208 -31 1210 -29
rect 1229 -31 1231 -29
rect 1245 -31 1247 -19
rect 1261 -21 1263 -12
rect 1266 -14 1268 -12
rect 1261 -31 1263 -28
rect 1266 -31 1268 -29
rect 1282 -31 1284 -12
rect 1298 -15 1300 -12
rect 1303 -14 1305 -12
rect 1298 -31 1300 -19
rect 1303 -31 1305 -24
rect 1319 -31 1321 -12
rect 1335 -21 1337 -12
rect 1340 -14 1342 -12
rect 1361 -14 1363 -12
rect 1377 -15 1379 -12
rect 1335 -31 1337 -28
rect 1340 -31 1342 -29
rect 1361 -31 1363 -29
rect 1377 -31 1379 -19
rect 1393 -21 1395 -12
rect 1398 -14 1400 -12
rect 1414 -20 1416 -12
rect 1393 -31 1395 -28
rect 1398 -31 1400 -29
rect 1414 -31 1416 -24
rect 101 -37 103 -35
rect 106 -38 108 -35
rect 122 -37 124 -35
rect 138 -37 140 -35
rect 143 -40 145 -35
rect 164 -40 166 -35
rect 180 -37 182 -35
rect 196 -37 198 -35
rect 201 -40 203 -35
rect 217 -37 219 -35
rect 233 -37 235 -35
rect 238 -38 240 -35
rect 254 -37 256 -35
rect 270 -37 272 -35
rect 275 -40 277 -35
rect 296 -40 298 -35
rect 312 -37 314 -35
rect 328 -37 330 -35
rect 333 -40 335 -35
rect 349 -37 351 -35
rect 365 -37 367 -35
rect 370 -38 372 -35
rect 386 -37 388 -35
rect 402 -37 404 -35
rect 407 -40 409 -35
rect 428 -40 430 -35
rect 444 -37 446 -35
rect 460 -37 462 -35
rect 465 -40 467 -35
rect 481 -37 483 -35
rect 1034 -37 1036 -35
rect 1039 -38 1041 -35
rect 1055 -37 1057 -35
rect 1071 -37 1073 -35
rect 1076 -40 1078 -35
rect 1097 -40 1099 -35
rect 1113 -37 1115 -35
rect 1129 -37 1131 -35
rect 1134 -40 1136 -35
rect 1150 -37 1152 -35
rect 1166 -37 1168 -35
rect 1171 -38 1173 -35
rect 1187 -37 1189 -35
rect 1203 -37 1205 -35
rect 1208 -40 1210 -35
rect 1229 -40 1231 -35
rect 1245 -37 1247 -35
rect 1261 -37 1263 -35
rect 1266 -40 1268 -35
rect 1282 -37 1284 -35
rect 1298 -37 1300 -35
rect 1303 -38 1305 -35
rect 1319 -37 1321 -35
rect 1335 -37 1337 -35
rect 1340 -40 1342 -35
rect 1361 -40 1363 -35
rect 1377 -37 1379 -35
rect 1393 -37 1395 -35
rect 1398 -40 1400 -35
rect 1414 -37 1416 -35
rect 333 -75 335 -72
rect 357 -75 359 -72
rect 1266 -75 1268 -72
rect 1290 -75 1292 -72
rect 333 -81 335 -79
rect 357 -81 359 -79
rect 1266 -81 1268 -79
rect 1290 -81 1292 -79
rect 353 -86 355 -84
rect 1286 -86 1288 -84
rect 353 -93 355 -90
rect 1286 -93 1288 -90
rect 342 -104 344 -102
rect 348 -104 367 -102
rect 1275 -104 1277 -102
rect 1281 -104 1300 -102
rect 333 -109 335 -107
rect 357 -109 359 -107
rect 1266 -109 1268 -107
rect 1290 -109 1292 -107
rect 333 -116 335 -113
rect 357 -116 359 -113
rect 1266 -116 1268 -113
rect 1290 -116 1292 -113
rect 101 -144 103 -142
rect 106 -144 108 -141
rect 122 -144 124 -142
rect 138 -144 140 -142
rect 143 -144 145 -141
rect 164 -144 166 -141
rect 180 -144 182 -141
rect 196 -144 198 -142
rect 201 -144 203 -141
rect 217 -144 219 -142
rect 233 -144 235 -142
rect 238 -144 240 -141
rect 254 -144 256 -142
rect 270 -144 272 -142
rect 275 -144 277 -141
rect 296 -144 298 -141
rect 312 -144 314 -141
rect 328 -144 330 -142
rect 333 -144 335 -141
rect 349 -144 351 -142
rect 365 -144 367 -142
rect 370 -144 372 -141
rect 386 -144 388 -142
rect 402 -144 404 -142
rect 407 -144 409 -141
rect 428 -144 430 -141
rect 444 -144 446 -141
rect 460 -144 462 -142
rect 465 -144 467 -141
rect 481 -144 483 -142
rect 1034 -144 1036 -142
rect 1039 -144 1041 -141
rect 1055 -144 1057 -142
rect 1071 -144 1073 -142
rect 1076 -144 1078 -141
rect 1097 -144 1099 -141
rect 1113 -144 1115 -141
rect 1129 -144 1131 -142
rect 1134 -144 1136 -141
rect 1150 -144 1152 -142
rect 1166 -144 1168 -142
rect 1171 -144 1173 -141
rect 1187 -144 1189 -142
rect 1203 -144 1205 -142
rect 1208 -144 1210 -141
rect 1229 -144 1231 -141
rect 1245 -144 1247 -141
rect 1261 -144 1263 -142
rect 1266 -144 1268 -141
rect 1282 -144 1284 -142
rect 1298 -144 1300 -142
rect 1303 -144 1305 -141
rect 1319 -144 1321 -142
rect 1335 -144 1337 -142
rect 1340 -144 1342 -141
rect 1361 -144 1363 -141
rect 1377 -144 1379 -141
rect 1393 -144 1395 -142
rect 1398 -144 1400 -141
rect 1414 -144 1416 -142
rect 101 -157 103 -152
rect 106 -154 108 -152
rect 101 -171 103 -161
rect 106 -171 108 -164
rect 122 -171 124 -152
rect 138 -161 140 -152
rect 143 -154 145 -152
rect 164 -154 166 -152
rect 180 -155 182 -152
rect 138 -171 140 -168
rect 143 -171 145 -169
rect 164 -171 166 -169
rect 180 -171 182 -159
rect 196 -161 198 -152
rect 201 -154 203 -152
rect 196 -171 198 -168
rect 201 -171 203 -169
rect 217 -171 219 -152
rect 233 -155 235 -152
rect 238 -154 240 -152
rect 233 -171 235 -159
rect 238 -171 240 -164
rect 254 -171 256 -152
rect 270 -161 272 -152
rect 275 -154 277 -152
rect 296 -154 298 -152
rect 312 -155 314 -152
rect 270 -171 272 -168
rect 275 -171 277 -169
rect 296 -171 298 -169
rect 312 -171 314 -159
rect 328 -161 330 -152
rect 333 -154 335 -152
rect 328 -171 330 -168
rect 333 -171 335 -169
rect 349 -171 351 -152
rect 365 -155 367 -152
rect 370 -154 372 -152
rect 365 -171 367 -159
rect 370 -171 372 -164
rect 386 -171 388 -152
rect 402 -161 404 -152
rect 407 -154 409 -152
rect 428 -154 430 -152
rect 444 -155 446 -152
rect 402 -171 404 -168
rect 407 -171 409 -169
rect 428 -171 430 -169
rect 444 -171 446 -159
rect 460 -161 462 -152
rect 465 -154 467 -152
rect 481 -160 483 -152
rect 1034 -157 1036 -152
rect 1039 -154 1041 -152
rect 460 -171 462 -168
rect 465 -171 467 -169
rect 481 -171 483 -164
rect 1034 -171 1036 -161
rect 1039 -171 1041 -164
rect 1055 -171 1057 -152
rect 1071 -161 1073 -152
rect 1076 -154 1078 -152
rect 1097 -154 1099 -152
rect 1113 -155 1115 -152
rect 1071 -171 1073 -168
rect 1076 -171 1078 -169
rect 1097 -171 1099 -169
rect 1113 -171 1115 -159
rect 1129 -161 1131 -152
rect 1134 -154 1136 -152
rect 1129 -171 1131 -168
rect 1134 -171 1136 -169
rect 1150 -171 1152 -152
rect 1166 -155 1168 -152
rect 1171 -154 1173 -152
rect 1166 -171 1168 -159
rect 1171 -171 1173 -164
rect 1187 -171 1189 -152
rect 1203 -161 1205 -152
rect 1208 -154 1210 -152
rect 1229 -154 1231 -152
rect 1245 -155 1247 -152
rect 1203 -171 1205 -168
rect 1208 -171 1210 -169
rect 1229 -171 1231 -169
rect 1245 -171 1247 -159
rect 1261 -161 1263 -152
rect 1266 -154 1268 -152
rect 1261 -171 1263 -168
rect 1266 -171 1268 -169
rect 1282 -171 1284 -152
rect 1298 -155 1300 -152
rect 1303 -154 1305 -152
rect 1298 -171 1300 -159
rect 1303 -171 1305 -164
rect 1319 -171 1321 -152
rect 1335 -161 1337 -152
rect 1340 -154 1342 -152
rect 1361 -154 1363 -152
rect 1377 -155 1379 -152
rect 1335 -171 1337 -168
rect 1340 -171 1342 -169
rect 1361 -171 1363 -169
rect 1377 -171 1379 -159
rect 1393 -161 1395 -152
rect 1398 -154 1400 -152
rect 1414 -160 1416 -152
rect 1393 -171 1395 -168
rect 1398 -171 1400 -169
rect 1414 -171 1416 -164
rect 101 -177 103 -175
rect 106 -178 108 -175
rect 122 -177 124 -175
rect 138 -177 140 -175
rect 143 -180 145 -175
rect 164 -180 166 -175
rect 180 -177 182 -175
rect 196 -177 198 -175
rect 201 -180 203 -175
rect 217 -177 219 -175
rect 233 -177 235 -175
rect 238 -178 240 -175
rect 254 -177 256 -175
rect 270 -177 272 -175
rect 275 -180 277 -175
rect 296 -180 298 -175
rect 312 -177 314 -175
rect 328 -177 330 -175
rect 333 -180 335 -175
rect 349 -177 351 -175
rect 365 -177 367 -175
rect 370 -178 372 -175
rect 386 -177 388 -175
rect 402 -177 404 -175
rect 407 -180 409 -175
rect 428 -180 430 -175
rect 444 -177 446 -175
rect 460 -177 462 -175
rect 465 -180 467 -175
rect 481 -177 483 -175
rect 1034 -177 1036 -175
rect 1039 -178 1041 -175
rect 1055 -177 1057 -175
rect 1071 -177 1073 -175
rect 1076 -180 1078 -175
rect 1097 -180 1099 -175
rect 1113 -177 1115 -175
rect 1129 -177 1131 -175
rect 1134 -180 1136 -175
rect 1150 -177 1152 -175
rect 1166 -177 1168 -175
rect 1171 -178 1173 -175
rect 1187 -177 1189 -175
rect 1203 -177 1205 -175
rect 1208 -180 1210 -175
rect 1229 -180 1231 -175
rect 1245 -177 1247 -175
rect 1261 -177 1263 -175
rect 1266 -180 1268 -175
rect 1282 -177 1284 -175
rect 1298 -177 1300 -175
rect 1303 -178 1305 -175
rect 1319 -177 1321 -175
rect 1335 -177 1337 -175
rect 1340 -180 1342 -175
rect 1361 -180 1363 -175
rect 1377 -177 1379 -175
rect 1393 -177 1395 -175
rect 1398 -180 1400 -175
rect 1414 -177 1416 -175
<< polycontact >>
rect 578 1740 582 1744
rect 615 1740 619 1744
rect 635 1740 639 1744
rect 673 1740 677 1744
rect 710 1740 714 1744
rect 747 1740 751 1744
rect 767 1740 771 1744
rect 805 1740 809 1744
rect 842 1740 846 1744
rect 879 1740 883 1744
rect 899 1740 903 1744
rect 937 1740 941 1744
rect 974 1740 978 1744
rect 1011 1740 1015 1744
rect 1031 1740 1035 1744
rect 1069 1740 1073 1744
rect 1511 1740 1515 1744
rect 1548 1740 1552 1744
rect 1568 1740 1572 1744
rect 1606 1740 1610 1744
rect 1643 1740 1647 1744
rect 1680 1740 1684 1744
rect 1700 1740 1704 1744
rect 1738 1740 1742 1744
rect 1775 1740 1779 1744
rect 1812 1740 1816 1744
rect 1832 1740 1836 1744
rect 1870 1740 1874 1744
rect 1907 1740 1911 1744
rect 1944 1740 1948 1744
rect 1964 1740 1968 1744
rect 2002 1740 2006 1744
rect 572 1720 576 1724
rect 590 1722 594 1726
rect 238 1707 242 1711
rect 275 1707 279 1711
rect 295 1707 299 1711
rect 333 1707 337 1711
rect 650 1722 654 1726
rect 608 1713 612 1720
rect 666 1713 670 1720
rect 687 1717 691 1721
rect 704 1720 708 1724
rect 722 1722 726 1726
rect 782 1722 786 1726
rect 740 1713 744 1720
rect 798 1713 802 1720
rect 819 1717 823 1721
rect 836 1720 840 1724
rect 854 1722 858 1726
rect 914 1722 918 1726
rect 872 1713 876 1720
rect 930 1713 934 1720
rect 951 1717 955 1721
rect 968 1720 972 1724
rect 986 1722 990 1726
rect 1046 1722 1050 1726
rect 1004 1713 1008 1720
rect 1062 1713 1066 1720
rect 1083 1717 1087 1721
rect 1505 1720 1509 1724
rect 1523 1722 1527 1726
rect 1171 1707 1175 1711
rect 1208 1707 1212 1711
rect 1228 1707 1232 1711
rect 1266 1707 1270 1711
rect 1583 1722 1587 1726
rect 1541 1713 1545 1720
rect 1599 1713 1603 1720
rect 1620 1717 1624 1721
rect 1637 1720 1641 1724
rect 1655 1722 1659 1726
rect 1715 1722 1719 1726
rect 1673 1713 1677 1720
rect 1731 1713 1735 1720
rect 1752 1717 1756 1721
rect 1769 1720 1773 1724
rect 1787 1722 1791 1726
rect 1847 1722 1851 1726
rect 1805 1713 1809 1720
rect 1863 1713 1867 1720
rect 1884 1717 1888 1721
rect 1901 1720 1905 1724
rect 1919 1722 1923 1726
rect 1979 1722 1983 1726
rect 1937 1713 1941 1720
rect 1995 1713 1999 1720
rect 2016 1717 2020 1721
rect 578 1699 582 1703
rect 615 1697 619 1701
rect 635 1697 639 1701
rect 671 1697 675 1701
rect 710 1699 714 1703
rect 747 1697 751 1701
rect 767 1697 771 1701
rect 803 1697 807 1701
rect 842 1699 846 1703
rect 879 1697 883 1701
rect 899 1697 903 1701
rect 935 1697 939 1701
rect 974 1699 978 1703
rect 1011 1697 1015 1701
rect 1031 1697 1035 1701
rect 1067 1697 1071 1701
rect 1511 1699 1515 1703
rect 1548 1697 1552 1701
rect 1568 1697 1572 1701
rect 1604 1697 1608 1701
rect 1643 1699 1647 1703
rect 1680 1697 1684 1701
rect 1700 1697 1704 1701
rect 1736 1697 1740 1701
rect 1775 1699 1779 1703
rect 1812 1697 1816 1701
rect 1832 1697 1836 1701
rect 1868 1697 1872 1701
rect 1907 1699 1911 1703
rect 1944 1697 1948 1701
rect 1964 1697 1968 1701
rect 2000 1697 2004 1701
rect 232 1687 236 1691
rect 250 1689 254 1693
rect 310 1689 314 1693
rect 268 1680 272 1687
rect 326 1680 330 1687
rect 345 1684 349 1688
rect 1165 1687 1169 1691
rect 1183 1689 1187 1693
rect 1243 1689 1247 1693
rect 1201 1680 1205 1687
rect 1259 1680 1263 1687
rect 1278 1684 1282 1688
rect 238 1666 242 1670
rect 275 1664 279 1668
rect 295 1664 299 1668
rect 331 1664 335 1668
rect 594 1656 598 1660
rect 638 1656 642 1660
rect 665 1656 669 1660
rect 710 1656 714 1660
rect 783 1663 787 1667
rect 356 1643 360 1647
rect 748 1649 752 1653
rect 239 1634 243 1638
rect 574 1636 578 1640
rect 606 1637 610 1641
rect 625 1636 629 1640
rect 681 1637 685 1641
rect 697 1636 701 1640
rect 724 1636 728 1640
rect 864 1663 868 1667
rect 1171 1666 1175 1670
rect 775 1645 779 1649
rect 802 1641 806 1645
rect 829 1649 833 1653
rect 1208 1664 1212 1668
rect 1228 1664 1232 1668
rect 1264 1664 1268 1668
rect 856 1645 860 1649
rect 883 1641 887 1645
rect 1527 1656 1531 1660
rect 1571 1656 1575 1660
rect 1598 1656 1602 1660
rect 1643 1656 1647 1660
rect 1716 1663 1720 1667
rect 1289 1643 1293 1647
rect 1681 1649 1685 1653
rect 781 1627 785 1631
rect 1172 1634 1176 1638
rect 1507 1636 1511 1640
rect 862 1627 866 1631
rect 1539 1637 1543 1641
rect 1558 1636 1562 1640
rect 1614 1637 1618 1641
rect 1630 1636 1634 1640
rect 1657 1636 1661 1640
rect 1797 1663 1801 1667
rect 1708 1645 1712 1649
rect 1735 1641 1739 1645
rect 1762 1649 1766 1653
rect 1789 1645 1793 1649
rect 1816 1641 1820 1645
rect 1714 1627 1718 1631
rect 1795 1627 1799 1631
rect 591 1619 595 1623
rect 635 1618 639 1622
rect 660 1619 665 1623
rect 707 1618 711 1622
rect 1524 1619 1528 1623
rect 1568 1618 1572 1622
rect 1593 1619 1598 1623
rect 1640 1618 1644 1622
rect 238 1605 242 1609
rect 276 1605 280 1609
rect 296 1605 300 1609
rect 333 1605 337 1609
rect 1171 1605 1175 1609
rect 1209 1605 1213 1609
rect 1229 1605 1233 1609
rect 1266 1605 1270 1609
rect 226 1582 230 1586
rect 261 1587 265 1591
rect 245 1578 249 1585
rect 303 1578 307 1585
rect 321 1587 325 1591
rect 591 1589 595 1593
rect 635 1590 639 1594
rect 339 1585 343 1589
rect 660 1589 665 1593
rect 707 1590 711 1594
rect 783 1587 787 1591
rect 864 1587 868 1591
rect 574 1572 578 1576
rect 240 1562 244 1566
rect 276 1562 280 1566
rect 296 1562 300 1566
rect 333 1564 337 1568
rect 606 1571 610 1575
rect 625 1572 629 1576
rect 681 1571 685 1575
rect 697 1572 701 1576
rect 724 1572 728 1576
rect 772 1571 778 1575
rect 853 1571 859 1575
rect 1159 1582 1163 1586
rect 1194 1587 1198 1591
rect 1178 1578 1182 1585
rect 1236 1578 1240 1585
rect 1254 1587 1258 1591
rect 1524 1589 1528 1593
rect 1568 1590 1572 1594
rect 1272 1585 1276 1589
rect 1593 1589 1598 1593
rect 1640 1590 1644 1594
rect 1716 1587 1720 1591
rect 1797 1587 1801 1591
rect 1507 1572 1511 1576
rect 1173 1562 1177 1566
rect 1209 1562 1213 1566
rect 1229 1562 1233 1566
rect 1266 1564 1270 1568
rect 1539 1571 1543 1575
rect 1558 1572 1562 1576
rect 1614 1571 1618 1575
rect 1630 1572 1634 1576
rect 1657 1572 1661 1576
rect 1705 1571 1711 1575
rect 1786 1571 1792 1575
rect 594 1552 598 1556
rect 638 1552 642 1556
rect 665 1552 669 1556
rect 710 1552 714 1556
rect 781 1551 785 1555
rect 862 1551 866 1555
rect 1527 1552 1531 1556
rect 1571 1552 1575 1556
rect 1598 1552 1602 1556
rect 1643 1552 1647 1556
rect 1714 1551 1718 1555
rect 1795 1551 1799 1555
rect 783 1531 787 1535
rect 594 1524 598 1528
rect 638 1524 642 1528
rect 665 1524 669 1528
rect 710 1524 714 1528
rect 888 1531 892 1535
rect 775 1513 779 1517
rect 574 1504 578 1508
rect 606 1505 610 1509
rect 625 1504 629 1508
rect 681 1505 685 1509
rect 697 1504 701 1508
rect 724 1504 728 1508
rect 802 1509 806 1513
rect 853 1517 857 1521
rect 1716 1531 1720 1535
rect 880 1513 884 1517
rect 907 1509 911 1513
rect 1527 1524 1531 1528
rect 1571 1524 1575 1528
rect 1598 1524 1602 1528
rect 1643 1524 1647 1528
rect 1821 1531 1825 1535
rect 1708 1513 1712 1517
rect 1507 1504 1511 1508
rect 781 1495 785 1499
rect 886 1495 890 1499
rect 1539 1505 1543 1509
rect 1558 1504 1562 1508
rect 1614 1505 1618 1509
rect 1630 1504 1634 1508
rect 1657 1504 1661 1508
rect 1735 1509 1739 1513
rect 1786 1517 1790 1521
rect 1813 1513 1817 1517
rect 1840 1509 1844 1513
rect 1714 1495 1718 1499
rect 1819 1495 1823 1499
rect 591 1487 595 1491
rect 635 1486 639 1490
rect 660 1487 665 1491
rect 707 1486 711 1490
rect 1524 1487 1528 1491
rect 1568 1486 1572 1490
rect 1593 1487 1598 1491
rect 1640 1486 1644 1490
rect 591 1457 595 1461
rect 635 1458 639 1462
rect 660 1457 665 1461
rect 707 1458 711 1462
rect 783 1456 787 1460
rect 888 1456 892 1460
rect 1524 1457 1528 1461
rect 1568 1458 1572 1462
rect 1593 1457 1598 1461
rect 1640 1458 1644 1462
rect 1716 1456 1720 1460
rect 1821 1456 1825 1460
rect 574 1440 578 1444
rect 606 1439 610 1443
rect 625 1440 629 1444
rect 681 1439 685 1443
rect 697 1440 701 1444
rect 724 1440 728 1444
rect 772 1440 778 1444
rect 877 1440 883 1444
rect 1507 1440 1511 1444
rect 1539 1439 1543 1443
rect 1558 1440 1562 1444
rect 1614 1439 1618 1443
rect 1630 1440 1634 1444
rect 1657 1440 1661 1444
rect 1705 1440 1711 1444
rect 1810 1440 1816 1444
rect 594 1420 598 1424
rect 638 1420 642 1424
rect 665 1420 669 1424
rect 710 1420 714 1424
rect 781 1420 785 1424
rect 886 1420 890 1424
rect 1527 1420 1531 1424
rect 1571 1420 1575 1424
rect 1598 1420 1602 1424
rect 1643 1420 1647 1424
rect 1714 1420 1718 1424
rect 1819 1420 1823 1424
rect 783 1399 787 1403
rect 594 1392 598 1396
rect 638 1392 642 1396
rect 665 1392 669 1396
rect 710 1392 714 1396
rect 864 1399 868 1403
rect 775 1381 779 1385
rect 574 1372 578 1376
rect 606 1373 610 1377
rect 625 1372 629 1376
rect 681 1373 685 1377
rect 697 1372 701 1376
rect 724 1372 728 1376
rect 802 1377 806 1381
rect 829 1385 833 1389
rect 954 1399 958 1403
rect 856 1381 860 1385
rect 883 1377 887 1381
rect 919 1385 923 1389
rect 1716 1399 1720 1403
rect 946 1381 950 1385
rect 973 1377 977 1381
rect 1527 1392 1531 1396
rect 1571 1392 1575 1396
rect 1598 1392 1602 1396
rect 1643 1392 1647 1396
rect 1797 1399 1801 1403
rect 1708 1381 1712 1385
rect 1507 1372 1511 1376
rect 781 1363 785 1367
rect 862 1363 866 1367
rect 952 1363 956 1367
rect 1539 1373 1543 1377
rect 1558 1372 1562 1376
rect 1614 1373 1618 1377
rect 1630 1372 1634 1376
rect 1657 1372 1661 1376
rect 1735 1377 1739 1381
rect 1762 1385 1766 1389
rect 1887 1399 1891 1403
rect 1789 1381 1793 1385
rect 1816 1377 1820 1381
rect 1852 1385 1856 1389
rect 1879 1381 1883 1385
rect 1906 1377 1910 1381
rect 1714 1363 1718 1367
rect 1795 1363 1799 1367
rect 1885 1363 1889 1367
rect 591 1355 595 1359
rect 635 1354 639 1358
rect 660 1355 665 1359
rect 707 1354 711 1358
rect 1524 1355 1528 1359
rect 1568 1354 1572 1358
rect 1593 1355 1598 1359
rect 1640 1354 1644 1358
rect 591 1325 595 1329
rect 635 1326 639 1330
rect 660 1325 665 1329
rect 707 1326 711 1330
rect 1524 1325 1528 1329
rect 1568 1326 1572 1330
rect 783 1321 787 1325
rect 864 1321 868 1325
rect 954 1321 958 1325
rect 1593 1325 1598 1329
rect 1640 1326 1644 1330
rect 1716 1321 1720 1325
rect 1797 1321 1801 1325
rect 1887 1321 1891 1325
rect 574 1308 578 1312
rect 606 1307 610 1311
rect 625 1308 629 1312
rect 681 1307 685 1311
rect 697 1308 701 1312
rect 724 1308 728 1312
rect 772 1305 778 1309
rect 853 1305 859 1309
rect 943 1305 949 1309
rect 1507 1308 1511 1312
rect 1539 1307 1543 1311
rect 1558 1308 1562 1312
rect 1614 1307 1618 1311
rect 1630 1308 1634 1312
rect 1657 1308 1661 1312
rect 1705 1305 1711 1309
rect 1786 1305 1792 1309
rect 1876 1305 1882 1309
rect 594 1288 598 1292
rect 638 1288 642 1292
rect 665 1288 669 1292
rect 710 1288 714 1292
rect 781 1285 785 1289
rect 862 1285 866 1289
rect 952 1285 956 1289
rect 1527 1288 1531 1292
rect 1571 1288 1575 1292
rect 1598 1288 1602 1292
rect 1643 1288 1647 1292
rect 1714 1285 1718 1289
rect 1795 1285 1799 1289
rect 1885 1285 1889 1289
rect 783 1267 787 1271
rect 594 1260 598 1264
rect 638 1260 642 1264
rect 665 1260 669 1264
rect 710 1260 714 1264
rect 1716 1267 1720 1271
rect 775 1249 779 1253
rect 574 1240 578 1244
rect 606 1241 610 1245
rect 625 1240 629 1244
rect 681 1241 685 1245
rect 697 1240 701 1244
rect 724 1240 728 1244
rect 802 1245 806 1249
rect 1527 1260 1531 1264
rect 1571 1260 1575 1264
rect 1598 1260 1602 1264
rect 1643 1260 1647 1264
rect 1708 1249 1712 1253
rect 1507 1240 1511 1244
rect 781 1231 785 1235
rect 1539 1241 1543 1245
rect 1558 1240 1562 1244
rect 1614 1241 1618 1245
rect 1630 1240 1634 1244
rect 1657 1240 1661 1244
rect 1735 1245 1739 1249
rect 1714 1231 1718 1235
rect 591 1223 595 1227
rect 635 1222 639 1226
rect 660 1223 665 1227
rect 707 1222 711 1226
rect 1524 1223 1528 1227
rect 1568 1222 1572 1226
rect 1593 1223 1598 1227
rect 1640 1222 1644 1226
rect 106 1205 110 1209
rect 143 1205 147 1209
rect 163 1205 167 1209
rect 201 1205 205 1209
rect 238 1205 242 1209
rect 275 1205 279 1209
rect 295 1205 299 1209
rect 333 1205 337 1209
rect 370 1205 374 1209
rect 407 1205 411 1209
rect 427 1205 431 1209
rect 465 1205 469 1209
rect 1039 1205 1043 1209
rect 1076 1205 1080 1209
rect 1096 1205 1100 1209
rect 1134 1205 1138 1209
rect 1171 1205 1175 1209
rect 1208 1205 1212 1209
rect 1228 1205 1232 1209
rect 1266 1205 1270 1209
rect 1303 1205 1307 1209
rect 1340 1205 1344 1209
rect 1360 1205 1364 1209
rect 1398 1205 1402 1209
rect 100 1185 104 1189
rect 118 1187 122 1191
rect 178 1187 182 1191
rect 136 1178 140 1185
rect 194 1178 198 1185
rect 213 1182 217 1186
rect 231 1187 235 1191
rect 250 1187 254 1191
rect 310 1187 314 1191
rect 268 1178 272 1185
rect 326 1178 330 1185
rect 345 1182 349 1186
rect 363 1187 367 1191
rect 382 1187 386 1191
rect 442 1187 446 1191
rect 400 1178 404 1185
rect 591 1193 595 1197
rect 635 1194 639 1198
rect 660 1193 665 1197
rect 707 1194 711 1198
rect 852 1193 856 1197
rect 896 1194 900 1198
rect 921 1193 926 1197
rect 968 1194 972 1198
rect 458 1178 462 1185
rect 479 1182 483 1186
rect 783 1185 787 1189
rect 1033 1185 1037 1189
rect 1051 1187 1055 1191
rect 574 1176 578 1180
rect 606 1175 610 1179
rect 625 1176 629 1180
rect 681 1175 685 1179
rect 697 1176 701 1180
rect 724 1176 728 1180
rect 106 1164 110 1168
rect 143 1162 147 1166
rect 163 1162 167 1166
rect 199 1162 203 1166
rect 238 1164 242 1168
rect 275 1162 279 1166
rect 295 1162 299 1166
rect 331 1162 335 1166
rect 370 1164 374 1168
rect 407 1162 411 1166
rect 427 1162 431 1166
rect 463 1162 467 1166
rect 772 1169 778 1173
rect 810 1176 814 1180
rect 867 1175 871 1179
rect 886 1176 890 1180
rect 942 1175 946 1179
rect 958 1176 962 1180
rect 985 1176 989 1180
rect 1111 1187 1115 1191
rect 1069 1178 1073 1185
rect 1127 1178 1131 1185
rect 1146 1182 1150 1186
rect 1164 1187 1168 1191
rect 1183 1187 1187 1191
rect 1243 1187 1247 1191
rect 1201 1178 1205 1185
rect 1259 1178 1263 1185
rect 1278 1182 1282 1186
rect 1296 1187 1300 1191
rect 1315 1187 1319 1191
rect 1375 1187 1379 1191
rect 1333 1178 1337 1185
rect 1524 1193 1528 1197
rect 1568 1194 1572 1198
rect 1593 1193 1598 1197
rect 1640 1194 1644 1198
rect 1785 1193 1789 1197
rect 1829 1194 1833 1198
rect 1854 1193 1859 1197
rect 1901 1194 1905 1198
rect 1391 1178 1395 1185
rect 1412 1182 1416 1186
rect 1716 1185 1720 1189
rect 1507 1176 1511 1180
rect 1539 1175 1543 1179
rect 1558 1176 1562 1180
rect 1614 1175 1618 1179
rect 1630 1176 1634 1180
rect 1657 1176 1661 1180
rect 594 1156 598 1160
rect 638 1156 642 1160
rect 665 1156 669 1160
rect 710 1156 714 1160
rect 1039 1164 1043 1168
rect 1076 1162 1080 1166
rect 1096 1162 1100 1166
rect 1132 1162 1136 1166
rect 1171 1164 1175 1168
rect 1208 1162 1212 1166
rect 1228 1162 1232 1166
rect 1264 1162 1268 1166
rect 1303 1164 1307 1168
rect 1340 1162 1344 1166
rect 1360 1162 1364 1166
rect 1396 1162 1400 1166
rect 1705 1169 1711 1173
rect 1743 1176 1747 1180
rect 1800 1175 1804 1179
rect 1819 1176 1823 1180
rect 1875 1175 1879 1179
rect 1891 1176 1895 1180
rect 1918 1176 1922 1180
rect 855 1156 859 1160
rect 899 1156 903 1160
rect 926 1156 930 1160
rect 971 1156 975 1160
rect 1527 1156 1531 1160
rect 1571 1156 1575 1160
rect 1598 1156 1602 1160
rect 1643 1156 1647 1160
rect 1788 1156 1792 1160
rect 1832 1156 1836 1160
rect 1859 1156 1863 1160
rect 1904 1156 1908 1160
rect 781 1149 785 1153
rect 1714 1149 1718 1153
rect 215 1134 219 1138
rect 239 1134 243 1138
rect 1148 1134 1152 1138
rect 1172 1134 1176 1138
rect 994 1128 998 1132
rect 1927 1128 1931 1132
rect 235 1109 239 1113
rect 1168 1109 1172 1113
rect 250 1101 254 1105
rect 1183 1101 1187 1105
rect 877 1095 881 1099
rect 914 1095 918 1099
rect 934 1095 938 1099
rect 972 1095 976 1099
rect 1810 1095 1814 1099
rect 1847 1095 1851 1099
rect 1867 1095 1871 1099
rect 1905 1095 1909 1099
rect 215 1086 219 1090
rect 239 1086 243 1090
rect 1148 1086 1152 1090
rect 1172 1086 1176 1090
rect 871 1075 875 1079
rect 889 1077 893 1081
rect 106 1065 110 1069
rect 143 1065 147 1069
rect 163 1065 167 1069
rect 201 1065 205 1069
rect 238 1065 242 1069
rect 275 1065 279 1069
rect 295 1065 299 1069
rect 333 1065 337 1069
rect 370 1065 374 1069
rect 407 1065 411 1069
rect 427 1065 431 1069
rect 465 1065 469 1069
rect 949 1077 953 1081
rect 907 1068 911 1075
rect 965 1068 969 1075
rect 984 1072 988 1076
rect 1804 1075 1808 1079
rect 1822 1077 1826 1081
rect 1039 1065 1043 1069
rect 1076 1065 1080 1069
rect 1096 1065 1100 1069
rect 1134 1065 1138 1069
rect 1171 1065 1175 1069
rect 1208 1065 1212 1069
rect 1228 1065 1232 1069
rect 1266 1065 1270 1069
rect 1303 1065 1307 1069
rect 1340 1065 1344 1069
rect 1360 1065 1364 1069
rect 1398 1065 1402 1069
rect 1882 1077 1886 1081
rect 1840 1068 1844 1075
rect 1898 1068 1902 1075
rect 1917 1072 1921 1076
rect 877 1054 881 1058
rect 100 1045 104 1049
rect 118 1047 122 1051
rect 178 1047 182 1051
rect 136 1038 140 1045
rect 194 1038 198 1045
rect 213 1042 217 1046
rect 231 1047 235 1051
rect 250 1047 254 1051
rect 310 1047 314 1051
rect 268 1038 272 1045
rect 326 1038 330 1045
rect 345 1042 349 1046
rect 363 1047 367 1051
rect 382 1047 386 1051
rect 442 1047 446 1051
rect 400 1038 404 1045
rect 914 1052 918 1056
rect 934 1052 938 1056
rect 970 1052 974 1056
rect 1810 1054 1814 1058
rect 458 1038 462 1045
rect 479 1042 483 1046
rect 1033 1045 1037 1049
rect 1051 1047 1055 1051
rect 1111 1047 1115 1051
rect 1069 1038 1073 1045
rect 1127 1038 1131 1045
rect 1146 1042 1150 1046
rect 1164 1047 1168 1051
rect 1183 1047 1187 1051
rect 1243 1047 1247 1051
rect 1201 1038 1205 1045
rect 1259 1038 1263 1045
rect 1278 1042 1282 1046
rect 1296 1047 1300 1051
rect 1315 1047 1319 1051
rect 1375 1047 1379 1051
rect 1333 1038 1337 1045
rect 1847 1052 1851 1056
rect 1867 1052 1871 1056
rect 1903 1052 1907 1056
rect 1391 1038 1395 1045
rect 1412 1042 1416 1046
rect 106 1024 110 1028
rect 143 1022 147 1026
rect 163 1022 167 1026
rect 199 1022 203 1026
rect 238 1024 242 1028
rect 275 1022 279 1026
rect 295 1022 299 1026
rect 331 1022 335 1026
rect 370 1024 374 1028
rect 407 1022 411 1026
rect 427 1022 431 1026
rect 463 1022 467 1026
rect 1039 1024 1043 1028
rect 1076 1022 1080 1026
rect 1096 1022 1100 1026
rect 1132 1022 1136 1026
rect 1171 1024 1175 1028
rect 1208 1022 1212 1026
rect 1228 1022 1232 1026
rect 1264 1022 1268 1026
rect 1303 1024 1307 1028
rect 1340 1022 1344 1026
rect 1360 1022 1364 1026
rect 1396 1022 1400 1026
rect 877 1009 881 1013
rect 914 1009 918 1013
rect 934 1009 938 1013
rect 972 1009 976 1013
rect 1810 1009 1814 1013
rect 1847 1009 1851 1013
rect 1867 1009 1871 1013
rect 1905 1009 1909 1013
rect 871 989 875 993
rect 889 991 893 995
rect 106 979 110 983
rect 143 979 147 983
rect 163 979 167 983
rect 201 979 205 983
rect 238 979 242 983
rect 275 979 279 983
rect 295 979 299 983
rect 333 979 337 983
rect 370 979 374 983
rect 407 979 411 983
rect 427 979 431 983
rect 465 979 469 983
rect 949 991 953 995
rect 907 982 911 989
rect 965 982 969 989
rect 984 986 988 990
rect 1006 984 1010 988
rect 1804 989 1808 993
rect 1822 991 1826 995
rect 1039 979 1043 983
rect 1076 979 1080 983
rect 1096 979 1100 983
rect 1134 979 1138 983
rect 1171 979 1175 983
rect 1208 979 1212 983
rect 1228 979 1232 983
rect 1266 979 1270 983
rect 1303 979 1307 983
rect 1340 979 1344 983
rect 1360 979 1364 983
rect 1398 979 1402 983
rect 1882 991 1886 995
rect 1840 982 1844 989
rect 1898 982 1902 989
rect 1917 986 1921 990
rect 1939 984 1943 988
rect 877 968 881 972
rect 100 959 104 963
rect 118 961 122 965
rect 178 961 182 965
rect 136 952 140 959
rect 194 952 198 959
rect 213 956 217 960
rect 231 961 235 965
rect 250 961 254 965
rect 310 961 314 965
rect 268 952 272 959
rect 326 952 330 959
rect 345 956 349 960
rect 363 961 367 965
rect 382 961 386 965
rect 442 961 446 965
rect 400 952 404 959
rect 914 966 918 970
rect 934 966 938 970
rect 970 966 974 970
rect 1810 968 1814 972
rect 458 952 462 959
rect 479 956 483 960
rect 1033 959 1037 963
rect 1051 961 1055 965
rect 1111 961 1115 965
rect 1069 952 1073 959
rect 1127 952 1131 959
rect 1146 956 1150 960
rect 1164 961 1168 965
rect 1183 961 1187 965
rect 1243 961 1247 965
rect 1201 952 1205 959
rect 1259 952 1263 959
rect 1278 956 1282 960
rect 1296 961 1300 965
rect 1315 961 1319 965
rect 1375 961 1379 965
rect 1333 952 1337 959
rect 1847 966 1851 970
rect 1867 966 1871 970
rect 1903 966 1907 970
rect 1391 952 1395 959
rect 1412 956 1416 960
rect 106 938 110 942
rect 143 936 147 940
rect 163 936 167 940
rect 199 936 203 940
rect 238 938 242 942
rect 275 936 279 940
rect 295 936 299 940
rect 331 936 335 940
rect 370 938 374 942
rect 407 936 411 940
rect 427 936 431 940
rect 463 936 467 940
rect 1039 938 1043 942
rect 1076 936 1080 940
rect 1096 936 1100 940
rect 1132 936 1136 940
rect 1171 938 1175 942
rect 1208 936 1212 940
rect 1228 936 1232 940
rect 1264 936 1268 940
rect 1303 938 1307 942
rect 1340 936 1344 940
rect 1360 936 1364 940
rect 1396 936 1400 940
rect 332 908 336 912
rect 356 908 360 912
rect 1265 908 1269 912
rect 1289 908 1293 912
rect 352 883 356 887
rect 1285 883 1289 887
rect 367 875 371 879
rect 1300 875 1304 879
rect 332 860 336 864
rect 356 860 360 864
rect 1265 860 1269 864
rect 1289 860 1293 864
rect 106 839 110 843
rect 143 839 147 843
rect 163 839 167 843
rect 201 839 205 843
rect 238 839 242 843
rect 275 839 279 843
rect 295 839 299 843
rect 333 839 337 843
rect 370 839 374 843
rect 407 839 411 843
rect 427 839 431 843
rect 465 839 469 843
rect 1039 839 1043 843
rect 1076 839 1080 843
rect 1096 839 1100 843
rect 1134 839 1138 843
rect 1171 839 1175 843
rect 1208 839 1212 843
rect 1228 839 1232 843
rect 1266 839 1270 843
rect 1303 839 1307 843
rect 1340 839 1344 843
rect 1360 839 1364 843
rect 1398 839 1402 843
rect 100 819 104 823
rect 118 821 122 825
rect 178 821 182 825
rect 136 812 140 819
rect 194 812 198 819
rect 213 816 217 820
rect 231 821 235 825
rect 250 821 254 825
rect 310 821 314 825
rect 268 812 272 819
rect 326 812 330 819
rect 345 816 349 820
rect 363 821 367 825
rect 382 821 386 825
rect 442 821 446 825
rect 400 812 404 819
rect 458 812 462 819
rect 479 816 483 820
rect 1033 819 1037 823
rect 1051 821 1055 825
rect 1111 821 1115 825
rect 1069 812 1073 819
rect 1127 812 1131 819
rect 1146 816 1150 820
rect 1164 821 1168 825
rect 1183 821 1187 825
rect 1243 821 1247 825
rect 1201 812 1205 819
rect 1259 812 1263 819
rect 1278 816 1282 820
rect 1296 821 1300 825
rect 1315 821 1319 825
rect 1375 821 1379 825
rect 1333 812 1337 819
rect 1391 812 1395 819
rect 1412 816 1416 820
rect 106 798 110 802
rect 143 796 147 800
rect 163 796 167 800
rect 199 796 203 800
rect 238 798 242 802
rect 275 796 279 800
rect 295 796 299 800
rect 331 796 335 800
rect 370 798 374 802
rect 407 796 411 800
rect 427 796 431 800
rect 463 796 467 800
rect 1039 798 1043 802
rect 1076 796 1080 800
rect 1096 796 1100 800
rect 1132 796 1136 800
rect 1171 798 1175 802
rect 1208 796 1212 800
rect 1228 796 1232 800
rect 1264 796 1268 800
rect 1303 798 1307 802
rect 1340 796 1344 800
rect 1360 796 1364 800
rect 1396 796 1400 800
rect 578 760 582 764
rect 615 760 619 764
rect 635 760 639 764
rect 673 760 677 764
rect 710 760 714 764
rect 747 760 751 764
rect 767 760 771 764
rect 805 760 809 764
rect 842 760 846 764
rect 879 760 883 764
rect 899 760 903 764
rect 937 760 941 764
rect 974 760 978 764
rect 1011 760 1015 764
rect 1031 760 1035 764
rect 1069 760 1073 764
rect 1511 760 1515 764
rect 1548 760 1552 764
rect 1568 760 1572 764
rect 1606 760 1610 764
rect 1643 760 1647 764
rect 1680 760 1684 764
rect 1700 760 1704 764
rect 1738 760 1742 764
rect 1775 760 1779 764
rect 1812 760 1816 764
rect 1832 760 1836 764
rect 1870 760 1874 764
rect 1907 760 1911 764
rect 1944 760 1948 764
rect 1964 760 1968 764
rect 2002 760 2006 764
rect 572 740 576 744
rect 590 742 594 746
rect 238 727 242 731
rect 275 727 279 731
rect 295 727 299 731
rect 333 727 337 731
rect 650 742 654 746
rect 608 733 612 740
rect 666 733 670 740
rect 687 737 691 741
rect 704 740 708 744
rect 722 742 726 746
rect 782 742 786 746
rect 740 733 744 740
rect 798 733 802 740
rect 819 737 823 741
rect 836 740 840 744
rect 854 742 858 746
rect 914 742 918 746
rect 872 733 876 740
rect 930 733 934 740
rect 951 737 955 741
rect 968 740 972 744
rect 986 742 990 746
rect 1046 742 1050 746
rect 1004 733 1008 740
rect 1062 733 1066 740
rect 1083 737 1087 741
rect 1505 740 1509 744
rect 1523 742 1527 746
rect 1171 727 1175 731
rect 1208 727 1212 731
rect 1228 727 1232 731
rect 1266 727 1270 731
rect 1583 742 1587 746
rect 1541 733 1545 740
rect 1599 733 1603 740
rect 1620 737 1624 741
rect 1637 740 1641 744
rect 1655 742 1659 746
rect 1715 742 1719 746
rect 1673 733 1677 740
rect 1731 733 1735 740
rect 1752 737 1756 741
rect 1769 740 1773 744
rect 1787 742 1791 746
rect 1847 742 1851 746
rect 1805 733 1809 740
rect 1863 733 1867 740
rect 1884 737 1888 741
rect 1901 740 1905 744
rect 1919 742 1923 746
rect 1979 742 1983 746
rect 1937 733 1941 740
rect 1995 733 1999 740
rect 2016 737 2020 741
rect 578 719 582 723
rect 615 717 619 721
rect 635 717 639 721
rect 671 717 675 721
rect 710 719 714 723
rect 747 717 751 721
rect 767 717 771 721
rect 803 717 807 721
rect 842 719 846 723
rect 879 717 883 721
rect 899 717 903 721
rect 935 717 939 721
rect 974 719 978 723
rect 1011 717 1015 721
rect 1031 717 1035 721
rect 1067 717 1071 721
rect 1511 719 1515 723
rect 1548 717 1552 721
rect 1568 717 1572 721
rect 1604 717 1608 721
rect 1643 719 1647 723
rect 1680 717 1684 721
rect 1700 717 1704 721
rect 1736 717 1740 721
rect 1775 719 1779 723
rect 1812 717 1816 721
rect 1832 717 1836 721
rect 1868 717 1872 721
rect 1907 719 1911 723
rect 1944 717 1948 721
rect 1964 717 1968 721
rect 2000 717 2004 721
rect 232 707 236 711
rect 250 709 254 713
rect 310 709 314 713
rect 268 700 272 707
rect 326 700 330 707
rect 345 704 349 708
rect 1165 707 1169 711
rect 1183 709 1187 713
rect 1243 709 1247 713
rect 1201 700 1205 707
rect 1259 700 1263 707
rect 1278 704 1282 708
rect 238 686 242 690
rect 275 684 279 688
rect 295 684 299 688
rect 331 684 335 688
rect 594 676 598 680
rect 638 676 642 680
rect 665 676 669 680
rect 710 676 714 680
rect 783 683 787 687
rect 356 663 360 667
rect 748 669 752 673
rect 239 654 243 658
rect 574 656 578 660
rect 606 657 610 661
rect 625 656 629 660
rect 681 657 685 661
rect 697 656 701 660
rect 724 656 728 660
rect 864 683 868 687
rect 1171 686 1175 690
rect 775 665 779 669
rect 802 661 806 665
rect 829 669 833 673
rect 1208 684 1212 688
rect 1228 684 1232 688
rect 1264 684 1268 688
rect 856 665 860 669
rect 883 661 887 665
rect 1527 676 1531 680
rect 1571 676 1575 680
rect 1598 676 1602 680
rect 1643 676 1647 680
rect 1716 683 1720 687
rect 1289 663 1293 667
rect 1681 669 1685 673
rect 781 647 785 651
rect 1172 654 1176 658
rect 1507 656 1511 660
rect 862 647 866 651
rect 1539 657 1543 661
rect 1558 656 1562 660
rect 1614 657 1618 661
rect 1630 656 1634 660
rect 1657 656 1661 660
rect 1797 683 1801 687
rect 1708 665 1712 669
rect 1735 661 1739 665
rect 1762 669 1766 673
rect 1789 665 1793 669
rect 1816 661 1820 665
rect 1714 647 1718 651
rect 1795 647 1799 651
rect 591 639 595 643
rect 635 638 639 642
rect 660 639 665 643
rect 707 638 711 642
rect 1524 639 1528 643
rect 1568 638 1572 642
rect 1593 639 1598 643
rect 1640 638 1644 642
rect 238 625 242 629
rect 276 625 280 629
rect 296 625 300 629
rect 333 625 337 629
rect 1171 625 1175 629
rect 1209 625 1213 629
rect 1229 625 1233 629
rect 1266 625 1270 629
rect 226 602 230 606
rect 261 607 265 611
rect 245 598 249 605
rect 303 598 307 605
rect 321 607 325 611
rect 591 609 595 613
rect 635 610 639 614
rect 339 605 343 609
rect 660 609 665 613
rect 707 610 711 614
rect 783 607 787 611
rect 864 607 868 611
rect 574 592 578 596
rect 240 582 244 586
rect 276 582 280 586
rect 296 582 300 586
rect 333 584 337 588
rect 606 591 610 595
rect 625 592 629 596
rect 681 591 685 595
rect 697 592 701 596
rect 724 592 728 596
rect 772 591 778 595
rect 853 591 859 595
rect 1159 602 1163 606
rect 1194 607 1198 611
rect 1178 598 1182 605
rect 1236 598 1240 605
rect 1254 607 1258 611
rect 1524 609 1528 613
rect 1568 610 1572 614
rect 1272 605 1276 609
rect 1593 609 1598 613
rect 1640 610 1644 614
rect 1716 607 1720 611
rect 1797 607 1801 611
rect 1507 592 1511 596
rect 1173 582 1177 586
rect 1209 582 1213 586
rect 1229 582 1233 586
rect 1266 584 1270 588
rect 1539 591 1543 595
rect 1558 592 1562 596
rect 1614 591 1618 595
rect 1630 592 1634 596
rect 1657 592 1661 596
rect 1705 591 1711 595
rect 1786 591 1792 595
rect 594 572 598 576
rect 638 572 642 576
rect 665 572 669 576
rect 710 572 714 576
rect 781 571 785 575
rect 862 571 866 575
rect 1527 572 1531 576
rect 1571 572 1575 576
rect 1598 572 1602 576
rect 1643 572 1647 576
rect 1714 571 1718 575
rect 1795 571 1799 575
rect 783 551 787 555
rect 594 544 598 548
rect 638 544 642 548
rect 665 544 669 548
rect 710 544 714 548
rect 888 551 892 555
rect 775 533 779 537
rect 574 524 578 528
rect 606 525 610 529
rect 625 524 629 528
rect 681 525 685 529
rect 697 524 701 528
rect 724 524 728 528
rect 802 529 806 533
rect 853 537 857 541
rect 1716 551 1720 555
rect 880 533 884 537
rect 907 529 911 533
rect 1527 544 1531 548
rect 1571 544 1575 548
rect 1598 544 1602 548
rect 1643 544 1647 548
rect 1821 551 1825 555
rect 1708 533 1712 537
rect 1507 524 1511 528
rect 781 515 785 519
rect 886 515 890 519
rect 1539 525 1543 529
rect 1558 524 1562 528
rect 1614 525 1618 529
rect 1630 524 1634 528
rect 1657 524 1661 528
rect 1735 529 1739 533
rect 1786 537 1790 541
rect 1813 533 1817 537
rect 1840 529 1844 533
rect 1714 515 1718 519
rect 1819 515 1823 519
rect 591 507 595 511
rect 635 506 639 510
rect 660 507 665 511
rect 707 506 711 510
rect 1524 507 1528 511
rect 1568 506 1572 510
rect 1593 507 1598 511
rect 1640 506 1644 510
rect 591 477 595 481
rect 635 478 639 482
rect 660 477 665 481
rect 707 478 711 482
rect 783 476 787 480
rect 888 476 892 480
rect 1524 477 1528 481
rect 1568 478 1572 482
rect 1593 477 1598 481
rect 1640 478 1644 482
rect 1716 476 1720 480
rect 1821 476 1825 480
rect 574 460 578 464
rect 606 459 610 463
rect 625 460 629 464
rect 681 459 685 463
rect 697 460 701 464
rect 724 460 728 464
rect 772 460 778 464
rect 877 460 883 464
rect 1507 460 1511 464
rect 1539 459 1543 463
rect 1558 460 1562 464
rect 1614 459 1618 463
rect 1630 460 1634 464
rect 1657 460 1661 464
rect 1705 460 1711 464
rect 1810 460 1816 464
rect 594 440 598 444
rect 638 440 642 444
rect 665 440 669 444
rect 710 440 714 444
rect 781 440 785 444
rect 886 440 890 444
rect 1527 440 1531 444
rect 1571 440 1575 444
rect 1598 440 1602 444
rect 1643 440 1647 444
rect 1714 440 1718 444
rect 1819 440 1823 444
rect 783 419 787 423
rect 594 412 598 416
rect 638 412 642 416
rect 665 412 669 416
rect 710 412 714 416
rect 864 419 868 423
rect 775 401 779 405
rect 574 392 578 396
rect 606 393 610 397
rect 625 392 629 396
rect 681 393 685 397
rect 697 392 701 396
rect 724 392 728 396
rect 802 397 806 401
rect 829 405 833 409
rect 954 419 958 423
rect 856 401 860 405
rect 883 397 887 401
rect 919 405 923 409
rect 1716 419 1720 423
rect 946 401 950 405
rect 973 397 977 401
rect 1527 412 1531 416
rect 1571 412 1575 416
rect 1598 412 1602 416
rect 1643 412 1647 416
rect 1797 419 1801 423
rect 1708 401 1712 405
rect 1507 392 1511 396
rect 781 383 785 387
rect 862 383 866 387
rect 952 383 956 387
rect 1539 393 1543 397
rect 1558 392 1562 396
rect 1614 393 1618 397
rect 1630 392 1634 396
rect 1657 392 1661 396
rect 1735 397 1739 401
rect 1762 405 1766 409
rect 1887 419 1891 423
rect 1789 401 1793 405
rect 1816 397 1820 401
rect 1852 405 1856 409
rect 1879 401 1883 405
rect 1906 397 1910 401
rect 1714 383 1718 387
rect 1795 383 1799 387
rect 1885 383 1889 387
rect 591 375 595 379
rect 635 374 639 378
rect 660 375 665 379
rect 707 374 711 378
rect 1524 375 1528 379
rect 1568 374 1572 378
rect 1593 375 1598 379
rect 1640 374 1644 378
rect 591 345 595 349
rect 635 346 639 350
rect 660 345 665 349
rect 707 346 711 350
rect 1524 345 1528 349
rect 1568 346 1572 350
rect 783 341 787 345
rect 864 341 868 345
rect 954 341 958 345
rect 1593 345 1598 349
rect 1640 346 1644 350
rect 1716 341 1720 345
rect 1797 341 1801 345
rect 1887 341 1891 345
rect 574 328 578 332
rect 606 327 610 331
rect 625 328 629 332
rect 681 327 685 331
rect 697 328 701 332
rect 724 328 728 332
rect 772 325 778 329
rect 853 325 859 329
rect 943 325 949 329
rect 1507 328 1511 332
rect 1539 327 1543 331
rect 1558 328 1562 332
rect 1614 327 1618 331
rect 1630 328 1634 332
rect 1657 328 1661 332
rect 1705 325 1711 329
rect 1786 325 1792 329
rect 1876 325 1882 329
rect 594 308 598 312
rect 638 308 642 312
rect 665 308 669 312
rect 710 308 714 312
rect 781 305 785 309
rect 862 305 866 309
rect 952 305 956 309
rect 1527 308 1531 312
rect 1571 308 1575 312
rect 1598 308 1602 312
rect 1643 308 1647 312
rect 1714 305 1718 309
rect 1795 305 1799 309
rect 1885 305 1889 309
rect 783 287 787 291
rect 594 280 598 284
rect 638 280 642 284
rect 665 280 669 284
rect 710 280 714 284
rect 1716 287 1720 291
rect 775 269 779 273
rect 574 260 578 264
rect 606 261 610 265
rect 625 260 629 264
rect 681 261 685 265
rect 697 260 701 264
rect 724 260 728 264
rect 802 265 806 269
rect 1527 280 1531 284
rect 1571 280 1575 284
rect 1598 280 1602 284
rect 1643 280 1647 284
rect 1708 269 1712 273
rect 1507 260 1511 264
rect 781 251 785 255
rect 1539 261 1543 265
rect 1558 260 1562 264
rect 1614 261 1618 265
rect 1630 260 1634 264
rect 1657 260 1661 264
rect 1735 265 1739 269
rect 1714 251 1718 255
rect 591 243 595 247
rect 635 242 639 246
rect 660 243 665 247
rect 707 242 711 246
rect 1524 243 1528 247
rect 1568 242 1572 246
rect 1593 243 1598 247
rect 1640 242 1644 246
rect 106 225 110 229
rect 143 225 147 229
rect 163 225 167 229
rect 201 225 205 229
rect 238 225 242 229
rect 275 225 279 229
rect 295 225 299 229
rect 333 225 337 229
rect 370 225 374 229
rect 407 225 411 229
rect 427 225 431 229
rect 465 225 469 229
rect 1039 225 1043 229
rect 1076 225 1080 229
rect 1096 225 1100 229
rect 1134 225 1138 229
rect 1171 225 1175 229
rect 1208 225 1212 229
rect 1228 225 1232 229
rect 1266 225 1270 229
rect 1303 225 1307 229
rect 1340 225 1344 229
rect 1360 225 1364 229
rect 1398 225 1402 229
rect 100 205 104 209
rect 118 207 122 211
rect 178 207 182 211
rect 136 198 140 205
rect 194 198 198 205
rect 213 202 217 206
rect 231 207 235 211
rect 250 207 254 211
rect 310 207 314 211
rect 268 198 272 205
rect 326 198 330 205
rect 345 202 349 206
rect 363 207 367 211
rect 382 207 386 211
rect 442 207 446 211
rect 400 198 404 205
rect 591 213 595 217
rect 635 214 639 218
rect 660 213 665 217
rect 707 214 711 218
rect 852 213 856 217
rect 896 214 900 218
rect 921 213 926 217
rect 968 214 972 218
rect 458 198 462 205
rect 479 202 483 206
rect 783 205 787 209
rect 1033 205 1037 209
rect 1051 207 1055 211
rect 574 196 578 200
rect 606 195 610 199
rect 625 196 629 200
rect 681 195 685 199
rect 697 196 701 200
rect 724 196 728 200
rect 106 184 110 188
rect 143 182 147 186
rect 163 182 167 186
rect 199 182 203 186
rect 238 184 242 188
rect 275 182 279 186
rect 295 182 299 186
rect 331 182 335 186
rect 370 184 374 188
rect 407 182 411 186
rect 427 182 431 186
rect 463 182 467 186
rect 772 189 778 193
rect 810 196 814 200
rect 867 195 871 199
rect 886 196 890 200
rect 942 195 946 199
rect 958 196 962 200
rect 985 196 989 200
rect 1111 207 1115 211
rect 1069 198 1073 205
rect 1127 198 1131 205
rect 1146 202 1150 206
rect 1164 207 1168 211
rect 1183 207 1187 211
rect 1243 207 1247 211
rect 1201 198 1205 205
rect 1259 198 1263 205
rect 1278 202 1282 206
rect 1296 207 1300 211
rect 1315 207 1319 211
rect 1375 207 1379 211
rect 1333 198 1337 205
rect 1524 213 1528 217
rect 1568 214 1572 218
rect 1593 213 1598 217
rect 1640 214 1644 218
rect 1785 213 1789 217
rect 1829 214 1833 218
rect 1854 213 1859 217
rect 1901 214 1905 218
rect 1391 198 1395 205
rect 1412 202 1416 206
rect 1716 205 1720 209
rect 1507 196 1511 200
rect 1539 195 1543 199
rect 1558 196 1562 200
rect 1614 195 1618 199
rect 1630 196 1634 200
rect 1657 196 1661 200
rect 594 176 598 180
rect 638 176 642 180
rect 665 176 669 180
rect 710 176 714 180
rect 1039 184 1043 188
rect 1076 182 1080 186
rect 1096 182 1100 186
rect 1132 182 1136 186
rect 1171 184 1175 188
rect 1208 182 1212 186
rect 1228 182 1232 186
rect 1264 182 1268 186
rect 1303 184 1307 188
rect 1340 182 1344 186
rect 1360 182 1364 186
rect 1396 182 1400 186
rect 1705 189 1711 193
rect 1743 196 1747 200
rect 1800 195 1804 199
rect 1819 196 1823 200
rect 1875 195 1879 199
rect 1891 196 1895 200
rect 1918 196 1922 200
rect 855 176 859 180
rect 899 176 903 180
rect 926 176 930 180
rect 971 176 975 180
rect 1527 176 1531 180
rect 1571 176 1575 180
rect 1598 176 1602 180
rect 1643 176 1647 180
rect 1788 176 1792 180
rect 1832 176 1836 180
rect 1859 176 1863 180
rect 1904 176 1908 180
rect 781 169 785 173
rect 1714 169 1718 173
rect 215 154 219 158
rect 239 154 243 158
rect 1148 154 1152 158
rect 1172 154 1176 158
rect 994 148 998 152
rect 1927 148 1931 152
rect 235 129 239 133
rect 1168 129 1172 133
rect 250 121 254 125
rect 1183 121 1187 125
rect 877 115 881 119
rect 914 115 918 119
rect 934 115 938 119
rect 972 115 976 119
rect 1810 115 1814 119
rect 1847 115 1851 119
rect 1867 115 1871 119
rect 1905 115 1909 119
rect 215 106 219 110
rect 239 106 243 110
rect 1148 106 1152 110
rect 1172 106 1176 110
rect 871 95 875 99
rect 889 97 893 101
rect 106 85 110 89
rect 143 85 147 89
rect 163 85 167 89
rect 201 85 205 89
rect 238 85 242 89
rect 275 85 279 89
rect 295 85 299 89
rect 333 85 337 89
rect 370 85 374 89
rect 407 85 411 89
rect 427 85 431 89
rect 465 85 469 89
rect 949 97 953 101
rect 907 88 911 95
rect 965 88 969 95
rect 984 92 988 96
rect 1804 95 1808 99
rect 1822 97 1826 101
rect 1039 85 1043 89
rect 1076 85 1080 89
rect 1096 85 1100 89
rect 1134 85 1138 89
rect 1171 85 1175 89
rect 1208 85 1212 89
rect 1228 85 1232 89
rect 1266 85 1270 89
rect 1303 85 1307 89
rect 1340 85 1344 89
rect 1360 85 1364 89
rect 1398 85 1402 89
rect 1882 97 1886 101
rect 1840 88 1844 95
rect 1898 88 1902 95
rect 1917 92 1921 96
rect 877 74 881 78
rect 100 65 104 69
rect 118 67 122 71
rect 178 67 182 71
rect 136 58 140 65
rect 194 58 198 65
rect 213 62 217 66
rect 231 67 235 71
rect 250 67 254 71
rect 310 67 314 71
rect 268 58 272 65
rect 326 58 330 65
rect 345 62 349 66
rect 363 67 367 71
rect 382 67 386 71
rect 442 67 446 71
rect 400 58 404 65
rect 914 72 918 76
rect 934 72 938 76
rect 970 72 974 76
rect 1810 74 1814 78
rect 458 58 462 65
rect 479 62 483 66
rect 1033 65 1037 69
rect 1051 67 1055 71
rect 1111 67 1115 71
rect 1069 58 1073 65
rect 1127 58 1131 65
rect 1146 62 1150 66
rect 1164 67 1168 71
rect 1183 67 1187 71
rect 1243 67 1247 71
rect 1201 58 1205 65
rect 1259 58 1263 65
rect 1278 62 1282 66
rect 1296 67 1300 71
rect 1315 67 1319 71
rect 1375 67 1379 71
rect 1333 58 1337 65
rect 1847 72 1851 76
rect 1867 72 1871 76
rect 1903 72 1907 76
rect 1391 58 1395 65
rect 1412 62 1416 66
rect 106 44 110 48
rect 143 42 147 46
rect 163 42 167 46
rect 199 42 203 46
rect 238 44 242 48
rect 275 42 279 46
rect 295 42 299 46
rect 331 42 335 46
rect 370 44 374 48
rect 407 42 411 46
rect 427 42 431 46
rect 463 42 467 46
rect 1039 44 1043 48
rect 1076 42 1080 46
rect 1096 42 1100 46
rect 1132 42 1136 46
rect 1171 44 1175 48
rect 1208 42 1212 46
rect 1228 42 1232 46
rect 1264 42 1268 46
rect 1303 44 1307 48
rect 1340 42 1344 46
rect 1360 42 1364 46
rect 1396 42 1400 46
rect 877 29 881 33
rect 914 29 918 33
rect 934 29 938 33
rect 972 29 976 33
rect 1810 29 1814 33
rect 1847 29 1851 33
rect 1867 29 1871 33
rect 1905 29 1909 33
rect 871 9 875 13
rect 889 11 893 15
rect 106 -1 110 3
rect 143 -1 147 3
rect 163 -1 167 3
rect 201 -1 205 3
rect 238 -1 242 3
rect 275 -1 279 3
rect 295 -1 299 3
rect 333 -1 337 3
rect 370 -1 374 3
rect 407 -1 411 3
rect 427 -1 431 3
rect 465 -1 469 3
rect 949 11 953 15
rect 907 2 911 9
rect 965 2 969 9
rect 984 6 988 10
rect 1006 4 1010 8
rect 1804 9 1808 13
rect 1822 11 1826 15
rect 1039 -1 1043 3
rect 1076 -1 1080 3
rect 1096 -1 1100 3
rect 1134 -1 1138 3
rect 1171 -1 1175 3
rect 1208 -1 1212 3
rect 1228 -1 1232 3
rect 1266 -1 1270 3
rect 1303 -1 1307 3
rect 1340 -1 1344 3
rect 1360 -1 1364 3
rect 1398 -1 1402 3
rect 1882 11 1886 15
rect 1840 2 1844 9
rect 1898 2 1902 9
rect 1917 6 1921 10
rect 1939 4 1943 8
rect 877 -12 881 -8
rect 100 -21 104 -17
rect 118 -19 122 -15
rect 178 -19 182 -15
rect 136 -28 140 -21
rect 194 -28 198 -21
rect 213 -24 217 -20
rect 231 -19 235 -15
rect 250 -19 254 -15
rect 310 -19 314 -15
rect 268 -28 272 -21
rect 326 -28 330 -21
rect 345 -24 349 -20
rect 363 -19 367 -15
rect 382 -19 386 -15
rect 442 -19 446 -15
rect 400 -28 404 -21
rect 914 -14 918 -10
rect 934 -14 938 -10
rect 970 -14 974 -10
rect 1810 -12 1814 -8
rect 458 -28 462 -21
rect 479 -24 483 -20
rect 1033 -21 1037 -17
rect 1051 -19 1055 -15
rect 1111 -19 1115 -15
rect 1069 -28 1073 -21
rect 1127 -28 1131 -21
rect 1146 -24 1150 -20
rect 1164 -19 1168 -15
rect 1183 -19 1187 -15
rect 1243 -19 1247 -15
rect 1201 -28 1205 -21
rect 1259 -28 1263 -21
rect 1278 -24 1282 -20
rect 1296 -19 1300 -15
rect 1315 -19 1319 -15
rect 1375 -19 1379 -15
rect 1333 -28 1337 -21
rect 1847 -14 1851 -10
rect 1867 -14 1871 -10
rect 1903 -14 1907 -10
rect 1391 -28 1395 -21
rect 1412 -24 1416 -20
rect 106 -42 110 -38
rect 143 -44 147 -40
rect 163 -44 167 -40
rect 199 -44 203 -40
rect 238 -42 242 -38
rect 275 -44 279 -40
rect 295 -44 299 -40
rect 331 -44 335 -40
rect 370 -42 374 -38
rect 407 -44 411 -40
rect 427 -44 431 -40
rect 463 -44 467 -40
rect 1039 -42 1043 -38
rect 1076 -44 1080 -40
rect 1096 -44 1100 -40
rect 1132 -44 1136 -40
rect 1171 -42 1175 -38
rect 1208 -44 1212 -40
rect 1228 -44 1232 -40
rect 1264 -44 1268 -40
rect 1303 -42 1307 -38
rect 1340 -44 1344 -40
rect 1360 -44 1364 -40
rect 1396 -44 1400 -40
rect 332 -72 336 -68
rect 356 -72 360 -68
rect 1265 -72 1269 -68
rect 1289 -72 1293 -68
rect 352 -97 356 -93
rect 1285 -97 1289 -93
rect 367 -105 371 -101
rect 1300 -105 1304 -101
rect 332 -120 336 -116
rect 356 -120 360 -116
rect 1265 -120 1269 -116
rect 1289 -120 1293 -116
rect 106 -141 110 -137
rect 143 -141 147 -137
rect 163 -141 167 -137
rect 201 -141 205 -137
rect 238 -141 242 -137
rect 275 -141 279 -137
rect 295 -141 299 -137
rect 333 -141 337 -137
rect 370 -141 374 -137
rect 407 -141 411 -137
rect 427 -141 431 -137
rect 465 -141 469 -137
rect 1039 -141 1043 -137
rect 1076 -141 1080 -137
rect 1096 -141 1100 -137
rect 1134 -141 1138 -137
rect 1171 -141 1175 -137
rect 1208 -141 1212 -137
rect 1228 -141 1232 -137
rect 1266 -141 1270 -137
rect 1303 -141 1307 -137
rect 1340 -141 1344 -137
rect 1360 -141 1364 -137
rect 1398 -141 1402 -137
rect 100 -161 104 -157
rect 118 -159 122 -155
rect 178 -159 182 -155
rect 136 -168 140 -161
rect 194 -168 198 -161
rect 213 -164 217 -160
rect 231 -159 235 -155
rect 250 -159 254 -155
rect 310 -159 314 -155
rect 268 -168 272 -161
rect 326 -168 330 -161
rect 345 -164 349 -160
rect 363 -159 367 -155
rect 382 -159 386 -155
rect 442 -159 446 -155
rect 400 -168 404 -161
rect 458 -168 462 -161
rect 479 -164 483 -160
rect 1033 -161 1037 -157
rect 1051 -159 1055 -155
rect 1111 -159 1115 -155
rect 1069 -168 1073 -161
rect 1127 -168 1131 -161
rect 1146 -164 1150 -160
rect 1164 -159 1168 -155
rect 1183 -159 1187 -155
rect 1243 -159 1247 -155
rect 1201 -168 1205 -161
rect 1259 -168 1263 -161
rect 1278 -164 1282 -160
rect 1296 -159 1300 -155
rect 1315 -159 1319 -155
rect 1375 -159 1379 -155
rect 1333 -168 1337 -161
rect 1391 -168 1395 -161
rect 1412 -164 1416 -160
rect 106 -182 110 -178
rect 143 -184 147 -180
rect 163 -184 167 -180
rect 199 -184 203 -180
rect 238 -182 242 -178
rect 275 -184 279 -180
rect 295 -184 299 -180
rect 331 -184 335 -180
rect 370 -182 374 -178
rect 407 -184 411 -180
rect 427 -184 431 -180
rect 463 -184 467 -180
rect 1039 -182 1043 -178
rect 1076 -184 1080 -180
rect 1096 -184 1100 -180
rect 1132 -184 1136 -180
rect 1171 -182 1175 -178
rect 1208 -184 1212 -180
rect 1228 -184 1232 -180
rect 1264 -184 1268 -180
rect 1303 -182 1307 -178
rect 1340 -184 1344 -180
rect 1360 -184 1364 -180
rect 1396 -184 1400 -180
<< metal1 >>
rect 559 1754 574 1758
rect 578 1754 610 1758
rect 614 1754 677 1758
rect 681 1754 706 1758
rect 710 1754 742 1758
rect 746 1754 809 1758
rect 813 1754 838 1758
rect 842 1754 874 1758
rect 878 1754 941 1758
rect 945 1754 970 1758
rect 974 1754 1006 1758
rect 1010 1754 1073 1758
rect 1077 1754 1093 1758
rect 1492 1754 1507 1758
rect 1511 1754 1543 1758
rect 1547 1754 1610 1758
rect 1614 1754 1639 1758
rect 1643 1754 1675 1758
rect 1679 1754 1742 1758
rect 1746 1754 1771 1758
rect 1775 1754 1807 1758
rect 1811 1754 1874 1758
rect 1878 1754 1903 1758
rect 1907 1754 1939 1758
rect 1943 1754 2006 1758
rect 2010 1754 2026 1758
rect 499 1747 598 1751
rect 602 1747 626 1751
rect 630 1747 656 1751
rect 660 1747 693 1751
rect 697 1747 730 1751
rect 734 1747 758 1751
rect 762 1747 788 1751
rect 792 1747 825 1751
rect 829 1747 862 1751
rect 866 1747 890 1751
rect 894 1747 920 1751
rect 924 1747 957 1751
rect 961 1747 994 1751
rect 998 1747 1022 1751
rect 1026 1747 1052 1751
rect 1056 1747 1089 1751
rect 1432 1747 1531 1751
rect 1535 1747 1559 1751
rect 1563 1747 1589 1751
rect 1593 1747 1626 1751
rect 1630 1747 1663 1751
rect 1667 1747 1691 1751
rect 1695 1747 1721 1751
rect 1725 1747 1758 1751
rect 1762 1747 1795 1751
rect 1799 1747 1823 1751
rect 1827 1747 1853 1751
rect 1857 1747 1890 1751
rect 1894 1747 1927 1751
rect 1931 1747 1955 1751
rect 1959 1747 1985 1751
rect 1989 1747 2022 1751
rect 568 1737 571 1747
rect 589 1737 592 1747
rect 605 1737 608 1747
rect 619 1740 624 1744
rect 628 1740 635 1744
rect 647 1737 650 1747
rect 663 1737 666 1747
rect 684 1737 687 1747
rect 700 1737 703 1747
rect 721 1737 724 1747
rect 737 1737 740 1747
rect 751 1740 756 1744
rect 760 1740 767 1744
rect 779 1737 782 1747
rect 795 1737 798 1747
rect 816 1737 819 1747
rect 832 1737 835 1747
rect 853 1737 856 1747
rect 869 1737 872 1747
rect 883 1740 888 1744
rect 892 1740 899 1744
rect 911 1737 914 1747
rect 927 1737 930 1747
rect 948 1737 951 1747
rect 964 1737 967 1747
rect 985 1737 988 1747
rect 1001 1737 1004 1747
rect 1015 1740 1020 1744
rect 1024 1740 1031 1744
rect 1043 1737 1046 1747
rect 1059 1737 1062 1747
rect 1080 1737 1083 1747
rect 1501 1737 1504 1747
rect 1522 1737 1525 1747
rect 1538 1737 1541 1747
rect 1552 1740 1557 1744
rect 1561 1740 1568 1744
rect 1580 1737 1583 1747
rect 1596 1737 1599 1747
rect 1617 1737 1620 1747
rect 1633 1737 1636 1747
rect 1654 1737 1657 1747
rect 1670 1737 1673 1747
rect 1684 1740 1689 1744
rect 1693 1740 1700 1744
rect 1712 1737 1715 1747
rect 1728 1737 1731 1747
rect 1749 1737 1752 1747
rect 1765 1737 1768 1747
rect 1786 1737 1789 1747
rect 1802 1737 1805 1747
rect 1816 1740 1821 1744
rect 1825 1740 1832 1744
rect 1844 1737 1847 1747
rect 1860 1737 1863 1747
rect 1881 1737 1884 1747
rect 1897 1737 1900 1747
rect 1918 1737 1921 1747
rect 1934 1737 1937 1747
rect 1948 1740 1953 1744
rect 1957 1740 1964 1744
rect 1976 1737 1979 1747
rect 1992 1737 1995 1747
rect 2013 1737 2016 1747
rect 225 1721 234 1725
rect 238 1721 270 1725
rect 274 1721 337 1725
rect 341 1721 553 1725
rect 585 1723 590 1726
rect 594 1723 618 1726
rect 643 1723 650 1726
rect 654 1723 676 1726
rect 225 1714 258 1718
rect 262 1714 286 1718
rect 290 1714 316 1718
rect 320 1714 353 1718
rect 357 1714 493 1718
rect 228 1704 231 1714
rect 249 1704 252 1714
rect 265 1704 268 1714
rect 279 1707 284 1711
rect 288 1707 295 1711
rect 307 1704 310 1714
rect 323 1704 326 1714
rect 344 1704 347 1714
rect 601 1713 608 1716
rect 612 1717 631 1720
rect 631 1710 634 1716
rect 659 1713 666 1716
rect 670 1717 687 1720
rect 717 1723 722 1726
rect 726 1723 750 1726
rect 775 1723 782 1726
rect 786 1723 808 1726
rect 733 1713 740 1716
rect 744 1717 763 1720
rect 763 1710 766 1716
rect 791 1713 798 1716
rect 802 1717 819 1720
rect 849 1723 854 1726
rect 858 1723 882 1726
rect 907 1723 914 1726
rect 918 1723 940 1726
rect 865 1713 872 1716
rect 876 1717 895 1720
rect 895 1710 898 1716
rect 923 1713 930 1716
rect 934 1717 951 1720
rect 981 1723 986 1726
rect 990 1723 1014 1726
rect 1039 1723 1046 1726
rect 1050 1723 1072 1726
rect 1158 1721 1167 1725
rect 1171 1721 1203 1725
rect 1207 1721 1270 1725
rect 1274 1721 1486 1725
rect 997 1713 1004 1716
rect 1008 1717 1027 1720
rect 223 1687 232 1691
rect 245 1690 250 1693
rect 254 1690 278 1693
rect 303 1690 310 1693
rect 314 1690 336 1693
rect 568 1694 571 1706
rect 589 1694 592 1706
rect 605 1694 608 1706
rect 619 1697 631 1700
rect 647 1694 650 1706
rect 663 1694 666 1706
rect 684 1694 687 1706
rect 700 1694 703 1706
rect 721 1694 724 1706
rect 737 1694 740 1706
rect 751 1697 763 1700
rect 779 1694 782 1706
rect 795 1694 798 1706
rect 816 1694 819 1706
rect 832 1694 835 1706
rect 853 1694 856 1706
rect 869 1694 872 1706
rect 883 1697 895 1700
rect 911 1694 914 1706
rect 927 1694 930 1706
rect 948 1694 951 1706
rect 1027 1710 1030 1716
rect 1055 1713 1062 1716
rect 1066 1717 1083 1720
rect 1518 1723 1523 1726
rect 1527 1723 1551 1726
rect 1576 1723 1583 1726
rect 1587 1723 1609 1726
rect 1158 1714 1191 1718
rect 1195 1714 1219 1718
rect 1223 1714 1249 1718
rect 1253 1714 1286 1718
rect 1290 1714 1426 1718
rect 964 1694 967 1706
rect 985 1694 988 1706
rect 1001 1694 1004 1706
rect 1015 1697 1027 1700
rect 1043 1694 1046 1706
rect 1059 1694 1062 1706
rect 1080 1694 1083 1706
rect 1161 1704 1164 1714
rect 1182 1704 1185 1714
rect 1198 1704 1201 1714
rect 1212 1707 1217 1711
rect 1221 1707 1228 1711
rect 1240 1704 1243 1714
rect 1256 1704 1259 1714
rect 1277 1704 1280 1714
rect 1534 1713 1541 1716
rect 1545 1717 1564 1720
rect 1564 1710 1567 1716
rect 1592 1713 1599 1716
rect 1603 1717 1620 1720
rect 1650 1723 1655 1726
rect 1659 1723 1683 1726
rect 1708 1723 1715 1726
rect 1719 1723 1741 1726
rect 1666 1713 1673 1716
rect 1677 1717 1696 1720
rect 1696 1710 1699 1716
rect 1724 1713 1731 1716
rect 1735 1717 1752 1720
rect 1782 1723 1787 1726
rect 1791 1723 1815 1726
rect 1840 1723 1847 1726
rect 1851 1723 1873 1726
rect 1798 1713 1805 1716
rect 1809 1717 1828 1720
rect 1828 1710 1831 1716
rect 1856 1713 1863 1716
rect 1867 1717 1884 1720
rect 1914 1723 1919 1726
rect 1923 1723 1947 1726
rect 1972 1723 1979 1726
rect 1983 1723 2005 1726
rect 1930 1713 1937 1716
rect 1941 1717 1960 1720
rect 511 1690 598 1694
rect 602 1690 626 1694
rect 630 1690 656 1694
rect 660 1690 730 1694
rect 734 1690 758 1694
rect 762 1690 788 1694
rect 792 1690 862 1694
rect 866 1690 890 1694
rect 894 1690 920 1694
rect 924 1690 994 1694
rect 998 1690 1022 1694
rect 1026 1690 1052 1694
rect 1056 1690 1093 1694
rect 261 1680 268 1683
rect 272 1684 291 1687
rect 291 1677 294 1683
rect 319 1680 326 1683
rect 330 1684 345 1687
rect 1156 1687 1165 1691
rect 1178 1690 1183 1693
rect 1187 1690 1211 1693
rect 1236 1690 1243 1693
rect 1247 1690 1269 1693
rect 1501 1694 1504 1706
rect 1522 1694 1525 1706
rect 1538 1694 1541 1706
rect 1552 1697 1564 1700
rect 1580 1694 1583 1706
rect 1596 1694 1599 1706
rect 1617 1694 1620 1706
rect 1633 1694 1636 1706
rect 1654 1694 1657 1706
rect 1670 1694 1673 1706
rect 1684 1697 1696 1700
rect 1712 1694 1715 1706
rect 1728 1694 1731 1706
rect 1749 1694 1752 1706
rect 1765 1694 1768 1706
rect 1786 1694 1789 1706
rect 1802 1694 1805 1706
rect 1816 1697 1828 1700
rect 1844 1694 1847 1706
rect 1860 1694 1863 1706
rect 1881 1694 1884 1706
rect 1960 1710 1963 1716
rect 1988 1713 1995 1716
rect 1999 1717 2016 1720
rect 1897 1694 1900 1706
rect 1918 1694 1921 1706
rect 1934 1694 1937 1706
rect 1948 1697 1960 1700
rect 1976 1694 1979 1706
rect 1992 1694 1995 1706
rect 2013 1694 2016 1706
rect 1444 1690 1531 1694
rect 1535 1690 1559 1694
rect 1563 1690 1589 1694
rect 1593 1690 1663 1694
rect 1667 1690 1691 1694
rect 1695 1690 1721 1694
rect 1725 1690 1795 1694
rect 1799 1690 1823 1694
rect 1827 1690 1853 1694
rect 1857 1690 1927 1694
rect 1931 1690 1955 1694
rect 1959 1690 1985 1694
rect 1989 1690 2026 1694
rect 547 1683 574 1687
rect 578 1683 625 1687
rect 629 1683 675 1687
rect 679 1683 706 1687
rect 710 1683 757 1687
rect 761 1683 807 1687
rect 811 1683 838 1687
rect 842 1683 889 1687
rect 893 1683 939 1687
rect 943 1683 970 1687
rect 974 1683 1021 1687
rect 1025 1683 1071 1687
rect 1075 1683 1093 1687
rect 1194 1680 1201 1683
rect 1205 1684 1224 1687
rect 228 1661 231 1673
rect 249 1661 252 1673
rect 265 1661 268 1673
rect 279 1664 291 1667
rect 307 1661 310 1673
rect 323 1661 326 1673
rect 344 1661 347 1673
rect 499 1670 572 1674
rect 576 1670 588 1674
rect 592 1670 606 1674
rect 610 1670 617 1674
rect 621 1670 623 1674
rect 627 1670 642 1674
rect 646 1670 679 1674
rect 683 1670 684 1674
rect 688 1670 696 1674
rect 700 1670 724 1674
rect 728 1670 740 1674
rect 744 1670 764 1674
rect 768 1670 818 1674
rect 822 1670 845 1674
rect 849 1670 899 1674
rect 903 1670 922 1674
rect 1224 1677 1227 1683
rect 1252 1680 1259 1683
rect 1263 1684 1278 1687
rect 1480 1683 1507 1687
rect 1511 1683 1558 1687
rect 1562 1683 1608 1687
rect 1612 1683 1639 1687
rect 1643 1683 1690 1687
rect 1694 1683 1740 1687
rect 1744 1683 1771 1687
rect 1775 1683 1822 1687
rect 1826 1683 1872 1687
rect 1876 1683 1903 1687
rect 1907 1683 1954 1687
rect 1958 1683 2004 1687
rect 2008 1683 2026 1687
rect 535 1663 599 1667
rect 603 1663 630 1667
rect 634 1663 652 1667
rect 656 1663 717 1667
rect 721 1663 735 1667
rect 747 1666 750 1670
rect 225 1657 258 1661
rect 262 1657 286 1661
rect 290 1657 316 1661
rect 320 1657 505 1661
rect 225 1650 234 1654
rect 238 1650 285 1654
rect 289 1650 335 1654
rect 339 1650 541 1654
rect 642 1656 645 1660
rect 669 1656 670 1660
rect 714 1656 716 1660
rect 756 1653 759 1658
rect 771 1660 774 1670
rect 801 1666 804 1670
rect 828 1666 831 1670
rect 223 1634 239 1638
rect 348 1636 352 1640
rect 364 1636 368 1640
rect 372 1636 574 1640
rect 582 1639 585 1645
rect 589 1639 592 1645
rect 582 1636 592 1639
rect 582 1631 585 1636
rect 231 1627 235 1631
rect 247 1627 368 1631
rect 589 1631 592 1636
rect 598 1641 601 1645
rect 598 1637 600 1641
rect 604 1637 606 1641
rect 614 1640 617 1645
rect 642 1642 645 1645
rect 614 1638 625 1640
rect 598 1631 601 1637
rect 614 1636 620 1638
rect 614 1631 617 1636
rect 624 1636 625 1638
rect 643 1638 645 1642
rect 642 1631 645 1638
rect 745 1649 748 1652
rect 787 1649 790 1652
rect 658 1641 661 1645
rect 668 1641 671 1645
rect 668 1637 677 1641
rect 689 1640 692 1645
rect 714 1641 717 1645
rect 658 1631 661 1637
rect 668 1631 671 1637
rect 689 1636 690 1640
rect 694 1636 697 1639
rect 716 1637 717 1641
rect 732 1640 735 1645
rect 756 1644 759 1649
rect 764 1645 775 1648
rect 787 1646 795 1649
rect 689 1631 692 1636
rect 714 1631 717 1637
rect 732 1631 735 1636
rect 218 1619 234 1623
rect 238 1619 301 1623
rect 305 1619 337 1623
rect 341 1619 553 1623
rect 634 1618 635 1622
rect 659 1619 660 1623
rect 706 1618 707 1622
rect 222 1612 255 1616
rect 259 1612 285 1616
rect 289 1612 313 1616
rect 317 1612 493 1616
rect 228 1602 231 1612
rect 249 1602 252 1612
rect 265 1602 268 1612
rect 280 1605 287 1609
rect 291 1605 296 1609
rect 307 1602 310 1612
rect 323 1602 326 1612
rect 344 1602 347 1612
rect 523 1611 587 1615
rect 591 1611 646 1615
rect 650 1611 671 1615
rect 675 1611 702 1615
rect 706 1611 735 1615
rect 747 1608 750 1640
rect 764 1639 767 1645
rect 787 1640 790 1646
rect 799 1641 802 1644
rect 810 1644 813 1658
rect 837 1653 840 1658
rect 852 1660 855 1670
rect 882 1666 885 1670
rect 821 1649 822 1652
rect 826 1649 829 1652
rect 1161 1661 1164 1673
rect 1182 1661 1185 1673
rect 1198 1661 1201 1673
rect 1212 1664 1224 1667
rect 1240 1661 1243 1673
rect 1256 1661 1259 1673
rect 1277 1661 1280 1673
rect 1432 1670 1505 1674
rect 1509 1670 1521 1674
rect 1525 1670 1539 1674
rect 1543 1670 1550 1674
rect 1554 1670 1556 1674
rect 1560 1670 1575 1674
rect 1579 1670 1612 1674
rect 1616 1670 1617 1674
rect 1621 1670 1629 1674
rect 1633 1670 1657 1674
rect 1661 1670 1673 1674
rect 1677 1670 1697 1674
rect 1701 1670 1751 1674
rect 1755 1670 1778 1674
rect 1782 1670 1832 1674
rect 1836 1670 1855 1674
rect 1468 1663 1532 1667
rect 1536 1663 1563 1667
rect 1567 1663 1585 1667
rect 1589 1663 1650 1667
rect 1654 1663 1668 1667
rect 1680 1666 1683 1670
rect 868 1649 871 1652
rect 810 1641 818 1644
rect 837 1644 840 1649
rect 810 1636 813 1641
rect 818 1637 822 1641
rect 845 1645 856 1648
rect 868 1646 876 1649
rect 762 1630 767 1635
rect 771 1608 774 1636
rect 801 1608 804 1632
rect 828 1608 831 1640
rect 845 1639 848 1645
rect 868 1640 871 1646
rect 880 1641 883 1644
rect 891 1644 894 1658
rect 1158 1657 1191 1661
rect 1195 1657 1219 1661
rect 1223 1657 1249 1661
rect 1253 1657 1438 1661
rect 1158 1650 1167 1654
rect 1171 1650 1218 1654
rect 1222 1650 1268 1654
rect 1272 1650 1474 1654
rect 1575 1656 1578 1660
rect 1602 1656 1603 1660
rect 1647 1656 1649 1660
rect 1689 1653 1692 1658
rect 1704 1660 1707 1670
rect 1734 1666 1737 1670
rect 1761 1666 1764 1670
rect 891 1641 903 1644
rect 891 1636 894 1641
rect 843 1630 848 1635
rect 852 1608 855 1636
rect 1156 1634 1172 1638
rect 1281 1636 1285 1640
rect 1297 1636 1301 1640
rect 1305 1636 1507 1640
rect 1515 1639 1518 1645
rect 1522 1639 1525 1645
rect 1515 1636 1525 1639
rect 882 1608 885 1632
rect 1515 1631 1518 1636
rect 1164 1627 1168 1631
rect 1180 1627 1301 1631
rect 1522 1631 1525 1636
rect 1531 1641 1534 1645
rect 1531 1637 1533 1641
rect 1537 1637 1539 1641
rect 1547 1640 1550 1645
rect 1575 1642 1578 1645
rect 1547 1638 1558 1640
rect 1531 1631 1534 1637
rect 1547 1636 1553 1638
rect 1547 1631 1550 1636
rect 1557 1636 1558 1638
rect 1576 1638 1578 1642
rect 1575 1631 1578 1638
rect 1678 1649 1681 1652
rect 1720 1649 1723 1652
rect 1591 1641 1594 1645
rect 1601 1641 1604 1645
rect 1601 1637 1610 1641
rect 1622 1640 1625 1645
rect 1647 1641 1650 1645
rect 1591 1631 1594 1637
rect 1601 1631 1604 1637
rect 1622 1636 1623 1640
rect 1627 1636 1630 1639
rect 1649 1637 1650 1641
rect 1665 1640 1668 1645
rect 1689 1644 1692 1649
rect 1697 1645 1708 1648
rect 1720 1646 1728 1649
rect 1622 1631 1625 1636
rect 1647 1631 1650 1637
rect 1665 1631 1668 1636
rect 1151 1619 1167 1623
rect 1171 1619 1234 1623
rect 1238 1619 1270 1623
rect 1274 1619 1486 1623
rect 1567 1618 1568 1622
rect 1592 1619 1593 1623
rect 1639 1618 1640 1622
rect 1155 1612 1188 1616
rect 1192 1612 1218 1616
rect 1222 1612 1246 1616
rect 1250 1612 1426 1616
rect 511 1604 573 1608
rect 577 1604 579 1608
rect 583 1604 587 1608
rect 591 1604 605 1608
rect 609 1604 614 1608
rect 618 1604 623 1608
rect 627 1604 646 1608
rect 650 1604 680 1608
rect 684 1604 695 1608
rect 699 1604 723 1608
rect 727 1604 740 1608
rect 744 1604 764 1608
rect 768 1604 818 1608
rect 825 1604 845 1608
rect 849 1604 899 1608
rect 239 1588 261 1591
rect 265 1588 272 1591
rect 523 1597 587 1601
rect 591 1597 646 1601
rect 650 1597 671 1601
rect 675 1597 702 1601
rect 706 1597 735 1601
rect 297 1588 321 1591
rect 325 1588 330 1591
rect 634 1590 635 1594
rect 659 1589 660 1593
rect 706 1590 707 1594
rect 343 1585 352 1589
rect 230 1582 245 1585
rect 284 1582 303 1585
rect 249 1578 256 1581
rect 281 1575 284 1581
rect 307 1578 314 1581
rect 582 1576 585 1581
rect 589 1576 592 1581
rect 572 1573 574 1576
rect 582 1573 592 1576
rect 228 1559 231 1571
rect 249 1559 252 1571
rect 265 1559 268 1571
rect 284 1562 296 1565
rect 307 1559 310 1571
rect 323 1559 326 1571
rect 344 1559 347 1571
rect 582 1567 585 1573
rect 589 1567 592 1573
rect 598 1575 601 1581
rect 614 1576 617 1581
rect 598 1571 600 1575
rect 604 1571 606 1575
rect 614 1574 620 1576
rect 624 1574 625 1576
rect 614 1572 625 1574
rect 642 1574 645 1581
rect 598 1567 601 1571
rect 614 1567 617 1572
rect 643 1570 645 1574
rect 642 1567 645 1570
rect 658 1575 661 1581
rect 668 1575 671 1581
rect 689 1576 692 1581
rect 668 1571 677 1575
rect 689 1572 690 1576
rect 694 1573 697 1576
rect 714 1575 717 1581
rect 732 1576 735 1581
rect 771 1584 774 1604
rect 852 1584 855 1604
rect 1161 1602 1164 1612
rect 1182 1602 1185 1612
rect 1198 1602 1201 1612
rect 1213 1605 1220 1609
rect 1224 1605 1229 1609
rect 1240 1602 1243 1612
rect 1256 1602 1259 1612
rect 1277 1602 1280 1612
rect 1456 1611 1520 1615
rect 1524 1611 1579 1615
rect 1583 1611 1604 1615
rect 1608 1611 1635 1615
rect 1639 1611 1668 1615
rect 1680 1608 1683 1640
rect 1697 1639 1700 1645
rect 1720 1640 1723 1646
rect 1732 1641 1735 1644
rect 1743 1644 1746 1658
rect 1770 1653 1773 1658
rect 1785 1660 1788 1670
rect 1815 1666 1818 1670
rect 1754 1649 1755 1652
rect 1759 1649 1762 1652
rect 1801 1649 1804 1652
rect 1743 1641 1751 1644
rect 1770 1644 1773 1649
rect 1743 1636 1746 1641
rect 1751 1637 1755 1641
rect 1778 1645 1789 1648
rect 1801 1646 1809 1649
rect 1695 1630 1700 1635
rect 1704 1608 1707 1636
rect 1734 1608 1737 1632
rect 1761 1608 1764 1640
rect 1778 1639 1781 1645
rect 1801 1640 1804 1646
rect 1813 1641 1816 1644
rect 1824 1644 1827 1658
rect 1824 1641 1836 1644
rect 1824 1636 1827 1641
rect 1776 1630 1781 1635
rect 1785 1608 1788 1636
rect 1815 1608 1818 1632
rect 1444 1604 1506 1608
rect 1510 1604 1512 1608
rect 1516 1604 1520 1608
rect 1524 1604 1538 1608
rect 1542 1604 1547 1608
rect 1551 1604 1556 1608
rect 1560 1604 1579 1608
rect 1583 1604 1613 1608
rect 1617 1604 1628 1608
rect 1632 1604 1656 1608
rect 1660 1604 1673 1608
rect 1677 1604 1697 1608
rect 1701 1604 1751 1608
rect 1758 1604 1778 1608
rect 1782 1604 1832 1608
rect 1172 1588 1194 1591
rect 1198 1588 1205 1591
rect 1456 1597 1520 1601
rect 1524 1597 1579 1601
rect 1583 1597 1604 1601
rect 1608 1597 1635 1601
rect 1639 1597 1668 1601
rect 1230 1588 1254 1591
rect 1258 1588 1263 1591
rect 1567 1590 1568 1594
rect 1592 1589 1593 1593
rect 1639 1590 1640 1594
rect 1276 1585 1285 1589
rect 1163 1582 1178 1585
rect 658 1567 661 1571
rect 668 1567 671 1571
rect 689 1567 692 1572
rect 716 1571 717 1575
rect 714 1567 717 1571
rect 732 1567 735 1572
rect 762 1571 767 1576
rect 771 1572 772 1575
rect 787 1574 790 1580
rect 787 1571 795 1574
rect 842 1571 847 1576
rect 851 1572 853 1575
rect 868 1574 871 1580
rect 1217 1582 1236 1585
rect 1182 1578 1189 1581
rect 1214 1575 1217 1581
rect 868 1571 876 1574
rect 1240 1578 1247 1581
rect 1515 1576 1518 1581
rect 1522 1576 1525 1581
rect 1505 1573 1507 1576
rect 1515 1573 1525 1576
rect 787 1568 790 1571
rect 868 1568 871 1571
rect 218 1555 255 1559
rect 259 1555 285 1559
rect 289 1555 313 1559
rect 317 1555 505 1559
rect 642 1552 645 1556
rect 669 1552 670 1556
rect 714 1552 716 1556
rect 218 1548 236 1552
rect 240 1548 286 1552
rect 290 1548 337 1552
rect 341 1548 541 1552
rect 587 1545 599 1549
rect 603 1545 630 1549
rect 634 1545 652 1549
rect 656 1545 717 1549
rect 721 1545 735 1549
rect 771 1542 774 1560
rect 852 1542 855 1560
rect 1161 1559 1164 1571
rect 1182 1559 1185 1571
rect 1198 1559 1201 1571
rect 1217 1562 1229 1565
rect 1240 1559 1243 1571
rect 1256 1559 1259 1571
rect 1277 1559 1280 1571
rect 1515 1567 1518 1573
rect 1522 1567 1525 1573
rect 1531 1575 1534 1581
rect 1547 1576 1550 1581
rect 1531 1571 1533 1575
rect 1537 1571 1539 1575
rect 1547 1574 1553 1576
rect 1557 1574 1558 1576
rect 1547 1572 1558 1574
rect 1575 1574 1578 1581
rect 1531 1567 1534 1571
rect 1547 1567 1550 1572
rect 1576 1570 1578 1574
rect 1575 1567 1578 1570
rect 1591 1575 1594 1581
rect 1601 1575 1604 1581
rect 1622 1576 1625 1581
rect 1601 1571 1610 1575
rect 1622 1572 1623 1576
rect 1627 1573 1630 1576
rect 1647 1575 1650 1581
rect 1665 1576 1668 1581
rect 1704 1584 1707 1604
rect 1785 1584 1788 1604
rect 1591 1567 1594 1571
rect 1601 1567 1604 1571
rect 1622 1567 1625 1572
rect 1649 1571 1650 1575
rect 1647 1567 1650 1571
rect 1665 1567 1668 1572
rect 1695 1571 1700 1576
rect 1704 1572 1705 1575
rect 1720 1574 1723 1580
rect 1720 1571 1728 1574
rect 1775 1571 1780 1576
rect 1784 1572 1786 1575
rect 1801 1574 1804 1580
rect 1801 1571 1809 1574
rect 1720 1568 1723 1571
rect 1801 1568 1804 1571
rect 1151 1555 1188 1559
rect 1192 1555 1218 1559
rect 1222 1555 1246 1559
rect 1250 1555 1438 1559
rect 1575 1552 1578 1556
rect 1602 1552 1603 1556
rect 1647 1552 1649 1556
rect 1151 1548 1169 1552
rect 1173 1548 1219 1552
rect 1223 1548 1270 1552
rect 1274 1548 1474 1552
rect 1520 1545 1532 1549
rect 1536 1545 1563 1549
rect 1567 1545 1585 1549
rect 1589 1545 1650 1549
rect 1654 1545 1668 1549
rect 1704 1542 1707 1560
rect 1785 1542 1788 1560
rect 499 1538 572 1542
rect 576 1538 588 1542
rect 592 1538 606 1542
rect 610 1538 617 1542
rect 621 1538 623 1542
rect 627 1538 642 1542
rect 646 1538 679 1542
rect 683 1538 684 1542
rect 688 1538 696 1542
rect 700 1538 724 1542
rect 728 1538 740 1542
rect 744 1538 764 1542
rect 768 1538 818 1542
rect 822 1538 845 1542
rect 849 1538 907 1542
rect 911 1538 922 1542
rect 1432 1538 1505 1542
rect 1509 1538 1521 1542
rect 1525 1538 1539 1542
rect 1543 1538 1550 1542
rect 1554 1538 1556 1542
rect 1560 1538 1575 1542
rect 1579 1538 1612 1542
rect 1616 1538 1617 1542
rect 1621 1538 1629 1542
rect 1633 1538 1657 1542
rect 1661 1538 1673 1542
rect 1677 1538 1697 1542
rect 1701 1538 1751 1542
rect 1755 1538 1778 1542
rect 1782 1538 1840 1542
rect 1844 1538 1855 1542
rect 535 1531 583 1535
rect 587 1531 599 1535
rect 603 1531 630 1535
rect 634 1531 652 1535
rect 656 1531 717 1535
rect 721 1531 735 1535
rect 771 1528 774 1538
rect 801 1534 804 1538
rect 852 1534 855 1538
rect 642 1524 645 1528
rect 669 1524 670 1528
rect 714 1524 716 1528
rect 571 1504 574 1507
rect 582 1507 585 1513
rect 589 1507 592 1513
rect 582 1504 592 1507
rect 582 1499 585 1504
rect 589 1499 592 1504
rect 598 1509 601 1513
rect 598 1505 600 1509
rect 604 1505 606 1509
rect 614 1508 617 1513
rect 642 1510 645 1513
rect 614 1506 625 1508
rect 598 1499 601 1505
rect 614 1504 620 1506
rect 614 1499 617 1504
rect 624 1504 625 1506
rect 643 1506 645 1510
rect 642 1499 645 1506
rect 787 1517 790 1520
rect 658 1509 661 1513
rect 668 1509 671 1513
rect 668 1505 677 1509
rect 689 1508 692 1513
rect 714 1509 717 1513
rect 658 1499 661 1505
rect 668 1499 671 1505
rect 689 1504 690 1508
rect 694 1504 697 1507
rect 716 1505 717 1509
rect 732 1508 735 1513
rect 764 1513 775 1516
rect 787 1514 795 1517
rect 689 1499 692 1504
rect 714 1499 717 1505
rect 764 1507 767 1513
rect 787 1508 790 1514
rect 799 1509 802 1512
rect 810 1512 813 1526
rect 861 1521 864 1526
rect 876 1528 879 1538
rect 906 1534 909 1538
rect 845 1517 846 1520
rect 850 1517 853 1520
rect 1468 1531 1516 1535
rect 1520 1531 1532 1535
rect 1536 1531 1563 1535
rect 1567 1531 1585 1535
rect 1589 1531 1650 1535
rect 1654 1531 1668 1535
rect 1704 1528 1707 1538
rect 1734 1534 1737 1538
rect 1785 1534 1788 1538
rect 892 1517 895 1520
rect 818 1512 823 1517
rect 861 1512 864 1517
rect 810 1509 818 1512
rect 732 1499 735 1504
rect 810 1504 813 1509
rect 869 1513 880 1516
rect 892 1514 900 1517
rect 762 1498 767 1503
rect 634 1486 635 1490
rect 659 1487 660 1491
rect 706 1486 707 1490
rect 523 1479 587 1483
rect 591 1479 646 1483
rect 650 1479 671 1483
rect 675 1479 702 1483
rect 706 1479 735 1483
rect 771 1476 774 1504
rect 801 1476 804 1500
rect 852 1476 855 1508
rect 869 1507 872 1513
rect 892 1508 895 1514
rect 904 1509 907 1512
rect 915 1512 918 1526
rect 1575 1524 1578 1528
rect 1602 1524 1603 1528
rect 1647 1524 1649 1528
rect 915 1509 921 1512
rect 915 1504 918 1509
rect 1504 1504 1507 1507
rect 1515 1507 1518 1513
rect 1522 1507 1525 1513
rect 1515 1504 1525 1507
rect 867 1498 872 1503
rect 876 1476 879 1504
rect 906 1476 909 1500
rect 1515 1499 1518 1504
rect 1522 1499 1525 1504
rect 1531 1509 1534 1513
rect 1531 1505 1533 1509
rect 1537 1505 1539 1509
rect 1547 1508 1550 1513
rect 1575 1510 1578 1513
rect 1547 1506 1558 1508
rect 1531 1499 1534 1505
rect 1547 1504 1553 1506
rect 1547 1499 1550 1504
rect 1557 1504 1558 1506
rect 1576 1506 1578 1510
rect 1575 1499 1578 1506
rect 1720 1517 1723 1520
rect 1591 1509 1594 1513
rect 1601 1509 1604 1513
rect 1601 1505 1610 1509
rect 1622 1508 1625 1513
rect 1647 1509 1650 1513
rect 1591 1499 1594 1505
rect 1601 1499 1604 1505
rect 1622 1504 1623 1508
rect 1627 1504 1630 1507
rect 1649 1505 1650 1509
rect 1665 1508 1668 1513
rect 1697 1513 1708 1516
rect 1720 1514 1728 1517
rect 1622 1499 1625 1504
rect 1647 1499 1650 1505
rect 1697 1507 1700 1513
rect 1720 1508 1723 1514
rect 1732 1509 1735 1512
rect 1743 1512 1746 1526
rect 1794 1521 1797 1526
rect 1809 1528 1812 1538
rect 1839 1534 1842 1538
rect 1778 1517 1779 1520
rect 1783 1517 1786 1520
rect 1825 1517 1828 1520
rect 1751 1512 1756 1517
rect 1794 1512 1797 1517
rect 1743 1509 1751 1512
rect 1665 1499 1668 1504
rect 1743 1504 1746 1509
rect 1802 1513 1813 1516
rect 1825 1514 1833 1517
rect 1695 1498 1700 1503
rect 1567 1486 1568 1490
rect 1592 1487 1593 1491
rect 1639 1486 1640 1490
rect 1456 1479 1520 1483
rect 1524 1479 1579 1483
rect 1583 1479 1604 1483
rect 1608 1479 1635 1483
rect 1639 1479 1668 1483
rect 1704 1476 1707 1504
rect 1734 1476 1737 1500
rect 1785 1476 1788 1508
rect 1802 1507 1805 1513
rect 1825 1508 1828 1514
rect 1837 1509 1840 1512
rect 1848 1512 1851 1526
rect 1848 1509 1854 1512
rect 1848 1504 1851 1509
rect 1800 1498 1805 1503
rect 1809 1476 1812 1504
rect 1839 1476 1842 1500
rect 511 1472 573 1476
rect 577 1472 579 1476
rect 583 1472 587 1476
rect 591 1472 605 1476
rect 609 1472 614 1476
rect 618 1472 623 1476
rect 627 1472 646 1476
rect 650 1472 680 1476
rect 684 1472 695 1476
rect 699 1472 723 1476
rect 727 1472 740 1476
rect 744 1472 764 1476
rect 768 1472 818 1476
rect 822 1472 845 1476
rect 849 1472 869 1476
rect 873 1472 921 1476
rect 1444 1472 1506 1476
rect 1510 1472 1512 1476
rect 1516 1472 1520 1476
rect 1524 1472 1538 1476
rect 1542 1472 1547 1476
rect 1551 1472 1556 1476
rect 1560 1472 1579 1476
rect 1583 1472 1613 1476
rect 1617 1472 1628 1476
rect 1632 1472 1656 1476
rect 1660 1472 1673 1476
rect 1677 1472 1697 1476
rect 1701 1472 1751 1476
rect 1755 1472 1778 1476
rect 1782 1472 1802 1476
rect 1806 1472 1854 1476
rect 523 1465 587 1469
rect 591 1465 646 1469
rect 650 1465 671 1469
rect 675 1465 702 1469
rect 706 1465 735 1469
rect 634 1458 635 1462
rect 659 1457 660 1461
rect 706 1458 707 1462
rect 771 1453 774 1472
rect 876 1453 879 1472
rect 1456 1465 1520 1469
rect 1524 1465 1579 1469
rect 1583 1465 1604 1469
rect 1608 1465 1635 1469
rect 1639 1465 1668 1469
rect 1567 1458 1568 1462
rect 1592 1457 1593 1461
rect 1639 1458 1640 1462
rect 1704 1453 1707 1472
rect 1809 1453 1812 1472
rect 582 1444 585 1449
rect 589 1444 592 1449
rect 572 1441 574 1444
rect 582 1441 592 1444
rect 582 1435 585 1441
rect 589 1435 592 1441
rect 598 1443 601 1449
rect 614 1444 617 1449
rect 598 1439 600 1443
rect 604 1439 606 1443
rect 614 1442 620 1444
rect 624 1442 625 1444
rect 614 1440 625 1442
rect 642 1442 645 1449
rect 598 1435 601 1439
rect 614 1435 617 1440
rect 643 1438 645 1442
rect 642 1435 645 1438
rect 658 1443 661 1449
rect 668 1443 671 1449
rect 689 1444 692 1449
rect 668 1439 677 1443
rect 689 1440 690 1444
rect 694 1441 697 1444
rect 714 1443 717 1449
rect 732 1444 735 1449
rect 658 1435 661 1439
rect 668 1435 671 1439
rect 689 1435 692 1440
rect 716 1439 717 1443
rect 761 1440 766 1445
rect 770 1441 772 1444
rect 787 1443 790 1449
rect 787 1440 795 1443
rect 867 1440 872 1445
rect 876 1441 877 1444
rect 892 1443 895 1449
rect 892 1440 900 1443
rect 1515 1444 1518 1449
rect 1522 1444 1525 1449
rect 1505 1441 1507 1444
rect 1515 1441 1525 1444
rect 714 1435 717 1439
rect 732 1435 735 1440
rect 787 1437 790 1440
rect 892 1437 895 1440
rect 1515 1435 1518 1441
rect 642 1420 645 1424
rect 669 1420 670 1424
rect 714 1420 716 1424
rect 535 1413 599 1417
rect 603 1413 630 1417
rect 634 1413 652 1417
rect 656 1413 717 1417
rect 721 1413 735 1417
rect 771 1410 774 1429
rect 876 1410 879 1429
rect 1522 1435 1525 1441
rect 1531 1443 1534 1449
rect 1547 1444 1550 1449
rect 1531 1439 1533 1443
rect 1537 1439 1539 1443
rect 1547 1442 1553 1444
rect 1557 1442 1558 1444
rect 1547 1440 1558 1442
rect 1575 1442 1578 1449
rect 1531 1435 1534 1439
rect 1547 1435 1550 1440
rect 1576 1438 1578 1442
rect 1575 1435 1578 1438
rect 1591 1443 1594 1449
rect 1601 1443 1604 1449
rect 1622 1444 1625 1449
rect 1601 1439 1610 1443
rect 1622 1440 1623 1444
rect 1627 1441 1630 1444
rect 1647 1443 1650 1449
rect 1665 1444 1668 1449
rect 1591 1435 1594 1439
rect 1601 1435 1604 1439
rect 1622 1435 1625 1440
rect 1649 1439 1650 1443
rect 1694 1440 1699 1445
rect 1703 1441 1705 1444
rect 1720 1443 1723 1449
rect 1720 1440 1728 1443
rect 1800 1440 1805 1445
rect 1809 1441 1810 1444
rect 1825 1443 1828 1449
rect 1825 1440 1833 1443
rect 1647 1435 1650 1439
rect 1665 1435 1668 1440
rect 1720 1437 1723 1440
rect 1825 1437 1828 1440
rect 1575 1420 1578 1424
rect 1602 1420 1603 1424
rect 1647 1420 1649 1424
rect 1468 1413 1532 1417
rect 1536 1413 1563 1417
rect 1567 1413 1585 1417
rect 1589 1413 1650 1417
rect 1654 1413 1668 1417
rect 1704 1410 1707 1429
rect 1809 1410 1812 1429
rect 499 1406 572 1410
rect 576 1406 588 1410
rect 592 1406 606 1410
rect 610 1406 617 1410
rect 621 1406 623 1410
rect 627 1406 642 1410
rect 646 1406 679 1410
rect 683 1406 684 1410
rect 688 1406 696 1410
rect 700 1406 724 1410
rect 728 1406 740 1410
rect 744 1406 764 1410
rect 768 1406 818 1410
rect 822 1406 845 1410
rect 849 1406 899 1410
rect 903 1406 907 1410
rect 911 1406 935 1410
rect 939 1406 989 1410
rect 1432 1406 1505 1410
rect 1509 1406 1521 1410
rect 1525 1406 1539 1410
rect 1543 1406 1550 1410
rect 1554 1406 1556 1410
rect 1560 1406 1575 1410
rect 1579 1406 1612 1410
rect 1616 1406 1617 1410
rect 1621 1406 1629 1410
rect 1633 1406 1657 1410
rect 1661 1406 1673 1410
rect 1677 1406 1697 1410
rect 1701 1406 1751 1410
rect 1755 1406 1778 1410
rect 1782 1406 1832 1410
rect 1836 1406 1840 1410
rect 1844 1406 1868 1410
rect 1872 1406 1922 1410
rect 535 1399 599 1403
rect 603 1399 630 1403
rect 634 1399 652 1403
rect 656 1399 717 1403
rect 721 1399 735 1403
rect 771 1396 774 1406
rect 801 1402 804 1406
rect 828 1402 831 1406
rect 642 1392 645 1396
rect 669 1392 670 1396
rect 714 1392 716 1396
rect 571 1372 574 1375
rect 582 1375 585 1381
rect 589 1375 592 1381
rect 582 1372 592 1375
rect 582 1367 585 1372
rect 589 1367 592 1372
rect 598 1377 601 1381
rect 598 1373 600 1377
rect 604 1373 606 1377
rect 614 1376 617 1381
rect 642 1378 645 1381
rect 614 1374 625 1376
rect 598 1367 601 1373
rect 614 1372 620 1374
rect 614 1367 617 1372
rect 624 1372 625 1374
rect 643 1374 645 1378
rect 642 1367 645 1374
rect 787 1385 790 1388
rect 658 1377 661 1381
rect 668 1377 671 1381
rect 668 1373 677 1377
rect 689 1376 692 1381
rect 714 1377 717 1381
rect 658 1367 661 1373
rect 668 1367 671 1373
rect 689 1372 690 1376
rect 694 1372 697 1375
rect 716 1373 717 1377
rect 732 1376 735 1381
rect 764 1381 775 1384
rect 787 1382 795 1385
rect 689 1367 692 1372
rect 714 1367 717 1373
rect 764 1375 767 1381
rect 787 1376 790 1382
rect 799 1377 802 1380
rect 810 1380 813 1394
rect 837 1389 840 1394
rect 852 1396 855 1406
rect 882 1402 885 1406
rect 918 1402 921 1406
rect 821 1385 822 1388
rect 826 1385 829 1388
rect 868 1385 871 1388
rect 810 1377 818 1380
rect 837 1380 840 1385
rect 732 1367 735 1372
rect 810 1372 813 1377
rect 818 1373 822 1377
rect 845 1381 856 1384
rect 868 1382 876 1385
rect 762 1366 767 1371
rect 634 1354 635 1358
rect 659 1355 660 1359
rect 706 1354 707 1358
rect 523 1347 587 1351
rect 591 1347 646 1351
rect 650 1347 671 1351
rect 675 1347 702 1351
rect 706 1347 735 1351
rect 771 1344 774 1372
rect 801 1344 804 1368
rect 828 1344 831 1376
rect 845 1375 848 1381
rect 868 1376 871 1382
rect 880 1377 883 1380
rect 891 1380 894 1394
rect 927 1389 930 1394
rect 942 1396 945 1406
rect 972 1402 975 1406
rect 916 1385 919 1388
rect 1468 1399 1532 1403
rect 1536 1399 1563 1403
rect 1567 1399 1585 1403
rect 1589 1399 1650 1403
rect 1654 1399 1668 1403
rect 1704 1396 1707 1406
rect 1734 1402 1737 1406
rect 1761 1402 1764 1406
rect 958 1385 961 1388
rect 891 1377 900 1380
rect 927 1380 930 1385
rect 891 1372 894 1377
rect 843 1366 848 1371
rect 852 1344 855 1372
rect 934 1383 946 1384
rect 938 1381 946 1383
rect 958 1382 966 1385
rect 958 1376 961 1382
rect 970 1377 973 1380
rect 981 1380 984 1394
rect 1575 1392 1578 1396
rect 1602 1392 1603 1396
rect 1647 1392 1649 1396
rect 981 1377 1001 1380
rect 882 1344 885 1368
rect 918 1344 921 1376
rect 981 1372 984 1377
rect 1504 1372 1507 1375
rect 1515 1375 1518 1381
rect 1522 1375 1525 1381
rect 1515 1372 1525 1375
rect 942 1344 945 1372
rect 972 1344 975 1368
rect 1515 1367 1518 1372
rect 1522 1367 1525 1372
rect 1531 1377 1534 1381
rect 1531 1373 1533 1377
rect 1537 1373 1539 1377
rect 1547 1376 1550 1381
rect 1575 1378 1578 1381
rect 1547 1374 1558 1376
rect 1531 1367 1534 1373
rect 1547 1372 1553 1374
rect 1547 1367 1550 1372
rect 1557 1372 1558 1374
rect 1576 1374 1578 1378
rect 1575 1367 1578 1374
rect 1720 1385 1723 1388
rect 1591 1377 1594 1381
rect 1601 1377 1604 1381
rect 1601 1373 1610 1377
rect 1622 1376 1625 1381
rect 1647 1377 1650 1381
rect 1591 1367 1594 1373
rect 1601 1367 1604 1373
rect 1622 1372 1623 1376
rect 1627 1372 1630 1375
rect 1649 1373 1650 1377
rect 1665 1376 1668 1381
rect 1697 1381 1708 1384
rect 1720 1382 1728 1385
rect 1622 1367 1625 1372
rect 1647 1367 1650 1373
rect 1697 1375 1700 1381
rect 1720 1376 1723 1382
rect 1732 1377 1735 1380
rect 1743 1380 1746 1394
rect 1770 1389 1773 1394
rect 1785 1396 1788 1406
rect 1815 1402 1818 1406
rect 1851 1402 1854 1406
rect 1754 1385 1755 1388
rect 1759 1385 1762 1388
rect 1801 1385 1804 1388
rect 1743 1377 1751 1380
rect 1770 1380 1773 1385
rect 1665 1367 1668 1372
rect 1743 1372 1746 1377
rect 1751 1373 1755 1377
rect 1778 1381 1789 1384
rect 1801 1382 1809 1385
rect 1695 1366 1700 1371
rect 1567 1354 1568 1358
rect 1592 1355 1593 1359
rect 1639 1354 1640 1358
rect 1456 1347 1520 1351
rect 1524 1347 1579 1351
rect 1583 1347 1604 1351
rect 1608 1347 1635 1351
rect 1639 1347 1668 1351
rect 1704 1344 1707 1372
rect 1734 1344 1737 1368
rect 1761 1344 1764 1376
rect 1778 1375 1781 1381
rect 1801 1376 1804 1382
rect 1813 1377 1816 1380
rect 1824 1380 1827 1394
rect 1860 1389 1863 1394
rect 1875 1396 1878 1406
rect 1905 1402 1908 1406
rect 1849 1385 1852 1388
rect 1891 1385 1894 1388
rect 1824 1377 1833 1380
rect 1860 1380 1863 1385
rect 1824 1372 1827 1377
rect 1776 1366 1781 1371
rect 1785 1344 1788 1372
rect 1867 1383 1879 1384
rect 1871 1381 1879 1383
rect 1891 1382 1899 1385
rect 1891 1376 1894 1382
rect 1903 1377 1906 1380
rect 1914 1380 1917 1394
rect 1914 1377 1934 1380
rect 1815 1344 1818 1368
rect 1851 1344 1854 1376
rect 1914 1372 1917 1377
rect 1875 1344 1878 1372
rect 1905 1344 1908 1368
rect 511 1340 573 1344
rect 577 1340 579 1344
rect 583 1340 587 1344
rect 591 1340 605 1344
rect 609 1340 614 1344
rect 618 1340 623 1344
rect 627 1340 646 1344
rect 650 1340 680 1344
rect 684 1340 695 1344
rect 699 1340 723 1344
rect 727 1340 740 1344
rect 744 1340 764 1344
rect 768 1340 818 1344
rect 825 1340 845 1344
rect 849 1340 899 1344
rect 903 1340 935 1344
rect 939 1340 989 1344
rect 1444 1340 1506 1344
rect 1510 1340 1512 1344
rect 1516 1340 1520 1344
rect 1524 1340 1538 1344
rect 1542 1340 1547 1344
rect 1551 1340 1556 1344
rect 1560 1340 1579 1344
rect 1583 1340 1613 1344
rect 1617 1340 1628 1344
rect 1632 1340 1656 1344
rect 1660 1340 1673 1344
rect 1677 1340 1697 1344
rect 1701 1340 1751 1344
rect 1758 1340 1778 1344
rect 1782 1340 1832 1344
rect 1836 1340 1868 1344
rect 1872 1340 1922 1344
rect 523 1333 587 1337
rect 591 1333 646 1337
rect 650 1333 671 1337
rect 675 1333 702 1337
rect 706 1333 735 1337
rect 634 1326 635 1330
rect 659 1325 660 1329
rect 706 1326 707 1330
rect 582 1312 585 1317
rect 589 1312 592 1317
rect 572 1309 574 1312
rect 582 1309 592 1312
rect 582 1303 585 1309
rect 589 1303 592 1309
rect 598 1311 601 1317
rect 614 1312 617 1317
rect 598 1307 600 1311
rect 604 1307 606 1311
rect 614 1310 620 1312
rect 624 1310 625 1312
rect 614 1308 625 1310
rect 642 1310 645 1317
rect 598 1303 601 1307
rect 614 1303 617 1308
rect 643 1306 645 1310
rect 642 1303 645 1306
rect 658 1311 661 1317
rect 668 1311 671 1317
rect 689 1312 692 1317
rect 668 1307 677 1311
rect 689 1308 690 1312
rect 694 1309 697 1312
rect 714 1311 717 1317
rect 732 1312 735 1317
rect 771 1318 774 1340
rect 852 1318 855 1340
rect 942 1318 945 1340
rect 1456 1333 1520 1337
rect 1524 1333 1579 1337
rect 1583 1333 1604 1337
rect 1608 1333 1635 1337
rect 1639 1333 1668 1337
rect 1567 1326 1568 1330
rect 1592 1325 1593 1329
rect 1639 1326 1640 1330
rect 658 1303 661 1307
rect 668 1303 671 1307
rect 689 1303 692 1308
rect 716 1307 717 1311
rect 714 1303 717 1307
rect 732 1303 735 1308
rect 762 1305 767 1310
rect 771 1306 772 1309
rect 787 1308 790 1314
rect 787 1305 795 1308
rect 842 1305 847 1310
rect 851 1306 853 1309
rect 868 1308 871 1314
rect 868 1305 876 1308
rect 935 1306 943 1309
rect 958 1308 961 1314
rect 1515 1312 1518 1317
rect 1522 1312 1525 1317
rect 1505 1309 1507 1312
rect 958 1305 966 1308
rect 1515 1309 1525 1312
rect 787 1302 790 1305
rect 868 1302 871 1305
rect 958 1302 961 1305
rect 1515 1303 1518 1309
rect 642 1288 645 1292
rect 669 1288 670 1292
rect 714 1288 716 1292
rect 1522 1303 1525 1309
rect 1531 1311 1534 1317
rect 1547 1312 1550 1317
rect 1531 1307 1533 1311
rect 1537 1307 1539 1311
rect 1547 1310 1553 1312
rect 1557 1310 1558 1312
rect 1547 1308 1558 1310
rect 1575 1310 1578 1317
rect 1531 1303 1534 1307
rect 1547 1303 1550 1308
rect 1576 1306 1578 1310
rect 1575 1303 1578 1306
rect 1591 1311 1594 1317
rect 1601 1311 1604 1317
rect 1622 1312 1625 1317
rect 1601 1307 1610 1311
rect 1622 1308 1623 1312
rect 1627 1309 1630 1312
rect 1647 1311 1650 1317
rect 1665 1312 1668 1317
rect 1704 1318 1707 1340
rect 1785 1318 1788 1340
rect 1875 1318 1878 1340
rect 1591 1303 1594 1307
rect 1601 1303 1604 1307
rect 1622 1303 1625 1308
rect 1649 1307 1650 1311
rect 1647 1303 1650 1307
rect 1665 1303 1668 1308
rect 1695 1305 1700 1310
rect 1704 1306 1705 1309
rect 1720 1308 1723 1314
rect 1720 1305 1728 1308
rect 1775 1305 1780 1310
rect 1784 1306 1786 1309
rect 1801 1308 1804 1314
rect 1801 1305 1809 1308
rect 1868 1306 1876 1309
rect 1891 1308 1894 1314
rect 1891 1305 1899 1308
rect 1720 1302 1723 1305
rect 1801 1302 1804 1305
rect 1891 1302 1894 1305
rect 535 1281 599 1285
rect 603 1281 630 1285
rect 634 1281 652 1285
rect 656 1281 717 1285
rect 721 1281 735 1285
rect 771 1278 774 1294
rect 852 1278 855 1294
rect 942 1278 945 1294
rect 1575 1288 1578 1292
rect 1602 1288 1603 1292
rect 1647 1288 1649 1292
rect 1468 1281 1532 1285
rect 1536 1281 1563 1285
rect 1567 1281 1585 1285
rect 1589 1281 1650 1285
rect 1654 1281 1668 1285
rect 1704 1278 1707 1294
rect 1785 1278 1788 1294
rect 1875 1278 1878 1294
rect 499 1274 572 1278
rect 576 1274 588 1278
rect 592 1274 606 1278
rect 610 1274 617 1278
rect 621 1274 623 1278
rect 627 1274 642 1278
rect 646 1274 679 1278
rect 683 1274 684 1278
rect 688 1274 696 1278
rect 700 1274 724 1278
rect 728 1274 740 1278
rect 744 1274 764 1278
rect 768 1274 818 1278
rect 822 1274 845 1278
rect 849 1274 935 1278
rect 939 1274 993 1278
rect 1432 1274 1505 1278
rect 1509 1274 1521 1278
rect 1525 1274 1539 1278
rect 1543 1274 1550 1278
rect 1554 1274 1556 1278
rect 1560 1274 1575 1278
rect 1579 1274 1612 1278
rect 1616 1274 1617 1278
rect 1621 1274 1629 1278
rect 1633 1274 1657 1278
rect 1661 1274 1673 1278
rect 1677 1274 1697 1278
rect 1701 1274 1751 1278
rect 1755 1274 1778 1278
rect 1782 1274 1868 1278
rect 1872 1274 1926 1278
rect 535 1267 599 1271
rect 603 1267 630 1271
rect 634 1267 652 1271
rect 656 1267 717 1271
rect 721 1267 735 1271
rect 771 1264 774 1274
rect 801 1270 804 1274
rect 642 1260 645 1264
rect 669 1260 670 1264
rect 714 1260 716 1264
rect 571 1240 574 1243
rect 582 1243 585 1249
rect 589 1243 592 1249
rect 582 1240 592 1243
rect 582 1235 585 1240
rect 589 1235 592 1240
rect 598 1245 601 1249
rect 598 1241 600 1245
rect 604 1241 606 1245
rect 614 1244 617 1249
rect 642 1246 645 1249
rect 614 1242 625 1244
rect 598 1235 601 1241
rect 614 1240 620 1242
rect 614 1235 617 1240
rect 624 1240 625 1242
rect 643 1242 645 1246
rect 642 1235 645 1242
rect 1468 1267 1532 1271
rect 1536 1267 1563 1271
rect 1567 1267 1585 1271
rect 1589 1267 1650 1271
rect 1654 1267 1668 1271
rect 1704 1264 1707 1274
rect 1734 1270 1737 1274
rect 787 1253 790 1256
rect 658 1245 661 1249
rect 668 1245 671 1249
rect 668 1241 677 1245
rect 689 1244 692 1249
rect 714 1245 717 1249
rect 658 1235 661 1241
rect 668 1235 671 1241
rect 689 1240 690 1244
rect 694 1240 697 1243
rect 716 1241 717 1245
rect 732 1244 735 1249
rect 764 1249 775 1252
rect 787 1250 795 1253
rect 689 1235 692 1240
rect 714 1235 717 1241
rect 764 1243 767 1249
rect 787 1244 790 1250
rect 799 1245 802 1248
rect 810 1248 813 1262
rect 1575 1260 1578 1264
rect 1602 1260 1603 1264
rect 1647 1260 1649 1264
rect 818 1248 823 1253
rect 810 1245 818 1248
rect 732 1235 735 1240
rect 810 1240 813 1245
rect 1504 1240 1507 1243
rect 1515 1243 1518 1249
rect 1522 1243 1525 1249
rect 1515 1240 1525 1243
rect 762 1234 767 1239
rect 93 1219 102 1223
rect 106 1219 138 1223
rect 142 1219 205 1223
rect 209 1219 234 1223
rect 238 1219 270 1223
rect 274 1219 337 1223
rect 341 1219 366 1223
rect 370 1219 402 1223
rect 406 1219 469 1223
rect 473 1219 553 1223
rect 634 1222 635 1226
rect 659 1223 660 1227
rect 706 1222 707 1226
rect 93 1212 126 1216
rect 130 1212 154 1216
rect 158 1212 184 1216
rect 188 1212 221 1216
rect 225 1212 258 1216
rect 262 1212 286 1216
rect 290 1212 316 1216
rect 320 1212 353 1216
rect 357 1212 390 1216
rect 394 1212 418 1216
rect 422 1212 448 1216
rect 452 1212 485 1216
rect 489 1212 493 1216
rect 566 1215 587 1219
rect 591 1215 596 1219
rect 600 1215 646 1219
rect 650 1215 671 1219
rect 675 1215 702 1219
rect 706 1215 735 1219
rect 771 1212 774 1240
rect 801 1212 804 1236
rect 1515 1235 1518 1240
rect 1522 1235 1525 1240
rect 1531 1245 1534 1249
rect 1531 1241 1533 1245
rect 1537 1241 1539 1245
rect 1547 1244 1550 1249
rect 1575 1246 1578 1249
rect 1547 1242 1558 1244
rect 1531 1235 1534 1241
rect 1547 1240 1553 1242
rect 1547 1235 1550 1240
rect 1557 1240 1558 1242
rect 1576 1242 1578 1246
rect 1575 1235 1578 1242
rect 1720 1253 1723 1256
rect 1591 1245 1594 1249
rect 1601 1245 1604 1249
rect 1601 1241 1610 1245
rect 1622 1244 1625 1249
rect 1647 1245 1650 1249
rect 1591 1235 1594 1241
rect 1601 1235 1604 1241
rect 1622 1240 1623 1244
rect 1627 1240 1630 1243
rect 1649 1241 1650 1245
rect 1665 1244 1668 1249
rect 1697 1249 1708 1252
rect 1720 1250 1728 1253
rect 1622 1235 1625 1240
rect 1647 1235 1650 1241
rect 1697 1243 1700 1249
rect 1720 1244 1723 1250
rect 1732 1245 1735 1248
rect 1743 1248 1746 1262
rect 1751 1248 1756 1253
rect 1743 1245 1751 1248
rect 1665 1235 1668 1240
rect 1743 1240 1746 1245
rect 1695 1234 1700 1239
rect 1026 1219 1035 1223
rect 1039 1219 1071 1223
rect 1075 1219 1138 1223
rect 1142 1219 1167 1223
rect 1171 1219 1203 1223
rect 1207 1219 1270 1223
rect 1274 1219 1299 1223
rect 1303 1219 1335 1223
rect 1339 1219 1402 1223
rect 1406 1219 1486 1223
rect 1567 1222 1568 1226
rect 1592 1223 1593 1227
rect 1639 1222 1640 1226
rect 1026 1212 1059 1216
rect 1063 1212 1087 1216
rect 1091 1212 1117 1216
rect 1121 1212 1154 1216
rect 1158 1212 1191 1216
rect 1195 1212 1219 1216
rect 1223 1212 1249 1216
rect 1253 1212 1286 1216
rect 1290 1212 1323 1216
rect 1327 1212 1351 1216
rect 1355 1212 1381 1216
rect 1385 1212 1418 1216
rect 1422 1212 1426 1216
rect 1499 1215 1520 1219
rect 1524 1215 1529 1219
rect 1533 1215 1579 1219
rect 1583 1215 1604 1219
rect 1608 1215 1635 1219
rect 1639 1215 1668 1219
rect 1704 1212 1707 1240
rect 1734 1212 1737 1236
rect 96 1202 99 1212
rect 117 1202 120 1212
rect 133 1202 136 1212
rect 147 1205 152 1209
rect 156 1205 163 1209
rect 175 1202 178 1212
rect 191 1202 194 1212
rect 212 1202 215 1212
rect 228 1202 231 1212
rect 249 1202 252 1212
rect 265 1202 268 1212
rect 279 1205 284 1209
rect 288 1205 295 1209
rect 307 1202 310 1212
rect 323 1202 326 1212
rect 344 1202 347 1212
rect 360 1202 363 1212
rect 381 1202 384 1212
rect 397 1202 400 1212
rect 411 1205 416 1209
rect 420 1205 427 1209
rect 439 1202 442 1212
rect 455 1202 458 1212
rect 476 1202 479 1212
rect 511 1208 573 1212
rect 577 1208 579 1212
rect 583 1208 587 1212
rect 591 1208 605 1212
rect 609 1208 614 1212
rect 618 1208 623 1212
rect 627 1208 646 1212
rect 650 1208 680 1212
rect 684 1208 695 1212
rect 699 1208 723 1212
rect 727 1208 740 1212
rect 744 1208 764 1212
rect 768 1208 848 1212
rect 852 1208 866 1212
rect 870 1208 875 1212
rect 879 1208 884 1212
rect 888 1208 907 1212
rect 911 1208 941 1212
rect 945 1208 956 1212
rect 960 1208 984 1212
rect 988 1208 997 1212
rect 113 1188 118 1191
rect 122 1188 146 1191
rect 171 1188 178 1191
rect 182 1188 204 1191
rect 224 1188 231 1191
rect 245 1188 250 1191
rect 254 1188 278 1191
rect 303 1188 310 1191
rect 314 1188 336 1191
rect 356 1188 363 1191
rect 377 1188 382 1191
rect 386 1188 410 1191
rect 523 1201 587 1205
rect 591 1201 596 1205
rect 600 1201 646 1205
rect 650 1201 671 1205
rect 675 1201 702 1205
rect 706 1201 735 1205
rect 435 1188 442 1191
rect 446 1188 468 1191
rect 634 1194 635 1198
rect 659 1193 660 1197
rect 706 1194 707 1198
rect 129 1178 136 1181
rect 140 1182 159 1185
rect 159 1175 162 1181
rect 187 1178 194 1181
rect 198 1182 213 1185
rect 261 1178 268 1181
rect 272 1182 291 1185
rect 291 1175 294 1181
rect 319 1178 326 1181
rect 330 1182 345 1185
rect 393 1178 400 1181
rect 404 1182 423 1185
rect 423 1175 426 1181
rect 451 1178 458 1181
rect 462 1182 479 1185
rect 582 1180 585 1185
rect 589 1180 592 1185
rect 572 1177 574 1180
rect 582 1177 592 1180
rect 582 1171 585 1177
rect 96 1159 99 1171
rect 117 1159 120 1171
rect 133 1159 136 1171
rect 147 1162 159 1165
rect 175 1159 178 1171
rect 191 1159 194 1171
rect 212 1159 215 1171
rect 228 1159 231 1171
rect 249 1159 252 1171
rect 265 1159 268 1171
rect 279 1162 291 1165
rect 307 1159 310 1171
rect 323 1159 326 1171
rect 344 1159 347 1171
rect 360 1159 363 1171
rect 381 1159 384 1171
rect 397 1159 400 1171
rect 411 1162 423 1165
rect 439 1159 442 1171
rect 455 1159 458 1171
rect 476 1159 479 1171
rect 589 1171 592 1177
rect 598 1179 601 1185
rect 614 1180 617 1185
rect 598 1175 600 1179
rect 604 1175 606 1179
rect 614 1178 620 1180
rect 624 1178 625 1180
rect 614 1176 625 1178
rect 642 1178 645 1185
rect 598 1171 601 1175
rect 614 1171 617 1176
rect 643 1174 645 1178
rect 642 1171 645 1174
rect 658 1179 661 1185
rect 668 1179 671 1185
rect 689 1180 692 1185
rect 668 1175 677 1179
rect 689 1176 690 1180
rect 694 1177 697 1180
rect 714 1179 717 1185
rect 732 1180 735 1185
rect 771 1182 774 1208
rect 807 1201 826 1205
rect 830 1201 848 1205
rect 852 1201 907 1205
rect 911 1201 932 1205
rect 936 1201 963 1205
rect 967 1201 996 1205
rect 1029 1202 1032 1212
rect 1050 1202 1053 1212
rect 1066 1202 1069 1212
rect 1080 1205 1085 1209
rect 1089 1205 1096 1209
rect 1108 1202 1111 1212
rect 1124 1202 1127 1212
rect 1145 1202 1148 1212
rect 1161 1202 1164 1212
rect 1182 1202 1185 1212
rect 1198 1202 1201 1212
rect 1212 1205 1217 1209
rect 1221 1205 1228 1209
rect 1240 1202 1243 1212
rect 1256 1202 1259 1212
rect 1277 1202 1280 1212
rect 1293 1202 1296 1212
rect 1314 1202 1317 1212
rect 1330 1202 1333 1212
rect 1344 1205 1349 1209
rect 1353 1205 1360 1209
rect 1372 1202 1375 1212
rect 1388 1202 1391 1212
rect 1409 1202 1412 1212
rect 1444 1208 1506 1212
rect 1510 1208 1512 1212
rect 1516 1208 1520 1212
rect 1524 1208 1538 1212
rect 1542 1208 1547 1212
rect 1551 1208 1556 1212
rect 1560 1208 1579 1212
rect 1583 1208 1613 1212
rect 1617 1208 1628 1212
rect 1632 1208 1656 1212
rect 1660 1208 1673 1212
rect 1677 1208 1697 1212
rect 1701 1208 1781 1212
rect 1785 1208 1799 1212
rect 1803 1208 1808 1212
rect 1812 1208 1817 1212
rect 1821 1208 1840 1212
rect 1844 1208 1874 1212
rect 1878 1208 1889 1212
rect 1893 1208 1917 1212
rect 1921 1208 1930 1212
rect 807 1189 810 1201
rect 895 1194 896 1198
rect 920 1193 921 1197
rect 967 1194 968 1198
rect 658 1171 661 1175
rect 668 1171 671 1175
rect 689 1171 692 1176
rect 716 1175 717 1179
rect 834 1180 837 1185
rect 843 1180 846 1185
rect 850 1180 853 1185
rect 714 1171 717 1175
rect 732 1171 735 1176
rect 761 1169 766 1174
rect 770 1170 772 1173
rect 787 1172 790 1178
rect 819 1177 853 1180
rect 787 1169 795 1172
rect 787 1166 790 1169
rect 93 1155 126 1159
rect 130 1155 154 1159
rect 158 1155 184 1159
rect 188 1155 258 1159
rect 262 1155 286 1159
rect 290 1155 316 1159
rect 320 1155 390 1159
rect 394 1155 418 1159
rect 422 1155 448 1159
rect 452 1155 505 1159
rect 642 1156 645 1160
rect 669 1156 670 1160
rect 714 1156 716 1160
rect 819 1163 822 1177
rect 843 1171 846 1177
rect 850 1171 853 1177
rect 859 1179 862 1185
rect 875 1180 878 1185
rect 859 1175 861 1179
rect 865 1175 867 1179
rect 875 1178 881 1180
rect 885 1178 886 1180
rect 875 1176 886 1178
rect 903 1178 906 1185
rect 859 1171 862 1175
rect 875 1171 878 1176
rect 904 1174 906 1178
rect 903 1171 906 1174
rect 1046 1188 1051 1191
rect 1055 1188 1079 1191
rect 1104 1188 1111 1191
rect 1115 1188 1137 1191
rect 1157 1188 1164 1191
rect 1178 1188 1183 1191
rect 1187 1188 1211 1191
rect 1236 1188 1243 1191
rect 1247 1188 1269 1191
rect 1289 1188 1296 1191
rect 1310 1188 1315 1191
rect 1319 1188 1343 1191
rect 1456 1201 1520 1205
rect 1524 1201 1529 1205
rect 1533 1201 1579 1205
rect 1583 1201 1604 1205
rect 1608 1201 1635 1205
rect 1639 1201 1668 1205
rect 1368 1188 1375 1191
rect 1379 1188 1401 1191
rect 1567 1194 1568 1198
rect 1592 1193 1593 1197
rect 1639 1194 1640 1198
rect 919 1179 922 1185
rect 929 1179 932 1185
rect 950 1180 953 1185
rect 929 1175 938 1179
rect 950 1176 951 1180
rect 955 1177 958 1180
rect 975 1179 978 1185
rect 993 1180 996 1185
rect 919 1171 922 1175
rect 929 1171 932 1175
rect 950 1171 953 1176
rect 977 1175 978 1179
rect 975 1171 978 1175
rect 993 1171 996 1176
rect 1062 1178 1069 1181
rect 1073 1182 1092 1185
rect 1092 1175 1095 1181
rect 1120 1178 1127 1181
rect 1131 1182 1146 1185
rect 1194 1178 1201 1181
rect 1205 1182 1224 1185
rect 1224 1175 1227 1181
rect 1252 1178 1259 1181
rect 1263 1182 1278 1185
rect 1326 1178 1333 1181
rect 1337 1182 1356 1185
rect 1356 1175 1359 1181
rect 1384 1178 1391 1181
rect 1395 1182 1412 1185
rect 1515 1180 1518 1185
rect 1522 1180 1525 1185
rect 1505 1177 1507 1180
rect 1515 1177 1525 1180
rect 1515 1171 1518 1177
rect 93 1148 102 1152
rect 106 1148 153 1152
rect 157 1148 203 1152
rect 207 1148 234 1152
rect 238 1148 285 1152
rect 289 1148 335 1152
rect 339 1148 366 1152
rect 370 1148 417 1152
rect 421 1148 467 1152
rect 471 1149 541 1152
rect 585 1149 599 1153
rect 603 1149 630 1153
rect 634 1149 652 1153
rect 656 1149 717 1153
rect 721 1149 735 1153
rect 771 1146 774 1158
rect 903 1156 906 1160
rect 930 1156 931 1160
rect 975 1156 977 1160
rect 1029 1159 1032 1171
rect 1050 1159 1053 1171
rect 1066 1159 1069 1171
rect 1080 1162 1092 1165
rect 1108 1159 1111 1171
rect 1124 1159 1127 1171
rect 1145 1159 1148 1171
rect 1161 1159 1164 1171
rect 1182 1159 1185 1171
rect 1198 1159 1201 1171
rect 1212 1162 1224 1165
rect 1240 1159 1243 1171
rect 1256 1159 1259 1171
rect 1277 1159 1280 1171
rect 1293 1159 1296 1171
rect 1314 1159 1317 1171
rect 1330 1159 1333 1171
rect 1344 1162 1356 1165
rect 1372 1159 1375 1171
rect 1388 1159 1391 1171
rect 1409 1159 1412 1171
rect 1522 1171 1525 1177
rect 1531 1179 1534 1185
rect 1547 1180 1550 1185
rect 1531 1175 1533 1179
rect 1537 1175 1539 1179
rect 1547 1178 1553 1180
rect 1557 1178 1558 1180
rect 1547 1176 1558 1178
rect 1575 1178 1578 1185
rect 1531 1171 1534 1175
rect 1547 1171 1550 1176
rect 1576 1174 1578 1178
rect 1575 1171 1578 1174
rect 1591 1179 1594 1185
rect 1601 1179 1604 1185
rect 1622 1180 1625 1185
rect 1601 1175 1610 1179
rect 1622 1176 1623 1180
rect 1627 1177 1630 1180
rect 1647 1179 1650 1185
rect 1665 1180 1668 1185
rect 1704 1182 1707 1208
rect 1740 1201 1759 1205
rect 1763 1201 1781 1205
rect 1785 1201 1840 1205
rect 1844 1201 1865 1205
rect 1869 1201 1896 1205
rect 1900 1201 1929 1205
rect 1740 1189 1743 1201
rect 1828 1194 1829 1198
rect 1853 1193 1854 1197
rect 1900 1194 1901 1198
rect 1591 1171 1594 1175
rect 1601 1171 1604 1175
rect 1622 1171 1625 1176
rect 1649 1175 1650 1179
rect 1767 1180 1770 1185
rect 1776 1180 1779 1185
rect 1783 1180 1786 1185
rect 1647 1171 1650 1175
rect 1665 1171 1668 1176
rect 1694 1169 1699 1174
rect 1703 1170 1705 1173
rect 1720 1172 1723 1178
rect 1752 1177 1786 1180
rect 1720 1169 1728 1172
rect 1720 1166 1723 1169
rect 1026 1155 1059 1159
rect 1063 1155 1087 1159
rect 1091 1155 1117 1159
rect 1121 1155 1191 1159
rect 1195 1155 1219 1159
rect 1223 1155 1249 1159
rect 1253 1155 1323 1159
rect 1327 1155 1351 1159
rect 1355 1155 1381 1159
rect 1385 1155 1438 1159
rect 1575 1156 1578 1160
rect 1602 1156 1603 1160
rect 1647 1156 1649 1160
rect 1752 1163 1755 1177
rect 1776 1171 1779 1177
rect 1783 1171 1786 1177
rect 1792 1179 1795 1185
rect 1808 1180 1811 1185
rect 1792 1175 1794 1179
rect 1798 1175 1800 1179
rect 1808 1178 1814 1180
rect 1818 1178 1819 1180
rect 1808 1176 1819 1178
rect 1836 1178 1839 1185
rect 1792 1171 1795 1175
rect 1808 1171 1811 1176
rect 1837 1174 1839 1178
rect 1836 1171 1839 1174
rect 1852 1179 1855 1185
rect 1862 1179 1865 1185
rect 1883 1180 1886 1185
rect 1862 1175 1871 1179
rect 1883 1176 1884 1180
rect 1888 1177 1891 1180
rect 1908 1179 1911 1185
rect 1926 1180 1929 1185
rect 1852 1171 1855 1175
rect 1862 1171 1865 1175
rect 1883 1171 1886 1176
rect 1910 1175 1911 1179
rect 1908 1171 1911 1175
rect 1926 1171 1929 1176
rect 811 1149 816 1153
rect 820 1149 860 1153
rect 864 1149 891 1153
rect 895 1149 913 1153
rect 917 1149 978 1153
rect 982 1149 996 1153
rect 1026 1148 1035 1152
rect 1039 1148 1086 1152
rect 1090 1148 1136 1152
rect 1140 1148 1167 1152
rect 1171 1148 1218 1152
rect 1222 1148 1268 1152
rect 1272 1148 1299 1152
rect 1303 1148 1350 1152
rect 1354 1148 1400 1152
rect 1404 1149 1474 1152
rect 1518 1149 1532 1153
rect 1536 1149 1563 1153
rect 1567 1149 1585 1153
rect 1589 1149 1650 1153
rect 1654 1149 1668 1153
rect 1704 1146 1707 1158
rect 1836 1156 1839 1160
rect 1863 1156 1864 1160
rect 1908 1156 1910 1160
rect 1744 1149 1749 1153
rect 1753 1149 1793 1153
rect 1797 1149 1824 1153
rect 1828 1149 1846 1153
rect 1850 1149 1911 1153
rect 1915 1149 1929 1153
rect 100 1142 484 1145
rect 499 1142 572 1146
rect 576 1142 588 1146
rect 592 1142 606 1146
rect 610 1142 617 1146
rect 621 1142 623 1146
rect 627 1142 642 1146
rect 646 1142 679 1146
rect 683 1142 684 1146
rect 688 1142 696 1146
rect 700 1142 724 1146
rect 728 1142 764 1146
rect 768 1142 807 1146
rect 811 1142 818 1146
rect 822 1142 833 1146
rect 837 1142 849 1146
rect 853 1142 867 1146
rect 871 1142 878 1146
rect 882 1142 884 1146
rect 888 1142 903 1146
rect 907 1142 940 1146
rect 944 1142 945 1146
rect 949 1142 957 1146
rect 961 1142 985 1146
rect 989 1142 997 1146
rect 1033 1142 1417 1145
rect 1432 1142 1505 1146
rect 1509 1142 1521 1146
rect 1525 1142 1539 1146
rect 1543 1142 1550 1146
rect 1554 1142 1556 1146
rect 1560 1142 1575 1146
rect 1579 1142 1612 1146
rect 1616 1142 1617 1146
rect 1621 1142 1629 1146
rect 1633 1142 1657 1146
rect 1661 1142 1697 1146
rect 1701 1142 1740 1146
rect 1744 1142 1751 1146
rect 1755 1142 1766 1146
rect 1770 1142 1782 1146
rect 1786 1142 1800 1146
rect 1804 1142 1811 1146
rect 1815 1142 1817 1146
rect 1821 1142 1836 1146
rect 1840 1142 1873 1146
rect 1877 1142 1878 1146
rect 1882 1142 1890 1146
rect 1894 1142 1918 1146
rect 1922 1142 1930 1146
rect 243 1135 352 1138
rect 535 1135 581 1139
rect 585 1135 815 1138
rect 1005 1136 1013 1140
rect 1176 1135 1285 1138
rect 1468 1135 1514 1139
rect 1518 1135 1748 1138
rect 1938 1136 1946 1140
rect 223 1127 227 1131
rect 231 1127 235 1131
rect 523 1128 825 1131
rect 1001 1120 1005 1124
rect 1156 1127 1160 1131
rect 1164 1127 1168 1131
rect 1456 1128 1758 1131
rect 1934 1120 1938 1124
rect 83 1116 211 1120
rect 215 1116 231 1120
rect 247 1116 1144 1120
rect 1148 1116 1164 1120
rect 1180 1116 2026 1120
rect 239 1109 484 1112
rect 559 1109 873 1113
rect 877 1109 909 1113
rect 913 1109 976 1113
rect 980 1109 996 1113
rect 1172 1109 1417 1112
rect 1492 1109 1806 1113
rect 1810 1109 1842 1113
rect 1846 1109 1909 1113
rect 1913 1109 1929 1113
rect 254 1102 484 1105
rect 499 1102 859 1106
rect 863 1102 897 1106
rect 901 1102 925 1106
rect 929 1102 955 1106
rect 959 1102 992 1106
rect 223 1093 227 1097
rect 231 1093 235 1097
rect 867 1092 870 1102
rect 888 1092 891 1102
rect 904 1092 907 1102
rect 918 1095 923 1099
rect 927 1095 934 1099
rect 946 1092 949 1102
rect 962 1092 965 1102
rect 983 1092 986 1102
rect 1187 1102 1417 1105
rect 1432 1102 1792 1106
rect 1796 1102 1830 1106
rect 1834 1102 1858 1106
rect 1862 1102 1888 1106
rect 1892 1102 1925 1106
rect 1156 1093 1160 1097
rect 1164 1093 1168 1097
rect 1800 1092 1803 1102
rect 1821 1092 1824 1102
rect 1837 1092 1840 1102
rect 1851 1095 1856 1099
rect 1860 1095 1867 1099
rect 1879 1092 1882 1102
rect 1895 1092 1898 1102
rect 1916 1092 1919 1102
rect 243 1086 353 1089
rect 93 1079 102 1083
rect 106 1079 138 1083
rect 142 1079 205 1083
rect 209 1079 234 1083
rect 238 1079 270 1083
rect 274 1079 337 1083
rect 341 1079 366 1083
rect 370 1079 402 1083
rect 406 1079 469 1083
rect 473 1079 553 1083
rect 93 1072 126 1076
rect 130 1072 154 1076
rect 158 1072 184 1076
rect 188 1072 221 1076
rect 225 1072 258 1076
rect 262 1072 286 1076
rect 290 1072 316 1076
rect 320 1072 353 1076
rect 357 1072 390 1076
rect 394 1072 418 1076
rect 422 1072 448 1076
rect 452 1072 485 1076
rect 489 1072 493 1076
rect 884 1078 889 1081
rect 893 1078 917 1081
rect 1176 1086 1286 1089
rect 942 1078 949 1081
rect 953 1078 975 1081
rect 1026 1079 1035 1083
rect 1039 1079 1071 1083
rect 1075 1079 1138 1083
rect 1142 1079 1167 1083
rect 1171 1079 1203 1083
rect 1207 1079 1270 1083
rect 1274 1079 1299 1083
rect 1303 1079 1335 1083
rect 1339 1079 1402 1083
rect 1406 1079 1486 1083
rect 96 1062 99 1072
rect 117 1062 120 1072
rect 133 1062 136 1072
rect 147 1065 152 1069
rect 156 1065 163 1069
rect 175 1062 178 1072
rect 191 1062 194 1072
rect 212 1062 215 1072
rect 228 1062 231 1072
rect 249 1062 252 1072
rect 265 1062 268 1072
rect 279 1065 284 1069
rect 288 1065 295 1069
rect 307 1062 310 1072
rect 323 1062 326 1072
rect 344 1062 347 1072
rect 360 1062 363 1072
rect 381 1062 384 1072
rect 397 1062 400 1072
rect 411 1065 416 1069
rect 420 1065 427 1069
rect 439 1062 442 1072
rect 455 1062 458 1072
rect 476 1062 479 1072
rect 900 1068 907 1071
rect 911 1072 930 1075
rect 113 1048 118 1051
rect 122 1048 146 1051
rect 171 1048 178 1051
rect 182 1048 204 1051
rect 224 1048 231 1051
rect 245 1048 250 1051
rect 254 1048 278 1051
rect 303 1048 310 1051
rect 314 1048 336 1051
rect 356 1048 363 1051
rect 377 1048 382 1051
rect 386 1048 410 1051
rect 435 1048 442 1051
rect 446 1048 468 1051
rect 930 1065 933 1071
rect 958 1068 965 1071
rect 969 1072 984 1075
rect 1026 1072 1059 1076
rect 1063 1072 1087 1076
rect 1091 1072 1117 1076
rect 1121 1072 1154 1076
rect 1158 1072 1191 1076
rect 1195 1072 1219 1076
rect 1223 1072 1249 1076
rect 1253 1072 1286 1076
rect 1290 1072 1323 1076
rect 1327 1072 1351 1076
rect 1355 1072 1381 1076
rect 1385 1072 1418 1076
rect 1422 1072 1426 1076
rect 1817 1078 1822 1081
rect 1826 1078 1850 1081
rect 1875 1078 1882 1081
rect 1886 1078 1908 1081
rect 1029 1062 1032 1072
rect 1050 1062 1053 1072
rect 1066 1062 1069 1072
rect 1080 1065 1085 1069
rect 1089 1065 1096 1069
rect 1108 1062 1111 1072
rect 1124 1062 1127 1072
rect 1145 1062 1148 1072
rect 1161 1062 1164 1072
rect 1182 1062 1185 1072
rect 1198 1062 1201 1072
rect 1212 1065 1217 1069
rect 1221 1065 1228 1069
rect 1240 1062 1243 1072
rect 1256 1062 1259 1072
rect 1277 1062 1280 1072
rect 1293 1062 1296 1072
rect 1314 1062 1317 1072
rect 1330 1062 1333 1072
rect 1344 1065 1349 1069
rect 1353 1065 1360 1069
rect 1372 1062 1375 1072
rect 1388 1062 1391 1072
rect 1409 1062 1412 1072
rect 1833 1068 1840 1071
rect 1844 1072 1863 1075
rect 867 1049 870 1061
rect 888 1049 891 1061
rect 904 1049 907 1061
rect 918 1052 930 1055
rect 946 1049 949 1061
rect 962 1049 965 1061
rect 983 1049 986 1061
rect 129 1038 136 1041
rect 140 1042 159 1045
rect 159 1035 162 1041
rect 187 1038 194 1041
rect 198 1042 213 1045
rect 261 1038 268 1041
rect 272 1042 291 1045
rect 291 1035 294 1041
rect 319 1038 326 1041
rect 330 1042 345 1045
rect 393 1038 400 1041
rect 404 1042 423 1045
rect 423 1035 426 1041
rect 451 1038 458 1041
rect 462 1042 479 1045
rect 511 1045 897 1049
rect 901 1045 925 1049
rect 929 1045 955 1049
rect 959 1045 996 1049
rect 1046 1048 1051 1051
rect 1055 1048 1079 1051
rect 1104 1048 1111 1051
rect 1115 1048 1137 1051
rect 1157 1048 1164 1051
rect 1178 1048 1183 1051
rect 1187 1048 1211 1051
rect 1236 1048 1243 1051
rect 1247 1048 1269 1051
rect 1289 1048 1296 1051
rect 1310 1048 1315 1051
rect 1319 1048 1343 1051
rect 1368 1048 1375 1051
rect 1379 1048 1401 1051
rect 1863 1065 1866 1071
rect 1891 1068 1898 1071
rect 1902 1072 1917 1075
rect 1800 1049 1803 1061
rect 1821 1049 1824 1061
rect 1837 1049 1840 1061
rect 1851 1052 1863 1055
rect 1879 1049 1882 1061
rect 1895 1049 1898 1061
rect 1916 1049 1919 1061
rect 547 1038 873 1042
rect 877 1038 924 1042
rect 928 1038 974 1042
rect 978 1038 996 1042
rect 1062 1038 1069 1041
rect 1073 1042 1092 1045
rect 96 1019 99 1031
rect 117 1019 120 1031
rect 133 1019 136 1031
rect 147 1022 159 1025
rect 175 1019 178 1031
rect 191 1019 194 1031
rect 212 1019 215 1031
rect 228 1019 231 1031
rect 249 1019 252 1031
rect 265 1019 268 1031
rect 279 1022 291 1025
rect 307 1019 310 1031
rect 323 1019 326 1031
rect 344 1019 347 1031
rect 360 1019 363 1031
rect 381 1019 384 1031
rect 397 1019 400 1031
rect 411 1022 423 1025
rect 439 1019 442 1031
rect 455 1019 458 1031
rect 476 1019 479 1031
rect 870 1031 991 1034
rect 1092 1035 1095 1041
rect 1120 1038 1127 1041
rect 1131 1042 1146 1045
rect 1194 1038 1201 1041
rect 1205 1042 1224 1045
rect 1224 1035 1227 1041
rect 1252 1038 1259 1041
rect 1263 1042 1278 1045
rect 1326 1038 1333 1041
rect 1337 1042 1356 1045
rect 1356 1035 1359 1041
rect 1384 1038 1391 1041
rect 1395 1042 1412 1045
rect 1444 1045 1830 1049
rect 1834 1045 1858 1049
rect 1862 1045 1888 1049
rect 1892 1045 1929 1049
rect 1480 1038 1806 1042
rect 1810 1038 1857 1042
rect 1861 1038 1907 1042
rect 1911 1038 1929 1042
rect 559 1023 873 1027
rect 877 1023 909 1027
rect 913 1023 976 1027
rect 980 1023 996 1027
rect 93 1015 126 1019
rect 130 1015 154 1019
rect 158 1015 184 1019
rect 188 1015 258 1019
rect 262 1015 286 1019
rect 290 1015 316 1019
rect 320 1015 390 1019
rect 394 1015 418 1019
rect 422 1015 448 1019
rect 452 1015 505 1019
rect 863 1016 897 1020
rect 901 1016 925 1020
rect 929 1016 955 1020
rect 959 1016 992 1020
rect 1029 1019 1032 1031
rect 1050 1019 1053 1031
rect 1066 1019 1069 1031
rect 1080 1022 1092 1025
rect 1108 1019 1111 1031
rect 1124 1019 1127 1031
rect 1145 1019 1148 1031
rect 1161 1019 1164 1031
rect 1182 1019 1185 1031
rect 1198 1019 1201 1031
rect 1212 1022 1224 1025
rect 1240 1019 1243 1031
rect 1256 1019 1259 1031
rect 1277 1019 1280 1031
rect 1293 1019 1296 1031
rect 1314 1019 1317 1031
rect 1330 1019 1333 1031
rect 1344 1022 1356 1025
rect 1372 1019 1375 1031
rect 1388 1019 1391 1031
rect 1409 1019 1412 1031
rect 1803 1031 1924 1034
rect 1492 1023 1806 1027
rect 1810 1023 1842 1027
rect 1846 1023 1909 1027
rect 1913 1023 1929 1027
rect 93 1008 102 1012
rect 106 1008 153 1012
rect 157 1008 203 1012
rect 207 1008 234 1012
rect 238 1008 285 1012
rect 289 1008 335 1012
rect 339 1008 366 1012
rect 370 1008 417 1012
rect 421 1008 467 1012
rect 471 1008 541 1012
rect 867 1006 870 1016
rect 888 1006 891 1016
rect 904 1006 907 1016
rect 918 1009 923 1013
rect 927 1009 934 1013
rect 946 1006 949 1016
rect 962 1006 965 1016
rect 983 1006 986 1016
rect 1026 1015 1059 1019
rect 1063 1015 1087 1019
rect 1091 1015 1117 1019
rect 1121 1015 1191 1019
rect 1195 1015 1219 1019
rect 1223 1015 1249 1019
rect 1253 1015 1323 1019
rect 1327 1015 1351 1019
rect 1355 1015 1381 1019
rect 1385 1015 1438 1019
rect 1796 1016 1830 1020
rect 1834 1016 1858 1020
rect 1862 1016 1888 1020
rect 1892 1016 1925 1020
rect 1026 1008 1035 1012
rect 1039 1008 1086 1012
rect 1090 1008 1136 1012
rect 1140 1008 1167 1012
rect 1171 1008 1218 1012
rect 1222 1008 1268 1012
rect 1272 1008 1299 1012
rect 1303 1008 1350 1012
rect 1354 1008 1400 1012
rect 1404 1008 1474 1012
rect 1800 1006 1803 1016
rect 1821 1006 1824 1016
rect 1837 1006 1840 1016
rect 1851 1009 1856 1013
rect 1860 1009 1867 1013
rect 1879 1006 1882 1016
rect 1895 1006 1898 1016
rect 1916 1006 1919 1016
rect 99 1001 484 1004
rect 93 993 102 997
rect 106 993 138 997
rect 142 993 205 997
rect 209 993 234 997
rect 238 993 270 997
rect 274 993 337 997
rect 341 993 366 997
rect 370 993 402 997
rect 406 993 469 997
rect 473 993 553 997
rect 93 986 126 990
rect 130 986 154 990
rect 158 986 184 990
rect 188 986 221 990
rect 225 986 258 990
rect 262 986 286 990
rect 290 986 316 990
rect 320 986 353 990
rect 357 986 390 990
rect 394 986 418 990
rect 422 986 448 990
rect 452 986 485 990
rect 489 986 493 990
rect 884 992 889 995
rect 893 992 917 995
rect 1032 1001 1417 1004
rect 942 992 949 995
rect 953 992 975 995
rect 1026 993 1035 997
rect 1039 993 1071 997
rect 1075 993 1138 997
rect 1142 993 1167 997
rect 1171 993 1203 997
rect 1207 993 1270 997
rect 1274 993 1299 997
rect 1303 993 1335 997
rect 1339 993 1402 997
rect 1406 993 1486 997
rect 96 976 99 986
rect 117 976 120 986
rect 133 976 136 986
rect 147 979 152 983
rect 156 979 163 983
rect 175 976 178 986
rect 191 976 194 986
rect 212 976 215 986
rect 228 976 231 986
rect 249 976 252 986
rect 265 976 268 986
rect 279 979 284 983
rect 288 979 295 983
rect 307 976 310 986
rect 323 976 326 986
rect 344 976 347 986
rect 360 976 363 986
rect 381 976 384 986
rect 397 976 400 986
rect 411 979 416 983
rect 420 979 427 983
rect 439 976 442 986
rect 455 976 458 986
rect 476 976 479 986
rect 900 982 907 985
rect 911 986 930 989
rect 113 962 118 965
rect 122 962 146 965
rect 171 962 178 965
rect 182 962 204 965
rect 224 962 231 965
rect 245 962 250 965
rect 254 962 278 965
rect 303 962 310 965
rect 314 962 336 965
rect 356 962 363 965
rect 377 962 382 965
rect 386 962 410 965
rect 435 962 442 965
rect 446 962 468 965
rect 930 979 933 985
rect 958 982 965 985
rect 969 986 984 989
rect 995 984 1006 988
rect 1026 986 1059 990
rect 1063 986 1087 990
rect 1091 986 1117 990
rect 1121 986 1154 990
rect 1158 986 1191 990
rect 1195 986 1219 990
rect 1223 986 1249 990
rect 1253 986 1286 990
rect 1290 986 1323 990
rect 1327 986 1351 990
rect 1355 986 1381 990
rect 1385 986 1418 990
rect 1422 986 1426 990
rect 1817 992 1822 995
rect 1826 992 1850 995
rect 1875 992 1882 995
rect 1886 992 1908 995
rect 1029 976 1032 986
rect 1050 976 1053 986
rect 1066 976 1069 986
rect 1080 979 1085 983
rect 1089 979 1096 983
rect 1108 976 1111 986
rect 1124 976 1127 986
rect 1145 976 1148 986
rect 1161 976 1164 986
rect 1182 976 1185 986
rect 1198 976 1201 986
rect 1212 979 1217 983
rect 1221 979 1228 983
rect 1240 976 1243 986
rect 1256 976 1259 986
rect 1277 976 1280 986
rect 1293 976 1296 986
rect 1314 976 1317 986
rect 1330 976 1333 986
rect 1344 979 1349 983
rect 1353 979 1360 983
rect 1372 976 1375 986
rect 1388 976 1391 986
rect 1409 976 1412 986
rect 1833 982 1840 985
rect 1844 986 1863 989
rect 867 963 870 975
rect 888 963 891 975
rect 904 963 907 975
rect 918 966 930 969
rect 946 963 949 975
rect 962 963 965 975
rect 983 963 986 975
rect 129 952 136 955
rect 140 956 159 959
rect 159 949 162 955
rect 187 952 194 955
rect 198 956 213 959
rect 261 952 268 955
rect 272 956 291 959
rect 291 949 294 955
rect 319 952 326 955
rect 330 956 345 959
rect 393 952 400 955
rect 404 956 423 959
rect 423 949 426 955
rect 451 952 458 955
rect 462 956 479 959
rect 511 959 897 963
rect 901 959 925 963
rect 929 959 955 963
rect 959 959 996 963
rect 1046 962 1051 965
rect 1055 962 1079 965
rect 1104 962 1111 965
rect 1115 962 1137 965
rect 1157 962 1164 965
rect 1178 962 1183 965
rect 1187 962 1211 965
rect 1236 962 1243 965
rect 1247 962 1269 965
rect 1289 962 1296 965
rect 1310 962 1315 965
rect 1319 962 1343 965
rect 1368 962 1375 965
rect 1379 962 1401 965
rect 1863 979 1866 985
rect 1891 982 1898 985
rect 1902 986 1917 989
rect 1928 984 1939 988
rect 1800 963 1803 975
rect 1821 963 1824 975
rect 1837 963 1840 975
rect 1851 966 1863 969
rect 1879 963 1882 975
rect 1895 963 1898 975
rect 1916 963 1919 975
rect 547 952 873 956
rect 877 952 924 956
rect 928 952 974 956
rect 978 952 996 956
rect 1062 952 1069 955
rect 1073 956 1092 959
rect 1092 949 1095 955
rect 1120 952 1127 955
rect 1131 956 1146 959
rect 1194 952 1201 955
rect 1205 956 1224 959
rect 1224 949 1227 955
rect 1252 952 1259 955
rect 1263 956 1278 959
rect 1326 952 1333 955
rect 1337 956 1356 959
rect 1356 949 1359 955
rect 1384 952 1391 955
rect 1395 956 1412 959
rect 1444 959 1830 963
rect 1834 959 1858 963
rect 1862 959 1888 963
rect 1892 959 1929 963
rect 1480 952 1806 956
rect 1810 952 1857 956
rect 1861 952 1907 956
rect 1911 952 1929 956
rect 96 933 99 945
rect 117 933 120 945
rect 133 933 136 945
rect 147 936 159 939
rect 175 933 178 945
rect 191 933 194 945
rect 212 933 215 945
rect 228 933 231 945
rect 249 933 252 945
rect 265 933 268 945
rect 279 936 291 939
rect 307 933 310 945
rect 323 933 326 945
rect 344 933 347 945
rect 360 933 363 945
rect 381 933 384 945
rect 397 933 400 945
rect 411 936 423 939
rect 439 933 442 945
rect 455 933 458 945
rect 476 933 479 945
rect 1029 933 1032 945
rect 1050 933 1053 945
rect 1066 933 1069 945
rect 1080 936 1092 939
rect 1108 933 1111 945
rect 1124 933 1127 945
rect 1145 933 1148 945
rect 1161 933 1164 945
rect 1182 933 1185 945
rect 1198 933 1201 945
rect 1212 936 1224 939
rect 1240 933 1243 945
rect 1256 933 1259 945
rect 1277 933 1280 945
rect 1293 933 1296 945
rect 1314 933 1317 945
rect 1330 933 1333 945
rect 1344 936 1356 939
rect 1372 933 1375 945
rect 1388 933 1391 945
rect 1409 933 1412 945
rect 93 929 126 933
rect 130 929 154 933
rect 158 929 184 933
rect 188 929 258 933
rect 262 929 286 933
rect 290 929 316 933
rect 320 929 390 933
rect 394 929 418 933
rect 422 929 448 933
rect 452 929 505 933
rect 1026 929 1059 933
rect 1063 929 1087 933
rect 1091 929 1117 933
rect 1121 929 1191 933
rect 1195 929 1219 933
rect 1223 929 1249 933
rect 1253 929 1323 933
rect 1327 929 1351 933
rect 1355 929 1381 933
rect 1385 929 1438 933
rect 93 922 102 926
rect 106 922 153 926
rect 157 922 203 926
rect 207 922 234 926
rect 238 922 285 926
rect 289 922 335 926
rect 339 922 366 926
rect 370 922 417 926
rect 421 922 467 926
rect 471 922 541 926
rect 1026 922 1035 926
rect 1039 922 1086 926
rect 1090 922 1136 926
rect 1140 922 1167 926
rect 1171 922 1218 926
rect 1222 922 1268 926
rect 1272 922 1299 926
rect 1303 922 1350 926
rect 1354 922 1400 926
rect 1404 922 1474 926
rect 99 916 484 919
rect 1032 916 1417 919
rect 224 909 328 912
rect 1157 909 1261 912
rect 340 901 344 905
rect 348 901 352 905
rect 1273 901 1277 905
rect 1281 901 1285 905
rect 83 890 328 894
rect 332 890 348 894
rect 364 890 1013 894
rect 1017 890 1261 894
rect 1265 890 1281 894
rect 1297 890 1946 894
rect 1950 890 2028 894
rect 356 883 484 886
rect 1289 883 1417 886
rect 371 876 484 879
rect 1304 876 1417 879
rect 340 867 344 871
rect 348 867 352 871
rect 1273 867 1277 871
rect 1281 867 1285 871
rect 224 860 328 863
rect 1157 860 1261 863
rect 93 853 102 857
rect 106 853 138 857
rect 142 853 205 857
rect 209 853 234 857
rect 238 853 270 857
rect 274 853 337 857
rect 341 853 366 857
rect 370 853 402 857
rect 406 853 469 857
rect 473 853 553 857
rect 1026 853 1035 857
rect 1039 853 1071 857
rect 1075 853 1138 857
rect 1142 853 1167 857
rect 1171 853 1203 857
rect 1207 853 1270 857
rect 1274 853 1299 857
rect 1303 853 1335 857
rect 1339 853 1402 857
rect 1406 853 1486 857
rect 93 846 126 850
rect 130 846 154 850
rect 158 846 184 850
rect 188 846 221 850
rect 225 846 258 850
rect 262 846 286 850
rect 290 846 316 850
rect 320 846 353 850
rect 357 846 390 850
rect 394 846 418 850
rect 422 846 448 850
rect 452 846 485 850
rect 489 846 493 850
rect 1026 846 1059 850
rect 1063 846 1087 850
rect 1091 846 1117 850
rect 1121 846 1154 850
rect 1158 846 1191 850
rect 1195 846 1219 850
rect 1223 846 1249 850
rect 1253 846 1286 850
rect 1290 846 1323 850
rect 1327 846 1351 850
rect 1355 846 1381 850
rect 1385 846 1418 850
rect 1422 846 1426 850
rect 96 836 99 846
rect 117 836 120 846
rect 133 836 136 846
rect 147 839 152 843
rect 156 839 163 843
rect 175 836 178 846
rect 191 836 194 846
rect 212 836 215 846
rect 228 836 231 846
rect 249 836 252 846
rect 265 836 268 846
rect 279 839 284 843
rect 288 839 295 843
rect 307 836 310 846
rect 323 836 326 846
rect 344 836 347 846
rect 360 836 363 846
rect 381 836 384 846
rect 397 836 400 846
rect 411 839 416 843
rect 420 839 427 843
rect 439 836 442 846
rect 455 836 458 846
rect 476 836 479 846
rect 1029 836 1032 846
rect 1050 836 1053 846
rect 1066 836 1069 846
rect 1080 839 1085 843
rect 1089 839 1096 843
rect 1108 836 1111 846
rect 1124 836 1127 846
rect 1145 836 1148 846
rect 1161 836 1164 846
rect 1182 836 1185 846
rect 1198 836 1201 846
rect 1212 839 1217 843
rect 1221 839 1228 843
rect 1240 836 1243 846
rect 1256 836 1259 846
rect 1277 836 1280 846
rect 1293 836 1296 846
rect 1314 836 1317 846
rect 1330 836 1333 846
rect 1344 839 1349 843
rect 1353 839 1360 843
rect 1372 836 1375 846
rect 1388 836 1391 846
rect 1409 836 1412 846
rect 113 822 118 825
rect 122 822 146 825
rect 171 822 178 825
rect 182 822 204 825
rect 224 822 231 825
rect 245 822 250 825
rect 254 822 278 825
rect 303 822 310 825
rect 314 822 336 825
rect 356 822 363 825
rect 377 822 382 825
rect 386 822 410 825
rect 435 822 442 825
rect 446 822 468 825
rect 129 812 136 815
rect 140 816 159 819
rect 159 809 162 815
rect 187 812 194 815
rect 198 816 213 819
rect 261 812 268 815
rect 272 816 291 819
rect 291 809 294 815
rect 319 812 326 815
rect 330 816 345 819
rect 393 812 400 815
rect 404 816 423 819
rect 423 809 426 815
rect 451 812 458 815
rect 462 816 479 819
rect 1046 822 1051 825
rect 1055 822 1079 825
rect 1104 822 1111 825
rect 1115 822 1137 825
rect 1157 822 1164 825
rect 1178 822 1183 825
rect 1187 822 1211 825
rect 1236 822 1243 825
rect 1247 822 1269 825
rect 1289 822 1296 825
rect 1310 822 1315 825
rect 1319 822 1343 825
rect 1368 822 1375 825
rect 1379 822 1401 825
rect 1062 812 1069 815
rect 1073 816 1092 819
rect 1092 809 1095 815
rect 1120 812 1127 815
rect 1131 816 1146 819
rect 1194 812 1201 815
rect 1205 816 1224 819
rect 1224 809 1227 815
rect 1252 812 1259 815
rect 1263 816 1278 819
rect 1326 812 1333 815
rect 1337 816 1356 819
rect 1356 809 1359 815
rect 1384 812 1391 815
rect 1395 816 1412 819
rect 96 793 99 805
rect 117 793 120 805
rect 133 793 136 805
rect 147 796 159 799
rect 175 793 178 805
rect 191 793 194 805
rect 212 793 215 805
rect 228 793 231 805
rect 249 793 252 805
rect 265 793 268 805
rect 279 796 291 799
rect 307 793 310 805
rect 323 793 326 805
rect 344 793 347 805
rect 360 793 363 805
rect 381 793 384 805
rect 397 793 400 805
rect 411 796 423 799
rect 439 793 442 805
rect 455 793 458 805
rect 476 793 479 805
rect 1029 793 1032 805
rect 1050 793 1053 805
rect 1066 793 1069 805
rect 1080 796 1092 799
rect 1108 793 1111 805
rect 1124 793 1127 805
rect 1145 793 1148 805
rect 1161 793 1164 805
rect 1182 793 1185 805
rect 1198 793 1201 805
rect 1212 796 1224 799
rect 1240 793 1243 805
rect 1256 793 1259 805
rect 1277 793 1280 805
rect 1293 793 1296 805
rect 1314 793 1317 805
rect 1330 793 1333 805
rect 1344 796 1356 799
rect 1372 793 1375 805
rect 1388 793 1391 805
rect 1409 793 1412 805
rect 93 789 126 793
rect 130 789 154 793
rect 158 789 184 793
rect 188 789 258 793
rect 262 789 286 793
rect 290 789 316 793
rect 320 789 390 793
rect 394 789 418 793
rect 422 789 448 793
rect 452 789 505 793
rect 1026 789 1059 793
rect 1063 789 1087 793
rect 1091 789 1117 793
rect 1121 789 1191 793
rect 1195 789 1219 793
rect 1223 789 1249 793
rect 1253 789 1323 793
rect 1327 789 1351 793
rect 1355 789 1381 793
rect 1385 789 1438 793
rect 93 782 102 786
rect 106 782 153 786
rect 157 782 203 786
rect 207 782 234 786
rect 238 782 285 786
rect 289 782 335 786
rect 339 782 366 786
rect 370 782 417 786
rect 421 782 467 786
rect 471 782 541 786
rect 1026 782 1035 786
rect 1039 782 1086 786
rect 1090 782 1136 786
rect 1140 782 1167 786
rect 1171 782 1218 786
rect 1222 782 1268 786
rect 1272 782 1299 786
rect 1303 782 1350 786
rect 1354 782 1400 786
rect 1404 782 1474 786
rect 559 774 574 778
rect 578 774 610 778
rect 614 774 677 778
rect 681 774 706 778
rect 710 774 742 778
rect 746 774 809 778
rect 813 774 838 778
rect 842 774 874 778
rect 878 774 941 778
rect 945 774 970 778
rect 974 774 1006 778
rect 1010 774 1073 778
rect 1077 774 1093 778
rect 1492 774 1507 778
rect 1511 774 1543 778
rect 1547 774 1610 778
rect 1614 774 1639 778
rect 1643 774 1675 778
rect 1679 774 1742 778
rect 1746 774 1771 778
rect 1775 774 1807 778
rect 1811 774 1874 778
rect 1878 774 1903 778
rect 1907 774 1939 778
rect 1943 774 2006 778
rect 2010 774 2026 778
rect 499 767 598 771
rect 602 767 626 771
rect 630 767 656 771
rect 660 767 693 771
rect 697 767 730 771
rect 734 767 758 771
rect 762 767 788 771
rect 792 767 825 771
rect 829 767 862 771
rect 866 767 890 771
rect 894 767 920 771
rect 924 767 957 771
rect 961 767 994 771
rect 998 767 1022 771
rect 1026 767 1052 771
rect 1056 767 1089 771
rect 1432 767 1531 771
rect 1535 767 1559 771
rect 1563 767 1589 771
rect 1593 767 1626 771
rect 1630 767 1663 771
rect 1667 767 1691 771
rect 1695 767 1721 771
rect 1725 767 1758 771
rect 1762 767 1795 771
rect 1799 767 1823 771
rect 1827 767 1853 771
rect 1857 767 1890 771
rect 1894 767 1927 771
rect 1931 767 1955 771
rect 1959 767 1985 771
rect 1989 767 2022 771
rect 568 757 571 767
rect 589 757 592 767
rect 605 757 608 767
rect 619 760 624 764
rect 628 760 635 764
rect 647 757 650 767
rect 663 757 666 767
rect 684 757 687 767
rect 700 757 703 767
rect 721 757 724 767
rect 737 757 740 767
rect 751 760 756 764
rect 760 760 767 764
rect 779 757 782 767
rect 795 757 798 767
rect 816 757 819 767
rect 832 757 835 767
rect 853 757 856 767
rect 869 757 872 767
rect 883 760 888 764
rect 892 760 899 764
rect 911 757 914 767
rect 927 757 930 767
rect 948 757 951 767
rect 964 757 967 767
rect 985 757 988 767
rect 1001 757 1004 767
rect 1015 760 1020 764
rect 1024 760 1031 764
rect 1043 757 1046 767
rect 1059 757 1062 767
rect 1080 757 1083 767
rect 1501 757 1504 767
rect 1522 757 1525 767
rect 1538 757 1541 767
rect 1552 760 1557 764
rect 1561 760 1568 764
rect 1580 757 1583 767
rect 1596 757 1599 767
rect 1617 757 1620 767
rect 1633 757 1636 767
rect 1654 757 1657 767
rect 1670 757 1673 767
rect 1684 760 1689 764
rect 1693 760 1700 764
rect 1712 757 1715 767
rect 1728 757 1731 767
rect 1749 757 1752 767
rect 1765 757 1768 767
rect 1786 757 1789 767
rect 1802 757 1805 767
rect 1816 760 1821 764
rect 1825 760 1832 764
rect 1844 757 1847 767
rect 1860 757 1863 767
rect 1881 757 1884 767
rect 1897 757 1900 767
rect 1918 757 1921 767
rect 1934 757 1937 767
rect 1948 760 1953 764
rect 1957 760 1964 764
rect 1976 757 1979 767
rect 1992 757 1995 767
rect 2013 757 2016 767
rect 225 741 234 745
rect 238 741 270 745
rect 274 741 337 745
rect 341 741 553 745
rect 585 743 590 746
rect 594 743 618 746
rect 643 743 650 746
rect 654 743 676 746
rect 225 734 258 738
rect 262 734 286 738
rect 290 734 316 738
rect 320 734 353 738
rect 357 734 493 738
rect 228 724 231 734
rect 249 724 252 734
rect 265 724 268 734
rect 279 727 284 731
rect 288 727 295 731
rect 307 724 310 734
rect 323 724 326 734
rect 344 724 347 734
rect 601 733 608 736
rect 612 737 631 740
rect 631 730 634 736
rect 659 733 666 736
rect 670 737 687 740
rect 717 743 722 746
rect 726 743 750 746
rect 775 743 782 746
rect 786 743 808 746
rect 733 733 740 736
rect 744 737 763 740
rect 763 730 766 736
rect 791 733 798 736
rect 802 737 819 740
rect 849 743 854 746
rect 858 743 882 746
rect 907 743 914 746
rect 918 743 940 746
rect 865 733 872 736
rect 876 737 895 740
rect 895 730 898 736
rect 923 733 930 736
rect 934 737 951 740
rect 981 743 986 746
rect 990 743 1014 746
rect 1039 743 1046 746
rect 1050 743 1072 746
rect 1158 741 1167 745
rect 1171 741 1203 745
rect 1207 741 1270 745
rect 1274 741 1486 745
rect 997 733 1004 736
rect 1008 737 1027 740
rect 223 707 232 711
rect 245 710 250 713
rect 254 710 278 713
rect 303 710 310 713
rect 314 710 336 713
rect 568 714 571 726
rect 589 714 592 726
rect 605 714 608 726
rect 619 717 631 720
rect 647 714 650 726
rect 663 714 666 726
rect 684 714 687 726
rect 700 714 703 726
rect 721 714 724 726
rect 737 714 740 726
rect 751 717 763 720
rect 779 714 782 726
rect 795 714 798 726
rect 816 714 819 726
rect 832 714 835 726
rect 853 714 856 726
rect 869 714 872 726
rect 883 717 895 720
rect 911 714 914 726
rect 927 714 930 726
rect 948 714 951 726
rect 1027 730 1030 736
rect 1055 733 1062 736
rect 1066 737 1083 740
rect 1518 743 1523 746
rect 1527 743 1551 746
rect 1576 743 1583 746
rect 1587 743 1609 746
rect 1158 734 1191 738
rect 1195 734 1219 738
rect 1223 734 1249 738
rect 1253 734 1286 738
rect 1290 734 1426 738
rect 964 714 967 726
rect 985 714 988 726
rect 1001 714 1004 726
rect 1015 717 1027 720
rect 1043 714 1046 726
rect 1059 714 1062 726
rect 1080 714 1083 726
rect 1161 724 1164 734
rect 1182 724 1185 734
rect 1198 724 1201 734
rect 1212 727 1217 731
rect 1221 727 1228 731
rect 1240 724 1243 734
rect 1256 724 1259 734
rect 1277 724 1280 734
rect 1534 733 1541 736
rect 1545 737 1564 740
rect 1564 730 1567 736
rect 1592 733 1599 736
rect 1603 737 1620 740
rect 1650 743 1655 746
rect 1659 743 1683 746
rect 1708 743 1715 746
rect 1719 743 1741 746
rect 1666 733 1673 736
rect 1677 737 1696 740
rect 1696 730 1699 736
rect 1724 733 1731 736
rect 1735 737 1752 740
rect 1782 743 1787 746
rect 1791 743 1815 746
rect 1840 743 1847 746
rect 1851 743 1873 746
rect 1798 733 1805 736
rect 1809 737 1828 740
rect 1828 730 1831 736
rect 1856 733 1863 736
rect 1867 737 1884 740
rect 1914 743 1919 746
rect 1923 743 1947 746
rect 1972 743 1979 746
rect 1983 743 2005 746
rect 1930 733 1937 736
rect 1941 737 1960 740
rect 511 710 598 714
rect 602 710 626 714
rect 630 710 656 714
rect 660 710 730 714
rect 734 710 758 714
rect 762 710 788 714
rect 792 710 862 714
rect 866 710 890 714
rect 894 710 920 714
rect 924 710 994 714
rect 998 710 1022 714
rect 1026 710 1052 714
rect 1056 710 1093 714
rect 261 700 268 703
rect 272 704 291 707
rect 291 697 294 703
rect 319 700 326 703
rect 330 704 345 707
rect 1156 707 1165 711
rect 1178 710 1183 713
rect 1187 710 1211 713
rect 1236 710 1243 713
rect 1247 710 1269 713
rect 1501 714 1504 726
rect 1522 714 1525 726
rect 1538 714 1541 726
rect 1552 717 1564 720
rect 1580 714 1583 726
rect 1596 714 1599 726
rect 1617 714 1620 726
rect 1633 714 1636 726
rect 1654 714 1657 726
rect 1670 714 1673 726
rect 1684 717 1696 720
rect 1712 714 1715 726
rect 1728 714 1731 726
rect 1749 714 1752 726
rect 1765 714 1768 726
rect 1786 714 1789 726
rect 1802 714 1805 726
rect 1816 717 1828 720
rect 1844 714 1847 726
rect 1860 714 1863 726
rect 1881 714 1884 726
rect 1960 730 1963 736
rect 1988 733 1995 736
rect 1999 737 2016 740
rect 1897 714 1900 726
rect 1918 714 1921 726
rect 1934 714 1937 726
rect 1948 717 1960 720
rect 1976 714 1979 726
rect 1992 714 1995 726
rect 2013 714 2016 726
rect 1444 710 1531 714
rect 1535 710 1559 714
rect 1563 710 1589 714
rect 1593 710 1663 714
rect 1667 710 1691 714
rect 1695 710 1721 714
rect 1725 710 1795 714
rect 1799 710 1823 714
rect 1827 710 1853 714
rect 1857 710 1927 714
rect 1931 710 1955 714
rect 1959 710 1985 714
rect 1989 710 2026 714
rect 547 703 574 707
rect 578 703 625 707
rect 629 703 675 707
rect 679 703 706 707
rect 710 703 757 707
rect 761 703 807 707
rect 811 703 838 707
rect 842 703 889 707
rect 893 703 939 707
rect 943 703 970 707
rect 974 703 1021 707
rect 1025 703 1071 707
rect 1075 703 1093 707
rect 1194 700 1201 703
rect 1205 704 1224 707
rect 228 681 231 693
rect 249 681 252 693
rect 265 681 268 693
rect 279 684 291 687
rect 307 681 310 693
rect 323 681 326 693
rect 344 681 347 693
rect 499 690 572 694
rect 576 690 588 694
rect 592 690 606 694
rect 610 690 617 694
rect 621 690 623 694
rect 627 690 642 694
rect 646 690 679 694
rect 683 690 684 694
rect 688 690 696 694
rect 700 690 724 694
rect 728 690 740 694
rect 744 690 764 694
rect 768 690 818 694
rect 822 690 845 694
rect 849 690 899 694
rect 903 690 922 694
rect 1224 697 1227 703
rect 1252 700 1259 703
rect 1263 704 1278 707
rect 1480 703 1507 707
rect 1511 703 1558 707
rect 1562 703 1608 707
rect 1612 703 1639 707
rect 1643 703 1690 707
rect 1694 703 1740 707
rect 1744 703 1771 707
rect 1775 703 1822 707
rect 1826 703 1872 707
rect 1876 703 1903 707
rect 1907 703 1954 707
rect 1958 703 2004 707
rect 2008 703 2026 707
rect 535 683 599 687
rect 603 683 630 687
rect 634 683 652 687
rect 656 683 717 687
rect 721 683 735 687
rect 747 686 750 690
rect 225 677 258 681
rect 262 677 286 681
rect 290 677 316 681
rect 320 677 505 681
rect 225 670 234 674
rect 238 670 285 674
rect 289 670 335 674
rect 339 670 541 674
rect 642 676 645 680
rect 669 676 670 680
rect 714 676 716 680
rect 756 673 759 678
rect 771 680 774 690
rect 801 686 804 690
rect 828 686 831 690
rect 223 654 239 658
rect 348 656 352 660
rect 364 656 368 660
rect 372 656 574 660
rect 582 659 585 665
rect 589 659 592 665
rect 582 656 592 659
rect 582 651 585 656
rect 231 647 235 651
rect 247 647 368 651
rect 589 651 592 656
rect 598 661 601 665
rect 598 657 600 661
rect 604 657 606 661
rect 614 660 617 665
rect 642 662 645 665
rect 614 658 625 660
rect 598 651 601 657
rect 614 656 620 658
rect 614 651 617 656
rect 624 656 625 658
rect 643 658 645 662
rect 642 651 645 658
rect 745 669 748 672
rect 787 669 790 672
rect 658 661 661 665
rect 668 661 671 665
rect 668 657 677 661
rect 689 660 692 665
rect 714 661 717 665
rect 658 651 661 657
rect 668 651 671 657
rect 689 656 690 660
rect 694 656 697 659
rect 716 657 717 661
rect 732 660 735 665
rect 756 664 759 669
rect 764 665 775 668
rect 787 666 795 669
rect 689 651 692 656
rect 714 651 717 657
rect 732 651 735 656
rect 218 639 234 643
rect 238 639 301 643
rect 305 639 337 643
rect 341 639 553 643
rect 634 638 635 642
rect 659 639 660 643
rect 706 638 707 642
rect 222 632 255 636
rect 259 632 285 636
rect 289 632 313 636
rect 317 632 493 636
rect 228 622 231 632
rect 249 622 252 632
rect 265 622 268 632
rect 280 625 287 629
rect 291 625 296 629
rect 307 622 310 632
rect 323 622 326 632
rect 344 622 347 632
rect 523 631 587 635
rect 591 631 646 635
rect 650 631 671 635
rect 675 631 702 635
rect 706 631 735 635
rect 747 628 750 660
rect 764 659 767 665
rect 787 660 790 666
rect 799 661 802 664
rect 810 664 813 678
rect 837 673 840 678
rect 852 680 855 690
rect 882 686 885 690
rect 821 669 822 672
rect 826 669 829 672
rect 1161 681 1164 693
rect 1182 681 1185 693
rect 1198 681 1201 693
rect 1212 684 1224 687
rect 1240 681 1243 693
rect 1256 681 1259 693
rect 1277 681 1280 693
rect 1432 690 1505 694
rect 1509 690 1521 694
rect 1525 690 1539 694
rect 1543 690 1550 694
rect 1554 690 1556 694
rect 1560 690 1575 694
rect 1579 690 1612 694
rect 1616 690 1617 694
rect 1621 690 1629 694
rect 1633 690 1657 694
rect 1661 690 1673 694
rect 1677 690 1697 694
rect 1701 690 1751 694
rect 1755 690 1778 694
rect 1782 690 1832 694
rect 1836 690 1855 694
rect 1468 683 1532 687
rect 1536 683 1563 687
rect 1567 683 1585 687
rect 1589 683 1650 687
rect 1654 683 1668 687
rect 1680 686 1683 690
rect 868 669 871 672
rect 810 661 818 664
rect 837 664 840 669
rect 810 656 813 661
rect 818 657 822 661
rect 845 665 856 668
rect 868 666 876 669
rect 762 650 767 655
rect 771 628 774 656
rect 801 628 804 652
rect 828 628 831 660
rect 845 659 848 665
rect 868 660 871 666
rect 880 661 883 664
rect 891 664 894 678
rect 1158 677 1191 681
rect 1195 677 1219 681
rect 1223 677 1249 681
rect 1253 677 1438 681
rect 1158 670 1167 674
rect 1171 670 1218 674
rect 1222 670 1268 674
rect 1272 670 1474 674
rect 1575 676 1578 680
rect 1602 676 1603 680
rect 1647 676 1649 680
rect 1689 673 1692 678
rect 1704 680 1707 690
rect 1734 686 1737 690
rect 1761 686 1764 690
rect 891 661 903 664
rect 891 656 894 661
rect 843 650 848 655
rect 852 628 855 656
rect 1156 654 1172 658
rect 1281 656 1285 660
rect 1297 656 1301 660
rect 1305 656 1507 660
rect 1515 659 1518 665
rect 1522 659 1525 665
rect 1515 656 1525 659
rect 882 628 885 652
rect 1515 651 1518 656
rect 1164 647 1168 651
rect 1180 647 1301 651
rect 1522 651 1525 656
rect 1531 661 1534 665
rect 1531 657 1533 661
rect 1537 657 1539 661
rect 1547 660 1550 665
rect 1575 662 1578 665
rect 1547 658 1558 660
rect 1531 651 1534 657
rect 1547 656 1553 658
rect 1547 651 1550 656
rect 1557 656 1558 658
rect 1576 658 1578 662
rect 1575 651 1578 658
rect 1678 669 1681 672
rect 1720 669 1723 672
rect 1591 661 1594 665
rect 1601 661 1604 665
rect 1601 657 1610 661
rect 1622 660 1625 665
rect 1647 661 1650 665
rect 1591 651 1594 657
rect 1601 651 1604 657
rect 1622 656 1623 660
rect 1627 656 1630 659
rect 1649 657 1650 661
rect 1665 660 1668 665
rect 1689 664 1692 669
rect 1697 665 1708 668
rect 1720 666 1728 669
rect 1622 651 1625 656
rect 1647 651 1650 657
rect 1665 651 1668 656
rect 1151 639 1167 643
rect 1171 639 1234 643
rect 1238 639 1270 643
rect 1274 639 1486 643
rect 1567 638 1568 642
rect 1592 639 1593 643
rect 1639 638 1640 642
rect 1155 632 1188 636
rect 1192 632 1218 636
rect 1222 632 1246 636
rect 1250 632 1426 636
rect 511 624 573 628
rect 577 624 579 628
rect 583 624 587 628
rect 591 624 605 628
rect 609 624 614 628
rect 618 624 623 628
rect 627 624 646 628
rect 650 624 680 628
rect 684 624 695 628
rect 699 624 723 628
rect 727 624 740 628
rect 744 624 764 628
rect 768 624 818 628
rect 825 624 845 628
rect 849 624 899 628
rect 239 608 261 611
rect 265 608 272 611
rect 523 617 587 621
rect 591 617 646 621
rect 650 617 671 621
rect 675 617 702 621
rect 706 617 735 621
rect 297 608 321 611
rect 325 608 330 611
rect 634 610 635 614
rect 659 609 660 613
rect 706 610 707 614
rect 343 605 352 609
rect 230 602 245 605
rect 284 602 303 605
rect 249 598 256 601
rect 281 595 284 601
rect 307 598 314 601
rect 582 596 585 601
rect 589 596 592 601
rect 572 593 574 596
rect 582 593 592 596
rect 228 579 231 591
rect 249 579 252 591
rect 265 579 268 591
rect 284 582 296 585
rect 307 579 310 591
rect 323 579 326 591
rect 344 579 347 591
rect 582 587 585 593
rect 589 587 592 593
rect 598 595 601 601
rect 614 596 617 601
rect 598 591 600 595
rect 604 591 606 595
rect 614 594 620 596
rect 624 594 625 596
rect 614 592 625 594
rect 642 594 645 601
rect 598 587 601 591
rect 614 587 617 592
rect 643 590 645 594
rect 642 587 645 590
rect 658 595 661 601
rect 668 595 671 601
rect 689 596 692 601
rect 668 591 677 595
rect 689 592 690 596
rect 694 593 697 596
rect 714 595 717 601
rect 732 596 735 601
rect 771 604 774 624
rect 852 604 855 624
rect 1161 622 1164 632
rect 1182 622 1185 632
rect 1198 622 1201 632
rect 1213 625 1220 629
rect 1224 625 1229 629
rect 1240 622 1243 632
rect 1256 622 1259 632
rect 1277 622 1280 632
rect 1456 631 1520 635
rect 1524 631 1579 635
rect 1583 631 1604 635
rect 1608 631 1635 635
rect 1639 631 1668 635
rect 1680 628 1683 660
rect 1697 659 1700 665
rect 1720 660 1723 666
rect 1732 661 1735 664
rect 1743 664 1746 678
rect 1770 673 1773 678
rect 1785 680 1788 690
rect 1815 686 1818 690
rect 1754 669 1755 672
rect 1759 669 1762 672
rect 1801 669 1804 672
rect 1743 661 1751 664
rect 1770 664 1773 669
rect 1743 656 1746 661
rect 1751 657 1755 661
rect 1778 665 1789 668
rect 1801 666 1809 669
rect 1695 650 1700 655
rect 1704 628 1707 656
rect 1734 628 1737 652
rect 1761 628 1764 660
rect 1778 659 1781 665
rect 1801 660 1804 666
rect 1813 661 1816 664
rect 1824 664 1827 678
rect 1824 661 1836 664
rect 1824 656 1827 661
rect 1776 650 1781 655
rect 1785 628 1788 656
rect 1815 628 1818 652
rect 1444 624 1506 628
rect 1510 624 1512 628
rect 1516 624 1520 628
rect 1524 624 1538 628
rect 1542 624 1547 628
rect 1551 624 1556 628
rect 1560 624 1579 628
rect 1583 624 1613 628
rect 1617 624 1628 628
rect 1632 624 1656 628
rect 1660 624 1673 628
rect 1677 624 1697 628
rect 1701 624 1751 628
rect 1758 624 1778 628
rect 1782 624 1832 628
rect 1172 608 1194 611
rect 1198 608 1205 611
rect 1456 617 1520 621
rect 1524 617 1579 621
rect 1583 617 1604 621
rect 1608 617 1635 621
rect 1639 617 1668 621
rect 1230 608 1254 611
rect 1258 608 1263 611
rect 1567 610 1568 614
rect 1592 609 1593 613
rect 1639 610 1640 614
rect 1276 605 1285 609
rect 1163 602 1178 605
rect 658 587 661 591
rect 668 587 671 591
rect 689 587 692 592
rect 716 591 717 595
rect 714 587 717 591
rect 732 587 735 592
rect 762 591 767 596
rect 771 592 772 595
rect 787 594 790 600
rect 787 591 795 594
rect 842 591 847 596
rect 851 592 853 595
rect 868 594 871 600
rect 1217 602 1236 605
rect 1182 598 1189 601
rect 1214 595 1217 601
rect 868 591 876 594
rect 1240 598 1247 601
rect 1515 596 1518 601
rect 1522 596 1525 601
rect 1505 593 1507 596
rect 1515 593 1525 596
rect 787 588 790 591
rect 868 588 871 591
rect 218 575 255 579
rect 259 575 285 579
rect 289 575 313 579
rect 317 575 505 579
rect 642 572 645 576
rect 669 572 670 576
rect 714 572 716 576
rect 218 568 236 572
rect 240 568 286 572
rect 290 568 337 572
rect 341 568 541 572
rect 587 565 599 569
rect 603 565 630 569
rect 634 565 652 569
rect 656 565 717 569
rect 721 565 735 569
rect 771 562 774 580
rect 852 562 855 580
rect 1161 579 1164 591
rect 1182 579 1185 591
rect 1198 579 1201 591
rect 1217 582 1229 585
rect 1240 579 1243 591
rect 1256 579 1259 591
rect 1277 579 1280 591
rect 1515 587 1518 593
rect 1522 587 1525 593
rect 1531 595 1534 601
rect 1547 596 1550 601
rect 1531 591 1533 595
rect 1537 591 1539 595
rect 1547 594 1553 596
rect 1557 594 1558 596
rect 1547 592 1558 594
rect 1575 594 1578 601
rect 1531 587 1534 591
rect 1547 587 1550 592
rect 1576 590 1578 594
rect 1575 587 1578 590
rect 1591 595 1594 601
rect 1601 595 1604 601
rect 1622 596 1625 601
rect 1601 591 1610 595
rect 1622 592 1623 596
rect 1627 593 1630 596
rect 1647 595 1650 601
rect 1665 596 1668 601
rect 1704 604 1707 624
rect 1785 604 1788 624
rect 1591 587 1594 591
rect 1601 587 1604 591
rect 1622 587 1625 592
rect 1649 591 1650 595
rect 1647 587 1650 591
rect 1665 587 1668 592
rect 1695 591 1700 596
rect 1704 592 1705 595
rect 1720 594 1723 600
rect 1720 591 1728 594
rect 1775 591 1780 596
rect 1784 592 1786 595
rect 1801 594 1804 600
rect 1801 591 1809 594
rect 1720 588 1723 591
rect 1801 588 1804 591
rect 1151 575 1188 579
rect 1192 575 1218 579
rect 1222 575 1246 579
rect 1250 575 1438 579
rect 1575 572 1578 576
rect 1602 572 1603 576
rect 1647 572 1649 576
rect 1151 568 1169 572
rect 1173 568 1219 572
rect 1223 568 1270 572
rect 1274 568 1474 572
rect 1520 565 1532 569
rect 1536 565 1563 569
rect 1567 565 1585 569
rect 1589 565 1650 569
rect 1654 565 1668 569
rect 1704 562 1707 580
rect 1785 562 1788 580
rect 499 558 572 562
rect 576 558 588 562
rect 592 558 606 562
rect 610 558 617 562
rect 621 558 623 562
rect 627 558 642 562
rect 646 558 679 562
rect 683 558 684 562
rect 688 558 696 562
rect 700 558 724 562
rect 728 558 740 562
rect 744 558 764 562
rect 768 558 818 562
rect 822 558 845 562
rect 849 558 907 562
rect 911 558 922 562
rect 1432 558 1505 562
rect 1509 558 1521 562
rect 1525 558 1539 562
rect 1543 558 1550 562
rect 1554 558 1556 562
rect 1560 558 1575 562
rect 1579 558 1612 562
rect 1616 558 1617 562
rect 1621 558 1629 562
rect 1633 558 1657 562
rect 1661 558 1673 562
rect 1677 558 1697 562
rect 1701 558 1751 562
rect 1755 558 1778 562
rect 1782 558 1840 562
rect 1844 558 1855 562
rect 535 551 583 555
rect 587 551 599 555
rect 603 551 630 555
rect 634 551 652 555
rect 656 551 717 555
rect 721 551 735 555
rect 771 548 774 558
rect 801 554 804 558
rect 852 554 855 558
rect 642 544 645 548
rect 669 544 670 548
rect 714 544 716 548
rect 571 524 574 527
rect 582 527 585 533
rect 589 527 592 533
rect 582 524 592 527
rect 582 519 585 524
rect 589 519 592 524
rect 598 529 601 533
rect 598 525 600 529
rect 604 525 606 529
rect 614 528 617 533
rect 642 530 645 533
rect 614 526 625 528
rect 598 519 601 525
rect 614 524 620 526
rect 614 519 617 524
rect 624 524 625 526
rect 643 526 645 530
rect 642 519 645 526
rect 787 537 790 540
rect 658 529 661 533
rect 668 529 671 533
rect 668 525 677 529
rect 689 528 692 533
rect 714 529 717 533
rect 658 519 661 525
rect 668 519 671 525
rect 689 524 690 528
rect 694 524 697 527
rect 716 525 717 529
rect 732 528 735 533
rect 764 533 775 536
rect 787 534 795 537
rect 689 519 692 524
rect 714 519 717 525
rect 764 527 767 533
rect 787 528 790 534
rect 799 529 802 532
rect 810 532 813 546
rect 861 541 864 546
rect 876 548 879 558
rect 906 554 909 558
rect 845 537 846 540
rect 850 537 853 540
rect 1468 551 1516 555
rect 1520 551 1532 555
rect 1536 551 1563 555
rect 1567 551 1585 555
rect 1589 551 1650 555
rect 1654 551 1668 555
rect 1704 548 1707 558
rect 1734 554 1737 558
rect 1785 554 1788 558
rect 892 537 895 540
rect 818 532 823 537
rect 861 532 864 537
rect 810 529 818 532
rect 732 519 735 524
rect 810 524 813 529
rect 869 533 880 536
rect 892 534 900 537
rect 762 518 767 523
rect 634 506 635 510
rect 659 507 660 511
rect 706 506 707 510
rect 523 499 587 503
rect 591 499 646 503
rect 650 499 671 503
rect 675 499 702 503
rect 706 499 735 503
rect 771 496 774 524
rect 801 496 804 520
rect 852 496 855 528
rect 869 527 872 533
rect 892 528 895 534
rect 904 529 907 532
rect 915 532 918 546
rect 1575 544 1578 548
rect 1602 544 1603 548
rect 1647 544 1649 548
rect 915 529 921 532
rect 915 524 918 529
rect 1504 524 1507 527
rect 1515 527 1518 533
rect 1522 527 1525 533
rect 1515 524 1525 527
rect 867 518 872 523
rect 876 496 879 524
rect 906 496 909 520
rect 1515 519 1518 524
rect 1522 519 1525 524
rect 1531 529 1534 533
rect 1531 525 1533 529
rect 1537 525 1539 529
rect 1547 528 1550 533
rect 1575 530 1578 533
rect 1547 526 1558 528
rect 1531 519 1534 525
rect 1547 524 1553 526
rect 1547 519 1550 524
rect 1557 524 1558 526
rect 1576 526 1578 530
rect 1575 519 1578 526
rect 1720 537 1723 540
rect 1591 529 1594 533
rect 1601 529 1604 533
rect 1601 525 1610 529
rect 1622 528 1625 533
rect 1647 529 1650 533
rect 1591 519 1594 525
rect 1601 519 1604 525
rect 1622 524 1623 528
rect 1627 524 1630 527
rect 1649 525 1650 529
rect 1665 528 1668 533
rect 1697 533 1708 536
rect 1720 534 1728 537
rect 1622 519 1625 524
rect 1647 519 1650 525
rect 1697 527 1700 533
rect 1720 528 1723 534
rect 1732 529 1735 532
rect 1743 532 1746 546
rect 1794 541 1797 546
rect 1809 548 1812 558
rect 1839 554 1842 558
rect 1778 537 1779 540
rect 1783 537 1786 540
rect 1825 537 1828 540
rect 1751 532 1756 537
rect 1794 532 1797 537
rect 1743 529 1751 532
rect 1665 519 1668 524
rect 1743 524 1746 529
rect 1802 533 1813 536
rect 1825 534 1833 537
rect 1695 518 1700 523
rect 1567 506 1568 510
rect 1592 507 1593 511
rect 1639 506 1640 510
rect 1456 499 1520 503
rect 1524 499 1579 503
rect 1583 499 1604 503
rect 1608 499 1635 503
rect 1639 499 1668 503
rect 1704 496 1707 524
rect 1734 496 1737 520
rect 1785 496 1788 528
rect 1802 527 1805 533
rect 1825 528 1828 534
rect 1837 529 1840 532
rect 1848 532 1851 546
rect 1848 529 1854 532
rect 1848 524 1851 529
rect 1800 518 1805 523
rect 1809 496 1812 524
rect 1839 496 1842 520
rect 511 492 573 496
rect 577 492 579 496
rect 583 492 587 496
rect 591 492 605 496
rect 609 492 614 496
rect 618 492 623 496
rect 627 492 646 496
rect 650 492 680 496
rect 684 492 695 496
rect 699 492 723 496
rect 727 492 740 496
rect 744 492 764 496
rect 768 492 818 496
rect 822 492 845 496
rect 849 492 869 496
rect 873 492 921 496
rect 1444 492 1506 496
rect 1510 492 1512 496
rect 1516 492 1520 496
rect 1524 492 1538 496
rect 1542 492 1547 496
rect 1551 492 1556 496
rect 1560 492 1579 496
rect 1583 492 1613 496
rect 1617 492 1628 496
rect 1632 492 1656 496
rect 1660 492 1673 496
rect 1677 492 1697 496
rect 1701 492 1751 496
rect 1755 492 1778 496
rect 1782 492 1802 496
rect 1806 492 1854 496
rect 523 485 587 489
rect 591 485 646 489
rect 650 485 671 489
rect 675 485 702 489
rect 706 485 735 489
rect 634 478 635 482
rect 659 477 660 481
rect 706 478 707 482
rect 771 473 774 492
rect 876 473 879 492
rect 1456 485 1520 489
rect 1524 485 1579 489
rect 1583 485 1604 489
rect 1608 485 1635 489
rect 1639 485 1668 489
rect 1567 478 1568 482
rect 1592 477 1593 481
rect 1639 478 1640 482
rect 1704 473 1707 492
rect 1809 473 1812 492
rect 582 464 585 469
rect 589 464 592 469
rect 572 461 574 464
rect 582 461 592 464
rect 582 455 585 461
rect 589 455 592 461
rect 598 463 601 469
rect 614 464 617 469
rect 598 459 600 463
rect 604 459 606 463
rect 614 462 620 464
rect 624 462 625 464
rect 614 460 625 462
rect 642 462 645 469
rect 598 455 601 459
rect 614 455 617 460
rect 643 458 645 462
rect 642 455 645 458
rect 658 463 661 469
rect 668 463 671 469
rect 689 464 692 469
rect 668 459 677 463
rect 689 460 690 464
rect 694 461 697 464
rect 714 463 717 469
rect 732 464 735 469
rect 658 455 661 459
rect 668 455 671 459
rect 689 455 692 460
rect 716 459 717 463
rect 761 460 766 465
rect 770 461 772 464
rect 787 463 790 469
rect 787 460 795 463
rect 867 460 872 465
rect 876 461 877 464
rect 892 463 895 469
rect 892 460 900 463
rect 1515 464 1518 469
rect 1522 464 1525 469
rect 1505 461 1507 464
rect 1515 461 1525 464
rect 714 455 717 459
rect 732 455 735 460
rect 787 457 790 460
rect 892 457 895 460
rect 1515 455 1518 461
rect 642 440 645 444
rect 669 440 670 444
rect 714 440 716 444
rect 535 433 599 437
rect 603 433 630 437
rect 634 433 652 437
rect 656 433 717 437
rect 721 433 735 437
rect 771 430 774 449
rect 876 430 879 449
rect 1522 455 1525 461
rect 1531 463 1534 469
rect 1547 464 1550 469
rect 1531 459 1533 463
rect 1537 459 1539 463
rect 1547 462 1553 464
rect 1557 462 1558 464
rect 1547 460 1558 462
rect 1575 462 1578 469
rect 1531 455 1534 459
rect 1547 455 1550 460
rect 1576 458 1578 462
rect 1575 455 1578 458
rect 1591 463 1594 469
rect 1601 463 1604 469
rect 1622 464 1625 469
rect 1601 459 1610 463
rect 1622 460 1623 464
rect 1627 461 1630 464
rect 1647 463 1650 469
rect 1665 464 1668 469
rect 1591 455 1594 459
rect 1601 455 1604 459
rect 1622 455 1625 460
rect 1649 459 1650 463
rect 1694 460 1699 465
rect 1703 461 1705 464
rect 1720 463 1723 469
rect 1720 460 1728 463
rect 1800 460 1805 465
rect 1809 461 1810 464
rect 1825 463 1828 469
rect 1825 460 1833 463
rect 1647 455 1650 459
rect 1665 455 1668 460
rect 1720 457 1723 460
rect 1825 457 1828 460
rect 1575 440 1578 444
rect 1602 440 1603 444
rect 1647 440 1649 444
rect 1468 433 1532 437
rect 1536 433 1563 437
rect 1567 433 1585 437
rect 1589 433 1650 437
rect 1654 433 1668 437
rect 1704 430 1707 449
rect 1809 430 1812 449
rect 499 426 572 430
rect 576 426 588 430
rect 592 426 606 430
rect 610 426 617 430
rect 621 426 623 430
rect 627 426 642 430
rect 646 426 679 430
rect 683 426 684 430
rect 688 426 696 430
rect 700 426 724 430
rect 728 426 740 430
rect 744 426 764 430
rect 768 426 818 430
rect 822 426 845 430
rect 849 426 899 430
rect 903 426 907 430
rect 911 426 935 430
rect 939 426 989 430
rect 1432 426 1505 430
rect 1509 426 1521 430
rect 1525 426 1539 430
rect 1543 426 1550 430
rect 1554 426 1556 430
rect 1560 426 1575 430
rect 1579 426 1612 430
rect 1616 426 1617 430
rect 1621 426 1629 430
rect 1633 426 1657 430
rect 1661 426 1673 430
rect 1677 426 1697 430
rect 1701 426 1751 430
rect 1755 426 1778 430
rect 1782 426 1832 430
rect 1836 426 1840 430
rect 1844 426 1868 430
rect 1872 426 1922 430
rect 535 419 599 423
rect 603 419 630 423
rect 634 419 652 423
rect 656 419 717 423
rect 721 419 735 423
rect 771 416 774 426
rect 801 422 804 426
rect 828 422 831 426
rect 642 412 645 416
rect 669 412 670 416
rect 714 412 716 416
rect 571 392 574 395
rect 582 395 585 401
rect 589 395 592 401
rect 582 392 592 395
rect 582 387 585 392
rect 589 387 592 392
rect 598 397 601 401
rect 598 393 600 397
rect 604 393 606 397
rect 614 396 617 401
rect 642 398 645 401
rect 614 394 625 396
rect 598 387 601 393
rect 614 392 620 394
rect 614 387 617 392
rect 624 392 625 394
rect 643 394 645 398
rect 642 387 645 394
rect 787 405 790 408
rect 658 397 661 401
rect 668 397 671 401
rect 668 393 677 397
rect 689 396 692 401
rect 714 397 717 401
rect 658 387 661 393
rect 668 387 671 393
rect 689 392 690 396
rect 694 392 697 395
rect 716 393 717 397
rect 732 396 735 401
rect 764 401 775 404
rect 787 402 795 405
rect 689 387 692 392
rect 714 387 717 393
rect 764 395 767 401
rect 787 396 790 402
rect 799 397 802 400
rect 810 400 813 414
rect 837 409 840 414
rect 852 416 855 426
rect 882 422 885 426
rect 918 422 921 426
rect 821 405 822 408
rect 826 405 829 408
rect 868 405 871 408
rect 810 397 818 400
rect 837 400 840 405
rect 732 387 735 392
rect 810 392 813 397
rect 818 393 822 397
rect 845 401 856 404
rect 868 402 876 405
rect 762 386 767 391
rect 634 374 635 378
rect 659 375 660 379
rect 706 374 707 378
rect 523 367 587 371
rect 591 367 646 371
rect 650 367 671 371
rect 675 367 702 371
rect 706 367 735 371
rect 771 364 774 392
rect 801 364 804 388
rect 828 364 831 396
rect 845 395 848 401
rect 868 396 871 402
rect 880 397 883 400
rect 891 400 894 414
rect 927 409 930 414
rect 942 416 945 426
rect 972 422 975 426
rect 916 405 919 408
rect 1468 419 1532 423
rect 1536 419 1563 423
rect 1567 419 1585 423
rect 1589 419 1650 423
rect 1654 419 1668 423
rect 1704 416 1707 426
rect 1734 422 1737 426
rect 1761 422 1764 426
rect 958 405 961 408
rect 891 397 900 400
rect 927 400 930 405
rect 891 392 894 397
rect 843 386 848 391
rect 852 364 855 392
rect 934 403 946 404
rect 938 401 946 403
rect 958 402 966 405
rect 958 396 961 402
rect 970 397 973 400
rect 981 400 984 414
rect 1575 412 1578 416
rect 1602 412 1603 416
rect 1647 412 1649 416
rect 981 397 1001 400
rect 882 364 885 388
rect 918 364 921 396
rect 981 392 984 397
rect 1504 392 1507 395
rect 1515 395 1518 401
rect 1522 395 1525 401
rect 1515 392 1525 395
rect 942 364 945 392
rect 972 364 975 388
rect 1515 387 1518 392
rect 1522 387 1525 392
rect 1531 397 1534 401
rect 1531 393 1533 397
rect 1537 393 1539 397
rect 1547 396 1550 401
rect 1575 398 1578 401
rect 1547 394 1558 396
rect 1531 387 1534 393
rect 1547 392 1553 394
rect 1547 387 1550 392
rect 1557 392 1558 394
rect 1576 394 1578 398
rect 1575 387 1578 394
rect 1720 405 1723 408
rect 1591 397 1594 401
rect 1601 397 1604 401
rect 1601 393 1610 397
rect 1622 396 1625 401
rect 1647 397 1650 401
rect 1591 387 1594 393
rect 1601 387 1604 393
rect 1622 392 1623 396
rect 1627 392 1630 395
rect 1649 393 1650 397
rect 1665 396 1668 401
rect 1697 401 1708 404
rect 1720 402 1728 405
rect 1622 387 1625 392
rect 1647 387 1650 393
rect 1697 395 1700 401
rect 1720 396 1723 402
rect 1732 397 1735 400
rect 1743 400 1746 414
rect 1770 409 1773 414
rect 1785 416 1788 426
rect 1815 422 1818 426
rect 1851 422 1854 426
rect 1754 405 1755 408
rect 1759 405 1762 408
rect 1801 405 1804 408
rect 1743 397 1751 400
rect 1770 400 1773 405
rect 1665 387 1668 392
rect 1743 392 1746 397
rect 1751 393 1755 397
rect 1778 401 1789 404
rect 1801 402 1809 405
rect 1695 386 1700 391
rect 1567 374 1568 378
rect 1592 375 1593 379
rect 1639 374 1640 378
rect 1456 367 1520 371
rect 1524 367 1579 371
rect 1583 367 1604 371
rect 1608 367 1635 371
rect 1639 367 1668 371
rect 1704 364 1707 392
rect 1734 364 1737 388
rect 1761 364 1764 396
rect 1778 395 1781 401
rect 1801 396 1804 402
rect 1813 397 1816 400
rect 1824 400 1827 414
rect 1860 409 1863 414
rect 1875 416 1878 426
rect 1905 422 1908 426
rect 1849 405 1852 408
rect 1891 405 1894 408
rect 1824 397 1833 400
rect 1860 400 1863 405
rect 1824 392 1827 397
rect 1776 386 1781 391
rect 1785 364 1788 392
rect 1867 403 1879 404
rect 1871 401 1879 403
rect 1891 402 1899 405
rect 1891 396 1894 402
rect 1903 397 1906 400
rect 1914 400 1917 414
rect 1914 397 1934 400
rect 1815 364 1818 388
rect 1851 364 1854 396
rect 1914 392 1917 397
rect 1875 364 1878 392
rect 1905 364 1908 388
rect 511 360 573 364
rect 577 360 579 364
rect 583 360 587 364
rect 591 360 605 364
rect 609 360 614 364
rect 618 360 623 364
rect 627 360 646 364
rect 650 360 680 364
rect 684 360 695 364
rect 699 360 723 364
rect 727 360 740 364
rect 744 360 764 364
rect 768 360 818 364
rect 825 360 845 364
rect 849 360 899 364
rect 903 360 935 364
rect 939 360 989 364
rect 1444 360 1506 364
rect 1510 360 1512 364
rect 1516 360 1520 364
rect 1524 360 1538 364
rect 1542 360 1547 364
rect 1551 360 1556 364
rect 1560 360 1579 364
rect 1583 360 1613 364
rect 1617 360 1628 364
rect 1632 360 1656 364
rect 1660 360 1673 364
rect 1677 360 1697 364
rect 1701 360 1751 364
rect 1758 360 1778 364
rect 1782 360 1832 364
rect 1836 360 1868 364
rect 1872 360 1922 364
rect 523 353 587 357
rect 591 353 646 357
rect 650 353 671 357
rect 675 353 702 357
rect 706 353 735 357
rect 634 346 635 350
rect 659 345 660 349
rect 706 346 707 350
rect 582 332 585 337
rect 589 332 592 337
rect 572 329 574 332
rect 582 329 592 332
rect 582 323 585 329
rect 589 323 592 329
rect 598 331 601 337
rect 614 332 617 337
rect 598 327 600 331
rect 604 327 606 331
rect 614 330 620 332
rect 624 330 625 332
rect 614 328 625 330
rect 642 330 645 337
rect 598 323 601 327
rect 614 323 617 328
rect 643 326 645 330
rect 642 323 645 326
rect 658 331 661 337
rect 668 331 671 337
rect 689 332 692 337
rect 668 327 677 331
rect 689 328 690 332
rect 694 329 697 332
rect 714 331 717 337
rect 732 332 735 337
rect 771 338 774 360
rect 852 338 855 360
rect 942 338 945 360
rect 1456 353 1520 357
rect 1524 353 1579 357
rect 1583 353 1604 357
rect 1608 353 1635 357
rect 1639 353 1668 357
rect 1567 346 1568 350
rect 1592 345 1593 349
rect 1639 346 1640 350
rect 658 323 661 327
rect 668 323 671 327
rect 689 323 692 328
rect 716 327 717 331
rect 714 323 717 327
rect 732 323 735 328
rect 762 325 767 330
rect 771 326 772 329
rect 787 328 790 334
rect 787 325 795 328
rect 842 325 847 330
rect 851 326 853 329
rect 868 328 871 334
rect 868 325 876 328
rect 935 326 943 329
rect 958 328 961 334
rect 1515 332 1518 337
rect 1522 332 1525 337
rect 1505 329 1507 332
rect 958 325 966 328
rect 1515 329 1525 332
rect 787 322 790 325
rect 868 322 871 325
rect 958 322 961 325
rect 1515 323 1518 329
rect 642 308 645 312
rect 669 308 670 312
rect 714 308 716 312
rect 1522 323 1525 329
rect 1531 331 1534 337
rect 1547 332 1550 337
rect 1531 327 1533 331
rect 1537 327 1539 331
rect 1547 330 1553 332
rect 1557 330 1558 332
rect 1547 328 1558 330
rect 1575 330 1578 337
rect 1531 323 1534 327
rect 1547 323 1550 328
rect 1576 326 1578 330
rect 1575 323 1578 326
rect 1591 331 1594 337
rect 1601 331 1604 337
rect 1622 332 1625 337
rect 1601 327 1610 331
rect 1622 328 1623 332
rect 1627 329 1630 332
rect 1647 331 1650 337
rect 1665 332 1668 337
rect 1704 338 1707 360
rect 1785 338 1788 360
rect 1875 338 1878 360
rect 1591 323 1594 327
rect 1601 323 1604 327
rect 1622 323 1625 328
rect 1649 327 1650 331
rect 1647 323 1650 327
rect 1665 323 1668 328
rect 1695 325 1700 330
rect 1704 326 1705 329
rect 1720 328 1723 334
rect 1720 325 1728 328
rect 1775 325 1780 330
rect 1784 326 1786 329
rect 1801 328 1804 334
rect 1801 325 1809 328
rect 1868 326 1876 329
rect 1891 328 1894 334
rect 1891 325 1899 328
rect 1720 322 1723 325
rect 1801 322 1804 325
rect 1891 322 1894 325
rect 535 301 599 305
rect 603 301 630 305
rect 634 301 652 305
rect 656 301 717 305
rect 721 301 735 305
rect 771 298 774 314
rect 852 298 855 314
rect 942 298 945 314
rect 1575 308 1578 312
rect 1602 308 1603 312
rect 1647 308 1649 312
rect 1468 301 1532 305
rect 1536 301 1563 305
rect 1567 301 1585 305
rect 1589 301 1650 305
rect 1654 301 1668 305
rect 1704 298 1707 314
rect 1785 298 1788 314
rect 1875 298 1878 314
rect 499 294 572 298
rect 576 294 588 298
rect 592 294 606 298
rect 610 294 617 298
rect 621 294 623 298
rect 627 294 642 298
rect 646 294 679 298
rect 683 294 684 298
rect 688 294 696 298
rect 700 294 724 298
rect 728 294 740 298
rect 744 294 764 298
rect 768 294 818 298
rect 822 294 845 298
rect 849 294 935 298
rect 939 294 993 298
rect 1432 294 1505 298
rect 1509 294 1521 298
rect 1525 294 1539 298
rect 1543 294 1550 298
rect 1554 294 1556 298
rect 1560 294 1575 298
rect 1579 294 1612 298
rect 1616 294 1617 298
rect 1621 294 1629 298
rect 1633 294 1657 298
rect 1661 294 1673 298
rect 1677 294 1697 298
rect 1701 294 1751 298
rect 1755 294 1778 298
rect 1782 294 1868 298
rect 1872 294 1926 298
rect 535 287 599 291
rect 603 287 630 291
rect 634 287 652 291
rect 656 287 717 291
rect 721 287 735 291
rect 771 284 774 294
rect 801 290 804 294
rect 642 280 645 284
rect 669 280 670 284
rect 714 280 716 284
rect 571 260 574 263
rect 582 263 585 269
rect 589 263 592 269
rect 582 260 592 263
rect 582 255 585 260
rect 589 255 592 260
rect 598 265 601 269
rect 598 261 600 265
rect 604 261 606 265
rect 614 264 617 269
rect 642 266 645 269
rect 614 262 625 264
rect 598 255 601 261
rect 614 260 620 262
rect 614 255 617 260
rect 624 260 625 262
rect 643 262 645 266
rect 642 255 645 262
rect 1468 287 1532 291
rect 1536 287 1563 291
rect 1567 287 1585 291
rect 1589 287 1650 291
rect 1654 287 1668 291
rect 1704 284 1707 294
rect 1734 290 1737 294
rect 787 273 790 276
rect 658 265 661 269
rect 668 265 671 269
rect 668 261 677 265
rect 689 264 692 269
rect 714 265 717 269
rect 658 255 661 261
rect 668 255 671 261
rect 689 260 690 264
rect 694 260 697 263
rect 716 261 717 265
rect 732 264 735 269
rect 764 269 775 272
rect 787 270 795 273
rect 689 255 692 260
rect 714 255 717 261
rect 764 263 767 269
rect 787 264 790 270
rect 799 265 802 268
rect 810 268 813 282
rect 1575 280 1578 284
rect 1602 280 1603 284
rect 1647 280 1649 284
rect 818 268 823 273
rect 810 265 818 268
rect 732 255 735 260
rect 810 260 813 265
rect 1504 260 1507 263
rect 1515 263 1518 269
rect 1522 263 1525 269
rect 1515 260 1525 263
rect 762 254 767 259
rect 93 239 102 243
rect 106 239 138 243
rect 142 239 205 243
rect 209 239 234 243
rect 238 239 270 243
rect 274 239 337 243
rect 341 239 366 243
rect 370 239 402 243
rect 406 239 469 243
rect 473 239 553 243
rect 634 242 635 246
rect 659 243 660 247
rect 706 242 707 246
rect 93 232 126 236
rect 130 232 154 236
rect 158 232 184 236
rect 188 232 221 236
rect 225 232 258 236
rect 262 232 286 236
rect 290 232 316 236
rect 320 232 353 236
rect 357 232 390 236
rect 394 232 418 236
rect 422 232 448 236
rect 452 232 485 236
rect 489 232 493 236
rect 566 235 587 239
rect 591 235 596 239
rect 600 235 646 239
rect 650 235 671 239
rect 675 235 702 239
rect 706 235 735 239
rect 771 232 774 260
rect 801 232 804 256
rect 1515 255 1518 260
rect 1522 255 1525 260
rect 1531 265 1534 269
rect 1531 261 1533 265
rect 1537 261 1539 265
rect 1547 264 1550 269
rect 1575 266 1578 269
rect 1547 262 1558 264
rect 1531 255 1534 261
rect 1547 260 1553 262
rect 1547 255 1550 260
rect 1557 260 1558 262
rect 1576 262 1578 266
rect 1575 255 1578 262
rect 1720 273 1723 276
rect 1591 265 1594 269
rect 1601 265 1604 269
rect 1601 261 1610 265
rect 1622 264 1625 269
rect 1647 265 1650 269
rect 1591 255 1594 261
rect 1601 255 1604 261
rect 1622 260 1623 264
rect 1627 260 1630 263
rect 1649 261 1650 265
rect 1665 264 1668 269
rect 1697 269 1708 272
rect 1720 270 1728 273
rect 1622 255 1625 260
rect 1647 255 1650 261
rect 1697 263 1700 269
rect 1720 264 1723 270
rect 1732 265 1735 268
rect 1743 268 1746 282
rect 1751 268 1756 273
rect 1743 265 1751 268
rect 1665 255 1668 260
rect 1743 260 1746 265
rect 1695 254 1700 259
rect 1026 239 1035 243
rect 1039 239 1071 243
rect 1075 239 1138 243
rect 1142 239 1167 243
rect 1171 239 1203 243
rect 1207 239 1270 243
rect 1274 239 1299 243
rect 1303 239 1335 243
rect 1339 239 1402 243
rect 1406 239 1486 243
rect 1567 242 1568 246
rect 1592 243 1593 247
rect 1639 242 1640 246
rect 1026 232 1059 236
rect 1063 232 1087 236
rect 1091 232 1117 236
rect 1121 232 1154 236
rect 1158 232 1191 236
rect 1195 232 1219 236
rect 1223 232 1249 236
rect 1253 232 1286 236
rect 1290 232 1323 236
rect 1327 232 1351 236
rect 1355 232 1381 236
rect 1385 232 1418 236
rect 1422 232 1426 236
rect 1499 235 1520 239
rect 1524 235 1529 239
rect 1533 235 1579 239
rect 1583 235 1604 239
rect 1608 235 1635 239
rect 1639 235 1668 239
rect 1704 232 1707 260
rect 1734 232 1737 256
rect 96 222 99 232
rect 117 222 120 232
rect 133 222 136 232
rect 147 225 152 229
rect 156 225 163 229
rect 175 222 178 232
rect 191 222 194 232
rect 212 222 215 232
rect 228 222 231 232
rect 249 222 252 232
rect 265 222 268 232
rect 279 225 284 229
rect 288 225 295 229
rect 307 222 310 232
rect 323 222 326 232
rect 344 222 347 232
rect 360 222 363 232
rect 381 222 384 232
rect 397 222 400 232
rect 411 225 416 229
rect 420 225 427 229
rect 439 222 442 232
rect 455 222 458 232
rect 476 222 479 232
rect 511 228 573 232
rect 577 228 579 232
rect 583 228 587 232
rect 591 228 605 232
rect 609 228 614 232
rect 618 228 623 232
rect 627 228 646 232
rect 650 228 680 232
rect 684 228 695 232
rect 699 228 723 232
rect 727 228 740 232
rect 744 228 764 232
rect 768 228 848 232
rect 852 228 866 232
rect 870 228 875 232
rect 879 228 884 232
rect 888 228 907 232
rect 911 228 941 232
rect 945 228 956 232
rect 960 228 984 232
rect 988 228 997 232
rect 113 208 118 211
rect 122 208 146 211
rect 171 208 178 211
rect 182 208 204 211
rect 224 208 231 211
rect 245 208 250 211
rect 254 208 278 211
rect 303 208 310 211
rect 314 208 336 211
rect 356 208 363 211
rect 377 208 382 211
rect 386 208 410 211
rect 523 221 587 225
rect 591 221 596 225
rect 600 221 646 225
rect 650 221 671 225
rect 675 221 702 225
rect 706 221 735 225
rect 435 208 442 211
rect 446 208 468 211
rect 634 214 635 218
rect 659 213 660 217
rect 706 214 707 218
rect 129 198 136 201
rect 140 202 159 205
rect 159 195 162 201
rect 187 198 194 201
rect 198 202 213 205
rect 261 198 268 201
rect 272 202 291 205
rect 291 195 294 201
rect 319 198 326 201
rect 330 202 345 205
rect 393 198 400 201
rect 404 202 423 205
rect 423 195 426 201
rect 451 198 458 201
rect 462 202 479 205
rect 582 200 585 205
rect 589 200 592 205
rect 572 197 574 200
rect 582 197 592 200
rect 582 191 585 197
rect 96 179 99 191
rect 117 179 120 191
rect 133 179 136 191
rect 147 182 159 185
rect 175 179 178 191
rect 191 179 194 191
rect 212 179 215 191
rect 228 179 231 191
rect 249 179 252 191
rect 265 179 268 191
rect 279 182 291 185
rect 307 179 310 191
rect 323 179 326 191
rect 344 179 347 191
rect 360 179 363 191
rect 381 179 384 191
rect 397 179 400 191
rect 411 182 423 185
rect 439 179 442 191
rect 455 179 458 191
rect 476 179 479 191
rect 589 191 592 197
rect 598 199 601 205
rect 614 200 617 205
rect 598 195 600 199
rect 604 195 606 199
rect 614 198 620 200
rect 624 198 625 200
rect 614 196 625 198
rect 642 198 645 205
rect 598 191 601 195
rect 614 191 617 196
rect 643 194 645 198
rect 642 191 645 194
rect 658 199 661 205
rect 668 199 671 205
rect 689 200 692 205
rect 668 195 677 199
rect 689 196 690 200
rect 694 197 697 200
rect 714 199 717 205
rect 732 200 735 205
rect 771 202 774 228
rect 807 221 826 225
rect 830 221 848 225
rect 852 221 907 225
rect 911 221 932 225
rect 936 221 963 225
rect 967 221 996 225
rect 1029 222 1032 232
rect 1050 222 1053 232
rect 1066 222 1069 232
rect 1080 225 1085 229
rect 1089 225 1096 229
rect 1108 222 1111 232
rect 1124 222 1127 232
rect 1145 222 1148 232
rect 1161 222 1164 232
rect 1182 222 1185 232
rect 1198 222 1201 232
rect 1212 225 1217 229
rect 1221 225 1228 229
rect 1240 222 1243 232
rect 1256 222 1259 232
rect 1277 222 1280 232
rect 1293 222 1296 232
rect 1314 222 1317 232
rect 1330 222 1333 232
rect 1344 225 1349 229
rect 1353 225 1360 229
rect 1372 222 1375 232
rect 1388 222 1391 232
rect 1409 222 1412 232
rect 1444 228 1506 232
rect 1510 228 1512 232
rect 1516 228 1520 232
rect 1524 228 1538 232
rect 1542 228 1547 232
rect 1551 228 1556 232
rect 1560 228 1579 232
rect 1583 228 1613 232
rect 1617 228 1628 232
rect 1632 228 1656 232
rect 1660 228 1673 232
rect 1677 228 1697 232
rect 1701 228 1781 232
rect 1785 228 1799 232
rect 1803 228 1808 232
rect 1812 228 1817 232
rect 1821 228 1840 232
rect 1844 228 1874 232
rect 1878 228 1889 232
rect 1893 228 1917 232
rect 1921 228 1930 232
rect 807 209 810 221
rect 895 214 896 218
rect 920 213 921 217
rect 967 214 968 218
rect 658 191 661 195
rect 668 191 671 195
rect 689 191 692 196
rect 716 195 717 199
rect 834 200 837 205
rect 843 200 846 205
rect 850 200 853 205
rect 714 191 717 195
rect 732 191 735 196
rect 761 189 766 194
rect 770 190 772 193
rect 787 192 790 198
rect 819 197 853 200
rect 787 189 795 192
rect 787 186 790 189
rect 93 175 126 179
rect 130 175 154 179
rect 158 175 184 179
rect 188 175 258 179
rect 262 175 286 179
rect 290 175 316 179
rect 320 175 390 179
rect 394 175 418 179
rect 422 175 448 179
rect 452 175 505 179
rect 642 176 645 180
rect 669 176 670 180
rect 714 176 716 180
rect 819 183 822 197
rect 843 191 846 197
rect 850 191 853 197
rect 859 199 862 205
rect 875 200 878 205
rect 859 195 861 199
rect 865 195 867 199
rect 875 198 881 200
rect 885 198 886 200
rect 875 196 886 198
rect 903 198 906 205
rect 859 191 862 195
rect 875 191 878 196
rect 904 194 906 198
rect 903 191 906 194
rect 1046 208 1051 211
rect 1055 208 1079 211
rect 1104 208 1111 211
rect 1115 208 1137 211
rect 1157 208 1164 211
rect 1178 208 1183 211
rect 1187 208 1211 211
rect 1236 208 1243 211
rect 1247 208 1269 211
rect 1289 208 1296 211
rect 1310 208 1315 211
rect 1319 208 1343 211
rect 1456 221 1520 225
rect 1524 221 1529 225
rect 1533 221 1579 225
rect 1583 221 1604 225
rect 1608 221 1635 225
rect 1639 221 1668 225
rect 1368 208 1375 211
rect 1379 208 1401 211
rect 1567 214 1568 218
rect 1592 213 1593 217
rect 1639 214 1640 218
rect 919 199 922 205
rect 929 199 932 205
rect 950 200 953 205
rect 929 195 938 199
rect 950 196 951 200
rect 955 197 958 200
rect 975 199 978 205
rect 993 200 996 205
rect 919 191 922 195
rect 929 191 932 195
rect 950 191 953 196
rect 977 195 978 199
rect 975 191 978 195
rect 993 191 996 196
rect 1062 198 1069 201
rect 1073 202 1092 205
rect 1092 195 1095 201
rect 1120 198 1127 201
rect 1131 202 1146 205
rect 1194 198 1201 201
rect 1205 202 1224 205
rect 1224 195 1227 201
rect 1252 198 1259 201
rect 1263 202 1278 205
rect 1326 198 1333 201
rect 1337 202 1356 205
rect 1356 195 1359 201
rect 1384 198 1391 201
rect 1395 202 1412 205
rect 1515 200 1518 205
rect 1522 200 1525 205
rect 1505 197 1507 200
rect 1515 197 1525 200
rect 1515 191 1518 197
rect 93 168 102 172
rect 106 168 153 172
rect 157 168 203 172
rect 207 168 234 172
rect 238 168 285 172
rect 289 168 335 172
rect 339 168 366 172
rect 370 168 417 172
rect 421 168 467 172
rect 471 169 541 172
rect 585 169 599 173
rect 603 169 630 173
rect 634 169 652 173
rect 656 169 717 173
rect 721 169 735 173
rect 771 166 774 178
rect 903 176 906 180
rect 930 176 931 180
rect 975 176 977 180
rect 1029 179 1032 191
rect 1050 179 1053 191
rect 1066 179 1069 191
rect 1080 182 1092 185
rect 1108 179 1111 191
rect 1124 179 1127 191
rect 1145 179 1148 191
rect 1161 179 1164 191
rect 1182 179 1185 191
rect 1198 179 1201 191
rect 1212 182 1224 185
rect 1240 179 1243 191
rect 1256 179 1259 191
rect 1277 179 1280 191
rect 1293 179 1296 191
rect 1314 179 1317 191
rect 1330 179 1333 191
rect 1344 182 1356 185
rect 1372 179 1375 191
rect 1388 179 1391 191
rect 1409 179 1412 191
rect 1522 191 1525 197
rect 1531 199 1534 205
rect 1547 200 1550 205
rect 1531 195 1533 199
rect 1537 195 1539 199
rect 1547 198 1553 200
rect 1557 198 1558 200
rect 1547 196 1558 198
rect 1575 198 1578 205
rect 1531 191 1534 195
rect 1547 191 1550 196
rect 1576 194 1578 198
rect 1575 191 1578 194
rect 1591 199 1594 205
rect 1601 199 1604 205
rect 1622 200 1625 205
rect 1601 195 1610 199
rect 1622 196 1623 200
rect 1627 197 1630 200
rect 1647 199 1650 205
rect 1665 200 1668 205
rect 1704 202 1707 228
rect 1740 221 1759 225
rect 1763 221 1781 225
rect 1785 221 1840 225
rect 1844 221 1865 225
rect 1869 221 1896 225
rect 1900 221 1929 225
rect 1740 209 1743 221
rect 1828 214 1829 218
rect 1853 213 1854 217
rect 1900 214 1901 218
rect 1591 191 1594 195
rect 1601 191 1604 195
rect 1622 191 1625 196
rect 1649 195 1650 199
rect 1767 200 1770 205
rect 1776 200 1779 205
rect 1783 200 1786 205
rect 1647 191 1650 195
rect 1665 191 1668 196
rect 1694 189 1699 194
rect 1703 190 1705 193
rect 1720 192 1723 198
rect 1752 197 1786 200
rect 1720 189 1728 192
rect 1720 186 1723 189
rect 1026 175 1059 179
rect 1063 175 1087 179
rect 1091 175 1117 179
rect 1121 175 1191 179
rect 1195 175 1219 179
rect 1223 175 1249 179
rect 1253 175 1323 179
rect 1327 175 1351 179
rect 1355 175 1381 179
rect 1385 175 1438 179
rect 1575 176 1578 180
rect 1602 176 1603 180
rect 1647 176 1649 180
rect 1752 183 1755 197
rect 1776 191 1779 197
rect 1783 191 1786 197
rect 1792 199 1795 205
rect 1808 200 1811 205
rect 1792 195 1794 199
rect 1798 195 1800 199
rect 1808 198 1814 200
rect 1818 198 1819 200
rect 1808 196 1819 198
rect 1836 198 1839 205
rect 1792 191 1795 195
rect 1808 191 1811 196
rect 1837 194 1839 198
rect 1836 191 1839 194
rect 1852 199 1855 205
rect 1862 199 1865 205
rect 1883 200 1886 205
rect 1862 195 1871 199
rect 1883 196 1884 200
rect 1888 197 1891 200
rect 1908 199 1911 205
rect 1926 200 1929 205
rect 1852 191 1855 195
rect 1862 191 1865 195
rect 1883 191 1886 196
rect 1910 195 1911 199
rect 1908 191 1911 195
rect 1926 191 1929 196
rect 811 169 816 173
rect 820 169 860 173
rect 864 169 891 173
rect 895 169 913 173
rect 917 169 978 173
rect 982 169 996 173
rect 1026 168 1035 172
rect 1039 168 1086 172
rect 1090 168 1136 172
rect 1140 168 1167 172
rect 1171 168 1218 172
rect 1222 168 1268 172
rect 1272 168 1299 172
rect 1303 168 1350 172
rect 1354 168 1400 172
rect 1404 169 1474 172
rect 1518 169 1532 173
rect 1536 169 1563 173
rect 1567 169 1585 173
rect 1589 169 1650 173
rect 1654 169 1668 173
rect 1704 166 1707 178
rect 1836 176 1839 180
rect 1863 176 1864 180
rect 1908 176 1910 180
rect 1744 169 1749 173
rect 1753 169 1793 173
rect 1797 169 1824 173
rect 1828 169 1846 173
rect 1850 169 1911 173
rect 1915 169 1929 173
rect 100 162 484 165
rect 499 162 572 166
rect 576 162 588 166
rect 592 162 606 166
rect 610 162 617 166
rect 621 162 623 166
rect 627 162 642 166
rect 646 162 679 166
rect 683 162 684 166
rect 688 162 696 166
rect 700 162 724 166
rect 728 162 764 166
rect 768 162 807 166
rect 811 162 818 166
rect 822 162 833 166
rect 837 162 849 166
rect 853 162 867 166
rect 871 162 878 166
rect 882 162 884 166
rect 888 162 903 166
rect 907 162 940 166
rect 944 162 945 166
rect 949 162 957 166
rect 961 162 985 166
rect 989 162 997 166
rect 1033 162 1417 165
rect 1432 162 1505 166
rect 1509 162 1521 166
rect 1525 162 1539 166
rect 1543 162 1550 166
rect 1554 162 1556 166
rect 1560 162 1575 166
rect 1579 162 1612 166
rect 1616 162 1617 166
rect 1621 162 1629 166
rect 1633 162 1657 166
rect 1661 162 1697 166
rect 1701 162 1740 166
rect 1744 162 1751 166
rect 1755 162 1766 166
rect 1770 162 1782 166
rect 1786 162 1800 166
rect 1804 162 1811 166
rect 1815 162 1817 166
rect 1821 162 1836 166
rect 1840 162 1873 166
rect 1877 162 1878 166
rect 1882 162 1890 166
rect 1894 162 1918 166
rect 1922 162 1930 166
rect 243 155 352 158
rect 535 155 581 159
rect 585 155 815 158
rect 1005 156 1013 160
rect 1176 155 1285 158
rect 1468 155 1514 159
rect 1518 155 1748 158
rect 1938 156 1946 160
rect 223 147 227 151
rect 231 147 235 151
rect 523 148 825 151
rect 1001 140 1005 144
rect 1156 147 1160 151
rect 1164 147 1168 151
rect 1456 148 1758 151
rect 1934 140 1938 144
rect 79 136 211 140
rect 215 136 231 140
rect 247 136 1144 140
rect 1148 136 1164 140
rect 1180 136 2026 140
rect 239 129 484 132
rect 559 129 873 133
rect 877 129 909 133
rect 913 129 976 133
rect 980 129 996 133
rect 1172 129 1417 132
rect 1492 129 1806 133
rect 1810 129 1842 133
rect 1846 129 1909 133
rect 1913 129 1929 133
rect 254 122 484 125
rect 499 122 859 126
rect 863 122 897 126
rect 901 122 925 126
rect 929 122 955 126
rect 959 122 992 126
rect 223 113 227 117
rect 231 113 235 117
rect 867 112 870 122
rect 888 112 891 122
rect 904 112 907 122
rect 918 115 923 119
rect 927 115 934 119
rect 946 112 949 122
rect 962 112 965 122
rect 983 112 986 122
rect 1187 122 1417 125
rect 1432 122 1792 126
rect 1796 122 1830 126
rect 1834 122 1858 126
rect 1862 122 1888 126
rect 1892 122 1925 126
rect 1156 113 1160 117
rect 1164 113 1168 117
rect 1800 112 1803 122
rect 1821 112 1824 122
rect 1837 112 1840 122
rect 1851 115 1856 119
rect 1860 115 1867 119
rect 1879 112 1882 122
rect 1895 112 1898 122
rect 1916 112 1919 122
rect 243 106 353 109
rect 93 99 102 103
rect 106 99 138 103
rect 142 99 205 103
rect 209 99 234 103
rect 238 99 270 103
rect 274 99 337 103
rect 341 99 366 103
rect 370 99 402 103
rect 406 99 469 103
rect 473 99 553 103
rect 93 92 126 96
rect 130 92 154 96
rect 158 92 184 96
rect 188 92 221 96
rect 225 92 258 96
rect 262 92 286 96
rect 290 92 316 96
rect 320 92 353 96
rect 357 92 390 96
rect 394 92 418 96
rect 422 92 448 96
rect 452 92 485 96
rect 489 92 493 96
rect 884 98 889 101
rect 893 98 917 101
rect 1176 106 1286 109
rect 942 98 949 101
rect 953 98 975 101
rect 1026 99 1035 103
rect 1039 99 1071 103
rect 1075 99 1138 103
rect 1142 99 1167 103
rect 1171 99 1203 103
rect 1207 99 1270 103
rect 1274 99 1299 103
rect 1303 99 1335 103
rect 1339 99 1402 103
rect 1406 99 1486 103
rect 96 82 99 92
rect 117 82 120 92
rect 133 82 136 92
rect 147 85 152 89
rect 156 85 163 89
rect 175 82 178 92
rect 191 82 194 92
rect 212 82 215 92
rect 228 82 231 92
rect 249 82 252 92
rect 265 82 268 92
rect 279 85 284 89
rect 288 85 295 89
rect 307 82 310 92
rect 323 82 326 92
rect 344 82 347 92
rect 360 82 363 92
rect 381 82 384 92
rect 397 82 400 92
rect 411 85 416 89
rect 420 85 427 89
rect 439 82 442 92
rect 455 82 458 92
rect 476 82 479 92
rect 900 88 907 91
rect 911 92 930 95
rect 113 68 118 71
rect 122 68 146 71
rect 171 68 178 71
rect 182 68 204 71
rect 224 68 231 71
rect 245 68 250 71
rect 254 68 278 71
rect 303 68 310 71
rect 314 68 336 71
rect 356 68 363 71
rect 377 68 382 71
rect 386 68 410 71
rect 435 68 442 71
rect 446 68 468 71
rect 930 85 933 91
rect 958 88 965 91
rect 969 92 984 95
rect 1026 92 1059 96
rect 1063 92 1087 96
rect 1091 92 1117 96
rect 1121 92 1154 96
rect 1158 92 1191 96
rect 1195 92 1219 96
rect 1223 92 1249 96
rect 1253 92 1286 96
rect 1290 92 1323 96
rect 1327 92 1351 96
rect 1355 92 1381 96
rect 1385 92 1418 96
rect 1422 92 1426 96
rect 1817 98 1822 101
rect 1826 98 1850 101
rect 1875 98 1882 101
rect 1886 98 1908 101
rect 1029 82 1032 92
rect 1050 82 1053 92
rect 1066 82 1069 92
rect 1080 85 1085 89
rect 1089 85 1096 89
rect 1108 82 1111 92
rect 1124 82 1127 92
rect 1145 82 1148 92
rect 1161 82 1164 92
rect 1182 82 1185 92
rect 1198 82 1201 92
rect 1212 85 1217 89
rect 1221 85 1228 89
rect 1240 82 1243 92
rect 1256 82 1259 92
rect 1277 82 1280 92
rect 1293 82 1296 92
rect 1314 82 1317 92
rect 1330 82 1333 92
rect 1344 85 1349 89
rect 1353 85 1360 89
rect 1372 82 1375 92
rect 1388 82 1391 92
rect 1409 82 1412 92
rect 1833 88 1840 91
rect 1844 92 1863 95
rect 867 69 870 81
rect 888 69 891 81
rect 904 69 907 81
rect 918 72 930 75
rect 946 69 949 81
rect 962 69 965 81
rect 983 69 986 81
rect 129 58 136 61
rect 140 62 159 65
rect 159 55 162 61
rect 187 58 194 61
rect 198 62 213 65
rect 261 58 268 61
rect 272 62 291 65
rect 291 55 294 61
rect 319 58 326 61
rect 330 62 345 65
rect 393 58 400 61
rect 404 62 423 65
rect 423 55 426 61
rect 451 58 458 61
rect 462 62 479 65
rect 511 65 897 69
rect 901 65 925 69
rect 929 65 955 69
rect 959 65 996 69
rect 1046 68 1051 71
rect 1055 68 1079 71
rect 1104 68 1111 71
rect 1115 68 1137 71
rect 1157 68 1164 71
rect 1178 68 1183 71
rect 1187 68 1211 71
rect 1236 68 1243 71
rect 1247 68 1269 71
rect 1289 68 1296 71
rect 1310 68 1315 71
rect 1319 68 1343 71
rect 1368 68 1375 71
rect 1379 68 1401 71
rect 1863 85 1866 91
rect 1891 88 1898 91
rect 1902 92 1917 95
rect 1800 69 1803 81
rect 1821 69 1824 81
rect 1837 69 1840 81
rect 1851 72 1863 75
rect 1879 69 1882 81
rect 1895 69 1898 81
rect 1916 69 1919 81
rect 547 58 873 62
rect 877 58 924 62
rect 928 58 974 62
rect 978 58 996 62
rect 1062 58 1069 61
rect 1073 62 1092 65
rect 96 39 99 51
rect 117 39 120 51
rect 133 39 136 51
rect 147 42 159 45
rect 175 39 178 51
rect 191 39 194 51
rect 212 39 215 51
rect 228 39 231 51
rect 249 39 252 51
rect 265 39 268 51
rect 279 42 291 45
rect 307 39 310 51
rect 323 39 326 51
rect 344 39 347 51
rect 360 39 363 51
rect 381 39 384 51
rect 397 39 400 51
rect 411 42 423 45
rect 439 39 442 51
rect 455 39 458 51
rect 476 39 479 51
rect 870 51 991 54
rect 1092 55 1095 61
rect 1120 58 1127 61
rect 1131 62 1146 65
rect 1194 58 1201 61
rect 1205 62 1224 65
rect 1224 55 1227 61
rect 1252 58 1259 61
rect 1263 62 1278 65
rect 1326 58 1333 61
rect 1337 62 1356 65
rect 1356 55 1359 61
rect 1384 58 1391 61
rect 1395 62 1412 65
rect 1444 65 1830 69
rect 1834 65 1858 69
rect 1862 65 1888 69
rect 1892 65 1929 69
rect 1480 58 1806 62
rect 1810 58 1857 62
rect 1861 58 1907 62
rect 1911 58 1929 62
rect 559 43 873 47
rect 877 43 909 47
rect 913 43 976 47
rect 980 43 996 47
rect 93 35 126 39
rect 130 35 154 39
rect 158 35 184 39
rect 188 35 258 39
rect 262 35 286 39
rect 290 35 316 39
rect 320 35 390 39
rect 394 35 418 39
rect 422 35 448 39
rect 452 35 505 39
rect 863 36 897 40
rect 901 36 925 40
rect 929 36 955 40
rect 959 36 992 40
rect 1029 39 1032 51
rect 1050 39 1053 51
rect 1066 39 1069 51
rect 1080 42 1092 45
rect 1108 39 1111 51
rect 1124 39 1127 51
rect 1145 39 1148 51
rect 1161 39 1164 51
rect 1182 39 1185 51
rect 1198 39 1201 51
rect 1212 42 1224 45
rect 1240 39 1243 51
rect 1256 39 1259 51
rect 1277 39 1280 51
rect 1293 39 1296 51
rect 1314 39 1317 51
rect 1330 39 1333 51
rect 1344 42 1356 45
rect 1372 39 1375 51
rect 1388 39 1391 51
rect 1409 39 1412 51
rect 1803 51 1924 54
rect 1492 43 1806 47
rect 1810 43 1842 47
rect 1846 43 1909 47
rect 1913 43 1929 47
rect 93 28 102 32
rect 106 28 153 32
rect 157 28 203 32
rect 207 28 234 32
rect 238 28 285 32
rect 289 28 335 32
rect 339 28 366 32
rect 370 28 417 32
rect 421 28 467 32
rect 471 28 541 32
rect 867 26 870 36
rect 888 26 891 36
rect 904 26 907 36
rect 918 29 923 33
rect 927 29 934 33
rect 946 26 949 36
rect 962 26 965 36
rect 983 26 986 36
rect 1026 35 1059 39
rect 1063 35 1087 39
rect 1091 35 1117 39
rect 1121 35 1191 39
rect 1195 35 1219 39
rect 1223 35 1249 39
rect 1253 35 1323 39
rect 1327 35 1351 39
rect 1355 35 1381 39
rect 1385 35 1438 39
rect 1796 36 1830 40
rect 1834 36 1858 40
rect 1862 36 1888 40
rect 1892 36 1925 40
rect 1026 28 1035 32
rect 1039 28 1086 32
rect 1090 28 1136 32
rect 1140 28 1167 32
rect 1171 28 1218 32
rect 1222 28 1268 32
rect 1272 28 1299 32
rect 1303 28 1350 32
rect 1354 28 1400 32
rect 1404 28 1474 32
rect 1800 26 1803 36
rect 1821 26 1824 36
rect 1837 26 1840 36
rect 1851 29 1856 33
rect 1860 29 1867 33
rect 1879 26 1882 36
rect 1895 26 1898 36
rect 1916 26 1919 36
rect 99 21 484 24
rect 93 13 102 17
rect 106 13 138 17
rect 142 13 205 17
rect 209 13 234 17
rect 238 13 270 17
rect 274 13 337 17
rect 341 13 366 17
rect 370 13 402 17
rect 406 13 469 17
rect 473 13 553 17
rect 93 6 126 10
rect 130 6 154 10
rect 158 6 184 10
rect 188 6 221 10
rect 225 6 258 10
rect 262 6 286 10
rect 290 6 316 10
rect 320 6 353 10
rect 357 6 390 10
rect 394 6 418 10
rect 422 6 448 10
rect 452 6 485 10
rect 489 6 493 10
rect 884 12 889 15
rect 893 12 917 15
rect 1032 21 1417 24
rect 942 12 949 15
rect 953 12 975 15
rect 1026 13 1035 17
rect 1039 13 1071 17
rect 1075 13 1138 17
rect 1142 13 1167 17
rect 1171 13 1203 17
rect 1207 13 1270 17
rect 1274 13 1299 17
rect 1303 13 1335 17
rect 1339 13 1402 17
rect 1406 13 1486 17
rect 96 -4 99 6
rect 117 -4 120 6
rect 133 -4 136 6
rect 147 -1 152 3
rect 156 -1 163 3
rect 175 -4 178 6
rect 191 -4 194 6
rect 212 -4 215 6
rect 228 -4 231 6
rect 249 -4 252 6
rect 265 -4 268 6
rect 279 -1 284 3
rect 288 -1 295 3
rect 307 -4 310 6
rect 323 -4 326 6
rect 344 -4 347 6
rect 360 -4 363 6
rect 381 -4 384 6
rect 397 -4 400 6
rect 411 -1 416 3
rect 420 -1 427 3
rect 439 -4 442 6
rect 455 -4 458 6
rect 476 -4 479 6
rect 900 2 907 5
rect 911 6 930 9
rect 113 -18 118 -15
rect 122 -18 146 -15
rect 171 -18 178 -15
rect 182 -18 204 -15
rect 224 -18 231 -15
rect 245 -18 250 -15
rect 254 -18 278 -15
rect 303 -18 310 -15
rect 314 -18 336 -15
rect 356 -18 363 -15
rect 377 -18 382 -15
rect 386 -18 410 -15
rect 435 -18 442 -15
rect 446 -18 468 -15
rect 930 -1 933 5
rect 958 2 965 5
rect 969 6 984 9
rect 995 4 1006 8
rect 1026 6 1059 10
rect 1063 6 1087 10
rect 1091 6 1117 10
rect 1121 6 1154 10
rect 1158 6 1191 10
rect 1195 6 1219 10
rect 1223 6 1249 10
rect 1253 6 1286 10
rect 1290 6 1323 10
rect 1327 6 1351 10
rect 1355 6 1381 10
rect 1385 6 1418 10
rect 1422 6 1426 10
rect 1817 12 1822 15
rect 1826 12 1850 15
rect 1875 12 1882 15
rect 1886 12 1908 15
rect 1029 -4 1032 6
rect 1050 -4 1053 6
rect 1066 -4 1069 6
rect 1080 -1 1085 3
rect 1089 -1 1096 3
rect 1108 -4 1111 6
rect 1124 -4 1127 6
rect 1145 -4 1148 6
rect 1161 -4 1164 6
rect 1182 -4 1185 6
rect 1198 -4 1201 6
rect 1212 -1 1217 3
rect 1221 -1 1228 3
rect 1240 -4 1243 6
rect 1256 -4 1259 6
rect 1277 -4 1280 6
rect 1293 -4 1296 6
rect 1314 -4 1317 6
rect 1330 -4 1333 6
rect 1344 -1 1349 3
rect 1353 -1 1360 3
rect 1372 -4 1375 6
rect 1388 -4 1391 6
rect 1409 -4 1412 6
rect 1833 2 1840 5
rect 1844 6 1863 9
rect 867 -17 870 -5
rect 888 -17 891 -5
rect 904 -17 907 -5
rect 918 -14 930 -11
rect 946 -17 949 -5
rect 962 -17 965 -5
rect 983 -17 986 -5
rect 129 -28 136 -25
rect 140 -24 159 -21
rect 159 -31 162 -25
rect 187 -28 194 -25
rect 198 -24 213 -21
rect 261 -28 268 -25
rect 272 -24 291 -21
rect 291 -31 294 -25
rect 319 -28 326 -25
rect 330 -24 345 -21
rect 393 -28 400 -25
rect 404 -24 423 -21
rect 423 -31 426 -25
rect 451 -28 458 -25
rect 462 -24 479 -21
rect 511 -21 897 -17
rect 901 -21 925 -17
rect 929 -21 955 -17
rect 959 -21 996 -17
rect 1046 -18 1051 -15
rect 1055 -18 1079 -15
rect 1104 -18 1111 -15
rect 1115 -18 1137 -15
rect 1157 -18 1164 -15
rect 1178 -18 1183 -15
rect 1187 -18 1211 -15
rect 1236 -18 1243 -15
rect 1247 -18 1269 -15
rect 1289 -18 1296 -15
rect 1310 -18 1315 -15
rect 1319 -18 1343 -15
rect 1368 -18 1375 -15
rect 1379 -18 1401 -15
rect 1863 -1 1866 5
rect 1891 2 1898 5
rect 1902 6 1917 9
rect 1928 4 1939 8
rect 1800 -17 1803 -5
rect 1821 -17 1824 -5
rect 1837 -17 1840 -5
rect 1851 -14 1863 -11
rect 1879 -17 1882 -5
rect 1895 -17 1898 -5
rect 1916 -17 1919 -5
rect 547 -28 873 -24
rect 877 -28 924 -24
rect 928 -28 974 -24
rect 978 -28 996 -24
rect 1062 -28 1069 -25
rect 1073 -24 1092 -21
rect 1092 -31 1095 -25
rect 1120 -28 1127 -25
rect 1131 -24 1146 -21
rect 1194 -28 1201 -25
rect 1205 -24 1224 -21
rect 1224 -31 1227 -25
rect 1252 -28 1259 -25
rect 1263 -24 1278 -21
rect 1326 -28 1333 -25
rect 1337 -24 1356 -21
rect 1356 -31 1359 -25
rect 1384 -28 1391 -25
rect 1395 -24 1412 -21
rect 1444 -21 1830 -17
rect 1834 -21 1858 -17
rect 1862 -21 1888 -17
rect 1892 -21 1929 -17
rect 1480 -28 1806 -24
rect 1810 -28 1857 -24
rect 1861 -28 1907 -24
rect 1911 -28 1929 -24
rect 96 -47 99 -35
rect 117 -47 120 -35
rect 133 -47 136 -35
rect 147 -44 159 -41
rect 175 -47 178 -35
rect 191 -47 194 -35
rect 212 -47 215 -35
rect 228 -47 231 -35
rect 249 -47 252 -35
rect 265 -47 268 -35
rect 279 -44 291 -41
rect 307 -47 310 -35
rect 323 -47 326 -35
rect 344 -47 347 -35
rect 360 -47 363 -35
rect 381 -47 384 -35
rect 397 -47 400 -35
rect 411 -44 423 -41
rect 439 -47 442 -35
rect 455 -47 458 -35
rect 476 -47 479 -35
rect 1029 -47 1032 -35
rect 1050 -47 1053 -35
rect 1066 -47 1069 -35
rect 1080 -44 1092 -41
rect 1108 -47 1111 -35
rect 1124 -47 1127 -35
rect 1145 -47 1148 -35
rect 1161 -47 1164 -35
rect 1182 -47 1185 -35
rect 1198 -47 1201 -35
rect 1212 -44 1224 -41
rect 1240 -47 1243 -35
rect 1256 -47 1259 -35
rect 1277 -47 1280 -35
rect 1293 -47 1296 -35
rect 1314 -47 1317 -35
rect 1330 -47 1333 -35
rect 1344 -44 1356 -41
rect 1372 -47 1375 -35
rect 1388 -47 1391 -35
rect 1409 -47 1412 -35
rect 93 -51 126 -47
rect 130 -51 154 -47
rect 158 -51 184 -47
rect 188 -51 258 -47
rect 262 -51 286 -47
rect 290 -51 316 -47
rect 320 -51 390 -47
rect 394 -51 418 -47
rect 422 -51 448 -47
rect 452 -51 505 -47
rect 1026 -51 1059 -47
rect 1063 -51 1087 -47
rect 1091 -51 1117 -47
rect 1121 -51 1191 -47
rect 1195 -51 1219 -47
rect 1223 -51 1249 -47
rect 1253 -51 1323 -47
rect 1327 -51 1351 -47
rect 1355 -51 1381 -47
rect 1385 -51 1438 -47
rect 93 -58 102 -54
rect 106 -58 153 -54
rect 157 -58 203 -54
rect 207 -58 234 -54
rect 238 -58 285 -54
rect 289 -58 335 -54
rect 339 -58 366 -54
rect 370 -58 417 -54
rect 421 -58 467 -54
rect 471 -58 541 -54
rect 1026 -58 1035 -54
rect 1039 -58 1086 -54
rect 1090 -58 1136 -54
rect 1140 -58 1167 -54
rect 1171 -58 1218 -54
rect 1222 -58 1268 -54
rect 1272 -58 1299 -54
rect 1303 -58 1350 -54
rect 1354 -58 1400 -54
rect 1404 -58 1474 -54
rect 99 -64 484 -61
rect 1032 -64 1417 -61
rect 224 -71 328 -68
rect 1157 -71 1261 -68
rect 340 -79 344 -75
rect 348 -79 352 -75
rect 1273 -79 1277 -75
rect 1281 -79 1285 -75
rect 76 -90 328 -86
rect 332 -90 348 -86
rect 364 -90 1013 -86
rect 1017 -90 1261 -86
rect 1265 -90 1281 -86
rect 1297 -90 1946 -86
rect 1950 -90 2033 -86
rect 356 -97 484 -94
rect 1289 -97 1417 -94
rect 371 -104 484 -101
rect 1304 -104 1417 -101
rect 340 -113 344 -109
rect 348 -113 352 -109
rect 1273 -113 1277 -109
rect 1281 -113 1285 -109
rect 224 -120 328 -117
rect 1157 -120 1261 -117
rect 93 -127 102 -123
rect 106 -127 138 -123
rect 142 -127 205 -123
rect 209 -127 234 -123
rect 238 -127 270 -123
rect 274 -127 337 -123
rect 341 -127 366 -123
rect 370 -127 402 -123
rect 406 -127 469 -123
rect 473 -127 553 -123
rect 1026 -127 1035 -123
rect 1039 -127 1071 -123
rect 1075 -127 1138 -123
rect 1142 -127 1167 -123
rect 1171 -127 1203 -123
rect 1207 -127 1270 -123
rect 1274 -127 1299 -123
rect 1303 -127 1335 -123
rect 1339 -127 1402 -123
rect 1406 -127 1486 -123
rect 93 -134 126 -130
rect 130 -134 154 -130
rect 158 -134 184 -130
rect 188 -134 221 -130
rect 225 -134 258 -130
rect 262 -134 286 -130
rect 290 -134 316 -130
rect 320 -134 353 -130
rect 357 -134 390 -130
rect 394 -134 418 -130
rect 422 -134 448 -130
rect 452 -134 485 -130
rect 489 -134 493 -130
rect 1026 -134 1059 -130
rect 1063 -134 1087 -130
rect 1091 -134 1117 -130
rect 1121 -134 1154 -130
rect 1158 -134 1191 -130
rect 1195 -134 1219 -130
rect 1223 -134 1249 -130
rect 1253 -134 1286 -130
rect 1290 -134 1323 -130
rect 1327 -134 1351 -130
rect 1355 -134 1381 -130
rect 1385 -134 1418 -130
rect 1422 -134 1426 -130
rect 96 -144 99 -134
rect 117 -144 120 -134
rect 133 -144 136 -134
rect 147 -141 152 -137
rect 156 -141 163 -137
rect 175 -144 178 -134
rect 191 -144 194 -134
rect 212 -144 215 -134
rect 228 -144 231 -134
rect 249 -144 252 -134
rect 265 -144 268 -134
rect 279 -141 284 -137
rect 288 -141 295 -137
rect 307 -144 310 -134
rect 323 -144 326 -134
rect 344 -144 347 -134
rect 360 -144 363 -134
rect 381 -144 384 -134
rect 397 -144 400 -134
rect 411 -141 416 -137
rect 420 -141 427 -137
rect 439 -144 442 -134
rect 455 -144 458 -134
rect 476 -144 479 -134
rect 1029 -144 1032 -134
rect 1050 -144 1053 -134
rect 1066 -144 1069 -134
rect 1080 -141 1085 -137
rect 1089 -141 1096 -137
rect 1108 -144 1111 -134
rect 1124 -144 1127 -134
rect 1145 -144 1148 -134
rect 1161 -144 1164 -134
rect 1182 -144 1185 -134
rect 1198 -144 1201 -134
rect 1212 -141 1217 -137
rect 1221 -141 1228 -137
rect 1240 -144 1243 -134
rect 1256 -144 1259 -134
rect 1277 -144 1280 -134
rect 1293 -144 1296 -134
rect 1314 -144 1317 -134
rect 1330 -144 1333 -134
rect 1344 -141 1349 -137
rect 1353 -141 1360 -137
rect 1372 -144 1375 -134
rect 1388 -144 1391 -134
rect 1409 -144 1412 -134
rect 113 -158 118 -155
rect 122 -158 146 -155
rect 171 -158 178 -155
rect 182 -158 204 -155
rect 224 -158 231 -155
rect 245 -158 250 -155
rect 254 -158 278 -155
rect 303 -158 310 -155
rect 314 -158 336 -155
rect 356 -158 363 -155
rect 377 -158 382 -155
rect 386 -158 410 -155
rect 435 -158 442 -155
rect 446 -158 468 -155
rect 129 -168 136 -165
rect 140 -164 159 -161
rect 159 -171 162 -165
rect 187 -168 194 -165
rect 198 -164 213 -161
rect 261 -168 268 -165
rect 272 -164 291 -161
rect 291 -171 294 -165
rect 319 -168 326 -165
rect 330 -164 345 -161
rect 393 -168 400 -165
rect 404 -164 423 -161
rect 423 -171 426 -165
rect 451 -168 458 -165
rect 462 -164 479 -161
rect 1046 -158 1051 -155
rect 1055 -158 1079 -155
rect 1104 -158 1111 -155
rect 1115 -158 1137 -155
rect 1157 -158 1164 -155
rect 1178 -158 1183 -155
rect 1187 -158 1211 -155
rect 1236 -158 1243 -155
rect 1247 -158 1269 -155
rect 1289 -158 1296 -155
rect 1310 -158 1315 -155
rect 1319 -158 1343 -155
rect 1368 -158 1375 -155
rect 1379 -158 1401 -155
rect 1062 -168 1069 -165
rect 1073 -164 1092 -161
rect 1092 -171 1095 -165
rect 1120 -168 1127 -165
rect 1131 -164 1146 -161
rect 1194 -168 1201 -165
rect 1205 -164 1224 -161
rect 1224 -171 1227 -165
rect 1252 -168 1259 -165
rect 1263 -164 1278 -161
rect 1326 -168 1333 -165
rect 1337 -164 1356 -161
rect 1356 -171 1359 -165
rect 1384 -168 1391 -165
rect 1395 -164 1412 -161
rect 96 -187 99 -175
rect 117 -187 120 -175
rect 133 -187 136 -175
rect 147 -184 159 -181
rect 175 -187 178 -175
rect 191 -187 194 -175
rect 212 -187 215 -175
rect 228 -187 231 -175
rect 249 -187 252 -175
rect 265 -187 268 -175
rect 279 -184 291 -181
rect 307 -187 310 -175
rect 323 -187 326 -175
rect 344 -187 347 -175
rect 360 -187 363 -175
rect 381 -187 384 -175
rect 397 -187 400 -175
rect 411 -184 423 -181
rect 439 -187 442 -175
rect 455 -187 458 -175
rect 476 -187 479 -175
rect 1029 -187 1032 -175
rect 1050 -187 1053 -175
rect 1066 -187 1069 -175
rect 1080 -184 1092 -181
rect 1108 -187 1111 -175
rect 1124 -187 1127 -175
rect 1145 -187 1148 -175
rect 1161 -187 1164 -175
rect 1182 -187 1185 -175
rect 1198 -187 1201 -175
rect 1212 -184 1224 -181
rect 1240 -187 1243 -175
rect 1256 -187 1259 -175
rect 1277 -187 1280 -175
rect 1293 -187 1296 -175
rect 1314 -187 1317 -175
rect 1330 -187 1333 -175
rect 1344 -184 1356 -181
rect 1372 -187 1375 -175
rect 1388 -187 1391 -175
rect 1409 -187 1412 -175
rect 93 -191 126 -187
rect 130 -191 154 -187
rect 158 -191 184 -187
rect 188 -191 258 -187
rect 262 -191 286 -187
rect 290 -191 316 -187
rect 320 -191 390 -187
rect 394 -191 418 -187
rect 422 -191 448 -187
rect 452 -191 505 -187
rect 1026 -191 1059 -187
rect 1063 -191 1087 -187
rect 1091 -191 1117 -187
rect 1121 -191 1191 -187
rect 1195 -191 1219 -187
rect 1223 -191 1249 -187
rect 1253 -191 1323 -187
rect 1327 -191 1351 -187
rect 1355 -191 1381 -187
rect 1385 -191 1438 -187
rect 93 -198 102 -194
rect 106 -198 153 -194
rect 157 -198 203 -194
rect 207 -198 234 -194
rect 238 -198 285 -194
rect 289 -198 335 -194
rect 339 -198 366 -194
rect 370 -198 417 -194
rect 421 -198 467 -194
rect 471 -198 541 -194
rect 1026 -198 1035 -194
rect 1039 -198 1086 -194
rect 1090 -198 1136 -194
rect 1140 -198 1167 -194
rect 1171 -198 1218 -194
rect 1222 -198 1268 -194
rect 1272 -198 1299 -194
rect 1303 -198 1350 -194
rect 1354 -198 1400 -194
rect 1404 -198 1474 -194
<< m2contact >>
rect 553 1754 559 1758
rect 574 1754 578 1758
rect 610 1754 614 1758
rect 677 1754 681 1758
rect 706 1754 710 1758
rect 742 1754 746 1758
rect 809 1754 813 1758
rect 838 1754 842 1758
rect 874 1754 878 1758
rect 941 1754 945 1758
rect 970 1754 974 1758
rect 1006 1754 1010 1758
rect 1073 1754 1077 1758
rect 1486 1754 1492 1758
rect 1507 1754 1511 1758
rect 1543 1754 1547 1758
rect 1610 1754 1614 1758
rect 1639 1754 1643 1758
rect 1675 1754 1679 1758
rect 1742 1754 1746 1758
rect 1771 1754 1775 1758
rect 1807 1754 1811 1758
rect 1874 1754 1878 1758
rect 1903 1754 1907 1758
rect 1939 1754 1943 1758
rect 2006 1754 2010 1758
rect 493 1747 499 1751
rect 1426 1747 1432 1751
rect 574 1740 578 1744
rect 624 1740 628 1744
rect 677 1740 681 1744
rect 706 1740 710 1744
rect 756 1740 760 1744
rect 809 1740 813 1744
rect 838 1740 842 1744
rect 888 1740 892 1744
rect 941 1740 945 1744
rect 970 1740 974 1744
rect 1020 1740 1024 1744
rect 1073 1740 1077 1744
rect 1507 1740 1511 1744
rect 1557 1740 1561 1744
rect 1610 1740 1614 1744
rect 1639 1740 1643 1744
rect 1689 1740 1693 1744
rect 1742 1740 1746 1744
rect 1771 1740 1775 1744
rect 1821 1740 1825 1744
rect 1874 1740 1878 1744
rect 1903 1740 1907 1744
rect 1953 1740 1957 1744
rect 2006 1740 2010 1744
rect 597 1729 601 1733
rect 234 1721 238 1725
rect 270 1721 274 1725
rect 337 1721 341 1725
rect 553 1721 559 1725
rect 568 1720 572 1724
rect 581 1723 585 1729
rect 618 1723 622 1729
rect 631 1725 635 1729
rect 655 1729 659 1733
rect 729 1729 733 1733
rect 639 1723 643 1729
rect 676 1723 680 1729
rect 692 1725 696 1729
rect 493 1714 499 1718
rect 234 1707 238 1711
rect 284 1707 288 1711
rect 337 1707 341 1711
rect 581 1710 585 1714
rect 597 1710 601 1716
rect 631 1716 635 1720
rect 618 1710 622 1714
rect 639 1710 643 1714
rect 655 1710 659 1716
rect 700 1720 704 1724
rect 713 1723 717 1729
rect 750 1723 754 1729
rect 763 1725 767 1729
rect 787 1729 791 1733
rect 861 1729 865 1733
rect 771 1723 775 1729
rect 808 1723 812 1729
rect 824 1725 828 1729
rect 676 1710 680 1714
rect 692 1710 696 1714
rect 713 1710 717 1714
rect 729 1710 733 1716
rect 763 1716 767 1720
rect 750 1710 754 1714
rect 771 1710 775 1714
rect 787 1710 791 1716
rect 832 1720 836 1724
rect 845 1723 849 1729
rect 882 1723 886 1729
rect 895 1725 899 1729
rect 919 1729 923 1733
rect 993 1729 997 1733
rect 903 1723 907 1729
rect 940 1723 944 1729
rect 956 1725 960 1729
rect 808 1710 812 1714
rect 824 1710 828 1714
rect 845 1710 849 1714
rect 861 1710 865 1716
rect 895 1716 899 1720
rect 882 1710 886 1714
rect 903 1710 907 1714
rect 919 1710 923 1716
rect 964 1720 968 1724
rect 977 1723 981 1729
rect 1014 1723 1018 1729
rect 1027 1725 1031 1729
rect 1051 1729 1055 1733
rect 1530 1729 1534 1733
rect 1035 1723 1039 1729
rect 1072 1723 1076 1729
rect 1088 1725 1092 1729
rect 1167 1721 1171 1725
rect 1203 1721 1207 1725
rect 1270 1721 1274 1725
rect 1486 1721 1492 1725
rect 940 1710 944 1714
rect 956 1710 960 1714
rect 977 1710 981 1714
rect 993 1710 997 1716
rect 1027 1716 1031 1720
rect 1014 1710 1018 1714
rect 257 1696 261 1700
rect 219 1687 223 1691
rect 241 1690 245 1696
rect 278 1690 282 1696
rect 291 1692 295 1696
rect 315 1696 319 1700
rect 299 1690 303 1696
rect 336 1690 340 1696
rect 352 1690 356 1696
rect 574 1699 578 1703
rect 611 1697 615 1701
rect 631 1697 635 1701
rect 675 1697 679 1701
rect 706 1699 710 1703
rect 743 1697 747 1701
rect 763 1697 767 1701
rect 807 1697 811 1701
rect 838 1699 842 1703
rect 875 1697 879 1701
rect 895 1697 899 1701
rect 939 1697 943 1701
rect 956 1702 960 1706
rect 1035 1710 1039 1714
rect 1051 1710 1055 1716
rect 1501 1720 1505 1724
rect 1514 1723 1518 1729
rect 1551 1723 1555 1729
rect 1564 1725 1568 1729
rect 1588 1729 1592 1733
rect 1662 1729 1666 1733
rect 1572 1723 1576 1729
rect 1609 1723 1613 1729
rect 1625 1725 1629 1729
rect 1426 1714 1432 1718
rect 1072 1710 1076 1714
rect 1088 1710 1092 1714
rect 970 1699 974 1703
rect 1007 1697 1011 1701
rect 1027 1697 1031 1701
rect 1071 1697 1075 1701
rect 1088 1702 1092 1706
rect 1167 1707 1171 1711
rect 1217 1707 1221 1711
rect 1270 1707 1274 1711
rect 1514 1710 1518 1714
rect 1530 1710 1534 1716
rect 1564 1716 1568 1720
rect 1551 1710 1555 1714
rect 1572 1710 1576 1714
rect 1588 1710 1592 1716
rect 1633 1720 1637 1724
rect 1646 1723 1650 1729
rect 1683 1723 1687 1729
rect 1696 1725 1700 1729
rect 1720 1729 1724 1733
rect 1794 1729 1798 1733
rect 1704 1723 1708 1729
rect 1741 1723 1745 1729
rect 1757 1725 1761 1729
rect 1609 1710 1613 1714
rect 1625 1710 1629 1714
rect 1646 1710 1650 1714
rect 1662 1710 1666 1716
rect 1696 1716 1700 1720
rect 1683 1710 1687 1714
rect 1704 1710 1708 1714
rect 1720 1710 1724 1716
rect 1765 1720 1769 1724
rect 1778 1723 1782 1729
rect 1815 1723 1819 1729
rect 1828 1725 1832 1729
rect 1852 1729 1856 1733
rect 1926 1729 1930 1733
rect 1836 1723 1840 1729
rect 1873 1723 1877 1729
rect 1889 1725 1893 1729
rect 1741 1710 1745 1714
rect 1757 1710 1761 1714
rect 1778 1710 1782 1714
rect 1794 1710 1798 1716
rect 1828 1716 1832 1720
rect 1815 1710 1819 1714
rect 1836 1710 1840 1714
rect 1852 1710 1856 1716
rect 1897 1720 1901 1724
rect 1910 1723 1914 1729
rect 1947 1723 1951 1729
rect 1960 1725 1964 1729
rect 1984 1729 1988 1733
rect 1968 1723 1972 1729
rect 2005 1723 2009 1729
rect 2021 1725 2025 1729
rect 1873 1710 1877 1714
rect 1889 1710 1893 1714
rect 1910 1710 1914 1714
rect 1926 1710 1930 1716
rect 1960 1716 1964 1720
rect 1947 1710 1951 1714
rect 1190 1696 1194 1700
rect 505 1690 511 1694
rect 241 1677 245 1681
rect 257 1677 261 1683
rect 291 1683 295 1687
rect 278 1677 282 1681
rect 299 1677 303 1681
rect 315 1677 319 1683
rect 1152 1687 1156 1691
rect 1174 1690 1178 1696
rect 1211 1690 1215 1696
rect 1224 1692 1228 1696
rect 1248 1696 1252 1700
rect 1232 1690 1236 1696
rect 1269 1690 1273 1696
rect 1285 1690 1289 1696
rect 1507 1699 1511 1703
rect 1544 1697 1548 1701
rect 1564 1697 1568 1701
rect 1608 1697 1612 1701
rect 1639 1699 1643 1703
rect 1676 1697 1680 1701
rect 1696 1697 1700 1701
rect 1740 1697 1744 1701
rect 1771 1699 1775 1703
rect 1808 1697 1812 1701
rect 1828 1697 1832 1701
rect 1872 1697 1876 1701
rect 1889 1702 1893 1706
rect 1968 1710 1972 1714
rect 1984 1710 1988 1716
rect 2005 1710 2009 1714
rect 2021 1710 2025 1714
rect 1903 1699 1907 1703
rect 1940 1697 1944 1701
rect 1960 1697 1964 1701
rect 2004 1697 2008 1701
rect 2021 1702 2025 1706
rect 1438 1690 1444 1694
rect 541 1683 547 1687
rect 574 1683 578 1687
rect 625 1683 629 1687
rect 675 1683 679 1687
rect 706 1683 710 1687
rect 757 1683 761 1687
rect 807 1683 811 1687
rect 838 1683 842 1687
rect 889 1683 893 1687
rect 939 1683 943 1687
rect 970 1683 974 1687
rect 1021 1683 1025 1687
rect 1071 1683 1075 1687
rect 336 1677 340 1681
rect 352 1677 356 1681
rect 1174 1677 1178 1681
rect 1190 1677 1194 1683
rect 1224 1683 1228 1687
rect 1211 1677 1215 1681
rect 234 1666 238 1670
rect 271 1664 275 1668
rect 291 1664 295 1668
rect 335 1664 339 1668
rect 493 1670 499 1674
rect 572 1670 576 1674
rect 606 1670 610 1674
rect 623 1670 627 1674
rect 679 1670 683 1674
rect 696 1670 700 1674
rect 724 1670 728 1674
rect 1232 1677 1236 1681
rect 1248 1677 1252 1683
rect 1474 1683 1480 1687
rect 1507 1683 1511 1687
rect 1558 1683 1562 1687
rect 1608 1683 1612 1687
rect 1639 1683 1643 1687
rect 1690 1683 1694 1687
rect 1740 1683 1744 1687
rect 1771 1683 1775 1687
rect 1822 1683 1826 1687
rect 1872 1683 1876 1687
rect 1903 1683 1907 1687
rect 1954 1683 1958 1687
rect 2004 1683 2008 1687
rect 1269 1677 1273 1681
rect 1285 1677 1289 1681
rect 529 1663 535 1667
rect 599 1663 603 1667
rect 630 1663 634 1667
rect 652 1663 656 1667
rect 717 1663 721 1667
rect 505 1657 511 1661
rect 234 1650 238 1654
rect 285 1650 289 1654
rect 335 1650 339 1654
rect 541 1650 547 1654
rect 573 1653 577 1657
rect 598 1656 602 1660
rect 605 1653 609 1657
rect 623 1653 627 1657
rect 645 1656 649 1660
rect 670 1656 674 1660
rect 680 1653 684 1657
rect 696 1653 700 1657
rect 716 1656 720 1660
rect 723 1653 727 1657
rect 787 1663 791 1667
rect 352 1643 356 1647
rect 219 1634 223 1638
rect 344 1636 348 1640
rect 368 1636 372 1640
rect 227 1627 231 1631
rect 368 1627 372 1631
rect 600 1637 604 1641
rect 620 1634 624 1638
rect 639 1638 643 1642
rect 741 1649 745 1653
rect 756 1649 760 1653
rect 658 1637 662 1641
rect 677 1637 681 1641
rect 690 1636 694 1640
rect 712 1637 716 1641
rect 720 1636 724 1640
rect 732 1636 736 1640
rect 573 1623 577 1627
rect 605 1623 609 1627
rect 623 1623 627 1627
rect 680 1623 684 1627
rect 695 1623 699 1627
rect 723 1623 727 1627
rect 234 1619 238 1623
rect 301 1619 305 1623
rect 337 1619 341 1623
rect 553 1619 559 1623
rect 587 1619 591 1623
rect 630 1618 634 1622
rect 652 1619 659 1623
rect 702 1618 706 1622
rect 493 1612 499 1616
rect 234 1605 238 1609
rect 287 1605 291 1609
rect 337 1605 341 1609
rect 517 1611 523 1615
rect 587 1611 591 1615
rect 646 1611 650 1615
rect 671 1611 675 1615
rect 702 1611 706 1615
rect 795 1641 799 1649
rect 868 1663 872 1667
rect 822 1649 826 1653
rect 837 1649 841 1653
rect 1167 1666 1171 1670
rect 1204 1664 1208 1668
rect 1224 1664 1228 1668
rect 1268 1664 1272 1668
rect 1426 1670 1432 1674
rect 1505 1670 1509 1674
rect 1539 1670 1543 1674
rect 1556 1670 1560 1674
rect 1612 1670 1616 1674
rect 1629 1670 1633 1674
rect 1657 1670 1661 1674
rect 1462 1663 1468 1667
rect 1532 1663 1536 1667
rect 1563 1663 1567 1667
rect 1585 1663 1589 1667
rect 1650 1663 1654 1667
rect 818 1641 822 1645
rect 764 1635 768 1639
rect 777 1627 781 1631
rect 876 1641 880 1649
rect 1438 1657 1444 1661
rect 1167 1650 1171 1654
rect 1218 1650 1222 1654
rect 1268 1650 1272 1654
rect 1474 1650 1480 1654
rect 1506 1653 1510 1657
rect 1531 1656 1535 1660
rect 1538 1653 1542 1657
rect 1556 1653 1560 1657
rect 1578 1656 1582 1660
rect 1603 1656 1607 1660
rect 1613 1653 1617 1657
rect 1629 1653 1633 1657
rect 1649 1656 1653 1660
rect 1656 1653 1660 1657
rect 1720 1663 1724 1667
rect 903 1641 907 1645
rect 1285 1643 1289 1647
rect 845 1635 849 1639
rect 1152 1634 1156 1638
rect 1277 1636 1281 1640
rect 1301 1636 1305 1640
rect 858 1627 862 1631
rect 1160 1627 1164 1631
rect 1301 1627 1305 1631
rect 1533 1637 1537 1641
rect 1553 1634 1557 1638
rect 1572 1638 1576 1642
rect 1674 1649 1678 1653
rect 1689 1649 1693 1653
rect 1591 1637 1595 1641
rect 1610 1637 1614 1641
rect 1623 1636 1627 1640
rect 1645 1637 1649 1641
rect 1653 1636 1657 1640
rect 1665 1636 1669 1640
rect 1506 1623 1510 1627
rect 1538 1623 1542 1627
rect 1556 1623 1560 1627
rect 1613 1623 1617 1627
rect 1628 1623 1632 1627
rect 1656 1623 1660 1627
rect 1167 1619 1171 1623
rect 1234 1619 1238 1623
rect 1270 1619 1274 1623
rect 1486 1619 1492 1623
rect 1520 1619 1524 1623
rect 1563 1618 1567 1622
rect 1585 1619 1592 1623
rect 1635 1618 1639 1622
rect 1426 1612 1432 1616
rect 505 1604 511 1608
rect 573 1604 577 1608
rect 587 1604 591 1608
rect 605 1604 609 1608
rect 623 1604 627 1608
rect 646 1604 650 1608
rect 680 1604 684 1608
rect 695 1604 699 1608
rect 723 1604 727 1608
rect 256 1594 260 1598
rect 219 1588 223 1594
rect 235 1588 239 1594
rect 272 1588 276 1594
rect 280 1590 284 1594
rect 314 1594 318 1598
rect 517 1597 523 1601
rect 587 1597 591 1601
rect 646 1597 650 1601
rect 671 1597 675 1601
rect 702 1597 706 1601
rect 293 1588 297 1594
rect 330 1588 334 1594
rect 587 1589 591 1593
rect 630 1590 634 1594
rect 652 1589 659 1593
rect 702 1590 706 1594
rect 352 1585 356 1589
rect 573 1585 577 1589
rect 605 1585 609 1589
rect 623 1585 627 1589
rect 680 1585 684 1589
rect 695 1585 699 1589
rect 723 1585 727 1589
rect 219 1575 223 1579
rect 235 1575 239 1579
rect 280 1581 284 1585
rect 256 1575 260 1581
rect 272 1575 276 1579
rect 293 1575 297 1579
rect 314 1575 318 1581
rect 330 1575 334 1579
rect 568 1573 572 1577
rect 236 1562 240 1566
rect 280 1562 284 1566
rect 300 1562 304 1566
rect 337 1564 341 1568
rect 600 1571 604 1575
rect 620 1574 624 1578
rect 639 1570 643 1574
rect 658 1571 662 1575
rect 677 1571 681 1575
rect 690 1572 694 1576
rect 787 1587 791 1591
rect 1167 1605 1171 1609
rect 1220 1605 1224 1609
rect 1270 1605 1274 1609
rect 1450 1611 1456 1615
rect 1520 1611 1524 1615
rect 1579 1611 1583 1615
rect 1604 1611 1608 1615
rect 1635 1611 1639 1615
rect 1728 1641 1732 1649
rect 1801 1663 1805 1667
rect 1755 1649 1759 1653
rect 1770 1649 1774 1653
rect 1751 1641 1755 1645
rect 1697 1635 1701 1639
rect 1710 1627 1714 1631
rect 1809 1641 1813 1649
rect 1836 1641 1840 1645
rect 1778 1635 1782 1639
rect 1791 1627 1795 1631
rect 1438 1604 1444 1608
rect 1506 1604 1510 1608
rect 1520 1604 1524 1608
rect 1538 1604 1542 1608
rect 1556 1604 1560 1608
rect 1579 1604 1583 1608
rect 1613 1604 1617 1608
rect 1628 1604 1632 1608
rect 1656 1604 1660 1608
rect 1189 1594 1193 1598
rect 868 1587 872 1591
rect 1152 1588 1156 1594
rect 1168 1588 1172 1594
rect 1205 1588 1209 1594
rect 1213 1590 1217 1594
rect 1247 1594 1251 1598
rect 1450 1597 1456 1601
rect 1520 1597 1524 1601
rect 1579 1597 1583 1601
rect 1604 1597 1608 1601
rect 1635 1597 1639 1601
rect 1226 1588 1230 1594
rect 1263 1588 1267 1594
rect 1520 1589 1524 1593
rect 1563 1590 1567 1594
rect 1585 1589 1592 1593
rect 1635 1590 1639 1594
rect 1285 1585 1289 1589
rect 1506 1585 1510 1589
rect 1538 1585 1542 1589
rect 1556 1585 1560 1589
rect 1613 1585 1617 1589
rect 1628 1585 1632 1589
rect 1656 1585 1660 1589
rect 712 1571 716 1575
rect 720 1572 724 1576
rect 732 1572 736 1576
rect 767 1572 771 1576
rect 795 1571 799 1575
rect 847 1572 851 1576
rect 1152 1575 1156 1579
rect 1168 1575 1172 1579
rect 1213 1581 1217 1585
rect 1189 1575 1193 1581
rect 1205 1575 1209 1579
rect 876 1571 880 1575
rect 1226 1575 1230 1579
rect 1247 1575 1251 1581
rect 1263 1575 1267 1579
rect 1501 1573 1505 1577
rect 505 1555 511 1559
rect 573 1555 577 1559
rect 598 1552 602 1556
rect 605 1555 609 1559
rect 623 1555 627 1559
rect 645 1552 649 1556
rect 670 1552 674 1556
rect 680 1555 684 1559
rect 696 1555 700 1559
rect 716 1552 720 1556
rect 723 1555 727 1559
rect 236 1548 240 1552
rect 286 1548 290 1552
rect 337 1548 341 1552
rect 541 1548 547 1552
rect 583 1545 587 1549
rect 599 1545 603 1549
rect 630 1545 634 1549
rect 652 1545 656 1549
rect 717 1545 721 1549
rect 777 1551 781 1555
rect 1169 1562 1173 1566
rect 1213 1562 1217 1566
rect 1233 1562 1237 1566
rect 1270 1564 1274 1568
rect 1533 1571 1537 1575
rect 1553 1574 1557 1578
rect 1572 1570 1576 1574
rect 1591 1571 1595 1575
rect 1610 1571 1614 1575
rect 1623 1572 1627 1576
rect 1720 1587 1724 1591
rect 1801 1587 1805 1591
rect 1645 1571 1649 1575
rect 1653 1572 1657 1576
rect 1665 1572 1669 1576
rect 1700 1572 1704 1576
rect 1728 1571 1732 1575
rect 1780 1572 1784 1576
rect 1809 1571 1813 1575
rect 1438 1555 1444 1559
rect 1506 1555 1510 1559
rect 858 1551 862 1555
rect 1531 1552 1535 1556
rect 1538 1555 1542 1559
rect 1556 1555 1560 1559
rect 1578 1552 1582 1556
rect 1603 1552 1607 1556
rect 1613 1555 1617 1559
rect 1629 1555 1633 1559
rect 1649 1552 1653 1556
rect 1656 1555 1660 1559
rect 1169 1548 1173 1552
rect 1219 1548 1223 1552
rect 1270 1548 1274 1552
rect 1474 1548 1480 1552
rect 1516 1545 1520 1549
rect 1532 1545 1536 1549
rect 1563 1545 1567 1549
rect 1585 1545 1589 1549
rect 1650 1545 1654 1549
rect 1710 1551 1714 1555
rect 1791 1551 1795 1555
rect 493 1538 499 1542
rect 572 1538 576 1542
rect 606 1538 610 1542
rect 623 1538 627 1542
rect 679 1538 683 1542
rect 696 1538 700 1542
rect 724 1538 728 1542
rect 1426 1538 1432 1542
rect 1505 1538 1509 1542
rect 1539 1538 1543 1542
rect 1556 1538 1560 1542
rect 1612 1538 1616 1542
rect 1629 1538 1633 1542
rect 1657 1538 1661 1542
rect 529 1531 535 1535
rect 583 1531 587 1535
rect 599 1531 603 1535
rect 630 1531 634 1535
rect 652 1531 656 1535
rect 717 1531 721 1535
rect 787 1531 791 1535
rect 573 1521 577 1525
rect 598 1524 602 1528
rect 605 1521 609 1525
rect 623 1521 627 1525
rect 645 1524 649 1528
rect 670 1524 674 1528
rect 680 1521 684 1525
rect 696 1521 700 1525
rect 716 1524 720 1528
rect 723 1521 727 1525
rect 567 1504 571 1508
rect 600 1505 604 1509
rect 620 1502 624 1506
rect 639 1506 643 1510
rect 658 1505 662 1509
rect 677 1505 681 1509
rect 690 1504 694 1508
rect 712 1505 716 1509
rect 720 1504 724 1508
rect 732 1504 736 1508
rect 795 1509 799 1517
rect 892 1531 896 1535
rect 846 1517 850 1521
rect 861 1517 865 1521
rect 1462 1531 1468 1535
rect 1516 1531 1520 1535
rect 1532 1531 1536 1535
rect 1563 1531 1567 1535
rect 1585 1531 1589 1535
rect 1650 1531 1654 1535
rect 1720 1531 1724 1535
rect 764 1503 768 1507
rect 818 1508 822 1512
rect 573 1491 577 1495
rect 605 1491 609 1495
rect 623 1491 627 1495
rect 680 1491 684 1495
rect 695 1491 699 1495
rect 723 1491 727 1495
rect 587 1487 591 1491
rect 630 1486 634 1490
rect 652 1487 659 1491
rect 702 1486 706 1490
rect 517 1479 523 1483
rect 587 1479 591 1483
rect 646 1479 650 1483
rect 671 1479 675 1483
rect 702 1479 706 1483
rect 777 1495 781 1499
rect 900 1509 904 1517
rect 1506 1521 1510 1525
rect 1531 1524 1535 1528
rect 1538 1521 1542 1525
rect 1556 1521 1560 1525
rect 1578 1524 1582 1528
rect 1603 1524 1607 1528
rect 1613 1521 1617 1525
rect 1629 1521 1633 1525
rect 1649 1524 1653 1528
rect 1656 1521 1660 1525
rect 921 1509 925 1513
rect 869 1503 873 1507
rect 1500 1504 1504 1508
rect 882 1495 886 1499
rect 1533 1505 1537 1509
rect 1553 1502 1557 1506
rect 1572 1506 1576 1510
rect 1591 1505 1595 1509
rect 1610 1505 1614 1509
rect 1623 1504 1627 1508
rect 1645 1505 1649 1509
rect 1653 1504 1657 1508
rect 1665 1504 1669 1508
rect 1728 1509 1732 1517
rect 1825 1531 1829 1535
rect 1779 1517 1783 1521
rect 1794 1517 1798 1521
rect 1697 1503 1701 1507
rect 1751 1508 1755 1512
rect 1506 1491 1510 1495
rect 1538 1491 1542 1495
rect 1556 1491 1560 1495
rect 1613 1491 1617 1495
rect 1628 1491 1632 1495
rect 1656 1491 1660 1495
rect 1520 1487 1524 1491
rect 1563 1486 1567 1490
rect 1585 1487 1592 1491
rect 1635 1486 1639 1490
rect 1450 1479 1456 1483
rect 1520 1479 1524 1483
rect 1579 1479 1583 1483
rect 1604 1479 1608 1483
rect 1635 1479 1639 1483
rect 1710 1495 1714 1499
rect 1833 1509 1837 1517
rect 1854 1509 1858 1513
rect 1802 1503 1806 1507
rect 1815 1495 1819 1499
rect 505 1472 511 1476
rect 573 1472 577 1476
rect 587 1472 591 1476
rect 605 1472 609 1476
rect 623 1472 627 1476
rect 646 1472 650 1476
rect 680 1472 684 1476
rect 695 1472 699 1476
rect 723 1472 727 1476
rect 1438 1472 1444 1476
rect 1506 1472 1510 1476
rect 1520 1472 1524 1476
rect 1538 1472 1542 1476
rect 1556 1472 1560 1476
rect 1579 1472 1583 1476
rect 1613 1472 1617 1476
rect 1628 1472 1632 1476
rect 1656 1472 1660 1476
rect 517 1465 523 1469
rect 587 1465 591 1469
rect 646 1465 650 1469
rect 671 1465 675 1469
rect 702 1465 706 1469
rect 587 1457 591 1461
rect 630 1458 634 1462
rect 652 1457 659 1461
rect 702 1458 706 1462
rect 573 1453 577 1457
rect 605 1453 609 1457
rect 623 1453 627 1457
rect 680 1453 684 1457
rect 695 1453 699 1457
rect 723 1453 727 1457
rect 787 1456 791 1460
rect 1450 1465 1456 1469
rect 1520 1465 1524 1469
rect 1579 1465 1583 1469
rect 1604 1465 1608 1469
rect 1635 1465 1639 1469
rect 892 1456 896 1460
rect 1520 1457 1524 1461
rect 1563 1458 1567 1462
rect 1585 1457 1592 1461
rect 1635 1458 1639 1462
rect 1506 1453 1510 1457
rect 1538 1453 1542 1457
rect 1556 1453 1560 1457
rect 1613 1453 1617 1457
rect 1628 1453 1632 1457
rect 1656 1453 1660 1457
rect 1720 1456 1724 1460
rect 1825 1456 1829 1460
rect 568 1441 572 1445
rect 600 1439 604 1443
rect 620 1442 624 1446
rect 639 1438 643 1442
rect 658 1439 662 1443
rect 677 1439 681 1443
rect 690 1440 694 1444
rect 712 1439 716 1443
rect 720 1440 724 1444
rect 732 1440 736 1444
rect 766 1441 770 1445
rect 795 1440 799 1444
rect 872 1441 876 1445
rect 900 1440 904 1444
rect 1501 1441 1505 1445
rect 573 1423 577 1427
rect 598 1420 602 1424
rect 605 1423 609 1427
rect 623 1423 627 1427
rect 645 1420 649 1424
rect 670 1420 674 1424
rect 680 1423 684 1427
rect 696 1423 700 1427
rect 716 1420 720 1424
rect 723 1423 727 1427
rect 529 1413 535 1417
rect 599 1413 603 1417
rect 630 1413 634 1417
rect 652 1413 656 1417
rect 717 1413 721 1417
rect 777 1420 781 1424
rect 1533 1439 1537 1443
rect 1553 1442 1557 1446
rect 1572 1438 1576 1442
rect 1591 1439 1595 1443
rect 1610 1439 1614 1443
rect 1623 1440 1627 1444
rect 1645 1439 1649 1443
rect 1653 1440 1657 1444
rect 1665 1440 1669 1444
rect 1699 1441 1703 1445
rect 1728 1440 1732 1444
rect 1805 1441 1809 1445
rect 1833 1440 1837 1444
rect 882 1420 886 1424
rect 1506 1423 1510 1427
rect 1531 1420 1535 1424
rect 1538 1423 1542 1427
rect 1556 1423 1560 1427
rect 1578 1420 1582 1424
rect 1603 1420 1607 1424
rect 1613 1423 1617 1427
rect 1629 1423 1633 1427
rect 1649 1420 1653 1424
rect 1656 1423 1660 1427
rect 1462 1413 1468 1417
rect 1532 1413 1536 1417
rect 1563 1413 1567 1417
rect 1585 1413 1589 1417
rect 1650 1413 1654 1417
rect 1710 1420 1714 1424
rect 1815 1420 1819 1424
rect 493 1406 499 1410
rect 572 1406 576 1410
rect 606 1406 610 1410
rect 623 1406 627 1410
rect 679 1406 683 1410
rect 696 1406 700 1410
rect 724 1406 728 1410
rect 1426 1406 1432 1410
rect 1505 1406 1509 1410
rect 1539 1406 1543 1410
rect 1556 1406 1560 1410
rect 1612 1406 1616 1410
rect 1629 1406 1633 1410
rect 1657 1406 1661 1410
rect 529 1399 535 1403
rect 599 1399 603 1403
rect 630 1399 634 1403
rect 652 1399 656 1403
rect 717 1399 721 1403
rect 787 1399 791 1403
rect 573 1389 577 1393
rect 598 1392 602 1396
rect 605 1389 609 1393
rect 623 1389 627 1393
rect 645 1392 649 1396
rect 670 1392 674 1396
rect 680 1389 684 1393
rect 696 1389 700 1393
rect 716 1392 720 1396
rect 723 1389 727 1393
rect 567 1372 571 1376
rect 600 1373 604 1377
rect 620 1370 624 1374
rect 639 1374 643 1378
rect 658 1373 662 1377
rect 677 1373 681 1377
rect 690 1372 694 1376
rect 712 1373 716 1377
rect 720 1372 724 1376
rect 732 1372 736 1376
rect 795 1377 799 1385
rect 868 1399 872 1403
rect 822 1385 826 1389
rect 837 1385 841 1389
rect 818 1377 822 1381
rect 764 1371 768 1375
rect 573 1359 577 1363
rect 605 1359 609 1363
rect 623 1359 627 1363
rect 680 1359 684 1363
rect 695 1359 699 1363
rect 723 1359 727 1363
rect 587 1355 591 1359
rect 630 1354 634 1358
rect 652 1355 659 1359
rect 702 1354 706 1358
rect 517 1347 523 1351
rect 587 1347 591 1351
rect 646 1347 650 1351
rect 671 1347 675 1351
rect 702 1347 706 1351
rect 777 1363 781 1367
rect 876 1377 880 1385
rect 958 1399 962 1403
rect 912 1385 916 1389
rect 927 1385 931 1389
rect 1462 1399 1468 1403
rect 1532 1399 1536 1403
rect 1563 1399 1567 1403
rect 1585 1399 1589 1403
rect 1650 1399 1654 1403
rect 1720 1399 1724 1403
rect 900 1377 904 1381
rect 845 1371 849 1375
rect 934 1379 938 1383
rect 966 1377 970 1385
rect 1506 1389 1510 1393
rect 1531 1392 1535 1396
rect 1538 1389 1542 1393
rect 1556 1389 1560 1393
rect 1578 1392 1582 1396
rect 1603 1392 1607 1396
rect 1613 1389 1617 1393
rect 1629 1389 1633 1393
rect 1649 1392 1653 1396
rect 1656 1389 1660 1393
rect 858 1363 862 1367
rect 1001 1376 1005 1380
rect 1500 1372 1504 1376
rect 948 1363 952 1367
rect 1533 1373 1537 1377
rect 1553 1370 1557 1374
rect 1572 1374 1576 1378
rect 1591 1373 1595 1377
rect 1610 1373 1614 1377
rect 1623 1372 1627 1376
rect 1645 1373 1649 1377
rect 1653 1372 1657 1376
rect 1665 1372 1669 1376
rect 1728 1377 1732 1385
rect 1801 1399 1805 1403
rect 1755 1385 1759 1389
rect 1770 1385 1774 1389
rect 1751 1377 1755 1381
rect 1697 1371 1701 1375
rect 1506 1359 1510 1363
rect 1538 1359 1542 1363
rect 1556 1359 1560 1363
rect 1613 1359 1617 1363
rect 1628 1359 1632 1363
rect 1656 1359 1660 1363
rect 1520 1355 1524 1359
rect 1563 1354 1567 1358
rect 1585 1355 1592 1359
rect 1635 1354 1639 1358
rect 1450 1347 1456 1351
rect 1520 1347 1524 1351
rect 1579 1347 1583 1351
rect 1604 1347 1608 1351
rect 1635 1347 1639 1351
rect 1710 1363 1714 1367
rect 1809 1377 1813 1385
rect 1891 1399 1895 1403
rect 1845 1385 1849 1389
rect 1860 1385 1864 1389
rect 1833 1377 1837 1381
rect 1778 1371 1782 1375
rect 1867 1379 1871 1383
rect 1899 1377 1903 1385
rect 1791 1363 1795 1367
rect 1934 1376 1938 1380
rect 1881 1363 1885 1367
rect 505 1340 511 1344
rect 573 1340 577 1344
rect 587 1340 591 1344
rect 605 1340 609 1344
rect 623 1340 627 1344
rect 646 1340 650 1344
rect 680 1340 684 1344
rect 695 1340 699 1344
rect 723 1340 727 1344
rect 1438 1340 1444 1344
rect 1506 1340 1510 1344
rect 1520 1340 1524 1344
rect 1538 1340 1542 1344
rect 1556 1340 1560 1344
rect 1579 1340 1583 1344
rect 1613 1340 1617 1344
rect 1628 1340 1632 1344
rect 1656 1340 1660 1344
rect 517 1333 523 1337
rect 587 1333 591 1337
rect 646 1333 650 1337
rect 671 1333 675 1337
rect 702 1333 706 1337
rect 587 1325 591 1329
rect 630 1326 634 1330
rect 652 1325 659 1329
rect 702 1326 706 1330
rect 573 1321 577 1325
rect 605 1321 609 1325
rect 623 1321 627 1325
rect 680 1321 684 1325
rect 695 1321 699 1325
rect 723 1321 727 1325
rect 568 1309 572 1313
rect 600 1307 604 1311
rect 620 1310 624 1314
rect 639 1306 643 1310
rect 658 1307 662 1311
rect 677 1307 681 1311
rect 690 1308 694 1312
rect 787 1321 791 1325
rect 868 1321 872 1325
rect 1450 1333 1456 1337
rect 1520 1333 1524 1337
rect 1579 1333 1583 1337
rect 1604 1333 1608 1337
rect 1635 1333 1639 1337
rect 1520 1325 1524 1329
rect 1563 1326 1567 1330
rect 1585 1325 1592 1329
rect 1635 1326 1639 1330
rect 958 1321 962 1325
rect 1506 1321 1510 1325
rect 1538 1321 1542 1325
rect 1556 1321 1560 1325
rect 1613 1321 1617 1325
rect 1628 1321 1632 1325
rect 1656 1321 1660 1325
rect 712 1307 716 1311
rect 720 1308 724 1312
rect 732 1308 736 1312
rect 767 1306 771 1310
rect 795 1305 799 1309
rect 847 1306 851 1310
rect 876 1305 880 1309
rect 931 1306 935 1310
rect 1501 1309 1505 1313
rect 966 1305 970 1309
rect 573 1291 577 1295
rect 598 1288 602 1292
rect 605 1291 609 1295
rect 623 1291 627 1295
rect 645 1288 649 1292
rect 670 1288 674 1292
rect 680 1291 684 1295
rect 696 1291 700 1295
rect 716 1288 720 1292
rect 723 1291 727 1295
rect 1533 1307 1537 1311
rect 1553 1310 1557 1314
rect 1572 1306 1576 1310
rect 1591 1307 1595 1311
rect 1610 1307 1614 1311
rect 1623 1308 1627 1312
rect 1720 1321 1724 1325
rect 1801 1321 1805 1325
rect 1891 1321 1895 1325
rect 1645 1307 1649 1311
rect 1653 1308 1657 1312
rect 1665 1308 1669 1312
rect 1700 1306 1704 1310
rect 1728 1305 1732 1309
rect 1780 1306 1784 1310
rect 1809 1305 1813 1309
rect 1864 1306 1868 1310
rect 1899 1305 1903 1309
rect 529 1281 535 1285
rect 599 1281 603 1285
rect 630 1281 634 1285
rect 652 1281 656 1285
rect 717 1281 721 1285
rect 777 1285 781 1289
rect 858 1285 862 1289
rect 1506 1291 1510 1295
rect 948 1285 952 1289
rect 1531 1288 1535 1292
rect 1538 1291 1542 1295
rect 1556 1291 1560 1295
rect 1578 1288 1582 1292
rect 1603 1288 1607 1292
rect 1613 1291 1617 1295
rect 1629 1291 1633 1295
rect 1649 1288 1653 1292
rect 1656 1291 1660 1295
rect 1462 1281 1468 1285
rect 1532 1281 1536 1285
rect 1563 1281 1567 1285
rect 1585 1281 1589 1285
rect 1650 1281 1654 1285
rect 1710 1285 1714 1289
rect 1791 1285 1795 1289
rect 1881 1285 1885 1289
rect 493 1274 499 1278
rect 572 1274 576 1278
rect 606 1274 610 1278
rect 623 1274 627 1278
rect 679 1274 683 1278
rect 696 1274 700 1278
rect 724 1274 728 1278
rect 1426 1274 1432 1278
rect 1505 1274 1509 1278
rect 1539 1274 1543 1278
rect 1556 1274 1560 1278
rect 1612 1274 1616 1278
rect 1629 1274 1633 1278
rect 1657 1274 1661 1278
rect 529 1267 535 1271
rect 599 1267 603 1271
rect 630 1267 634 1271
rect 652 1267 656 1271
rect 717 1267 721 1271
rect 787 1267 791 1271
rect 573 1257 577 1261
rect 598 1260 602 1264
rect 605 1257 609 1261
rect 623 1257 627 1261
rect 645 1260 649 1264
rect 670 1260 674 1264
rect 680 1257 684 1261
rect 696 1257 700 1261
rect 716 1260 720 1264
rect 723 1257 727 1261
rect 567 1240 571 1244
rect 600 1241 604 1245
rect 620 1238 624 1242
rect 639 1242 643 1246
rect 1462 1267 1468 1271
rect 1532 1267 1536 1271
rect 1563 1267 1567 1271
rect 1585 1267 1589 1271
rect 1650 1267 1654 1271
rect 1720 1267 1724 1271
rect 658 1241 662 1245
rect 677 1241 681 1245
rect 690 1240 694 1244
rect 712 1241 716 1245
rect 720 1240 724 1244
rect 732 1240 736 1244
rect 795 1245 799 1253
rect 1506 1257 1510 1261
rect 1531 1260 1535 1264
rect 1538 1257 1542 1261
rect 1556 1257 1560 1261
rect 1578 1260 1582 1264
rect 1603 1260 1607 1264
rect 1613 1257 1617 1261
rect 1629 1257 1633 1261
rect 1649 1260 1653 1264
rect 1656 1257 1660 1261
rect 764 1239 768 1243
rect 818 1244 822 1248
rect 1500 1240 1504 1244
rect 573 1227 577 1231
rect 605 1227 609 1231
rect 623 1227 627 1231
rect 680 1227 684 1231
rect 695 1227 699 1231
rect 723 1227 727 1231
rect 587 1223 591 1227
rect 102 1219 106 1223
rect 138 1219 142 1223
rect 205 1219 209 1223
rect 234 1219 238 1223
rect 270 1219 274 1223
rect 337 1219 341 1223
rect 366 1219 370 1223
rect 402 1219 406 1223
rect 469 1219 473 1223
rect 553 1219 559 1223
rect 630 1222 634 1226
rect 652 1223 659 1227
rect 702 1222 706 1226
rect 493 1212 499 1216
rect 587 1215 591 1219
rect 596 1215 600 1219
rect 646 1215 650 1219
rect 671 1215 675 1219
rect 702 1215 706 1219
rect 777 1231 781 1235
rect 1533 1241 1537 1245
rect 1553 1238 1557 1242
rect 1572 1242 1576 1246
rect 1591 1241 1595 1245
rect 1610 1241 1614 1245
rect 1623 1240 1627 1244
rect 1645 1241 1649 1245
rect 1653 1240 1657 1244
rect 1665 1240 1669 1244
rect 1728 1245 1732 1253
rect 1697 1239 1701 1243
rect 1751 1244 1755 1248
rect 1506 1227 1510 1231
rect 1538 1227 1542 1231
rect 1556 1227 1560 1231
rect 1613 1227 1617 1231
rect 1628 1227 1632 1231
rect 1656 1227 1660 1231
rect 1520 1223 1524 1227
rect 1035 1219 1039 1223
rect 1071 1219 1075 1223
rect 1138 1219 1142 1223
rect 1167 1219 1171 1223
rect 1203 1219 1207 1223
rect 1270 1219 1274 1223
rect 1299 1219 1303 1223
rect 1335 1219 1339 1223
rect 1402 1219 1406 1223
rect 1486 1219 1492 1223
rect 1563 1222 1567 1226
rect 1585 1223 1592 1227
rect 1635 1222 1639 1226
rect 1426 1212 1432 1216
rect 1520 1215 1524 1219
rect 1529 1215 1533 1219
rect 1579 1215 1583 1219
rect 1604 1215 1608 1219
rect 1635 1215 1639 1219
rect 1710 1231 1714 1235
rect 102 1205 106 1209
rect 152 1205 156 1209
rect 205 1205 209 1209
rect 234 1205 238 1209
rect 284 1205 288 1209
rect 337 1205 341 1209
rect 366 1205 370 1209
rect 416 1205 420 1209
rect 469 1205 473 1209
rect 505 1208 511 1212
rect 573 1208 577 1212
rect 587 1208 591 1212
rect 605 1208 609 1212
rect 623 1208 627 1212
rect 646 1208 650 1212
rect 680 1208 684 1212
rect 695 1208 699 1212
rect 723 1208 727 1212
rect 848 1208 852 1212
rect 866 1208 870 1212
rect 884 1208 888 1212
rect 907 1208 911 1212
rect 941 1208 945 1212
rect 956 1208 960 1212
rect 984 1208 988 1212
rect 125 1194 129 1198
rect 96 1185 100 1189
rect 109 1188 113 1194
rect 146 1188 150 1194
rect 159 1190 163 1194
rect 183 1194 187 1198
rect 257 1194 261 1198
rect 167 1188 171 1194
rect 204 1188 208 1194
rect 220 1188 224 1194
rect 241 1188 245 1194
rect 278 1188 282 1194
rect 291 1190 295 1194
rect 315 1194 319 1198
rect 389 1194 393 1198
rect 299 1188 303 1194
rect 336 1188 340 1194
rect 352 1188 356 1194
rect 373 1188 377 1194
rect 410 1188 414 1194
rect 423 1190 427 1194
rect 447 1194 451 1198
rect 517 1201 523 1205
rect 587 1201 591 1205
rect 596 1201 600 1205
rect 646 1201 650 1205
rect 671 1201 675 1205
rect 702 1201 706 1205
rect 431 1188 435 1194
rect 468 1188 472 1194
rect 484 1190 488 1194
rect 587 1193 591 1197
rect 630 1194 634 1198
rect 652 1193 659 1197
rect 702 1194 706 1198
rect 573 1189 577 1193
rect 605 1189 609 1193
rect 623 1189 627 1193
rect 680 1189 684 1193
rect 695 1189 699 1193
rect 723 1189 727 1193
rect 109 1175 113 1179
rect 125 1175 129 1181
rect 159 1181 163 1185
rect 146 1175 150 1179
rect 167 1175 171 1179
rect 183 1175 187 1181
rect 204 1175 208 1179
rect 220 1175 224 1179
rect 241 1175 245 1179
rect 257 1175 261 1181
rect 291 1181 295 1185
rect 278 1175 282 1179
rect 299 1175 303 1179
rect 315 1175 319 1181
rect 336 1175 340 1179
rect 352 1175 356 1179
rect 373 1175 377 1179
rect 389 1175 393 1181
rect 423 1181 427 1185
rect 410 1175 414 1179
rect 431 1175 435 1179
rect 447 1175 451 1181
rect 468 1175 472 1179
rect 484 1175 488 1179
rect 568 1177 572 1181
rect 102 1164 106 1168
rect 139 1162 143 1166
rect 159 1162 163 1166
rect 203 1162 207 1166
rect 234 1164 238 1168
rect 271 1162 275 1166
rect 291 1162 295 1166
rect 335 1162 339 1166
rect 366 1164 370 1168
rect 403 1162 407 1166
rect 423 1162 427 1166
rect 467 1162 471 1166
rect 600 1175 604 1179
rect 620 1178 624 1182
rect 639 1174 643 1178
rect 658 1175 662 1179
rect 677 1175 681 1179
rect 690 1176 694 1180
rect 826 1201 830 1205
rect 848 1201 852 1205
rect 907 1201 911 1205
rect 932 1201 936 1205
rect 963 1201 967 1205
rect 1035 1205 1039 1209
rect 1085 1205 1089 1209
rect 1138 1205 1142 1209
rect 1167 1205 1171 1209
rect 1217 1205 1221 1209
rect 1270 1205 1274 1209
rect 1299 1205 1303 1209
rect 1349 1205 1353 1209
rect 1402 1205 1406 1209
rect 1438 1208 1444 1212
rect 1506 1208 1510 1212
rect 1520 1208 1524 1212
rect 1538 1208 1542 1212
rect 1556 1208 1560 1212
rect 1579 1208 1583 1212
rect 1613 1208 1617 1212
rect 1628 1208 1632 1212
rect 1656 1208 1660 1212
rect 1781 1208 1785 1212
rect 1799 1208 1803 1212
rect 1817 1208 1821 1212
rect 1840 1208 1844 1212
rect 1874 1208 1878 1212
rect 1889 1208 1893 1212
rect 1917 1208 1921 1212
rect 848 1193 852 1197
rect 891 1194 895 1198
rect 913 1193 920 1197
rect 963 1194 967 1198
rect 1058 1194 1062 1198
rect 866 1189 870 1193
rect 884 1189 888 1193
rect 941 1189 945 1193
rect 956 1189 960 1193
rect 984 1189 988 1193
rect 787 1185 791 1189
rect 712 1175 716 1179
rect 720 1176 724 1180
rect 732 1176 736 1180
rect 766 1170 770 1174
rect 806 1176 810 1180
rect 795 1169 799 1173
rect 573 1159 577 1163
rect 505 1155 511 1159
rect 598 1156 602 1160
rect 605 1159 609 1163
rect 623 1159 627 1163
rect 645 1156 649 1160
rect 670 1156 674 1160
rect 680 1159 684 1163
rect 696 1159 700 1163
rect 716 1156 720 1160
rect 723 1159 727 1163
rect 861 1175 865 1179
rect 881 1178 885 1182
rect 900 1174 904 1178
rect 1029 1185 1033 1189
rect 1042 1188 1046 1194
rect 1079 1188 1083 1194
rect 1092 1190 1096 1194
rect 1116 1194 1120 1198
rect 1190 1194 1194 1198
rect 1100 1188 1104 1194
rect 1137 1188 1141 1194
rect 1153 1188 1157 1194
rect 1174 1188 1178 1194
rect 1211 1188 1215 1194
rect 1224 1190 1228 1194
rect 1248 1194 1252 1198
rect 1322 1194 1326 1198
rect 1232 1188 1236 1194
rect 1269 1188 1273 1194
rect 1285 1188 1289 1194
rect 1306 1188 1310 1194
rect 1343 1188 1347 1194
rect 1356 1190 1360 1194
rect 1380 1194 1384 1198
rect 1450 1201 1456 1205
rect 1520 1201 1524 1205
rect 1529 1201 1533 1205
rect 1579 1201 1583 1205
rect 1604 1201 1608 1205
rect 1635 1201 1639 1205
rect 1364 1188 1368 1194
rect 1401 1188 1405 1194
rect 1417 1190 1421 1194
rect 1520 1193 1524 1197
rect 1563 1194 1567 1198
rect 1585 1193 1592 1197
rect 1635 1194 1639 1198
rect 1506 1189 1510 1193
rect 1538 1189 1542 1193
rect 1556 1189 1560 1193
rect 1613 1189 1617 1193
rect 1628 1189 1632 1193
rect 1656 1189 1660 1193
rect 919 1175 923 1179
rect 938 1175 942 1179
rect 951 1176 955 1180
rect 973 1175 977 1179
rect 981 1176 985 1180
rect 993 1176 997 1180
rect 1042 1175 1046 1179
rect 1058 1175 1062 1181
rect 1092 1181 1096 1185
rect 1079 1175 1083 1179
rect 1100 1175 1104 1179
rect 1116 1175 1120 1181
rect 1137 1175 1141 1179
rect 1153 1175 1157 1179
rect 1174 1175 1178 1179
rect 1190 1175 1194 1181
rect 1224 1181 1228 1185
rect 1211 1175 1215 1179
rect 1232 1175 1236 1179
rect 1248 1175 1252 1181
rect 1269 1175 1273 1179
rect 1285 1175 1289 1179
rect 1306 1175 1310 1179
rect 1322 1175 1326 1181
rect 1356 1181 1360 1185
rect 1343 1175 1347 1179
rect 1364 1175 1368 1179
rect 1380 1175 1384 1181
rect 1401 1175 1405 1179
rect 1417 1175 1421 1179
rect 1501 1177 1505 1181
rect 807 1159 811 1163
rect 833 1159 837 1163
rect 102 1148 106 1152
rect 153 1148 157 1152
rect 203 1148 207 1152
rect 234 1148 238 1152
rect 285 1148 289 1152
rect 335 1148 339 1152
rect 366 1148 370 1152
rect 417 1148 421 1152
rect 467 1148 471 1152
rect 541 1149 547 1153
rect 581 1149 585 1153
rect 599 1149 603 1153
rect 630 1149 634 1153
rect 652 1149 656 1153
rect 717 1149 721 1153
rect 859 1156 863 1160
rect 866 1159 870 1163
rect 884 1159 888 1163
rect 906 1156 910 1160
rect 931 1156 935 1160
rect 941 1159 945 1163
rect 957 1159 961 1163
rect 977 1156 981 1160
rect 984 1159 988 1163
rect 1035 1164 1039 1168
rect 1072 1162 1076 1166
rect 1092 1162 1096 1166
rect 1136 1162 1140 1166
rect 1167 1164 1171 1168
rect 1204 1162 1208 1166
rect 1224 1162 1228 1166
rect 1268 1162 1272 1166
rect 1299 1164 1303 1168
rect 1336 1162 1340 1166
rect 1356 1162 1360 1166
rect 1400 1162 1404 1166
rect 1533 1175 1537 1179
rect 1553 1178 1557 1182
rect 1572 1174 1576 1178
rect 1591 1175 1595 1179
rect 1610 1175 1614 1179
rect 1623 1176 1627 1180
rect 1759 1201 1763 1205
rect 1781 1201 1785 1205
rect 1840 1201 1844 1205
rect 1865 1201 1869 1205
rect 1896 1201 1900 1205
rect 1781 1193 1785 1197
rect 1824 1194 1828 1198
rect 1846 1193 1853 1197
rect 1896 1194 1900 1198
rect 1799 1189 1803 1193
rect 1817 1189 1821 1193
rect 1874 1189 1878 1193
rect 1889 1189 1893 1193
rect 1917 1189 1921 1193
rect 1720 1185 1724 1189
rect 1645 1175 1649 1179
rect 1653 1176 1657 1180
rect 1665 1176 1669 1180
rect 1699 1170 1703 1174
rect 1739 1176 1743 1180
rect 1728 1169 1732 1173
rect 1506 1159 1510 1163
rect 1438 1155 1444 1159
rect 1531 1156 1535 1160
rect 1538 1159 1542 1163
rect 1556 1159 1560 1163
rect 1578 1156 1582 1160
rect 1603 1156 1607 1160
rect 1613 1159 1617 1163
rect 1629 1159 1633 1163
rect 1649 1156 1653 1160
rect 1656 1159 1660 1163
rect 1794 1175 1798 1179
rect 1814 1178 1818 1182
rect 1833 1174 1837 1178
rect 1852 1175 1856 1179
rect 1871 1175 1875 1179
rect 1884 1176 1888 1180
rect 1906 1175 1910 1179
rect 1914 1176 1918 1180
rect 1926 1176 1930 1180
rect 1740 1159 1744 1163
rect 1766 1159 1770 1163
rect 777 1149 781 1153
rect 816 1149 820 1153
rect 860 1149 864 1153
rect 891 1149 895 1153
rect 913 1149 917 1153
rect 978 1149 982 1153
rect 1035 1148 1039 1152
rect 1086 1148 1090 1152
rect 1136 1148 1140 1152
rect 1167 1148 1171 1152
rect 1218 1148 1222 1152
rect 1268 1148 1272 1152
rect 1299 1148 1303 1152
rect 1350 1148 1354 1152
rect 1400 1148 1404 1152
rect 1474 1149 1480 1153
rect 1514 1149 1518 1153
rect 1532 1149 1536 1153
rect 1563 1149 1567 1153
rect 1585 1149 1589 1153
rect 1650 1149 1654 1153
rect 1792 1156 1796 1160
rect 1799 1159 1803 1163
rect 1817 1159 1821 1163
rect 1839 1156 1843 1160
rect 1864 1156 1868 1160
rect 1874 1159 1878 1163
rect 1890 1159 1894 1163
rect 1910 1156 1914 1160
rect 1917 1159 1921 1163
rect 1710 1149 1714 1153
rect 1749 1149 1753 1153
rect 1793 1149 1797 1153
rect 1824 1149 1828 1153
rect 1846 1149 1850 1153
rect 1911 1149 1915 1153
rect 96 1141 100 1145
rect 484 1141 488 1145
rect 493 1142 499 1146
rect 572 1142 576 1146
rect 606 1142 610 1146
rect 623 1142 627 1146
rect 679 1142 683 1146
rect 696 1142 700 1146
rect 724 1142 728 1146
rect 807 1142 811 1146
rect 833 1142 837 1146
rect 867 1142 871 1146
rect 884 1142 888 1146
rect 940 1142 944 1146
rect 957 1142 961 1146
rect 985 1142 989 1146
rect 1029 1141 1033 1145
rect 1417 1141 1421 1145
rect 1426 1142 1432 1146
rect 1505 1142 1509 1146
rect 1539 1142 1543 1146
rect 1556 1142 1560 1146
rect 1612 1142 1616 1146
rect 1629 1142 1633 1146
rect 1657 1142 1661 1146
rect 1740 1142 1744 1146
rect 1766 1142 1770 1146
rect 1800 1142 1804 1146
rect 1817 1142 1821 1146
rect 1873 1142 1877 1146
rect 1890 1142 1894 1146
rect 1918 1142 1922 1146
rect 219 1134 224 1138
rect 352 1134 356 1138
rect 529 1135 535 1139
rect 581 1135 585 1139
rect 815 1135 819 1139
rect 1001 1136 1005 1140
rect 1013 1136 1017 1140
rect 1152 1134 1157 1138
rect 1285 1134 1289 1138
rect 1462 1135 1468 1139
rect 1514 1135 1518 1139
rect 1748 1135 1752 1139
rect 1934 1136 1938 1140
rect 1946 1136 1950 1140
rect 227 1127 231 1131
rect 517 1127 523 1131
rect 825 1128 829 1132
rect 990 1128 994 1132
rect 211 1123 215 1127
rect 243 1123 247 1127
rect 1160 1127 1164 1131
rect 1450 1127 1456 1131
rect 1758 1128 1762 1132
rect 1923 1128 1927 1132
rect 1144 1123 1148 1127
rect 1176 1123 1180 1127
rect 211 1116 215 1120
rect 243 1116 247 1120
rect 1144 1116 1148 1120
rect 1176 1116 1180 1120
rect 227 1109 231 1113
rect 484 1109 488 1113
rect 553 1109 559 1113
rect 873 1109 877 1113
rect 909 1109 913 1113
rect 976 1109 980 1113
rect 1160 1109 1164 1113
rect 1417 1109 1421 1113
rect 1486 1109 1492 1113
rect 1806 1109 1810 1113
rect 1842 1109 1846 1113
rect 1909 1109 1913 1113
rect 484 1101 488 1105
rect 493 1102 499 1106
rect 859 1102 863 1106
rect 211 1097 215 1101
rect 243 1097 247 1101
rect 227 1093 231 1097
rect 873 1095 877 1099
rect 923 1095 927 1099
rect 976 1095 980 1099
rect 1417 1101 1421 1105
rect 1426 1102 1432 1106
rect 1792 1102 1796 1106
rect 1144 1097 1148 1101
rect 1176 1097 1180 1101
rect 1160 1093 1164 1097
rect 1806 1095 1810 1099
rect 1856 1095 1860 1099
rect 1909 1095 1913 1099
rect 219 1086 224 1090
rect 353 1086 357 1090
rect 896 1084 900 1088
rect 102 1079 106 1083
rect 138 1079 142 1083
rect 205 1079 209 1083
rect 234 1079 238 1083
rect 270 1079 274 1083
rect 337 1079 341 1083
rect 366 1079 370 1083
rect 402 1079 406 1083
rect 469 1079 473 1083
rect 553 1079 559 1083
rect 493 1072 499 1076
rect 867 1075 871 1079
rect 880 1078 884 1084
rect 917 1078 921 1084
rect 930 1080 934 1084
rect 954 1084 958 1088
rect 1152 1086 1157 1090
rect 1286 1086 1290 1090
rect 1829 1084 1833 1088
rect 938 1078 942 1084
rect 975 1078 979 1084
rect 991 1078 995 1084
rect 1035 1079 1039 1083
rect 1071 1079 1075 1083
rect 1138 1079 1142 1083
rect 1167 1079 1171 1083
rect 1203 1079 1207 1083
rect 1270 1079 1274 1083
rect 1299 1079 1303 1083
rect 1335 1079 1339 1083
rect 1402 1079 1406 1083
rect 1486 1079 1492 1083
rect 102 1065 106 1069
rect 152 1065 156 1069
rect 205 1065 209 1069
rect 234 1065 238 1069
rect 284 1065 288 1069
rect 337 1065 341 1069
rect 366 1065 370 1069
rect 416 1065 420 1069
rect 469 1065 473 1069
rect 880 1065 884 1069
rect 896 1065 900 1071
rect 930 1071 934 1075
rect 917 1065 921 1069
rect 125 1054 129 1058
rect 96 1045 100 1049
rect 109 1048 113 1054
rect 146 1048 150 1054
rect 159 1050 163 1054
rect 183 1054 187 1058
rect 257 1054 261 1058
rect 167 1048 171 1054
rect 204 1048 208 1054
rect 220 1048 224 1054
rect 241 1048 245 1054
rect 278 1048 282 1054
rect 291 1050 295 1054
rect 315 1054 319 1058
rect 389 1054 393 1058
rect 299 1048 303 1054
rect 336 1048 340 1054
rect 352 1048 356 1054
rect 373 1048 377 1054
rect 410 1048 414 1054
rect 423 1050 427 1054
rect 447 1054 451 1058
rect 431 1048 435 1054
rect 468 1048 472 1054
rect 484 1050 488 1054
rect 938 1065 942 1069
rect 954 1065 958 1071
rect 1426 1072 1432 1076
rect 1800 1075 1804 1079
rect 1813 1078 1817 1084
rect 1850 1078 1854 1084
rect 1863 1080 1867 1084
rect 1887 1084 1891 1088
rect 1871 1078 1875 1084
rect 1908 1078 1912 1084
rect 1924 1078 1928 1084
rect 975 1065 979 1069
rect 991 1065 995 1069
rect 1035 1065 1039 1069
rect 1085 1065 1089 1069
rect 1138 1065 1142 1069
rect 1167 1065 1171 1069
rect 1217 1065 1221 1069
rect 1270 1065 1274 1069
rect 1299 1065 1303 1069
rect 1349 1065 1353 1069
rect 1402 1065 1406 1069
rect 1813 1065 1817 1069
rect 1829 1065 1833 1071
rect 1863 1071 1867 1075
rect 1850 1065 1854 1069
rect 873 1054 877 1058
rect 910 1052 914 1056
rect 930 1052 934 1056
rect 974 1052 978 1056
rect 1058 1054 1062 1058
rect 109 1035 113 1039
rect 125 1035 129 1041
rect 159 1041 163 1045
rect 146 1035 150 1039
rect 167 1035 171 1039
rect 183 1035 187 1041
rect 204 1035 208 1039
rect 220 1035 224 1039
rect 241 1035 245 1039
rect 257 1035 261 1041
rect 291 1041 295 1045
rect 278 1035 282 1039
rect 299 1035 303 1039
rect 315 1035 319 1041
rect 336 1035 340 1039
rect 352 1035 356 1039
rect 373 1035 377 1039
rect 389 1035 393 1041
rect 423 1041 427 1045
rect 410 1035 414 1039
rect 431 1035 435 1039
rect 447 1035 451 1041
rect 505 1045 511 1049
rect 1029 1045 1033 1049
rect 1042 1048 1046 1054
rect 1079 1048 1083 1054
rect 1092 1050 1096 1054
rect 1116 1054 1120 1058
rect 1190 1054 1194 1058
rect 1100 1048 1104 1054
rect 1137 1048 1141 1054
rect 1153 1048 1157 1054
rect 1174 1048 1178 1054
rect 1211 1048 1215 1054
rect 1224 1050 1228 1054
rect 1248 1054 1252 1058
rect 1322 1054 1326 1058
rect 1232 1048 1236 1054
rect 1269 1048 1273 1054
rect 1285 1048 1289 1054
rect 1306 1048 1310 1054
rect 1343 1048 1347 1054
rect 1356 1050 1360 1054
rect 1380 1054 1384 1058
rect 1364 1048 1368 1054
rect 1401 1048 1405 1054
rect 1417 1050 1421 1054
rect 1871 1065 1875 1069
rect 1887 1065 1891 1071
rect 1908 1065 1912 1069
rect 1924 1065 1928 1069
rect 1806 1054 1810 1058
rect 1843 1052 1847 1056
rect 1863 1052 1867 1056
rect 1907 1052 1911 1056
rect 468 1035 472 1039
rect 484 1035 488 1039
rect 541 1038 547 1042
rect 873 1038 877 1042
rect 924 1038 928 1042
rect 974 1038 978 1042
rect 1042 1035 1046 1039
rect 1058 1035 1062 1041
rect 1092 1041 1096 1045
rect 1079 1035 1083 1039
rect 102 1024 106 1028
rect 139 1022 143 1026
rect 159 1022 163 1026
rect 203 1022 207 1026
rect 234 1024 238 1028
rect 271 1022 275 1026
rect 291 1022 295 1026
rect 335 1022 339 1026
rect 366 1024 370 1028
rect 403 1022 407 1026
rect 423 1022 427 1026
rect 467 1022 471 1026
rect 866 1030 870 1034
rect 991 1031 995 1035
rect 1100 1035 1104 1039
rect 1116 1035 1120 1041
rect 1137 1035 1141 1039
rect 1153 1035 1157 1039
rect 1174 1035 1178 1039
rect 1190 1035 1194 1041
rect 1224 1041 1228 1045
rect 1211 1035 1215 1039
rect 1232 1035 1236 1039
rect 1248 1035 1252 1041
rect 1269 1035 1273 1039
rect 1285 1035 1289 1039
rect 1306 1035 1310 1039
rect 1322 1035 1326 1041
rect 1356 1041 1360 1045
rect 1343 1035 1347 1039
rect 1364 1035 1368 1039
rect 1380 1035 1384 1041
rect 1438 1045 1444 1049
rect 1401 1035 1405 1039
rect 1417 1035 1421 1039
rect 1474 1038 1480 1042
rect 1806 1038 1810 1042
rect 1857 1038 1861 1042
rect 1907 1038 1911 1042
rect 553 1023 559 1027
rect 873 1023 877 1027
rect 909 1023 913 1027
rect 976 1023 980 1027
rect 505 1015 511 1019
rect 859 1016 863 1020
rect 1035 1024 1039 1028
rect 1072 1022 1076 1026
rect 1092 1022 1096 1026
rect 1136 1022 1140 1026
rect 1167 1024 1171 1028
rect 1204 1022 1208 1026
rect 1224 1022 1228 1026
rect 1268 1022 1272 1026
rect 1299 1024 1303 1028
rect 1336 1022 1340 1026
rect 1356 1022 1360 1026
rect 1400 1022 1404 1026
rect 1799 1030 1803 1034
rect 1924 1031 1928 1035
rect 1486 1023 1492 1027
rect 1806 1023 1810 1027
rect 1842 1023 1846 1027
rect 1909 1023 1913 1027
rect 102 1008 106 1012
rect 153 1008 157 1012
rect 203 1008 207 1012
rect 234 1008 238 1012
rect 285 1008 289 1012
rect 335 1008 339 1012
rect 366 1008 370 1012
rect 417 1008 421 1012
rect 467 1008 471 1012
rect 541 1008 547 1012
rect 873 1009 877 1013
rect 923 1009 927 1013
rect 976 1009 980 1013
rect 1438 1015 1444 1019
rect 1792 1016 1796 1020
rect 1035 1008 1039 1012
rect 1086 1008 1090 1012
rect 1136 1008 1140 1012
rect 1167 1008 1171 1012
rect 1218 1008 1222 1012
rect 1268 1008 1272 1012
rect 1299 1008 1303 1012
rect 1350 1008 1354 1012
rect 1400 1008 1404 1012
rect 1474 1008 1480 1012
rect 1806 1009 1810 1013
rect 1856 1009 1860 1013
rect 1909 1009 1913 1013
rect 95 1001 99 1005
rect 484 1001 488 1005
rect 896 998 900 1002
rect 102 993 106 997
rect 138 993 142 997
rect 205 993 209 997
rect 234 993 238 997
rect 270 993 274 997
rect 337 993 341 997
rect 366 993 370 997
rect 402 993 406 997
rect 469 993 473 997
rect 553 993 559 997
rect 493 986 499 990
rect 867 989 871 993
rect 880 992 884 998
rect 917 992 921 998
rect 930 994 934 998
rect 954 998 958 1002
rect 1028 1001 1032 1005
rect 1417 1001 1421 1005
rect 1829 998 1833 1002
rect 938 992 942 998
rect 975 992 979 998
rect 991 994 995 998
rect 1013 992 1017 996
rect 1035 993 1039 997
rect 1071 993 1075 997
rect 1138 993 1142 997
rect 1167 993 1171 997
rect 1203 993 1207 997
rect 1270 993 1274 997
rect 1299 993 1303 997
rect 1335 993 1339 997
rect 1402 993 1406 997
rect 1486 993 1492 997
rect 102 979 106 983
rect 152 979 156 983
rect 205 979 209 983
rect 234 979 238 983
rect 284 979 288 983
rect 337 979 341 983
rect 366 979 370 983
rect 416 979 420 983
rect 469 979 473 983
rect 880 979 884 983
rect 896 979 900 985
rect 930 985 934 989
rect 917 979 921 983
rect 125 968 129 972
rect 96 959 100 963
rect 109 962 113 968
rect 146 962 150 968
rect 159 964 163 968
rect 183 968 187 972
rect 257 968 261 972
rect 167 962 171 968
rect 204 962 208 968
rect 220 962 224 968
rect 241 962 245 968
rect 278 962 282 968
rect 291 964 295 968
rect 315 968 319 972
rect 389 968 393 972
rect 299 962 303 968
rect 336 962 340 968
rect 352 962 356 968
rect 373 962 377 968
rect 410 962 414 968
rect 423 964 427 968
rect 447 968 451 972
rect 431 962 435 968
rect 468 962 472 968
rect 484 964 488 968
rect 938 979 942 983
rect 954 979 958 985
rect 975 979 979 983
rect 991 979 995 988
rect 1426 986 1432 990
rect 1800 989 1804 993
rect 1813 992 1817 998
rect 1850 992 1854 998
rect 1863 994 1867 998
rect 1887 998 1891 1002
rect 1871 992 1875 998
rect 1908 992 1912 998
rect 1924 994 1928 998
rect 1946 992 1950 996
rect 1013 976 1017 980
rect 1035 979 1039 983
rect 1085 979 1089 983
rect 1138 979 1142 983
rect 1167 979 1171 983
rect 1217 979 1221 983
rect 1270 979 1274 983
rect 1299 979 1303 983
rect 1349 979 1353 983
rect 1402 979 1406 983
rect 1813 979 1817 983
rect 1829 979 1833 985
rect 1863 985 1867 989
rect 1850 979 1854 983
rect 873 968 877 972
rect 910 966 914 970
rect 930 966 934 970
rect 974 966 978 970
rect 1058 968 1062 972
rect 109 949 113 953
rect 125 949 129 955
rect 159 955 163 959
rect 146 949 150 953
rect 167 949 171 953
rect 183 949 187 955
rect 204 949 208 953
rect 220 949 224 953
rect 241 949 245 953
rect 257 949 261 955
rect 291 955 295 959
rect 278 949 282 953
rect 299 949 303 953
rect 315 949 319 955
rect 336 949 340 953
rect 352 949 356 953
rect 373 949 377 953
rect 389 949 393 955
rect 423 955 427 959
rect 410 949 414 953
rect 431 949 435 953
rect 447 949 451 955
rect 505 959 511 963
rect 1029 959 1033 963
rect 1042 962 1046 968
rect 1079 962 1083 968
rect 1092 964 1096 968
rect 1116 968 1120 972
rect 1190 968 1194 972
rect 1100 962 1104 968
rect 1137 962 1141 968
rect 1153 962 1157 968
rect 1174 962 1178 968
rect 1211 962 1215 968
rect 1224 964 1228 968
rect 1248 968 1252 972
rect 1322 968 1326 972
rect 1232 962 1236 968
rect 1269 962 1273 968
rect 1285 962 1289 968
rect 1306 962 1310 968
rect 1343 962 1347 968
rect 1356 964 1360 968
rect 1380 968 1384 972
rect 1364 962 1368 968
rect 1401 962 1405 968
rect 1417 964 1421 968
rect 1871 979 1875 983
rect 1887 979 1891 985
rect 1908 979 1912 983
rect 1924 979 1928 988
rect 1946 976 1950 980
rect 1806 968 1810 972
rect 1843 966 1847 970
rect 1863 966 1867 970
rect 1907 966 1911 970
rect 468 949 472 953
rect 484 949 488 953
rect 541 952 547 956
rect 873 952 877 956
rect 924 952 928 956
rect 974 952 978 956
rect 1042 949 1046 953
rect 1058 949 1062 955
rect 1092 955 1096 959
rect 1079 949 1083 953
rect 1100 949 1104 953
rect 1116 949 1120 955
rect 1137 949 1141 953
rect 1153 949 1157 953
rect 1174 949 1178 953
rect 1190 949 1194 955
rect 1224 955 1228 959
rect 1211 949 1215 953
rect 1232 949 1236 953
rect 1248 949 1252 955
rect 1269 949 1273 953
rect 1285 949 1289 953
rect 1306 949 1310 953
rect 1322 949 1326 955
rect 1356 955 1360 959
rect 1343 949 1347 953
rect 1364 949 1368 953
rect 1380 949 1384 955
rect 1438 959 1444 963
rect 1401 949 1405 953
rect 1417 949 1421 953
rect 1474 952 1480 956
rect 1806 952 1810 956
rect 1857 952 1861 956
rect 1907 952 1911 956
rect 102 938 106 942
rect 139 936 143 940
rect 159 936 163 940
rect 203 936 207 940
rect 234 938 238 942
rect 271 936 275 940
rect 291 936 295 940
rect 335 936 339 940
rect 366 938 370 942
rect 403 936 407 940
rect 423 936 427 940
rect 467 936 471 940
rect 1035 938 1039 942
rect 1072 936 1076 940
rect 1092 936 1096 940
rect 1136 936 1140 940
rect 1167 938 1171 942
rect 1204 936 1208 940
rect 1224 936 1228 940
rect 1268 936 1272 940
rect 1299 938 1303 942
rect 1336 936 1340 940
rect 1356 936 1360 940
rect 1400 936 1404 940
rect 505 929 511 933
rect 1438 929 1444 933
rect 102 922 106 926
rect 153 922 157 926
rect 203 922 207 926
rect 234 922 238 926
rect 285 922 289 926
rect 335 922 339 926
rect 366 922 370 926
rect 417 922 421 926
rect 467 922 471 926
rect 541 922 547 926
rect 1035 922 1039 926
rect 1086 922 1090 926
rect 1136 922 1140 926
rect 1167 922 1171 926
rect 1218 922 1222 926
rect 1268 922 1272 926
rect 1299 922 1303 926
rect 1350 922 1354 926
rect 1400 922 1404 926
rect 1474 922 1480 926
rect 95 915 99 919
rect 484 915 488 919
rect 1028 915 1032 919
rect 1417 915 1421 919
rect 220 908 224 912
rect 328 908 332 912
rect 352 908 356 912
rect 1153 908 1157 912
rect 1261 908 1265 912
rect 1285 908 1289 912
rect 344 901 348 905
rect 328 897 332 901
rect 360 897 364 901
rect 1277 901 1281 905
rect 1261 897 1265 901
rect 1293 897 1297 901
rect 328 890 332 894
rect 360 890 364 894
rect 1013 890 1017 894
rect 1261 890 1265 894
rect 1293 890 1297 894
rect 1946 890 1950 894
rect 344 883 348 887
rect 484 883 488 887
rect 1277 883 1281 887
rect 1417 883 1421 887
rect 484 875 488 879
rect 1417 875 1421 879
rect 328 871 332 875
rect 360 871 364 875
rect 344 867 348 871
rect 1261 871 1265 875
rect 1293 871 1297 875
rect 1277 867 1281 871
rect 220 860 224 864
rect 328 860 332 864
rect 352 860 356 864
rect 1153 860 1157 864
rect 1261 860 1265 864
rect 1285 860 1289 864
rect 102 853 106 857
rect 138 853 142 857
rect 205 853 209 857
rect 234 853 238 857
rect 270 853 274 857
rect 337 853 341 857
rect 366 853 370 857
rect 402 853 406 857
rect 469 853 473 857
rect 553 853 559 857
rect 1035 853 1039 857
rect 1071 853 1075 857
rect 1138 853 1142 857
rect 1167 853 1171 857
rect 1203 853 1207 857
rect 1270 853 1274 857
rect 1299 853 1303 857
rect 1335 853 1339 857
rect 1402 853 1406 857
rect 1486 853 1492 857
rect 493 846 499 850
rect 1426 846 1432 850
rect 102 839 106 843
rect 152 839 156 843
rect 205 839 209 843
rect 234 839 238 843
rect 284 839 288 843
rect 337 839 341 843
rect 366 839 370 843
rect 416 839 420 843
rect 469 839 473 843
rect 1035 839 1039 843
rect 1085 839 1089 843
rect 1138 839 1142 843
rect 1167 839 1171 843
rect 1217 839 1221 843
rect 1270 839 1274 843
rect 1299 839 1303 843
rect 1349 839 1353 843
rect 1402 839 1406 843
rect 125 828 129 832
rect 96 819 100 823
rect 109 822 113 828
rect 146 822 150 828
rect 159 824 163 828
rect 183 828 187 832
rect 257 828 261 832
rect 167 822 171 828
rect 204 822 208 828
rect 220 822 224 828
rect 241 822 245 828
rect 278 822 282 828
rect 291 824 295 828
rect 315 828 319 832
rect 389 828 393 832
rect 299 822 303 828
rect 336 822 340 828
rect 352 822 356 828
rect 373 822 377 828
rect 410 822 414 828
rect 423 824 427 828
rect 447 828 451 832
rect 1058 828 1062 832
rect 431 822 435 828
rect 468 822 472 828
rect 484 824 488 828
rect 109 809 113 813
rect 125 809 129 815
rect 159 815 163 819
rect 146 809 150 813
rect 167 809 171 813
rect 183 809 187 815
rect 204 809 208 813
rect 220 809 224 813
rect 241 809 245 813
rect 257 809 261 815
rect 291 815 295 819
rect 278 809 282 813
rect 299 809 303 813
rect 315 809 319 815
rect 336 809 340 813
rect 352 809 356 813
rect 373 809 377 813
rect 389 809 393 815
rect 423 815 427 819
rect 410 809 414 813
rect 431 809 435 813
rect 447 809 451 815
rect 1029 819 1033 823
rect 1042 822 1046 828
rect 1079 822 1083 828
rect 1092 824 1096 828
rect 1116 828 1120 832
rect 1190 828 1194 832
rect 1100 822 1104 828
rect 1137 822 1141 828
rect 1153 822 1157 828
rect 1174 822 1178 828
rect 1211 822 1215 828
rect 1224 824 1228 828
rect 1248 828 1252 832
rect 1322 828 1326 832
rect 1232 822 1236 828
rect 1269 822 1273 828
rect 1285 822 1289 828
rect 1306 822 1310 828
rect 1343 822 1347 828
rect 1356 824 1360 828
rect 1380 828 1384 832
rect 1364 822 1368 828
rect 1401 822 1405 828
rect 1417 824 1421 828
rect 468 809 472 813
rect 484 809 488 813
rect 1042 809 1046 813
rect 1058 809 1062 815
rect 1092 815 1096 819
rect 1079 809 1083 813
rect 1100 809 1104 813
rect 1116 809 1120 815
rect 1137 809 1141 813
rect 1153 809 1157 813
rect 1174 809 1178 813
rect 1190 809 1194 815
rect 1224 815 1228 819
rect 1211 809 1215 813
rect 1232 809 1236 813
rect 1248 809 1252 815
rect 1269 809 1273 813
rect 1285 809 1289 813
rect 1306 809 1310 813
rect 1322 809 1326 815
rect 1356 815 1360 819
rect 1343 809 1347 813
rect 1364 809 1368 813
rect 1380 809 1384 815
rect 1401 809 1405 813
rect 1417 809 1421 813
rect 102 798 106 802
rect 139 796 143 800
rect 159 796 163 800
rect 203 796 207 800
rect 234 798 238 802
rect 271 796 275 800
rect 291 796 295 800
rect 335 796 339 800
rect 366 798 370 802
rect 403 796 407 800
rect 423 796 427 800
rect 467 796 471 800
rect 1035 798 1039 802
rect 1072 796 1076 800
rect 1092 796 1096 800
rect 1136 796 1140 800
rect 1167 798 1171 802
rect 1204 796 1208 800
rect 1224 796 1228 800
rect 1268 796 1272 800
rect 1299 798 1303 802
rect 1336 796 1340 800
rect 1356 796 1360 800
rect 1400 796 1404 800
rect 505 789 511 793
rect 1438 789 1444 793
rect 102 782 106 786
rect 153 782 157 786
rect 203 782 207 786
rect 234 782 238 786
rect 285 782 289 786
rect 335 782 339 786
rect 366 782 370 786
rect 417 782 421 786
rect 467 782 471 786
rect 541 782 547 786
rect 1035 782 1039 786
rect 1086 782 1090 786
rect 1136 782 1140 786
rect 1167 782 1171 786
rect 1218 782 1222 786
rect 1268 782 1272 786
rect 1299 782 1303 786
rect 1350 782 1354 786
rect 1400 782 1404 786
rect 1474 782 1480 786
rect 553 774 559 778
rect 574 774 578 778
rect 610 774 614 778
rect 677 774 681 778
rect 706 774 710 778
rect 742 774 746 778
rect 809 774 813 778
rect 838 774 842 778
rect 874 774 878 778
rect 941 774 945 778
rect 970 774 974 778
rect 1006 774 1010 778
rect 1073 774 1077 778
rect 1486 774 1492 778
rect 1507 774 1511 778
rect 1543 774 1547 778
rect 1610 774 1614 778
rect 1639 774 1643 778
rect 1675 774 1679 778
rect 1742 774 1746 778
rect 1771 774 1775 778
rect 1807 774 1811 778
rect 1874 774 1878 778
rect 1903 774 1907 778
rect 1939 774 1943 778
rect 2006 774 2010 778
rect 493 767 499 771
rect 1426 767 1432 771
rect 574 760 578 764
rect 624 760 628 764
rect 677 760 681 764
rect 706 760 710 764
rect 756 760 760 764
rect 809 760 813 764
rect 838 760 842 764
rect 888 760 892 764
rect 941 760 945 764
rect 970 760 974 764
rect 1020 760 1024 764
rect 1073 760 1077 764
rect 1507 760 1511 764
rect 1557 760 1561 764
rect 1610 760 1614 764
rect 1639 760 1643 764
rect 1689 760 1693 764
rect 1742 760 1746 764
rect 1771 760 1775 764
rect 1821 760 1825 764
rect 1874 760 1878 764
rect 1903 760 1907 764
rect 1953 760 1957 764
rect 2006 760 2010 764
rect 597 749 601 753
rect 234 741 238 745
rect 270 741 274 745
rect 337 741 341 745
rect 553 741 559 745
rect 568 740 572 744
rect 581 743 585 749
rect 618 743 622 749
rect 631 745 635 749
rect 655 749 659 753
rect 729 749 733 753
rect 639 743 643 749
rect 676 743 680 749
rect 692 745 696 749
rect 493 734 499 738
rect 234 727 238 731
rect 284 727 288 731
rect 337 727 341 731
rect 581 730 585 734
rect 597 730 601 736
rect 631 736 635 740
rect 618 730 622 734
rect 639 730 643 734
rect 655 730 659 736
rect 700 740 704 744
rect 713 743 717 749
rect 750 743 754 749
rect 763 745 767 749
rect 787 749 791 753
rect 861 749 865 753
rect 771 743 775 749
rect 808 743 812 749
rect 824 745 828 749
rect 676 730 680 734
rect 692 730 696 734
rect 713 730 717 734
rect 729 730 733 736
rect 763 736 767 740
rect 750 730 754 734
rect 771 730 775 734
rect 787 730 791 736
rect 832 740 836 744
rect 845 743 849 749
rect 882 743 886 749
rect 895 745 899 749
rect 919 749 923 753
rect 993 749 997 753
rect 903 743 907 749
rect 940 743 944 749
rect 956 745 960 749
rect 808 730 812 734
rect 824 730 828 734
rect 845 730 849 734
rect 861 730 865 736
rect 895 736 899 740
rect 882 730 886 734
rect 903 730 907 734
rect 919 730 923 736
rect 964 740 968 744
rect 977 743 981 749
rect 1014 743 1018 749
rect 1027 745 1031 749
rect 1051 749 1055 753
rect 1530 749 1534 753
rect 1035 743 1039 749
rect 1072 743 1076 749
rect 1088 745 1092 749
rect 1167 741 1171 745
rect 1203 741 1207 745
rect 1270 741 1274 745
rect 1486 741 1492 745
rect 940 730 944 734
rect 956 730 960 734
rect 977 730 981 734
rect 993 730 997 736
rect 1027 736 1031 740
rect 1014 730 1018 734
rect 257 716 261 720
rect 219 707 223 711
rect 241 710 245 716
rect 278 710 282 716
rect 291 712 295 716
rect 315 716 319 720
rect 299 710 303 716
rect 336 710 340 716
rect 352 710 356 716
rect 574 719 578 723
rect 611 717 615 721
rect 631 717 635 721
rect 675 717 679 721
rect 706 719 710 723
rect 743 717 747 721
rect 763 717 767 721
rect 807 717 811 721
rect 838 719 842 723
rect 875 717 879 721
rect 895 717 899 721
rect 939 717 943 721
rect 956 722 960 726
rect 1035 730 1039 734
rect 1051 730 1055 736
rect 1501 740 1505 744
rect 1514 743 1518 749
rect 1551 743 1555 749
rect 1564 745 1568 749
rect 1588 749 1592 753
rect 1662 749 1666 753
rect 1572 743 1576 749
rect 1609 743 1613 749
rect 1625 745 1629 749
rect 1426 734 1432 738
rect 1072 730 1076 734
rect 1088 730 1092 734
rect 970 719 974 723
rect 1007 717 1011 721
rect 1027 717 1031 721
rect 1071 717 1075 721
rect 1088 722 1092 726
rect 1167 727 1171 731
rect 1217 727 1221 731
rect 1270 727 1274 731
rect 1514 730 1518 734
rect 1530 730 1534 736
rect 1564 736 1568 740
rect 1551 730 1555 734
rect 1572 730 1576 734
rect 1588 730 1592 736
rect 1633 740 1637 744
rect 1646 743 1650 749
rect 1683 743 1687 749
rect 1696 745 1700 749
rect 1720 749 1724 753
rect 1794 749 1798 753
rect 1704 743 1708 749
rect 1741 743 1745 749
rect 1757 745 1761 749
rect 1609 730 1613 734
rect 1625 730 1629 734
rect 1646 730 1650 734
rect 1662 730 1666 736
rect 1696 736 1700 740
rect 1683 730 1687 734
rect 1704 730 1708 734
rect 1720 730 1724 736
rect 1765 740 1769 744
rect 1778 743 1782 749
rect 1815 743 1819 749
rect 1828 745 1832 749
rect 1852 749 1856 753
rect 1926 749 1930 753
rect 1836 743 1840 749
rect 1873 743 1877 749
rect 1889 745 1893 749
rect 1741 730 1745 734
rect 1757 730 1761 734
rect 1778 730 1782 734
rect 1794 730 1798 736
rect 1828 736 1832 740
rect 1815 730 1819 734
rect 1836 730 1840 734
rect 1852 730 1856 736
rect 1897 740 1901 744
rect 1910 743 1914 749
rect 1947 743 1951 749
rect 1960 745 1964 749
rect 1984 749 1988 753
rect 1968 743 1972 749
rect 2005 743 2009 749
rect 2021 745 2025 749
rect 1873 730 1877 734
rect 1889 730 1893 734
rect 1910 730 1914 734
rect 1926 730 1930 736
rect 1960 736 1964 740
rect 1947 730 1951 734
rect 1190 716 1194 720
rect 505 710 511 714
rect 241 697 245 701
rect 257 697 261 703
rect 291 703 295 707
rect 278 697 282 701
rect 299 697 303 701
rect 315 697 319 703
rect 1152 707 1156 711
rect 1174 710 1178 716
rect 1211 710 1215 716
rect 1224 712 1228 716
rect 1248 716 1252 720
rect 1232 710 1236 716
rect 1269 710 1273 716
rect 1285 710 1289 716
rect 1507 719 1511 723
rect 1544 717 1548 721
rect 1564 717 1568 721
rect 1608 717 1612 721
rect 1639 719 1643 723
rect 1676 717 1680 721
rect 1696 717 1700 721
rect 1740 717 1744 721
rect 1771 719 1775 723
rect 1808 717 1812 721
rect 1828 717 1832 721
rect 1872 717 1876 721
rect 1889 722 1893 726
rect 1968 730 1972 734
rect 1984 730 1988 736
rect 2005 730 2009 734
rect 2021 730 2025 734
rect 1903 719 1907 723
rect 1940 717 1944 721
rect 1960 717 1964 721
rect 2004 717 2008 721
rect 2021 722 2025 726
rect 1438 710 1444 714
rect 541 703 547 707
rect 574 703 578 707
rect 625 703 629 707
rect 675 703 679 707
rect 706 703 710 707
rect 757 703 761 707
rect 807 703 811 707
rect 838 703 842 707
rect 889 703 893 707
rect 939 703 943 707
rect 970 703 974 707
rect 1021 703 1025 707
rect 1071 703 1075 707
rect 336 697 340 701
rect 352 697 356 701
rect 1174 697 1178 701
rect 1190 697 1194 703
rect 1224 703 1228 707
rect 1211 697 1215 701
rect 234 686 238 690
rect 271 684 275 688
rect 291 684 295 688
rect 335 684 339 688
rect 493 690 499 694
rect 572 690 576 694
rect 606 690 610 694
rect 623 690 627 694
rect 679 690 683 694
rect 696 690 700 694
rect 724 690 728 694
rect 1232 697 1236 701
rect 1248 697 1252 703
rect 1474 703 1480 707
rect 1507 703 1511 707
rect 1558 703 1562 707
rect 1608 703 1612 707
rect 1639 703 1643 707
rect 1690 703 1694 707
rect 1740 703 1744 707
rect 1771 703 1775 707
rect 1822 703 1826 707
rect 1872 703 1876 707
rect 1903 703 1907 707
rect 1954 703 1958 707
rect 2004 703 2008 707
rect 1269 697 1273 701
rect 1285 697 1289 701
rect 529 683 535 687
rect 599 683 603 687
rect 630 683 634 687
rect 652 683 656 687
rect 717 683 721 687
rect 505 677 511 681
rect 234 670 238 674
rect 285 670 289 674
rect 335 670 339 674
rect 541 670 547 674
rect 573 673 577 677
rect 598 676 602 680
rect 605 673 609 677
rect 623 673 627 677
rect 645 676 649 680
rect 670 676 674 680
rect 680 673 684 677
rect 696 673 700 677
rect 716 676 720 680
rect 723 673 727 677
rect 787 683 791 687
rect 352 663 356 667
rect 219 654 223 658
rect 344 656 348 660
rect 368 656 372 660
rect 227 647 231 651
rect 368 647 372 651
rect 600 657 604 661
rect 620 654 624 658
rect 639 658 643 662
rect 741 669 745 673
rect 756 669 760 673
rect 658 657 662 661
rect 677 657 681 661
rect 690 656 694 660
rect 712 657 716 661
rect 720 656 724 660
rect 732 656 736 660
rect 573 643 577 647
rect 605 643 609 647
rect 623 643 627 647
rect 680 643 684 647
rect 695 643 699 647
rect 723 643 727 647
rect 234 639 238 643
rect 301 639 305 643
rect 337 639 341 643
rect 553 639 559 643
rect 587 639 591 643
rect 630 638 634 642
rect 652 639 659 643
rect 702 638 706 642
rect 493 632 499 636
rect 234 625 238 629
rect 287 625 291 629
rect 337 625 341 629
rect 517 631 523 635
rect 587 631 591 635
rect 646 631 650 635
rect 671 631 675 635
rect 702 631 706 635
rect 795 661 799 669
rect 868 683 872 687
rect 822 669 826 673
rect 837 669 841 673
rect 1167 686 1171 690
rect 1204 684 1208 688
rect 1224 684 1228 688
rect 1268 684 1272 688
rect 1426 690 1432 694
rect 1505 690 1509 694
rect 1539 690 1543 694
rect 1556 690 1560 694
rect 1612 690 1616 694
rect 1629 690 1633 694
rect 1657 690 1661 694
rect 1462 683 1468 687
rect 1532 683 1536 687
rect 1563 683 1567 687
rect 1585 683 1589 687
rect 1650 683 1654 687
rect 818 661 822 665
rect 764 655 768 659
rect 777 647 781 651
rect 876 661 880 669
rect 1438 677 1444 681
rect 1167 670 1171 674
rect 1218 670 1222 674
rect 1268 670 1272 674
rect 1474 670 1480 674
rect 1506 673 1510 677
rect 1531 676 1535 680
rect 1538 673 1542 677
rect 1556 673 1560 677
rect 1578 676 1582 680
rect 1603 676 1607 680
rect 1613 673 1617 677
rect 1629 673 1633 677
rect 1649 676 1653 680
rect 1656 673 1660 677
rect 1720 683 1724 687
rect 903 661 907 665
rect 1285 663 1289 667
rect 845 655 849 659
rect 1152 654 1156 658
rect 1277 656 1281 660
rect 1301 656 1305 660
rect 858 647 862 651
rect 1160 647 1164 651
rect 1301 647 1305 651
rect 1533 657 1537 661
rect 1553 654 1557 658
rect 1572 658 1576 662
rect 1674 669 1678 673
rect 1689 669 1693 673
rect 1591 657 1595 661
rect 1610 657 1614 661
rect 1623 656 1627 660
rect 1645 657 1649 661
rect 1653 656 1657 660
rect 1665 656 1669 660
rect 1506 643 1510 647
rect 1538 643 1542 647
rect 1556 643 1560 647
rect 1613 643 1617 647
rect 1628 643 1632 647
rect 1656 643 1660 647
rect 1167 639 1171 643
rect 1234 639 1238 643
rect 1270 639 1274 643
rect 1486 639 1492 643
rect 1520 639 1524 643
rect 1563 638 1567 642
rect 1585 639 1592 643
rect 1635 638 1639 642
rect 1426 632 1432 636
rect 505 624 511 628
rect 573 624 577 628
rect 587 624 591 628
rect 605 624 609 628
rect 623 624 627 628
rect 646 624 650 628
rect 680 624 684 628
rect 695 624 699 628
rect 723 624 727 628
rect 256 614 260 618
rect 219 608 223 614
rect 235 608 239 614
rect 272 608 276 614
rect 280 610 284 614
rect 314 614 318 618
rect 517 617 523 621
rect 587 617 591 621
rect 646 617 650 621
rect 671 617 675 621
rect 702 617 706 621
rect 293 608 297 614
rect 330 608 334 614
rect 587 609 591 613
rect 630 610 634 614
rect 652 609 659 613
rect 702 610 706 614
rect 352 605 356 609
rect 573 605 577 609
rect 605 605 609 609
rect 623 605 627 609
rect 680 605 684 609
rect 695 605 699 609
rect 723 605 727 609
rect 219 595 223 599
rect 235 595 239 599
rect 280 601 284 605
rect 256 595 260 601
rect 272 595 276 599
rect 293 595 297 599
rect 314 595 318 601
rect 330 595 334 599
rect 568 593 572 597
rect 236 582 240 586
rect 280 582 284 586
rect 300 582 304 586
rect 337 584 341 588
rect 600 591 604 595
rect 620 594 624 598
rect 639 590 643 594
rect 658 591 662 595
rect 677 591 681 595
rect 690 592 694 596
rect 787 607 791 611
rect 1167 625 1171 629
rect 1220 625 1224 629
rect 1270 625 1274 629
rect 1450 631 1456 635
rect 1520 631 1524 635
rect 1579 631 1583 635
rect 1604 631 1608 635
rect 1635 631 1639 635
rect 1728 661 1732 669
rect 1801 683 1805 687
rect 1755 669 1759 673
rect 1770 669 1774 673
rect 1751 661 1755 665
rect 1697 655 1701 659
rect 1710 647 1714 651
rect 1809 661 1813 669
rect 1836 661 1840 665
rect 1778 655 1782 659
rect 1791 647 1795 651
rect 1438 624 1444 628
rect 1506 624 1510 628
rect 1520 624 1524 628
rect 1538 624 1542 628
rect 1556 624 1560 628
rect 1579 624 1583 628
rect 1613 624 1617 628
rect 1628 624 1632 628
rect 1656 624 1660 628
rect 1189 614 1193 618
rect 868 607 872 611
rect 1152 608 1156 614
rect 1168 608 1172 614
rect 1205 608 1209 614
rect 1213 610 1217 614
rect 1247 614 1251 618
rect 1450 617 1456 621
rect 1520 617 1524 621
rect 1579 617 1583 621
rect 1604 617 1608 621
rect 1635 617 1639 621
rect 1226 608 1230 614
rect 1263 608 1267 614
rect 1520 609 1524 613
rect 1563 610 1567 614
rect 1585 609 1592 613
rect 1635 610 1639 614
rect 1285 605 1289 609
rect 1506 605 1510 609
rect 1538 605 1542 609
rect 1556 605 1560 609
rect 1613 605 1617 609
rect 1628 605 1632 609
rect 1656 605 1660 609
rect 712 591 716 595
rect 720 592 724 596
rect 732 592 736 596
rect 767 592 771 596
rect 795 591 799 595
rect 847 592 851 596
rect 1152 595 1156 599
rect 1168 595 1172 599
rect 1213 601 1217 605
rect 1189 595 1193 601
rect 1205 595 1209 599
rect 876 591 880 595
rect 1226 595 1230 599
rect 1247 595 1251 601
rect 1263 595 1267 599
rect 1501 593 1505 597
rect 505 575 511 579
rect 573 575 577 579
rect 598 572 602 576
rect 605 575 609 579
rect 623 575 627 579
rect 645 572 649 576
rect 670 572 674 576
rect 680 575 684 579
rect 696 575 700 579
rect 716 572 720 576
rect 723 575 727 579
rect 236 568 240 572
rect 286 568 290 572
rect 337 568 341 572
rect 541 568 547 572
rect 583 565 587 569
rect 599 565 603 569
rect 630 565 634 569
rect 652 565 656 569
rect 717 565 721 569
rect 777 571 781 575
rect 1169 582 1173 586
rect 1213 582 1217 586
rect 1233 582 1237 586
rect 1270 584 1274 588
rect 1533 591 1537 595
rect 1553 594 1557 598
rect 1572 590 1576 594
rect 1591 591 1595 595
rect 1610 591 1614 595
rect 1623 592 1627 596
rect 1720 607 1724 611
rect 1801 607 1805 611
rect 1645 591 1649 595
rect 1653 592 1657 596
rect 1665 592 1669 596
rect 1700 592 1704 596
rect 1728 591 1732 595
rect 1780 592 1784 596
rect 1809 591 1813 595
rect 1438 575 1444 579
rect 1506 575 1510 579
rect 858 571 862 575
rect 1531 572 1535 576
rect 1538 575 1542 579
rect 1556 575 1560 579
rect 1578 572 1582 576
rect 1603 572 1607 576
rect 1613 575 1617 579
rect 1629 575 1633 579
rect 1649 572 1653 576
rect 1656 575 1660 579
rect 1169 568 1173 572
rect 1219 568 1223 572
rect 1270 568 1274 572
rect 1474 568 1480 572
rect 1516 565 1520 569
rect 1532 565 1536 569
rect 1563 565 1567 569
rect 1585 565 1589 569
rect 1650 565 1654 569
rect 1710 571 1714 575
rect 1791 571 1795 575
rect 493 558 499 562
rect 572 558 576 562
rect 606 558 610 562
rect 623 558 627 562
rect 679 558 683 562
rect 696 558 700 562
rect 724 558 728 562
rect 1426 558 1432 562
rect 1505 558 1509 562
rect 1539 558 1543 562
rect 1556 558 1560 562
rect 1612 558 1616 562
rect 1629 558 1633 562
rect 1657 558 1661 562
rect 529 551 535 555
rect 583 551 587 555
rect 599 551 603 555
rect 630 551 634 555
rect 652 551 656 555
rect 717 551 721 555
rect 787 551 791 555
rect 573 541 577 545
rect 598 544 602 548
rect 605 541 609 545
rect 623 541 627 545
rect 645 544 649 548
rect 670 544 674 548
rect 680 541 684 545
rect 696 541 700 545
rect 716 544 720 548
rect 723 541 727 545
rect 567 524 571 528
rect 600 525 604 529
rect 620 522 624 526
rect 639 526 643 530
rect 658 525 662 529
rect 677 525 681 529
rect 690 524 694 528
rect 712 525 716 529
rect 720 524 724 528
rect 732 524 736 528
rect 795 529 799 537
rect 892 551 896 555
rect 846 537 850 541
rect 861 537 865 541
rect 1462 551 1468 555
rect 1516 551 1520 555
rect 1532 551 1536 555
rect 1563 551 1567 555
rect 1585 551 1589 555
rect 1650 551 1654 555
rect 1720 551 1724 555
rect 764 523 768 527
rect 818 528 822 532
rect 573 511 577 515
rect 605 511 609 515
rect 623 511 627 515
rect 680 511 684 515
rect 695 511 699 515
rect 723 511 727 515
rect 587 507 591 511
rect 630 506 634 510
rect 652 507 659 511
rect 702 506 706 510
rect 517 499 523 503
rect 587 499 591 503
rect 646 499 650 503
rect 671 499 675 503
rect 702 499 706 503
rect 777 515 781 519
rect 900 529 904 537
rect 1506 541 1510 545
rect 1531 544 1535 548
rect 1538 541 1542 545
rect 1556 541 1560 545
rect 1578 544 1582 548
rect 1603 544 1607 548
rect 1613 541 1617 545
rect 1629 541 1633 545
rect 1649 544 1653 548
rect 1656 541 1660 545
rect 921 529 925 533
rect 869 523 873 527
rect 1500 524 1504 528
rect 882 515 886 519
rect 1533 525 1537 529
rect 1553 522 1557 526
rect 1572 526 1576 530
rect 1591 525 1595 529
rect 1610 525 1614 529
rect 1623 524 1627 528
rect 1645 525 1649 529
rect 1653 524 1657 528
rect 1665 524 1669 528
rect 1728 529 1732 537
rect 1825 551 1829 555
rect 1779 537 1783 541
rect 1794 537 1798 541
rect 1697 523 1701 527
rect 1751 528 1755 532
rect 1506 511 1510 515
rect 1538 511 1542 515
rect 1556 511 1560 515
rect 1613 511 1617 515
rect 1628 511 1632 515
rect 1656 511 1660 515
rect 1520 507 1524 511
rect 1563 506 1567 510
rect 1585 507 1592 511
rect 1635 506 1639 510
rect 1450 499 1456 503
rect 1520 499 1524 503
rect 1579 499 1583 503
rect 1604 499 1608 503
rect 1635 499 1639 503
rect 1710 515 1714 519
rect 1833 529 1837 537
rect 1854 529 1858 533
rect 1802 523 1806 527
rect 1815 515 1819 519
rect 505 492 511 496
rect 573 492 577 496
rect 587 492 591 496
rect 605 492 609 496
rect 623 492 627 496
rect 646 492 650 496
rect 680 492 684 496
rect 695 492 699 496
rect 723 492 727 496
rect 1438 492 1444 496
rect 1506 492 1510 496
rect 1520 492 1524 496
rect 1538 492 1542 496
rect 1556 492 1560 496
rect 1579 492 1583 496
rect 1613 492 1617 496
rect 1628 492 1632 496
rect 1656 492 1660 496
rect 517 485 523 489
rect 587 485 591 489
rect 646 485 650 489
rect 671 485 675 489
rect 702 485 706 489
rect 587 477 591 481
rect 630 478 634 482
rect 652 477 659 481
rect 702 478 706 482
rect 573 473 577 477
rect 605 473 609 477
rect 623 473 627 477
rect 680 473 684 477
rect 695 473 699 477
rect 723 473 727 477
rect 787 476 791 480
rect 1450 485 1456 489
rect 1520 485 1524 489
rect 1579 485 1583 489
rect 1604 485 1608 489
rect 1635 485 1639 489
rect 892 476 896 480
rect 1520 477 1524 481
rect 1563 478 1567 482
rect 1585 477 1592 481
rect 1635 478 1639 482
rect 1506 473 1510 477
rect 1538 473 1542 477
rect 1556 473 1560 477
rect 1613 473 1617 477
rect 1628 473 1632 477
rect 1656 473 1660 477
rect 1720 476 1724 480
rect 1825 476 1829 480
rect 568 461 572 465
rect 600 459 604 463
rect 620 462 624 466
rect 639 458 643 462
rect 658 459 662 463
rect 677 459 681 463
rect 690 460 694 464
rect 712 459 716 463
rect 720 460 724 464
rect 732 460 736 464
rect 766 461 770 465
rect 795 460 799 464
rect 872 461 876 465
rect 900 460 904 464
rect 1501 461 1505 465
rect 573 443 577 447
rect 598 440 602 444
rect 605 443 609 447
rect 623 443 627 447
rect 645 440 649 444
rect 670 440 674 444
rect 680 443 684 447
rect 696 443 700 447
rect 716 440 720 444
rect 723 443 727 447
rect 529 433 535 437
rect 599 433 603 437
rect 630 433 634 437
rect 652 433 656 437
rect 717 433 721 437
rect 777 440 781 444
rect 1533 459 1537 463
rect 1553 462 1557 466
rect 1572 458 1576 462
rect 1591 459 1595 463
rect 1610 459 1614 463
rect 1623 460 1627 464
rect 1645 459 1649 463
rect 1653 460 1657 464
rect 1665 460 1669 464
rect 1699 461 1703 465
rect 1728 460 1732 464
rect 1805 461 1809 465
rect 1833 460 1837 464
rect 882 440 886 444
rect 1506 443 1510 447
rect 1531 440 1535 444
rect 1538 443 1542 447
rect 1556 443 1560 447
rect 1578 440 1582 444
rect 1603 440 1607 444
rect 1613 443 1617 447
rect 1629 443 1633 447
rect 1649 440 1653 444
rect 1656 443 1660 447
rect 1462 433 1468 437
rect 1532 433 1536 437
rect 1563 433 1567 437
rect 1585 433 1589 437
rect 1650 433 1654 437
rect 1710 440 1714 444
rect 1815 440 1819 444
rect 493 426 499 430
rect 572 426 576 430
rect 606 426 610 430
rect 623 426 627 430
rect 679 426 683 430
rect 696 426 700 430
rect 724 426 728 430
rect 1426 426 1432 430
rect 1505 426 1509 430
rect 1539 426 1543 430
rect 1556 426 1560 430
rect 1612 426 1616 430
rect 1629 426 1633 430
rect 1657 426 1661 430
rect 529 419 535 423
rect 599 419 603 423
rect 630 419 634 423
rect 652 419 656 423
rect 717 419 721 423
rect 787 419 791 423
rect 573 409 577 413
rect 598 412 602 416
rect 605 409 609 413
rect 623 409 627 413
rect 645 412 649 416
rect 670 412 674 416
rect 680 409 684 413
rect 696 409 700 413
rect 716 412 720 416
rect 723 409 727 413
rect 567 392 571 396
rect 600 393 604 397
rect 620 390 624 394
rect 639 394 643 398
rect 658 393 662 397
rect 677 393 681 397
rect 690 392 694 396
rect 712 393 716 397
rect 720 392 724 396
rect 732 392 736 396
rect 795 397 799 405
rect 868 419 872 423
rect 822 405 826 409
rect 837 405 841 409
rect 818 397 822 401
rect 764 391 768 395
rect 573 379 577 383
rect 605 379 609 383
rect 623 379 627 383
rect 680 379 684 383
rect 695 379 699 383
rect 723 379 727 383
rect 587 375 591 379
rect 630 374 634 378
rect 652 375 659 379
rect 702 374 706 378
rect 517 367 523 371
rect 587 367 591 371
rect 646 367 650 371
rect 671 367 675 371
rect 702 367 706 371
rect 777 383 781 387
rect 876 397 880 405
rect 958 419 962 423
rect 912 405 916 409
rect 927 405 931 409
rect 1462 419 1468 423
rect 1532 419 1536 423
rect 1563 419 1567 423
rect 1585 419 1589 423
rect 1650 419 1654 423
rect 1720 419 1724 423
rect 900 397 904 401
rect 845 391 849 395
rect 934 399 938 403
rect 966 397 970 405
rect 1506 409 1510 413
rect 1531 412 1535 416
rect 1538 409 1542 413
rect 1556 409 1560 413
rect 1578 412 1582 416
rect 1603 412 1607 416
rect 1613 409 1617 413
rect 1629 409 1633 413
rect 1649 412 1653 416
rect 1656 409 1660 413
rect 858 383 862 387
rect 1001 396 1005 400
rect 1500 392 1504 396
rect 948 383 952 387
rect 1533 393 1537 397
rect 1553 390 1557 394
rect 1572 394 1576 398
rect 1591 393 1595 397
rect 1610 393 1614 397
rect 1623 392 1627 396
rect 1645 393 1649 397
rect 1653 392 1657 396
rect 1665 392 1669 396
rect 1728 397 1732 405
rect 1801 419 1805 423
rect 1755 405 1759 409
rect 1770 405 1774 409
rect 1751 397 1755 401
rect 1697 391 1701 395
rect 1506 379 1510 383
rect 1538 379 1542 383
rect 1556 379 1560 383
rect 1613 379 1617 383
rect 1628 379 1632 383
rect 1656 379 1660 383
rect 1520 375 1524 379
rect 1563 374 1567 378
rect 1585 375 1592 379
rect 1635 374 1639 378
rect 1450 367 1456 371
rect 1520 367 1524 371
rect 1579 367 1583 371
rect 1604 367 1608 371
rect 1635 367 1639 371
rect 1710 383 1714 387
rect 1809 397 1813 405
rect 1891 419 1895 423
rect 1845 405 1849 409
rect 1860 405 1864 409
rect 1833 397 1837 401
rect 1778 391 1782 395
rect 1867 399 1871 403
rect 1899 397 1903 405
rect 1791 383 1795 387
rect 1934 396 1938 400
rect 1881 383 1885 387
rect 505 360 511 364
rect 573 360 577 364
rect 587 360 591 364
rect 605 360 609 364
rect 623 360 627 364
rect 646 360 650 364
rect 680 360 684 364
rect 695 360 699 364
rect 723 360 727 364
rect 1438 360 1444 364
rect 1506 360 1510 364
rect 1520 360 1524 364
rect 1538 360 1542 364
rect 1556 360 1560 364
rect 1579 360 1583 364
rect 1613 360 1617 364
rect 1628 360 1632 364
rect 1656 360 1660 364
rect 517 353 523 357
rect 587 353 591 357
rect 646 353 650 357
rect 671 353 675 357
rect 702 353 706 357
rect 587 345 591 349
rect 630 346 634 350
rect 652 345 659 349
rect 702 346 706 350
rect 573 341 577 345
rect 605 341 609 345
rect 623 341 627 345
rect 680 341 684 345
rect 695 341 699 345
rect 723 341 727 345
rect 568 329 572 333
rect 600 327 604 331
rect 620 330 624 334
rect 639 326 643 330
rect 658 327 662 331
rect 677 327 681 331
rect 690 328 694 332
rect 787 341 791 345
rect 868 341 872 345
rect 1450 353 1456 357
rect 1520 353 1524 357
rect 1579 353 1583 357
rect 1604 353 1608 357
rect 1635 353 1639 357
rect 1520 345 1524 349
rect 1563 346 1567 350
rect 1585 345 1592 349
rect 1635 346 1639 350
rect 958 341 962 345
rect 1506 341 1510 345
rect 1538 341 1542 345
rect 1556 341 1560 345
rect 1613 341 1617 345
rect 1628 341 1632 345
rect 1656 341 1660 345
rect 712 327 716 331
rect 720 328 724 332
rect 732 328 736 332
rect 767 326 771 330
rect 795 325 799 329
rect 847 326 851 330
rect 876 325 880 329
rect 931 326 935 330
rect 1501 329 1505 333
rect 966 325 970 329
rect 573 311 577 315
rect 598 308 602 312
rect 605 311 609 315
rect 623 311 627 315
rect 645 308 649 312
rect 670 308 674 312
rect 680 311 684 315
rect 696 311 700 315
rect 716 308 720 312
rect 723 311 727 315
rect 1533 327 1537 331
rect 1553 330 1557 334
rect 1572 326 1576 330
rect 1591 327 1595 331
rect 1610 327 1614 331
rect 1623 328 1627 332
rect 1720 341 1724 345
rect 1801 341 1805 345
rect 1891 341 1895 345
rect 1645 327 1649 331
rect 1653 328 1657 332
rect 1665 328 1669 332
rect 1700 326 1704 330
rect 1728 325 1732 329
rect 1780 326 1784 330
rect 1809 325 1813 329
rect 1864 326 1868 330
rect 1899 325 1903 329
rect 529 301 535 305
rect 599 301 603 305
rect 630 301 634 305
rect 652 301 656 305
rect 717 301 721 305
rect 777 305 781 309
rect 858 305 862 309
rect 1506 311 1510 315
rect 948 305 952 309
rect 1531 308 1535 312
rect 1538 311 1542 315
rect 1556 311 1560 315
rect 1578 308 1582 312
rect 1603 308 1607 312
rect 1613 311 1617 315
rect 1629 311 1633 315
rect 1649 308 1653 312
rect 1656 311 1660 315
rect 1462 301 1468 305
rect 1532 301 1536 305
rect 1563 301 1567 305
rect 1585 301 1589 305
rect 1650 301 1654 305
rect 1710 305 1714 309
rect 1791 305 1795 309
rect 1881 305 1885 309
rect 493 294 499 298
rect 572 294 576 298
rect 606 294 610 298
rect 623 294 627 298
rect 679 294 683 298
rect 696 294 700 298
rect 724 294 728 298
rect 1426 294 1432 298
rect 1505 294 1509 298
rect 1539 294 1543 298
rect 1556 294 1560 298
rect 1612 294 1616 298
rect 1629 294 1633 298
rect 1657 294 1661 298
rect 529 287 535 291
rect 599 287 603 291
rect 630 287 634 291
rect 652 287 656 291
rect 717 287 721 291
rect 787 287 791 291
rect 573 277 577 281
rect 598 280 602 284
rect 605 277 609 281
rect 623 277 627 281
rect 645 280 649 284
rect 670 280 674 284
rect 680 277 684 281
rect 696 277 700 281
rect 716 280 720 284
rect 723 277 727 281
rect 567 260 571 264
rect 600 261 604 265
rect 620 258 624 262
rect 639 262 643 266
rect 1462 287 1468 291
rect 1532 287 1536 291
rect 1563 287 1567 291
rect 1585 287 1589 291
rect 1650 287 1654 291
rect 1720 287 1724 291
rect 658 261 662 265
rect 677 261 681 265
rect 690 260 694 264
rect 712 261 716 265
rect 720 260 724 264
rect 732 260 736 264
rect 795 265 799 273
rect 1506 277 1510 281
rect 1531 280 1535 284
rect 1538 277 1542 281
rect 1556 277 1560 281
rect 1578 280 1582 284
rect 1603 280 1607 284
rect 1613 277 1617 281
rect 1629 277 1633 281
rect 1649 280 1653 284
rect 1656 277 1660 281
rect 764 259 768 263
rect 818 264 822 268
rect 1500 260 1504 264
rect 573 247 577 251
rect 605 247 609 251
rect 623 247 627 251
rect 680 247 684 251
rect 695 247 699 251
rect 723 247 727 251
rect 587 243 591 247
rect 102 239 106 243
rect 138 239 142 243
rect 205 239 209 243
rect 234 239 238 243
rect 270 239 274 243
rect 337 239 341 243
rect 366 239 370 243
rect 402 239 406 243
rect 469 239 473 243
rect 553 239 559 243
rect 630 242 634 246
rect 652 243 659 247
rect 702 242 706 246
rect 493 232 499 236
rect 587 235 591 239
rect 596 235 600 239
rect 646 235 650 239
rect 671 235 675 239
rect 702 235 706 239
rect 777 251 781 255
rect 1533 261 1537 265
rect 1553 258 1557 262
rect 1572 262 1576 266
rect 1591 261 1595 265
rect 1610 261 1614 265
rect 1623 260 1627 264
rect 1645 261 1649 265
rect 1653 260 1657 264
rect 1665 260 1669 264
rect 1728 265 1732 273
rect 1697 259 1701 263
rect 1751 264 1755 268
rect 1506 247 1510 251
rect 1538 247 1542 251
rect 1556 247 1560 251
rect 1613 247 1617 251
rect 1628 247 1632 251
rect 1656 247 1660 251
rect 1520 243 1524 247
rect 1035 239 1039 243
rect 1071 239 1075 243
rect 1138 239 1142 243
rect 1167 239 1171 243
rect 1203 239 1207 243
rect 1270 239 1274 243
rect 1299 239 1303 243
rect 1335 239 1339 243
rect 1402 239 1406 243
rect 1486 239 1492 243
rect 1563 242 1567 246
rect 1585 243 1592 247
rect 1635 242 1639 246
rect 1426 232 1432 236
rect 1520 235 1524 239
rect 1529 235 1533 239
rect 1579 235 1583 239
rect 1604 235 1608 239
rect 1635 235 1639 239
rect 1710 251 1714 255
rect 102 225 106 229
rect 152 225 156 229
rect 205 225 209 229
rect 234 225 238 229
rect 284 225 288 229
rect 337 225 341 229
rect 366 225 370 229
rect 416 225 420 229
rect 469 225 473 229
rect 505 228 511 232
rect 573 228 577 232
rect 587 228 591 232
rect 605 228 609 232
rect 623 228 627 232
rect 646 228 650 232
rect 680 228 684 232
rect 695 228 699 232
rect 723 228 727 232
rect 848 228 852 232
rect 866 228 870 232
rect 884 228 888 232
rect 907 228 911 232
rect 941 228 945 232
rect 956 228 960 232
rect 984 228 988 232
rect 125 214 129 218
rect 96 205 100 209
rect 109 208 113 214
rect 146 208 150 214
rect 159 210 163 214
rect 183 214 187 218
rect 257 214 261 218
rect 167 208 171 214
rect 204 208 208 214
rect 220 208 224 214
rect 241 208 245 214
rect 278 208 282 214
rect 291 210 295 214
rect 315 214 319 218
rect 389 214 393 218
rect 299 208 303 214
rect 336 208 340 214
rect 352 208 356 214
rect 373 208 377 214
rect 410 208 414 214
rect 423 210 427 214
rect 447 214 451 218
rect 517 221 523 225
rect 587 221 591 225
rect 596 221 600 225
rect 646 221 650 225
rect 671 221 675 225
rect 702 221 706 225
rect 431 208 435 214
rect 468 208 472 214
rect 484 210 488 214
rect 587 213 591 217
rect 630 214 634 218
rect 652 213 659 217
rect 702 214 706 218
rect 573 209 577 213
rect 605 209 609 213
rect 623 209 627 213
rect 680 209 684 213
rect 695 209 699 213
rect 723 209 727 213
rect 109 195 113 199
rect 125 195 129 201
rect 159 201 163 205
rect 146 195 150 199
rect 167 195 171 199
rect 183 195 187 201
rect 204 195 208 199
rect 220 195 224 199
rect 241 195 245 199
rect 257 195 261 201
rect 291 201 295 205
rect 278 195 282 199
rect 299 195 303 199
rect 315 195 319 201
rect 336 195 340 199
rect 352 195 356 199
rect 373 195 377 199
rect 389 195 393 201
rect 423 201 427 205
rect 410 195 414 199
rect 431 195 435 199
rect 447 195 451 201
rect 468 195 472 199
rect 484 195 488 199
rect 568 197 572 201
rect 102 184 106 188
rect 139 182 143 186
rect 159 182 163 186
rect 203 182 207 186
rect 234 184 238 188
rect 271 182 275 186
rect 291 182 295 186
rect 335 182 339 186
rect 366 184 370 188
rect 403 182 407 186
rect 423 182 427 186
rect 467 182 471 186
rect 600 195 604 199
rect 620 198 624 202
rect 639 194 643 198
rect 658 195 662 199
rect 677 195 681 199
rect 690 196 694 200
rect 826 221 830 225
rect 848 221 852 225
rect 907 221 911 225
rect 932 221 936 225
rect 963 221 967 225
rect 1035 225 1039 229
rect 1085 225 1089 229
rect 1138 225 1142 229
rect 1167 225 1171 229
rect 1217 225 1221 229
rect 1270 225 1274 229
rect 1299 225 1303 229
rect 1349 225 1353 229
rect 1402 225 1406 229
rect 1438 228 1444 232
rect 1506 228 1510 232
rect 1520 228 1524 232
rect 1538 228 1542 232
rect 1556 228 1560 232
rect 1579 228 1583 232
rect 1613 228 1617 232
rect 1628 228 1632 232
rect 1656 228 1660 232
rect 1781 228 1785 232
rect 1799 228 1803 232
rect 1817 228 1821 232
rect 1840 228 1844 232
rect 1874 228 1878 232
rect 1889 228 1893 232
rect 1917 228 1921 232
rect 848 213 852 217
rect 891 214 895 218
rect 913 213 920 217
rect 963 214 967 218
rect 1058 214 1062 218
rect 866 209 870 213
rect 884 209 888 213
rect 941 209 945 213
rect 956 209 960 213
rect 984 209 988 213
rect 787 205 791 209
rect 712 195 716 199
rect 720 196 724 200
rect 732 196 736 200
rect 766 190 770 194
rect 806 196 810 200
rect 795 189 799 193
rect 573 179 577 183
rect 505 175 511 179
rect 598 176 602 180
rect 605 179 609 183
rect 623 179 627 183
rect 645 176 649 180
rect 670 176 674 180
rect 680 179 684 183
rect 696 179 700 183
rect 716 176 720 180
rect 723 179 727 183
rect 861 195 865 199
rect 881 198 885 202
rect 900 194 904 198
rect 1029 205 1033 209
rect 1042 208 1046 214
rect 1079 208 1083 214
rect 1092 210 1096 214
rect 1116 214 1120 218
rect 1190 214 1194 218
rect 1100 208 1104 214
rect 1137 208 1141 214
rect 1153 208 1157 214
rect 1174 208 1178 214
rect 1211 208 1215 214
rect 1224 210 1228 214
rect 1248 214 1252 218
rect 1322 214 1326 218
rect 1232 208 1236 214
rect 1269 208 1273 214
rect 1285 208 1289 214
rect 1306 208 1310 214
rect 1343 208 1347 214
rect 1356 210 1360 214
rect 1380 214 1384 218
rect 1450 221 1456 225
rect 1520 221 1524 225
rect 1529 221 1533 225
rect 1579 221 1583 225
rect 1604 221 1608 225
rect 1635 221 1639 225
rect 1364 208 1368 214
rect 1401 208 1405 214
rect 1417 210 1421 214
rect 1520 213 1524 217
rect 1563 214 1567 218
rect 1585 213 1592 217
rect 1635 214 1639 218
rect 1506 209 1510 213
rect 1538 209 1542 213
rect 1556 209 1560 213
rect 1613 209 1617 213
rect 1628 209 1632 213
rect 1656 209 1660 213
rect 919 195 923 199
rect 938 195 942 199
rect 951 196 955 200
rect 973 195 977 199
rect 981 196 985 200
rect 993 196 997 200
rect 1042 195 1046 199
rect 1058 195 1062 201
rect 1092 201 1096 205
rect 1079 195 1083 199
rect 1100 195 1104 199
rect 1116 195 1120 201
rect 1137 195 1141 199
rect 1153 195 1157 199
rect 1174 195 1178 199
rect 1190 195 1194 201
rect 1224 201 1228 205
rect 1211 195 1215 199
rect 1232 195 1236 199
rect 1248 195 1252 201
rect 1269 195 1273 199
rect 1285 195 1289 199
rect 1306 195 1310 199
rect 1322 195 1326 201
rect 1356 201 1360 205
rect 1343 195 1347 199
rect 1364 195 1368 199
rect 1380 195 1384 201
rect 1401 195 1405 199
rect 1417 195 1421 199
rect 1501 197 1505 201
rect 807 179 811 183
rect 833 179 837 183
rect 102 168 106 172
rect 153 168 157 172
rect 203 168 207 172
rect 234 168 238 172
rect 285 168 289 172
rect 335 168 339 172
rect 366 168 370 172
rect 417 168 421 172
rect 467 168 471 172
rect 541 169 547 173
rect 581 169 585 173
rect 599 169 603 173
rect 630 169 634 173
rect 652 169 656 173
rect 717 169 721 173
rect 859 176 863 180
rect 866 179 870 183
rect 884 179 888 183
rect 906 176 910 180
rect 931 176 935 180
rect 941 179 945 183
rect 957 179 961 183
rect 977 176 981 180
rect 984 179 988 183
rect 1035 184 1039 188
rect 1072 182 1076 186
rect 1092 182 1096 186
rect 1136 182 1140 186
rect 1167 184 1171 188
rect 1204 182 1208 186
rect 1224 182 1228 186
rect 1268 182 1272 186
rect 1299 184 1303 188
rect 1336 182 1340 186
rect 1356 182 1360 186
rect 1400 182 1404 186
rect 1533 195 1537 199
rect 1553 198 1557 202
rect 1572 194 1576 198
rect 1591 195 1595 199
rect 1610 195 1614 199
rect 1623 196 1627 200
rect 1759 221 1763 225
rect 1781 221 1785 225
rect 1840 221 1844 225
rect 1865 221 1869 225
rect 1896 221 1900 225
rect 1781 213 1785 217
rect 1824 214 1828 218
rect 1846 213 1853 217
rect 1896 214 1900 218
rect 1799 209 1803 213
rect 1817 209 1821 213
rect 1874 209 1878 213
rect 1889 209 1893 213
rect 1917 209 1921 213
rect 1720 205 1724 209
rect 1645 195 1649 199
rect 1653 196 1657 200
rect 1665 196 1669 200
rect 1699 190 1703 194
rect 1739 196 1743 200
rect 1728 189 1732 193
rect 1506 179 1510 183
rect 1438 175 1444 179
rect 1531 176 1535 180
rect 1538 179 1542 183
rect 1556 179 1560 183
rect 1578 176 1582 180
rect 1603 176 1607 180
rect 1613 179 1617 183
rect 1629 179 1633 183
rect 1649 176 1653 180
rect 1656 179 1660 183
rect 1794 195 1798 199
rect 1814 198 1818 202
rect 1833 194 1837 198
rect 1852 195 1856 199
rect 1871 195 1875 199
rect 1884 196 1888 200
rect 1906 195 1910 199
rect 1914 196 1918 200
rect 1926 196 1930 200
rect 1740 179 1744 183
rect 1766 179 1770 183
rect 777 169 781 173
rect 816 169 820 173
rect 860 169 864 173
rect 891 169 895 173
rect 913 169 917 173
rect 978 169 982 173
rect 1035 168 1039 172
rect 1086 168 1090 172
rect 1136 168 1140 172
rect 1167 168 1171 172
rect 1218 168 1222 172
rect 1268 168 1272 172
rect 1299 168 1303 172
rect 1350 168 1354 172
rect 1400 168 1404 172
rect 1474 169 1480 173
rect 1514 169 1518 173
rect 1532 169 1536 173
rect 1563 169 1567 173
rect 1585 169 1589 173
rect 1650 169 1654 173
rect 1792 176 1796 180
rect 1799 179 1803 183
rect 1817 179 1821 183
rect 1839 176 1843 180
rect 1864 176 1868 180
rect 1874 179 1878 183
rect 1890 179 1894 183
rect 1910 176 1914 180
rect 1917 179 1921 183
rect 1710 169 1714 173
rect 1749 169 1753 173
rect 1793 169 1797 173
rect 1824 169 1828 173
rect 1846 169 1850 173
rect 1911 169 1915 173
rect 96 161 100 165
rect 484 161 488 165
rect 493 162 499 166
rect 572 162 576 166
rect 606 162 610 166
rect 623 162 627 166
rect 679 162 683 166
rect 696 162 700 166
rect 724 162 728 166
rect 807 162 811 166
rect 833 162 837 166
rect 867 162 871 166
rect 884 162 888 166
rect 940 162 944 166
rect 957 162 961 166
rect 985 162 989 166
rect 1029 161 1033 165
rect 1417 161 1421 165
rect 1426 162 1432 166
rect 1505 162 1509 166
rect 1539 162 1543 166
rect 1556 162 1560 166
rect 1612 162 1616 166
rect 1629 162 1633 166
rect 1657 162 1661 166
rect 1740 162 1744 166
rect 1766 162 1770 166
rect 1800 162 1804 166
rect 1817 162 1821 166
rect 1873 162 1877 166
rect 1890 162 1894 166
rect 1918 162 1922 166
rect 219 154 224 158
rect 352 154 356 158
rect 529 155 535 159
rect 581 155 585 159
rect 815 155 819 159
rect 1001 156 1005 160
rect 1013 156 1017 160
rect 1152 154 1157 158
rect 1285 154 1289 158
rect 1462 155 1468 159
rect 1514 155 1518 159
rect 1748 155 1752 159
rect 1934 156 1938 160
rect 1946 156 1950 160
rect 227 147 231 151
rect 517 147 523 151
rect 825 148 829 152
rect 990 148 994 152
rect 211 143 215 147
rect 243 143 247 147
rect 1160 147 1164 151
rect 1450 147 1456 151
rect 1758 148 1762 152
rect 1923 148 1927 152
rect 1144 143 1148 147
rect 1176 143 1180 147
rect 211 136 215 140
rect 243 136 247 140
rect 1144 136 1148 140
rect 1176 136 1180 140
rect 227 129 231 133
rect 484 129 488 133
rect 553 129 559 133
rect 873 129 877 133
rect 909 129 913 133
rect 976 129 980 133
rect 1160 129 1164 133
rect 1417 129 1421 133
rect 1486 129 1492 133
rect 1806 129 1810 133
rect 1842 129 1846 133
rect 1909 129 1913 133
rect 484 121 488 125
rect 493 122 499 126
rect 859 122 863 126
rect 211 117 215 121
rect 243 117 247 121
rect 227 113 231 117
rect 873 115 877 119
rect 923 115 927 119
rect 976 115 980 119
rect 1417 121 1421 125
rect 1426 122 1432 126
rect 1792 122 1796 126
rect 1144 117 1148 121
rect 1176 117 1180 121
rect 1160 113 1164 117
rect 1806 115 1810 119
rect 1856 115 1860 119
rect 1909 115 1913 119
rect 219 106 224 110
rect 353 106 357 110
rect 896 104 900 108
rect 102 99 106 103
rect 138 99 142 103
rect 205 99 209 103
rect 234 99 238 103
rect 270 99 274 103
rect 337 99 341 103
rect 366 99 370 103
rect 402 99 406 103
rect 469 99 473 103
rect 553 99 559 103
rect 493 92 499 96
rect 867 95 871 99
rect 880 98 884 104
rect 917 98 921 104
rect 930 100 934 104
rect 954 104 958 108
rect 1152 106 1157 110
rect 1286 106 1290 110
rect 1829 104 1833 108
rect 938 98 942 104
rect 975 98 979 104
rect 991 98 995 104
rect 1035 99 1039 103
rect 1071 99 1075 103
rect 1138 99 1142 103
rect 1167 99 1171 103
rect 1203 99 1207 103
rect 1270 99 1274 103
rect 1299 99 1303 103
rect 1335 99 1339 103
rect 1402 99 1406 103
rect 1486 99 1492 103
rect 102 85 106 89
rect 152 85 156 89
rect 205 85 209 89
rect 234 85 238 89
rect 284 85 288 89
rect 337 85 341 89
rect 366 85 370 89
rect 416 85 420 89
rect 469 85 473 89
rect 880 85 884 89
rect 896 85 900 91
rect 930 91 934 95
rect 917 85 921 89
rect 125 74 129 78
rect 96 65 100 69
rect 109 68 113 74
rect 146 68 150 74
rect 159 70 163 74
rect 183 74 187 78
rect 257 74 261 78
rect 167 68 171 74
rect 204 68 208 74
rect 220 68 224 74
rect 241 68 245 74
rect 278 68 282 74
rect 291 70 295 74
rect 315 74 319 78
rect 389 74 393 78
rect 299 68 303 74
rect 336 68 340 74
rect 352 68 356 74
rect 373 68 377 74
rect 410 68 414 74
rect 423 70 427 74
rect 447 74 451 78
rect 431 68 435 74
rect 468 68 472 74
rect 484 70 488 74
rect 938 85 942 89
rect 954 85 958 91
rect 1426 92 1432 96
rect 1800 95 1804 99
rect 1813 98 1817 104
rect 1850 98 1854 104
rect 1863 100 1867 104
rect 1887 104 1891 108
rect 1871 98 1875 104
rect 1908 98 1912 104
rect 1924 98 1928 104
rect 975 85 979 89
rect 991 85 995 89
rect 1035 85 1039 89
rect 1085 85 1089 89
rect 1138 85 1142 89
rect 1167 85 1171 89
rect 1217 85 1221 89
rect 1270 85 1274 89
rect 1299 85 1303 89
rect 1349 85 1353 89
rect 1402 85 1406 89
rect 1813 85 1817 89
rect 1829 85 1833 91
rect 1863 91 1867 95
rect 1850 85 1854 89
rect 873 74 877 78
rect 910 72 914 76
rect 930 72 934 76
rect 974 72 978 76
rect 1058 74 1062 78
rect 109 55 113 59
rect 125 55 129 61
rect 159 61 163 65
rect 146 55 150 59
rect 167 55 171 59
rect 183 55 187 61
rect 204 55 208 59
rect 220 55 224 59
rect 241 55 245 59
rect 257 55 261 61
rect 291 61 295 65
rect 278 55 282 59
rect 299 55 303 59
rect 315 55 319 61
rect 336 55 340 59
rect 352 55 356 59
rect 373 55 377 59
rect 389 55 393 61
rect 423 61 427 65
rect 410 55 414 59
rect 431 55 435 59
rect 447 55 451 61
rect 505 65 511 69
rect 1029 65 1033 69
rect 1042 68 1046 74
rect 1079 68 1083 74
rect 1092 70 1096 74
rect 1116 74 1120 78
rect 1190 74 1194 78
rect 1100 68 1104 74
rect 1137 68 1141 74
rect 1153 68 1157 74
rect 1174 68 1178 74
rect 1211 68 1215 74
rect 1224 70 1228 74
rect 1248 74 1252 78
rect 1322 74 1326 78
rect 1232 68 1236 74
rect 1269 68 1273 74
rect 1285 68 1289 74
rect 1306 68 1310 74
rect 1343 68 1347 74
rect 1356 70 1360 74
rect 1380 74 1384 78
rect 1364 68 1368 74
rect 1401 68 1405 74
rect 1417 70 1421 74
rect 1871 85 1875 89
rect 1887 85 1891 91
rect 1908 85 1912 89
rect 1924 85 1928 89
rect 1806 74 1810 78
rect 1843 72 1847 76
rect 1863 72 1867 76
rect 1907 72 1911 76
rect 468 55 472 59
rect 484 55 488 59
rect 541 58 547 62
rect 873 58 877 62
rect 924 58 928 62
rect 974 58 978 62
rect 1042 55 1046 59
rect 1058 55 1062 61
rect 1092 61 1096 65
rect 1079 55 1083 59
rect 102 44 106 48
rect 139 42 143 46
rect 159 42 163 46
rect 203 42 207 46
rect 234 44 238 48
rect 271 42 275 46
rect 291 42 295 46
rect 335 42 339 46
rect 366 44 370 48
rect 403 42 407 46
rect 423 42 427 46
rect 467 42 471 46
rect 866 50 870 54
rect 991 51 995 55
rect 1100 55 1104 59
rect 1116 55 1120 61
rect 1137 55 1141 59
rect 1153 55 1157 59
rect 1174 55 1178 59
rect 1190 55 1194 61
rect 1224 61 1228 65
rect 1211 55 1215 59
rect 1232 55 1236 59
rect 1248 55 1252 61
rect 1269 55 1273 59
rect 1285 55 1289 59
rect 1306 55 1310 59
rect 1322 55 1326 61
rect 1356 61 1360 65
rect 1343 55 1347 59
rect 1364 55 1368 59
rect 1380 55 1384 61
rect 1438 65 1444 69
rect 1401 55 1405 59
rect 1417 55 1421 59
rect 1474 58 1480 62
rect 1806 58 1810 62
rect 1857 58 1861 62
rect 1907 58 1911 62
rect 553 43 559 47
rect 873 43 877 47
rect 909 43 913 47
rect 976 43 980 47
rect 505 35 511 39
rect 859 36 863 40
rect 1035 44 1039 48
rect 1072 42 1076 46
rect 1092 42 1096 46
rect 1136 42 1140 46
rect 1167 44 1171 48
rect 1204 42 1208 46
rect 1224 42 1228 46
rect 1268 42 1272 46
rect 1299 44 1303 48
rect 1336 42 1340 46
rect 1356 42 1360 46
rect 1400 42 1404 46
rect 1799 50 1803 54
rect 1924 51 1928 55
rect 1486 43 1492 47
rect 1806 43 1810 47
rect 1842 43 1846 47
rect 1909 43 1913 47
rect 102 28 106 32
rect 153 28 157 32
rect 203 28 207 32
rect 234 28 238 32
rect 285 28 289 32
rect 335 28 339 32
rect 366 28 370 32
rect 417 28 421 32
rect 467 28 471 32
rect 541 28 547 32
rect 873 29 877 33
rect 923 29 927 33
rect 976 29 980 33
rect 1438 35 1444 39
rect 1792 36 1796 40
rect 1035 28 1039 32
rect 1086 28 1090 32
rect 1136 28 1140 32
rect 1167 28 1171 32
rect 1218 28 1222 32
rect 1268 28 1272 32
rect 1299 28 1303 32
rect 1350 28 1354 32
rect 1400 28 1404 32
rect 1474 28 1480 32
rect 1806 29 1810 33
rect 1856 29 1860 33
rect 1909 29 1913 33
rect 95 21 99 25
rect 484 21 488 25
rect 896 18 900 22
rect 102 13 106 17
rect 138 13 142 17
rect 205 13 209 17
rect 234 13 238 17
rect 270 13 274 17
rect 337 13 341 17
rect 366 13 370 17
rect 402 13 406 17
rect 469 13 473 17
rect 553 13 559 17
rect 493 6 499 10
rect 867 9 871 13
rect 880 12 884 18
rect 917 12 921 18
rect 930 14 934 18
rect 954 18 958 22
rect 1028 21 1032 25
rect 1417 21 1421 25
rect 1829 18 1833 22
rect 938 12 942 18
rect 975 12 979 18
rect 991 14 995 18
rect 1013 12 1017 16
rect 1035 13 1039 17
rect 1071 13 1075 17
rect 1138 13 1142 17
rect 1167 13 1171 17
rect 1203 13 1207 17
rect 1270 13 1274 17
rect 1299 13 1303 17
rect 1335 13 1339 17
rect 1402 13 1406 17
rect 1486 13 1492 17
rect 102 -1 106 3
rect 152 -1 156 3
rect 205 -1 209 3
rect 234 -1 238 3
rect 284 -1 288 3
rect 337 -1 341 3
rect 366 -1 370 3
rect 416 -1 420 3
rect 469 -1 473 3
rect 880 -1 884 3
rect 896 -1 900 5
rect 930 5 934 9
rect 917 -1 921 3
rect 125 -12 129 -8
rect 96 -21 100 -17
rect 109 -18 113 -12
rect 146 -18 150 -12
rect 159 -16 163 -12
rect 183 -12 187 -8
rect 257 -12 261 -8
rect 167 -18 171 -12
rect 204 -18 208 -12
rect 220 -18 224 -12
rect 241 -18 245 -12
rect 278 -18 282 -12
rect 291 -16 295 -12
rect 315 -12 319 -8
rect 389 -12 393 -8
rect 299 -18 303 -12
rect 336 -18 340 -12
rect 352 -18 356 -12
rect 373 -18 377 -12
rect 410 -18 414 -12
rect 423 -16 427 -12
rect 447 -12 451 -8
rect 431 -18 435 -12
rect 468 -18 472 -12
rect 484 -16 488 -12
rect 938 -1 942 3
rect 954 -1 958 5
rect 975 -1 979 3
rect 991 -1 995 8
rect 1426 6 1432 10
rect 1800 9 1804 13
rect 1813 12 1817 18
rect 1850 12 1854 18
rect 1863 14 1867 18
rect 1887 18 1891 22
rect 1871 12 1875 18
rect 1908 12 1912 18
rect 1924 14 1928 18
rect 1946 12 1950 16
rect 1013 -4 1017 0
rect 1035 -1 1039 3
rect 1085 -1 1089 3
rect 1138 -1 1142 3
rect 1167 -1 1171 3
rect 1217 -1 1221 3
rect 1270 -1 1274 3
rect 1299 -1 1303 3
rect 1349 -1 1353 3
rect 1402 -1 1406 3
rect 1813 -1 1817 3
rect 1829 -1 1833 5
rect 1863 5 1867 9
rect 1850 -1 1854 3
rect 873 -12 877 -8
rect 910 -14 914 -10
rect 930 -14 934 -10
rect 974 -14 978 -10
rect 1058 -12 1062 -8
rect 109 -31 113 -27
rect 125 -31 129 -25
rect 159 -25 163 -21
rect 146 -31 150 -27
rect 167 -31 171 -27
rect 183 -31 187 -25
rect 204 -31 208 -27
rect 220 -31 224 -27
rect 241 -31 245 -27
rect 257 -31 261 -25
rect 291 -25 295 -21
rect 278 -31 282 -27
rect 299 -31 303 -27
rect 315 -31 319 -25
rect 336 -31 340 -27
rect 352 -31 356 -27
rect 373 -31 377 -27
rect 389 -31 393 -25
rect 423 -25 427 -21
rect 410 -31 414 -27
rect 431 -31 435 -27
rect 447 -31 451 -25
rect 505 -21 511 -17
rect 1029 -21 1033 -17
rect 1042 -18 1046 -12
rect 1079 -18 1083 -12
rect 1092 -16 1096 -12
rect 1116 -12 1120 -8
rect 1190 -12 1194 -8
rect 1100 -18 1104 -12
rect 1137 -18 1141 -12
rect 1153 -18 1157 -12
rect 1174 -18 1178 -12
rect 1211 -18 1215 -12
rect 1224 -16 1228 -12
rect 1248 -12 1252 -8
rect 1322 -12 1326 -8
rect 1232 -18 1236 -12
rect 1269 -18 1273 -12
rect 1285 -18 1289 -12
rect 1306 -18 1310 -12
rect 1343 -18 1347 -12
rect 1356 -16 1360 -12
rect 1380 -12 1384 -8
rect 1364 -18 1368 -12
rect 1401 -18 1405 -12
rect 1417 -16 1421 -12
rect 1871 -1 1875 3
rect 1887 -1 1891 5
rect 1908 -1 1912 3
rect 1924 -1 1928 8
rect 1946 -4 1950 0
rect 1806 -12 1810 -8
rect 1843 -14 1847 -10
rect 1863 -14 1867 -10
rect 1907 -14 1911 -10
rect 468 -31 472 -27
rect 484 -31 488 -27
rect 541 -28 547 -24
rect 873 -28 877 -24
rect 924 -28 928 -24
rect 974 -28 978 -24
rect 1042 -31 1046 -27
rect 1058 -31 1062 -25
rect 1092 -25 1096 -21
rect 1079 -31 1083 -27
rect 1100 -31 1104 -27
rect 1116 -31 1120 -25
rect 1137 -31 1141 -27
rect 1153 -31 1157 -27
rect 1174 -31 1178 -27
rect 1190 -31 1194 -25
rect 1224 -25 1228 -21
rect 1211 -31 1215 -27
rect 1232 -31 1236 -27
rect 1248 -31 1252 -25
rect 1269 -31 1273 -27
rect 1285 -31 1289 -27
rect 1306 -31 1310 -27
rect 1322 -31 1326 -25
rect 1356 -25 1360 -21
rect 1343 -31 1347 -27
rect 1364 -31 1368 -27
rect 1380 -31 1384 -25
rect 1438 -21 1444 -17
rect 1401 -31 1405 -27
rect 1417 -31 1421 -27
rect 1474 -28 1480 -24
rect 1806 -28 1810 -24
rect 1857 -28 1861 -24
rect 1907 -28 1911 -24
rect 102 -42 106 -38
rect 139 -44 143 -40
rect 159 -44 163 -40
rect 203 -44 207 -40
rect 234 -42 238 -38
rect 271 -44 275 -40
rect 291 -44 295 -40
rect 335 -44 339 -40
rect 366 -42 370 -38
rect 403 -44 407 -40
rect 423 -44 427 -40
rect 467 -44 471 -40
rect 1035 -42 1039 -38
rect 1072 -44 1076 -40
rect 1092 -44 1096 -40
rect 1136 -44 1140 -40
rect 1167 -42 1171 -38
rect 1204 -44 1208 -40
rect 1224 -44 1228 -40
rect 1268 -44 1272 -40
rect 1299 -42 1303 -38
rect 1336 -44 1340 -40
rect 1356 -44 1360 -40
rect 1400 -44 1404 -40
rect 505 -51 511 -47
rect 1438 -51 1444 -47
rect 102 -58 106 -54
rect 153 -58 157 -54
rect 203 -58 207 -54
rect 234 -58 238 -54
rect 285 -58 289 -54
rect 335 -58 339 -54
rect 366 -58 370 -54
rect 417 -58 421 -54
rect 467 -58 471 -54
rect 541 -58 547 -54
rect 1035 -58 1039 -54
rect 1086 -58 1090 -54
rect 1136 -58 1140 -54
rect 1167 -58 1171 -54
rect 1218 -58 1222 -54
rect 1268 -58 1272 -54
rect 1299 -58 1303 -54
rect 1350 -58 1354 -54
rect 1400 -58 1404 -54
rect 1474 -58 1480 -54
rect 95 -65 99 -61
rect 484 -65 488 -61
rect 1028 -65 1032 -61
rect 1417 -65 1421 -61
rect 220 -72 224 -68
rect 328 -72 332 -68
rect 352 -72 356 -68
rect 1153 -72 1157 -68
rect 1261 -72 1265 -68
rect 1285 -72 1289 -68
rect 344 -79 348 -75
rect 328 -83 332 -79
rect 360 -83 364 -79
rect 1277 -79 1281 -75
rect 1261 -83 1265 -79
rect 1293 -83 1297 -79
rect 328 -90 332 -86
rect 360 -90 364 -86
rect 1013 -90 1017 -86
rect 1261 -90 1265 -86
rect 1293 -90 1297 -86
rect 1946 -90 1950 -86
rect 344 -97 348 -93
rect 484 -97 488 -93
rect 1277 -97 1281 -93
rect 1417 -97 1421 -93
rect 484 -105 488 -101
rect 1417 -105 1421 -101
rect 328 -109 332 -105
rect 360 -109 364 -105
rect 344 -113 348 -109
rect 1261 -109 1265 -105
rect 1293 -109 1297 -105
rect 1277 -113 1281 -109
rect 220 -120 224 -116
rect 328 -120 332 -116
rect 352 -120 356 -116
rect 1153 -120 1157 -116
rect 1261 -120 1265 -116
rect 1285 -120 1289 -116
rect 102 -127 106 -123
rect 138 -127 142 -123
rect 205 -127 209 -123
rect 234 -127 238 -123
rect 270 -127 274 -123
rect 337 -127 341 -123
rect 366 -127 370 -123
rect 402 -127 406 -123
rect 469 -127 473 -123
rect 553 -127 559 -123
rect 1035 -127 1039 -123
rect 1071 -127 1075 -123
rect 1138 -127 1142 -123
rect 1167 -127 1171 -123
rect 1203 -127 1207 -123
rect 1270 -127 1274 -123
rect 1299 -127 1303 -123
rect 1335 -127 1339 -123
rect 1402 -127 1406 -123
rect 1486 -127 1492 -123
rect 493 -134 499 -130
rect 1426 -134 1432 -130
rect 102 -141 106 -137
rect 152 -141 156 -137
rect 205 -141 209 -137
rect 234 -141 238 -137
rect 284 -141 288 -137
rect 337 -141 341 -137
rect 366 -141 370 -137
rect 416 -141 420 -137
rect 469 -141 473 -137
rect 1035 -141 1039 -137
rect 1085 -141 1089 -137
rect 1138 -141 1142 -137
rect 1167 -141 1171 -137
rect 1217 -141 1221 -137
rect 1270 -141 1274 -137
rect 1299 -141 1303 -137
rect 1349 -141 1353 -137
rect 1402 -141 1406 -137
rect 125 -152 129 -148
rect 96 -161 100 -157
rect 109 -158 113 -152
rect 146 -158 150 -152
rect 159 -156 163 -152
rect 183 -152 187 -148
rect 257 -152 261 -148
rect 167 -158 171 -152
rect 204 -158 208 -152
rect 220 -158 224 -152
rect 241 -158 245 -152
rect 278 -158 282 -152
rect 291 -156 295 -152
rect 315 -152 319 -148
rect 389 -152 393 -148
rect 299 -158 303 -152
rect 336 -158 340 -152
rect 352 -158 356 -152
rect 373 -158 377 -152
rect 410 -158 414 -152
rect 423 -156 427 -152
rect 447 -152 451 -148
rect 1058 -152 1062 -148
rect 431 -158 435 -152
rect 468 -158 472 -152
rect 484 -156 488 -152
rect 109 -171 113 -167
rect 125 -171 129 -165
rect 159 -165 163 -161
rect 146 -171 150 -167
rect 167 -171 171 -167
rect 183 -171 187 -165
rect 204 -171 208 -167
rect 220 -171 224 -167
rect 241 -171 245 -167
rect 257 -171 261 -165
rect 291 -165 295 -161
rect 278 -171 282 -167
rect 299 -171 303 -167
rect 315 -171 319 -165
rect 336 -171 340 -167
rect 352 -171 356 -167
rect 373 -171 377 -167
rect 389 -171 393 -165
rect 423 -165 427 -161
rect 410 -171 414 -167
rect 431 -171 435 -167
rect 447 -171 451 -165
rect 1029 -161 1033 -157
rect 1042 -158 1046 -152
rect 1079 -158 1083 -152
rect 1092 -156 1096 -152
rect 1116 -152 1120 -148
rect 1190 -152 1194 -148
rect 1100 -158 1104 -152
rect 1137 -158 1141 -152
rect 1153 -158 1157 -152
rect 1174 -158 1178 -152
rect 1211 -158 1215 -152
rect 1224 -156 1228 -152
rect 1248 -152 1252 -148
rect 1322 -152 1326 -148
rect 1232 -158 1236 -152
rect 1269 -158 1273 -152
rect 1285 -158 1289 -152
rect 1306 -158 1310 -152
rect 1343 -158 1347 -152
rect 1356 -156 1360 -152
rect 1380 -152 1384 -148
rect 1364 -158 1368 -152
rect 1401 -158 1405 -152
rect 1417 -156 1421 -152
rect 468 -171 472 -167
rect 484 -171 488 -167
rect 1042 -171 1046 -167
rect 1058 -171 1062 -165
rect 1092 -165 1096 -161
rect 1079 -171 1083 -167
rect 1100 -171 1104 -167
rect 1116 -171 1120 -165
rect 1137 -171 1141 -167
rect 1153 -171 1157 -167
rect 1174 -171 1178 -167
rect 1190 -171 1194 -165
rect 1224 -165 1228 -161
rect 1211 -171 1215 -167
rect 1232 -171 1236 -167
rect 1248 -171 1252 -165
rect 1269 -171 1273 -167
rect 1285 -171 1289 -167
rect 1306 -171 1310 -167
rect 1322 -171 1326 -165
rect 1356 -165 1360 -161
rect 1343 -171 1347 -167
rect 1364 -171 1368 -167
rect 1380 -171 1384 -165
rect 1401 -171 1405 -167
rect 1417 -171 1421 -167
rect 102 -182 106 -178
rect 139 -184 143 -180
rect 159 -184 163 -180
rect 203 -184 207 -180
rect 234 -182 238 -178
rect 271 -184 275 -180
rect 291 -184 295 -180
rect 335 -184 339 -180
rect 366 -182 370 -178
rect 403 -184 407 -180
rect 423 -184 427 -180
rect 467 -184 471 -180
rect 1035 -182 1039 -178
rect 1072 -184 1076 -180
rect 1092 -184 1096 -180
rect 1136 -184 1140 -180
rect 1167 -182 1171 -178
rect 1204 -184 1208 -180
rect 1224 -184 1228 -180
rect 1268 -184 1272 -180
rect 1299 -182 1303 -178
rect 1336 -184 1340 -180
rect 1356 -184 1360 -180
rect 1400 -184 1404 -180
rect 505 -191 511 -187
rect 1438 -191 1444 -187
rect 102 -198 106 -194
rect 153 -198 157 -194
rect 203 -198 207 -194
rect 234 -198 238 -194
rect 285 -198 289 -194
rect 335 -198 339 -194
rect 366 -198 370 -194
rect 417 -198 421 -194
rect 467 -198 471 -194
rect 541 -198 547 -194
rect 1035 -198 1039 -194
rect 1086 -198 1090 -194
rect 1136 -198 1140 -194
rect 1167 -198 1171 -194
rect 1218 -198 1222 -194
rect 1268 -198 1272 -194
rect 1299 -198 1303 -194
rect 1350 -198 1354 -194
rect 1400 -198 1404 -194
rect 1474 -198 1480 -194
<< metal2 >>
rect 219 1638 222 1687
rect 219 1594 222 1634
rect 227 1631 231 1774
rect 235 1711 238 1721
rect 242 1681 245 1690
rect 258 1683 261 1696
rect 271 1668 274 1721
rect 338 1711 341 1721
rect 278 1696 282 1700
rect 279 1681 282 1690
rect 234 1654 237 1666
rect 275 1664 276 1668
rect 285 1654 288 1707
rect 291 1687 294 1692
rect 300 1681 303 1690
rect 316 1683 319 1696
rect 337 1681 340 1690
rect 336 1654 339 1664
rect 219 1579 222 1588
rect 103 1209 106 1219
rect 110 1179 113 1188
rect 126 1181 129 1194
rect 139 1166 142 1219
rect 206 1209 209 1219
rect 146 1194 150 1198
rect 147 1179 150 1188
rect 102 1152 105 1164
rect 143 1162 144 1166
rect 153 1152 156 1205
rect 159 1185 162 1190
rect 168 1179 171 1188
rect 184 1181 187 1194
rect 205 1179 208 1188
rect 221 1179 224 1188
rect 204 1152 207 1162
rect 96 1049 99 1141
rect 221 1138 224 1175
rect 227 1131 231 1627
rect 344 1640 348 1774
rect 493 1751 499 1765
rect 493 1718 499 1747
rect 353 1688 356 1690
rect 353 1681 356 1684
rect 353 1647 356 1677
rect 493 1674 499 1714
rect 234 1609 237 1619
rect 235 1579 238 1588
rect 256 1581 259 1594
rect 272 1579 275 1588
rect 281 1585 284 1590
rect 236 1552 239 1562
rect 287 1552 290 1605
rect 293 1594 297 1598
rect 293 1579 296 1588
rect 301 1566 304 1619
rect 337 1609 340 1619
rect 314 1581 317 1594
rect 330 1579 333 1588
rect 299 1562 300 1566
rect 338 1552 341 1564
rect 235 1209 238 1219
rect 242 1179 245 1188
rect 258 1181 261 1194
rect 271 1166 274 1219
rect 338 1209 341 1219
rect 278 1194 282 1198
rect 279 1179 282 1188
rect 234 1152 237 1164
rect 275 1162 276 1166
rect 285 1152 288 1205
rect 291 1185 294 1190
rect 300 1179 303 1188
rect 316 1181 319 1194
rect 337 1179 340 1188
rect 336 1152 339 1162
rect 211 1120 215 1123
rect 211 1101 215 1116
rect 227 1113 231 1127
rect 243 1127 247 1131
rect 243 1120 247 1123
rect 243 1101 247 1116
rect 227 1097 231 1098
rect 243 1093 247 1097
rect 103 1069 106 1079
rect 110 1039 113 1048
rect 126 1041 129 1054
rect 139 1026 142 1079
rect 206 1069 209 1079
rect 146 1054 150 1058
rect 147 1039 150 1048
rect 102 1012 105 1024
rect 143 1022 144 1026
rect 153 1012 156 1065
rect 221 1054 224 1086
rect 159 1045 162 1050
rect 168 1039 171 1048
rect 184 1041 187 1054
rect 205 1039 208 1048
rect 221 1039 224 1048
rect 204 1012 207 1022
rect 96 963 99 1001
rect 103 983 106 993
rect 110 953 113 962
rect 126 955 129 968
rect 139 940 142 993
rect 206 983 209 993
rect 146 968 150 972
rect 147 953 150 962
rect 102 926 105 938
rect 143 936 144 940
rect 153 926 156 979
rect 159 959 162 964
rect 168 953 171 962
rect 184 955 187 968
rect 205 953 208 962
rect 221 953 224 962
rect 204 926 207 936
rect 96 823 99 915
rect 221 912 224 949
rect 103 843 106 853
rect 110 813 113 822
rect 126 815 129 828
rect 139 800 142 853
rect 206 843 209 853
rect 146 828 150 832
rect 147 813 150 822
rect 102 786 105 798
rect 143 796 144 800
rect 153 786 156 839
rect 221 828 224 860
rect 159 819 162 824
rect 168 813 171 822
rect 184 815 187 828
rect 205 813 208 822
rect 221 813 224 822
rect 204 786 207 796
rect 219 658 222 707
rect 219 614 222 654
rect 227 651 231 1093
rect 235 1069 238 1079
rect 242 1039 245 1048
rect 258 1041 261 1054
rect 271 1026 274 1079
rect 338 1069 341 1079
rect 278 1054 282 1058
rect 279 1039 282 1048
rect 234 1012 237 1024
rect 275 1022 276 1026
rect 285 1012 288 1065
rect 291 1045 294 1050
rect 300 1039 303 1048
rect 316 1041 319 1054
rect 337 1039 340 1048
rect 336 1012 339 1022
rect 235 983 238 993
rect 242 953 245 962
rect 258 955 261 968
rect 271 940 274 993
rect 338 983 341 993
rect 278 968 282 972
rect 279 953 282 962
rect 234 926 237 938
rect 275 936 276 940
rect 285 926 288 979
rect 291 959 294 964
rect 300 953 303 962
rect 316 955 319 968
rect 337 953 340 962
rect 336 926 339 936
rect 344 905 348 1636
rect 368 1631 372 1636
rect 493 1616 499 1670
rect 493 1542 499 1612
rect 493 1410 499 1538
rect 493 1278 499 1406
rect 367 1209 370 1219
rect 353 1179 356 1188
rect 374 1179 377 1188
rect 390 1181 393 1194
rect 353 1138 356 1175
rect 403 1166 406 1219
rect 470 1209 473 1219
rect 493 1216 499 1274
rect 410 1194 414 1198
rect 411 1179 414 1188
rect 366 1152 369 1164
rect 407 1162 408 1166
rect 417 1152 420 1205
rect 423 1185 426 1190
rect 432 1179 435 1188
rect 448 1181 451 1194
rect 469 1179 472 1188
rect 485 1179 488 1190
rect 468 1152 471 1162
rect 485 1145 488 1175
rect 485 1113 488 1141
rect 493 1146 499 1212
rect 493 1106 499 1142
rect 353 1054 356 1086
rect 367 1069 370 1079
rect 353 1039 356 1048
rect 374 1039 377 1048
rect 390 1041 393 1054
rect 403 1026 406 1079
rect 470 1069 473 1079
rect 410 1054 414 1058
rect 411 1039 414 1048
rect 366 1012 369 1024
rect 407 1022 408 1026
rect 417 1012 420 1065
rect 485 1054 488 1101
rect 423 1045 426 1050
rect 432 1039 435 1048
rect 448 1041 451 1054
rect 469 1039 472 1048
rect 485 1039 488 1050
rect 468 1012 471 1022
rect 485 1005 488 1035
rect 493 1076 499 1102
rect 367 983 370 993
rect 353 953 356 962
rect 374 953 377 962
rect 390 955 393 968
rect 353 912 356 949
rect 403 940 406 993
rect 470 983 473 993
rect 493 990 499 1072
rect 410 968 414 972
rect 411 953 414 962
rect 366 926 369 938
rect 407 936 408 940
rect 417 926 420 979
rect 423 959 426 964
rect 432 953 435 962
rect 448 955 451 968
rect 469 953 472 962
rect 485 953 488 964
rect 468 926 471 936
rect 485 919 488 949
rect 328 894 332 897
rect 328 875 332 890
rect 344 887 348 901
rect 360 901 364 905
rect 360 894 364 897
rect 360 875 364 890
rect 485 887 488 915
rect 344 871 348 872
rect 360 867 364 871
rect 235 843 238 853
rect 242 813 245 822
rect 258 815 261 828
rect 271 800 274 853
rect 338 843 341 853
rect 278 828 282 832
rect 279 813 282 822
rect 234 786 237 798
rect 275 796 276 800
rect 285 786 288 839
rect 291 819 294 824
rect 300 813 303 822
rect 316 815 319 828
rect 337 813 340 822
rect 336 786 339 796
rect 235 731 238 741
rect 242 701 245 710
rect 258 703 261 716
rect 271 688 274 741
rect 338 731 341 741
rect 278 716 282 720
rect 279 701 282 710
rect 234 674 237 686
rect 275 684 276 688
rect 285 674 288 727
rect 291 707 294 712
rect 300 701 303 710
rect 316 703 319 716
rect 337 701 340 710
rect 336 674 339 684
rect 219 599 222 608
rect 103 229 106 239
rect 110 199 113 208
rect 126 201 129 214
rect 139 186 142 239
rect 206 229 209 239
rect 146 214 150 218
rect 147 199 150 208
rect 102 172 105 184
rect 143 182 144 186
rect 153 172 156 225
rect 159 205 162 210
rect 168 199 171 208
rect 184 201 187 214
rect 205 199 208 208
rect 221 199 224 208
rect 204 172 207 182
rect 96 69 99 161
rect 221 158 224 195
rect 227 151 231 647
rect 344 660 348 867
rect 353 828 356 860
rect 367 843 370 853
rect 353 813 356 822
rect 374 813 377 822
rect 390 815 393 828
rect 403 800 406 853
rect 470 843 473 853
rect 410 828 414 832
rect 411 813 414 822
rect 366 786 369 798
rect 407 796 408 800
rect 417 786 420 839
rect 485 828 488 875
rect 423 819 426 824
rect 432 813 435 822
rect 448 815 451 828
rect 469 813 472 822
rect 485 820 488 824
rect 493 850 499 986
rect 485 813 488 816
rect 468 786 471 796
rect 493 771 499 846
rect 493 738 499 767
rect 353 708 356 710
rect 353 701 356 704
rect 353 667 356 697
rect 493 694 499 734
rect 234 629 237 639
rect 235 599 238 608
rect 256 601 259 614
rect 272 599 275 608
rect 281 605 284 610
rect 236 572 239 582
rect 287 572 290 625
rect 293 614 297 618
rect 293 599 296 608
rect 301 586 304 639
rect 337 629 340 639
rect 314 601 317 614
rect 330 599 333 608
rect 299 582 300 586
rect 338 572 341 584
rect 235 229 238 239
rect 242 199 245 208
rect 258 201 261 214
rect 271 186 274 239
rect 338 229 341 239
rect 278 214 282 218
rect 279 199 282 208
rect 234 172 237 184
rect 275 182 276 186
rect 285 172 288 225
rect 291 205 294 210
rect 300 199 303 208
rect 316 201 319 214
rect 337 199 340 208
rect 336 172 339 182
rect 211 140 215 143
rect 211 121 215 136
rect 227 133 231 147
rect 243 147 247 151
rect 243 140 247 143
rect 243 121 247 136
rect 227 117 231 118
rect 243 113 247 117
rect 103 89 106 99
rect 110 59 113 68
rect 126 61 129 74
rect 139 46 142 99
rect 206 89 209 99
rect 146 74 150 78
rect 147 59 150 68
rect 102 32 105 44
rect 143 42 144 46
rect 153 32 156 85
rect 221 74 224 106
rect 159 65 162 70
rect 168 59 171 68
rect 184 61 187 74
rect 205 59 208 68
rect 221 59 224 68
rect 204 32 207 42
rect 96 -17 99 21
rect 103 3 106 13
rect 110 -27 113 -18
rect 126 -25 129 -12
rect 139 -40 142 13
rect 206 3 209 13
rect 146 -12 150 -8
rect 147 -27 150 -18
rect 102 -54 105 -42
rect 143 -44 144 -40
rect 153 -54 156 -1
rect 159 -21 162 -16
rect 168 -27 171 -18
rect 184 -25 187 -12
rect 205 -27 208 -18
rect 221 -27 224 -18
rect 204 -54 207 -44
rect 96 -157 99 -65
rect 221 -68 224 -31
rect 103 -137 106 -127
rect 110 -167 113 -158
rect 126 -165 129 -152
rect 139 -180 142 -127
rect 206 -137 209 -127
rect 146 -152 150 -148
rect 147 -167 150 -158
rect 102 -194 105 -182
rect 143 -184 144 -180
rect 153 -194 156 -141
rect 221 -152 224 -120
rect 159 -161 162 -156
rect 168 -167 171 -158
rect 184 -165 187 -152
rect 205 -167 208 -158
rect 221 -167 224 -158
rect 204 -194 207 -184
rect 227 -208 231 113
rect 235 89 238 99
rect 242 59 245 68
rect 258 61 261 74
rect 271 46 274 99
rect 338 89 341 99
rect 278 74 282 78
rect 279 59 282 68
rect 234 32 237 44
rect 275 42 276 46
rect 285 32 288 85
rect 291 65 294 70
rect 300 59 303 68
rect 316 61 319 74
rect 337 59 340 68
rect 336 32 339 42
rect 235 3 238 13
rect 242 -27 245 -18
rect 258 -25 261 -12
rect 271 -40 274 13
rect 338 3 341 13
rect 278 -12 282 -8
rect 279 -27 282 -18
rect 234 -54 237 -42
rect 275 -44 276 -40
rect 285 -54 288 -1
rect 291 -21 294 -16
rect 300 -27 303 -18
rect 316 -25 319 -12
rect 337 -27 340 -18
rect 336 -54 339 -44
rect 344 -75 348 656
rect 368 651 372 656
rect 493 636 499 690
rect 493 562 499 632
rect 493 430 499 558
rect 493 298 499 426
rect 367 229 370 239
rect 353 199 356 208
rect 374 199 377 208
rect 390 201 393 214
rect 353 158 356 195
rect 403 186 406 239
rect 470 229 473 239
rect 493 236 499 294
rect 410 214 414 218
rect 411 199 414 208
rect 366 172 369 184
rect 407 182 408 186
rect 417 172 420 225
rect 423 205 426 210
rect 432 199 435 208
rect 448 201 451 214
rect 469 199 472 208
rect 485 199 488 210
rect 468 172 471 182
rect 485 165 488 195
rect 485 133 488 161
rect 493 166 499 232
rect 493 126 499 162
rect 353 74 356 106
rect 367 89 370 99
rect 353 59 356 68
rect 374 59 377 68
rect 390 61 393 74
rect 403 46 406 99
rect 470 89 473 99
rect 410 74 414 78
rect 411 59 414 68
rect 366 32 369 44
rect 407 42 408 46
rect 417 32 420 85
rect 485 74 488 121
rect 423 65 426 70
rect 432 59 435 68
rect 448 61 451 74
rect 469 59 472 68
rect 485 59 488 70
rect 468 32 471 42
rect 485 25 488 55
rect 493 96 499 122
rect 367 3 370 13
rect 353 -27 356 -18
rect 374 -27 377 -18
rect 390 -25 393 -12
rect 353 -68 356 -31
rect 403 -40 406 13
rect 470 3 473 13
rect 493 10 499 92
rect 410 -12 414 -8
rect 411 -27 414 -18
rect 366 -54 369 -42
rect 407 -44 408 -40
rect 417 -54 420 -1
rect 423 -21 426 -16
rect 432 -27 435 -18
rect 448 -25 451 -12
rect 469 -27 472 -18
rect 485 -27 488 -16
rect 468 -54 471 -44
rect 485 -61 488 -31
rect 328 -86 332 -83
rect 328 -105 332 -90
rect 344 -93 348 -79
rect 360 -79 364 -75
rect 360 -86 364 -83
rect 360 -105 364 -90
rect 485 -93 488 -65
rect 344 -109 348 -108
rect 360 -113 364 -109
rect 235 -137 238 -127
rect 242 -167 245 -158
rect 258 -165 261 -152
rect 271 -180 274 -127
rect 338 -137 341 -127
rect 278 -152 282 -148
rect 279 -167 282 -158
rect 234 -194 237 -182
rect 275 -184 276 -180
rect 285 -194 288 -141
rect 291 -161 294 -156
rect 300 -167 303 -158
rect 316 -165 319 -152
rect 337 -167 340 -158
rect 336 -194 339 -184
rect 344 -208 348 -113
rect 353 -152 356 -120
rect 367 -137 370 -127
rect 353 -167 356 -158
rect 374 -167 377 -158
rect 390 -165 393 -152
rect 403 -180 406 -127
rect 470 -137 473 -127
rect 410 -152 414 -148
rect 411 -167 414 -158
rect 366 -194 369 -182
rect 407 -184 408 -180
rect 417 -194 420 -141
rect 485 -152 488 -105
rect 423 -161 426 -156
rect 432 -167 435 -158
rect 448 -165 451 -152
rect 469 -167 472 -158
rect 485 -160 488 -156
rect 493 -130 499 6
rect 485 -167 488 -164
rect 468 -194 471 -184
rect 493 -208 499 -134
rect 505 1694 511 1765
rect 505 1661 511 1690
rect 505 1608 511 1657
rect 505 1559 511 1604
rect 505 1476 511 1555
rect 505 1344 511 1472
rect 505 1212 511 1340
rect 505 1159 511 1208
rect 505 1049 511 1155
rect 505 1019 511 1045
rect 505 963 511 1015
rect 505 933 511 959
rect 505 793 511 929
rect 505 714 511 789
rect 505 681 511 710
rect 505 628 511 677
rect 505 579 511 624
rect 505 496 511 575
rect 505 364 511 492
rect 505 232 511 360
rect 505 179 511 228
rect 505 69 511 175
rect 505 39 511 65
rect 505 -17 511 35
rect 505 -47 511 -21
rect 505 -187 511 -51
rect 505 -208 511 -191
rect 517 1615 523 1765
rect 517 1601 523 1611
rect 517 1483 523 1597
rect 517 1469 523 1479
rect 517 1351 523 1465
rect 517 1337 523 1347
rect 517 1205 523 1333
rect 517 1131 523 1201
rect 517 635 523 1127
rect 517 621 523 631
rect 517 503 523 617
rect 517 489 523 499
rect 517 371 523 485
rect 517 357 523 367
rect 517 225 523 353
rect 517 151 523 221
rect 517 -208 523 147
rect 529 1667 535 1765
rect 529 1535 535 1663
rect 529 1417 535 1531
rect 529 1403 535 1413
rect 529 1285 535 1399
rect 529 1271 535 1281
rect 529 1139 535 1267
rect 529 687 535 1135
rect 529 555 535 683
rect 529 437 535 551
rect 529 423 535 433
rect 529 305 535 419
rect 529 291 535 301
rect 529 159 535 287
rect 529 -208 535 155
rect 541 1687 547 1765
rect 541 1654 547 1683
rect 541 1552 547 1650
rect 541 1153 547 1548
rect 541 1042 547 1149
rect 541 1012 547 1038
rect 541 956 547 1008
rect 541 926 547 952
rect 541 786 547 922
rect 541 707 547 782
rect 541 674 547 703
rect 541 572 547 670
rect 541 173 547 568
rect 541 62 547 169
rect 541 32 547 58
rect 541 -24 547 28
rect 541 -54 547 -28
rect 541 -194 547 -58
rect 541 -208 547 -198
rect 553 1758 559 1765
rect 553 1725 559 1754
rect 575 1744 578 1754
rect 553 1623 559 1721
rect 582 1714 585 1723
rect 598 1716 601 1729
rect 611 1701 614 1754
rect 678 1744 681 1754
rect 707 1744 710 1754
rect 618 1729 622 1733
rect 619 1714 622 1723
rect 574 1687 577 1699
rect 615 1697 616 1701
rect 625 1687 628 1740
rect 631 1720 634 1725
rect 640 1714 643 1723
rect 656 1716 659 1729
rect 677 1714 680 1723
rect 693 1723 696 1725
rect 693 1720 700 1723
rect 693 1714 696 1720
rect 714 1714 717 1723
rect 730 1716 733 1729
rect 676 1687 679 1697
rect 693 1680 696 1710
rect 743 1701 746 1754
rect 810 1744 813 1754
rect 839 1744 842 1754
rect 750 1729 754 1733
rect 751 1714 754 1723
rect 706 1687 709 1699
rect 747 1697 748 1701
rect 757 1687 760 1740
rect 763 1720 766 1725
rect 772 1714 775 1723
rect 788 1716 791 1729
rect 809 1714 812 1723
rect 825 1723 828 1725
rect 825 1720 832 1723
rect 825 1714 828 1720
rect 846 1714 849 1723
rect 862 1716 865 1729
rect 808 1687 811 1697
rect 693 1677 745 1680
rect 573 1657 576 1670
rect 599 1660 602 1663
rect 606 1657 609 1670
rect 623 1657 626 1670
rect 553 1223 559 1619
rect 573 1608 576 1623
rect 587 1615 590 1619
rect 605 1608 608 1623
rect 624 1608 627 1623
rect 630 1622 633 1663
rect 646 1615 649 1656
rect 652 1623 655 1663
rect 671 1615 674 1656
rect 680 1657 683 1670
rect 696 1657 699 1670
rect 717 1660 720 1663
rect 724 1657 727 1670
rect 742 1666 745 1677
rect 825 1674 828 1710
rect 875 1701 878 1754
rect 942 1744 945 1754
rect 971 1744 974 1754
rect 882 1729 886 1733
rect 883 1714 886 1723
rect 838 1687 841 1699
rect 879 1697 880 1701
rect 889 1687 892 1740
rect 895 1720 898 1725
rect 904 1714 907 1723
rect 920 1716 923 1729
rect 941 1714 944 1723
rect 957 1723 960 1725
rect 957 1720 964 1723
rect 957 1714 960 1720
rect 978 1714 981 1723
rect 994 1716 997 1729
rect 940 1687 943 1697
rect 957 1680 960 1702
rect 1007 1701 1010 1754
rect 1074 1744 1077 1754
rect 1014 1729 1018 1733
rect 1015 1714 1018 1723
rect 970 1687 973 1699
rect 1011 1697 1012 1701
rect 1021 1687 1024 1740
rect 1027 1720 1030 1725
rect 1036 1714 1039 1723
rect 1052 1716 1055 1729
rect 1073 1714 1076 1723
rect 1089 1723 1092 1725
rect 1089 1720 1093 1723
rect 1089 1714 1092 1720
rect 1089 1706 1092 1710
rect 1072 1687 1075 1697
rect 823 1669 828 1674
rect 885 1676 960 1680
rect 742 1663 787 1666
rect 742 1653 745 1663
rect 760 1650 780 1653
rect 777 1631 780 1650
rect 680 1608 683 1623
rect 695 1608 698 1623
rect 702 1615 706 1618
rect 723 1608 726 1623
rect 573 1589 576 1604
rect 587 1593 590 1597
rect 605 1589 608 1604
rect 624 1589 627 1604
rect 573 1542 576 1555
rect 599 1549 602 1552
rect 573 1525 576 1538
rect 583 1535 587 1545
rect 606 1542 609 1555
rect 623 1542 626 1555
rect 630 1549 633 1590
rect 646 1556 649 1597
rect 652 1549 655 1589
rect 671 1556 674 1597
rect 680 1589 683 1604
rect 695 1589 698 1604
rect 702 1594 706 1597
rect 723 1589 726 1604
rect 680 1542 683 1555
rect 599 1528 602 1531
rect 606 1525 609 1538
rect 623 1525 626 1538
rect 573 1476 576 1491
rect 587 1483 590 1487
rect 605 1476 608 1491
rect 624 1476 627 1491
rect 630 1490 633 1531
rect 646 1483 649 1524
rect 652 1491 655 1531
rect 671 1483 674 1524
rect 680 1525 683 1538
rect 696 1542 699 1555
rect 717 1549 720 1552
rect 724 1542 727 1555
rect 777 1555 780 1627
rect 788 1591 791 1663
rect 823 1666 826 1669
rect 823 1663 868 1666
rect 823 1653 826 1663
rect 696 1525 699 1538
rect 717 1528 720 1531
rect 724 1525 727 1538
rect 777 1521 780 1551
rect 788 1535 791 1587
rect 795 1575 799 1641
rect 783 1531 787 1534
rect 776 1518 780 1521
rect 777 1499 780 1518
rect 680 1476 683 1491
rect 695 1476 698 1491
rect 702 1483 706 1486
rect 723 1476 726 1491
rect 573 1457 576 1472
rect 587 1461 590 1465
rect 605 1457 608 1472
rect 624 1457 627 1472
rect 573 1410 576 1423
rect 599 1417 602 1420
rect 573 1393 576 1406
rect 606 1410 609 1423
rect 623 1410 626 1423
rect 630 1417 633 1458
rect 646 1424 649 1465
rect 652 1417 655 1457
rect 671 1424 674 1465
rect 680 1457 683 1472
rect 695 1457 698 1472
rect 702 1462 706 1465
rect 723 1457 726 1472
rect 680 1410 683 1423
rect 599 1396 602 1399
rect 606 1393 609 1406
rect 623 1393 626 1406
rect 573 1344 576 1359
rect 587 1351 590 1355
rect 605 1344 608 1359
rect 624 1344 627 1359
rect 630 1358 633 1399
rect 646 1351 649 1392
rect 652 1359 655 1399
rect 671 1351 674 1392
rect 680 1393 683 1406
rect 696 1410 699 1423
rect 717 1417 720 1420
rect 724 1410 727 1423
rect 777 1424 780 1495
rect 788 1460 791 1531
rect 696 1393 699 1406
rect 717 1396 720 1399
rect 724 1393 727 1406
rect 777 1367 780 1420
rect 788 1403 791 1456
rect 795 1444 799 1509
rect 783 1399 787 1402
rect 826 1402 829 1653
rect 841 1650 861 1653
rect 858 1631 861 1650
rect 858 1555 861 1627
rect 869 1591 872 1663
rect 876 1575 880 1641
rect 885 1542 888 1676
rect 1089 1673 1092 1702
rect 913 1670 1020 1673
rect 847 1538 888 1542
rect 847 1534 850 1538
rect 847 1531 892 1534
rect 847 1521 850 1531
rect 865 1518 885 1521
rect 847 1516 850 1517
rect 882 1499 885 1518
rect 882 1424 885 1495
rect 893 1460 896 1531
rect 900 1444 904 1509
rect 680 1344 683 1359
rect 695 1344 698 1359
rect 702 1351 706 1354
rect 723 1344 726 1359
rect 573 1325 576 1340
rect 587 1329 590 1333
rect 605 1325 608 1340
rect 624 1325 627 1340
rect 573 1278 576 1291
rect 599 1285 602 1288
rect 573 1261 576 1274
rect 606 1278 609 1291
rect 623 1278 626 1291
rect 630 1285 633 1326
rect 646 1292 649 1333
rect 652 1285 655 1325
rect 671 1292 674 1333
rect 680 1325 683 1340
rect 695 1325 698 1340
rect 702 1330 706 1333
rect 723 1325 726 1340
rect 680 1278 683 1291
rect 599 1264 602 1267
rect 606 1261 609 1274
rect 623 1261 626 1274
rect 553 1113 559 1219
rect 573 1212 576 1227
rect 587 1219 590 1223
rect 573 1193 576 1208
rect 596 1205 600 1215
rect 605 1212 608 1227
rect 624 1212 627 1227
rect 630 1226 633 1267
rect 646 1219 649 1260
rect 652 1227 655 1267
rect 671 1219 674 1260
rect 680 1261 683 1274
rect 696 1278 699 1291
rect 717 1285 720 1288
rect 724 1278 727 1291
rect 777 1289 780 1363
rect 788 1325 791 1399
rect 823 1399 868 1402
rect 823 1389 826 1399
rect 841 1386 861 1389
rect 696 1261 699 1274
rect 717 1264 720 1267
rect 724 1261 727 1274
rect 777 1235 780 1285
rect 788 1271 791 1321
rect 795 1309 799 1377
rect 858 1367 861 1386
rect 858 1289 861 1363
rect 869 1325 872 1399
rect 913 1402 916 1670
rect 1024 1670 1092 1673
rect 1152 1638 1155 1687
rect 1152 1594 1155 1634
rect 1160 1631 1164 1774
rect 1168 1711 1171 1721
rect 1175 1681 1178 1690
rect 1191 1683 1194 1696
rect 1204 1668 1207 1721
rect 1271 1711 1274 1721
rect 1211 1696 1215 1700
rect 1212 1681 1215 1690
rect 1167 1654 1170 1666
rect 1208 1664 1209 1668
rect 1218 1654 1221 1707
rect 1224 1687 1227 1692
rect 1233 1681 1236 1690
rect 1249 1683 1252 1696
rect 1270 1681 1273 1690
rect 1269 1654 1272 1664
rect 1152 1579 1155 1588
rect 913 1399 958 1402
rect 913 1389 916 1399
rect 931 1386 951 1389
rect 876 1309 880 1377
rect 948 1367 951 1386
rect 948 1289 951 1363
rect 959 1325 962 1399
rect 966 1309 970 1377
rect 783 1267 787 1270
rect 680 1212 683 1227
rect 695 1212 698 1227
rect 702 1219 706 1222
rect 723 1212 726 1227
rect 587 1197 590 1201
rect 605 1193 608 1208
rect 624 1193 627 1208
rect 573 1146 576 1159
rect 599 1153 602 1156
rect 581 1139 585 1149
rect 606 1146 609 1159
rect 623 1146 626 1159
rect 630 1153 633 1194
rect 646 1160 649 1201
rect 652 1153 655 1193
rect 671 1160 674 1201
rect 680 1193 683 1208
rect 695 1193 698 1208
rect 702 1198 706 1201
rect 723 1193 726 1208
rect 680 1146 683 1159
rect 696 1146 699 1159
rect 717 1153 720 1156
rect 724 1146 727 1159
rect 777 1153 780 1231
rect 788 1189 791 1267
rect 795 1173 799 1245
rect 807 1146 811 1159
rect 816 1139 819 1149
rect 826 1132 829 1201
rect 848 1197 851 1201
rect 866 1193 869 1208
rect 885 1193 888 1208
rect 833 1146 837 1159
rect 860 1153 863 1156
rect 867 1146 870 1159
rect 884 1146 887 1159
rect 891 1153 894 1194
rect 907 1160 910 1201
rect 913 1153 916 1193
rect 932 1160 935 1201
rect 941 1193 944 1208
rect 956 1193 959 1208
rect 963 1198 967 1201
rect 984 1193 987 1208
rect 941 1146 944 1159
rect 957 1146 960 1159
rect 978 1153 981 1156
rect 985 1146 988 1159
rect 1001 1140 1005 1376
rect 1036 1209 1039 1219
rect 1043 1179 1046 1188
rect 1059 1181 1062 1194
rect 1072 1166 1075 1219
rect 1139 1209 1142 1219
rect 1079 1194 1083 1198
rect 1080 1179 1083 1188
rect 1035 1152 1038 1164
rect 1076 1162 1077 1166
rect 1086 1152 1089 1205
rect 1092 1185 1095 1190
rect 1101 1179 1104 1188
rect 1117 1181 1120 1194
rect 1138 1179 1141 1188
rect 1154 1179 1157 1188
rect 1137 1152 1140 1162
rect 994 1128 995 1131
rect 553 1083 559 1109
rect 553 1027 559 1079
rect 553 997 559 1023
rect 859 1020 863 1102
rect 874 1099 877 1109
rect 881 1069 884 1078
rect 897 1071 900 1084
rect 910 1056 913 1109
rect 977 1099 980 1109
rect 917 1084 921 1088
rect 918 1069 921 1078
rect 873 1042 876 1054
rect 914 1052 915 1056
rect 924 1042 927 1095
rect 992 1084 995 1128
rect 930 1075 933 1080
rect 939 1069 942 1078
rect 955 1071 958 1084
rect 976 1069 979 1078
rect 992 1069 995 1078
rect 975 1042 978 1052
rect 992 1035 995 1065
rect 553 857 559 993
rect 867 993 870 1030
rect 874 1013 877 1023
rect 881 983 884 992
rect 897 985 900 998
rect 910 970 913 1023
rect 977 1013 980 1023
rect 917 998 921 1002
rect 918 983 921 992
rect 873 956 876 968
rect 914 966 915 970
rect 924 956 927 1009
rect 930 989 933 994
rect 939 983 942 992
rect 955 985 958 998
rect 976 983 979 992
rect 992 993 995 994
rect 1013 996 1017 1136
rect 1029 1049 1032 1141
rect 1154 1138 1157 1175
rect 1160 1131 1164 1627
rect 1277 1640 1281 1774
rect 1426 1751 1432 1765
rect 1426 1718 1432 1747
rect 1286 1688 1289 1690
rect 1286 1681 1289 1684
rect 1286 1647 1289 1677
rect 1426 1674 1432 1714
rect 1167 1609 1170 1619
rect 1168 1579 1171 1588
rect 1189 1581 1192 1594
rect 1205 1579 1208 1588
rect 1214 1585 1217 1590
rect 1169 1552 1172 1562
rect 1220 1552 1223 1605
rect 1226 1594 1230 1598
rect 1226 1579 1229 1588
rect 1234 1566 1237 1619
rect 1270 1609 1273 1619
rect 1247 1581 1250 1594
rect 1263 1579 1266 1588
rect 1232 1562 1233 1566
rect 1271 1552 1274 1564
rect 1168 1209 1171 1219
rect 1175 1179 1178 1188
rect 1191 1181 1194 1194
rect 1204 1166 1207 1219
rect 1271 1209 1274 1219
rect 1211 1194 1215 1198
rect 1212 1179 1215 1188
rect 1167 1152 1170 1164
rect 1208 1162 1209 1166
rect 1218 1152 1221 1205
rect 1224 1185 1227 1190
rect 1233 1179 1236 1188
rect 1249 1181 1252 1194
rect 1270 1179 1273 1188
rect 1269 1152 1272 1162
rect 1144 1120 1148 1123
rect 1144 1101 1148 1116
rect 1160 1113 1164 1127
rect 1176 1127 1180 1131
rect 1176 1120 1180 1123
rect 1176 1101 1180 1116
rect 1160 1097 1164 1098
rect 1176 1093 1180 1097
rect 1036 1069 1039 1079
rect 1043 1039 1046 1048
rect 1059 1041 1062 1054
rect 1072 1026 1075 1079
rect 1139 1069 1142 1079
rect 1079 1054 1083 1058
rect 1080 1039 1083 1048
rect 1035 1012 1038 1024
rect 1076 1022 1077 1026
rect 1086 1012 1089 1065
rect 1154 1054 1157 1086
rect 1092 1045 1095 1050
rect 1101 1039 1104 1048
rect 1117 1041 1120 1054
rect 1138 1039 1141 1048
rect 1154 1039 1157 1048
rect 1137 1012 1140 1022
rect 992 988 995 989
rect 975 956 978 966
rect 1013 894 1017 976
rect 1029 963 1032 1001
rect 1036 983 1039 993
rect 1043 953 1046 962
rect 1059 955 1062 968
rect 1072 940 1075 993
rect 1139 983 1142 993
rect 1079 968 1083 972
rect 1080 953 1083 962
rect 1035 926 1038 938
rect 1076 936 1077 940
rect 1086 926 1089 979
rect 1092 959 1095 964
rect 1101 953 1104 962
rect 1117 955 1120 968
rect 1138 953 1141 962
rect 1154 953 1157 962
rect 1137 926 1140 936
rect 553 778 559 853
rect 1029 823 1032 915
rect 1154 912 1157 949
rect 1036 843 1039 853
rect 1043 813 1046 822
rect 1059 815 1062 828
rect 1072 800 1075 853
rect 1139 843 1142 853
rect 1079 828 1083 832
rect 1080 813 1083 822
rect 1035 786 1038 798
rect 1076 796 1077 800
rect 1086 786 1089 839
rect 1154 828 1157 860
rect 1092 819 1095 824
rect 1101 813 1104 822
rect 1117 815 1120 828
rect 1138 813 1141 822
rect 1154 813 1157 822
rect 1137 786 1140 796
rect 553 745 559 774
rect 575 764 578 774
rect 553 643 559 741
rect 582 734 585 743
rect 598 736 601 749
rect 611 721 614 774
rect 678 764 681 774
rect 707 764 710 774
rect 618 749 622 753
rect 619 734 622 743
rect 574 707 577 719
rect 615 717 616 721
rect 625 707 628 760
rect 631 740 634 745
rect 640 734 643 743
rect 656 736 659 749
rect 677 734 680 743
rect 693 743 696 745
rect 693 740 700 743
rect 693 734 696 740
rect 714 734 717 743
rect 730 736 733 749
rect 676 707 679 717
rect 693 700 696 730
rect 743 721 746 774
rect 810 764 813 774
rect 839 764 842 774
rect 750 749 754 753
rect 751 734 754 743
rect 706 707 709 719
rect 747 717 748 721
rect 757 707 760 760
rect 763 740 766 745
rect 772 734 775 743
rect 788 736 791 749
rect 809 734 812 743
rect 825 743 828 745
rect 825 740 832 743
rect 825 734 828 740
rect 846 734 849 743
rect 862 736 865 749
rect 808 707 811 717
rect 693 697 745 700
rect 573 677 576 690
rect 599 680 602 683
rect 606 677 609 690
rect 623 677 626 690
rect 553 243 559 639
rect 573 628 576 643
rect 587 635 590 639
rect 605 628 608 643
rect 624 628 627 643
rect 630 642 633 683
rect 646 635 649 676
rect 652 643 655 683
rect 671 635 674 676
rect 680 677 683 690
rect 696 677 699 690
rect 717 680 720 683
rect 724 677 727 690
rect 742 686 745 697
rect 825 694 828 730
rect 875 721 878 774
rect 942 764 945 774
rect 971 764 974 774
rect 882 749 886 753
rect 883 734 886 743
rect 838 707 841 719
rect 879 717 880 721
rect 889 707 892 760
rect 895 740 898 745
rect 904 734 907 743
rect 920 736 923 749
rect 941 734 944 743
rect 957 743 960 745
rect 957 740 964 743
rect 957 734 960 740
rect 978 734 981 743
rect 994 736 997 749
rect 940 707 943 717
rect 957 700 960 722
rect 1007 721 1010 774
rect 1074 764 1077 774
rect 1014 749 1018 753
rect 1015 734 1018 743
rect 970 707 973 719
rect 1011 717 1012 721
rect 1021 707 1024 760
rect 1027 740 1030 745
rect 1036 734 1039 743
rect 1052 736 1055 749
rect 1073 734 1076 743
rect 1089 743 1092 745
rect 1089 740 1093 743
rect 1089 734 1092 740
rect 1089 726 1092 730
rect 1072 707 1075 717
rect 823 689 828 694
rect 885 696 960 700
rect 742 683 787 686
rect 742 673 745 683
rect 760 670 780 673
rect 777 651 780 670
rect 680 628 683 643
rect 695 628 698 643
rect 702 635 706 638
rect 723 628 726 643
rect 573 609 576 624
rect 587 613 590 617
rect 605 609 608 624
rect 624 609 627 624
rect 573 562 576 575
rect 599 569 602 572
rect 573 545 576 558
rect 583 555 587 565
rect 606 562 609 575
rect 623 562 626 575
rect 630 569 633 610
rect 646 576 649 617
rect 652 569 655 609
rect 671 576 674 617
rect 680 609 683 624
rect 695 609 698 624
rect 702 614 706 617
rect 723 609 726 624
rect 680 562 683 575
rect 599 548 602 551
rect 606 545 609 558
rect 623 545 626 558
rect 573 496 576 511
rect 587 503 590 507
rect 605 496 608 511
rect 624 496 627 511
rect 630 510 633 551
rect 646 503 649 544
rect 652 511 655 551
rect 671 503 674 544
rect 680 545 683 558
rect 696 562 699 575
rect 717 569 720 572
rect 724 562 727 575
rect 777 575 780 647
rect 788 611 791 683
rect 823 686 826 689
rect 823 683 868 686
rect 823 673 826 683
rect 696 545 699 558
rect 717 548 720 551
rect 724 545 727 558
rect 777 541 780 571
rect 788 555 791 607
rect 795 595 799 661
rect 783 551 787 554
rect 776 538 780 541
rect 777 519 780 538
rect 680 496 683 511
rect 695 496 698 511
rect 702 503 706 506
rect 723 496 726 511
rect 573 477 576 492
rect 587 481 590 485
rect 605 477 608 492
rect 624 477 627 492
rect 573 430 576 443
rect 599 437 602 440
rect 573 413 576 426
rect 606 430 609 443
rect 623 430 626 443
rect 630 437 633 478
rect 646 444 649 485
rect 652 437 655 477
rect 671 444 674 485
rect 680 477 683 492
rect 695 477 698 492
rect 702 482 706 485
rect 723 477 726 492
rect 680 430 683 443
rect 599 416 602 419
rect 606 413 609 426
rect 623 413 626 426
rect 573 364 576 379
rect 587 371 590 375
rect 605 364 608 379
rect 624 364 627 379
rect 630 378 633 419
rect 646 371 649 412
rect 652 379 655 419
rect 671 371 674 412
rect 680 413 683 426
rect 696 430 699 443
rect 717 437 720 440
rect 724 430 727 443
rect 777 444 780 515
rect 788 480 791 551
rect 696 413 699 426
rect 717 416 720 419
rect 724 413 727 426
rect 777 387 780 440
rect 788 423 791 476
rect 795 464 799 529
rect 783 419 787 422
rect 826 422 829 673
rect 841 670 861 673
rect 858 651 861 670
rect 858 575 861 647
rect 869 611 872 683
rect 876 595 880 661
rect 885 562 888 696
rect 1089 693 1092 722
rect 913 690 1020 693
rect 847 558 888 562
rect 847 554 850 558
rect 847 551 892 554
rect 847 541 850 551
rect 865 538 885 541
rect 847 536 850 537
rect 882 519 885 538
rect 882 444 885 515
rect 893 480 896 551
rect 900 464 904 529
rect 680 364 683 379
rect 695 364 698 379
rect 702 371 706 374
rect 723 364 726 379
rect 573 345 576 360
rect 587 349 590 353
rect 605 345 608 360
rect 624 345 627 360
rect 573 298 576 311
rect 599 305 602 308
rect 573 281 576 294
rect 606 298 609 311
rect 623 298 626 311
rect 630 305 633 346
rect 646 312 649 353
rect 652 305 655 345
rect 671 312 674 353
rect 680 345 683 360
rect 695 345 698 360
rect 702 350 706 353
rect 723 345 726 360
rect 680 298 683 311
rect 599 284 602 287
rect 606 281 609 294
rect 623 281 626 294
rect 553 133 559 239
rect 573 232 576 247
rect 587 239 590 243
rect 573 213 576 228
rect 596 225 600 235
rect 605 232 608 247
rect 624 232 627 247
rect 630 246 633 287
rect 646 239 649 280
rect 652 247 655 287
rect 671 239 674 280
rect 680 281 683 294
rect 696 298 699 311
rect 717 305 720 308
rect 724 298 727 311
rect 777 309 780 383
rect 788 345 791 419
rect 823 419 868 422
rect 823 409 826 419
rect 841 406 861 409
rect 696 281 699 294
rect 717 284 720 287
rect 724 281 727 294
rect 777 255 780 305
rect 788 291 791 341
rect 795 329 799 397
rect 858 387 861 406
rect 858 309 861 383
rect 869 345 872 419
rect 913 422 916 690
rect 1024 690 1092 693
rect 1152 658 1155 707
rect 1152 614 1155 654
rect 1160 651 1164 1093
rect 1168 1069 1171 1079
rect 1175 1039 1178 1048
rect 1191 1041 1194 1054
rect 1204 1026 1207 1079
rect 1271 1069 1274 1079
rect 1211 1054 1215 1058
rect 1212 1039 1215 1048
rect 1167 1012 1170 1024
rect 1208 1022 1209 1026
rect 1218 1012 1221 1065
rect 1224 1045 1227 1050
rect 1233 1039 1236 1048
rect 1249 1041 1252 1054
rect 1270 1039 1273 1048
rect 1269 1012 1272 1022
rect 1168 983 1171 993
rect 1175 953 1178 962
rect 1191 955 1194 968
rect 1204 940 1207 993
rect 1271 983 1274 993
rect 1211 968 1215 972
rect 1212 953 1215 962
rect 1167 926 1170 938
rect 1208 936 1209 940
rect 1218 926 1221 979
rect 1224 959 1227 964
rect 1233 953 1236 962
rect 1249 955 1252 968
rect 1270 953 1273 962
rect 1269 926 1272 936
rect 1277 905 1281 1636
rect 1301 1631 1305 1636
rect 1426 1616 1432 1670
rect 1426 1542 1432 1612
rect 1426 1410 1432 1538
rect 1426 1278 1432 1406
rect 1300 1209 1303 1219
rect 1286 1179 1289 1188
rect 1307 1179 1310 1188
rect 1323 1181 1326 1194
rect 1286 1138 1289 1175
rect 1336 1166 1339 1219
rect 1403 1209 1406 1219
rect 1426 1216 1432 1274
rect 1343 1194 1347 1198
rect 1344 1179 1347 1188
rect 1299 1152 1302 1164
rect 1340 1162 1341 1166
rect 1350 1152 1353 1205
rect 1356 1185 1359 1190
rect 1365 1179 1368 1188
rect 1381 1181 1384 1194
rect 1402 1179 1405 1188
rect 1418 1179 1421 1190
rect 1401 1152 1404 1162
rect 1418 1145 1421 1175
rect 1418 1113 1421 1141
rect 1426 1146 1432 1212
rect 1426 1106 1432 1142
rect 1286 1054 1289 1086
rect 1300 1069 1303 1079
rect 1286 1039 1289 1048
rect 1307 1039 1310 1048
rect 1323 1041 1326 1054
rect 1336 1026 1339 1079
rect 1403 1069 1406 1079
rect 1343 1054 1347 1058
rect 1344 1039 1347 1048
rect 1299 1012 1302 1024
rect 1340 1022 1341 1026
rect 1350 1012 1353 1065
rect 1418 1054 1421 1101
rect 1356 1045 1359 1050
rect 1365 1039 1368 1048
rect 1381 1041 1384 1054
rect 1402 1039 1405 1048
rect 1418 1039 1421 1050
rect 1401 1012 1404 1022
rect 1418 1005 1421 1035
rect 1426 1076 1432 1102
rect 1300 983 1303 993
rect 1286 953 1289 962
rect 1307 953 1310 962
rect 1323 955 1326 968
rect 1286 912 1289 949
rect 1336 940 1339 993
rect 1403 983 1406 993
rect 1426 990 1432 1072
rect 1343 968 1347 972
rect 1344 953 1347 962
rect 1299 926 1302 938
rect 1340 936 1341 940
rect 1350 926 1353 979
rect 1356 959 1359 964
rect 1365 953 1368 962
rect 1381 955 1384 968
rect 1402 953 1405 962
rect 1418 953 1421 964
rect 1401 926 1404 936
rect 1418 919 1421 949
rect 1261 894 1265 897
rect 1261 875 1265 890
rect 1277 887 1281 901
rect 1293 901 1297 905
rect 1293 894 1297 897
rect 1293 875 1297 890
rect 1418 887 1421 915
rect 1277 871 1281 872
rect 1293 867 1297 871
rect 1168 843 1171 853
rect 1175 813 1178 822
rect 1191 815 1194 828
rect 1204 800 1207 853
rect 1271 843 1274 853
rect 1211 828 1215 832
rect 1212 813 1215 822
rect 1167 786 1170 798
rect 1208 796 1209 800
rect 1218 786 1221 839
rect 1224 819 1227 824
rect 1233 813 1236 822
rect 1249 815 1252 828
rect 1270 813 1273 822
rect 1269 786 1272 796
rect 1168 731 1171 741
rect 1175 701 1178 710
rect 1191 703 1194 716
rect 1204 688 1207 741
rect 1271 731 1274 741
rect 1211 716 1215 720
rect 1212 701 1215 710
rect 1167 674 1170 686
rect 1208 684 1209 688
rect 1218 674 1221 727
rect 1224 707 1227 712
rect 1233 701 1236 710
rect 1249 703 1252 716
rect 1270 701 1273 710
rect 1269 674 1272 684
rect 1152 599 1155 608
rect 913 419 958 422
rect 913 409 916 419
rect 931 406 951 409
rect 876 329 880 397
rect 948 387 951 406
rect 948 309 951 383
rect 959 345 962 419
rect 966 329 970 397
rect 783 287 787 290
rect 680 232 683 247
rect 695 232 698 247
rect 702 239 706 242
rect 723 232 726 247
rect 587 217 590 221
rect 605 213 608 228
rect 624 213 627 228
rect 573 166 576 179
rect 599 173 602 176
rect 581 159 585 169
rect 606 166 609 179
rect 623 166 626 179
rect 630 173 633 214
rect 646 180 649 221
rect 652 173 655 213
rect 671 180 674 221
rect 680 213 683 228
rect 695 213 698 228
rect 702 218 706 221
rect 723 213 726 228
rect 680 166 683 179
rect 696 166 699 179
rect 717 173 720 176
rect 724 166 727 179
rect 777 173 780 251
rect 788 209 791 287
rect 795 193 799 265
rect 807 166 811 179
rect 816 159 819 169
rect 826 152 829 221
rect 848 217 851 221
rect 866 213 869 228
rect 885 213 888 228
rect 833 166 837 179
rect 860 173 863 176
rect 867 166 870 179
rect 884 166 887 179
rect 891 173 894 214
rect 907 180 910 221
rect 913 173 916 213
rect 932 180 935 221
rect 941 213 944 228
rect 956 213 959 228
rect 963 218 967 221
rect 984 213 987 228
rect 941 166 944 179
rect 957 166 960 179
rect 978 173 981 176
rect 985 166 988 179
rect 1001 160 1005 396
rect 1036 229 1039 239
rect 1043 199 1046 208
rect 1059 201 1062 214
rect 1072 186 1075 239
rect 1139 229 1142 239
rect 1079 214 1083 218
rect 1080 199 1083 208
rect 1035 172 1038 184
rect 1076 182 1077 186
rect 1086 172 1089 225
rect 1092 205 1095 210
rect 1101 199 1104 208
rect 1117 201 1120 214
rect 1138 199 1141 208
rect 1154 199 1157 208
rect 1137 172 1140 182
rect 994 148 995 151
rect 553 103 559 129
rect 553 47 559 99
rect 553 17 559 43
rect 859 40 863 122
rect 874 119 877 129
rect 881 89 884 98
rect 897 91 900 104
rect 910 76 913 129
rect 977 119 980 129
rect 917 104 921 108
rect 918 89 921 98
rect 873 62 876 74
rect 914 72 915 76
rect 924 62 927 115
rect 992 104 995 148
rect 930 95 933 100
rect 939 89 942 98
rect 955 91 958 104
rect 976 89 979 98
rect 992 89 995 98
rect 975 62 978 72
rect 992 55 995 85
rect 553 -123 559 13
rect 867 13 870 50
rect 874 33 877 43
rect 881 3 884 12
rect 897 5 900 18
rect 910 -10 913 43
rect 977 33 980 43
rect 917 18 921 22
rect 918 3 921 12
rect 873 -24 876 -12
rect 914 -14 915 -10
rect 924 -24 927 29
rect 930 9 933 14
rect 939 3 942 12
rect 955 5 958 18
rect 976 3 979 12
rect 992 13 995 14
rect 1013 16 1017 156
rect 1029 69 1032 161
rect 1154 158 1157 195
rect 1160 151 1164 647
rect 1277 660 1281 867
rect 1286 828 1289 860
rect 1300 843 1303 853
rect 1286 813 1289 822
rect 1307 813 1310 822
rect 1323 815 1326 828
rect 1336 800 1339 853
rect 1403 843 1406 853
rect 1343 828 1347 832
rect 1344 813 1347 822
rect 1299 786 1302 798
rect 1340 796 1341 800
rect 1350 786 1353 839
rect 1418 828 1421 875
rect 1356 819 1359 824
rect 1365 813 1368 822
rect 1381 815 1384 828
rect 1402 813 1405 822
rect 1418 820 1421 824
rect 1426 850 1432 986
rect 1418 813 1421 816
rect 1401 786 1404 796
rect 1426 771 1432 846
rect 1426 738 1432 767
rect 1286 708 1289 710
rect 1286 701 1289 704
rect 1286 667 1289 697
rect 1426 694 1432 734
rect 1167 629 1170 639
rect 1168 599 1171 608
rect 1189 601 1192 614
rect 1205 599 1208 608
rect 1214 605 1217 610
rect 1169 572 1172 582
rect 1220 572 1223 625
rect 1226 614 1230 618
rect 1226 599 1229 608
rect 1234 586 1237 639
rect 1270 629 1273 639
rect 1247 601 1250 614
rect 1263 599 1266 608
rect 1232 582 1233 586
rect 1271 572 1274 584
rect 1168 229 1171 239
rect 1175 199 1178 208
rect 1191 201 1194 214
rect 1204 186 1207 239
rect 1271 229 1274 239
rect 1211 214 1215 218
rect 1212 199 1215 208
rect 1167 172 1170 184
rect 1208 182 1209 186
rect 1218 172 1221 225
rect 1224 205 1227 210
rect 1233 199 1236 208
rect 1249 201 1252 214
rect 1270 199 1273 208
rect 1269 172 1272 182
rect 1144 140 1148 143
rect 1144 121 1148 136
rect 1160 133 1164 147
rect 1176 147 1180 151
rect 1176 140 1180 143
rect 1176 121 1180 136
rect 1160 117 1164 118
rect 1176 113 1180 117
rect 1036 89 1039 99
rect 1043 59 1046 68
rect 1059 61 1062 74
rect 1072 46 1075 99
rect 1139 89 1142 99
rect 1079 74 1083 78
rect 1080 59 1083 68
rect 1035 32 1038 44
rect 1076 42 1077 46
rect 1086 32 1089 85
rect 1154 74 1157 106
rect 1092 65 1095 70
rect 1101 59 1104 68
rect 1117 61 1120 74
rect 1138 59 1141 68
rect 1154 59 1157 68
rect 1137 32 1140 42
rect 992 8 995 9
rect 975 -24 978 -14
rect 1013 -86 1017 -4
rect 1029 -17 1032 21
rect 1036 3 1039 13
rect 1043 -27 1046 -18
rect 1059 -25 1062 -12
rect 1072 -40 1075 13
rect 1139 3 1142 13
rect 1079 -12 1083 -8
rect 1080 -27 1083 -18
rect 1035 -54 1038 -42
rect 1076 -44 1077 -40
rect 1086 -54 1089 -1
rect 1092 -21 1095 -16
rect 1101 -27 1104 -18
rect 1117 -25 1120 -12
rect 1138 -27 1141 -18
rect 1154 -27 1157 -18
rect 1137 -54 1140 -44
rect 553 -208 559 -127
rect 1029 -157 1032 -65
rect 1154 -68 1157 -31
rect 1036 -137 1039 -127
rect 1043 -167 1046 -158
rect 1059 -165 1062 -152
rect 1072 -180 1075 -127
rect 1139 -137 1142 -127
rect 1079 -152 1083 -148
rect 1080 -167 1083 -158
rect 1035 -194 1038 -182
rect 1076 -184 1077 -180
rect 1086 -194 1089 -141
rect 1154 -152 1157 -120
rect 1092 -161 1095 -156
rect 1101 -167 1104 -158
rect 1117 -165 1120 -152
rect 1138 -167 1141 -158
rect 1154 -167 1157 -158
rect 1137 -194 1140 -184
rect 1160 -208 1164 113
rect 1168 89 1171 99
rect 1175 59 1178 68
rect 1191 61 1194 74
rect 1204 46 1207 99
rect 1271 89 1274 99
rect 1211 74 1215 78
rect 1212 59 1215 68
rect 1167 32 1170 44
rect 1208 42 1209 46
rect 1218 32 1221 85
rect 1224 65 1227 70
rect 1233 59 1236 68
rect 1249 61 1252 74
rect 1270 59 1273 68
rect 1269 32 1272 42
rect 1168 3 1171 13
rect 1175 -27 1178 -18
rect 1191 -25 1194 -12
rect 1204 -40 1207 13
rect 1271 3 1274 13
rect 1211 -12 1215 -8
rect 1212 -27 1215 -18
rect 1167 -54 1170 -42
rect 1208 -44 1209 -40
rect 1218 -54 1221 -1
rect 1224 -21 1227 -16
rect 1233 -27 1236 -18
rect 1249 -25 1252 -12
rect 1270 -27 1273 -18
rect 1269 -54 1272 -44
rect 1277 -75 1281 656
rect 1301 651 1305 656
rect 1426 636 1432 690
rect 1426 562 1432 632
rect 1426 430 1432 558
rect 1426 298 1432 426
rect 1300 229 1303 239
rect 1286 199 1289 208
rect 1307 199 1310 208
rect 1323 201 1326 214
rect 1286 158 1289 195
rect 1336 186 1339 239
rect 1403 229 1406 239
rect 1426 236 1432 294
rect 1343 214 1347 218
rect 1344 199 1347 208
rect 1299 172 1302 184
rect 1340 182 1341 186
rect 1350 172 1353 225
rect 1356 205 1359 210
rect 1365 199 1368 208
rect 1381 201 1384 214
rect 1402 199 1405 208
rect 1418 199 1421 210
rect 1401 172 1404 182
rect 1418 165 1421 195
rect 1418 133 1421 161
rect 1426 166 1432 232
rect 1426 126 1432 162
rect 1286 74 1289 106
rect 1300 89 1303 99
rect 1286 59 1289 68
rect 1307 59 1310 68
rect 1323 61 1326 74
rect 1336 46 1339 99
rect 1403 89 1406 99
rect 1343 74 1347 78
rect 1344 59 1347 68
rect 1299 32 1302 44
rect 1340 42 1341 46
rect 1350 32 1353 85
rect 1418 74 1421 121
rect 1356 65 1359 70
rect 1365 59 1368 68
rect 1381 61 1384 74
rect 1402 59 1405 68
rect 1418 59 1421 70
rect 1401 32 1404 42
rect 1418 25 1421 55
rect 1426 96 1432 122
rect 1300 3 1303 13
rect 1286 -27 1289 -18
rect 1307 -27 1310 -18
rect 1323 -25 1326 -12
rect 1286 -68 1289 -31
rect 1336 -40 1339 13
rect 1403 3 1406 13
rect 1426 10 1432 92
rect 1343 -12 1347 -8
rect 1344 -27 1347 -18
rect 1299 -54 1302 -42
rect 1340 -44 1341 -40
rect 1350 -54 1353 -1
rect 1356 -21 1359 -16
rect 1365 -27 1368 -18
rect 1381 -25 1384 -12
rect 1402 -27 1405 -18
rect 1418 -27 1421 -16
rect 1401 -54 1404 -44
rect 1418 -61 1421 -31
rect 1261 -86 1265 -83
rect 1261 -105 1265 -90
rect 1277 -93 1281 -79
rect 1293 -79 1297 -75
rect 1293 -86 1297 -83
rect 1293 -105 1297 -90
rect 1418 -93 1421 -65
rect 1277 -109 1281 -108
rect 1293 -113 1297 -109
rect 1168 -137 1171 -127
rect 1175 -167 1178 -158
rect 1191 -165 1194 -152
rect 1204 -180 1207 -127
rect 1271 -137 1274 -127
rect 1211 -152 1215 -148
rect 1212 -167 1215 -158
rect 1167 -194 1170 -182
rect 1208 -184 1209 -180
rect 1218 -194 1221 -141
rect 1224 -161 1227 -156
rect 1233 -167 1236 -158
rect 1249 -165 1252 -152
rect 1270 -167 1273 -158
rect 1269 -194 1272 -184
rect 1277 -208 1281 -113
rect 1286 -152 1289 -120
rect 1300 -137 1303 -127
rect 1286 -167 1289 -158
rect 1307 -167 1310 -158
rect 1323 -165 1326 -152
rect 1336 -180 1339 -127
rect 1403 -137 1406 -127
rect 1343 -152 1347 -148
rect 1344 -167 1347 -158
rect 1299 -194 1302 -182
rect 1340 -184 1341 -180
rect 1350 -194 1353 -141
rect 1418 -152 1421 -105
rect 1356 -161 1359 -156
rect 1365 -167 1368 -158
rect 1381 -165 1384 -152
rect 1402 -167 1405 -158
rect 1418 -160 1421 -156
rect 1426 -130 1432 6
rect 1418 -167 1421 -164
rect 1401 -194 1404 -184
rect 1426 -208 1432 -134
rect 1438 1694 1444 1765
rect 1438 1661 1444 1690
rect 1438 1608 1444 1657
rect 1438 1559 1444 1604
rect 1438 1476 1444 1555
rect 1438 1344 1444 1472
rect 1438 1212 1444 1340
rect 1438 1159 1444 1208
rect 1438 1049 1444 1155
rect 1438 1019 1444 1045
rect 1438 963 1444 1015
rect 1438 933 1444 959
rect 1438 793 1444 929
rect 1438 714 1444 789
rect 1438 681 1444 710
rect 1438 628 1444 677
rect 1438 579 1444 624
rect 1438 496 1444 575
rect 1438 364 1444 492
rect 1438 232 1444 360
rect 1438 179 1444 228
rect 1438 69 1444 175
rect 1438 39 1444 65
rect 1438 -17 1444 35
rect 1438 -47 1444 -21
rect 1438 -187 1444 -51
rect 1438 -208 1444 -191
rect 1450 1615 1456 1765
rect 1450 1601 1456 1611
rect 1450 1483 1456 1597
rect 1450 1469 1456 1479
rect 1450 1351 1456 1465
rect 1450 1337 1456 1347
rect 1450 1205 1456 1333
rect 1450 1131 1456 1201
rect 1450 635 1456 1127
rect 1450 621 1456 631
rect 1450 503 1456 617
rect 1450 489 1456 499
rect 1450 371 1456 485
rect 1450 357 1456 367
rect 1450 225 1456 353
rect 1450 151 1456 221
rect 1450 -208 1456 147
rect 1462 1667 1468 1765
rect 1462 1535 1468 1663
rect 1462 1417 1468 1531
rect 1462 1403 1468 1413
rect 1462 1285 1468 1399
rect 1462 1271 1468 1281
rect 1462 1139 1468 1267
rect 1462 687 1468 1135
rect 1462 555 1468 683
rect 1462 437 1468 551
rect 1462 423 1468 433
rect 1462 305 1468 419
rect 1462 291 1468 301
rect 1462 159 1468 287
rect 1462 -208 1468 155
rect 1474 1687 1480 1765
rect 1474 1654 1480 1683
rect 1474 1552 1480 1650
rect 1474 1153 1480 1548
rect 1474 1042 1480 1149
rect 1474 1012 1480 1038
rect 1474 956 1480 1008
rect 1474 926 1480 952
rect 1474 786 1480 922
rect 1474 707 1480 782
rect 1474 674 1480 703
rect 1474 572 1480 670
rect 1474 173 1480 568
rect 1474 62 1480 169
rect 1474 32 1480 58
rect 1474 -24 1480 28
rect 1474 -54 1480 -28
rect 1474 -194 1480 -58
rect 1474 -208 1480 -198
rect 1486 1758 1492 1765
rect 1486 1725 1492 1754
rect 1508 1744 1511 1754
rect 1486 1623 1492 1721
rect 1515 1714 1518 1723
rect 1531 1716 1534 1729
rect 1544 1701 1547 1754
rect 1611 1744 1614 1754
rect 1640 1744 1643 1754
rect 1551 1729 1555 1733
rect 1552 1714 1555 1723
rect 1507 1687 1510 1699
rect 1548 1697 1549 1701
rect 1558 1687 1561 1740
rect 1564 1720 1567 1725
rect 1573 1714 1576 1723
rect 1589 1716 1592 1729
rect 1610 1714 1613 1723
rect 1626 1723 1629 1725
rect 1626 1720 1633 1723
rect 1626 1714 1629 1720
rect 1647 1714 1650 1723
rect 1663 1716 1666 1729
rect 1609 1687 1612 1697
rect 1626 1680 1629 1710
rect 1676 1701 1679 1754
rect 1743 1744 1746 1754
rect 1772 1744 1775 1754
rect 1683 1729 1687 1733
rect 1684 1714 1687 1723
rect 1639 1687 1642 1699
rect 1680 1697 1681 1701
rect 1690 1687 1693 1740
rect 1696 1720 1699 1725
rect 1705 1714 1708 1723
rect 1721 1716 1724 1729
rect 1742 1714 1745 1723
rect 1758 1723 1761 1725
rect 1758 1720 1765 1723
rect 1758 1714 1761 1720
rect 1779 1714 1782 1723
rect 1795 1716 1798 1729
rect 1741 1687 1744 1697
rect 1626 1677 1678 1680
rect 1506 1657 1509 1670
rect 1532 1660 1535 1663
rect 1539 1657 1542 1670
rect 1556 1657 1559 1670
rect 1486 1223 1492 1619
rect 1506 1608 1509 1623
rect 1520 1615 1523 1619
rect 1538 1608 1541 1623
rect 1557 1608 1560 1623
rect 1563 1622 1566 1663
rect 1579 1615 1582 1656
rect 1585 1623 1588 1663
rect 1604 1615 1607 1656
rect 1613 1657 1616 1670
rect 1629 1657 1632 1670
rect 1650 1660 1653 1663
rect 1657 1657 1660 1670
rect 1675 1666 1678 1677
rect 1758 1674 1761 1710
rect 1808 1701 1811 1754
rect 1875 1744 1878 1754
rect 1904 1744 1907 1754
rect 1815 1729 1819 1733
rect 1816 1714 1819 1723
rect 1771 1687 1774 1699
rect 1812 1697 1813 1701
rect 1822 1687 1825 1740
rect 1828 1720 1831 1725
rect 1837 1714 1840 1723
rect 1853 1716 1856 1729
rect 1874 1714 1877 1723
rect 1890 1723 1893 1725
rect 1890 1720 1897 1723
rect 1890 1714 1893 1720
rect 1911 1714 1914 1723
rect 1927 1716 1930 1729
rect 1873 1687 1876 1697
rect 1890 1680 1893 1702
rect 1940 1701 1943 1754
rect 2007 1744 2010 1754
rect 1947 1729 1951 1733
rect 1948 1714 1951 1723
rect 1903 1687 1906 1699
rect 1944 1697 1945 1701
rect 1954 1687 1957 1740
rect 1960 1720 1963 1725
rect 1969 1714 1972 1723
rect 1985 1716 1988 1729
rect 2006 1714 2009 1723
rect 2022 1723 2025 1725
rect 2022 1720 2026 1723
rect 2022 1714 2025 1720
rect 2022 1706 2025 1710
rect 2005 1687 2008 1697
rect 1756 1669 1761 1674
rect 1818 1676 1893 1680
rect 1675 1663 1720 1666
rect 1675 1653 1678 1663
rect 1693 1650 1713 1653
rect 1710 1631 1713 1650
rect 1613 1608 1616 1623
rect 1628 1608 1631 1623
rect 1635 1615 1639 1618
rect 1656 1608 1659 1623
rect 1506 1589 1509 1604
rect 1520 1593 1523 1597
rect 1538 1589 1541 1604
rect 1557 1589 1560 1604
rect 1506 1542 1509 1555
rect 1532 1549 1535 1552
rect 1506 1525 1509 1538
rect 1516 1535 1520 1545
rect 1539 1542 1542 1555
rect 1556 1542 1559 1555
rect 1563 1549 1566 1590
rect 1579 1556 1582 1597
rect 1585 1549 1588 1589
rect 1604 1556 1607 1597
rect 1613 1589 1616 1604
rect 1628 1589 1631 1604
rect 1635 1594 1639 1597
rect 1656 1589 1659 1604
rect 1613 1542 1616 1555
rect 1532 1528 1535 1531
rect 1539 1525 1542 1538
rect 1556 1525 1559 1538
rect 1506 1476 1509 1491
rect 1520 1483 1523 1487
rect 1538 1476 1541 1491
rect 1557 1476 1560 1491
rect 1563 1490 1566 1531
rect 1579 1483 1582 1524
rect 1585 1491 1588 1531
rect 1604 1483 1607 1524
rect 1613 1525 1616 1538
rect 1629 1542 1632 1555
rect 1650 1549 1653 1552
rect 1657 1542 1660 1555
rect 1710 1555 1713 1627
rect 1721 1591 1724 1663
rect 1756 1666 1759 1669
rect 1756 1663 1801 1666
rect 1756 1653 1759 1663
rect 1629 1525 1632 1538
rect 1650 1528 1653 1531
rect 1657 1525 1660 1538
rect 1710 1521 1713 1551
rect 1721 1535 1724 1587
rect 1728 1575 1732 1641
rect 1716 1531 1720 1534
rect 1709 1518 1713 1521
rect 1710 1499 1713 1518
rect 1613 1476 1616 1491
rect 1628 1476 1631 1491
rect 1635 1483 1639 1486
rect 1656 1476 1659 1491
rect 1506 1457 1509 1472
rect 1520 1461 1523 1465
rect 1538 1457 1541 1472
rect 1557 1457 1560 1472
rect 1506 1410 1509 1423
rect 1532 1417 1535 1420
rect 1506 1393 1509 1406
rect 1539 1410 1542 1423
rect 1556 1410 1559 1423
rect 1563 1417 1566 1458
rect 1579 1424 1582 1465
rect 1585 1417 1588 1457
rect 1604 1424 1607 1465
rect 1613 1457 1616 1472
rect 1628 1457 1631 1472
rect 1635 1462 1639 1465
rect 1656 1457 1659 1472
rect 1613 1410 1616 1423
rect 1532 1396 1535 1399
rect 1539 1393 1542 1406
rect 1556 1393 1559 1406
rect 1506 1344 1509 1359
rect 1520 1351 1523 1355
rect 1538 1344 1541 1359
rect 1557 1344 1560 1359
rect 1563 1358 1566 1399
rect 1579 1351 1582 1392
rect 1585 1359 1588 1399
rect 1604 1351 1607 1392
rect 1613 1393 1616 1406
rect 1629 1410 1632 1423
rect 1650 1417 1653 1420
rect 1657 1410 1660 1423
rect 1710 1424 1713 1495
rect 1721 1460 1724 1531
rect 1629 1393 1632 1406
rect 1650 1396 1653 1399
rect 1657 1393 1660 1406
rect 1710 1367 1713 1420
rect 1721 1403 1724 1456
rect 1728 1444 1732 1509
rect 1716 1399 1720 1402
rect 1759 1402 1762 1653
rect 1774 1650 1794 1653
rect 1791 1631 1794 1650
rect 1791 1555 1794 1627
rect 1802 1591 1805 1663
rect 1809 1575 1813 1641
rect 1818 1542 1821 1676
rect 2022 1673 2025 1702
rect 1846 1670 1953 1673
rect 1780 1538 1821 1542
rect 1780 1534 1783 1538
rect 1780 1531 1825 1534
rect 1780 1521 1783 1531
rect 1798 1518 1818 1521
rect 1780 1516 1783 1517
rect 1815 1499 1818 1518
rect 1815 1424 1818 1495
rect 1826 1460 1829 1531
rect 1833 1444 1837 1509
rect 1613 1344 1616 1359
rect 1628 1344 1631 1359
rect 1635 1351 1639 1354
rect 1656 1344 1659 1359
rect 1506 1325 1509 1340
rect 1520 1329 1523 1333
rect 1538 1325 1541 1340
rect 1557 1325 1560 1340
rect 1506 1278 1509 1291
rect 1532 1285 1535 1288
rect 1506 1261 1509 1274
rect 1539 1278 1542 1291
rect 1556 1278 1559 1291
rect 1563 1285 1566 1326
rect 1579 1292 1582 1333
rect 1585 1285 1588 1325
rect 1604 1292 1607 1333
rect 1613 1325 1616 1340
rect 1628 1325 1631 1340
rect 1635 1330 1639 1333
rect 1656 1325 1659 1340
rect 1613 1278 1616 1291
rect 1532 1264 1535 1267
rect 1539 1261 1542 1274
rect 1556 1261 1559 1274
rect 1486 1113 1492 1219
rect 1506 1212 1509 1227
rect 1520 1219 1523 1223
rect 1506 1193 1509 1208
rect 1529 1205 1533 1215
rect 1538 1212 1541 1227
rect 1557 1212 1560 1227
rect 1563 1226 1566 1267
rect 1579 1219 1582 1260
rect 1585 1227 1588 1267
rect 1604 1219 1607 1260
rect 1613 1261 1616 1274
rect 1629 1278 1632 1291
rect 1650 1285 1653 1288
rect 1657 1278 1660 1291
rect 1710 1289 1713 1363
rect 1721 1325 1724 1399
rect 1756 1399 1801 1402
rect 1756 1389 1759 1399
rect 1774 1386 1794 1389
rect 1629 1261 1632 1274
rect 1650 1264 1653 1267
rect 1657 1261 1660 1274
rect 1710 1235 1713 1285
rect 1721 1271 1724 1321
rect 1728 1309 1732 1377
rect 1791 1367 1794 1386
rect 1791 1289 1794 1363
rect 1802 1325 1805 1399
rect 1846 1402 1849 1670
rect 1957 1670 2025 1673
rect 1846 1399 1891 1402
rect 1846 1389 1849 1399
rect 1864 1386 1884 1389
rect 1809 1309 1813 1377
rect 1881 1367 1884 1386
rect 1881 1289 1884 1363
rect 1892 1325 1895 1399
rect 1899 1309 1903 1377
rect 1716 1267 1720 1270
rect 1613 1212 1616 1227
rect 1628 1212 1631 1227
rect 1635 1219 1639 1222
rect 1656 1212 1659 1227
rect 1520 1197 1523 1201
rect 1538 1193 1541 1208
rect 1557 1193 1560 1208
rect 1506 1146 1509 1159
rect 1532 1153 1535 1156
rect 1514 1139 1518 1149
rect 1539 1146 1542 1159
rect 1556 1146 1559 1159
rect 1563 1153 1566 1194
rect 1579 1160 1582 1201
rect 1585 1153 1588 1193
rect 1604 1160 1607 1201
rect 1613 1193 1616 1208
rect 1628 1193 1631 1208
rect 1635 1198 1639 1201
rect 1656 1193 1659 1208
rect 1613 1146 1616 1159
rect 1629 1146 1632 1159
rect 1650 1153 1653 1156
rect 1657 1146 1660 1159
rect 1710 1153 1713 1231
rect 1721 1189 1724 1267
rect 1728 1173 1732 1245
rect 1740 1146 1744 1159
rect 1749 1139 1752 1149
rect 1759 1132 1762 1201
rect 1781 1197 1784 1201
rect 1799 1193 1802 1208
rect 1818 1193 1821 1208
rect 1766 1146 1770 1159
rect 1793 1153 1796 1156
rect 1800 1146 1803 1159
rect 1817 1146 1820 1159
rect 1824 1153 1827 1194
rect 1840 1160 1843 1201
rect 1846 1153 1849 1193
rect 1865 1160 1868 1201
rect 1874 1193 1877 1208
rect 1889 1193 1892 1208
rect 1896 1198 1900 1201
rect 1917 1193 1920 1208
rect 1874 1146 1877 1159
rect 1890 1146 1893 1159
rect 1911 1153 1914 1156
rect 1918 1146 1921 1159
rect 1934 1140 1938 1376
rect 1927 1128 1928 1131
rect 1486 1083 1492 1109
rect 1486 1027 1492 1079
rect 1486 997 1492 1023
rect 1792 1020 1796 1102
rect 1807 1099 1810 1109
rect 1814 1069 1817 1078
rect 1830 1071 1833 1084
rect 1843 1056 1846 1109
rect 1910 1099 1913 1109
rect 1850 1084 1854 1088
rect 1851 1069 1854 1078
rect 1806 1042 1809 1054
rect 1847 1052 1848 1056
rect 1857 1042 1860 1095
rect 1925 1084 1928 1128
rect 1863 1075 1866 1080
rect 1872 1069 1875 1078
rect 1888 1071 1891 1084
rect 1909 1069 1912 1078
rect 1925 1069 1928 1078
rect 1908 1042 1911 1052
rect 1925 1035 1928 1065
rect 1486 857 1492 993
rect 1800 993 1803 1030
rect 1807 1013 1810 1023
rect 1814 983 1817 992
rect 1830 985 1833 998
rect 1843 970 1846 1023
rect 1910 1013 1913 1023
rect 1850 998 1854 1002
rect 1851 983 1854 992
rect 1806 956 1809 968
rect 1847 966 1848 970
rect 1857 956 1860 1009
rect 1863 989 1866 994
rect 1872 983 1875 992
rect 1888 985 1891 998
rect 1909 983 1912 992
rect 1925 993 1928 994
rect 1946 996 1950 1136
rect 1925 988 1928 989
rect 1908 956 1911 966
rect 1946 894 1950 976
rect 1486 778 1492 853
rect 1486 745 1492 774
rect 1508 764 1511 774
rect 1486 643 1492 741
rect 1515 734 1518 743
rect 1531 736 1534 749
rect 1544 721 1547 774
rect 1611 764 1614 774
rect 1640 764 1643 774
rect 1551 749 1555 753
rect 1552 734 1555 743
rect 1507 707 1510 719
rect 1548 717 1549 721
rect 1558 707 1561 760
rect 1564 740 1567 745
rect 1573 734 1576 743
rect 1589 736 1592 749
rect 1610 734 1613 743
rect 1626 743 1629 745
rect 1626 740 1633 743
rect 1626 734 1629 740
rect 1647 734 1650 743
rect 1663 736 1666 749
rect 1609 707 1612 717
rect 1626 700 1629 730
rect 1676 721 1679 774
rect 1743 764 1746 774
rect 1772 764 1775 774
rect 1683 749 1687 753
rect 1684 734 1687 743
rect 1639 707 1642 719
rect 1680 717 1681 721
rect 1690 707 1693 760
rect 1696 740 1699 745
rect 1705 734 1708 743
rect 1721 736 1724 749
rect 1742 734 1745 743
rect 1758 743 1761 745
rect 1758 740 1765 743
rect 1758 734 1761 740
rect 1779 734 1782 743
rect 1795 736 1798 749
rect 1741 707 1744 717
rect 1626 697 1678 700
rect 1506 677 1509 690
rect 1532 680 1535 683
rect 1539 677 1542 690
rect 1556 677 1559 690
rect 1486 243 1492 639
rect 1506 628 1509 643
rect 1520 635 1523 639
rect 1538 628 1541 643
rect 1557 628 1560 643
rect 1563 642 1566 683
rect 1579 635 1582 676
rect 1585 643 1588 683
rect 1604 635 1607 676
rect 1613 677 1616 690
rect 1629 677 1632 690
rect 1650 680 1653 683
rect 1657 677 1660 690
rect 1675 686 1678 697
rect 1758 694 1761 730
rect 1808 721 1811 774
rect 1875 764 1878 774
rect 1904 764 1907 774
rect 1815 749 1819 753
rect 1816 734 1819 743
rect 1771 707 1774 719
rect 1812 717 1813 721
rect 1822 707 1825 760
rect 1828 740 1831 745
rect 1837 734 1840 743
rect 1853 736 1856 749
rect 1874 734 1877 743
rect 1890 743 1893 745
rect 1890 740 1897 743
rect 1890 734 1893 740
rect 1911 734 1914 743
rect 1927 736 1930 749
rect 1873 707 1876 717
rect 1890 700 1893 722
rect 1940 721 1943 774
rect 2007 764 2010 774
rect 1947 749 1951 753
rect 1948 734 1951 743
rect 1903 707 1906 719
rect 1944 717 1945 721
rect 1954 707 1957 760
rect 1960 740 1963 745
rect 1969 734 1972 743
rect 1985 736 1988 749
rect 2006 734 2009 743
rect 2022 743 2025 745
rect 2022 740 2026 743
rect 2022 734 2025 740
rect 2022 726 2025 730
rect 2005 707 2008 717
rect 1756 689 1761 694
rect 1818 696 1893 700
rect 1675 683 1720 686
rect 1675 673 1678 683
rect 1693 670 1713 673
rect 1710 651 1713 670
rect 1613 628 1616 643
rect 1628 628 1631 643
rect 1635 635 1639 638
rect 1656 628 1659 643
rect 1506 609 1509 624
rect 1520 613 1523 617
rect 1538 609 1541 624
rect 1557 609 1560 624
rect 1506 562 1509 575
rect 1532 569 1535 572
rect 1506 545 1509 558
rect 1516 555 1520 565
rect 1539 562 1542 575
rect 1556 562 1559 575
rect 1563 569 1566 610
rect 1579 576 1582 617
rect 1585 569 1588 609
rect 1604 576 1607 617
rect 1613 609 1616 624
rect 1628 609 1631 624
rect 1635 614 1639 617
rect 1656 609 1659 624
rect 1613 562 1616 575
rect 1532 548 1535 551
rect 1539 545 1542 558
rect 1556 545 1559 558
rect 1506 496 1509 511
rect 1520 503 1523 507
rect 1538 496 1541 511
rect 1557 496 1560 511
rect 1563 510 1566 551
rect 1579 503 1582 544
rect 1585 511 1588 551
rect 1604 503 1607 544
rect 1613 545 1616 558
rect 1629 562 1632 575
rect 1650 569 1653 572
rect 1657 562 1660 575
rect 1710 575 1713 647
rect 1721 611 1724 683
rect 1756 686 1759 689
rect 1756 683 1801 686
rect 1756 673 1759 683
rect 1629 545 1632 558
rect 1650 548 1653 551
rect 1657 545 1660 558
rect 1710 541 1713 571
rect 1721 555 1724 607
rect 1728 595 1732 661
rect 1716 551 1720 554
rect 1709 538 1713 541
rect 1710 519 1713 538
rect 1613 496 1616 511
rect 1628 496 1631 511
rect 1635 503 1639 506
rect 1656 496 1659 511
rect 1506 477 1509 492
rect 1520 481 1523 485
rect 1538 477 1541 492
rect 1557 477 1560 492
rect 1506 430 1509 443
rect 1532 437 1535 440
rect 1506 413 1509 426
rect 1539 430 1542 443
rect 1556 430 1559 443
rect 1563 437 1566 478
rect 1579 444 1582 485
rect 1585 437 1588 477
rect 1604 444 1607 485
rect 1613 477 1616 492
rect 1628 477 1631 492
rect 1635 482 1639 485
rect 1656 477 1659 492
rect 1613 430 1616 443
rect 1532 416 1535 419
rect 1539 413 1542 426
rect 1556 413 1559 426
rect 1506 364 1509 379
rect 1520 371 1523 375
rect 1538 364 1541 379
rect 1557 364 1560 379
rect 1563 378 1566 419
rect 1579 371 1582 412
rect 1585 379 1588 419
rect 1604 371 1607 412
rect 1613 413 1616 426
rect 1629 430 1632 443
rect 1650 437 1653 440
rect 1657 430 1660 443
rect 1710 444 1713 515
rect 1721 480 1724 551
rect 1629 413 1632 426
rect 1650 416 1653 419
rect 1657 413 1660 426
rect 1710 387 1713 440
rect 1721 423 1724 476
rect 1728 464 1732 529
rect 1716 419 1720 422
rect 1759 422 1762 673
rect 1774 670 1794 673
rect 1791 651 1794 670
rect 1791 575 1794 647
rect 1802 611 1805 683
rect 1809 595 1813 661
rect 1818 562 1821 696
rect 2022 693 2025 722
rect 1846 690 1953 693
rect 1780 558 1821 562
rect 1780 554 1783 558
rect 1780 551 1825 554
rect 1780 541 1783 551
rect 1798 538 1818 541
rect 1780 536 1783 537
rect 1815 519 1818 538
rect 1815 444 1818 515
rect 1826 480 1829 551
rect 1833 464 1837 529
rect 1613 364 1616 379
rect 1628 364 1631 379
rect 1635 371 1639 374
rect 1656 364 1659 379
rect 1506 345 1509 360
rect 1520 349 1523 353
rect 1538 345 1541 360
rect 1557 345 1560 360
rect 1506 298 1509 311
rect 1532 305 1535 308
rect 1506 281 1509 294
rect 1539 298 1542 311
rect 1556 298 1559 311
rect 1563 305 1566 346
rect 1579 312 1582 353
rect 1585 305 1588 345
rect 1604 312 1607 353
rect 1613 345 1616 360
rect 1628 345 1631 360
rect 1635 350 1639 353
rect 1656 345 1659 360
rect 1613 298 1616 311
rect 1532 284 1535 287
rect 1539 281 1542 294
rect 1556 281 1559 294
rect 1486 133 1492 239
rect 1506 232 1509 247
rect 1520 239 1523 243
rect 1506 213 1509 228
rect 1529 225 1533 235
rect 1538 232 1541 247
rect 1557 232 1560 247
rect 1563 246 1566 287
rect 1579 239 1582 280
rect 1585 247 1588 287
rect 1604 239 1607 280
rect 1613 281 1616 294
rect 1629 298 1632 311
rect 1650 305 1653 308
rect 1657 298 1660 311
rect 1710 309 1713 383
rect 1721 345 1724 419
rect 1756 419 1801 422
rect 1756 409 1759 419
rect 1774 406 1794 409
rect 1629 281 1632 294
rect 1650 284 1653 287
rect 1657 281 1660 294
rect 1710 255 1713 305
rect 1721 291 1724 341
rect 1728 329 1732 397
rect 1791 387 1794 406
rect 1791 309 1794 383
rect 1802 345 1805 419
rect 1846 422 1849 690
rect 1957 690 2025 693
rect 1846 419 1891 422
rect 1846 409 1849 419
rect 1864 406 1884 409
rect 1809 329 1813 397
rect 1881 387 1884 406
rect 1881 309 1884 383
rect 1892 345 1895 419
rect 1899 329 1903 397
rect 1716 287 1720 290
rect 1613 232 1616 247
rect 1628 232 1631 247
rect 1635 239 1639 242
rect 1656 232 1659 247
rect 1520 217 1523 221
rect 1538 213 1541 228
rect 1557 213 1560 228
rect 1506 166 1509 179
rect 1532 173 1535 176
rect 1514 159 1518 169
rect 1539 166 1542 179
rect 1556 166 1559 179
rect 1563 173 1566 214
rect 1579 180 1582 221
rect 1585 173 1588 213
rect 1604 180 1607 221
rect 1613 213 1616 228
rect 1628 213 1631 228
rect 1635 218 1639 221
rect 1656 213 1659 228
rect 1613 166 1616 179
rect 1629 166 1632 179
rect 1650 173 1653 176
rect 1657 166 1660 179
rect 1710 173 1713 251
rect 1721 209 1724 287
rect 1728 193 1732 265
rect 1740 166 1744 179
rect 1749 159 1752 169
rect 1759 152 1762 221
rect 1781 217 1784 221
rect 1799 213 1802 228
rect 1818 213 1821 228
rect 1766 166 1770 179
rect 1793 173 1796 176
rect 1800 166 1803 179
rect 1817 166 1820 179
rect 1824 173 1827 214
rect 1840 180 1843 221
rect 1846 173 1849 213
rect 1865 180 1868 221
rect 1874 213 1877 228
rect 1889 213 1892 228
rect 1896 218 1900 221
rect 1917 213 1920 228
rect 1874 166 1877 179
rect 1890 166 1893 179
rect 1911 173 1914 176
rect 1918 166 1921 179
rect 1934 160 1938 396
rect 1927 148 1928 151
rect 1486 103 1492 129
rect 1486 47 1492 99
rect 1486 17 1492 43
rect 1792 40 1796 122
rect 1807 119 1810 129
rect 1814 89 1817 98
rect 1830 91 1833 104
rect 1843 76 1846 129
rect 1910 119 1913 129
rect 1850 104 1854 108
rect 1851 89 1854 98
rect 1806 62 1809 74
rect 1847 72 1848 76
rect 1857 62 1860 115
rect 1925 104 1928 148
rect 1863 95 1866 100
rect 1872 89 1875 98
rect 1888 91 1891 104
rect 1909 89 1912 98
rect 1925 89 1928 98
rect 1908 62 1911 72
rect 1925 55 1928 85
rect 1486 -123 1492 13
rect 1800 13 1803 50
rect 1807 33 1810 43
rect 1814 3 1817 12
rect 1830 5 1833 18
rect 1843 -10 1846 43
rect 1910 33 1913 43
rect 1850 18 1854 22
rect 1851 3 1854 12
rect 1806 -24 1809 -12
rect 1847 -14 1848 -10
rect 1857 -24 1860 29
rect 1863 9 1866 14
rect 1872 3 1875 12
rect 1888 5 1891 18
rect 1909 3 1912 12
rect 1925 13 1928 14
rect 1946 16 1950 156
rect 1925 8 1928 9
rect 1908 -24 1911 -14
rect 1946 -86 1950 -4
rect 1486 -208 1492 -127
<< m3contact >>
rect 96 1181 100 1185
rect 353 1684 357 1688
rect 352 1581 356 1585
rect 96 201 100 205
rect 485 816 489 820
rect 353 704 357 708
rect 352 601 356 605
rect 485 -164 489 -160
rect 564 1720 568 1724
rect 604 1637 609 1642
rect 615 1633 620 1638
rect 638 1642 643 1647
rect 662 1637 667 1642
rect 677 1641 682 1647
rect 707 1637 712 1642
rect 736 1636 741 1641
rect 691 1631 696 1636
rect 720 1631 724 1636
rect 762 1630 767 1635
rect 568 1577 573 1582
rect 604 1570 609 1575
rect 615 1574 620 1579
rect 638 1565 643 1570
rect 662 1570 667 1575
rect 691 1576 696 1581
rect 720 1576 724 1581
rect 677 1565 682 1571
rect 707 1570 712 1575
rect 736 1571 741 1576
rect 762 1571 767 1576
rect 567 1508 572 1513
rect 604 1505 609 1510
rect 615 1501 620 1506
rect 638 1510 643 1515
rect 662 1505 667 1510
rect 818 1636 823 1641
rect 677 1509 682 1515
rect 707 1505 712 1510
rect 736 1504 741 1509
rect 691 1499 696 1504
rect 720 1499 724 1504
rect 762 1498 767 1503
rect 568 1445 573 1450
rect 604 1438 609 1443
rect 615 1442 620 1447
rect 638 1433 643 1438
rect 662 1438 667 1443
rect 691 1444 696 1449
rect 720 1444 724 1449
rect 677 1433 682 1439
rect 707 1438 712 1443
rect 736 1439 741 1444
rect 761 1440 766 1445
rect 567 1376 572 1381
rect 604 1373 609 1378
rect 615 1369 620 1374
rect 638 1378 643 1383
rect 662 1373 667 1378
rect 677 1377 682 1383
rect 707 1373 712 1378
rect 736 1372 741 1377
rect 691 1367 696 1372
rect 720 1367 724 1372
rect 762 1366 767 1371
rect 818 1512 823 1517
rect 843 1630 848 1635
rect 842 1571 847 1576
rect 903 1636 908 1641
rect 867 1498 872 1503
rect 867 1440 872 1445
rect 568 1313 573 1318
rect 604 1306 609 1311
rect 615 1310 620 1315
rect 638 1301 643 1306
rect 662 1306 667 1311
rect 691 1312 696 1317
rect 720 1312 724 1317
rect 677 1301 682 1307
rect 707 1306 712 1311
rect 736 1307 741 1312
rect 762 1305 767 1310
rect 567 1244 572 1249
rect 604 1241 609 1246
rect 615 1237 620 1242
rect 638 1246 643 1251
rect 662 1241 667 1246
rect 677 1245 682 1251
rect 707 1241 712 1246
rect 736 1240 741 1245
rect 691 1235 696 1240
rect 720 1235 724 1240
rect 762 1234 767 1239
rect 818 1372 823 1377
rect 843 1366 848 1371
rect 842 1305 847 1310
rect 1020 1669 1024 1673
rect 925 1509 930 1514
rect 900 1381 905 1386
rect 934 1374 939 1379
rect 931 1301 936 1306
rect 568 1181 573 1186
rect 604 1174 609 1179
rect 615 1178 620 1183
rect 638 1169 643 1174
rect 662 1174 667 1179
rect 691 1180 696 1185
rect 720 1180 724 1185
rect 677 1169 682 1175
rect 707 1174 712 1179
rect 736 1175 741 1180
rect 761 1169 766 1174
rect 818 1248 823 1253
rect 806 1180 811 1185
rect 865 1174 870 1179
rect 876 1178 881 1183
rect 899 1169 904 1174
rect 923 1174 928 1179
rect 952 1180 957 1185
rect 981 1180 985 1185
rect 938 1169 943 1175
rect 968 1174 973 1179
rect 993 1180 998 1185
rect 1029 1181 1033 1185
rect 867 1071 871 1075
rect 1286 1684 1290 1688
rect 992 989 996 993
rect 564 740 568 744
rect 604 657 609 662
rect 615 653 620 658
rect 638 662 643 667
rect 662 657 667 662
rect 677 661 682 667
rect 707 657 712 662
rect 736 656 741 661
rect 691 651 696 656
rect 720 651 724 656
rect 762 650 767 655
rect 568 597 573 602
rect 604 590 609 595
rect 615 594 620 599
rect 638 585 643 590
rect 662 590 667 595
rect 691 596 696 601
rect 720 596 724 601
rect 677 585 682 591
rect 707 590 712 595
rect 736 591 741 596
rect 762 591 767 596
rect 567 528 572 533
rect 604 525 609 530
rect 615 521 620 526
rect 638 530 643 535
rect 662 525 667 530
rect 818 656 823 661
rect 677 529 682 535
rect 707 525 712 530
rect 736 524 741 529
rect 691 519 696 524
rect 720 519 724 524
rect 762 518 767 523
rect 568 465 573 470
rect 604 458 609 463
rect 615 462 620 467
rect 638 453 643 458
rect 662 458 667 463
rect 691 464 696 469
rect 720 464 724 469
rect 677 453 682 459
rect 707 458 712 463
rect 736 459 741 464
rect 761 460 766 465
rect 567 396 572 401
rect 604 393 609 398
rect 615 389 620 394
rect 638 398 643 403
rect 662 393 667 398
rect 677 397 682 403
rect 707 393 712 398
rect 736 392 741 397
rect 691 387 696 392
rect 720 387 724 392
rect 762 386 767 391
rect 818 532 823 537
rect 843 650 848 655
rect 842 591 847 596
rect 903 656 908 661
rect 867 518 872 523
rect 867 460 872 465
rect 568 333 573 338
rect 604 326 609 331
rect 615 330 620 335
rect 638 321 643 326
rect 662 326 667 331
rect 691 332 696 337
rect 720 332 724 337
rect 677 321 682 327
rect 707 326 712 331
rect 736 327 741 332
rect 762 325 767 330
rect 567 264 572 269
rect 604 261 609 266
rect 615 257 620 262
rect 638 266 643 271
rect 662 261 667 266
rect 677 265 682 271
rect 707 261 712 266
rect 736 260 741 265
rect 691 255 696 260
rect 720 255 724 260
rect 762 254 767 259
rect 818 392 823 397
rect 843 386 848 391
rect 842 325 847 330
rect 1020 689 1024 693
rect 1285 1581 1289 1585
rect 925 529 930 534
rect 900 401 905 406
rect 934 394 939 399
rect 931 321 936 326
rect 568 201 573 206
rect 604 194 609 199
rect 615 198 620 203
rect 638 189 643 194
rect 662 194 667 199
rect 691 200 696 205
rect 720 200 724 205
rect 677 189 682 195
rect 707 194 712 199
rect 736 195 741 200
rect 761 189 766 194
rect 818 268 823 273
rect 806 200 811 205
rect 865 194 870 199
rect 876 198 881 203
rect 899 189 904 194
rect 923 194 928 199
rect 952 200 957 205
rect 981 200 985 205
rect 938 189 943 195
rect 968 194 973 199
rect 993 200 998 205
rect 1029 201 1033 205
rect 867 91 871 95
rect 1418 816 1422 820
rect 1286 704 1290 708
rect 992 9 996 13
rect 1285 601 1289 605
rect 1418 -164 1422 -160
rect 1497 1720 1501 1724
rect 1537 1637 1542 1642
rect 1548 1633 1553 1638
rect 1571 1642 1576 1647
rect 1595 1637 1600 1642
rect 1610 1641 1615 1647
rect 1640 1637 1645 1642
rect 1669 1636 1674 1641
rect 1624 1631 1629 1636
rect 1653 1631 1657 1636
rect 1695 1630 1700 1635
rect 1501 1577 1506 1582
rect 1537 1570 1542 1575
rect 1548 1574 1553 1579
rect 1571 1565 1576 1570
rect 1595 1570 1600 1575
rect 1624 1576 1629 1581
rect 1653 1576 1657 1581
rect 1610 1565 1615 1571
rect 1640 1570 1645 1575
rect 1669 1571 1674 1576
rect 1695 1571 1700 1576
rect 1500 1508 1505 1513
rect 1537 1505 1542 1510
rect 1548 1501 1553 1506
rect 1571 1510 1576 1515
rect 1595 1505 1600 1510
rect 1751 1636 1756 1641
rect 1610 1509 1615 1515
rect 1640 1505 1645 1510
rect 1669 1504 1674 1509
rect 1624 1499 1629 1504
rect 1653 1499 1657 1504
rect 1695 1498 1700 1503
rect 1501 1445 1506 1450
rect 1537 1438 1542 1443
rect 1548 1442 1553 1447
rect 1571 1433 1576 1438
rect 1595 1438 1600 1443
rect 1624 1444 1629 1449
rect 1653 1444 1657 1449
rect 1610 1433 1615 1439
rect 1640 1438 1645 1443
rect 1669 1439 1674 1444
rect 1694 1440 1699 1445
rect 1500 1376 1505 1381
rect 1537 1373 1542 1378
rect 1548 1369 1553 1374
rect 1571 1378 1576 1383
rect 1595 1373 1600 1378
rect 1610 1377 1615 1383
rect 1640 1373 1645 1378
rect 1669 1372 1674 1377
rect 1624 1367 1629 1372
rect 1653 1367 1657 1372
rect 1695 1366 1700 1371
rect 1751 1512 1756 1517
rect 1776 1630 1781 1635
rect 1775 1571 1780 1576
rect 1836 1636 1841 1641
rect 1800 1498 1805 1503
rect 1800 1440 1805 1445
rect 1501 1313 1506 1318
rect 1537 1306 1542 1311
rect 1548 1310 1553 1315
rect 1571 1301 1576 1306
rect 1595 1306 1600 1311
rect 1624 1312 1629 1317
rect 1653 1312 1657 1317
rect 1610 1301 1615 1307
rect 1640 1306 1645 1311
rect 1669 1307 1674 1312
rect 1695 1305 1700 1310
rect 1500 1244 1505 1249
rect 1537 1241 1542 1246
rect 1548 1237 1553 1242
rect 1571 1246 1576 1251
rect 1595 1241 1600 1246
rect 1610 1245 1615 1251
rect 1640 1241 1645 1246
rect 1669 1240 1674 1245
rect 1624 1235 1629 1240
rect 1653 1235 1657 1240
rect 1695 1234 1700 1239
rect 1751 1372 1756 1377
rect 1776 1366 1781 1371
rect 1775 1305 1780 1310
rect 1953 1669 1957 1673
rect 1858 1509 1863 1514
rect 1833 1381 1838 1386
rect 1867 1374 1872 1379
rect 1864 1301 1869 1306
rect 1501 1181 1506 1186
rect 1537 1174 1542 1179
rect 1548 1178 1553 1183
rect 1571 1169 1576 1174
rect 1595 1174 1600 1179
rect 1624 1180 1629 1185
rect 1653 1180 1657 1185
rect 1610 1169 1615 1175
rect 1640 1174 1645 1179
rect 1669 1175 1674 1180
rect 1694 1169 1699 1174
rect 1751 1248 1756 1253
rect 1739 1180 1744 1185
rect 1798 1174 1803 1179
rect 1809 1178 1814 1183
rect 1832 1169 1837 1174
rect 1856 1174 1861 1179
rect 1885 1180 1890 1185
rect 1914 1180 1918 1185
rect 1871 1169 1876 1175
rect 1901 1174 1906 1179
rect 1926 1180 1931 1185
rect 1800 1071 1804 1075
rect 1925 989 1929 993
rect 1497 740 1501 744
rect 1537 657 1542 662
rect 1548 653 1553 658
rect 1571 662 1576 667
rect 1595 657 1600 662
rect 1610 661 1615 667
rect 1640 657 1645 662
rect 1669 656 1674 661
rect 1624 651 1629 656
rect 1653 651 1657 656
rect 1695 650 1700 655
rect 1501 597 1506 602
rect 1537 590 1542 595
rect 1548 594 1553 599
rect 1571 585 1576 590
rect 1595 590 1600 595
rect 1624 596 1629 601
rect 1653 596 1657 601
rect 1610 585 1615 591
rect 1640 590 1645 595
rect 1669 591 1674 596
rect 1695 591 1700 596
rect 1500 528 1505 533
rect 1537 525 1542 530
rect 1548 521 1553 526
rect 1571 530 1576 535
rect 1595 525 1600 530
rect 1751 656 1756 661
rect 1610 529 1615 535
rect 1640 525 1645 530
rect 1669 524 1674 529
rect 1624 519 1629 524
rect 1653 519 1657 524
rect 1695 518 1700 523
rect 1501 465 1506 470
rect 1537 458 1542 463
rect 1548 462 1553 467
rect 1571 453 1576 458
rect 1595 458 1600 463
rect 1624 464 1629 469
rect 1653 464 1657 469
rect 1610 453 1615 459
rect 1640 458 1645 463
rect 1669 459 1674 464
rect 1694 460 1699 465
rect 1500 396 1505 401
rect 1537 393 1542 398
rect 1548 389 1553 394
rect 1571 398 1576 403
rect 1595 393 1600 398
rect 1610 397 1615 403
rect 1640 393 1645 398
rect 1669 392 1674 397
rect 1624 387 1629 392
rect 1653 387 1657 392
rect 1695 386 1700 391
rect 1751 532 1756 537
rect 1776 650 1781 655
rect 1775 591 1780 596
rect 1836 656 1841 661
rect 1800 518 1805 523
rect 1800 460 1805 465
rect 1501 333 1506 338
rect 1537 326 1542 331
rect 1548 330 1553 335
rect 1571 321 1576 326
rect 1595 326 1600 331
rect 1624 332 1629 337
rect 1653 332 1657 337
rect 1610 321 1615 327
rect 1640 326 1645 331
rect 1669 327 1674 332
rect 1695 325 1700 330
rect 1500 264 1505 269
rect 1537 261 1542 266
rect 1548 257 1553 262
rect 1571 266 1576 271
rect 1595 261 1600 266
rect 1610 265 1615 271
rect 1640 261 1645 266
rect 1669 260 1674 265
rect 1624 255 1629 260
rect 1653 255 1657 260
rect 1695 254 1700 259
rect 1751 392 1756 397
rect 1776 386 1781 391
rect 1775 325 1780 330
rect 1953 689 1957 693
rect 1858 529 1863 534
rect 1833 401 1838 406
rect 1867 394 1872 399
rect 1864 321 1869 326
rect 1501 201 1506 206
rect 1537 194 1542 199
rect 1548 198 1553 203
rect 1571 189 1576 194
rect 1595 194 1600 199
rect 1624 200 1629 205
rect 1653 200 1657 205
rect 1610 189 1615 195
rect 1640 194 1645 199
rect 1669 195 1674 200
rect 1694 189 1699 194
rect 1751 268 1756 273
rect 1739 200 1744 205
rect 1798 194 1803 199
rect 1809 198 1814 203
rect 1832 189 1837 194
rect 1856 194 1861 199
rect 1885 200 1890 205
rect 1914 200 1918 205
rect 1871 189 1876 195
rect 1901 194 1906 199
rect 1926 200 1931 205
rect 1800 91 1804 95
rect 1925 9 1929 13
<< metal3 >>
rect 563 1724 569 1725
rect 563 1720 564 1724
rect 568 1720 569 1724
rect 563 1719 569 1720
rect 1496 1724 1502 1725
rect 1496 1720 1497 1724
rect 1501 1720 1502 1724
rect 1496 1719 1502 1720
rect 563 1689 568 1719
rect 1496 1689 1501 1719
rect 352 1688 568 1689
rect 352 1684 353 1688
rect 357 1684 568 1688
rect 1285 1688 1501 1689
rect 1285 1684 1286 1688
rect 1290 1684 1501 1688
rect 352 1683 358 1684
rect 1285 1683 1291 1684
rect 1019 1673 1025 1674
rect 1019 1669 1020 1673
rect 1024 1669 1025 1673
rect 1019 1668 1025 1669
rect 1952 1673 1958 1674
rect 1952 1669 1953 1673
rect 1957 1669 1958 1673
rect 1952 1668 1958 1669
rect 604 1647 644 1648
rect 604 1643 638 1647
rect 603 1642 610 1643
rect 603 1637 604 1642
rect 609 1637 610 1642
rect 637 1642 638 1643
rect 643 1642 644 1647
rect 676 1647 712 1652
rect 637 1641 644 1642
rect 661 1642 668 1643
rect 603 1636 610 1637
rect 614 1638 621 1639
rect 614 1633 615 1638
rect 620 1633 621 1638
rect 661 1637 662 1642
rect 667 1637 668 1642
rect 676 1641 677 1647
rect 682 1646 712 1647
rect 682 1641 683 1646
rect 707 1643 712 1646
rect 676 1640 683 1641
rect 706 1642 713 1643
rect 706 1637 707 1642
rect 712 1637 713 1642
rect 735 1641 742 1642
rect 661 1636 668 1637
rect 690 1636 697 1637
rect 706 1636 713 1637
rect 719 1636 725 1637
rect 662 1633 667 1636
rect 614 1628 667 1633
rect 690 1631 691 1636
rect 696 1631 697 1636
rect 719 1631 720 1636
rect 724 1631 725 1636
rect 690 1630 725 1631
rect 691 1626 725 1630
rect 735 1636 736 1641
rect 741 1636 742 1641
rect 817 1641 824 1642
rect 817 1636 818 1641
rect 823 1636 824 1641
rect 902 1641 909 1642
rect 902 1636 903 1641
rect 908 1636 909 1641
rect 735 1635 742 1636
rect 761 1635 768 1636
rect 817 1635 824 1636
rect 842 1635 849 1636
rect 902 1635 909 1636
rect 735 1630 762 1635
rect 767 1630 768 1635
rect 818 1630 843 1635
rect 848 1630 849 1635
rect 735 1609 740 1630
rect 761 1629 768 1630
rect 842 1629 849 1630
rect 899 1630 908 1635
rect 568 1603 740 1609
rect 351 1585 357 1586
rect 351 1581 352 1585
rect 356 1581 489 1585
rect 568 1583 573 1603
rect 351 1580 489 1581
rect 95 1185 101 1186
rect 95 1181 96 1185
rect 100 1181 101 1185
rect 95 1180 101 1181
rect 484 821 489 1580
rect 567 1582 574 1583
rect 567 1577 568 1582
rect 573 1577 574 1582
rect 567 1576 574 1577
rect 614 1579 667 1584
rect 691 1582 725 1586
rect 603 1575 610 1576
rect 603 1570 604 1575
rect 609 1570 610 1575
rect 614 1574 615 1579
rect 620 1574 621 1579
rect 662 1576 667 1579
rect 690 1581 725 1582
rect 690 1576 691 1581
rect 696 1576 697 1581
rect 719 1576 720 1581
rect 724 1576 725 1581
rect 614 1573 621 1574
rect 661 1575 668 1576
rect 690 1575 697 1576
rect 706 1575 713 1576
rect 719 1575 725 1576
rect 735 1576 742 1577
rect 761 1576 768 1577
rect 841 1576 848 1577
rect 603 1569 610 1570
rect 637 1570 644 1571
rect 637 1569 638 1570
rect 604 1565 638 1569
rect 643 1565 644 1570
rect 661 1570 662 1575
rect 667 1570 668 1575
rect 661 1569 668 1570
rect 676 1571 683 1572
rect 604 1564 644 1565
rect 676 1565 677 1571
rect 682 1566 683 1571
rect 706 1570 707 1575
rect 712 1570 713 1575
rect 735 1571 736 1576
rect 741 1571 762 1576
rect 767 1571 768 1576
rect 735 1570 742 1571
rect 761 1570 768 1571
rect 818 1571 842 1576
rect 847 1571 848 1576
rect 706 1569 713 1570
rect 707 1566 712 1569
rect 682 1565 712 1566
rect 676 1560 712 1565
rect 736 1543 741 1570
rect 567 1537 741 1543
rect 567 1514 572 1537
rect 604 1515 644 1516
rect 566 1513 573 1514
rect 566 1508 567 1513
rect 572 1508 573 1513
rect 604 1511 638 1515
rect 566 1507 573 1508
rect 603 1510 610 1511
rect 603 1505 604 1510
rect 609 1505 610 1510
rect 637 1510 638 1511
rect 643 1510 644 1515
rect 676 1515 712 1520
rect 818 1518 823 1571
rect 841 1570 848 1571
rect 899 1542 904 1630
rect 861 1537 904 1542
rect 637 1509 644 1510
rect 661 1510 668 1511
rect 603 1504 610 1505
rect 614 1506 621 1507
rect 614 1501 615 1506
rect 620 1501 621 1506
rect 661 1505 662 1510
rect 667 1505 668 1510
rect 676 1509 677 1515
rect 682 1514 712 1515
rect 682 1509 683 1514
rect 707 1511 712 1514
rect 817 1517 824 1518
rect 817 1512 818 1517
rect 823 1512 824 1517
rect 817 1511 824 1512
rect 676 1508 683 1509
rect 706 1510 713 1511
rect 706 1505 707 1510
rect 712 1505 713 1510
rect 735 1509 742 1510
rect 661 1504 668 1505
rect 690 1504 697 1505
rect 706 1504 713 1505
rect 719 1504 725 1505
rect 662 1501 667 1504
rect 614 1496 667 1501
rect 690 1499 691 1504
rect 696 1499 697 1504
rect 719 1499 720 1504
rect 724 1499 725 1504
rect 690 1498 725 1499
rect 691 1494 725 1498
rect 735 1504 736 1509
rect 741 1504 742 1509
rect 861 1504 866 1537
rect 924 1514 931 1515
rect 924 1509 925 1514
rect 930 1509 931 1514
rect 924 1508 931 1509
rect 735 1503 742 1504
rect 761 1503 768 1504
rect 735 1498 762 1503
rect 767 1498 768 1503
rect 861 1503 873 1504
rect 861 1498 867 1503
rect 872 1498 873 1503
rect 735 1477 740 1498
rect 761 1497 768 1498
rect 866 1497 873 1498
rect 568 1471 740 1477
rect 568 1451 573 1471
rect 567 1450 574 1451
rect 567 1445 568 1450
rect 573 1445 574 1450
rect 567 1444 574 1445
rect 614 1447 667 1452
rect 691 1450 725 1454
rect 603 1443 610 1444
rect 603 1438 604 1443
rect 609 1438 610 1443
rect 614 1442 615 1447
rect 620 1442 621 1447
rect 662 1444 667 1447
rect 690 1449 725 1450
rect 690 1444 691 1449
rect 696 1444 697 1449
rect 719 1444 720 1449
rect 724 1444 725 1449
rect 760 1445 767 1446
rect 866 1445 873 1446
rect 614 1441 621 1442
rect 661 1443 668 1444
rect 690 1443 697 1444
rect 706 1443 713 1444
rect 719 1443 725 1444
rect 735 1444 761 1445
rect 603 1437 610 1438
rect 637 1438 644 1439
rect 637 1437 638 1438
rect 604 1433 638 1437
rect 643 1433 644 1438
rect 661 1438 662 1443
rect 667 1438 668 1443
rect 661 1437 668 1438
rect 676 1439 683 1440
rect 604 1432 644 1433
rect 676 1433 677 1439
rect 682 1434 683 1439
rect 706 1438 707 1443
rect 712 1438 713 1443
rect 706 1437 713 1438
rect 735 1439 736 1444
rect 741 1440 761 1444
rect 766 1440 767 1445
rect 741 1439 742 1440
rect 760 1439 767 1440
rect 862 1440 867 1445
rect 872 1440 873 1445
rect 862 1439 873 1440
rect 735 1438 742 1439
rect 707 1434 712 1437
rect 682 1433 712 1434
rect 676 1428 712 1433
rect 735 1411 740 1438
rect 567 1405 740 1411
rect 862 1411 867 1439
rect 862 1406 905 1411
rect 567 1382 572 1405
rect 604 1383 644 1384
rect 566 1381 573 1382
rect 566 1376 567 1381
rect 572 1376 573 1381
rect 604 1379 638 1383
rect 566 1375 573 1376
rect 603 1378 610 1379
rect 603 1373 604 1378
rect 609 1373 610 1378
rect 637 1378 638 1379
rect 643 1378 644 1383
rect 676 1383 712 1388
rect 900 1387 905 1406
rect 637 1377 644 1378
rect 661 1378 668 1379
rect 603 1372 610 1373
rect 614 1374 621 1375
rect 614 1369 615 1374
rect 620 1369 621 1374
rect 661 1373 662 1378
rect 667 1373 668 1378
rect 676 1377 677 1383
rect 682 1382 712 1383
rect 682 1377 683 1382
rect 707 1379 712 1382
rect 899 1386 906 1387
rect 899 1381 900 1386
rect 905 1381 906 1386
rect 899 1380 906 1381
rect 925 1379 930 1508
rect 933 1379 940 1380
rect 676 1376 683 1377
rect 706 1378 713 1379
rect 706 1373 707 1378
rect 712 1373 713 1378
rect 735 1377 742 1378
rect 661 1372 668 1373
rect 690 1372 697 1373
rect 706 1372 713 1373
rect 719 1372 725 1373
rect 662 1369 667 1372
rect 614 1364 667 1369
rect 690 1367 691 1372
rect 696 1367 697 1372
rect 719 1367 720 1372
rect 724 1367 725 1372
rect 690 1366 725 1367
rect 691 1362 725 1366
rect 735 1372 736 1377
rect 741 1372 742 1377
rect 817 1377 824 1378
rect 817 1372 818 1377
rect 823 1372 824 1377
rect 913 1374 934 1379
rect 939 1374 940 1379
rect 913 1373 925 1374
rect 933 1373 940 1374
rect 735 1371 742 1372
rect 761 1371 768 1372
rect 817 1371 824 1372
rect 842 1371 849 1372
rect 735 1366 762 1371
rect 767 1366 768 1371
rect 818 1366 843 1371
rect 848 1366 849 1371
rect 735 1345 740 1366
rect 761 1365 768 1366
rect 842 1365 849 1366
rect 913 1365 918 1373
rect 568 1339 740 1345
rect 880 1344 918 1365
rect 568 1319 573 1339
rect 567 1318 574 1319
rect 567 1313 568 1318
rect 573 1313 574 1318
rect 567 1312 574 1313
rect 614 1315 667 1320
rect 691 1318 725 1322
rect 603 1311 610 1312
rect 603 1306 604 1311
rect 609 1306 610 1311
rect 614 1310 615 1315
rect 620 1310 621 1315
rect 662 1312 667 1315
rect 690 1317 725 1318
rect 690 1312 691 1317
rect 696 1312 697 1317
rect 719 1312 720 1317
rect 724 1312 725 1317
rect 614 1309 621 1310
rect 661 1311 668 1312
rect 690 1311 697 1312
rect 706 1311 713 1312
rect 719 1311 725 1312
rect 735 1312 742 1313
rect 603 1305 610 1306
rect 637 1306 644 1307
rect 637 1305 638 1306
rect 604 1301 638 1305
rect 643 1301 644 1306
rect 661 1306 662 1311
rect 667 1306 668 1311
rect 661 1305 668 1306
rect 676 1307 683 1308
rect 604 1300 644 1301
rect 676 1301 677 1307
rect 682 1302 683 1307
rect 706 1306 707 1311
rect 712 1306 713 1311
rect 735 1307 736 1312
rect 741 1310 742 1312
rect 761 1310 768 1311
rect 841 1310 848 1311
rect 741 1307 762 1310
rect 735 1306 762 1307
rect 706 1305 713 1306
rect 736 1305 762 1306
rect 767 1305 768 1310
rect 707 1302 712 1305
rect 682 1301 712 1302
rect 676 1296 712 1301
rect 736 1279 741 1305
rect 761 1304 768 1305
rect 818 1305 842 1310
rect 847 1305 848 1310
rect 567 1273 741 1279
rect 567 1250 572 1273
rect 604 1251 644 1252
rect 566 1249 573 1250
rect 566 1244 567 1249
rect 572 1244 573 1249
rect 604 1247 638 1251
rect 566 1243 573 1244
rect 603 1246 610 1247
rect 603 1241 604 1246
rect 609 1241 610 1246
rect 637 1246 638 1247
rect 643 1246 644 1251
rect 676 1251 712 1256
rect 818 1254 823 1305
rect 841 1304 848 1305
rect 637 1245 644 1246
rect 661 1246 668 1247
rect 603 1240 610 1241
rect 614 1242 621 1243
rect 614 1237 615 1242
rect 620 1237 621 1242
rect 661 1241 662 1246
rect 667 1241 668 1246
rect 676 1245 677 1251
rect 682 1250 712 1251
rect 682 1245 683 1250
rect 707 1247 712 1250
rect 817 1253 824 1254
rect 817 1248 818 1253
rect 823 1248 824 1253
rect 817 1247 824 1248
rect 676 1244 683 1245
rect 706 1246 713 1247
rect 706 1241 707 1246
rect 712 1241 713 1246
rect 735 1245 742 1246
rect 661 1240 668 1241
rect 690 1240 697 1241
rect 706 1240 713 1241
rect 719 1240 725 1241
rect 662 1237 667 1240
rect 614 1232 667 1237
rect 690 1235 691 1240
rect 696 1235 697 1240
rect 719 1235 720 1240
rect 724 1235 725 1240
rect 690 1234 725 1235
rect 691 1230 725 1234
rect 735 1240 736 1245
rect 741 1240 742 1245
rect 735 1239 742 1240
rect 761 1239 768 1240
rect 735 1234 762 1239
rect 767 1234 768 1239
rect 880 1235 885 1344
rect 930 1306 937 1307
rect 930 1301 931 1306
rect 936 1301 937 1306
rect 930 1300 937 1301
rect 837 1234 885 1235
rect 735 1213 740 1234
rect 761 1233 768 1234
rect 568 1207 740 1213
rect 806 1229 885 1234
rect 931 1238 936 1300
rect 931 1232 998 1238
rect 568 1187 573 1207
rect 567 1186 574 1187
rect 567 1181 568 1186
rect 573 1181 574 1186
rect 567 1180 574 1181
rect 614 1183 667 1188
rect 691 1186 725 1190
rect 806 1186 811 1229
rect 603 1179 610 1180
rect 603 1174 604 1179
rect 609 1174 610 1179
rect 614 1178 615 1183
rect 620 1178 621 1183
rect 662 1180 667 1183
rect 690 1185 725 1186
rect 690 1180 691 1185
rect 696 1180 697 1185
rect 719 1180 720 1185
rect 724 1180 725 1185
rect 805 1185 812 1186
rect 614 1177 621 1178
rect 661 1179 668 1180
rect 690 1179 697 1180
rect 706 1179 713 1180
rect 719 1179 725 1180
rect 735 1180 742 1181
rect 603 1173 610 1174
rect 637 1174 644 1175
rect 637 1173 638 1174
rect 604 1169 638 1173
rect 643 1169 644 1174
rect 661 1174 662 1179
rect 667 1174 668 1179
rect 661 1173 668 1174
rect 676 1175 683 1176
rect 604 1168 644 1169
rect 676 1169 677 1175
rect 682 1170 683 1175
rect 706 1174 707 1179
rect 712 1174 713 1179
rect 735 1175 736 1180
rect 741 1175 742 1180
rect 805 1180 806 1185
rect 811 1180 812 1185
rect 875 1183 928 1188
rect 952 1186 986 1190
rect 993 1186 998 1232
rect 805 1179 812 1180
rect 864 1179 871 1180
rect 735 1174 742 1175
rect 760 1174 767 1175
rect 706 1173 713 1174
rect 707 1170 712 1173
rect 682 1169 712 1170
rect 737 1169 761 1174
rect 766 1169 767 1174
rect 864 1174 865 1179
rect 870 1174 871 1179
rect 875 1178 876 1183
rect 881 1178 882 1183
rect 923 1180 928 1183
rect 951 1185 986 1186
rect 951 1180 952 1185
rect 957 1180 958 1185
rect 980 1180 981 1185
rect 985 1180 986 1185
rect 875 1177 882 1178
rect 922 1179 929 1180
rect 951 1179 958 1180
rect 967 1179 974 1180
rect 980 1179 986 1180
rect 992 1185 999 1186
rect 992 1180 993 1185
rect 998 1180 999 1185
rect 992 1179 999 1180
rect 864 1173 871 1174
rect 898 1174 905 1175
rect 898 1173 899 1174
rect 676 1164 712 1169
rect 760 1168 767 1169
rect 865 1169 899 1173
rect 904 1169 905 1174
rect 922 1174 923 1179
rect 928 1174 929 1179
rect 922 1173 929 1174
rect 937 1175 944 1176
rect 865 1168 905 1169
rect 937 1169 938 1175
rect 943 1170 944 1175
rect 967 1174 968 1179
rect 973 1174 974 1179
rect 967 1173 974 1174
rect 968 1170 973 1173
rect 943 1169 973 1170
rect 937 1164 973 1169
rect 1020 1141 1025 1668
rect 1537 1647 1577 1648
rect 1537 1643 1571 1647
rect 1536 1642 1543 1643
rect 1536 1637 1537 1642
rect 1542 1637 1543 1642
rect 1570 1642 1571 1643
rect 1576 1642 1577 1647
rect 1609 1647 1645 1652
rect 1570 1641 1577 1642
rect 1594 1642 1601 1643
rect 1536 1636 1543 1637
rect 1547 1638 1554 1639
rect 1547 1633 1548 1638
rect 1553 1633 1554 1638
rect 1594 1637 1595 1642
rect 1600 1637 1601 1642
rect 1609 1641 1610 1647
rect 1615 1646 1645 1647
rect 1615 1641 1616 1646
rect 1640 1643 1645 1646
rect 1609 1640 1616 1641
rect 1639 1642 1646 1643
rect 1639 1637 1640 1642
rect 1645 1637 1646 1642
rect 1668 1641 1675 1642
rect 1594 1636 1601 1637
rect 1623 1636 1630 1637
rect 1639 1636 1646 1637
rect 1652 1636 1658 1637
rect 1595 1633 1600 1636
rect 1547 1628 1600 1633
rect 1623 1631 1624 1636
rect 1629 1631 1630 1636
rect 1652 1631 1653 1636
rect 1657 1631 1658 1636
rect 1623 1630 1658 1631
rect 1624 1626 1658 1630
rect 1668 1636 1669 1641
rect 1674 1636 1675 1641
rect 1750 1641 1757 1642
rect 1750 1636 1751 1641
rect 1756 1636 1757 1641
rect 1835 1641 1842 1642
rect 1835 1636 1836 1641
rect 1841 1636 1842 1641
rect 1668 1635 1675 1636
rect 1694 1635 1701 1636
rect 1750 1635 1757 1636
rect 1775 1635 1782 1636
rect 1835 1635 1842 1636
rect 1668 1630 1695 1635
rect 1700 1630 1701 1635
rect 1751 1630 1776 1635
rect 1781 1630 1782 1635
rect 1668 1609 1673 1630
rect 1694 1629 1701 1630
rect 1775 1629 1782 1630
rect 1832 1630 1841 1635
rect 1501 1603 1673 1609
rect 1284 1585 1290 1586
rect 1284 1581 1285 1585
rect 1289 1581 1422 1585
rect 1501 1583 1506 1603
rect 1284 1580 1422 1581
rect 1028 1185 1034 1186
rect 1028 1181 1029 1185
rect 1033 1181 1034 1185
rect 1028 1180 1034 1181
rect 867 1136 1025 1141
rect 867 1076 872 1136
rect 866 1075 872 1076
rect 866 1071 867 1075
rect 871 1071 872 1075
rect 866 1070 872 1071
rect 1029 1013 1034 1180
rect 992 1008 1034 1013
rect 992 994 997 1008
rect 991 993 997 994
rect 991 989 992 993
rect 996 989 997 993
rect 991 988 997 989
rect 1417 821 1422 1580
rect 1500 1582 1507 1583
rect 1500 1577 1501 1582
rect 1506 1577 1507 1582
rect 1500 1576 1507 1577
rect 1547 1579 1600 1584
rect 1624 1582 1658 1586
rect 1536 1575 1543 1576
rect 1536 1570 1537 1575
rect 1542 1570 1543 1575
rect 1547 1574 1548 1579
rect 1553 1574 1554 1579
rect 1595 1576 1600 1579
rect 1623 1581 1658 1582
rect 1623 1576 1624 1581
rect 1629 1576 1630 1581
rect 1652 1576 1653 1581
rect 1657 1576 1658 1581
rect 1547 1573 1554 1574
rect 1594 1575 1601 1576
rect 1623 1575 1630 1576
rect 1639 1575 1646 1576
rect 1652 1575 1658 1576
rect 1668 1576 1675 1577
rect 1694 1576 1701 1577
rect 1774 1576 1781 1577
rect 1536 1569 1543 1570
rect 1570 1570 1577 1571
rect 1570 1569 1571 1570
rect 1537 1565 1571 1569
rect 1576 1565 1577 1570
rect 1594 1570 1595 1575
rect 1600 1570 1601 1575
rect 1594 1569 1601 1570
rect 1609 1571 1616 1572
rect 1537 1564 1577 1565
rect 1609 1565 1610 1571
rect 1615 1566 1616 1571
rect 1639 1570 1640 1575
rect 1645 1570 1646 1575
rect 1668 1571 1669 1576
rect 1674 1571 1695 1576
rect 1700 1571 1701 1576
rect 1668 1570 1675 1571
rect 1694 1570 1701 1571
rect 1751 1571 1775 1576
rect 1780 1571 1781 1576
rect 1639 1569 1646 1570
rect 1640 1566 1645 1569
rect 1615 1565 1645 1566
rect 1609 1560 1645 1565
rect 1669 1543 1674 1570
rect 1500 1537 1674 1543
rect 1500 1514 1505 1537
rect 1537 1515 1577 1516
rect 1499 1513 1506 1514
rect 1499 1508 1500 1513
rect 1505 1508 1506 1513
rect 1537 1511 1571 1515
rect 1499 1507 1506 1508
rect 1536 1510 1543 1511
rect 1536 1505 1537 1510
rect 1542 1505 1543 1510
rect 1570 1510 1571 1511
rect 1576 1510 1577 1515
rect 1609 1515 1645 1520
rect 1751 1518 1756 1571
rect 1774 1570 1781 1571
rect 1832 1542 1837 1630
rect 1794 1537 1837 1542
rect 1570 1509 1577 1510
rect 1594 1510 1601 1511
rect 1536 1504 1543 1505
rect 1547 1506 1554 1507
rect 1547 1501 1548 1506
rect 1553 1501 1554 1506
rect 1594 1505 1595 1510
rect 1600 1505 1601 1510
rect 1609 1509 1610 1515
rect 1615 1514 1645 1515
rect 1615 1509 1616 1514
rect 1640 1511 1645 1514
rect 1750 1517 1757 1518
rect 1750 1512 1751 1517
rect 1756 1512 1757 1517
rect 1750 1511 1757 1512
rect 1609 1508 1616 1509
rect 1639 1510 1646 1511
rect 1639 1505 1640 1510
rect 1645 1505 1646 1510
rect 1668 1509 1675 1510
rect 1594 1504 1601 1505
rect 1623 1504 1630 1505
rect 1639 1504 1646 1505
rect 1652 1504 1658 1505
rect 1595 1501 1600 1504
rect 1547 1496 1600 1501
rect 1623 1499 1624 1504
rect 1629 1499 1630 1504
rect 1652 1499 1653 1504
rect 1657 1499 1658 1504
rect 1623 1498 1658 1499
rect 1624 1494 1658 1498
rect 1668 1504 1669 1509
rect 1674 1504 1675 1509
rect 1794 1504 1799 1537
rect 1857 1514 1864 1515
rect 1857 1509 1858 1514
rect 1863 1509 1864 1514
rect 1857 1508 1864 1509
rect 1668 1503 1675 1504
rect 1694 1503 1701 1504
rect 1668 1498 1695 1503
rect 1700 1498 1701 1503
rect 1794 1503 1806 1504
rect 1794 1498 1800 1503
rect 1805 1498 1806 1503
rect 1668 1477 1673 1498
rect 1694 1497 1701 1498
rect 1799 1497 1806 1498
rect 1501 1471 1673 1477
rect 1501 1451 1506 1471
rect 1500 1450 1507 1451
rect 1500 1445 1501 1450
rect 1506 1445 1507 1450
rect 1500 1444 1507 1445
rect 1547 1447 1600 1452
rect 1624 1450 1658 1454
rect 1536 1443 1543 1444
rect 1536 1438 1537 1443
rect 1542 1438 1543 1443
rect 1547 1442 1548 1447
rect 1553 1442 1554 1447
rect 1595 1444 1600 1447
rect 1623 1449 1658 1450
rect 1623 1444 1624 1449
rect 1629 1444 1630 1449
rect 1652 1444 1653 1449
rect 1657 1444 1658 1449
rect 1693 1445 1700 1446
rect 1799 1445 1806 1446
rect 1547 1441 1554 1442
rect 1594 1443 1601 1444
rect 1623 1443 1630 1444
rect 1639 1443 1646 1444
rect 1652 1443 1658 1444
rect 1668 1444 1694 1445
rect 1536 1437 1543 1438
rect 1570 1438 1577 1439
rect 1570 1437 1571 1438
rect 1537 1433 1571 1437
rect 1576 1433 1577 1438
rect 1594 1438 1595 1443
rect 1600 1438 1601 1443
rect 1594 1437 1601 1438
rect 1609 1439 1616 1440
rect 1537 1432 1577 1433
rect 1609 1433 1610 1439
rect 1615 1434 1616 1439
rect 1639 1438 1640 1443
rect 1645 1438 1646 1443
rect 1639 1437 1646 1438
rect 1668 1439 1669 1444
rect 1674 1440 1694 1444
rect 1699 1440 1700 1445
rect 1674 1439 1675 1440
rect 1693 1439 1700 1440
rect 1795 1440 1800 1445
rect 1805 1440 1806 1445
rect 1795 1439 1806 1440
rect 1668 1438 1675 1439
rect 1640 1434 1645 1437
rect 1615 1433 1645 1434
rect 1609 1428 1645 1433
rect 1668 1411 1673 1438
rect 1500 1405 1673 1411
rect 1795 1411 1800 1439
rect 1795 1406 1838 1411
rect 1500 1382 1505 1405
rect 1537 1383 1577 1384
rect 1499 1381 1506 1382
rect 1499 1376 1500 1381
rect 1505 1376 1506 1381
rect 1537 1379 1571 1383
rect 1499 1375 1506 1376
rect 1536 1378 1543 1379
rect 1536 1373 1537 1378
rect 1542 1373 1543 1378
rect 1570 1378 1571 1379
rect 1576 1378 1577 1383
rect 1609 1383 1645 1388
rect 1833 1387 1838 1406
rect 1570 1377 1577 1378
rect 1594 1378 1601 1379
rect 1536 1372 1543 1373
rect 1547 1374 1554 1375
rect 1547 1369 1548 1374
rect 1553 1369 1554 1374
rect 1594 1373 1595 1378
rect 1600 1373 1601 1378
rect 1609 1377 1610 1383
rect 1615 1382 1645 1383
rect 1615 1377 1616 1382
rect 1640 1379 1645 1382
rect 1832 1386 1839 1387
rect 1832 1381 1833 1386
rect 1838 1381 1839 1386
rect 1832 1380 1839 1381
rect 1858 1379 1863 1508
rect 1866 1379 1873 1380
rect 1609 1376 1616 1377
rect 1639 1378 1646 1379
rect 1639 1373 1640 1378
rect 1645 1373 1646 1378
rect 1668 1377 1675 1378
rect 1594 1372 1601 1373
rect 1623 1372 1630 1373
rect 1639 1372 1646 1373
rect 1652 1372 1658 1373
rect 1595 1369 1600 1372
rect 1547 1364 1600 1369
rect 1623 1367 1624 1372
rect 1629 1367 1630 1372
rect 1652 1367 1653 1372
rect 1657 1367 1658 1372
rect 1623 1366 1658 1367
rect 1624 1362 1658 1366
rect 1668 1372 1669 1377
rect 1674 1372 1675 1377
rect 1750 1377 1757 1378
rect 1750 1372 1751 1377
rect 1756 1372 1757 1377
rect 1846 1374 1867 1379
rect 1872 1374 1873 1379
rect 1846 1373 1858 1374
rect 1866 1373 1873 1374
rect 1668 1371 1675 1372
rect 1694 1371 1701 1372
rect 1750 1371 1757 1372
rect 1775 1371 1782 1372
rect 1668 1366 1695 1371
rect 1700 1366 1701 1371
rect 1751 1366 1776 1371
rect 1781 1366 1782 1371
rect 1668 1345 1673 1366
rect 1694 1365 1701 1366
rect 1775 1365 1782 1366
rect 1846 1365 1851 1373
rect 1501 1339 1673 1345
rect 1813 1344 1851 1365
rect 1501 1319 1506 1339
rect 1500 1318 1507 1319
rect 1500 1313 1501 1318
rect 1506 1313 1507 1318
rect 1500 1312 1507 1313
rect 1547 1315 1600 1320
rect 1624 1318 1658 1322
rect 1536 1311 1543 1312
rect 1536 1306 1537 1311
rect 1542 1306 1543 1311
rect 1547 1310 1548 1315
rect 1553 1310 1554 1315
rect 1595 1312 1600 1315
rect 1623 1317 1658 1318
rect 1623 1312 1624 1317
rect 1629 1312 1630 1317
rect 1652 1312 1653 1317
rect 1657 1312 1658 1317
rect 1547 1309 1554 1310
rect 1594 1311 1601 1312
rect 1623 1311 1630 1312
rect 1639 1311 1646 1312
rect 1652 1311 1658 1312
rect 1668 1312 1675 1313
rect 1536 1305 1543 1306
rect 1570 1306 1577 1307
rect 1570 1305 1571 1306
rect 1537 1301 1571 1305
rect 1576 1301 1577 1306
rect 1594 1306 1595 1311
rect 1600 1306 1601 1311
rect 1594 1305 1601 1306
rect 1609 1307 1616 1308
rect 1537 1300 1577 1301
rect 1609 1301 1610 1307
rect 1615 1302 1616 1307
rect 1639 1306 1640 1311
rect 1645 1306 1646 1311
rect 1668 1307 1669 1312
rect 1674 1310 1675 1312
rect 1694 1310 1701 1311
rect 1774 1310 1781 1311
rect 1674 1307 1695 1310
rect 1668 1306 1695 1307
rect 1639 1305 1646 1306
rect 1669 1305 1695 1306
rect 1700 1305 1701 1310
rect 1640 1302 1645 1305
rect 1615 1301 1645 1302
rect 1609 1296 1645 1301
rect 1669 1279 1674 1305
rect 1694 1304 1701 1305
rect 1751 1305 1775 1310
rect 1780 1305 1781 1310
rect 1500 1273 1674 1279
rect 1500 1250 1505 1273
rect 1537 1251 1577 1252
rect 1499 1249 1506 1250
rect 1499 1244 1500 1249
rect 1505 1244 1506 1249
rect 1537 1247 1571 1251
rect 1499 1243 1506 1244
rect 1536 1246 1543 1247
rect 1536 1241 1537 1246
rect 1542 1241 1543 1246
rect 1570 1246 1571 1247
rect 1576 1246 1577 1251
rect 1609 1251 1645 1256
rect 1751 1254 1756 1305
rect 1774 1304 1781 1305
rect 1570 1245 1577 1246
rect 1594 1246 1601 1247
rect 1536 1240 1543 1241
rect 1547 1242 1554 1243
rect 1547 1237 1548 1242
rect 1553 1237 1554 1242
rect 1594 1241 1595 1246
rect 1600 1241 1601 1246
rect 1609 1245 1610 1251
rect 1615 1250 1645 1251
rect 1615 1245 1616 1250
rect 1640 1247 1645 1250
rect 1750 1253 1757 1254
rect 1750 1248 1751 1253
rect 1756 1248 1757 1253
rect 1750 1247 1757 1248
rect 1609 1244 1616 1245
rect 1639 1246 1646 1247
rect 1639 1241 1640 1246
rect 1645 1241 1646 1246
rect 1668 1245 1675 1246
rect 1594 1240 1601 1241
rect 1623 1240 1630 1241
rect 1639 1240 1646 1241
rect 1652 1240 1658 1241
rect 1595 1237 1600 1240
rect 1547 1232 1600 1237
rect 1623 1235 1624 1240
rect 1629 1235 1630 1240
rect 1652 1235 1653 1240
rect 1657 1235 1658 1240
rect 1623 1234 1658 1235
rect 1624 1230 1658 1234
rect 1668 1240 1669 1245
rect 1674 1240 1675 1245
rect 1668 1239 1675 1240
rect 1694 1239 1701 1240
rect 1668 1234 1695 1239
rect 1700 1234 1701 1239
rect 1813 1235 1818 1344
rect 1863 1306 1870 1307
rect 1863 1301 1864 1306
rect 1869 1301 1870 1306
rect 1863 1300 1870 1301
rect 1770 1234 1818 1235
rect 1668 1213 1673 1234
rect 1694 1233 1701 1234
rect 1501 1207 1673 1213
rect 1739 1229 1818 1234
rect 1864 1238 1869 1300
rect 1864 1232 1931 1238
rect 1501 1187 1506 1207
rect 1500 1186 1507 1187
rect 1500 1181 1501 1186
rect 1506 1181 1507 1186
rect 1500 1180 1507 1181
rect 1547 1183 1600 1188
rect 1624 1186 1658 1190
rect 1739 1186 1744 1229
rect 1536 1179 1543 1180
rect 1536 1174 1537 1179
rect 1542 1174 1543 1179
rect 1547 1178 1548 1183
rect 1553 1178 1554 1183
rect 1595 1180 1600 1183
rect 1623 1185 1658 1186
rect 1623 1180 1624 1185
rect 1629 1180 1630 1185
rect 1652 1180 1653 1185
rect 1657 1180 1658 1185
rect 1738 1185 1745 1186
rect 1547 1177 1554 1178
rect 1594 1179 1601 1180
rect 1623 1179 1630 1180
rect 1639 1179 1646 1180
rect 1652 1179 1658 1180
rect 1668 1180 1675 1181
rect 1536 1173 1543 1174
rect 1570 1174 1577 1175
rect 1570 1173 1571 1174
rect 1537 1169 1571 1173
rect 1576 1169 1577 1174
rect 1594 1174 1595 1179
rect 1600 1174 1601 1179
rect 1594 1173 1601 1174
rect 1609 1175 1616 1176
rect 1537 1168 1577 1169
rect 1609 1169 1610 1175
rect 1615 1170 1616 1175
rect 1639 1174 1640 1179
rect 1645 1174 1646 1179
rect 1668 1175 1669 1180
rect 1674 1175 1675 1180
rect 1738 1180 1739 1185
rect 1744 1180 1745 1185
rect 1808 1183 1861 1188
rect 1885 1186 1919 1190
rect 1926 1186 1931 1232
rect 1738 1179 1745 1180
rect 1797 1179 1804 1180
rect 1668 1174 1675 1175
rect 1693 1174 1700 1175
rect 1639 1173 1646 1174
rect 1640 1170 1645 1173
rect 1615 1169 1645 1170
rect 1670 1169 1694 1174
rect 1699 1169 1700 1174
rect 1797 1174 1798 1179
rect 1803 1174 1804 1179
rect 1808 1178 1809 1183
rect 1814 1178 1815 1183
rect 1856 1180 1861 1183
rect 1884 1185 1919 1186
rect 1884 1180 1885 1185
rect 1890 1180 1891 1185
rect 1913 1180 1914 1185
rect 1918 1180 1919 1185
rect 1808 1177 1815 1178
rect 1855 1179 1862 1180
rect 1884 1179 1891 1180
rect 1900 1179 1907 1180
rect 1913 1179 1919 1180
rect 1925 1185 1932 1186
rect 1925 1180 1926 1185
rect 1931 1180 1932 1185
rect 1925 1179 1932 1180
rect 1797 1173 1804 1174
rect 1831 1174 1838 1175
rect 1831 1173 1832 1174
rect 1609 1164 1645 1169
rect 1693 1168 1700 1169
rect 1798 1169 1832 1173
rect 1837 1169 1838 1174
rect 1855 1174 1856 1179
rect 1861 1174 1862 1179
rect 1855 1173 1862 1174
rect 1870 1175 1877 1176
rect 1798 1168 1838 1169
rect 1870 1169 1871 1175
rect 1876 1170 1877 1175
rect 1900 1174 1901 1179
rect 1906 1174 1907 1179
rect 1900 1173 1907 1174
rect 1901 1170 1906 1173
rect 1876 1169 1906 1170
rect 1870 1164 1906 1169
rect 1953 1141 1958 1668
rect 1800 1136 1958 1141
rect 1800 1076 1805 1136
rect 1799 1075 1805 1076
rect 1799 1071 1800 1075
rect 1804 1071 1805 1075
rect 1799 1070 1805 1071
rect 1924 993 1930 994
rect 1924 989 1925 993
rect 1929 989 1930 993
rect 1924 988 1930 989
rect 484 820 490 821
rect 484 816 485 820
rect 489 816 490 820
rect 484 815 490 816
rect 1417 820 1423 821
rect 1417 816 1418 820
rect 1422 816 1423 820
rect 1417 815 1423 816
rect 1925 784 1930 988
rect 96 779 1930 784
rect 96 206 101 779
rect 563 744 569 745
rect 563 740 564 744
rect 568 740 569 744
rect 563 739 569 740
rect 1496 744 1502 745
rect 1496 740 1497 744
rect 1501 740 1502 744
rect 1496 739 1502 740
rect 563 709 568 739
rect 1496 709 1501 739
rect 352 708 568 709
rect 352 704 353 708
rect 357 704 568 708
rect 1285 708 1501 709
rect 1285 704 1286 708
rect 1290 704 1501 708
rect 352 703 358 704
rect 1285 703 1291 704
rect 1019 693 1025 694
rect 1019 689 1020 693
rect 1024 689 1025 693
rect 1019 688 1025 689
rect 1952 693 1958 694
rect 1952 689 1953 693
rect 1957 689 1958 693
rect 1952 688 1958 689
rect 604 667 644 668
rect 604 663 638 667
rect 603 662 610 663
rect 603 657 604 662
rect 609 657 610 662
rect 637 662 638 663
rect 643 662 644 667
rect 676 667 712 672
rect 637 661 644 662
rect 661 662 668 663
rect 603 656 610 657
rect 614 658 621 659
rect 614 653 615 658
rect 620 653 621 658
rect 661 657 662 662
rect 667 657 668 662
rect 676 661 677 667
rect 682 666 712 667
rect 682 661 683 666
rect 707 663 712 666
rect 676 660 683 661
rect 706 662 713 663
rect 706 657 707 662
rect 712 657 713 662
rect 735 661 742 662
rect 661 656 668 657
rect 690 656 697 657
rect 706 656 713 657
rect 719 656 725 657
rect 662 653 667 656
rect 614 648 667 653
rect 690 651 691 656
rect 696 651 697 656
rect 719 651 720 656
rect 724 651 725 656
rect 690 650 725 651
rect 691 646 725 650
rect 735 656 736 661
rect 741 656 742 661
rect 817 661 824 662
rect 817 656 818 661
rect 823 656 824 661
rect 902 661 909 662
rect 902 656 903 661
rect 908 656 909 661
rect 735 655 742 656
rect 761 655 768 656
rect 817 655 824 656
rect 842 655 849 656
rect 902 655 909 656
rect 735 650 762 655
rect 767 650 768 655
rect 818 650 843 655
rect 848 650 849 655
rect 735 629 740 650
rect 761 649 768 650
rect 842 649 849 650
rect 899 650 908 655
rect 568 623 740 629
rect 351 605 357 606
rect 351 601 352 605
rect 356 601 489 605
rect 568 603 573 623
rect 351 600 489 601
rect 95 205 101 206
rect 95 201 96 205
rect 100 201 101 205
rect 95 200 101 201
rect 484 -159 489 600
rect 567 602 574 603
rect 567 597 568 602
rect 573 597 574 602
rect 567 596 574 597
rect 614 599 667 604
rect 691 602 725 606
rect 603 595 610 596
rect 603 590 604 595
rect 609 590 610 595
rect 614 594 615 599
rect 620 594 621 599
rect 662 596 667 599
rect 690 601 725 602
rect 690 596 691 601
rect 696 596 697 601
rect 719 596 720 601
rect 724 596 725 601
rect 614 593 621 594
rect 661 595 668 596
rect 690 595 697 596
rect 706 595 713 596
rect 719 595 725 596
rect 735 596 742 597
rect 761 596 768 597
rect 841 596 848 597
rect 603 589 610 590
rect 637 590 644 591
rect 637 589 638 590
rect 604 585 638 589
rect 643 585 644 590
rect 661 590 662 595
rect 667 590 668 595
rect 661 589 668 590
rect 676 591 683 592
rect 604 584 644 585
rect 676 585 677 591
rect 682 586 683 591
rect 706 590 707 595
rect 712 590 713 595
rect 735 591 736 596
rect 741 591 762 596
rect 767 591 768 596
rect 735 590 742 591
rect 761 590 768 591
rect 818 591 842 596
rect 847 591 848 596
rect 706 589 713 590
rect 707 586 712 589
rect 682 585 712 586
rect 676 580 712 585
rect 736 563 741 590
rect 567 557 741 563
rect 567 534 572 557
rect 604 535 644 536
rect 566 533 573 534
rect 566 528 567 533
rect 572 528 573 533
rect 604 531 638 535
rect 566 527 573 528
rect 603 530 610 531
rect 603 525 604 530
rect 609 525 610 530
rect 637 530 638 531
rect 643 530 644 535
rect 676 535 712 540
rect 818 538 823 591
rect 841 590 848 591
rect 899 562 904 650
rect 861 557 904 562
rect 637 529 644 530
rect 661 530 668 531
rect 603 524 610 525
rect 614 526 621 527
rect 614 521 615 526
rect 620 521 621 526
rect 661 525 662 530
rect 667 525 668 530
rect 676 529 677 535
rect 682 534 712 535
rect 682 529 683 534
rect 707 531 712 534
rect 817 537 824 538
rect 817 532 818 537
rect 823 532 824 537
rect 817 531 824 532
rect 676 528 683 529
rect 706 530 713 531
rect 706 525 707 530
rect 712 525 713 530
rect 735 529 742 530
rect 661 524 668 525
rect 690 524 697 525
rect 706 524 713 525
rect 719 524 725 525
rect 662 521 667 524
rect 614 516 667 521
rect 690 519 691 524
rect 696 519 697 524
rect 719 519 720 524
rect 724 519 725 524
rect 690 518 725 519
rect 691 514 725 518
rect 735 524 736 529
rect 741 524 742 529
rect 861 524 866 557
rect 924 534 931 535
rect 924 529 925 534
rect 930 529 931 534
rect 924 528 931 529
rect 735 523 742 524
rect 761 523 768 524
rect 735 518 762 523
rect 767 518 768 523
rect 861 523 873 524
rect 861 518 867 523
rect 872 518 873 523
rect 735 497 740 518
rect 761 517 768 518
rect 866 517 873 518
rect 568 491 740 497
rect 568 471 573 491
rect 567 470 574 471
rect 567 465 568 470
rect 573 465 574 470
rect 567 464 574 465
rect 614 467 667 472
rect 691 470 725 474
rect 603 463 610 464
rect 603 458 604 463
rect 609 458 610 463
rect 614 462 615 467
rect 620 462 621 467
rect 662 464 667 467
rect 690 469 725 470
rect 690 464 691 469
rect 696 464 697 469
rect 719 464 720 469
rect 724 464 725 469
rect 760 465 767 466
rect 866 465 873 466
rect 614 461 621 462
rect 661 463 668 464
rect 690 463 697 464
rect 706 463 713 464
rect 719 463 725 464
rect 735 464 761 465
rect 603 457 610 458
rect 637 458 644 459
rect 637 457 638 458
rect 604 453 638 457
rect 643 453 644 458
rect 661 458 662 463
rect 667 458 668 463
rect 661 457 668 458
rect 676 459 683 460
rect 604 452 644 453
rect 676 453 677 459
rect 682 454 683 459
rect 706 458 707 463
rect 712 458 713 463
rect 706 457 713 458
rect 735 459 736 464
rect 741 460 761 464
rect 766 460 767 465
rect 741 459 742 460
rect 760 459 767 460
rect 862 460 867 465
rect 872 460 873 465
rect 862 459 873 460
rect 735 458 742 459
rect 707 454 712 457
rect 682 453 712 454
rect 676 448 712 453
rect 735 431 740 458
rect 567 425 740 431
rect 862 431 867 459
rect 862 426 905 431
rect 567 402 572 425
rect 604 403 644 404
rect 566 401 573 402
rect 566 396 567 401
rect 572 396 573 401
rect 604 399 638 403
rect 566 395 573 396
rect 603 398 610 399
rect 603 393 604 398
rect 609 393 610 398
rect 637 398 638 399
rect 643 398 644 403
rect 676 403 712 408
rect 900 407 905 426
rect 637 397 644 398
rect 661 398 668 399
rect 603 392 610 393
rect 614 394 621 395
rect 614 389 615 394
rect 620 389 621 394
rect 661 393 662 398
rect 667 393 668 398
rect 676 397 677 403
rect 682 402 712 403
rect 682 397 683 402
rect 707 399 712 402
rect 899 406 906 407
rect 899 401 900 406
rect 905 401 906 406
rect 899 400 906 401
rect 925 399 930 528
rect 933 399 940 400
rect 676 396 683 397
rect 706 398 713 399
rect 706 393 707 398
rect 712 393 713 398
rect 735 397 742 398
rect 661 392 668 393
rect 690 392 697 393
rect 706 392 713 393
rect 719 392 725 393
rect 662 389 667 392
rect 614 384 667 389
rect 690 387 691 392
rect 696 387 697 392
rect 719 387 720 392
rect 724 387 725 392
rect 690 386 725 387
rect 691 382 725 386
rect 735 392 736 397
rect 741 392 742 397
rect 817 397 824 398
rect 817 392 818 397
rect 823 392 824 397
rect 913 394 934 399
rect 939 394 940 399
rect 913 393 925 394
rect 933 393 940 394
rect 735 391 742 392
rect 761 391 768 392
rect 817 391 824 392
rect 842 391 849 392
rect 735 386 762 391
rect 767 386 768 391
rect 818 386 843 391
rect 848 386 849 391
rect 735 365 740 386
rect 761 385 768 386
rect 842 385 849 386
rect 913 385 918 393
rect 568 359 740 365
rect 880 364 918 385
rect 568 339 573 359
rect 567 338 574 339
rect 567 333 568 338
rect 573 333 574 338
rect 567 332 574 333
rect 614 335 667 340
rect 691 338 725 342
rect 603 331 610 332
rect 603 326 604 331
rect 609 326 610 331
rect 614 330 615 335
rect 620 330 621 335
rect 662 332 667 335
rect 690 337 725 338
rect 690 332 691 337
rect 696 332 697 337
rect 719 332 720 337
rect 724 332 725 337
rect 614 329 621 330
rect 661 331 668 332
rect 690 331 697 332
rect 706 331 713 332
rect 719 331 725 332
rect 735 332 742 333
rect 603 325 610 326
rect 637 326 644 327
rect 637 325 638 326
rect 604 321 638 325
rect 643 321 644 326
rect 661 326 662 331
rect 667 326 668 331
rect 661 325 668 326
rect 676 327 683 328
rect 604 320 644 321
rect 676 321 677 327
rect 682 322 683 327
rect 706 326 707 331
rect 712 326 713 331
rect 735 327 736 332
rect 741 330 742 332
rect 761 330 768 331
rect 841 330 848 331
rect 741 327 762 330
rect 735 326 762 327
rect 706 325 713 326
rect 736 325 762 326
rect 767 325 768 330
rect 707 322 712 325
rect 682 321 712 322
rect 676 316 712 321
rect 736 299 741 325
rect 761 324 768 325
rect 818 325 842 330
rect 847 325 848 330
rect 567 293 741 299
rect 567 270 572 293
rect 604 271 644 272
rect 566 269 573 270
rect 566 264 567 269
rect 572 264 573 269
rect 604 267 638 271
rect 566 263 573 264
rect 603 266 610 267
rect 603 261 604 266
rect 609 261 610 266
rect 637 266 638 267
rect 643 266 644 271
rect 676 271 712 276
rect 818 274 823 325
rect 841 324 848 325
rect 637 265 644 266
rect 661 266 668 267
rect 603 260 610 261
rect 614 262 621 263
rect 614 257 615 262
rect 620 257 621 262
rect 661 261 662 266
rect 667 261 668 266
rect 676 265 677 271
rect 682 270 712 271
rect 682 265 683 270
rect 707 267 712 270
rect 817 273 824 274
rect 817 268 818 273
rect 823 268 824 273
rect 817 267 824 268
rect 676 264 683 265
rect 706 266 713 267
rect 706 261 707 266
rect 712 261 713 266
rect 735 265 742 266
rect 661 260 668 261
rect 690 260 697 261
rect 706 260 713 261
rect 719 260 725 261
rect 662 257 667 260
rect 614 252 667 257
rect 690 255 691 260
rect 696 255 697 260
rect 719 255 720 260
rect 724 255 725 260
rect 690 254 725 255
rect 691 250 725 254
rect 735 260 736 265
rect 741 260 742 265
rect 735 259 742 260
rect 761 259 768 260
rect 735 254 762 259
rect 767 254 768 259
rect 880 255 885 364
rect 930 326 937 327
rect 930 321 931 326
rect 936 321 937 326
rect 930 320 937 321
rect 837 254 885 255
rect 735 233 740 254
rect 761 253 768 254
rect 568 227 740 233
rect 806 249 885 254
rect 931 258 936 320
rect 931 252 998 258
rect 568 207 573 227
rect 567 206 574 207
rect 567 201 568 206
rect 573 201 574 206
rect 567 200 574 201
rect 614 203 667 208
rect 691 206 725 210
rect 806 206 811 249
rect 603 199 610 200
rect 603 194 604 199
rect 609 194 610 199
rect 614 198 615 203
rect 620 198 621 203
rect 662 200 667 203
rect 690 205 725 206
rect 690 200 691 205
rect 696 200 697 205
rect 719 200 720 205
rect 724 200 725 205
rect 805 205 812 206
rect 614 197 621 198
rect 661 199 668 200
rect 690 199 697 200
rect 706 199 713 200
rect 719 199 725 200
rect 735 200 742 201
rect 603 193 610 194
rect 637 194 644 195
rect 637 193 638 194
rect 604 189 638 193
rect 643 189 644 194
rect 661 194 662 199
rect 667 194 668 199
rect 661 193 668 194
rect 676 195 683 196
rect 604 188 644 189
rect 676 189 677 195
rect 682 190 683 195
rect 706 194 707 199
rect 712 194 713 199
rect 735 195 736 200
rect 741 195 742 200
rect 805 200 806 205
rect 811 200 812 205
rect 875 203 928 208
rect 952 206 986 210
rect 993 206 998 252
rect 805 199 812 200
rect 864 199 871 200
rect 735 194 742 195
rect 760 194 767 195
rect 706 193 713 194
rect 707 190 712 193
rect 682 189 712 190
rect 737 189 761 194
rect 766 189 767 194
rect 864 194 865 199
rect 870 194 871 199
rect 875 198 876 203
rect 881 198 882 203
rect 923 200 928 203
rect 951 205 986 206
rect 951 200 952 205
rect 957 200 958 205
rect 980 200 981 205
rect 985 200 986 205
rect 875 197 882 198
rect 922 199 929 200
rect 951 199 958 200
rect 967 199 974 200
rect 980 199 986 200
rect 992 205 999 206
rect 992 200 993 205
rect 998 200 999 205
rect 992 199 999 200
rect 864 193 871 194
rect 898 194 905 195
rect 898 193 899 194
rect 676 184 712 189
rect 760 188 767 189
rect 865 189 899 193
rect 904 189 905 194
rect 922 194 923 199
rect 928 194 929 199
rect 922 193 929 194
rect 937 195 944 196
rect 865 188 905 189
rect 937 189 938 195
rect 943 190 944 195
rect 967 194 968 199
rect 973 194 974 199
rect 967 193 974 194
rect 968 190 973 193
rect 943 189 973 190
rect 937 184 973 189
rect 1020 161 1025 688
rect 1537 667 1577 668
rect 1537 663 1571 667
rect 1536 662 1543 663
rect 1536 657 1537 662
rect 1542 657 1543 662
rect 1570 662 1571 663
rect 1576 662 1577 667
rect 1609 667 1645 672
rect 1570 661 1577 662
rect 1594 662 1601 663
rect 1536 656 1543 657
rect 1547 658 1554 659
rect 1547 653 1548 658
rect 1553 653 1554 658
rect 1594 657 1595 662
rect 1600 657 1601 662
rect 1609 661 1610 667
rect 1615 666 1645 667
rect 1615 661 1616 666
rect 1640 663 1645 666
rect 1609 660 1616 661
rect 1639 662 1646 663
rect 1639 657 1640 662
rect 1645 657 1646 662
rect 1668 661 1675 662
rect 1594 656 1601 657
rect 1623 656 1630 657
rect 1639 656 1646 657
rect 1652 656 1658 657
rect 1595 653 1600 656
rect 1547 648 1600 653
rect 1623 651 1624 656
rect 1629 651 1630 656
rect 1652 651 1653 656
rect 1657 651 1658 656
rect 1623 650 1658 651
rect 1624 646 1658 650
rect 1668 656 1669 661
rect 1674 656 1675 661
rect 1750 661 1757 662
rect 1750 656 1751 661
rect 1756 656 1757 661
rect 1835 661 1842 662
rect 1835 656 1836 661
rect 1841 656 1842 661
rect 1668 655 1675 656
rect 1694 655 1701 656
rect 1750 655 1757 656
rect 1775 655 1782 656
rect 1835 655 1842 656
rect 1668 650 1695 655
rect 1700 650 1701 655
rect 1751 650 1776 655
rect 1781 650 1782 655
rect 1668 629 1673 650
rect 1694 649 1701 650
rect 1775 649 1782 650
rect 1832 650 1841 655
rect 1501 623 1673 629
rect 1284 605 1290 606
rect 1284 601 1285 605
rect 1289 601 1422 605
rect 1501 603 1506 623
rect 1284 600 1422 601
rect 1028 205 1034 206
rect 1028 201 1029 205
rect 1033 201 1034 205
rect 1028 200 1034 201
rect 867 156 1025 161
rect 867 96 872 156
rect 866 95 872 96
rect 866 91 867 95
rect 871 91 872 95
rect 866 90 872 91
rect 1029 33 1034 200
rect 992 28 1034 33
rect 992 14 997 28
rect 991 13 997 14
rect 991 9 992 13
rect 996 9 997 13
rect 991 8 997 9
rect 1417 -159 1422 600
rect 1500 602 1507 603
rect 1500 597 1501 602
rect 1506 597 1507 602
rect 1500 596 1507 597
rect 1547 599 1600 604
rect 1624 602 1658 606
rect 1536 595 1543 596
rect 1536 590 1537 595
rect 1542 590 1543 595
rect 1547 594 1548 599
rect 1553 594 1554 599
rect 1595 596 1600 599
rect 1623 601 1658 602
rect 1623 596 1624 601
rect 1629 596 1630 601
rect 1652 596 1653 601
rect 1657 596 1658 601
rect 1547 593 1554 594
rect 1594 595 1601 596
rect 1623 595 1630 596
rect 1639 595 1646 596
rect 1652 595 1658 596
rect 1668 596 1675 597
rect 1694 596 1701 597
rect 1774 596 1781 597
rect 1536 589 1543 590
rect 1570 590 1577 591
rect 1570 589 1571 590
rect 1537 585 1571 589
rect 1576 585 1577 590
rect 1594 590 1595 595
rect 1600 590 1601 595
rect 1594 589 1601 590
rect 1609 591 1616 592
rect 1537 584 1577 585
rect 1609 585 1610 591
rect 1615 586 1616 591
rect 1639 590 1640 595
rect 1645 590 1646 595
rect 1668 591 1669 596
rect 1674 591 1695 596
rect 1700 591 1701 596
rect 1668 590 1675 591
rect 1694 590 1701 591
rect 1751 591 1775 596
rect 1780 591 1781 596
rect 1639 589 1646 590
rect 1640 586 1645 589
rect 1615 585 1645 586
rect 1609 580 1645 585
rect 1669 563 1674 590
rect 1500 557 1674 563
rect 1500 534 1505 557
rect 1537 535 1577 536
rect 1499 533 1506 534
rect 1499 528 1500 533
rect 1505 528 1506 533
rect 1537 531 1571 535
rect 1499 527 1506 528
rect 1536 530 1543 531
rect 1536 525 1537 530
rect 1542 525 1543 530
rect 1570 530 1571 531
rect 1576 530 1577 535
rect 1609 535 1645 540
rect 1751 538 1756 591
rect 1774 590 1781 591
rect 1832 562 1837 650
rect 1794 557 1837 562
rect 1570 529 1577 530
rect 1594 530 1601 531
rect 1536 524 1543 525
rect 1547 526 1554 527
rect 1547 521 1548 526
rect 1553 521 1554 526
rect 1594 525 1595 530
rect 1600 525 1601 530
rect 1609 529 1610 535
rect 1615 534 1645 535
rect 1615 529 1616 534
rect 1640 531 1645 534
rect 1750 537 1757 538
rect 1750 532 1751 537
rect 1756 532 1757 537
rect 1750 531 1757 532
rect 1609 528 1616 529
rect 1639 530 1646 531
rect 1639 525 1640 530
rect 1645 525 1646 530
rect 1668 529 1675 530
rect 1594 524 1601 525
rect 1623 524 1630 525
rect 1639 524 1646 525
rect 1652 524 1658 525
rect 1595 521 1600 524
rect 1547 516 1600 521
rect 1623 519 1624 524
rect 1629 519 1630 524
rect 1652 519 1653 524
rect 1657 519 1658 524
rect 1623 518 1658 519
rect 1624 514 1658 518
rect 1668 524 1669 529
rect 1674 524 1675 529
rect 1794 524 1799 557
rect 1857 534 1864 535
rect 1857 529 1858 534
rect 1863 529 1864 534
rect 1857 528 1864 529
rect 1668 523 1675 524
rect 1694 523 1701 524
rect 1668 518 1695 523
rect 1700 518 1701 523
rect 1794 523 1806 524
rect 1794 518 1800 523
rect 1805 518 1806 523
rect 1668 497 1673 518
rect 1694 517 1701 518
rect 1799 517 1806 518
rect 1501 491 1673 497
rect 1501 471 1506 491
rect 1500 470 1507 471
rect 1500 465 1501 470
rect 1506 465 1507 470
rect 1500 464 1507 465
rect 1547 467 1600 472
rect 1624 470 1658 474
rect 1536 463 1543 464
rect 1536 458 1537 463
rect 1542 458 1543 463
rect 1547 462 1548 467
rect 1553 462 1554 467
rect 1595 464 1600 467
rect 1623 469 1658 470
rect 1623 464 1624 469
rect 1629 464 1630 469
rect 1652 464 1653 469
rect 1657 464 1658 469
rect 1693 465 1700 466
rect 1799 465 1806 466
rect 1547 461 1554 462
rect 1594 463 1601 464
rect 1623 463 1630 464
rect 1639 463 1646 464
rect 1652 463 1658 464
rect 1668 464 1694 465
rect 1536 457 1543 458
rect 1570 458 1577 459
rect 1570 457 1571 458
rect 1537 453 1571 457
rect 1576 453 1577 458
rect 1594 458 1595 463
rect 1600 458 1601 463
rect 1594 457 1601 458
rect 1609 459 1616 460
rect 1537 452 1577 453
rect 1609 453 1610 459
rect 1615 454 1616 459
rect 1639 458 1640 463
rect 1645 458 1646 463
rect 1639 457 1646 458
rect 1668 459 1669 464
rect 1674 460 1694 464
rect 1699 460 1700 465
rect 1674 459 1675 460
rect 1693 459 1700 460
rect 1795 460 1800 465
rect 1805 460 1806 465
rect 1795 459 1806 460
rect 1668 458 1675 459
rect 1640 454 1645 457
rect 1615 453 1645 454
rect 1609 448 1645 453
rect 1668 431 1673 458
rect 1500 425 1673 431
rect 1795 431 1800 459
rect 1795 426 1838 431
rect 1500 402 1505 425
rect 1537 403 1577 404
rect 1499 401 1506 402
rect 1499 396 1500 401
rect 1505 396 1506 401
rect 1537 399 1571 403
rect 1499 395 1506 396
rect 1536 398 1543 399
rect 1536 393 1537 398
rect 1542 393 1543 398
rect 1570 398 1571 399
rect 1576 398 1577 403
rect 1609 403 1645 408
rect 1833 407 1838 426
rect 1570 397 1577 398
rect 1594 398 1601 399
rect 1536 392 1543 393
rect 1547 394 1554 395
rect 1547 389 1548 394
rect 1553 389 1554 394
rect 1594 393 1595 398
rect 1600 393 1601 398
rect 1609 397 1610 403
rect 1615 402 1645 403
rect 1615 397 1616 402
rect 1640 399 1645 402
rect 1832 406 1839 407
rect 1832 401 1833 406
rect 1838 401 1839 406
rect 1832 400 1839 401
rect 1858 399 1863 528
rect 1866 399 1873 400
rect 1609 396 1616 397
rect 1639 398 1646 399
rect 1639 393 1640 398
rect 1645 393 1646 398
rect 1668 397 1675 398
rect 1594 392 1601 393
rect 1623 392 1630 393
rect 1639 392 1646 393
rect 1652 392 1658 393
rect 1595 389 1600 392
rect 1547 384 1600 389
rect 1623 387 1624 392
rect 1629 387 1630 392
rect 1652 387 1653 392
rect 1657 387 1658 392
rect 1623 386 1658 387
rect 1624 382 1658 386
rect 1668 392 1669 397
rect 1674 392 1675 397
rect 1750 397 1757 398
rect 1750 392 1751 397
rect 1756 392 1757 397
rect 1846 394 1867 399
rect 1872 394 1873 399
rect 1846 393 1858 394
rect 1866 393 1873 394
rect 1668 391 1675 392
rect 1694 391 1701 392
rect 1750 391 1757 392
rect 1775 391 1782 392
rect 1668 386 1695 391
rect 1700 386 1701 391
rect 1751 386 1776 391
rect 1781 386 1782 391
rect 1668 365 1673 386
rect 1694 385 1701 386
rect 1775 385 1782 386
rect 1846 385 1851 393
rect 1501 359 1673 365
rect 1813 364 1851 385
rect 1501 339 1506 359
rect 1500 338 1507 339
rect 1500 333 1501 338
rect 1506 333 1507 338
rect 1500 332 1507 333
rect 1547 335 1600 340
rect 1624 338 1658 342
rect 1536 331 1543 332
rect 1536 326 1537 331
rect 1542 326 1543 331
rect 1547 330 1548 335
rect 1553 330 1554 335
rect 1595 332 1600 335
rect 1623 337 1658 338
rect 1623 332 1624 337
rect 1629 332 1630 337
rect 1652 332 1653 337
rect 1657 332 1658 337
rect 1547 329 1554 330
rect 1594 331 1601 332
rect 1623 331 1630 332
rect 1639 331 1646 332
rect 1652 331 1658 332
rect 1668 332 1675 333
rect 1536 325 1543 326
rect 1570 326 1577 327
rect 1570 325 1571 326
rect 1537 321 1571 325
rect 1576 321 1577 326
rect 1594 326 1595 331
rect 1600 326 1601 331
rect 1594 325 1601 326
rect 1609 327 1616 328
rect 1537 320 1577 321
rect 1609 321 1610 327
rect 1615 322 1616 327
rect 1639 326 1640 331
rect 1645 326 1646 331
rect 1668 327 1669 332
rect 1674 330 1675 332
rect 1694 330 1701 331
rect 1774 330 1781 331
rect 1674 327 1695 330
rect 1668 326 1695 327
rect 1639 325 1646 326
rect 1669 325 1695 326
rect 1700 325 1701 330
rect 1640 322 1645 325
rect 1615 321 1645 322
rect 1609 316 1645 321
rect 1669 299 1674 325
rect 1694 324 1701 325
rect 1751 325 1775 330
rect 1780 325 1781 330
rect 1500 293 1674 299
rect 1500 270 1505 293
rect 1537 271 1577 272
rect 1499 269 1506 270
rect 1499 264 1500 269
rect 1505 264 1506 269
rect 1537 267 1571 271
rect 1499 263 1506 264
rect 1536 266 1543 267
rect 1536 261 1537 266
rect 1542 261 1543 266
rect 1570 266 1571 267
rect 1576 266 1577 271
rect 1609 271 1645 276
rect 1751 274 1756 325
rect 1774 324 1781 325
rect 1570 265 1577 266
rect 1594 266 1601 267
rect 1536 260 1543 261
rect 1547 262 1554 263
rect 1547 257 1548 262
rect 1553 257 1554 262
rect 1594 261 1595 266
rect 1600 261 1601 266
rect 1609 265 1610 271
rect 1615 270 1645 271
rect 1615 265 1616 270
rect 1640 267 1645 270
rect 1750 273 1757 274
rect 1750 268 1751 273
rect 1756 268 1757 273
rect 1750 267 1757 268
rect 1609 264 1616 265
rect 1639 266 1646 267
rect 1639 261 1640 266
rect 1645 261 1646 266
rect 1668 265 1675 266
rect 1594 260 1601 261
rect 1623 260 1630 261
rect 1639 260 1646 261
rect 1652 260 1658 261
rect 1595 257 1600 260
rect 1547 252 1600 257
rect 1623 255 1624 260
rect 1629 255 1630 260
rect 1652 255 1653 260
rect 1657 255 1658 260
rect 1623 254 1658 255
rect 1624 250 1658 254
rect 1668 260 1669 265
rect 1674 260 1675 265
rect 1668 259 1675 260
rect 1694 259 1701 260
rect 1668 254 1695 259
rect 1700 254 1701 259
rect 1813 255 1818 364
rect 1863 326 1870 327
rect 1863 321 1864 326
rect 1869 321 1870 326
rect 1863 320 1870 321
rect 1770 254 1818 255
rect 1668 233 1673 254
rect 1694 253 1701 254
rect 1501 227 1673 233
rect 1739 249 1818 254
rect 1864 258 1869 320
rect 1864 252 1931 258
rect 1501 207 1506 227
rect 1500 206 1507 207
rect 1500 201 1501 206
rect 1506 201 1507 206
rect 1500 200 1507 201
rect 1547 203 1600 208
rect 1624 206 1658 210
rect 1739 206 1744 249
rect 1536 199 1543 200
rect 1536 194 1537 199
rect 1542 194 1543 199
rect 1547 198 1548 203
rect 1553 198 1554 203
rect 1595 200 1600 203
rect 1623 205 1658 206
rect 1623 200 1624 205
rect 1629 200 1630 205
rect 1652 200 1653 205
rect 1657 200 1658 205
rect 1738 205 1745 206
rect 1547 197 1554 198
rect 1594 199 1601 200
rect 1623 199 1630 200
rect 1639 199 1646 200
rect 1652 199 1658 200
rect 1668 200 1675 201
rect 1536 193 1543 194
rect 1570 194 1577 195
rect 1570 193 1571 194
rect 1537 189 1571 193
rect 1576 189 1577 194
rect 1594 194 1595 199
rect 1600 194 1601 199
rect 1594 193 1601 194
rect 1609 195 1616 196
rect 1537 188 1577 189
rect 1609 189 1610 195
rect 1615 190 1616 195
rect 1639 194 1640 199
rect 1645 194 1646 199
rect 1668 195 1669 200
rect 1674 195 1675 200
rect 1738 200 1739 205
rect 1744 200 1745 205
rect 1808 203 1861 208
rect 1885 206 1919 210
rect 1926 206 1931 252
rect 1738 199 1745 200
rect 1797 199 1804 200
rect 1668 194 1675 195
rect 1693 194 1700 195
rect 1639 193 1646 194
rect 1640 190 1645 193
rect 1615 189 1645 190
rect 1670 189 1694 194
rect 1699 189 1700 194
rect 1797 194 1798 199
rect 1803 194 1804 199
rect 1808 198 1809 203
rect 1814 198 1815 203
rect 1856 200 1861 203
rect 1884 205 1919 206
rect 1884 200 1885 205
rect 1890 200 1891 205
rect 1913 200 1914 205
rect 1918 200 1919 205
rect 1808 197 1815 198
rect 1855 199 1862 200
rect 1884 199 1891 200
rect 1900 199 1907 200
rect 1913 199 1919 200
rect 1925 205 1932 206
rect 1925 200 1926 205
rect 1931 200 1932 205
rect 1925 199 1932 200
rect 1797 193 1804 194
rect 1831 194 1838 195
rect 1831 193 1832 194
rect 1609 184 1645 189
rect 1693 188 1700 189
rect 1798 189 1832 193
rect 1837 189 1838 194
rect 1855 194 1856 199
rect 1861 194 1862 199
rect 1855 193 1862 194
rect 1870 195 1877 196
rect 1798 188 1838 189
rect 1870 189 1871 195
rect 1876 190 1877 195
rect 1900 194 1901 199
rect 1906 194 1907 199
rect 1900 193 1907 194
rect 1901 190 1906 193
rect 1876 189 1906 190
rect 1870 184 1906 189
rect 1953 161 1958 688
rect 1800 156 1958 161
rect 1971 205 2027 210
rect 1800 96 1805 156
rect 1799 95 1805 96
rect 1799 91 1800 95
rect 1804 91 1805 95
rect 1799 90 1805 91
rect 1971 33 1976 205
rect 1925 28 1976 33
rect 1925 14 1930 28
rect 1924 13 1930 14
rect 1924 9 1925 13
rect 1929 9 1930 13
rect 1924 8 1930 9
rect 484 -160 490 -159
rect 484 -164 485 -160
rect 489 -164 490 -160
rect 484 -165 490 -164
rect 1417 -160 1423 -159
rect 1417 -164 1418 -160
rect 1422 -164 1423 -160
rect 1417 -165 1423 -164
<< labels >>
rlabel metal1 96 232 99 236 1 Vdd!
rlabel metal1 97 175 100 179 1 GND!
rlabel metal1 98 168 101 172 2 ~clk
rlabel metal1 96 239 99 243 4 clk
rlabel metal1 228 232 231 236 1 Vdd!
rlabel metal1 229 175 232 179 1 GND!
rlabel metal1 230 168 233 172 2 ~clk
rlabel metal1 228 239 231 243 4 clk
rlabel metal1 360 232 363 236 1 Vdd!
rlabel metal1 361 175 364 179 1 GND!
rlabel metal1 362 168 365 172 2 ~clk
rlabel metal1 360 239 363 243 4 clk
rlabel polysilicon 217 152 217 152 1 0
rlabel polysilicon 241 152 241 152 1 1
rlabel polysilicon 237 141 237 141 1 2
rlabel metal1 96 92 99 96 1 Vdd!
rlabel metal1 97 35 100 39 1 GND!
rlabel metal1 98 28 101 32 2 ~clk
rlabel metal1 96 99 99 103 4 clk
rlabel metal1 228 92 231 96 1 Vdd!
rlabel metal1 229 35 232 39 1 GND!
rlabel metal1 230 28 233 32 2 ~clk
rlabel metal1 228 99 231 103 4 clk
rlabel metal1 360 92 363 96 1 Vdd!
rlabel metal1 361 35 364 39 1 GND!
rlabel metal1 362 28 365 32 2 ~clk
rlabel metal1 360 99 363 103 4 clk
rlabel metal1 360 13 363 17 4 clk
rlabel metal1 362 -58 365 -54 2 ~clk
rlabel metal1 361 -51 364 -47 1 GND!
rlabel metal1 360 6 363 10 1 Vdd!
rlabel metal1 228 13 231 17 4 clk
rlabel metal1 230 -58 233 -54 2 ~clk
rlabel metal1 229 -51 232 -47 1 GND!
rlabel metal1 228 6 231 10 1 Vdd!
rlabel metal1 96 13 99 17 4 clk
rlabel metal1 98 -58 101 -54 2 ~clk
rlabel metal1 97 -51 100 -47 1 GND!
rlabel metal1 96 6 99 10 1 Vdd!
rlabel metal1 360 -127 363 -123 4 clk
rlabel metal1 362 -198 365 -194 2 ~clk
rlabel metal1 361 -191 364 -187 1 GND!
rlabel metal1 360 -134 363 -130 1 Vdd!
rlabel metal1 228 -127 231 -123 4 clk
rlabel metal1 230 -198 233 -194 2 ~clk
rlabel metal1 229 -191 232 -187 1 GND!
rlabel metal1 228 -134 231 -130 1 Vdd!
rlabel metal1 96 -127 99 -123 4 clk
rlabel metal1 98 -198 101 -194 2 ~clk
rlabel metal1 97 -191 100 -187 1 GND!
rlabel metal1 96 -134 99 -130 1 Vdd!
rlabel polysilicon 334 -73 334 -73 1 6
rlabel polysilicon 358 -73 358 -73 1 7
rlabel polysilicon 354 -91 354 -91 1 8
rlabel polysilicon 217 112 217 112 1 3
rlabel polysilicon 241 112 241 112 1 4
rlabel polysilicon 239 123 239 123 1 5
rlabel polysilicon 334 -114 334 -114 1 9
rlabel polysilicon 358 -115 358 -115 1 10
rlabel polysilicon 353 -103 353 -103 1 11
rlabel metal1 566 683 570 687 3 clk
rlabel metal1 566 690 570 694 3 Vdd!
rlabel metal1 566 631 570 635 3 ~clk
rlabel metal1 566 617 570 621 3 ~clk
rlabel metal1 566 624 570 628 3 GND!
rlabel metal1 566 551 570 555 3 clk
rlabel metal1 566 558 570 562 3 Vdd!
rlabel metal1 566 499 570 503 3 ~clk
rlabel metal1 566 433 570 437 3 clk
rlabel metal1 566 485 570 489 3 ~clk
rlabel metal1 566 492 570 496 3 GND!
rlabel metal1 566 228 570 232 3 GND!
rlabel metal1 566 221 570 225 3 ~clk
rlabel metal1 566 162 570 166 3 Vdd!
rlabel metal1 566 235 570 239 3 ~clk
rlabel metal1 566 294 570 298 3 Vdd!
rlabel metal1 566 287 570 291 3 clk
rlabel metal1 566 360 570 364 3 GND!
rlabel metal1 566 353 570 357 3 ~clk
rlabel metal1 566 301 570 305 3 clk
rlabel metal1 566 367 570 371 3 ~clk
rlabel metal1 566 426 570 430 3 Vdd!
rlabel metal1 566 419 570 423 3 clk
rlabel polysilicon 830 201 832 204 5 reset
rlabel polysilicon 812 192 814 195 5 D
rlabel metal1 768 162 772 166 1 Vdd!
rlabel metal1 769 228 772 232 1 GND!
rlabel metal1 939 294 943 298 1 Vdd!
rlabel metal1 849 294 853 298 1 Vdd!
rlabel metal1 768 294 772 298 1 Vdd!
rlabel metal1 940 360 943 364 1 GND!
rlabel metal1 850 360 853 364 1 GND!
rlabel metal1 769 360 772 364 1 GND!
rlabel metal1 939 426 943 430 1 Vdd!
rlabel metal1 768 426 772 430 1 Vdd!
rlabel metal1 849 426 853 430 1 Vdd!
rlabel metal1 769 492 772 496 1 GND!
rlabel metal1 874 492 877 496 1 GND!
rlabel metal1 768 558 772 562 1 Vdd!
rlabel metal1 849 558 853 562 1 Vdd!
rlabel metal1 918 529 921 532 7 Y
rlabel metal1 768 690 772 694 1 Vdd!
rlabel metal1 849 690 853 694 1 Vdd!
rlabel metal1 769 624 772 628 1 GND!
rlabel metal1 850 624 853 628 1 GND!
rlabel metal2 913 685 916 690 1 select_out
rlabel metal1 568 767 571 771 1 Vdd!
rlabel metal1 569 710 572 714 1 GND!
rlabel metal1 570 703 573 707 2 ~clk
rlabel metal1 568 774 571 778 4 clk
rlabel metal1 701 710 704 714 1 GND!
rlabel metal1 702 703 705 707 2 ~clk
rlabel metal1 700 774 703 778 4 clk
rlabel metal1 832 767 835 771 1 Vdd!
rlabel metal1 833 710 836 714 1 GND!
rlabel metal1 834 703 837 707 2 ~clk
rlabel metal1 832 774 835 778 4 clk
rlabel metal1 964 774 967 778 4 clk
rlabel metal1 966 703 969 707 2 ~clk
rlabel metal1 965 710 968 714 1 GND!
rlabel metal1 964 767 967 771 1 Vdd!
rlabel m3contact 565 740 568 743 3 ctrl_reg
rlabel metal2 742 695 745 700 1 select0
rlabel metal2 825 694 828 701 1 select1
rlabel metal2 885 694 888 700 1 select2
rlabel metal1 829 162 833 166 1 Vdd!
rlabel metal1 818 228 822 232 1 GND!
rlabel metal1 819 221 823 225 1 ~clk
rlabel metal1 822 169 825 173 1 clk
rlabel metal1 700 767 703 771 1 Vdd!
rlabel metal2 544 782 544 782 5 p_clk_b
rlabel metal2 556 782 556 782 5 p_clk
rlabel metal2 532 781 532 781 5 f_clk
rlabel metal2 520 782 520 782 4 f_clk_b
rlabel metal1 228 734 231 738 1 Vdd!
rlabel metal1 229 677 232 681 1 GND!
rlabel metal1 230 670 233 674 2 ~clk
rlabel metal1 228 741 231 745 4 clk
rlabel polysilicon 358 661 358 661 1 CB2
rlabel metal1 344 632 347 636 1 Vdd!
rlabel metal1 343 575 346 579 1 GND!
rlabel metal1 342 568 345 572 8 ~clk
rlabel metal1 344 639 347 643 6 clk
rlabel metal1 349 607 349 607 1 D
rlabel polysilicon 241 653 241 653 1 CB1
rlabel metal1 867 129 870 133 4 clk
rlabel metal1 869 58 872 62 2 ~clk
rlabel metal1 868 65 871 69 1 GND!
rlabel metal1 867 122 870 126 1 Vdd!
rlabel metal1 867 36 870 40 1 Vdd!
rlabel metal1 868 -21 871 -17 1 GND!
rlabel metal1 869 -28 872 -24 2 ~clk
rlabel metal1 867 43 870 47 4 clk
rlabel polysilicon 1019 6 1019 6 1 CB4
rlabel polysilicon 1007 150 1007 150 1 CB3
rlabel metal1 998 399 998 399 1 out
rlabel metal2 495 783 495 783 1 Vdd!
rlabel metal2 507 783 507 783 1 GND!
rlabel metal1 1029 232 1032 236 1 Vdd!
rlabel metal1 1030 175 1033 179 1 GND!
rlabel metal1 1031 168 1034 172 2 ~clk
rlabel metal1 1029 239 1032 243 4 clk
rlabel metal1 1161 232 1164 236 1 Vdd!
rlabel metal1 1162 175 1165 179 1 GND!
rlabel metal1 1163 168 1166 172 2 ~clk
rlabel metal1 1161 239 1164 243 4 clk
rlabel metal1 1293 232 1296 236 1 Vdd!
rlabel metal1 1294 175 1297 179 1 GND!
rlabel metal1 1295 168 1298 172 2 ~clk
rlabel metal1 1293 239 1296 243 4 clk
rlabel polysilicon 1150 152 1150 152 1 0
rlabel polysilicon 1174 152 1174 152 1 1
rlabel polysilicon 1170 141 1170 141 1 2
rlabel metal1 1029 92 1032 96 1 Vdd!
rlabel metal1 1030 35 1033 39 1 GND!
rlabel metal1 1031 28 1034 32 2 ~clk
rlabel metal1 1029 99 1032 103 4 clk
rlabel metal1 1161 92 1164 96 1 Vdd!
rlabel metal1 1162 35 1165 39 1 GND!
rlabel metal1 1163 28 1166 32 2 ~clk
rlabel metal1 1161 99 1164 103 4 clk
rlabel metal1 1293 92 1296 96 1 Vdd!
rlabel metal1 1294 35 1297 39 1 GND!
rlabel metal1 1295 28 1298 32 2 ~clk
rlabel metal1 1293 99 1296 103 4 clk
rlabel metal1 1293 13 1296 17 4 clk
rlabel metal1 1295 -58 1298 -54 2 ~clk
rlabel metal1 1294 -51 1297 -47 1 GND!
rlabel metal1 1293 6 1296 10 1 Vdd!
rlabel metal1 1161 13 1164 17 4 clk
rlabel metal1 1163 -58 1166 -54 2 ~clk
rlabel metal1 1162 -51 1165 -47 1 GND!
rlabel metal1 1161 6 1164 10 1 Vdd!
rlabel metal1 1029 13 1032 17 4 clk
rlabel metal1 1031 -58 1034 -54 2 ~clk
rlabel metal1 1030 -51 1033 -47 1 GND!
rlabel metal1 1029 6 1032 10 1 Vdd!
rlabel metal1 1293 -127 1296 -123 4 clk
rlabel metal1 1295 -198 1298 -194 2 ~clk
rlabel metal1 1294 -191 1297 -187 1 GND!
rlabel metal1 1293 -134 1296 -130 1 Vdd!
rlabel metal1 1161 -127 1164 -123 4 clk
rlabel metal1 1163 -198 1166 -194 2 ~clk
rlabel metal1 1162 -191 1165 -187 1 GND!
rlabel metal1 1161 -134 1164 -130 1 Vdd!
rlabel metal1 1029 -127 1032 -123 4 clk
rlabel metal1 1031 -198 1034 -194 2 ~clk
rlabel metal1 1030 -191 1033 -187 1 GND!
rlabel metal1 1029 -134 1032 -130 1 Vdd!
rlabel polysilicon 1267 -73 1267 -73 1 6
rlabel polysilicon 1291 -73 1291 -73 1 7
rlabel polysilicon 1287 -91 1287 -91 1 8
rlabel polysilicon 1150 112 1150 112 1 3
rlabel polysilicon 1174 112 1174 112 1 4
rlabel polysilicon 1172 123 1172 123 1 5
rlabel polysilicon 1267 -114 1267 -114 1 9
rlabel polysilicon 1291 -115 1291 -115 1 10
rlabel polysilicon 1286 -103 1286 -103 1 11
rlabel metal1 1499 683 1503 687 3 clk
rlabel metal1 1499 690 1503 694 3 Vdd!
rlabel metal1 1499 631 1503 635 3 ~clk
rlabel metal1 1499 617 1503 621 3 ~clk
rlabel metal1 1499 624 1503 628 3 GND!
rlabel metal1 1499 551 1503 555 3 clk
rlabel metal1 1499 558 1503 562 3 Vdd!
rlabel metal1 1499 499 1503 503 3 ~clk
rlabel metal1 1499 433 1503 437 3 clk
rlabel metal1 1499 485 1503 489 3 ~clk
rlabel metal1 1499 492 1503 496 3 GND!
rlabel metal1 1499 228 1503 232 3 GND!
rlabel metal1 1499 221 1503 225 3 ~clk
rlabel metal1 1499 162 1503 166 3 Vdd!
rlabel metal1 1499 235 1503 239 3 ~clk
rlabel metal1 1499 294 1503 298 3 Vdd!
rlabel metal1 1499 287 1503 291 3 clk
rlabel metal1 1499 360 1503 364 3 GND!
rlabel metal1 1499 353 1503 357 3 ~clk
rlabel metal1 1499 301 1503 305 3 clk
rlabel metal1 1499 367 1503 371 3 ~clk
rlabel metal1 1499 426 1503 430 3 Vdd!
rlabel metal1 1499 419 1503 423 3 clk
rlabel polysilicon 1763 201 1765 204 5 reset
rlabel polysilicon 1745 192 1747 195 5 D
rlabel metal1 1701 162 1705 166 1 Vdd!
rlabel metal1 1702 228 1705 232 1 GND!
rlabel metal1 1872 294 1876 298 1 Vdd!
rlabel metal1 1782 294 1786 298 1 Vdd!
rlabel metal1 1701 294 1705 298 1 Vdd!
rlabel metal1 1873 360 1876 364 1 GND!
rlabel metal1 1783 360 1786 364 1 GND!
rlabel metal1 1702 360 1705 364 1 GND!
rlabel metal1 1872 426 1876 430 1 Vdd!
rlabel metal1 1701 426 1705 430 1 Vdd!
rlabel metal1 1782 426 1786 430 1 Vdd!
rlabel metal1 1702 492 1705 496 1 GND!
rlabel metal1 1807 492 1810 496 1 GND!
rlabel metal1 1701 558 1705 562 1 Vdd!
rlabel metal1 1782 558 1786 562 1 Vdd!
rlabel metal1 1851 529 1854 532 7 Y
rlabel metal1 1701 690 1705 694 1 Vdd!
rlabel metal1 1782 690 1786 694 1 Vdd!
rlabel metal1 1702 624 1705 628 1 GND!
rlabel metal1 1783 624 1786 628 1 GND!
rlabel metal2 1846 685 1849 690 1 select_out
rlabel metal1 1501 767 1504 771 1 Vdd!
rlabel metal1 1502 710 1505 714 1 GND!
rlabel metal1 1503 703 1506 707 2 ~clk
rlabel metal1 1501 774 1504 778 4 clk
rlabel metal1 1634 710 1637 714 1 GND!
rlabel metal1 1635 703 1638 707 2 ~clk
rlabel metal1 1633 774 1636 778 4 clk
rlabel metal1 1765 767 1768 771 1 Vdd!
rlabel metal1 1766 710 1769 714 1 GND!
rlabel metal1 1767 703 1770 707 2 ~clk
rlabel metal1 1765 774 1768 778 4 clk
rlabel metal1 1897 774 1900 778 4 clk
rlabel metal1 1899 703 1902 707 2 ~clk
rlabel metal1 1898 710 1901 714 1 GND!
rlabel metal1 1897 767 1900 771 1 Vdd!
rlabel m3contact 1498 740 1501 743 3 ctrl_reg
rlabel metal2 1675 695 1678 700 1 select0
rlabel metal2 1758 694 1761 701 1 select1
rlabel metal2 1818 694 1821 700 1 select2
rlabel metal1 1762 162 1766 166 1 Vdd!
rlabel metal1 1751 228 1755 232 1 GND!
rlabel metal1 1752 221 1756 225 1 ~clk
rlabel metal1 1755 169 1758 173 1 clk
rlabel metal1 1633 767 1636 771 1 Vdd!
rlabel metal2 1477 782 1477 782 5 p_clk_b
rlabel metal2 1489 782 1489 782 5 p_clk
rlabel metal2 1465 781 1465 781 5 f_clk
rlabel metal2 1453 782 1453 782 4 f_clk_b
rlabel metal1 1161 734 1164 738 1 Vdd!
rlabel metal1 1162 677 1165 681 1 GND!
rlabel metal1 1163 670 1166 674 2 ~clk
rlabel metal1 1161 741 1164 745 4 clk
rlabel polysilicon 1291 661 1291 661 1 CB2
rlabel metal1 1277 632 1280 636 1 Vdd!
rlabel metal1 1276 575 1279 579 1 GND!
rlabel metal1 1275 568 1278 572 8 ~clk
rlabel metal1 1277 639 1280 643 6 clk
rlabel metal1 1282 607 1282 607 1 D
rlabel polysilicon 1174 653 1174 653 1 CB1
rlabel metal1 1800 129 1803 133 4 clk
rlabel metal1 1802 58 1805 62 2 ~clk
rlabel metal1 1801 65 1804 69 1 GND!
rlabel metal1 1800 122 1803 126 1 Vdd!
rlabel metal1 1800 36 1803 40 1 Vdd!
rlabel metal1 1801 -21 1804 -17 1 GND!
rlabel metal1 1802 -28 1805 -24 2 ~clk
rlabel metal1 1800 43 1803 47 4 clk
rlabel polysilicon 1952 6 1952 6 1 CB4
rlabel polysilicon 1940 150 1940 150 1 CB3
rlabel metal1 1931 399 1931 399 1 out
rlabel metal2 1428 783 1428 783 1 Vdd!
rlabel metal2 1440 783 1440 783 1 GND!
rlabel metal2 1440 1763 1440 1763 1 GND!
rlabel metal2 1428 1763 1428 1763 1 Vdd!
rlabel metal1 1931 1379 1931 1379 1 out
rlabel polysilicon 1940 1130 1940 1130 1 CB3
rlabel polysilicon 1952 986 1952 986 1 CB4
rlabel metal1 1800 1023 1803 1027 4 clk
rlabel metal1 1802 952 1805 956 2 ~clk
rlabel metal1 1801 959 1804 963 1 GND!
rlabel metal1 1800 1016 1803 1020 1 Vdd!
rlabel metal1 1800 1102 1803 1106 1 Vdd!
rlabel metal1 1801 1045 1804 1049 1 GND!
rlabel metal1 1802 1038 1805 1042 2 ~clk
rlabel metal1 1800 1109 1803 1113 4 clk
rlabel polysilicon 1174 1633 1174 1633 1 CB1
rlabel metal1 1282 1587 1282 1587 1 D
rlabel metal1 1277 1619 1280 1623 6 clk
rlabel metal1 1275 1548 1278 1552 8 ~clk
rlabel metal1 1276 1555 1279 1559 1 GND!
rlabel metal1 1277 1612 1280 1616 1 Vdd!
rlabel polysilicon 1291 1641 1291 1641 1 CB2
rlabel metal1 1161 1721 1164 1725 4 clk
rlabel metal1 1163 1650 1166 1654 2 ~clk
rlabel metal1 1162 1657 1165 1661 1 GND!
rlabel metal1 1161 1714 1164 1718 1 Vdd!
rlabel metal2 1453 1762 1453 1762 4 f_clk_b
rlabel metal2 1465 1761 1465 1761 5 f_clk
rlabel metal2 1489 1762 1489 1762 5 p_clk
rlabel metal2 1477 1762 1477 1762 5 p_clk_b
rlabel metal1 1633 1747 1636 1751 1 Vdd!
rlabel metal1 1755 1149 1758 1153 1 clk
rlabel metal1 1752 1201 1756 1205 1 ~clk
rlabel metal1 1751 1208 1755 1212 1 GND!
rlabel metal1 1762 1142 1766 1146 1 Vdd!
rlabel metal2 1818 1674 1821 1680 1 select2
rlabel metal2 1758 1674 1761 1681 1 select1
rlabel metal2 1675 1675 1678 1680 1 select0
rlabel m3contact 1498 1720 1501 1723 3 ctrl_reg
rlabel metal1 1897 1747 1900 1751 1 Vdd!
rlabel metal1 1898 1690 1901 1694 1 GND!
rlabel metal1 1899 1683 1902 1687 2 ~clk
rlabel metal1 1897 1754 1900 1758 4 clk
rlabel metal1 1765 1754 1768 1758 4 clk
rlabel metal1 1767 1683 1770 1687 2 ~clk
rlabel metal1 1766 1690 1769 1694 1 GND!
rlabel metal1 1765 1747 1768 1751 1 Vdd!
rlabel metal1 1633 1754 1636 1758 4 clk
rlabel metal1 1635 1683 1638 1687 2 ~clk
rlabel metal1 1634 1690 1637 1694 1 GND!
rlabel metal1 1501 1754 1504 1758 4 clk
rlabel metal1 1503 1683 1506 1687 2 ~clk
rlabel metal1 1502 1690 1505 1694 1 GND!
rlabel metal1 1501 1747 1504 1751 1 Vdd!
rlabel metal2 1846 1665 1849 1670 1 select_out
rlabel metal1 1783 1604 1786 1608 1 GND!
rlabel metal1 1702 1604 1705 1608 1 GND!
rlabel metal1 1782 1670 1786 1674 1 Vdd!
rlabel metal1 1701 1670 1705 1674 1 Vdd!
rlabel metal1 1851 1509 1854 1512 7 Y
rlabel metal1 1782 1538 1786 1542 1 Vdd!
rlabel metal1 1701 1538 1705 1542 1 Vdd!
rlabel metal1 1807 1472 1810 1476 1 GND!
rlabel metal1 1702 1472 1705 1476 1 GND!
rlabel metal1 1782 1406 1786 1410 1 Vdd!
rlabel metal1 1701 1406 1705 1410 1 Vdd!
rlabel metal1 1872 1406 1876 1410 1 Vdd!
rlabel metal1 1702 1340 1705 1344 1 GND!
rlabel metal1 1783 1340 1786 1344 1 GND!
rlabel metal1 1873 1340 1876 1344 1 GND!
rlabel metal1 1701 1274 1705 1278 1 Vdd!
rlabel metal1 1782 1274 1786 1278 1 Vdd!
rlabel metal1 1872 1274 1876 1278 1 Vdd!
rlabel metal1 1702 1208 1705 1212 1 GND!
rlabel metal1 1701 1142 1705 1146 1 Vdd!
rlabel polysilicon 1745 1172 1747 1175 5 D
rlabel polysilicon 1763 1181 1765 1184 5 reset
rlabel metal1 1499 1399 1503 1403 3 clk
rlabel metal1 1499 1406 1503 1410 3 Vdd!
rlabel metal1 1499 1347 1503 1351 3 ~clk
rlabel metal1 1499 1281 1503 1285 3 clk
rlabel metal1 1499 1333 1503 1337 3 ~clk
rlabel metal1 1499 1340 1503 1344 3 GND!
rlabel metal1 1499 1267 1503 1271 3 clk
rlabel metal1 1499 1274 1503 1278 3 Vdd!
rlabel metal1 1499 1215 1503 1219 3 ~clk
rlabel metal1 1499 1142 1503 1146 3 Vdd!
rlabel metal1 1499 1201 1503 1205 3 ~clk
rlabel metal1 1499 1208 1503 1212 3 GND!
rlabel metal1 1499 1472 1503 1476 3 GND!
rlabel metal1 1499 1465 1503 1469 3 ~clk
rlabel metal1 1499 1413 1503 1417 3 clk
rlabel metal1 1499 1479 1503 1483 3 ~clk
rlabel metal1 1499 1538 1503 1542 3 Vdd!
rlabel metal1 1499 1531 1503 1535 3 clk
rlabel metal1 1499 1604 1503 1608 3 GND!
rlabel metal1 1499 1597 1503 1601 3 ~clk
rlabel metal1 1499 1611 1503 1615 3 ~clk
rlabel metal1 1499 1670 1503 1674 3 Vdd!
rlabel metal1 1499 1663 1503 1667 3 clk
rlabel polysilicon 1286 877 1286 877 1 11
rlabel polysilicon 1291 865 1291 865 1 10
rlabel polysilicon 1267 866 1267 866 1 9
rlabel polysilicon 1172 1103 1172 1103 1 5
rlabel polysilicon 1174 1092 1174 1092 1 4
rlabel polysilicon 1150 1092 1150 1092 1 3
rlabel polysilicon 1287 889 1287 889 1 8
rlabel polysilicon 1291 907 1291 907 1 7
rlabel polysilicon 1267 907 1267 907 1 6
rlabel metal1 1029 846 1032 850 1 Vdd!
rlabel metal1 1030 789 1033 793 1 GND!
rlabel metal1 1031 782 1034 786 2 ~clk
rlabel metal1 1029 853 1032 857 4 clk
rlabel metal1 1161 846 1164 850 1 Vdd!
rlabel metal1 1162 789 1165 793 1 GND!
rlabel metal1 1163 782 1166 786 2 ~clk
rlabel metal1 1161 853 1164 857 4 clk
rlabel metal1 1293 846 1296 850 1 Vdd!
rlabel metal1 1294 789 1297 793 1 GND!
rlabel metal1 1295 782 1298 786 2 ~clk
rlabel metal1 1293 853 1296 857 4 clk
rlabel metal1 1029 986 1032 990 1 Vdd!
rlabel metal1 1030 929 1033 933 1 GND!
rlabel metal1 1031 922 1034 926 2 ~clk
rlabel metal1 1029 993 1032 997 4 clk
rlabel metal1 1161 986 1164 990 1 Vdd!
rlabel metal1 1162 929 1165 933 1 GND!
rlabel metal1 1163 922 1166 926 2 ~clk
rlabel metal1 1161 993 1164 997 4 clk
rlabel metal1 1293 986 1296 990 1 Vdd!
rlabel metal1 1294 929 1297 933 1 GND!
rlabel metal1 1295 922 1298 926 2 ~clk
rlabel metal1 1293 993 1296 997 4 clk
rlabel metal1 1293 1079 1296 1083 4 clk
rlabel metal1 1295 1008 1298 1012 2 ~clk
rlabel metal1 1294 1015 1297 1019 1 GND!
rlabel metal1 1293 1072 1296 1076 1 Vdd!
rlabel metal1 1161 1079 1164 1083 4 clk
rlabel metal1 1163 1008 1166 1012 2 ~clk
rlabel metal1 1162 1015 1165 1019 1 GND!
rlabel metal1 1161 1072 1164 1076 1 Vdd!
rlabel metal1 1029 1079 1032 1083 4 clk
rlabel metal1 1031 1008 1034 1012 2 ~clk
rlabel metal1 1030 1015 1033 1019 1 GND!
rlabel metal1 1029 1072 1032 1076 1 Vdd!
rlabel polysilicon 1170 1121 1170 1121 1 2
rlabel polysilicon 1174 1132 1174 1132 1 1
rlabel polysilicon 1150 1132 1150 1132 1 0
rlabel metal1 1293 1219 1296 1223 4 clk
rlabel metal1 1295 1148 1298 1152 2 ~clk
rlabel metal1 1294 1155 1297 1159 1 GND!
rlabel metal1 1293 1212 1296 1216 1 Vdd!
rlabel metal1 1161 1219 1164 1223 4 clk
rlabel metal1 1163 1148 1166 1152 2 ~clk
rlabel metal1 1162 1155 1165 1159 1 GND!
rlabel metal1 1161 1212 1164 1216 1 Vdd!
rlabel metal1 1029 1219 1032 1223 4 clk
rlabel metal1 1031 1148 1034 1152 2 ~clk
rlabel metal1 1030 1155 1033 1159 1 GND!
rlabel metal1 1029 1212 1032 1216 1 Vdd!
rlabel metal2 507 1763 507 1763 1 GND!
rlabel metal2 495 1763 495 1763 1 Vdd!
rlabel metal1 998 1379 998 1379 1 out
rlabel polysilicon 1007 1130 1007 1130 1 CB3
rlabel polysilicon 1019 986 1019 986 1 CB4
rlabel metal1 867 1023 870 1027 4 clk
rlabel metal1 869 952 872 956 2 ~clk
rlabel metal1 868 959 871 963 1 GND!
rlabel metal1 867 1016 870 1020 1 Vdd!
rlabel metal1 867 1102 870 1106 1 Vdd!
rlabel metal1 868 1045 871 1049 1 GND!
rlabel metal1 869 1038 872 1042 2 ~clk
rlabel metal1 867 1109 870 1113 4 clk
rlabel polysilicon 241 1633 241 1633 1 CB1
rlabel metal1 349 1587 349 1587 1 D
rlabel metal1 344 1619 347 1623 6 clk
rlabel metal1 342 1548 345 1552 8 ~clk
rlabel metal1 343 1555 346 1559 1 GND!
rlabel metal1 344 1612 347 1616 1 Vdd!
rlabel polysilicon 358 1641 358 1641 1 CB2
rlabel metal1 228 1721 231 1725 4 clk
rlabel metal1 230 1650 233 1654 2 ~clk
rlabel metal1 229 1657 232 1661 1 GND!
rlabel metal1 228 1714 231 1718 1 Vdd!
rlabel metal2 520 1762 520 1762 4 f_clk_b
rlabel metal2 532 1761 532 1761 5 f_clk
rlabel metal2 556 1762 556 1762 5 p_clk
rlabel metal2 544 1762 544 1762 5 p_clk_b
rlabel metal1 700 1747 703 1751 1 Vdd!
rlabel metal1 822 1149 825 1153 1 clk
rlabel metal1 819 1201 823 1205 1 ~clk
rlabel metal1 818 1208 822 1212 1 GND!
rlabel metal1 829 1142 833 1146 1 Vdd!
rlabel metal2 885 1674 888 1680 1 select2
rlabel metal2 825 1674 828 1681 1 select1
rlabel metal2 742 1675 745 1680 1 select0
rlabel m3contact 565 1720 568 1723 3 ctrl_reg
rlabel metal1 964 1747 967 1751 1 Vdd!
rlabel metal1 965 1690 968 1694 1 GND!
rlabel metal1 966 1683 969 1687 2 ~clk
rlabel metal1 964 1754 967 1758 4 clk
rlabel metal1 832 1754 835 1758 4 clk
rlabel metal1 834 1683 837 1687 2 ~clk
rlabel metal1 833 1690 836 1694 1 GND!
rlabel metal1 832 1747 835 1751 1 Vdd!
rlabel metal1 700 1754 703 1758 4 clk
rlabel metal1 702 1683 705 1687 2 ~clk
rlabel metal1 701 1690 704 1694 1 GND!
rlabel metal1 568 1754 571 1758 4 clk
rlabel metal1 570 1683 573 1687 2 ~clk
rlabel metal1 569 1690 572 1694 1 GND!
rlabel metal1 568 1747 571 1751 1 Vdd!
rlabel metal2 913 1665 916 1670 1 select_out
rlabel metal1 850 1604 853 1608 1 GND!
rlabel metal1 769 1604 772 1608 1 GND!
rlabel metal1 849 1670 853 1674 1 Vdd!
rlabel metal1 768 1670 772 1674 1 Vdd!
rlabel metal1 918 1509 921 1512 7 Y
rlabel metal1 849 1538 853 1542 1 Vdd!
rlabel metal1 768 1538 772 1542 1 Vdd!
rlabel metal1 874 1472 877 1476 1 GND!
rlabel metal1 769 1472 772 1476 1 GND!
rlabel metal1 849 1406 853 1410 1 Vdd!
rlabel metal1 768 1406 772 1410 1 Vdd!
rlabel metal1 939 1406 943 1410 1 Vdd!
rlabel metal1 769 1340 772 1344 1 GND!
rlabel metal1 850 1340 853 1344 1 GND!
rlabel metal1 940 1340 943 1344 1 GND!
rlabel metal1 768 1274 772 1278 1 Vdd!
rlabel metal1 849 1274 853 1278 1 Vdd!
rlabel metal1 939 1274 943 1278 1 Vdd!
rlabel metal1 769 1208 772 1212 1 GND!
rlabel metal1 768 1142 772 1146 1 Vdd!
rlabel polysilicon 812 1172 814 1175 5 D
rlabel polysilicon 830 1181 832 1184 5 reset
rlabel metal1 566 1399 570 1403 3 clk
rlabel metal1 566 1406 570 1410 3 Vdd!
rlabel metal1 566 1347 570 1351 3 ~clk
rlabel metal1 566 1281 570 1285 3 clk
rlabel metal1 566 1333 570 1337 3 ~clk
rlabel metal1 566 1340 570 1344 3 GND!
rlabel metal1 566 1267 570 1271 3 clk
rlabel metal1 566 1274 570 1278 3 Vdd!
rlabel metal1 566 1215 570 1219 3 ~clk
rlabel metal1 566 1142 570 1146 3 Vdd!
rlabel metal1 566 1201 570 1205 3 ~clk
rlabel metal1 566 1208 570 1212 3 GND!
rlabel metal1 566 1472 570 1476 3 GND!
rlabel metal1 566 1465 570 1469 3 ~clk
rlabel metal1 566 1413 570 1417 3 clk
rlabel metal1 566 1479 570 1483 3 ~clk
rlabel metal1 566 1538 570 1542 3 Vdd!
rlabel metal1 566 1531 570 1535 3 clk
rlabel metal1 566 1604 570 1608 3 GND!
rlabel metal1 566 1597 570 1601 3 ~clk
rlabel metal1 566 1611 570 1615 3 ~clk
rlabel metal1 566 1670 570 1674 3 Vdd!
rlabel metal1 566 1663 570 1667 3 clk
rlabel polysilicon 353 877 353 877 1 11
rlabel polysilicon 358 865 358 865 1 10
rlabel polysilicon 334 866 334 866 1 9
rlabel polysilicon 239 1103 239 1103 1 5
rlabel polysilicon 241 1092 241 1092 1 4
rlabel polysilicon 217 1092 217 1092 1 3
rlabel polysilicon 354 889 354 889 1 8
rlabel polysilicon 358 907 358 907 1 7
rlabel polysilicon 334 907 334 907 1 6
rlabel metal1 96 846 99 850 1 Vdd!
rlabel metal1 97 789 100 793 1 GND!
rlabel metal1 98 782 101 786 2 ~clk
rlabel metal1 96 853 99 857 4 clk
rlabel metal1 228 846 231 850 1 Vdd!
rlabel metal1 229 789 232 793 1 GND!
rlabel metal1 230 782 233 786 2 ~clk
rlabel metal1 228 853 231 857 4 clk
rlabel metal1 360 846 363 850 1 Vdd!
rlabel metal1 361 789 364 793 1 GND!
rlabel metal1 362 782 365 786 2 ~clk
rlabel metal1 360 853 363 857 4 clk
rlabel metal1 96 986 99 990 1 Vdd!
rlabel metal1 97 929 100 933 1 GND!
rlabel metal1 98 922 101 926 2 ~clk
rlabel metal1 96 993 99 997 4 clk
rlabel metal1 228 986 231 990 1 Vdd!
rlabel metal1 229 929 232 933 1 GND!
rlabel metal1 230 922 233 926 2 ~clk
rlabel metal1 228 993 231 997 4 clk
rlabel metal1 360 986 363 990 1 Vdd!
rlabel metal1 361 929 364 933 1 GND!
rlabel metal1 362 922 365 926 2 ~clk
rlabel metal1 360 993 363 997 4 clk
rlabel metal1 360 1079 363 1083 4 clk
rlabel metal1 362 1008 365 1012 2 ~clk
rlabel metal1 361 1015 364 1019 1 GND!
rlabel metal1 360 1072 363 1076 1 Vdd!
rlabel metal1 228 1079 231 1083 4 clk
rlabel metal1 230 1008 233 1012 2 ~clk
rlabel metal1 229 1015 232 1019 1 GND!
rlabel metal1 228 1072 231 1076 1 Vdd!
rlabel metal1 96 1079 99 1083 4 clk
rlabel metal1 98 1008 101 1012 2 ~clk
rlabel metal1 97 1015 100 1019 1 GND!
rlabel metal1 96 1072 99 1076 1 Vdd!
rlabel polysilicon 237 1121 237 1121 1 2
rlabel polysilicon 241 1132 241 1132 1 1
rlabel polysilicon 217 1132 217 1132 1 0
rlabel metal1 360 1219 363 1223 4 clk
rlabel metal1 362 1148 365 1152 2 ~clk
rlabel metal1 361 1155 364 1159 1 GND!
rlabel metal1 360 1212 363 1216 1 Vdd!
rlabel metal1 228 1219 231 1223 4 clk
rlabel metal1 230 1148 233 1152 2 ~clk
rlabel metal1 229 1155 232 1159 1 GND!
rlabel metal1 228 1212 231 1216 1 Vdd!
rlabel metal1 96 1219 99 1223 4 clk
rlabel metal1 98 1148 101 1152 2 ~clk
rlabel metal1 97 1155 100 1159 1 GND!
rlabel metal1 96 1212 99 1216 1 Vdd!
<< end >>
