magic
tech scmos
timestamp 1607766592
<< ntransistor >>
rect -7 462 -5 466
rect 19 458 21 462
rect 24 458 26 462
rect 74 462 76 466
rect 100 458 102 462
rect 105 458 107 462
rect 47 454 49 458
rect 128 454 130 458
rect 19 428 21 432
rect 24 428 26 432
rect 100 428 102 432
rect 105 428 107 432
rect 19 358 21 362
rect 24 358 26 362
rect 98 362 100 366
rect 124 358 126 362
rect 129 358 131 362
rect 47 354 49 358
rect 152 354 154 358
rect 19 328 21 332
rect 24 328 26 332
rect 124 328 126 332
rect 129 328 131 332
rect 19 258 21 262
rect 24 258 26 262
rect 74 262 76 266
rect 100 258 102 262
rect 105 258 107 262
rect 164 262 166 266
rect 190 258 192 262
rect 195 258 197 262
rect 47 254 49 258
rect 128 254 130 258
rect 218 254 220 258
rect 19 228 21 232
rect 24 228 26 232
rect 100 228 102 232
rect 105 228 107 232
rect 190 228 192 232
rect 195 228 197 232
rect 19 158 21 162
rect 24 158 26 162
rect 47 154 49 158
rect 53 119 55 123
rect 71 119 73 123
rect 87 119 89 123
rect 103 119 105 123
rect 126 119 128 123
rect 131 119 133 123
rect 157 119 159 123
rect 178 119 180 123
rect 198 119 200 123
rect 203 119 205 123
rect 221 119 223 123
rect 19 112 21 116
rect 24 112 26 116
<< ptransistor >>
rect -7 480 -5 488
rect 19 474 21 482
rect 24 474 26 482
rect 47 480 49 488
rect 74 480 76 488
rect 100 474 102 482
rect 105 474 107 482
rect 128 480 130 488
rect 19 408 21 416
rect 24 408 26 416
rect 100 408 102 416
rect 105 408 107 416
rect 19 374 21 382
rect 24 374 26 382
rect 47 380 49 388
rect 98 380 100 388
rect 124 374 126 382
rect 129 374 131 382
rect 152 380 154 388
rect 19 308 21 316
rect 24 308 26 316
rect 124 308 126 316
rect 129 308 131 316
rect 19 274 21 282
rect 24 274 26 282
rect 47 280 49 288
rect 74 280 76 288
rect 100 274 102 282
rect 105 274 107 282
rect 128 280 130 288
rect 164 280 166 288
rect 190 274 192 282
rect 195 274 197 282
rect 218 280 220 288
rect 19 208 21 216
rect 24 208 26 216
rect 100 208 102 216
rect 105 208 107 216
rect 190 208 192 216
rect 195 208 197 216
rect 19 174 21 182
rect 24 174 26 182
rect 47 180 49 188
rect 19 92 21 100
rect 24 92 26 100
rect 53 97 55 105
rect 71 97 73 105
rect 87 97 89 105
rect 103 97 105 105
rect 126 97 128 105
rect 131 97 133 105
rect 157 97 159 105
rect 178 97 180 105
rect 198 97 200 105
rect 203 97 205 105
rect 221 97 223 105
<< ndiffusion >>
rect -8 462 -7 466
rect -5 462 -4 466
rect 16 458 19 462
rect 21 458 24 462
rect 26 458 27 462
rect 73 462 74 466
rect 76 462 77 466
rect 97 458 100 462
rect 102 458 105 462
rect 107 458 108 462
rect 46 454 47 458
rect 49 454 50 458
rect 127 454 128 458
rect 130 454 131 458
rect 16 428 19 432
rect 21 428 24 432
rect 26 428 27 432
rect 97 428 100 432
rect 102 428 105 432
rect 107 428 108 432
rect 16 358 19 362
rect 21 358 24 362
rect 26 358 27 362
rect 97 362 98 366
rect 100 362 101 366
rect 121 358 124 362
rect 126 358 129 362
rect 131 358 132 362
rect 46 354 47 358
rect 49 354 50 358
rect 151 354 152 358
rect 154 354 155 358
rect 16 328 19 332
rect 21 328 24 332
rect 26 328 27 332
rect 121 328 124 332
rect 126 328 129 332
rect 131 328 132 332
rect 16 258 19 262
rect 21 258 24 262
rect 26 258 27 262
rect 73 262 74 266
rect 76 262 77 266
rect 97 258 100 262
rect 102 258 105 262
rect 107 258 108 262
rect 163 262 164 266
rect 166 262 167 266
rect 187 258 190 262
rect 192 258 195 262
rect 197 258 198 262
rect 46 254 47 258
rect 49 254 50 258
rect 127 254 128 258
rect 130 254 131 258
rect 217 254 218 258
rect 220 254 221 258
rect 16 228 19 232
rect 21 228 24 232
rect 26 228 27 232
rect 97 228 100 232
rect 102 228 105 232
rect 107 228 108 232
rect 187 228 190 232
rect 192 228 195 232
rect 197 228 198 232
rect 16 158 19 162
rect 21 158 24 162
rect 26 158 27 162
rect 46 154 47 158
rect 49 154 50 158
rect 52 119 53 123
rect 55 119 56 123
rect 60 119 66 123
rect 70 119 71 123
rect 73 119 74 123
rect 86 119 87 123
rect 89 119 90 123
rect 102 119 103 123
rect 105 119 106 123
rect 121 119 126 123
rect 128 119 131 123
rect 133 119 134 123
rect 155 119 157 123
rect 159 119 160 123
rect 177 119 178 123
rect 180 119 181 123
rect 193 119 198 123
rect 200 119 203 123
rect 205 119 206 123
rect 220 119 221 123
rect 223 119 224 123
rect 16 112 19 116
rect 21 112 24 116
rect 26 112 27 116
<< pdiffusion >>
rect -8 480 -7 488
rect -5 480 -4 488
rect 16 474 19 482
rect 21 474 24 482
rect 26 474 27 482
rect 46 480 47 488
rect 49 480 50 488
rect 73 480 74 488
rect 76 480 77 488
rect 97 474 100 482
rect 102 474 105 482
rect 107 474 108 482
rect 127 480 128 488
rect 130 480 131 488
rect 16 408 19 416
rect 21 408 24 416
rect 26 408 27 416
rect 97 408 100 416
rect 102 408 105 416
rect 107 408 108 416
rect 16 374 19 382
rect 21 374 24 382
rect 26 374 27 382
rect 46 380 47 388
rect 49 380 50 388
rect 97 380 98 388
rect 100 380 101 388
rect 121 374 124 382
rect 126 374 129 382
rect 131 374 132 382
rect 151 380 152 388
rect 154 380 155 388
rect 16 308 19 316
rect 21 308 24 316
rect 26 308 27 316
rect 121 308 124 316
rect 126 308 129 316
rect 131 308 132 316
rect 16 274 19 282
rect 21 274 24 282
rect 26 274 27 282
rect 46 280 47 288
rect 49 280 50 288
rect 73 280 74 288
rect 76 280 77 288
rect 97 274 100 282
rect 102 274 105 282
rect 107 274 108 282
rect 127 280 128 288
rect 130 280 131 288
rect 163 280 164 288
rect 166 280 167 288
rect 187 274 190 282
rect 192 274 195 282
rect 197 274 198 282
rect 217 280 218 288
rect 220 280 221 288
rect 16 208 19 216
rect 21 208 24 216
rect 26 208 27 216
rect 97 208 100 216
rect 102 208 105 216
rect 107 208 108 216
rect 187 208 190 216
rect 192 208 195 216
rect 197 208 198 216
rect 16 174 19 182
rect 21 174 24 182
rect 26 174 27 182
rect 46 180 47 188
rect 49 180 50 188
rect 16 92 19 100
rect 21 92 24 100
rect 26 92 27 100
rect 52 97 53 105
rect 55 97 56 105
rect 60 97 66 105
rect 70 97 71 105
rect 73 97 74 105
rect 86 97 87 105
rect 89 97 90 105
rect 102 97 103 105
rect 105 97 106 105
rect 121 97 126 105
rect 128 97 131 105
rect 133 97 134 105
rect 155 97 157 105
rect 159 97 160 105
rect 177 97 178 105
rect 180 97 181 105
rect 193 97 198 105
rect 200 97 203 105
rect 205 97 206 105
rect 220 97 221 105
rect 223 97 224 105
<< ndcontact >>
rect -12 462 -8 466
rect -4 462 0 466
rect 12 458 16 462
rect 27 458 31 462
rect 69 462 73 466
rect 77 462 81 466
rect 93 458 97 462
rect 108 458 112 462
rect 42 454 46 458
rect 50 454 54 458
rect 123 454 127 458
rect 131 454 135 458
rect 12 428 16 432
rect 27 428 31 432
rect 93 428 97 432
rect 108 428 112 432
rect 12 358 16 362
rect 27 358 31 362
rect 93 362 97 366
rect 101 362 105 366
rect 117 358 121 362
rect 132 358 136 362
rect 42 354 46 358
rect 50 354 54 358
rect 147 354 151 358
rect 155 354 159 358
rect 12 328 16 332
rect 27 328 31 332
rect 117 328 121 332
rect 132 328 136 332
rect 12 258 16 262
rect 27 258 31 262
rect 69 262 73 266
rect 77 262 81 266
rect 93 258 97 262
rect 108 258 112 262
rect 159 262 163 266
rect 167 262 171 266
rect 183 258 187 262
rect 198 258 202 262
rect 42 254 46 258
rect 50 254 54 258
rect 123 254 127 258
rect 131 254 135 258
rect 213 254 217 258
rect 221 254 225 258
rect 12 228 16 232
rect 27 228 31 232
rect 93 228 97 232
rect 108 228 112 232
rect 183 228 187 232
rect 198 228 202 232
rect 12 158 16 162
rect 27 158 31 162
rect 42 154 46 158
rect 50 154 54 158
rect 48 119 52 123
rect 56 119 60 123
rect 66 119 70 123
rect 74 119 78 123
rect 82 119 86 123
rect 90 119 94 123
rect 98 119 102 123
rect 106 119 110 123
rect 117 119 121 123
rect 134 119 138 123
rect 151 119 155 123
rect 160 119 164 123
rect 173 119 177 123
rect 181 119 185 123
rect 189 119 193 123
rect 206 119 210 123
rect 216 119 220 123
rect 224 119 228 123
rect 12 112 16 116
rect 27 112 31 116
<< pdcontact >>
rect -12 480 -8 488
rect -4 480 0 488
rect 12 474 16 482
rect 27 474 31 482
rect 42 480 46 488
rect 50 480 54 488
rect 69 480 73 488
rect 77 480 81 488
rect 93 474 97 482
rect 108 474 112 482
rect 123 480 127 488
rect 131 480 135 488
rect 12 408 16 416
rect 27 408 31 416
rect 93 408 97 416
rect 108 408 112 416
rect 12 374 16 382
rect 27 374 31 382
rect 42 380 46 388
rect 50 380 54 388
rect 93 380 97 388
rect 101 380 105 388
rect 117 374 121 382
rect 132 374 136 382
rect 147 380 151 388
rect 155 380 159 388
rect 12 308 16 316
rect 27 308 31 316
rect 117 308 121 316
rect 132 308 136 316
rect 12 274 16 282
rect 27 274 31 282
rect 42 280 46 288
rect 50 280 54 288
rect 69 280 73 288
rect 77 280 81 288
rect 93 274 97 282
rect 108 274 112 282
rect 123 280 127 288
rect 131 280 135 288
rect 159 280 163 288
rect 167 280 171 288
rect 183 274 187 282
rect 198 274 202 282
rect 213 280 217 288
rect 221 280 225 288
rect 12 208 16 216
rect 27 208 31 216
rect 93 208 97 216
rect 108 208 112 216
rect 183 208 187 216
rect 198 208 202 216
rect 12 174 16 182
rect 27 174 31 182
rect 42 180 46 188
rect 50 180 54 188
rect 12 92 16 100
rect 27 92 31 100
rect 48 97 52 105
rect 56 97 60 105
rect 66 97 70 105
rect 74 97 78 105
rect 82 97 86 105
rect 90 97 94 105
rect 98 97 102 105
rect 106 97 110 105
rect 117 97 121 105
rect 134 97 138 105
rect 151 97 155 105
rect 160 97 164 105
rect 173 97 177 105
rect 181 97 185 105
rect 189 97 193 105
rect 206 97 210 105
rect 216 97 220 105
rect 224 97 228 105
<< psubstratepcontact >>
rect -19 442 -15 446
rect 5 442 9 446
rect 59 442 66 446
rect 86 442 90 446
rect 140 442 144 446
rect -19 342 -15 346
rect 5 342 9 346
rect 59 342 63 346
rect 86 342 90 346
rect 110 342 114 346
rect -19 242 -15 246
rect 5 242 9 246
rect 59 242 66 246
rect 86 242 90 246
rect 140 242 144 246
rect 176 242 180 246
rect 230 242 234 246
rect -19 142 -15 146
rect 5 142 9 146
rect 78 135 82 139
rect 107 135 111 139
rect 143 135 147 139
rect 182 135 186 139
rect 59 76 63 80
<< nsubstratencontact >>
rect -19 492 -15 496
rect 5 492 9 496
rect 59 492 63 496
rect 86 492 90 496
rect 140 492 144 496
rect -19 392 -15 396
rect 5 392 9 396
rect 59 392 63 396
rect 86 392 90 396
rect 148 392 152 396
rect -19 292 -15 296
rect 5 292 9 296
rect 59 292 63 296
rect 86 292 90 296
rect 140 292 144 296
rect 148 292 152 296
rect 176 292 180 296
rect 230 292 234 296
rect -19 192 -15 196
rect 5 192 9 196
rect 59 192 63 196
rect 86 192 90 196
rect 176 192 180 196
rect 75 83 79 87
rect 107 83 111 87
rect 143 83 147 87
rect 182 83 186 87
rect 5 76 9 80
<< polysilicon >>
rect -7 488 -5 490
rect 19 482 21 486
rect 47 488 49 490
rect 74 488 76 490
rect 24 482 26 485
rect -7 466 -5 480
rect 100 482 102 486
rect 128 488 130 490
rect 105 482 107 485
rect 19 471 21 474
rect 24 472 26 474
rect 20 467 21 471
rect 19 462 21 467
rect 24 462 26 464
rect -7 460 -5 462
rect 47 458 49 480
rect 74 466 76 480
rect 100 471 102 474
rect 105 472 107 474
rect 101 467 102 471
rect 100 462 102 467
rect 105 462 107 464
rect 74 460 76 462
rect 128 458 130 480
rect 19 456 21 458
rect 24 453 26 458
rect 100 456 102 458
rect 47 452 49 454
rect 105 453 107 458
rect 128 452 130 454
rect 19 432 21 435
rect 24 432 26 435
rect 100 432 102 435
rect 105 432 107 435
rect 19 416 21 428
rect 24 426 26 428
rect 24 416 26 418
rect 100 416 102 428
rect 105 426 107 428
rect 105 416 107 418
rect 19 406 21 408
rect 24 403 26 408
rect 100 406 102 408
rect 105 403 107 408
rect 19 382 21 386
rect 47 388 49 390
rect 98 388 100 390
rect 24 382 26 385
rect 124 382 126 386
rect 152 388 154 390
rect 129 382 131 385
rect 19 371 21 374
rect 24 372 26 374
rect 20 367 21 371
rect 19 362 21 367
rect 24 362 26 364
rect 47 358 49 380
rect 98 366 100 380
rect 124 371 126 374
rect 129 372 131 374
rect 125 367 126 371
rect 124 362 126 367
rect 129 362 131 364
rect 98 360 100 362
rect 152 358 154 380
rect 19 356 21 358
rect 24 353 26 358
rect 124 356 126 358
rect 47 352 49 354
rect 129 353 131 358
rect 152 352 154 354
rect 19 332 21 335
rect 24 332 26 335
rect 124 332 126 335
rect 129 332 131 335
rect 19 316 21 328
rect 24 326 26 328
rect 24 316 26 318
rect 124 316 126 328
rect 129 326 131 328
rect 129 316 131 318
rect 19 306 21 308
rect 24 303 26 308
rect 124 306 126 308
rect 129 303 131 308
rect 19 282 21 286
rect 47 288 49 290
rect 74 288 76 290
rect 24 282 26 285
rect 100 282 102 286
rect 128 288 130 290
rect 164 288 166 290
rect 105 282 107 285
rect 19 271 21 274
rect 24 272 26 274
rect 20 267 21 271
rect 19 262 21 267
rect 24 262 26 264
rect 47 258 49 280
rect 74 266 76 280
rect 190 282 192 286
rect 218 288 220 290
rect 195 282 197 285
rect 100 271 102 274
rect 105 272 107 274
rect 101 267 102 271
rect 100 262 102 267
rect 105 262 107 264
rect 74 260 76 262
rect 128 258 130 280
rect 164 266 166 280
rect 190 271 192 274
rect 195 272 197 274
rect 191 267 192 271
rect 190 262 192 267
rect 195 262 197 264
rect 164 260 166 262
rect 218 258 220 280
rect 19 256 21 258
rect 24 253 26 258
rect 100 256 102 258
rect 47 252 49 254
rect 105 253 107 258
rect 190 256 192 258
rect 128 252 130 254
rect 195 253 197 258
rect 218 252 220 254
rect 19 232 21 235
rect 24 232 26 235
rect 100 232 102 235
rect 105 232 107 235
rect 190 232 192 235
rect 195 232 197 235
rect 19 216 21 228
rect 24 226 26 228
rect 24 216 26 218
rect 100 216 102 228
rect 105 226 107 228
rect 105 216 107 218
rect 190 216 192 228
rect 195 226 197 228
rect 195 216 197 218
rect 19 206 21 208
rect 24 203 26 208
rect 100 206 102 208
rect 105 203 107 208
rect 190 206 192 208
rect 195 203 197 208
rect 19 182 21 186
rect 47 188 49 190
rect 24 182 26 185
rect 19 171 21 174
rect 24 172 26 174
rect 20 167 21 171
rect 19 162 21 167
rect 24 162 26 164
rect 47 158 49 180
rect 19 156 21 158
rect 24 153 26 158
rect 47 152 49 154
rect 87 131 89 134
rect 131 132 133 134
rect 88 127 89 131
rect 132 128 133 132
rect 157 131 159 135
rect 203 132 205 134
rect 53 123 55 126
rect 71 123 73 126
rect 87 123 89 127
rect 103 123 105 125
rect 126 123 128 125
rect 131 123 133 128
rect 158 127 159 131
rect 204 128 205 132
rect 157 123 159 127
rect 178 123 180 125
rect 198 123 200 125
rect 203 123 205 128
rect 221 123 223 125
rect 19 116 21 119
rect 24 116 26 119
rect 53 114 55 119
rect 19 100 21 112
rect 24 110 26 112
rect 53 105 55 110
rect 71 105 73 119
rect 87 117 89 119
rect 87 105 89 107
rect 103 105 105 119
rect 126 114 128 119
rect 131 117 133 119
rect 157 117 159 119
rect 122 110 128 114
rect 126 105 128 110
rect 131 105 133 107
rect 157 105 159 107
rect 178 105 180 119
rect 198 114 200 119
rect 203 117 205 119
rect 194 110 200 114
rect 198 105 200 110
rect 203 105 205 107
rect 221 105 223 119
rect 24 100 26 102
rect 53 94 55 97
rect 71 94 73 97
rect 87 94 89 97
rect 103 95 105 97
rect 126 95 128 97
rect 131 94 133 97
rect 157 94 159 97
rect 178 94 180 97
rect 198 95 200 97
rect 203 94 205 97
rect 221 95 223 97
rect 19 90 21 92
rect 24 87 26 92
rect 157 90 158 94
rect 87 87 89 90
rect 131 87 133 90
rect 157 87 159 90
rect 203 87 205 90
<< polycontact >>
rect 24 485 28 489
rect -11 471 -7 475
rect 105 485 109 489
rect 16 467 20 471
rect 43 463 47 467
rect 70 471 74 475
rect 97 467 101 471
rect 124 463 128 467
rect 22 449 26 453
rect 103 449 107 453
rect 24 435 28 439
rect 105 435 109 439
rect 13 419 19 423
rect 94 419 100 423
rect 22 399 26 403
rect 103 399 107 403
rect 24 385 28 389
rect 129 385 133 389
rect 16 367 20 371
rect 43 363 47 367
rect 94 371 98 375
rect 121 367 125 371
rect 148 363 152 367
rect 22 349 26 353
rect 127 349 131 353
rect 24 335 28 339
rect 129 335 133 339
rect 13 319 19 323
rect 118 319 124 323
rect 22 299 26 303
rect 127 299 131 303
rect 24 285 28 289
rect 105 285 109 289
rect 16 267 20 271
rect 43 263 47 267
rect 70 271 74 275
rect 195 285 199 289
rect 97 267 101 271
rect 124 263 128 267
rect 160 271 164 275
rect 187 267 191 271
rect 214 263 218 267
rect 22 249 26 253
rect 103 249 107 253
rect 193 249 197 253
rect 24 235 28 239
rect 105 235 109 239
rect 195 235 199 239
rect 13 219 19 223
rect 94 219 100 223
rect 184 219 190 223
rect 22 199 26 203
rect 103 199 107 203
rect 193 199 197 203
rect 24 185 28 189
rect 16 167 20 171
rect 43 163 47 167
rect 22 149 26 153
rect 84 127 88 131
rect 128 128 132 132
rect 153 127 158 131
rect 200 128 204 132
rect 24 119 28 123
rect 13 103 19 107
rect 51 110 55 114
rect 99 109 103 113
rect 118 110 122 114
rect 174 109 178 113
rect 190 110 194 114
rect 217 110 221 114
rect 87 90 91 94
rect 131 90 135 94
rect 158 90 162 94
rect 203 90 207 94
rect 22 83 26 87
<< metal1 >>
rect -15 492 5 496
rect 9 492 59 496
rect 63 492 86 496
rect 90 492 140 496
rect 144 492 163 496
rect -12 488 -9 492
rect -3 475 0 480
rect 12 482 15 492
rect 42 488 45 492
rect 69 488 72 492
rect -14 471 -11 474
rect 28 471 31 474
rect -3 466 0 471
rect 5 467 16 470
rect 28 468 36 471
rect -12 446 -9 462
rect 5 461 8 467
rect 28 462 31 468
rect 40 463 43 466
rect 51 466 54 480
rect 78 475 81 480
rect 93 482 96 492
rect 123 488 126 492
rect 62 471 63 474
rect 67 471 70 474
rect 109 471 112 474
rect 51 463 59 466
rect 78 466 81 471
rect 51 458 54 463
rect 59 459 63 463
rect 86 467 97 470
rect 109 468 117 471
rect 3 452 8 457
rect 12 446 15 458
rect 42 446 45 454
rect 69 446 72 462
rect 86 461 89 467
rect 109 462 112 468
rect 121 463 124 466
rect 132 466 135 480
rect 132 463 144 466
rect 132 458 135 463
rect 84 452 89 457
rect 93 446 96 458
rect 123 446 126 454
rect -15 442 5 446
rect 9 442 59 446
rect 66 442 86 446
rect 90 442 140 446
rect 12 432 15 442
rect 93 432 96 442
rect 3 419 8 424
rect 12 420 13 423
rect 28 422 31 428
rect 28 419 36 422
rect 83 419 88 424
rect 92 420 94 423
rect 109 422 112 428
rect 109 419 117 422
rect 28 416 31 419
rect 109 416 112 419
rect 12 396 15 408
rect 93 396 96 408
rect -15 392 5 396
rect 9 392 59 396
rect 63 392 86 396
rect 90 392 148 396
rect 152 392 163 396
rect 12 382 15 392
rect 42 388 45 392
rect 93 388 96 392
rect 28 371 31 374
rect 5 367 16 370
rect 28 368 36 371
rect 5 361 8 367
rect 28 362 31 368
rect 40 363 43 366
rect 51 366 54 380
rect 102 375 105 380
rect 117 382 120 392
rect 147 388 150 392
rect 86 371 87 374
rect 91 371 94 374
rect 133 371 136 374
rect 59 366 64 371
rect 102 366 105 371
rect 51 363 59 366
rect 51 358 54 363
rect 110 367 121 370
rect 133 368 141 371
rect 3 352 8 357
rect 12 346 15 358
rect 42 346 45 354
rect 93 346 96 362
rect 110 361 113 367
rect 133 362 136 368
rect 145 363 148 366
rect 156 366 159 380
rect 156 363 162 366
rect 156 358 159 363
rect 108 352 113 357
rect 117 346 120 358
rect 147 346 150 354
rect -15 342 5 346
rect 9 342 59 346
rect 63 342 86 346
rect 90 342 110 346
rect 114 342 162 346
rect 12 332 15 342
rect 117 332 120 342
rect 2 319 7 324
rect 11 320 13 323
rect 28 322 31 328
rect 28 319 36 322
rect 108 319 113 324
rect 117 320 118 323
rect 133 322 136 328
rect 133 319 141 322
rect 28 316 31 319
rect 133 316 136 319
rect 12 296 15 308
rect 117 296 120 308
rect -15 292 5 296
rect 9 292 59 296
rect 63 292 86 296
rect 90 292 140 296
rect 144 292 148 296
rect 152 292 176 296
rect 180 292 230 296
rect 12 282 15 292
rect 42 288 45 292
rect 69 288 72 292
rect 28 271 31 274
rect 5 267 16 270
rect 28 268 36 271
rect 5 261 8 267
rect 28 262 31 268
rect 40 263 43 266
rect 51 266 54 280
rect 78 275 81 280
rect 93 282 96 292
rect 123 288 126 292
rect 159 288 162 292
rect 62 271 63 274
rect 67 271 70 274
rect 109 271 112 274
rect 51 263 59 266
rect 78 266 81 271
rect 51 258 54 263
rect 59 259 63 263
rect 86 267 97 270
rect 109 268 117 271
rect 3 252 8 257
rect 12 246 15 258
rect 42 246 45 254
rect 69 246 72 262
rect 86 261 89 267
rect 109 262 112 268
rect 121 263 124 266
rect 132 266 135 280
rect 168 275 171 280
rect 183 282 186 292
rect 213 288 216 292
rect 157 271 160 274
rect 199 271 202 274
rect 132 263 141 266
rect 168 266 171 271
rect 132 258 135 263
rect 84 252 89 257
rect 93 246 96 258
rect 175 269 187 270
rect 179 267 187 269
rect 199 268 207 271
rect 199 262 202 268
rect 211 263 214 266
rect 222 266 225 280
rect 222 263 234 266
rect 123 246 126 254
rect 159 246 162 262
rect 222 258 225 263
rect 183 246 186 258
rect 213 246 216 254
rect -15 242 5 246
rect 9 242 59 246
rect 66 242 86 246
rect 90 242 140 246
rect 144 242 176 246
rect 180 242 230 246
rect 12 232 15 242
rect 93 232 96 242
rect 183 232 186 242
rect 3 219 8 224
rect 12 220 13 223
rect 28 222 31 228
rect 28 219 36 222
rect 83 219 88 224
rect 92 220 94 223
rect 109 222 112 228
rect 109 219 117 222
rect 176 220 184 223
rect 199 222 202 228
rect 199 219 207 222
rect 28 216 31 219
rect 109 216 112 219
rect 199 216 202 219
rect 12 196 15 208
rect 93 196 96 208
rect 183 196 186 208
rect -15 192 5 196
rect 9 192 59 196
rect 63 192 86 196
rect 90 192 176 196
rect 180 192 234 196
rect 12 182 15 192
rect 42 188 45 192
rect 28 171 31 174
rect 5 167 16 170
rect 28 168 36 171
rect 5 161 8 167
rect 28 162 31 168
rect 40 163 43 166
rect 51 166 54 180
rect 59 166 64 171
rect 51 163 59 166
rect 51 158 54 163
rect 3 152 8 157
rect 12 146 15 158
rect 42 146 45 154
rect -15 142 5 146
rect 9 142 80 146
rect 84 142 139 146
rect 143 142 164 146
rect 168 142 195 146
rect 199 142 228 146
rect 12 116 15 142
rect 48 135 78 139
rect 82 135 107 139
rect 111 135 143 139
rect 147 135 182 139
rect 186 135 228 139
rect 48 123 51 135
rect 98 123 101 135
rect 117 123 120 135
rect 127 128 128 132
rect 152 127 153 131
rect 173 123 176 135
rect 189 123 192 135
rect 199 128 200 132
rect 216 123 219 135
rect 75 114 78 119
rect 82 114 85 119
rect 2 103 7 108
rect 11 104 13 107
rect 28 106 31 112
rect 60 111 85 114
rect 28 103 36 106
rect 28 100 31 103
rect 60 97 63 111
rect 82 105 85 111
rect 91 113 94 119
rect 107 114 110 119
rect 91 109 93 113
rect 97 109 99 113
rect 107 112 113 114
rect 117 112 118 114
rect 107 110 118 112
rect 135 112 138 119
rect 91 105 94 109
rect 107 105 110 110
rect 136 108 138 112
rect 135 105 138 108
rect 151 113 154 119
rect 161 113 164 119
rect 182 114 185 119
rect 161 109 170 113
rect 182 110 183 114
rect 187 111 190 114
rect 207 113 210 119
rect 151 105 154 109
rect 161 105 164 109
rect 182 105 185 110
rect 209 109 210 113
rect 225 113 228 119
rect 207 105 210 109
rect 225 105 228 109
rect 12 80 15 92
rect 48 87 52 97
rect 75 87 78 97
rect 98 87 101 97
rect 117 87 120 97
rect 135 90 138 94
rect 162 90 163 94
rect 173 87 176 97
rect 189 87 192 97
rect 207 90 209 94
rect 216 87 219 97
rect 48 83 75 87
rect 79 83 107 87
rect 111 83 143 87
rect 147 83 182 87
rect 186 83 228 87
rect -19 76 5 80
rect 9 76 59 80
rect 63 76 91 80
rect 95 76 120 80
rect 124 76 145 80
rect 149 76 209 80
rect 213 76 228 80
<< m2contact >>
rect 28 485 32 489
rect -18 471 -14 475
rect -3 471 1 475
rect 36 463 40 471
rect 109 485 113 489
rect 63 471 67 475
rect 78 471 82 475
rect 59 463 63 467
rect 5 457 9 461
rect 18 449 22 453
rect 117 463 121 471
rect 144 463 148 467
rect 86 457 90 461
rect 99 449 103 453
rect 28 435 32 439
rect 109 435 113 439
rect 8 420 12 424
rect 36 419 40 423
rect 88 420 92 424
rect 117 419 121 423
rect 18 399 22 403
rect 99 399 103 403
rect 28 385 32 389
rect 36 363 40 371
rect 133 385 137 389
rect 87 371 91 375
rect 102 371 106 375
rect 5 357 9 361
rect 59 362 63 366
rect 18 349 22 353
rect 141 363 145 371
rect 162 363 166 367
rect 110 357 114 361
rect 123 349 127 353
rect 28 335 32 339
rect 133 335 137 339
rect 7 320 11 324
rect 36 319 40 323
rect 113 320 117 324
rect 141 319 145 323
rect 18 299 22 303
rect 123 299 127 303
rect 28 285 32 289
rect 36 263 40 271
rect 109 285 113 289
rect 63 271 67 275
rect 78 271 82 275
rect 59 263 63 267
rect 5 257 9 261
rect 18 249 22 253
rect 117 263 121 271
rect 199 285 203 289
rect 153 271 157 275
rect 168 271 172 275
rect 141 263 145 267
rect 86 257 90 261
rect 175 265 179 269
rect 207 263 211 271
rect 99 249 103 253
rect 189 249 193 253
rect 28 235 32 239
rect 109 235 113 239
rect 199 235 203 239
rect 8 220 12 224
rect 36 219 40 223
rect 88 220 92 224
rect 117 219 121 223
rect 172 220 176 224
rect 207 219 211 223
rect 18 199 22 203
rect 99 199 103 203
rect 189 199 193 203
rect 28 185 32 189
rect 36 163 40 171
rect 5 157 9 161
rect 59 162 63 166
rect 18 149 22 153
rect 80 142 84 146
rect 139 142 143 146
rect 164 142 168 146
rect 195 142 199 146
rect 80 127 84 131
rect 123 128 127 132
rect 145 127 152 131
rect 195 128 199 132
rect 28 119 32 123
rect 7 104 11 108
rect 47 110 51 114
rect 36 103 40 107
rect 93 109 97 113
rect 113 112 117 116
rect 132 108 136 112
rect 151 109 155 113
rect 170 109 174 113
rect 183 110 187 114
rect 205 109 209 113
rect 213 110 217 114
rect 225 109 229 113
rect 91 90 95 94
rect 138 90 142 94
rect 163 90 167 94
rect 209 90 213 94
rect 18 83 22 87
rect 91 76 95 80
rect 120 76 124 80
rect 145 76 149 80
rect 209 76 213 80
<< metal2 >>
rect -17 488 -14 501
rect -17 485 28 488
rect -17 475 -14 485
rect 1 472 21 475
rect 18 453 21 472
rect 18 403 21 449
rect 29 439 32 485
rect 64 488 67 501
rect 64 485 109 488
rect 64 475 67 485
rect 18 375 21 399
rect 29 389 32 435
rect 36 423 40 463
rect 24 385 28 388
rect 17 372 21 375
rect 18 353 21 372
rect 18 303 21 349
rect 29 339 32 385
rect 18 253 21 299
rect 29 289 32 335
rect 36 323 40 363
rect 24 285 28 288
rect 67 288 70 475
rect 82 472 102 475
rect 99 453 102 472
rect 99 403 102 449
rect 110 439 113 485
rect 117 423 121 463
rect 126 396 129 501
rect 88 392 129 396
rect 88 388 91 392
rect 88 385 133 388
rect 88 375 91 385
rect 106 372 126 375
rect 88 370 91 371
rect 123 353 126 372
rect 123 303 126 349
rect 134 339 137 385
rect 141 323 145 363
rect 18 203 21 249
rect 29 239 32 285
rect 64 285 109 288
rect 64 275 67 285
rect 82 272 102 275
rect 18 153 21 199
rect 29 189 32 235
rect 36 223 40 263
rect 99 253 102 272
rect 99 203 102 249
rect 110 239 113 285
rect 154 288 157 501
rect 154 285 199 288
rect 154 275 157 285
rect 172 272 192 275
rect 117 223 121 263
rect 189 253 192 272
rect 189 203 192 249
rect 200 239 203 285
rect 207 223 211 263
rect 24 185 28 188
rect 18 87 21 149
rect 29 123 32 185
rect 36 107 40 163
rect 80 131 83 142
rect 92 80 95 90
rect 120 80 123 132
rect 139 94 142 142
rect 145 80 148 127
rect 164 94 167 142
rect 195 132 199 142
rect 210 80 213 90
<< m3contact >>
rect 3 452 8 457
rect 3 419 8 424
rect 59 458 64 463
rect 3 352 8 357
rect 2 319 7 324
rect 3 252 8 257
rect 59 366 64 371
rect 84 452 89 457
rect 83 419 88 424
rect 144 458 149 463
rect 108 352 113 357
rect 108 319 113 324
rect 3 219 8 224
rect 3 152 8 157
rect 59 258 64 263
rect 84 252 89 257
rect 83 219 88 224
rect 166 363 171 368
rect 141 267 146 272
rect 175 260 180 265
rect 172 215 177 220
rect 2 103 7 108
rect 59 166 64 171
rect 47 114 52 119
rect 112 116 117 121
rect 97 108 102 113
rect 127 108 132 113
rect 155 108 160 113
rect 184 114 189 119
rect 213 114 217 119
rect 170 103 175 109
rect 200 108 205 113
rect 229 109 234 114
<< metal3 >>
rect 58 463 65 464
rect 58 458 59 463
rect 64 458 65 463
rect 143 463 150 464
rect 143 458 144 463
rect 149 458 150 463
rect 2 457 9 458
rect 58 457 65 458
rect 83 457 90 458
rect 143 457 150 458
rect -3 452 3 457
rect 8 452 9 457
rect 59 452 84 457
rect 89 452 90 457
rect 2 451 9 452
rect 83 451 90 452
rect 140 452 149 457
rect 2 424 9 425
rect 82 424 89 425
rect -5 419 3 424
rect 8 419 9 424
rect 2 418 9 419
rect 59 419 83 424
rect 88 419 89 424
rect 59 372 64 419
rect 82 418 89 419
rect 140 396 145 452
rect 102 391 145 396
rect 58 371 65 372
rect 58 366 59 371
rect 64 366 65 371
rect 58 365 65 366
rect 102 358 107 391
rect 165 368 172 369
rect 165 363 166 368
rect 171 363 172 368
rect 165 362 172 363
rect 2 357 9 358
rect -3 352 3 357
rect 8 352 9 357
rect 102 357 114 358
rect 102 352 108 357
rect 113 352 114 357
rect 2 351 9 352
rect 107 351 114 352
rect 1 324 8 325
rect 107 324 114 325
rect -6 319 2 324
rect 7 319 8 324
rect 1 318 8 319
rect 103 319 108 324
rect 113 319 114 324
rect 103 318 114 319
rect 103 297 108 318
rect 103 292 146 297
rect 141 273 146 292
rect 140 272 147 273
rect 140 267 141 272
rect 146 267 147 272
rect 140 266 147 267
rect 166 265 171 362
rect 174 265 181 266
rect 58 263 65 264
rect 58 258 59 263
rect 64 258 65 263
rect 154 260 175 265
rect 180 260 181 265
rect 154 259 166 260
rect 174 259 181 260
rect 2 257 9 258
rect 58 257 65 258
rect 83 257 90 258
rect -3 252 3 257
rect 8 252 9 257
rect 59 252 84 257
rect 89 252 90 257
rect 2 251 9 252
rect 83 251 90 252
rect 154 251 159 259
rect 121 246 159 251
rect 2 224 9 225
rect 82 224 89 225
rect -5 219 3 224
rect 8 219 9 224
rect 2 218 9 219
rect 59 219 83 224
rect 88 219 89 224
rect 59 172 64 219
rect 82 218 89 219
rect 58 171 65 172
rect 58 166 59 171
rect 64 166 65 171
rect 58 165 65 166
rect 2 157 9 158
rect -3 152 3 157
rect 8 152 9 157
rect 121 153 126 246
rect 171 220 178 221
rect 171 215 172 220
rect 177 215 178 220
rect 171 214 178 215
rect 78 152 126 153
rect 2 151 9 152
rect 47 147 126 152
rect 172 156 177 214
rect 172 150 234 156
rect 47 120 52 147
rect 111 121 160 122
rect 46 119 53 120
rect 46 114 47 119
rect 52 114 53 119
rect 111 116 112 121
rect 117 117 160 121
rect 184 120 218 124
rect 117 116 118 117
rect 111 115 118 116
rect 155 114 160 117
rect 183 119 218 120
rect 183 114 184 119
rect 189 114 190 119
rect 212 114 213 119
rect 217 114 218 119
rect 229 115 234 150
rect 46 113 53 114
rect 96 113 103 114
rect 1 108 8 109
rect -6 103 2 108
rect 7 103 8 108
rect 96 108 97 113
rect 102 108 103 113
rect 96 107 103 108
rect 126 113 133 114
rect 126 108 127 113
rect 132 108 133 113
rect 126 107 133 108
rect 154 113 161 114
rect 183 113 190 114
rect 199 113 206 114
rect 212 113 218 114
rect 228 114 235 115
rect 154 108 155 113
rect 160 108 161 113
rect 154 107 161 108
rect 169 109 176 110
rect 1 102 8 103
rect 97 102 132 107
rect 169 103 170 109
rect 175 104 176 109
rect 199 108 200 113
rect 205 108 206 113
rect 228 109 229 114
rect 234 109 235 114
rect 228 108 235 109
rect 199 107 206 108
rect 200 104 205 107
rect 175 103 205 104
rect 169 98 205 103
<< labels >>
rlabel metal1 9 192 13 196 1 Vdd!
rlabel metal1 10 242 13 246 1 GND!
rlabel metal1 10 142 13 146 1 GND!
rlabel metal1 91 242 94 246 1 GND!
rlabel metal1 90 292 94 296 1 Vdd!
rlabel metal1 90 192 94 196 1 Vdd!
rlabel metal1 9 292 13 296 1 Vdd!
rlabel metal1 9 492 13 496 1 Vdd!
rlabel metal1 9 392 13 396 1 Vdd!
rlabel metal1 10 442 13 446 1 GND!
rlabel metal1 10 342 13 346 1 GND!
rlabel metal3 -3 452 -1 457 1 a0
rlabel metal3 -5 419 -3 424 1 a1
rlabel metal3 -3 352 -1 357 1 a2
rlabel metal3 -6 319 -4 324 1 a3
rlabel metal1 91 442 94 446 1 GND!
rlabel metal1 90 492 94 496 1 Vdd!
rlabel metal1 90 392 94 396 1 Vdd!
rlabel metal1 115 342 118 346 1 GND!
rlabel metal1 159 363 162 366 7 Y
rlabel metal3 -3 252 -1 257 1 a4
rlabel metal3 -5 219 -3 224 1 a5
rlabel metal3 -3 152 -1 157 1 a6
rlabel metal2 -17 497 -14 501 4 select0
rlabel metal2 64 497 67 501 5 select1
rlabel metal2 126 497 129 501 5 select2
rlabel metal1 9 76 13 80 1 Vdd!
rlabel metal3 -6 103 -4 108 1 a7
rlabel metal1 67 135 74 139 5 GND!
rlabel metal1 75 76 78 80 2 clk
rlabel metal1 75 142 78 146 4 ~clk
rlabel polysilicon 53 106 55 109 5 D
rlabel polysilicon 71 115 73 118 5 reset
rlabel metal1 72 83 75 87 5 Vdd!
rlabel metal1 180 192 184 196 1 Vdd!
rlabel metal1 181 242 184 246 1 GND!
rlabel metal1 180 292 184 296 1 Vdd!
rlabel metal2 154 496 157 501 5 select_out
rlabel metal1 231 263 234 266 7 out
<< end >>
